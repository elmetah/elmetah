MPQ    �(#    h�  h                                                                                 ��A=,ʵ�w��1��}匍��$T���b�)`FV���&J��:����ֹ�h��l�~a�\	!�=A=C`�q�H�DH�V���B�7&�N6�ݓlhM�yƹ@0�z��������0�X2O���o���lnJ�X���<��5qP�<.�O��jy�ғ����z���N�W��=�����][�P��R\�C��@{��!��3T�˝��X�ru��0����:
�
�l�Y��$��y��$)X��G�N�'E�\��5�4i�&��3�a)��*�7���څn��G�����K�Q�`_!�\�W�I���^m� {.���2?�/
63`/�"�J�|�Xo��-K`�0�(Xݫ�0-�92�R���"��so���B�w*�}гh싧Gn���'vW� ���"D���B��˒A�c����	��MfôﹸFB���~�E-��K���?�ҍ��Q����c8��A�t�9Kj4[l_;.�U|��4��٩�B�no>d�QƗ'�w��`���O�f����%B���@eUA�V��s:�#m4[�(�;>�К"�[;���]@�u�3����¢�x��iw��M�GpZ�)3T���v8�vJ'�Q~��9��u�S���F�ʬ�.Fi�Қ��Ǡ3l㕬,��&�y�S�����I���>����膚k*[ɥ��g�@�����������-1�G�;]��Bձ�w�Vu�\4�㒵:N��*��*@m%�ۀ�/|'
��F2�4��r���hp��Rr<晡���?_4���}�$�l�p�豨�׵�5
jq���OeOs��D�������-���9�E�# XV��T>�$��ߧ�a�-�:��G���&p�J�qy���οG�5z��%6D�����ï+�;s��A4;',hz�v]��le"V�~����/\�0���,]m��!�y�q
3	�@�fLK�"��fQ��&�D{���=V�6����_��JT�����s��]�:/��8�RBal����=�J�[�J������2���+�sˤHQ���I�}�k��G>z���=F)�������0�a����p�%_/�_&5�,��Y<*���f�^'*:�3+�kq���X?�Y3<ܲ��K� �)�@!��C�'��((��a$����J��WC��9h�T�V�HM^7����rjU,�b����>�c�t����CWU��o�b'���
#��He6���\������Z����]٤]�wٽS/���9��^I �TlS��mNd���G����L�og��x��Q���#�sE�}�Zu�ٷ��(֣� �ٹ�љ v�߳�3���C����dOp)���鹀�|ޠ��������E��M�4�A_���9&��1��*8��4��:&�US�fh��do���"��+⩑�aˀ���>�Z�1���tH'��ߘ�2�nwT.nG�W,��B�A�����7}�A��Rƙz�u���aU��8[�-n_@y8"<�j`�L�R�{�5��I,�{'/v��2�=aq������+P!,�^ �hR#�D�r�p\Qm4D�|vb�N��N�MI-mk���>g�p�U�'!�~La��Y���{~]nN5
���9D��d�8����q�X�	B��izo������E��|��:��bv�$�%ǀC�R#{L�ݕ9B�8u^�s?$[�6�9]�A1�>�S���&���0��X�g6�II���MX&5G���Z��T�p������N����;�z_8Sb�~�f`��$vN��]3�!���	�O+������E���׋��{�?�P�!�����50�L�~�9}ۂ ��7K���+�}&7Ո#�<@+����?}��.ǜI�D��^
�࿇�g��~g��vz_��3_��7rj�ng%�5^�H��KQ�Ud&L͓LoǊ���Q�)�XC��/��[e (Fx5�t����[���yW���������j�9�c�>7p����n�S��d���~���!��-�g��?��G�s�����֎qd�0�ף��V���l=	��P#�L?���َ����8������B�<Wq��#G*��I��@/�<= ��K��������}�*�5�r�ᝮ�9Q]}]{�ʖ�	{���s($��$Ʒ�Q�q�ip̫�7�^�T9��I#+��%;�����5�ͥ|�������.%CU�$��Sf�J�9�� ��5� �S��E�G�=��ln 8�T�*k��gI�t�A�f�cr�6����\!�Ŀ��wI*Y2��d@h�8W��=��Ѐ-sE�ϒ��"Ԛ�^u��/+��c�B���?�SG7��TC-��!oP��;��D�����s�/֗��%Ot17���H@�U^/���zZ?%��x����6�^���A�v)�;۱s���c�w������b�#�=�G6 Aq��in�C�2�~qo�6'�n	D�����:]!��UXeA���\�(���I7�{�����pv�1��u��6�1���(����mɟG^�R砾�ڒz�P�otG������E�X�ut\���)��"N=(���[WkE�Q��棑�����sW�뎟�M&=�`���\�h�˲�̩����= í���M�R ������נ���uwlLo�Ⱥtշ�i�[��.�/޴ڂ�Y���m�yË~d���M�%G�f8�4�/c�D+��r?�yg�ߛ Jn+c*���Y"����y��u둚��$�.#�u,����j��Le��$E�=Z��Җ��#E��c�5�bAB�oWP\V~�{�QrYG9FQ׻Gs{�F�:���1������|$i�_\��a�x8�`g�\�tu=�}�߳�12�Bn�/�7;�b�s�Zՠ������S��F1$u�)OsLK�T���ڟ�	b��<�#_v|�A����k��P��?4���U�1�O��*��
i�F�//�V-�σ�KVW4���8���+���+*��		�=�E)#i���t!�0s����c�
7x�9p��C�>(֫b/�u>�/�c���=��(�<dH͆�9��0#ܩ���Q�R�X�g��=����V�a����R(���UB��rW��>��P�}#ۄ#� �C���lM/��Ž@�g0C�$�x�����~��,��i�>]cz�p���l��ە&$��2����v�n�8\bj��}�d/���j��hn\�ؓ��
 %(��яG?�5������}��}�cG�g����թ5�A^H"��D��b�W⠑��F�~O\�	�_~&U2:tiA��|���V)���4��]�~���+�(O)u퍍V��j 묦*nAUF<Ts�pe���M� �i�w�̋!�Ii�F
a~����V�i�1�AsA�N�����cy|	Z�Ap�q�owiI�1�M������Bzx~�:p-��\K�=z�CV��m� �!��mf�c�<�A��9ƿ�[Gd�.���|�!�tB���o���Qᔻ��9`l�aO�z�B�E%=�>Ǜ����]V���%4#H�B[��νֻ"Е?O�lU.;��1)v��3��8 �*�=�{�e׏��MG+AA)N��d8o'^'�[���p���J�-��.a/�Mg����L3��&�G�}�!]�s$��\�*�}�-�s�i�-�_�TPɠ�?gS=�eA��	�
[z�#��ׄ]|s�լ<w~��G.M����pe8�m���|�k���-�O#t���2�_p	�C�r�P���t?�����B��?C�l"�K�[�����5�?�����O�����o�2f�%{�p���*SVEAd�XQ��T��1ÊO�|����d��"�P�a�:J�C�y���)�����e��&�DB���3m�f��։��<�'���zS���X�e�}	���»��X���0��],����y��Oq�텓�I�f��;"�ĤQ|_"����B�1�Q\�j�����Շ�{��d]��<�U�FR�V���Y�=�*[^���O7�Z������ �s�%�Q�nI]yk��>���yk�)������<�a�{���{p�W�_j_�O��5�[�,��*�3\f����k�3ዏk�a���B��T���kK�"�)3 �!=��C�3i�d�j������c�W�1�9���ֶH(Ԉ7�a���LP9"��i�>�IP�4�>l�C�����^D�:��D�C#����P��$��~��(��c��ٟ fw4��/h �(ٟ�p ch��Nm�~�廵v����*@�h^�̅�����B}=������.7���Ԫ��_��h��n���d4@���+Oˬ.ڟ>��F�|Y*����&�+��EB'?�/i^_�:����!��L�l�ɻ����uAU�_�h�fd�]�����1�>�R�[���(tZmc�����'j���SH����[T�ذ��ÿ�7
��ڕ��p7��ư�ƴ�u��<�i�s[�-�u�@t3�<�!�q?��=��J٣V7|v+�2~��a�O��ҷձ_�F��,���C�����:�m/Ս�&�b�
ܞɁTM���k�狣y>Ch�$P�p���9�Ja�&Y�5{YngNpB*
��i9?/�׿´�_t�q��a6���%�o5���|ԧE����� �:�E�v�g%|>/C���{�F��0ô�32"�Λ_[s89x��1$�Sdь&���t{�ٯvߗg�'�I����|X��G�:���DJO=Ϳ��l��NJL�;��UǖS���+e����5;�3�����	<��+w���C'��; ���5�?�d!����8��0l
��`}v#�����n�]�&8���]/���+�%t�ڈr�����r���8�y{��[D��{�ֹ�̒�b�
�_�H�-���茰-��Q���VU��͎a�o"?_�W,�lژ��0����H�,�e�taxet���P&���-��v۴��7RWjJ�8�^N57��h��ػ�n��d0���Y��\s-����:6�GI���Y�f֩i9���K��HJ���=���Pd�L�	(��E���`��ӯ���#���wB�5fq�����ǈ@F�[��<��\���:�)C�}�ox��rcc����]�Y�{�6��Db��V^(2�$!����q83i���o^K�'��I���G��B�;�Pe'H�gD �P����U�\�����Ju\7�;5s�@SsX拂���|� 3b�� �kv?I��6A+oLcM T6���$��!����g|�wc�YMo���aRh���W�2�r�-nފ��W`"�^@^�SCcΒ+^Fvc�kyŎ� �N��F8�C�I`!�2�sݓ;�7�2��}�"��]\�V�qO�M�1R��&�@�p/UX�#��:��4�����6�Z��Z�KQ�M;�:��*�r�n��w6b}��>�����x�Z�$�����<�y��oMƙ'��	_�#�'�q8���e�!���)�D�����R��ZO'�K�l	2u��숞@^��w��q���Yi����-'��P�zG�]��_�GL
�y΅�sI�t׀��⾞��[=��Y��=�Wڦ�����b)�N����+�M�P'`�q�\;ϫ�m�
��X�zʱÈ�d���R����1S0��[������L�F�ȕ;����fE��K�/9qk�F���3�ymr���Yֹ�/�.%��8�^4�,������i�y���<�nF�*1oMY^��a�u�E�i���$O篠P���+��6�e�x��;hZ��D����E��cl�P����
�R�f��0{��2Yb$QR
�sV �F���1�׹�xz~�7#�i�5���x��gI����=�\����2�h�n5���uo;���s�;�6蝿��w֔S;�1?!4)ʢ�Kɧ�ک��:�	]�����_1^AN����P�y?o����7*�����0�
$JRF±�������K�g�tv���F~z+�O�	$�"JV�#D����<�������1�d�73VyT���۫(�v�U�uٴ�����&�}��W�b����Ԧ�#�(��齘M)P�vL�B��AR�Ѽ����΍d{�d߹�N�W��=i��<��ز ���	�M��ŸB�g�E������9��y����b]�;p��rl�U��PM��z�an�Q�n�s� b/�xt�/$�-�N���BU\����n��s�%ÀW���?�9�INΘ�}y̠�BD�:I�5ObH�zD�ǳ{������h���~a��:�b
i<�;c�=�hz*�:s�4v�6�Yu
�V)>����u�Qg�:�j���E��U��s��O��s���� ����-����Xi� a�R�VWJ�_�EA��ߩ�����y�eQn!S�Lr�w��a��$M���O�7B5X~��#-�xKз�~��'�����U�c�KA�79A5i["�	.U�����/����o�Q���m��`Gk9O��K��'Q%8}����9��HV��Zi1�##
�[,��qY�А�x��Ł;���)$��3�3[�i�ؽ��S�OdMG�G4)i�6�u�8J�!'X
F�� ��ky럥R��@�3.|۠��S��}xU3��>��ɔ���\j���E����41�h�,����ɛZVg�Y� �P޸甅ݳU�&����](�է��w\�Q��y_I�E�0�����(�Pvm[���$�|����S�m�j���h�X�:��~�rr�f��R'?O��a�?�Z��l���g.N�+�5@5���6DO�D�ḻ�}⍠)�K	��e��E��,XLi�T����E}����s�0^(��ϭ���<JK�y{����ϫ���GHD�L&��篡 �q�օ7(�'�ڇz@X��dWe)��[Ի3-�eY0�t^,6$�?�y��q Ȏ��s�f���",�zQw��������21�l>��Θ�ԇ�rg�a�]�����=R�lȎ�&�=�W[9*	�A������d:��sA��Q	:�I���k�T>���6){���y�Wh7a��7p�-_��ٽ갡5�'ׇ��*j�f�Z� �$3�Fk��A͎f��OA=�h��KKdS)N�I!��Cv_&Wu�_�H� {W��9��O�L�H��73��3FJKfͯf��$QD>����]G��C�]��/ñ�2�����#]s��,��7�Y�x�c�h��ZyٚÉw��K/#�C�ͤ��b >��tm��M�C?�Mf���8��x�G���mR���}؅���I
�ަJ�v���寧я���C Ʃ����D���O&Pv��z��,J|��d��q��f��Eݢh�*X�_<	��9r�����t0�nU�F�h� �d%WAӘDQ�L���F��6���2�Z����^�'��l��C���<T$c����i�M�>����;�73\���~cu�a��?Nˮ{P-B��@oN�<t?#��6p��� ��jR�1gvMV2C}a�
�k;귐l�a f,|���T������7?m*�`2��b[�����M?z2k�m���"�Kk��ڃ��a�Y���{4�N���
2�"9:vX����fHq&��܂~�yFop9���E�Ϙ�8r,:=v-%��ICu@{¨��l��.b�)�[.&�9���1��>S?�&t
�RPvL8�ц�g��vI���CC�X��G.�r���RJ��Ge'�N&q��z0OES؎)�����LĐ8�3pS�m^	�hf+R+��~�'�{���I���?F��!�L鴳��0G����^}������^hP�}2&SCy�~����1�+���u�z�L����f�*������m�����r������t_W�薧���+m������U�	�͉��o}������1��Nk{˽�r��eV�x
�tv�?� �!ޫ���aۏ'�r"Uj��Y�7&�t�NMщ�pd�f_�4_CϗN�-+ͧ�5��G��Κ܃�ā��&ë��ӭ�I��=?4pP�KL����e����Ց.:ų�+����B&N�q��=)�CW��v�o<3cB��셧u�(���}��v���r��	�4]V�{k§�i�0E�(��$|�t����qS�if;��S/^���oN�I%���s^��Hg�k�ê�B&[���d�@U����	��J0��V�5�uSN嶋����(� .:o�
�Mk1�I�^RA���c(8e6F��,!����)w��.Yh��Z�PhգbWI'����-i�<�H0I"JBD^���ތ+9�yc���)?�I/�ԡ;qC��}!�x����;kp>�����	������}O�Gw1m����z�@p�Q/?�v����59/�k��6w���`!,'�;Qf��2�<�mk��@�Q�v�Y���=�G����_4��y���t[�o�u5'[�	z�h��3U��=61ew���2Q��ҕ�m�!���9�&v����uC�2���b��|��"��"Mɕ�+�=��z��ͩ�ppG�;�4
J��tR�y𽤣�BE�=8�/��]W5z��Q��٭p��qk�)Yc��M\��`�#\�U}�(���8��v��c���6�RS2k�������qg��?�L
>��p"�PyTOm�ȈQ/�M��	[�NL�m���4h��j��%}�A8	�F4M��𝁨��y]�֛�y n��*�N�Y1������ Q,��0$ʿ�+��fj���b�e�����ZC���jE��cG;0���q��d+Mmo{TYwY}/�Q�x�s1>�FG2M�j1����-���A�i�+�����x�i g���Ūl�=�[Z�i|2��nP�]%z�;bj�sN���ů蘉}���%S���1Z�,)E�K��Ď��i^	X����_���A2��a��P�cC?�㔝����U����
ߔF�S��L�M���K̗�=k��秼��+�%	?��ņ#��w��f�"��Z:7o@(�9W(�a�؛xut��j�_k��8�Qr
��|a�<#R,c�PbB�H�c�x��R���+�G�L�s��Cg���$�������WH��j��u��5� g�:�qMe>�ųdg榿�����C�������_��e{]��ap��plW�x�6z� �J��`��,(��69b�/W�s,"/f��	�X� =�\�@�I�T�K��%^���ux?u� �2�γ�}�Tƛ��uܨ5�>H��D>Ì��3
�Yډt�_��P�~�q3:IȘi7ږ����#���U.!4��4c������^�u�5]�}jvh�`��U<�s`��(uC֓ ���-�O��J,i"I?a�b�ZU5V�	��^MAG���0�E��y��� ��'a�wߎn�g�M=G憎�B�ǎ~�^-�!K�Q̓��壣g�!1�#eLci�A/
9�ʅ[�͸.���겋��
��S3oo��Q�;��ڎ`"[aO5�q�xz4%3#��Q5<r�V���\�#��	[g�x�Ћ��"VU;C#�D7ly�3�R���<�s���돪�G�n�)����8%�'�8�����f��� 9;��aw.��Z�C`��X.3�*�}���Q�)'�%�`e{�#k"[{�ޣ��<�ɖ��g	��۰��wN� ��0�9��S]��>բ�Xw�,�ʍ��d����pӻ7ۈrm�O=��W�|8p>���Ʌ-���7K��+���|r���P'?p���6�u#�l�H�B!S�fR�5�J�����Ov��'�w�8�f��(�&����@EwE�XG��TO�+� ����'S��w�����<�J��Qyv`v���fЉ���=D8���]�0��o5m�2RJ'=Dz�ԫ��e������ջn�� A>0�i�,n�?�� y��kq{�#���f�z�"���Qr���UY/���T��@j`Z����i�Z��D�]�{���tRs�܎�h=�O[�̓Df����&�5���s��;Q$6IS�2kvf>+>$��&�)v���_�=a�m�.�p�#�_�E����5�/��;�*%��f���.}3���k"�|�)���J���$KƷ)i2:!3ٺCQ��aZҠ����[�Wt�19������Hޡ�7n�g��_�F�������r>���*	"=�C;v��G��Ju���#v���H�՟4$m��Jٕ�iw�$(/�g^CĤ�! �Oh0m���㇨��ڠQ+٨�����j���}sK0����9?��1/��
�z�
<�i.��Ђ�uڱ�1O�^P�Z�
30|O��[jv硾(Ex>ʽ%gL_��R�j��݃\�bһO����#oU$M�h��Kd�p��S���g_0��v�Ş2]<Z�&����' *3������l�T�(Ц� �G�"�v�����7���<Fc��0�u
W���b���-��@j��<��d�}��W�����v���2���a���� b�Ksܙ|��,��J��╗�J7�AU�m%W/��b���G�M�P�k������-F�&�����a9BY
�s{�iN��|
�z95�g�u/��w�qA�WT�co���ͲqhE����J:�^|va�%r��CP�k{�*#�f6�)섴�[�M�9��e1�VSU�&L-��M�q3�,NggmCI�*ܾ�XX��aGiK��+dEC���W|�T�NA^�1��CS2��7 �0���US3+�+M�	2L�+-~���L������?�#!��.S0"�/�O}�����������[&n�e��/
����+1�O� ��	�Z��u��鯝Y�Q��H7�/u�G>r� �_��
���������,r����pU5+
̈́�o�A��7�������˘*�W�ke�m`x5Ct�������<@ҹy�T�j|b���j��`�TW7�:��L�"Ѥ�d&W��_��Id-�/w�0��G�s����߹������k~�ۄ��=��P	F�LP*ϻ }����R���法�8�3�B���q�gBX	���t���<�4T���ѧ���_j}��.��r��B�$Œ]�r�{Fnh�����S<(֛$׻��?�qn�{i�1�Ȫ�^��
��I� �6�ğ� �����>]f�()�43��r#U�,��dl�J��qb�5i�VS)����0����� )}8�eE?k��I6A!�0c��6W�m�Z�!������wz4�Y�oX��h;h���W��y���3-dp�ϣ(�"F�^�)LYk�+�c>��đu�D����^�C^G?!�ޱi(;Fɣ���ʳ|(���FJODa�1�5��u�.@K/z3i�YN0s}�ꄥ�&++6#���P c�P;��ͭݰhph���mؼ�th�ˢ��u��� �o+"oE�'?T	��U�����lx��eQ���49H�PI �� �Pp�&��?�u��P���B�B���Y�p�1
��t�㗃�H��z}i6���G����e���Xt��G�8�}3=Ӂ��W�}���8���k�X�ٳ
��?�M��K`�ߛ\����ө��͡pC��>][���R����	�$��m����L�U��K)��[��xM���6/�I�����i�tmhA��å��%�8��4�E�u́��y�/ԛ���n��#*gN�Y$��R.���2��q
$E�-��ۏ�m=�l�te��HV�Z��T��L�E���c"����@:3H�ogX{@Y�Z�QHqs�F�&T��1�_��.N���HiB����x�r�g����E�=�z��z62H��nk�-���;=�s�?�q܀�sq�-	�S�7]1uٍ)�a�KEiP�f�p�=	Sb�MXv_��{AM�l��n�P�m�?�(��&���o��;�
���F�R���y`B?K�a�����2 ����+[�	Z2F@�F#�j��%�ݲ[����_t��7�7Z�����J(gl��u�|�KU��kx���Z�����G����#��1���ޘCa��Ӭ�P��F�d���>�|���=��� ����W�^������d���� BA�H�FM ��Ů��gA(N�U9��)��/u�ýƴ���]4� p���l��4��m��;Ң�Ws7������eb;t�n�/�=���R��W\|C[�$ֺǆ��%��؝�+?������Κ�}o����VAӰ��5�1�HkD�𱳈Ց8I ���C���6~�/�:�Mi2�%:��!��p	W4l@�q��̛����u�9og!�j1W��{`�U�xs;;5�N��1p �vK�j��R��i=��a����5�,V���%�A��6�_��� �ly�}xd@]�p�wyo�H�M�+��B�W ~0p"-UK����ժ�>@�Q<�~��c$-UAJ}�97�N[�2�.˖s�M���u��k�o*;�Q2L(�c�`�j�Op����%.�'Ǭ��-KV�a�_�6#�_�[��{���kІ���}�;�ޮ_j��3����ѣ�/����,G\�)�W�k�8 ��'�Bޅ,H0�a�s�[?b�3.��\ݾ���3��3X0��ʨ����X��q>�{Y���6���1��א ɑ��gd�w���W=�{B��\�3_�]M�m՝tfw���H?ZK��&ħӖ�)�m��x���c|�"���}�ɠ�r�^�	��G���N3r�P��}n?�����|�ِ�[l�>��4�ס��5v�����OѰ�����Ss��F�e���^�E�XB��T��û��͝Z�&�軳�x��]J�yqߒ:yx�!����zD�5��8K�����[�-�'��tz���0�Ke���t�ǻ�A��"�0�~�,�~[��`�y#Fq��D�~'Zf8 t"bJ�Qm���8��s����b�ۿ�[�{�����߰�]�&��f��R.�4�!�=�L[�'�!S�+�0��%�@�s�g�Q?
vIΫqkQ� >f�J�)qF��/����a7�E�
u�p�99_sE� �}5�h�=��*�sf���3rn�k]�k��X�E�.���K�G�)��r!��
C,���;�j}l�����W/�19ԩ��B�H���7��ŕi�
A ����`�>��H�~@���CC8T�e�T��ǴU�#Әp�^�������ٻ��4Zuِ�wE�D/��y������ ��;?{�m��嬿d�av�[�����= ����1�f}1���[��������%�]х�W������<�5�˱��)O���,��%Y>|ʆ��6�����[E�c� �_�J�%�_���P��<H�*���&cDU�sJh��md۩#��}��[ũ}%��쀉�m��Z>�Z��Ȗ'{��߄�e��S�T�5Ё�翂��ts�;Z7�Z���[��u�l�ͨ��$�-xL4@e�<*��8"����}���&Dv��2O�Va���!�9����0K,rL����F�0��ܒm H����b��0��GM5G(kxٺ�*bP9S�A�u�N%�j'�aT��Y�$U{�`sN!��
h�<90d��Е����q\�e�{�/Ro�Gz�M�LE�S%��tI:�Mv7��%�d�C+��{8�)� ��$)V��p[��E9���1��S���&��c∢�l�ɯ�5�g"@4I)�5�9��X���G�¥�#�@�J��i#��eN\)��]]澒SN�$��J=����F�(3� FM�	�O.+�q�������;��F]�?�_�!�U��k�0�j��}G�����"�o��Zx&��z�tɹ�|+lrK��k3��u��M*0Y��^�̑�#w��jd:��~���%_�f^�u��W��!\�pF�7z�U�l��`�o3�����?�D@��s�����e�Dx u�t,8"�FN�W ��f��E�ٮ�"�j���O�7ܤM��<ѿ�Id�gO��~3�e�-a��+X/GZ	���=���)�Z0�FI�ۿ˨=u�;P�L��b��H���ؑ$g�p��n�NB\�#q�ӄ���ǹ���'�<)&��mΧ��t�-�}�F;��r����?�8]��9{!:����Zf�/(��$2���=�Kq��Ji\*ዣ!�^�^Y�a|I���,+�sˁ�ҧ�/w��ITё�ݚw�U�ħ��J��/��<5���S_�3�.�^k{ $���qk�wI.��A�HUc�x6�N���!{	Ŀx��w5��Y��Ph��LW�˵C'�-_i���@�"�i�^����iZ+�O1cy���_B��?�!�W�KC��!�d��Y�;!B�0���N���W�g��O���1��T����@&%�/��/��Գ+�h�E����T6>����⤺;ǚI�h���c����d�����J��3��lhB��~d��|��j@o^4�'��	��ꜘ������e�������3��������0�����LuyG��r�������f�L�ɋ���Z��sqz����\G]�����^��´tH$"�s�]߸��=n�#��1�W�/�=?��JƕӔt��ڐ�z��M�K2`��P\L�`˞^�T���//�َ�9?R���z��d�׌�g���L ���&P��]7¥��b�/Jf�w8���j�m��p�����ª%��|8�)�4�G�06�ާnyS�}�|S�n��v*nGY7�r��v�}��$������ܐ��X2e�����'Z�2��PE�UKc��?�N:r��/3C4n��+{���Y���QõAs��F�_
�zM1���ω���hߞi3x����Xx��`g�Y���=�����2ƕn��E��;�esĎ^���}��R�Sl��1��V);�mKZĥ�X3���	N7,���<_b�Ahӡ�WI�Po��? ����������
U�F���BR;KBX٭E~���W}�+1t	u���G>#���`Ns��=����@���7d�`����/�|(B�	N�!u�=��L�������0��rN�e�@#�.������>-ߔ.��� �a���BQ6�W%z�>ٓ�5$����W��/n�d��Gx�NV 3�M�;�ũg�ɼ�+�D낥�\�Ø���U��]Ϡp���l[�ہ��V!��ҥ!��Ц$��b��o�i�O/55��5:�6��\��!��Q��kV%�����ۙ?+�N�z���x}��u��.���b�5 l~H� D�=7�C�SY�j��u6	~:�i-lAt�����F���4�
��U������Hu�]����j�e�F�U2"bs0���ly�� �e��8Ӌ^iX˔a
�h�=�V�P0eA���ߺ�藻�7y�9����ݞwU�d՝�~M�&��`��Bf�~Kn-�	Ka�`�/����.�������Nc�gAe�9�U�[���.�s���� ��	�Ko� QM�����J`ؚ�O������%)�-�`a�ibVʦ�e#�:�[���B��ЁC����|;���z�b�3^>��©�x�p�`�G�)�J#��a8�*�'	�8����\�eI�q%K.����9�j��O3����%���ߩw��Q�m�z�i*��L�r:�Ɍ��g�n^Q�f/V���$���n�q]�5՘wm[����5�����q�rQYm,/l���|���넛�ɻ������ώ�/�=rC;�x��?&���%R٫�l���f���N?5ֲ���GO,ٿ����n���p��B��{E��tX=��TP��vYU��3���
��
�Me|J2 yl~������C��0k D.���C5�R��B$��(!'�v�z?^��KI�e�{�O�����6$p0�I,$Sw�p�Fyz�qq�Y��fs�Y"���Qh�)�8�.�����VE��6��Ђe�z��]|����̢R�mю0N�=	�[�iғ��Y��?�APK�Osrh'QZ"�IIǜk,\�>��o��ad)l��Ǌ@���aR�%�۳pao&_Vdٽ���5�K�טr�*���f�4�q�3MO�k���_�Z�@Ɓ�y��K|��)���!)��C������ʘx.���W�$9�mT̽4�H��7����<���w 'U�>FV� ��C~UF� ����ٵ��<h#��T��y�p������ω�ً�]w�	�/T���-	��� �+xz�bmU)B姭��^q��gi[Ÿ���j��l�Z}�60����υ���$�@WI� ����d��Z=��6ձ�aO7�ƚ�@�t|E������GCE��5��*_M4�����ƌ�X�
�h��a��UZ�h��d6e��r걝w©��K��>���Z�in�˭ '���?����ZT����\8���L��~���7D
b��[x� �zu ������_��-�u@`_<�n���G�������¶�v���2꺇a� d�|�q���陲��,����8h�kWT�w�hmY�C(fb�9 �5��M�]�kS��e}��<�Oܩ:�%�tao^�Y �b{��,N\3�
9+;�+&�K�#qwM(��
Uo!���莉E����I&(:n�vR)8%h\"C��{s�$ݜ)0�f
�:MN[_��9�T&1K+S�X&�{��#ug���<'g�2IID:�ܴ��Xm%�G��7�a�;ɗ�X�
X03Nw^��'6���1S�ؠ�m�5�L�ġ�]3�am�	(st+�|�/	�LR骤I���?w�>!��$�M0�A ���}��'���^�o"��Iy�&�ŷ���+�v��F����7�,,붖��?��G��
�֥s\�}����_h���2��#����KB��r�ZUk�6�z�Jo�P#�Ckb�������j�N�O��e'�x�ԑt����<��rd�oL>� ���#S�j��h�J:i77/��o���bd�y�ž��H� -�T��&N�G����E�3������T�!4y���=��P��*L�v��45�se��-N�K����?B�W�q�_� ��t[3��u<�7��HOz�&A��[}ڝ��erO�ڮZ']w�{�%Z�0?��z(��$�^���8�q��i����~�^7��@�I
�6�츑�.0����4"�Ӌ�f�5��U�|���Ja'u��65_S�KI�n!����� c����kb6%II�UA�Ec��y6͟���!vWj���>w��WY�������hfjW����ތ.-Z�:�Yy"{�h^�uO�
+�=�c�P���+�:{bԲ�C�Į!�
_�l;��~kC/�����YΗ�B#O���1�7��k8�@i�/�ʍ�{�&G����2���b6Y���F�*��;e����^�R�QI�N|3���,�@�G�TԢJ�U�e+�o�C�'�,	�Q(���9��v�eH 6��b0�m���4Y��v�F:۷�X��um�����L������g:i���뙭���i�z����c�G���e}����tÚ�N���Z=	�A��m�WF�y��e��*H��NV;���/뵜cM-�P`��A\��r�YƬ�,=ϡf<���t��t�R$�p�u�o����Gǽ��[�L{������\�+v���u/����2 y��)�m^fz���P��%N��8���4^���눔��Q�y��ӛW��n2�*���Y	jP��V�1��!|$;	ܠ�ST�����e��q�Zt���-�Evيcسo�����vE+>�h�{��]Y��Q>�s·hF��T��1�g'����#^�iN�>���x�g5}��{�s=�(�zפ2��n���GH;���s��qէi+艧m��S'A61��)���K5c����ڦNe	I,��a_۩A��^��CPJ�0?[2�\*������m1
54F.����H�)K}脭ࣛ��(弲g�+�f�	��6�#������\�7@���O�*�Q7���h�����(���.$uE�3�m�p���ic�����t��@�8#���!�`�9G��c!��2�|9ٽ�Y�2��y�Y��g���j�WYk)0���ӄ�
% �~��fRM6�(Ť��g�����Q�_o��%dZ�s�0��|}]j��p�SlhG��<=�q��M��ӽ��_n�bq]`�dQ/�L��:8��Q�\r^���O��S�%/:����?�A֒5{s��}e����&�&V�5���H	�DO�����n���ЫP�K~M�:�i(��57�TIX���4b��쎟B�Q�/uԡ��Uj��ۦ�LEU���s�۫�wI� }t�>'���?is��a��]����VC��uA�t����v��y@Z����
w��M�8�M��h���B!�O~f�A-��bK<�B�j ��t�v��'�4S c���A��q9-K�[�\�.A�����[C�d�8o��QhfY�Y<[`��O�IܭI2�%$��b%����V#R�U�#�5�[A޽� �|��3��;t���0/ݜO39�Gt.�D ��1]���GҢi)ը�a��8�{'D�F�b��WU����,7�.�?9ݴEF�駘3���N�a�g�:AV�I��1����T�$ɇ��gE� Ju��q'��8���Y]�:�Փ�Uw�"�ʾ���?��?�L����m������|I��?��֬Z�T���w��ju�r�E"�s
P?���M�u��c�l��.�ӹ��>5�K����O�!�X[�މ�$��#���@�Q��EH�gX8y-T`���181����Y�i���)OJ�}+yg=��ϗ�~�K�D��d��﯍}���@�#��'N@�z�R��f��e���*�{��(�E�0�;,G��+@�y8�q�q+�4[f��S"�C�Qc�1�fW�靘��&�께h0�s"���]w܄��R���K��=�[�i͓����a����V�-s-��QuZ�I��k�>��C��/�)g(�����CWiam�� b�p<ţ_�u�Vӹ5ӗ.��={*V�f8ӯC�3(PkӮe��4��;��ԧ#K7�})���!�ΎC�N�4�q�sߟl�JW�q�9
R&�8��HoFp7^��l�7ZS��L8�>-���S��UC��L���X��Q@��A#I>]����m����O,��j�Qنrw��=/�-��W�x1' ���zm��C墻�������[*���3'c�E�Q�;�}D\�����Jș�bڷ�[�<�{w��ƕqтk������O���)��[�|�����R��EI�?�Tt_��x���]�.����k��AkU� Mh�H�d�|�ӄ;���'�s�Xˢ���Zt;��Ʋ&'1��������T���7�����]�̣���W7��Ȋm��;�u{�����˚<.-�{o@[�3<�h����܉���s,0��f�v9Cq2�͐a���
�|������,h¨������n�m���x�bG�S�Pa�M+�Nk.Ū���=op7�E7%�����a��Y{�{���N��?
�79&��׆�b�m�q����尞o\�Y̓ME�W"���:)��vm��%�s�C�%{�q�7S���:�I�[��9��R1���S�
W&�h⾫�b,̯=d�g�E�I_�D�/9�XH�lG����6�����1�DN�����.q�� S��p� �
���m�3\6F|��	���+�6��j���'�-����?2�!49ᴟh�0������}}&x��O������N&���j\��^��+�_��̠�6�k*����� A2�º�پ���R�"���mG_�׾�)��ӌ
&�D��νUP�u�eo餔��J���;�:�}�)�G1e���x�T#t�������&6��Q5��:Y�^�UjQ2�E�7��&�}e<���Bd��o�dσ��-���!d�G�ٚ ��0"��qe��>��5x=�*�P���La�
�Q@I�"�����&C���mB��q�^i+��/����<i��#�֧a��0S}��?[lr
�̮up]]��{�1��k�+�?(<�$�����:q�G!iR���Yo�^rc���I���Ge���g?����4=����G����\U�T3�u�J�ކ�P�5�qS�Xڋ��_픪� ��v�k�Id��A�yc�W�6S�+�l!q��.w�^-Y��R�F�hAo�W5`ʵy�-U��ϴ��"6}^[���+�K)c��ŕ��5����C��\!�|�LQ;ד��\ʄ/���(���/Ounh1������@���/+q9�*B�!�S���I�W�T6t'������^;=Om��␰Y?���M�	���8[�)��"��KIX��X�`[Pos�'G/�	����I���)wTe�m��]HJ��ҁ�[�Mν�}ے���u�߻����Sҟ�%т��Ɂ,��thW��zN�@���9G=� 9����t>1��)|X�.
M=��w��ɱW��d�����Ef���7.���~��ȔMȒ�`��n\�D����GF<��h���0f��SR��"�p�e��$��PvL�[�����<m������/ �@���5���m�(����V=�%�8� 4�{����.��yI�՛2�nm\�*8�Y�B�(	$��ߑ<1J$�ae����R7�=�5e��)gN�Z/$\�7��E�|�c�����B�{9�_x�S{@�Y雙Q�rs�uoF323���1���?;6���7iiD��}ڮxZM�gp���=�����5�2y�Wn�KN��;��s:�Y�B���u�>E+S��x1�]!)1p�K"�m��A0�	DA8�^�_�GA�!��M^�P%K�?�����v����LM�
���FI^�8�� fK��d�{[q���q�r�+���	��W���#�J<�֤���b���ŗ�/7�y��`c�%��(�L,���u�8�퓮$��,4�$ώ��_�h�?���#>����E�4%˔��&>�����8T���Mδqӊk�8��A7W�!����w��? ��3��M�MѸ�ş,[gRl:���\�z����[�N�V��nf]��p�}Al�Sh���W��ܱ�j�Әoa��kdb�_L�/�A��Z��le�\��ص��7\�%ʎ����?ᣝ��('�j}�U��>��ai�5VAHu�D�8b��V�����`dx�+��~�*�:���i#~�*�����Z)4ݻ)��ZX�}�H��R�u�Nxk�jb�j��r�U(�qs�%6��85�V x���5W���"i��
a ٞ�Ƥ�V~F=f9�A�ni�p� �1`zy@�^��\�w��*�ӜM���[mB���~�ŝ-x~;K�4��u��V�����cU=�A���9�`�[i!W.|W�jöD��:eo[�FQ�#��Ԝ7`�Z"O!�R��3%��ǽ
^k�V>�a�J�#jP�[S�=�xMn�w̎פ;/�$��HX��3����Q��ȇ��e�M�G�I�)�&4���8��F'�	��"��R܂�lX��h/.��/�m��ñ3	�$��1�i&����H%���W�	���+ޏ�{����ɂ�gu�+��e�:��If��&���]��Վ�7w#
��yW��i���U�'�ǩlmb�{��c�|����6����z��Y�?2��8Oryp-�n��?�A[�����c2l�S�,��R˲5Gᕭ�c�O≒�ϸޤ�ɍr髒^�㌊E�rX3��T�V���6���a��ԻD|ю��JR�ybQKT��R7�f��D$�2��
z��l�x�7�:h'�)�z�g㶁�Ge���=�Z�.l��0�}�,�[����yS�qg��%�f��a"3�Q^��������L��_L�%���҇F�尗]r���w��R_�֎f�=�+[���0d��$`��9�js�ɣQ���I?^�k��>��)bɮ�@��"�a�.��{�p;�_̦���+�5���N)�*\PfSS�4�3q(k�p͕��6��/�UK��)���!�C��M{6��n���oW`ފ9%V`̳#@HJ�;7Zo��:02'k�-�I��U>H
��/��C��f�6�����f�fK;#��"�K�����b��I�فrBwVn/ʒ�ʗn�� ����t�m�����Ɇڌ�4E��Ů�� �)⹟}ߡ�������-����vm8��u��������x0���$O�`><�D�v�Y|;`�ǍW�O.E�쁽��_�V��I�ݝN�s���p���U���h���d���?�o�����c��}�w�F>Z-���ר'�{MߵF7�+əT������3�DE)a����7��O�(��V9�u�l�^������-IC!@V�<;��i�a�8*��쥣x6�vtY2  ra���2V�7v�����,�¨e����A��m�C��8b+�kT�M���k	���ۥ�
a2�W��E����a���Y��{{s�N��
9�9!����_����q��dC�ɀ�,�o�͇�,E�	����:�v�q%^�$C��C{�s��Ҝ>�@���e�[�,x9s100S�ܯ&8v��Y`�]t7����gSx�Iz.Hܪ#X#�zGU쿥�"G1�e�a�΋�N�(��G-w�_S���������T�W�3��i	�+�	���E��������WV�?�zj!O�3�y0����}�����+�%���&����U��9��+�w�|n��Fp��Hpaj^�b��=���������X���w�_!���Y�+���� ���(U��C�p�oD¹J���^��o�4C��e]�x��Pt=�f㲆"����ew���a��Xj�Q�@�k7�s�8{"���dY2�{�tϾv�-2�%��Gk�������K�A��,b��i1�p��=Fx2P��VL���l�=�����#�B[B-��q����v�ꨂ��qQ<��T��0㧜Y.�8�}Ы$��3r������]m$>{�]���mR7�(�($C�3�n��qګ(ìx�4F^� v�I �<�1_�����_�*g�o6�i��kE�U�L��Љ�J��l�݊�5U�S�����F�/z� ɶ���k��MIؕAB�co/m6C&����!lSK��l?wfWgY������h��Wp>x��	-P{�JW"�^2V�E%�+�y�c*��0A�0�8�h,DCJ®!,�U�a;�l�=�����p�x��O0�1��)�a6@�P�/fp|��(��S�V�@��*6���<^�sј;xY�94�T�-�r�Ļp����5����^�R��[�Boo�!'j�	V��	�Z#6d��e~/\��x�B%�<�����<2��m%��,[uJr:���]��w�Ev�ѝ�Y�����OC~�4�z韉�ߥ�Gn�����\�t����.�iK�=?dƵ�E�W���n��`��D9M�p~�+zMcf6`�;�\]���ω��bo�\�Yê
�� RZ+-�k��u85׽��2ddLq��ȷ�{�w$�_����/[{҂������mT2�{!�Ñ��%���8���4#��a��/)y�%����n�Ԩ*ӌ�Y�/���۠�����WE$1ں�rC�����ط{e�-�KHZ��&�R��El@�c�����Y���4�R���{��YG�Q4��sxSFn˥T\V1��Ϛ�n���zi��K��3�x5�g��9ű�=�63�0�24C_n��>�p�;�-5su<��v6�[���S�ʟ1��")�_�K� �<'Q��1m	?v����_�z�A�xq�ȘuP �?�}����x��Ϸ�L?
���Fd^���3��U�K�hx�3��Ӟ��h�+G2�	�&�,Y�#f*��,�m����[��B7�z��x�����(����څu{���b�&���Z��٪��!���	�#y�4�W�B�/Qk�?����D��kٳ%��g?��m�O&��8�W��S��:sc��� �vz�4U�Ml�Ś�g�mI�A,L���ȥ���)�l��C]�M-p�
�l�$۲�����T�C�(�sQ¦Ո�b��	�Z�'/Fۥ簝�ɇ��\h�}ؐI4�r��%e�|���N?<&�����:��}[�w�dv�Ӝ��5��3H�b�D��t�鑤I�����!~�h&:P��i7$��4����ܵ4XzK�{豟� ��e��uʉ��n[jR���_U��;s�^A�:��J� s�C�c��>��i���a{-,���+V��q��A�2��Q����y9.�P���n��wb��nNM�u��q��B�֏~�́-�h�K�27���W�����P����c�A���9#�*[D�.�׬��>�1��oOQ� ��O�`i��O\@��N%Ah��VY�Ky#E�%[�M����r���;���vjө�3����	�z�3�Ɋ�q�mGH])�x�Wof8l}+'�3���V�M�U�ǘ�G.26ݪ~�����3DM5���X���A��]t�$���i� ������z�C�'�}�gУ�w��J�g�aw<��Զ]�ՉԵw~��4J�!�:=�(n�mm�m���6Z|�+�뵴���b�J2��\'���Vr��i&?7�;��������le艿�׍��5�{���(O=���b޿�v���7�m���ǃ�E~��X.�T
çUա9�	��z�eO��J�t*y]^�2���K���AD��L���ԯ|M����'3�zp����Me�	Ń��ﻕ�(�0��,5�˛��"yn? q�B��f$��"μ�QY_��k�_%�+AǕ;��q����8�K��]m-��IR�?���(=zN [[ɳ�kNg����~��\Vs�*�Q�*�I�٦k���>R]H��*K)]��Ǜ���a�����Νp��N_����V5ɏeש4�*�ҌfnOF�3ޱ�kIG0�0ܲ�1k�܊�GK��+)�'!�gCC�*��?ҧV3i4��"msWk9@z�.�&H%T�7��ƕտ,-���E[���>c�푈�iFC/m��Ѿ���)��U#�c�=������{���������|��w�P7/��[�|M�n"� `�+�m&���7�o֡�G��`y��)����rX�}zu���� B��Ajّ(<�q���e�������H���e�OH�F��Y�1|�l���&H��2E(����_^��tl�d��N�������U+N�h}�dG�i������*�ic��X|��YaZ�>z���'�_�p���F0�TB����nl?ॶ����7U������q�{uqғ9����U-�*�@Q��<��n�$y+�SI$�i��S&[v���2�R+a�z���Z����,^:��@�l����H�KmL�Tybb�����gSM!a�k�0ۣ�{�5j-��{;�V�a��Yqj�{VdzN��
�9�:�<o�|��q�k���V���+o��͹*PE�ۏ�Z�:�Nyv�E�%��C�	R{$���m����K�[��;952D1��Sa�&s���4�X�>���g�`I����%�CX���G�$ҥ2b�,�i�@�i4NȽ����R�S:B�>5/����Ĳ�>3�����#	���+t�<�����3�雟&��>�?�nF!j�� 0i�4V1�}�a��W������z��&�g_�`o1��+XCD�ZF���!��t��6���c���5�Va��N����_y��J3��FH��Z�ܾ�#�`U<���kto��w�tjB�)܆�0jG��[�~1�e��x�t�uh�m1\��
l��'۱��ԣ�j�AZ�;{�7H� ��L�+{\d����V>���b-��-��'Gƞ��v�h�f�o�K���5۫�&=��tP��L,��Ƿ��X\>�AD��F�Z��Bȁrq�ç�)ǥ�� *<,C��џ��f|�}�b��g�r�o�����]���{��]��4M�|m(��$�B-�)��q�/�iH�؋=c^���I����Ɵ_7ā����3�d��F���{U�d/�+��J������5Ќ�SpҌ�za��i
 �,�,Q�k��I�bA�*�cJ'_6~�al3!g�����w!pY
 -�<*�h��bW�<���}k-K��j�@"�82^Mqp��c+[�ace���D��+�����C�!G��п�;�e� �ʺF��&��ӭ�O���1�����@���/����`/�u������B�6���巽N �;��a�ԥ�OiU�b������P���؏�����/&�V�o�1~'��~	ќ��5Ƞ�מew�곬 ݼ���-hս�rg�Hu�	xu�$��{ʊ�	=�� �'Ѹr��w#��*>�o�z��ʩ�vG������0�ut4��ߧ�ߤ��=��,���WW��)�H�{S��Z��K^-�f�M�Y�`��}\�)ˊ�1�}���! Å~�%"R����f�eЩ��x=�M��L��Ȓ+/�����(�����/�d�c���&6m���Vsk��7%�8뉅4o�-�AЁJby?sޛ�&n�l�*n,QY��[���]�b�Q�r�$�rܠM�a��]��se�jiZ��U�mm�E�#�ciL��:3��GF�/B.A|{�o�Y�Q���sSQ-F����<41����G�T�ai���s��xbg�i��LR=��ߋR�2�*n�mw5J;��s���x-��z�����SX��1�U�)'oQK���w��wS�	:�4��W_N��A����C�yP�~�?c��-p���"�l�
A��F���.�k��pK.Y���*E�Ή����+ȉ	�sL�I#A*8�L{�Y��_;��7P�d�q��|(��:��u�
퉐���M��F���^����_�#�����W�*�'��e�!D��R�.����h��*�㊡�K��O�Wj�"Z��Ul����Y �"��o|�M�sŕ�$g�8��x�����:��9s�A�];�$p���ly���md߹U���C�NS3��rbB�U�/�R*�k �ɢ�\����k��ǭ��% 2��'�?���f�Z�U��}�'f�?δ���5�� H�pD`��/(����W�Vk��ၴ~��:��Iih������0�4�Xy�V����i�� T�u�-o.��j��u�)U2s����u��� na�O�ۋ�7i�O�a���|�3V�$z��A��W�&�ٗ��MyTjx˽Z�I��wA���	 �M�z��̃PBR6~���-ns�K͌I����E/��� ��Ea�c˒fAї�9��O[�.�w}�T�#��{�uo�W�Q���ʽT`D��O��;�
C%���s5-��Vt���X# ��[�Y��(��mG-�DX�;�i]�I�N�W3ʕ��WU�z���ˏ�#�G��)&����j8G.�'����3���HJd�"?g�],$.9۠�%K��z[T3$�`ب�l��K/��!���6�Q}���]{�� ��xE�g+��=�g������R���Z��]T�BՄ��w�8I��\E赍���݄w=z�m�mk��)�|Z~j�pR��'L��*��7/��r�%̡d�5?�|�~:���l�Ob�dr�����5}lY��U�O��e�����
,��n��H�i���E��X)�Tq��b���T�ٙ��M��m}�96 J� �yX:�1�ȪX����D���R��>����-��'_\�z+�W��9Meuyك�S���$�ju0���,���\�y��q]A ���f_:�"i��QT���wuا~!�)��B����&������&\]h]�-� RՄ쎜Bt=���[6)������2�yٓ�+s^��Q��OI5u�k��J>��x�QX�)Xkx���t:a���q��p͆|_Bi�'=�5�;+�`*�imf��}w.3��k�ã��ߕ�,�&��J�Kh�()i�!�Cs��i�B��dvߟ}�WW��9[�̩�yH �7�s�p��(!���lA7�>~B����D��Cj
إlS��y��ڎ#z&OX����%�V��� �Ѫ;��w�wS�/@Y �����Y ;K�f��m��Y哥·����{i�Ť��ց*X�}�ѐ�8،[q�����٬H��҂�@�V�Fm�<9챓iXO�G������|1���}�����E���a�_�-_�����N�D#�q7;�M�U��hx�}d��+ӵŅ�	(ȩ��3�q���wZEpn���!'Bd��+F��a�DT�����_���aN{B����f7����Tƌ��u�0�a��K�7-2�@L�(<�1��9�n������.6)v�%2Vża�x:��@�����Y�,م��dN�W���㦇mݶ�)bxhf���*M��bk��K�Q��@~�(O�HWуI�a��Y�KQ{1u�NH$X
o�S9�חu��7�q�t�90�v�*o`�TI�E����+d:Z��v�9�%Tz�CrpP{_ؘ��-�����>[K�9P	1��eS<��&���)�Sd�N��g�=I��GܠX�X(G�|����'U$�ĥ(DgN�rV��	-��Su�ٵ�����]���3�pn�-�	A�+O�ߺ�h�閈h�G?c��!�z���0Dyf��}N����i��/�54_&�<�ۨ���o�+��č�eנ�$��|�ם6�Q��3�Nj��֑�-��%����,_�T��a����)o�}K�^=�Uה1�f��o�a��/���D7����˺�X�֫e�Y�x甀t�T��(����,��["#ی�T�j"��6&_7������F��d��1���4�*-h�fG!��1aBց���� �����j(=|s�P��rLr�ǻ�#��s?쑋����$�����BczBq��vzm��`vb�3�*<��]�������}�9BPr;�;��;�]c��{h��mK(��$�#���q�oiï���S�^#��A�I�3�X*-���(^  ,�?��C�ݡn�U����؄JM��_�5KJ�SK?��Z���ey: �^���+kN-�I���A3c%?�6�,����Z!bϜ�?g�wܨY%pv�}h�W@W�Z0�Jc�-F&��Ś�"g��^h�);BD+65Vc�5W�f���&K��_C�??!b�K�;h~vWT�U}��U�.��O���1*�u�WJ@m�B/��~��U�og�������6Ż��2=�)��;��ɝo7}�J.���:{����C��2���\��+��Q��o%��'x?�	7ڮ��)_�;�7�e��b���[��Ҳ��*%��2��#�rD�	u����v�d"	�w�����Έ�Y���|z���ghG$��Q,�Kb�t���m���-�=u�����XW���@{斀ڕ:��&ό�aM�m�`�)_\�;�E͐��!4�R���`$`��R�J�a#p+;��3���h�xLg�k�m�ҷ�H>i����/���_��f(mJ0�1����`%�1�8�q�4�����ׁe:Cy���ã�n%$*	�Y�u��9�Z�A��$'+ʠ(��!���e���x�>Z`~薈m�Eb'�cD���u���ۼ*a-���{q��Y:��Q*�
s.o�F�]G�=*1��V�P�����i�f���F�x�G[g!N���\=��.���2�6�n/���;_��s�����u���O��Sԙ1^)��XK����~��U	5@�o�_	�7AԾm
P�HO?Gh��T��]��
�XF�BS�����>Kii<�LBC�ɔ��Q�+�}�	��r"Z	#J����L����������7�_,	լ�7K(�M�u�u��B�1я�q�U�g/@Y��Nf�չ#��.��.��%	 ��P�ox���1`٩Ƞ���3�e�y�<������W� �:�p��v<Y d�w��ZM��<Ő�gc������˿�����߯i�|�]�`�p���l�8��(\)�݌ޱ9���)u��K#bݯ�P�n/����&��ɽ�0\^�F���4/%�}�����?�t�!���pY0}Q� �F��c5'q�H��hD��s���̑ډ�������~9E�:��i	�;�2�@ȡ�D4NW��1d�.���u��)���j����U�QTs]0h������4 i�� ���>gi���aq6+�W�V/�V7m&A��߁d��bN�yoưF���$iiw|�{դxM䟴�'H�BV�~�:�-�K�l�V5'������N��Pc�m�A��-9a![�/�.-8���`������)lo��+Q��E~�`j<OҶ���<%-1��z��ݴV��GA##�`[��I�)�h�7̟�!;`�?=��6�3��H395°����(�'��G���)Aaz�M��8"�'0쉅�Q�C1��}���.T�Sݠ7��U��3�ӕ�>������ (B>����OSX�6�@_�yj�s�~g�����2�1�]q�-����Ξ]�L�D�w4��ʪ��!�V��Ӹ�x�m3����<�|��|�+ �B���@C>�W��VB`rJ�_�_�:?��9Q��2$2lu�K�?E����5b/���UO󂏢D�T��U�x��#x��=֯E�I$X$��T�����	�oҙ�L�Ֆ[�tz�J#�	ySy,\OEσ�)����D��d�Z&��y�#I�,��'��>z�e��E�e�Z���$��=�0Ȝ�,�X�ty��q����BGf��"��QOk��e��B�D����k�}�ڇ�s偞�]c������R��ݎ��=po[�ړ�$j��l(t!dsL�Q�z I�0Jks�	>�I�쥽)SlW�Q��/F�aٷ����p�\:_}�j���S5��_�'*B �f�K-�Ȼ3���k�_��f��'y��@�lK#��)&�!��(CN>�����S�_ؗ�؏W���9v"�$z8H��>7& ���#N��>�~��+>�����*C��.�h���q��w��#5	�s�r�w�1���;�C��W��r[wgu1/�{��c�d�� #W�� m\��3x�%Q�ڽ~��y���r�S���}�2&���������N)-���[�g1�
VƁV��In���O��7m�o����|��n�X�9�>�UE����P�_�ֲ����L�L�X�~�Ua�shsp�d����p�f�$�ͩ_����֞��Z��ډ�'������-�|^fT�6У9��vq�)�~;�7W��YA%Ƨ��ug�;���6ˆ�M-Z�@G�G<L�3��䊉�#q�_�ϣ	fGv%0	2�W&a�^��C�+�h�9��,T�J��>���&��~��m�j
�5b3Dʞ��	M�,k�L��	
���#�6�R�̯�a�T6YgM;{�N�p�

��9.g��֏�s�q����fU�Q`�oHs
���E��m�}�:(�v�M�%�SCM�>{�:Xݣ9��w��{{[��9kV1wwRS&�]R�*>�N"��A�g���IˌC�/�X�5�G���hA{"��xP��4N�G���P*�S�(��t���A��h�
3HD��P	��+*BC�V���S��鑑��ho?��!�%[���0W(�C}�h����1�6�����&+tB�Vv����+�k��M����Ç��cw��H�l��ᮌE���̟t������U�_/����B�| �i�\�����Ur���a��oU6[��	��_jo�&�A˕O���e.�x│tNT����;��nB�֧��gN��J$�j�Г�1��7���30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�%ڜ4�z^��2�Z�n�;:�|͚�<���͟E9F�_6���(�(F��Z$����8#lfuP��Դ�I��O����Ŭ[:v�,�82�B'�l�(�,YB��F�2�%xd4��o����C�ƶ=wS�%һL>[q
�\�������� �1}?M6�h0&�	 Ic[:������  Ll|�A5E�Rv�/�h��]��
���Y�������le5H>�Q�핥r)�Z�Z��7�O�S�h�՟ހ���Ii�}��ϥ@ʼ�n|�̕�U����ֿ%���T{�OL�Z��m�:f�"�S�T*����	Z��?gj��f�LoM��J-"m��<4�Ӎ�y|����Ձo�3t�A���' �ՖI��G
cG|�jS!�#���W�֐��7�N�In��:���OԚQ!�#�q.$�֤RѻB����:�0uϹ�Q4 �yZ6����?E�>|�tG?���
�9�|��_��g�e��ːT�g�u���G4�xL�ȉ�%��>�!U�����TqHb������M��|�_�P�1Izp!�:�f�
��.r��e����#����T��UIa�c�P�A���I穼���j ���M��i�s�ř�c/�ߒ-�Kv����}9bx%1Cg1^�h�O���B���d�Сy� �0�bX}��g�Tt�X��D�����S���L��	5@oL����J��c��NaÀ�N���-[�U�V�wa�o��v��ݨ4[����c��<d���P��U�f(q��G��*p�aX��lc�C7�{�T�tQs�=��~اp�OΕ����ka�U��ޫ7��=F���������r�����8ʣ��/ ��܁��{#us$�?�Eu��7���i�����?j� 8$Pje�W��b3���~H���N�>O6 +ÂKQBA��ˤ��� ��~SkBc�2���T�&�`�7oOy�E�݌'P��@_ܩ�� ����"�-r���Tj�؜�ƭ2��<xۥ��fj88w�_v�.'3.� �QQ2_���H�~D����(��������)����ѿG[ :Y]�R�沌g;;1\�>���g�r�&�G�WYD�>�Ґ+���-�x3�i4�b���2"˦�`��#D�s>@���M3?�/�(���w�Dr?}�S�N�/n@��_e�6K�2x1�H���S{(��Q�v�u_Nߋt��m�d�dN�h�w�������8�\KX|O��->���xV�9�9�¢x��p��Ke�%&��a'����?�Qe�9�N����JCW��#k��Ǔ�������N���+N���3�IK`9�z�jF�v��I.�/��M '� �f�ج�~nu;z����<g[�ԫ�:�L��w���/��H�u~!3:P��G��KF�I5O��в�P&+�g��r���I\�R}�O�i�T���V����:)�H��lg\�}����a�4�	,�#
�)�Ţn������4zV\Da�dp��Y����a��f�EI�>�����URA��w[U���Sy�����d��y�5q����gλ�j�[�K�1��I���~�J~�C��|8�j1X��a�|�MzM�9�+1L决ڷ|�\�h�	J��H񎣑U��R�Zf�M/]i	v�V�]05C���kL_��Pt։��c �����k*�NlZ�)����0D�7O0��xu�k��k߇�s|�M��|k��Eㅆ��Jxrʝ}
�F�i���\�k�٭�E)�)
UB^R������W���Ҭ�7J����:��,:Mc˃�($��6q�$ڰ����2���t��,%���7��W���(��0g8�#�M��e.>�y����(J?���c����ˆ�vWk��>��)۷�<���S�����$�`X� u%i_��� A��e;�x������?Ar�e/���:`��J�c���r�0��~_k������-:������1LR%-��G�zJ���c��C���ـUx��a�@�"o�:�lһ9}.&�C������H�OL�;a�ߦ�~�3�"�[w�;��<���q�Ә� [ U��H4�韅�;�����$���L����lV��H���m�B��ƨ9q\7����*�#�����簝��3(���T�pLOբ�k��'��S�Xj�I��l�����)�cA�Ü����=M��QU�#+��僎���m�V؀��7�ɔ�V1{$��z��0�&5!��6PV���;�h����MD��%�Q:1���(�������T6�}&')��hV�	�N�B�&B�ġ�ۺ
�r��z&�}�lB$hyO�lNx�tW����Jl
��o��Lm���včd�y���W�q`\g�w���E1kS���dKK�	���wo��2ƾ��b��1�"v�^���_����5پ._+�	��Й	J�9�^����-)H�M�l][�-:A��>&k��ȿ=C��R˟	
r
r�S;�徎j��ô��]��'�DسH
/��#���wb�=�~Ec*�������b�8�ost3nG�wp���a*�����j<������$ǥ��w��_|G�UɒJ�Rq�Q���{X�����)��k���3�t��h�?��7Q-�_�ڮQ#��M��y+�~�,��މ�\�Ț��<A6�8�$z�G�+\5հ�=t}� �<|�7�F��c8�� ]~3ʥ�`)��Q�s:����Z��R�����ֻi��q�/`�1���~�j�R�%�nC@��샪2�W��~���]��1v�qp�� �+�z�*��M��}~<��]2�HF��:��=��rm���x1�ȸ&
@�s�|����F=�+�:�Xj�]w`��ŉ�A\������_�q	�^�m�FĮT�U�1�z�I2/�C�{/0�(E�*G�m��q2�t�?�,3>��G㹸�.S�� 0_C���$�ҵ6Tc��u��^G�,bL�$����j�b�=!������#T���?�}�Š�����mS3!(8�f/���w�rܩx��d�G��`�ԓym����eQ�]�ɩ�������oM}6�Gl�i_���?�Q`-��b�(�����b�LC�����	��=B�YP��ɯ�]�0=sb�Qǋ�t`�6Ն�������ک����� �B�@�h�6�&J�$�L9�a��N/�-����w�ă�M�'��[�9��@Sc?��di��C�y��(s�G ��pd���c�/��~9��x/tul�=_!�~)�prfŕÑj���a8�V���[�=�s�5N1;	�u�SK����G�/Dg �%v�{G�$r�E�I���pȦi�zG�3�����D�$���{���P�|��|�~�<4�1����u6Dc'�&��Be��H�%�D��~��Ec����Ð�J
��y�y9�ˁЛP�=����l���,�;"G���V�X+jk�\�>bb2SЄ�7'�7�9j/Ffwx2��8�����J���lw��U�S��6!Ar����k�Q��:�(�@ϱ��Q�o�ƔBX����(Rz�<���6�!;p��䲑�$T�K:����)a �h�  ��D�r-8���������v���U��>׫��/�s=�����Ne> ��9.��MRi>�##әP�]�o��[�\�9ҳ��2��������ߜƬQe�k]�dC�'��hf�*�Y׉�i8����TD�eFq*d�7y�6��?�$��5��ck�W�4@�����!Lb*1m��^?u�dD �����O�|��R��w?L�M���ޒȽT9@�'��+��"�^���f�Fj���2f��s�b�/ߋ�m��PD1�͢� �"��&���T�x�3�E��\5l�*��g�� bc<%�,����񽰿Z��;�"�Eꁒ�����o�*aܧ��>(ѠZ2ܿ��Zl{��S����՚!�@o��O��	8}���_B2X+����Y��F�W%$����o�{���o���� SVI ҆H[�>\
�oH�S�� .D?X��h���	��[eT��>g��&l��/5�v�r,h!E�QF���6VY$����ţ%��5�I�\�rXu����۲ΐk��*F�'�hGԦ��s�h��'=�%eeGa/�������H�\�n�n�q�7�Y�!N�v�8��?�b�S�.�-<���:ӹ��u���xvB��[�DU�{�çR����ѿqk��&F;Hh������7W�%\޻=��Pl��mSAb��1����*�rP6!g��vb'�Foo��n���wl����4M*�G�~� <�1�ۙ;���3�Զw�˼|ÚNɎ��aQ�?[��˄��i)F��g����W#��sd?N�Q)���V��#�ٔ��ޥ+��7,�;ޅ���D���8]��t8�����+X�p�`Q�}ң�<��\�i�F 8�x]��Yʡ�^)A����rs����/x�a�v����7��m�`����֍��	A�!m(C�����`���z���ߗ1rZp�'��z���IG�����~8e]���F�x�@��n�1�H�[��I�
�V��xT�m@�F9�+e�tXf�w�}͠�VSA؋Ɠ�}�/�+�me���{m��Ʈ�Y���
B���{2+��f��$l1ۦMgm�y|2
?�qK>�/G�-�ȪF���x_�S��N�T_u,`jG���L`��ņ���3�!��Y�{�T�f�>�1�y7������鍷!$��f�ce�s��rX�M��3���k�\�����������EY�֩\a��
2�m�jMyV�	���eaC���-co�$����b%UC%�=r�&;��Uƿ�pe.��9�0�� b�F�t\`Q@�pk�h�ᯝ�I�V{�I�@O��2W�Jf�V�H^Uac��N+7�-��l�6�wg�I�H�}�X[��;�d�$c;�d����������(��G�� p`�	Q:Hc��z��ҵ�3�t�=[�U~�Spn?%�?����<a��Q�{�c�ק�=���-P@5*����7��C/����!X}{�0�$no:E���s��K:i��I�������q��j�$�9m����L�m�I��~��C߉;���#6����"�~B����D� ���;~��cff���Y���_`��~By����}P:��>:�I�������3T��!����jg��ɺ�S2O/�v2�3��j�;wt�cvirO�� &��2���_DWy�x����"=uD�A\*���l�v�B+ ���K�̊"�~��c����������<y�����xP�����ܓ��JS������A��8rj�yɄ��2YCLbݥ��ju#�w~��v��w]YA ��t2	�<�2��Dᡈ�o���&?�{X,
��]7�i��
�tY���Uf��@1FNh��ѷ��L�zG�>�Yn�ў<��+,H=�"\3H��41Q��p��ː|�r�+��@ɒ���H3iڟ�����E=�D\�� ,UN@�$�e���:�1��-��P�{�o{Z�����5	��W�玵KhN�ʚ4�N������K��5�F����#j��S9}�zx�JE��Ă�ae��
=���ֆi8te qNH�j�4����#K_�����mt���1�&�G�NT��3�6�`c9�5:� ��I���:b� �j��p���ue�����-��-;G:�e�����P;��2Eu��:�!G]o	Fl/�O0C)�Z�@�gӷ���#���\V��}?�O��]TZ�� ��zOa)ea�9d�\�b��S��k{͞�^��Ui�)��n��z��z@ 7�N��|#���������0�b��/� ��
|ۧ����UL��=l&��Y��|�5[l ��8��js�ZK�n��E�Т���î𽪷A��8[G�j۩��KB�|!�������G��p��������	���H�_c���RT^��OKi�V�P)5�<����Ug��ɦ��IxcʮG�|\�kT�lĹ�ki���0n��O���x�I�P�k-����{��J�|U~aE@og�+�]x��?�g$.
�׸i��I�)T�æ�ES�A
�y��b�O8�r�	(/�V�?74,�5s�Y�O,�]MMs�T�$3�qW�����\�?���>,�rJѷ)���|�+=���������f>f�!ˉFJ)�\Ӎ���*�놞"�kr��h��?���d�ZG�N"^X,�%:�݋��-�mEh�Dj��"r�2*�4_�:
l�4J����r�^�sb>~I����Tg(HZ:B�Ο���L|[�k1�$�'��Z+��$��*)��"Da���"��{�k"9�*h&Ϯ3]�&ᓚ*ӉؚpIP�P����������eQu:�8 d(Pd���/�5�}'�M��m�J� գ�-Bz��(��
x��[�e}�BIBE�iOI�oN�j�W>�&���
�e�o�rn�˻��dʄr��z�WCQf\��(�8�	��1l����d��	V���?,�}*�s�B�4�1�E�vX��D�EuJ1Do5'`����К���Z���|�Yx�����]qSi7�������!���av����{u�\�^nY�b���<���I��"����+_���L^�C��p]C5�q�S���Y�p嫼��0U���V�2��� �o���BDJ��C��NJ�'(�������J;���gJ�BW;:gVV�_�=%� U�6l�w�O$�u���lD�<����__ںdN��v��V�9LS>��l��__Q��:ݢ���9+�'U�9Q~}О�?���]T!�<T�=P����؊z��K�+ �u��-8^Zi�#�e��$� ��[.)� ��EK6J�&Wl��z)p�[;ҵ�����2䌾�>��CC]H�z�����dE��%�+��2�#�^���?ǸNh�Ԃj��XsQ���b0���U�y˱f�S�E�Q.uL\��7�Ȯ�����s8���b<{�ޞ|8�.a
��	@(K_��E��=�)1N\{o� bV;��Hl�=kU
��7E҈CcF��(	f6y��x��nÛtIU-���'�#J&Ek/%�g���o�|��G�W� ���s*<s
O]��8/��z4��ρ�1���7	WRi���<��F�7�Ώ0���� e��	��WN��J�W-oZ����j���
̖��x{�}��5U�P��� 4�%r���-vhI45y����k��[���8H�2�z��̂r�$�(J+J��j+l�ɽ
�-�e�֏q�u�	{��vD,��J�ꍯԠC\��}��2��i�
��;��1���<�(D�6q��2uU)�4{I�>g6�>>�2�;7f_�{5q�f���C�8��5*�K)�L5����vH���O�8/{#	X���9�K���.{ʝd�\^�V%e�f��X���}�Y�K*@I/H��St���[Q%XH��_������=��7���ෲ�Z�����-�c���b#4-����d�	�@Qd�"�TF��!7�?x�L���=Q�B?}���f�@�ǖ�Vو Y�nq��ie*"{���n��7fkiEK���x���x�Ra^D��CG/8���J��&wg�:�,�n&��ak��4;R��g�����p$�\ຍcBR�"�_p�1^���gi�*�xу�w)��P,�C0�,��t8V��%g~�lN�q�wks�ԮVA��zat�ȬE@>Do��*,���׫/�,/A�C@�� AV`+�~?�U��c��NY��+�����`�([��ɢ2������m���,_A���v6a`Q(��Mɴ��Nt:����JJ�c}��Bw꺤�1Ǘw/��>��
D�PG"C�J��睈'����3��,�Ҡ�q��
]���!�Α`łA��Hj$�P�ʏ��)�Xn��;M��+6.�}��~9��Д�[J'{5���J$��&}�x`*6����H�;�g����"�1W�)�V��*ζ�ƹV�ǣ]5����T�P��e(�"x[��W�m�!�,^]�$O"�,//v.{�7���r��U:O�A�;KD�!�CD���e{ �7��<+�A��D�%bLͮ�>͐D2���}ϋ֖�˵�l��	.b�L�9G�V^���b��W�"�n�m�e�N�;�Ŋτ:Y�Y�V�{95��p>�=r%J���Z�o�zr�oD�r/��D騚�R�33��ߊ�渗6⛖o�����# 4b�R����vZd1}o��ԬJ�WC��j%i��/��QN0���y���:�M��	~YQB��>�J{V|ZU-�g�4�y�F��Ѓ�KD$x�3��S��T��:�Y���&�G�7��`����S)Kz�V����d���-�?|nؚ`�l˅�i1��$Q�e4�H��~��-k���Ӷ������Ӂd��ʈR�/��2MW��̖�.k�߃� �5�y�D%��*�Y%�A�6���DP[�õ�Q对v줦���D��n:�� ٍ�3pt&����sp2PS���㿼���n<�S��N��cퟩ��.�iNj����@����̠�p���f֊�E���/��wZ��Թ���"x�g_#k�X�Zn.Tg�"�f�Io�9�Z�+�<���a�z<�c�A��L�����4����n)�'pmIAV��@���\�e�&"e�/� �w��N��V<R�;��7hm��������QE}�%I( #f����2|}��ؾ���%��s%�BJ����?
H=��+C}�<Bu�O>�N�ժW��ػ/Z
P��oT�7>���g2?d����ɵxW�\�����1(1<���d\��	�`^�Ȥ��M{�C���',1{��v�>g�A�P3ys�꾿-u��B�j�A�*�����)#z����K,]��{��n�ܝ$&\����=@uZ��Co	��r�BUS����摒��ʶ]���Oя@*X�r�������HZ#�;�I��e���<Ez��I�,��P嵙٭HZ��f���jqp��^ڪ�=��J&OR|��� ��PDkNy��w�s���t+�x&�f���8�xWES�+�!~�ss[���S�����&A�M2�<�^oրI�ϥ|x�m��quPC�^�����M�ȹz?�U�̹'�ɨ@�6�u?%�Ŏ��<�4i�ZUr �'֥1,��^y����d��©�4�R��d��["��:BC�ʯ�����<�F�8l�=v�R^^�c����mώ��s����`N��K���o�B�u۬hZ`K۟-ka�ޡ��o���W�Q)�az��a��B��I#����zÈzԏ�������=�"f�W��BR�x��p�T��"������~���Y�ߧ��� ���A��{bp_�x��Z���u�	�+K�eʬ	{S�e�T�rr;!�A�(7R�`Z�>��S�k�A`�f�.d��u-	�n�`Xܑ�g���wDQ�BI�ݻG�w�G-��e�H�p �LE�(�N��o<P��̯��k�p8Z5����"�YwY��(�/���]0�����/���B�|����n�V����LY;&�ߞ��A2�Q׻*���d3�n�S�V���U�����q
(i��1�Sޓ@����̙x!��&��P�W���SH/Z-y޹>s#"QhX�p�q
�Z��Fg��f!��o��\"��!d4�j�ӑ��|����7o&8Ct����A�� ໱I^�
g~�|a�N!�kt��[g��y�7��CI��>�l�`�U-�#D�O$�#X�(��Fr��y���0�����Y#U�¨�iu��F4����A>�uj0ǩ�U�?r�\�!U��4Dk�'��Γ�±j��E���e� �ZWX��~��	~�P�7�ʎ�;�<��F��}��P`���b)�+�h =�H��rA�<�j���vT�U*�H>�64��iñ\� �փ{X{R<\��칌a��>��'#7�PwF�o��<��H�9����Ʒ%���X�<�ڦOei��xx��إ�|JY*p�H�ۢ��$��h�e�֛*,7�6I�?����CH��|W����ܸ��@JL��hm�_�?	��D4���Аm��E�ڋ_�L Ⱦ�,)��&u[�h�?���v����^3� ���j�Z��t� ���-�����$���s Xx��:�S�^�x��_E4�#'�;1B{Ɛ ��%�o�9F���TZKB�;����r��+�D���>_�M_(�Z�٫�kl����<���dծ���Fˬ�w,����8�'+��?fBF�6�'{5Y!=�F�K%�!72o��}���`���wS�B:Қt�[0.�\Q�� �g�6 ��?l�h/��	�ߺ[�VB�'����l��75�Dv�1�h���e��r��Y8��~=��9J�5���pv%�j�Ӝ]o]�3h�¾�s'����:t�s����B=+��c16�a�"�M��p��p���#����0����5�@v"�5�S�����.�<~�I :���	��$?�v֚G[�R3��c�fdS�v�q3caú@�H��;~�����u���-����b6����*"��Jצ��7�b;�Loףn׋�w -���)�*J����%O<@��ۭ����y�H�w%�X|�ci�"\�}RQ^`xɌ��aQ)Z�u� ������}��?�#Q����j��#�2��� +Su�,�|�����XǱ��ذ��A8.�P��	r+�ްt��}f�G<�̮_�^F"�78�
Y]�r�5��)U��5Ls�/2�R�u�׊�E�K~n�n` ���Ef'�����1dC�<`��=t�����	1�p2Z���Ɨz�����㑞�V~̧�]�uAFITF�T:��k�\��X+%
�j@��#����F�P
+y�LX�ܫw�P��U�A�sד�h�C��淤�z*mt�O�� W���b�
��2�+$�x����ۺ�m/��2 �?�O�>0Gs��Ⱦ+����_�͛��۫bV�T�H�u@ęGh��Lt���YbF��!��n�TT��R/>�@��0���a���!�&�f�ZH��rl���5����e[���	�^��z�����өpA<����M.Nĉ��m���D�-w#���V�1��b�P�C��՜��:����l���u�T�	0ͫJb�����7t��e�G�B��|?�1�]�j�
*@#���_,Jz�����aw�VN�i�-v�0^{w���Α�f['l�x�jcϚ�d�Q�����	�(�Q&G�Zfp��ec ֘�/�����tI�=�F~�� p�i�S6�"'�a��������==zr��u��I�8�$�K���׋�/�c�ܵ�{�o$�GE)BkJ����iP�u��3��sҾ��}�$��������İ�]5?~K�ߝM��rxZ6��ö��B��������~�7czL�"C���k�yɆn��jPN�tG�]���T�(���P�a����\j�����i2�Jy,��� 7j�vwu�v}��g`� :�P2������>D��㹯݌1�i�EЫPQ���s��ʯ��Y����y��8�1��r� ����֝	G��EYx�'��++��g����3R�i4{7����^�Z�*�,Hu��@S�	�>Q3s����.��ֶD&�*P�NN��@1s�e\6)�D(1EQ�&�G{ܵJ����)Vb߿As�!NQ�8Qh�����2����߬� �K�x���k�%��-Wb�홥9�xT�t�$݂���"���X��s��eJRjN�����X������3p�oB[혁&��q�|���.cU��^�@�^6_Xx��9O)s�>{�C $���u1�_
�U�|m��j%�EA���ƾ��]yT2���	��cFU�V>��'���&�+�/��ưot��~y�G^���ϓG�D<u��]���/S0�}�u�j��������x���5:r¢���ׯ(j��K"L�݄G̢#�M��_Ʈ�2� ��8�o�jZ�Ϫ�|`
��*q�ԫl�O�
�ed��NK	s8{H:X���1Rso��B~i��>V{��5L��S)�\�]�	�:c�0A�[�kWlcoA�Қ1��0�YeO�c�x)ЁQk�2��|�K�vÏ|��E��J�=x�P#�Fą
vsi��҅���"�E�Yc
����*j�^%�]���j���647�n��Ug�x&J,�eM,�ύZ$���q�a��
qa���e��(%,ο�і���/��݆�Y�8�l�X�"�>��2ˈ"JJH�Loc�ɵن�;k���Z�����Ͻ�d%��I�X�Ǳ%���<�C����{��Cd&�I�r��ӌ�:�Mm�[�E6rD�r�~(.هs�Ǥ�:������L��늙b�#�xr��8����٩(GK�a遺"���9˱�&�9���5�O�4aX>k�gf�3�Y��$e?;�/<��P��v���4 xN���H�S��h,w;�0������� L5�>JV?^�HC�m��=���9z�1��GB�s����3ڢF��YA���@�Ԇ�pU�E� )�`A���3S$��˗5������2 3A�,Y����ɦ�^�b�;���١op����m,V@Z��-���[C�8��WvT�Y��Q�搘V�$�;b�hϼ��̰d-3Q�6�����(�]��ƴ�o}��ӾaM����o�B�v;��' 
�?��Øk}Z(
B��GO���NA7oW�E,�SW�
踓o�2ֶ/��e�d2L��a/�W��B\E�������1��@�<8ad���	��"�`iG��i�����6ŏ1�v|�(g�����U1�ed�W��R���)L��G\� ���(�p�VӇ]�dHv���t�&�IF��:=�N��;P�	,�r3��S����'`(�'�,�x-����f���@�zr#�ה�τ���#b��������#�ԁ��oM�m�P����qvZ��̋Iq��^r��=$�&�,͇�&{��sJ�Q�QS�z�����G�%����e���-������
X��M�H����6��N;�c�yLuѱ-�\��7s�;7Q�D�G�}�t�
��2p_��Cq۞�}/�}fZ�ǉk���S|Z,���ݪ*�q|�u��vf��|K��
x�.���u��a���/�8�n�Ss	�����:�!��t�n��;Rh�w����*|b�O^��h�1R}�]_�?�^Ug<�5諹�Bf����,�"���U�t8����~gQ�|l�F�
=��ǲ�A2�-�\t�+"�`�&�]y�U�r/�s�AQi��|�Ki&����
_�9%����j\�Pԯ��2 (n���~��6��mv�,R����
66s(�oM<ë�!Q��I��ݧ�cp ����W�[Ǫf��i���COPz@��"o��K�	t�3�ɱ�#$������,��7%!���`����Upj�r���D��=�n�LM��D6�����W��6�)�,[{HԆ��1׃������65���3�H�tgMn��5^	1ʁ=�)2]�7�Y����%]�:�vك�c*���r"K
��(I� QD� ��]3�"�U/BC�.��7�ุ~�����O	�����	��t�D�5�e�F�7ԛa<^s������m���DE�����i���
󞜆9��r��V�㗇Eb�Nl�T��A_���r��Ȱ[1��71��l~�����=�p;V}=D���,ŭ�ItZ��t��a[��č��5�R�3gD�@���\㌗Iu���S�pu� g��Rd۷��3d��ww�笒����f�=�q��Ч��h0��yJ��:|PI�מQ�r>�4{��W��!g�1eyQ�6���KW�Bʦ�S�ڂT��,���)Y	�D7�K`����#S�z�؉7� O�d�-C!�n��Y`﹅a.��� �Q����N�qk*-�P��������F	�bX%���غOiJ����k����H�5�E�)��YY��[�)J�b�vʭd�����ܦ|]B�w�n�6V��g%���&f뱳�~�2�#ۻd���k�n�^�S����&t�\���+��i�������@HN�G�̓6�Hj��=���Q�M�{Zg����_�"}�R{#��\�Z!O�g�Y�fcSo����["���no4�V#�|��Z��?�o`�gtq:V���� �b�IU�
���|��!��K�����J��B}7��-I,���D%&��O�#~��$%x!���{�@��賛���0��.��2#�	��v�>u���4�VG��\>`Q0���U���P=�!ϻȊ�[�k�6�����+ ���K��_�Nה��X��v;��J��>;��v� r& ��f��W�)�w�h�A���Ir���B���ȩvO�U�A?>j�������A��z5ȃ5�LF��6��Sz>fF�#1p�P���oA���9�'�� ��X��~��w�e��)��	e�`�1�vb*�=i�U��Aص�b=ye�`�*��P7�26a�?֩��A���W�[�� �`�L��Nm��*?C|�D�a��ҽ�ЊLX 8��@L����&���`���⠳�u�����D^�]��9/j�D�� ���S�Y��J�T�[�L ἡ4`a��ݸx#��E�2�������� ��'%���s_�K"Z��;�/���\����P��8EQ��P(_�ZZ]C޿�l߳F3��ϰ�ը'�ܓ8�tlC�e!w8�"с-��B�<G��KZY%�F���%��:�do�����O]�S�-�Ҕ�4[j��\�����
�axW ��?��h���	�{.[3r)�P�9�l�ˬ5�lvga�ho*�_c��B�Y�li�8)m�3�5�ʛ�������m�����?�x�^'��4�tБsu�A_HN=%��LA�FcaiB���cP�	3�ꛜY�[��Ů�.K���&vܹ��MR��!..b����:�;p�C�MĞv��}[�4�I�}��ղ�0��q-c����H�S)����>͝�DK�I@�О�o�{1`bV�,��F3*�=rDVޕ8b��Co��n���w: �k|+*�Ə���<z�4�'�I�^S��w_Gi|Q������ܰpQ��\���@j�)T	5 ��=���7��?�Q�&G��b$#��v��t�+�.�,]���vS�R�����KT 8����)+&���P�} ��<����F��8>a�]���o�)�Of��os���l����D��D	<�E3�;�i`���������h���>CJX��͇n���H#�g��1�</p,������z����y��	~c�]<�9F�B�N㣹<�K�֨���
� ��F@�����F��Q+sʅX4?w%�"�eXA�cm��WE���廋Ĥ���m���^�àM�_��H2��(��(��r_0۴�Dmix2��?<\>*�pG��]�8�"�j��_��;��}�܍�T�owu:�mG��QL��y�V~���!ðr�	&�T_^!�L�E�G��ŪTŮ>F�t!�Jf9F���3�rf���o���Q~D��������x��og=�{��jM���q��	�M�o�=��3��)F��6-q�	��� ��p�bf��C�����R��'���D�~�����:0GR�bF)��Ct*�����\D�vYدk���I�׬�@� ��J��|���Daq(�N�\-�Ѐ�qwb����M[�b��r�1c	(:d��>���%(��^G*<�p���_:�cZ�����B�ft�ݸ=)Ī~3�p�㫕M� \��aB�0�����,'=�@8?�8{bC�7�t���m�ʑ��/άz��l�{Q��$���E#Dr�?�K��i
�>��֐�ԁ�N��$>(�����T>�׫~~M*ߗJ|�16NL�p�B��k�>��N]m~A~Dct�̐\8'�T��%I�y�ʎ�K��P�@�.���WZӥ���E���Z����Xj5t>�Hς2�޲&�k$j9(�w�U�vw���Wh ��{2M6��\�D%"��3;��Ǥ�?"FN�5�!h�ѭ��μ%Y�|�s+�UM�1
Ug�������G�ΰY��� k�+p���3���4��h洙��T-��I���u@@�ᗞ�3���V[䅉�5D Rid�iNȥ�@��	eV�<�~!�1�%;��v{��>��Eң#��y�F�b�����h�ؚx|����l!�����}��B�ܴ�r�Yo&
F�%�E.�(�oI�z����ƣ.Sx�����[>o�\������� �4�?:��h�0.	M��[Ƽ���M���l)W5��v�9�hC�鍳M��*�YO*�VJ��t�5�|w�>l_z!>�}(J����L��'�c�H�sɳ�3S=y4�\��P&a=���OS��~㿪>��-/���qD��Ҙ��(v��סU�����.����׹�:5�,����5'vdk9[�4_���4��q��1��ÔH�%����Qj����Wޝ�[�r����b*�w�ܠ�*��������b	o���n%�Ywh���q*عڏ�Q*<N�:�{�2���e�w3�|�4ɰ�|0�QlD��.���)� h	<.���k��?j�9Q���8P#����y^+a�,i�ާk�æ=:��H��8�B��%��+�R�Bv}��<�7m�F�ފ84]\Q�C�9)#"�Ì>s�@<T�C!��p֙Gb�a�`�ߵ��T��HL@���C�H�졂�3��#o��K1���p��Թɾ;z����kf��r~���]���Fמ����/�"V�*���1
~ȓh��OȃF[I(+��)X1*wy&���A:����w�Q双T���[m�w����Ǡ!���Xs^2���r��F���ڔm=�[2�6�?;S>~q0G��Ȍ��>�_!" ���0��T���u���Gv�HLBd`��3�@D!��I�]��T3e���h���H���ҮaK��!�`�f�����Er�uu�CS���M�~��W�����`���{�*��V������O��M���k�[����4���-Ŧ��ƥB��2b:��Ci=�ժa����w����ޮ�b�`0�(�b�U�ist�Y3���G��ʞn�?�m�84$��p@q���6JH��j7aŁ�N��
-�����LwcE��h�_�h[�uK�� 0c�?dl����Wq(��ZG~X*p��K���c.����+���AtS��=�9~�ִp�{��M�0(�a��ʝ{��9L=�JE���O1��/��Hd����e��/"����
�{�7a$�R^Ew1y�|��	iލ�V��3�$K�Y^���OY�+"�~ٍ���m��M6���D��BC����Ͱ̢��~S[c���0�F������g:yď���P�#�eܫݘ�b���B���^��j	,�ɜ�:2q�`z�����Dj���w���v�'u�� o�2!��J�D�7��錿�୓W�"�ӄuBDс��"|_Y�&%mWҌ)�H1^�X��2��t��d8G�Y�U�Tc�+D�ê/Q�3`��4I����t˨
��C��@�����3����q�]͛DtM�8"�N�7@� \e�u��RQ)1Pɚ�x�{*� ��I��W�M}0�o��福Khf�ŚL����V��.�K��)�^�: A��;ܑ���9��Cx��9�,�D�����������2��BUegsN`p��Lٌ��ySw�����VۛIN�_t�Nlw�3���`{'nM먨8{�I0?4�R�� ����(
����u}��������6W:8��h���J�u��B:��Gus;F��OH���4���g�
���>��9�\n�#}^�OŘ�TrA�)��:�)*�|�Qu\�����`��@Ͷ�����_%�b)���n	Aa���OzXo���Z�񲶿�<�����H8���$ �|���#��͈�zUd~�U��20wq�e�xC5s몢5��P[j��uK۹;�]lޢU������Y��8s��j�W�c%A|9�+�� ��s�NH���}8k�R��rW����S��(DA-���L}��9ܜ�'��Pc�m�/CǡMȲ7��gTT��g�4^�q�PQ�u~E�tA+em��0�����q��Z������S&���x�U��v~�O�߼��[�@tx�%�)��0���I�H)�7��*A��g�Us�9���f�tu`��^������	 4G~���m�"��ɫ�lެ�e�^ƓlC�i�p�ª�-�x�VlYTv����0I���1�X#߅������ظ���
1J�`�qM��!<��ȅ��J�OvWwpV�SJ_�j༱�r`3w�˗$iWì]�l�9܍p�k_�d
�	����n��9���qpBl���3�صZ�^E'�u�'c�9O<	~9#)Ű�̝��}����y�^��$.�����J B�~�hf��T��O�e.r]$a����>�.�s�  cE x�KGB(ze��[�9����l�|L�n3��$	��H[M�z�o�ߏ�c�� �+?�x�_`m�<�!��g�̐�K\�X/�K�U��b��ԑ�yϨGf�E���.� h���t��2�{st9��h<�{���|�D�.�Z�F@d��_R�Έ�K|)�#{���m~�<�5�����u�V�4v��[�#���f�V1��f�q#,)ê'zHz�+�l���~��_0޿�D��`�q��b�����*	*:�s��b+6	o�!�n�40w����γ*:"Y���u<0��۝7��Q��wyy|����8���QN��Ue�v�;)Jx����y��m�j?�Q����Z,�#	�P��s�+C,����	�:�H8��g�3�8Ғ��r�+�Bϰd��}V�u<�-�OFB8t�]���%WP)Eђ%?�s���"U�eP��z���;���Ԕ`�7�5I]��������C�y��؋d5��X!���D1���p"�ҹ��z(E�͟����~���]��F9D�D[Ϲ�:��L���H�*
�����!��q�F�T+i��X�.w�]e�E7�A�|֓}��3����=��{dmdʮ����/���|�2�Bt��lr��2�۪�dm�,2r�?r��> �hGc�^Ȯ@���m_î���R3AT��=u0��GX��Ldb��I���R�!y�p��T��;�B����&
� �Įte6�p!��f�>��3�r\�#�%�j��Ʈ�괓��J��Ie��N��Q�`�v����q�mM�p�e���,�'�-g���o��!9:b��WCTPՌL��*;H����tvD�Dk�0�0�b|���t��Uu�2���l�j�!=�Z>�0�@׉��Jj"T���agyN��b-��6 a�w���͙�΁0P[g�hc��d��t���:(��'G���p�� U[Ac=��<��x�et���=��~�'�p�v�CoA~5a�[��ѓ��n=j��K ���9�B�`s�;����N/Ą�ܥCf{ǌ�$�KE'�[���	Wi@h���DA�c@�ĊH$tZ���)����M:�~;��ߍN��b��6��>æ�B��z��+���|~w�'cj=������['�y�o`�ޙP>��d�S�M�:�D�a滟��Q	��5#j�Pɾ��2ӽ��ѥ��7j�C.w�߼vm��WG{ *��2�멗��D����l��!(֭5��'@��d=���Į)Y��5��󌋃�1 R_b���|����G�V�Yh� �v�,+����ц�3B��4k̡����JK�����eZ@C"r�Ǿ3c0ø̙!���D���N>/�@!�~eL�H�4�$15z2��W{�&]uw-���߯L3��爿?h�@��5m��H��[K�CA���?�~E�� ���29��VxD���݂�Q��Ιt���c� e:��N¤>����N������S.�=�+�Ɯ���N���3��`]�Do^R��RtI��4� ˷e���N��u_m��0v��`�M�x|�:�1R�D����Su���:�i�G��IF&~�O*i��V��Jͽg��o�k0����\�0 }��O�T�H�z���4��)Rf�s�8\
v�Y����E���Ԁ�-�qǸ�)�Hon+�P���.z��y���0��!���[	��*[����bX�����viG�9�,U���?����5=I�7r��j�qK}�?��>�U�n׮��-�;�8���jUR���|aj�X,�O���*�I�������	no^H�1��y��R�6��q�i��V�F25���	U�S��,��-�cD���6��kNb�l������0hQ�O�R�x�����k'����ɽq[�|�E:�نe�x/n��!��
���i8&�Ҁ޳}�EMg�
���v�q����*�CE���da7�[�� ��֍,?�M
O$Q�(q�Z�e��Vܔ��8,I�|�q���o�e�؆T������ݘ%>���l�J��\Ӈ��d�3�u�k,u �Aշ.8��@d0�?IE�H�XfNO%�A��G]��`���p�C���r�Ra�n~:�r���ʔ�r#���p~�臮��bV:��A�F�nLv���z��f��S������Wr�٤�I�,�a��W"9]���/9��"&��8TJ����O�y)a/���n33e���X;1K<;)���d�<� 3����HX���CR�;���$���KL��#�DkVZ<�H�>�m�so�3$9F��.Z��j��;�ڽ��-��׼��~�p�J���R��K��S(�U�m����,���I�A��V�H�aL6�}5�G\:�JB~���m��V;���Fɸ�����C����J
H���QV�7�;��h��*�3���EQ�^��۬/(S��v���}JҔ�|x7�-�Q��A�B���+#
��\�a}�yB�۱O,{�N��W�~���=
�, oG&����Ad�EK�<X�W��r\�Ʃ�MN�vՍ1���WY�do��	_�
���)Հ�־�ր��1�WQv��t�Ђ�x[ԯ�8��Reˣ�l0н(����ַ���MYH���K]��h��/�'&,%%�=�#��v��	��r.@VSߢ&��u&�B���e��0��"qK@]��r�+�ﵚ�F��#}� �\����Ͽ��
g��nbP&�,��Z�D��Ppq�r^���=�z�&��{�	r�S*����:ka1[��17s͖�t^�n&F�sV�8+>�W��؀>��!�s.�}���,�Z`��@TM�i����\P2��t@��q�y����L���M I-ʶ+6V�ϒ'���,�~��
p��}i���r�����*��]��6'����H��g�B�'F\1�g탛��z�K��,�:]��k�(�U9�
��"�������� �2�]��<"T��/4��. �7a�k�j����zO;��� ̛���D���e c�7F>�<d��s:�Jo��~�ң��D7#��"����ﵼd��_��D���V�
㉉�b,�����SV����A��`���N �^R�� ���L�}p��0=���D�d�c��#�t�Ʊ�V���n<R�f�33��Ų���%��;툐Q>xꌂ��U�F
c�M!�9gq6x�rz�~9<��:X���W��
e�9�N2��^�
�M�	⤓�I�Nf��Hh��a���c���� 4��Q���Y섘�)�����b���/ޏ��?n�4QO+��<�#+`���9!+�,m���+]�ê_��^{��|8@V��){=+~W�F�}xSV<�?F�U;8���]`[����,)'{@�G&s,��& �G\�לo֝S�ߓ�f`��L�W�L��G*0C�G��%b��?ߠ�J�ġ1��p��&�M1�z�b��+���~^�]�KaF[�`��̅���j�.H��jtM
"�q�����S1�F��t+ˋX�+�w}q�g�>A> ��M��ZD��pEm�ɮ�����N�\S2Q�ϑ�cB��e�m��2�	�?�n_>��G��ȐɁ��r�_%(�-S�4��TZ�u���G�`>LF��k�$�D0!��a�T� ;�����OP�Ю�>�On�!J�2f�����er�e���C��)��w�[�h�)uK���/����
��0���S}�MN�o�_Ջ�2鈖%�-��J���2b�b`Cmu�.|C�_���fݦ� ���0�ub����m�t�e$7�&�TW��Ξ-����<E�/�@uM��X"�JL�����a�EeNQ%�-��BFywgk��oO#�c��[9��ʈVca��dp1�����[�(7�*G���pj���c�u������tW��=���~��p>Օ�]u�8�a�#D�!���=�~=�����Ӕ��(8�������;Z/&��G�{��x$�nE{�V�?U���ibWo���A�����$�
=�]�ֶr,t�/�o~]�7��c3�Y�6��.����BG�?�j�̦X~���c̔S��T������}��y�^ˣ"_P �;�~|ܯ#��濜�=�s���|j���ɠ:i2��f~�E�Y7'j�w��v�o���) �c2���N֡D}Ƣ�jq�C�t�����u�y�,��&\Y#��qz;��?�1b��/��y����
G��nY
ly�XJ�+ȻN�3	�3�U�4Mof��_ˬ.R��*^GS�@e����3�۸��C����Dx+?���N 5[@CP�e����֑L1�T�8�{.���a��������s���*�hj���:����m�"U�K�Ͳ���$	A翤�쿙:9�Sx��H���8���^�4�]��m�O�e�N�ٯP��(<{���7k���u�͞ �c�N���3�s:`�OQ.����I4S��0F ����_��N�uK�D�������:����x��m�N�5uDX :ֽ#G��aF�RO��K�8`�lޤg�98M ��ȟ\�o} �WOI�zTvҡ������p)��f�U�E\,J*��k�v��ͺ��O�J)r�)e.�nX ���z\W�'iX��m�C�V��'���������0P��^�]�rU���Y-�ݶ��u2�2�K5w[â���T�j��KߋT��~� �9���6�	���P�8wɒjwo�g��|�N{��Z�q{��F��B�ܼ��f	��H�4o��+Rp��ē_Ri��VX�25�v�+v�q�[����26cf��☻�k�T�l�O����0
�O�:�x��T�k����������|qg%E�{��GT�xQT���;�
SҦi��Ң:����E�ޣ
��{�Æ_I5�%�����7P�v���u�,a�}MiB=�$39*q�7�����W7���*,k����T:��K�G�#�v�m�)�+���>���%Z�JEs��)"�F�j�:��k��7�����<�bT���=���hNXH�%�rV�����qb��Y��5� Oer\U��P��:���P�c�lr��
�~e /�PS�D:��ʟ�rL�뇅���\-��Qᇅ�6�9M���HaFo�"��픲��9~�&ke�6��1�,OR��a�8z�d��3U_��a�;��<����XӞ�P �U.��nHz�!��^;|�d����:R�L�mPwR4V<��H�<�m�5��9�(x�nS�0��Z�&ڟ����-��9�l��p�AE�9�q�/����S
���Vr��-����A
��b�����_=��i`���V��F�m��4V]稷�/��Z�������I�\�� E�c��V�~P;�Xhb$6��p�NWQkI�}E�(5R��5��Zz}���^��O	��H��B�����
�3���}���B��?ON�N~E�W�	���4
z�o��33��mJd�Sn��HwI�q<-a0@++�����;�9(<��7�2�]ӓ� j��HO�:�R�;�J��������L�rÜVq�=H�&maZ6����9�>7�n:��%�� m��{��{殊T���p�<E��Df3���S?k4�d��炟��V��d�A_ö��ɘ�{�����>Y!�!�D��ȦmI��V�B�������(]����Gc4�茤E2VF_�;�jh�m��J���P�Q�ȑ��Q�(����$��O�u}��������$eս��B�����/
R�uE�}LkFB�1O#�XN���W���؅As
Z�o�q���0�1�d�e��w�W���\KA۩�	�͇�1Ƨ��n��df"�	6���Ry]�x��M���'�1�Tv�y��յ�_e��7�υ��ɶ���������4���s������J]��P(P��f{&&EZa�=�ޒ�-ִ	Ip�r��IS6���o�Y�Y���Y�����M\@�e�r����Fk��}��#���S5�^�ƫġ�6�{P^7m�cI�Z��;����q�^d��=V<&Y튇`��;����kX�-�ˈTs�Ȼt�5=&�ke@�8bscW�G�5\!�?�s����	J��bQ�p��M��;�(���S����z���q?0��h^ƻf��MWD��"�����'�{Ѩ�I	�@�]?_���f�4s�aU�ٟ'`��,h�y�DT�^�Rq$�sl4u#Y$�ʆ���Q��`m <��2ը��~ �D�VO� ��s>���iV�O���*�5GV��YS�E�@����1���4]��&��G��Y:\ ��@$+�wr�cK73��4}���<$f��#��JJwy	@�����359<�޼���D�5��\NP��@sl�e�WI�z:1G���h��{^��GKh�+j�]rޣ�3�Z,�h�� ��\|�R�K��,kT����%����9Ix�iv����ۃ[�dv���ކ5�xeL�N�ͯ�����8R����gG�����F���tN m03-n6`/Z��t���*�Id�ݛ	� ݆�܈6��x}u1��B~b�����
э:��-G���~Q�ut��:d�G) F�D�O�V�h���g��h�О�\"�.}P�
Oya�T��֡��z�ƶI)޵V��5\\�>v�B��k�&Y\�)�^'n=��F|Cz��(W1�h�sS�����"���V�\3�P�Hʼ�KpNU���w�����KbT�5�=��!�
�j?��K
�?v�P~6��n̮<з��8�'�j���ϗe�|�>��ġ7G弈6�r3��b�	�� H'��K�R��V��KZi?!�V�o�5�4*[�F��.��m.�?��c��K��]8k =l>j7w���0:E�O���x��=�wk���){��d�|�ѦE,W�w
Ex����=D
��iJ?K��N����E�W
 H�'1�H��=�UP��"��7�sf��	����,���M��fܮf$c�4q#�����(���*�@,����������w}Q��RW�YJ���>�9o�U�Ju5%�Y
��v��jx�k��4��`��@R�������/:���Xx!%�v��)'���2b�����0qr��?рC�:��+�q����r5��?�;~�r,���t��:>���\�LH�뷻���X���e���K�i����&8bravϔ"%7���E980�&�]if�
�a�=O�!�a��̦�B^3��첑 �;9<M���A��5y f��H�2J���;����6)��jv�L"��B�Vl��H�mx����9'�R�I��`h����Ϲ��&l�i3e����p #�iw���u��S:t���!r�������ߞ�A:�Ӏ蜽�3`G���;���ߡܜ͎�^Gm��V�ˠ���ɊTA�Bd�$Ʋ_��i�����V!�A;OTlh���EkӰ1�QJ������(eЭ�e.��Dd}�¾��*���x��B�g��=:n
-��
�}���B�1�O~�uN�םW��.� �
5�o�A6c�Ļ,��d������W��d\����pe�c�1a��i�d�wo	��V�m��Ւ�>�(,�#�1�I�v���4V%��E�:�J�)��쒣?��Џ����2�)���.�������]ѽ�cLV���&!<�_7�=E�ЪH��	�l�r�+Sq���}��T�V�E��b�@��7@o�!rp҂ׁ}ՄTK#��+̮Cw�jh��Z��Z�bP�T0��Z�*;�X��qu`C^�u=��&4z7��/�%H>�۩�k���V�s�M�tp^%&����s�8�~W
����	@!��Is  ��}�ŬE���ϸMW먎#�΀��Х����q���C쥻��kM�|?x9}�.�Jy'��x�MS��4�?���=�V�aj�4��IUwӍ'{�s,�E�y�(���kE�n)�4`΋�i��� ��?Z��Ux�h��#F~P�Ӣ��Rc/q�Bm����Wsp����h���X��g���G��Q�r`���-�:��cn��a*���~�m��.VPzKB!� `�Bw��#B6���uMz���$�K�Y1�Ǣ2�X�B7㥧"�ZTӱu����]����÷���۔GK�Pz 
::i��W*�/T�יA�1�.������^PW܎di��!��nV;g꺯�C�&D�Ω�۰@a(}O'���P��)�{!pCȟ�~'���=|T��yR �^xg�P��	uJ�;���}A�`���/�R�,���c\
�;���XUcxZ]֪���u�؞�[VN@]? %��0���l���I�a��m�vQ6�3���O���G�S�u,��^�4&��0��U������L1"l�Ы+O�����^9�Ca��p��
��޸f�wY Kx�D&�0�KJ���Y�$~��h�����<�P���gJ[-�=�N.����!ۅJ�jJ���W��6V�@�_Zy�����Lw�>�$N5��x�dl�Hэ<�_��d�7B��XO�:M�9���=қl�A�l�$T��*����x '��79� a~�}�����&��j0�ť[�����R���h� ����48��٘��ez��$-/|�;�.��� L�E�H_�����Uz���[���Gx�H�����xY��ˮ�H'�az)��[��3+��ԫ���
��@�E�\g�Ry�X�w.����b��O���py���ff�mE���.��%��f�P���g��s��n�4��{b�|� .�"�l@�R�_}P�%G6)��{�$ �R�ͅ�O��{�U����Eq��tŭ?kl���y 5�)��#�U��[c��'"=f&͵�/���5��&�G�C)�����<�+�]E�/
��4S�Ӂ��+�g	�y/ʢ'<�4����ܮ�w3 ������:~	vqN:���^�ZAT���/8�|�i{䔨������^�,:��ܣ�x�Jh�u�5Ou������ai������J��~J{�+�8����o���a���g���ٗ������JP��\I\N13�/��E���Y<�C�TM�H�(�/�q�O�2��䤼ԣIT�69��5����_&
7q�C�|�Co�½��K�znL�-F�\7�I;�J/|X�"z���Kj��ж�^����\�ft%�i�ft�X
�}h�����I����iӓ4I%࿔��%�@\��Ÿ�������LD�X���ă�ycb2%ꤡ-�������R�Q�����4٩�����
Ԁ��X���)�}�7=fON��u���/n�t*�=��*��c��f�~RKc��x(-����3���~a�[��b�8E�HhVĮE���!�������g�$AR(�-*��{�����
�RR�_�K0^j��g�y� n�7���,)�˴,nt��	��wOg�il�����4�\�>A7g���t[���*F̪���|�J�/��A��Q� �!�2{��z��֞A���m������?(�S��*-�I��C�mI�,�?��c�6� 1()��MQ�����L�[�ҟ�c�@��N��,���Qd�~Idϒ��P��?��?i�%���>����=��z��Wx;��W@#"��r�.�9�C�O֘�U���2�h��Z�â��q"F�i�ҫ���QZ|�~gcO$f6$o>=|��A"�����0�4�lc�f�F||����o�LhtLEj�6y u�IP�
<�Z|���!���)���=�	��7'��I'N��p��Y�j�#��)$ �m�pT�������<�0n��9#
���Q�_u�T4������	>��E0<�+U�%���c!�r9�)�=k=�����Ϻ��z���X��V���^��K2���A;Y���4�)�הß�2��)�ih���}J7r�(��Ps����vʫUU��>�Ov�/�H�<>���b����Zg6-��)�����>�#��RP��wo�_�ey�9�"�{ٍ�eA�MJ4�oh3e��v�M�R��Ͻ�ν*%�=�0�l�|�����0e�/o*�M7���6/�?Q~$�[�����|W�"������!Lk�0m�mM?��&D�p���%~QiW�`�LL���A|���*u��Z����q�K��7�^���oT�jӶa�{�n��N���9�,&q�\׶)T ͆��O���\��x�`E)'��~��%P_� k��%�*����&ݼZ@�.;.�*����֟�v�Sx���2(:&�Z�d���T�l�6��m������E�Wu�O}���M�8&��(��BC	��]Y6.�F]�%l[�,�o�1���ڗƪ��S_��ү��[�&�\s`���:��� �gV?A;�h�ɖ	[x[�4��|'��t=lp��5��dv��h*x��z�;�'P}Y�)��s���15�~�E2:a�F衐${���³N�'/���o�sА<Ѥ=@QGa�\�Y�a��$���0���E�`�������N$���v3������.�q��%X:���þ��yl�v�rc[=)ʈDwէ;4����qH|��o|�Hkg^0{�Ԙ����Cޤɽ�Yu���}�b�V��c@*��7��٪lbc�ox�n�. w�2��F�*?&�'Kp<u�?ۂy��Е�,0Xwڬ�|,���qrwh6Q��������)o���p�� �rD�?�/�Q�Ж?��#��5��ld+*�,����=���;�����y8�o����\+�U ��f#}[fV<1���F���8�W�]#�Y��^V)���*Lps_.�gq��J�Y���_�`��߶�t`ue�:�/��O��g	C�9�숔	��D��J �B 1�.p�⃹�a�z����R6����~���]ZzF>Û���7���1�����
�z����ϔ��F��+ںX/B�w�\ڠ��AɆ�B`���������9R�m��خ����F�2t��`�W��}+�O��mdA2��[?��>E�G(�c�$����_h/�Bԫ7q�Th��uU��Gj�L�
řN�,؇�3!��~�d4cT8��g������Ņ�yO���h!턧f���|�fr�|���2u�   �  C  �  �  �*  g6  B  �M  oY  .d  �o  �z  W�  ��  ��  F�  ��  >�  ��  Ҽ  �  ]�  ��  �  t�  ��  1�  ��  ��  o�  � ?	 � � � �# a* �4 �= �C `L &U �[ b Yh �l  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+a��6 \��	�<4�d5h��'�B�'���'	�'/�'�B�'��I2w��5Kk����e��U�D܃��'�b�'A��'���'}��'��'�>��5�\ h4tIR �>���'l��'��'���'2�'���'b�Iz�k�fVЂG�[�x.(���'���'/2�'��'"�'"�'�^�qs�S%V��c߁Lb>ıf�'��'@r�'���' ��'h��'J����b���@�3MTV<q�'�B�'�'���'���'^��'��`�$�͡9Ql�#[�=�"���?i��?����?!��?9���?A���?P�Σ9<�x�
�&�+K[�Jъ���O<���O��D�O����O���O��DLw�eȴ���ŢW�2(�'��O0��O���O"���O�d�O&���O,���ƏX���K�8�n͊���OP�$�O��D�O����O����Oz���OL,���0�"&�:3�f�j���O����OD���O����O����Or���Oؕ����JT�
�G�Oݨ��Ԣ�OT��OF�$�O���O����O����OH�0t�ʰ[O�XbQd|�^4�G��OP�d�O@�D�O����O���Lئ��iީ�ć/TF�U�ՁN�:�Z�34�ڂ����O��S�g~�h���%k�2�8�!#$>=�B��PX
`��	��M���y�'a�S�)� @���@-\��r���'�R��5Ǜ����'r|�Ę~��!O1*�E� � �͛z��?�.O>�}�1�A%��D�(�����6뛦����'5���nz�)����Kp�D��ě�D&�!�����	�<Y�O1�N��ƌs���	�3��2�,yp����	�>���	�<��'�@�G{�O�2eʝ9f-�F�@1�=�3"�.�y�Q��$� Y�4+�(�<ɠ�L���(�&K�	H�JU�,��'�(��?)��ybQ����J۔Zx^�`��F�t���01
"?���j�l8�aB�ḑj�n�d���?)V�Ѣ�lG�M:9��0���#��D�<9�S��yR
�M�Q0EJ�h�*A��-�yR�|�8�[��`�4����4.��";���1��3B�ڰ�@:�y��'�b�'n!�T�i����|*��O�l�b�}-bCVBŕJ�(pن%�f�Uy�OF2�'b��'��lS?^��U��F��X�f�ھY��	*�M��J����O��?aQ!!�(AV��"�#E�>9�wI���d\Ц1�ܴ!������OQ��#�S��` `�&{�J����Ӹat-�A��GDҫ�N8��������@≾��?;hdTY�PM~n�¿葊D�'R��'����P�\ڴd��Az����P&�Z��ya���"#d����1d���CY}��iӌIl�M��4	x�AҫA�K�^��TL��F"��۴�y"�Q�R����@ek:ظ��'��t��0
B篂�E�X�S�ꑈ!����k���y��'���'�b�'����f;��5I�:}�HL:TI%^q�$�O����ꦉSrn>��	�M�K>��]69yzѦkڞ.Qy"3���+3�'P��Bb�2��[�j�7-������12�n�y��@r��1}�*��C�rʚ@y�%p�0��|����?	�x"n������{����Ęj2>:���?-O)lڍ|D��I�D��u�4�$9d�͹H��j���bU������T}R�t�Ȧ��N<�O��å�ކV}�#W�
�T���S�)�/\M��3vF�2���º���O��!.O�N O��A���c�a	�*��w�f���O����Ob��i�<���i��AC̈6䈍� �:PH:t�a�[�4�R�'p@6�)�I���Ē���� �'��	Q�Ƞrl��wKÿ�M�ճigܘ���i����O<��D�
��c��8���3^ra���Xz ��g-�Mc.O����O$���O�$�Onʧ9�����f׃!�*��D�j��P��i�f�sT�d�	^�ϟ�R���+r`�&��y!wf�"u�iQP�ƶ�?!�sd���O�\�0b�iY������� �t�2�C�$���M/	,�	�>ʓ�E�ey�O���8�t�bA�.�p�ĉ��Q��'s�'���!�M�bM�?!��?	�
� |lMJ��L��b���(��'����?I����'V5{Ei�-a0��q�²)7����'�����١B=��$Iƺ+���O�A2���.��r)�ezDd����y������?����?)����F�n�������1� �x��\R|�'"vj���ͦ�8�� �	��M��w2I����- E*�懌x��@�'���p���l�
�lZ�<�7<��;p�0|!D��G���z4�>;X��Ǚ��D�Ԧѕ����'��'��'���F��yt�)m�L 	]�0�޴c��m����?����O�Bp��-,"!�s�]!gj>���	�>��iw�7g�i>����?�ط��,Ws�� `�,5y���喽Z%~�r��/?	�'�-p�@�d��ަ��'��t��U������9Q�E���'���'}�����X��0��Z�8��\^|}���2R�FȂ7Bњ@g�L����Mc�2��<���M���i>~0��͕!l2%��
>�h��q�ܪyk�<O��D�>T�H��.C�I��u���� �l!$K�Y�Q�t�Sh��2O��d�O\�d�O����O��?��`l�$���#֊ 
@#G.�ٟ@����؉�4f(���'�?��ir�'��M��L�����Sd	
er�y�|b�j�R�n��������!̓��a��٭ho&����+���A!$бg뾌�F2A�֑xƻ<����?����?���Кl�B��!GKG��)A�G��?����$
Цq+�L矀����0�O�02Ŗ0l����N���O"��'���'Tɧ��y��ჯG�8��-pGCI�w*z����:�>����[p��y�ɃHQ�0���\(�`��!Ɛ ����ş\���`�)�Suyb%u��V�[rR�u��FږM|pt�BN��E���d�OFim�O�o[��֟�т'�='�r� ��	�����mџ��ɰ+�f�l�<a�xN��07��Hi�'��a���*��2BYf�D'*�I����I����	̟���b��MÏ�Ƙ:��ݗ���,/�D6�C���d�O���;�)�Od�lz�5#ǟ�Hl�3��J�Xp���A3�?�����?I�S�?-�EE��)ΓQ��g��8�����
/�H�͓}fލ�p��O0��H>�(O,���O�q��`h���E~��3��O�,#�i�O
�d�<�ǰ��Z�$�O���O���A���r���cJ�S8tq���(�ɱ�����}��ē*?"���
�Do p³b�Lah͓�?1��&;`Q�� ���D������ب��A�H���+u�G.h�Ѥ䈦�4�d�OR���O���'�'�?qe�Ə8����O���/߈�?qQ�i
 ��#�':2�f�P�杣]����V.<Vpz]E�ž<|Z�	��M���'��6o�>��6��Lŀ�8>s��,� ���֏֑ H\Q�'��k��$�D�'(��'vr�'6��'�2ԋ�g��	2�(Ade��Bk�pP!^����4SH�z���?�����Odn�j�/۩l�|��R�ò"�[���>����?	I>ͧ�?y�%z�kQEC#g�~��1l�\f�eЖĎ�M{`X��2�(4$t��9���<���M,JA8�!�6W�u�c&��?i���?Y���?ͧ��D榅SE�@͟,��JS`��oW#�
�!w�S�8�4��'HL듼?���?	T�R����`J9�!�Q��$b��A`ܴ�y��'
	��PIR.O�i���|8�ㆊ(c��b�ǿ~���@A7Ol�$�O����Oh�$�O�?���"!-���AB�'����˟�	`�۴'����Oy�7:���~S�e� ׶k�Z!��B�NF�O���O���"7Mm�P�	=T���)��E�*=ބ�����:'-B�r�X�]y�Ol��'AZ���Zs����X�C�̑a��y�����'�7�J�n� ���O4���>�)��o�ƉscÅ�`<��E.�ɔ���O���<�4���d)J� �I�(m�����)G	(�"6t���F��X��(1��W�	S��Ţ�gH�W�Fx�FP=qw�Q������I����)��pyR�s��%b�ɬjں9��F�<eZI0��k�����O��o�k����ɛ�M�2��)q�c�.ޛ- �����9��f`nӆ�Q�n���I͟\��(\�v��� eyr���$���(*��m�ZaJ�Γ��D�O^��O����O��$�|�'��D�HU�0��*4)����-G��_
B�'���T�'x�7=�QS`C�y���6�K�o�ʨ;�!L���������|��������M�'�\�����8-A
�"Ĝ~�Ș'Ɍ����pq�|�U���I�X���ה{"�H��oE�%�R�ğ,�	ş���yy"�y�0�j���O��d�Od�C�R�I�A��� �UC�n'��+���ƦM����3�0��3"k ����W�a,�'@� 8���{�d0����X0p�'��0���Z ��s�����'f��'���'��>���!U��Q2�c�R��8����Q��(�	3�?ѣdΟ|�ɾ�Mk��w�p�$OЇeF8�e�J'mn�,[�'2"�'t򼔸��4�y��'0�4ӦǊ�?�Ħ�8��%SU�'Mh�=+�/m�'k�i>���ޟL���P���c\œ��J|�&�y���1K��̖'D�7M,^����O��#�9O�M)\@Yk �\��Zq
��I�'�x6mY즡�H<ͧ���'&��ɠ�˝�r@��b��&(��+֎�M�ȁ�'HP�����蟸E�|�]�p�TJR7l�Y��K�rnx��K��0�	ϟh�	���Iy2,b�X�[1�O�8�3�� �@8zŃI3 '�-zB��O��m�ʟ4%���O�<oZ��?a�4|4MStO� %0f�ځM�0�@a*(�M��'�b���b,�S�l��?����3����4��}1(Z�K��I����	ݟt�Iݟ��I{��,�,�Z����Y�C�������?y��	�V������'y>7M"��=X�ڰ���
"������Qzx�'��n��M��'�Rq��4�yr�'8�A�p�A�&E����M07��Q�!OڶK����<n(�'��Iʟ\�I����	>)"�a�d 5g��4s�JE)o*��	ן�'T�6��^����O����|��j2>��#��"9�q��k~�+�<����?�L>���?�+@ج�L�Fk�h{Qm����@8n��'����̟��R�|U-�@�T�@=0��(@�îw���'2�'o���Q���ܴ&s0鲴�S�^��m &�L=\.�xk֢߮����ئ��?Y&V��`�4~\2���u��ip���1*[��Bҵi��7mA	M�6�h�p�	�y���G�O���S�?  1؅#�l�\)�`��n
<S:Ot��?��?���?i�����ȳ B�q�EИhJ��jE�QE><�oڤ��'�2��4�'�86=��۰�J0t\�|���9N
*ac���Y�4=]����Oj��H�8��F;O6�[�����5�?�@��2OJH��+� �?��(�d�<ͧ�?�B)�2s)rt���N/|MHh��>�?����?!���dPĦ���������ӟ`B�ۆIdp����A�|^@A����B��V�������IL�;P����8f�d�gML7N��h�c�	�Pr�ԣ$?���.����F��?��j��FL�)�u Ι�ĩ�@@��?���?���?Y����O�@Ҵ�ԙ2[:D)6LN�z�
�G�O�}mZ�NH����ϟ���4���y���BK�1���U�G6��H��y��'��1O@a�¹i�iݩ`��Kj�޸B*��`�K�D��{a�������O|�d�O^��O��$V";c��cJ��U"إ4�Z>/�˓U����q���'�2����'���˵�ұ_k�5rE]�e��xҀL�>Y���?	L>ͧ�?��8� q��,!1|͑2OT�q�EBE���M��P��#�.�*��d(���<!T��4j� ɳ�҇n�b�
���?a���?	���?ͧ���즭��k��0��)Ţl�:�����A�V�1�����޴��'����?���?q�l\Y�X�y�M֧`��r1/�/Yz�Q�4�y��'1���LYx:,Od�����0�Rd�%� ���s���8#4OD���Oh���OP�D�Ol�?M� �Р|&���lϭ[DV����ԟ�Iܟ�{�4WG2tΧ�?9��i��'@J�xmΝ.J�\�IS4`�B��$��){ܴ�u���M��'�R�D�w�B���O�~Gh�x!����^)ZJT�\�g�|2Z��S�4�	�DP�����h�(�I5�ҟ��	[y�#r����`��O��d�O�ʧIv�i�	�#�șX�IN�dq�Y�'c��$p�6�nӊ|&��
*�٤ꄹW�"��� F�)�����2�ր��i�H~�O~���I$v�'i��PŃ0FtpPs�fȏ|�n3��'c2�'J"���O|�	��M�S$�UK0��W ��ut�U���F-"���A��?�T�i��O���'��K�{$����$�����W/r�'Dh�!�i}��OD�r��J���W�W�WL�k�nȠ\e���n�\�'���'s�'�B�'-哥:نUp���0^R�`D��Ed<kڴB������?��䧟?����y���H�dh�!
��Vd���A���'�ɧ���'���	N#�F:O5�F�F������)d�:w:Oh�`��x��I���'u�i>q�I���E�Ɏ
(TB�"ƿe�����<����$�'�6��  �D�O���F�a�Q3	O�&�u�Ga�� �~�XٯO���OԓOb���M�I��/������=�y2�'~�}�������O��)���?���OD�Iф��0��F�	�x�H@p���O����O�d�Oң}2�]� ��ܟ}�*�s�,�1Zt���d���u���'��6-9�i޵R�*F�Z���)d4AK3�m�Ъڴ,*��j�,dpaz�j�IğH��OS25d���	m֘�hC�]���,�'R4?(�$� �����'�R�'���'bb(��7y��q��G	��8�R��K�4R�P��?Q���䧗?)�:9�t�S�U9�@�`�W< �	��M[��i(O�����ɕ,l�A�$�ܐ.��������b������Hp�Im^65)w�'���'�8�'+> P�J�0Ju����O�9Be~i��'�R�'�R���X� �ڴZ�H0@�:�q�6h�.U>U��X�V�z,���V�����`y��'���GcӤ���k� O�4�pm_�	�TQ�4��6�f����#*�,���O�h�����3�b�+hH�8V@ES�B� /�b���?����?���?y���O�D�h�I�
-�������nT��B��'�b�'|6;��I�O�mE�	�rJ4M�E,M�l(�LA�݊y$��:O<���i����O��y��i��	�r�4IQ�-�;�bUb�B����v�͓7����{��Ry��'c��'Z�P5"�JxH��G�]6dţ��3|V"�'m���M��
H�?A���?�+���R��E�8�-�b��/w��"����R�Ox�nZ��?�O<�O�F��bE�BXΌ; '�((����mZ`&�����B:�i>��0�'�
�%�D꓌��)�ܩ�v�%*�\}"QO�㟰�Iݟ<�I��b>9�'Ȋ6ML
"~nL"%�'H���
�%tO|��g�O.�D�%�?9�Z�x�4�5��c� ܁�
(UX^I3żi��7ʇ]cf7Md�0��5v |#��O�@��'��ܳ����R��ң/5X耟'I�	ϟ$���t�	���I���A�J�Όa��k13,K�l�n6M^.����O��=���O|amz����<1��)��D�g/���J�ɟL��^�i>e��ٟ�Ce���͓�άX-I	�pX�r�ʈ5:�Γt�2����O��PK>1(O�i�O�%XXM&(m���~�>�.#���'���'��I��MS���?����?Ɇ%̯O�6(�W.��x�W���'Ҁ��?�����'��l� ��$ �����WH�H͓�?Y��S�U�8��4h�	�?�J��O���ٖ@#��֭_� �@��Y���$�O���O��D<��[�k��=&��e�A\S:���%_<�?Y�iKZ ���'�b%w�D��c��=:��ۀN;��7�Y�^q���ßH�	��p(��¦%͓��Ԡ�^s�� ��2���NY�b�G3/��a9��"��<����?����?���?Ѳ��`k2���U� � ��텶����զ�ZЁݟ��I���*� 9	��]�U��*̀H	��,l��	�����`�i>��	柌c�/Rt��BFL�g�.�ɒ�Z�r�J�o���N�[�B�k�'��'��	ۮ8B �%Ml4Q3נ�&��I���	ݟ��i>і'-�6�\m������5��\�Q�m��p�,R��lJ�',6m-�ə���ߦ	�4՛V�#x����Y%8_ؘ�gӬJ�P)�i>�I�M(*1*1�O�q�,��D3~!h�;-4�!@�՝w����O"�d�O*�$�O�$0��1��v	U7��ysb2Sꌕ'~"�j�X��A7����ۦ�$��#�ر"^��Ɣ�:�`�C��O8��w��He�J�i\v�|7�d� �	;J�ac��� �i��'Ԍp(�7�O�Wor+�V�Ipy�O��'�bA	��,Uӡ-G�,$�cN�0< B�'���/�MC���?y��?/�Ќ;�/�5)2���Ε�C��3�����OB�o"�?�N<�'�ZFGI"�b@��7t��G�N�lt�%b�퐯}���3)O��)�7�?9F�-��5;a�uyaa[�X{��PDĻV����O��D�Oh��	�<I�i#@� ���6|��l ��'hE*52NA�R���'��6m(�	,��d�¦e㠄�K��ð�$ N�E���MC��i�ʜ���iC�$�O�,�_�
,�<94��5!��Ђ/-I���"��`���d�O���O����ON�d�|j����78J����J)^�-r��/:��vd,U���'eR����'�6=�8ʱ�6����ҡn���a��s����|j���
�/	�M��'sH=3���C��q`a�
=*-�y��'\��3�J�ğ�B�|�Z����՟�۲�46)b "�y����I���I��`�	Zy�j���q��O����OL��\���y�o�52Ҹ�2�4�	�����O��<�dKN
he�QŖl⨅c@�ٿb���O�%�K�N17��Dy��OW�|��?y�h� ��8*� ��4UGi	�?���?	��?���)�O��Ұ��+:���i�����ְ�?Iq�i�tF�'��v�^��]:V$��-D:�E�l��I⟸�I�$җ��馥Γ��4C �l���I�y��M���T�:�d<{��7 �Onʓ�?Y��?y���?��%-ؔ�� �m������<��X@(O�nڙ�~��I`�	v��TQ����p���b5G���U���	˟�'��S��h���*j�a��³s�ܨ�WLX) �B8���ɦU:,OLyb��~�|T�l�a��?����rS�VZX����˟d���$�	���Cy�r�X�+�/�O�Y0�/.������ �Bzf5 �M�O��n�P��I��IٟL�����S�� d�B��D?��P�5X'��Im��<���g�������'����wS�\����S,�$[�凭:s�h�'��'b�' ��'�p-8R=i�l=�	c�K.)����O.�����0�Ap>�����M�L>ID%L��%�-ܹw���� ���䓧?����?�˴�M+�'���J
����T� �� Ĺ_���u�
͟� �|R^��͟��	����m��fa�]�aِ#F(���ߟ�I`y��hӈ �$/�O
���OHʧ3�~XBAظ94��	�"R*�M�'��?9���S�FQ<jD����+�(��Ř6b�B��27����O��A(�?y:����=���X�/]�D���ȕ+T����O����O���I�<��ip���!�Hz�D(�2�@�Ȇ��80��'��7�;�	����O���BH�>u��su���q*�I�v��O,�$	6X�65?��O��'�V�)=�b��QJԇ&1S������y�Z�H������I埤�	ڟ`�O�XI��D�v� wK*�	�0�r��q�C��Ob��O"��`�$�����$ih5sd�L�sﰁ��J�_LL�Iӟ�'���������Xl�<y���WD�1�@C
?3���3���<iE䋞	>�$_,����4�4�dR�:���7DE)�� ޜdu��d�O���OJ�1ޛc�{;r�'��m��c�PX8`ύ�uJ���)0���|b�>Q��iV�6M}�I�2I�{��/6������&]z�I�l�Ҋ\
6z�hr�7?���o����/�?A�>m�f��8,�����+�?y���?i��?��I�OĜ�E�C�X����[�Z�ZU�W'�O��m<�}�	�|0۴���ywM�*tJ�����1O��E8e����y�h{Ӑpl��MK�ׇ�MS�OR�St�Ӎ��N\H"��Z1��� �j|	4��T)ƓOl��|����?y���?���hK�6s,&D&$�d�"My�g�2XX�@�Ob���O�	�|���mhR�*��?�2u����e3�V������8K>�S�?����>���
ZTi���9�E�go�H�L�Csa[4/�OޙZH>A,O��i�"M�xj���#ȸArSF�O����O*�D�O�i�<aƼi֞- �'uLAG+�7!$t�v��&ZT�YG�'��7$�ɯ�����C�4>�f�N"M6$�G�F�d�.JcbV�YT��	�ia�d�O�̒5�ݚ�;^����?U���W�(�����wz�� ����X��۟T�I͟������	V�'>Y���bJG�:���ħ�5Q�d���?���eD�6������'Bv68�����u5b�y�NU�
H�� �[��M#���.ôh�֖� p#n.� �5P$��H>��wkG�&���XR,���?���*�D�<�'�?Y���?��	�SS�X �J�3i���Ñ���?���?���M��E$E��?�-���lz>=�e�;n�a�s�S�U6����K2?)�W�(�ܴW�f�;�4�D�I�8j�2V2Ch�œ�L=*��`�Cɸy��%c�����p�bH�y�	�ntܠ��	�����'�8dFQ��ߟ���Ο��)��\y��x�@��(ӓ=d@Ę��:/,�?(l5����?ɴ�i;�Oȩ�'p�6���;�@����Ts>��7��>U�z$n��M��b��M�'lB���ɖ��ӿa��Iy�`
�ڗK�Mp�R�Z,��	gy"�'���'�r�'�RX>�A6I�8�����5M=���
�Må���?���?�K~��9���w&�H���B}P�cs�E(Km�D(`m��\�IR�i>!��?y7%U̦�ngDLKg'x��xѢ*��ǮΓv֠pjGI�O�AK>I/O����O襹b�A&(���R�ֶ6gd�+�g�O8���OH���<)�i����'���'r�%��e݊v�l1�Z4���c��V}�}Ӭ���u�?��#g��/!l�Ǆ%��������V�}&�,����my�OU���	�v����ҝ�2	�Z�z@n��h*��'�R�'�R�s�%��B�#��y���B֒��2MП��47��%8���?���i�O�N��$���eK�O,�sT�ӥ3���O6�D�O8ܹf�{��	NWi����� �)4�-
�J��<+�dܨ?A�'��	П��Iԟd�	ԟ��	�|ǐ9�eT���Q��N�A����'  6M�)9v�D�O��$.�i�O���bA	N�J#`�;v�˒d|}R�'��|�O��'C�YS��^)6�g�#v�j��R@��RC���<�U˖���{�By�F�	)VK�bp���e/�N�B�'���'��OE�	��M�r�A��?�@��=a�,a�ܩ#�*Aqv��<i �i*�O���'�R�i�6W�����<��0`%�C����m���韬�AR(�$�-?q��ݿK��Ո��̨C��v���n�<����?���?���?	��TCŝEOF�" h#ބ3�f��E6��'�2�j��P���<�'�iD�'0@be�P�L���0�+H��s�A#�dL�!��|J�e���M��O����GH�,3Q�@�w�Z�x�6��I��?aE)�$�<ͧ�?q��?᠊��ID�ժW�E?t��q %
��?�����ڦ��nF�������(�O������N(KVX���ӕ�1?��R��)�4v�v�.�4�P���,'6�T��v�M�vI�.��̪fc��*�T��A����S�R"�q�I(�
ZQ A?��=��O��������	����)�|ymӾT���?e��Y1c�u��u��kݒnK�ʓb����A}�Di�|D��E�>0`��G<��F�Ħ��ߴ(���ڴ�y��'�����?���O��K'MX�4�hS�`F?¨��8O���?����?���?1�����Y9S����bG0c��T�@�ӧ,uoڳ&�X���ԟ\���?��OQ2�s��	�O�6��3�Jz�0G�ٲM3P�d�O��O���O��D�3gdT7-v�ti��֖\�32	�s����j�`9!�N�#��$>���<���?��(�JZ4p�Zpm��U��<�?����?�����ܦ�a�L����Iʟ@����0�L	Q�̄�%�yJs��E��qh��ȟ�I~��\C(]��o��B��U�ϧx�R�����-Ė��oڊ��埠 H�'jbV��l�0ß�t��9i�׶�R�' r�'2������A͞F�Di�a�M*X|<(&��۟���4a&�i��?��i"�O�N�m>��f�DJO�d c�U/z/�D���Y��47�v*l��;O�$�t&n���'j>XI{�ˍ;PDr�NL`�܍�e�<�Ĭ<!���?���?���?�po�u�f5C,�3gFb�JA�B:��$V��9`C�W˟�	���'?�	WҔ�Z0-m@^�`���\���y�OmoZ��?�M<�'�:�'"�xtag�]qQ�Ұ5즐-^����@�Ty��62*����W�'.�I�:��x�ǎ�	������u�~��͟��	����i>��'�@7���j�d�$�������o��Q0��}���d�y�?��Z�ܳشw2·iq8y�nٱ$fP1�)	j�p@�eE�����$Á�L��,IS����	 �A<fT}���"^���x1�w��������؟��I�L��G�\!x�JV�{�j �?����?�s�i���	�O�/u���O�asP�R�i�$�A�
�6�A�8�D�O��d�O���jo�&��~S�I�.y�mӠk�c����`�!ڈ��'B�'@�i�MC��?��H�z	��@��;�8D�dk?mImB��?i*O�m�{(�x�'��]>�"`D!?�8߱ri 	��6?�Z����П�$��)��2�����\E"Ř��MN`t�7E��?�h�5e_}���B%��O&��H>�1+�37B����Z]�Vt�R�؅�?a��?A��?�|�,O�,n�#Ğ�HD�Z�)�v�F�	� �R���˟`����M��2H�>���(\��!HƄJ��Q��l�+���?�����MӜ'���K��SQy�!�j 4�&˘4O��;���*�y2R�8�����Iڟ�	����O��Y���r^ڹ��͋�
K�U���}Ӏ�QP��O���Od���|���w%�4�5�>KFȰ���
��XU�h�f�l����|����®�MK��� �uA�&F��%sbAFD��:O�i�����?A�@$�d�<�'�?���KpH�ps+W!z���&fC-�?I���?Y����ܦ�K���I՟����f�*����B82�E+"�~�VD�	�M�R�i��O.�p`�5:>� 1`Fi�X�#�;O2���Nf��$(?G>�	�?���'�|X��'k����`ޭ���pK8BP�I�����ɟ��I`�O���W�J�,-�gO#�<�c/�
���uӆ0�`��<��i�"�|�w;��` 8�0�Q.C�+z,��'�6-զ���4�&M��4�y��'�6(�2��?�`�*����S���F�r����B�|�X���x�I���I���$��S����af�>ĎD봮W[y�a�@�zdd�O��D�O��?��w�N�_���Pn��v�@�)������Ol��,�4�����O ��A��'-1�J��w�ى��T�jPm�P��8� �-(�`��ly�(R2^�:s�b��TLs�*� ���'2�'��O�剂�M�E�Y�?ѷ&�5�P��ꄾ6	Bqrb�	�?a��ir�Ob`�'�"�'�r���bȠ���
y��ȫ���`�qJ!�iV�D�O����S����ߡ��N��@j����?2��I�u������ ��̟x��������(]uf�a�	�-	�:,+����?����?a2�iX���O�GsӖ�$�<!qg��9!P�ެ���������?����?����M��'������=�4��+�Ѕ�zv&mꡏ��x$���'2�'���'���[dH�g�ݨ1!��^��$�'�rU�`�4s��(���?����i7��x��X�zf�S֠�9)��.����O���,�4��dX�V�N$6�Cjh��%F�|�V�ݭ2��7_yB�O�l�����w�j�����n���4ȹ�()����?)��?��S�'��Ė�q�%�"b6 �td��~����7u�B$�'�T6m.�ɦ��������‮MH���Z,UD)1�m���M���i��u�'�i �ɭL��u�t�O_�' x�|J�Ӡ1���Q�nW�,
�1ϓ��d�O����O����O��Ģ|ꕏ^7]��j�9'xщ��-r��f��� ��֟�&?��	�Mϻ~uVQ�`���p����O��q����v�i8���0��iLq1.7M� R�!��eSa"�bk�����y� B@��)B��X�	py2�'��.Ԯ]9Z���KH�4}PB���e���'��'^剑�M��]��?���?G�Y�CZ�d���? Bf�pEh���'�
˓�?���ēe�,l�I�q_��T-�3Ǫ8��?�%�=�ذ�pL������VH��*��X�l��lƶ䚼��] ����O(�d�O���1ڧ�?�r�I}~��� �ȌD5�A<�?)e�i�L��':��j�F����h2�j׀
�"UqgF� >��>�M{r�iL�7�T�F��6�x���Iv�l��O��,5&�5|p��fO������a�P��sy2�'��'�"�'Q�̓�~B�� ��N<8a�y",T�&��	��M�G���?y��?�M~r�)(��a�W�C�`iQN׌L���؂R��	�t&�� �	�X/�x���j3��ڀ�K*P�m��B�7C��U�Zj&��O�[J>y.O��HA��Ͳ�Ő�j����qf�O����O*���O��<af�'���Q�S��1�$�� i)GkL].u9��w3�F�D�L}R�'T2�'yX�`�
q��+��{w�T��GM�p�6Or���B[� �����	�?��])�4}cӪ�`�I�ǿ|�n�����Il������	U�''��q�U�=�XX��W�h.pR��?���( ���������'p7M*���!4N8���W*`M,�J�U�{3��O,���O����&9�7�y���'��)�z��DD[,Xnx�&���~�|�\�D�����������*��y������/(���1��_ɟ��IoyR�k��8Q�<�����ͨ<���ɗ�U�\5��D�9g��ɰ��D�O���,�4�r�d�T�9�DgX�|�~D�EcͰ/�RP��-	�rU�w�����J ��O�&~pH�B�)^	r��e#�(��1��������l�)�Sy2�xӎi�@�Q/z�d;5���7��{�h��H���O��n�^������� 9��ÐVlP)*�g�l�����ܟ��I���al�<�OP"�ן`�B��jP�[$)~�����l]���d�OD���On���O���|ruc�28����-?��E+�B�{��^|'�	���&?��	&�Mϻ^3J,�pk�"��)Pr��:
H|�����?9J>�'�?9��B<��C�4�y".�":��F����Fj}�	�N԰����OړO���?���ohP�0O�JiCi¬��
���I�����^y��jӢT���<���h�$Ӂ�z{bI����)S �5�����m�ޟ��Ik��HtDj_�ųիR�W�v���'�6B�J�{�,�FyB�O���	�R�k.!:l�	�d7p/��%A�B�'�'W2����ks� �2��E�hm*�2�n�ޟ���4�v�����?i �i!�O���o{�C�m�A��ɈC/ֽ0�� �	�ݴx0��Ϟ8D��?O��$�|�P�s�'h{.a���%)����W�f�h�{��;�D�<����?���?����?)Ak�)y^������0^>�{�g�#��DԦ�����꟤�I���&?�����\t�'��wM��,&��h@�h
D}"�}��(�	F�)��@zl� n��g�P�d"e#��{T�kGI>V��˓b�D��N�OF�SL>�-O`eceK��w���VBѫc���8���OD���O|���O�)�<9w�O�ԩ��ߎ��G�	.M$>1H���)�����D�����e}��'3�'K��"�B[�y��0���Q�s���C�m������n(���4����&��k۶O��J�,�$K*4��&=O����Od���O`���O��?��Q�I)+��lʱcT(�i}y��'�z6�O�
����Oz�o�g�I
~<����h�{v��AE ���$���Iğ擕9�Em�q~ZwR�țO
-C�mI��'TQ�-G`>Y��D"���<���?A���?a�*�Ft��Y/���3N�r��	��'�H7�Bx�$�O��|25Hίa�����U)T�$�PD�L~� �>Q��?N>�Op2a�sd��%L<A:�ğ=��3'�>S��"�i����|�2���x&���E`�i�����2a���;��
ޟ�	��`���b>E�'= 7-�"(e�DX��H|Hd$�`�B��P�Af�O����a�?ɑ\�t�޴��i�eՓ$>)1F�-�<<�i<�6��'*�7-;?�!�(=�	3���T�7ʊ�9�Ĉ�e��lP�aV��y�\��������	���I�X�Oy,X���@ pT�E'O({z}!�eӶm���O���O����� ��]�Re�vm��s�,�z��Ģu�VTPٴlқf�<��צDn6-u�l�B̄D��5!D(y/li�F!x�l@D�ݕC�R��v�	Uy�O�2(17є�[$kUy���ׁ@�P���'�r�'U�%�M[R��?����?	R"D�=!�P� �e���C���!��'p�] �-|ӄ&�ܲ�$��~�ĩC�u�L�c�~�0�I�H:� Dm�9�����qh�O,ѱ��^UB�D�)I��U��0��P���?����?1���h�|�75T�)@'-,Jf�9W*8�D�ӦAr��\�I��M���wd���t��mO �p�jU�%C�r�'b�'��䎄x�V1O���ժBK�4��'T���	;y�Ҩ�0G�IJ���Щ:�D�<ͧ�?A���?���?��c�ŀ�Q��\��Q������d�̦A�����\��Ɵ$'?Y�Ʉs��0�D��+�w��7*�1�O(���OP�O��O���',rPjת����W�%�q�m�"'�I� $ /�?qpB7���<QA��6*��WN�1[$�
��q���شHk�s�J5\u�#��(,5������α���C���ĎP}�'�b�'���Aq���b�Ppc��@�&mY�m��v����Tc��pq�	:�	��6%1E��;G���Kx��A�:O���D��-Ɉ�x2���h �(��Ć�.�����O�����+M3
4�i�'�뀘�"C�a����b �!j�	ß��i>)q�����u�?}#�a`'m��^T���Pa��_�����O^�O����'�蔐�߻J>���PӪU����A����j����	ӟL�O?�ä�
����.T�a�l�s�O���'���'iɧ�)���P��Aɒ��)YQE�<o��n�3�86�Aey�O������}JD��)͍������{J^���Q6�v�� ��y4�kd�X�'�P�x� ��'�oӈ㟴��O��d�0�����}��P@  7Stv�d�O���a��Ӻ��O����T�|�1E�o��D���U��ڽ��`�X�'��{��Š&i20L@�JW͸å�z,6m�����O���)�S�M�;�~��!\�l�� ��8��A����?�I>�|�����M��'� �	��ȍDW|�B��\���`�'<�dI��Ag?!L>�*O
�K���RF�*6i�36�,�ra�ቀ�M�$*�<�?	���?�qƙ�0��X�%#��
�Q�Un7��'��듐?����!�\LPAb�z�>p����%Q���'�P��V�D9E/��K!�釉�~2�'߈�hE#*2�� �3��ͣ�'@�x����g	��c0��A��+��'�7-��;���OzDmZD�Ӽcg�X�ed���g�9[P�֤ �<)���?��b�t۴���������?�Ѐ��&KDĬ��-s�]KQK_�IRy���!3�~|
`��LԮd��$�/	 r�'�b�iÈ{#�l01	A,sH�K���j̈�'�B�'ɧ�O8����]�V!�Iک~<�)B��(u�����<9�AC'�@�	s��RyүC�ya�ܰ��&��@)�#���0>��i�Ͱ��'�L b�ڤ&��MXb�A�{����'2�7m2������O���OhI2B�ːv��Mp%D�:PB��$Cٜ7m ?�K��]���k�S��E����b����Uf��G$��jd�e����� ��<p'�]�p���h�HZ:P���ß��	��MC��VJ�D|�ԒOzP����7,!��[
&��"�'��O,�4�\�s"i���Ӻ۴cڗ��A�a�.`�@��`��:��y��'��'��	|�l^�L�<�(	��D�>'��Ex��cӴ���O���Oʧ`��	��P+^X��+Z�=���'�$꓍?	����S��  8�цWŤ����_�P`��n�gn��ɤ	x������$e�f?!O>��O<GD�8��:鸸��nDz<q��i$���X�Z	Z!��.�)h�xCmĒjE��'�@6�-�I�����OҸ� 	����%E�B�O��jq#�O��3p7�9?��5��!�O�"O��`J.2P10�	q�<I��?	���?A���?Q.�re:����<����JzR�zQ\��r��,��ȟ�&?)�	�M�;6�t���m9�Z��S�y�r�bF�i��D=�󩃦B��6d��:��ֳ!�6�ƌX��ؤm�,RbÍCoR��X��Ly"�'��cҖ'����b�0��s`M�$B�'��')�I��M����?i��?���T�[Į�b�cLb�U���Z���'���{ƛ���O�O,)+@�J&m0��n�����\��&��P��Ih�C�w�R�rC�埄��aJ=S|@(+FiȤn˸Ղ���`����Vr����1�'�?�m�"?�~�A���Z���tK�$�?qa�i<���'��o{�N��]23��A�0F��\���dT�#n��	̟��ݟTh�I�צ-�u��-#l����D�!���l�t0۶�^d��O~ʓ�?I���?���?q�'%��چG�-g��z��H�{y���.O|m�*9�������H��W�S����'F��ԃ:6�	�ɋ
7j�%دO��D�OR�O1����Q�^��Ba��"���TQ����6mFzy��
u.������G�QS�P�����K���q@��p�a|�
i�(-b�+�O�M�!�]���|8�L�xd����O0�oZX��r���ܟ�����XD��>����e�EK*��P�Pm�}n�U~��ʑCY����䧩��'�G��@H�I��9&�Q�<q�@#$0�����7pȘ{��W<7Fr8"���?1�xg�����IBܦ�'��z��(e��x��j�40�Ĺ[�h��8�i>
'C���u����Z�V�@�Iߖ�+" Nq����Op�Oʓ��'Br*e�+;�ċ�D�{X�PC��$�Цɒ����8�	Οx�O�%!��TqjK�rჇFH~�Ŵ>���?	J>�O�0qU�M��H��^�f����
Wq|+аi���|��+��x$��S��aڊ�J�(�C�d�3j/���ڴVf���q��,*�ٍM�L��G0�?�������Il}��'����N�%Fr��~��B��'����旟�ݥ%I�'���,^6�� g�V}\x;.�2n��Ī<���?����?	��?�.� �C���+�	��ܨ@���[!Y���yeG�ៜ��ԟp&?�����Mϻ
bL�I�*(�B4��
h���?�J>�|�t�
�MÜ'���qH�s�L�t��2���r�'��a8� �ş� Ú|�P��S��bH�?��-z��[����l�؟�����`��_y��h��D��M�O����O�� �N!��\`d�@�nV�42e�;�	����O��$ �Ĝ"?Fz]ؤ!�)&\t��&ۙ&��ɊSdL
�	�3G�b>MA�'M���ɩ\.���Q�
\.XL�7*Ӗ��	�����\���O��`F@��d�V�M�v�P�VOD�sӜ����O���F��}�?�;#��3���1I��$���	9r	����?���?醬��M��O��@���O�1X��������u�@�0���#gf�O���|���?a��?�����9����h�q1oS�4�*O�o��z�'����$�'^�`�t%ȒTNB�xU'��+� %H5b�>q���?YM>�|*2�
�?Z�hP�M�B0k�Jɍs��7��o~�����\�I+_�'��ɇ�n�JР��ch"y��L׻�4i�I����֟��i>��'�6�<}�:���M�B!��J����Q�Yr�U T�'�6 �I+����O��$�O�����I��d{��G�T��q�&�)�N6�!?!��WmBb�)3���U�3������uǉ6m4jD���i�$��ݟ �IƟ<�I���󯍋%}f4��n��a��P�J���?i��?	��ib섻�OL�j}Ӑ�O6�3Sj�/-斄�B�ךt������3���O<�4�丣�L}�L�L�l�
�*�oH�Ҕ�c�v�J�J��X��U��䓊�4� ���O��DՊa���eѻU�2a��jE�=5����O��9e���0�r�'�R>��.Ź��xi��b%���J#?�V���	蟌'��a�.D�@�Ҏ2�,���ʝ.�N���H�&�B�9��o~�O[ȑ��%^@�'�<3Fn�S^<�DdER(�˰�'���'^��O�I5�M����!�r��E9T�a���	�Z����?�&�i��OHM�'r���H86�*r�(�Xb,�%���'���90�i����M��0W�O�n���Ά�&H	ʃ����E+^�D8h����J�(�A�C�8a�̃�;v�ɅɄ��bA��!{L�Ie�&?�t���`�u���$Fـ^�V9��T��(���WVν��K��"�q�Ë�G�!�Ŵiv��L�h��A�͜8�9�p��ܼ�av�M^���!#��SP� N�|����DΛ6&�����
^�\0GQ�Gt����Y2d$&��y08��4�D0Z���\���g`�g@9uEB&v�QQ\��C���m
"0��kC'1#z��@d�A�4]t��6�4	�4�?	��?A�'Gb�O��( %��f.� �֌J���ݦZcD%�S�OAB�1� �!Z�n�O� �c&�c%���i���'|rj�
V+�O����O�I���@�5E
>1����į��{��b�P��o0�	⟜�	�x�#/�:.xڭZ�ƍJB���C)�>�MK��e5n�1u�x��'Kb�|Zc��w��;��}�t�)
�䚯O��9f��O����O�ʓe��8�ް:��L�h�p7D�˓��'���'*�'��	�Nخ�y��!;/�%�sj�(���`��7���,�Iҟ�'C�0z�m>m�1��,?�r��a R�+ 9@@$�>���?)I>�/O���T��"�:o�`�b"��9Fļi��>I��?�����%L4&>�򃟁?���M�?����,��M3������$%Y��OΩ!uJ��
�
$C���6D�Uz_��L�I˟��'Q,|PÄ4�	�O����)I� �+i�����J�2wBd0	a�i	��tybN������s�ƭ�.�0RN�A*�i�2<AHT��i����ڴ!o���h�S����M.C|��hE(h�Qd�H6'N�vX���h*�S�'B��9�d�1�Tպv_�%"mZk_�� ޴�?����?���zǉ'ψ	o=�9���e~"�����)S�n6��c��"|���tɕ�52��Yɠ�@�:��Uɑ�i�R�'Rh_.*�Tb��It?!��?6D�VOϺږ�QL�D�V�jt�<���?���86���ńBXp=���!a>����i�R�4��OF���O.�Ok����S Қ�>ѩ������I����	ey��c�<��)һv4��3�A�'R�9ƥ3��O���/�$#}�#gU�0.�|��3mK�����}��'���'��I%FB�X��O�P3 ��J��Oӵr ��h�4����O�O����Ot����Ŵoq*H�C�GjLE`sh�>	���?����$ݦv���O����xI+��e_hE�v�Q�E�7M�O�O��d�O�t"0k+�ɛh~��)`�ahN�� �+�06��O:�$�<Qc	R4KF�S۟(���?y)b ҰR�鹖'Kc`�g�ˊ�ē�?!��	{�M��ҟ�u"أJ��(H�h]+c� `pP�i��I8Z �4�?1��?��'d��i���6��+Bav�U<��m�����OZ5�$��O��Oh�>!;AM^�'Xx�d�<W04�q�~���Q���˦	�	͟�	�?�a�Obʓr��QHg��ag\e�ˇ�g$�DI��i9,Y��'��'�����U�*Ab��#�h�"�聪U�o��p�I͟\ A�ʀ��$�<���~�g˅^�8(�S�UO��F V���'�0���y��'���'ze��J�s��m�抒6�}�4�zӒ�d2��\�'v�П%��X�O��=a@��Xo.���_���x+�Y;�����O����O��$t:�㌓�/q��@�:sM��[�B\(T��ILy��'��'���'	�E��/3�ƨ��� 3!;�-�cM�~��X�,����	by2��?>B�Sj ��3��K=>`���d]���io�	��%���I�PRk��X�0i�;o;x�h�Mߢ�,=X�#6���O���O��PCL��Q?u��;o���aB>ao��sk7���P�4�?�N>	���?YA]���'	�%2���*3���@��)\@8��4�?�����Ĝ6{���O;b�'�������),WQ\��Ϥ_����ƝxB�'��|%��?��OϲT���,(��IC@+<;�p��4���%��m���)�OZ�)^~�!�/��+!��*2L�%f��M�)O����O>�'>�'?7��)�ĕ�1�rZr��#�k!Q�iRP�"	hӖ��OB�D��%��S${w�e��J�yܠWA�%&}��i��qSe�'��T�d'?�	ݟ����� $��.֔��@���M���?	��>枌�x��?��'�zճ ɜ@�{�A�V��ݴ�?�)O4�rZfb��<)��?�z���d��>db!��,ݏ��`hD�i�ң��d��O��'�ɧu7�ʷA��Y����;�aǟP)��_�(!�����?i)OP��֚'/���Ʊ7�ZYsC�:$p�����<����?ɏ�'��<-P��h�c�~4������`�j1��'�2Y� �ɠx=>��'^����&X"��9J�H��8���o�ٟ@�	f���?����4�`HڦA�IH6�#�) f����8��OV��?q�ʸ����O�A �[N~�0�AT�R�]�F�e�?Y��?�Ʀ]�.���'��ÁƓfKDu(�FֱD��
�r�H���<���"��(�����O8���8=�3H_/o�����D�#Bp�@�x��'G��>s���y�����CN��@��F��*@���_�X��,,��������ǟl��XyZwe�Q`�`M,_1씳��/¬!�ݴ�?�����ҬGJ�S�m�ks Ϭ &����I��@��n�="`��4�?Y��?q�'����4ЃO�
ႁcU�R����K/@��ș�V��'U�	g�3?q6�
>V%K�Me�a�@$ϧ|{�&�'��'>0���_���ɦ�"�*U�ގw��}`�)�
-48���y���-�������O��U�JP�(�//l��RW��6/(Z�o���*p����S�	N�I*���� �*xD���G<V��tk�O�:&�O��Or���<��a�� `Y0��^5���a�E�dzn��S�܅����O���'�����	�T��6��>O����吠g�n=���#�c�<�	wy��'�&u��ܟ^���b�nv�QQ*�76_Q����?I����'��'�<j�b4�M��j¼R�bt��(�/6���I}�'[r�'&�IR���M|�0�_s,i�f�:]]�U��
�f�'��'?�(�`�Id�iW8ی�OT?E �0��d���'6�W�$�E�
&�ħ�?I�����;$P,;�$��a�^Y���}�	Jy�ą$k2���џ�Z��N�Z�E��ܚdܤ&�i��	{�Ԡ��4J������ ��dF�3�h+���n9����
��R�t-�̟L8H|�N~n>�� +�?�h���N�%d_�7mЈOD8���O��D�OV���<�O���S��E�l������	)���5g�$ț�HɈB#1O>)��a�q6B�'8o2���C�Vv�!`�4�?����?Ibn�1x���gy��'��DW�p	��!�4[)&@u"�^���|Rj��yʟ���O,��(4�ݡ$�8��` -�z+�9m���\�Q��=����<������Ok��IZ���R�׼顒!C�I$;�"�?Y��?I����DF�D��TmҨW��i��� 6�����Ni}^�P�Ify�'�R�'��D�ɾ�����N�  
|��K�#�yr]�d�I៨��uyȉ�WR�ӽib�<�d�F+�Ⱒ��ÆpeJ6M�<a����d�O.���O���D9O��q��S/0��Iu`�>i��8��jѦ}�	��	؟h�'�Z�3��~��O��L{1��V�P0E�f����iNS�4�	��<�I
R������jd����3E��PG�ڌcP]m��$�Iuy�C ?Z���?������T�	/�ЦĀ�b��iH6��G������	�\9j�d��qy�؟����I)�����2i���9��i��ɮ
���ݴ�?����?���C��iݑ�$�.W�DB ��=�bU3v�p�����Oj�C䐟ȗ'!q�԰xQ���IA�dܽe�v<�%�i�܌�aJq�D�d�Ob��$�'��Ʌ����A�5��uIf�ޑV�J���43�*�͓����OR��7/#�2�EV6º�`0�Z-o�X6M�O��d�O�x�-�K}�U����N?1agR��:��B��ȰⶤU�A�	Gy�Ь�yʟ����Oj�DR�eV��lN�S.<�Jv(K�X04`n�Ꟍ�%��$�<�����Ok,�c{��BfF�0��<8�'���I�D��	ɟ����� ��ݟ��'g`��Eb�N���hgD��h�"����Y� �����O�˓�?Y���?��œw��H��d-�К���m��?A��?Q���?�)O0�j����|�"�J�%nlyR��U�����ئy�'u2\�|�����I�a�N�	��!{ş"����� w�p@�4�?����?�����D�C�,|�O��5d'd�)�`$#iP,�@A�x6��O4ʓ�?����?qU���<QH�l˱�֗��`��!���e�e�6���O�n��v[?�	ȟ0��Z�p�Q�g=tlp�	m�����O��D�OJ��L���	Vy�ןz, �m�o�X�I@��aoej�iA�	�/�$l`۴�?I��?���qo�i�	���Ǣ��Js���\4��B�wӔ�D�O�#9OP��O���,����e�� �;o����ǔP�D7-� &��l�ޟ��	��������ħ<�LM?���5%G!HK���3$��J^��yb�|����O�ܲǭ-g�E�N�F�x�笙�������������(�O�˓�?1�'��CK�H��5��%�5>���ڴ�?Y��?�VO��<�Ow��',�B´%}*�����>BV�*c,!Bf�6��O�)x�GJ}�V���Ijy���5f�ʕ06rĨ2�ːl*`҈��A+0�$�OD���Ov��|Γ{*�5�E���"�i����yA�#$��	y�'[�I����	П\�B�_�Z���Cb4�Ĵk�m�}7V�	QyB�'���'E�Ic�D���O�R��b.�$NR���h�*�jڴ��$�O���?���?Yq�L�<��N�"J�aˆd��e��#
�v%��'���'��^�$��@C�����O 0��\4�T��ձ��#�Ħ�Iny�'5r�'�^�A�'c����Ѕ���&�L���ix��o�şD��Iy�P�l�'�?���*RC�l�X:dk�>@�0�hj� 8����	�Q�$��4���2|� !��N �dǇ��M[(OnX[�`E����������?M�O�NK�8�IÇE��Y�/" �v�'hR����Ĳ<I��4�A�Um��!��+A�xh�띯�M# ��d'�F�'��'����>�(OJ�:�jJ�C����P�n�0Q#��������w�'�@�:�
՚�@��l���ۑGݫu��m���i��':�B�$m�����D�O<�	��l8����
AB<c��7�O��#����S���'T��'�lDA�eYU\R���Hٍ6����zӴ���8Yv�$�'��I����'�Zc��)h�KC�L!��a���%��M��4�?�J��<�*Of�$�OP�D�<Qe�0NbMjVc�@�h���l�����T�$�'��X� �	ן��	�xB�%���F�)S��Ό/
��ce ~�$�'�2�'��T����L�����N�����<I<`E���M�)O$�D�<���?���Q����'���K�a�)�y�
�G�t�Hܴ�?����?�����MR��O=Z� �qp�|���֧���a�io�S���I˟��	�-]�IO��.��q(FaQ��������= 7�O���<)�bA�zىO?R�O������Ђ��ҭ�tl��!=�$�O �$� 5�<��?�Z���au�"c�Q-<� g�{�V˓3�-8ֱi��맸?����O���v�����l�R�9XXȶ�i���'�P�R�'��'Rq�T�3�)Y�m�"��$D�����w�i�@�`}�<���O��d��'����8NO4����H.��9�Q���?�`��4|j0 ������Ob�G�o�s�����I`�`\Z�6��O��d�O�|��@TT��?��'?����
^�J��a���<��
ݴ��v0�������O����OkZU��Pwɀ����g�î����'�V(���3�d�O���<A����@(D�H��i�#8�J)d�i}�)��aZ����D�Ihy��i���7�T:12���B&A!�Q�F%0����%������ث���	a����jDHhr��'F=,�	@yr�'���'剈x;��y�O!~	7�ز@A��@!�0���B�O��$�O��O���O�!�51O���Qb�
6Bb�zi@9��1��-P}B�'-b�'��I � �sH|����T�贈�,�(g�����k)���'@�'���'y�p2�'7�04dI��Aèt�AY#�J8��8l��h��`yR��Z������DI��-��Oֶp�J�<;�\r��A���L��9y���W�	KB��	$���`�g�VR��X٦=�'��m
w�@p`��~�����#��|
%� ,"y(̐`)Ț*L:,ӑ��f��O������OޒO.�>�c5�l�~�N	�7(0�~Ӛ1)��ϦU�	ş �I�?u��}B�?r�$X�烚�an0� �@!�7��A��d-��4��ɟ ���\�r� k҂�Y��XT�ʈ�M����?��{�Q��x2�'���O�]��'C>[���PK@5"nX����i��'ު�
B�%���O���O���ec&z��!V#N�w�����G���"Ih$R�}��'�ɧ5օI�v϶�#!A���#� �����ȥx}�d�<A���?����^�zĐV�M�Z!�Y��Gǜ+,�Z���L��Ο\E{b�O��Z�o� @��� ;r�;#�i%2Y���ҟ���dy�훽u�b��57��Pa�X2�m�@B��,Y>��?Y��D�<	�?Rx��gB7d��Ѻ���~2�U��Z�$���P�I֟��	�j��	��p�	<�⁢��  �vHJ��"+��3ݴ�?�K>���򤍥Sb�'�0!�,��G3���KŶ��M��4�?������AR�'>}�	�?E!'��3&�ܙ:�jZ�@IC��M{�«-����i �l�e��,<g�r� x��+�4�?���J� �"���?�,O:���O�������$�\�85X܊�9ŵi�2R� ��2�S�1:[ЩP�)@?CK� 4(�Xg�iL�YwF`��d�O��$��>�'@�	t1$!h�͘b��u��e�>�]p�42!�Γ�䓅�O-ҡ��D~�(�m
�,2< {�耉w6��O��d�O8%��n]B}�]���	~?Y�a��1�V�;�&	�_}�-�G��æ���0��>J��)����?��eND��9q����b:�2�p��i�"K��JP���d�O�ʓ�?�1��x[�m7�J
��39 ���'�v���'��'Q2�'nbQ� �ddZ�;P���P�
4-+,� �ȏ�;���O�˓�?�,O��d�O��D\#PĐ�ꀳ�����уT�h$�q��0��ퟄ�	ٟ�'/��c�Mi>}q��R���)-�-��	͛��7-�<a�����O����O��9rU�D����X���C�� }� ��G|Ӝ�d�O��$�O�ʓL�X�a�[?��i��i�j�y�^鰔��Mq\H�0�{Ә���<���?i�h�(ϓ��icB��֔�~p�c��~TD��ٴ�?�����ď��O��'��$ �Jt�g��B":@	�B�#3^��?���?�PN��<!/���?)��	�\L�t�K�k)`�y�(c��ʓ�X�6�i�B�'���O,`�Ӻ�V���<���0��Of�H���d�Ȧ�Iٟ�*�~���������_�']�}K`g](y&����ƨ8�n�J\�TP�4�?����?y��vI�IMy���=7� h�	�!���0��'z��6�� '���Oʓ��O��
� ��\��GN�w ֠�o�7��O����O:l)��u}�W���	y?у�Ӆ.�z@��Y<w��'��Y�	ϟ,͓�0�)����?��O$isS �W��e���Ӛ:$,�бio⋏,L��꓍���O>��?��?{v�˧@I�;��Рk[�j��m�̟4K7 q�L�Iޟ���៨��t�4E˥Q�h�%oX�`$�@J]� (� �[���I�$�Ik�	� �%:^�аi�zS���,�.LM��m�a����?)���?/O�qs��D�|2fĄGkZ탧��<�&�E@}��'n��',�O&�[�]?i@�%�(�r��儀h*��k�&�>���?���?����&�����?y�'Y�@j���NmAE��#os��ݴ�?�J>A���ԕC�'k��A�		2��*�֭���e�>"]�O��}� ��k �@�M��Іȓ�H�@��ԗFjN\a2�ݸp�l��a.��G�\U1dFE�!s�œJD/�z��4LWIJ�ysdY1c�<��,�F�? 0@�� ��d�h�JS@�#��eɀ�	~:X��	�q�<Q�Q�����!&��P��Ћ�E��pŉ�V���$��4X�*A�}�f�!�(� %<$X�І}�����P)w�X�[���?Y���?���u�[�q��E:��M��i�f�9rf�f	�����oV�o�.l� �;擒��I1H8ؐR��ȃ,N4C�ٵZ�����D�5�Z����ȯ*�����4��w�|i��'� 0@UH�L����/�R��(2��'���$�4�4��=q0qF�(��Ȏ_ђ=��N\@�<�6�@I��,B� <	��� .My~rI>�S��P��b6��!�}�K֭8�0h�"�#1X\��"��ӟX�	̟|�I�u��'�5�d�ж��;*iFy�&΍#���`䌤*"F �c���g>X��ɜw ���w�@q�5#J ��ғJ�Y�c���=Ab�Z7'6� v͏�+@ɇ��'s����ޟ�F{���2bưtc��9c��4h[69�!�d�
=A��
A�>[j���\g�1O�%�'*�I�k  K�O0�D#7� ��5Jk�9�qgK�_�V��O0%I��O��di>�i�*��K,�ˠC��~���b��+�Xm^@��-�p<	���4g 	H"�#D��DҋJ`&q�w�9�&�S��".��x��߉�?	�����/a��Y�nݱ%�$@eF�i1O���$�37�i�B�I�)�$���F-g�!��\�B1	�)m�D]��oqU0eG"x���'xd�ʷE�>����)֟l�`�$�9���*D@͗0����3b�6:�2���O�<pp(S���2���T>��O�f�J�a��f��w�	*2�CL�(�t�c,�PVLZ7먟��@펅���1�*3<}y�>�Ac Ɵ��IL�O�?h�Ԭ�Eӯj�8�p�!�y¢�t���җ�vx IJP)�0<����<RUv�Z� �8ts|�0��ٸ.�(�#�O����Ol0ApfʇQ;n�D�O����O��ʉ7 ^�P�H���n,��JO8gpy�F	#���6J�&8�p�*�3�$[�c�i6��7��Y�DD�(l�9'��P
�-�	B8������|2A�Ey��K������٨!ҝ������O�=ړ.�����+uwf\X$��h�I�ȓӞ��D�x��Do�x�t�'�#=�O�I�G*�a�E��8����7Ac��@�W�dL&��f�'���'d­g�i�	��8ͧ�L���M�E ����,o�ta���12��f��XXdXkE�!O@t9�E>e��\a�i�� N������*0d]b�ʅP�Lx��3�p<�E���n��	?�P�c�/ITH6����M�w�i��O���~��J�$�� �-[J@���j�_�<y��J�RB�hI��NÈ�{�g]�1��Xy�P�\&z7��O���S+); ���G�y��iy�gۿIWJ��O:�! I�O����O"��-^�V�x�`V'~;b��M�pS�Uy�#O6
z:�z�F_J1�xB�^�,��haC͍�IE��`P�		� qiV�O,,8�W���XÓ~b���۟h�ܴ�?Y7N�?ɢ�AA���j��Ig.ъ��D�O��"|2�N�al��
�C�~��$d�hO?�޴c���Iab�� �8��֊G8Mx��hOV�=9�#]*=���0T��FD�E�&#�E�<�V)�7j?��h�E?����*�B�<9���*6F됢 
��\r'|�<�F��&$-��i�B�d��A4c�]�<i�'�*;Ϛ9х�A�p���o�E�<�b�.:֜{����Q�x�$��}�<��O��������W��В��R�<	�1Hl:(*C-�2�l�p�P�<��NI33���j@� ���E)�J�<�Gkߕ[�ԍ��)_�},����C�<��G�It��Q�`�07�~��Q��B�<�	���
�!��N��,��a�E�<����L���AY�a+x�õj�C�<��*&g,	�i�6�-Be�@�<A��g��q*T�8�!l�G�<9��-=�dD��k<0�xQ��f�x�<9 ��9�"{��^���:�B�q�<���;��u#���~I��j�*�E�<9&�Un�}
aD��� �P��k�<q�ܓ1W � a�߇a7�}��Gf�<�5k��	�;�`\-j�܊DUe�<�'I�8'@�-Q��ʭI�����|�<� �g �d��Kt��5EkB4�2"OF���� 4�l�"O��t���06"O�I�gƼ>��{�nD"~��`��"O�`�Ǖ�}#J����{Ŗ] "O =@e���L�S@��P����"O*)�A��ꁻ��[2^L.�0�"Ox�y��V�����`L)aG�y"O8���"��N��X;�.3#nyR"O0;��j����6
P\Kr"O�8ѩ�w�p\l���Z"O�=�cJ�'!�� X%��"�<��E"O4!��Ή�fF���
��4���"O�tЗ$J�a��բ�]�)���Hq"O0�)C%��?[>�#ǩ\6q碀�D"OL)C�)��]����K!�*�
�"O�P��,G}�n���U� �8�"O�c�E�g�]�G�W�?���"O^�a��Ҍ�<�Z�`K31E`H�"O��LH����p�N�v/��"O����/�=~��4O+�2��U"O��b��L����Ĩ� �`p�"OXYyW��o*��.���A��"O~�x�@�q�uY�-�4l�\�ap"ONQ�0���9��T9B�� �R���"O�<�B��)S��ۥ��c>!iG"O�H����EA2�9��A�P�&0u"O"q���%]�� Rg
�)�4�j"O���S�Y�����#t�H<�R"O��ZՁ8�h��L���u"O�\K�Ƌ�t������S�"��m�"O|@�,='����.^��7"Oz��Ҏ\�PBn�#rl��j�8?�y���M<�x�c(S�\��ixg`���yrg�=̮lz!%��BZvl�G��y"*Y=n�����h�$�#����yI\�F��:4f0Yi���%�+�y��e�fC%kI�JH�4 ң�y�h͋2}�lz�';9:Uq���y2��z�صjBZ�-���vL$�y�D�23J��u��z�+P2@:*������39��/�B#��e�<)��2�Đ�ǥx�	�'Cb�<�¡
3zO��*b��v�v�pt]�<ɓ-&1�����M�cJ\��e�Y�<YЏ�0\&�I׆ϵ�r=�'R�<�J:���'�'M-�գdI�W�<٥��� �v�kdr��˄��J�<�1AB/��D���")	&�	r�<���n��-B5+��en8�T*	g�<��<S6F���Ǔp�Ę�3�e�<�F���t���!ɹ}����fă#j<)
�}b���U�+�z��p��46�p�y�9D�����u�8�b"�� ���)&��OzpW�R/��>�Ag]�e���0�%e�@� 3��h��pv
�6��	�GK�����%B���b0$W�W�B�
#��8(�n�i<⁩��1�⟼�f���4��
6z��"$K�<`��y��"O�<R��"'����j��Y�A�O ���)�'�$����ö�SK$>u����'��BO�;j��u�Q�ӠRَ��OƉ�$�5lOf̹�"�: g"٫Pi� lؐI�g�'��yڱ�iKFE�Kk��[��_��5�'h��@o��V��H���@:��FK@�y*�Od�7���'P��47�H���?E���qg#P<s���d"O� �2�%.-u����.EWF�05�@(7Wr��?����.g)�6���*�S��ʱ~H���"Ñ�]��09�M@=�0=�aH٬`b�������<郎&��� \�e+N��r�ί>(�@�F�<}��%6R���'|�1J��˿0�.���ؽl^.��<�e�ٿhV>��@ga��<�;h��{7!�;*)%�G���*iΓӲ���H�d���d�
^�l�d!��A3�Y9'��)S`6����W:D�	W��b>��B-3fPM[�gw=h`5�� `��"1��B�I:yy�C#�*���2�Z�l�d���90������� FN��� ��>�O�xD�8Z�bEz@%�>jT � "LO2��a�
=:�8�1O�TJs��)l(\�* T�L�l�Q-V�T�ȹ� Ν��?����P���'�Ҷ�T�o�,���ވWYxP�y"�ߊSQh!so�"�(��,4E��#KJCȺ��`�*�@UȂ�_r$Es��=�F���L�z��WƏ�x�8}x�@�)�����tm��2
[6�ӛ0�|���˷w�p�4�T�:�TZf�[+�F�;�+�P'\��@"ORQx!́�XT�U����:G���/��h�ŅZ�\�p�l��*5�P{'����M��g:��1���ʊ�?�|�g�_8a���DݝP��sF/����d� K���Ţ�5_��asC�$H6�6Ȁ>8�JX��4,�(���9�3�$́���C����r��5ពc�1Ob���។g��<0�ӡD+�����;8�!���*%<5�V>a�,�Їo�~���ד�|�*�(]#-����G��_24���I����p�˗*o�iK1숿QE���]C��C���$ֺ|�	�'~�l{B���cI��(���&hjH�N<Un��PՓ"����0�����!M� �h�h�YZr%��j�d�!�Ćb �P�iαM��	��@���&

>%]f��'>���>)��D�PF4�I'��]�����Oh<IUN�#�АB � 	T(y�Μ�d�$7�Q-z��a�.�:�p=iG��M��Q�bö%�ЄťW8��@��Zl����)�ꟴ����F �m�BC�	����QV�fP��s'�>]4\B��*q�t��dKP���;�]��'��U
f�	S{�%�͞�8;����'���37�Г}��a`A����J�	�'Z��3��	W�"�����0��P
�'V�k W"�<T���%&�<a	�'���2W�ʔg]��Q1�H4�	�'ƖQ��G� ���ql3���yrj�O�	{P�C'�}:���yR英QX̸Z$M xw �C��'�yʉ�^���E��>>;J��ϙ;�y2-�?KEj$�@?J�h��p)��yb+�X��Mc�%M�v֞1�P
��y"�Q):��)�ƚo�I"�6�y�R�~� L�8m�.�E�ɏ�y2ㆀ>t�h+b��d؊��W�P��y�ă�8����oĕ&&�|pW��P��|��� h)$d"a�=aA��D+X���'b�lR"�L	��B�χ)l�z<(����q�O24١������I�.���)�"OtE��c\���M���	���6剞j�deË�I֗h1@�h��4P_JȂc��0�!�d�����ɦN�D  �J&%�6��� ��ا���	מ1���ɟ#Cb�*Ud?�yb������R�L%V`�������d�^ma}�O0g�XP���
�$$�{a�ڕ�y�k+~�I�f�h�|݁0��y�,�����.�<�vlή�y"�8"~T�bD� tB�H[v�P��Ċ���|
�5p�<�� ȴv�T�rp�u�<�',چW���)����P�,��Oo�	X���ɚ?<��f�������$�]dR��$Ԙ;4��r�A��^�tI�툅&�6��P4D��p�I
x��v*#y�I:T�=�#!�]P��	�(T&��b�ѕY���D�!�dF�����j[&[�Z��3�剨i�|��?E�� `4{�+V<�:`:�*��[�z$"O�u	��=\�"�
RJ��	4
�|�J��<azr�	%Oj��@Ч^�O� A�PI̛�p>A�aB'5g�}9���?ð0;��0g2f\R4�� m�(B�ɫ
�b�I`� ^�RT0خ�<q �۩�r#~"��K�� ���/oc����D�H�<Iq�C�~jhL�)خX�����H�o(d�'��F�S��?�����ۑfM4a_|i!b��(t�C�	�u�n|�t���X�&��R� &��I�Ou�䢷�'��m� n@�IX9p`��������B>v��R�v��%���@i2���HE�`_�<���5D��v*�79��(��U��z�`R#3�"="-��*$�NF�H��'r�$��g�"^�x$��/WrݳQ��*"IE!�A��
t��%�?}(��=E���jRD�V�H�9��9�gԓ�����T�����d8EB�< �l��~E����&"�O��A�;4���3���)��'o�a���d�P�O�}�F(s惝:T�0K'G$D�s�ŖRB��1<|����4D��5��|yB�0ʜ�t�h��5D��SQ�R.ٓ���9����BE3D�4�c Ϲ<�F�C��>��xka�$D� r� �i�1��ܥ}Ǭt��"D�$�2�۽U)�����d�%D� �4$� 9�h�Z_]z�jg"?D��P�f�K��t	�Zb�"�%?D�,�q��}��]�щ��o,ZH�<D����@5T��̀Q�ѡU�d�9��;D�,����&r�"$)��>IzB��SL%D�(��X w�@�(��4�t@�&� D�8��#�2uET� D����i1B D���#W� q�`)p���2R�>D��+��D�T�u0t���U�� 	<D� S��
D,����l�6�۶�Q?�y��H�^�>;���\�\����yBK�	QF���6�A�M7���S���y�%/GN�Q�
/JI���RM���y�a�qT�A�b�%A�\XX7o��y�'�f�HX�i�=��lJW��y�E_e0*{��
>Dˠ��M��y�d�h��M�$�Ԇ�t��%��9�yR]�m�t�u�N�6�6�x"�J��y���(0� �
.���e���y�l]�nn�x㴧M�Ü4���ް�y�,֊M2��1f�J����d��y� ϑkm�Q�f�.%�k 9�yb��2�b�jṕ� HluO��yb��5y�<���N	SX4%J$K��yb�)Rn��Pp-R�~�>�&+^"�y�O�Pn�
1
Y>Lͨ��V�M��yBnSM��dXJ�;IB��RcmB0�y�G�6N�eb�Έx"���=�y2"�]4&=�1#ոwG��ID˻�ybe�mql=�b�Ib�.X��W�yBȜ ������Y A�R�y�OT#']u�2��R�a�#0�yB�{wl���\)`��mZԧI'�y"�I�K#���z�B�o��5�ȓX�"�@�c��Q9�(�����E:����8���1A��Q(N�B��Q~>���8����F��1�ΰRA-��0)t�ȓyx�)����W�T��'�%D��̇ȓ+���;`�܆+�΄�7�P$V��%�ȓ_����)]q�hY #�U@�����S�? �QC�朮yJ)�2&	<.u~���"O�Ec#��yX�Ɣ�kӤ�2�"OҀ@E��<������%O�J ��"O@�8Gk
9i}b �nˁu]��"OF�C�MJ
F^z%�'G�p[Ҽ)�"O�1@�U?L��g��EI�S�"O:���	j��5�&搓j!"�"O�<R6El�N|�ŤL"Lz���4"OH�LO<��$�c�5b��	�"Ol��c&d8P�8�M�j4T$�"O��ꁭ��� ��S�3�`&"O�Xz�LY"8� ����8�"O13��dG �s̛6q0Y� �+\O�e�w���}�׉�	���2�"O��v J_F����A��j�;�"Ov#�ɇ;�
#�ӯ�d��"ONݻeO@/1��PeA?8z�"O�EcЂ�<=ɪ-��O��ӑ"O��q�`@��@h��
�s"O�Luo7I� ��J��)V��A"O�3���#H^�c�H'�"��7"OV���2CP�Xh��"<�l\xA"O�hRe�C�:8�F@��o�`%"O�1P�M�A��`aq�_!�����"OV�;��B�i�AHT'ͤaM��P"O�9���V�	�PQt��?��XP"O�  ��N:�j�p���\>��P@"OJ��%�B� �>��v��z:pͩ�"OF��a�B�&���Fђ	)D���"Ob@:��3R��H[1@�"$
D�"O,	Z@�U+���Qn�3}�~���"O�0j���w=���0�5K��&"Oz��%�ߎs�-�S��"/�X�"O����ԗ����3�C�K	.)�՝|��'�MiS�0i �Ie^�v?�(��'q�Ȉv�֧JQ���"�ʠ^�%��'�Դ�N�>�١�'K�nQ��'$���� �m�)�� 9
��D�� ����
�3{V ��ȴM����ȓp}$�1VS�R��Q��� ���Pj��C4���d)@���F�~|A��oY08��c)%vD]A$�	�ޒ5��TM2�D�2j�}óCʜ�b��"�Ȑa!�_�*P���E��)��̇ȓQ�@];F�%)1t��3��1�:Y�ȓ@{�X�)F���њb�#�dՄ�`P0E!!��r��
��G8�̄ȓ8h$����( �FԻ�g��^� Y���]i�H�-���y���j&r���u�0��t-�e���k�
�{����}�މ2��F�Z�kV�/#��y���t�M�|Jtͱ��-��Ą�U\�꒱���Ō�>U�@=�ȓq�X���0;6�`���7�X��ȓh��b,�B`
�f�"�^�ȓb��8rW�Y�5��m�#� �}�\%��rf�H�PV, �.8�f*�r9�ȓX�.�_}�(�S`�4$��b��y�C-t;�R�
=(sd�v�<�δqZD큃j��f'���
r�<��&�3$���f�N�%�l�KOp�<Y�ٝn,�.C G�9Jǘw}��)ҧE��03bO��*�$���94�P�ȓ93�`bdX�̔;�Ѥ ��S�? X:A
�,���۴*�MȆ��6"OJ�a6�V��u�QɚU��P!"OX�Y��R�QOp�9�Wx�|���"O��vk�6X�0,�Ь'��`2�"O�� ���s�n�ꃱ�R��"OY��G^ C?��p�,9Z&����"O�9*e ǎd=옱ա�{k��#�"Oh����0=�����ߑ�$��"OT��#�[��I*��=����"O`\D�� /'T�*�E�?�b�C@"ON�aP�՟F�2��n�Q��u+�"O~ {�QA��kW�@> ����"O`E�$�I�P�,�c�n��2E"O.�҆6��{�׎/8Y�"OR���Ƒ6���F�ۑ#кE��"O����E�NZ���rI�"��T��"O�Q��[- ����Ԋ]��F"O�Y���ɗ'���0I��U����'�󄗰`�� �!�t�^�ؖ��~�!��)#��A%A
�3~j���&K)�!�D
�nR��c�ڀb�ѯʶ�!�䋒*�nql+m`�%I��r!�$(Jz�rd`�!���c�H�!�$��I��Ȕv�*Lq�aZ�S�!��M#��s
��	��К��F-J!���
r�}Kn�|��U��/��XH!�C*T�$34@]�,Ue�&,C!��s��E��4K�������^Q!�䍨^K�� �CB
m�`e3ĀG�Nf!�A�fX�B�0mk�`{���HJ!�ē�B��sB�8|O�$�2<!�ă��E�D�Quj���Gb 	7�!��6G^��ǥ\�hb�󃢍.+P!�D� o�Kħ˺Hy$Ă��ݐ3!�D�	$�K5��L��m�揊�_!�K,r6���Oėac�Ԭ�	G�!�J?h�~T���^�^���3�A�*q�!�d �v��Rce9C�A�'�C%!�	�\^���%D-l�]��c�@}!����B�.áGј�k����l!�:2R�B�!</ΆH�+[d!�D�0/�6ѢEo�nV�J&���t�!�����fgM�Z��L���5f!�Ĝ"_�>cQf�4
 F�;2�!�DT�u�����=�X�k��ާ:C!����q ��ǹ
2@U�G��Lb!򤖮ClX�8�f	xY�@9&9!�B�j3(���Ȩ$H0�#4�C�A!�d	s3"h�Ƌ�o/&1���H�x!�$��J��p&Iʙ[L����)"^!򤊝O�e��oZ���d�ư`6!򤔕x�b��'K fƉ����)!�D�AkZ�Q�eS�e�D?
v!�D�LMx�j���' 2�!�	N^!��ד��jb�
D��	As��mz!�ޥ��E�"���{O֍�"�v�!�䓢Q��hd�R�\�(Hk%� �P�!�$ʲ3V�׋A)o�H���J�6j&!�dN�oHf�S��	<�ĝJ��g�!�dϠI-DE��l���԰{a	֧_�!�DJ5:�0��-�.����nԶ�!��Z%H��(�Q�O��I`��κLr!��~$8iF�0?*�X��M� c!򤋾\s����j#jzn	(��E�'!�� .E�t�b���4g #7}Z�"O�e��M�&W��T
Q�Q+(�I`"O�U0��Q3%�ąQ�ԭ3�؉a�"O�9�H�B�L�A�ݕ[ޘ�B"Oh�ň�Kk�Р�l��B��v"O�Pv/�bN���0kFx 0р"O$�� Z����d�d�P����C>�[v���I�R"³>�Z�;R�5D���`@��F]^�0tK_5x�<u#��1D�t*�đ7o�,���b���D%.D�����ei�y�T �B��0��F0D��
�Gڲv�l�J����g��+��3D��c�ƘJ4��ʲ�R8Y�Z�;"m�<��y/ mj�������O�
$FV��}=���/�4��:P�G��x��B�����A#v(�@^b��Ey��'�J���+z��p1��98�P�'�f-K�Oߢ:˦�P瞣 �pI�'Ӏ@cF>�xQZ�J���0�'�F7]�ޅP�N�#A�4��"OR|j��PKH�Sh
�G�h��"O*`Ŭ`�({�'�%7���"O`����2)�*1�tD�.���"O8Ui��	uRp��F�r�`���"O \�E��g�8��'L���"�"O
\ 
���,���^u���"Olգ�▔*��y��ݹ
��ӂ"O��(�e�*$�hQPc��Kf2���"OT�["���)Tx���#˿0S�tbs"O.kpiM�q:JEbr�J�[M6�3�"O�́&$�>YRᓇ�ę�"O8U2��N�6����-����'"O�T��B���L��1C	;?|�x�"O�ġ��6Ph�	X�P� "O�p���D�z��q��1r���pp"O$����[)tg�@CgM�R���"O��XWdB f5	�eV16rd��"OxY2��Z����D�u
�)�"OF02�Ϩ|�p��ף��5�ĵ�e"O*ERg�4"V�[#�#f����P"O\u�6CT:]���0�B)b�l�{U"OЌې�^�*�h%�D`�t��y�w"O�1`a*L1y��cpȋ� ��"O(�q$H�</��Q�U炔GV�"O���]Z��WOb��� n�#�!�D�2@�" 1�.(�F	�jQ<,o!�D@%0s���F�O�-z��J�9i!�.P6���JL�"��ƛ�'�!���1Q(�
V��}j��^&'%!򤜰g -���L�.�aƔU!򤏢]��k4�E�8�4`�ʏT�!�Y9tw�MQg�'�(�fJю�!��@F�ʦ�A(]p4�)`ό�j�!��� ��xܬOj�͚�DDC�
OZlt򢟈��X>Ή��"O�Y��
� 갭D�Y�J��*=D�L� _ "N����3y�H4rl-D���O[.�l��FVj.dH��'D���Dǒ5�t���!ԑX�����#D����O�[-��; O;sVƐ(�=D��rnO�-'Ft1P�A'>װ8+2e;D�095�üV�|��#"��v��D�8D��X��@�;�\�؂%��
٬q��7D��ke@�}E~h��
C�=��91 5D�� (�w�A�7qde�a�&I��-P�"O"�#�$��2�p�)�Fۅfۂ�Q�"O�!0i�,���
����SӀL�"O�� "��$1�"�_

�Ñ"O�T�r�/V ha�V�C��!��"O�屠�q�:���J9I��"OJ� ��V (�RI�"!��ᓤ"O�I �^p�(���nx�@"OR�ss$&T*U²e�pn�[�"O�%r�O%2������4ZP�E"Oܵ��J,1bx�e�٥{g8��2"O�*瀖�C �⁋�t\`1$"Ot9� �T��2G�W�x�8��"Otș���sw�8z���03�H-1`"O)��Z<?p���g���?mj�.�y�b�'r��2ӛ��JSG���y2�ƾ)N�����|
�X3R
��yG�a�t}Y��ؐ���BE��yR.�4=�,R�FťiX຤hم�y���6��-��b/�@����;�y��
xp�X(��\!��u�L��y���9�600îC��P�����yԫE(��8��P8��U�$끱�y��}��'/Y:y~h��!T&�y�MWJ�*6Ɨ)$B�2¬��yBAp�J]��F�yH�%I��8�y�HHSpR�.qXB
�.�k�$���Z:M��k��S於qa摍*��Q�ȓ��		�ۧh��Y9�O��ȓ�� 3��O�kEi��lƂ90t��1(~VQ�Uz��u哅�A�D"Of�3��!x�2TY�U�$"OΔ�C�!gy| �c�ΚKT��2�"O*���d�Ǩ�+�(W�YBr�*"O�1�oE�$�d�'׋v�z�y&"OT����'��h�(� �xe��"O�d��Ԇ4ƀ�@�`�� 
&"O�<[�h�	�^�����28^�c6"OZس�A�*�.b���rۈ�[�"Of����n�xm�2�T���8�1"O�X�RB���$$@S�IaP 4"O�x��M߉6<J�0��,sB�@	�"O�M���0I~�5�tgő$�a�"O>��
��-:��]�$&��PB"O@�	"���$`�Aכ%@-�"OR�!��E��2�fd=�X5�d"O���	[	_�R@ա'-���"O�bf�K� ���1iK;e&�$�G"O��񋈵i�L��.S�E9r"O&HP�e\#G��0B��O�H�Kd"O"t��G&|$���C�=6¤)R"O"���j�<|�HH���*!��2""Od$�wN�:m�s�ܸ"*��`"O�hJ����W8�yBW�2]�(��"O�@w�j� �`��=&QpzU"Oh�!R�^%O����@._NX��"OP�*�GӥmF�h����=18	��"On�����iQ~��ʟ��`�C"O����L����ǟ%K��4�P"O���2�R� �X�b��3J�u��"O`;1�P/q,�yqAG1e5n��"O�9�0JPD�X��闙S"�A��"O���0���/��C�46���"O�ԑ��0t�[Щ� � h��"O� ����fا�H�!���Nڂ��"Oi�lL�\�u 5�
��1��"O,\R6��u�tm�uX��)��"O���rG��0����%�r��U�"O���'cΫG؞R��K3 8zU"O|��9:�vM6��$E؜!�"O����E�����S���-��9�"ONY��B[�T�n�q'�� ��"O���kF/t�8� s�6��"O����+��;�I�1;b��"O� Qʍ
Et	S����+RK��yH];*\
t[Z��` EI�aw$C��+9�b�R5�W3p>�H0�Gy �B�	
;�Ќk7#RL�6�c�F�͢C�	(5��R��7�jY���	�]�DC�		�@hQi�X�R����O�C�Ʌt�d0�V��9D�2]s�/�8	ЌB䉇$��0��!{�j\ G 
U��C䉕M���ZP�Z���"�[7zB�� N�4�����;�.�;���7qT@B�	/w��pX���W�FU3��,"�8B��AV���,Ƃ0&JPx���"B�b jY���7n������*�B�0��c�ĩ8	�LB�R�)7�B�	.���Y�$ұ�Ag�Q�|B�I�Z�ڤ1���3>�d���k��B��(V��`��U�@��� 4@U�2��B�	)Rʬ8b���/gA@5��>,�FB�	*@��P��FٚF��R$j�D�B�	0E�����3�ٸ�`بf�TB�	�C�<à-		���sJ�|�HB�	O�dq��(���  l��B�I�l*��`U��U�[d�8B�|B�	������ˏVޚ䪖C��b�^B�I�4�P4����,�D*�扰[bC�ɺ+�ũ�)ٺ�n\�W'C�q��C�	�T�`�i�n�g��x�� �C�(�NA+���.m%!�X$nC�ɆT�v�ؔs2`rC�p���ȓ�t �%� )b�4R�W8mJV����k�mW����bLA�ꬅ�e�l���G
{r4k��ˬ: q�ȓ4d�
A���r�Ȋ�*��8���ȓ!Uj�pA	 �&��*�n
�s� ��ȓD��a)׽Fڰ����VX�&��(�a���^��J��P���Z[����~�-��ʆ"��q���W2�	��Z��qѢ�$H��-�����ȓPSV�����f�hTE��0�����?� ���Ї6���&�?5X؄�)�4�#�&�4X�r�$��p)��?����g
u��=`�'�$j�ȓ'��W"��n�;W��s�rԇȓ*;8]�@�N(iPԍ�T��2��i��-E��9UȚ,M�XI�g�5.�^�ȓ^"`Q�J�!R���L��1D� i�Cن�/�w�Tt��ɊV�<3��5\B���*�3p��|��LJ�<��h�A�|����R�y��zy��'Z����T�kl �{%�IO��'���`�8d��H� �*��y	�'"^̳r�Ʃ4�lE�� ͝#j ���'ʺ!aWk�>��i� �m��'��p"��6��[�/,qf���/O���� ���C��Lp��S�$Ť@��"O���3,B���i6m��v��]��P���Id��a�_+�5��ƙ�v�6��C�<���0>��ơ*�tb%H��~!���p�<ahV�wm�%�T3�Ig��p�<1ӌO[|���䂗Pոiy��h�<٤�
�
Ѳ]��Gזf�"9��E�Ly"�'��`�눜-{"��Q'l\��'#ƀ{4��o֞�ȳ(� 8\�O>��%��;Ӗ�Be�ɶL�4`�Ì��$�˓�0?Q��B&>:��A�<}F�9��v�<Q�I[�D��P4k0b Kq&W�<)�H]����Ɲ��v��J�<i� ^����d�ҧv���BE~y��'j��x�c�|�waH����ϓ�?y�yBDC�?����v�\1w�<��J���y���"�hm�pM��r�r�ٰmɶ�yb	D�~�*ذ�Vj&�� 	#�yi��ҾC��M�v�H�NϽ�y�BK4Nv�h��P�
�l��©��y����m�I�m����!�"B��y�';+FMP5�Z��te���>��=i�y"M�UjTF�&��M㭊�y��
���*Z�L�]�w�R7�yB�M�vw4�;�!��X���i2��y҂��x]zT�Y�V�� ���O��yI�<S��ېGP�YQ�}yD�
�y��f4�3g����p��g�8�y�Aݝ�j��Di�'�lb�$���yr*�&f��J� ��R#���y�CY�/bp�3��׳"� ����=�yB�:0_T�!,�8����J�yB��pCP����µ� ���;�y�#3al��b�d)Q� �y�iW �|Q�"f�;��͂���S�ѹ�V�[��� b	 ^�\����3K��vp����툱�ȓW�R�@�B؉B���*ѵ0�L`��.g���QJ��1��L��͖�J���X�|�`4�H�2��<"t�Q�z�D���0-r,hd�p%4ɡ�O�N��`��[����#�D(�t�,M�	��(�ȓޅ�3*]P3x	n��u"O�X(7'��v[b��$ۮ����D��I�'|,m�0F\+r�� t�ٶH�����"Ov�I�n��AQ�@�K�5j�{B"O��R�6��ɦ�({��m;U"O��{��Z��\���L�HIa�"O����	m�`��'��J�W�P`�<�R���]�Si�.v�b�����\�<��]�|9��x'���W���{p&ch<	C�*FB��*Qn�����8�?��'��y3a�͞e�v1p���>%�R�;�'����J��H�p��5,\��'ØEJ� Q/Wj%�M?!p.�I�'-$���[6#8\"����`��'h�Pc�n��zHp�#�9��y�*OX�=E�ĂӟuI�Mc#O�%�<kė
�y���ġzᎽT|-���ۢ�y�c�9:$DP��	@�)pa1�y�h�#<��lq���!c��iI��L�y�!X�4�8�'��Y$��Z��y2�^'0G@cW�R'%!,��yr��X+E���
�h�����y
� 
e��H�2w����X"x��`B�"O�B��1OAC%O$<��U&"O���[>m"0�qa�::�&��"O���S�W����-��"O�A�d�<��M�R��R���2�"O"���^�
�����ss
mۆ"ObDHWc�M�8H!�2m,�����d>m�'��	��@�iG�b�����J9D���aK�a��r�cB�;�Dx2�*D��sΈ��[o��Y�� �
,D�t�QJ�_��L��Vn�,��+D�t;�- ZD����?{I���5K)D�����>�sQ	V�"�̋&E2D�� ��C�/�
Qc��3`��0�;�I_���S%�� j9@:tyge�:$H�C�InGH �!k�f��(���Y�k�r�O�<LO���*�Nz<c��/[��t��"O��q�ی\�:���M�#�2��S"O`��4��G~�(�M�B���"Ohd��N\�T߬��ҎF?|�؈#P"O4����Ѿ}��%餬��O�� ��"OZ,x�ʕo�Ό8ŋ�3"l�y��'��n �X`��҈_���V����'�a|b])��s1 E�Z��M� ̓�y��ʂ"�����I�K�<,�!ҷ�y�ÔL6�І"�H��§�yO�0H \;�J��oBH�t�2�y��|�| ��@6p���j�D�y�h
G�P\��� V<��z�gH���x�/�n�꽓�	@.d|�Dɷ�Y�to�Ip��`�K�!z&�#'nC$�\;a�5D�� 0��*e�4ĨQɟ�IV�8d�&D�Ȃ��ō?���7���%�@a�`(?D���!�ج5�����F�*�+�=!�Dɤ�D���dx���@$^!�$Z�d��C�
A�u���u}!���y���;�ԃRDa3u,[�a�!�$�.�bX
��$�K9J�`}��' ���0n��&�6Qr�ǌv�t���'|I�@���X�qe��V�.�'�8��B�I�B�b5ʗ�%��Y�'��P ��R*5��Uؔ������ߓ�?��O�b�#Ք5� �)窆,u!Z�B"O��1DF0���/R4CmpA�"O`9��ᓠs#����D�6]jt"O��u&ڮe���G���i� "Od�A���<�գ'� }rޔ�C"Opk@��-3���!v%W�OY�I�c"Oޔ2Ŭ�o��|å�I2;���T�'$1O�9�o6�f������e�1"O��#�!1u4�@���\��=��"Ol�r��Αe6��F���P̊�"OL�-�.<b�xx@/ʬV��I�W"OމR&K�3����P�K&�� jW"O��(�ԕ����b\	y`$�AO�T���0t�}���F��$i�� :D�(p����-QW���Z��t��7D�䒱�� t���'FD.K!z 2�"D�\i'�
zG�q�(mc�A�  D�@jC� �S�*����!F���1�M*D� ���ҔF�(�iFA��B �wm)D���㨜5s5��8&)W�;�2L�Gg#D�� �H� byz-chէ6״����>D�pc�N�d������{蚈�>D�� b���G��ZB氂���9U��%��"O�x �w�p0��6��	R"OL���/�]�z�k��LX�y"O�4si�s����a22���c"O���1GQ"�h�9��Y@P�90"OB1���Y+0$b��:�I��"Of��A�M����΃TvT"O$P24� �L�|;e��N�Da5"OP8�d���fi��O�|�p��"OBɹ��Xha�t��5�zT�a"Ox���qpdM{�m��V����""O�8����#U��P�:2Ƞ�a"O\�(tKa����(�"��q"O���h��K�\c�-N%<���	"OLIt�<cr<�;�I��J&p�ʑ"O,�1��7kA�c�N��Y�"O�D�Ů�r16}H��LD< �a"O��!wO��;��9[F��N:t���"O�,P�Z�<�£�ݞb &=��"O�P���>6�h�k�o���!Zr"OsPH�q*4k��K8�|�DR����{�"�9ᜀ,��J���'*B�IvO��JS�Z)hb����C3��C�	:��L�D��^�IȂn�Co�C�ɐ�(��A�2��钔��0�B�I(��#n_�hw^]�%FP�CΰB�	�6�8�7L�2�4x�͛�A��B㉀��A�°M3�:v�Q8S��'�џ�<�	�9�IBC�n{$K+d�<p�9`���ۄi�1�v+�`�U�<�&"�6fHH�$�8ʸT떃[X�<� c@�V���'
:XG����V�<�Ѐ��$�A
ҋC�V ���m|�<q��/ӨQiSCp�T��pl74�p��`K�[,��BE\2r6�� ��X��b�'P�L�b=b�j�;�hP�,5��i�
��ta��3���F�3fi���b�ʹ��	�^�V�("-�N���ȓ:��=M�>~qq��r|�y�ȓ����VJZ�!<�I��ώ��\�ȓ��}""D���(�!!@��p�ȓ:�V�2�
��ci�E��܈�\�ȓl���&*�t��S*C�ǒ݅�S#عk��Z	u�,�z�� +�P؅�mܨ9����<��"B�t����C�h�����,�Zے Μ0jI�ȓo�@�S���#k��,�q&VC����ȓ�hy���)�%�1'��>����0����&�۾'v�Z�g�&�|���u��h��ĕ;.�"�J�N7C�蔠�d�'N��I[��H��O��Z���kƜ�r�"x��6D�0��'O��	�uj�;S�Zi2.1D�tc#���1���b��Z�<�F�(�0D����&L3J/����AD
|2m)$/D��b蔃v���I������k+D����șP����� �`��Y�p-/��0<y#��#r�)��k�M�б3w�I�<1G�G;�>�ç��c��1�#��A�<���ej,T��KݏJ�E`b�~�<�5��<+s��`��H'tNZ�#S��`�<q2%��\z�
�jȹG����"��Y�<�n�>[�Hi��aH�f����W�<�'@�i�2̃`� +(�L�ua�T�<q]ڈ���M"�k�OƎՌB�)� �����
mt�a�aG	f,fH�7"O$��6� k�� Wm	�(��e"O��bti�v˾D�R�O~��lSB"Oĸ0�X�2�`l�Q�,��9��"OZL����0��<0 ����� 7"O�����A�#�b�s!
�F���Aq"O���̞;`9����� ��8C��-LO��,7O�H��cM1_R�K�"O���+L,<��(��ǫo ��P"O�lI�!�;���A#I Tk�H�%"O�YI�e�8]�B@�v`L+j���"O"��Ī��y�Ibsb�0W�eR"OL�i�\�p5� 7UcB9�@�'!�$��Xy�צ"pW����'!�DͲv���9P��[>x]�	��J!�d^��,�%��,p�՛p�],!�ɽ3����ŢAq��Z��2�!���9�P$ta�2R�U3�P�E�!��0�H���ӌ6̠̒T��:W�!�$PZJQ��-�,4�P��%ّ/��}���,�3�	�JT�"��(�t�3D�@�Tm5W��u�`��}.�dI��3D�(�W���F���sgK�?@*�ۑ�<D�,��iF�A��1.MˣI;�O>˓@�f�k��BVi�5+�i��J/$�#�'�x�!�̥,�x��c�S3 	�'Iv�c2�ý>�va�C�S�xl$� �'��5��%2!.��Ӎ�sgT���'���:�L�{�8���˟�R�Y�'��P�b�>�p噳X�]m>H�
�'�\� �N�	���u"WZ��8���?ye�r� �L	}�<)E�ǵ\��L��'�ԈW��1|
�tI����Sn�<{�Ƙ'�PCAI:o�T�L�W�(�'�p���*�LiA6σ�W���;�'O(𘗏�q0����8��E�'5���c�m���� D�)W����'ɰ��g��m� yp���*��
�'|��	�G+���'��	*���	�'�k�$����r Ə/l<��"O6e���Ėx�5��rQFds�"O� 3�c�N�J��[HOj��'"O�����S�y���T9b6Ĭ)�"OmK��Y�f=~�J�i�:xm�p"Of$:2��27a6����½=(t�H�"O��S��= �fi��%�;`1QU��,�S�i:t��A$h�R`��@c07�!�$A��0�dI�	`��oF!W,B�ɢW�H5 ԌB-2	�$���ߛ �C�I�"�Ha�N-p &�J6��
h�pC�	 >�f㕵���iA-HY_�C�I���јėu@��E�]�C��+�*U(A�E���;q�:GO&�O,˓�0|�wD�A[�w�,�N��bC�<�wOݟKTؑq�/L�a-�#֦�{�<q��ND�� �=x�d�sK�9�!�	t�b���#NO$�q�,��s�!��&xf�,(��q�&X2Dk���!�߆ء@uGQ�1�xUb隅y�!�$�:5����.��9���X��@�l!�dŏ0�QCED��A����F�/U!�d<q��p�A@�uWz%#��ST]!��ڃ����cE��h��T�9�!��M�tA��7��,X@����g�?]�!�� ��S.D�8n�e�g����!d"O�ym�1��ӅᚑR�T��"O��B�V2T����AL�x�8�"O��У_����:�B�=CQ$囒"Od���nZM��Q�r�̷�%k$�	m�O�x�7¹R�&���І	�>��'���pq��/[�r� 5��JE@��
�'����w�J�4ʖ+�nĎC����	�'�� 㰎�l���C�A܂A����	���' �)�m�'6�\���9H����'A��R@V<�b��@E;9V�)I�'Ȩ|�D*_�c��@���2-n�C�'G2�1!���@�tؙ�O�2ٜ4�
�'\`�2�C.BD �;����*&~p�
�'�d����@�J�7埲��[�'k��V/Ȫj���hvK��D���'�j��v�C������ڄ�H+�'��fC��%�hda�H�:F(i�'�����GĂEI�G�	�0$)�'�����Lʍx�2\��ҽte�0+�'��y	�.�*�M���aDʠ��'qL���춀�+�j��\�Ƅ �'J����-�$#�nh�aF��Q28�!�'Ҙ�@ �" ���	�Nݪ1��'��3��R1xlz���t\ݘ��d?���:S�M�)�Z��g`IuN]�F"O48�C�V)a*A�6f�3k>@X��"O��1�N6c�I�OSa'���"O���"o۩U~�����V�%"Oހ@d22"�j& N&4�m��"OXAٶ�
�?1��:��	��bq"O@=P��FJ%ЖA�j���	�"O��HƎ1p�j�8�o3y���;�"O����C� �n����S����"O*�X�,ƁL`v@�C<[4�c�"O@��6Ƃ�i=�B�!K6,"Υ3"O|1��Y�u���)3'A�FE�$�'��ɱ{6����P�d � Z'��k�0B䉱^#*�q��M:$�X��Y/2��B�ɚ9��PX��2���[� �B䉂&�H����w���B
HC�I0�lqA6A�e?��A5hW(C�	5@P�L�&G�mw��d� 
��B�ɟdt �Kv ��&d���oZ�p����8?� .�8!8�I�gP4_rB<+�mFM�<Y���+ �XA,Ąd��-sŏ�I�<A� 'ix�k���y�6M�bA�E�<�)Ɩd�Fe�1�<	�89��Fy�<�(��p)V�`�66��dq��Lr�<���Vw%����H�X�����k�<����8e��! �}��Ҥ-j�<q�Y2�@PIZ3"8��JP�<����[�6S���2c�4*R%HH�<q��e�D\���-$����$*UC�<	Q�V]�9˗/G5	h<�N�d�<���r����`�z�Q�q��^�<����u�Ы�DEL^��Cc[�<�����<|�Ah��m���T�<9�|0�z� �g�ֹ@F�O�<JO�.��b�d��	e�<�Ǉӿy�C�C�V�,�+�� d�<q�֝kb����
F���i��	�^�<	�o�8~>ݳf�Ǩ'�e�b�q�<���D�5a��"C`��w�J܁0��m�<� =��BM*�`;�k��3Yr��"O.ݙG�
��@��*�FX��q]�З'0ў�O.@��@KI�c�5j
J))v@�x�'ǎLcS�@&x�1:VJ�����'����X��蜒bNP$���'��� ��S�|��J�L̜l0�Q���x��D�&p��Al@+oo�`j���yr�üq֎-�1 Ϙ`:|��iP�y���t���(ƻb��y��O��yr�-:���:&#��A����X�yߌXI���A"آM�0���&��y2&ٜEު��Ԫ�Jnf!��k ���'~ў�O��t	@�Y( �N��-0Z����'��p�͈(,�|A��ڹV�A�'-����s�E
����k��Qc�'�?��j]<V��q+��@,<K�x��$D�4ze��=~�� ,m��kы-D��Ök�
� \0��\([@��7�,D���Ѓ6]�v�����{=V��a*(D�@�C��Yw`%;D�D 3� ��&�9D���FӢer���0Pi�a�;D�|�&�z�A�!���\A�"�$<O�#<�P�ȹ�n�K$�ЛR���y���G�<	��Rh���N�u\�7�h�<�V@>:� �'��h�V�R�l�<Ɂ�L�1����^ k���R�<�DôM��x��X�G�p��EO�<	$/�3T�h����bA:�D�t�<!!�I�4/�9I��]�4�Z�g�Jf�<Y7��]���3���fIԁ���ܖ'~ў�>]80#�B�Z��Ũ9X9�D��1D����z�0�ԀCE:j|P��,D�xbp)^.C���ns���J+D�@���O�6![�a�@��@��(D�d1����UzT��I 
����&'D�|�wkZ"jlPr#&CC�ZU#ҁ&���/§C�x��A7AL$a�	�bT������	�6\¬(׵?�\�2�K(>B�	�O���M�3.�6��`	J�B�,}؊	pC�4�l�Y�Q�g�B䉓%���q��|�ub�-ʇɲB�I� 2����6�J�`r�&�TB��&u�ؙ�3g�W��dQ��I�a����$8�w/�C�k�2�r�H%gr��E{��'���97���X��R��4D��=y
�'��<QOP=SI�]HPC˅_h�9�'�N�)�&~g��� ��0�l��
�'��u��ɜW�y���*U�l�
�'�<���#������Y+�e�	�'���au�8%�Dj �T�](
���'%~��&�):�>p�'��7� PQ	�']J0�0m�z�ĩ��P�!�\��'(���I�d<�F����,���'�2PSqjD�J�,�P�&'	�x!�'G�Mhq�O�X��8��EV�y�p0�'�&��IE�W��$�ta	2[tm9�'X��W��b3�D!�
TI��Q�
�'B�Y3���st*�!����r2��z	�'l�aKr,�5t����qa�W�pA��'�`��.��`��蓯,�8E��'x�l�d����RQ`c����X���'�ڈ�����p�"�*���'���c'"6}&x��.lx���'\�<��ؚu������L3������ E�C#In�<pg��IM�h���|��)�x5��5�<o��A�ʔ<�XB�ɺKfp����F﬽� bHJZ�C�ɻ2,�H�f�ܷg�vY�w�ǆh�C�ɓ��\K ĚdXv�i�K��C��T��a�[i!����/S��]�	�'��y��n,Q� �1����'O�فoP�X"\Đ"�-{��p�
�'B�)Y��F:e�v�P�F�l�� �'qv�;�h���*��Mg�'�O�%c��J��ѭМ���1�f��U��q�Ɛd�(e������k{�X��"�ܹ���	<���>T-�u�X	U;L�ʄ$x8�m�ȓU�Ry��!��QY��$>+�`�	˟��?E���7�F
�� ȷDY�w�ڥ��"OB�Z�o�!S�	�C[��4�'�ў"~�gd9h0�yj���:�x���y���E:�!L�s'(d#$͗�y�"�>ֶ�"!d�#��e��o��y�E�'-� �J����k
S��Py�����^�qv�Є���s� Bb�'��'t���Hr�BX�ҁ��� T|┐cK�wh<����� ��D�iGpc3��?i����O.牌,��"Q���s�ˉu��C�I�=��!$��#!� 0�d�$g�fC�I0Z���A0�L��Ɗ��HC�I�PެP���9)r���E�*G�LB䉽9�ЈZw�3�@���[9zv�C㉂�ة�RCL�K��]�5��Næ���n�Ey�fG�1��#�r!����'B��C7b�7�Y0��š#<hL`�'�H��/îZ��mkaHڡH�'���S+P4B�������ƕp�' pI�!g�n�bB��'�}��'�h�H�N��L)ңG	Y^,����y"΂�O^rH9BJI0&e��
�'R�˧H��)P��e�?�l����'�P�#�s<��3�{�D�s	�'j��`"&Nn��S�C?�j�'u.p#���~ Hd�+f��S�'�b�j$o�T
�öˍ+���
�'+����O�v9�!�$�L�
�'�|�j&UL��K�k�Ji��'l�K�B�>ʁ`���*�q�'�bh�d;�zԺ���7[�����'�� ���J�.D�pg��R��u �'�Ea�ٝ�x\S�N�Qӌ��'"p]��-s[���+מr���'�u���K}�Mq�b��
�����'¥I��V� }>��,�r�,�����'h`�YD�фD���s�
��3�N`��'�$�w
^oA
�Y��S,�ذ��'�������>q���f_��X�'�p�ǨA�}r�53��T��S�'��|{�Z7r��Tj�� Y3n5��'jh���W	!�^�[3��O3����'�4�SCʮ4P�A�g�үC>6HP	���ć�K5�q�7�T$K��qP&�g}!�&���&�� >���1&M��!�$�����"6AǞo% l[�))�!��2S���R�h�P��)�&Y�a!�d
7�$F�ϘU`*�y"�PFP!�$�0C�V�@T/_��4�vjХmc!�� ���Soq۴���t��l�Q"O��×��2����ȺY�8��"O:uS��W }�vi�� M��E"OD��.ǧ.��<���Ֆw��#@"OD�h�J�b�B%i��]�q�"&"O=�.Z�.I����9Ϡ�Z%"O�A���ƕ2���D�8�j͘�"O�us�%>�X{���b��Ȣ��'1O�I G�9*�@��	�"O<�#T M�F|~�Qe�C���"OLh�b�ׯ-|���%*�Da��"O$��T�	�!�h�AӒH�6u��"O�Y��ၛ<���xѠ!0����2"OLX��#� <���ɇ=+|&��"O��*0	��s��y�����QE���q�'�I5K�\����	6KanA��#3>jB�I�!�T����)�0�9'��GDB�	�%�\���R�%Z�刷.֮��C�I:����D=wM �7o��C�ɨF0�PTi�(J�P�eFTAw6B����sc�َm4�(�V��"B�ɲr�,�*!�Q�kXE��Ɏ�p����d�O��	&�(
 c�)B�"�S�΍�#��˓��<!�Ob�� %�=������/* �5 �"O ���K��d���@'�?�`X��"O�ՑDAO�a/,1uc[�C*��"O�x�A��)qg�4!'�I �����"O����IN���r�ڥ5T]��"O��ѩ������G��Ҁ"a�'�$Wj��"Bg�+f��Q _�qZ��'}a~�ꔱa\J�hc��92�0H�����<�O:�Q��K����E_k��T"OQ�C�_C��Vƕj^E{�"O ��`A�4{��ChD�	UhPg"O����m�2�~��'R;RȀ�"OJ0��X1J�8 VA�N=���U��H�O�}�%R� ��aC�;@���'��'�J�H����@j� ���^f� ���?Q�vB!���6I�!��i�Mg$��|͔$*�*M_L��Ytc�t��ȓH)h�KH��C��%��/@"la��H�lm���S |���H
� �Ɠ�@̓���:G��Pj�BJ?�İ����O�#|�`T 0�r�^�:&�4$��������p~���n舷b�1�\����� �?Y�'�pH�wJF�c2 
�Ճe�L�
�'q�H#��+t]rT��nU�Xi�'�QQG��s�tи!��|(
�'��#��Ͼ,j�[��X>4	�	�'u�<���ãM��T��F�<sx�S���O�˓��DG1,JQz��3i˾��5O˨f5^B�<a8�!�ŘX���*�!��B�0>���ʄ�ӻ ��=C�Ǆ�&C�!��q�����FقA����5K��C�I��:��J1Ti��mF�D���-\āf*�$�<��؍��}���G�^��PA�!���XS�{�<SL!	P���F-��O
oF!�D QC��EE�1��}r�/�K/!��Em,� ��<M"z@�!�G!��/��p!i���q�l��?;!�%�ܭ����&	�"�L�.r+!��F+t^��tAֈM0�����&�{�D�4; ^��bn�
*��eBğ8b!�� ����Mƪt?��J�܇D������'���X� �����P��Q1Q	$>�!����};Ɓ88�" 2��A'>�!�$�0��J��Bm8�s�C��!򄟗7�ZP	6n�.[N��2iA9[�!�D���g��N8�l!�(�2!�!�d�@�v+E�6.�`5�G�=�!�� k�4�"#��l�:CEԞ`�!����P��Ȅ�h�9	�m�}}!�d��c���i�_r��aR�!��D��4�h��+8��(%g�!��V�d�P����v%�zҦ�$�!�$�4b,�EM�[<�����R�!��������*3�b�z��ߤ|�!���/��1p ���6��ɘ2d��:�!���I�B�ى&��Iq�V�!�Đ=o��\��Iřh%s7)Z�r�!򄔧RAR��&���JX��iJ�3�!�0f�2����Kg�P:&�Ȏ5�!�D���2�*��\�.�@X�eٮ!� �?�)i�nF�x���+7�
T�!��NJ�C���N���ӵ���;�!�$\�Q�����1�b�
z�!򄙍T��Q�B��/s�VI��`��!�J�NR�q�ѤS�c}Π��M5s!�dZ���� ��%}��D]2k_!�D�8wp ht^m��%E8ci!��x�4Prf���T 5{��F"c!�D�u5��pc�=8�	���(!��
�<�braР	�IP��"OP�K�m�5��](Q��6#t�9�"O|����6l���.�:���0"O�@�瀷d;�q����d��R�"O��3��9�\��%�37����"O�Y��t��=�bDG�B� ��A"O�ih�`�?�� �#�Q#Dؘ=�"O~bdڌs�*A�%�8E� �Y�"OJ��LO�^�ҌY�� �#���� "O��O�@�>0&����E�g�<��C܆;.tS*O�NQ��h�Fb�<��&��?�0T��-^��l�T�Qa�<�!ܢ���8��2([�<9$�N�h��-�VI"�"�Q�<	f$�%�zu�W�%
��.�c�<ieJ�o|�K��
A�\� g�c�<�3�D>t �E�0-[�V�t��!HW�<)Ra��7���DJRM)���P�<����|B7	�/R�Aц��u�<�rɁ�*z��af�ެPd��X�<�! ���½A���L�r	J��U�<����_O��S4���I�t́f�TT�<Y0	JPcp�ue��ϲ����e�<!㊚�2�.�P��B�\>��͔Y�<�f���"ʮ�;$@Qs��	',U�<�N]2\�����B�?hp-y�N�<٦c�2ܴ��t"K����R�F�<�&�@3tz
��󢖕sEp��p�~�<Y���5����[���P�6�\��ȓH"@�ԌU�&�Zth$�P�t_X,�ȓm�V ��Z V�l��A�
[�p��"/^�#э�8�(�5���MɘM��b�V�����U�E�;:�ڰ�ȓ,��1�aBQKҰ ;𧝶CV����}r�����>�$���}�⡇�S�? ڝ�R�J�sS�$��*N=+��`"Ol����+D��+Ӛ�\Y�"O܁yI��Y䴈q7e�3f��� "O����Q mx�Xq�#ݍ�B�S"O��� ͌�����j��-C"O���g�X��H� Ę|�bT�"O@ͳe �l��p��N	so��0�"O�i�4�مL�Zu ܽ 54I�4"O�� a�j�� A`�ճoޜ�R"O�e+�cձh�\�D�څx0$26"Oh���O���34f֧�(�K$"O�8!�F?0(P@U%8`�p���"O��1�Β�8%0��Չ%۸��"O�2��J��xH4��:u�"OȅA����<:�(�0^�*��""O&�a���e� �(@@E��"Oe�V�q "���S0#�6��"Ot}��lቝ�&o���V"Oލ��mY�O�$��vI:u�f��V"O�
T�D�RMY�H��g
�H�b"O�\	jܥL�!ز[��RX�b"ON�%!a�~�X�J�za#�"O@D"�R2OO�50�������"O(�����1�j]�ť�I��	��"O��"/�7X/&�:���+X�N�*7"O�V�؊��s�L�>�0BC"O��[S� 9��AM]���A�R"O"$�1��I��M����)�ֵ�P"O`��Bϊ���!�C�y�0X�A"O�Lq�3u^�) *�<�\ �"O@��(��dr�Ȱ�b29h���s"O8�规Y#P�ЁO��8"O�L�%'�$u�Aڳmڞ({�"O%�Ff�]���z� ȿ:��Y��"Ob��hV8��ysΙ�����"O�9���`�`�;���G"O���Wcܳ&&� �1���Q�F"OLp����z%hUeD�3s"O�qS*��h�,��b��xGV��"O�i��×,d���x�[+?b|�F"O�m�BN4:UY�	;%��"O�|�p���r]b(����^�r���"OD��L��6��P�tL5y՘A�!"O���g��T�Ѝ� *T�#�|Xx�"O�5�#�ij�Yቔ�o�N4ڄ"O - 5)_%Z�:�Ш�0$��`H�"O�QFnT6,B>�AA�t13f"O�M��h�:��E+3a�$i����6"OH�XЎȯ{�p�	"�ҷ1Y�}��'�6��d�ƑA�r93�b]�LH��X�'��A�։^&^E ��sJ��H��9�	�'��@�2�)��D���A��-�	�'����aDL҄�.;����'�����-��Q��	#jR�c�'�<m̒s��|!@�
�Ni�}"�'Ě��e��Lڼ����T��4��'��]�������R�>�f���'~P��@kؕO^j�Q�H >d�q:	�'!&��N�5��� S7?.=K�'��9��2��EAB� 0����'S�<��W?E���1��T>0�')i!蓡d�.Ա�
F�D]�	�'���$߰NQ���b'OE�!K�'��u��l���pP+���:Q0MP��� �H(B�^����'Ꮃa�h��"O��Se
A]0��� T
���"O�A�I�69m���O�"�2��s"O���i��g�Y���'�]Q4"O��� KD4F��2�,��	�$��"O�ɂB\�CX�9F�P�z�n�"O�i3�Vm�YR*���<" "O����n�,+2�PA��6l�����"O>��W�	A�@́�a١-C��sA"O����͈#"�X�A�/�2PC�q+ "O6	�P���8�s�H�/6L��%"O�I�R���L鹐^%7@J��"O[k��,O�2�R6>7�c"Oz5�3Ȟ�=�p&��Z/��S"O�z��"CV\�B���$Z���"O�a�C����0bh���)D"O�����b���{��1J�>��"O�Cq�܃�J�#al�"Q�i�"O���,_ �*���I����"O�-�ǊV8#ˤ���N��KB"Oؐ�S�Ŵ4����N�,���"OPX���g'iʴ�O�!&���"O�!��Iz���K_	�E#7"OL����
��Hb�A��t.�:r"O �!Q�8��ɱ�%SgZL�"O<�IX�|�bp/̎<Y:��E"O���f�>t
9���	7#�Uц"O|�B&N �}�����Ta�"O�C�
i��"�5`�Q�&"O�)Z���1٪���K;Y�B%"O�����\�H�L��FEB@����"OR(2nI�j�"���A�;M.y��"OZh����2�t��C�I���	�"O�y5��!x�iB'�9�:�"O�˥���%E�A��&m���%"Oh4�
�b�J�U�%���i�R~B*��<ɍy��������Ɓ?�n���NN[a!��ъKu0A�_�R�S�� /+�5��R��cAH@it���l�
�� c4�4$�,���&�R�Buh�.<��)���5��Y�'��	�%�1��|�S��@�`9*	�:���䎁X(��ul�
n��)���("�!�d���\��cג|U��`��1�� ����?��O^"t¼�Z��(i��d�;D���p�Gyy��2��բP����&,$��{؞(�3�]�Sl}�w��mTȻ��6�Ov�ͺ��L�&ڜw�_�FP�ȓc�:!�'���t����aA,h�TG{��O��I�LS�!l:�A	5L5�%��'@�D3Vn̥ �ZDk�C��2K�e���'q���S�0���N�*.��{�'}�tXr.��g�$��͍��D-��y�Z�,E��'�A�PH�&Q*gJ�0�!��'�B�1p��CU�!���Z\~ ��'ߐ���m ��q���֕G%|��
�'�L� �T���aE �B)0a�
�'�h$"��=��M�O��=�. �	�'�>T��H��zAj�A���l^���'yDa�qb�O�
�y�I)rT��'.Y�Н2��0��P_ ]�'�ܘy�nן@����`�
�n���'���R�#NP�Z�8��7Fк�'�FIv�/��Lꣃ�H+<D��'6�H�뒑�$q:��3M�<`��� l@¦�]�y~x8P&F,�8��f"O�"G���;�M�1pq�(��"Ov��t��Ԙ��M�*Z�q��"O(�8qlP+I|-B�Rx�kU"OH���!ڽ}�=�@���%P�}I�"OD�à�N�:a� I��x���a"O�L�lQ#9t�g"��,Y�"O.�`'��u�а�A�f�ܨ��"O\��`o΅&���r(Լ9�@�KC"O�a�Ӂ\3R�NȢUh��K��]�$"O(3�+Ei����2-��@D��(O?�Ɏ~bj��+2l�����?C䉠7���2wI�w��)Qf�&m��B�ɉ��5[�m��@%
�`��B�		h�H����/K-ԀA��ȕQ�&B�I�X�B�
�� ��g�iYR�<ٍ�T>co[�>RT��*�e#8���m8D��@��^��b�䘸kM��1e"D�D
��W�B��4#Z9ִ\c�@>D�iŧF�@�P�3�-𰼈��>D�|�0��82� ���"��%�rh1�OBʓj:�)rKĩ6�P"@�18fX1�ȓI�@C��V?@�mF눴N�� ���������Qo(�����L�ࠄȓHX&�I3�V�t9�$SU	X�H1�ȓ1�v���FU�f�t����1B,��ɨF��:|�����dڝx:�]ے�5Tu�B�I�?�l5����E�|�@� Τ+��<q��T>�XfO�,c�`�&b^=�4���'D��#4�;BLd}#��֢ ��p�pFF:�(Of�}�� �*�z��T�r� b�^$�xD}b���֜�����/Rt�p딋�E�Ksa~GJ�d�l�eY41���#Ŋʵ���=��|�0�|��$���(���/����ڙ�yb@+Y�1�#�ٖ1�~K�n���~B5O�b��' �h�9D���ipTQ�E��~��ȓx�$i�X�P��ÇݳA�>-��L���h����f���A��Š:�JA�˞G�ay����.h�ޑ1�����Jm�#�^ C���yO<yq��>E��'���4ȇ�l�Jx���C�.��!��'L��Be�h^���IX\$�����'nay"i΃4tmiM��m��U�1��
�ē�HO��D�|�����9�T�i�V��ce��yb�Z)$�����ϛWE�8p3������y��d3���/��:6�)�J��t@�NZ B䉣.jm ��/�TŃ�ͳ\nC�ɇ"�~�Y�^�� cq����2��������ҟD�#(��7ՌE ��/v4@U�d�,�>�O����da��c  �u���ە�I�1�O����9dH�����$|�q�G�V�<�JB�I�qN ��w�P�9��RDB�V}f6�%�Id?�O-��MS#�XA��`���)�T�"�C�<@FE	�F�ђ�Ш/�r��vD�<�������b��b���Q����P��#J�!��"O�,c�LޙMʘ#,߸E8�q��$1|O�J��+��ZVJ�0�l �8O������Q��$"���1A�Pka���zRnL_̓kn.`���
a��=��XM�Zą�iܓdX�Q$��hj�li�-g��>	L��F���S�&T�qcN�x���1��y��Ô9��@b�m�p�e�R������6�S�O��iɀ��O���)g�q��Ě�'"�%z�DE5^[FY��ɩ_�m�'�t��$�$.QH�[��H��`Y��� �Q3 ��wIX�a�p����"Ol�eL �BL"A��@��HȶOL��T(kt��d�� ����aM��J�#�'21O�32C��7É=d �F��t2���]��~��)ŗ�h���`�t�e �R���p?)�%ҢX��	�/��\�~@�f �Z?Ip�H���'<��|�g$�/���O�.s�����5�O���OP�A��L����d�q�.�S��y��Q��м�cdea�%@��+�(O�9�c#2�}S���Fm�.b��ۣ��}��t�ȓ([�=� �ɍ;D��A�D��4���E��k҃^R��]�4��(�(0�ȓ{�hE��&��?�ʵr f\~6P�>y������ة�*|h�/�X��)+�C���y��ݨu��1ԀۜS_��q(��HO���Іr��@��Ϝ+N�����M�A|!�IP��[�I.}B��0ˉ}!�+B���M�!0I�TgSQ�XG{*��1;7l!.f��Qw�طޞ�h5�4�D3�O�P:���*d~�rn_�(t-��L~��H���I�zh��	¡�`4�vc�HB�I�u$Y`��N)I�<��$��<Ki|� �'�ўH*�5jt}�UA�=}�����P�<!�,���5��@�0����P}�|ri(�g}�-D�2\��g*"����3��,�y�`T(a`8����ݹ�Zi��D ���mX��2擩}��%@r�W�Z^�xk�#>D����_��a�0�V\�X�o1D��r"�)*��	���F�,T.ES�c5D�(��U�N��A�n�<7  %!�	5D�Ĩ뙏 U���9p`�9�D5D����ļi<](c���R\JC1���	�0daC�.XLU�$A�\�$���� 1�s���7����$Z$���IZ��(FH�8Bǟ�U|��fD�J�\��JQ�gD�f��䅁�f�)�ȓN�ș�� H�PB,c�b(Q ���M�&|3P��(U�|M(t�F�O���ȓ|�xYBA��jS�'/��?�	�� ��]��!J1g��;`�����P��x$�����7p�X� ��v�4�ȓD�����Ҹ��5#^�PE����o�e(�dM�.�l��%��!@����ȓ&E4�ć��B9j @�	�ȓs��$�ׁ�.���Ig��I~��0f(��7OLîUS�a��8��ȓZ<��ɖ6/��B���^�|ɇ�O��6�#!/Ρ�$�X#z�N�ȓU�����K�@��PV��5�ȓt�D�hGN�,������
y����pNI[��P
����C	���ȓ@�f�����L���Bڰ�ȓcC�X(T�
Z��pTh�8�.��ȓ	��`������=)�9�"y��z.ݸD
����@���A���	=���ĩF�O�2����<&6�ȓs�*��Λ;NJ���� BF���ȓT����$��O���f�S�W��ȇ�1;\	ZR .�$����+r���ȓ/�j�j�グ8� ��U��~��$��0�tl���-� h��I��xd��!{:�	6-�C�\0��I��C�L�ȓR$@�U��%m�fl��'�A@8���r�ز�ʆ}��Y��A7!����S�? j CT9L=����|c�h�1"O��Pg㉡@�wH�&=Z�H(D�x�Ӆ�)$�$qp�Ϯ�#��;D�(Ĥ� �A0��Zq<�A��6D��z�-�4D(U�qǜF��h�Q/D����k�>9��`wM^=QS���@�,找V\�����)o���`�؉q��c�@`�L��.�'���'��Q�b(D�l����Ld�i3ÚI!�*�$D�t�0�זU�Ƹ)ËL���1�g#D��j��4���T��3A�-��� D����`�+Q�$�qٮv��uG?D�,�sdW~ ��v�ٕe���S;D�\re��+pޠ�q'�!y��5a�;D�,���͈9�r]�dg*.r��6�/D���D ���-�����v�"�'+D�\���a~aSVA�#f^Zٻ�a/D�t�te�=F{|��`D�[���"/D��iw�	�tq��>P�Q�J/D��`���'rn.��$�ā\��(7D�����m���M���B'L7D���t�J<,���%^��ԋ�D>D����a��hߞ�yu�9n�2��+D�D����	�>�Y�g-�taE�)D�L�'��G�s�EZC��l��#%D�l�w��=F�d��f[�lڢx(B$D����,¥����&(��{3Z�˶�.D�d�q���z��DJf�Ȩ�:i��(-D� �G��@�����Ia>-ӵM*D���Q�Q��`}��j[�R%�H{��>D����~����غ��lÒ�#D�H��
��S�н���> �j����#D����aM$�F��L��
�id�#D���f�\�
�D<��ˉ|=8<0�i+D����g]�_�f��2"yd�vo&D��+ �,c^Xu�#�͘>&�Г�2�ɟ�X��?%?e�w)H�H��$O�0T�R�0D��if�ΕmD`ɢfM->0�:���d�qOl	B%�3?��B��ҝ�Ӂ�R]��[焚T�<�"�W�l�\aI��I%Sƚ Z���+l9���5�O���ug��+ƪ�V��15��D��'�qSs�[�D��/h�Lxv���uΠV�Ռ=�!�$�$_�Z��%��b�eCQ)�)`�1O�y�i �ḧ�O~ ��C�'t}�Y�ud͏F��B
�'|��GC**1 N�6��]��a�zܓK�QD��O ����4<&eO�4J��9W"O��N�*�)�d��?x��.
�b��I Kfd08�A�F�X���KF�����.rh�.�eP���2��$@�c�%�!�ȓ�<MxG��V��]�Ңϊ � �Dx2�ځ:�qF�Ώ/]�%! +�=O��� �)�y©�	�j`*�C>9 �0�W�
�4p�pI�f�S��y���X�Q���:z��ɔ����y�����SƧۗ�t%�ㄞ��y���bw�m���-u�|���*� �b�Y�����^�.�`�'�2��oV�2|��5�w��}q�'Y�Y1p�˼d��p�!EH5dh �H��DM�μl����ʨ#���z�J�-$��UA��!�$�?1rb�� Ί�O��J�.�<5���cG�J�S��?�� /��h+$������Fl�w�<1�@�QqBtʢ�޾[��(c��K�<�dm�kw���Kڿ\x�:�g�B�<�De�<��A1F�H;1J@͢��Gx�<QG�� NrK��f� d��|�<�V∋q��P5K�48��	�x�<� �X{g�ԱB�M�`)��<Ȣ�s"O��7���BLl�r�W�=�����"O��ɢM�+4�2�@&�x� Xq�"Ob�"���i�$�+dEs��H�"Ot	�Ѻ	�|P�㗖(���3U"O�)
�՚\�" �QD �J�$����ݥA���&m1�'P�d�d+�(ҢJ�G���ȓ�J���
1�nt��lC�>!�c�	��b"z�'|F9��x"H����jr��'^b�|���74�LA��T���1Q B@?g`��9G���D	�Q��% ���I.u�\E����
��t�6I
�%���D��	��\��	�&��	�W��ڷ$��a�H �-	���B�	�@D���1K�(5�qْ��a7��O�e�2(�g;��1d+���5�l8�' 2�Q{��N f-(�q��� ��[_r�$���bt��4���5�HEP��'�^$�F0����X�Oi�]���ș(Ҹ�(v [�>1�͹GL 4�q&�1���d�U�7�� ـK�e��!C�M�DP]��Z0�A,��P��P�'��Z���d��S��� ug��Y���h*�8�E,{��(��#m��B䉃�Ryb���ejR٢��d�OPъ�фg� Pp5��P
0!�"�Lu�0}1Ǝ�v!򤅤h�J9��@��Q����V�7kP\��(3��I�k�"|�' �r�NY�@�q�?] Ľj	�'Rx](-�
����3*�+O�ء!��D,��J)�I��F(�����
�:����=-K"��2'�U�!��3fx��Ш�AU�iI剘��9���	d��p=Y׉�1Q����jE�<ce�5��E؞� ���.��a��Γ�mh�/�79N5�a ��.9r��h<a�x4Jٰ�I���8�"�Pئ��B��i}2IL.v�IA��x3Hՠ�)̏7�e�AT�;�<���B�4EF�z�I�-`��'�����!���6��I��R�P�A+9�a�����$��(���7)�I��Z\Ҳ/ްjw$�d��78a��  U@�ʄ#<L�P��Kx�$�AP���<�lx�'�� ��IN�"!�tFA!4�D�b'B�D�Y��2�	���ӡ5�N�Z�bC	�E��R�ט �Ad�K��D�C>7'v%@P
O��s��ۡ ��p�T�ț[�s����TB�520�'䊰��
Q�C�����[� ��|�D�D:.��\j�N�g�ʬ����7��z�b:1�.��'B�)Q��Nfz�!a��	O�mz���(�Ć�8И������O�� ":�bH�3�u6)Ҏ	��)��}�B*f�>+� 5�I~*2���$O,��2�ֲvY*��b��9�FEk�$B*�rG%-^t��sN4O|1�3*��p���� �����uZ��[en�����O0*��|�$r�#�2V�V�2���� �7N^��c"2z�P�?�O���gϟ�h��Q0���;*��tYT�V�z������� xܼ��.�B|p�ڗ�.m��M ��)��lqt�v>}��������g�$k�`��7,O��ɏ?bK�8��^�Y�Z�%G�yT�m���E&��uGגeUn ��E�G(�SDےX}d5ƥ�b����mJ�	>5[r�A�ԑY%r��7%�.5���d6�L�u�W�T|�z��ٿ6]x��IUZ v�'e��D��㛵#��됅N�X�V 0d(5�q�M�R���%j�@E`�:H<a�	���9�p��d�D�`�|�4��O�xУ�.H�\�X�,�N���Q��?���Eg�h�d!H�u�A�6���!�ȇ-<��Z�R�@�"�����A�6�B��,�|3�Q�#��! ׏N`{�a�!L-3&�[윀s��@Y�Ǚ�`���#û!��'��gp�IkV�ͯ|6"�s�j֥������cW�0۶�cZ�|��O |h�f#�-~�m!�ڞGFl��v�H�"Z���r�+*�A��E�r#f	᥯��$�:TX�Sf�T��O���&�9�n�����AS`�ka�`BG�s�ֱ��b^�6j ¢�MI�0Ez�$�9/�	[��`��)��vk\���$EY��K��I�sz�u{A%ŭYLT$�� Y=f���#�'w�g����g�<�v(3�"�k��X�Z�HĉJ��n+�bs,Ӹtx���+ĝ<��ͧ3�*�C�'�F��[/@���7�	U��@�ӥ�
'�,p*#嘅27�c�@!&�LM�S�TU,[ʄű��A�c�9�g��\فլ�>��k���|Ӣ�ˡ�U�YΌ��SI`�>�[���5q?�'^T 9����UzhV�_�yȢ�'�p��c�3����Mh�1Fq��4
���F��e��kT�Q�<�0��hn�>�O��awC�_2�� ��ͼb�j�+�|��M�c�f�d��w�Q>�I��";`�92ER�^[>pq ��{�LArC!Qa~��(PK���Տ��_"��s�g�*��~���D��{���"`�\~2F�<D����נD1V��P@ʹ�y�H��1A"�Ϳ\K|�s�bM��?�p��% ���D�;Q'� :K���~� f��P�Qd8�}�iޯh\`�t"O�<)q��@�
�j3'�c`�	�2�L������C�%+�3��՚sY��i����	w&���EƏ4qOL@��ǈ���Ԕ��Ԗx�|�i�+?�丫QMU�&gDq�gk��0?q��ܡ0o4�Je	�.tVT���V��K>��iq���T�IU|����>�����5*��;�ɜ(3G8����\hh<��l�q:�g��Ϭâ�տKʼ�!�A�?rdb�CЌ�0-X\��>�Q�ϵ�l
�C[i���E3<Oh:5�l�� �O,I{A*C*̦%Q�͖�ER*I�"O�Y�5�і&�͋u+N�n���[7�|R���k���G*E�Oz�ň�d��j޴�����~��B�'�b���
�rѳ7ؾl��eqF��/O:��'�a�"��>!É	v0���)��V�pâDJh<�%�Ҹ��`�hL��%��?|dxr�	(��o�|� 0�2O �!!�A2��'����ТT:B����X�X�P��	ϓU>N��w�Y�[�T6M]^� �iр�f�4 �����P����:7������r4�7LO���C)K
\!�f����*�|�&���@�
�Z8p��� n"��qI�+���CVV��Yd�ګ/_�)Ja�� >fC㉠�nT���Q�x��t��гBb ��5*u�^�K�hRV�B����Ѣ����!	�<[d���Z@}�R�G6�!�$��|��:��,l2���CS�wJ8���߮4����VA�\3,�)�$ӫ}��*��O0�O�H�b�A{�v(�7����|�9��'��T��@d��@J���V��ؔ�|��ώ�uܴP U�N����<˥,U�MеC���Frџp8�l��Re"h�N>,��I"���AGl�bʟ�R`�h����&��	�'���3���JJQz� 6����*O.uũ�Q�h���K(&��<�U
�F�'h{�AYW�ȗ: �%�P�C��D��
^�z�DD����H�
j:*���E� 4B<�!���O�����c�[�)9��'&|�B E]	W�V���
���
���2bG�^�� ��A�h�|��MF�~���(��J3;,�VȆ��t��',�2W��=�f}X��,!�:d���d��J�����F�:�lZ, �6x��b� rn�HrG_��D99�"���O�@����m!��0gΑG9p���i<V��mE��)��'��Pё
�l ��k��)vj���E�G/i��h"�e��`!�$��9@�=�G�M�H��*࣐�A�^3�̀�4Iݣ9 1ԧu�o1�qOn7gY�n@��RKQ�	?z�k�O"�Ox��g`�\��1��ĉZ�<��"�@0tt�:,�oN!�D�,"�>�R��T�$��v*�\����2խ�dR��j/��~��g�L n�DC��.��C�I���� D3:{�-!��n���@.>T�3����)�'O�X"�
�G>��f�0�v9�
�'#��I�b{B�� �N+R��*O��!զB87j�@˓q��!�Y7������
���	�}�� ���P�z�Lc��/d��Ya���P�Ɠ<��2�A�+E܂��AP� �E}ң�-2PE���Q<7�
���Y�R��!�7)���y".�=#�向���UP�y�ƀW-�yr��e���ر�N�8����ǡ["�yb�1]+FY�m�=�P�P�%�y���#���e���6P�w'ߓ�yb����a��-��'Fm`�nG�yb�ɤ�.�#����m�J�۶�1�y"�I]���R`�(MX����M��yҧhVh����<E=>uqP���y� }a�	��@R��`�ę�yҥă9@��A/»JXi��"׸�y"/�@6�cǌ�?P�X(7*2�y�l�"�Ys�S~T����Ɓ��y��Wڲ]k0�[�t�����ɨ�y�ޞljm+�
_�u9mh��*�y�oڒ�d�R� ^�>#������y"g�"M�nx
vE g�Mx��9�yr���X-b7��o�T�Ң���y�oBVLū��9I�1 )�y
� ���H���!//W�r�"O�����y����&(�	LFIZ1"O��'�-���͑3mJn0�Q"O�%�ꑐ4�>[�[�#�D�6"O���%`��k��u�Z�8��٘t"O
�)��>T*�EC�%�ά "Ozq� ��.wNY��͒.?���"Oz��5*���{GkR"x+�]9�"O����)�"�� �A.'�,Q�"OB��HU�E4�J�'�#I��"O��r�*�m�'�"���"O���t�ڲ$A�j����pT"O$��Y'b�6���׏t^Ĺ�"O�Ƭ��T��#��@��ۧ"O�yy�A�� � ʒ�9I<y�"OH���&�dt
	Pd�͟g[>%�"O�ȥ���mf�!F�@Gd�d"O��`u�Q�0' ���O�@�"O.�׈L21�*�	����Xq+P"O�5�$��9(�����o)� x�"Oj��a ��@�`��1����"Oz��0��h�RM*`K�NA�"O(�襤��	\�ЊF홗)�Ĉ��"Ob�"p'��4x�g+Є� s�"O���S��$Ir�U�2���C`"OD��O>Vv!r�Voj0�3"O.�PbM�JD��M��M �H"O�Y1��1�$��˄�H(�f"O�-��oF�/RH%Y%�d.����"O �؃P�~�f�he(u0.�)�"O8�;%o�0���J+Y)B�)&"O.��cꙵ ��- #Û�<,�4�Q"Oh����z��Tza�_D=^��&"O���施9�NXxWMM(m-©P"OJ�c���t����T-�5P��[$"Op�Cq,ފlw�X�T�.s�06"OM��S=$�|��_	ʥP�"O�:��_5af,���Gc�~8K#"O��@w��/{P��F��>T�M�Q"O8��b�@%>�D�hǂ�:l���"O*�)�jU�Q/"y�ׂ@�7s� �"O��q�[1F����ψ�N% �"OĴ��ȷi���eoʹM����"O�Y(" K���Y{D,�.8����C"O�t�6σ�S ٫�f��~��"OV�R2�G�\�����%��^IJ�
s"O�9��D�zyd(c���95$�Z�"O�e��
�>�j�޵b���"O��Ѭ���@�c
�F���c�"O:q�'΃�'Wd�(��u�,��"O6��T��%(P&�@7ƃ/(�2(��"ON)��OU`���ֻf�����"O�����>����"O䩀I_�N`QZ��޶+���H@"O���jf(�jE+�frD@S"O*���n�] �+t+D�H�"OY�j>
�@9h1C�>U2h@�"O-a���A���R� �?^���6"OL�b���!j��m�8K�@(�"Ob|(U���D��8�l�EO8�)"O�٨E���CV�P�k;a(Ղ�"ORmqҏ:���B��Z%>�i"O�1[�S�(�9
 ��8�^���"OxuC6+O �$���G�`2 "O� ��;F�dY4h�b*Ώ~�$��"O�4rG�
RF�I�[�Ws���p"O�i���0w��!�$Lakd,a�"O�l���T?PK�պ4��;sS�](�"OZ�C�HR�v>� RA�N�[�l`"Onh87��K�pm�6HXZ3d��"O��׃T3�� �琝t'4Ht"O.D� AԕQ1^ūpF��}���`"O���KݱK}.D�#O76�r�"OL} N�&�N5�d(�*�����LH�C�#�Sdd ��:@@��qSiP�yͦ��ȓw9X��g�<p�v���'Y j��R�#ř{D�'��1��P�b��jJ|S�,�9�x1�&4�h�U�*c�a�Q,^�5N<�Q$0T\�BF�'�桇�#_;����D�����BOy�V��DD����[CNz�R�I�/u&�3ǟ�
B��"�8�BC䉛R��-`�Ѥ�4��v`\p�8�O0����]v� �=�R�n,`6h�/Қ)�Q`-a��Յ�a֢ R�`�?w���2����i��#`
�P�'h���>�5�¶��Hhr Tk�9���gh<��*ܛ6㎙�©�|�L��^>*�̕	�n�:(�����kj8�2M�.'�0�S�&Ͻ&����I.%� �ffN�"����D �AJ�f�s.%� �FRQ�ȓ9k�Ձq.��L`�p��i��M��p%�t���N��l���]�O�@��A���ԩ�!���4 	�'V� T��(&{�����<��0�O�B���O�q:��3?�BB�kB�ԉ%͗; ��HX���H�<��*�!�JA�7���S�8 �j�i��"�Ba}�+�C��4��A�U���'�� �y�L�0c��!w�
�Oq��"��J��y�)�gƪ� W%�Vf=Rq�M��y��݂pf�yrkߧE��S�D��y�'�=����H�P�1b�X $X���ȓ(��ai���5KT
u)񅛵LkP���v�h=P�NN�H{9!�&�3H�V��ȓ��E�AiY,H�t��b��*Ʉ�:���aa�UwJf�`t�( '���|�����̑X�Ă�
�)��\�ȓk(�(t$
9Z�.T�m֍WbP��ȓv��l ��x�:�Ȁ�U�q�`͇ȓ��Q;ᨕ�_BX�v)��HM�ȓrf\	y4�Y�����<��`�ȓ&��jq���N�K��?h�G2�E��Z�&�`�+B�B$���ְ�� ��d&|�1O,D��GG�;:.dAU�.SE2q�%P���1�K+`,r��Ov��CV�R��6���*�Y^d���E�8�;O^��d_�T6�,Dm)nf��A¥D�J���AEcɲC���v�&^H�%�Y�#j[`j��/�x�`Hʉ��q��	��Dqڼ��ɔ���d��	��I��J)�T�%�.�.��nڌ�Px�P�H���d��j;V@a�C���O괉fg�������>�k&�>�ūی/z6�3���5��d���^���'p�l�#��S{���K�k�jP��`Q����G(�Oꖂt��a�4�Z*(�,�5쟽}�uwO�L����Bi�[������u��I��Jۨ+�,	�-O�M�M_��2��ʐ1~A၍6�Y�ƀ�9Hp	�ǌ[��q��±/�(���Ŗs�t���4�2��Z��Q����yb�@� \�`8�*Үn7Ĵa��3U�� �d1O��(s-:T�|Y�]Fځڄ� �Ȭ"��>��hbR��Gt )O��#�ȗzX�q��d��G/�8H��ϸvh��@�*J��p ��xGK/R���WŕN��1w�|Җg]"�h9�% �I&���@4'�~h��k�_����\�Tt�H�\��4B�b�;��)�E�5�|��ejO�/�i��:�V|3��7��}�琧y+��S�$U��*C�Ɉ?Urc7M�q?H��/	5���s��G�uԀ�p7#�y���x�(�9v��j��m3�Fѕ��I��W�T!��>7(�K`� �$aT���	pydD p?䌋2;�� Ix��3��P%mg�#�d �1���L�<R'�HQiq��'�2�*^�y�Mr����n�T��K>y��>l�Z����Z��(��	
� ~%Xb�ܧU0��k��t�\���V�#�ar��'�Z9SA�B$8�,ŭ�+�x��b
ղ�,@&����O(��0�+kºU�'��uѴ���x�VI���B�.��<��'��=��Ĕ}4�bC�r90��8NHqp�'��5��������F�GL6�#^U�+����T��Q"O5�׊;��,8у�/�vD{U'т{��Z��V�/�3�d	�L�d`�IX�!�E�󁕢PXqO ���
Ѩ����l���� ��yb�%W�lR����
IV9`���0?i'k��NY���Iv6�� ��t��1H>� %�S�d��)�^\���>)6���!���ʿz�R��w	�Ah<y��A�o|�FH�w� �ٳ�_;{��!�&�0sm��p�K<I���>�HP,ą��ЈB�c��0fH<<O����Xf�� �O��8vl�0K3��a�@�!(+d��"O�Ec���
h|LEa�\p��w�|b�LYh���t�O`^��4�Q�v����A�R�~:PS�'���ęb�`�Eh�7y��}X6
M#BK��'�(�p��>���W?J;L��7m�Q���+"DErh<��L
�b�lT���T�I�4���J��Ȫ�I�G'�N�l�&^�\� 1O���D#W���'�z-x��a�`q���:��8q�`�lQ�w�9��6-د�
,	g���f��q$2,��I9���rt~6�Q,|<��a��1LO��(!n��9��D!��[�x� �|�D�X�v��p���2��Ӫ�AJT]�u,	e�� .�4s���Č
z�"�D�fS`B�ɧm�,�c��#+�rq�Cʇ�kri�6�b���K���,kzD�0m�K�vq�!G�}�����yG(^t��ŀV�H��-��y�낳 ��  ��N�Vt�Cb� �(83"n�1�h�٤�ŕ8(�90���!��(�'O��'��T(ƂM< r��fg�"7�|\����|H���/[O~�;�Ě�ilZ��j@o"Պ��91I�Y���*��y2��/(�0���U�Z��!� \���O�T��
�QSdm2w$�uq��耫�g�F$��$�*=���T��\-�Յ�U��&�7v���J2�^��~)�'��%��kH���m���:h��!˒�=��SB���P7<CF�ir�S?�B�ɩ[/L�1�I��DQb���*ݎ���b�V���9���t��<��M(��`(��!!��p���8ڸMR�㇗a������0LAz!��N����C�ܴ3.�f�[>G�D�Ä�،?�U[���>e ���	�/{����j"N�h&K֣�<�=��@K�82�t��M�KQvd�CGA�'��!��'j�F\��k[>B�!/����A��-��,k`�R����[(|�Q�"ϳ�~⅐��@��0��D�.����9pU�d���F�2C�	���%4F�U�p ��aPSG��	2Aa�1yU��JA �O���I+�'w�x���5wPh�S�(�8��	�)�6�с��h�9tl�'S��J$OL������ $�� ȇF⊄/�qq�B;Fjў�1t�@�	��	!'�I�{9��U	�X�²@�S!�$�1m����`��p�d�TN�(D�
��9
� Hg�@��+x49�&C�A�xl��4��0���2l{wL �|.Ba#�ϑx]ą�'=��8�m\>D+�q��I�I�P�B�R r�r�r���d1���Ѳ��Y�ʂ`�H�V�Ž[�
qz�j@,w.B�ɿZ��%z�oWF�^E;�L�$O̢>���ܢF�t#|e��:bv�Z$�F *�V	�4"[�<��93�����M!
h~h�k�R�<���S�JslՓ���" ��pJN�<Ѷ鑷�����F�
�4�(c�
J�<�"�޴��J��.sȠ�`D�l�<q�I�y�VI�ɩZ��!X��k�<y�Ȋ^ԍg�9�Z|����z�<!H�>i�:Z���?��1
Z�<ɀ�Ӵo<�� �)ԲI2_Q�<�e�Ƽ3O��(#� �Δ�i
�M�<���x|B �"a��%��!)���B�<��cχ6 �#��x?^���N|�<YC�#ɰ�Ao�8r�>��	~�<��R%^���*��ɴHT�X�m�~�<Q���-߲��Q�˳#�8, skb�<� X"E��`�D;`��O�v���"O��`V$dIs0
f�p�'"O����)�����_�o��A�"O��KjƸ0���ƀ6�P��"OԬv��{��xքo���JԞ�yBF�2�V�'k��`�� ����y�C��K�V�8��.U�N�� �Z��y��;^! 	1�B�N�� ��*�y2� P�:)����B	���w@ӝ�y����1�b���
��1�\s�!��y"��~iֆއ+��qg9�y��H)8�<���$��5Yea�?�y�F�;g�����o���h5�C��yb��7@Ĉ��@�70*�4��/�'?4(���m	0@{�l3.���ybk�A��b�i�'w�,����yB��b�`"���Y�M�#�Ê�y2�$�\{V*:� 9Y����y�P�o�e�K�]gV}9E��0�y�)^�`<jAb(тM��T��G��y���b|1��R�=�:�!PC?�y"	^c�(��e!��8#&u���V��y��KbP�f���D����^��y	\�,�r����Q'�tH�����y�8N@��0��:g�@Ɗ��ăP��(����f#R�R�&A#BC��ru�)o7 Q!U��[�	X�m�#r���Z�'��n�Ve���0}��k�F���S3ae���tT�-���ξi�"�'� S�gW}�A���gUbh���%\� 8�ጘX�R�>�.应 ��fɧ(���3��ִ{��9ʴ��<\�,�`�'�nI��#L�ɧ��x��P
�&��8KWk_��a�HūƤ�[���b�.�����֡�:_���H>D���7HشC�~��I� Ov���h<D�|�.�8�qAw+A,x��`�.D�HK!�B}�M�&�"H��Pd:D����`۾G��*�=U���##!8T�H�I9��rM�~@�DK3"O��:P�U?muh��skD�+NM)&�i���iQvG�8*�,J(�R!�a
�j!�D�2NS�iHB�.(������.F�!�dT�-���)��P���Dt 1 �'Y��AH\�z�6qkc-��65��i�'���� ���X`����ލ-c�@��'�4 ��=Tj\��oD�!�̜0�'�h��+�4j��c�!S�W��'��Eۆ��>)�� &T�e�LK	�'$���b�.�y���4�DEj�'���c��?#�ް����F��Z�'�`�# �<"��Q #]�p�����'z�����Utt	�Bp�Z��
�'�u:b%��?�j P��ٝZ����'v(�#�4e���V��L� Q��'�*��8���5)C*B P=C�'xLe)ǎ'4E�4����NHAa�'�<<��a�)T�x9`��-M�By#�'Vy8E�ܖP�@�S&�J�K���	�'G���c�kH<*�F�oS���	�'t2���Ս��iBƈx�B%��'ݨ�J��D>H���k�����'�
�[pM�-X���aJ�_3����'�0���"3
&�0,G� C���'��=�'�'i��W�	�Y�1Z	�'J4C��ɸ5|�L�7�óy����'E>���|c�(QV�8!��k�'�v��%���C��Ԋ��^�{t0���� �0Sfd����a�jX^S�I�"O�А�M�A�b��a�<4��e"O�a��GMs�l4�4�D�8���"OVi�d�4N���؅'�z��dI�"O�H����(�4����+�t4:3"OL���Ȳo�`��T%2>�L��"O,�*�b>Z9"��ř�٦!!�"O`���� ���d*�t IS"O��)��*H[V�����-�9R"O8�b�gӧ~��X�g��v�%;�"O\�C�L�3b��teΎF
�A�"O6�c�ՒF^$T:���J<"b"Op=A1쎒%���{���H����E"O�}s`�ˑHP-�#�f�:q�A"O8�(�֑+�d��vg�(��u"O����F�R`E�F�Q�m��Y"O(9�ލA�>}sq�3�\("6"O0�� ۸W㦙:`$�!w���s"OQh"�y����J�"O�X��H�z2�h�C��rN6a��"O֐���M	1����,����"Or!�v��JF��K��!����w"O�M`g��P���_iƭk�"O&9��D��m)c��fV� �"O���9L������'>%��Ñ"Oj|9q �?j�TZ���_ <�`"ON}AtG�bhq�7��i�"OČ�ƥā]��CE��xl�0�G"O&�z Oȍd�ڭz��۾O��y�"O`Hh�5nfblzÆ������!"O4��rON�W���� Kc����"O�p�Q9�DY�B�$-�8a�"O���O�:p�T������z5"O�����R����S#D#"҅r�"O�t1��\>a<�Ƀa_6� ��c"O��ÇZ6>�pP�ے!��d �"O�|�B���6���h��&�r���"Ot �S��Pvh���@���6�[�"O�CU�X�p�9�`��<�H4�3"O2l="��#��R)x
R��c��'�yR'��Z�(��CK[i.�1f�-�y�o�O�RD�� d�LJ��C��y��ߺKѢyj�AL4EFq���1�y"O�<���J�g���`�*��yr��0s��f�W�	Q�,��J��yjU6Nn3p �{���R�(0�Py�|��u����4(�6EP��j�<�FB�b�>��C��B'�t�҉�Z�<����P⚽���ݭ��); �Jm�<�fdح(A�4a�*
�5���XM�<"�E"�%φ�Z6�� ��BL�<y�(�� jb����6(\�HBI�N�<�K��8!�D
�J�.}���z�I�<Q�� V�i���#O�8) ��Y�<��E�i�
�.Ü1_�}�G�<9���!(U���T�<΂���|�<��m�*�:��q葻{q��c��]R�<� .�-��u�I7�mS���s�<Ƀ>=�ɨB�0b�ܘ�"�t�<�/�tw�\�4�.E���*�"E�<aAҔH@�!E��!]A�iR��D�<�� ��ő�"�6/����r��x�<���9U�؉��i�?9���m�]�<����{���P��g*�E���D[�<� :��wA� 2��R�F9J�� "O�a���'(&8 +��>װ)p�"Oa�3���ga��&���(�� �'"O %�%��r� T*vd�5|�j �"O��!�(!(0�p��S�t��{"O�=��CB%�	��Ndb�l�v"OB�Y�$�{�p| ��CW��Ʉ"O�5�v菈$P\��&�T�F2\ �"O&��:w�E����2A��o,D�hPSȃ�cvРc'|�r� D�ܢ�Oo��}�4h�7"���#�>D��h���"*�pȣ��
#,�iX&�<D��S�b�*��!y�g�- ��ɶ�<D��A@ЪS��y#A��!�E��L D�����Ϋ���U�rɺU
2D�4���xતy��f�8�QB""D�d�3E�Z^���!`W�Ip  �?D�ġ�l���d�6�±=��Д�7D��A�M��G,:a󆀖T.����:D��h�+ňV;�Ԁ'i�2\��X���9D��P���
E��8�����c�
:D���M��H��,�#�*�(´�%D�,pa�_V:� e�#h骐��#D�(����QI̞,}�81aԮ#D���'どSyp݂g���xB�!���!D�H�!��#��r�F�=��A1��?D�DyХ̷IU�I���{�
�p�,+D��o	��r�����'
g�H� M>D�xz#�~�e1Ң�5Hа�V<D���FN��S�!�6�|:�L$D�X%)_$C�(�CE�x��b!D���U�Ƽ|�\K�D�Ò%Yp�;D����@�I��c�T3Y���'.;D�(
FF�L�+3%^,�`��:D�sAf�
�8I��hϭtS4y�k>D��#�WtI Q����2��DH2D��A�D��I��18��@))��K:D�p`� ҙ,7��Ӧ	]84l�����;D��I���-����f��*G� Q��9D��C����R�Ύe��P���$D�p�sO�j\�9�dM�\2�i�� D�Ġ'�s�ƽ��'J[9���	<D��ŉH�5��U�G��6 ��Ym9D� s&fF�H��D�	�$"��Y`�7D�8�'�u�T��3d�3�T����'D�L8��x�	�JI�DTD98b�&D�Բ�n_�m������ž@yh�$#D��
C��:(n�i�Ў�Y�z�%D������J��h��?d"i @�!D���O�+��d�dBG�"9H�z�;D��1��P�c��U�E=%<�1�9D�����E�+��X&��L:D�pX�n����a���9���q�*D�,��A�0����Ԯm���#)D�y���
6���H�w�`4��O%D��* �N���Ҥ-|�6��ҥ!D�h�1��?��H1��
�N�$�8u3D�T��̒NzƸQ_�$�T4W��C�I=[�x-5�։j"�=z���p"O�8R�ͼ
J��L7(��"Op�*�F	T��u��悖$:��"�"O�;�E�N4ά��/�O�F�G"O�!�#�V�&9vL����&m�hb�"O`��@&E=*Q҂c�b���Z&"O� \%�c��*"�%�a4>�@e+�"O�I���p����p�jL�g"O�0��._�;���礐�$.�y�"O��7˘J�m�D��J6��""O�L�h΁���7�7?|�"�"O�b&�wP����� 8�DY�"OV<Ɇ�\5`����P���r1"O��THݵj����Ј3�N��"O^-;�G�&�<��û&��!��"Oac�oG�J���&�
|�:�k�"O�mÁNY)Q �H�\ 3�2e�"OP%ipg
q���2$ڕW��=A"O�@A���8Ed	VC�f�}J�"O�AQp���#�СT%qH<S�"OrS�T��6����TZb	;�"O����֙_���y��1I����"O�|��5�6�h&	�,3�a)P"O�(r�@As��`��Q)�Y��"OJ��BdZ�7Z�L��o��>��0�"O�l�%�:t��9���ƀ`�f�#"O���ƣԍB�0��Եa�:��v"Ot,@w�O�L�$I	��
$�dL�@"O�zԫK�[f�����B�_�~��"O����i9L��0z&��,���Kq"OP}�+	�` ]`�O�&H�t��"O4)ɱ�֓*^�	����j+>�au"O�x�ՎTBT�s4�޺o8`q"O���Β�d�����#48"�z"OT#b]1L�^�����/d2@���"O�!�!� ���k��QRn�B�"Or�
�Nʖ>���o�&�Q�"O�%B�!S@��A��a)+�a �"O�� ��9��l���T�OR-��"O�%!�!��T�*幕���oZ��SS"O�Pᦩ�|"Hi�A�.�`D�W"O��q3�V����U���r�=�5"O��RN�m������'mEP�S�"O��`�W�S�A���R,�吳"O$���G0.�n� 1f�4v���"O�i�wE�>��b;<����V"O��;��ˊt��W�#~b�:w"O�2�(T�s�P s�E�5z:Ĺ6"O�� ®�L|�,WG��Փ�"O���G   ��     �  B  �  m*  �5  yA  	M  �X  ~d  7n  �w  ��  ͋  g�  ��  �  o�  ��  ��  b�  ��  '�  ��  ��  '�  k�  ��   �  B�  ��    �
 � � �" �* z1 (: B J OP �V oZ  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p���hO�>U2��F1C4ӡ%B�>��eW�%D�����9]����"8�
mS�#D�th���*��6��4��$#D�\��2~F��u
�!.���sA D����ýe������[�<�����?D�@�w%��&�f�SS%D��8a!�(D�HY&N�1V�ȥ���V&D�A�`!�	�#��yr�C>s|D劥o^2;#y�Qk��Px�K�{�T�:���(8��+�#$����>iS�'lO�m���KTѐsF�W�ճ��'�铤�$ũN���rć:5�@3"��)rm!�P-s�h3eH�r�xb⪙�j�!�䈾�Bl�*ݎzp��a2c�1Y�!��8$�N9�%�D#f?��
�#��y�!�$R*l���2�Ɵ�1���8cǈV!���+ D�
�dV�e"⼐Fip!�$�8p�,�7�֐:$��`H�;�!��vM��­�@�0��/Et!�ĚYゼY@!҃&���K�f��l�!�� ,.�T�%rd$�4�]<~!�䛱���kah�f\삑�M<+`!���8�e��2G,%s�FS�gI!�� ~��d�)b4��ci��.�2�"O�a�L�I��=@Dg�0��TP"O�1���F�nؘA�5^�
���*O��(�NB4)�xt�θNy�:	��Ms�O�ݒ��hҊ�Q Ў!�ZM�"O�������@K�ux6Q���{�O˦�l�+E�x�Q�đ2 Na�	�'٬D9e��91��p�X$>��a��'�б�Q����i�&D ;? $��'͢\"�b�^�@!`�A70uش�~"�Pc8�@SD�?(31���T�j	���?\OB���$�`s8�Xt�����I�f�!�D_�)��#��R8�$=[���F��'Mў�>]@EÜ� ��9z#Ï1�̐ .?D�X�h�%;��hK�ɚk���F D�*$J�)" � I�3*�q'�9D�L��l�K�d<�7�1<�5xү3D��q3O��%pafӀ)R��p�/D���f��J������Ib"���-D�L� R.أ#�	�D�*u�7@+D��8R&R�2���B*^,�Tk�k5D���3
L0�,��f�1(��xC��t��=E�ܴe����Q�0�Z�(�N˖|���ȓ[��}(�h�0"��_�Y �0��j��s&�O @�B�I���@p�P���F~���`F��%�^�7��H�ӳ�y��9P�����:Dql9�F���y��N�'�4[�IE�%ߘ��E�̥�y" h�^�ڇ��5�-�'�yR	 ����P�S?`*y�����ySc8P�{��`���'��y"�U�S$�R�$b��z�K&�y��X�rm��"��\}&�I� +�y�)>1��E���O�H���؟Ǹ'�ў���a"QF�D�A$���;�"O����7��<�2��5c,dts�~����BAH�8�YPg�rhR����y�$�ޘcF�U�n���^��?qQ)=�ONa����ph6��F좱pe"O�e�/���Ukֶc�I��"O���茰+�j|����vp�d4�S��z��X�W {E4�(�&�DhC��2z��iH4�l%��7|�\C�	l��2�利@��MR���z'HC�I�)r�(z���$㠝c��+�FC�	�L��<�����Wl-s�D�$2C�I�]��%��� �X!�BE��ybgH�(�L�g�� �&�Prm����d*�S�O�<��� ({��Ar&�T
#��t`
�'�<M2�g��h5�����	�'�0`!�(��&��`ժ���� 	�'%���7�L�RE�Q$FB��"�'��h�Wl�B��	�qO�+K��ea�'O��Ȱ�H�j"�y��W�>��z���'*fՉ�Q*y������gӄq�'6Ȍa��5��Y2nϤTTh�8��Dp�ޣ}�qb��T�6(��Ob��u.P^�<a!��Vp��ᨕIF��S�GbK$P��O?��B��*h�w�ۿm U�6(Y!�\s����?s��!��$�����>��M�+�����*@�Rm�#�e�<�b�5q�������1�|0'"O4t�2�մer2�/�(i���"O������<4}B���M��!C����2<O� ʅ���^#7
��bQ��];bOx�����&PP�,[��=��( �� $���`8��2����7Z�����>+��;W�=�O��A�'^�}��(�d�X7��<wR�52��HO���&��&X+�c"�r��$I�"OJ��`S�l�1O�
���W<O��=E�t�܉k�Z(ˉX��0Bd	�:�y�: +d��)ɰ\�`�� )T���Cݟ̇���	7G�I�<}���������<IR.��h1����%"�&���n�p�<�u��0Am���4�D�e���yĊ�e�<�W�J�I%�a���
BRV�١AF_�<aTE�TԤ)���=0�U!7�x�F{��逯L`�!#$�˯[�&e��	�"|�B�	j��e��޳�-SET��ɧI��I��~��hO����Ǆ�$L�rs�<8oڅX�'�d��'�4��b�d0Q.Y�f��n�W������m� `�z�nZydN�V��0=A7�%��$o��<Rŕ�,��K�肍M��듚p?���	c����e�E�mhb`а��}X�ԦO�<q��ѷa�pz�X�L���"O<p��C�	R���y�-*g�|B�'��O�c���Tyƚ����Z4�����0D�x#� ��@�:��������d1D��!�[����g��r%p%��/D�� ����7x���ʕ3Y����&-�	��Q��O��좷��'>i�`��o"��	�'
�A4i_�f�\ѓiD�3L�ّ�A,ʓ�h�����t��|f)*>z���t+�m�!�:�1gI�>} e����)�Op��r옺i��h�&ԠXw
"O�p�A/EJ��E&��Wg�-i"O8���R A�	&e��d?N$	0"O��C	qȜ8p�!1`�V"OlUAR �;I����.	�(h��"O6�$�ܻZqd8S4�L(��e�F"Oڥ"`��?bH����t�(5�s"Oй�&ǝ5n$�`vkA�"O2�Q�!�Z�|�o>1���"O� �r�E�1ಸ��͔�/�1�"O`,b�m؜��H�&��8�`��|M��jȞU�ƍ���Ǿ^o�8�ȓRBL�j��@>A>qKv�N�pńȓP�0Z��E�
C�s��!9����ȓ�Tڰ�š<����s�T7R���ȓ-ъ�J0�O,B4^�#�a0|�ڴ�ȓ5� �+�!;ЌS0e��Smf���G�\���
U���dO��&�h%�ȓS�Pe�4DTJ�Ve����*p��m�ȓa@�����[��q��G)�,��ȓSIl��+m{B�ѳ���H
�ԇȓm*�U�#�>;�`p��S�y(�������Q@M��}��-S%ƻ'*Ra�ȓt8����������P�>� ����@�A�A�7#O�S7D��+	���JR᳢G@q`�[��\B��ȓR��;�n�iP��J�:{ņ�?x$I�6	E���L�ES�2.���ȓk�`��3Oĉ�7G�p�4Q�ȓlA���Mլ9�ɳB���$4l��l�*��T B�Rf�P�̇+D�$Ņȓ[z�akFk�7tv��C޲C4|�ȓZ��5��^;d��;A��+��|�ȓ���G��%Lժ���[vhɅ�S�? ,�T��5M�<���"8=�"O���Aٓ8.�ᡧ�7B ���"O�%�X�F�+��B�/�F"O�T� �/f��\u`�89��Q"O��(q��uJ~�	6k��&���0�'�B�'U��'�R�'�b�'���'arP�$@�[��9�,�95����'C��''�'�2�'NB�'���'��lX7F����ȣ��ͷn��H��'+��'���'�R�'���'���'�ik��4+*��'C�|/8DF�'���'���'�r�'���'%��'�t��I��[���LV�+-�?A���?q��?q��?!��?y���?q��ؽ�����K�MX�O'�?Q���?����?����?����?)��?���N���p$̂�s�:��D���?����?����?����?����?q���?�B��*�~�i��Z+Z�Ő�����?9��?A��?����?9���?!���?�S�F�)�d9�C�ab��A�����?����?q��?���?1���?���?�0E��g��A�Q]0,-p̙q�� �?9���?����?A���?��?���?��!3,KHI�4��/M.������4�?9���?	��?���?A��?���?I��=�X���R�;rr�$E���?y���?a���?q��?����?����?	P��)n��LS�ĕ5>F���6)E��?���?9��?A��?���aG�6�'n�x.�3��|��p��@�-8���?�*O1��	��M�#�?q������¦Fr��,/`,4��'�6m0�i>�	��p�v��.E����w��`Ǐ�����-��5$���';��đ>�R�ӂdY��N��Tf̓�?�*Oj�}�0�^.8�����֘{78�R7m̋H��$�'��'�Hnz�5�Т_v�x�ĉe�n����Bӟ��I�<A�O1�����<1.� ��Y���ؑ���<��'^��D��hO���O֡� Aհ_���xZ9��2uʑ�<Y-OX�O.aoZ�,2b�4A�DZָ�b�뜂&S^Bo S��Z �Iݟ����<�O�4c@o��d�lS�_�W�d\ ��	�6�>��P�>�'Tl������dTC���i��
����]
�,i!Z���'��9O��Ђ/�?X�ań�.�Xh�:O��m?Ϛ�3|�V�4�8B�` �j���H aDc��R�9O���Ol���2�6�Ot���J� Ҹ;��I�&˔n!Z�(�B��}�"�OX�S�g̓W�� S�
*��r]
,n(�'h�7͟Z(��D�O��D*�Sxê�q`l�8#�jyxG&�	 �H��ODm���MC0�x��d.Ёx
z�h˕��\�f!P�:�p�B)A�7�剄@��R�u��|BR�T�e�O�m��}K�/D�
jK	�*Da|�a�}V$�O�t���^�l}v�k���9|�Tu�p��O��lZN�u���pnZ�M�It�4���Wt�L](��H9XZ�K>��R�1��^�S�ߙxr�	g�V�"P`#	�0��Oe�����3g^���W�=F��peC�TRj(��ϟp�	�M��AM�dBg�t�O4����՛@2DmJ�+�
'
�:�!#�$�O��4���3�''���4=b�G	�Y�����k�iM�A�"�P#|��IO��Py��d�/Rʦ�:�A��pd	%�� N��,�ܴ9	X,���?�����	T l�
l(#�
$1n����l�62������d�O��� ��?p͚���-Z�͊'+vi[����YP*�ş�����D�i?QI>!g�S\:�\��FU�C"�L�1�?I���?����?�|J.O�5mZ�[��DC.0A�IGA��@$ND_܆�$�Oڍn�F�/��I�M�N9M�ea@AE�S�d�	O�i�Ȅ��%3��œ@X^\0�'w���B�N�2�c��H-HјV��	ܼ����D�Ol���O��$�O��D�|�D(��r#.���̕c���u�ˎT��V�G P�I�t&?5�	�Mϻt3�E�ǋ�^x���Y�1��H"�i��6-�g�)�}���'������ wP ��ֆK���ٙ'L�A��&C?�N>q+O��C���Щl�6�i �O@�̄�I1�MK�d�?����?!Sb�"7��+�蘔)�.��@?��'� ��?)���J<�s��[�x�0�ȇm��)�'6������1C�t�E?���v��ْd�E1=�����������?���?���h�����|��ֆ�+��`�'eŦ]���d��e��۟��	��Mc���4���Y�Zφ�j��� AV��g��q�d�5�4A�����?X�Iퟴ���\�P	��B>9�,�W#T�x���ȓl�)a��O����O��xcaE�7�|K�-�JiP��0&i�n�r�'""�I[�p�P�����l	�@Ґ�'%�6�Ц��I<�|b��<ک:� 1wڄEJ�>,������/{��@��'&�'A�	<��T���*7.����N�f��ݟ��	ϟ�i>��' V7���F2v���C�pc�$F�&h��
E�g2��d_���?A�]���	�0sشp��U�7$��]����Ŋ�Q����d�,��Q0��w�����>��=� 4�y��^�d��Rd�T�{�2�+`4O���ć�K���+�gT 9@C+-�t��O,�DU��)�a�3B��i��'3�Ы��wP`���ܨB�Jt�(�d���� ��|�G�)��Ax�s�l�2T�:��,�z���O:I��ӟ�����O����O�dКk7���T�`i���w�W�\��O˓)��AC"C��'��V>uQ4HC<uhe��bݪ(3 �-?Q7^�����CO>��?M+��Ohf��wb	,k�v�x�eL�b�̓0���"��*��O�.6�D"Zz2��@�},��SC�Z�P���O����O��I�<q0�iC�pbQ�x�U�e	O,-�m�5vR�'.r6�$�I'���b�P���l��=޲C �0o�� F+�ڦ��ݴC��1�(OP��ޚk����	�0{�b7�=����r��O���	hy2�'92�'���'n�U>�Q���%f�8)�N�)*f�œd�ې�?�� ӟ��I���%?�����M�;rߌ�bgd�fL��צBTD#��'u��1���tꖎ{��I�1&��F�΃q����աbgt�� j�� �'X'���'�r�'��l�!�T�4⣣K��Mˆ��O����O�$�<���i ���'���'4.��k�=+h�{���;S�D ��F}��'�"�|r�\/D�*%�qZ�
��DT"0
8��f?�4�H<��'��NײO�a��L	�V�����l�"�'���'t��S�����'�0s 6@�&�6/|Xزg	�ޟ���4hb�����?��i��O�� ]Yܙ���Y<I�2�@ڄW����O�7-�A��ÝF�@���O���խ�.T>��q�)YO��!�Z͟��'C�i>�Iȟ���ϟ8�I23�(B��8~�bM`����Q�ba�'��7m�'z�"���O���<���OD��d��YЄ�tO���D�*Bx}��'B�g2��!j�����e�Z6���n���(�1�J]���	4-[��3��u��|P�P���="���'\�0lni� Hɟ��ɟ �	���pyBKo������O,��W�#Nm�'mD	O
����O~<o�A�F��������ğL��g�&"�ht�S�ը��̚$�*>O��'�bo�<k&��`���� ��/ N9���-%�9��;>����O��d�O*���O
��,��@�R�	�p؄Z aH�#q ��	џ���&�M��C�|*��!z�֙|"A�_������^�&��1
g2@O�o/�M[�����,O �����$��ԭYA��x�v*üZi:��5E�+�?�h'�$�<����?!���?��I͸�	���J'�@����)�?����d����#v@\Ο��ßt�S�?�V��QI��H ��<@��1?�#]�<b�4cܛ64�4���ɒW�v@��	(4��Z2#@�,���V�L�M#���ch�<Y�'"�.����O��C�ǝ@r��[�l�&a�(�ON���O���O1�(�*]���U�l��Pa����v5B�B�:0��f�'��E�X⟤ۭO��oږ�B� 6+_%��U`�gE?:��ts�48ƛV��\$��柌0F��$��dfEoy�Nٜy�Y�s!�nQ��x���&�y�]�@��şp�	���ӟ�OO4T��+�&a��}�f� fy��1'`�,U86L�On���O����D�Ц�*2��(!O.g�j��$C�K\b�)۴{$���9�4���i�����d�<A6f�'BK���� �I� \�0�	�%"l����']$'���'�b�'Զ����Y�]`�T5i�~4V�@�'#B�'�rQ�|��4C����?�����)��/�4*&�I�4����H>y��Z��I�M�i�FO����F�N%�ƨ�8����8O�Q��4Aa���O˓���<�I�q9��rC�¸i��(p�@�,[��\�����ʟP�It��y�&�=Oն�1�ɓ8�,��d��`�h���O�$즥'��s����]�o8��w�J
oT�*vOf����43����{ӆ�y@4���7N�0��'T�}�c��FG�q�"�M5<�TRd�9�d�<q���?y��?����?D�Mo��(�I�t�}�Q	J���$�঱�'ŃLyr�'���^>q��H��IR��K����+"����OXn#�M[��x�O���O��a�g��1�&�[���1;SNöm�RU�<"��L����#���<YAZ�{��piEzH�!)��=�?����?	��?ͧ���ԦA�C����s��I��P��Ô|J`Ѝ��H�޴�?�J>	3Y�H�	֟���15({P���0�����:I��D� y��'�$�[�l�E�+O��I�Ԣ�%P$,��qH��+�(p�78O��$�O��d�O��d�O�?tm]�R��J-+���������ٟ(j�4ydyϧ�?���i��'����S�m܄��h��ƞ|��'���'���X�^�0�'40��b�O&[�n,Hf�&h%�Ɋ'"�-�~�|�\����������� ����?�;Q�/N��ek�����	~yreu���!p%�O����O��'+M�=�c�
��ل{�(9�'����?������|���_���A&�f�@����q\1���4���O���M��D$��S񆁠s?���b�Σy�Ib�A��D�Iԟ��I��b>��'�b6-հyT|H�4��[
�/A�>����SE�<�զ�?a�[���I"0�4��B�6$�
0۾e��t��ȟB��ny�П������?͖�� �J+��R�M�싽;vL�x17O���?A���?Q��?����	A�ߒT�$,�a���JgfW)?^h�nZ'�U�I՟��I@�՟  ����3�"Z5�|�B�(�CJ�?������|���?��&��
�(C��b�Ꭺ&��$y�b&.�d�*��z�'��'x�����I(��h��DU�|c2=0Q���T\ @�Iݟ0�	ȟt�'IN7��D�D�O��$H���0���!��<��� 
�xH�O���O��O���&^�e���[ÇQ�~$�-PĞ��鷃O;�tZ �>ͧw:�����Č�~�JDy��gyt-��?v����O �d�O ��.�'�?�'��:�t��-g�8��2�G0�?Y�i�� h��'_�dhӒ���q�:@P�a��LH��L+�~�	��`��ş�p��D�I�t����O�:�`-���N�[�h�`�ny�O�R�'���'�RJ��y�~�a�Ԧ<0�T��.l�剆�M#����?���?QI~�� @�T �Ϟ
g�"���[�5�tq�P�������%��Sޟ��	��nXP�J/BN��We�3�ZM�PJ�
��Yg��
��O�7��<1�ΕT?��q1��/|@����ׄ�?����?���?ͧ��$�֦��qLȟ �iP�5�Pё�Q�����Sҟ�P�4��'��ꓦ?1���?)DJ��h��p���2.��CG?+%�M�(O���Y�"�z�'���?�]"L(,	�ًkV�b�䍈#H�ҟ$�I���柰�IO�')ҩ�"���`�RЈ�U]X����?�����& ޜ��I��$��:F�<^ ���S�p�xb��h�I՟��I���Lny��'�����ӳp׆(�U/Y�F�(@��kʄ7n2)�	�[��'l�i>��	��\�ɰy9,}�oX<}�8�4%	U��l�	�T�'b7mP�3�N��O��d�|rs��<Y�T�g*��!�4�H�a�O~��>I��?��xʟ�(��A�0R�2�8�.[9x����"1�dP�����i>m����u��|�M�~l|�!�Y^�����U�1��'��',��Z��۴j�X��s/�7@��:p��-5*�+SHΊ�?)��_�����i}R�'��9H@Z�����A��^N�"7�'?�7��%g���?Y -C�|}T��,}r�ӱo��y�s���L�
�P�yb[�H��ȟ��	���	ȟ �O�te�V�:�^E�!��?I3I�/tӲ�"Q��<�����?T��y�%w���ibm�
0T�ك�G�R���'ޒO�I�O���ʀQM��2�>��U�)t�l5��ĕG�ϓ^�����o�OV�yL>�/O��O6E�F�Xp˶�$I�Z{�1�J�O��D�O��Ŀ<A��i. q���'��'��㳧ߙ3w�2�Z.�����ĆC}��'�b�:��σ7�hal�2tp�gx���Ox(�'D>�p�O���Ӎ9Zw2�AK~��Ʈذ,���ä,�7I���'���'�"�S����a�T rjP�E�(|c^)��OʟԪ�4Z����?��i��O��;/���ȇ�
h9P*�z\�o��l�1�M[恏����O�R��:�����E�`��[dIsQ(���UK>Q,O��Op���O��d�O",����x��X6��_� ;q(�<�g�i,�4�'8"�'��@�"b�}�Q�C.˜.!�{e�\D}��'�2�|�Ou��'���ÈؗEے��%jRj1�A���V8*��U�Of�d�-�?�;�䓶�d5a��6�W�o�t�(Ѝِh>D���O(�d�O��4��ʓO0�v&ƣ�R
A�3�B�h%HƵg)~��b��� l���
)O|�Dt�^)lڒ[B6Nq�}8�Č� ��J�m�S�I� ��}) �O$q���.�i'���ᣏ�:MP �bV�r����O`���O���O��)��?qT�7��D����ԏ՟y��e��ԟ�	2�M��*�|���<ț�|��&)8�a����%����l̢Y��O��o��Mϧ"��!M>�u��0��S�nZ����Պ�#h\Q2���O�%�J>*O�⟨��\4c,E#q �lgF�x5`>����U
r�"�'�2S>	`�EO2��惀 5b$ 5�=?1$X� ����('��'��A�"E�����6,j*�낺�dq�����4�FԂ�' �'5XL��S�D� ���c`�q:�'*�'����O��I��Mۗ�Q�;�.yU��-�*u:�n	�U ���?��i�ɧ�4�>Y��*Tf
`�z��1�
 @F� Y���y2��
��Ӻ3��ٹ���\���D��~���(�֫@v ��os�T�'���'Ub�'��'�������N�i�$�*O�b4R��Wf60������o�S�8"������Ir��Q��,�h`��@��?�����|���?1������$��\`=K�l�0C ]�"��:L0�dֳC�b�'e�'��	ٟ���r�x؁"��q0<l��� `���ԟ�����Ȕ'n�6-\��d�O����<i��[��$�U��j�5|LN�`��O����O�O^�� ��A�Pr�M�
���P����L]�.�����y�1.����O���B�#�6�J�Ĕ�LF$�p��Ob�d�O��D�O,�}���0���Td�ȡc���J�h��[ʛ$�;��Ŷi��O��X�B$�'(���yRA��$5��$�O��D�O��!H�<I�k���H$��v�� ��@��T9�^E�Ď� GD���.�$�<ͧ�?����?����?�"�Z/|�y�4E��tp��k����$Ҧ�B�@џ��I��l&?���9'�̨�*�.�\��V�I�y<T��O����O�O���O��䙐4���)E��D+�"�xd����/�O��P>���K���$�ԕ'�(���C8������4���ar�'Z"�'Br���tW���۴m�p4��`:�{ Ϛ<eVX`"GcO�~�+��ܚݴ��'���?��e8��\57�ءx��ՍR���`b�����|Rb�
�A�SK�'��{#h�f~�P���I#?ӄ�i�j��<i���?a��?���?����ٝ)���J�֣�e�r�ݎ/�"�'��#~�>d���<Y�i?�'�b�Hq�[�"��`E���`����|B�'R�'D�*�^�8�'&)|]�pΐ�J�lsԣП,D0RR��%�~ґ|[�p�I�D�I埀��Rx�<�`@A\?�9�M��t�	my"x�v�d)�On��O��''�N �Gџ@���`�� �J�`�'2�듊?q�����|��\��A��R�6�`҄T3~|P���Ñ.��L�����������'M�'c(I��)����� Oh *!z��'��'B�O$�ɗ�M�(KDȔ�ՎM�l�dY�M	�Q1܅����?AW�i�ɧ�D��>�ir��R�P�?�VTi��O:"�|�)��p�zn	Sح�'�2�І?�TD�'��̕���[`NC:O���⃋/[L�D�<q��?���?A��?q(���1��(<fb9j��]�0 U��\ަ���l���I�H'?���M�; A$5w��¯�I*�����?	K>�|
��E���ĉ�nMj`LP�U�D u��>7.�֤5�@�j�'G�'��i>��I�O��S+]�;�1p1`^4]x��	���ʟ̗'��7m
�@�\��?V��"g욐hՠ�`�+���.���?	�T��hߴ&��� ��*:���`'��(9N(8��D�W�IQ�r�*�噠j�0�%?�2r��u��'e�R\tZ 5(���)���y��'�"�'���'I�>��I�~x�qJ�#�2qoD`��&��y�I(�M�)ƈ�?I�3���4���S'�/'O�US��Ҕ��<J�5O����OpEm>K<0�'$�)JX^1��:���b�#֭?�r���	�O�D+�|�W��ǟ��Iן(���x�I	d��82�߁7n
̓W�cy"�oӞ<�G��O���O���d������ƾ �� q�'T9Mi ��'�7�JЦ�"O<�'�*�'"(8dSte�[�I��Ǩ�W,D��?�/OphؖC��~b�|�^�8!�ǘ#"G4X2�Ӫ���w�ڟ��	ş<�I���jy2�b����N�O��Fgӻ8�*�pf(?bƴ3=OB�n�D�I��I��MŲi� 6�ߕQ��!@vC�		���qƈ� u%�P�*�<1�Lp� g�?�'����wj�Hq�P�l�{DJߩZ�}�'��'���'2�'���䁤��1~F���-Nd̑p���O8�D�Oʽn������'�\7�<�$
��(�d���2���a��P�T'��mZ)�M��'(1���*O���
�jϨlY3��$j�����Y����/���~R�|�T����ܟ��Iڟ`C�$��-�� �0gÌd�����Dy��hӤ�҆C�O,�D�O�' �q���� nQrܫ���(_G�y�'o ��?	�4�ɧ���|0p���mS��ɞ�&�FQ�8u���[���p�>�Č<	gDe��\k_Ft31�
�+����O����O���i�<ђ�i��a򉞤tǾ�c�͒&���i� ��&�B�'�R6M>�����Ħ��s/=*����E�
�TARRk�2�M�W�iw���0�|"���4ڬd�'���@4Pak�.��7.������t��<����?)���?����?a(�.� �K��	�F9� b/W�����lE˦	�Q��iy��'�O�R�w��n�Rtɸ���dn�P�Q��xͦdn���M+`�x����*I��	�x�F pG�G[�)�����I��ps��O��O���?��AB<��⏬c�ԁ��_x�a���?1��?�.O��l�E0�@�':�-ϝ*(�xFEM�I^����"��'�$�>Qc�i�6�K�pФ�EF�
 I6�(�ȑ7 b.�@mh�J
8>@�\2I~��j�O���O���F׾R�9���J�a���8��O2���O��D�OҢ}λ}���+^Z�9��5,Ҙ`Jwa������4�������?���i�ɧ��w�Z���iKL��K�m��X�5�'x�6M���eܴ"f�HK>�&�U#ʈ�i&A��a��`�����4J���^�YN>�,O���Ol��OL��O���V$S�q�X�X��<� �i�l�OB���"��T� ��s����̙q^�U�#l}��'���|�O1��' �	k�Ô� ��,��`	�.bv�U�6Q�'avm5&w?9M>1+O���H�P~biK�Ŗ�!.t��PJ�O�d�O$��O�ɤ<qջi�M"%�'|�i���&C8H��)�#%����t�'�,7&�4��\�'���'Bn�$�r���<��eQ�x�X�0�|�eј딹����'r�"��0E�:
.���q$�8e�е�I	�O|���k�<��[A�찙�G�0�	!�'�6q���K�/̸:��!#0�Af��@d������-�l���rzf�r��S�<aX��C�ί82Z=�G�5?��ǘ�]w�HsG�=[��ژAN�eٱf�3}p� X�D�O��]�%�]�_����f�4�ߒUf��3c�%р ��Su�@�,��A{W�-.Ş��B
=["4h���a��B�o�57`� ��G�0͠����':��	�� ��oO�TkvcH�Cd��C�9����i���'aB�>T�����O��Ɉ*,2H)7��z�D�p��LNxc��1ӦS�	���	�ȰN�|x���HW�<VP�!���M���%5 슥W�<�'�"�|ZcDX��'����O]$	4���O^�8%��O�˓�?���?y/O��!�ǎU�u��o��r�@E8D \3���'�	�P'���I��@v��:/���F�@��5q�-�(�$�����x�IKy��4KF�S�>Q��ҵ-�W;6���A8)&6��<�����?���?���'!��W��E�&�!Т̙�@�"�O�d�O����<��Č�E�� �G-�5�P�@GDˎ|��dP���Ms�����?y�
� 5Љ{B� %�>�S �ڙC�<1�W��M���?1+O1q�]R�$�'���O �Hl�l2l�!��ͼkq�qq�&-���O��H�
�㟨��3p���%=A.L��خ}>�nZAyr��p7-�O���ON���n}Zc
�}
Q�]��V���]S�LE��4�?��y��(������:;��T/M&}ؖ}�E��//țf�\�7-�Ov���O���R}}�[��%I�u�Q�e!�?u�rH�j�M��K'��'T��������bdW
h�&�L&c�>�l���I͟��$���D�<1��~�c��y�	k�g

v�T!�0	Y���'�D�Xd�|��'�b�'��u��hԹPT4�h%d[�z?v��(l����U�a�'��I���&��؇#6��PAK9���ZPh�=Ȭ�A�yq����d�Ox�d�OʓA]����1F �
� B%
$�1�&gJ/U�	ay��'��'��'ި��F�r#�Q  �F0L�x��J�sh�' �'9"R�@�ˉ����C�!�
��'�
u|�z!���M�/OR��4�D�OP�Ē�8��0�޸s�BN��ҡH�����ꓖ?����?�-On=B"��z�S�7�����SX�س��0G��ٴ�?�I>*O��S��O��O6rl�F�'F�
�IRM�}���4�?���dó+8�@'>����?�؆p}����b2|Ollq�^CRH6��<q���?�qk	��?	H~����aπ	��!@WMD�=G��{@�����'��i0r�}���O��O���gޤ�ɱʣm-��H��E1Pp�l�Ty�͋�&Rb'�i<��iy�Ȃjԕo��$_�V3�5I�4S���2ǽi�B�'I��O�O��G�9�0�6��91/��	c���t���nZ>3v���ٟ���ߟ��S��R>Ya���N�� �#�����hۛ�M#��?y�Lبis+O�Sv��ma(�e�̆:
j0�C��H��m�<)Em�7C�Ow"�'\�-�a@��V&F���E�� 8��7��OH-��(N@�i>���ܟ��'�)���%�v�`f$єpm:-���t�<�$_�k����<ͧ�?�*O���8�d�b��=�Di��.��b�o�<���?Ɉ�'b�i��(��ˌ	`uѕ$�=D ؠ��P��d�O����OTʓh�,%B�6��Ly׏\n�}��@'PRF0PtS���	�����by��'��! �" ��s޼,�U�N�$x%eH0IN���?9�����O�s҉�|���h^L*u-�&Q6��C��bU�БB�i��O����O�rB��9��'m.��EC�A�>��B�
-X���4�?�����D��&>����?��	xqv�# N�0ia�-v��#X7�<��?I�E���?IN~���C6[��^Muf�o%�hJ��Qަe�'�B�"(sӒ��O���Oh4�A9��gB��`A�S&@':7UoZ��I�t@T��ɫ��'�(����>v��1���X�m�>4cT 
9�M!�9?����'�r�'��d�2�4�k��YP�!1�ω�e�|12G�H�DK��'k�'��X������N�2�A�����RQ4��yo��8���@���Ҍ���|����?�vLU����4��Ri��!B��Wś��'�B�'I�	3��~�'��'�*J I�pk��	)^�"��A�i�F�$N�S��5%��̟���{yJ��,����$�F]�W��%t6��O��9]��|��'��\�XX�(�	`�\�{#"��Ԁ�?~� �I<���?Q������O~��QBv�� ���I������ӡR�E�G'�ONʓ�?����?1)O
�!v��|�e�]�K�FX��+��s�9Y�fBD}r�'(�'�ɟ����9 "��ie\H��G�l����B0Z�؜��*�>i��?Q.Op��:ns��'�?�ҐM�i�D�E$1-I"fJ������O~�@6"�:I�xR�[8�NP�p������C�M����?�+O���-�D�S�� �s�	[a╕zzݰ,C�N���17�!�$�<�C%	�?�J~��O����B
I�0�ֱ0)^0��O2�DO����D�O����O��)�<�;l�
<3�ʑwRtJ��lRTIo��D���N�D�u�5�)��|G�d�A�F� �̠x�I)U�7��%\<��l�h�����S����|*��+�s"�	aa����,D)r̛&O[*{`��'��IN�4\�x����tC��8�b0k��K Q0"��ݴ�?I���?IT
n���xy��'�����eJ�h�A�5(�rU�wn�&Uۛ&�'��'׆���)�O���O�)��cת��2��N�%|q��o����	w�<r�O�˓�?�,O����� DQÊ����p{#f^�-���a�i����y2�'!2�'F��'R� x�.����>Af��A�ԅl��E���°���<������O,�$�O]i6i�)���aj����lP*6���OB���O0�D�O�ʓ^��[�:�v�b��&+k���ab
Ѻ �iU�֟��'Tr�'[�'��yb��1�Y(e�8.�����W�V��7��O�D�Ot�d�<�6�Cc������<�:�I��1X��%5����7��O���?����?IwF@�<!���~⁘����!ȒO���r�A��MC��?Q*O��2T̑D��'y2�Ov"� �aš@˪���4�v��!"�>Q���?��v����Om�IH�QjK�V�J�mǉag� S�i̦i�'j�P2�oy�(�D�OT�D� קu��P&a�ƠCf�ӚW�,y���M����?�F���<	���-�ӟbr�� HW�V�y�rE�5QX6��<J�n���p�	ԟ��S7���<ɒI��8��ńL��i����֏C�y��'l��O���?��Гr����a�Ǚ}ۨ�CFbR�9 ���'8��'��#�h�>�)OB���4pg�Np�,�����yd�2�`����<���<�O��'�r��9j>��s�]�B4֭jc�v��7��O~��D�z}�[�x��wy���5��E
1�~�����gc�K��,����T,���@�Iٟ��	|y�k�hdr���O�0Y
�I��E���F�>�.O ��<����?	��S�!�����Q���ly�H�<)��?A��?i���$˪pF�1�'F�œ6g���ة��B�6v���lZ{y��'��	��(�	��@CM{���WÁ?RӨTã��211�Q'X��M���?���?!+Oz�hrjDX���'�H}٤�C��Ai��N�^���O`��d�<a���?Q��&S�@̓��i���j��B%��t:���+x�^�r�4�?A���L�в8�O���'���ɁD�R�RuGS� ����4�~��?����?�����<�K>Q�O�	HU.ř9��G*��o)0ݴ��č�y�HqoƟ,��ٟ�������Z@B�k�v��l0&_6v�z��i���'l�@ �'��'q�X�k��)����g$)�v�j��i3����Os���D�O��d��I�OX���O��"WMV!��;���>�h$��n�˦�A����p��͟ s�������^�]�^IӐ �8-~Ъ�4T�n�����ϟ�pT�
 ��$�<1���~����ov�y��. �@i����Ms���dɢ:�?	��؟���o�D�������3�D'CzX�"�4�?���A��ky�'��֘)f}�)�5��I��iЁ~���F�����?����?!��?�,OԼ{!���֤��R���	���b��>�,O����<���?���2��"`%ܰRn�)����QX�dꄦ��<!-O4���O`��������|���ʛ�j��?
	�౱�Aئ}�'>bV�x��ٟ��I�`~��I�76�-j5�<�p�g�4��0[�4�?I���?�����W
���O�Zc���$�
�3�~uv���@���hٴ�?9)ON�D�O��d�b����Op�Ċ������.��r�pcw���dZ*�n���|�ICyBl�K�h꧂?���"r�J(�H�ʰ�
T!�iـ$	*6�	Ɵ���Ɵ(���z�@�'��֟\�cUR)�@2�NW3zARb3�i��Ʌ[�=ڴ�?)���?���[A�i�A{�A9O�$rp&\�>)(��Gu����O�0OΠ��yB�	�t���	���%���
�j�����%2��6��OR���Ob�i^}R�@S��L�1S��C��E鹄�	��M�ah�@~�W���R��vc ����#�� b#O�C�^����i���'M�ҭ�������Op�I�	�����H ��6��S�$�6��O˓w��S���'ur�'�� 0W��4H�r��7�a4jx����(\~��'���۟��'�Zc��a(�'�
N�x�k��?ɲ��ON5:O��d�OB���Ox��<��	ǐZ @dE�Z��@��Vo�iBQ���'��U�����4���6O��@�1`�j�nQb�:�
`�c��I����	���	qy��2NR����p"�Fr��)Ë&?�7M�<Q����d�O��d�O�ыR7Obi��V�F�\��B �d(\Ij7����	ԟ�������'�S�n�~2��+��m��L�1U��p�7a��9�	QyB�'��'AD�'G�s���P�'����@ ��&z[�9�@�i#r�'	��d7n�����O��IC�p�K7#�;�����F.syR��' ��'cr�������#�0�y4��+A�$Z&7��(nZFy2h67�O"���O��)f}Zw�B,�K��vü!X��Y6=S��i�4�?���S���ϓ�䓅�O��0���p`�g�N�4���۴&|��Xưi���'���O3b�� �!(T���Ͻz��}+�'��MKD�<�O>)����'ц�Eē�\}�1�f�	�Iz\x��m~����On�DM:�H��>Y���~B-_�[X6��֛7��cI8�M�J>q���?�*O��d�O����TmZ��D�D,Lh�C.:h��io�I	5xO���OH�Okl�?��e�'+�-���2��?��I�4�i�	ay��'���'���r��HZ�m�/�luva� <��Z&�����?����䓟?��=6Fd���)/1����q�*�2�䓊?����?�*O���@��|
���%(��`��5ne��L�h}b�'�|r�'��h��$� ZuX��ՍO��Z��%i�x�qY�d��ҟ4�INyr�S���t���ЁF����a�}�Bm�Wn�ߦ��	t��	�����i�$A<���2�ݷI�x4���qu�f�'"Y�������'�?)�'�d[� �	,�����Px+���f�xR�'���߮�y�|�ݟ�,K��7"P�B��M%j2��i(�8�v�0ٴXJ�П8�����ÑzdJ}���B�@����&�G,(7�F�'��%��yb�|�iV�J��pI�CR9i� �F�(8��( �.jp6�O���O��I�N�I���B�n�z$�[%"�d�XŴi.\<��'��'�Z�$E�֮5��oW:-����E�8m����	�����-��'�R�Ov�ꖤG\�  & 9eX��ӳi��'���b5�'�i�O��D�O��'&U�8Ј����G�F#"�Ǧ��	#q�:���}��'�ɧ5F�Z�J�q��/{��,٦�Ǯ��$�2+��ĩ<����?�����$� P��J�>Am:�a�50���1��j�I����Iy�	�����<ruC�%���w�99���r�v�@�'�"�'�Y�0�1�$��$��5U��"/\����C�����?�O>����?�ъٯ�?���B$9<IC�л_��Pr%�+�I�\�Iß\�'`�,sw% �i��F��P��$̠|��@�bJ�?A�doD�'�g)m�B�'N�$ْLЙ��F�e�*՚��$13���'�\��fHI��ħ�?���ö���`rDE�k�5�\0bǧE쓗?)C�ߔ�?����T?�%y����h:�>e!G��>���rA���ʟ��I�?���u�]�Bm]�MIq)G-� �4�?��Lݸ�Q��l�S�q$�M�LմN����B��M|�o������4�?���?���OӉ'��m
�j"���/�#���6Ɂij�7��������	�9�v�ݍ{�04q�f�ZP� RG�i�b�'JR'��DnO����O��;��M�fg�	�i�^]0c�ЊFJ0����ܟ�ۆa�A�T�I$*Z�v�&]��P��M���X�D�,O��O��|�iP�N�T�!�NYe-X��.q2�:q���v/�z~��'#��'��I�V���*�ڶYF*Lywd�$J��m�4+�����O>�d�O��D;�ɹ
�6dy���VT������@�D5@���S����T�	؟��I蟈` F�C��O+y�F�q)�e��}��'Wݦ��'��|"�'��E`
6�=\ Z��f
ܞ]L���&��$n����|�I�� �'����3�~��\ ؐ0r`�3N�x���9*k0u�s�i'RW�T��ܟ��I3D��Iן��I�� ��!z1�i�`N��]X��M#���?�(Od)���H��'{��OB�A�*iT���OA�a�	�%�>A��?���V����9O��ӵ9{,9߻D��}�%W�6M�<��-W����'r�'��d�>�;jP&xC�L�}�d�!�"^}��o�ğ���u���	|�Il�'G�������E�,�AR�2g��n|Az#�4�?���?���g��dyR��!I�P��$fʜрӫC�xl7m�%���9��3�SП�Bd�v����_�a��iB���MK��?��i池�_���'�r�O��	Q���
�����HA�Sp�"&�i'�'ϸ��S�T�'�2�' 
%�B��]i!�/t:H�b�
b���D��g��i�'���ڟ�'�Zc������w�H���47ڒ�!�O��h>O���?����� �e	$��+u7���iT%!� !��<��Ify�'j�	��	П�ap��-f:���ڗHrƜ���
e5��	Yy��'��'e��'϶�1�ҟ�y�wi��*�&�X���7-���E�i�r�'���|b�'���\��ݴ���3�i�P�z���&H{8��'�R�'U�Y���/0����O����	�Tt"1�Ye$��`��@��?����'��x�&�$]�d_�����Dku8L�t���Ax�F�'�r�'�"��l���'��'�����(Ⱥ��W����@
���(��Ob���OҬ
�(a1O��;�Є���LaK:tH��	�Q�6-�<ɤ�*XO�f�'���'����>��u�f̩PhÑ(p���皍m�To�̟h�I�nט�ԟ�����0�}
���� �ڜ w��>r��8AU�y�`��/�M���?I��:rR�X�'7�������@z ���
%eh|�tӢ�<Ov���<y����'�4f녺K�H�G���r�2���&u���d�O��_v.��'K�I���;��Qi��XA�ă���rc�4n����'�x�����)�O����O�Q��#Ρ?WVx*�
4r�Lh�&JEަ���a򐠚�OD��?�-OF��Ƅ	�n]�Mu>�B���5hXpek4V���oy�\�	���	ß���uy����^��d33(��Z�~p15A
>��%g�>�.O��$�<���?��"8L��[2.j���Պa_��٥�L�<�OB�8 F�
I̠��ooj	;����BlV�:��x�	�;�U���+9|(��O�-���"]͂��U���������K
K��q��n��@4��l��k7T��l0�.���H�_�(J�+ؓH��:��י��	�D��j��m)NQ�5ŔMx3M�?7|�e-׍t�<���ڃ9�<�Q����4��� � 8�4�
#"�].���SJ�X2�P"�j��1N2i@��� �PY&�E:��{�N;dM'�"��A�E��p���m�X`R�'N��q��
����W �j�r�X�.�� `ts�L�-%Z3�� �z}Y��>����n�I˱D^^�D����T	*�CC�~2��ƚE�P��Q�Ӷ.��p�t�D��m}R�'4�>��>	|k�$�J:�"�F��=��C�	�]t��Af�	�����R�r�h��$p�'�V@��`:�6�X;�*��ei�>���?I�BS�>��pQ��?����?ͻ �����H�} e��ѿ�@z��:X�F����&P�g��83� ��Aj�7HC<Ds$̀v�1��.����:���|�� �~�%fX3=�BH��Z8}�����O�	=ړR���vbZ�<��	tEW:7?���ȓ*K�Ĳ2��4Rc�NQ�;����'��#=�On�ɶ�*�zs�۬2�Q.SZ�Y!w�*Q���Iڟ ��џ�z_w���' ��b��C[�[��Q'�]"{6|�8��K%JQxe�׏݄A,��ā>p�D���C�-��
�cD� XJ�g�{��t� K�24W���{}֍Is�]6�V�8�]�=`(���'�r�	}���Y��bT?d�5�WN	'�8�ȓ�� ��=)�b��ë��h���<)4T�Ԕ'd�x�HhӮ���O�<��t_����AN��Da�`%�O��d�����O��B0�m�_�"6	BW�n�4�;��B����$T�'�lc������8Y:��1��9�E?O 0�4�'�rT��" ��oDP�`��,�k��~���	ş��?E��a�[�*I� \1�qrwJE�xR�~Ӣ,h��_6�@x�$��*%�AJQ9O��?T��Q�|�IO�4gŷJA�(қo�@�DH�V0��I��I���'P$ȖEV�D��٦� [���T>��OH�@!���",U���T[R�r��H�b�í��}s��F��/�Myt#Q A�"h{%�����ɛA�P��O��}���X��p��ؕ��]�%�O�S��d�ȓ@
T��"F�����oֺ8� 0����HO�<S��&0��� �<8�@�Ӧ��I�|��.~�yR�
����	ğl�i��C�LX�
B�K'` �]dFc`7>�\c2�	 Mk���I(����|&��1"g�=D"���Q@�.V�de�O		>I��� l��Z�[?{�X�>�O�)H�� �`��oǬ?�"�#�?�	�=�*���|��ī9�,`�Z�q&��`�`���y"���e��	@%�,�9�V�������8�t��cM�Y�JVW��\�^7Af��$�O��D�O��dB޺S���?Q�O�������=2�:i��j'	@9���O}�|��Щ:[˸�3�}Ѵ���I��m�L���X�*���qB�X����p�M	�$E�q�A�@A�p�'%��6�"ؘ���-%�����m�e���$!�O�!�X+y�6DhCJ������"OF�Z�ĵd���(ЭQ������R�*�PÓ�i���'���e^2~^����.�#0d�����'NbڑM���'<�	*O�j7M<��V|"<��'�1a��}p"j �_i�x���Y��O�A�W�Ǎ^��a����F���"u�'6x�����?���?iwkʱUD�p@�,��I["�W����Ob�"|z��T9T�q���A�p��B�n<�`�i:p���F�a����Д
�-c�'��+kP�ش�?�����[ �`�$�#D��+��F4� @�O�&ky����ONX:��O�b��g~�r!���c �j(f�������	�C��"<�*tnW��@* ���dF(��'�S��@.c������~ԉxu��b��T���ɯB!�$.l�~8C�^�b #̘6.axd?ғ��%��ףiʐy
0ş�j�YгiX2�'1bA"-x�H��'��'�w�J���âS��a#�
c�-��
U��yV�en`��%"&X��ǝ���'Tr��ϓ8?�`��(S65[������5��yr$���?�}&���1B�w�LE@v�#	�hX�0�<D��&U?,V	Ѓ�@�^�[#�4?���i>}$�T���@�r�P���o8$s��/.k0� �@����I柼���u��'�?�6��B��8D�����՜y �xk㄁TN4���'�O���r�*s�p��'.ؕ����QcL$�'�pA̡�A'QTX��hF)б�B��&?]8'��u�
��,�O�iSPOB��15��	�����'w�'B4�BO��n����l��]~���yB�p���OꄹaJFA���'��P��DO+>���I�,Ȏe<��3P�'_2��D��'��)�3�r�K��ĆMYNz��`�p� � ��m�(�	AD4N�jP��'p�7�Y�&�x��Rk%kV�� ��������wB����#$�'C����?�)O^���C�;�� ����m�|[6��O����68ƅ;l�*)��qr��+H��G{�O�7�D�#��Уu�ݵv#V(2��"0N��<�f�Ʈ}@�&�'	�]>u�1�ʟxX��=5�"caD��ȩk��ğX���w����z�S��Oڐy�%])*OpAi���[~�)3�>��ȍN���O�� R/[���eNoo�٫N� �j�ON��O��� �ӓ��1���&�h���p�c�X��ex�hK�Ď�Y�,Hu,�}����<O�1Ez"Iӧ]���Fcý+rp�w��^�66��O��D�O.�K�4�����O$���O�N�y����˹e9�L�*�2$��@����v�h��4
�uSF"�F�g�I�0 ���B���f��s-9`?�: �=D-���i9p�l�h�g�I4n'���E,��Oǘ��UhV�i���<�hV̟�>�OȜ�Ѩ�+q�bU@�d�<|��t"Olp� ��dG$�K'Cˌ�F�w���Y����~?^� �l\ �N,�f�+sH��A��Ň 8�a������ݟ�^wS�'���]�!"LQ�Cn1:��l�r.���aO�퉐��M��� Y�)��(���!�d�M�N��B���jS�,+ᡎa��y�'���-��C�Y��suB�y�o0E�����ѡ8p :V�[���'ǎc���!�O0�Ms��?--4*\[R&�:;&�)�a�A"�����,��\����|b���+{����b�ȹ6sb�HѤW��#G�Xr���"���9 l��d�"T-+�4q	h���F��<.��hi*9��@�-ڕ=u�m@�%5OF���'@�'*IC��	@�bSń*tq���'>,+тL61�kbLǰ�|��'��7�+|<�,�cݤ-�aj�"��u�1OV4�t��ʦQ�I˟h�OQTp T�'L8�S��l3�Q�w�ݪ�����'�2"�.MCb�T>�9iX���̏�2����"oF 7zrȥO8Q��)���Q(�)�N�=E����#�_#.t�'�����Θ��O�.��cZ	��Ҷ,͡q$�'�Ƶ��nI?1R�%�Q�@|��A
�
����KUA�k��X���٘/ΈtK���?�MS��?��e�q˖B��?����?��Ӽb�Y�S��[f匤y2 @Ǐ)��'>� ϓi� �ӶT�܉`�	�Tm�=��	^x������+�f���d�p��m:S �G�s��}�)�3����c=�(��/�(�  �ߥZ!�$8k��DA+ׇ)�D�ؒnY&2
���HO>qj��À;�� ƃ��a���^.Y|x��Ο|�	Ο4��q�$�'X��C�/\R@�e��!1��Ų�A�:u�x�Ɇ�)�O�&h�#!��3Sh[\:�T;7��i�<��r�ݡ�l���'�^}!��!��=bh��3� ��	1�?�2�id7��Oʓ�?ы� ,�0���QU<�a�Z��Oʣ=�O۾�P�F]�e���_�T8�����|�i،T�7��<���	�A���O��7i����0+T��͘w�R��z�D�Or@��	�O6���O���C�K�C��O���0䘘t)f88)�K~\h"s�'&9���V,sal98������'ǊPv9P�C6j�d��Q8�D�� �O���W˦Q�I.aE�l���Y�F6��En��_�<��'����SJ�����Y8?T�x��]�-�T����O$�n�:" d�Z�L�4��`A��G�j8ڴ��d'@,8n������b�D�R�[�t�k�oD
0�l3iͳZ(��'�� 9R�'�1O�3?FթZBR�g雁E�Z}�CmZg�d��2���?59�� �
�h4��:w��I3n/}�Ĺ�?a���?�����OT�qi�OV�Nt:)H���.(,�ˈy2�';�y�h��\1�^΢�E�՛�J��ቆ�HO��I<%[��ht�+�����Z�e����@���I�h�)� �՟�����8�����r5L�a��F!� ,L���k���)D�0�)�l�g�	�Y��M�톫"��5(�*yV=!N>�B̒Cv��>�O����lԍS���j_���'7�����,O<��=��F�N�uŶ�ʴ-�-aTC�W+jq�Kϲ^V�����������?I�'���c���>( J��$�[$K6dr�@�G����'��'�x�	�I��<���D�� �奇;T.�Hk�b��1��XQɓ�e~���ũ@A�3 m�/'� ���S�]���1�C�7캵SF��f��X��h��p��"u�N�HH�a�D#<a3�7� �����W�t�ʳ���z�D��Dg�O��DW릱��iy��'�����Q<�Y�'J4 @ׇ��8�)
��H�h��h+�'w��#]�,�&��_��H�y��;�,X0ņb�P�dTL}"[>�2��)�M����?)$+��.�n1���Lui��c��H��?i�P851���?i�.춵aS�i��'⢱�ק���ڤK#*Еm]J�zǓO��4B�� �P-|���O��X&
�%� \X���jʌ-'�'�Z������f)pӚ�DL�!zh�U���s$3��!>�ʓ�?����4�'+��ED�P�j�Ȳ�Yޮ��	�'Ԯ68i48�E B9���qs*�	520�o�[y"�]�{eNБ!�'ARS>!(&HF� z��� 6�
�F;�\����^㟰�	%I�)�,ؤO8����0t|૭���'I!f%�$|1���KJ���O��rRL�3B�A�2o
5v���B�(��Md��gdK6V�����<V�'����l#���'w����'>�z1�u��if�H�eت��'���'p��'&� @��ҽ�Vg=R��a�=O��FzR��%UН��&�3o�@���C�p�z6��OR���O�=��I�SJ��d�O�D�O��;|Ϟea�Z�1e�P	�� �l%�s�yrB�_�ʏ�D��<
J\R��	6&��g��.!�Zc���J�& �q��'*�Xj��ÎG�*�
�!�ͅ�:G��'��aZ�:�)�<1��7�;�)�,-@bJS��b
�'�U��.��}��Y ��2��p�O$�GzB�AZ?�*O�4ш�D6��"��Ҽ��J�ݢ9F��O����Od�$�պ����?)���̒B#(Ť%��B5)'*pC�'���<��+p�1PÌ�N
�0��R�~��A�4S�8{���g��uR/�E���b�=(�l�cڂ5ڊ,�Lɭj�,�$�O�	lџ0�'���D���|�tjW�L�n	ī'd��*�ODyХ/�z5���������6,4��^��j�l�Ky"�M�1�םퟬ�ɶ;V�2���>lg8��*T�n�����	������|�b&����z�*]^�Ԥ�4J�d����Rr �C�#*h�	��6\�����؁o�b$�F�����Q�I)	,4�P���]p�4���:O ���'���'��ҳj�Ё�A`DR�&�8��T5L��ß �?E���O�LM#s�_�G���-�xR/p������()��1�᪖�Fk�s<O,�R�Ցb�i��'��S:/W���	�@��� W8E��!_R�
T�I؟��wgިB:v=��)ML~*�@ʧ3tހ����PYb&k��(�bQ�O~����*V>�ŢA���r�"}�U��� �|LXC�$]���2g�Jl�Ĉ;H�"�'��'o�Dly�bI���Tԡ��o������O&��8B�$CG�U�}�h�j`ߦ�ax��&ғiq�Qp��Un(�%"3�F�-@�\�'V�}R,]	g�2,�WF]�/�ثMN�y�m�dL�f�� 8Ā	ǎ_�yBKBJ��%�3���[���3�C0�yb��}&��zO��|�d��R��y��Ғ^�(��"��� ����y �)>�I�5-Cy�qF�=�y2���]��uB�oW�Nf~������y�d�b��ҝK�r8��k�<�e��(A�ਇ�!� i2F^u�<IT��L��u�R'w���cǞu�<�@�N�ꕁ��H:���P�Yi�<��  B���9tA��J�~�<i��ڪg|�ӆ�����a�x�<�SA=w ���s�߁~��s k�<�udJ�Gt��1SA��P�$��r�M�<1!]�&����`J_	"`�-
��F�<iP�ӟh6��.���x���@�<�c��	��M����%0�(QI�o�F�<qKοyDUi�-آ-8�@���w�<��պA�H`�r!�a<]����r�<Y"��4V�} �L��8�*ݠF�X�<�"G 0{+�P�$%B�Z�������N�<)D=Q�\�Go�
{N  K��u�<�"�\�q$J�䔂^՜�Z�L�<Qp��=�^��d�N����W��M�<iGN�9=���(T�0L���I�<� N��E!A�6T��/Ir�y�"O�lÇ�D&�xi�Q�ǙX�T	�"O"}�����r�D$�J�'�x� 7-�j:9�'>�����O�Ϙ'*�@4�U�3<~��e�M�/L=Q��g�T��@ҊH�.�rբ�7��"��1'g$����zxs�&[ʠq.�6/m�t86�Ś#��G~R��0a�xk��Ñy����ן~ ��؆�H��L�h��
�"O�8�B瓔M�r ��cI�(1N�!1�O�m���_��E�q��Y�]G��%P%��f��ՎlI�*1�yb���"�`���G�x�<�kT��".�Hh�8`��S��u�-�媘�&�p�э���Lyp�:�㝑2 ƀ��v�azr�Ɍ� #��Q���dȥ��4���� ��u`�K1�V:�L�5}�RiKU�'�2]H&�_i"�	5n ��x���y�n��hỗ/҇`j�*Z�caɴ��?q�$�K%<؉P]�R�d�I�H�)�y2�6�� s�F�.�S2/V	2{ � í2�h2�.B e{r�b7�-vT�O�r�`�w��Lan�k����F�.�
�'�20�I[=l��hjw
��'D �X#!;��r��r/�{D��U�"�7IZ?h��b�����M�����ewV�#��0LO�UI@��?��税� hP�� � "Ϣt�փۖH�.��s�0j��!�$Z�*��l�דT����&hA��"F�ǡ|^���<aƆƣxV��i������`������عBԸ��u�Й��=JF/T)��ywA�U�<g�>�ژaӠl�H,�5xF`����+R���0��"zAo�~��O�����wFp���Ev�M����O�DY0
�'b��B�έn�`Xاj�6+�U�J�>h����� ��"Fh�D-D%/j�ϯj�px�=�qB�{D��ՂȈl��9z!kAO���*�dE4`���5���w��M�@O�k�\([R0�43Kє!�t�pǕ�eՀP��'��l��j� ^�f��42 (H�y��0:�I�x#��
䩙�ֺ�J'�����;�x4���{����Φ=�C�I��l��vy��eOB�D��S$�A?���R0 ��M�f9�#2�Z�8	����'b*����n����(�%ޜ�s���t���+9܌��AK�?���|皕h�q8���!��1;�`<���X�R4�Qc�8b���38o��*A15����'��{���3M�8��@�[nP1�%�G ��'�4�H�@b��7�F�~�Ad�Z	���D�>zm����F[���k���-D��2O���q ���:!�I�������ɩӮ���MоYW�tsm�~M
����K�(�͛u�]'qW�i�Ӭ��_S����E��9�qOz�i��E�#�:��`�X�B\J`�Ǧ��F�^;ƦӉ�p>arfԽl!��p�� w5ԈpOf�F���*��L��,2QO%�3������m�Nĳ{����ҡ 3>��2|Os`#�<�:M�FT�&o�X� ���J
�"�H�1�ax�Κ$ ŜUP�� �R��� "A�w�r���?$�h�k�m�&�$�G��� ��Q	(�6�b�D�d�P(J$�P.U����]��@�g�H�Oq:hiv�<)m�b->�뤭�= j5�1OD�'��qħ^6�xH��U\|���]Ct�E��')X����^�<���s��NE��yH�y2�D�NUPa��Ό0N�& �wJsN��P6Om�	��	;&���! `��kd:)������aF?F���®��MS6j�ߺ�O*C����Zc}ܰ��eB�w��,#t�9&p>�;�'��c ƵG
XA�AY�T�T���b���~b֕�X@�II�|��.q�|��ʒ�r�����H2uMVAS�y��h{e,��f+�(	�#� xAcЅO����!;Q�8� tY���"�  4lD\�@��x@aԍ_���'(�P�@D)I��PX��3��y��sB���R(E�D��	���'����,��:Q���v�ɐ^(ljSg��~M�9�M�/'�{"oK%,?�I��ݗQ�r��FOY<9r�U��+�@�|��9��'#`䔧��c�� DY�!�#��c���C(<�T���sR��p�aK�&��EЅ˚*2�#<QA^����-A3_"��a���0PuF�t� �ƍ�4�U���%�)��.$���t�Z,(h�-C3EQF� x�e*$ @�H��zt\ݲ��!}���}u蹸a��#���@��$��'dTX�]�h��u�*[�1F#�O���v%E�"�b�0B`��J+8���'_Bdi򘟼*Ճ��(8�Hr��W��D٘#BӋ�X���7�|���V�my@�f��/#Dq�"��-aj�ے��!F�Y�6�'���0��OqP�Z挍++TQښ�y��GeB��@V�ytt�ڷ�V�*�!��7�l=wl�j��pY�O�7Chh(5�Ǳ5O6X�Rf�Qt4�9����V��t�'m�q[�G�w�hi*�O�B$�O�u��1�C�T�U����I������P?'�h�d�'IH �ELh��E
穑���g[R�T��N柨QЭ�Ey�1�M<�=�Rd����v�ԻJv�]�6��U~"��3���DeZ	k܊�0��
��M#���=5��Z�n�eS�������G�ŚO����6�M!�zx�D��==�a|�J�e���#ŗ�
���r�.-�(R2�^�|�|��ϓ�y� U��Q 0�
�H1"����HQOT��Z�9a�4hcZl�Z��v��H��2�'�5jkJ5,Z��r��`!�Rb^8^#2��[��Г��2U(f�Er�ؘ
�n��H_:bJT��1�����c$ұ7|z��邟h�(rT��	}���X��E��M��jN�]�#���Dy2m3<�p!fiB�����õ�����tr���t��4�2�� ���}���K�i�J�&�VX�$3oo���i�&*$m���:<8���r�@��b	�shJ�G��`�SFq�O�����>H����D�z⚯o�8�����������t�.}���V�yv=�=��F�^�v<�0OlPK���7K����8�% �E3���Pk��WZҠ�%��U�'D���NS�=�^hK��x��$=6��e���;"~Ͳ��W�]˲�a'�Mv?�`��?���|�<�Q���h��)�Dٳ\ff�tn�L���'9�d�l�3}��3�vU+�K�no��	F�D�D�Z�@�dG�?$����M~���]�BVz�f< \���R��69��7�:���<��H��v�� ���Tw?�ӥ`�u@ᢕ,1[hё���M2�$3��,Od���H��ܸ'�ȅ��!z98�C�MP<�ez�)H�H�����tX��g)���?ex�w�2%!'g�X���s�P;4x�J�O�L��������T�ߩJ��&䇡Hr���у|?ϐa�E����u��Q��Z�;yx�ܪ1n׉��@��a;�ɩWF�A���|2f�|�rcY�[�t����Cj��ap��f���DǏ�x�;�N=lO�N˰gf����e
�����$솃��yJ>� 䖣B'�d�I;hۦ�)u"�Ο�'o4����(X'E�����E��R J3�	697�^h7�� �(���o��%rV��흋P�.��gU�yz�Y&oE,\޸
�ү>�V��S��y�h�5~��Qcs�>+
���j ^vXᓄ6�n�㷪�;)(F ���e�D3y�,0b�ݳcMp���#
�?����"c�<9���<��ם�SMў�9���&��01���<)��y�@�q�{�虼�?i6f3���Ӽ#BG�.qK�u�ӎ˿)��$㊜b�D��,J��hO���gZy��� c=��Ѹ� �C��,�ݖN�����'F1x��ڲ�l�O�1`��#��*H*6�n	d"V��J�cE�U2�؀У	Rh�r ؁ҧB� �b+4�D^dc��J~��}$pB��_\��0��"��$�+IB&]s�r��"�T?	��� l�UZ 9O�չ"L�IB��5l��`�H�kB�p�  DzhQ��f�"r�O�-�ED��Q;�b\�r�8�(Ѓ��e��?Y��jL�28�*ԋ�B����s& hT���e� Dvr<�5��	=o��T�I���yc��!Q��Z�`P<�B�)E�?8��(���e�"=��8�Ȅ�W�.?��nѰU{�M�UDޝ~�̍pbϓ�2�'����ۦ�9�iʂ!+����$'h��kנ�*c*��#)�	�j�*��+��1jMp��Y�6ZA궦#?A�i\�DT0ūҀ���4F�k~�V�qODUrA�âF����0N�4�z���V�!r��Q#*���iX����ja�G�4��c�8{���?˟����C[}�< qd�R�#O&�p��|b�B�c�&�r�+����Dӣ�2��'�Ƥ�!
D��Fx��֗/x��� e\
��'��>�I�՘Ł��E� d� ۥb���xT�I<Z\u
D���qO�Ӑq�2qϻ���$+w쉷M
�F�h�����O���{��}��6b>(4��E�YfH�ӌ��y�1OH�ׄ��9�a!�R��t8����\oA,}��jӕ2�^(��΅�Q��y�bõrS^)��ƕ�u���,G� ��EpjU�gLؽ#/�$U�rU��O$'!V�{�b��IP���?���`	�x�D�$,h4Li'Kݡ^<��螧T�I��FӴ62����$ˍEQ �p��F�7��t�al�+���Z�DWAj��>�Ą���&�u�'bJĊG�N9-�\����0xj�#�T�8���&�U)/�.��=�O��� P?��YK���-6�䋃M��O�^�"a���d���`w�L�xXy���Rf���O��PS�k�*\_Ȳ� G#(����/�I-c�����u8f���M�+�rc�<�E��l@&�pB���q�z4 b`ΓQ��l�<ӣW#`����9#P�;��F�`��(��Oߒĭ�9���+R�n�
�A�"*z�,K 薼S~�xR#��>dV�Y�GQ�}��(���0d(���5����/�)�'(rpd 'jV*�=i��Ζ&�:e�㉊��e��zۚ��	�O�8�(�Ν���Y/;�ڙ;qI^����e�̉]����{*�j�1s�b�����]4��p�@��F�\pȷ�!}�=x���gQ#�޹E��F6�l�ÅD�*=�މB��zi1OވF��:��aa��V�t��w�ĜN� J3,C�Pɦ��	F�y���� ��tC�$�'���A(��dJ"ɔx,�h��bX��E([
R*���gy&�B.��z�Z���(U�"��ys��'��` o:_�1�I�)���GS2Bx��a���1S�@�Ƃ��4$!����y2AK�v�V�9$��+E]X3W i�铗�' F�{���+�X1S
6�y�ρ�`IV�+C�����97)�UV�$e��6��H�'g��]*i$,�ƅ��1*�kW:g�d�DàjT�A���F:v�qRGF�?-�&��'j�$�3u"���tt "��|$���#����%EW'��	'�?� ���J��� 䲀O�H]�͸v!�p*QOp$L��Mʬ+��I��A��� O�T�S+r2"���	G,	���sF�ޝ!���I�=pŐ� X'$�S�?Kd�)žith�R7�+!q�9Qt�8)F}"G�5CN�/�3E��郗j���Ϙ'αؑJC�;J�1U�ì' ưX�O�Aa$�Ƨ�@�c5��;3BI�=Y���]qΡC��l]&%�,�v���Z���@��mBH"qF}R��yg%�B$���kX�6���&)	ֲ�"4AC;��c�l�T���!��-�'D�$�-{b���dS��|�y����#>�aG�Au�m�j#�S�u�������Ov�p ��ϔ�'��H"��(+�f����|�uH�~]�"R��<���<���5>�"d{��3}��I�<>c��c��)YH�k#ɉ\��ϡvn�{����	Ь����-��鉠!�4��g�L��IS��<)��
r����b�#۬e*B"�b�������Ğ�,��٢�	�4{��CvW!�D<M����p �+x��T��F!�$I8|ڄ�[=&�|`:�%R9K=!�d^�%M@lkW�A&L�y@1CL�E�!�č�3�֕�K[�0�+�G� %%!�H�F-hD���y�8bU�B5);!�dI/lX��X��ıyjt xI �!�D͊њ�ҧ%�sc���! �!��
 �Iz�MN����i���MY!�0sY �ф� �z�@�b�ƞd7!��d��X�(�!U%���R�Bg�!���0����� �.\""�ԁr��C䉠>���3%�W�F���e�?VFC��(_ƹҧ���v�t�#Q�˧��B�ɯH�zY�'�ץFVJ�b֝��B�I2jݦ5!pJ	%&I�H��һ��B�@�NVR�@ L0㣞$��=��'u��M�;P�'fG;�H�'r�k���|�1	�Z�2�yr����$y4L��afe���>�y�ϚWS��7#& �:��1�yo�$:�R|�Z-!� ����yN?i�<��(\�D�nH�f(X�y�'�2��i{`"�9�� �T��yB�͜e�,Y#Ç�$�pq�b��yb(�Q4�Ԉ^��Xly1���y2)�(K�fG���D��s-�y��
�]y\e��!��h��T=�y�`�*j7����l�j��e��y ���Ȩ����^�dA���y���0P4uC#�� VIЃ�D5�yB^�N�F���@�p���iC��y�$��O�L��E�Μc�y�s	�yүD�dļ!�dj��X���S��L�y��=�����|��$�B 	��y�dN/f摸e��:{�q�򭑭�y2DT�,�R蛺)'��� L��y��YR�*�H�"�v8���4�yr��	�F���K�o� Us�̖�y���U�h��O��|�\��R@���y��	�&v����\�r4����Z=�y2I��o(杀��"m�ƙH�چ�y��
�`��q��bܘQ8��	�y�Q��1"O��H�%�����y2(L�X|��JBC9N�����mė�yR"���V���_[��$̎�ybO�eޔ�5j�&(sR���S��y2�Y�R��:BM� �d�Kt���yba�V� �"p�ˬGҰ�j��J��y"�M2B� ��@��iA�H����/�y��Ɉ0����3���54`Q��P#�y�%*��t��Y$��)��͈�y
� D���B�Kz����p�T;r"O�Z&�0-���P鞗o�,��"O }���}��� ��Q����W"O�\�q��(D�����w��E"Oʠ�䯗�� �#7!DV���"O�Y�s�W�Nfh�����>*&"O%����q{��S���$D8h�6"O�ա�����e ʕ8#B`R�"O`���#2)�}k�,v��cA"O$q��*li2�K'lh�\����y�n�2f����%@m�9@�П�y"��d�����$�pTcB ���y�@V�.$xh�Y�s�J����yRH�;��e0!�;3�}C����y�J�'
	Н�!G�@r���D��y��o�ڳ��"1��1��(���y��=qL�c0�_%�>��@$��yr�Ɣ�^�hdȜ#����e�&�y"�/+X,io�p�t��H@��yҫF�9�q�Ҿ~u���	�!�yR�H�g$�C��R�w���dg��y#�?�|L�V���&!9
����yR��	i�tS���6zB���Ǖ��yB` /ZS��)%�ě1�1���4�y��9KIҥ�'��<$5ڽ�����y�� �Ʊ���Ѿs��bDE��yBe֯*0�%Y��\(�u!���y	�*[�֡�D��#N6��9b� �~b�)ڧtZ�`�E�"�Iҵ)��~�P��=9������A�NDf��3M�3�+!%����R�t�8}i���|.=��Ɩ-!�d��� ӃǍSQZ��A�@8!�QPd��P`��S�PKR#n!�D�;B,�LǪG� ���U�!��=��Ȁ�[(������q�!��-�ASbə4������;�!�D�~����u)(�ڤ��a��!�DR�d�̌ "��x��#�b��!��.�N�RH�R�����L��!�$v�i��MH�;�@ȑ�O�	m�!��3d
.��߽|��H�CC�B�!�D�8a����׬�Ш:em�,F�!�D�C#���e ˶c�p 6�[�Z�!�$+f�����3|�G�8
��*�S�OZ|�1��t>��n�D#Fy�
�'�m�T�9S�<��敕D��̳
�'�N h����{-2E���8*c
�'*�`cM��G�zd�G��2&��S
�'݀�c��)D	�	@�2ŀ���$+�r��(�x�9��E�(,(AQ""O:I�3��0�F\��₈{��F"O�˰���c�4��p�v�
 "O�����L|
��1�8X�P�"O�����2A����M;���Ж�M����ú>]�0�U'@�lN���$D���'GR�݂���R�t����'�d3�Sܧl���M�P�,�bΕ�|�XL�ȓah8{�H
k���S"L�����ȓt����p�ƥ��I�D솴e����<�* {�팈��x1�@������X��0iT+�R�:Ԯ�0( .q��	�I֨#<I���]��I6�űM��В5��_�<)�bص#@x�HS/YIx���	UyB<w���Ӟ|��)�Xo|�9�BR5F��Icҩ.I�!�� �� S�[%:͊�2�iĢ1�
�zF�d�z���C�G� Q�N�����D��UG�+D��)�(��ؽ��Y�mz� G�.D�P87��&��M��-�0m�k"c.D��HU�N+b�D�	�Ɨi ढ1m0D�,A�с;~�j6�%4w��f*OZ�i��R鄘sc�0/���t"O�)z���Q#�t�&��&�q��"OTLɆ'7B`~	砗(WiAu"O�yI炙ȩ5b�w$iAG"O��x�h��C�K��A�$*�"OR�R���-&��ka!�!�R���"O�m;j_9�܄����-?�<ĒB"O��g�$
�f���F�-x� ���"OV�c�jD�y���s"����@&"O�DC�l^�/R,!�%"۱8��Qr�"OL���~�T�aR��1,�����'#!��%J�ҹ)U,Y &�hi��	�!��	�AT��l�3	�n����v�!�D��0H(�S�G?,��ۑ��Nz!�77h��ǬR�N�~:�B(�!���$&��+��yY�a�Y�s!��^%X� ��S5x�`p����V!��*A�R���Rp$�x�C8)F!���1#
���`y���(��ךW�dB�I/Q�~���fՈ�¸ʶK�(�NB��0w��$ N��h���ϐ|����hO�>)0Sd_8e>2a
ɺw��Xe@.�O����5�M;y?��h�A�7m��ȓ=��9�?|�2���ȓ|�p)R�f�(\����M���JX�hC:�����ǁQe���x���hp�����k�M�1��Ia̓=9P@��6|�t`ۡL�)z܆�V3R�fж�*@���ӄ	�����ܛ�S�a� �z�J�Mn̔�ȓgV��	�-!��vAۊ���Ol�=�������`�B�5(v#�]�<Y&P�v���	aę=1�Vū��]�<�%$ɫ�də�K���rY{#���<�*���L]�u�ڿTtNȋuIU@�'��?��yz}3G��OފU[�>D��"SD�h'~e)�.^*4�hU��C���F{���_=s��QCu�U:"8��S�[�lN!�$���֐p
H�k��xc�Ӑ$!�$N��=
��@$p1ˤ��z��	h��H����-
��y��n7�!�v"O��rPi�xr,I�l( $�"O�X#2��<����	.0�#"OHM�fՠD� +�B �=�L��"O�6�N�&��;��Y>Ӑ�"O܅i %	{~�C5l�JWPC"OPʗ/Ɯ3'*����M�sT�Љ�"On!c�`��pHx����ZS(�b`"O�#%���d/��m4LJ�H!�"O�MҡI^?���0F���N8�&"O��{4C�h�8��=��"O@,��-��N-�DIH�X���S�"O��b �Ԋ  �T�a�ƹb���N�<I��_,��x���R24���b��K�<1�}hB�#���9/R�Җ�_P�<@��>���@��;I����kQ�<����#�����X�3� �O�<��ʛ�Z�����Ψ��Pw�d�<� m��j�:a>&	ۓ�c!ƍ�"Odth�/3�P��A+܁3
�ػS"O�̒2̅�Jr�Ջ�»2�B��"O&H�A�9%�B��
	w -��"O�HFȏ	 ��8&�Z��A`�	F���i��1� DҲ�!�����	 ]�!�dǋn�Ҁc���8A�~b4a��"O`���+@6�u�cD�ߒ�K��y����^��S@E(!*���'���yb�]�"�d�'+��r�y�Wo��yb�GP��DcQ�4���b�-�y��\e�ᙦ'ŗ~=0�I"���y�΂�z[��Ҁ�$qU �k!E���yB���.�Y��탻j�:]Y���y2č ����rW	�<�A���y�F�\��<xw�ðG!���B��y�R�إS&��Ȑ�A���yr'= :���I[;|�b��yB W0R� Kb.M�)��!�GH�y�JIDz14A��~T�ȃ�y�H�6��}
g)Y)�s�F���yb�Nb�|b@v8`���ylFL��H�V�6��`'�,�y�W��*d(s  [��AW(�y���&���"j���zqB��̞�yr"�
SG`��#��f�8TLI`�<1�oqP��`��ˁR�f�iv	�M�<�``��3}@��f��@��R��M_�<aB�ya7�s`�i"CH�AJ���2��t��;|�[�mޅ>ȓ_��<�3$�5$�p�YL��~��T�ȓ�4d8��T��Ixģӽ��m��\���J��''�r ���:@�hD��JB�$̭ k�4�(ŵzhZ �ȓD��x��b��[�
dC��ȓc���H�p/ZQ�ABY ά�ȓf�,`[�@�6WU& �6͹-|�!�ȓJ���q硆"&δu:&d��V�Đ��F a�Cc�,A�6�`�Δ�$5<�ȓ?�V���n�1�$	�	����C��A9���h�VY���S�+�̤�ȓ'��m(�Nަc�&���A�[�L�����ـ6D*hsj�27�DTK�AZb�<I����6a5�[2��]�,�v�<�U-Ørb�����Y�8 !	�^�<����M!������+S�U�%Z�<i�e3$��ts�A[)��4�HZX�<q�a��J�*p�c��%��:eόi�<Y�ˇ:p�aB�L�!Є���M�j�<��hX��n�*�E�a�ޜ*lD|�<� %�f$jj��__��{��\�<�!�.~ap�k��Vp��j�Y�<1$fU�^I�e���Y�p�v��'DM�<م�O�z��ǀ7n�����E�<P���(ǆi�&��4��1�� �C�<qԥ|����̖!fw���$Rv�<�A��2�x��h�c�����X�<�`��(���P�E1XB�)��c�X�<�i�7�<��a‸{HдeWT�<�E�1�}2��_����V�O�<a�lGt�X�ŕ	+�XT�@/�G�<IaǲT�ȸ���C:ӂ
���E�<��I�OO����%AzX��P~�<��C�ۂ�(�%��#��mIT�{�<� .� �+���he��WKS�X+'"Ox1��KIn ���!*�',B�!qS"O��*�+��g�X��G6++�-b�"O0��⊌$�=�d���iA"Ol[��?VXb���&�$66��2"O�A�mQ�]�)M�m��B �>�!�d=>Z�qN�2~��py�Z?}\!�D�#�`��Rl��B�����C+\P!�d�.qZ0��HE�[�@pj�V�?6!��J�?����&��%�Xy$�L�.*!�$W�∹3A(+��9��ܦ !�$Q
A|��p��&!���c�Ǆ!��֚Q;E.�B����!Y#!�D��K�Ɗ@���@,Y!���0d��ؐ��R�4��xH��U"�!�Ӕߢ�ƅ�Rt�r@E�.-w!�䆹W�@4��e�zM
Up*�`l!�$�~9�������b/\i�j[$yh!��ѹW��X�D. @#�i2iQ#K!�d�@*M�&�P>-��Q�NW 
1!�$��V�X�k�o�<b����ؙ'!�Dϭ����k�$�t�v�	!�d��6�Ѐ I�f��<�iV�%*!�Ċ�S�4YҡŀM�Duا(��R�!��[�8Y�ɖC��i��@0g薵&M!���VONA��8t��P�u爡qC!�$Z1,���@kmb���+5!�Dܗ[�|Uh��#O���/xO!��F�Q�rD�ud˵e� ��ƦFD!��]y")Q�-
�%|h(H�ʈ�3=!�\�Y��h�턮;g>U�Dǐ�!򤚼0x����j]#+�\!�ǙMe!�V�bz�uˀ�¬}8���Gғf5!�DV�\�@lS���"��E$��"�!�D[m��p��ίJ��IjD,R#4�!�D�J{r��LYP��}Q���!��T>)���:����X5!�d��VNQ��K�' $	"j��z�!��K5F`0!m'f�8�wBM'!��A�t`Y��;b`jq�۶�!�D�j��!�'�N�(����!�8Gh̙�l]�p�ʙ1��œ1�!��>AS�8`�:h�blxu�9	�!�$���H��]>'�С҅��!�bݎ��&��(c��E�n!��/^�Y��!��;$+h�!��L���� �	�88	����,�!�D��/H�,�-8zp��JD�o�!�䈕��0�$�B�%��X�S<u�!�ǞIQ�M�����'aD�Pn,|�!��X���f�ݟ+X�چ�џM�!��1�)����BK J�F�c�"OD}+�4$BHCq!�8�h��1"Ol�9f@ϲ��ԩ�@ r��A"O
��'�8|�H����J�h�"OȄ/��80�E�Zv��o0�!��	�(��9"�ӭ$0*�$��O�!�Q�Lxt��fG�s�|"CMY a�!��|{�s�@E�a�vI����p�!򤋞
Ș� Ö(2��t�7�^	�!�[�j�h���	o,V�� ��,:!�dD-� ��J�	 q���r�!���:+TTK�O�Y�`ɰ�M�S�!���|5LHdO�#�&$Y���!�� ����q�ظV	Z�N����t"O��*�&�	7V�T�EW�i "O�=X��� '��E�ӊ�O�Șt"Oօ�U��lf�)5�X9z�d�u"O�h�*��'v��[L�L��Ȁ�"O���c�M� `^@�sDɉm j	iV"O~\)�(M�<a�r�b�`���"OXc�w:�$�c����y�"O,d��`V?1!�	�BP�[T2	%"O�h�dY�dhʡ�� ǹ=���	�'I�%q'E�,���� @A�',h�Q�l�h�"u!�yx�"�'�d�¥ꉴE2iP��`��
�'���bC��$ h:`%���	�'��h�@t�-���V�h��'� �� �_�h!uŖ:#����'i$�P&:����Q9�<��
�'�T����.�PC�!a���
�'g�|����|Xp\�C�Y�J(֠�'A{Ã/mj�Q6�<�� �'ڗ��q��� 8%,R
�'�]`e�]";E\��B9-�"�	�'�$Ԑ!�W���h�--j�,��'x���w�I�XfȁY�+��T�r�'ٺ]�2�]�[f��a �7V �"�'��SȖ�G��t!�POA "�'�da�B��(��Qg�"D���
�'rbx�q�	`ܦ���<���
�'������#�)��)�.1��'
�4��	F1�p8sFG&�K�'��TH��Ư7���s
U<�Z��'�ν!��tt���mY .�L���'54`mX+�����6r�> ��'\��Q��,30L��%ߊl� q�'��!�D�F�Ja�H��W�/5Li��'�l��Y86$<3�D�-/^��	�'�2YK���|���f�s�&H��'#l�$%Ό,�8`FLÇ6ZE��'�>����W�Q������,yJ� ����Op��0§�
�ۣDZ:<|��
Г6�T�'�2�'P���O|�J%�u����"j������.28HC䉺E�R�͗]7�(�GeD�BC�I==Bpiu��	���Q/�	,�(C�	�9&�z�@ӊ͌ �F-��}"C�ɜ=ٺ=bq�Nt��OǴ)��B䉮a��h9R-��R����'��l��?A��iO�B`�c�b]<���"I$E�S�h&��gܓe�F�PT,�P��X���	9�ȓd�m��
�GƠ���5�Ň�8��%�g��#ae� F.�&kyR0�ȓE�>��JU$8���M�O�xT�ȓ�=�fÓ >̱2��rWb��ȓV���8E��G���Y��jJ���T�����؞�i�@\<"EL��?�ӓ^^��5��5�
-q��ȓ\� Ȑq@� x	p���>���ȓ`:���Ț '�\� BJ/M,��bu�pv�Q�3�h��4G�)��(�ȓ���RE�Y�8<3�l�4����>�l���H7�DQ+c-��PӤ��FL���"�Ё�Z���<�'����Э�0@�0h)���)`�C�ɮZ\"�[���7�b�1��[x TC�	�	!	��d�>�)Q�k�tC�)� dX���ȹV$A�q�ʶ�̲�"O�|���YT= ������ʵ"O�`��G�_��)�C�/����f"O2}��j�uN��d��={�4�C"OT�[���`
�[�Ⰼ�Q�^J�<�!�]mAP���WrNS�TE�<��oՕ;
v}(�/�e4�]����|�<�w�.{��L�%��<H���s�d�p�<Y�e�\��9�d��?lV|k���m�<�A��k�z�CF����n,#e �O���,��@>y��%F4?J�=�"��Y�h�"E1D��*穕/L���k1�[13���P5D��P[���0,�4[U�HQa�0z�,C��/n�@X�\�{̼��C�.O�B�I&���(��t]�M!�,5�B䉃|R,�pn��!�Y����ra�C��	9�����O� #�œŮڙ'^⟬�	D>e�`�z��D�Dم=m�\ۀ.1D�4³�R���E�w�ظ�ĲRD$D��I�J��(򖨪��*2D PQl!D�$�u�� eU�2\���
���y"�2v^�Ԡ$��O~5+�J��yR���%v��X�H?2��HEj�2�y�GG�6��qCNY��q�gDP���hOq�lI�!D� U|� ��e���C�"O�dpQ
@p:�X���G+P�-"3"O$"�+�\
DF�0���X�"O�UB��X�R��ɂ�D��]��<��"Ol) �l�)f����������X�"Of�c�J�1'¬�T�Z	
�~� c"OR�����бo�Ќ��Y�xD{��N�R����Bo�L���9��]�!��>Q����Մ��fy섂�KڂZ!��S���:ce�qL�A�j��!�$� V��ѐ�Ί#$:"�7��7!�$�1d��VC��<�����U�Q!� k��``N���
y��־�!�D�g�.Ӏ+�)"�`��A�P+�2�)�'E]0����@�j�,�#�%Q����'2��⥝�'��ccOW+6!X���'U�K7�0=B�$C9����'�TMec�X��9� �95�v�!�'TV ��e�0b���۳d�+.�����'�r,a�"Jb@H�83	Y�z���'|��.@�T��D�c8n��'���+s���W����U�9#&�
�'�z�IQ�Y�r���3���7�zi�'/��W!U�v�PLE꜁k�� A�'`L�HA���>d���#{F�l��'�	2e�g�5�H4��GaU��y̋&/���hH�Bj�Y�����yr��6N�F I��Ǩ?�I�G��?���'J��i�^}�� 5Z���t!\k�<A�D< O�-#Rjͫue^��7D�c�<9�����n�*�o�L���&g�G�<Y3��2[�8�	�5P}NdZ�A�<��B�q��tG(c{"xB  {�<���A���	�,�����%�x�<Q�  �-�$������r�(��q�<����bl�xp���9��4��E�n�<3�Ͽ�J�2��-C�����j�<qe����!׭5jK�bK	f�<�"��;4j���¸iJ��V��V�<�䪙x�Hu��1��ݺ�.T\�<� ��" FP�9�Ty�5l��w�b@ Q"O&��$�� �YzKF�(��)y�"O�|��Oլ��Lq������Q"O�$22�ݭn����� г/D��J"O@಄�>�<pzr��?"��t"!"O.��P�̅#
����ŋ:�R�a�"On�k1c�0hOh�rg�<(��(1"O�� ��V`��&�\��"O���dl0%ۗNu6�iY!"O��h�0o�,+��ӏ ���"O��"�L�#h"��K̠X��YV"O�5c�PE��H{j^/Y�Hc�"O�pxl[u�dhPF�Q�*Ժ�"O|,R���o�4���G�����"O�u�D��-�@-	UB;8h��A"O�`Z�aEK
��D���3�
r���O���2���"!o��5v�1���ص�N���%��i88����N\��m��P��Ș��53\
�����X��!��y�t�D�֛	�B�R��*)q�-��:j8��ƀ�<d�d
�.'zj�l��'���Q�K�2M����j3r��JP�!��h��D�93�oO�d��0�?�-O#~��XK����	t������H�<Ib��Eh�Q����B$4���j�<�צ�y©��͇�l�jۤ�EQ�<�ȃ1B���u*�1��ݪqL�X�<9� \$Ei0�y8�z���V�<�T'W�>
ʵ���B/lI9QGJ~�<�C�U
����A�M�z��$�TO���?���ň�b��cO	�T�A�'KE;�&��"O�i�D��
.������[�]��Ma�"O�$ѵ�̥d����H�A����"O�-���Ȁs�J�s2�89j�"O�!ff��.���EC
Eiy��"OΌ�U#I�_���C�֒C3teA�"OV�J�"�"%��<[Ċз	-�`f"OR8T�6Ÿ�Z ��2�P� "O�Ak��K�|A�D���R�D@!�"Oܜ���܉���Cd�$�g"O�H����(u�\�s�E�vn	��"O��ë]����b��N��Ʌ"O�%-R)%=H%���@Y���;�"O�9�qN)q�9Pˋ'0l�aA"O� �%�2�-Ѕ�];�N�U�|R�'�az"'�,ph�V�����p����yҤ�$/VP�Q��&�|+����y�-�I�d[�E({�YY'�;�yR�J�{������ku6]oJ��y�g�JN���s!ɏ]n��S�	ŵ�y���25V�1�B� \NZeb�-�y�AX�4tZ\p%��#D�ROF�䓥0>	D�7���Qև�c�x|�uJ{�<W!�{j�)v��	o`���'Xs�<��'?i�!�4+�-	P�@ K
{�<Q'�v	��(S�|w�(H�u�<�se��D��p� [������J�<i���:̜D�A@Rlơ��A�<Q C�kG��P�gV=Byv��`�	~�<�4IהX���Ygė6k�B=c��{�<iH��	&����C�6F)�y���t�<���I�X��h��m�R�ҐH!+ Z�<qA�+K��X�Nź��a((�q�<a�Yƒ�w�
�bڌ��Uw�<� ���	\y���z��g�2%��"O0"�d�n	���GMkJ��v"O0Aڂ(f�ɲ��>DёR"OF�DE�6u&hS��R�Ftb)yw"O��c�/Q� ���k,L-
�q�c"O�H���!���Q�/�����"O��X��
�>�*M1ʃ)��S�"O��8 �0/T�J��E7t�Hp7P�,��ɴ]�J�Ƈ4�l�сF!��C�ɉYU��{����pe	c��C�I�O���XbH"AX�W�.6^zC���,��� ڼu9�����̄.��B�I�6��qq`��#d�9`l�,_��B�ɂd���c���OT�����"Y)����g�(*�����ćU�%�h��8D�,ʄm�-�:���KR�2�` ��5D������2S#2l)u+R/]���hp�&D�\���{<q�&!\�?3����$D���hG<얥&�@Y��$D���  �w(��#,V��(6 !D����M��e�`�q@�, ���
?D����?k�l�!6I�-�ހ�/D����)<(Ķ ;�KH�}�l���.D�X&�ٔP����c�)
�����-D�<;a�2բ|�oF�R|xz��*D���U���	yn�H (EBh��b@,D����Q�U$���- �A=�}Jm4D�<Ah�4i�~,��X�Z-���&�O��d�i�B�L��@����R&�	�ȓA��0��N_8]X0�;�C�,��ԄȓNDzz��C58q$�;p�~U��+�Z(є�?$��(��7hm*U�ȓit䉻v���Qx�����X5���ȓ
�]��,B�+��3E��2cؐ�ȓ:RƸ�4o�l�Y��g�� �����I����I�<�6���p��(hf��We�B��I�<��L�$����g���W��l"�E]�<1U�ڔ~c�݁�n�&R��Ѣ.�\�<)�a�V�&0�Ԉ�1o)�I9��m�<�EgK2p/�����2A��!��u�<!�CWd��L��'�08����&�q�<��Z���pht�N$j�b�B	�Ex���'��Pő�:X����gO.Z�^ #�'{Z���ǉ��(������W<$��'X�y�tCD��\Rd�I�b��'���蟶9��T)�([�x���'Le�e�RD�PX�cC�Ԩ�'2�����t�U�GJ��R���'4D I�A�a*�X�%�$E�Ɲ��L�H���KP��z��W!d��݇ȓ�xq�s��ee�ݐW HqX$��:�X�2�#�~$�V���{b�Є��.� �,���S �	�t@��U����h�Ly�mS�h�`�ȓb�EJ�&�U<��=��ȓ	C�=
��I�v�*'�@�����ȓ�Tإ��u�TM�@�d& |�����c��	k����W��z���$��,a�R�n�"m�v��H����Z&�;'W�d��ʔN&M�JЕ'�a~�Iϛw����O?`ϖi�c昚�y�g�3e,à\�OjL��3d�?�yr�Y��lk�A:���q�@��y�-\'A& ��b��2�b\y��E	��d�Oj⟢|� Ɓ��d/y�@�RԤ�-�,*�"ONR@��,4�3��CY{�	�""O��cT!>�arD��Ef��"O� �� ��%���`,�o�����"O����@1NڒD�kg�`�X"O�x���+)V��L.`�\�R�"O���S��2))�	�> � x��D>ړ��D�3xX��ڄt���yA F�Y4!�>桠�
�W��p��ˎf!�d�^n�k�&�?U�j�Т� �.���'�a~��J)C��أ&�� E<�+V؁�yBc�%f�ډ���K�S?40q��ݷ�y�չ&�
<`T���PӞ1걉��yb(@�1���`)]�EL �с�A��hO*��I��~�5	��	������!�d�
8�K0�D�cLa�v���!��8d��L`r��.�^9�p&��!�D��L��֪M�v�.T�4��+]~!�M�!���RQ�Eln���eC�/�!��D��8"�i̝Wax�@�ݸ
n!��[�_�	i��K�riq�8 �Ox�=���
5���v�d�mX�@�VxA "O���2�������b'.�ȷ"O`U{��OB�E�F\��R"Od��¢�8�U�-Q���ʇ"O�-�Հ�%
��d���VF���"OYZw�Ƚ&��#�f�*T��I�"OD�����L�qY���_�D�#"O�s��Q�<��l�7P3`Ⱝ��"Od�q�O1.2-�W�-OB>��G"O�}�g �)����_%z�c�"O愻$i*aP�¡N�!rb��"O"���F��>Jb�rB>8S�la�"Ox�ke���U��p�a��w�8�"O�q�<#VV*�O���y�"ObX�G�E�2x���Ņ-�`a�a"O�V����������o�` �"O�XfNԸa�X5 ��.��Ы�"O���+~,����n�1a����"O�IQ��>K~d�Rc�L��Tz"OX �@�0 H���ޜU�r�C�"O"�xw�C�-˶���6�4%��"O�(S��AD2Re�ٽd��0�"O��A"]�h�� 9��)FBE�"O�!�nS�9	��B���8�my�"O���+�zh�#�oTA H)k&"O�S3���=��������C
2��"Oƭr2�٬'/h�p%�#e�� ��"Op4�@/�-[���A��%Ҝ�
�"O�S�R���a��D�1"OгũW� ��|:��σD��h��"O��Yd�����w��0�.��"Ot�;�Ǉ�1�
̀���?Y����B"O���FA)栰PL�Ny��&"O숑d�!w$��q`X�5[$���"O���U(۹l7�0&m�}<�Ix�"O��rf��,�OKֱ�r"O��p���Lq�3���f5�tXV"O��rc�l۲	r �C�Y2lQ8�"O*�[�o�s YKi�0"2mJ"O\�ȴ�
��@��f��>�#7"O�Z���+e&"I���
����v"O$���n�<1Q�1Q��Xjt"O�*�g��t�f	;�#�<w@@�d"O� Q��g�V�� ��A_�qY�"OF,��Aڲx����g�*+"�x�"O��9惞:��P1��@��^��"O>03f+�*m`B}��Ř��D7� D����W/����H�"?l�I�m"D�4cU��8H5�C�XÚk-D���2녫b.���@N�;W���ɴ�*D�P��E��y;D.�9rFIե(D�����ptj��]��%ʜ�#!�dԺk~ )�@�·dFN�HQAQ=}�!�I����A��92J0ء@I�-�!�d�o���W�ǿo� ʗJ��!�$D2J�*)F����R��!�K�4�f����W�=�f�r�	�!�D	�F)���	�w���8�LD/n�!򄜶�n-�W�G�G��D`r�˱�!��Ly@.���JX'Wm�(�Q�[l!��"�R�dؠQ\��;b�]�!��@j��@�L^!ONH��5�Y�[{!�(	���%4���� {�!�M�F�xQBCމu�n1��x]!�ĔJ��h�#:���#�V'Z1!�dM�kҌ��.L3_��-`�&�#!��?�P��D�c���Q�E &!�1��+Zo�n�бNR�!��>�:1P��Ύ&R��Q�l�-�!�D�(���4��'.�m�Pl��X�!��s�p�D��L)80�Ʀ�!򤛲U*.�"�.u��x���=MX�C�I1.$�أt�@	aw�5cBØ�_��C�Ii|�=j��Ԍ<�!�'"�?�C�I�E����u�x���߲V��C�I�u �yQa&�|�F�����1U�B䉫!_���.qL��Ǉ�dxrB䉊H�
t�E��<e:حkV@�>�lB䉌O�.�
��XS~ĽK���oJ�C�	5rȍx7 P��^]sc�˷Nr�C�-c2J��I�B�2�Y� �&^�tC�I�='b������N�X�Z����q�RC䉙\���&	N�$J]ʑ� &2fC�I}*B1�#�D��x��BU�JjB��
zT��%��[�P��"O�RN�2?��$�%�7mD���"O��s�jֆt�Y�'�E�j��b"O� +�
���`��@
�&hXM:�"Ob�0aL�-���ToT�R*t��"O�A�Ҋy$�`QTI�~b\�w"O2i#���B���(�G�>B�]R�"OJ��_�2�p 4FK�uX���"O�!�P�ZR�=q��R��y�g"O�9��	�t�����!z�l�؆"O�|�s�]�|V�G:N�
��"O�p`�IY�}R鐧�A���$"O��0J�:o��a�GVi���2"O� ��jS�+Č������`��As"O@�Ґ$B7b)�5�0���'���*2�'�'�B��>!a�X�<(�0�Y�1~<2E
�x�<�SF��j��Q��2���#�u�<��	&yx@��(Գ+O����V�<yf
��|�,�EN�/�@!�mSO�<��!K:v��erC���[�x��E��D�<��J�y��R�٩-�\���
@�<�J*wr=P!J�;�v)��~�<Qs�Xf�}�Ɂ;U+<񨇅�y�<� ��+Tc
������m �=���s"O\�8t��9=�ᰱ&�,<&P�k�"O�qq�ZB���AS�=�$"O�5B�,�S�~teɌ*.؄��"O|�����:S�5�v�K���2"Oh4롊@�Lj%H�r��3"Ot9H$�ˤ$δ`
Pi�/L��څ"O�8�'����D�"�K'�( �Q"O����!]7�QÇI�R�"O�)2�Ĝ�^��5���&K
�ٓ"O�бc�����F�_`����"O&��BÏ�g��u�Ȑ�A6%��"O���5��1���皱w����"O^�sCoY�Yz��YUg��HFY�"Oj��f��a�f�a��Q,�!�"OX��"ْ|�� ���*G;ؐ1�"O.9�ǖ�p�ū0��0���"Or)	5-G�tMq�%��G"O.�;5̞J�"���ܠ)i�"OԽSĭ�=<�����X (�6"OT%��d�CV�S�쌸j�= �"O&���Ϙ[1���j��y����"O�|Ҁ�h��*�X���
%"O��Ti���T����[�A t"O>���_T� G,�&��II%"O|�ja䁐j ���ʇ�D�j	y�"O��2F�ֆg�Ȥx2G�0�(�Q"O��AF���_f�ak�*4EJ�!�"O(,�*:&�D��P:
�@X$"Or�+����#M"�8vcAI�zEr"O̴8�O$P������1]��Rw"OtU2i��ZR�D���A}�zD�"O��ҋH�[��:��T�Hqc�"O�qPP��=>ߘ@A��)�N	��"O�t"F'O#w��[E��y��D�3"O���DҤSB�i&.�dv���"O,q�
�*-j񀃂CYj�q��"O���T� `b6�[�yp��ۓ"Ov�"V)��.p�5Z�Ŗa!zb"O`ui#\{&�k㪈�bRR��"O���cDJ�^��#�g�3@E���"O֔[w�=ԁ*cF��WAưK�"O�ЛhW-�e�d>6�D�'"OХYPV"\y��r霅"��B�"O��TeF@�\H���Ão?���""O����@�"9&DrV�3
���&"O�Y�Ӌ�^�P�����&в5rR"Oެ��+�,5V`C4�)�d� �"O4!�M (�j��/P<�8���"O�A	uF	�y�x�2,�"n����q"OR����@�X�	S� ��\��"Ob�zV�I_V��������7"O6�� �$eEV����J�^� "O
��C
�Fp�`�Mӓv�p|y@"O��ѐ@�Y'�Չ��Q�KEr!��"OʙӲcZ49|�T��K6_�%R�"O�țB��*R���pNI[Z|1�"O$J2m=X�4I��qR�T�p"OD��4�ɹ��E�m�6:H�� "Oȩ�6�B��|i���J�2��0"O���"N�ܔ�eB�)HՒ��V"O�9�%N�J���c��9�f}i�"O�$3ǅU�c���p��	/�.g"O�a�G����9HT�#j���&"O� F0�m�i.�h��_T�@aI�"O�tP�C�ď�A�Y�e"O��b�.J�=��+a䛡5qP""O,,R�J��-����0K1��b&"O0� ���Gr=���m��PX�"O� Cs���;pd���Y|@D�#"O.�c�%{�xaS5�� �U��"O�Ē�,�Mv���!$A��"O|D��,i+ !��w�ڨE"O5��$[�+䦑*ԏ$d?���"O���@B$+��Mx��@�A��� "O���H&?�05� �(8+F��"On��D�ǥB'@����:z�H�"OHZ�E�m�HX�H��Q�	��"O�fG9	��9�F�=.���"O�Eu�G,Az
�d�@/��0�"O�E��lQ 4�N"� �`��"O�I�G4B�<��!մ���"Ot�Д/U-$��]Ɂ!�:~$"Ov%: 	M�|�x�!���**�J!p"O�𠲨�q�����7�8 �p"O0HǮN =��b��պ
�v�"OZ%{T,՛5(��rƄ�@k�T��"O� ׏�!z��c%�A>���"O��B�a�(l[t=�ă-(2�Tau"O���� ~ִ;�Y�!�zR"OV�X0%��ab�-9�]8;/����"Oδ�T�5 �jG��HoJͣw"O.0��#u^�dn�"md|�q�"O���u�_�BUR����	|X�0"O�%�n! �u�q�%hV0Ա6"O49S`Ç�	�&��_C4X�"O疴�B��IװZY�a�"O^�S��2-�Xq0��H�=�%"O� �g�X!Ct���65�Zt"O�1g�-�4�� ��.(�"O�x�ĦC���
Jt��%"Ob-�$I�3TJX(p�I���C�"O�D#�# �*Q�G$��t�"O ���	;v@-Pn�����"O���edǣW���Ҍ�E��B�"O�!��ںH�ܳU�'"�m�"O��!"M�p�pykSǮD-�U"O
0�4�{�Bo�L�"O�Q8 ��	0���j�m_�A�b�H"O��X�W� '���$7M(�"O�i�0g�&@#e�ˢV�+"O~Y�0�W��)�U���|��=�A�|"�'g���1�%'��	�ΕMff1�	�':���qȕ&F:����:V�$�k	�'KP�7䆪Ob�4���0R��]��'��SSL��rN0'��K�.�R
�'s�ى5��(s�<��Aqx$�	�'���� �*.p�]rT.�7C�5 �'r���r���@Ϻ�#�/�?���K>�
�c��ܣ�K֎��FEY�[ ��3>��U�ݽ����̀) ���ȓ`��I��1m�j�"B�?u�J��ȓe=�-�$�?*�Mqf�>>��!��p��Y��#<U4���ȱ� ��W���b�<]Ԅi���)U,���Ed���d�Z��yi��ܧ�d �ȓ���Z�@�q?:$�DdԊm��(�ȓ\�" v��c���@�炬r2���S�? "�P�'Y������#Ϛ=��Ī�"O�	��ْ���RF�K�/C��t"O:UZfm��n08�� �v6���s"O�B0�K6�٠�^4"�3�"O�pG�W�Q���+Q���I5��"O�����;"����KׅxX$2�"OȽ�#@әH�N�P��]k�Yk "O�3h�(0hY ���<<�qzV"OB��&n�'�rdQ4aW�h��d"O8�@�-a`�Ж��5-"@|ك"O�ap�H�7���vN� �U+�"OJ�3v�?42�ӊ�\�4��"O��P����a�ԧ	vø�r'"O�}Sw�F�x*�@� T�"w"O������:��1aۀ[R�e�"O��b���8�� ��^)6���"O�(�5��Z]2e�uo[z�@"�"O���u,A+.\������Ig`u1�'���q0�-�.ē�7 ƌ���	3D�(���9?��&�ۜ �e�1�1D��C��F4?�%$�s�1S���	�y�&M�.>�@XA�K�RD�rv�1�y2Ak �u��'\�N��@�B�Ɖ�y��I'B��kH�AT�ٳ!"�y���+@��X�k�&=�h�Cϐ��x¡]7Rp7�N:d
�Ea��&�!�&N�TPVa�� �)ai*`�!�DH7T�݋��X?�48�h��{\!�$D�f��)0P!�?m�<��)9A2!�NBw�#e�׏Bp�xҳ�SF&!��t�J��%kX�4Z֕!)��!�� �{�<�g��::jh���x���1Oj�P��O2v���I�o�0��"Ol�A�&�8{bp(�(,B�)(�"O"t끅��(���bK%K� ��R"O�|#��S![��@Xfg�@�N��"O���D
4(��`�����k��3"Ox�l� �qf#ة	�Ԥ��"OF,b���⎽��"��u
"O��JE��2�@�	ʦhQt"O0�����k9А�ԏK1.���"O>���Ρ�	��OE��m�"OKF�>���3�E�d
��K �L6�yR�Ɋ^^^�K�e�]��%
��y�a��xS�nR�b�3�cK��y�؉�TCw�}�2������y��V8bNw����_ �y­��l,�g�oi *!�L#�y��O�R�����jG�Pjp��ʁ�y�D�t��H6GR6��A�W'�y2�˕~��"���'��ţѥ9�yb
ڼg���X�
�	B�۠Dߎ�y䖌?*p4���ܜ_z��`�!�y�W�9����u'�+4V�� �@�y�%�0� �0ŏ�niq��U�y�4	���)q��H��,rɕ�y2�� ]���aJX�m=�q�v�C��y�՚Kb�|q��/\A�( ����H�<9��`����Ջ]D.�ȓreva��� �h�2���)Ȝ��6����Z6j��f�w`X��ȓ����`#.���Ĝt�8���iVʕ3D�ԖX+1� E��d�ȓn��U@��K� �G�G�����S�? �);s�ىR�FU��h��	%�Qȁ"O���iJ(ZX�$+�ߧf�!R�"OF�Q��z)N�[�k^�s�VQ��"O�Y�#�̋@_��j��
>a��b"OF��@��W�,Cb
Ee�����"OșdF.��<BlS1^�N�t"OܠPs%W:xh�%!�l� ��c�"OR�` �Z
	�H�s�I��r�,�I�"ORՒ ��k#��ZT#�^pbذ�"O �`]���yyС�:j ���"O�1��@	+l�@g��b����"OYW�O�R��yG�� �D�*C"O��� W�JB�����ԕQ���3v"O�p���)X�%J� P .�X��"O
L`�K&J�
ШP/Q'��j "Ox�U��1pT�MX�/W�&�F��"O�-���ݼ4P,�D��mwT8B�"O��ǫ�E� Ô ��[P�X"OH!�vj�36�b ��(ƩkCBI��"Ot�%̘�9s��²g�+jasA"O����^,sZ��� ���d"O���P._�fgi����H��"Otʂ��f��p��S:/e�&"O�-;��[�n�|�C��l��1��"O�8�"#\�m�ހ�oE�v�t���"O`����F�p�C��C����"O�1�j��������\N��)f"O�Y�cK!,=�e���\��}I%"O�`@�_h0`+w��Y����Q"O��ض�؇Q�D�чF�s� ܪu"Ol);&�� /��5)�̞���"O�m�%fL}��Gk�- R��"O��H���i(6	 ��O�<��1w"O�±�\1o��ɸ������`Q"O
F���w ���f�4���s "O2q��#Ǝh��I�4c�Fd�Ҕ"O������nX��9EKW�xӲHJ�"OX�U�Ӹs�b)`
�Ϩ�0P"O昂�e#6e��3cT*_�م"O��3�IF�F�T���Ѝi<|d�%"O��� ���U��4��"Q"
#P"O��F�c�����f�B�X�"O�-9��Q-aFH��l�J�:$ g"O�l����HHBv�օK֌�05"OE�����h���Sv��j�\̨�"O�Z���4�fu��/��\c�"OTU P�'������ Z�6x�t"O�9��9+���ňBKL}*�"OⰂ��+�1�3:�3�'���EF����,�P�(>�<��'�u:W�ȏmc�Р)X�;^4�[�'�F�SA��S�)s�!�=5��ɚ	�'xj�A�^�h�u�;+�4��	�'&�����+�$�H&e�>L���"�'ʄ�d�Դm�Xha�LB�Iun�x�'����K�~=�Y���A+^)�	�'�R�!Pj��5�ޘ*���:.�J���'+��o�Q�[�|TKa��U��'/���!�E�!�ry�'�Dd���'"��a�L�Vic�/� ,�|�
�'�.�T�UnUr����9�	�'�̫� R�r}��uGHuC	�'����d^�F̩��I/g'�ث�'���B�+82��X�)��Y�@�8��� �|�+JT}����٠m�င"OH�X�F�9�vMk��Ro�x�`"ON0	Ł�� ^��#DB|�|��"O֡����@���C+�:�Ӥ"O���c̥E�Z�׆Y'."O�`!��h]���2�\#"���V"O�ـ&/,I�M���,X*��a"O8�f�ɖ5�r9ZE	J+ބ��"O����0��gƟ<;����B"O>��. �ri"0����h��"O�9 ,��'���"c��8؈��D"O<�C���% �D��s���,�$�`�"O��KA��c���QE"�=	P��"O�Yr�oE��s!�J�
Yiu"Oy���X)oj� �7!�mި�Q"O��y�J�E��F"�o;�98f"OjX��f��U��k�斋 ��	�"O�����
c��J�.p8�"O�@CE�Q���@5�Q'89#$"O�9�u�V�+6�Xۥe�?i�!)"O����l��T����ì7�����"O�H�$I���y;&�����s"O���ă5�֘"@���v�r"Oށ�d.]�x=�D���!7��z�"O�l�ԗ.�2ԑV+��>�X@�@"O��X�*N-;3�k kB���:b"O����a?F�����D\Q�"O0���3uO,���.�Eh�"OT�5"�4&�dL�6G�w�Y��"OI�+\�ѷ ݣ0�
�i"O��3iD��IpT�N`n� jt"O�x%��[����Tm�.Y�"�"O�y�$�J3�T��NwT�i�"O4ɠ����LL�	V�*fj8I9�"O����xӨ�YCG>��� �	1D���g�Q�as�U2C�!_���"��<D���"�G�/y"�9ϕ=�t��ą5D�iF�6yjĳC�)Z�r�j4D��B�A��J�!I"K��E�α�4D�@��`A0I���`��Fm��%�d<D� � J߮*�ȸc�����i��9D��:�nC�~m��w��71oؑ�b7D��A�4��1F�Bs�U:sG3D�P�4mٻcì$�2'U�d��jq4D�4ɡ��)}�B�f�my��xw�0D�@���? ��\��E�'*p@ Hg�4D����BB��^�a1*A�B�>�2â%D�
G�ݫs�N��_9�8�K�o1D�8�p��zY�T�^)��Đ��-D��#��ӷ3�4���!��p�s�+D�D;�ʷ7͌My�΃-?h�,/D�hxv��<}P�ܩ�L9� �kD�,D�Љ�b��I�Ƙ�PF����U�D D����oU�)�T[�DI�E��UR��(D�`�¡H_�Xz�b�2p�\�J��<D�@Q2b�'��q)AJ��~  ��j;D�$���'.��1�u"��F �1%/8D�8[�
\f��ؔ B''��ca�5D��!�ʍ')�6\��!�N�Jp��I/D�TI��a��iP�D��>�:��(D�x�ꈿJ̀J�<Sg�X'�$D���an�)#��fG8.=*�s�"#D�Ђ�\q��蕦32�&��6D���	M�j#BmЦ��}_^���(D�� ��Y�A#n������GP8�a"O�)bQ�E01���j�CN~��Q"O%ꇋQ68�^̉�a^5i�� �"O���W�he�B�P	o��ܹB"O�5Sq��9R���H%����<D� +��L��t��ѧp�P��<D��s4sV]��O]0*�����&7D�`�1��1BN\�G\)&����J*D��8eFM<-ab-+�NZ�2�d!�)D��ūW�^�eGbR�l\,�;1�&D���c�	f (Q�5"�_j��� D���b ��&���r��0|Fc�"D�l{� %A���R3��#�J��>D�$
�hO�`��2�@��s������/D� ��85�PT҄拣L�ȉ8g&)D�����H�z>�)�/�4bU�A�'D�|Sb�:2�%��2P(4H!D����G��\f�L���0���4�,D�$�`�N `n�(T)F�*��̢��<D��y�%Q�(�9�G�sa.�q�<D��9�!դl�=x2Ƈ< ��k:D�$8�GB�\�ȼB�*
a޴�4D�i��Y��6N�o��@@�%D��C0J��=� �c��cN�QN!D�$I�$͇6>��3$R�/<R��#!D��Zplө�6�$�ĭ%�hQ�w+!D��c0$�>ɔ19vLC�3j���t!D�|@W��n�RM���b�(0 �=D�$��i�l�h43K#�q��<D��4�n(�UY)R� dx��>D�p�4(	��lx���Z���ҡ�;D�d!�-�d�L�����B�P!�7D��R1� �����?da�qs׀;LOH�@�7��34�XQ��A��sF���v�;D�L�A��)�  ���@�"��m�!'�IF���ON��XV�N.\�*��W�P!��'ŢMX����zd� ;��N�z��M�
�'��]��/p|d�A6���\_�,��'	T���Y�IdA&Є[�(�c�y��)�ӑF:���CZ�F=TX��M�-q C�I�k?$`�	K�LP�8��)9��C�	�IE�9�qL�|:lY��lC�ɸR�࣢G��e���{"�Y9�pC�ɭ�pYqU)�.�m���2Zd��'(1O?�	?gr�2�H���9����Y�JC�	�m�j��T�'S��UT$Ԙ�<�Ip��໔ϋ TTB5�
�;]��� 1D�T1�o	�t��؃��g���e:ʓi�xˎ�=���9��� K������y��]*v"�M�|�Y�с�
E��i�|FlA��&�1e�֙Hg�"��	I���,�ɯm�-�Ӄ�@����󄁹b��B�	 /�Q:�c��բ$��W|���u؟�i�����=�1�����)5�'D�(V�j�Hw��,Yt\�P`(D���U�^3��}PA/U	v�ڰ$&ʓ�hO�&Z�����X�X� (#��RB�	/\\�Aj�
Z$D6�Cb�ϭS�����.�DJ�L�
 D�92� ���u�!�R�ԤI�+"]:��4:�B"�}�'����+�!�&��'a��%�x�� �)D��(���~B4ق$��zl��E�&D�abΝ �|l���J�QMh�&�/D�8� �_.���֕7�F<yv,-D�� ���2դ��!��t�"%i�"O�!C
�[�.�z4*B��
<$"O�[�aԾ'�d)׈*qX^�8��'�(�<Ad���sp�P��	?|��8�HF�<	�8z���@��$(����JM~'?�S�O[6�	�A�^�r�ƋD�1��H��)��<��Ʊ�΁�C�K:sn^ ��RB�<q�ᔚ�^�Q�+W�I�A��ʔ�<�
��,$8�Z@.���bcم�FX�$�O�3R�K�)}�5�%E§Z��@��'��'�i�v����`�`cW)F� q���'�S���C9K��Yy�E��|7�Уa�X��OF���k�-�d��fj�@�|�q�DyX� �O��9U΁�0^j����p����7"O�%��ގ+��	��NNF�4%I�O&Ͱ$/� Fn�8���70�yy��#}"�'������,D��݈��++�X���O������}�j'�� / �CP�D?C�a~U����ꏩ\+^:�H F�Z��v�>�
��P(&$��7��dB�"
���g	�p����'l$��'���
H���ӮeH&��[�PE �[4w;0�ȓTAf("V���/j8`���f���'�a~��>mP������qT��а=9�{r��_�i#��ݰ,[���D�	��y�b��+@p���0k�y�G�D���'���FyJ~UC�0`c���R�����`9&�UV�' �O��'źl��"G���@���WB1Dy��Q�ܪ��%���`Bǀ2Yݔ���g���?i���CRU���
Ul�i7�X8,�V
Oޅ���?#�V-#Ü	Щ�|2�)�Ss �LIe�j( ��z���'&n����|m��:�,J�}, hs�y"�'�,ѺצT�t��E	{��k
�'��X��1�v4��ũ:N��	�'�>��6�L'h�~PZ�C��5�ޡ��'0��@"Q|�4{Ҡ֟*8%��'������YX�P���ة�	�'A�Q�#�.<[�0��w;d`	�'�`�
љdxȅx���Eb�{�o�'<�'�� ��N�"8�
�K)"��
�'�D�(�#�#y�(�_�Hٖ�u"O���e9>���ҧ3*\IJc���'�ў��,!A�<F�
ё%���T�RX8"O<1���x�&@s�Q<Q�T=3"O�ݪ��-3[jX��F!z�޹C3"O4p�2��7 *a��F0e(���"O�h�q�S�0%KkL6y���"Ox�)�b�1V���P�I�;θk��$8|ODZ�(ג(cؙ�È.Hn���"OM�5�οc�\a:#h��+�yqP�'�	D
4��a-��%�Ш��iN�*����q���qJ�5��{��]�g�ȻM>�������|����0$� � (ɳ"O�i�'��*3�`1C�X,m�*�PA�6�SⓥS"�d�a��Q(��Q#k u�jB䉰 �>�u�SM��yc�n<�C�}"�i5>�C@��V��9J�M[tM�o)����f?i�� |��<��ů?���Q��M[�z�Z�RK�4Di�Ӹx���_�O�h[�j�p?��j�d����,�١FN�e����!D���'͈�-pʥ�QbȦ���C�=,O����Is�
W���Hءe̼8�p5�M<�O�Ϙ'�����%X���kg%��7��MQ���1�g�? ���`��:d�� pQ�R�a��٩�:O����� �慪e�>����&+�44y���$>�ĝ2$�+ٽ-�2��K�[D�~P�d�fعl|X�s���'�L=���*}��'�6�S3V� � ��]۩OVc��D�T���lU�U����8�#�eΞ�yR�T�s[>��eC�-��)���'�ў�	�䂔��y�B۠_��"G"ON}�!�Ʊ?����4��*^0���	g8��A��\��$�!ԩ�Ah�c3D��ذ'
�p1�y:��71��9�2�(�	a�'�N���'֒�܀s�Q6=��,P�'�EyZw(�'~��P3��!�S��km3G�!����`�v��I�r��w.E�l��I.�yR�/ғV�Pa���(ƈD��-WO\$�ȓ$4&��#��$r�V��)W#�6}�O�=�bE��(�Gb�C�АbJ^H�<��:`�Xh3���		���)�o�Fܓ���hO�%;F��2����L/x�O��Z�b9�X��.�E�"����6`�!�D�51I�SFD̢m��LPw����'��'��?I�Dd�"�bAJC��)&�aT�.D����d��b��AwANh �G�O�7�<�S�'��^!+d�2�C[�xp�uΕ r�!���`��0U�?�jq�U5=��o-�|�DؖtoH<�a��)#�y� hӶ�0?�,O��1@�Z���X�.A�W6!��"O���-�;+����gKD2(��+�"O�� �'l�}k��N.
�f0" "O8���LUdy��̐t�"O���&C6��5��J��b�I��"O�s��T�y�9s ��e(���"O��sASB>4�!��S1C� ��s"OT(gl��\� `¥�7�Q��"O`L)2�/aH��Eg�&���"Od!�W�s�Q��E�	w,}�t"O�e��Q7)����پ���!�Ó\uԩ�fɑ�)+�Y �ժ!9!�$���p�I�`O������˿3!��=��@R�J��߀{�,��<!�K
{6V���-�*�}SҊ��&!�$�CJ�k�	I�P�0�)���q!�ѹ+&�	ԠE&D�
�:D�`!��ϫ	�����#5.ʒ���<U!�$���֌�@�E)t�.�ʆ*k!��;y��H�R����ZL;׎4cb!�-p�qu� �<�ܥqQ(�7jI!�d
`�L�����$�28�pD(:!�DZ9:�8p�!��{��t��E!�dA�Ww��J3C�1O�Xc1�	�p�!���;8�����;]d^����D�0�!�dŪM�p� �&��uKv���
�9.�!��N	P����/eI|��)ġR:!��@v�LBf��n�\�q��<_�!�dP�`Dp��Ð_� Չũ��!�D�7ij��)��A�PD�v��?�!��'>�[�D��S�� �Vh�>W�!�d�9=�M�#H��w�T4҄M�2�!��	1Rk�5���	PE�����H�!��9��)���i;�t+u�	1D�!�d��Cdlu�B��>u�V�7�!�$Wp�dʥN#�
�Q��%J/!�H�Ʋ�����l�FY(�g��9�!��R;êm*͎� �Zh�F��i�!�� 4���&:rVѹ�LT�!jp��"O0�`�䕃l&��+˄�s�N��P蒌AF@��J9%�R�A�'�&�PnU��"�5a�.�@��'�*��4[����eQ�����'Ȁ�#�
ϫ�N-�U H�}U��[�'h�Q��ނ\��6���jy����'���"��5C������:g��9��'�1�V��&��!�^�g�T��'&�������9qV=i�ԜZC�I#��"��^|!@�̀��C�	;3S���F�A�%��1m�� q�C�xo�$�GW�:�=s2/� 0�^C�ɞSY��s-J�NΑ����7�C��0����BtI�hh�NI�*C�ɒN�0eqehAL�Lp��:*C�	}�ܐ���˨:�oʔz�C�I�s�b1됎��8�$�¡L��C䉿Mf��� ).p�؅�BڈB䉯(\P�,I�d���P��(	�B�Ɏ����Ǚ�0:��J7�X�	/�B�I���Ī&D��c��ʦ�ܮY^RB�I0���2C�=Cf��#�e�(.��C�	2�x�g�ʚJ��'F�8��C�8��Ei��ܤcq�2�K�	ntB�I�d>B)y�j�h� ��d�/�C��&8v��1eT01�Ԡ��'��Ms B�IZ�a�&� �`��NB�I�p�j�1GM6og�l��`� !�$߼pݐű$�֢5|�i���fe!��'Rc�)(��3|
����Z�W!���7<�� 5+	P9K���!�DM�i�x���W�,�|���ϋ6/��~���5��q�!dF�OS8�9C�.s�T=Xe��u�<IA��4PTL$+n�=�E�S��Z�'jV�rmԕ���~��L��p���m.N���Ya	�W�<1�������+kRl��b�#.Lȑ*\_z����Y?E���[��@�,#[@U�ҌD�i�Ʉȓn�HA���H�q�dh���.Ԕ��:��8���'I:���� ͉��O��(�-��O|0*`�C�S=�H��'��1�
��N���u�hY�Cʌ	B�M��oXI�'+�Ȩ@`V.t �lK�"�#��I�r��"�Z��с��X�H���\�Ӑ8$�u�S���M��a*��B�I[~X\:#		K�t����葵G�7�����J�&U���+�g?1��x(��s+�':�p��L�<��%�$Bm I+#k�
\"���B XZ�D:��R�6�����a+,,��;��O�|#�o2k�*�!A!\76c��'24 ��dg�ę��޼�rE.ƥK��]+e� =?���Q�ȠV��~��PxfHa@l�u���C��4��'��1�p��J Z�����r����>�8�Æ�E*'�NKA�Z�G��B��?=��ZqT2�A�5�� _U���à)\iQ�N��\4��UE,�'�~�o	�	BN��㜠G-T�Z�n���=���X���]�ȁ�7�G�{���U�	:������(~�v4�W^���c/�̺+���ã�؉q����]�eA��D5sKqO��s7ڸ'�]�qq'�ŷvG"bA)��4V<QK��8?���q�)� 9x3E�5�p?�򈇇}��xz3`��uӃm�#*�v`���<���7d���Q^,"���Q�n��hs�8�Ī�"Ϫ0���Y@��0p���SG"O��{do[=Q�����b���ŝ?F���u��<I0E`f�
)]��K�/�?T���˟�D�4u:����$ljݐJ�~;azrb�3�vx�r�?i`�u�jd0��K�̬{������A) Z�t�`��Ե5�ϨO��Rb�
�HEZ6��-ߜ�{���E.Մ�d����	�_�-q�h�5YF�z�n�S��1;S)i�9+�G�U쀉��	�$��DBR��1�
d�5ə#xX�)&��F1��"�$JM �����?a4��B�4J��}����<Y�
=��cRk�<�wf�6x��,�vн`,���n̸yb@�׉�o��� �Rk?�@�>OHh�'���S�? �)"�d��3CoK�f�d�I��'񈍑�Ř2B�Ҡ���2�a5�6�� JZ!s����'�`��3��h����	0�<��ФI�z(vu���['���\¢ʒ]�,��z�+X�0�>�@�'���vg�;V	�e���9D��R��Jnʰb0fU�%��A�IW,dJ���=ф�<�`LS�[��Ijâ�3X��8�5D��H�)�)w0� �Dʂ;=>�9��'�K��W}B�P;��9C��CO�<9e��1�d���:f����@��H�<)6�,lhP^ؔS��/`c�!��b���+sC�UY��XKA$;#FA��p9��%�B9�Ó@�'@N��ȓ@�|m;uH��|���#7��2������R�`q��j�x��	��,2Uy�#%�
ap `�!�YÊ{"���c�� uX` �ޟH!wI�;IQ��P�ᖩR�D��)D��C���:�>i3w�,�us�q�ܼ�G�&o��7��9a� [��5:��S�S9i�ȵ��_�-��A#������DK�o�T���C#�ybOK�����G�� ��{�+[��|;���~�ʓA``�|�'���6bʠS^*!B�χ
�yX�{�gC�(�"T�Ht�O�p8r ̞v0�a��a�e��NǢd��١ǀ��t��d�O�iP(ׇ0���ٕ�"���O��09��O�lj��V�mf��T�i'lz��F�4H���F�����y�'���:#��*�@��-�VSB�-p:z��� ]��R�T3#���:��<%?5��l�6Z&q`��¸	�t����=\O%����(���q�'" 1�$�6wW�ٛ����{Z�y�B��D�IC7��<�r$9�gy�_��8�T��33�Jt�'�����''2��@�Mt���D�DJþ,� 1���+~,p�1d�\;�6�� Γp����"7lOtac'���t��U��n��'f�	s�׷u���[�߅z��d���'{�^,R2&�3`v����S�T�	`$
e�T�� � X!�Đ�B>}1j�67�ZŢ�nC�"�F��&-&L�æF*Z��a�t�!V�8�O�i�O_����j�#-R$)��Ϥc���3�2��D*I�pX���EE��IبD���4+���9F_0vV�B��!X�ԲS�_�h�qFBC�^�=�3�/��4��7�����%�܇y��LI�@!$ވC�	�Ѵݠ�I�)8�$��T�+�z���y�\��ӫ���)�'m�.%���a� �r�A��6��dJ�'g���	�
����ï�&�tC-O,�{3�μp�h˓0�~�C�k��Nd	����'ꖡ��ɭL`��	%킑j��V�?�H�&�	d�ʉ��NX3����SO��sꛭ �*�r�A'(���*Q�x򂃋LU�ţE��9kZU��X$��O�ԍ$���0����,[����	�'s�|�fo�"}��=R�B�c��TgK�i�1�'H\�� ,�.�¸O�'k���(͖[7�W�.E�.�3B�,�<�sc��rr�-F���o�8O��A��ߟ(O���@d��<�����8���HB�p_69�R�ZAA��"qh�c|����	h5y�� Kd���K\�LOڤ�S�@���(
QE:�C֛��Q�����z�D�@T �b���H�D�!�4��ɧ}� h�Ֆj�>�ڢ�S�?VP0��dm��ɔ�o�RH�gA3D�t6�C�	`�/�FL�wC�(-y���>���WV�d!�k�.
dqO�n
�)ڬQ�n�;�j��c ��S����n�v!����A����O9jN��*B.��תE	���q�jҶ(D�D�M�Ffh��I�w�����6�p<��M�9$��!��.?9r�Ƞf�Dh���Nv�D����R~B��>��x��4\��dc:���H�e	�8NO�œ�ċr�O�ӆ#�mZ#3���C�T]©"C�1	LxB䉕	�r�ڂ�	���8g��#L�JP��{b��&d'��vј�a0+��l���@19���ȓ�J4�6�ޟB�����N����'�F�����yWl�b6����@9����'q�����<To*��UďE@jP	�'��Z�՚$;�p��dC�9V��y�y��)�J�%��Dߠca�haJ�	�C�	JZ�(Q����L���Uƅ|#<�ϓ��]��F�$7�T �h\Z����S�? B�Pvnڽe��˔ �k���@b	$4����=>�2D�u�U�iz!F!$LO���r�� ����'�QS��� D�����Q\n=S£B.^����T$4D��K�Á=g$&����D��DO5D�LPT��u�Yp5j�'Y\(�b�>D�D▩^ w���6��0�p�B9D���u� j�ʇ�͇o��Y"*=D�p�L�M���wI	48���S&8�O�	���~��Ɇσ�f�@1'£X ��'�EhS9e�j� �#3>�iN>�#�~¬@�@��9�D�|��J�4dA‒=�d0:W��/�$��	a��u���>S� ���9�$=*����!�"�LKpt�s�c���� �<D���5f�=��c2�"ԣ�+K��O��`C����O�@أ���lx)@"ȧ`ͤU��O�����ŒJɖY� ��yq��!�@>�4��m�!�SvNi�A�H�n��0�t_���êqA�'�e E��F��'Ѥ~�.���J��E�6��HMw�H5:e�P�&��QQ��C�,��LY��4}��i��|���K��^'��\2��Q2�V�\�R,�'�3J�����cPꙠ�OŒ\|:5���4+ĳL�T|h���8���%
���Q�P� HB�@���Od�e'#l�P	��	�'�^�c��L�s��#��K���,ľn��Q?���X�x*֌!@��xH��Bg/"������E�
ܱD:8qb�>1b�����(vv���$�';�L� �+ĸ1��,�e��.5F"a��8OF�#Ӊ
]<��BC��'<�R�P��y�ԟ��j&��||�Q��>$�����,d�i���F�7l�D��"1��
�n�R"���A�$�N�=Zq9�/�)zB��F�ŀ�@ӧ��Dx`�Z�J�I���Mh8@�∥�\r�>`4�tj�1O8�1��§p�(�k���l\):��m𕌂���ɵe���W3	~Vp"��חа<%E]�� �p�Ax�y�� �<!����`�A�$xɦ�J!�o´I��u�
;v��z�ɇJ԰BI
�VoB]���>�OFM�b�_�2�m���8IP�-x���;?�Xh�-��~B-�gr����i�m��A�9HQɧ��ʟ2��y��E66\���AF���O�!�Y�_^�ih�O��H���F6%y��V���JU�"TDy`�'��xu�Ii�S�O��	�X�;�1�t,�%5G&X0�O����/�a�.�O�>��s⒂'����OϘi�l��)1D��y����)�y$JT�V�G�.��U�R�˓
g:��`��~8��C�E[
B>��ȓF=� ņ�F�>�[e*L�Z��ȓ~xA,D�!%D��!�6�T��ȓH������N����T� �T��чȓSY���a0W���P"��%��+X8��l�S~d#B�нB+�!�ȓPvN��O�&��ђ��	?-FH��	���+4��->�d�:p��9Xh�ȓA���ȉ��cP,F�_�,���x�#ef�^��'Ɯ.r�0��*}d��;?}�գ�@�f��h��I��+��S}�J�;�H�`�(�ȓh�Di��F��=�a�
|I�ЅȓqW� ���	���UxD�B&(��ȓ:��p�W'Yc������%���A�U(��M�1�`Q!��& B剪;n�$!���2=Jؙ�,��l>D�؃����{���"��Dq-�1;�?D�X�d��Z��d{d"!z=i�H)D�$"��ǚ<�X����U�52����;D�������4xG�9�J�@�ȗs�<���#oߌ��*�ilpyPcBD�<cn�)c�����[)o�>�3�+�H�<�5La�ͫ�Q!
jl�I K�<�c��26qpb+W����Б�FG�<!�g֜N��f�ܙd�	P4	OA�<)����\�Ru!O�1�8�+P�@G�<�o�t|3'�Z}Z�I�u�F�<�%s���ʑ�(Wx$�2��z�<Qï�
�����JH&�����
r�<� �p��2��p�f�:K��M�"O,�1@��P��s��K��ҡ��"Ol��N�o��t�s�!|��b"O��R�AX)f�ؕq!
%��"O
yK�Z*L!F%27;_�2�"O�m�2́)h�hbi�	�j��A"O\�����,�@�]1Ko(�(�"Od��.�Y�֌ �eD�uAd���"O����+��Pw$�&OW�0)`"O�-��G?%y�L�`c�:A4��"O��%O�}=@�C�!0�a(�"OX�S$H�25�`��"�)(ȡ�"O����%� ��U���k��"O���6�aO�h#�[�M&��!"O�T���_-)DxD�Ԭ�!%n�*�"O�ju�W�mKE� #څ����yR��.0oyR%W,'�:��ꃤ�yb >(/�JF,/Xnij6O���y���}6� ����w��&���y�%�)� l�b��)�ċ��ɢ�y�1]��C.A�O�t�%��8�yr�ʫI����k���Q�@[�yB" jDޱ��tݲ�U� ?�y"'Д8Q�2F��n��DY�%��y��E�&4�aJG ^�)"�H�^8�yR�ٿS�&5!c�%�8��2�y"ɖ�~\��@i��x�+�)�y���5�V���۝| @���O�yBɏ+&�ԋ2O��v�,l�K�yR�ԑ޴�x���r0佚�d)�y2掼nR"����]x��2�A�7�yb)�L� l��̋9�D���C�yRgɀ=��<1	"Q���yb�/n�h��%%�l `��y�π�y�r�7'D�y,�ා�2�y���4鰁%Jެsxʝ $�y��E��,B�B�4Y���:LI�y2�Sbd(aR3M/]��i2�o��y���	Y�2�3�à �fpI��9�y���=w-Ra�i�Bm�!-�"�yJ��F[p���ԅc��U�`g��y".��)M2� �ҟc¹�0-P��y�[4����C�g����铏�y�k\�;�|�@�
�
���ؤH� �y���*��10��U�t��8˳e�y�D��:Qbad���z?
!C����ybK�$h���VM֏h���X���y��	K�@9�i�4l���#t!��yo �CFT�2�$E"�����y��(tnpM�ѷ"���R���
�y�,G��ٛ@Z%V���J���yҪ�� �\�V�Y�<99��Q��y-��D:��CN�9�0���yH�l��LN��$=Y$C�2�yr�W�;UѰ��t�H��s�@��=�N��;|�W���N�n4D3�͖��X��	��c��!9>���L�2�6��=iDHtZ@؍���B����M�1x�ȃ�	]!���9wK6�H#I�x:�
t��XyP�K�����	��"|�'2��)�$ׂ5NL� TY ̌0�'�0ژu��� ���$�0}U�� %�����@x8�TY�kU<�:���	O3���&�6LO�L�$'����Y��'�)RЬ ���D�0j0�P��'�4%e�b��<��g����y¤�
b�ꅳ���p�π �I���'+�z�Ç���:��"O"��*��S� %h&��6K�(�0��O�\\+M�X26!?�g~��˰��M��ʠs��;�fʉ�y"j�!*18�f���,}��J:L��ePrᓁ7mα��IN�p�R��}��2� �%|x���D�	<KT�c�B���~2���q�0�S��Ҏd�H=`��С�ya�0W����C��P&��A������'Nְ�m�	��?�:��:��)
E��E�޸��j/D�X��,��I���
E�C��(3_�X�="�>�#Wa!�A%���yI:D�gM
a�<���9��E��K�s~8m3�]i�<I�ر\�z�*��7`t��Zg@�k�<���_m�N}p�A�&�@�;���I�<a�D��2��u�۸X�:��^�<F��<2��)������P�Z��B��z��)1 �Ц���x!��
%�B�	�w�h0���M�#�����%�;`�~���*��+�)+�Odq+�DXTB%��C�?b��Yc���s3H��=�O|���Ⱦ`��MC�o�O��y��"Fc����Z1ex�4�b"O��Fj���jL����Y
��c�i�L]��bV�Hs��(փC��D�#�ڨJ��)�	�$*��2c�lH�I���z�`[�z�H�˲-��<A�HЉrOؙ��K� #�r�ˤA�1@��xW����	�Q>�n���Zfj�0d�("�.C2��H�=q���rt�P�t4�'��l�"�@����-��زp�'y,���$Ș�a{�3?a D��.�8O��i�,�V�X ��� %��ɠf��-2�AW'��G�Z9�4Em��X��۶tg�|hm�{60��ȓ�~}j$��
����0 pm��h�I�C>@�� �L��}P�L��`}�S���~�1R��������ҧl��H�'��(�4��-9	�R��4���Y�$,�"��="D�aU.�4��Y��0��<A�#Į*w� h�l��?��0���W�@j�T�ժ
�%r#~��oF!<�H}Bre�1Z�%p�L�h�b �3o�'P����'w2��d�!5D��H��-��U��C�MO\�qĜ�~��D�P�h�b�aa�'��}aB+�!B�E5�[0�&�8�'���q�@�b�x���+K+%m�!C�4��-0I>�d��%U7ǔ�)dMc�	��T�+
��$i��_�FD3����{k�{�(�4b:��F��(���B�C�F]���%N+&��b@mH<9rm�o ����0rj@�+w��_�'}�D���`(5�~Z�
W�pw�U)�\$�����X�<)t�ô-��X��C�\�2-�R���D��k�.�⥚>E�4-�0_��i���-7�����%ϐ�!�J��e��苄?��]����7��$��
u")�V'���<	B�F�x@�$B���R�]x��h`O$C���"���6<4�x�H!mY[��X�f���їȁUn!�dQ�t����s�ҍ|.K4 ��y�'��L2��@%8�<Z�ޖwt�A���d��=%p�A�CEV���ʦ���y2� p�)а�fA�6a���U��p�1��"F#.h;��+ܸO�' <8�va��'v��`�U�g ���'�q��<T_H$��3u�8�Rr��9hz���Ĳ :�({�����<� 
��[�.5��#V(і�j��{8����
�^� Xs֪��c�:��3f �|��y�2��	�ň�?�!�Ė
Hf��t-.y漈��\�	Y����#�>���қ���!�E�f8(�����!�;
_*�`C���=�rq�e �>��Е>��J L��>�O��b�'!���S�ٖoIb�;�
O�U���^�G[&l��Q�R�6�J�샵k���(4��'�0?*����k��1�
��D��v8�L:�o��e��:𓟔��L�R 8U{P-��{N�p�*O�����AO���R$�/ �Ǖx"�H�4Z
(F�|��d�ߗq���0lK#$�(pN-�yŔ�L&��B����v������$�DL�g�D��z|DM��KM�:֍îY�!��:F��t��,�Y����P�>�!�
*1I�5C��?.b��m�!��̄s|�UG�3z�f� ��0�!�� zM�r�
�����Ƙe2Lk'"O��S&l4;�б���	*�5��"O`��[�Q��́1CT8s���"O.8 tD�	�vH2�HlbD�"O�t��VEӺ�SF�'dN8�"O.�)�h��M��P�#kM�$]zD��"OA�cC+-9b5J�*�* ���"O|H*�E�<
p"_�]u`)Ic"O��L�r�FE���dPl�U"OP5IbCV"r¬�P�C@pP��"O��R1��5�t�u��v�j�I�"O��b�Z�����S^����R"Ot�k5,;v��rF��o�Ԕb$�'����*��x/��2g�yI����O���{�	��j�WN���ٗ2�
\E}2.�!)��a��i�9,��)�9�Cr��TX!�D2k+Z����Lp�"�T�2H�	<�l`k�7��)��3J0)��Q�Hؤ<���  �2�U��!
%!�PΔ��(S
{E��A��V�ɦ�4#f�!�2��Aj�3?�i&���>cG� ��,Q= ��{��-L\�?�#�E�:�[���l�Z���(6c	+7j��U�!HR� �E��c6��J�`��\�S�O1ƹA��]�w����@@�b����]��U�/���pk�D�i�*klv�>�r�N;Y�|���ڱ �Xy'n�<�%��1o�f��"�=,O����Y`.�e�1S6�يT4O4���f�X�Z�۬ID�'�F�jF6Z���[��K�v 䨀*�h�"5sfm0�P z�1�\ *@�� ��(�%�%/E#�G�H"�:RHk� y�"Q�6d��`�, ����^����?��*J�<t�+䨘�n�\x���<�{��|��'�3A���i�_ (�gj2N1h�s `�0�4�{��B�0�=�4�ƺ.jC����)�'	H��5�L�rb���闩KB��'d�y���D?K�F%̓ ��J�fX:�T�>����(L�����ٯC&ȕ��Ƣ<�S�Ra��*/,OBi�S�_��EK�G�}:Z��!0O�����5�n��g� �il��Hw�F�38��P^���Y����[�|���F#"ܽC�&НP�����	Ň��l2�ǟ0X�����h ���}8��m�����BI�G�i>�X�ŤM���q��C�4V�`*��!�5ZZT℩ܟ{>�DT�Ѣb
%(G�!�F�F8<�Z����S���Ij�l�����S[B��"Pa@t����-�2�
2����]���S�O	�0 E�b���"AE�yf��1�'v�ECv��J[�A���r]���N>�šs_���dB7`�������{�蚃A~!�$�(2�D�R���^�,��uA1k�!�D'7=pTKr�����A
�W�!�$�{�tZ� %aɂ@B�V�!�	�"%�wOZ/�0�o��!��6cSB�QA�_6f��Q4��6�!�dE8H{t9��T>a����햤�!��7O�6p���	qgDh�K9:�!����(��&WR�����Y:G�!��a=,�� ص6w��#�#�yM!�DL%�����C�xt��2$��'#!�ė<g�l7� �G3��XP㗘o)!����(�P�H��8���b(�0d!��O0(FA����2:���S�A��!��P�8�B@'�u̔��Ꮛ;�!��?y�Ȭ�$kĉ ���RV �e�!���<{F@�buC�� ���`!'�!�d�L2ޑ;��[�4��� ��S�hq!�51j�P7劔H(����@�
l!�d��P}�E��
�qR��C�N��!�D��2�2��4�Q�	$I��nH3/�!�ϖ}���h���#4�������N�!������bo^S,0Tr[\�!�DE �p��J.>A1w��!�!�$��K,�$qw�y�i���+i�!��Fg>�Y�ׇ.L��LS!�!�� ��dsK�9��F�%h�$�"�"O�󀝶K�L����,���C"Oj���)F�;�Ta�O��v�P1"O�1B�g![��U9Pm�{��л�"O�q�6`"*�X<J��L�h�:<�"O4���.���˧צ\�)�"O��i��Ƌa�@0��HI��.���"O �p��"w�.@�Ԫ$��"O@�1�kL�Je�A��A$�"mc0"OV�b��w\mi�#��
'"�9$D��lA<<����a)Z$Q"p�;Pb�0{��O�SU����2(U�Ah2����4L$ Y՚>�Ƀ�!i�L�|M~�iLeRr��ӏ�-M�.��� RB��_�[��YH��A$�0|b���T |����&Ul�j��|?	�C��6�:p�6}��� �5	Z�iA)��,���J��+<�S��U�@���>E�t�J��S+��Q�d҄ș%1F��j�$>� <�M����.6Mp5�ᓬL-dD����=�����#!9����b$M�-�JK�8�C�~z��)ϵ�n� �J����Q��%8�X���R�V�q��]�>+bDP�S?�F��ɜ[����R*
 IZt�	�I@��?��

�,����e@��)�GҜ-{�L�\%x�	���X�Xp4�2�}�E��p���"�f�[6�K4xB"l���Ǩx�A�>e��@�7�V?1V���L�$��@�"�lT�MNR���P�@��� ԭb�D����t@�~�	&�I�|��)FT|���umn)�1_�4���/txY�۴R�a@�J?֝ݟT�l�a��}��JV/s��!@�J~Ӕ�)!��`j� e��]I�O��Sm��T��	��լx@>�O<AJ�+Y��xn�:�PG��)h�*Tk@�@6>�"@�� l0�	� ���i��Ȏ���d��B��4,�j�N�gBҊ��	�nԛ<�?O��AH�<t��wl_�)o�Z\�|��h~�a��F�"D�E'��t�>ɍ����D�<+�(z��%O���k�����0>��fķGpe9��A�0�,�`i0.kDx�a��+� ��C��S���`E��j=:E%2�ɚA�LU��S�w��eZc��;���bP
F(�O��'� ��Hv˧V�$��o&b$V�V #����F��8;Jr�'�l:���l�����>﨟輨�.۾4�J��b��6i>B7�'��CÍ�*,�ʤa�Ɠ�t"a���ֵ
��t٣�M�h��y�Ҋ����h��}�
�Jf�qP��ˁB�xS6͇�D1xu��?N~Lb��؊lZ����)�d���ujJ(�A2)lZ}�ۍo2Ɇ�����r�˖���P�AS�6u��Lj�
�dV�Wy����
?�D��ȓ^��)c����LW�T8+��C�fD��`q�I��O$�P���	;>/&���OD�@�-�8��d�7�2%��]z����&`M��PîB�Tơ���e+��H �0�kG�!��Ćȓ]��'�7l��Ҷ��gt���>�\�':SeL�F��?^z��ȓUa����Ί�p�H�fE
��@`�ȓ�H�SSi�zP� �P::���C�^�CtH�M�����A]2.8.Y�ȓ���'�ӭz'&X�cҵQ�J9�ȓ \�}��Gεw�ACA�\�p�ȓu#jm!#�1v��DCƇFK(�ȓ	���{Q�Z�3�`4�p��o�,��ȓ]���Al %ˁ#J�%.���p���cI):�n���"R3�d�ȓ���0�ˋ�t�Υ�t%��-��b��]8q��XDpS$�]	�͆�L� '��p�������Xc"��ȓc��,�"�ޞ+�<I1$��,ex��ȓ�e�a�FH}����fV�]jņȓ"�H'�J�Jf���uL�:F����X���)��#(�!�"GW< �&̈́ȓ3��\*�k.���� xp��S�? (�#`:6���ِHƌ.�ͪ"O��vE��A��QBBH@0��i�b"O`�[��PP��eSe�*���d"ON{���a~,H�W�+jd�i�"O�av�)=��V��-�BIx�"Ov5����a��*��w�����"O��a� �`=(���	�.[3�y���r����c	H4�l����y¢�'`��
�ʝt˨1ᓉ��y��@�������aI�U�r�T>�yd��L��H��� B��8Â�̖�y�'[��D��ʒIU�8C��yr�סp^��d�A�@�$��a����y�j��7BPh1��7h�ݛ!l_��yR�҇!�8�0��_�,a�9@鏁�y"^!8�tX�G)���,(�Pn�0�y���IHbY�T�D&z�vؐu�M��yb91�\[�b��ZD�o
�y��>`
Ⱥ����"�L�Ys�ʊ�y��</�Չ�E	.n<pg���y�&r�� A'ȸ_�$�	U�H��y�3s�1��	͔,Y�<����3�y�tb��!�������/]��y2� ��l��	��n�n�94� �yr�}�B�1���f\Ą�I��yrǤdL���K�O8�))`����y��P�鰤��HB'L�h	ڒ.@��y�g��g9X�pK�:���/W�y"*Z" s@X;@�RW-E"�y�OL�p��{��Iw���y��	G�&N�z��|���_+�y2B�h�r�3��=��2&���y�'M�>�2I`�O�3;��P�Iȭ�y�޹Jf
�x�䈧%@���Vg�,�yrj���s�J}�)�����y҄��7��1�!�;�@� Dᘰ�y2�M�D���0M�70�E@���yR���Rd(J�+إ�u.�$�y��K��<� P(T�o+�Up5Ȃ��y�"�k�F9Jq�C�c?j$)ƦO��y��!�viI�⁻*�2�զ���yB���`�|xҠ+hH	E%���yb��{>��H�ۺo3�m��*�yB�o9Ry�cM�9j�H�C!���yB�@_u�U���aݮ��B��y�6x��`�LU�x\	abD�*�yRhӆf2���eӺ6g����dҥ�y�X;����BC#,�(!���\.�y�8m�������e�֬܈�y��:��A���t4����y��O"�R
� �-`�N5�A����y"M�*R�8�x ��
D�Q�1)E!�y�Cբrj��6�Rx��(��y�`%2]�����(�$�I�K�'�y�mN��������Z�qa'J,�yb�6�|s�DX�0��s�̏�y��ܮKN�	@�1�6U:�bP�y�J�^��'�8?�jXB���yҏXK6��(�hC=n�x�Æ�7�y�L%M+�;�/�Z� H �́��yr�It�.� �ũW2���*й�y��\����MKU :�������y��څEl<C&�E#}J��'̔��y�	�R��%��'S8xܔy��	��y
� $b���X��k��[9�ִ1�"O>�iP\A�5k�C-\n�a��"O�R�e��h��䡕���t\��1"O��;P�؎zMĝ�6(K�H �d� "O]�3l��&�zI��ң"O�kS���+|��s���4)��"O��rf'�'LBtɂcfR��U�&"O��(� U�C�Tu�S	��
�"O�qSV�����W��~����"O�����8�P,�6�	��9�"O������%���g���*�I5"O`�4�G���٠�bD�w���5"O�}�5�ٶ[L��y2�)�y�"O��"ca��2l9vaӼ)V)�W"O~���M&R?.����T�z�"OfH)W)N�S��d D������"OU�2%C vm̅����%�^��"OɛN�5H4��3�]�TAn�w"O +r��PJ؅�b�ݭ1�42s"O�q
�扝w;K嫐��Z�"O�`�V�Ӏ7�d�4���*�dL"O�u!��Xh��aM�G��`"Od�B�">
Za�j��b;V���"O�E���  Dz�oL+N4�u�"O*����.'�:���Ͼ3���""Op=��� �9"�m�JR�$C"O���`��b[�,�
K'h�Q6"O:h�U
��W��$�P�̴ 9\�@"O�<����¥�T��RP��S�"O�U�E�Z/T�M�Pb@�5����"O8�"�n��`bZ�q�BX�`9��"O4=�0▐V)2$c���p�8�s"O�d:�BƸw^
���]6[Vvݐc"O�\� ��S ,��E�+p���"O�[�c߄)}Ȩ��c��X0�"O\U��[��	�bB[�8�=X"OP���bOزE�G}ܝӣ"O�����������%΀�}oVB�"Oh<�Eo�$�@��*�3r_(\�5"O$��r C>����@	 
�x�P"O�4`�Jͤd�ء���6�@G"O��``��)A��B7��k5�(�"O��x�ǅ��2ex�L��w����"O^���Z�T�ܤaQ�V�uV��c�"OD��bH�}�r�P1��j=T��P"O�A�ի�1�riQgFC�uG:�"�"O�Ir�lF 1��d�
C+!��i�"O���+ X1������b"O��l����ɶ)U)%�
i�5"OR!g��0:H@�
Ȭo��D�Q"Obe��섳�����]�wκe:u"OT���#�*Yv�����N��x�"Od��gݨ�l}HA��<q��Cq"O�Dz�E!fY���fd��k��y�$"O`�җD��<�\0��ɽd���b�"OHɉ'f
3���t�̡in�� �"O|����׽9��[�ɓ.[�Xp%"O6��F#V<I�j\ң'�/@Wt���"O
�+CK�F%�PF�]�8YS"O���� ��q�"yq(7~Q+�"O����P���F/$�yV"OZ�r��J)&����&��7��D+E"O������|e�4y��pwAk�"O�#�_T�q���˯FEu�Q"O� ��k���qh)����04QXd"Ot5
W	M�(��q�[,#��H1"O�9��є&�vh�&�pe�t�"OTxf�:��	�� 9J��Q"Ox�)A͏�y�赩����"7��W"O� A��Y��
ҋ_	��R�"OV9@,B~���sT�N.��	�"O�ų���:F�1�D!��!��"O �A��̈A
������Q"O�|8��J�i�p�!��O=	�N!Z�"O�RpEPvA`���(*l�܉�"O�=���k�P��凗)>�-�"OrqRf��+: 4����08�iD"O��,M�i��+U
&��6C���y���$j��	��Ӆ*D\1'��y��ռ
EP�R�'l���5��(�y�7f�H�2큼m60��,��yb�^8VVb�b)�0d |�	�b
��y���̚%��Ƹ���O� �y�(�eL�	���Ѩ�3�Q�yB�M�L	�)RL�< h�"��y"�x\��0%�!a>e�!!G��y�̎+�n��c��щ��yRP���H��bW�I��ba�-�yb��ZZ�C0+*FKJ �E�:�yb��6hW��C�DJG1���c#��yr,�:�h�c�B-P$!���8�yb	�*2D�7 ��At �����y���";gT�X#�_�c2��� g�2�y")F:Uľ(P!(�_��R���yҩN�7x<�bo��Q{��( g��yR�N��x�A X+�d�I�,S�y�m�Pز�k��`���X��y�Ό�1&�`j�g��+	��RW�M$�yrD��zNR��!�FaA��yҮ����ӥ��򩂀O�.�y"�C�>���
�$�����,�ybo� ������R���Rb埂�yR�?�Թ2�E�8S���f
G��y�HG    ��   �  i  �    �*  �6  UB  �H  �Q  X  J^  �d  �j  q  Zw  �}  ��  _�  א  1�  s�  ��  ��  <�  �  ��  ?�  ��  ��  �  ��  �  L�  ��  ��  ��   ^   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.�T�DxB�'��PnS�8�2 �f6Q��$��'#j��G  �?�	{7�>� %k�'A�)0�˲e!>�i���%��ə��(Oz�J��_�c�q7(�4GW�ȱ"Oр�Hr�́a6-�E�	f��E{��i�dI�hSm�?�4��Ń�	O!�?�[5)ɂPɌIP��vY!�D+q#b��@^����A�芢
I!�� ���2iR�7�`���R�/PFxe"OP���]���A(�1�4AV"OPձW
�=~�����T�Z�[c"ON!)�fi�	5 �H�4 ��d,�S��:6T�����x�d@�PoxB䉆��i�7�Ʌ4�0�sl."J�"=IǓ�VUP�͎
#nDc���0���ȓu���Т�1�Рxԋ��B�J�<�指�$Ҏ�3�Kh|Y��B�<)��ݧ|@�����E�D��v�<��胹����g��>6X]tg^n�<a�B��m����w)�C�ɟ��b/��C��Y(�r4b�O�����7� ���I��&�PU8�.�x�!�F�3@(�Q�K?<�X�pG+1��	@��̫7�\�Mİ��nW�_UTyKa
-������~¶��k�%^��L �f K"1m�O(<���S��3F��e�h`WGK?i����n�NQ��N��a����$�@=c�C�	�EP
���cJ�z�̀�C��_;J���<��'����O�3�I9Hj)�.@P��5��8<�DC�	� �y�cbN*B�{����M�C�	o�������9��%Bm��Z%�>��)�#Q�����g�^,ц��[!�Q/�$�p1��6a���F���!��1&�̉�"��'�zDBcFM�	!��H��Q��Q�qc�;�$�%7c�'�a|�O$�4��&�Et�2�	/�y�F\�r8bf��st�4�p. �y�G�2:Ѯ�15�a�2,@�I��y!U�p�n��7��3Zcb@c2ب�y�K��*��U�N�`V<������'�ў��ȍ�E�Z(
��2�Pc"O���R(�/(�z���_�{��hB��0L��x��;Y�ȍH�*W��4����y�GO1�DՃ ��2�j�# 3�y"GL5~X�"�<��H��yR%�|����!5��H�숝�y�埕t�\�ƥ�GfU!���y�&֗���9 �O+D'��R�b�y��<s�|y�T
E�?���rʔ0�y���lV(-����%ېP���	�y�f<V��v�T#�����2�y�윖t}HI��/0_|l�e���y2'   ^"���*E#h�RqoI��y� �60 ijQ�>�>���H�yB%�s��h�V���=�V�Rd���y�G�7<0��!�mS(*B�PDB^��y���xQ�D����a��Q�y���9P�Z�����ty�F��y�M�'e�\���R"����w���y2�.+��LyV��~�@`�!B��y�b�2���zb�3.qj���)��y�C�=F�o�#S88Y6�Ƴ�yRE�t/�@��<U@����U�yr�٩,HY9�#I4W ֨�d�ݰ�yrB��Cl��uiO,{����ʑ�yܑ*vp3%'��K��P���	i�fO@LD��0��ƛA(��ȓl���ce�}�ZP pʘ1q�Q�ȓ4 xI���c�,��D���A�ȓ *�m�(�� ���
66m�ԇȓAW^�2e���5A=a!�� ���J��!���l��������S�? H�ق��"c�����s��!�"O
����M��HP�� +t���1"Ot��c��'O��	�B � ��kg"Oa�4G��T���dI�$2�2�"Ol��Q)sN�c����'#�-�t"O k���,b&��5<��t"O���T�#$?bl�g��1��� 6"O� �pa¼�0|Sp��03��Y"O"����|�����V�	���%"O.P�b�ۯ/v�����k��c!�ڂ/ov�AFl����I��+@�6�!��u��x��d.ƘUʏ� �!�dW!=~ �����]%0�(��:�!��C�j�C$)Pa�G	�1�!�D��w�6���p���(���C䉆��x���X�	�ε�b�EV��C�ɷ<}��;0EL�j�	I3(ޗW�C�	�|���v��g��-���APC�ɭ\���C�͊�4����˸ PXB�I�(u"���dDP_|��R�ɋJ&�C䉊5���*���T�DmKJD|� B�I�t�xMz&��8�.ٺ�IA��^C䉡/�n�.6d%*e�@> }���sSD3¥�O�q�/	=z����ȓp�\I�E�P\�сN7n�� �ȓ4�zPP� ,"�|����.]�(��V��VE�$��2�%
!}��`�ȓ�2�36g�"v,��*		W����t-jv�1�2����񎔇ȓk��
�eׂ5�����J��X��Yv���N�w�
���Z�;{X�ȓg�Zx�5�N3�f���#L�%����#�����J�J�b�{�K�3g8���Bq��t�	�=�N|k�H$fK�H�ȓ
�B�Ba�D5r�(e٠$�B��ȓ\}L��Q
K�G^��Xp��#��$���8-Q��جJ��U�¢n'�y��`��@�#�^!v$�7e��(&���K�ɚc� �N\;g,�<a�$����,��Ǡb\�ď��s.���S�u��O��^��=����?q]�݆�!.���U���җ<:U�Іȓ�6���	���R���;y��L���������h��e�tQ�ȓS�H�2�c��Y�!`Za��)�ȓ���)�I4�"7ɔ #��Ԇȓs�~�#�/a��┘U�|�ȓO����Ȓ��)c��>Y.�ȓO��|��]��`q��5�de��k��x��LāG1�LI n�Gp�X��\�V5kd�L�6�:©ݾ='����\�T�؁ŃO��P�$�Y�?�Lx�ȓ���ů�*~Pek�f�6;�D��ȓ1����`^�zt�	[u��(�>��,3,=i�ą�\�*���-�=��G(a�7�ݑ+���2M 0��!�ȓJv���I;�q �ϗ9kx]�ȓ�4hr�"=C��A�Iʑ=͆��N�|�H�j�hD>�����^��ȓ5��{���1(��v�˪d)�ȓ�Pm eƇ���T'$i����y(�13��3\uT�iĤI H��X�ȓp�<E�V�-�0A�MtK6��ȓ�6�A+�T���KW�ü=�~���S�? P�k%H1�輣�+C�B��"OV���U)%�"EhD�Ow�l�'"O����OB�UVE���!�|Q�w"OD%Z��l���&�:k�<tH�"O���0k�����aH ������'���ٟ����	韨�����I,tvɲ�NE�E����'�|�I�`��۟��	柠����	ɟT�ɨ =���V�Î[�`�Ƈ�*N-vd�I֟�	ҟ`��֟���ǟ����X�ɕ#ﴠ�w �4#p��螄p}��ݟ8�	��P���$�I����Iğ���_�
 �t�M!���b�G��]O���I����	���	ϟ�����P��ߟ|��9}B��a7�Q�l$X�����z��$��L���\���8�	����	��I�0P�ea
1� z&�T<}8���ڟ������	럸�����������I�PA�q�ӧa��]+jD,�������	� �����I�������I3�$AQ���-B�m;�W�8 �9���,�	ȟ�I��	П����I(c3�qS��^�B�@��W*�=_'(�����	����������I����I�)u�T)vB<";��fLħ.+RT��ڟ4�Iǟh��䟼���@�I�|�	�w��)�Ɏ6(��1�M�ff���	ן��ş����d�	�h��ϟ���	V���6f��(�,@+12>�	Ο���ן��I����ڟl"ٴ�?9�}D�K�n H� �ON�-�QWT��	y���O,�n%�^L���ܮ*����EK�0�RP�"�%?���i��O�9O����-t<���C$m����EL�d�O�$r�r����$��$�O_�h���4j���RɀF�b0�yB�'��V�O������^�q$V]*B=h_�1A�l�f�s#��4�Ӟ�M�;U�"M����-V0���L* ��P��?љ'-�)��8'y ilZ�<��!�=�e�APht��d��<��'�$A��hO�)�O��Ѣ�АsaZ���v-���0O˓��ji�&�2Ę'������fڶ����"${<�����e}��'��=O,�)9�<���Єum�u�Q��Ar�$�'���,p��,���#��(5�'�F��7gş ��=��L؍cT���]�<�'U��9O�Til�*�~����Y;��q�:O@�l�!x�x�=_��4�F|	�"R.r�����X��-A7O���O��D�>Y~6�(?��O�B�	��|<� ���f���``�[�3}\qI>i(O���O����O��D�O��G� ���[r艎K�~��pį<�0�iG��;�[����S�ߟ�qGJX����Aȓ�c�4�jQ��DLΦ0�4g=�����O��t���<siZ�CZM�d��=8&И�iB����ZX���1BL?�I���R�a1��icr�k�b�=a�d����؟�����@�	՟�SOy"}��	g%�O�a��d5���A��9v>]Y�$�O�yoW�{��	�M�R�i�47��J>�!OE�v���� _
�)C'`�6物9U���̋#���B�<�+H�����VQ8l8!/�6g��1A!�U����Ɵ���֟��Iџ��	s��%�j]#��Z3X��P�Lު6	��y*Oz�����4m>��	��M�M>Y6iAD>*�k�Tx�.�d��'J�6���i��(} �l��<��f�A9��K�5�*�A�^�-����臬rO��D������O���O���6�:����$�A��		�~���OF˓r���PA2���ЖO��� ��P�XsF܀�oD3o޾���O���'~�6�Ҧ� L<�'�Z!'�*?���y��[�1�H�`C�?r��Z%Fݓ�M�R���S�1��D,��ol�J�G}&�Y��1>mV���O��$�O����<�&�i����ƀI04 ��
�U�~(�R�.�&m�'D7m%����$�ަիF(��M~mGte����	��M��i�u���i���O�`b���R�o/?C��4T"���ڻ��-	��|�@�'���'bb�'��'Q哚o�� `�`RV!�9����4���4|9�H:��?�����<����y�R�^d~Y
�Oڔ%�F�:�ʐ8�(7����N<ͧ�r�'%�f b�4�yB.Dh�u������gj�Γ{�����On��K>�,O��d�O��qSa�y��P�����򄬩���O���O��D�<1T�i@�B �'X�'��t1�QN�|1�Ϸu���s��$�^}2�q� �n����]B�)R9�Q�����J�Γ�?IC�
o��Sp�4���
�a��R�F��$m�"x�)֙c3�����N�d�O4��O���2����*�V	XTJ��P�L�*I�vL��?�7�iو���Y�d8�4���y-�K�)�5KJ3Wߪq�ACP/�y��q��LmZ#�M���M��'s����-��'j��<�u�ʁ0M�p�M�-��L>�+O8�$�O��d�O\���O�0	�EȚ'�S�i�I%�h����<���iw~9#A�'T��'���y�C׭���'����yFJ�.n`��?Y�4S8ɧB���br�D<	�c��sօXKE�NP C1AК��A�Q�xQQ��Fk��O|˓˜L��`��U���"fCY�}.��j���?Q��?���|�,O`ql�Y�z=�I4)�x]�w@eY�����4lK�;O|�og�M��	��do�4�Mۢ�s(=f��0��5��y�|L��4�y�B��V�������?mz�8O����he�=� ���^��Ea�M ��8Ѡ:O��d�O����OL�d�O��?��-[+l&�+g�
�\�H���-�Jy��'3&7M A����M�����^�n��$Q���!dW�;�h�~y�'��o$�M���*cI��4�yZw���G��e�H�B�@9l2Y�g!�!Y�x���'�&�|�.O^���O����O���!˦j�n-	�=I�]�Aj�O��d�<�ջi�dh���'��'��>U�|��� Q�i���I���n7��S�ꇱY��P[WCB�u�2X��+�z�~P��H�
em�&ȵ<ͧJ�\��y�ɢk��y��� �Iy�N*�t�	��h��ݟ��)�Qy��Ӭ0��&~�HI�cnG�

�I8CË�a������DF|}�ak�l!@��P�>�J�C����3�A�֦9�ش4k�iߴ�y��'�,�f�Us�,OT	��f � ������5��?Oʓ�?I���?	���?����) ���}�7��շ���m�Y��ij�&�'�2�'��y��l��&4XdрS�8�˄�X'3�mn+�MӴ�x�O���O̬*�it�Č�6�2HXW�T�.����D>>󤃄85ڴy�o�ؒO�ʓ�?	��S���r�.�'E@wc�����?9��?q.OvhnڛFv@�I� �I�	C�5�5��&�%��h��w��I�?�T^���ݴ}���"�>��������'�<�I�"���O(�V(��h��Qͽ<Y�'7���H��?)%,K+Q�$ec�6p`��e�E��?	���?y��?1��i�O&����0o#ȸ�׋M=&�2u\0�$���q���Zyr�d����,=l+A�r�P�1�m�,T=b��ɦ�1ߴ#'����b��=On��Ή�T���O��u؆���]r4�9E��;I\�qs�|rR���	��X��Ο������wg�3��3�T;`�N
$dUyr)i�J��p��O����O��?�R��	�P�Ԑ��%�/?�@�V%���T����4cՉ����O���Z�):>�P���)z0@�&O�(:��Z��E�=xbO�y�Sy��W�.����6f�_�X1�,\�&F��'F��'��O����Mˠ���?��!����Ʃݩ"�����?Ɂ�i��O:��'�¾i�26�$(�ҭI4V�5�l�#�ݣg-��Qw�x�4�	ٟ{d�JZ�dh�~yB�O��
�0�,`��K�\6l`A3E�%�y2�'�2�'L��'���iJ�Y�m Sa��B�N��V@s&����O��䦩�t��Ty�"d��O"];Q�צ�c*R�+�|�XbRu�I<�M�ǳi�����s|��<O���ҵ^��4�6I	�|`�h"*��q"����?�&��<����?y���?Af�^B��A�DW$N:vD�����?�����dXЦuh��쟼�I�`��?���	�=�u"� �I
�!�a"'?��X���ٴ`q�F�%�4��I�;U�A��c��s�n(0��88��G%=
�HCǪ�<��''���+��L:T�2@N��F�F���u��T��?���?��Ş��DĦe0�R�Jo�lV�.+���V�I�,��'��6m7��-��$��is�"��Nh!��)�5h��r�թ�MK�iV�x�e�i��D�O�|D������<1��D�e��3��O�s�꼓4��<y.O����O��d�O��D�O@˧.�TS�*!_���%l�1tHdx��i:p )��'���'W��yr�o���]��CW�S�+F���#{N|m��M�t�x�Ou���O��}�Ѽid�Ĉ=�1�nC"bTڸ`W�~,�d3�(��t%�O
ʓ�?I�WE2�����t���"W�QފI@��?����?),O��oZ$kBܗ'��!��u��u$�$y�u�6J^��O�'��i{�O�apR�˦UHe��@Ct�S=O�$Q�bT99�'�:�@˓����O��Z��%�A�>��L���1u�� '�������㟀�Iş�G�T�'�<��n#
m�ݛ���,!�I��'��6�DS��˓` ���4�P����ݰo� �d�Tk@���8O�o��Ms4�i��ƹi6��O@�`Ҍ���Ŗ2	�m�$N�)�Ht�"�)@���O@��?���?����?a���X�a���^.��	�OibT�)O��m��i�u��͟���A�s�x�1ߧN݈HTO�E0�Ǘ����̦AIݴ	������O;��#[L����+A6(-��٣�Z|F���Y:�� *j�e�'p��&���'`yP��Z�X����@�U��`S��'V�'������W�`r�4a��,Q��s@0�j�.�'2�b,�j������'��'��k����~��	mZR��0���9!�v4��厏]�b�sG)�Φ�͓�?�+�!���釅���䟸��N�R
,J���H�}�7���e'��O����O�i\��'��hy���zv$ȕ�^�.���"�O��d�OB�n��6@��'�6�4�Ď0*^V��u&�Ȳ��$��'��شZ�6�O1Vp*�iO��O�3䥁=�v�hՍP�nn�%�(J,ܣ�'��'�	�t����	<�֝���&m��T��b��p�I����'d\6m�&�E�'���'1�S�?.0ɘ��>n�f �� A�mX�o��I��M�ѷi0�O�	���y�@''�:Ǉ�\��A�5�3٢@i�- t����C��O�UhL>�0j��i^��i��_(Ҧ@������?9��?y��?�|�+O�$nZ)}T�):�/��lahZ�/��9Úcyboe�h�H�Or�nZp��@�ah��c��P�[�����4E6�&O&�v;O��Ē*s�8�Oq�)� ����%�4ֈ%�0��?��\��;OJ˓�?q���?����?)���?iMI�|�:�Vj6��2խ��Fl�E/9a���.O�ܦc>�`�4�?a1.^'Mv�C�@��i28`�"[6⛦c�<$���?M�S`�d-l�<�d�<o���B�.̽	}�����<�V
�/J����H
�����Ov���/��E2�K��Vyps!�.$���D�O��$�O��H��&HҨl���'����o�Ayw�BiE( Շ�^[�O���'S7�Ŧ�H<i���0��e�H�%JЋ6K��<���W���0pa'u��M;(OR�ӄ�?�7��O�I�3��/�Ҹ��b� #�Ƅ"�N�O����O����O��}
��w^p���P f����E�5o`��!ۛ���	W���2�M[��w��0Ư�>�9#ժP%Xp �'\�7M��:�4v�I��4��$�!������jp���/��Րg��
+��"��/�$�<���?���?��?�b�\�lp�pB��,9��Ӗ��$Iæ1��BIџ�I�L�SG��'����?x�F�*� ��0yk���>�%�i+�7��f�i>����?ɪ�A^<����5���Ť{�R���LayR�ߪ�����2��'���$F����D��Q���Ba퇗1z��	ٟ�����i>=�'�6-�#�"�$ݓm�
E1���̚����e�?AfX���	���cڴD�&�#&�˥5i�h���X�v�1�۠�M�'6t4+U�%d�8�'L܆K%�O�4ט� F��tO�VPI���r�f�	ϟ��IɟD�I�����s����AQmR s��� ��C��)���?Q�Z4�v��e3剰�M�M>�".L�l���+5�qk� "M��)��'b�6����ӭM��oZD~REܾ
������V�s
��[>�I�����!P�|�^��	⟰�	�x�U�H�fji�0cK�u�"x;!�Zڟ��Izy¨a�ҡ�b��O����O�˧4�Ҽ�2�-<.��#�X� `��'l����{Ӵ%����?��HI"F��ru`�$	a�Y룪ѭq���U�=W�e�'�������&�|R�
�J^����%*�Բf�@+M�'���'����_��۴m�5�R� ��aL6��q��?1��k���d�F}��hӬ�1��7�	��e	�&�<X�L���޴D���ش�yb�'뺽*����?	�EU�4kv��4~��X���YV��``|�@�'��'���'B�'哈U��KRcX�x���	2ǈ� A��Yش}����?����䧽?Ѵ��yg�K�q�n�C'�G�:G0=�Q��,;�6mKͦ�I<ͧ����)&A�۴�y��G;=vȘÅD�71Ѽ4Y���-�y�̛\j<P��� �'k�Iȟ�	�W�)�b*��y�� �Z"�%��՟�IןĔ'R6���zV����O �d��XA�p@�Zj�"ǀj�lوr�<����Ms��x!�a�Z���m � �!P�@� �y��'�H
۩Mi��*�<����F�	ğ4)���B� �H�aĩx��D�&ߟT�Iğx�	���E���'��PRW�Ʋ�А0� ;2�	+��'�<6�\�_b˓hh�v�4��x�h�g�������"����O�7�E˦I�ߴ�^M��4�y��'��i����?�
d�9BZ4Q�#H�|@H����΄G=�'B�	ϟP��ßP�	۟���1vQ�i�aD	+t#�`5��-��ԗ'��7�4f���O��d5���O|�����a��".�q �$ �G�\}�n�b�l����|*����EL�S��l��+��P�
� ݂,{��wO������0
�����6���O�ʓ^���a�� 
w�E �.��7޵)��?!��?���|�+O\o�U����ɾ�^�ᑍu��e�7e֫D����	�M{��>�g�i7m�ɦ�@��]y��re�`w"� G+Է�,�l�<y��:�z���h����/O������=y��A?W'^(8�c��&���Jt>O���O���O����O>�?��G �'`��	Ck����A�bJ�Οx��ß��4~���)OL�ml��� ��V&�Aī��c��P(I>Q�4ś�OXYt�ih���O �0T�˥,�3r�ؑqK<�0U�ņi�L���$��O���?����?���xt<���x'`�Dʳh�4	���?).O�mZ7Lfl���<��B��8��p5��7f�@٥�����{}��~���l�5���|"��H����s��,	�8�*҄ũ}cE��	!�l�bjR������F���N���O��4�؏}EΩ*L��9����e��O���O���O1��˓,��&�I��r-X����St�s�d��_�%���'҅pӎ��q�O�AoZ<��Y��"��Z��P���W�&�,�A�4_��V�M��'1")V(xab���1^��I�=N��Ӻ%`���3�6�IHy��'r�'7��'�RU>��+s5R�h�%M"Mb����M#��¢�?Y��?�K~Γ[&��w�N��f��]�궧 
=	�@Ӄ�d��1l�����|2�'�ZD䕗�M��'��%A��֚5�,9�j<Q��ؚ'Kl�Z��S?�H>�(O2�d�O���)A�}����G*֕d���'��O"�d�OR�ľ<r�i�t�*��'���'�N�C�"%_~�;d�כZ�*ͫ��D�g}�HzӼ!n%�ēQh�H!�ȅO��0��'�;e���͓�?��_��fa
Ԉ��������iD�D�4@Z�ЀJY�
qx'�֜n����O����O^�d*ڧ�?�Ō;l������N��I��o��?IT�i��I�Y�d��4���y�CG�d���ӧG.H�X5H����yB��Ox6��립��k�ܦy͓�?Y��R�:]��	�M�? ��B�5%�.�@A��P	�y�F�9���<i���?1��?Q���?a�ē(X=���~�:@��X���D�Ħq��$Jhy��'K��e�W��C��]��%�536PT���tyb�'֛��:��O��$�OkҰB��[FH`���V�= ̳Mþq(gU�H�V������*��)-�uГ�IX�P�;��O�=��O\�9m��8$�H�s��ܢ�1D�lx�� $0]Ft�##گ�D����;�	�y��l�	�Lj�����G0W'T�8�j�1��`��K
�nk����e
C 8�di�	���H�'Z�E�RW�٧��3�P�5�U�;1v�A���w�&�ѳ� Ԃ-�@̇-,*H���'�\�a����T�"b�!%]���\�.���c���L��1�Q<�Rxl��Z��r��^��ڱ �!خ�Y�O����O��O����OUʴ��ON9	Bk�2F�m��Eьc5�A�q}��'��'.�*+���I|�CΆ^��̨�CL1|/������iכ��'��'���'����'�� �*9���W��hg@H�m�x�IAy2�OC}���d�
9��HJ��EҲ@́[�&E��Xt��؟H��>�`A�	`�Ip���ǌ�� b���v�l)D�զ��'�T�J�!i�\��?��'sJ�i�%�v��?h���c@N�k�Ҹ#A�r�,���OlI���O��$�O��?��T���:Q���&JМ��DL�~�D6-�&F�nZڟ�	�Ӗ����<I�'��N@*���? :�=����>R
�f(N0xW�'}��'��Oq"�'��F�\33���p��	
E%�=JRE ���	П4�ɸ ��ۯO�ʓ�?I�'�
]p�R>'¤��A�En�3�4�?����?�cBX�~��������۟H��I��	��F64���JR*�dK"o��*%�Ҧ�ē�?�����{�EEX������0Cv�@0�Uo}��Ѓo�[���	��t%?�0��A6�ZE���f�Y-�(Qj���}"�'0�'x2�'*f��%Ҁ=4��j�F��c�]JB]���I���Iuy��˽:>��U�~��ӎљ
Ш���LOK����?�����?���k��K��W?��Hbf��ԃ�㎎ah�u�gR���������~y��Bzx��?Ab&�'e�`�F� 0b��p�S�,���'�	ş`�'�f"�P>]�I�ϸ��s L>,P, � D�'����4�?a���?	���t��W?�	؟\��;>�$`R�jL�C����GI_/t.�9�O���<�@-���	�Ol���?!0F�V�WnR٨1@�CTx@�сs�J���OX�`��Ϧ��'lr�Ox��k$Ǳp�<��"ͭk\-x�#U���Iß`Q5K��I˟t�	Z�cr�C���e*L!i�-\+:�)�4s��Z��i`B�'f�OÖO�)�A��)"�ֺ~�V)�����mڥ)gzh��������h�m��W>���Nj�pił�%{J����ż�M��?�3�ཐ/O��I���# b��``�� =4���#��L�O�������./jQ�J�&I<���+�M�l�H���Gy��~��B�?���Xŀ��aQ�@5w�7��On@����ܟ��'v�C�P~D�!^�C��e� 6F��m�W�D�	����?)��?1��[(Z�$��G��l҄�V)g�4�ۈ�')��h����s"�_6S<�䒧�ϡ�6�������ڟ��?Y��?A���]}򊕘h�>��PbY�>@@%{�Oŧ�ē�?�/O��ŧ4��ʧ�?y�U��p	V�״ k�x���"2��F���O���ւ*� �O� s'��K|��*q,qi�#��I㟀�'` �bc(���O���Ƽ�#Lx�8ę��N�k�=`��x"Y�� #�ӟl'?=�'d�LJ�J�&`भ�7�$ �bL�'#"�U/y�R�'y��'��Z���07�n�S��N;�(x��P�<�`7��O���G�\��b?ɐw�1,�!0�=)8�ȉ'IxӚq3�P���IΟX�I�?��N<�'J݂���_�W't�SCڭN\4����i8H�'P��'R�O��s������+d�̴��h�
_����rΟ�&z0��'�ʼ�2y`0���b� _�ݙ��Fv"
���3W�lx)D������6e5'I�uJ��T�@����vo��2��9K���ŉ���м��g�)�OO/'L�+�䝱?)�l�숎,A��Q2C��Te��[�a���hS�_3<h�皿+� ��.�7������,�5y�#�y0�	�"�0��	ޟD�	ڟ`���ɟ��I�|��dЍ?Sp$���� p��#��\�d�ް��ݟ��%�Q�\�Bp��DV�N�X�f�JQm�����PXt1c��~\��bG@8n����Ǔ<�u�	��M�G�4<�M�0��<V���DbҼby���dZ^��yB�(���n�y_��"�y�b٪@"t2fa�<6��f��y��>9+O6HC�d���M�Iߟ��O�
p�CD�:e�MkƇܥps��▊B�2��'2��_�� �[C�24`�kT�K�$��O�jY��܁t�vi��� �lo�4Î�D�]���Yb
=�6c��;iT�'!NB���)X6ɂš�	@�HGy�a���?���䧡?9b�rV8�y��KL���r����?����9O0��6k@$^АYsV-<(S$`�'�O~]�)�|T��*�?q4�#�<ON�[�Mզ	�I��<�O�X5�'���'��d�Ȇ�d>�٥,�"����H�=�l H��{�^�ԧ��'��O� ����ԭ$ܜ�3�L3E>܃&K[)���:�/�&#��J�O?�H�$R *�q�x��5�	����i"��OZb�"~�	*hu�l�g��}<��,&C�5J��H�����1.}����v�2"<�$�)*G!OV=�+*�����K�<ivG�Q�|DK�G"J�����`�<1�HXc�ԑr2큞8����Y_�<��fW���������kB*��\�<���ڂ4�!�D�iB����D�W�<qfd9qH��R�P��=�F!�L�<��:�P�Gg��S���`��G�<a�G�J� XA@�^�^A����G�<�V$�8iF8u���GCT�`#$�]h�<�GOO?��< �J
�\V +��a�<1��ۀX� @:�.۴e������`�<�6�ҟLt�k#�
e��X`�r�<)DLK0[Q�=�qB�{�RdrQ��j�<�^XS �D-fuz����>u�h�ȓa���z�Ʈ+���	��&\lΡ��u^�d�S�ͧ>6� �Ӌ��~p��0_��*�Eǲe��p��]�5����%��F�3F,^�]¹�ȓ(��cE��,)����1�B':��ȓ'�
)Y�%ٯnL��PB�~$�ȓ�U`�.��<����8�"O�q�F/�X��)P�T�����"O,��Ӄ��F��I�&Ne��9��"O��â˘,<��waA�i����"O���"ۍ	��̉A'�XJ��h�"O �,E���i`�"5y(�i���y�aJ& �� ��`�3% �Cdc��y��W��ճ�>~��E��y�"ݏj2J��0ꋦfFN%�b���yr�'Z3ZQ�gƣfK�@rE �yr��3{�(�JT
�Z�����y��ɑ{�H�{��E�Q�=��ԙ�yg�0H��Òk6D�$��3a���yR�)H�HsS�^�5����w�ؓ�yBf��v<��V#L�`�lI��O�yRN�AK8�����Q=bܺ7mT��yBgR
$p�XQ�fF�P&��ö����y�eŖ�R��s`X-=�0Yj&�R�yi�J��4�P$Ω+'��K! �yb�&���(Z���Ӂ����y����mx�t�%�PC���F]��yH�8�84�-��ҽ��c��y�
�zx+�.�-?F��#f�y"jK8�x���	�2�y�֎�y���w\p�E-ājy
�Z�L� �y@^�6x���"�4��������y��ԑp���Q��%e�@�J�y2�W����-�T�\�3�kD:�yR�A�\}B��3M-�ݙ���y�e��	�g�I�H"���Pl���y��0V��)Qh��>ּ �"��yr���$N=A5ِ0Z:��r�K!�yB"�75P�ȴ��!�@4�2`�7�ybW�W3�u��n�R��R/��'F(SR�2S8ҽD��-�Lx�z���3*�����y�n�)��"� ������k5yl����B��	�]T�"|�'���"o�?�rq��A�  Te��'Ѹ���� �)�ȟ�����Q���uP�1�{��0�>�!���B�AYvIP��p=񷌀�Ж\P.F؟D����Ĉz%.�9-�����.(D�� \�0���<����@�F2
b�S���VD�b�Q��E)i.�}��l���(!$&����d��	XC�<�3��0h�F�"dI�Ϯi��g��~s��rc��򄞾%
>�snm"e�ܙYv�͛�`�Ʈ,�ȓ,Df����ވG��)@'� ���Bl�<L;�z��"��='I '2a�DÞ[I��FG�gX��9օ�`�)+>�� �C���&l�A�N&�y"�]00��ގf��<+�ֺ�HO�\ ����h�V�SR��C���3��B6ȣ�"O����y�~��K]�q��ȁP�iS"��%'�o�S��M����Tas"X�i^�qS��h�<�c&�!WlQ���ܼFx�D��Pv��}���i��Q���V`OR]QC�
��z��R� lOh\C�hI��J'�АRi���/С	A�(�B�Ԧ[%�Y)I��S
�.�$d+j��_�f�hDO)�~T�>QEB�_պ]���P�5�~�����'�j��	:S�t�� ���M�x��	�'�L���t�vT�0�x�\%Kp��$X<BsfW�N���	bӼ`@��Y�)I����^>�$���"�;&R�{Q��[؟8y�CO�P���+e�G�"`��Ytd���1�4P���	R ��Q�k� qf0 S�F�@��!ӷ�8��է'{�Y�S͹��0���QmQ�|x�o��y5Н�����A��ю�O^؈���{��8`��Kݺ�`앭��'�.��)7�J���<i��P�vi""N
j�0�NSW?i��X3Q�9RT#�95��Rs�H?��̙�:�L��ҩ��S���K��!�� �n��>}�Pڒ�&4���&,G:)..�!��b�~�#�DE�(Br����z?A��jZE�/�$wWP���A��s�:���"P�ADj���o_�_�����'=�m cL
(M",H�(�<V8�D:A-�8#L�@q� ʒD��b�gE�3TB�1�$G�"-J� ���E8M>����=h/�R�e�u�S�_v�'�݁���e�*IRb`@7|��d��0�Z�� �X9P^$���M�%�$7�E8kR
� �Iʋ=�XQϓ"���+D��.8���G�2��'�z��q�ɷ�Z�+��H�/��|�O>��צT�'
}f���wdT�1�N�)Uʠ�C�:�JB�ɎN�<L3b� ݢ�{��"q���`��cV�	��%�[?�1b_�&��t�)����g͌f�����:#`drc�x�<Q�I�D��E��;�޹��dE�!K�lٲH����72�I��D��[�)��p�Ç�	���1QF�_v쑆�	t�ʩ��Þ���f�Y�8��_2;w���*A�;6����+)4��S�ăC� U�X�p�O� )�	�{�Rizq�4�']��
���_�f!j�l���q�Z�!P M�j��2 ��l�MlZ+{�
�+R��s�h5*��֒g̾|�e�n#6�I`"O���)Ki�=���&����^�H�T�ɸ05�{B�P�"IV�R�z���K��G�>��(��v\��$F�D?PcW��@�CF@֚a9!�Jr=�=;�]}0)�Ta^:*ב�P�R-�^K�>�t@
9D<�ȅ�T�[�9�);D���sI*P�2�ҤӦi�j�r`�e�.hA�E��������چaD��suo�*-\x-��cV;�y�kM9^L���hrI��Ί���d�x�D��-+B!��F]�V�`	1���Y��u��I9G2n���'$n���@�2�0�aX/.'Θ�'
A�2dA�=y\��#-��r���2��䅩L y��	$?EjH(3�3I��PN�rg!� n2ܱ`�N��ꐓ_���]�{�LX�=E�ܴh�&�ց׌#s|`�%N՝*?�����كN�x_|���ޱ*��(�'<�|���'����׫wO�m�1D�c�����'L2ء��o�l���)��S�'Y�!ÑdP<�$����wm��y��Ip�%;�Q█b`��!�yҮ7�D���J9L� q;��,�y�\LLEZ���K*�pL�/�y�ĈA��rԩ��N@���f)�y�˶Jtd ��M;I��10#0�yR�H&B�&�)��>�^�4�y�]<�
��a��f9`���޳�y
� �(yta�Ml���L#l�m��"O@�ѲaB7AR��BCI]�¡�"O���7Μ7����+խ�t�2V"O�y�.�A3` ۖL���݋s"O,�����	(q�ņ�Ȍ9"OH}z�A����h+�� |�8��"O��`ή1���Y�d�Z� tP�"O�\۳��e̼P��@ج��A��"O��g!��9�RAW��� ��1�"O�����"bBh	�-�
u��a��"Of����� �/a�Nm�"O@d�ꚝm�H0ӥ䋸%z\h��"OVH	T��.'w���D �JF6�Q"ORܢQU�H� �H8���"Oh@��ү~�*%&�-!R���"O��W̋�,o6�Y�,��	d"Ol(�/��Z�tIժL�H�=��"O�ݓ�䔡O+\�D�� �$��y� �����[�6>.8(�KG�yR03��$*����'��[�	ޡ�y⢜�s�`*-���n�0Č,�y���xEK���J̘Ӧ���y"'��w�T���)�$����<�yr��*K�\�H�2i)"o�:�y�ʭN�*���<R)�L]&�y���m�R���>�P��h��y����_> �Y�V
�(чل�y��CKl$I4!�~���4�y<a�y�&�&8�9����y���'���QK(`����U��y"�޵��m����/h^�tٶh[��y�-�|�6�KW늓*�p��P&���yb���Q� ��-��R���'�y䆹-B�yӐ�M .r�(d԰�yG_+6����G��~9 
$�C��y���:c��NH>he���y�f��#�Ip�m�,����y�B��VMīW�C�f�aÀ���yR�$ֈ� K��;ʞD�RB�9�y�n	�ʬr���!=*�#�(_��y"�L�\�`�A�$�fU�D���y��
7(���BQ+{�zQ��:�y�H��[]����]��Xk�=�y�ǀ� ���P'[?$��� q�Q�y�C@+	�5��K-kMZ5�͟%�y2!����)��K�K~������y�&�JV���B]���q����yZP� �D��t!"T)���"C�Ɂb9��xS	G��ݣ�v�$C��64����Λm����s�f��C�I�R�rm{pN�W&��ifi�	<"C�	� �P@�g�D+1`ŋ4�{UC䉦P��С���DYn�?V;�C�	�x��I	6�� TI�u�P�~èC�	#Z��a�M�H7��� ǟ:z��C�f�E:�+�L�!I�_QC�C�	�r �L�`�X<�,(�C��7:82���@�.�F����6zC�I=X�hF@�*h��6�V�j{2C䉍`d怣PjJ�)����G�7^C�I�t�� b©F#�i%F�O��C�I���c��.����DY+ǂC䉋]
�bD�Ǧ[�~Io�3Sw���ȓdl]��&�<&�yg��6f�H��S�? �C�mH�B��{��q"OI��`T�2��Lp�"O�a�'�� �r�ل@�T�V�S$"O�����B��
E^� �"O��ឥ_A`a���P��<��"O�Q"_�M�!����:�&��"Oҩ	g��J�05�P/��h�"O�TU�ا$H�:���l�ĵ��"O�����о3��ſw�\D�"O8Ա�hK5�
�&��L����"O>:w�J�sXr�EɧcX-�"O���eoL�:Pes��Te�C�"O~X����!l�촩f��;F��g"Ot�+�N
�HRm ����Y80Xҗ"O�!�"�O*���sr�R,Na��"OݓTK�BT����˜ �A3�"O>��QKP;<4,��ᒖ�X�"Oh���ÒH/ ��P ��v<ͺ�"O΅X�A�s/.��#NJ�2H���"O�����a<r�,W�5��c"OH��䎣|�(�;�I��0Jh�"O2�j�,_<A�z00�G	cW��p"OH��e�9]ʄ��V��[4R ;�"O�(Ś�eV4�(�Ћ#�Ft��"O�t���*0VY��蕤ɘ �b"O(����҇nl>����X�b�T��"O��(û)|.\	�,��	�j0��"O��A�腰L{�D)UkQ�`�c�"Ol��*�3
��`�	E�T`��"O��SGB�ma��S�G%�U%"O`�X���KP@�����/0x��G"O���p�J�@��FB�]v�"O����dޥ7��ᅌW�ez
�@"OR�el��d`�X�ą(uU�t"O�逕杵t�Nl�"�6qY�s�"Ov��p��r�vpd.ƄlV�] �"Of5�O���}��.�9��"O�{���~�Tl�����q�"O��Wj�/4u8�B��b�K7"O����Ȫ��y�S�g����'"OI��U�n6&� �=u����s"O�)1�ω'A��I���^�0ؓ�"O��Y�d��]{��rn�	�`i�"OVt*�ˋ*�P�mW�Q
�� �"O�s񣃒b/�Ål��Sb�q�"O�����n���Q�LlAn�V"O E�udԞ~2ȀG�w"$D`�"O�����<q�xcDmXsx(�"O�01���6���d��lb�Cw"O�(�#�"e T�`oY7EX��r�"O^����ҖBRHre�I.�0h��"OL���8����E��tk^iKu"O&��Ƈp�m҃�
����"OЁ�p<]l�ԓG��f��9�"O�J� ԟ4��[A�"~ŔXA�"OV�Ar��=;�U��1W
�͋U"O�x�����r̆!���;Ljd��"O��e�	<���AAŸP��E��"O��ۺG���q���6�B�8d"O�$r@�ѻ^��`��Fz�
#"O$�"ed�-~��bD���d~��"OΈC��\ jnh�C'ׁ;��u��"O��V��(i:-��ƀ�|%���`"O��c��O/c��r��;j��Bw"O� *�j�E)��xDS**�ٓ"O�\k��30+�Z��W��h��"Ob ����
ir��Y�6���"O�P��g�*^<�D�=P�p� R"ON�і�߱LAZ�ȕ:\s��y�"O8}EK�U�M(Gk��"O>��6㝸'.�V��HS�H�"Oꀀ�kUM�ipb�rƝC""OX4��r���i�b�(NS�� 	�'�p�� �ʦJ�$Ո���:W[Ą)�'���[�ˎ���1�B�NU�Ir�'p,����_�hse�M�K��@*�'������Q\ ���сm�����'V�i�#�w/��0�L%̴���'bd�aĝ�c�R����Ŏ �U�
�'_�4Yf�o ޥ����.%�e��'���nT�*f`( �� sJ��;�'�aᦩ�� fm���d�✈�'Vt����);�j�H�%����'M�U��a�'.���&iS��4)��'E�H�GHh�q��J���6Eh�'�@s5�ҿ%� ��&N�uZ����'���$�	BJ5Q�h�'�l��'�1c��;�i�V��Cn�ӓ��'��(7C�0:�jٸe�6\!Y
�'�.9�F�,Np���&���P�'�h$�a$CFl�l�7J]�u��(��'���	���$>�B$��,>����	�'������`���N_�NXy�	�'w쐰S�BBԀ��o�.����O�왕��`�$_'uFn���"O��qR́1=.�84dY�\��z�"O��K%5Dv<�EH���� R"O �B���?<ÄHH���v3�=�4"O����$ޮ
�	���Iq24�#�"O�T���S;?��E[ŀM/w0�l�d"O��h�� ������4J�J�"O����<F��ER���]f��"O��u)�%!vq)��F����!"OJ 4HܕC��@(4/H/I�@%��"O8h�6�׉0�(�0�N��y���� "O���΄�N�{f$��B�XX�b"Oި` �u3<pCp�F
�0�a#"O.X�U��(͈�`?
h2���>A
�CPbE��f���e�F��A�r݆ȓ07r�A�)�]���Y�*�	�"\�ȓ'�����	p�)�MJW�V|�ȓ=��uaU��t�#��9��1��;k��GE��H�\���x^Ty��b��Rf��(��u�k`~���7@�,Sd[7������?t��(��P;!a �ǚU�.yDÔ�BF�� ������)���ĉ�t��WRv@gŃ��d{BeQ�'�-�ȓb�KE@���֪q_���y�@�NΈ�!���S�`h���Í�y��ʠ<�
�p�J�A�4����y�F�:/�^\h�ئ©@K/�y��Z�{����@j�|l���yb' N�E��{Ҕ����:�PyR�	&S���R�dn�pƧ\A�<I����!0��?g���XƊt�<�P�L01E��xR��V�����Hr�<i���+��r�KQ�{Zn�"�h�m�<� Zu��� m|�5�ԃ$3��\(�"O��G�� ��]���4^��=��"OM��*K<
x��aU�S�Tq�s"O��C�.(�V�Q�+�����"O���E�z��x!`Ȉ1�t��"OH`
��us��3��tm�� 5"Oqj%Jڛt�l�)�*R�{:�䣧"O�]yw'�":!�\d��/.Yb}�"O�2�->dz�i�4b�l�"OHY7 }�Rm`i�"�����"O�0RG\�Y Z͐�CBJ�m��"O��؅V�yr �r�8;+ᚒ"O<��`]M��` ݫ%^� "O��s6AS ���r��	:�1"O1�E(ѐ�2��$d4��s�"O*��3(ڒ^�B�x��q��_��y¥���L����i|�P�͉�y2
 f�%� ��X�$s�� �yD��(�
pxą
:�X��Y��yR	��*��p
�c[�	�<���yR�)8��1T���+�0%Z�,E�y�(S.ϤdP�'O<veH����]�yb���B ��8�ɀ+qh�� ����yR&U�a�p,˷�͸Ln\/�y�.֎K��b�h1Nؠ#tmԳ�y�."�u��'T�!E�a��5�y�B �QE0��Ą1!��@�;�yBkL<"Җy��F�rT��G���y��Z']���2)����#���y���)���󀀿�D�(�n֝�y�E�J��i�������Y�y� б��(�uC�$�Duy��	��yr���D-a��єLz�ݲ�#(�y�JɎH^,\X!��<��<+����y�EN�3��/Q�-:������4�y��1����dF�3$�}1�<�y�(�]�0�j͡`Z�H35�I �y��)K��U��,Yb�b���y���b�˴��O"�ġ���1�y�	�3C����Ą�J�%�R�Ȱ�y�+�A�<�����::��)ǀ�
�y��̝i�̜�&U�H�����\��y���B��QR���o�؉X E���ybŉ'�
���� 'dĺP����yr��6¼�뇁עW�V(H�a��y"C7By���q��6Y��uK��Ņ�y�S�7�V`Y��A�LISw@I?�y���@1��ȁ�69�	P�HT2�y����Ґ{�eL�vE�?�y"K�_��Y�CK���rqp ����y��S;�~�Pte��w���2�-�
�y��YO���k��R�D� ��&O��yr��{߈  �nR2;?��)����y�Vj��Y�k�3����mĤ�yr`]�a�4��< t 2��y��E�$$�w`�&���I�yҥ	.\�����z�tT���yi�@�S!L��'uܝ��F��yREس�p:JV����I���y2B�m����'�4���$���yr��0/ �{O�j-�8#��9�y" �!n�Q�I�*hT��!��R�y��|����,�M��DjX��y��f
�۳�O�O|�وt� >�y
� ���3'���i�&Zt�$ v"O�m;E`�0g���P�=:��("�"O4�*��d�^���ăRS
�E"OD<�.��8��a�Lt0��T�<AЎD(~.Ź�3@ ��
�Q�<qdnթ�!z0H
/W!������V�<qR�;P����l�g�<A4(G6n�|c�Gӓ�j�u��l�<q%hș��-��ܦ��EQ�Qs�<a�K�Eh��Z�&��k"����W�<����Q�a��D
Q�1d��J�<��c7ms:�K$�("�,1B�JE�<1�"J9*q��j�#(&B�H�l�G�<���6D�48�vjRIܒ���#NF�<a�N��Lsd�H���:h`pQ+��<iE�b���a�lN��K�b�f�<��n��D~Z�(��ŵR�"��A�a�<��-q7&a�DW�d����g�w�<���U�j��B�6�4��F�h�<aT,�W���q�E��5����y�<y��Vn|JE@$iȹj�V����x�<a�-Q?=��k�B�?�,)�d�w�<����(؆���*X<1%N\��l�<I��FTn�XzdJ�8�l�p�@@�<I��Z�JlXI^�b�p�}�<���K/B
�yF�M�,^�u�uÝO�<A�ɛ�LXūQAlJv}�7JXJ�<Y�#j��RPpC��A��G�<ARaD�lQV�!aT�M&�t"�`HE�<�b蓘o\D�+��T��"�&�C�<��[=gˈ�儒35>�f�x�<Y���>*�q�c�':�{�ii�<�tǖ�{(�h;���A���ӭ b�<�6 
 T��@������@m�a�<�4�ɱX����2DԐzf/a�<�.���i���ܞ:d��PG�[�<�᥈>�V�Dg�0���7/�\�<Ia��=;�����\T	��0�(�|�<��֥^)�R��$�؀��Oy�<y#�^*z���d��D88PT��u�<Yuf�8 "l i����$0x��G�<9���n��A�J�8`���^�<�r���=<6�@�B�6d�	�mFW�<Y��-7����˻`�ʉ��]O�<!�� 0Q�U��M�8;f��b��L�<)&$�=�z�ۇ�*u2^4c`#LF�<i�B�q����-K��D äh�D�<i����7g�x�%,׉_����G@�<���۶/Ct��B́�ZQ�Q�7�GW�<	�L*k��m�F/�e��)P�T�<��ӎ�v�aq���Ƭq �v�<!��N�=�����79Φl�.J�<Y�)1����[�y��!QWH�<Q�LG�pM�q�(D�N�_�<��C��J�L�9cNˢ)<����r�<RMF�w������Z�Z��W��r�<�pkE����Lː�BDڥ�Z�<Y6� �<_�����=J�u ��YT�<A�,�� ��P��@Z!"�����eR{�<�!!�`�D��S!�r�<l�d��y�<�ҍ�_r�6��z�ިAF�a�<��l�u�ș�-ōM�E��O�h�<��쐾o=�4� H���S	�M�<�d�6*��H1셅�,�̈́`�<� 0L���ЗZ5��C@C8$�h��"Ou��D��T� ����4��Æ�^�<၌�J�nq`UG�>����_�<A���Ŵ�b �Đ<�*(e�W�<���	z�Yr�-�5h1��h�V�<q再/0P5�G�	X�4q�3��g�<���AϤ����Y��т�f�c�<�q-@�J9{Po��7�����k�<�4/�<CJ�A�a[�n�X���&�g�<����w�nI�CO�IL�*W,	L�<�$KB,H@�D�]4'U��Ba�<Ƀ��97jʰ`%ШTl�B,_H�<�����d��x��$��1��Yy�<)wh)0z�4����	B!ڴ	�)�o�<!r�[c�mR�K�;�ai�"�S�<�2(S%L�KӮ2��w��V�<V�ͫq �)@�N�d�����CH�<ye$Rx�Uk��
8 Z�Hd*Y�<A
oa�/��q����T�A�$q���{ȴ�I�$ˎ���KV�X�n�.M��iֵ𐄐�GJ��7��5U���ȓS;M���I�lTL;��� �:���-�T�PR!;n?����l,K<�,�ȓ\��=IR�^$sF��Wj��LVL�� ��(R戠��q"Š5�q��J\�ej2-�:d��OɁ	�ԇȓjr�(r�%�=�Z򇋇{�H�ȓD��l	�B�0>�ة��L���NL����u�Ѕ�G�, <�������q�R'4� 1	ƫU+0t�-��"�8 ��)9 �u�!��Eb�'>�@��F�S�H��Q@I^|���
�'���Jʝ~�
 a��?hFp`�'P�E�1%�7.F�[�œ9�E�'D6��ec�?\
����K�)�����'!.!j��]'M��Mۧ5
Vp�
�'�(��ѫ� 3�> a4��=6``a
�'��;���}(���ˌDy�ٸ	�'fn�	�&�y"8�JQ+�>�ʘ�	�'3��"��4d\H����ȓP%�-JBER�E���rGE@����]�R�b�"K"�\س�ļM�,܆ȓ"q���Ð(8�u�V��!1�e�ȓ{��u�����T����H氅�}�����żrt��B7>������d�Έ�j�i��]'Fn�ȓd����KN�����iZ�]sH��+��B�,b�@���8���ȓL�@��#!�b0���7h<���\y���A4�����2g@HI��#]��#ϗ.�8��A�(bx���}�����!�9;�%��F��m�H	�ȓ/�ZlRT�ѲZz���C�?���ȓSV`�q�%B�aԈ��EJN�%j��Fh��O���'�P,<��]�ȓ�ؔK��4�D�ӕ�̦|Z�Ԅ��j)�a���	��i�"���h|M���Ԓ!W~A�1��Z�@`�ȓ�(�Yb����T��ȷ_�t`�����cG*G])�C޻E�@8�ȓR(pP]y��(cQT�2ئ$��"O �Ic�I�e�Mh�!�!M�ʹ�f"Oذ�6W�����֋3{�d��\�<A�KJ�3�hi@(�]���J���B�<� n�#e�J#:�^ �i�w��5q�"O��I�`.���w����䐓"O1�m\�cޢ�1'_1d��dQ%"O�Lk�'�59:45jwK@m�"O2����r$���f�� f�h`�"O�9)rN�c�(�:p� {ʥ��"O�a�!�4��šp%�"+`���"Ob��C��Xa���s�7�b���'�(��!�5�Xa`0%T+�J���'��e���#�x�K�Qh���'��+�`�i��2ք��'�|��ubZvA�tX��A!��\��'�`["��xt��D	�ܚ��'f,�ch�7@m�V�(�bT��+��= ��G'H�mA4�	�ȓz�����-ѷ9\2���&����|��@a��>-Tj��w(���i���CX1�Z@��o��@���ȓB="M�s�'&$��`&$�%����ȓI{�@���$�]PC��ä���%��"lڽ1���Ɔ�P^Շȓ,�1!g"̺[�&h� �"O��ȓ>R��W��$r�BA���%#�4H��!�8Ê:v�@��Ս^Ϯ�ȓ2É�Z^��Wg5��a��v,�!!�u��v&�>:��ȓ@����P�ȕ:�~�2��G:p#̵��*�Z`{���W�$��+�4z�"��r���Ru`Fk[xDBh9=�Їȓ3�R4�FBǺ�E��gӴc��̇� 1������7R�5lU%F0���l��̰��@$�"��$`�����oQ�q�d����!uE������D�d����l�j��3 �3e�LՅȓ�2P�u`�	t�|9�)̭iKȘ�ȓ �<�d�^������,(>���e�s�+�1S�Xq�C�)�Ć�QX�Qr�7S��0�B��B����ȓfR �f�W-3ޘ 1�T�=��ԄȓpŊ�0���Z� ��<l��̄ȓh��<XB�5�]2�H�Y9��ȓ,r*i�ghly��] 1�,d���� X�>pH���ǿT������{�,$"!ZR��;/�r=�ȓ��0�K�^�NL3�(ǾM�p��ȓ+_�����i�t��a\?|�m�����B��P�pd:� ��v��نȓ"_�u#��Q�F��\�;�R��	v�������.���� �L]d4�-�;D�}��<D�p�H�eR]B��K';	8�q��/D�P����'ZR�����\7I0����+D�4R���xpnEX�+V�m�9��)$D�D�򢔀4t�
�\� Ai4-/D�lc��LE.��fO^�3�����,D�`�V$'pd+��9,E��Q�?D��D,P�
�ɫ6B*
t� C#c?D���獢1�mф�@,^����<D� �4C�/6��� C߽#�:���9D����LØ2��g&_FP��+D�d�0%��O"�Q�°$�N��D*D����U+&�@�+�ø+D�z�h2D��@!#E	\��9h����D��i�O@�=E���&&K�0�B)��\4�e�R�,n!���[��z#� �y�Æ!;P!�� ��Y�~�<uǚ4pY^��"OtX�V��
7ܞ�a�����"OE(҆�-��Q���ļF}JT�e"O��#�R�3�n�"6|��
�"O�H8�����Xx�MHSqfi[��d�O���Oj�;w��J���HE
^�*��)��'�f���o��'R�;Uo��z���'���vNȝM�f`�A�ϝw>l�B�'��ҍ�~@����}'���'��ybEAV�0���*�v�r��'l�lR���<E<��۠=F�8�'�l1���I���H�� ȄʓB���`u��u�fZ2)�A��ȓ� )�S_ N?2(��н]�bH�ȓ.��-��
Y�*�hѓ"U�I��`��w)��
'.ƕDڬ	�#��}�X\��e��c��ͣ~�$|pփ�)C�����!��!�Q�ld8�b�*H��'����ԔȠ�ϔr< ��"�4؉�EK�"�I��T�Q�Xi��:��o��8�ұ$%�@���v��%�@�L�~�J�z�W5�F���G�Z8�ǩ��_r�
҅	'o�9�ȓy�ع��,q��)�ACT�Н��FN^��$����Kw'�G�ńȓzLnMI���-+���E�T�9�*��ȓ+/ u+A�L�_�̱�MƎ%,B��(�����#ƫLR�1�JF
6�0y�ȓh�ɒCU�3��pѠcɜt|d�ȓ-���!��T�P:|�6��(��`�ȓ����݊a�RZ�KYT�d��ȓ5�d*D�H^d��ɲ�#F�rp��/��Mң���X,yA�X�F�h��!���Gɋ&r@��x!"\08a*Y��af������<Ft�H�c�*nN��ȓR���E�4%Cf ���>K�4���3&hy���	�c���ӀO�;gH���ȓo�X�9S�БOs���զ�7s�4�ȓ�*PbG���OCL ��O�/O�>��[8���5�b ���.t�61�ȓ?N8=�P�S4(�ڔ)���&)� ��-�09�`/R�Zd��OH�Rt�Ȅȓ3�P�Q�`��n[�$r4GҊw��l��V͖�9���%(�pm�.R@���ȓ�(���۳_fB�i�CX�ZR���i�����טPÎU��<�Ե��/֩�Vb��6e԰i2jF�%���,��+0'�'wV&��t��P �8�� >%9��ɿ/�0��M��5�ȓT8��r��';��p���cq�]���r\�`�_1I@H��I܁p��ȓCӰ��rLI;F*�s�&A?yVv=�ȓ�⭃�K%P�Fh3H��(�ȓC�|��$��!h�-��dQoR�!�?9���0|
֠R	3����G.!�H!���d�<����K� x�4Ę�r�DXaHa�<��	1o�4	1�b��*�[�<I�쎀e8�m�T"D�F^bh�L�<1A@�1)����#u���(7�P�<y�*�^������S�
�8��[W�<i����>�|��X�u������m�<��%\�J!�Th�"��� ����g�<��ģ,�, ��l�	2@ +w�]e�<�Ύ�kT�(F�ֶW����BCEd�<� ���ĕ!%@�h��J�q"O pAPf�o�J��P�!s��0��"O�ݻQ	�e����m�x�c"O2P�[6~-6��cϜ-O�� x��$�O���IB�+�
� ƕ�v� �X�aȋqў���I�+(6Qi�E	�:ؙ�l­w]B�IX�D�KEN̋} ��P�E�1"2C�	�K\1�rO��hXN���l�<47C�ɪEEr8�ǃҋq�,* �R�B�ɷ^k���$K*d���J_����$h�P��f�.1 4��$D�)�t��'&)D�(�f=R�|��%��g�(�4n(D���t�:WF,�aw.^�
$�(�E!"D���r�TyG��`�%юyK~@h�B>D��	h����Q5R��K D��2�J/��aJ�P.t�t��g�0D��!�I7s��PǪ1Kz��/.4�x��Z3(�$��9	�����ψ|y��'��83�.i��a�FĔD�FHH>I�
tC�O�z�V�ZP�òY��X�ȓjɖ��p�O�D�4-Rd̗�~ނD���"�z���vp!:A�"Fв$��AIEK��kr�ꏢG�Ω�ȓO�f����?����MJ�!-�=�ȓB���)Q�+B�Eт�	�hh��7<�h��C�>���!$��bٕ'�a~b J(�4�^�����%�K��yb�E�'����,�X��� �!Ƅ�y��FD\q�߃}z�A�'�5�y��Υ���G�6f�\]b#�'�y2�~n��;)U2�� R��5��x�V?z�� �#Z$�("F�V w!򤚧zh`a[�j�-%V�E��MS!�$O"S���e�*h��%`TJZ?!򄞂<6{���8}N��FI>X%!�E�m��L+�  �(�V����A�!�d�-!`T��V�=/ڬ�1��
�!�dD�l2�����X-�\J��n�!�Ę<Z��}����;��S@����!�H�xX��)'�_^*�k�B]>�'a|�!�2�	�B���ta���C�y��firAk�,Y4��`V�3A�����2U���ȈDp��#��2<(�%�ȓV �@e|o2e�b�+NZ����}K����:b0�;���*"݆�Bs��2�2�b���lI?��5E{2�'}Hq���"ŜQB�&ɶ&錐i
�'�r�Y��u9�	Bo�H@��	�'h@�5��7\��A2��F_��I�'�6������^)80�7C�<KHb)a�'�L�G�Cz���V�š7���P�'$b��ˋ*k�"!3����0�ȓ�(���̔�_���Pk@�6!�M���g~"�E0��]����8G2\������y�#��^dɁ�P�A��qS�;�y2���J5(i�H�#���y��č�y2ⓞ)V��3��Уl}̵{D���y���g�\��]�9�S�^�y2�L90���YS��]�b�s�I�!�y� P�f��$IfU�0�7�y��2n$f��*	�����ꘕ�y��N�4U^����*����V�y�e
)W��!*2+$�L
w��5�y2�K$Fh��R�#'�𐖠��y
� <�i�f	�����S��}�"O�ʅ�^\Y ��BjR��ܸ��"Of�1GO��V3*�0G��-t+����"O����l١�(H��Z��"O<āGA�$Қd��C�h��"O�=0�G�x��A�U�Ț��Q�"O�l9��'E��P��n�L��졤"O6�I��);�O�	ƌ��"Oz�ە@O薌I mηP���E"O&H	�
<u� =�a��$4�؁y�"OL��u��>�n
����HC�'��Q��Y�lA&C#�T�C�'����	�+�<h� �ن�p�J�'8�"V��',|���k��?�Y��'�p�iVn��3#�U��c�;}@�r�'�$���ʠDSB,3��i{	�'jN�̏-;9��0�mK((qx$q(O��OZ�}��0�����,h�V	�0�
� �vm��~R>�C�֘[�n��%�E�5��i�ȓ��WH 5���x��4 7 L�ȓb�p�kaF�W~�`A�%6�ؠ�ȓ^�zYi�P�.��$��F9W߈X�ȓ�r�t��Q}¬�U���ȓ@�D��'�S&4�TMIV�ͅy�����|����z��# �|�@IAL�
�<�3�8D�0C�;>�:���� 3LLu"��!D��R��%CW�y�aO�"g��)�&%D���F 9ig����М�,u"��?D�\���ڷF��PY�G�%n�b99+?D�dK��!`�S�MO�3�P�<��Vy��58fFE�2�ҒUݲ���(	�˓���h��d����%�ʎvevP���K3�!�&!�T�� ���Qba괧�&�!���K�>�[�ށ�l�b��R�!򄖉}vޠU�3>�p 
�e�2k�!��R����d-N�5δ��E_:Kp!�$�q'.��E��� �T<c%�H~4�O����|
�O7�H�gl����Okux1�	�'*H|� Ɛ�j(�%�>s��A"
�'8�q�������T���d����	�'qt��e�\�N��Q���Z	�'�������z�3�o P���'�
D+���Xn�a�PH�y��er�'14��G�^;\N��w�FgD��[��'����|:P���<AހI��>'#�0�t�YV�<���4f��kd˼Q��¡)�{�<����96pMb'�ܶ�J��db�a�<��c�gb��(1-b���֍a�<���
�%� �It�S�|{�$Z���E�<���I�Lø�1��V!:�)��\�<a��^+Y��W�&XZ�Ы���X����$2�
S4�'	�*IwA�A)�v����L�H9���ߍ~Tb��v�4I����족�˙',�e��/Hz�u�ȓiU*y����P�b��,��v;Q$/r�A+�.5Qsv��v�`-�2L��1xz��f��<{j	�ȓPa�� @�	<؂�
f/5Hp6��wwr��-� �N�ʑ�J Dx��	{~r/��FF��.֬z�b,�Eg���y��� *)R�["Z�m�}�u��yb�޻#�L5���ߢ<�"���Ԅ�y�h�)��X9 �K	0�@ѣ�T��y�@�L���K+��<��^��y
� T���D]D=�� �r��D"O�r���:R
�q�N�O�8EQ'�P���pO״�8��ݫZVP(U�"D���#@�=5"��P�`	t�*��Ӌ%D���3�I�yn���#�9v�u�1D��x��ޑO� |�F�\�Wn$��e�;D�Xx���'_[�y�CN�q��AIt�.D�,y��L+XB=#�M־�� pv�,D�p�ć&-������T��`�!+D�|�W�S�(��,�rL�+�\\AF*6D��`�D.\��4��H��I���a�9D�\I@e	�B��z5��n��D`F�7D�<R�n]4䜌���D �Ԍ��+D��R����d2Pܨ���#�b��7 &D�䨆�E_E���~R��ĥ$D�XQ�
Y�V�l���I����O�OC��<^�:PR4k�*�@�
\abLʓ�?��_�l�i��J�6�bF�J6s�����;-Dp �kL<6H@�鰦P3v[��ȓ`�|%�E/\���m-X��9�ȓ~��ɢ��Fa�LA ��"\�Ru��%5�łBJ�V<�F(	H�.5�Ɠ|6L��*��n$BD��z9�X�-O���΄k̥��&,�)��r���d��@��g�P��m�4�PCY��j>D��0j��m��p�Z�~�t��i<D��ئM�q�H��$��`)ҥ��.D�� Eǫb�\�.�!�E��c&D�)3Ï7�tA9��x���P�P����
|�i�E� ��`Ѝ��/�B��ȓlt��ࡗ0Wit$z���>K����?����hY ��>ju���|�x��ȓD�t� �N����(c���P��Մȓ%�x��$Vy�4¤h[�e~ƀ��ON��s��ܿ4���)ѦC���d��9\*E� b͌Z�,�	�G�*3$���;2Hy���Ѻ>�lX8�m�K��<�ȓb��h�F�!M�`��fL;I$^��ȓ�T8��M�NV�����P�x,Ԑ�ȓ���b��8��t#S�l\|(��nވ�G*��.���#!S�i��V�qr
ز�L�@�&�n��ȓw��!��C�":瘈�g�U	��ȓ&6����� Z���t��+���2A̽����%�p���<s��J0,`#  W.:� ���$ȦspD��tY��"<�&����8t4��)Z�L�����35���k*l�&u��8bPia(߂?1�ET�/���ȓ)�]Y��CQ��bǂ�@�f��ȓ-ty���¶ckZeK�(6X�l��B-�A�R�Ń} ��f�浆�b�����V�zAƠ��(��9����P�c!�( �<�p�®E����!����J��~R�*E��O5��ȓ?��bQ�ԌZ�푫l}�	��=D�d�"יTg���O<n㸑�Ԇ<D�Tz�G���1:��M#<�X� D�� �J�U�݊0e^�{�6���@3D����НK����U^4,�;D��zTĐ�?�y��[M]���p�<D����fG,F�i���x���:D����@_ �4�����<���,D�T���̃ ��R2*S�z�����'D�� \5b�gZ,��H�!��W��X&"O��jq��kײx	Ȍ<�Eb"O��aW�؈��\
'���`E!�"O���`�kE�Ih�+��f�ni�"O0��&H���B8�d��H�@T�%"O�Y*gؗA_N�[��#q�(��"O��b� �1��3��;����"Oʽkw���4R�J� �F&�"O�M�f��bӾ���	=$#f�:�"O"�A�38�С��)��0����"O =�W@!~)�acwȌ0Q��
�"O  �e�.|�LqP�G�n}ހ�"OĜ�p�[�&���K�M��ڜe"O�`Q�i���R޶	up"Ol��7�H>4��D��ܦP��qxV*O,h����n�ؓBX�[����'K�0P�� �% 2J�K�^)0�3
�'�!���:��@�$O�L���A�'�\EH����x@ C���{��a�'�=�7ˇ5�V�*7�ԅ!E��'��h�ӧ�1A�����o��ɒ8�
�'��0��K8��pHV��&Җ��'�fi��8pB��u�N���9��'Uz����+&�����c<�����'��l+���g`�(Ί�}�`�
�'�� 1K�洂�'� z�j��''�<�vn� l���e
V�>��9#�',�Q5鏕KA�c�[�3��l{�'�r�YG��N���k�ȇ0��
�'�M�$c��7]�(��7��i;
�'ؚ�P�ٌ
z���Bҿ�0y��'b.U`���@���N&u�K�'�r��a�Q�n!�E�į@$���"O�� ��Hq��d AP�F��""O�@�ZR`��8��Im�� r"O�p���E�f�z���N9vɠqx6"O��؃E�Dj"u�U�����"O���GcX��u��&؀|�����"O��0���!�Ba�䐫+|x�!�"O�����Py����7�E�x�FY�W"OV����x)�!�!{��[�"O���W���-� ��0����@I0"O�,��*ޭ*�)�Yp���"Or�Av�?�8��l�-�j��"O���/F�e����V',���.�!��	��hc��.h �� �ϑ?2�!���FC��"�Nꄝ�A��~!�D��tE�,ƥ�;u��aVMV0,i!�d!ݴ�ㄨ~�$�� ��vq!�$a�l%�foR$a���c#$�>5!�Ę�@�\�� �S�>��DIO��!�$B�pU0���g�rYR�']4B�!��-
�x���k���AL�4�!�$2X7����ÓXʰ]��do�!�DF�tT�"��\R��p䋋!�$Q's3�!�hY�RV"�#��Ppg!�C� _�yjflN��񁓠S�-Z!�$~�"H6K�8I'V�!v���A!���0t�z��-�>'�U�r�Z�9'!��DQ��e�G!2�~$8���!�ė�5;A�#�a����!t�!�d^��R��J�NҀ�U��'�!�7k�
1���N�Y�amG�r�!�	��&�9�L�m+������!�� ����APT�,b"D�ar��S"O\�
w��=+ؼ�@@Ǥ8�Y��"O
T�d*�3L��9Ơ�[o�	�'"OP]�q�Yw�l�UF�u˄b�"O&��3 �<�ly+�D�_��P%"O�)��,� C����PW�Yl*ȑF"Ob���")4G��;��zb�"Ol��r	[^u�À]|�: a�"O�ڠ� �{v���Z�{���"O�p�q���������C�"OL��Z3�RܪԢS�Hֈh�"O"����2����'�b*P�� "O�*Q�.w�DY��f�.I�=�"O�{�䁚0A�2�f4<кm "O��be\�4��kA��:�N��$"O�E�C\Khp��@��z�n�g"OI�'�\"��q�" �p�r��"O�<"����5H���-���H%"OPdud��
$�Qɀ�˵>�j4I�"O �3�HЬO1t�a��1m`NT��"O8`ꡈZ,0G
(e�$S.�(�"O�𑬁J�t!oD�"CP��A"O�qREʴc/0�nV���.!�dг<U�eB���F�b�͌�Ar!��4�L��É&�R�X2J	�4t!�dP������#�l�&�"?n!��Û:�:� Њ��z���ɶG�!�ʶ#������9�Nݪ��W�J�!�d+�J, �dG�?�����9�!�dڍ]������#5�I�|ќC�I"�����ŉg�Z�A�41ΞC�ɽ"H���i�-PFDxD,��yP�C�<T���c!�̀<�D Z��̨u8JB�I;x?�Y�K�;m���g�~} B�I%d�x��_9Y�������,B�ɯ�ua��	y��qXE䋳R��C�	U��M���LI]�1�E�՚5�C䉪wU�x�&�M�	%�� �m�(#M�B�	8�t�5(F��X-]P�B�L��K��	.Ek�y
���9d��B�F4�	F�42|��1�jB��,th���z����^�KDB�I\��T�h {��ȆB�I�lݪ�+�-�(b�.�B�C�>��C�	+-�ʩ�Ն�d��8�PkT|��C�ɚ4!����P������L�<B�#E�Q�%]�NR�q"a�1o�B�	�^�HC3������Y�W�p�
�'"���[b��h�こ�L�RU�
�'�6b�![�?��`c�o�(}`
�'�ؐ�tgY�`R��˂�:gI��'��R$�=,���Ɨ4:����'�H���Δ_����"Õ%g}1
�'.l�3BƆ�.�v���l�P�*P3	�'b%�aR�y��i@>'�1��'y���sD4)aLa��QQ0pZ
�'U��R��6c������)�'����4�_�.F�asA��-@{�y�'�����RA]�0��j�6�P�J�'<����X?m���uHU�𲈘�'s<��_�$�z�c�
(��'6j�X���	��d��|�~��'��I�C$[�j I4�;?��k	�'��mȤK]?D|8�� &������� $�F�&� ����p7���c"Ox���|C�\�#�Z p��e"O���1NO�,L��Џ!���"O6D"�ƿw"�A�t`��-�!�s"O�ڰ��IPB�ޤR�`hw���yB�<����i�}��|��K�y zIr��D�ܼy�A+�䓶�y2��bY�!������F,�y�'�<.R��ˑa�,
�R%*����y����d��P��4�����G܁�y"j,1���6��*2�2����ԅ�yR(@6�^��d΋�3:�ٻ��O2�y�H�sP($jsl�#�2���e�yr��/{ )����!v�8�a&X��y�K��N�LMP�΂��	8dJ��y���0:�u�P�E,	o@�ϙ�y���6��2��(w]`Px�R�yR�&����Իpx	��!�y����1�Jv����1���y���y�v�9P/	��\<2�*�3�y�c��x�0�D�ا'��p������y  n��p�SZ#:�$��	R��y�D�&<��qɇ`
�P�V��)�y2.5�ś�G���h�㛵�y���,&"X���ҹK�-ڤ��yb+M�e�j��emw�ޥT�� �y2��rȤq" D4m��v�R6�yƃ�?��8���7���p$�y@�sV ɷ�"6���qť��y��]�v� �!����3���;�F�2�y����m� O����ˤ���yr��i����)
#*�&�Db_6�y�
J53�̸�b�&4����ȅ�y�Mߖ2�L���Z'O��9��]>�y"fX!¡��Τ��Ȣ��yrK��IZIzw�:��l�bJ��yn�@�I`��{�l	�c��y"kC�	a����\VU�vJR��yb�%AY���3N�조ࠋ��y)$���I�<�������yb�D )Լ���������#�yb�u�ƅ�'pq��E�y®�6�tzt�+��� ���y�$A��Y��I�|t�u��bX#�y�d�2 �R�FP�pN��xv%�1�yb�V�o�h�&�e��� K�y¨J��ġ�N?aI�]pS��yR�;A45�J�.��H��E��yB#�u�xpG��[` {�n�"�y�3a�:AY�C��y&�)�	�y��ߖ5����&a�����SsϚ�Py�
�T�#���J?@Z�ώV�<A�Cӊ_Ȩ���<�l�f S�<Aw*�'��C�B
_�i�T�GZ�<��	+,���xRe�2[�j帆��n�<1�Dk�V���o�+���`&Âi�<����*������'t%�� ���N�<�P�^z 4j�l��>?"ٳ�L�L�<y$��H33�Ě
K��1G�@�<�s�ɻBa�3հ!G���%�Js�<1C` 3>&@Bb�ߑg�ج��Gt�<9dKI2)�B	���P������m�<��ǌ=ҡ���D���ف�h�<aD$���B��Q;y�L9�&Qe�<� L�3��֢R���%Η�
IDE؅"O�m8p�N�<8��l��@��Q�"O��2U"Ѥ	|�ja&�T�~��c"O�򓇙�Im|b��w� "O��V��˄�0t*_2|�*��"O9��m��ZEkħF��"O�8�6�ƷJc$���L�D�N�	�"O���E�^jr��&�L��,+!"O��sՎ�q�܄(c �[�N�0�"OZQ��iT�����l�
�zW"O�-Y��9
�&IU��'Q��8�u"O� �Ů�d�[���2ܼ*�"OR��d+ݐ-R�ݲ�o��e�r%��"O��	e�׆\�Pq�`E�-�j�:D"O����e��d�t�p��Ђd2P=�2"O�ZW�P[�j�H�)S�Z.1H#"O���2혇�XE9Ї������"O ����F.���>T�N�yt"Or 9BOS�7�H �D�gODm��"OB4!�F�ґ��B8`>ʹ�s"O�X1�Ŏ�$� �JD��|�`B"O�1�U����f	�:R�`�G"O$�[pkȕFLFHq� 9��5"O���e-�M�,�zfCH�K�8�"O�]a��D/j���DN�+�dՉp"O.���
c��#�⚣2|nثS"Oh��pG,<���7Bd؆7�&D���G�V
��Z�LX���ŉ&D�h�ǧ�P��rT��G�\5�N#D�pQ¢�J�� � ���i�$"D��)�$�2,��9A��M\Ҵj!D��uj�*��؃�ɑ�jH�V�)D��&��>64�HD�.;ht	f�,D��ą6Kn킓�ěl��H7�)D���L��Ҡ��3-X^���!D�@ e߇��Baf�
I���0( D��Q��A�<�+�j�9�q��+D���.R�}ɲ�Q�
H��|�6"$D����9��׀�8W����*"D��ba��+�M���8D�|b'�-D�ԑGc�H�h�X4�7V�q��-D���sR9v��ԁ�`Q*kV�ԈS`*D��P���	X�5�'P4
z��J0&+D���#!Wy؞H�!�_j���'D�8	Aa� E����HL� �P��&�&D���gBf=�P+�.��%������0D�@�w/�>O�a��D#tb�9���0D����P6�T��g�]*j'�d�G�-D�@���\�*��K�k,X�!�i-D�Tf���|��e�4]�py�%D��n��m놵�P̙�GN�b&A#D��@���:UM���T$�2R�� D� X�c#iB��Yf#O;�
���I>D�\�#fS�/�b��F�8򶀙�'>D��H�@ע;�H�qFE�j��ؒJ?D��@V��]A��[1���r��(8�d>D��(���N4��(����,���׮?D���&b��Ea0,�㥚 +��q`�=D�عdMۛV6�� T�>r���EN=D�@[*ǜg� �I�K�fR*m��.:D��B0�V3��h�$�MO�`�,8D�� �#�6
P8x�j��|���0�6D��h7c��5�F�H���L�F���B4D�|3S,�"|`� �D����$7D�� �l s�3�)����za|�XP"O�� �AJ.#>��cd\C��0�"OZ�&�Љ�IZ1��.s9�=�e"O4�8a'V�v�Z��ŭѠ`%
I�0"O^$�%�Q5n��騶��:F,6M�p"O�Y����.5e�5�������"O�m�f���
��j4bf"O�0��H��d��$��l��T#�"O|�z�B��W<a
�dߔNE2�"O� ��'�#?�0�I��=���{�"Of��"S&㎙ѓGA���[4"O�p���F�lL0�Z$�T�gB��SD*O�1�J�6B��h�\��TmC	�'����o>en���M���M�	�'�՚���P/D�ITc�
�����'��LA㤉 �v]Q����xI�	�'v����H`�c�E49��S	�'r�p�b�A
pyF��� �H�!	�'��@%I��q�E��	ML��'\�	����1��t���3l��'��aP�ڹu�u�4�ъ}%��:�'t�-p�ɔ�<�|�n�M�r���'J�8���iz�$���\9���'��tXF�=�А�6k��5;�<�	�'��D qH� D�pt�f$My^� 	�'D��A��-@�}a�c�.E��,��'�|�(��OHL8TK*�\�B�'���8/Aqzļ!�g�-/j��	�'�l�����-V���4>�`�y	�'�H;��:4�H*�P�:hq�'c.@P���]¨������`�,t�
�'t��*��F>?�!gnQ��j�
�'�F��&
�)ف�@]Y�@h
�'֘񐎓7jԠ�-I�]O�]��'/p��`���krmTaj�A�'�H܁ө 6pA��a�I�2���'tx��S
7Z�Y�pk!� i�'ڤbv#ݨSܨ�B�����lQ�'\xQ륉��/�$1�RDΕ|40���'`���2�O�+x�IKrdO�c7�%��'Gt�J�'mrf q��V��<�']\��#���9�a㐿�\���'�h)k��X2,��0ao�v��A��'�P��D�U���KA j��=a�'�:l�T���Y��03�Փi�Qs�'D�9�r�ݘdB�P�NZ�/��(I�'�,PA ��!^�Z�Q�L#.�l��'=�H�,S Q"n�HRA%-���
�'���¤ �;�H��dȮ(��@�
�'�-���L�h�x���A%$0L��'�D��&��'�%�O/�x{�'�D��ĕ�9s��[�iH��RU�
�'}� (��G��aJ����9
�'_PX���U_:Mr�ɔ��i	�'���N�$�q��	*G� �'ւꕏ�=jA|�b��F�#�X�'�(p�Ë�'�XcP˅�+��I�'�N��C#N�.��;n�'��9c
�'*V-�D �vY�A�Ҫ-Y�5�	�'�F\35�� ڢs� ���%��'h���4,%�(�H33�`��'~6lke��+$��pt��W��Q�
�'f%� K2aG�ir��D��
�'�1�L�E�D�) [�Er	��� $D9R���^����cd��H�K�"Ob����V�b|�P��l�^L+�"Op�q�*t�~�p��[�X�����"O ���d�(< ��@�Ə7��"O*@ b��f
�5k�e�:"�C�"Oм	�E�h�X�d��r���@"Os���"[֡j�?Pь0�U"O\�����$ie�F�W3H�F���"Oޜ���=���Xя�2u��`�"O�hQ�B��m���`�K�v�pu"O4&l��y��T9�8~c���"OF�Я�%���K�lL�]_�"O�]�&K7Y�%���&Qhj��A"O����p肶�J^��5"�"O�XZ5lW:sT�ö���	���r�"O�@ NB����C��4�=z"O���ȇ%S8��j3&�75|�(�"O�!F���#s�	��'�3��V"OKB/l����Ť��A�N|���C	�y"�K#�Z,H���=Z�t;vLS
�y"�E��vȩw��0�,��#�y��4;#���!&è�j!ZBOC��y2'M�|��D�A��pp�NP��y��N'̙��W�4����,F.�y҂גt2�K-t��o,�y�$O.��I��GW u-��ꂨ���y�+Ғ2�p��R�یv�J$XŠD��yRHqQfE�RAP��9�CNH��y2�߉T���CK��J��FS��y��P�u�� ƌS>��QT	�7�y"�+D�@�JV�H�j�@�B̈́�yr �@9�F�O�dX�y�	ͽ�y��QA�4���Y�[�\m�wO��y�d"��K&��/T��12����yb�N.l��ty���9�@�i� ��y��>Z�y�N#Y$=��Z��y�Gpa�J�A	�Q3���0�����'��dEGP�(�s�ٶ%�ȉ�'R�܋��.G�&e�EVlk��K	�'1�d[6h�zb@X�A�*f��<��'������(2us'M�9[lʄ�
�'%�<���4aꈙá��`���	�'X�H�!��1_	&XB�j�_c2�R	�'�z\�-��։ipN&Q2�uI�'i���$�n����<J��<�'@밉P�}�d��sĒ B�v ��'f�Ʌ�K%	k�!S`E5f�Qb�'��E"�A���6���](bEZ4X�'�� �)
5d&��{�LP=h+ ��
�' ���&�[�ΘkQ�20\q��'�*@�ۡ;��uh�C?�����'��(㠜��|�"�δ]a X��'�\�qj�< �"lY�ט��'�z5�A�0��*�W�x��
�'$��!��A�/��d���.�x���'F���qd�$W�,�֏N}kt��
�'�X���e\�1T����'�����'�
lva�Gv�@�@3�:�	�'�,d��*[6���!0x�n1�ʓRH���uØ1���$b9?�Ĉ��H	�u�%�:n딴ZfB۹S�Bx�ȓj6���b,N�|�£oV�T����DVN�x�bH@C���n��H��D�ȓn�Tz��D�m� !��=����S�? @ pBa��IB �ajM���52�"Oj�J��!�R���h�5̢M�"Of�P��q��S��N�@��15"O�$@I c���3���>Ԫ�"Oʙb��O,W�	�*]m���"O���a�"C]�H`wV���qa"O}"v�� 1���sa�E��@��P"O�)s�O�e�:i[�
 !q��"O�w˝$Lo��롄G�un���4"O �Zp�2�`�գ��S1V]���Q@�<��M�2eZ�z���[���U
%]��	O�)�?��b��X����j:�PAc�<!D�L�m���a��LFʌ,a�F�C�<�)^�B^x���WP�\8eC�|�<��bҭ&�n��F"����c�y�<y�+�:�ly��/�\��� &��\�<��@��g���
1?�| �e�Y�<�Eg�>��w�V�Y�`�U�<�����D\����� W�����H�<A- ko�4�G�� m$���	P�<���
v��-�P�K�K)-���f�<�E_(X{D)��8�`8�w��m�<!pN�;�ʗ�#�~�A#`m��X�>�f��>~�(��� 5�����)�D�<i���A�T䛧�H<_\	�'�Z~�'�?u�q ��;\���>](���(D��8#R	n��|��4#�:�>���"�0� Ƅ8P����^#V���ȓs0p���%'�J�#/Ou44D��:�jՈD����d�c/X,��4E{b�'�� ���v����!C?']$+
�'X<@2�j�#�n<At�0 �E��'�F�G٤�p�:��#%z�=R�'�.����G�4�TM[��đr�u�
�'Q��B2G�0lZey���&J���'�
0h��ٓf�����aT\"u�H�,��IC�xT����}q(]e�@L,�C�	9R� b��D�G�1 v�D/CC�I�}<: �aΊ�p4u:��ś0H8c����ɐ(|�4�q�Q11gh���	7�C䉬[��]�aN�6c�Zٙ$G(��C�ɻJD]`w��~8�ڴep�d"Oؙ��F�0��
�J��*iY�<����=��,(x�0�K��7�(t��^�<�Ph_�Q{6؁v �	a� ����V�<�r�\�ju��e"�_����-�x�<��o�N�Ը�b�?u��Y��	t�'�?%���)I��M��o�2H��R��7D�P����=@ 岴	��1���2�A1D�@@�K�TVH�����{B`$D�(XS��`8�������E(�=D����H����qS�L�M��ݰU�-�O,�I,Ph�P����6(%��2�bWv�v#=�'��>IBt�=C���酦�n�`�)�O��'ޞ#!E��-�L�(bPc��J
�'�(���C \�A�
K�0l�*O�"=a��5g5~!q�L>��r��@�0C!�D�-3�����cŊ��1Ԥ7<Lў�P��K�M
"�tQ���W:^�b�"OJ���A�ܨ� Z>:�a
P��z�OY�R�X	p1W�.l�(h�'�6��1�E�$�����kK�a��%�'�@�a@�2��A��gָ�^x��'�@�Z�Bž�8Y���0?����� �I��%[q��*�ʇ�H٨��"O���ːf=����G&8J��"O���1��/�"�+�ɜ�>y6,��"O��c�P�Hy"Ƞ�*��8a:�"O��zҢ��u��5�
�R��!�:O@�=E�dI��WJ*�s�l	�d�0m
@��yb�ԴP-ܝ���NmY�A)���y2kT��D{g�?b����p��5�y��ܧ8���pg�Y���P`Eگ�y�⛈�2�౪؍PR�pp( �yr͐��d;D�.CR渒P`'�yr��1p�T�Ö��2@� m˗FD"�y����Yi<a��%3}C��:�y�'�M�1R�KĐ��L�R�yb$��������x2�wLG�yrnI���J�E��aNQ�&E��y�%�\ҔQQDS�^DI�a�Q��y�7l�U���T�aF���pM���y""��(���3��5H����@4�yrfA W�F�2���X�N܁�@��y��_�	���tFK�ebl�p!!F��y�ELhml0B�nͧF��؛PR�y�B�m.IZ�+��=�D�6(U�y���*�Z���+��4+��%i�4�yR.v�� l�&3@4���F��y�H6X4�i� *��Յ�y5L�b1��0�xk��Ǚ�yRD��~$b"$DC�l|�:��\��y��/	�܍�S,U&]��������y"OǜC�\8������P����yR ���K� �>3H �� �y"���2:6����C�#9��r&^�y�BV� j�E*@�[�6kvF���'5.t*��Y�$�-`F�+\��y��'��͑S���g���'`�L���(�'�H:��(GZ�1;���<�<��'�؈�h�� � 
$�A/EU���'E~�����1��`�*����'e�9Q�Α4z޸�VLO�$ê�'~p���ς
��ӕ�$n��	�'�dkAZ�8`�M)��V.�,�Z�'�L�qa-�t�j�r(S)��<��'���Ѥi_�$��`2�<I���#�'l��{�X
7#�-p���?�l2	�'Nlآbu�h9�Ƙ<���y�'r�}�2�L�æ��,�+,Wn���'{�y@e*�G'���ƥ[0$D���'#JM��,ޘR�,�8�dYs�8C�'�>Uq�0@��F�s�((8Q�m!�'W�ŉ�ڨ�@��Lϓ5z(P	�'�А���:!hF�Y�.��,��'@\ݨ���<t�B'� $�<X�'$�<�5&	�#j� ���s�<Qh�'O����]�x�8���N� �`���'G ��aG߃t�i��V� ˒���'�<�#��A�	}�Z��ي��tq�'H>\�UDN'%�(�v�]5xj����'��بp�J�s��`���\t��p[�'���O^H>,	a�Èw��	�'��#�X+�$)��-�0�X�	�'���ˢ��798`kL�%;�Q(�'���òˋ5E��!Z#�� 2����'h�����5Z�U�+���`��'IvA�cM�9~p �`)ڜ6|L���� �!:��@�7H �4��	h��"OdXB@��N�X`�0��J��݉!"O��J�-$n�¨S�៮h��@�"O�ݘpk�P����E���"O���c@�w���P'�S:f"��"O��8�+JF#���5�/h��z�"O�E���E[t�8B� ۱*��� �"O�0�Y�y��]	dbƧz��D�"Ot���%O�JDH��c,� "O<� ��T�h'Z���f�<U����"O,<x�c�# ��5pƜ�|FPd"O���$ 0�С���'xY��"O�a�eJ0L�`(Qe�ޢB`�V"ODЂ�A�y�F�©���l°"O�q�r	�'�05Cc�F�!��I�W"O��Z����� �h��JN��y"A�'z����U�f��}�����yB�+YbY���ϕe���Y��� �y2j_@�hf��g�Q�î�;�y���}�nK T�S�V���,��yҪ�������F@�P�`�!�y�Sl?������g|������'�yb`J����J����O�\���L� �yb(ˎ@�9�#@�B�b��E���yR(��9?ꈡ'��3;������y�Yd�%� Ђ;a�l��m7�yB˘�A��7KP,7I�T�����y���+9v�����+��0B0��y�&F�tb��	Th�VU(�B�O���y"L���I��o˳L;pࡃ��y�:]�q�CX>y�H�z b��y�kޚ��I7`K�x���h��A��yB��#��p�ړ�-�ge;i���`�M��0?ɵ��w��h���N�5@ihqC�r�<a��	o�t���-=B����j�[�<a�-�	�(Y����6����DKl�<�F��Q�B pT꟠��y�m�<�REW�P�@,�G �!#�N�0G&Md�<1D M.��R�[�o� ���c�<) ��S�U����0`�|�R��Z�<�E� F����\2��U�#�Q�<���){`��G/ݯ-�Z�Hu�<1��)G�8��uj��W��Mbd'�o�<a1C&oh�0�`��nE\�Z�fCe�<�eAB2+m"�����'Z��a�z�<A�n��,AȪ�'B�i;Z�֥U]�< ���/߀��g�E_
#%mLg�<i��	�L�f�A%��m��=��ȚH�<�Vd �1ؐ%Z	L�X"��D�<y�I�J�T!!J\�:�@]�GA�<�՗��\��8R��j��K�<�ը�Nutt�"�8� �q0� ^�<�@J�$�xe+��YoܠYe�c�<��f2s�x� �� �c���1�KZ�<y�eN#n>�C�Hv�\�Q�I]�<�R/Q-D>b���WQ�6|�f'w�<�3��#>���`T+~� ݀a$^s�<!D ۙ(&P�"�\.:��aYD��g�<�K�3Eǐ��dl�Z��Ѐ�j{�<iCP*dM�e	�ɝU"�}BC�j�<�g�Y��\*E��2��"�%T�D���ƲM�fT��`�LZ�YQ�2D�����Q�{Ĉ�Ivx��7�.D�<����eْ�����|�\"�f/D�� �t{���4lxw�(�,� Q"O~2�O�@N8��O3T{�D��"O�aY&cݮς�;���)hQ(�"O
HU`�kî�� -ú,D2H�C"O��BW�@�qR �1���9@�5є"O���B/�6�
�)�yF<��"Op0�5�F3E�R�K�ОB��ɰP"Ov`
S�S���Iʗ'�?ky��"O� rc��"�6,�����f���"O�4+��B�Sy&�"F ��]�����"O�`!�aû*B 9�O;k���2�"O��ńG�*7�{R�N�n�(�B"O�\�F��8!ƍ�A�� (`���"O�$���J`��i$B9J"O eG�<w:d��O��`���"O��R�K���eX��J?��ܒ�"O:Lũ^�M�=�F����"OP�����Xul���ڛ@�x�5"O$511��\�tU�2E�O
 A�"Ob1�!7D�Ȱ"���)#"O��8��X�X<"��D��-�F�W"O�!�3�F]E!���1v��5*2"O�9"!�O)���A`��uҜ��"O8A�-M�k�1���k96�"O�j�1S�x�NG�/p��"O��I��H5���с���)��'��P�G�a�S�O�P̛�O��vo���1dK�`Z~��a"OX�b lA �����cV-2�Ĳ��O���>�ny�	�*�f	�d0%h���㇃&�l�E}�IJT�	=|>d�I(�`YcT	"�~Q�w�N�6`��ЁL "E1!�TD<`!��)"]����dR��� �Ԃ��:�X[҂VA62�4ZR1������Ǜ2AK��G\��́]I!���m�(�"��x����~+�,���ۀQ.��ߴy���? �BO�z����O�@�&94�v��&坴2���"��$�O���EV�_#�� ȏ�F�dp�dF�
dÎ��1'!a��y��FMa� ���vz��'�D�@k� �`�5f��Z�l<��P�E����w`��M�!���z9�QH^4U� !��Y:=�����'�DŐ��\`��C�ɵo����`�-	��S �7H��jk��d`�)��CE�K�u�Af�+K�(�`Y|��<�
�p��K16�@�Ѭ͉ �3�"O�|K�K.r�dm� �҉, �T���50��j�W&�2��2"�%X��4�K�p�jM���S( ��x�A 9?�=�V�M0�^���I�F�ੑ��\	5��m#�B��������>zF��p�](©��J$`��c���uY��	�lj$����:A��!�b�;f7�c���.Y~���Q��)�]��
Z����ˁ��`�QC*�o�(�v	��A�"݋f�֟4����I�D�W��.d�4"�aP�~�d|�0dN{;@�B��A�@��M��E�l�'կe������+��� �n��"E��^Dt	(qDGw�'��@铨��l���,����"����P�v�۟,�|�3���C
`ם�"��Fg�-�T��Z�h��&<s����w`�Eu�l"UEa�����yqO���ɡ�U�T:�ɐ�K�oX�Ѷ(,b�~a�����q���Зf��i�4�z������ɱe����g��*C	4��AD���T�D�QlC�&ds�^���7m�
=�uP$��mΆ��@ҖW�I�Pf΅��(��耩k,a��G Za{�Kp��(�"ѤyXǏL�2���Q�6�t�x�{����FO9\�X�Ѧ��@�A������;`�F�H2���:C��)g��Z��F|2\
C�D�TK� �uC�eO P`���	M��" �sU�<B��ʟ��\w��{�ܔ8�X�y��>q �ݘx0!�F��2�đ���<�W��#l���;��h ��6%� 4
7F�=qeL�C@':VEpf Ԓ��6�L�|��g�+
�
�J��'>F�;[Ԗ�ȅn�5w���խI�D
i�$����:4P�K���<��B��eKB�xe"��$`�`�`�nJ�TB$#��_H<�p�X*J�a;�l�8m�qʒ��b�_�$��S��p�gLU	$��.eͻ|��:Bn�!n^�˦.	�%�l���%N��G��Y�`A�� ONj�n�	^��t��k�.n�h�'�6�� C�b�e�&9���h,H����R&�ȸ��I	Y�L�C䗛R�6er&
�%�μ�ߔ=�61���g�!��U
|m�%�p���DkSD��Ola
�H�)$� Њ2�3� � �%�*X���#�! ��͓�"O���d�D�]���#���35��X��Z?J�B����I9��d9�g?ٗ� G<�z�{��('O�U�<q�]�N�Liq�F�K��	u/���?����AdX���[R�*�p��j"&h�㤝#�� 7�Z�&:a|b@�8(Ҹ!�Q�M��q��+�~���ʇ�	'.b���q�ѧM���Lek��ضC�Y�����H��(O��9�,go����ޑ٘O�j�!⟝j?��q�dI�X,�2	�'9��s�B@>=�Ҩ���n��0z��( ��KM�xӧ���aG�b�F$b���E��q�A	"D� !⊂!����)G�"D��"}2����A�鉉h�� �uh��h&����B�|�C�$����O�<,��AJ0G7�C�I�L:`0�!עd�����2c��C䉔W#����a��@�c�Q�C�ɸF�>)��̴X��\KqA�8]�C�ɞ4�������M��Xx�IP�2��B�I t�<�9#���P9���4%�9u�C�ɦpo�D�V(�&�����I1:�B�I0v9�i�V�?7��4���	�mO�B�	\u�%�%��>Mv����>L�C�	������h10L���ǂc�C�	�p��؈��	�ӃEPۤC�	T,�]�Q&$W��%���Q��C䉱Rm�Qb`�
1���2��+.�C�	�*4c�Y6�����!�>*�B�I��\��݊1��̘'��_޲B�Io+|1�a��b�̬P�c� -ԂB�	%��Ш&OBF{�D:�a�I�PC�	�jP�#V�X��$�ӏXwKtB䉅.����n�#��qP��*�B�I/i�u8!�]Tȸ@�cۮ0V�C�	 v��`s��<"+�]�sFU-w�C�ɴ���S��4�pm�Ӭ	dC�	 ��ʀ�׸G�^�b3.N�OA�C�I9ĆT��#�R����}n�C�	�n�(��Uj5�\Ej��W�g� B䉀<7�zU&W�GO���K�Q["B�	�<!>��#��84�eP�d�4B�I0�dE,�!l�t�i��7��B䉳)S&��D�G ~��0*�>)�B�I?g�:������5Bqx�g_�ٲB�I�#�rhkq/&n��JBn�'m�\C�ɑ�B�a�X8M����ca��"�(C�	i��	82c�K����F�+�C䉜��u�Q�	�b ���䇓��C�	�|OZ[!%�=�$�ۦL��}��C��6��	��.�;*�w�0>N�C�	!VY�����GG>���M7(��B䉊<>6�@��O���m�� �:2�$B�,j�j�R��F�D�hj䌷?\��D�.6j� (�OB�N4� dE�aW!�d�G��颖&ģ��[��]�!�]/DS��ȖLL��Fс`ˡHw!�D�5,7�QVL����@����!�֐y�PH`C�H�`�\�A��k�!�e+�<*�p��L*5��@�!���8`-��/F��쵙�#1!�$Y�m/�h�W�'�n� �Q��!��� CU�d0vQ�)��A7M�j�!򤑻h��5� �;+?V	��@;y�!�Ԏ.�@�ŋD�f�J��
j!�d״l8!��*���"q�Nz!�$��tB�y'@� �Y�~!�� �x�@4it$\Z���C��P��"O�uce�T;iN�9s�eյ ��'"O��82#�	K�~t���P�)�"Ot���ŭ���c���L�
�"O���aB�W�	aw5�]*2"O�u1���I�d��4 �7�ڌZ"O�l�fOG� Y�1��A�
?Ѳ��p"O�d��j�;n�)s)�(q��K�"O@�#�W�Q����^>�b=;`"O���tę'ir�es�:0�>-��"O
��ѫ�&s��8�G�[�´S"O.��̛$c(u�"E+3�`5`�"Oް�%��E��J��P.�7"Oܤ"7@.2�"9 ��/C��7"O�L�wΜ:�ٹ�d@.g0���5"O�D ��S�[g���wC�%A)l�; "O�T�&MX��Q7�J�EL��"O����$�1m�+*$&1�\QG�~�<�bK�+��P�5eU=?�1��t�<1$"U��zs���J`��PC�k�<Q�'�	3zB� "��1'B][��3D�� �O��������J=�G0D���7h�$j����(�O�<5���/D�X��`3./�	��&I�/�)�r@ D����U�me����X�frrx+a�>D�4�g�ڿptdI1Mݩ"n���+?D�t[U�&w88�P�[�R�r��/D���wB�+W=*��H̽7Ur��9D�L��ގt�ŉ�
�&�`���1D�@��K�j�@����?ht���("D��9��F�1�p��&�=�|��n.D��X��`b>dI����b=����(D���&�8IF��g	�t��ru +D�8��"��b�"���-���1�)D�@1e�h�����M�8��F�3D�l�&�U~�b-k����dճ��.D�lC�IE��xT��![bO�)SA�(D�<�!)� =|DH!�d�!O�ƅ�bb=D�D�S��&Hb�9jқ{�B$[��:D�jW͞�H�T��`�R�d���t%2D��𒁒#W16����kT��E�4D��$`��e�#ច3�$�À$D�����m��A�I�m�� �"D��[5�� =/��c��ض[/���I%D� SM�C���PQD�6'�p�r-D��K$I�j[��.1�&�(C��
4C!����d ��e��~j��
�Iܫ)C!�ٻNO�ԩUoځE�X��t)!���9­�V#�(��9�m��7!���>O (��ц]�Bz�C��׏=`!�
,���p���bǄ���I&@r!���w�P�o�q�2�1�@�#_!���6\��+�3I��@���&J!�$�f�X�P�`���S�hJ!�đ2,`J����BM�ZXB�g�!T!��
��H-Q"��bؔ�БE�*4.!�J�`��$��l�3�N�)���Y!򄁽o�&�+�H�H���@��#c�!򄒳4S�$����q�*l�UfR$ j!��fu:E�D*`���f#��E�!���Y�%L�\�D;�b��_�!��1a�F�R� Q���J�O�A�!�A�lr���4`TBw�*�gM`!�DM(�4��ūN	h�3\!�� ����G)?B5�F���+��#"O �cgV��м�p��j��\��"O��@G�@�@A�o]M��r"Oƴ��Ũ]�"Xh���<-'�yav"O�qA�W	F�0:%��	Q&ò"O�� �Ŗ1h��iku/������"Ox�� �_� p����� E���F"O"Q��i1��<��J(c�&d0�"O�E�W��8��/+�8ˆ"Op��S�E��:'�pJq
F"O��`�aA"F�����jZ Y}D��"O��0Ğ}�� b0�FO����"O%��L�6X�ʩx�ㄇ2��,	C"O��:'�?�h��њq���`�"ORq�QF������Sȃ�N�"�w"O��1�mΑP��)P�� >h���"O��s� �`�����E��"O8L���;%�b�Y�%ހ���"O�������$I��E��}�2��"O�, p'
]��R��	1�ڭ�"O��*�,C��$#m�025"Ot�vf�����,�)�$-�`"O�|���+i<��jły�"@G"Oh��#��<�%[B(�1:��}��"O���v)ȓ )lQ �gB4,xz!6"O�@�`@ΑD%�6Ǘ+�x��"OR�[���h�p)�E�90�0�{D"O��$&�o3&@  � =L��"Ov�I���W��E)�OKN��9P"Op�����:2B��"�]�;���u"OlZu�^�P�}��X/*I�"O4pA3���(Ы��d�=�U"O����D��r�n$H��A ���i"O�����Q�`��S��t��"O��c%S�p@�3�	Z�vy��"O�m�-�m��Qg��;	q@"OT�P��7��U�2��k�̐�$"O�v�ۑ]d���gԸ\4��U"O��!�أ!�T0�E��]����"OP�䙈uP��# �� ;=�U�w"O�5Q荙�^��Ղ^9Z;��Ң"O~�4 �,,�L�I��2"Oxiu��=~3|�cΞ0;� �"O��)��^
������ >"e.��"OL piУ��<` �O
"B����"O��+7+�F�<���͒�pNBE��"O����x��,��J�1)��0�"O&�Aa�)�����J̻L�h1"O�M�w��:X`��d��<6|��"O�s҄�:5 �B�.4�䱘�"O"M���#��yc��O�f( "O�$s��@>T�0Z�c4[���Bw"O��Y�`�,-8�`b�-h�^}�"O8��8=��ᢌ�_[rMB%"O�P��`��*'�%� �ǉOM&��"O���&����EۚV:Q��"O��##F�U����aM�;�rq@�"Ot(���sL���<��-��"O�}r�����`���&��%YU"ON�[��cD$#Vb��Da0h��"O���5�ʁ$�)��B��C�����"O���RI�hXN1!A�ҫ	�
3"O E��E�S������g'�,�P"O��(6���7�ʔ���R� `���"O� ���Bس1݆���Օt�,���"Or��E��5��%��Ż�"O������(A�gjI�O�P��"O>�"����cƊ2$4��"O �J�V�wU�H�.� �Ț�"OZ4���R&��f��O�#�"O(�� ��A*B��� p8t�r"ON�ё�0T�,�R�Y�d����"O"Aᢍ��U�V1 wI�n��G"Oz�����H4��!�h��Vi~!�"O�0�@WK���S��(ED7"O~���4rw�-âM��H@j�b"O�@8�	��H��͘�/��Ka"O�i��E� �e�wPD x�"Oрb��/����J&j`SA"O��'��(Y��X �G�T\���V"O.�0�Q7��h�	�15���"O��b�.�L@8�C#>&���"OfԠ�*��IJ,� fE&0b�yg"O<tk3��>4��"#	h԰ې"O�P�$���-�@jf-�}>�s"O�4�+��R����A-^;���"O�41��s���ɀ���_&8P�F"O41��wG�p�c
`����"O,��Ƥ�Ada9ǣ�) 
th�S"O���c�Ae \("!ĺ\��"O�q�ă�4�ԢU���b�,%2�"O4���h`�MK�l�:��A.�yr���i8�o�[��A����y��3rq�S�	��M�`!T�_��y�iT�{�x���i��K4.C��y�,�2w��87TX��r��ȶ�y��qx�cVp�"c
��y�gS/wі�Hi�Kc֙3vG�yB�RD<t(��ډi���⩌7�yB�:5<�<ѷΌ�{r|ݢ/ϱ�y�,�v!�p�AE�ioP���$�y�����߉\���s�+�jfh��`����J��f   �?ɸy�ȓ{�~���l���Z��剓!���ȓ~Z���F�)DԶq{�_	[��ȓ-�Ό��ҴEt5�'@W�Y�ȓk*�8a&B�3�����D�{V4��jz��giַͶ�p�An�A�ȓW?^�:֦T)w�����6B{N\�ȓ2�t�@�Ț6|؂2��j%zL�ȓC�H)��k[/��K)8�)�� W��@�G�z��J�
� mȅ��*���tb
$[���
�.e�a�ȓEH��k4� �\:uO֍H��i�ȓl�d�Rj )zp�2h2[�Q�ȓ�.���l� xN$Uy��� �V0�ȓ?�A fb�	8���b�@_F̇ȓ�J���	lB��3c^�}r	��
�H����Rt���FG5(A�����E����%VR�s�E1���ȓ��q�S�II�ʁ��i�)=����{�hs��P&V`�˃�B�PX�U�ȓ���Tk�:b���Q�A�x��ȓ P���"���F�1۶��`F����IR�|Y�����r㩁�x�bІȓ \�(���Ӡ�~"u(�%l��m�ȓ+IT\J�#Ȧ|�9�aS�<V���ȓ3����j�8&���!bm��cm�P��S�? D�&h�&���� �Y/T�w"O�0���D�@1�4`�#7*i��"O䀲jG���@bo�2��s"OL��Ba�,{:ܡ5Ė�~>�I�s"O�L񦣛�^���9�39>��W"O����3(D,$ Kӧ%z��v"O���Y�VP5�ʬY��Z`"O�]�rn�Iۀ�����$
��f"O���1�ݢ"S���,N(t+d͊�"O�ų ��)��T�����`*x�4"O�CIM��V4��#*Dv9��"O��Ibo�)X�tZ#�·a>���"ODP��LH�h� L#�ɋ�S�Z��"O tإ
�
m����Ǉ2u$;�"O脐��=LԹ�ɢ'���B�"O������,Ȧ��
�*g���K�"O��	'i&mVu�D	���5ӆ"ODXJ�+����;�fЦG�4 �"Ohp����Ӡ��e��o�\��"O�u�3�\�*أ���z]��
&"OqQ �,. u���I�P)
"O���Ԩ�6}>9�sϑM��-�"O��(��Ru~��CD�<�I�"O���R��l?��+#�/9�jܘ!"O�� b� v�,�©��eٌ�@g"OfE��'%���au��� Ƙx:�"O4����p�
&]�q@ ��"O��S4oZ*=�|U�f�-RƌK�"OHd�g�]DN�
B<7\Q�"Ob$!6c��^�@4��Z� `���"O��R4B��Q&��֤	�}�t"O$p`#hE�R����mH��6+ "Of��P�&| �O�62x�Z�"O ��^_���`��<Z�L��"O,�ڥ�W<�2���%U��3"O���s���>��#lZ�i�"O���ӤL	��+P��-V����"O�sP-ԊG	։q����O�<P(�"O0�+�N�lF�(���1v�b-)�"O qr��/?����Eй�b`�"O���20gK����R&mn�I1�/��<F�''
8��D�2H1��@BDY<��3�'X�8�@�U��ē!H%,����'��-� m7Ux�+!	� <D��'p0�*
�c�*Q��=�jI>��ν��<�}��m\>@}�rG���]�~hqr��Gyb�]�v�t)�y��)]�d���B+�:���μf��ɷ>l����.�)�,vZ�"֋ .R��AeN�X2��r�Ũb�
�*��T��)��� ��)p�m�qv#C�lRl��q�Ȕ8���6Q�<���v*���Z�"�0���IE������#<ب�"b+���`YdoX<[�<ʓ�Oc~�������mV2R��m�&�Ǹa�R$���Ͻm�d!+����0|b�I
�k�Me�N�uv��:ZR|��4%5����q��;{H-"����~�K|�uJY�P��Ͳn4}�X�֎˕Z���U,����S��M�;j6�Pt	^�1َ�I��٩t=�$i�F3�	�0|2�K�MlY�׎]{f�J�B�Q��P�X�J|j%N��l3�Da�м��D�P��	2ê��?�~��f�,1�U(���:^�2H��TV�<9��=A7��hS����H�{P�BR�<��,ܭl���3%�}�!�Wn�r�<�.ՓO|���&B[n<HU��n�<�r`��	u�0+ �Z�~�v��C��l�<��Q/b��
3鄷#z��3���e�'~ay�*�Hx<��MՋeB������y�F7&,� ��'����FL5�y
� ����$�T=k�iV�y��Mb�"O��1C��7( ���0(���"O	��"�9:��]��m�6$�	�@"ON�)�'6���(�i�'n��0�v"Öq��^z�l�	H�<@����d"ONm���ߓ{��q,J�|d�Q�"O�� �,�#`FH��̗vY�b�"O���S�ƞDj~��ɍ-s<���"O���c���	������y0�Ub"O�TI��U)1XP��9x�@1"Oȸz�Y(�2��)��5Be"O�]b.mjn0ڳmL�0K�H�"ON�
ce�@z2�C��,T/ܬ2�"O� P�'G�8�4"xJ,{"O2y��s/��Jo��&���'"O �q��N>P��MC�" ����"O�Pk��%���P��e��H7"OL�0�(]��9R����E��"O �҉ZU�����
�%
�}��"O
��AEߤ>����
-M�|"OD@��gӼp�¬��J4z��bF"O,��6 ��t|�أ���Hx9K""OB�@��}�^Q8j4��B"O�Lk2���\�s0g],+`P�{�"OV8�քS� ��P��8PL�(�"O�UYUb��U~Ri��'���Q�"O�)P�Z
7�P�M:l͞�8�"ON%q@�"/��J5�>�A)�"O����hM�C��XX����_Fl
�"O�1C�]�S	b�c��B#��K$"O<܉6�B cr@A CdB%�
m�e"O��؂Kώ�6l�K���|5"O�q����_p�(�2a_����36"O:0�5䉻i;>�ɤ"')���q�"OpK���8�D����GQ��yТ"OȐJU B��I`#��|T�"OtL�� ߏt9Z9I�O�D}A�"OL�ySG�&8���q��|�䲄"O�<X$N��]�t�igʀ�{�L���"O�$Y �ØR#`I ʙ�;~x])�"O�5���-�� !B�%>�I��"O��� >:���Q�m�|�uzF"O"�x3,c�P3ƥT��;f"O([�DU�@NA��g��\����"OP�C���<ʄ���L>@m�Ts!"O�qY"�ߕ#"V��ܼP\��`"O����+ S�TpWʝ9.바��"OhE �+ѦZW��(P|�*h�R"O��eRP�=��7�hI!�"O cC��%#�B���eڼ5�����"O,�(�=G��� ���L�(@H�"O�$�2d�h�4dw�r{̅:�"O�x��O�t]�
��* ��y��_=�89QʔS�ڐ� ��yB�K<F ��ʧ*�2OKZ��rͲ�y�m2Yih#)� I��9b`ݶ�y�J<��0�:qb��a�@��y	��k�0��a��,`���Ja���y2F~�F�p���S��AY`�վ�yr�L��� d��a1��q�ӽ�yˢ&u�����C/`�P$� $E��yR�Tbj�!��T0ڄ��,�$�yҭ�P�Y��c�%QP���s�O��y���=8��;��	�8BY0�}�<� <���׊q������JFp4�c"O�,���ŷs�ވ�����3.�5ap*O���e�9Ea�
��\`�'"�����&M���ˌE�@�C�'� ��!Q<r�� Hg��9.m+
�'�p�����7�^�&�?*ݖ`Y�'��=����-ub�	�#�z�����'m�Y��A�k���E��xO-��'8�$qJ���t�vl�4_bΩY�'�J�0�Ł��aBG�W��m`�'dp��FK��Q���H�>�E�'  4����>��Y��(:,\���'�z)1�cȧ��*UJޡ!/Li��'�E�'�§j���HD�^�J2Ʃ��'�fٹS	��,�æ�xa��{�'I�m�u��6����E�o�p+�'\X�7ɇ�ow�9*���`��AS�'�h�K��4���F�A_�d���'rh��.��x���LC%V}8��'�8� �Kګ��!P��G�M����'�REHq �/4P��gX�L��L
�'rn�`oV�ܳ@��H��
�'���b7�ٹ#U�g L�9�|��	�'6���KBt|}p��2��	�
�'�8m�sKB(���4�69N�z�'����1�E�MRp���3�(9�'��d�V��M���E;�}�	�'�N}��
�l^�Y�GL+ Q�t��'�.y��G61u���	�1u��1�'�`P!�R�l�L� �o��k����'i�h��ɍ,�~3�/ݖa�@��'�ny�E�H5*�@fk�l�����'�B�y���5b�K6�ːz���;	�'K��q�jNx����]G��q��'O>!B�l
�M����"��<��`2�'W|���/����5�ʑ4	�(�
�'h<|q&¥@�� Vk�#�f��'�J4��Ǉ*_��3���*`��'tlQ U��-��Lha�1�N�2�'ld�I `ԫ\��S�iY�_�����'� m#d�݊�b��g�5H�p���'W�|��$Ō`]n���I���'S���ǧ ��cM:q� :�'ʦ�qn�3Tea@��
0��)"�'�n=+uL�;#/��bJ�$ݺ��
�'����qe
Or�0���L���ȓS�<��`D�/t�1t��C�Z��ȓK����&\ ���Q�@e�x��X\I:+��s���AQC�=����K�>���C^~x�ۂ蜝}Kꠇ�[C*Sh�� ��X� �K��x�ȓ9O�IRp�2qV�%{�A� 40��L(Jxg��j~lx;eNb;�y��y�0�t�%�P�kE�F�|���ȓm;D���>8�r5�1�O15Be�ȓ��<��bD�o�^�SP�4~.�Y��eH����X �Qs3�-� ��M�r�-�I���� �*�z��$���a�郯9����XBT�A��5�n�EE�'*XD�@'�3������f0I��2/"Y��/Gmp���'G�<Hb�͘^^3#��1I$ʕ�����2�X��X��$��1E��I�ȓS�ư+2a�� ��oC���S�? u�A�ħ+� KO�_j�Z"O�IYB�ߢl<��Dt��tY�"O8�	3�¹h��z�.�.9��]b3"Oz �6A�H]�b�,�ɒ�"O�ظ�n��,ش��Eg��V^�"O����`�3�p�2�(�Vيc"O2H�S`�a��f�LP��e"O�	���e
�� �+�%b��d(!�$��&�Dd���~�:��T�U�R%!�.Ex���֎�'�,���2!�
.u (�#�>R��`P��I2ko!�ބW��\�AѠ��}0��֎!��D�~	,4�������r����P�!�ߓ�n����$u�3��ي?�!�w��Mp����>�* ��� (�!�D�	\w��@f'�=�X�� �!���,�t�B�'�ܽv
�h�!��E:�ج[V�g�M�T�R4�!��T!8��m�r��m��U�7�E�g�!�׉�DI�]�}��(6��Q�!�$�Ixy���t�Z�j�1F�!�%\�f�a�Q�y׊z��L5t�!�DU�0�t�QT��7<]����A$�!�D�H����Лf2̲Sל"�!�d��^�4�6EIv0�7ki*!�$1I"�A�F8F�Ī"-��8!�d��&tv��WgM/E��Ȧ�Py�ءa?�)�M��'&y*d�ڮ�yrf�
���DF�l8�֒�y�B[9viM����H�r��:�y���r�ة8B��6QE�k�E�y������Іޡ2� ��� �yR(�)o�UH���h��@���y�i�-@�(
�*	�j���3C�y�����҃��2��pi ��,�y��K6y�(!t1>�'	���y"V�8|	�S�� �@�뀍�y�<8;�q�Dqm;&��d�!�ߜR�~ٲ���%M�*�'@'�!��5G3^E�G�%�n  �hB�	�!�$֘�ȡ��d��B��mI�Y�!�dJ�!.4��+�?��(;u��SX!���Q��
0��+�����;F!�D�yw�E��̊�yl��H��!�P3slZ��«V -s�e�JJ;S�!�$�:��CS�N�ȤٳC��>�!��:wݎ�*����_HU���sx!򄄯{�����^'BR��%��Qj!�<L�
�+�n)G�(�k��p�!�d�*0GB�{��O�cj�P���6QO!�\�=�6d�C�r�"Q��aV8R�!���X�. �e���X�r�A�&�5!�$�O;^�s�m 5S���9���!�D��2HB��A�_M��; n32!��˰EK�T��ϫ.� �I�ķ	!򄊵I�D�C,�	��b!����!�DL�6���W#��*`��F�U�!�^&V��*�
��]�U` �.L�!�ҏf�fDcK�lYfx�n F!�DA#��%�V@��x��V!��X)
�jIJ'g��?0d�F+��!�䎙�]�CkW�	&h������!�J�+��h��_v��*��E�XV!�DB� ���^)2
_(��"O� �Q�N�r�% C>��`@�"O�t�Ώ{'R]�ph�FHXe��"O�t�$���u���Y���}�"O���A��	g~a�Qχ�"��@
�"O�}`��g�mIԤ�.b�e9�"O�qC#�5�]�2ꆾ�M��8D�|2�
   ��:2�
f�<C\�b<�(�%�2�$ �cm�m�<)��<Ȝ��2��;*�@��i�<��՟*'�Ii�b�B�I^�'��&��h��\��:���>{���b-D����E��w� !-8��y4
�i�O ��)�x��&%5�n)�Ə�|�bYq�'ғ������3���8v�|G�����-�#=i���O�,��L�G)2��d�D��4�'��OԢ}�A<%q�	��@�A�9\���ɕY��݅��a�f0H�� 48'���fڋo�C�Ʉ,c��(��8��3C�юC�I�Z>}Hf�s+�j!�R�D�.C䉴U�b1u�P�l�9׌C��C�	lL�`�
}tlzҀ@0q>�"�S�O&�!�"\�h��ke��Pq��'�qOn���i�HJ1ʵ�
�m����"O� i�)@6M�Ib0iL]�nԣA"O�!�	͘;�&�!'���S�2(bD�D �S�)B!G���g�i�����X�X��D{��v�!���:(fN0����*̪��{����>deh"�&9e5\yp��v��=E�ܴ�x���,̱L�����(c�rԆȓU��,hE��.�4x��/��DІ�(�$�1��e�(됎X*���)���;G(H�@2� �^R�8Ub#$��
���&x�"�D�Lc���C�#�~�'��)�Cۃ,�HX�R� "/�����(On���B 2��T���N,s<mH�"O���]�w��]�s�]/W#����'3!��_�7=t8AoB�>���`��H�!�D�$_��xmʠ3��y��l˿)q�}�������
�9���@�U�<�؜!�-D��a�%�|����+�n������7D������^L�(3䎁�z�Xa7D���
�R�$��kY�>GZ�;2 4D�� �BΜ7
ոu�FNJ�\�yP�"O6t
s&G�X��	Q4-X%S���P"O��[p���B��� Q���V�OH��D]2z���H�<Vre�e/	�!��ʦBo4qҷ��'����FB7{qO�����
n�:�#]�-�v(�SQ�!򤆪xIriYց��(�DXH�a����^x�������w���G�[@B�e8OPJ��dI�i�d��H�]p���\J�!��\�'����� �	��m��m�1O,�=�|⡁A�U����1��i<���'�I8��$���.ƅ;�,�ЦE�f&���#D��K��7
�y�s�a�0�F�!D��8�l�/
ր�W�K�b�&)A�	?D�Xr�
������$T�B�E����<��'�qO�2
��Q��ν:�>���Ġf���$1���  Q��q��r��i�@�R�9֬����<��OdU�'/@<��t�hPR��<��"O2�0@ I�+1�xcDHQ�:�P*a"O��!��ABtH��,**���!�'��'w�K�j�@��"���JA
�'P2ԑʙ' ����b���m 
�'a�A��E��S��s�hTBH8�
�'�0ɘed���h�'n�3��B�IX	�m�� z�:98RF��Ƥ�����	�Z����Ǖ�{����?q�E�IY�!���7g&�����D��&�����ʁl2��y��ڢ ��u�e;D��Xv�Q
_�|Z��F�QJ�y9ņ�>�I���O���$խ0�ġ�	u� �XPB@�r�!��[�n؎����O��t��#	+9v��:�O�ܨ�$H4}�4x�)ڃL0��� "O 9Q,��r*����&!S��c8��hR�9�vE��Ѻ/��K��!4�����& ,�c�"�e=~�r����x� �R�nQ�q��D��k�h���<a���$"L��1@�4+d�ȳ�ӹO�!��	4јP��B9oI�4����'�:�IR̓i���5�.Y����8d�0�ȓDIB�[�BV"+'n�H�	'V�j�IDO9k1F�,^<2i��KY�B7�4p�"Oր�6��0�R �b�S�����"Ob �M
�5��\HQL3R��U $"OH�0e��btF(��(Y: ��|�c"O��h�+�0/�Ѐ��%8Y�`]�"O�M��jƠ7�Z�S@��.��%A0"ObES�$ۖ O��БL��/�U� "O(�Kd�:R�#$L���,��s"Oʬ���C[���,]���@�"OR,P0)y5nU K�!=Խ�C"Op!S�(�Q��UA���~�#A"OdMh&fZ�$�8Ep��9��Ѻ�"O�}iѧ߽f�0� ��1N��ZD"O�a�7�Z�x���{�lM9�Y�"O<�Bu���"��|�P+X�4��1��"O�-˶���,(��#K�8"s.u�P"O��YG�D-T`J�j?*r����"OzI���ߦBwR���Hęo.���"Oxt�A��%HX�!0����Ya&��"O�r��΍0֒���@�s1�<0b"O�L�/ݶD�tY���^�@B"O�mqP`ŕ�~�	� �Lv�yP"O"Y��iʜ@�FJ�X�0�T"O  �&xY��߶�X}:�"O� ��U	�&1X`˗ǒ#M�v �"O88IS+��v>"�0�fI��,U0�"O�9"V��N��u)$Gº8�F$�V"OF 9�d�<v���@[:7�FY�"O 4*�+�1�2���ԕc_�4�"O�5 ��#?�:	��B�S*�Xq"O�%P�	�?`��(��A.�`۷"OZy)� �g�<�p��)`����!"O��J�D�.	��`A��5n[�="u"O���GU'xPV �B�W��"O�U"p��Rz8�H oRD��2�"Ol8��K
�A.��IQ�:r��A��"O��(����5S��D�t��|�"O�9)$A��0�b'I�p���{�"O0ђ�̐�M�<�l]�p�0"O��P��U�M�����+�����"O^�Ԩ�3<�hY�$(���Z�"OX�82%V��T�q�C�(���(D"O��G�5�%I�ȊY�v# "O�t�$�O�4�l��NI}��#"OFa�TO�@��DIc�+ `���"O�Z�  ��iU�b޶� f&�	\!�S�)r�� ���%�����>}!�d�2cA�T�%.�
C�B$�a�?!��Hm٦Lxp�<`�F�{���!�ד'"�PsH�Wݜ��b監Z�!�D��Ag� *  ������ �j !�$�y�tz�N8��Yo@š�1l�A��Ӹo8��(�n��y⡉9Y�y7YW�mѣ�yB�]B�L
�C��e�� �=�y"c12"h���0,,���e��y2a:7��ȹD��'9������y���m�8���-������yb&˽�jM5M�<1:��f���yb뉽^4��H]
,S.������y��7]��4��D�1^�Bh�P%�y�ET>-l,PȖÅQFI�g�G5�yro֪Z>����'I�z��ŉ�3�yr�ޣ.���l�%�� BE�E�y��.5lP�Ƈ��$�,��7�,QJ:�B�F����h��ߨ|��92�k� &�,�C�O�!�$K	F
�:lD�8����zH�ݴF���-�E�r��	$��ze`�!�`�	�f+JE�z�8r��J%�ƭ�~��Ԣ��F�(KalH��y�#����jg.�B�2��B2˸'��3�a�l�f铯6�`���oZ
]��$��bA�7��B�I�[��B �I�GD�h�!"6��څ��#ʒ k,O���Y�@��mµjI>��bd��%�&C)D�8�e��E�@q�ʧwFT�� �Y�D5 �D���hj�^�H�A��>�����¯*춱��*9�l��0+�h�r�oڻ������M'	�����z.�s�<��j�v���N���+���Kܓ{L���t��$Q���`���`�`r��1et��˦�T��!�d%+�4����&< :ʓi�]�L��� 9K�i�'er1G�,O����ƌ"�R�JЯS�����"O����H��fQ�14���P`���Q�i�9���J!��Q��I��(��Si�B��a�g@W�i���d��zp���&|�c������#"/�>i�)��O&D�,C�~��K%�Q�@�N��dj$D�� D�Ρ]Y���N�<���O�ʵeZ* �&�O?ա� �9E�����* �t�>Ա�O�h�<Q0d�#E�2l��>#><=H��l}�![�r��١�Bx���"��9���%�"����@.:�O���V+�8k>��� ���r�.W�j���O��R�8䀑�LlH<� !4���3�EIےiD�Xn�'ւ���@�#1�������(��L� � LQbhiWI�>�!��ȲHx�R1[�7<t�󓆗�;q�$��"��*���yy���'(MX�@E�+�,[@/kKX�<�j�`���DWN'(	��N?�ՠ�5!��LZ�H̰<A��44�峳�N�,5��� �HE8�܀b��$ȱ�S��%v��2��v��@�4�Y�ē�nDb��ݗ):��
!���m��EyB!���zl2�\�+8��M�,AU�آ�Y<|Xl1�"O�\1�R�[p��Cs���]R,��I,?�+��<E���)� $���4���5*��v�Ʌ�T���@c�[�Z�d���"���'�6Ųv˗�:`D���	?v]�H�e�5I3.�Bs�C���������s��m�`�ե֬U�N� ���Cf�C�	s�� �$�تښ9�� 8�C�I~��(P��}���вq�x�)܌�	�n���R�x��צ�F�ء��I�{j�B$\�غ�IV478�.U/aDN�Z�%D��Kg#G�rtP��(���9Ԧ �ɾ>��<���:z2�M3̟�v�)��.ɪ�t�^42���P*^X�H���$t~4�R�Y�bt~��6b@<��Qb�{r0�$���I��H�R��kM6�~bÒ[�Hl���[�"ʒ��l��y�e��Q����/��&tLx�ǠS<�?e�
+�n�Xg�6|6�[����?��O&vHp�瀳~z���
?��d��I�Au�͉�E�\��9�& M>���-�,��ÅT�"�x�R�|����N���� �o��4k$���>x����U��3�.'���K��P�l���E7$�`��h{��U(/8�5�t�Wyu�9�h 7}哌_I���̜����H1��^����X��؅�ahڎT�h���]�*��!��3D3b���C�m�<������Ǽn�2����.���A�B;jĻ�ꂘl�>東<^���%N�{��1°k^0F���Dކ1E�/Z�jQ"!�N�P���x#�U�l���S�@�$��8[EJ[�7�P��fOʺApQ:Q�'���(S�T�j�{�0��ʁ�H!`92M)���;庄����>�z�2ٌIY�(ДG:)��� S6�	�����H
��v��8��
i 1��O�-PW@[��6!���|�=�@]�	�����L�8U<������䦭{�z[��rg
F�7��T�� 8���ge�)��Iү�T���C��11���jZ1D��
g#�>N;�q!c��B����D�03,��J@(
���#/��a�sc�H��*M�P��6�Hza6���z ���`�O $�~�F�l}���t�S�Y2���u���p>YV+�$P㾈A���#j�
�)��x�\=i$�	;Jh�f���A��L��(�D�@������Ğ�UI�K"e���te��DM@1���J�J�4i��(O@Q&�� @GV�"�!N�F�*d��fS�<`�`î.Ghj'�w�����֖g2�o��,�u�F$4>�8A`I������#Xpxl#�����4��,n��(�U��$5?�Ͽ+�C�/����ҕD2flKAB�m�<Q�(Ʋs%��)��<0I�MK�N&�h<#W�Zp��[S�#�"H�'�HO��(7+[�z᳠(�38�2z�'��4� ��&x5��r�jȴ{�2�Hqj�4|ր�Gg\�!��d�����a}�6r
Kŗ%��d�C,hаEy�fr ���Д#��@�v��i�S I�����
a�ݪ"V�h��B䉊F�0�Y��Z�B�te�&�A�Z�֨`�h��ay4,�ik��
�h����5dA�s����P,jݸ�k�)�y��)y����'g6�؀Wꐃ4+j����ɑ1��aJ�}�p����@�q#�& t���,Ta���*B,+�OPA�$ؗk4~�8VH�#^�����C~��q��P��M�#DK�5�}�ș*gQD�1�Y +֐�T�+�hON,R�j��r�Xvh�4&5 �'W�����ݑJ����&ɜϒe��y|!��'�� �(5�$�_�B	�I"{� P*Mw�U�Qm�@�O�b�:0�!&���2I	�;�<�"w"O���/�)eڄ�;"h	=�H2�l
��~2�]�@p�X�!�R����� e�t쑁��?��J�ы.wl����@ɬ���������&)$	W蹹c(��/������6T�ܣM�
�hH���ax≚�m�T�=IP��;���Cޢ��}k���B�<�&h���t�Y��ܚ�r��J}�<ِ��e����T��:��8��+Tl�<A�k�Iy���b��!Mt����L�i�<� >DЂ�̤?=�@8����~�U"O�A��O���+��p<t1�AE�l�����Ox<rc��R�R� �҃yu�y3T"O"E���I�Ro�(+�*A��H�2�>O��	�&ϳp����B	z�z��� �U��d�E&)�{�,X�}"��ɦ�#A��Ayz�r %U�z�J�
,#D�``P�O!0q$���
 ,�$�!���G�4�`�Ϟ@b�>	Y@�I�I� �҆���Gf#���` ��i��@'ȭya��(�hA֍�x��Y�ݙB��O8�}�exz�i�F\")�d�E�Wc` x�G�TnqO�}��_ՠ����Z:Hq*ĩȯk�Ե���{<���e��&@�a{R��(TT�X`H�,��D��,�	�?Ye Č �>��8�����|Ӥ	���+ra���"F�W0�h��'fj����g}2�X
0�,��D���"��@������'2� �/G�fQD�$M�pZ���ń�/'�����!K���'Q8Lq��Zj�OVhYݥ!���Ao��W��+A%�V��E�1b=}B��PS/?�Zu`l��F�	�Ξ�6���È{B���MK3ym�EW�� t�fE��k�0����s�.	��I�e�H�P�R#62������Vn�	�.=�቗E��2`3O��u 
Q9��ƍA!�*1"O�IH�Bܙo-���"M�r�
��"O��h��4r)zU��E6��"O������P�9���P%ڭ�"Oh�adM�n�,k�KI�q3"Ot�k��2QT���U=.		P�"O�����Q�N��G�([�m8�"O:��虸Fш��ǂ�'����P"O�t�7EԾn����\"�� j�'@�����ff�Ɇe�j$��H�'*�t�1A]�l�^�)��?S����'0J���L�2��HF�e�����o�~�I<)���;g�	9 �iȘ:D�]�<�U �G<��$UlXb��XF�m] Zä8�)��\� P��aP?z0A��[	A�B�I�)�T�c�֪�0�sK�2���䍘Y>�S8,AD�Ǧ�:�����97��d1TvGζH�m`0$�;��ycf#�dp����Ťg��L�`��{�(����a�az�L?
f�O�e��g�^��"���jS�4ڠ"O�l�^�G���E
?G����DT�<@���{���'�k�f�Y2&E�$�i��յ�ycP#g�a����%&%��˞�}2�Ћ��<aUa�#S��3��5�{Pw�<y�i�)v\i��M�:K�V�p Z�<��c�VX�)�5T4���T�<vNf�A�ɰn8:qtcP�<�'nTL�Q؂	��v�Z��e$�Q�<�hΒ8F�D���	~B�XJu��W�<a��8|�0�8��w�:�BV M�<�FI�B��aB��tC�Uja�a�<���K�>��u�q*�)l��Ka��Z�<��n��a�P���)|]؜�e��M�<i���E>D<�2l�?��m�/]f�<�f��m���PT'W=9��*��k�<�" ����㦊F"28k�z�<��Ή"l(Z]Z���t��b�w�<���ɬj�J3�9ݐ=�4GH�<��j1>�=("�K�lp�KG�<9�n��H̰�O���kf$�A�<����/z�����1+e����}�<�	Y*�6�����6�5I�V�<�3	��Cp�(�Qۿ/���(�Sk�<���X�U��@�YW<��rN�~�<!�AM]wx��	ĨT
2`�R�<� ��Rqe¶��CN���@"O�0���1x &J��ڱ��"O�=X�`_�$H�+P��8�"O@iKw	D+;�4x�@
</�(YIp"O�A�C�9-�� 8!���
�+"Ob�aT@;ϐ9�s���P����"O��ʧBI+<DCU�MO$��b"O�q2�o��jH6 ۝`j�*�"O�z���7$��LcD��\	�V"O�!�!C t���⑳b$��"O&�y��#P�9���4���T"Oʄ��Q� Hs�Q&#�Ll"O�ؒb�]/P��h&1�B��"O��ɀ�j$l����A�Z�t"O"�9���/�M���F�c�$ٗ"O���0�!;I��3uJ�?]����"O���,��iX~���)8�Б"O��вj�R�(!⇇9H�3 "Oڌ�D��_�
��Vƅ��V<�7"Op�j�(I�!}�*%�B$l&�T��"O�����������l yط"O�xv- �m�ff�"'ŲW"O�$P����{F� ��Ä!�X�`"OdBv������^, r8f"O.L	��T��~�."Vv�XPS"O�X���2I�z�C7	b�|*�"OJ�X�dZ,b�:	ԍ� F�ѩ�"Ozi����^��iSmG�	���"O�ԙuj��V�t a��_&��3�"O�-��%:~�bq�T1<6f�"O�!��wY�Ͱ%'K�Zq�hK"O���A ��_���FT ��<��"O�Pj���.|R9�ৌӲ��`"O�AKv揯
����V#�VQ8a[r"Of����
�3�蹐���qW�<(�"Oڄ�F�msX����N���"O8E��O�\4R��,N����"Oj9�E�V��$�����<a�"OJ�J��}�	�0-�=˰�
f"O89�!��"3�]��T1cĜ�"O@�!��2G��H�6�\�$�:|��"O��1��ʑ<J�b�G�mf��@"O>L���DJP�5O̹\t� "O44��j՛X��1��eS�+L���"O����У2�)�r��3i����C
5:C�|����#Eȶ�b��ķH�l(0�$D�����*2�$����>~��9�RDl��trf�x:��ߓFu�u����:����۔Z�\��I,~0p��FEֵR�m�м3���rx����0��B�ɉPF�Т�努W��}��I�$��XI��y�Z�r��U�O�Z�O��Zae�S�^�C�'�P�C�1a�.is�i
~~i�S�D#?��8+���<���/�gy2$M$sn4E�D�0J�����#�5�yꄃ_�|�\�}�����Դn�J,��!40���J/lO� �"2!-��B�t�|����'�4�Ӑ�(� e"�i�E@�D�<���R�Ϗ�xthQ��'P����Uqm�4�]8dR�h�{®�6#v���`�=u��>Us�T�y�@i�$�'���	sm/D��y�.;|�� G�8����Am��̬��I� ��5�(���n`���AbĄp���0�W��dC�ɺR�p%�B�Km$�@�/P�*�6��*�D� )��=9��ȹ{�`|r����en��a�c�u��LH�f�W;�]�E��;�̐;T� 4�����4��Q�҄��"m�3&��й��S�? 1xu/4SNA�S.�
J8T2�'F��R���;�ɧ�����5(]��Hh2��21x:`�a9D�� �
�*Or]P҃ϓf<�%�G�>��k�y� �!1<O]i!��8x�ޠ�`�=�!���'c�3���DPVܠ�OW'b>43�N_�h���x�FU{�!�D�2klj� �/� a�=�Q��qM0	aD*���z�' ���&�[�yԚI�eN��c�v���*%�\��!�1,�%��[�:�P�rb�=�(� ��3N��)�������|O ��oE -��f%D���/�y�|�xD�G�z��奟����Š-0�Up�˟~X�����M���1#΅�anH3��5�ON���M�Q<���' L�HEUP3�����dM-&A��'��E�M�./���ꓨ��u1��X`��m�#�,,��b?��e�K�.Z$l2��Ϡ?���ӌ(D� �# �'�Y�L�޸Ã��< X�I⁎���2(O?�d�$^�ZH���=/h؅¯+A�!�d�ML�����3[DR�F������r��3i6�y2A�+"��L���<(M����W#��>����#u��*"�ώ&;����!��3%���y�݁<PA�JO�:�`D��y�D�}��A����To(Q5�ז�yrO�z����� e�P�e��y�I�o }�����d�+u�;�y"nI;K���*e"	��,�ٔl��Px��� ,n���;)D�Z����F�Fi⢆�Z����R�'A�"D[�e��}KD_N8�DXÓ ��9�o�"`��d����%
EU*�X��j�nc1s��*D�C�D	kT$8���-t*��5+,-B��ΟJ{pp�#IX'K��#������V���Ի1<�#׫�	=Aڕ��0>�Q��/F�(�i3J��i��]0� pp� �T*Y�Ne��_�������X����շk���g�~�hHtmG�U����F��$X�A�OtM�͌'I(����o�����p�����IJ�z,�b�a�T��RеG�<��F�ʓL*�p���)�����ʾtȅ)T#
#>YkAn��0� �ʅX�R���t���Oȴh�E�U $(a3ю����N�c=Z�⥈\H��:��8���34U���@L(����-�:�|;Nߑ�8u�2k^�K��3ǳ#��%�@,�ǟܐdm;�d kb�_�|2fNI�.��pqGˈ~�4[GUV�'_�\�cmE)%���Q^��+e��?ݪ}��"T9/�tʦ�I<Rm�S�[.ҢΦhP�qѤ#T=��3�	.Hzh�iH����@VF5˓ �DL(P��Zx� ���$Pz2H���)��,NthB�� 8��|@��C�7�dq�q�S�w�ȹ�HK�V<��D�i�����VS�� �jݠfqn�ѶHσk�~�`*Kf��=:f7��ؖHQ��(iV
\#�~R����*a-^�M>������?	m��^գ�K�$���	��O��je;GmԿY�>9s��s���j0LV6r�D˓sfȥ�c�A0X���(y�����K2N#����i��s���?��"-t�,�G�'{����f�^�}ڰ�2(�o��E�PE�4 s��R�M�A(<� ѭI�Z
�KM(hJ\Q1c�Ojy"hD/6��5A�́?�|	Xd+��W�F��~���:.7�����B�����.�Y�<�����P1K�N:b2n�䈂���b0f��U�g�v�
��JG�	�X��ԡ�� ��D��F���W���r����tm��u)*�XBh�,x�jC�	2R���c�m�#�-{'&S6�C�ɭ7�P���G:]��A����8n�C�2fĥ)v��;;jN���K!r԰B�	0,d 8 F%ܫc����6��1bZTB�	(W*�ѐ�B�P݌�7k�*d��C�I.yJ�A� �JPE���ğIcC䉐-�*X(�g@�%�6U��4��B��?��Ѣ�����R�^	��B�	%m4p�)���>c�ؑq�݁�LC��(K����!9?,�ZH��SdC�	1J��1+�1jw�\R�o���hC�	 �x���"�I��
�L�!��B�	�Z��2Gm�aF<4���=J�$B�I�c~X܃�Lz�B�b�
�W'6B�I�o=9᥎��t�K�
G���C�)� 6<iP��w|C鈷T5��i�"O���r�\7�6p8!)[=s86�Q%"O�áN�*,�T�ƏYC��"O�|+��R�RwH�QZ�C��c�"O\I	bR�&�6%���04�11"O"�b0��P��X�kǂB�]��)�)*�����O�]��j@v��Тi�!?��e��"O���Z�,�j	@�b��w��p�0O����V($���Z*�HػP%��PLjR&D�1��{bA��%bL�(3���8�i�<2�(�W��0u�Ҹ��g%D�����0f䮡`�����p� �ɗ@>90�,s��Ɂ?1^-��K"8�$�Q�N�j�!�ě�EBm��˾(S��Fb�:?��D�Յ(Z��Oz�}����X�`��r~�0u�I	O��ȓ,�f�{ЦاK�9x���d��I;j�M�tAXE�a{�lS�z�P-c�ρ���d�` ����=�`o�	
��P�,sӔ��U��U��ÕB?M�q�V"O��`�f#~}�3=�2��`�dY�0�A	�H��s0$	�bĥ�e���N�І"O>�
�HG?PN]�&b�y����C��z�P��U�$6�g?�5k�����Z����A�2x��Ke�<YINX�hbƭ��-�����<���ϧd����
�i�P��r( Z��X����*shh���>�ı�1O�!"�F��������R"Oz|� �V2Gw��1fɎ~�4� "O:\�C�O�d���5�[���`��"O>m���\�̚�(�Ă�1�9 S"Ofqha?[p4��"�{7dRR"OFMSEiӌ+��Țt��1A=��;�"O�����^3-��p�p@�+�0��F"O^���f��"q����Mѧ�y*�"O~�*Z
Ep� eW&H��"OF$ꃆ��06`�� �:_�& h�"Oʹ�ѡܳ]��8�.,[L��#"Ov��?�D�1e�<&1�q�"O C��B.�s���%_ͬ��"O�A�"n�.��i��54�V�I�"O�T��>�nܰSLGL �"O:ѓ�)P�i^Q��ɍ�9�v*�"O�`{S[�16��bF?����"O��8�J�6LH���	 �Ȁ:2"O��@�E6���g�݃/�jl��"O`Ĩ!��114������}��,h�"O���RP�*��)�!u�L�t"O�m�F̎0n<�uf�{kZ �"OvŻc�V6�\{f�����2W"O���M�>q�Y�b�ђ!�<��a"O(Xf�J9h��5�:�,3"O�5�u�	j�V)���)&:P%"O��`pfıE4dx���kϖ��&"O���dA�7���2�]0(�\�1w"O��v�h��Ѓ'#U��ҕ� "O�E��I�<{�)"U/-�TLs`"OP {���j��  `��Fp�9�"O,=�ׂϘ9�8xiW�@Bur���"O�d'��	ؖ�rP?Hij�b6"O�i�ᡃkW���2Ͷ��G"O�P	�N��N�t�q�W�I��h`"Of R��	�&z�	3��F�{�
��"O�aV�ɢ��PH� ���K�"O�E2CJW�>�xm���.Gw��"O����Fބ/���UIֲ1s\i��"O \ʔ	
^�n�CRj�j1"O�L��C"|��L��C�3Rnu�1"O� ,��i�=u�Z��B�=xZ*}H�"Ov���L��58ș�ƇoO>=�2"O��3T�Ќ5>J�#�)/%<���"O��aj��	�Ti�ǈȖN��<�"Od	b7�L,p"��ѧ�ܕtz �W"O�yђM�����c���+j�X�"O�����^&�`c��x0N�q@"O�5��B��Q< �Z&�ӅM"d�Z"O����+��\ǨtzV��/'*ijs"O��J�T�2'����^�!�xz1"O���̊�	�h�q���/P6Y�"O6aS1�Nm�&qw
ߑA\ђc"O2���:FܱahD�L0��"OMR��=k�܊6�J�j�v@�"O8M��,�p�5��E��"ɸ�"O�H���D�Ei�JG�.�be+Q"O���A�oi��e�N��`�
6"O�D��Ò��8I�C� eT	��"O�e����4��PbDl�sEnYbv"O�u�	O0Cz�|�%��'J�	(V"OH���[�m;��h�%L�Y8lЪ�"O�,!e��\����Ć/GZɹ"O�܈2��F�t�R�#;.��a�"O���!I��u�8���ßg/����"O��9� �\�L��O�)+,a "O� �p�p)H7I�m �:�"Ol2�GG�^2�Є�G���HC"O�lJ��I�8¬43���i����&�&$~���
�s~�$��(���Ӗ-&��8�]�䬐��ϱ:��i�r��c;���-O�<�O|"47O���Ov��D拪+�&|+td
>�&��AOe���')� �D�?��Ģ��Xv�k�c��)r�����ZA�u���s>	S'�D<5@����=d�nuѶK3}2iC#{ɠ��Mצ��H����Q3@�4�����B��@�O����G��T�>%?�'B$�F0f�1q�%D>?�$�b�4D��� �⌵&o���/O�?��R�A;��u��ػ^��<���/+d��`
����L&�)"ҧ`��M2Ԍ��+$ ��P-�;T�ulZ9I��$�O�����O��sӘ�6��(�VA��d���B��i�Y���(�TO�?�R��<�H�if��4j�B��J�+��I�s�$�ĕU>��QlY�G�- �G�����I��Ĕc�ā�i*�Zȹ��Nܪòh;H�x��V���5�p$��A�Z>FL��Ș���� <`���]�a��䜶n�#�H�a�+�kq�Qf"�"�4�HDK���y_�e'�(�Ak�D���çU�4�7.Ջ~�@U�擄jF�Xe 	3~�P���* m�)�' �~���Z��n�{���;
{L���ǘo��a�Y��9��OlZ��ԃ�u�x8�S��r�Y��'����d #y�{�&�
k��m �'�
q���[�Oʨ=a�� �f!j��
�'�F�j%�-�h���IQ�Q���y�'�" Z&�[?x@C�g�'z)�s�'�,���U�7�|\�L]/R�y�'y�4�"kCo6z�;�NM����'/���W����dAfE�0,��'jvP�,�0s�0qq��N�e8^H8�'�R��0}�~��g�ۼJ�p��'�: �%f�58<�a�O�T���r�'�����Ί�U�=Y�D�����'>��.�`�h�ɽ>��4Z	�'��ٙ��9��13��	8;���'�^0 �@�#����࡜8-��U*�'E�bH.)WΠ1�	�8M>��'gx�	Gn̶$V�i������Y�'�&t���͞E���dIΠ��A��'�,���ZFU:X��!̄����
�'On j$*!%4չ�N�LPҼ��� �� ��� _��*P�9{����"OP��3��Y�Z��f�U	z�� 0"OzM�4D��?8<�\T��*�"O��k6��`�MBc�ͅPJ�D�"OJq)��;=���/;p,�X�"O�!��7~hi3�n �yH�"Or�C� I����S.D�i�l��"O��Cfj�9_,ez��j�>���"O�jE��o�V�C�
K>�zS"O�ሃdȆ?��8�䘍Q��-i!"OBD���ߤP1��aj�-,~�HÓ"O޹�t�D>g����:zk�(0"O �2�Һ�&�P�oMV4|��"O�PD'ؒo�`@	�n��80�Z"O��B��Zm|x�!��#Н�"ORE�U�ћ1�ތ��J̲�6���"O"���h��k���:�L 5R���"O�A���w�A*�o=�0��"Odl�4`I}
��
��y(Z0��"O�1ˆ��`�����B	h22�z "OD�cu�ځ-��4 0aґJ<`�"OnY�D�/�V��בr
:D�`"O��X��\�	�ҁ���(p   �"O�-[`�݅a��2�J氨s"O���6��*c_��p5J�)���P"O����9�l q0jv]P�"O�5A��$JO�Iqc�!dZ���0"O�1¶Ҷbg�,��A�$\I�\ˤ"OD0�A�S��� ���]5��z�"O"ic�I�1 �Y�,�,�m�B"O���X�M��i��i�3av�4xf"O
����;@ob���G /l\ր��"O� *�d�Y��F���<��mQS"O��V$Z*��B���v@J�"O��!�Oӗr��������l3va� "O����Kb� @�ŉ�%yJ�� "O�,�PI����HՉ�EbXQ��"Oĭ�f/�6{��5s�Yd)N;�"O�|s�RI�R�P0A"��"OJ�9�&��P��4"Q�+ x3G"O�}k`�R�RU*�!�;���#Q"O�=�dC	_PT	S%;4����"O�$���١l
�%2�̿A&U��"O*d¶�Q3Ҕ�"`�>&�=IP"O�I{G�3�q��;! ��r�"Or��GHV:��B�Ǻ'��A�"O��5I8e�Z�3��~�,\�"Ol�� ���
\z���9���	�"O��!�ǹs�>�9w�H^J�Ū'"O��@ĳo#ؼ@�
^C�$��"O��b0�W;��p��w}.(�D"O@��"�ɒr��!��3_Z�M�C"O�`Y0�%[{����$o���Q@.D�p1��СM�|�a�C��b3����/D����A� Űg�B�I��{%c9D����ə!H/`��pg
$�DYa��8D�\ڳLE^
�|�tF�"E��
�*"D�d�2���7��$� )U����("D��Q�]?j!�WD"j�%x�.D���cc��h���Ui����d+��,D���gC�+y�4SA�v�[$,D� 0%ɟYApD���٭Bt2}�s/=D���5*�qy�Ī��53���*Ӂ(D�x�5��lp�MyЇ0M �ZW�8D�� ʥj���Eo.�s�%J�8<�"O<x���1"�aA�
��9��qpq"Oa�C˝�o�FD+�AR�"ܣ�"O��3�.N�Qp��� 6.$Ч"O>��lO�@���6 H��)�"O}6�Ia
��!��/�JA��"O�\�kɡkG��2ӦɴCKb�{s"O2]V���L���$UK��I "O�Ƅ�F������;e��}D"O��1�M5�*�Ǥ[m*]��"O>�h�ص?�X�9���!-x��h�"Of,I��@h����#-\L\��"O$��`�%E�@;��уpH�D�!"On,�UhZ�kC��H�ƕ�n6��"O�Hq ��;s,���E��k$�j�"O��[dC�ݠ,!�@\��r�"O�2$��eI���p�T�$��QCC"O��ҳ��*�͚wɔ�d4�<j�"O,�ZN*ea^a�����=��Q�"O�t�S�vyf��牖�{�V�C"OPPЇ��H���R/�v��"O�z���^�)�w�ǀf'��
"O�
�H*���c�b	z2��@"O�u!$��!g<���G��t��e"O��(T ^�t����o͉1��h�"O ̣��,�8$N׭&�H��t"O~��$E�-+��K��_�?�	��"O"�8�)�)8a�b7�΃p:�Q""O*�C�A�=�48�D�;B� �"Ox�J�B�2
�N����t��YC"OƐ�W?(@>\Z�ޤ�l��y�F�h�!�ԋYC:84
@�y���4?������W�MCS悫�yr	C�$��˴c����]��윸�y��'�d(���^��uz�ꇝ!�D�P��i�W��]Z~�(�	�!�$߂ �����D�##Q@��)_!�G�,U�]"t�D��l��EJ��T!�Q!���`ĩ��L�Ԥ�b.9�!�dڈ&)Hsҏ-I���;�&{�!�ː֘0r f�n&�%#�OD�!�$S$+��P��V�F|�5P�Ͽ8�!�$ƬJu��k���Q[��pD��9m�!�$�-�p] �HDZ��!��bH~P۳f�P1��8P  pg!��= 8ᓆ!�2� �R�"k!�$Z�f�%�N�g����Q��@	!�$���Ȅ�FªP�\�s&��76#!�$F�4�\[�ז����ԇS�!�$A�gL	�Iܩ/������G�{�!�ė
o&��s,h{��)b��!�d��S�F�b��`���d!�K����#jO���\�� �>y�!�Ě�O4�m�$u��hT
Ǭ$�!�H;Z�(�:�eA�-k���ܞ-�!���o���@T�oL�k� 
xq!��"Y��	�#��7����,f!�D5��q��D�H6�%�GW�N[!���5Wx�
�J1?lH�e�V!�V�'fڕ�,�=sPt��n�,�!�ǼD9,�AnR�7���g�>�!�Dڅ8-A
�Y�B��%��x�!�$�?j��I+���L�$�� �ݘfp!��ҺH>���C/z��ɕ�_k!�� ����ՆOJH�A���<OL �"OXZ�؍+�5�&T�#(���"O��z�`
�~#D�#�$�`¬�z "O�L�a��Ǣ<�g��d�ޙ
%"Oĵ�G����P�9�00��q��"O�hc6/�?1����J�Y�҅2�"Op]��/�0���#c)˶ELt�s"O8����ԉ|{b `��V�9S��Z�'�R���F��T�:Q1'L��$e(�
�'Y��z�/V!p�NT��hZ�!���'�DEbwV�4�H0��♺D�RD��'�����\�s�L���H� Dz�'��bQ,ע��1Q���x���x�'�h��(B���F�C��h0�'�6��REf���g/�k>��'��Ŋ϶D�� ���ҁw��@	�'���Ԃ	גYQ��Y/��T��'���Q�+=a��X�.W�+n��
�'Z�|sDf��s��hß.r*�	
�'�~��#ڸ57Fp��#� dR�X��'�%�&#�:27��S��_S�-��'O���n]��@j�!Ef)�"O>͋G�Dm�i��dM!p����'"OFL@�b�=B�`��f�� ~^�&"OLuHP�0���$Y�\�k�'r
����փ
�����(�	�'H�ܨ��E�#g8(Q�Mc�����'���-ـ_�Ѻc$mӪ��"O���ӥT6����D�{��("O�X��-Y�I����E�W� �H"O���a��C�4,ӃN�a��(u"O�(�@*�C'��z�L�HW�H��"O:�p�(U;nJzQ�֯�14Z�=�T"O�P����43�p:��/X����"OH�OH?CF�@9��O�VT. PS"O��s`�>U�ԣf�\�B�� �"O,�Su��=+̪�@�S��3!"OX���4p�T�Au 8Z͈�"O��aLQ�V�tYqM�=��R"OJ��K)�6Y!q��|�
1@�"O �I�P0H ,8;�Ӑ:S:M�"Oν0EN������^T�8��"O���A�'&!����i�9m`U"O�,�Ge�vH�����^�PȆ"O��Rg㗭����x�$�u"Oɱ֢�'H�4A�c�����"O"�A� �5 �*AH�ݖO���A�"O�I��͛hNx���K?���6"On]c�	   ��     K  �    +  �6  �B  N  ^Z  -f  �q  4}  e�  O�  ��  �  ׵  x�  ��  ��  !�  q�  ��  ��  ;�  ��  <�  �  : � ; � "! s' �- 4 ; �A H sR <\ b �k �t | B� �� S�  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O��jg�=Pz�Aa`�#�h��!\��̇��#=B8#���fB8%pS��H�����fȉ'�$!q!c�	^+F b�ǂ!3�v|��'��EK%�ݵXF|ԲBER�/�f�ٌ��#�
ّ���5�`��'c�6vH��C$"Ox}e��N&}A�A�3Z`X�"OJi1�Hճ,U��I�	� 4Ft��"O�D�tkI:��͠�(A�Iddi��eOuH<YS@҂+2��p�T�w޵����h��\�>y���BdlcL
�g?x<����d�<7�5�)�늁yD	�`��J�<�"]2����ܿf:����G�q�<I&��d�ɓq�:Ρ����X�<񥮀�8TΩ���y\^P3�N_�<	BdJcV�����P2.�"�J�,�v�<i��1i��#P��,+=hR ]q�<���	4M\���#���:�����o�<i���3ZJ���5Y�%ԞU��g	h�<i�-
�Z����&��U@�ɱF�DM�<����+�|�h�O��i�ʤY�h�K�<����u�
� R?
Kv ça�<���.-���4��*��ZVŀY�<��ꈍ[����Se��e:��Q�<�%��$f��F�S�r��TeXX�<��(g��K�GįDlz�iU��P�<�w(]�>c�r!�*8`9K�"O���T�W���!G�Q�R-�"OHXB�X( �i#B��)^i"O"5K!h�5��В��+B
p�Ia"O��Y�Xr�-���,�ِQ"O���j�"�U��-�~��"O&���Ǚ7�l��t,�V (�"O�a 2]`��:G���ya]�&"O2K��ƹEέ�F�� F��QS"O�%�⋖�s�J�y"nԵ'��ۣ"O�Yk��z��i�`�@�p��"ODY�̙<RE��NK�l/2!��"OJ�jv�۽;�P;"�̼#j�P"O\I�/���Y�	I����q"O�D�$j�4F  �H1e��N@b�"O� ��
�/q:��W� �!��Ժ"O깚��
=%dU�f��3���7"Oba�6� "j0]H"�sΑJ�"O촁LTf�䍐ANL�r�4 T"O�LU�]�FP���2�xX�!"Ou���]�9��]ao��)��"O
�H3 ��Y��Qo�)I����"O�u�wƓ-r��@�7c��_���"Oz9T�ȧ&u�h�IK��< D"O��!�5�6���\�f�"�"O��k�eK-fCu����:���ar"O� >��sc���5S��	�C"O���I�8-��4�nO�G���"O��X �].8pw�R�u|�#"Ob�[h>S`�b��C"4]��!"O"-���[T�]!u�v%���Ĉ�?����?!��?����?1���?����?�C��J$d�bbT*v B��?���?���?��?���?y���?ٱ@�&i��(^@i���ز�?���?9��?���?��?����?i�f�	2J�x+�QEr�5����?���?���?���?���?���?���)rev\IQo�Z��=��2�?���?y���?y��?���?���?�� A�7{��9��+X,�ᑓ�?���?y��?����?���?I���?�jȍaBN��3�N����S��?����?���?Q���?����?����?��BL�`\��ߑ�v +p.���?���?Y��?���?)��?y���?��ᖚ͜�C�\�mHP�$�?���?��?����?Q���?y��?�U΋�@�Bi@rdݭn�����A��?���?1���?���?y���?����?���<��� ���m�BE�CG��?1���?���?����?����?����?AR ��d ʽ��  T�6��'f�+�?���?����?Y���?)��?���?�֋Z.1P�u�#PR��a���?����?����?���?��dQ�6�'
RgE/\\PC񋄇6\v�{�eN"�Tʓ�?�)O1�����M����]xb�� B�av@ ��ŕ�P8%�'2�6m&�i>�I��q���S� @p�f5�T���K�����	3�Pm�[~?�ڱ�S}��[�#�d�b��-�,��`�1O.�D�<���IĆz#B-��N�:%��y�D��b�&�lZU'�c������y�ǔ���1��D	7�����J ?2�'I�Ĭ>�|B�E���M#�']
��s�R�F�>e�㣕�m���'�����6�i>q�	�9k& �`��a�����+t�J�IByғ|��w�|�kv��n�����Nd18��U&���p��O���O6�|"�Z6D��ؠ�TU�#����Ot�����G�1�t���G�J�$�(w��x� $�<{�v=j���� ����O?��6fH�ً���y\�a����Z�牱�M�&��u~��yӎ��Ӱe�p,�'e�Np����42���ҟ���� Ӣ�
����'��i��?-��"M�SD�K�D�2T��h��?3*�'�i>)��ڟ<��ٟ��	G�9c��*H6��A�F�]��P�'�\7�g4����O��D4�9O�)��L�e�=�"�Hqǀ�<����?�ش2r��T�O!�t�ϸ!.�
�A�:_�:ӎ�) ��R��By�l�3��� AC�8/�Ɵx�!dʓ2�r��M�v�"$�O(
�����?���?���|�)OFqm�)z�r��	!��s�=|�j
�NC D�J��?�M����>9��i�7��O�uʒ V��q��o��5@�iM4x7�v�l�CԦ\8E��$A.�i�	�?Mj �S���nϨ{���h�A]�n���H��d����ȟ���˟ �I���Jg�̊&\�c��NF��5JE)��?A��?��i1���^���۴��S��2��	�0"cnL�c��b�yB�i�,6-�O���eӐ������ך���b�	B�+��@b��)r".ͱ��'� Ȕ'��7��<���?q���?��M��A�}p��Q�:�.L�֪���?	������ l�ȟ��IޟH�OpA������,ѢJ�j��ON<�'In7����%���?�8�h&�,5�N$yn�`C��3�I��N�?hl�'}�֝����dy��wa~����Co��!J�@ ̀��'?b�'���O��	��M#`o�S�k �%a�AXa��j*�+-O|�oZJ�g��	�MK�/M�vK6��T��:}#�< �B�I����'.��Y��iK�$�O�-	 ��1���@�<!��8]jV�����;��=@pE����[���	ğ��	�d��ϟ�Oz`%
C��t�<�:�"V�l|J��q�8����O^��O����|�4��w�����:V�\E�6	]�OS&�z"�O�6m<���I�O��6Mb��jP�sG4�"�J�d��#���I?��X#�'N��'P�6M�<a���?q1�����PCP�����K��?1��?������F�J��O�|���|*�I�q���kH-��2dK�C��$��	���o�L�ɞW���Ԧz�\8Zӈ$���I�h�7�Ŋ(.��AB�ULy��~�͐��'�X��I�F7d]1`H�U����T�G�=�e��Ɵ �	���Ic�O�R �OOz$��jS*�3��I�:��Z�Wo�I=�M��wLz���
(a7z�:�E��@J��'T���g���U6�c����q�"x1�O��̉�l�AP���tL�&N9FE�&l
Ny�s�:˓�?��?!���?��?*�6�o�Ā���ܫMr�)Oܙn;�\e��̟<�	w�s��kT���W[�����K��� �������ĝ䦅iٴ���|r�'�?Y _�(��G�;�dܡ��D�+���Ӈ!Q��򤖺_u��k�Fy��X뛖T���r΂;`��t�M0�݉�E[����ܟ��	ϟ�|yb�k��5K���OBl�&i��/�6	�/�9'� 0t6O�Qn�f����I �M���i*��⠴IQ�$���0��,ɶ8�q�im��ݜ�`�����B��e���MA[N�� �s� m��0⡈S)~v�h��4Ox�D�O����O����O�?]�it,��M�	�E�WcT՟����l�ش�Ĉ�*O��l�E�I|��@ o��Y.f���XZ���%��[ٴ@���Om3E�i��)L|��Scg�L �0��7	;\Y��j�0L��i�ЛÂ�'���'@"�'J��'�@e���R�fR�y��#R��S��'�Q��j�4�d����?9������C$�r��#|6݉ jH�W����'���w��v�a�T�O�"^�������T�k��C$
9�U��1�@}h���oyb�w�}��'����y��Y�><4
TD�[D��	�'���'B�'�bc�<����<�'��Zj��Mz<��'�[�7AYʅ�;]^�ʓ;�6�'��'�r�䛶�ͣ��D9��/'N�`�,̯e+�6��O�p��`ӎ�H\L�xd��r,OHx�#�F��Y #�������K�צ	�'�'h��'�2�'	哵u}B��j�.T�P$	���3����4_\����?���:.��A٦��:pz��%o\�;M���7�ˑu$�q����M+�yJ~R�"�M�',h�ٕ�-`��9  ��$#*���'��FPޟ�H"V���4��d�O���ۓ¼�����&�A�h�8���O���O4˓Z��G�����'��$� Y��L�I9���C�]Vk��|Bͽ<����M�I>�7��p&�d��I�����u�x~bMS�B|2����H)R�剷�u�E�ݟ�"�'F�ԁ߳~��HsǗ (`�4�'^"�'4"�'Z�>�]�q�Q�w�5Y ���Ь��5�����M�U�
��$Q����	m�i�iA,�J�2D ��;�4q@�H��tnڐ�M���q��ܴ�y�'q����c��?u˔-W<lN%d�݃x�\q��Ԇ��	6�M�+O2���O6���O���O
�3r�U-��9���L�q��L��B�<��i&����'F2�'���y���;x��s'��g�9g�@�wz*˓�?��4�����'�?���$�"�s���SV(�N=�V4 ��.��Dѻj��;��H���B�vP�3cƠV�j-!��:��b׀���'�R�'k�O��	��M[1�
�?	�F�CX�(ŅVyH0����<ѣ�i�R�|��<����M+�SS܄+�`Ʃ~n�^ x���R	�9�M�'��,B�{������S���1�u'�w�r�8Aj\G��hs���0�
��'�r�'K"�'���'��e���#=<� �g�^�R/D���.�O����O�MoڤJA�-�'�7��O$�*܌�wJ��tOT��ˊU=��aH>	C�ijj6=�@1"��t���*2��D% H�q�k�o�d�{�`��]W*������$¦��'N�'��'̒�Ӑ`@4T���C�m���P"�'6�W�Hr�4K�m��?i����	݈)��黦D	f2kMPX��Ot)�'�p6�̦�'����?�	&�@��)��
� �L�;�NQ� ���R��#a�"��	=2�����q�\�����k�A�A�XiS��E?v�>q *��?a���?���?�|�.O��l��8x��������ѓc,���3?��iI�OLL�'�6m(	�q�4��Q�Lsf_(Z�n�|ʑm�ݦ�̓�?	���!�V���Y~2���rD�۲�M>R�0�d��6m�<����?����?Y���?�+� ѐ�K?/��p@1�fK����/�¦� %�s�L��� &?牍�M�;d��ͨ�IȌb��6k��@��i547�9�4�N���O��@�goӊ�	$��SP�Z�&�(2"�9a*��I������',���'�6��<�'�?�����4��%���B	V��?���?A���d�5j��2?�����:A�x\�8�e�%��Mj��k�>9%�iq6�)�d��6�2�H�U�6��(ՙ=;��O6�r�ƈ@�����,B_wD$�ɞ?rb޹h�t�ȴ@�ԆhcՅǨ2��'B�'`r�ȟ؀��D5x¡��\������ϟ��ݴ&e�5�'Ƥ7�7�i�u�P��^m	��M�eki��㶟�n�M[�GV\�s�4�y��'���t/��?i⠥��2��	��� /T����JRS[�I��M�*O�i�O����O:���O.b��V�G7]R'f�!i��C��<���i��A�'���'���y�K����M߮{6@}ځj��FJ0�M��fgt�F�O�I�����= ����e��#`p�A����8@*E�s��k�I�M%��$�'�0��'z47�<��2&L�\#�K7.xޜ�ũ��?��?��?�'��D�Ѧ���i���`)�&2��d����32�>f��1�4��'���'`�6�|����$	��P⑬�.6@��1`N'NuN�0/f��:�˔�I�4�~"ù���NYIe�	��S%.��yj���OF���Ob�d�O���5���vx(�E�^�~��,�bϛ�#�������I?�MӦ��}~�����Ob�YP�X(MT����B�S����UO'���ŦѪ۴�?Y�n��M[�'�b�"h�d	ԈX%M�4R�nWZX�!��Nԟh��^�<1޴��4�����O��䚂6��h��' l���kQj��kG��$�Ox�YT��J��y��'��X>u ��V2*��}���_�V�E@%?�q}��tӺ�l�p�i>���y�*�ce�� [ K0hW�:�0���o�^Q�E�*?�"���|���T�˓��[�"�9ʂ�I �qeb�*⧟?�?i��?���?�|r.Ot\l�
�;�MO~��A�s��bD�Aqy� lӨ���OdhnZ�5o`�cWl�,FD�O�"�~Y��4P���f6O|�	#\�J�(�"�վw"��$��� �-�cg�^ۜy�gA��hĴit栗'+��'�b�'�R�'h�'@�N�eT�ٵꋄp.x4q�48Yٹ���?������<7��y�
�����D@'v�Za����6�ԦXK<�'�"�' 8zy"ܴ�y�˞(*h$�Ө�r��t�6(ъ�yҢF(:�`e�� k��I�Ms-O����O��2�
�A�ЍA�(�+�K�OR���Od�d�<�d�i��0��'
b�'@BM��`5���.V���2��'!�'y�˓�?�޴r�'�Sǀ�p�^yhw"_+pY<屚'2镍wRܨ5��	W��.�u'gM���p�'��ez��:jn 9*�g�N8��z5�'[�'\r�'��>��2[���,��'�ܭQcȖ�I��	&�M�ܻ��d�ɦM�?ͻ<T�%�,E�4XN����Vg�&`�̛��k��oZ6:�\�lZs~�ݧ'�.q�S�D��G�8W�X�cꍸi�R`DU�jٴ���O���O���O���:�
��	�qNV8���
"�VʓLe�6��L>��'	���'ʄ0��Z)�!B�������<9���Mc��|J~Q��!��A��fR�H���` �
#�(��i��$�ph����~Th˓�vS�����@�8k����_K��Z�kZџ�����������Dy)p��IZ'�O�!	�ϭA�����J�t�U�F;O�n_��8��I�M+ŵi˒6�C�<�����b�ZX�4@V"IPry�akh���ΟJ�Kʸ:����Gby�
q���Q�`�R�V�5Þ�P���!0��I柤�Iȟ(�	۟��I^��XF��IX���`�ƒQ�m����?y�؛���7-���4�MI>�w�>W���S ��!y&�L�zV�'�R6M����� $čl�g~��
#�T� �8����!�Z"�t䪴��֟0�C_����4���Of���O����'0���b��.3h(A�EI�&����O<ʓ=כV
 ����'8�T>��Æ�&�)��Fؼ7֞L!V�:?��]�8�	ݦ�hJ>���?�gQ��xW�]((~�H�"�p��X��^�wKV��'f��]'2ReKyb�w����D�E��@+"��E4n��4�'���'�b�O����Mk�B�)CP6��ߊ$H>��'ϩr�Ҝ",Oj)m�_��"H�I�Ic#�\+*�T�Q� W�����8�M�T�iJkG�i��D�OBUq�"ɫ����<Q��$-	�
�5�<��RE���R����ݟ���ٟT�Iٟ<�O
F��&��N� yȀ��C!6I���cӜ|��9O���O���$Z��]�$�mޓu������UX�41A�FD=��J�"6�w��#$���r�l8����-x����$�|��+g�)K1��	K��hy�O�� H�6�-Q�9�"(��A��?���?Q)O��n���	ʟ(��#?QL���O& <I�F�q�)�?1^� �ݴ\��i;�D� �`���E1�X�:�Fį+�I1$6�q�6��_
�b>���'����<!X��A���f��!b�G�]�����П���H�Ip��y�E,B�Vb�#�H�v���D٧QW��rӐ�p���B�4�?IN>�;|�0H��E	�i��$JS�ۇP���kX�6�r�b�mڜ<ln��<���2ty`��.Hಌ�'M�0m1t�מ��	�BJ��䓙�4����O����O6��, �M�'�yuJ�sE�s��L����2���'�����'1rD�2n�7���z����`	�S����4f�f�7�4�6���:��A�.D�xqA�ƴ�X1t
 b`�����<a`��)3��� �����G��%K����N�A$�
Ae���O`�D�O��4�d˓UM�fŞ,2=2 �Z���ڭ5�&h)��	��yr�q�|�`�O�HlZ2�M��i��|�q� ..�H���χ�4��a,�/R��1O���^" a���^\$����;S]�L(`C抍SU@к3����?���?��?����O1���<*�����L�^�ej7�'��'��6픔T�b�8�֚|ҍ��"��X��Ӑ]Qܸ��OB�q��O"�m��MK�'OZAQ۴�y��'��*b��;q�8�&�c�\�!�6p~>��ɒ&�'x��ɟ���˟���3<�0����( _�؂� 6�����T�'26�(C`���Op��|��H���zh���ukr�kCm�l~�J�<���M��|�'��S���/��i�`Rtڵ:#�ɢ�.ycq'��S	<0q/OB���?���4�D�w�Zr̓1Id=@i��8z����O��D�O���	�<���i V��$A�a�x,��i�1��|�^&^K�ə�Mۏri�>��iB�3 ��+v
�!Ǐ�2/�d�� t�r	mZ#N��Qn��<��rBH]Ac�y�-O��x&��G��i� �U�>y��as4O���?��?���?������O�48���L:�MZ�&���m�h�@1�Iȟx��u�s�������JS�6� v�
�͂Q�������`ӄU$��S�?i���#yv�o�<�I�o�0����4��
�<�VNн2��dL�������OT���ET�xՁ^�<n�@'kގE-&���O��d�O�˓+8�6���B�'��l���'^��=K5�;�Of��'�6-Y¦͛O<�ਘ1gR���񎉄*�4JϤI̓�?��p��2􌙕��u3�iV>�� �1N����A4��`@2���Or���OJ��'ڧ�?I��I�	.��� �R�@���H��?!�iJr�2@Q��H�4���y'狇[3��Ek��t�)�nJ��y2j�� lګ�M�TИ�M��'T�.�(ά���ۀ �ၧm��]� ��ٳ�ᐵ�1�d�<a��?9��?����?Ѳ.�:�xi�BȴR�.��� ���Ħ��@ܟ���̟�$?��4'4P:��:[��A��	�+0�r�P�OT�n��MS5�x�O��D�O�>�J�i�
g�0�r����b�����9���P[�x��"�1i��BQ|��py®]bV0�DlұUN�)��ĝ ���'��'m�OM�I��M���J�?��L�1��Q"TeĢ;k��!҇A�<�i��O���'W�6�Lަ�Q޴<_fAS��f��5��[�5a�	�1HO��M��'2B%̧Z���S���?����4!9�leYU��9������Пt��֟��Y���6�x�mE�8����2F�1K۾�k��?��4]����q�I �MsK>�p�#L�%PrM9Z��"g!Ѱŉ'46M�Ŧu��(2pt�l�<!����1�@���H��b�����\���H$GT�$9����d�OV��Oh��GwB����11�B$�DǞ��L���O�ʓc@�栕;���'-2_>E@g%v����Fό4��(���O�p�'�*6-N��ipO<ͧ�
�А"���&�Gh�k�I���:1`Ơon��*O��C��?	p�"�D��|2�a�@lOd�<J�$4����O��D�O`��<�i����N�ʔ�qW� 
̼�q�'�<!M�I�M{��Π>с�i����Έ�V�B *��"$쬰�ha�Zm0p���l��<���tD(��&��	p+O�ӓ��t�v$�5��+���3O���?Q��?����?����iX�4�DjQ���IJ ��ei��?��Ml�,%h<�I��\�	r�s������37�͝C$���
�B�5���33��v�`Ӌ#��ɞ4u�7q�7nJ�-,p��"F�%��3�
w��b��'Nb�	my��'���
��8:]����7�]�Z������?���?I-O��m�/x%�������bTN�Y��r�N��)L7{���?iA_�$@�42�6#�=BR�@�h�*qRmB`�!n��OI`�~1آ��<i��jXp�D���?�Gd���������4����?���?���?э�	�O&0���^���Q�gS����Kg��O��o�v��d�'�6�8�iޙ�VD[w1���r?�J�n��Rߴ ����|Ӧ��եj�<��.<x�$���hc���"@��1&M� �Byq�O�䓡��O����O�$�O���T�,��ъ�c(�2��0d��uh�	*��G�!�'���$�'_�� �R�7]�Y���H�����<)���M{%�|J~����N��j^�BL�9�l!���p�ʗ:��гU� H��S���O,ʓ#�����j-i%�Ò:h��?����?9��|R,Od�nډa-64��5Nl���� ��@R�D�"��I��MC���>���i�B6���q��8��T:G6h� ��CpmZO~2D�#���ӿ<%�Og��>��� g�Ӷmo*�0���y��'("�'=��'���)�-����p���I� C�3��D�O��$Ԧ��BFvy�v�ΓO�<(�×1���B�*	�MR��:caJC�I��M��i���~���>O��ʃ:tE["��P��L0SQ�yQ䴩B�4�?!�i#���<����?����?�kSS�]��GԊr�\uZ@MT��?Y���D����(�#O�t�I��8�O��@g��$�!�B��]�v���Ov4�'�t7���*K<ͧ���J�4�n��&K>�x�����a�3Ǜ�Tk�ԁ+O>�I��?�Rg'���O0�r&E�&�[� ��5(��$�ON�d�O����<�c�i&�̈�M�2��]�%ON]=�<��"h���MÉ�O�>qҽiV�ܠ�E>N�e��I�&� �9g�m�t�lZ�^BL�oB~"�E4O�Y�S&��ɣa�J`8���~d��1�ȧqTX��Fy"�'�r�'6��'�r\>���eųzD�� I�70�|8�f��M�ń��?���?�I~�?=��w���&��Z�{ .�*��i`�zӚ�nZ-���|B���j�͊��MK�'��97ɖ!Gj�(piڪ=La�'���	rϟ��3�|BV�����ĉ��)aFЉb0�\.&
��*�ɟ �I��\��Zy����d��O��D�O����?ݺ��̈�m�v����;��2��X�����4!��'�����mx�X&��gmP���O� Z��R�.�*��:��^��?����O `!��'���ʓ]���1���Ol�d�O��d�O��}λ��p	�͍)�12�"�S�B)K��k�6
��F��I=�M����Ӽ��/K���afK�kwB����<�q�i��6mݦ���M�����?�F'� O�����e�u����;���p� �|~�-�K>�(O���O����O����O�YZq��y���5EEaX8���<�g�iR�E���'���'���R>�,A���9S%^(w3rP�P)�E�R�O�o=�Mc��x��4��/mdZE�QCZ�2���$+�'U��*��Փ?t剮l�PmK��'Q��$�|�'�t��e'G+\;�eLR-x�|X!��'b��'�����R��bݴSV���A����E/[N( j�\.k�\�"���'��'���ӛf�|��o��{Ϟ�y��^�T��lr ֟SD���HC�����?�qjƾH���������l��?pa�Ɲ?M 9��	BS��$�Ot�d�O����O���5�S�h� 3`��iz{�ƙ=��}�����ɿ�M�6!����ʦ�'�r�׈9X��"��	�is*�z#C� ��0כ�imӚ�)�t�7a��I '�z� 8��TC&��D(���^���aRcG>�?���&��<����?��?q���{��	�&�/2�%zȝ�?!����ėǦC����	ڟ8�O�m"��%'|���A��<���r�O���'װ7m����M<�'��7G\-OgJ����Z�'_0�)�șYs*����/C��u{(Oh�	߇�?���)�䓯K����,<N��D���(k����OF�D�O���i�<q�i+V�z��;��K
: j̘ӳ��>w	�I�M��K�>��i�p���Ö:m܄���D���-X�cg���nZ`�>�lZ�<��:%pҦ��ص�.OJ؆�O��i$S<#<T��0O�ʓ�?����?I���?A����<*��sF�ֻd�D��$p�j4o�=F�K�OB���O���$�Ȧ�]?1�����7C��[�FU�u���	۴����0�4�*���܈Io�,���hL�WA�#$�r�C@��(j=��I�xb�Zr�'��'���'��'���U
��H1�4� G������'�2�'�2Y���ٴYY�PΓ�?!��E�L!��ϳ<���y�Onx y���>���i� 7��o≉;{�٢D��$|�@�D7���蟬@�N�Cn�sè#?a�'Q�$�dP��?�@�&Q����\n9��0s��8�?Y���?���?���9�����R�0T20�qC��R!�\33M�OX�mZ�Ssl��'~�6�4�i��bC~��E1O�;�.Y�r�p��4,&���nӜԺ��~�l�Iğ<���m��B޹N�4m!�fE�o2
l)`�K $��&�x�'�2�'#b�'���'�V s�ҝ>W|��g�ڒ'��Q�]���4w��8͓�?q�����<iDgE�_Cn�	��E o>L �g�H�>v�I �M��i��O1�t�I��
�b^�����4�sDO
<_�1S���8h�pRL�r��Uy�ДR+��C�&�wmɁ�$u���'q��'��O�ɟ�Mk ���<1��")���q���'(��	A�I�<Yſi��O���'�ҳi� 7m�>"�=��T X��Sa��&*�&� ��o�\�I��@��xu��L-?a�'���ݱ_���#�ė�47~�07�S�<���?���?���?����؄v�-�3��>�`@�^��yR�'���v�@�J���L��4��Y'� �oZ�,�*���C��$��e�xb!g�B�n��?��������?�u�F����`�4;&h8*'e�2���p/�OM�K>1(O��O����OV��ۿ-���PC��$�f��G�O>�d�<d�iJB5��O��D�|�h،B�)Ď0�r)j�E@~RI�<���Ms4�|�'�.Ll}:w�
H��r1�_!Șm�FC�'l8,y��i�p~��O�rx�	�a/�'S��(�*�Z��U2�I�A����P�'���'�B���O���M��V7
܈��)TQ��qyC�����a+O�n�Z�W��I �M˳䚡G_8�bCt�a��7J�F�k� ݱ4 l�8�I֟$�b�����my�!�/>z���$����q+C!��y�Q����֟��	ԟ��	韼�O16�;���V.h0�q�
'M�i�t�|`Њ�O��$�Od��������W�����$_.��&��)iv�@X��M�ě|�'����j�Z�xٴ�y�b�(V�Uk c��^������y���(���I�'�IƟ�I�fN��i�薏.�N��a/Q�P��	֟��	˟��'i�7���R&^ʓ�?ѣD��f�j``���E��h0Ц��'��V���x��'�\صfV6�H�jT�B�V���Y�y2�'���0�ܱweddtU����q�@�ş��!�7Tk�!)´q� �#ҏR�?���?Y��?��)�O`�)F��2�U4!ݏ+��9���O�o�=d�$��'@�6�;�i޽���߷dþJ�C�z����"l�|B޴t���~����r�d�t��🬻��M6o*���M�b�9/ٶ�a2ؽ'x�l$�x�'�'�R�'��'*��"���.j�M��
*Z�.�#Q�ly�4Z�0����?q�����<i��ߚ�$���Ǽ�ܠ
����nN���MK�iC4O�i��(�	K0q,eb5M����`9f��V{f��Ґ)�%��$�{V���V���OZ˓)�%��՘-4֭#��P�bx�J���?!��?���|*/O^�o�`�\E���_`�Qf��ԁ`��,)y�I��M�n�<i���M#ӻika�k�t�",P��1\�P[����=��:OH���'��4���N�˓�j��_�����E�}o<1:d���bo�D��?��?���?Y����O�<�@a�P-Qʱc4m	r�4� ��'���'��6I���˓P�&�|��G�?i`�(B�S�}�ëܯa�zO�n�+�M�'0_bQy�4�y��'�~<�3���yAp,�F�D���p�'Xi�����A"�'���ȟ0�IΟ ��,��)��EĂ)�E gN��jy��ǟ$�'�J6�-^�8���O:�d�|B��Á��u�P��1N��0c"Tn~r�<)��MKa�|�'�j @K�	֩�v/ǵk�9��H$-��c�^
/�@L�,O���-�?�1�:��O�=���*���yANH!����O�$�O���<q2�i�[��I:������B4?-ȱ34�4Eo�I��M[��<��4�B��5"��L��&�A�x�A��i�B6͒�[m�6�$?�b��O�������^u�`�4&p�Q0�E�_`�d�<����?���?���?�)��9(���+H�L��6v-捋�̦}BvL�������L'?�ɀ�M�;'�Եт�HO��9���%{��r��i�6Me�)擝Aڜho��<� ��*5`�7M��c���t�4�8O�xk�HJ:�?���$�Ī<9��?Qª� 7p�ke�/��vO�?���?����d�˦�sr�ܟ�	֟ s���x;G�F#+Qqi��Kr���O��l���MKD�x�c�A V�X��Nu|L@RI��y�'_A`��7�	Q�W�d��4��Eϟ�6m�KJ]�ס�UQ���W���	����I۟�G���'Dq��ʬ��jǌ
�a�2�I��'��6͏t�˓y����4��Ha��؜MH)��gQe�&���O�6�R¦Y۴d�r���4�yB�'������?U`¢ޣ;�~aţP�0�t��dAP�vm�'��	۟��ȟ\�I ���LP���t�G�Axʨ�a��ה��'�z7M�$#j ���O^��5�9Op	{b�W�|��̹v%�=�l5$	pyr�''�&�9��O��t�O�l�qSf]=ta��"���$�	��r�ֱcR���V#��U.R�X�y�hF�_�daS4�'���т�H>9���'=r�'F�O�剩�M����?Q��ۘ�:,���S��h�U�<9ָi��On<�'7��ܦ9kߴO��]2�eI%E����R�X|�0I�M]��M��'f�&�J����J���?u�]J�P���j��`;�-C�)��}���	ʟ��	����՟��I_��ܚ�{�n�{�d�1��	TU�}p)O��d�զ��U�#: �i��'�Фs��
���s���!̰���i-����1���|�r���M��O"���D�*C��a�K�Rd��֩_y|�R��Ox��?a��?���DR�}�-L,4�t���*�xlř���?�)ORm�_�����̟��	D���Xb,д1FIDT�Խ"AL�����H}B"v�>o���S����3����g
VZu�`�BOFJ�2��зMZ`���T���A���C�oD�`	$��F��	��N2Q;"!�	ğ0�	۟�)�SHy2.|Ӵ�U⋉���P�M��)��G΂s$��d�O�	m�|�@����M��eǅ�l���'r\���@[�fu�6-���o���ퟠ@A�%#�ĮXxy���H�����}�
Bt����y�\���I��X�	埸�����OÒA�k�:E�V���Cj��9"�~�T�b���O���O��?i������,��E`�u���mт�)0Mϛ�fl�T�$��S�?����E(pn�<Ir�ׅq tCF.]-�f	���<!7 7j���D�0�����O ��u��1�J�;S:��	�+F�V���OX���O��[B�ƫ ���Iß� '� ��y���ƹvŎ ��Z��x��	��M�c�i��OH����$��0�QBZ%ei6���8O@���$����!��������O~$+�o Q�BaD�jH]ef�*!�Xr��?���?a���h�*�d�%���{�K Zn�@ #�~���i'�My2�oӊ��]8X/8�Dc&R"�d��	����8�M{r�i�7m�u��6{����=A������O68��I�*f60��cг� AH�&@Q�IsyB�'���'�B�'�N�-A*��6Cɝ3��s�L�j�� �MC�.ֳ�?q���?�I~Γt���� T<hNP�/$%�4���\����4>�&�=�4���i����S�eP�B"�	i�<���V�]^�>��d��<Qv#�y`�������Ł\�f���FR�}��`��ZS��$�O@�$�OL�4���|�f�9).���*���p�*ަX�
�j�Q/�y"m�^�R�O\l��M�Ŷim�̚B:QyTY��
N 5�1e�|��f>Ob�d�27�x��'{�pʓ�r��Sxx�@`ƾrV����E9%���̓�?i��?��?����OL�9&	H�-&]�U��f(,�S�T� ����M��B��/r�h��<��JN(+��IU�E7}�`�GV=)��'��6��ަ��?���lZ�<a�/�����e�!N���xND&Ѣ�!_8�$ލ�䓚���O����O���@�y2�EX�MM3H>��H����:wd���O����&%	����'y�S>�ka�ٱ1�=3��L��O'?�!V����4i)�6,�4�f��=xW���X�M�/C�^$ʳ"=lU`<ʡ-ѴN��ʓ�����O��H>���W��E ��\+q�,�[�͊��?����?���?�|J-O��mZl*Ip�@Q:o�u���֫kP c�Dy�b�R�� �$�E}Rnl���1��d|��ԇ3d�֡jV���MK�4	����ڴ�yb�'�R�0��?Y��Z�䛒�K'35����,A<���p
p�x�'��'�r�'���'��z��:1�'i��Rq����hQ޴U� 8����?������<a���yG�̲E@�B�>'tfa��%�9~D�6���i�L<�'�J�'tq���4�y".�n���h��^%��|��)�y�.^��i�I�<~�'��ߟ�	J����R�k�(�zQ��#{u�Iǟ�����8�',�6�J���O��䎽" �S�_��Z����5_i��"��u}�xӸ�mZ���(�E��/ϡ$XL��P�N'b�ܕ̓�?��Ł�`�J42�^�����R�waB����$1R�̖($V�z��O�^���D�OR�d�O���'ڧ�?���3(r��@(�A؎0�녶�?�b�i9x�X X�޴���y�(4y��p�aj�~ڒI��d ��y��o� n"�M;��5�M��'&bM��No���3yU<�#/�Vʴ<C$)�8K^8�W�|Y�P�	��,���L�������J@�Q���P+"h���pyRBiӒ����O��D�O:���$��n� I��VT�h�PhI��!�'��6�Ǧ=�J<�'���'12z\� ��G����I&��Y����bʘ���6:41��.�O�
L>�/O�=@aL�4E�VDD�ְBdV8���OJ�D�OB�D�O�<�Կi�F<���'"T�
��ȋB<a��*]=4��ۙ'1�6�&�I���$E���Y�4�?����5�����P #��i�2	ʍTU�T�ܴ���$N6m��'��O�>�،#@�I�g��;v�=�!�
� �H��ԟ��I���Iڟ�	M��
\�����{P��$ڒE�t	����?���Ư6�a��M;M>�����4��&�a��@6���y�Z��(�4tW��Oe�A��i�ɵ�j�b_�*����"�^�(g�,#"`�\�Ily�O-"�'�b����qh�m�@�r<�#��CO��'�剂�M�2���?1��?�)���#&�A�k��K'N�fi~�ps��0�O��lZ��M;`�xʟ�hfhܭH� 81������e%O�j����3N��]|��|j7��O�u�K>��d 5\��D�����Y:����?��?	���?�|�+O��m���:P�.��4��k�4K��+�iycr�����O�l�k�0�:�G�8�d �5/�/$�|���4q囦��.�V3Ol�$U9M<~���'{q��{��u�@�+z�IwJ��.En-����O��d�O����O���|r$b�R��
�뀱iVT��tЁ_�V��9U���rS��y�S �<	�� S�����J{�27��Ǧ��K<�'����-$����4�yb�Hn�����܁T����2��y2��Jx���.)��'~�I�4�I�yva�׎��*�I���rK�M���d�Iޟ�'�7-X"�����O��D	)IL���m[*6|�y���-R]�⟴��O�m�>�M{r�x2�L�nO*�#Q%�e^$!�+�9��$J2Mˤ5 ѠBqlҒ��98��slD�D@�n�;�O9?[�!ʕ��. �0�$�O����OX��*�'�?A!O|*$0�0��R���?A�iV� h!V�`�ߴ���y�"��oLd=�gQ7�F8Q4���~2�'���*d��i�ҍp�6�V!�)�@ �}��K�;[�����
%g�P� '���'���'���'/�'ŘM!Ž1|l��Ǝ1�P�BY�� �4�L�	��?���j+��<]䚙`�f V��ф� O��'�7m�˦�SM<�'�J�'y��K1nԳS\P����y�I��O�B�L-j/O��"���?��4���<0G��/�@T�Ձ��1�����?����?��?ͧ��d��q�(��t���5ڽ�*�#cE�m�C�h��K�4�?yL>9�R�<޴m��%~��!�V�ۖ�D��ЁÏz&��t�i��6�w�H��t�h[@�O:���']���wS��9E�'L낌�@�
J�t�'���'"��'ER�'���:FB�1���d�F��$�3e��O����On�O��'��6��Oʓd�z=���P�n�����5\��xh�x��q�n�o�?��6��㦝��?y�K��@�so�E�>Pz�a����0�g�OԙYN>-O����On�D�OЬ;��ƿMt�6Қ!
"�� ��O�d�<E�i?��e�'o��'��S�(�y�t��c�����D_rd�p��I��M�#�i�,O���R	�?;�܉����f�YP�jȠ�d�*�-��2z˓���+�O�T�O>14�ֹ1^�����3�L���K֤�?���?����?�|j*On5nڶ2X�P���.
=�=D��٨�j�@^@y2Cp�|�d4�d`}2�a�̤� `Qc!2C��!b��{�l������4a:H�*�4�yb�'�,Tj��?usTZ����F�'b�a��U�41@���
t� �'<r�'2�'D��'��S�(z��q�5*��C��!����4)U�x`���?Y����<���yl�_�8GA�:;�8�W���7��A�I<�|Z��@.�M�'����@�/ >�y�A�m��2�'�P!��C؟4�֘|�U�0��쟸#���7,?t5��@V�X�x���@ퟸ��՟���Wy��l�,��2��O��$�O�42����B�CĀ[�F�0�.������զ��4�'����s��
R�Ju{v홮<m��1�'����*gl:m*�mXq��	�?-�t�'h�E�	;Aҥdm�0X%��H��:� ������ܟ`��J�OwaR�'6��Ԡ��l�	p��#;2�d�ʕJ���<	�i:�O�Nդkl��I�J&�p��e� vq�ݦ�ܴ@2��CB$��2O��D��d�x��B�БuUIs�č�(^�Zϟ���OV˓�?����?����?��l��0�mJ�)W��{ŋ�� ��/OĤmڧ	�U�I��<�	V�s��q�Hͮ3�|!�3%	10�P�S"��'��Mܦ�۴uH���T�O����C�5�1���M�����B�lEY�^%J��2,
���'�(u'��'�l=s�lH>�����O����'�"�'����^�8	�4/P����x�����'Z*lCf��w�!���}�����_}��z�F!lZ��M�Md�f��pF�IQn@S������۴�y2�'SJ��4���?���U�T��ߥ��T�&��a��E�;鲐��r���I؟���4��⟘�Zk�3R�Ҽ�'�� �E̚��?���?!�iHXڳ\� ݴ��s,D��
�O
�8��Y���L�|��'���O͂�J��iJ�I8Ubi# "�'E䌱�`,x
� ]�,��X{�I~y��'*�'�ҡ�SՎ��v���wS �£N	�?9r�'g��6�M�ӧΩ�?���?y/�6�h@�{��y6mvK�������*�O��n��M#E�xʟ� Ne:��˱)��]Ȳ� P��JV,T&8/��@U�� ���|Z���O�|�H>�k��3��w(Ld��#�,)�,���O���OL��<��i�fQ��9A����q��0cS�K���*��ɲ�Mˊ��>a�iQ�t��b�8`��-!�*F�+�"���n�Pm��3h�El�D~�"`��1��+��%k�0�1$�Ҏ�t��,H+ ��Zy�'��'Y"�'��R>�{�'�&p��s��,
蒰���?�&�hyb�'��O}�b����F�@�E�dx@�0�Z���Qm�M��x����Ǉ@i��<O����2@F�8�]�2�ꈳP5O>-��ǋ�?�s�&���<����?!@���Z]Z N_%xb�:�Y��?a��?�������p���ޟ��Iğ����Q�|#���J7
"	�#�Q[�yu�I�Mc�i�BO�H���˼B�T���}B������8�4

�w5�Iӂ�C��u9B��ӟ�#Wc[Yx� K ͅ�k��a��F��L������ݟ�G��wk�����[-?�� Ӑ ��6G\�p�'�7�#G���O6io�F�ӼkS��#�������@M,dY4JF�<��i��7-�Ӧe:����-�'��8�R��?�x�m�VZ�֬� ��ԁc�U-T��'��I矜�	�����㟰�ɹ0ˮ1������љ��<&\���'�N6�ɇkG����O��0�9O��� �A+[Y�$��Á/DxՊ��Uk}�Na�\�n-���|j���R"��$/q�-����.d�X�a
wehP�����Y)����wO��O���H`�СEDQ�x� jUo7XlP���?����?1��|Z)O(pn��mj4���.N
�����P-���_2*��7�M���>!ƹiIB6m��5Z7�/L��K!0%�͑6Q�кi��D�O�92�fһ��a*�<9��ǿs����f�L�T���/8t���?����?���?y���O�F=�<$��TC?B?��3t�'!��'L6�^&X�h�j��F�|���fN�!0�1j5�9�b�K�2�O��oZ��M��d6eh�4�yb�'=��bȂ���Qs�j�7_-���2G�,�$H�I3��'����p��˟��	^c�c��8����m�)]4vd�Iܟ��'�7-\�'���O���|�4�����Er%e
�J�}0��WG~��>1��iu�6u�)"�)M/`���3�Ɛ2Nn^u�엩1�z��Ƃ�j9����ǟrԙ|�dX!q�h��N�9V>��ǭ��r�'3b�'����Q����4E*Z)�'+�&AD&�c�+�;n��al�"����y�?�[��*޴1��!YS �s�'��!Ό��is$6���&6�/?�#!\�	����DȊm�8*�\
&�,k����d�<i���?���?���?�.����Rf���-S�4��N��:�E��L��ş(�RG��y7�����x��S/Wh�ي� �*�Dj�Hu&���t:E�z���	c|���(z�F�s��E�&�.�;l� A�'�'�\`'�H�'���'��D1u/�*@��������I��'�B�'�_�:�4R��TZ��?)��q(�(��"b�H�"U�PwXi!���<i���MSВx�Ǹ_��t�CF6�ʅLT����^̓φ(|��f��������'	�qv*��`8:���A����OF�D�O���/ڧ�?����e<hi)��T�u�q8�ˁ�?�'�iMD���^�,��4���yJ��%5Z%z�� c #;�yRG|���n �M��E�M{�O��րE5������P�5��!>᪜ �o��G�|rU���	ȟP��ğ��I��L�QG����0#�ćIq�E��Cy� k�n���N�O�D�Oz���$���څ��L�z�t0 �� +�B��'F�7M¦�L<�|��	� d�=@�o�>��7kG/ T�G�����ެx�0��wKҒO��5�l��Q 2}*AX%l�-������?����?	��|.O�oZ�@,^)�I�Y��xH��/g�4�!7�Q(5�X牸�Mˍ"!�>��i��6m�O��"g�p�N��R.\qJ�胉�g66�>?i�#V&4#��)9�Ӗ�5@Z9 ���`�	Cx��N��y"�'���'���'���	�!�b�����?V�$L`q�t���O�$D˦��b�ryB��F�O��
Ѩ\�pn�Y ���0�`D��{��'T�6����Z��Dl^~MU;F_�Y��o�8�I!��mMt���������|�V��S៤��ʟ�0F��&ٰ�����1&z�	ş`�	Eyc|ӈ��I�O,�d�O�'%If-*���:K���%�-"�i�'f&�2���i��$��'bu��¤� ��q���O-FxJ}Vg.XW� 9�����4�.Q��vt�OD@�d"�n�~��O�o�r�KG��O��$�OR���O1�˓	���i��lt
�h��غy+\h��&�E� �fW�\cٴ��''\�Qg�vML`��KSL�!<���1�O/?w�6�֦��$�����'b� Bc.��?��1Z�d@5'�0��q@j�0|$��zQ�o���'���'?R�'�r�'��;]�p͚$�*��xц��-��t#ܴ�
�H���?������<9���yW�B�<���7�#QQ ���mu$6-M����H<�|2��Ҏ�M��'h�)���'9�J��ǥGP}��'�j�����ٟ$qt�|�]�X��˟	���.1�B�(���R��nٟ�������tyaӜ ��O�O���O��%�\�k�>��� I�@�*�P�h.�I������k�4&���� 6�2�ٵlԸ�p @3	[�����h�	���P�q��V�ӏ�⏌Ɵ��V(Y�q8T���� -�t�	"������	ҟl��ԟ�D���'혅�$�,~���)f%A(�%�OBxo�2)�Q�'�7m$�iޕcEۊ=<b�Y���96���ȧ������Y��4s�ʡq�4������ �'-��X7��\�>�C�M9xu��Q%C(��<��?���?)��?񥡚�	��uAkҽ�%� �P
��$�㦭���Dy��'�x�ӂ
^���)GN߹&.Ѕ*��W}bAm�t�o���Şv�
I��"��Ү9���J�9����+�_/0�Z*O^���_��?	 J!��<�,��ZH$fu�j �7���?)���?����?�'����=ۓ-ȟD��ˋK��Y��݊c`�Bob���4��'6,�5Û��hӪamZ�NF(�c�n?� ��qP
���m�Ϧ!�'ĝ `ɓ�?b@���w� ���.h���'�Y�w��eȟ'�r�'�b�'���'��fmX�g��9�xA��Y'q�8�I�.�O���O�n� ��͖'L$7�?�$�&����TKK�&	���3��j�%����4^x��Ox���E�iM�ɭ;;1�'HғE��%���,~�)�	ъz�"�B��Ky��'���'7b�ȫy���c��*s�B	�͌D�'Y�	8�M�4�<�?���?�.���C���'�8$��́�}�X�[đ��[�OؼoZ��M�%�xʟ���nE�51��(͇��@g@ϬJ��l���3U�R��|z�%�Of-CK>a�lΖS6\����z$�0���?����?����?�|
/Oz�o�33I�13�+FP#VN�S�rs��sy��xӘ�`#�O5l�-ot����œ�1�l�+��@����޴3s��AJ>4�F������S50����{y�Q�ɀ�r�j���yA�,Ұ�y�\�\�I៌����`�	���OZ���CnB�|�3^��U��͂�5��pM�I�|�IW�s������cvl��o��I�A� �l��:věրm�x$�b>�i�C���Γ~���#�?v�>�	 ��`�ϓZ:*�#���OI>	.O��O �PA�֔�v�h�!E3.&���tL�O��$�O���<Qֶi}؄ј'\��'J&I��A�q5P�#g�В����r}�w�*lZ��}�D��7mK;z�Q���(P \�'�`��l�qr@���dNܟ4���'��NO�i��#�
r�`�'�B�'�B�'��>��?���Qq�ͳ�nZ�:�(�	�M��G�b~2�oӖ��ݨr�и�'���&�AW�&��牳�M�V�i�6-�>9��6�%?���@.$Lr��A`� �6��$R�!����-
PL>�.O���O ���O@�d�O����	b ��%�̲8���2��<	�i�,u��'A��'���y�IN�[9��R�f�wy��+�dl��di���|�
�'�b>�z�	X`et4 �]�D �aD�F\����/?�"R<=������䓿�D�� R*�H悆Bj��Д�[R�t��O���O��4��˓V�v���y�EC�r��yђK�;'�b��n�8�y@x�z���O��lZ��M���i�v`�ͷY�� �/N�^�ꍺ"'�9�v���w�J1P������h�I�0 �\���8%��)�&3O����Od���O����O��dI�ZV�9�<��A���.UfDE���#:ҥ�K�Of���O�mZ��tA�'R&6�-�D!%o�a���$.�NxZb钄@��&���4z���O��◺i����O���&[:0�a�	�&E��l��
'~ ��+��d�V�O���?!���?��8<�,��(ɟNN�Q,�$Qs���?�`:L0B�,�
w�(�,O�����瓰j�2A[�CP
�b�T�S$*Y~�t�I��MB�i�RO����@��.�<2YP���Rd9p�kge&�@9�d5Y��˓��դ�Onq�L>!S`�C���B+�#[?��x���S<���i����@ο:��u�vF�%	���+�$����&�Mˍ�F�>i �i�^А	�>?k
�ض��	e�0��eӒ�l�.�x�n��<I��O:���c��D�x)ODi��M������T!ztv5ʠ>O\ʓ��=�,���$�k#LK14:ZI9��K�$���ɀ�qo��ʟ������y�⌓jt�H��*gV�9���ZL�6�ѦM�N<�'�b��E�d��4�yb�Y�8��$rVLR����kRFǸ�y�/�g�"y�	�&.�'���Ky�̌q�,D`ê�#� 4WǕ5�0<���i,l�� [��	�a�:���d�(+b��&��?QFQ����4yQ�fl(�$_�NV�EIu��4^����	;m�$�O�)��e�'D�.���d�<���9��D��?�a@R�6�f=4�\^��d:��Wg�<)� �1)�>ɪ� P\�n�{�-���?1ÿi���b�[��{ش���y���{0��P`O�%P��y�D��yR"c���m��M�4�[�P#;OJ�Ċ6~�^����7���8�%��s/aK5���*�|��!�D�<I����*�,�:�*��(I )6%��	=�M[)G���D�O��?)k!�:���+���'�N�#������O�6m�I�韴����x"� z�%@۰d�@5I$��y8���c�<!�d��6q����䓵��>�H�92�z�AB��a|r�w� �H���O(u�� �Q�`}�Gl�0Zk����;O�IlZm����4�MCտi�>6� B���h2̊b�Xa����
N� ��7�k���		X�Z�"��O�2L�' �t�wrl:��l���cgɏ�&��(�'A�2��/�-+01t*P��Vɇ@�����x�ش2�^ �O�6m#�d� �]�S�*i�Mi.��Ro¹'�Hm���M���q&l��4�y�'��m����"m�����%J�gH �b��:p�5�I/�'v�IE�.�1��NW�]�$S7*C�$}Exr�rӸ�X׬�<1�����T ��M �HY�"��!X"
��ra�������O 6M\D����i�<�V��%�
A<q@�)�6Jx�c5��	7�Q��<���o$���D���U�N����ܸ~�DdsA�r�x���M�˱�p�3�L�g/��Zp:
�C Q�L��4��'#����Vl�/~H��(?v2��J0�:�6M	���
5N���5�'N���I��?�J�Q����F-�~ݐ��Z��srk�̖'=�{��_��ѥ�O��'Ţy��7�G;�p��?���$Be��>@Tc7n�.*DD�b$^	V�@�m(�MK��x���f֑ �6;O�ܒ��K,[��@0��h�4O���K��?)Ӡ7��<����?aB�A�}�z�{�.G-O���C���?����?�����礪���ty��'�(њ��

���� �Q�p����f�Mw}�/j�fo��ē6?Ԍ)_��pq��N�����;?���M�1Dl�(B�X&��"A�mZ�Ll���H�D��7BM�)��DZ,SJ���'0��'���S�$��֕��@	C!^v���П���4<p`�'��6�,�i�)�����RxBu�}�����l�Hj�4/��v�d���a'}�t� 'R���|ם ?M��3�@�5L�����&]j C|�R���͟���Ο��I֟r�ɄS�ܔ��E�u9Ī�hyBai��]��8OJ�D�ON�����Cԍa@�Z.]�����
M9Aθ�'�v7MP���!O<�|*�,;�r�"�Y�"gVA�&y6`���i~B�L�n��IRB�'��	�*�� ����x" ���ϟ#�`t�I���I��\�i>y�'��6m�~1󄌌&�2�B�l
��`8� 'W�H=��U�?�`[�4��尿��4ev"Ń��G4i��2���<�U���M��OxR��ܝ������wt�x�$Nٔo'zd�#�3��1��'�B�'�']�'�(�Lڄb
Ak���m/|�y�1O����OTm���>�:қV�|2d�a�@�ځe�Z6"�� BI�Ht�O$�$i�󩎪7|7>?!��0:c��{�� ,3`$Bk_>d�l��"��O�	�J>�*O���O����O����\h�� ��L�;7��x�n�O��D�<ц�i0@�'W2�'��S�?�RoB!u�:=����$
l�:�����M׷iȄO�SG�h���1�H����1r�Y`0!�j߮�<?�'xԮ�����J�0J@���NF�:"�G"����?����?��S�'��ݦ��$�~�t!�D������Ǐ)fc��A�&�D�A}b�y�Dp�wbFj��)��I*e�ftʢGT�� �4��2�4���@��i�����SԐ�f�9,x���c�6��Yy��'��'A��'
�P>�Cc�CǮL���Z"��ܘ�@�1�M��&��?����?�O~���c��w��:'��/}ء V�T�v�����z�D�nZ���Ş.o���ڴ�y��ƴN�pAH�+U�R���6B���y�	T�Z���mb�'���؟��	�rUĜR���"-�V���}\v�����,��럐�'�(6m¶^�Z�$�O���R>M؜���(T|~��P�ԥ�:�X��OܼmZ��M�A�x"�="d#j��i��d �hU?����:u�P�d��*rΤ��h	���~�&�-5����R"&5"F�J"*"���O��$�O��D3ڧ�?qc�>-`H|z�o	�[���;0m�
�?	�i7 4�A[�x�ܴ���y�n	4}�Ҽ#�+��X�\2�d@��yҥm�xtl�M�����M��O� yt�ʁ�J��֣0c��X��B�tX|�� :n��O\ʓ�?q��?a��?��I4i!3,E�^R���C��[@�-O�lڦh4&x�	�	n�s��s��>3֐j���?j6��v	����X���47Љ��OCF�"g�8,���;e��!g�DPs N�w�&���_����`:12�Co�IFybh�ZA\�ۥ	D=%p*h������'�B�''�O�I��M{�<�A`Ժʌ�Z�N�C�82�i��<a��iI�Ox(�'��6͈��(�4-���81M �	�%��ܤm�DZ�, �M��Ol����/�j����w�-���3��C+���a��<	��?Y���?i��?���� T	\:b�M�KW�	��X��y��'�"Fz�Bl�!�����4��1HZ4�$&3\3��s�#_�� I��x� g�<�oz>%���զ��'e��a���'�l�,� df�%���eRX�	�`��'T�)�s�H��J�(�xq򰢁2?���� �!�j%�&�X+W�񟀗OP�������T�br Y o����L}Kx� po���S���^�"$2`H �[��d
DgS�&=�=8am߄i���[��3|�b^|�䈸�������P��8B�ɕ�M��f��3� �*Cj�|�0Y���U7_�f)+O`o�v�z���'�M� ����	F���]�pb��U�Ϧu�ݴu����4��$�DF(�+�'rbDʓOb�0�I�0�0T�v,ڑ�z�Γ���OV���O���O���|�Q�=f�^h�ɍ����7�B�:��D�O���&�9O>�nz��3��?B��RqטrH4������?	�4�yb^����PXŁ���	�_y6ċ�k��^4p}����d���I�hq����'1*,$�������'Q�ES�%�`�R��$�:60����'L�'U�V��9�4������?)��8�Q�G�>&�P��1Hi=�%/�I����O`7�s�8�'�����k���r@G�*�q�O�ӵ��3��TТ�Ɏ2�?���On8����|���E%�M��� �O����O����Oޢ}��j��I��f��T	f�M�z~l���GP�6E *��		�MK��w)�ht,����8R
������'�J6��Ԧ����t� hoZr~�
�� ��ӃF��1 ��3{����8z��+��|T���P�I՟P�	����g.	�EID��7����U��ny�{� �'�Ot��O�����F
h���"G�E� ��ȉ�<Ҏ��'�7���!��H����P�?��U�5�6���Ǉ�%u��仢��
ǣ�-v��-d@ԣ�N����[�GQ"t×(څO|A+�V-趥�����[�"�$Q�a!�Ӆ`Gr�Y�JۥCG*!�Q/>���5���C�l�4%�9(�r-�2��h�cj���T�T&f�B�ѓ+K 2�.��m��I�@qRf/8��0P��h�Ը;$� k�z���Iң֢��e��Ԑ[�U�|�m*!��7$AnA� �c<��jtL߹,�r��Qc��'h$p���X�H�ܑ1F̔�2&΁�ƈ�,�R���`u�d9�#c�c�@�ҡ��/^��D�خD赎�6"����q�6�G�\"E�(v����5��^}��'v�|��'w�J^�$��!Q�Z1��S�h@L��%ài�6M�O��d�O6��O��`kC�O�������c� ./�̩�3� �0L5�'	k����>�d�O��H�RV���x ��]�Ȼɉ����%��MK���?9���?y��	$�?���?�����ͷDrr�!vl�#0�R疭6�'G��'���8f����������c��)G��8W��Сp�Z�X��f�'�c��:*��'��I�?������0��y����eR��4�67��O��D�[i���f��I͖+8@�f�<|�����8z����N�cr�'�	�?���џh�'p�Y�b6�u����e�,Tk�{�ˆ�B�n��y����O�=��T	�Ԙ���A�r2��J!�˦e��[y�_�)���Zy��'��D�U����SHD�}:�5ae�ͼb�*��<y��?��'�?���?QE,�Oꂝ���@+�ԋ�2;���'?$a�R��q����'�ē�?�I��+k�@�f-E:t1�'��.�^�H�O����O2��<ɦ"�\�H��B��FpR�*c��$ ؉�cX� �'�2�|B�'���ݪ,Y@ Vh��֠0ǁ�&�|��':��'��	~���K�O .U·�4jT��Hrb��b�x��4���O��O����Oz�9#����p��+$U4�ЄR�2�j�B�>)���?����^J]�O$�	�-BY1`K�>���� c�ws�6��O�O����O���>�I�@��ȡ՟$�
1-�@� 7��Oz�d�<)��ZT�����H�I�?��v�l���J�/�ưH׋߱�ē�?i���N���Bܟ�8�G��0���U� �2��i���
t
�L�޴�?���?��m��i���w�C(Ɉ�+G2h���J�z�,�D�ORd�,5�	nܧ X�@�$�9#`�hƠC0Tۮ oZfd\Zٴ�?���?���/(�	Gy6GJZ`��?VQtu�Ҧ+�T7M�e��$>�$)���h���e��lTB£cR8A��ʝ�M����?q�<��]��[�h�'���O�R�ς�m$��qC��saf�`��i��'K(b@L/���O����OV���Rg���b��B76�4u�$�TצE�ɸ�|q�OF��?�O>��+�R�cm(=���l�&Z���':`����'��IƟ0�	� �'�H���9 ����0��,x��Jq�ī�x�����Ob�O����O�p)UFͮR^e[F�"C�%��΃=_ВO��d�O��$�<�'�N�I�bڭ`�(ÖYtA�E�x��\���Ig�Iӟ��I1����4LX{����� �C���r��O����O0��<Aɏv��\{sdX�m��ܸ��Ǣ8m�Y��-ǂ�MC����?I�}A�Xq�{r [��"|�ũ����"�� �M���?y+O��R���K����s���M�xjq��a޲E��qÊ=��<���L��?1I~z�O�z��bE��*��D�p�L��޴���6;*�oڐ��i�O��x~��5��}pS��.%�v�����M�)O��`Ť�Oܠ&>�&?7�[1. ��8Ō�%y@�x[i�<nZ76zx޴�?q���?���v̉���@�}\� A!OZM��q)G�t 7�ҷd`��$�O,˓���<	��$S�1H���N��J$ȒD@2����i`��'���q�PO�	�O~�ɕ���Di���H��։cF���4�?I*O��p�J�}��'5�'!`�����#ϩX��x��^�v��7��OJ\P�L\�i>��IY�i݉ rG�h�r���Eʎ5���9�#�>3@��?M>i���$�O�i����2�i�e5�t�dj�-1�ʓ�?����'^��'e:5��N6Hdx0���Y;V�i4�GHf�x�y��'H�IʟLHƃ�X� �8�&Υ*5������hйi=r�'�O����O���CF�;ϛ�
�5	�N���������?.O.�D�^�r�'�?	X�ډjɂ$�����)R���nk��?i�d�:T���q�I�w��ժW�	�Vy�h��ұ��6�O*��?�E���i�OZ�D��klC�=K&8�%��wcN��aJ:7�'�R[���.6�Ӻ3'`�p1���� wx)�L}��'�I���'��'���O��i��Aw/���uy�7�0d~���D�<� Jz���'L ��a�Yj�|� c�	HL$�mڹ���	�	�<�S}yʟ��iqD[ 0�Ƭ�CΗ�H����\}J��O1�h�dP (�:	zr��=�T��b	��l�꟔��ӟLQ�dٛ���|���~�F��2��A�`M�>=�6�j���.�M[����$�S6(���y��'Y��'�ʄ��+0 IX#/�:+�4pf�vӰ���?j4h$��ڟd$��݈Z`|��	�x�lq��F�x�F����$�O����O��e�()wJ�X��	�O��&� �ےk����'L��'�'M�	)*��5s�@�	b-��P�B�XJ��d�Z��0�'"�'��P�0�������d�ƕCa.�#��,;� ���
�byr�'���|b_��2����9�%���lyF	<7ص*T�����$�OV�d�O>ʓ�,�Ж�A�5�Ι�$H�Ex���P�L�u�$6m�O�O ˓RV�в���(h�d*P���#@n��sǉ`$6��O��$�<���L@I�Ou"��5F-����0{g�۹d�&�QHR����O�˓}`��B����'���욿g���mݕ/:b�AGU�����O��HC�O.���O���⟶�Ӻ3u$�Y��&�=J�P\�)G���'Y��-u��y��Gӊ	�u�4�W?v^��;PL��Mg[!�?���?����
/O���	O�D�"�%bk�E(p�S3ga,|�ݴZyܝA���N�S�OW_��xJ���$uԅ��I�:|T7��Ob���O�����<�O��p�&!B4��+܈����f#(`���Hg'֝&>�	؟���$DLڸ�ЍC�N���#�#:���ܴ�?y���	dщ����'��QZA�O i����p�0Y��$�eL�j}b�]#QRT�������	Qyb��!z2$PE�V��B�ÀS�nY"I#�$�O��$2��<���9� 03�FΗHF`��B]�B��?Y)O����O�D�<i��+��	A�AF��C�H0 ��@�J֩*��I� ��J�	by"�hy��H`�Z�I#���)�����N8듅?����?q(O�ѹ#e��d�'�Z( �Ŗ�g�"�����cV�hV�e�p�Ĺ<���?���~�d\ϓ�?1�'���c�l��Lg�*:�XU�ߴ�?����֔i�^U�OZ��'�t�R�a� ��I4���Ef�����?y���yҊ�m��^��'"N�T�C��q�ܸ4
Ncu��l�_y��3Q�d6��O����O���DL}Zw�[!�� ���H�&(i�ش�?i�dK~H͓�?.OB�>ʂ���)����HB�M�Ԩ` a��08$e��������I�?�ʯO|�P�^���GĎ\�|0d �B�y9P�i�
�a�'��'��z����dQ���S�Ūbi���֊#���o����I�ԫ6D�����<����~BL�~<`����T:n���g_1�M���?���x�~5�S��'�r�'}�E�3�?�>��!�� �H��j��dS70���'����$�'�Zc�,1�O	�_�2]�b�[PK<t��O�`�e;O����O����OH�$�<��·RY2���g�,B�a�o�IF�x�U�D�'��T�@�I�����-4Ad8H�b��t�9�<�I�4�Iܟ��'|J��u�x>qh@a#p)�NT.���.v�8ʓ�?�)O:��O���U���
jx���(͘}�r����;rՔ��'���'f�\�PX&J^���i�Oz��6�H�p�<4#�Dj;����䦑�ICy"�'1R�'�^���'��7��4��N֏N�t}����F9D�m؟t��ny2D�D���?y���2�H,%�޴u'�-XUNGJ�"lu��������8§�q����ly�ݟ8!"�
�9���#��� q��2��i��	F�y�۴�?q��?!�'3q�i��#k߬� @掍	���ȓg�b���O���t3O��d�<9��$�W"���#�ɑ7�L	��k�MCCj5���'���'�����>.Ob1x��/
HUaQ���h�������R)h����џ,��B�'�?B� �Fn�֮X�i�&a���}I���'�"�'y��(5@�>�.O0����[E�Y3C�e ��
4��]�!�fӘ�D�OL�D��OM�?���ΟT�I1g�&��#�*��ϒ0P2��ش�?��.�A��Ly��'���̟�(3G(�a�ǚ����@�]�uD�`cb���?1��?I��?	*O>�b�OѵBע�bkROx�PrX��!��>�,OB�$�<���?����|Xg��%��`Ȱ �P�a�# V�<i*O0��O����<�C!ZL�i�| 섹��W�f���wJ�W�_����|y�'v��';��!�O���V%BXTE _�(�b����M���?��?�*O�����\����5��
�H`,����/�ހ�sBO��M����$�O���Of����?�q`d��j�w���`!]z�m�ş���Ay��Z8�4�'�?A���� ��k�(�-����4��28^8V�h�	䟐�	[��T���'���
�G�-KSe�&	�,܀w$Ρ`���X� �#�F�M����?A��JvT��ݪn�B�# '�}�\)�AH�d7��O���M�\��,�$7�Ӑ[t���d�*��DlF�7T7����.�nП0�	ğ��ӛ����<a��>C�� Y�%�4����h�t@�6$0�y��'@�Ia���?ae˄N�>�"�H�C��������P5�&�'Lb�'m�y1�Ŧ>!*O�D����GL�+=��Y�D
�n� �Bp�>�/O&�2����ݟ��	���]20�e1�N�#��L� l��MC��p�l�YUT���'��[���i�u��AU�RPBa����#k&�x�&�>���M�<q���?���?Y����d� zS"�q(�<U��Uȓ�ԫ>��dj%%�[}B^����^yR�'�"�'�q�� uZ0�X�gA�b7|]�E���y"U���	��TybĂ�Y��,P��5��(G��Έ�l� CE7M�<!���d�O���O<�(�:OL����:�����R�
1���Uܦ��Iܟ�������'���Q�G�~2��C�*�/XtUUC�'oI\ɱ�զ��Ijy��'���'Q�:�'�s�#��R|�T��)��O�&�i�B�'��M�α鮟6���O6���70��a�
eq�lҁ�Y,j̕�'Z��'�B�� ���<)�OҠ��� �i�m�3��&{
�*ش���BK���o������O|���}~`M�~˘�9se��4sJ�S���/�Mc���?�����<�M>َ��ۿQ��!���,7e�!� -��M����.��6�'���'��T�>�ɾQ�4�#@%�ts2���HRC��ٴ��͓����O�⌀�_k��wA�i�'�?L�l6��O,��O�R��BM��?1�'���$�)fB��LӄD�F�Aٴ��M��M�S���'���'�>!R��EN��店$:PI�ԙ��d�����<v�b)�>a�������7X�����>'��i9b�C}2͇�A�_��I���y¨��
��U�S��\p���Z��EQ�0�D�O���*�d�O���Q�/�ҁ:�EO
)��@�B�M�WpSU�O�ʓ�?����?�+OH�����|:OP!�&r�"��	� ����l�	��$�H�I���y��f�*cŚ���9�%�� ��b#b���$�O<���O�ʓ[�l x&�������y��E��~H�%,�
)��7��O��O>���O�uJ�c�O��'v$�$�5=v�1Q�&E��=�4�?9����$��4&>q�I�?��MܵZ ��(]tڸ������?!��&Ix�����䓂����
9N�X�E�G-s(�`��!ǻ�MS)O��	���Ŧ9���.�d���Q�'�� W GhBGÑ�1�}�ڴ�?��*h�����OH��"� Q�/���
�?)����42n�$��i�r�'0B�O�b��"��I%L�<4��G�&�EQa�-�M�%��?�L>����'�0�R���
u� ��h� Q<V�r�Is�����O��S�}/�d&� �I�����]՜�Q!�>tv�Ab��2aB&@ns�	;/����sy��'���5�Ԉs)3�Ё/*�l+�ğ��M;�r/�Ǖx"�'��|Zc,����.t^�1ՠ�7R�h=�O�E�3��O���?���?�.OR��ǂIx� ��H�$�`����6Z-H��>)���䓘?!�� �ڨ��d��S3�-b¢�eҵ�.�<-O|��OP�$�<��L$��3,��J��/'ԍ�uF��r1�	��xD{��'��@{�''X�"d@�W� ×�O��1�cӆ���O���O`ʓ5�6勵��d�)J��0 �ص�<$���1M�6M7ړ�?᧡L��?Q���~ªJ(vH1���(<��lʠ�M����?	+OLh�G%IB�ß��s���# 1N�
#���$�1׌=�I��l���Rǟd��ly��np�u�2<&X�S�L(�|pz��i���'����'��'z��O2��5&I߇[�Υ�@(�:d��H[��
��M���?A&�F�Ԏ��<�~Rg"O�8����Q��UD:���W�����X��M���?����J@�x�OG2096GJ�t�b�{�c�v�Dx�t&x�Jh��	>�	�?c����)�J����� '�Y#�ʰ8%z��ݴ�?	���?Y�#�?!����I�O��ɦJ��`�fʆp���G��*?ԐQ�yB'<;�*�`��O��D�`t�IA���RAP�ǅ�La�en��T�V���'t2�|Zc
��K�'�f\�Q�G�g,.�A�O.l���d�O����O"�S`�q�!M	y��m@�JTVn�� ��ē�?����?�dpaKe8_�,D�D���>�`��q��?q��?���?�o����œ �p�pg�*'ZL$�L��M[*O��d(�$�O���	U,��i����W�ˊ�����+�$�8�ЯO(���O���<�2��4�Op��E�5JH�1�@�����c!�}�H�d�O⟘�g�2�ӄ�liH���A�JT�F��(>	�7��O����O*���/˧���&��#��!0�0�BwNKZ�bQ��U��柰��t����i �~BAD�k3P�A��:����@Ц�'`*DZ�i�꧔?��i<���#ў ���ą���n�:7�O\�Ĕ�"9� �}bq��"��]	"d9'�R�Z�����c�զ)�	ʟ�	�?�J<1��r�� >���c[-0)C0 + �A��iv����ğL��D�='��r�}@�p�F���M����?q�~�,S����Or�	(O��gi�n	�!���H�b��5�9�Iҟl���d#���UzL$`��0jת8{��7�M���B�Q�q�x��'H��|Zc�z��q� ���Cq��>�A��O
����O2���OJʓ<�Љ��d��4MfͲC�įNc�`$�FN��_y��'���ߟp�	��;�I��� )��焗 -�QPEBo�@���|�I��	���'�hU�P�{>)Q�3t0�e� H&�t��+z��˓�?�)O��D�O|�DH@���I)K45y��A#��[f/U{}r�'�2�'��I?@lfȪ�F�K�%ij���Y�w|�ٳi�	^٨�m��l�'�R�'��K��yr�>y���80�vi+rj�y���T��ܦ������'�7�x��'L��Of��Sp(	�Nࠤ?e�:,����>1���?A��`��	̓�?I*O6�/���i�䍪sF�1��ÖaѾ7;<���%�V�'���'�4�>�;-�ʼ�e�ȁIӾY�#�V>Zt�1oٟ��,/�#<��d���}��Ayr*�7fJ*��U.�M�5�]�RL�V�'���'���>1,O��K�G%��uQ��A�>Y
o����St�4�'3��)�OLP2!�Z�� ��i���[ڦq���X��0���P�O˓�?��'e��Z��A��Mq!A�!?@<�2ڴ�?�*O<p�4O�ǟ,�	y���$�>�����1N��s�R�e�ɻoKPq�'�"�'�?yH>���I?H��nA(w��+3����I�fUbc�h�����	ٟ���9Q&���#
~�V` @���A�Ly2�'S��'#�'R��'G6p���w�ҼBBC�/"`�P!gJ�N�\��O<���O����<c��
MP���6 Yĭ��-�:ot|�!��&L=�f�'���'��D].<��ɭ,c�
�a�'���@�Q���?y��?���?�fFH��?a���?�
0�8� �02���i���C���'�'�P�lr"A1�$W.#�Xȣ����$ш��!��k��~"�ֽ)����%�4
�ƫ�y2�%@\&��m�{���! �X5tp�M2�e��M���w�KQV�G�#MG�{�l�j��Q�R?`X��r���DMle�k׭wdD�{�(�LvB|��CY9D̞���Q�z�i$�� p%���mܻ[<��t- �X^ܠF�[�5x�%��W�`7@�s~�`�aA#>�ʑC��Cư,�aӪ]6�$�OJ��Ov��;;6�0�؛67 �1S�̘	�Ę��fW�10R @�
�\������Oe�'Ő�ҶL�x76�+2�I;��Ҧ�U I��\ɔ�:`֠S�]�I�x=��+�|�E�%K���݉W���2⦋�W���G/!�U�Ie~b�^>�?�'�hOYPv��:)���s�㗶U��p�"Ob��V?M�(I+�!����|�����i���?�'�\5'��xה�W�C/-؜�f$��S�
��w�'�r�'Vr'p�Y�	㟜ͧi����N�~�#���~����`D���\8�V�R����ϓ&�l����ڇ'�`٪��$utt�# m���I��4
B��;
ϓn��(�����8���?�(țt(������o�'��Ol髧K� n�6YYg�
^QQ@"Oq�����Ii& Q�1˂��M}BY���������O��cegK�?D�fN�l	�7��O��D !��D�O��S֬Sb�|K�j��5�
T�OgF�8&'N�����b,6O�!���(V��u,�*l#����#>.i��C߳.��i7��>�p<���Ɵ�Ity�Yr�j�!��*�4ੵ*B#Ϙ'��{���O� �	mj�\9j	�xb	r��Px�Bǻl���嬂��xtC$8OD�B>��ڴ�?y����݌?�����gW���V��L�+�)��P&��Or��P/B�l�v@�7�~�[>��OG�l*׋^�+�:���;2�O�P����S[����L�~ŞU��ڼS�ҹa��?�ɱ'�.(�tj�퐈aN�A	(}��ۡ�?y��i�\6��O(�?90%�
&}Yd,a�T82h���p�H�'B�^��g�S���Th�OvP�鐄Z�;""��<Ɉy2�iv�6M�OV�lZ�4R��@ ѩ��ª3yD1AaT��M����?���cF6�FC��?����?���ҿ!�B!]L����V�x����N
'Dh ۶縟��׍� v�$?c�Z'׆z4����K@/�y�GչD�m�T\�s���s�̒Q[��>5 a�<ɖ��x��#ՌX�_dT��$�^��?��i�r��*���,O����5V�\iBA$	8W��i�.Z�����>y@�D9��ɒ5G\m`��c��B��q�X�m�]��h�DP� ȲB�0G��G�� )���� D��Ћ��u����f(�ZMD�>D��2tdѦd/�=k���%8V�"�7D�,�v�A1��t
&��2M|���:D�(q� K	i(���JJE�AKk9D��;EJ��N�$ܩ&����Y�c�6D�� $�WB����#��<�D���"O�i�M�
�!�`ԌE�~��"O$˃��L�ddO�mrx$"O��.CҶ��Ʈ* �����"O�1s  �&����N˨<˄��E"O�XQЌ�^)ld��k
;Pj2-;1"O䍨C��BI9��U�-N�T�D"O& "��_�9r�"�'"I�}*�"O��щϺCd
1��=v+�ѡ�"O �J�m�#Z�|���	]�vA��"O$��H�<P�P���nH>�X��"O�J���T�f�
Q�e����"OH�!b��kj�lZ�
���@r"O�-�q`�3�L�
��a�h�i�"O����]c�>�; �T�X~z%+�"O
I�G@���@��@�s�%��"OF]�0��=�(���A�"`[d1�"O�Z�GL�?�(��`�:n^2P�"OP�p�̓.hNt)���
��ґ�"O�ْ�5�u�MP���"�"O<(J&)�6N��Y�V��yS�"O|m(�"�'o�*�Ɔ���"O|EC���+�f5�Re&k�}CA"O<�i�>/Vt!�qi҈N�^�y"OR�Qd.��Hb��kt�<�dղ�"O.C�I�\���:���,�<9kS"O�4Y!G�.y%�Ī���-sBdؤ"O\�p�ۂ/�Q@�n�3Wp|�A"O�)��#r��! �ѫ"�f4� "O�=�R"�w����KƝl�\��"OP��Nٛdv`��Ȣ��#�"O��7��פ���F&$�J(kA"O�����#&��A�"�����c"O�A@��r��B���̌�R�"O�Y�%�5R2��넏C�<��"O�0a�_9G����G�#|<��\��s�j2�S�OU��+���H0̴��Ȑ�zR,���'�D ���F�/:�W*(-]>�I>Q�**�0=�գ%���kC�V8;�A�!��M����U��Un���ŉ�
TȽ�����n8��&u�u���Ca� ��v���u�ER��i>s�'�>׶<�p���y�6��� 9D���v�C�g���O�A�>!����<�Go>���(�xIT(�<W�
Y�R���y�$"O j�jӷ?B�R��E)r�n��2�|B�D+v�az���/W4j�S'�V�lh7�{����9�n�bc*�0���\�j�L�A�<Q�"5X���#��.Q�	Y7���'�pub6�S,u$.=���޴%�hI�N3�C�ɱ��@*�Fɠ"4<	�A̘
v<�!�����i=Q�p��F�K�%n�0�7f��x�!���pf�Q+I�,�f ��PXq�'�v � �'S�Y��(�x��&į�~I��'[�0����`y��,�.i�b@�ˎ�y2�"L�ű�l�rvl\�F�G�y����2^������,� f ��y�,[�x��q䝰ZL������y��t�~����C!? �A@Ȓ�y�H�(�B�k���\r�g�H��y�e�$N��	4��� ��H���y"Y�D�y�%Q
hݢ��Ѕ[!�y�+E�<l*=c�e|��A��R�y&/wU�t�AÝV}��'�R!��'�txjL<��T0�.�fY�W�O+.7��{WJ 	����S"O� ��qG�*$:E��i��\�tԁ1@���!�0���(���)^�6�yr�Z H�����h�DB䉱T�<,��F2V�0�O�}85�'d�'+����!���R7C�&X��Ub�4=<��C�;|Ofh�C�>եJ��M����UZ| u-PU�$�1��a}R�J'<'b!��i��\�j$a#���')|��L<e&������� �|ՠ)�J(Y	`"O�̱����u^|��.��R��Eo���' ��P3��H���]5��u@ӂ��c���hQ-\�"��C�I]6�iE�<F;��h���$�打R<������6ZX����Z�'񾠻冈�i}!�$O#R)� �@�7��-B��$~X!��[=��t;�V�yL�(�A*�!�$�(K}:="�%N@f	�e�N[�!��$s\�}������|℅�/�!�$ܽP�\s�JE��U����T�!�D���t�6��%�s���X�!򄊫U� ��V��c0J!�D -i�to��V��a�O�<<!�dO�e�5k�i��,��l'��6!�ϗD�:ibpE.2�<5!�e�72#!�P�;�`���20�B1�J����y��P 1O�a����RJF;E��)��"O ����k�x`�IO���z��>� ���X��x��$��y����ӳDLd����yr���qB��Q#��G�NP���0gxQY�<�r�����'?� c�Ο#�Z "��|�J]Q�� �O�!`���Z��A�Մ;�l�%"�:��3̓- �Lڵ�'и"A�=�aې�/9�"�{��� i�n�s�öd��bE��|:P�B�B����59�Փ��x�<�{/�Q+��7�����uyB�X&\��Q��3��B̮~���`��3"��(�.!W�&��UmN��!�D�k�3���(	���u�(K ���V#L<�n��~z^�Z�e;��ON�c�O֨)���1D�z�x�oז^D$�QOV�*�̇%-(�:�h��`rJ�e��V �Ԏ��J6�	 �D�y���8ŨO�)xH�7kIzQh��Pb1h�;��'�<XT�[�XE"�G��M���P�X<BH�'R�<�x�Sᗴ�?�E#�B��l�V_8�2KY�_a��b�o)?�Ei��twRɢ��ǢM
��F��}�f	Kq+-�d�J>i�dI �LG�HxZ`*H�y¤@(ּ̉���?��1Ҥ�̚z����g�Ӭ����7�-�N���4�iR���'<�!��,��X��T2[LD����u<� �[\p�A*�P+���`�X2	VRL��	ߎxd����W�K�$�d�i~(�����G�	����
`NI�S��X�ax�C�035 qCuF��n>���+��,��K��ِJ�yA�fޤt{��;u�/$�Ař?4RjdA�@J�����-4?Ʉ@��j��p �)B� �(9�NZ���O��9��b�m.���c 6e܄8�'Wf<�� m��prF�"G��(ui�YH��	��)Yb�P#req��'R��Xr�M�[8t�P��9��- M�'C��i�a*��~�d��r^:EI��s#L ��,�G^�J`�P�,ыz��zҮ��T�!tK�����΢���/9`2p8�{�.TѨ=(�ȭ�����ݶOR�tK���-�@�b⃏,�!�$�wo&�+�
u�jЩu��%��'�z����ERs�n��~҃O�_50�z���Qn9��p�4�F���5��I�~� ��3��,���ELi7��	���Z�A��J�/.���I�9~@"|
����?�Al�9n*�!�W&Q�7��C��Q�c1�4��"'NV�_�J�b�F��)ݸ1 �cG;"d��A��f���	:�ʐD{kH�>>A�w9����*�0=������A��Ò��m��[����R��cL�sì�<X_�����i��8��ɴ+/�M���R�2b Y�*\=8�O X�"Lx�M��jj��r�E9q����o��ih-�@m;�8y�  ��{�!�D��τkEx-�6���d��\Q�K߂Δ<+�x,�2���$�|K4?�OҮ�˙w���(��&F0��E��D��	�'���Tݒ(�@��&�ݤ8WTH�0�dB�k��x�D��h�E��Tm�'�T\�,]0F����a$9o�p��ۓ<��� �% �|��2� ��a�l�'u̦�bT _'<��!P)�;&IFxP�d�
��t�ī�{X���'�N�vr̈s%��'D�So/��)rT�ٗ�4z���3'ƅ�s�FO\��C��� Mc�eg�V�؇�`H<QSF�??�@�`$��-R�`1U��=u�����+��P�&�6UޓO駻y���.�Vز�oA�7�&��怽�y�o��
N��`��[�	Z��F[|&)%���NK6���L�*v���ɕ�5��d=��p�)n��D��F�|-���,�1 �cA#|IzY�4��+[D����Ȍy��3E����
��AO XH�͚HM_x��s��dY8���8�l���H8Y��#�'k#K��1�
��<���}�T\�/�,K�u��"@>g%F�a�'c�hǈ�jxB��`��c0�*1��6h��/�J�> ;kـR��)���E�#нp�8W�>�l�r1"O4=Jd��=�҅�wa�RuBUFÃt�&�KK�tj������i�4a��t�תX�L����ҏҧ-N�tf0�O�u� ܀NpZ�i]N��[��?<��{� M�t�@cˑE����	(\O��ʲ�J"Z��������1@�� L@d�T-X�L@Z.r��M<h|B�BF�#"��a #A��N]�ȓ4���b�J�W�����؜h|J���lF��{�b�!k��̋¯ľtv����94�-�"��$2햰#A�e��?�"��#8`�?mB��YP��2��0'������͔%^хE�
S)�q�9���'!#�O�� �
7�4�j����
�^��1�A���b��E��̬}��|��H�����0��	������9�x��X�0: )lOD
�KT�ì�w�T�J� �sp�'�TU���+�DD�1TT���[>Xe�D�9?T%��)+�Q�A)�Zg�;P�[1jU�@��I��5�.OD�8���h�P��խL�_UܽCcP�@��͎.�J��b�*V<;��'ҧs��#�H�	!�5�U���*4�?�pV�b�?�.%��0Z��X�4:y{"�ڟ	�~VG��,S:]
�<�U�ߤ��g�*�2x�d��:*���I^�d����+����'��>���#�7��H�ܮu�ޠ��C]u1�l�t���G��'�(7a{�*��}�19g�ؗW�쌳��D��y�i�w��#<!��O�/��Y�!�t�L�m�{���ST�
s�8�jSM�PټB�	�?���,��C64�:s�jM����׭<w��qf�S�|4L{�c]�b"��:��\T,C�	�i��@ ����6͘�bZ���6^f0��CFY�)��<c	]�Br�	�B�����U Y�<�v��-�!1r�L�<Szeʀ	]V�<I4�p��@�A�U3Ut�D��J�<!���  ���!Z.��|�T��A�<9�kA9g�J�s��(2@=ʣ��z�<)��?a�pX9 ��*U��!B[�<�v�A�<8��ZSG�.�ʘ����V�<�bE�#T�j���O�806L0���^R�<����`C�ţ�
�5�̠ä�B�<)�"��k�P�9�E��-�mpF@�<���X�N��� &ׄ�@(��Xb�<	�*&c���e&xP� �G�<� O[]+L�Bf V 8��3U��Z�<9���!������O��t�aZ~�<!�*�7h�4�g��dǲ��NA�<	Pi�j	LCe�YQ�%�H�@�<ArER�0t�ܡ�!@�.�m��z�<������nx�i�>�jTq��\t�<�R�2eC*�{�/�R=��X��n�<�'��WLy��=+
�1r "T��	BKɫe{�)���f�P{`�;D���F�fR��Ef9#��@�S�&D�����ۼ^��tqD��4V1A�2D��q�D]�Pyd˵$�+�B�:D�+D���!�@:��0��HT�0�H(D�P�c��P�N�*�Η�C��Qw�2D��J�#��rtQ�b�+OD�<a�:D�@2�D�C��#��G���B�,:D�@y#`��t>mh�gN�|���*ǎ9D�Ԩ6��!�4��JM���`�f9D�� �5�����QZ/݄DZ���"Opt�#�35��	w.ɔT-H r"O(�"$��	lL�$�[#H50$"O�	��W
7u@�3�kD�@�T"O2���"FS� ���@�dXQE"O !oU�D�'�Ⱦs��X* "OT�:Ff���ȉd����"O8T9@�� �ġa�"���"O����&��}���@�S�s�Z�s�"O1����.�q��E�F)J�"O&e��	�Z
�Q[£Ǐ?��1"Or����=$H�#����F�`%�t"OBeS��ӫ��8V�	�C�n�"O(Qh�1�~aS�+�$d�x���"Of	ɕ�̺h�dH��%f��"O�@ȁ����֨��CW+�L�"O�aG(T7n �K��àl��B "O��a -��8��q//r�V"O�l�c垞!zR�3�M�aՐ�"O�!� C��k�(�A�Q�&D�D"O��^ �j���^Yڰ�"O�!'B����Ȅ-S�K��A"O"�aaXU:���m��>��e"OD�bC��
���I��;_��"O�kg�
5&DP�I�8i�"O��J�f� "E:S������Y0"O��A�	�RW,�맩�1-�`�"O�`�FX2o�����gS�)��!�G"O�x�t�J1q��"��X�d���'��%��+�R�`QI���0�'x�"�ڥ4O�1,Ҿ>
ZE��'�.eZ�j&WnJ�9��/>�J���'yHl�#�L9b����Ŕ;<z��+�'�N��.VS�^��G�#9�V�I
�'�~���h7m��|q́�>�,�1�'��w�Qei�I���%1v����'-T���n;FKX<P�Z�R�Z�'# 10S(_*j�kWeW4NL���'.H�F�!h�pegn�?l`��'G
���I�m�F[Fl�*'��#�'Wb�%�߇S�T�dH
�i�"E:	�'kZ@rw�%��@D�C�s#����'���УO\�.�lx�Β9p��$��'d���.��	(x�`�G�=�
Ւ�'�\LQA��l��4"D�/:4�8��'^�@i'�N�/��%"��܇5�
@�'������Xb
})#N�3,��q�'R�bI�1XHi��]�.>�Ɉ�'��h�FH��?0���\�����'s~tQF�
&wiB	��m�$P�������*��)*m�o]*��p�P&.�!�D[�c����o�+G|�2#�5.�!���dHl��j��\��a�k̑IK!��&ytֵE�S�_�a�TDT$�!�DA��9��އ9k޹�q"�?&!��#�J�$��:HUX��b��V!�DL<�.������/�����i!��f��{7��@�de#'��5K�!��2D7�}�EC�&<�Z���E��~�!��<H��en�7��m�U�m!�ď&e�Qq�B�<T#�X��
�e!��HJ���F;zr�x�cP��!�$U5'�1� Jjo��ҩĭ)@!�$?[E�8��g��y�����N͝F!!�� 4�ʖ�
>m1
�x�J�,� �I�"O���j��J� �3�G�>�D�§"O�iҗ�X����G
1�`����Iu���	��&
�����W��ECb�V'!�d���Zx��dC�R����g(�!�d�
�4\s��M�4���fN/L�!�$بs�`�,�6�@Ec4�P�]�!�d��O��h& X�G��E���8/�!���ʪ0(0,��r���J��Ҥ�!�����'�
�V�z1`i�!5�!��s.����O%Y�F@���U�	�!�߻��x��ށz͜Yxa�R1k�!���B��h��ޯ,X���9k!�	4r��3G.�5j��	��!2{!���a��8c*��:YR q�
"Fl!��o>XT�T :��!+��W ^!� ,r쵚@�N�@��1dˏ_!��@&�`��n��1(ZA��h�=6X!�V aw(qc�,ԅ3q'��!�Ps��S���T���oZ	�!�d�Z�f'��!��aSU@�[�!�$�2>�P0�0�/N��A1ae!��O�E��B4̘,i� ^7(:����"O6������O�ب!�Yi,�$��"OL�!hG�k�n�yŨ̬w�D�:�"O���a�W�*HE��҄%"O Q{ӌى\�,$C�M9~�>ŘV"OrQ;W��*H~|��q�.-�-H"O"�1�&7O�PjU��%�6L�"O�Hy�%՟z��4	Rˊpڦ��"O�I�v�ڬA�&9��J^���"Ox�6��o�~e�b������F"O�9� b��F$0�U�2��\��"O4X"%E�lԮ�3.Ǝ�2�i�"O8ŋ��NG���GB4���"Ov�J'f�qnD�F����I�"O�z��´��`R=6����"O��0�;�|P9�[)",X��0"Om����tm��Ԭ�;��U+v"O�% "�˅��m�	��l�"OHM�懌(��j��FG�bF!��y!���w�l��7�=�a|��|�#yUD9�B�?q��-�`H�y"�бad�  k�,3�|]9ceˮ�y�ś%�p� ���(U��(�A%�y2��M�V� Aj��k��Uң���y�Ʈ��!%' i~��뒋6�y2�]nAi����c�N��b�U��yR��Y ��T̀?/��Xy��
+�y��M)&8�X��O4s�̈�y� �*;[|�0�U�n`bwo��yB�O�AȾ����T�
3Hy��+3�y2e_&i��8z`m\�{��)c���yb.�8]��Me��f�2�
SG���yR�\<}6�@��?6�y ��%�y��3����)��t  B��yBA�b�j�Cu*�4�S��N��y���[p�9�&��fP[�N���y�ǘ����(�a�H��:!��yr�Ɨv��� �;=8�}���V;�y��3��� �i�#,���˥+݁�ybA'=X��5@�=�8���G��yrj�	l&��&L+}s�y���yrui��w8��*V(���p?q�O� ���Z"kY��Y��дY��9�"OV�ڦ�͛?|Պ�C�
* ��"O.I���J�V�%C�#�>\��A�"O���k�,"�x� �$
X�+W"O�\�Ǣ\�3��tC���*ɜ}3a"OJ�;f��XJ���2D�ih��Q"OXq��f���p�A!r��Y�"O
T����"�N��$E�5a���"OT��P���z:(�I��QU�h��1"O8�`$��=i��\4u���"OL���艥L������^ ,�a;�"O>��p�L�\g�i����@�)�"O�	�g��Q�X�36�h�!p�"O� #^�ZG��3 y�b��"O����(Q!�`M`q�E�ش�`"O�$�'!�A���"�!~�y�"O��Xv˝Tb�`�p!�P��9#2"O�I�� �:>�,�!�	h��x��"O|H�*?B�p��b V�2�"O�Qs��!���V��!��Y "OQ�2��'�쭁 ��,_�� g"O��`�ǅ�0����A��&дx3Q"OĤ$�ׂ?�Lz�LQ�*����a"Ob� ��x��Tp���X;���"O<AY'�T3hX�dx$���f1�P3�"O�M�OM#��� �'��+ hi�&"O��!�FYF��;�E�.5ٖ"OT� �C�-����&W\��"O�CEj��T��j!/��@�D�3"O<qb��#LŦ�"�nC�v`��"O�h��^�N��B�]��� s"O�z�$�&GS&�Y�KށE��2�"OR 2󋈾`��d럊,}3�"Ov}�0K� En�x���{�xyYA"O��IwE�=D�,="�����E�!"O��iS�s%�� ��^,z�(�"O�3 h 0i�Д7cO���e�"O�ع@C)#0TŪUG��p��!"OP�٠�ы�HJ`F7n���;�"O��� ܛ$��$�T�Hx��!�"O�ݻ�C
,{��I��.�"i��m+�"O.)�t�s��(1G�?X�2��"O$��ɒhI��r�K �8� �p"O*lhe�͊Z��eH�o�
@�9��"O<��N9L���j6ُ@+&$�&"Oz�pl��n�Њ%�¹}6��"OX�2���Y ֌
siѰf����S"O�$
�Aڒ{��|0`"���"Oā�P\8j�	��ሏ�h0�d"O\�������n��$�s3"O�����D��\Y��NI��s"O¥��E���:��_�%���"OXDY�%�(:��-soO 9�T*4"O�5cK�H�Ҍ ����(�m3"O�嘕��?�^�tOګCfH5��"Oh���IC
W�1��@"d��"O�p5�T�/	l�:Ө�� �"O�Xf I}�<4	�g�O�2Yrd"O���DaB���z����C���!U"O�B�!'&�c��$z|1(B"O�l ���	ca�)r̊���T"O�I#W��9W�R�ӄ텃����"OF�1�l�T�n�%�����"Oj`IE���̼�X�BԨYz��"O� ������3z`�H�qcC	���"O.�aw�ʡ(�+���_� ��"O��FBL_��QP+ɰG��a��"O
 	�B?�ĐuiD�c�XI�"O4l�6�@�.Mx]X@/�=VI�@"O8�x2�P�F��!QM��Y� 5�"O�(���A���땟%̌Ej"O�0��<�9��,��ȯ�yD˄�`���MD�Y�h��I�#�y��I�E�~X�#�T��prД�y2��|q���T�4u9�t !�D��y�-L)Y&���e�7��m��W �y���Hk�uB^{���$	 �y�X:c`Бh�A-		6=q�F%�y�h�m՘<�R���-��l
d��y�"I��BU��9}\��*C��7�y�J���tEJ�(t�D#�I!�y�Nn��@ '�'rO:4�r
���y�3`
�L��Ϊf$s2
��yb��*;,��J �`"(B�i[��y�KA�J���V�b�����I�;�yrlҖ(�x|��ȋ9X봴����y2*6K|:���BM�?����,��yr��"{~(ەl=m�\�r*��y"+�,2 6� ���%c��QAG�y��A�:d�9��_�f!Ӂ����y«A ,(���*ǺP�ȴ:�a��y�CH;/��ق�Ԭ(`q��j��y�ǝ���Xw��#�XH[�����y��ϛar�����{ؼ���F��Py��Kԉ�W)դk�H��[�<i3�ч3�� e�J���E��S�<�eo�) �n	���L�T�@a?T�4�G�O"��8��)A��A��#!D�<�u�Z�疝pʅAФ�#!D��H&)FK�P��P V��"*D�*2���\U�$9PiΑiX�Cj)D����րd��� �o#7��Bֆ(D��(�6q����
�_��IQ�8D��B�� �f5 c>v�����i3D�h(�Rl�TP�ڪ	�8L�R$D�Hsg+&��$�e��1 ah�
G"D�`�����;�%�R 
Su�%k��?D��c#��6�����L�y��>D��swI ITZ�Mިa���i��&D��rŃ��Lp�Ы/A�5�`ш��$D�zD��K�Ⱥ�(�=:ƈ�;e -D�,��o�3, �H5��C~Z1��9D�(��h�%3�޵���<�4Qx��2D���rm�6����'kY;>i�/D���#�.&�HjS�-	Z���(D���SE_�X��dI�f V$�m�+4D�h`!�ߍ%�����2T+�ءF�3D�D�($�%�+ɺ?X�̸p5D��	���
�����Z-|��rU*3D�$��#��'�<%��D�.�D���n0D�$ke�ȽR�Fp�0��G����k.D���E�PTX �G���b����6�-D��A 	�?K0\ �(J�ts����c,D��	݊r���8��U?S)�m+b)D���B�^�:>��Ժ��	2�'D�����/5���k�0?cz�kF%D��T
T�<DM�VMʒjA8�3��8D��Ça�o~��1��A:�L�q�:D�� Z�� �_�i=ԁ�"!|T�Y�"O\	��?"�z25"]�fE
m�3"O�0p�&E�A}�1P��Ύ+�01"O�*R�M}0�j�!\�}� ��"OTdf�5AP@mR�ÈW�D=:�"O ����4�d�K%�<� b"O�`��Kґ!�$e���T$��x��"O��3*��H�h�A�	�H��Q�3"O��"��^-n���YOF-+�"O�,�bBW�N`񠮆�wK܈��"O6HksB��D���G�nCH�6"O���,�:<���l�*1U"O��v�K��J1�&�H��\��"O�ГaB3����I�%f6I�t"O�)0K�V(@�!���m�x01�"O�5;��R?�q�07��1�"OH��5N�'`V���;fj�,X
�'�� x��Bm��,9E؉+���
�'\h`�G�9Q^Y��c�3 � ��'�`��$D|U��(�C�J�'�<9�E�':F��+g�,��`�'�pؒF��-U�+�%�"#t0<��'#$QS��[&[�.)F�k�t�k�'8�E�U�U�tƊK�y���'&|��m�aI���X't�B���'v"$b�搭}~�Xv��v��	�']�ĻBn�	�¡�U���bVؑ��'::��AS�, jI%T&D�r�',ƭ�V��l-�Xu�N
PO����'Ր��#Ͼ�3b³O��<z	�'��m!�j9�
d��˳?�8�	�'^��[g�F�oF4l(wgҜv�~݆ȓp�P5C�%xB��#1���A��l��zh
]pl��lJF-���X��Ň�C�&�@AZ+�����.ɖk��B剤�n�F��4NSr=��m�.p�C�ɕy.��� gK�C,p����gP�C��!gjt�`A�&|heE��lC�I<<9���n�;�>�7�_�d�B䉓iP9xw�!��P0SG]d�B�	�+P�}�%�U�R�,�b��B�	�pԥ7,�96�\��V�e�B�+k��a�2���ep ������NB�I�U�.���P<Ҵ�H�f��+�$B�	����]�S��Uzd	�c6B�� 7��xc��^B�~�"Ƀ�cG�C���@��ym0�!G"_܂C䉇!~��oTv�Uf�ZH�C�I$C�J�;���@J���D�١5O�B�	�Ilp�g�2���e-�#;/
C�	�#��h���"*)���.�8�B䉭L��9���"_3`�ċR��B�	)��#�'ڬ%q2��Sa�)��B䉷�Ԉᷫ�*{��tHJQ+��B�	b�m�W��8��4�	ۯb�C�I.F9h�h���9��q�D��N��C��>x��$� -��*A�q�	�#s��C�I��(}[ī�]���T$�![(rC�	�(f,��|����/��wdB�I�t��ڡ(s��2Ӗ{��C�I,V�����8��Xp�O�J��C�	�^d�)U�#��"�� ]���0?фo�-פ���M���a�s��t�<���҈G�|�҅ܓ�0`�"�p�<� ��I$�ߚyw�4�D�&"22:�"O�%��ՠؐh�b
]�0"O��)���w�^�)f�\� Ӥ�8T"O��T�	�^T�9��"��{f�	�O���e�	#�였��ޠSf ���'�
��gS=X�(��`ьJ7�{�'7Ĝ�ӧ�(���i*+B)��'�4���9�x��)�$"�9	�'���3�۔H��!N_/	��p�	�'<&,ۓ�� �b�f%R��5��'^�U�aã.EbP�G3BXTq{�'E�T�JA1@�9 ���6��q�'�ΔȁHԭS Q�#�n[�'7dI���^hxs���P	�'�.�r� ɁXHT�+H��(L�h�'$�qYƬۢp�"�z��%���@�<�QG�	��<����j��Ԡ"�c�<��!$|��0�
�z�f�p7�]�<y��R�S�� 4��N�<���d\�<ËU�V`�#D@4Md nY�<Y��D���!��l{�] ��HX�<F�בt�����51�X�dQ�<���6x�M�uH)l�d��7��x�<�%J��>����ċ�;3�C
l�<���Y4z��Dn
�K���bD�Q��y"���%�z=��J��ɘM3t���y2%�:8��B o�s�UXI̐�yr�aBE��ā��4X�.��y�d�p��Y>�Y��W"F�=�ȓ&{� G�/dC�0S�lK)&�f���e�2��_��n��7m�
�p��,b�,٧N��f:�� NW�bX\��	ϟ�����C�}R�n��i���rrB_{��O��=�}��cw�p��Kp����!^|�<Y��0d�D�!��6H����I w�<��͕$�ڝږEK�G�By0p�[�<��N(f�>R�N#O��S��]~�<ٕ�ՐO�A+pKC�b�\�cWR�<!0�I�M�:��1���|�R͡a%��T��\����+?��I!)��Y�¥B�i��$�Ŭ�N�'a���94�˴&��w��8ǌ/�yBѽ'o<����A,ı*�,�9�y"%�O��(#��:ݺȁ�*�y2KN*\�~���%�*���p��yb���\���&���ġ*@'��x1x3>�9�늕	T,�҄�R[�0��*n��e�c"M�%��C������d5�S�O���05O��c����4M�7"O�����;}�4�0��6s���sF"O�� �#�?.H诏B0d
���U�<� �4$4Ѩ��7�Xr�,Gj�<)��Bl�*�!����D��`\p���hO�'ca\E�f�:n),1�ƩɸS��ؖ'o��'/��$+��a�.%���v(�:��zR��A�<�'�:A�@�9e�[#@�y���A�<1�b�<&lj�
#7���i�<��B��1�Nh���R
��%�d�<��O�� �B�Ύ�|0ش�%a�<�� �P��©��"�\�ro�^�'�?)YC�ŪTJ�<Qw�H,c�
hz��,�d�O���<�����k����J?i�1Qj9"��1;�D%D�0롂U�v��(��Y�e&�`�"D�t�aG�<4��h1j�w$Q�
<D�`Yh[�RDIQ��
!H���m%D�� @�����g�V�3t�Q>.� �"O4�:�oN�[D�I*!�XC���b��|��'�t���l@&1:�kIe���1�'����%��3K�2H�nFX��J
�'��9���S�n웅g�K�"�{�'T�H9�ƠK�d��%F��6��}A�'�Fј��>zƬh;U�9.���"�'D�<�rB��?SDT��G���Ti!
�'M��s�͏?������6ظpH�'5�k4��h��(��.ۋpA�P		�'O萲����ڪ�2�@�<i$��'t���E����2Cۚ1ܭ
�'"�����0 9TXA�+"����'R���sfЬrܱK'U���`i�'	2@�Pϝ=�B"a_!D�ȡ��'5�-����N+�̬f
�}�	�'��37�*x&��#�^4	��в	�'
|��f5X�"�xCX�z��'.�	���:Z���b��Cjt���'M4!I&cäu�DyҌ�=5���	�'cq(�*�0��P��у/�T���'jD�� �p���j:*G���'e4����:H�\��t��7%��`�/O�=q���z����H�}�ȺN�w�h0{�/D�8�B��izr5���KK\\��N-|O�c���D���+!vXٔ��=c%d��*D�h��k��j��B��3s&����)D��X�`�'!:0("�����Q)&D�SħS�S[��[4�N��!Yҏ6D���D�;<a� ��E�|#�=���OT�=����,7��'f�*P�:��th�Ȗ�L��l�*!���p���F�_.�0Q�!��!��5n�mbfK	��Hyr
��o�!�d F� �£�@$l�0�kb*V8Jk!��S�F�J������\�1p���ZZ!�Ƕ[���"�M�7s�b�@�ʊ8Z!���2�6�;kJ�V�ڴ��O��i���'�
uY��ɝhϠ��W��9����'z!�Ğ�W,�B�ˏ$/x����8!��0va"�J�ԇ]p8��+B�H!���.��U���>2��a���|5!�$ێ� ���_mҦ����O�!�� %�:�k��>�D�sr!�ב?���Jr�7�(��K!mM��P:!����7X�����^�WP��0?���׿d+@���A|
��6�Ay"�)�'E���R4+�	q%L��ES�:C��`��:�C&?�V��遌xc`T�ȓRsT� H!x͘���l�Z��D��IIZ�:G��jC�����F�DrN���e��=�5A�C�u��.K/�����.	Yש�3��0�%��:��(�'�ў�Fx�&c��ҡ�
�����K��yR�1���A@�<3B��v&���y���g����-
��Zf�
��y�-N�[l�;'/֛nG�)��'��y�`�F:N; A�<�p(+��-�yR��,70�j�W�;g��(�.ɿ�y���;U�ȍ���(. ɤ���y�>A��Ƀ��4�&���g��y"%�)I��37nH�1%��+��#�yR�¾�R@�5�W9S����'���y2S�0�ؕ��X$E����"���y��[�h<\U�$aX9>�x1K��y
� ��	�mW�Ex�Az X�
rZ��B�|�'az����`D㊛O܍���@��y�_�0�b6�$|��I҆���hOq�
(	Ƭ�%/T��O����=�"O@ݛ�'6�H�p��Lp~��"O�E{t�]�_��tҕ��-B](�r�"O2ap!Â-V�K3�VN$�+""O��X7A�lӀ��YB�-���|b�'���#5J���O�9����6͐��!�CoI fFw�`@�Q�߼ y��I��(�L�Q�/�(D���p"�y�"Op����_ ���JˑEW8̐�"O\Dk�iU�qz0<a&I8r���*�"O5�Ί�P@����ҁb���'�:����{�&�ZG�2]�B)C�'�2���N�Ԝ�f��7V����/O��=E�䀪�f\��MU.1F�P����?���?��<�š�&EvL\�p�F&'j�{i�Z�<A���iX<��FOА)��I��K�<�Ӛ34�J��V�fPb���E�<�D��$-\��D��xU��"�Ln���?��o\XGJm\�pV��1N��5��ئ�C�mצW��X��,+�PA�ȓW��	�茳3�% VD�Gt���ȓOT�!��*B�JaL���VNm^؄ȓ)'�P�sB�r�H����KѺ��K}T�Z(���Eg��~�21��Ӓ'*�<�x�J�+[%O�2t���O�=E���/U8L#��7D���'�өQ5�'ў�>}8p
�=l�!Э[b:H4�L7D�x���KB�Z8T-E,hFLs66D��DJQE<b�ȠJ�C�Zh��2D�`��e[&�p�d�U�^�)�,3D��!B�.tY���F��$A,D�p
�呠n���i��Yʨ��$��O|�O����O��=yd�P$O�B��4L^"��}h#���?i���'p��`��ǲ�̜�`�L"]�ȓe�n��#�,hkn4diE;1��ȅȓs�D�qp���L�.�{��S6���ȓ�|\�ĤٝZ�x\suK�1{ؑ��9�.�A�g;�<u�G�ǖW1>��P<��'��"֖}k2쐎n_>�ȓ�������B�Q�"�(�H��'*�':�\"��O�1�&����hR�'��Y�t^�0�4�#���"�
�'�P�0N��_(�٣�N��y��Az�i��t���F!!�y�Gb��å��
w���K���y��H:\Y�)R��'p_��TbL1�ynH�t;e�Y�dlL��!f���y"
P��YeÖ,XZ`�Å��y��!
�h�x1��Wդ�3B*ׯ�y�	W1�s� '^�^0�1E��y�@
tH�DلbU�XO<`Q�+�yb`���lp�G�D�U�`�����y"�ʭ%H��[�K�29G�9��F�7�y�l�f�N=�E�]?,�	q���y��'c\�8j��B�bF�S!=�y҈
fi�x���tI.(á�R�yr�˨@C�9u�<j��Z�"V�y�A].����2FJ�`�@1���yb셍c��P:�(��-6��HK��yr+�1�R�`����$*~�"L��y��D!2�]a!+�$0LHM"QJ�y
� ��I֏
��3G\� ~h�0��'��3)J�9���P��8�e��g��B��%k<(�14���壌7"�C�I���ۀ"A�a�
��d��7g�B�I�wj�J�<MµJ1,�7@�B�;�*�y��(@�U	D�)c�C䉵D�@��h`�!�ʈk���H��	�j�2����Bw�B�T�J� ��B�I�'�����bv�9x7K�,���ȓaF$��B��<r�S&��t��8���pQ�F�D�����'�ń�	;��+b�8g!�ӫ7/*U�ʓ*�‡G�F�8�ird�<D�jB�ɑ*R� � W�&+8�0��1�VB�	)o�U�!)]3K���	1GđQ�����O�a0��ׯ$ʆ)W'��X6 D��%/�*B���aL�;'Ф�;D�,I��Ʃy��"�F\o���b�i$D�a�N� s�����3W\ Z�K'D�(Zq��+R�` �B�6"#X��� D��%�3/"<�p7-��S��	)D��"�a��W�@1/I	����%�O��D�O���F�1/d���T�G6`n~���&!D�����$=Ob�hA��99�n���,?D�\˓B�M�� Q)��m$X4�w9D�,Q���T��]���V^F0�D�!D���o�`�v\�ec3r��*6� D� 	a#`���� Q)Y5p�`�D4D��P���"N����iХ9X���?�O��d�Z��	Y��^l�|+@(����C�	g��\�!_�0l.i���?P�C�ɤ��H�4��\���%��v��C�	�~�h��5,Y�A�ؘ�bB�+_�^B�ɑ�y�
��M~���j�*G	*B��$>�FMa2a��M�t�B6�*$*B�7L���O�U�&����
W����z�`;�!�(�h5k���+J��	�$=��K���T�'b�QV:qM���Ê�{5ja�u"OT=��݄>�Z4y�@�$t�:�"O����4gp"��n�E�H�"O<�*@�֨�ȑ	5M/.�6(��"OL� H�h�8��%�˃�ע$H!�$�T���7m��R�*H!�I��d�!�s���	�E,q��˦EL�N��Oz�=�+O4�jU�(�| +���80K�hs�@�OrC�		���P� ٣6kbБ�FǛb�.C�7@^6Lr!/�_�Z|�����C���̘���S�S�p�1G�Ήv�B�	�O�Lzi@:2*�8Y��L6HC�so>E����?�p�Ŋw�*C�ɥ�̔Q�G��l��T3A��=�H>����J9""��ۅ`�Z���8������$�Op��'gǚWB]q�u��C"O8�k ��g(M�sI�!j�|@�"O�I���Z�zU��)�Iy�@"Oƹ�BO�����лd
>��'Բ�s���:��L����v�1R
�'�0��Ņ�\FeP��\�h ����*��p�΄�N'2�a �@�z��'w!�d�DZ.�( I�q�9��]6W�!���9�����ƘV<��	C}!� �ᤅ[����S�^�Y���]m!�DS�L�zd��܎H���aţ o!�ʳ`�b=���'`4޸XPb�t^!�� F�J�l�]6���VO^2��9��IH>y��6L����D�Z���bv-:D�����r�ԭ��>c�ĩ�Q#;D�@3fðzD�h��K�Ab1*:D��� N�}��"�疓b좥�e�+|O��<?�4�/!(�'� ����'i�i�<a�J5�h�f"_�Nn�|�<I�ϋ"dڅ*R͟1�D��a'v�<Id�(S`��)E.��v�.}@R*�J���hO�-��̘��Ņ��YD(� ��ȓvH\m
���w�r;��QRч�Ej��y�i��֝:Ao�;Lr�1���v~b���n���G�NH@�1W��1�y��Z7f��Tb�?w>�`&.��yrO>s+j��昤8a4݋e�;�yR ��	�nX�F�ڠ[�����?���0|"�$֣z�tQh�" �@��5`�I�<Y�l���x�Z`JA�(:�M���Q�<ђ�29*F�[`eڜP��x#Du�<q�J \�\�yA OH��IS�z�<�#���D0.�HU��3A���f�u�<E�Ń>�	��%4��rA�^����?9���O��2S�8"��Y�H��y�J!�DL�@! D�|}̘�rmU}8!�$RSG�Yd�r
x<��L��x�!򤀉f!01� Eי#M�r��<(�!�D/�dH2MD&=��lS���Rv!�Q�2����J�*
,"�FО1S!�-}>�`K���u&
�Ge!��Iy�ԉ�� �M�BdΟ6!�d��zU��wD�ٔ��:�!�_I����ŕ���h� ٶX[!�$�+�p�	��Att0��
�8^!򄜚R�(=�Q��xT8��f���!�d�F��)�cO/-�� ��Zk�!��úq�>@a�	�	[�`:��*m����#?(��G��="��D��\f�B�ɉj�v�Z��[�sVD�T�,�B�ɟ\&}��.ٔT��Ce[V��$Åa�M!��)�¨�!fĀ:(�'vў�>y+�&Q&eF`k�ɚ�`�R8y�a#D��5D�Xb��T+��u���qN.D���C
Ō6�Z):F��&~�����L+D��+�]��D"�RYpƁ1�.D�����N�8o���ǐ�G>Hr��+D��H���5Zz,Z�jN�~wE��3D������s$e��J�@��q %��9�S�'A�荛aa\2R!8l�5H�2�̵��~8��(�(T��X]:R	�6B�ȓ�h�uʉ��n�(���*$fŇ�S��p׭�N�������7�ɇȓ.�⁹7�G�!�D�
��(��`��c��İg�F�.�t��˷Mg���ȓ;*i$����԰�C5'#'���IS�Sܧ=|��J�g�.����l��ȓU���0���+k�D�4��TqBh�ȓ	F��+/�<p���4"4~5�ȓ%�ؐ�g,�;^�$H҄%M%�����;1"���Z������T$\��h�ȓ;�Ȩ��KX��X�▥״st������Cɸz�@��!E��q29&��$�@��m�O�,;%��2�TAy��ջX_,��'0�1ѕ�C���3-9ϐm��'S`�i��S������!<ޖ�B
��� ����A�|����bT�
�3"O��A�ӤI>~���V�O�%�"O*X���3M���Q�^�Y4q�"O���6.��"rؔ�Cb]i�l��u��m�'���9g	߯@ޤ��C�����0��"OYx옲v��(X������q "O��Z�AA�h% -��쎜G�V ��"O��k�?,(��C�ۜl|�z�"OHa򧤃�t숍+���zV��"O���"�$�p(��+
/EH�Y�d"O�	9�i565�8�aɳvA:�@���S�'u�D�I�܉g��3 \���LoRO�`�ec�urqɔ���:S"O���4�����I��]�p�	q"O�A:P�ل�F%��I_�k���2�'�ў�I�<&�T��J�y��l��M�ul�-{`�Og�<	����(�� ����"^X�<Qo˿w��� 5a�!g�Q�<��i��}��Bh�c�\*6AhB�	�K�x}0Ī�)����P�%XBB�I�/��7GB�X���Uh_�3 |B�I��m�2-ۈz`H��Aʎg�0��d�<�O��e�D���Ub��"Ӫ�q"OB�˶*?� �['����i�"O�r#Q蜄�1�_�9���"O�"C�L8��`�8���y"OZ5*t��
�h3��?ﲔ�C"O x��K/΄I䀀>Z:��9"O2Up ���x|r�+K'rf� �E�|R�'.b�'��O���<J��湊6�*����B�4P�	�'�:x���1wO�p��ʊ!ON��C	�'*�"3��n���[�OF�K��p	�'�pD�)>�<E�CP�(L��'ָTx���$���*M��d�r�'("`M&qb���g��nL�'le�A�ʅ0e�؇�ܞx��S��?Y����OJ�S�'��x��!�4A�^xa�!��E)��	�'ڲ���쓊5t]�S�C�EI�'Vf��Ej	#}Lh�n��?V�@B�'�̝��ؼ��a�*=�2H@�'@��i��χ#���%���5�$���'�T��ԍ�w��M�+K�3��"Ov�Q%*  �xP�7B>Vn�H��D&�S�I�=�֌����5o��h�ԩ3�!���!Op(�Mx%.�&ɋ�B�!�dHR |�G 
6$����Y?3�!�$�7f݆a���U���"H�^!򤝖o�h�2'��[����i.cA!�u�mi��JN��\��
cC!�$�O���QW�wh�pZ�@Ɲt5ўX���e��<	t˒�D�h��'K_>�|B�I�,#hH�7�Ù,��U"��DB�I�Rw8�#�|r�_)O:4B�	J�0�;BbJ)�P�v ���2B�I*��u��C#�)�\>(�4C�I�{V���	W�r����L#9,C�I9H���V$�K��(I��O�d|6�?щ�IS+: z��O?D��H&f�j�!�D��5k���(��eƕ"�!�E�H8p`A���aŠJ�H9�C�;y��׭��_ ��
�BC�%aG�#�-G�f���#��-�fC�ɦ"�H<���[�� TC�I6o�p�UG�
�D��w�I�T�?��� ��W%B:A h�3��ݱyL�YAD"O�1�č,�V������3D��"OЅ`��ЕM�F-��@M=!����"Opl�C��ڲw>�!���7D�k�B9g���+��b��7D����gGK�[��l��P��7D�L�Df�(�J�٥�H�@E�x�v3D�tKפ��:�SB�k�t�"	6D�<db��A��݉Uk����(��g!D��b�K���|aJ�q�r���"D��Yj��GL�%A��B�!D����=jv��a'���l�`�S�2D����]<}�⸂�dƤFJ�g�-D��cPGC =� �0���.cd \��9D���C��9�����Y9���c �8D�`���+W���&B_���ɲi5D���P���ZyI�
ԇ{��1!�@>�Ȉ�n����VWz<܂s����u�0"Ox�?Cv-��Q�L��Q���y)˘��	0�
�	����gN�#�y�HV-;�r庥��Ut�e[��O�y"j��N��W���i�y�W!-�yB��`��Ly@FU!S�q�'��y�	�\"��EL>~�ά�6b�9��'���O
��D#Ҙb��8'���BP����yRjjcuyq��&fld�qЊ��yBh�>T�<����]f�!�d����y"���v8�9ӎA�Z)���g΢�y�.�UH9cS6{8�LK�F7�yb�Sd( ���y����Dm��yr[��pe���m~�Dh�&����?)���dL܄M��J�h߼[��K���?Y�'����U�)`�ɹ���.��-*�'0B�@�fAg�C��
���'nf ��V���1AdÇ �t��'ֲ�s�4g��	�3�C%O��Q��'2D	0DŖW 40A#����Y��'ͨ���Y	M!ތ��ˏS���+H>����?açQg�	��A���fȨ���E�L���I~"d�)9�\)c�%ʁ_J:m�C�D��y���'L�:���=Y�`i��$���yҧҸk �� s
��`d�!H&C���y�C��v�R�H�`���`���y��. !,���I��/�8qеJ���yboϣh�zA+�-�D4�u� ��d ��|b�y��L*�1���\�}1�yb�;)^M��`^]l(�x�����yB�I�X�S���bM��+=�y��� ��X7�f��TQ&���y���a�$P%g۫g��x2v#P��y��r�i#$Ğp�[FJqI�ȓɔT2��C�y�f��O�D����}�$d��)Ȧn�5
 �>�
��9�ecK�%oYp���J�8aC,|�ȓv��bs � I��]�d��"4��ȓqe�%����8wT8Q!�"B=FeP�ȓ���"��Y2R	!��t�]�ȓ@
��F�RKF���%R�m�h�ȓwD��{�^'8�� [V%��6r-��Y �y�ʴ��#rE {f��ȓ���e���A�4��Տ��̄�I�֩ڵ 5��9Bd�\�0��	�ȓNӂك��:V?�hZ�ϕ�DT��[�|��#Q*�i�MǘQ�*���S�? ��"�'D�@���BL�X�a"O�����6zW�Ȫ��޼D�N���"O6���ε%�u��kQ��N�!�"O�Qi ƕ5@�� �EQ$+��ٙ�"O���ÍH&qA(�U'�B�`pq�"O&9�$��w6c��F+��'"Old�%e "�9Q�qS"Op���g����$� �5�"O a��H���3�T�P$bq"OB���M�R��M
GZ�|�b `�"O��	�����,As�D�I5�"O���N+��#T�_�e��<��"Ov�{F�2"l6�;B)C�k�*m�T"O޴Ƞ�J�>ȕ@B*��D��#s"O��CP]:� 	��(�I�HI�"ON`!�ߊS��*���=�H��R"O��ŏ�;z��I$@��XӺ�
"O������/ +���0�$����"O�%���T7y�����fRfn~4��"O>�ʠEO��
�BƳC! a"O�8#'QbN9�jܡ!Ŵ��"O&�t����V��ɳ�"O:3�b=9��(��.B(vy�Ԫ��	ϟt�'�1��tF�q���c��BQjPHCt"Oĸ�'�/l��EDH���"O�QsS�
 ��eÃY�D���"O�P��2z��usT��B�j�"O��� ��E7@���3� 5��"O\���
$Gc�xb�Ԧ�
�P"OT�q��$��0� ]�
��ȵ�'���+�Տe2����	��1d�%9��$�O���B���IP�$S���$4W B�I�tW�1�'6�j�'F�
B�"B9'�
���7�[�O7�C�I�R��ĉg�/T~�%A�AFxXC�I�9��dZUf�'��1�����>��C�ɹ*����t�\�=10����Q�zB�	WR��ضM�N%"�i���#H�B��Dl�l������YWϠe[~�K3�'D�pQ���p9���L=}NL	f%:<O�"<q ����'�=g��MR�� [�<�B&��{��q!b�_���r�j�U�<��nY
��0CAM���@���y��V	,������4��T�"3�?����h����%��B�R/_�b�j&$�?4�}����a,��#�\��d�N"���C/D�$j�*�?�} �o
.�m8��2D�k�`�^�̨+YD��)Ƅ#D�h���֜ua4�Z��pI��;D��F�0x.^m����YY�U�d�8D���/_mj8&�	%��q��<YH>Q���O$��D�b (�'�An|����'R�I :���I"O�aG�m2EA�2EC�ɺ@x��������v� 2�?a����#;�H}Qg&$�i����I�!�䞨w��*'�<y�,L�Ҋ�q!�D�t��$�fc�9��ثA@�y4!��0��n�u��<���Μf�"�'/�'+�>���l�����W2r�\��@O�t�0B��Eh��5��I�)���:�*B�	�K��b� � 9�"${r.
�btz��8�I��G{2@ѓ.D��G�h�(�ZW�B:!�D�VG�,�G��$���� �-!�d��Q�����,xpnH3Chȅ�!�� �e��L�FҤ	�+�� Ja"O`�@��C�$���r���}�$i0#"O�qya��MR24k삠�(���'z��'N�ɱp�b����H߇T�#��',axb-��W�}�D�]�V�x���Z��y�����e;���P,d��g�ǭ�y���z^d��� ٿOZ����	D��y�lQ�!��b�K��5�j�a4��!�y2��[9�3�W��PTsc�+�y�Ѿ�s'�Q
�Ε�!����2�O���bQ�t�f�0��<(��Sc"O�C�i�!�h `Uм`�>�4"O��X�f�=�
$�0���	r�!HE"O���J�v�4rd�kLԺ%"O2�9��?�"͓"��Se�T�"Oxe'ǋ^�n���S/XyA�"OJi��&��T�f�t
��K"l@�X�D��	�8��B����x���qs�A�4�C�h|��� g���x�Ã�$C䉼qI�P����喍��CƶG|�B���YcGIP
�fq�5A��B�	"h���Em_�3�(�Z/�)�C�Y-���f��:8 c��-�vC�	2�(݂f*X5/�Ӆ��n�2B�ɎZ�h!c�:Mb�$+b�2"B�I ���+��ݾ��ISu�d�B�I�{IZ$1�&o]��{����C�%9���V�F��e�`"� \�zC�|�X Ggj�N5��۫+�PC�ɒP��C&��5�2M��Y��B�I���Y*�Ʌ�欣�?A�<B䉆c[x�e-���s6�¤	<B��6����G����C�E��tJC�	�#Gi'jbx�KEᐐ!e.C��	)V�XFX�Q��i�Ȑ�`,C��^�h@q�I!;�¬#W!ٴ}�C�I�>Nl	�`�4����LH��yb��#�.=A�$%{r�,��Cގ�y2���v��*m�>���ز�yr��WZ�A�b��3��(�0O�9�y�ŏ1-8j܊QȀ�Ɛ�5�א�yr%�T���K�h�՘d�Ϝ�y"�G�H� ���`+2�z�M�'�y�#��P[���F������"D����,PK4��q�qU�y��	�0(��h�-�&lxQ�N;�yRd�	#�9!�F.1RDp��5�y�II����j�n�'�e�p�˙�y�\�i�q�Ug֯z��X`�A��y�
�3{�iq�H�<	v�QcN���y��O��z)#>Tx]�rL�6�yB�Ha��݁5
�N����
��ybl~�8|�䌝�?C��	ՀE1�y�T�X\FՋc�PE�4�d����y���\G�@yu�?DL]����y�Jt��� ��.1�������ybnZ ]C�l;�Ӫ�΅:�.9�y��ΠQ��yw)�}�&���yraܙ%����c5���F��0�y"�ʌv�B�Kq����^i��ۍ�y�LQ����+Z�W�j=#�n+�y�B'OP"���m� WP�p5H-�y�B�q���E�pTX0��y"΋:Yj�D�Pl�(<����*��y
� �lz���/䀢�ŉ�T*"O�12�C&o�`��`c� w��YBT"O�4R�T�Z��uxw�ތth��&"O�x��]=Ib����֐����e�<����	5�a�e���Y(����y�<9��)+6�xa0%��k
J���c�l�<�F"(h��5� ���x5v���$i�<�@d��H��ܑF'�"�#։�M�<�[+0�4PBခƀpsEƖH�<�P`Ls�����ʢ�l�{ �D�<A��G)�%�AB��F��"�A�<Ѡ-C8U@y�q�ɾO�r !hM{�<���1��pa&Ȁ�1Й굋m�<�v�O*GV�;q��0r�
 ��M�<��?t0-����K��m�+W�<q��.- d��hȩ9��@��B�<!�A�>3���KA��jn��zpk��<�`�a5���W�ݧ"~�ҦD�|�<�Z$~:.���s&YBծ|�<Q��4�xe-N�
�|͢eLC�<�a@2�u�$ꍀg�,TzwB}�<��oB�:��Qi%-k�pb�Ey�<��U5!�d���S�{��i�C|�<��B� b9��Ν�At��F�^�<�4�@2V\��"Ӝa!Lh� g�E�<Ih2����G=�!6��D�<�5�R�A8��{���<N���PP��B�<��EB�A�7aҴY�^U�<�%�(%@��Hs.A63�>�H5�CP�<��>8'�� ��&t{ �H�L�<��a�NkH��h�"u�>�s��OE�<�Q��'vb���l�"	2ܓ��e�<)�� �?q���(A�րYa�[�<�`l��(ؾ5\4\Bth�Y�<1��K���RB�T�>�+���A�<�E��v��Qa.S5h�@H���]@�<I���1岬k�n5!
�|b4��~�<A5k�>nE�e��R1f��(:�~�<��-m�����F��-l�c�%u�<d@���r�C��TB�r��l�<q	�-oR:�A�酿c����@�e�<q�)�xFJ4R�� ��������`�<9Ԉ���	`P��F&��ֈ�E�<!#��$Q＄�c)��<� �h	@�<�rD��&#����;Ș���a�<q�A�L60PS⍞8��1��M�T�<�.�	�9 B/�;�ݫ�)�i�<��B�1�� � ��%"�+d�J�<�'c����2 �P,E��Y� ��]�<�V��(�e9 �ϼY��r�<���݃U攠#�KK�\��b���w�<qv��3^�\a�T��>�v� c��<)2O[�{�
abFďtr2��`Lt�<I��T/D�|��F�D�
�@�&�Y�<���"���H!k��U"�遅W�<�T�L ���ll��EלYlA�ȓ%ff�0�ߡ#��uq&�ʢh{�����(it��y�ެ:�ܵQ���ȓho慡"�"��� ��/?�����N�d�X���"����!�\���I����ւK��mK"�#VX�ȓPR����.��{��k��٠R�5�ȓ%���J��$%R��
�L�`�ȓW^(p�ѿel�ч���xP��S�? �@�iWrE���Ҝ1���`"O���O�4�xqC��L�HX"OV�����\x̹#Q�ܧ3�E��"O���f�#Z,�Р%�'�>�0q"OFB"/�5^�d�h�F�!z��E�""O����A8Jt�X��%�)|���x�"Oz����vZ,jQ�������"O����$J�2< ���V��"O�C"j�@�vQ���J0\a`"Oz�q��5}��!q��BA4Dc"O�0�(����i�ЍN�2F�s�"O�X�El���5fJ�'<�0"O
�8��H�^r�y�B�s)��'"O.�P�惙_���z�а��W"O���L(>p �B�%�|Ը�"O҄��/˘u2El1�䤀�"O �:�D+jԬ���d�� @�"O6I	�Ș]t\��$�łe�����"O��؄�Ѐb⦠K�CF;����"Oz�3D�D�)������"�x��t"O|��g���j�.�CU!T�`�"O�L)aAԸq��)�B_��(h"Oh`s��	*ot�09�O���Q��"OȀ8����1�fDa[�E�l�n"D�0��矄&��L:2A�`n�ͨ��8D�x��
Q�)��e��E䪕�D�5D�	Q�� �p�;p��	���x5O D�B�a;(�(�c�I$}JX�u�#D���E�(|D�c���C;2l�!D��ʗ��;9=d�@lA-P8P��>D� S�H۴_:�:�+��Uv���B-;D�Ȑ�N��L,�&��><��dm-T�����:$h�r�,O#2�dp4"OR�X�UF+ @���[�*B�Q؀"Oʴ����%gj��,A>���*O*aࢃ�ot�<[CG1n�%i
�'NJ��EOw�颓��\j�d
�'qb�{�������G��
�'�N�H�ʞ���X�BI:���Q�'�����i[�9��膋ƫV�Ex�'����!���s���2��#I h9	�'�:`HsbHɀ(	 nԕ?:����'*"�b���:s�h��º;vQJ�'`��X�,��2q�I�%ۈ��'�}�F+��C@\�k�@Z5#<�x�'�����mA��-�g�K�J�<x�'�2����������g˙L�Z�'��A �=\+D�Pf&�&	�Zx@�'������Gt\9v�	�|����'n1K eh~ĸ%1r	:�"�'�n�h� ϛn��H���k�4��''���tC_ 6���p� ܾgI�DS�'��as�C=:زlP�@	L\��
�'}椋Q-]��v@!�e��L�}�'(d@�.��t�ҡ!�d��K��}�'�BU��O�QmX����A�1	(ِ�'���Y���]�$��]��'�V�Ӯ�v�h� ��^4��e\���<����*H��� ���L���i�&G��}���������@��A��I+^ك�7D�HCD�\9kT�T&иul"I�i3}R�)��9v�LIq� �qWH��f��c�؄�I\�����q�ӥE�F�����a?)��P1��1�D
iC�W]�<� ��E�?W��R'��\0�!t�'>ў4�n3Wтl��N$5 ���!D�<��E�=z�t���b��I��"D��j�&B��ܨA�%%fN�x�G>�OP˓���1��_i���!��Q."(�'>R�'�x�(���*R����P���;���y�>�`�3$ -�D��?�y"퉲Dr��ᗉ	�(y�@��.���OD#~s��	#*�ؑ��,"�����D�<��eV#F�Q4g��f�+ph�}�<af�U fB�<۵�C"]�n�EX� �O>��Q�
o�Q�whۗ��݈[���� S�2e�����HP��I2���5���<�;�(�2u�$�I�e�`��&�-q85���:D�$"a��[\�E�a	�6@�8�9"�"D���@[�5��1��Y�\�ڡ��H D���gNY^����?�~T���3D�ԨQƁ#`����ޱ@�L|���0D���*W)H��)��
ۗ# ` �7
,D���ƙ.
�zE ��\��'+)D�\s�n�1g���t�V�
��*�"'D�����C� �l3C*�2 �:ykP�$��hO�S]�:�k1e�\-�8�ƊP�kb������`��J��\v�6� A-C|C"�n�ş(�?E��4q����7/�)a�����?�LFz��~�b�;mQ�Di�D�<H�
ف6�[?!P�O:��dOC��n�Ix��[E(5P��r��1O\��?���JA��P�%br��⤗pH<I$LV2?,(	�mB>� !J>.��	h��,��+����x��.&�S�A6LO�⟬z&�D�K���pL�Ȝ�S�N�>)�>ъ��wn�q� ���2[Q~���[j��&%^Ni�!�@���s��p�>�ۓ�����+��s��9K���,[�B�I'R�6�!4���{�\Q ���6Y�C�	?/����bED���$��eɘ�DUz���I$�I�n��E���4(�$��"^3�bB�I,$��I��ȞZ�K'��ŰS���4�L	Qr,@.��c�Ƚ8;f8��N?I���ϙU���� E�a��-�&�)���<)�d��NْC�L�I�.L� �d�''@8Fy�Q���F4�D$�7"�6����bO>��xB�. ]��ᇌ�S%��VA�$D��o�P��h��q����T
�+4D
=b� ��'�qO�"�O>�"�'��fȅ�t"O�Pc�	ͬ|׌ԁd�)~d���&�>ъ��)�	<����s#�'.��{���fF!�D�A5��5�Ȁuwe�592���)���`vn�*T`JD�L�~�p0/9D��`��_H��;��ؙ|�@���!x� �?1�ט'Z�S4K�:���@&�Z��ML2#���m�H&��ib�́53Xg��h#��!�v�8	1H�S�O����SnS%,��rO0uf.��'k<C�Ϲ��P� U,q�ZTA�'����Ȅ�V�Jm#�B�<��1�'�s��6�P)��A�
#|uy�'�����	 0uL
q�-o�{�����&eT-Oc4x�f	r ��#��y2荿~_nT�#%[oD���&����<�OR�Ђ�*I�����m�3.8D�(��	D���	K�1[��'�+�6ذvCN\$!�����+�C���� �0bA�1�k��ħ��I�"xRa`ff�;_�썀3'��Ɠ5*r�j� fPfru��Vٖ��	�<�5�)�~�H?��S�? h�ℏǣ\ŠMC7�C���S�'��̧>iCH�h��$�T�R� ћ�l�[y�'�Jy���'��5*膤XJ`�CU@�)b|����D#��?��ɷ1�rϒ`�$��S@�; )�U��!8���s�Ж*a\X���y��C� I�#N�E��ܐRLL���M�g�Z5���?NIt�Y�!Ewar�O�q�g���̦��Q��j���'ԛ���{���U`ި Y�yA�g�,sK�B�I"1��tS�&�)a�z8 ����G���<E��B2	 @L��ѱ`EN�T��y2�>x��sLŖ_��I`�lÌ��'�$܅�I<#�n}�fi�'	L%��e�5|ߐC�-)�H|ˇ���`�`���^%A�NC��uV�}'��9iE�� �Z�RC䉃B�ja��۝'��*v#�
yvC��3k�^tz�T+D��x2�LK���⟬E{J?����o�B�+k��^�(���:D�� d�!"�jLAS�R�J�X�{Q#7D�������J*`t ���t�v�	�A6D���U���x�TykR*�oF�tm(D�04E~�U����9XM�%D��@�e��Fpd3�eݣ{��l���"D�T��E#p��� �'r����,�$��1z�%�$��}0�Y�A�=H���p?!��܄mD��[�F%Rݓ�
y�<AA ��`� ��2k_R`��I�<9I��h�݃��	�@��(*���o�<�g 'i��xjgk�
{\z��Jk�<����(>��SSÔ��ZÔ@�<	Ď̂qp�أLN��X��c����?����:%T�a;��E�}}��3�O�X�<a�B�'6�L��gG<l����`̓ט'�0�|�JH�f�PdIp懸F��]9�/IY<��85�a�Q�p܀3cPD���'�ў"|*��-,AD��KF�΍0E��v��D{��� o������:�KebK���'���$�&
I\x��BMD�9�&O�GR!�4���2�*G*>�	i�M��!o!��ڶI7l��%�+g�RD��ƛ5���gy��'� �ca!���\��BL�4�
�'��d�`�ͪ�t|Yʈ)t�p�b��$<�S��b���&��Htb8 �jɛ�y"��]�@����%,�q���mZ�Q�Q�"~n�$2. I��ژ!�4���H�P��B�I*�v�jA�Z�rrE/��.�B�!�T��N��&��YS��h���	v؟�k�%�;9B�]��-��kM��#5D���1w��үO�=9�'�J�<��.�
"�9��K^j	.��#ꓢ蟂�3�@�$v����$9�(;�"O�l؅���.%.(z�OD�+�aЇ"ORT��oÞS;�uZP��fQ�"O� �[�v�`��P�Åh�au"Ox�Z�)ǈ{��K�%*�@}J"O���P��	4�H*����^`A�"O��GLΟAJa�s	; �h�"O�ț'30PTH%ŏy�nppE"O �qf �z,Ȅ��m_�N� �;�"O`\#�#X\4(P�ވ(b���"OR���������wϞ-T��"O�P�T�*8��i���8�<���"O�1Ɂ�7k�vd�qDH#h6bUc�"O�T�q,V���-�Y�
� �"O� �Q����4X�HJt��"3r0���"O0�pqBD�D2E�sѱII\�
�"O�L GlL�Y��M����RJ7"O��`�śH��Г�+�:^$��"O����Z�0�٠�, �2�"O��s���d� 0���(�n��"OmS�Z�&z:Uб��\~�\R�"OL���ώ�k�6	�ݳjl8��"O`�x5Ș'd��"dH�N��s�"O� K�G��d�"�� �k�V\@�"Oh��AN^��y8)^-1�<i��"O�A�a
�$��
"G��\�\H�"O�Y�W���]L	���U��P�"O�Q�EW|�P���!8,Y±"Ol:s��2_��d��I�%}���"O�Hb%*�>����e,z�x��"O�օ�Aײ�� ["l��p�"O�<���7Lr�m�`�,	�"�`�"O�	A	������Ώ�ʆ��`"Ot����DZf��\1���"O���uk�m�F���<d�p��4"O�E{�%F�Y�e��.C�f�(Ɂ"O H�#R�_u�d���ƉC�V`3�"O
���A'+���Y3$^H0��"O���gJ. ����~��Y�"O�L�"e�X��Q��F�-5bΔH�"Ozm��)VT�bd�3�W�Z	�p�"O ��Aǋ��4X�m��E�  *!"O�ya�/5$�p��6%��i����"O�=�`H�6ލ��ж�`�"O�I!`��5yC0$���Z�2���"O��b�S�)F=��I����9�"Ozi����S�ڕ*0j��A��Ը7"O� R¯ײU0��ɧI�E��tV"O��	001@�0���"2�X�"O>���Y�+�2� ��=g�T�"O�]���T6~l䱁�ѕ*{~(��"O� DȢ3fA Ӎ��`��!�"O4���D<Hf�a̙{�rܙ�"O8I�!͈�c�f���i��t�$)I�"O���c��_�����G�2p��"O&�s�B$_��=A��:X�ƕ0�"O�l�1"A�RXÀKL�[��|qu"O�4��I 4E2z��'I�����"Ot9Xc�T�s�,�y��6$�*���"O����/I�z�Icg��$���0""O���Ǚ�3 ���Gm!3*5D��;��l#��3W��v2��t�Nm�<�"M�A�"�QQ"PM����c�w�<��J"f��e�Ň�"4��x2�	Y�<�`C�8�J��U�E8�| "�c�V�<I��R�qf��IG?Pxyn_P�<�ևp�Lڦ�;?�B@[��N�<Yw.&bǘ��G��81'�L� j�R�<1�eD�GcX��%I0M)x�����A�<1((�~�S蛲�Z���&C�<9�$DOǠ*5aγ+�~a�''{�<鐏ߗa5nА��)�H��g��J�<Y�H�|,Lp$`�{�2�Q��\n�<u̖�3yl��т��T�1�G�<!��DNl�i�R��\|�<Ac�2|C�E%�	�ڨIIwL�}�<a�i �E��r�]�	i�U��";T�����Ԟ�&�q0k%c�ˤ�u��I1,B�qO?� t�9�aH:�d('��
޶��P"O�q�H�;l֌@��lJ�Q��X �Q�\#B%3+BY��Ʉg<p9@�գh�Q���P��N��$!@ȁ��,��!A��"7�s�Ԋ0���u
�'�mq�)_�y���k�͇8<�J�+���_�u�����Խ��OvĔ�K	"����s��3�����'O������9���F�� "U,���4:��B����lӧ�����UDX�z�	u�D����p<qQj]'��'#Mi$iJ�7�f�h5��\=X�OީI�ㄨ/����
ϓg�Dj�˂D�i�ᇏ�z�'�����CO�S��c��r��h�������n���x�"�=n��7H@h<��	L�q�����Y.�( !�B�W̓�<,q�b��ؘx�k�*��IN���۴H!�Qr�dH�hݤd����D<���x����ϨEMv�"w���Y�����iO�:$�:t��/��I^��M�p+ҭ���rƯ'�xy:ed������}�qO���/VU\�!���C.���c_�����4 R��'"e:�ΈO���AM��~ (�Ofe)PfÛ鸧�	ڎ|9[p�S�RO��`�*�2Mӄ�9��ʄBoRT �'&j��� O�������'j��0D�P㡎 N����5
Qt*P��p�g}�O�fI@�ƅQ-r�8cC�Lp�˓	�R��!fB�D+"�\"��$�۸D�� �R��RJ�ϓN���kĨ-�)�'$��YS �
Z�4l�J�qM���Oa�b�U��D{��;�c����#�����p�O$�3R��,�0=����T�upR�Դ!�����O&g�yiP�x�B$�;�q��N�L3������#_Z���-a����$�Ԋ�Px�@\��` �H� �X���n��<��i� �(!Ҝ|��@��8�=�S$FFykD�$���KEI�7����-+��7���2��_�ZT�Q!��5�L�#�N�.��)�θ�!�����S�O�Z�"rQ�`p�8Q���-In"�
I��YҬ
]��t�eB�k�OZ�]�W�C�p��܂�m˝Bd{L���u%9��8Ǔ2B��H5��E�
��SM�K=�lx�dڋV���5GT<٨2��l(�g}BaLn.�J�	��80�$ՁH^���됯%^���ɯ$	N1���s�0��4g��X�G`���t�䓻�ē�Mki֑K�6��D��z}���5{�B�+_2\��a����L2�p��	�e�h�Do�(��DO"S�@��%l�|����!e��O�1Mo�\¦��(5!v�	A"Ц�~RF�7`9\�Y���	���c�4q �W���S�ȁ�g~�O��C��	e|�	f�}YK�;&����&!a�:yh��	+D�a�D�I:I�e�IOw�����I�y��h�Hp2�S��ɪ��};�옮�P 2�)L?s�c�\�{q(�'23��Qt*�7{ڀc�����N�P!��C�+�8L�h]����(�)�F�"a�:��t,Vu���1Ï#y[L�S��M�N��,��쎳9��%Թ&Uƈ���H�<���q�!|QX�3�N�����|0��38�@fF�)RK��H��'	�``r�Z1 �(1���`͚���B�,�%S��S�v�Tc�L�/>(��%�� x���eʐȂC���TmD���x�A� �J(u��'���O�BEƎ�X �$��r�E3!�X���0�%�M
xs��ڑE��m��o�>!p@ۂNў�tl���$�n�,�����$�.Y�h��<���ޑ~�|I2�"PH�2��Kƥ(���O�q�!ݝ@N���/_ *�>���Oil��1� ;�a~���!��!��;����U��;_s��A��0�F�5�>=8�[?%��Ϟ8����O.�X��"MT�A�hD�[N�p�C�'�*�hr旇A�:��raĹl��X�pe(Tk.H��v��2�E�=�P�5���+]�E��k�Q�2�[�|yaxboZ�kZ<@Ҧ�v ޟ]�6�Q>?�B����@>Z�YV+Z��yRJޡRm&i$ğ;��e0p��1��$Ȉ>tZ=�P@�
f�R�k$
Md�O2\4���]s���9����r�� �'(�Q�%���]�������a��lyע�']� �㵨���1�Jȗ��g�O�<�aᏠ����'ʨ2����I g�:��Ab�V� �Щe0mXQ	̖�p�ɕU=�� �SF؞hR�M�Z."�Q��׿kNɻG�;�ش����F�t�f�~��yBYw6��t��9bJ�`����7���+�'�h�؀��B!8e �.�*�Y��'ٸm
DB��b`��Z�f���;ҧ'*Q(���Q�H��e�e��N���bÂH�� �?-\���O� )3$�رd�(3͠s�j���D��f)QԊܓL���'�N�:��}2�?8�Z�!V  2sh+2oG���kp��+B�<y��4!�,`��TH����7���� �x�}0AK�}ў�)AB�15H�� ��u�\��˃�'�� 4ږ#�"�"��'׽�<+QL�cH<9��� _>}B�x�2}�l���E�%.�����d�v��E�U(U#�;��Q�R��c���=�!M<+L���'�b�[քD؞$����AH�iZ�iC�E�� ".yX�h�����_�V*��'Dh��.[~�P� � �
H�������w|�����"�Rap�"�ZuH#J/D�܊F N4.϶I�Ն��i���Õċ�n�dۢ�[Xf���/��^O��҆��6��	>����S>Y�x ��� M՞�y��I��hO�%�ďV��R�$�7#l��BbX�L�z�h��.]HQ�&M0YI"�#҃Zd�<ɂ%D�k�0�'ʰ#}���rb昪� �r&>��CG&]��D){\%a��T2`@�5 �-qh�`�q%1��$�'탕{���m=Q���������@ݽn��j�'˴@�$��O�y�
�7 ��2���K��AȔa_71��T���΃��Ƀ?meZU��� Y�u���bMV�����-\U�T0� NIa~B��&�	+R�ɼ4�6�1�&��Y�����C������A"lY��05�pɽ6�4�I�h�OE0u�4gX-~����8v����$�Mw����MQ0o7���Pg�~�s�Y&K�ɠA�Y+co"�S�+�?e�� $Ҕ��O?���|Ν�����,�R��1��-<��Č/��q9�"�Xd�Q�#%��� C�!�, �%ʀ�A�v%h����}9��чnp��$�E�i�e�fm���R��-*�epA��4cCg���fA�L|Γ)n٪©�EBy��G��Yeq�3b�a*�m"�O@q��g-d�`�r�|r�`���+?F���R�Ȇ�M����n�?9�lN�3�^�{�	_\������_�r":}�
�֙��G�OF|�v`�*u�d���ʲ��4���{�(j `�8�8�1���p>��D�*޽�$iT�%��񃦚�'�@=	�GC�t�2M
��I"b��?�� ���Hs��!�n'N��4�b"Oj�YD�� �`2�
�R �!�'vD�H���$7��P.� Hz�yd�����Â�V'Ҝ��[?��\�ȓ$�p�F)�2W�tm���ָ�v�4j��)[�ֵ�~�S!̗a���I0h@\7���y�@��ƚ64�8�F��q�S�'j��D�䌛�Tͮ@+���h���"bJ����Q��J5q�T����,�0>��3Ŏ��F���f��L ,e�`#�kV�p�Np��ƙ�?a�p�W�.�� �O�t}[�dY�@�A��5=t��Rߓ(Dq�3��>����� :���0H�I��f����j�ቢv����*�,f20���j�O��X!`��.���c�@G�օ���;8�%���ɀx*��@a�Լ5���g�M	#� t��b��N�� ~�ؐ �^>�Gx%U������o��Xs GWF	j��.�Ic�O�a@T�U�n �3�ϳ?�@9SGH�R�\X�@8B��(ӓH�s8�P����3A"yҢ�V�Dn��d��OL�	c��&��8�H�C��On�XT��9���&8���t�M��|CH3]!a|��C��l���jJ:f�{5��,&�؉��E� �G�`�!g�����#-�^H��yB��$�>;V�ٟ?����S@0X��MC�b$�0�>�wt�n��`	�Q�7��S}�y��#��LhuO���%��7U
�0Ђ��oe,��׭���ft[�-� (@��Ų'������k<���I/%��IF���.���o�$$��g�=@�]�Df�6&C�	�s����Ce��XX�MJF�E�0|�,���Q8�ЬKv�^�O���5�ѕ�jQ�Ю�0V:l0
�'� u�W�߈r���GL���|�a����� qG�<��'�gy2��[x�{����ju!jq��y��J�b��y0M3:��P�\�h���	��O�\#�#lO��A!�ԱX�z��Ƭ�<���'$�)��gξ!����i-ҽ:P���
�L��b�.*�����'���P�b�{���җ��,/�ő�{B(֖��T�GDċ��>]IGh�/Ip:��%Dq|��w�-D���$A� D�1r�K�8�pH���N�Q@ Z��l���DɩIG�M�r�H�i@:03�P��!������j]:�Q:ǧ�6b��
)!�����'3�X���޳f���뀈Þc���b�'�P�aG%G%3�Se�!	]М��'��A�A�j�5�Tm�rؖI#�'w� ��s`�Sd��#cj�'l�@�0�����A��0E#
�'�(FY%G��=+2�
�|���Q
�'�`�I���}M`�J�M�z�1)&D�� b`��ȉ(p�V����ߎ�h42�"O �����n�qo�H��y`@"O�DB�fǧ�T�)�.WA�Xis"O ���U��Jݓ��
~DI�"O^��:��лC�08���"ONb���10�r��5n���ab"O��y��!g�nd����z�
q"O<�)��X��L�W�G"r����"OT��g>#1&�{W�Fd�1�"O�I��nE�i�������=�A`�"O���@�W����3\���Qs"O��Bc�1n��0��
x�2�"Op�d�Y'/�p��N�*>�����"Od+��c#ߡCϨ�q�j]!�](4�`��pF��2� =���W]!��'Q�ȣkC-{��H�"D�!��M�,
|| ��O>�e���7�!�d��-�d�$HԛB!b�צX��!���^CJ��u+U4
�-�t�.Q�!�P7JD������a�ٌ^�!�d�r�I1�ح&���r�� 0)�!�$S�6ư��P�
(`��ip!�ޡ!�ټE~�!���	~ö��EG�`]!�䙺HwB�;%�M��ơ҈&k'!�dтV�b<h'$6y���� k!��ޯ��Yb��%s�M�K\�	�!��
.C�B�k�(��01B2�D9!��X�&-��!�������,�=?.!�D�>>��xᤈ$~����+P�t
!��>�k��X�S$ԂT̗�!�$	�"��\y`��s0J-���8$!���A�pH+1·$)�d	Q�X �!�M�0,���EnA�5a��MV�!�$��F$�I@Jj��CVfLz�!�Ā7�^E8F�|i�1��Le!�$R�#t��C�"����ac���q�!��JqZ����:�%�M#�!�DN��J��s��+s�f�s�,$~p!�䃂8���0r�q��5iJ�`f!��}���s3k9D0��8ǊT�!���F����vK)>�rt��&�!�D��<��<a� O��0	�LBT�!��2I�yg�<5��yh d�.|�!�E�JO�Uh��� i�V�[�!�D�n�"pCp�6qdV��q�b�!�
8� ��.�C���'(d�!�DR>Mcp��dk@�[:2$��g*�!򤅘Q�dMHC�z��0�+Q=:{��������$͙�Fr�Y��	���A0-2���8u�1H�V�&�P��u�!S֭ـ8M���ʀ`�@���QP����v$�􂇸{�����\��D�R6�A��,�(��ȓ>�@R8 |%�T��Q�$q��cg�M�4��� ;�)� CR���Ɇ�锡`�H�"�4W�[|X��"J�Z`A�0+%�R�i[+����ȓYi� �	@��ԎL�<�,��ȓ^Ԑ횇�͠�5��@G7Ype���ԝ�VjR��qk�!E�"nЅ�U����,R:x�2�ô�Ɔ"Q�M��4��-�U!�$.EV��O(����pI�F�Ͼ�(A�(I-���ȓ��Pa&)�$Y�!䄊*e�FH��S�? �E�*���i��էP���{�"O�r�b^�I���s���=T�4�;�"O���CS�����e��}�n�q�"O@�7؆���j�P�jhAz4O�e�1�L-Ƹ�������A��zy���V>P::!"Od;�V�+�6%�&-S*A����^������5N�T ��ɓ85B����� �f���E
���2 0@rƨk�zM*4�1L-��H�$���'��9�"���=��m� 7H�0��D��h�EA���O�4�Z�n7b���#"ƓyֈD��'( ��MM�8�X��,]Pn�xشbж�I�ǖ�?g�ӧ����dۆV�����2��YQ���y"$��Y�,�Z��A5a��s����d�#U�5[���
��<1VnG9�����A,�
�r�vX�xE�U<j���Ṅ29����E^jtEԇ�!Z�񄔚b�<��.o��c�*L�,���l!5
L2kv���	3t��Q����A���rS�L�V�!�$�)��xP/S5D��R�O�wɛF�W �U����@��s� ��P$�?�>��HɀG�,8D"O⍚7�T��͊�g^�V�t��W���l�&;�����'�f��᫁8cS@(��L��!7�H�	�Adp���V�u8�1Q��]�A�>-H� %:L`PQ3�>$���a!�$������ɝ,+�,����f�Yb�x�ɏl�q"�S�)��:��ɘ��A�tT,__^��DE�3�ɫPi�(����^���[����R Iy7�d�+����{�����(�蔊��Ȉu�~ŠQ�"M$����1C �G�B8���I<jZ���$E�X��R Q�!�$�dr<��@R�B��Ö́"⦩;!�GsyB�?1���}&�,�$h�!1mL4�T*�vz��V"9�`:D� �R�3��X4��� ���ZȄ�h��9V\�M��ɠ�H��� �
	8��A�Mƒ��$T�\�@@J�`�`2�
_J�
3$�	G�i�̈́H�q�' I��	T�S�O<�Rv�	Ad̬�PP�=�
��I��q���.w�%�u�G�O��{�C����&�
7Rj�qN<4�k����p��1j��F�()\�z@(��-�LQ�꟢d�剡*T���E��I?�.�N�[���왁BW�r4�9�#��� y��>�O�Qp@�Q�f�hA�ߏl5�[���� �D �.�W�O6m95Dxɧ�[@��I�
��t��)��q�p�c��ҷx4�r7�'�p�@�ě$m�ld�.0�-�"и�aFؘQRF��QK° ��9��(l��)U���&�	oR� s,�hⓅy������V�V3c�FZ �OT#C��X"��A�IU)�10nx��!ł��M�� �#z��H�<�4���
�5��y���A�  b2���'f� C~���q�B�6%�(O�	CR'����i�4d��<�kH~���<Ĉxp�\ g*�l5��Bm����ʂ��-H��/�O<H�b�P,C,����H%iN��K�&+��"AdB�9M�L�FĞ� �<@���.I8��	�oF��wZ�Ċv	XL�L�����wxQ�0_�����֗����W%��R_,Mx	�*cvUA��Z�z_tm)Ӈa����'�N��ҋ�(-��O�~]�W�_	2�aфG�R݆����|/Ќ$��+pP]K�fK��u��q� �@�E�C�. �d��9� �O�%��'��$>c��Xrc�6ˠ4(�A�\�9���<�F�P�
8�K�g՘#��0�-��Ij��g�I�`�u���y��`��P |���AQMV_��T�5�.J�@���j��r�h��GP]y\���O�3���4���O�D�Ҡ���p��~
��#�� %Ǻ9Y���ob���	{���Գ,�)IP�Q�dQ��F<"�B)۱Xr�X�)kqO.�N|rD���Ua0��+!�*���:O<�S%�=@����D��.n��lZ�%�,�y���8A2�OB�6��C�8R9���s�8<9/�w�0�'��yhRD޼"�Q2���E�>����1H����&s�ԉs�O4D����˜�N�t$�m�s�P���>��u���#��L��~R	O (���C�D�t&��q�g��y�)U1\&�'\�m��u�7��?ё���*}�]�&�<lO"��B��0.;&����but ��'�x9j��*W*�lZ�z�1#��;h�6��P �m|�B䉈}X6	1� )��ƯڔpBV�P�B����x"�S�Z�l35b����qb��C�)� N	q�V'.�~�QqJ�7{�.5VȔ�"ba�"�'��s��c&a��<��E(ϒ�G�\ ���$D�x��.��$�ӏ�7j"�ٶ��p��dI���q#.<O��z�EM�$+4hg������'j8���~�8��Hҵ`���L�G[��O���R�1&�&�2W�F�V�ЈO����d�#�(�"��Dc^0n���80�ذ
���� ����@c�.��
ۓn�p�v���*"���q	|�i�6O�A��eȔ�x	<}J|�@�$m��z���3��݈�Qg4�R��nB!�� �@p�`���?`����[5��*|����-a�` �e�N�~�'�f� ���GE�	?k����2ֈ���ٌnKV��:���	�Jv��)S�+Լ��1�ȜU��IA�>y���O��:�m�Ê�
��� ��AE��:Y��
��3Q"q�(p��aǬ(�|�I�J�O��r��ObQFkN1Pxh�ӓ�xA�e��K���@DHŠ�`a̓[C䌂ꋏG�Pҧ����~��E���\RV����a1�� �L `�L�0"Oj��+�l��)N�\�M�%�>yӏ��3 �t�p�ί_Nf���B#}Q?Ys�MT�W=dl(�E	8������"D� �f�/�����%A:�,B���zd�؂���J�Zҧ���ǺY��$9���P�uP�.
<�y�B� >��`��n��_>�p����~bFt���aǓf��K��=~Ozh3� ��	��t�R�;�O�����c��������Q���YE��'��EQ!m�<�3o�R�P8�m��X��I1P�/<�ri;�'�21����T�'��P�x����3)�
�J! W[>'�a~�m��H�@�+w��O��\X����H���0�"J�C��E���n\<��I�|�$��q��.45.!�"���w��=9����
�rB�+�I��H��F���to�W� ��F^D8�(3����y��
+��h8r�^2E�
��ף��?�Bʊ�&=�c�y5>Pq!K
�h�����Z7��!��p��M ��%D���vB��}�,ъ� �6d@��DF�:n+�P�G�R,K�X#�D�@a:�'�O����ݳ6m��X�;x~l�U�'|fѕ� (?�v\R!$ěh,�D����U�
�q>*�(�b�7&�S�aKH��Wȇ�R:(��J�hG{����%�QL������ӆ/��	�_&lP����b+^��h���!����^(��<sD\����6h��l*��s��D5z��AӶ͑���>-�#a���RR��n>�S"�Z�<q�g�V�X���W;]�XHkСtz�[U�U,a�v��5Hŵ�O����dMjzH���G!V" a O-�O� ��'i���8�XL "a���x���12 i�	E��p>����-hj���0�2U.�:Q�W�'ZВ�f�ϟ48s�ҮT�ӅJ�F9Ж��A7�I�gΎ�HvB�	���04
�uj�� ^5��{��A
�}E�d��<f��m�F�p�j� 7��
�y2 ?�0�����?e��!� �I��a�Sk
���>�p�d�`�W�NBt@��i�b�∇�q��l�����UaA�U��	g̎��>5ـk�a{r$R�>8$��'Ĥ}r�r��W��p=q��Y�HD�զא�M�VCD��	��s'F0��
f�<I -B��f��
f�Yx��N�2�"��2�F�Fr}����<"����J1sa���_r�!�$D=EY$�"���(�ҳ���V�+T��-G��'ft@F�,O$,��
.rb Iu�3'���#"O`���mZ�A���VlW�v��	�3�)޲U{�/�n�|��ɗG�|c�KY�,L8�XӅ[/l���dM5�\�v�$[7��U8-ƬXͦ�z�j��5wjB�	�[� ���ZNZ=�R��w�*�@9�@�@�Z E�W�O"T�si��{�������@��% �'�\�.4:��)�b��hP�5��j��^�xP�s�>a��>qB�}�H��CbO�x���E�m�<q�Ԁv�lD���7;�2�)C��x���.��}���)L�d�� �\�,�BL)���W�NC�IE7)�vk�i�*��㇨O~>C�ID��������T���i��G.(kC�)� ��JS�W)�PQK�Y�"O\yEC 2�<����@�[B"OZě�f��OT(NO�;��l(�"O�R����v�8�㵣��D�B��"O�x�@� M�B*����bD@��"O�� .�A	�!��{���!�*OlТ"�\<w��}Z���h�����'0�%�D�	G�D�04cBd! T2�'�DYp��
/F�d�+PȢ�)�'}p�;�o�6`#�|Cm�]���P�'������L�=i2�""�6�F9	�'�ɪ�"�YɄ�p,s�z��'|-X�
://�ѱ��Ĝ>cpez�'����I�5�����I��*S�4��'��1"A�,T
���1�G%]j�8�'X�)e�1����𭅇^_֝q�'hR�����<�`!��W�DM��'e����Cp�\�{�R�LU4��';t�j䫅�!�`�t�����'���9 e�K����ƛU8�'?�����شW�~p�UI!w�d;�'z8e��c��|��e��/;^t���'����e[�.H�e�SF�:ި	��'kJ��Q B�z��񭒄 ��,�'̒�4b�D�t����z��	�'K`m��Ϟ�V%��hG6"�<�'��q��� \�n���l�S����'�
��M&>��%���]�Ț
�'f#�ԧ&i8��"V�p����	�')<|+�#��b�@AL<$r"���7BB�*B��zO���F�9q[�X�ȓ,{��+��_�is��F�-m� ��bYJ���"Y7@Pj@ lG���ȓh��)	ʃo�ݓ��ttx}���̱�q�ͅE�IK�����ȓ]� �r��-~�d�w�Θ1V:���m�D�+Ui��.L���f�C�R��ȓk����eT�/ޖ�k� �4�:��ȓ!(ȂD��O�N�A�_#A�*���_���$�O�֬	�HR�(M��+:���'�0*���;eń����aN��B�7+7"���(L�?"n%�@J���ا�O��2�]7�v̛���c����'逼A�C�,-&ɧ��L���(u�)��
��r9�<)��>;����%�Pe9G'���X�((Ů���z\�S��-l�5 �R툜�O,܄ᓴxޢX#�"H#�0tzO�+\�DL���u��W�^��}rN|�K�)Hm&\�A)Y	t�j]T�A�	�t�hY	D�R��M0���M�K(�9[@��H�,;�f�.
�`�� ��@b F��6�tX���R
��W�G�R8ap��0�����p$xШ�œ6H�	 	{>�9�FM�^�����M�){��\���H#h� ���ݖ���M��<E�D�J��:U��
�$̞�)��
5�pq�좄B��OFT��Ӊ)3�HP��L6jR0�A�1j�Ƙ�"#τU��ʓ.Ū}�'G�ά�D���țg���7'ytΌZy2O�!~{ܘ S��4_?�1��@��%��y<0��#ƘO���OzdPG#&�)�SU(�i��m�r vă��Igw��o"����G'L'����T�:j�X)�^�!�d�<�PL�"A-�hKf�P��!���N�>����Z��0U'ݿ4l!�dޓu	VyfD+�4 pƟ�%h!��޺!����n C���P:R!���@���IaO�M0�����+8R!�D�653�M`�%�$~-p�`��~;!�$řu����o�� - p{�N+!�B�=C���n�|�������#"+!�� �`
)NM��M��H�%�Na�"Op9���U��}��[$`x��6"O.�3eAؗ>K�%Ju���zG�� "O��	؞����e�4n;�q"O$���Y
U��r�� ,��Yh�"O
�{��H���Q�M��V�"OH�r�/ '$��ɴi�6Y@�v"O�<锠� sPb=���o����"ON�c��$Sx�-�A"Q9���qa"O����Ċ�4��(Q O�y?���"Oz� %e�";��Ѳ�78 Q�"O�L�oa�̀i=�L#6b$\�!���0�6���H�(�y �]M�!�d��u��;$/A!F PD�<+�!�d��~�+��� 	����Dw@!�X�;Z墳��IPu��Ǚ�%!�D��Bܠ� �*�n��sl�A!�D Ft��kݐkB�A�&˂��!�d\�4\X2l�.`��3C�<s�!��+f��u��#�~�(��D�!�d^=Ƽ3f���B���#�^�/�!�dα��+���sâuq�I+�!�$��`z,����[�^��=Y!��)�!�����2+0�Ь��^�7S!�ďL͢iR����܁NI!�$�I��m,b���Ҩ�=	=!�Đ�k`P� �o�X�Ah�#M!�D�9(�����\�Xy��@X�M!��[�M "����\$4l�U�􅖒*1!�$G ��	��OȯBk��P�;$!�$ʷF\��*�K��#fqx��=!�d�Q�4c��.{Z�%afn�=$!��g�z�cq�E��|���͆�2!�D�4U�0yIUH=�H)�uc=r�!�d�0e�P���n�">�ҍ�hP;F�!��P�h�%F�G����eh\�Gq��$ʷW�茒����M�`O�6�y� N�?��$Ӈ�3D��!�ehO��yR��k<V4IRDǣ":�3u���y��B�,y+@�Ps
�P���!�g��VB�T���c�}!�d�1>�,���D�Y�� �Eˮ@!��Čt�I��	!�d���%�;!�䈐V���3IF�$|$��#Ε!�P�s�l��gY�*f9K ��7!�$�:���q�N�~��r�-�K�!�
K�MB�FR3q�N)�e,xd!��	cܸ�S`�2Z��(ru�οc!�DY.��x*c@�5!� �Y�,C0)K!��B<F%���"�ʙ�U���JE!�\�,��p��"9��4C���:y5!��ư�U��M_��D��a���Py 48"0hQ�LZ�~m`�T�yҨ�/u��I���OFx����yboD�?�F���H�&=�v�;PI��y"�E�I�l���"G:�LQ�����y2�H����Z5�?9���؅ �3�yb9
�8�)&DӬHL�a�C���y��ήW��M3� A�<��mM>�y�ўD�P�Ь45f<a1�]��y+0"���$�	�3mt9���8�y�'�n�!�9_+l耵�8�y$ڎ�xp:*
M� �ڤN��yb�PV?��kD� C�ڠ��	��y
� �q�&�8,T-qpl� R{����"O8q2�I�Z{�l��n��ɫ�"O`�hI��@�,�2艛w�"��"O��Rq��^
�t��D�Kk (`�"O�0�fd|(�)�I̢F���"On�Cщ�.���r�=fy�h�"O~H��h��b5$߄[e��i�"On�e ��I\�-��(	�,�F"O��r�%-RT�!��~D�q҄"O~�2�f_�?A����G҈Z�7"O.d�Ή'�\I�p�ϦN�A �"O�i����-��"�H��)LH��e"Ol-aw�P6_	�Yh�F *~Sr]��"O" �V�Z�p��T2 &9`�"On��삛t�����D�MuLMBq"O�`)𪅬]Q���/��L_�A "OT�X���Ze8�W�@�w�XX�"Oa!�gG�L�@9�� Y�(!�"O���*ʈr��C��L*�F��p"O�q������Ү����d"O�Y���n9jí�`Y�"O��J�C�*(��!�":ڎ��E"O`����R� ��p/ɐH�&��"O
��2��F¢�U��;�Ҕ�f"O�L*�
��g0��M�M���"O�����#c����c��b�5"O�� R	���&0����!����"O��:r�;p���1Q왉z�d�Q�"O���0�Ɠ.v��I�#��;U"O��3g�?�VA:"��.3����4"O\�UC��5-��cV�Z�ƨ�"O�S�✎U��P�مo�0��"OX)��'�86j0�"���9�d��"O���/])S���P�@��r$��"O�Hr�(�@����m�?KL�!"Ozq[6n���@Aw*��)и�!"OZV�Y�Z�� �B����"O:� ǋȡQR�Y ��X��"O��q��J�O0�@y�d���Y<�yR�v� �Td��{�Vy�5���y�F�3<��`ȎF������yB�u9���s��8�ir�g�0�y����?�M�͖4�ʩ 4G���y2"��YĒ�:�(O&)����T�ט�y�˥p��CB����~u�f`�9�y2��[��D��+ O��y��;�ybH��Ux&�S��n�x4���y�L���j�����0����(��yR'��Q�]ѣ�đ~yp1��gא�yb�Q"7��"鎤	�
Qx3����y���g��9�!"H .���Ac�y�"%>��q���1ɒpɡ�� �y2G�4;�%�dK݌(��k�:�y"@O=$<*ŋ%L�4�e,���yr�6	<��	���+0�8�#��;�yrMՈ,�u]/#��X-B9�y"%L�yv���Ch_�d٤͟�y��L7o8R`�!Cбe�z�4k���y,�N�|� ��>e�x�yC.�yr���c������g�I�C/\��yb�ǡN�rM�4'�R���5��(�y��N�����FFE��i�d���y�M@�
$	��d��Cv�E�T6�yR��(Xp��]*?h����+�y
� �˃*�&�e��(Q	Y��h "O�}�B��<{Ҫ�*�'	7�p�Z5"O"��o�1~���� HkʬC"O�]��ݝ\�"M{S�R�t]�� "Ot����j?xM�ʕ.3A|Q��"O��&j�"K��©[�K9�x��"O&EH��P?S��4H�B�&�^]�W"O,��m�5Pr"�
3AQ�\�F`!6"O�$�ƩsӠ��Ǡħ]f��	'"O|��T/3FƁ�C@�1&c���"O�a��ͧA	�ȶ&E����"Oj���H�(}�b��BRR�؂�"O����j6>z����Q.�v886"OĥE�9[����Z������"OB�!P�C�\�t̓����"�[g"O��
7�U�@⮨bP�L;l� +�"O9���ݳO����1�߄im,�u"O�����qڸr��
0l`�@�"O���`�ۚo^��J-ɛ �H���"O�|{��/����Vk��J���[V"O����僮�pA+�lh ��"O� ��菈GԸ��dʁ��F3�"O96�7RN�Z�	�E��|��"OFD�s�ιXݘ����H6�dP�"O�A�(��Jg|�JB��'늬{d"O5��	`����%���p`S�"O6ͺ�O73����l�}�B�X�"O$t��#�* �Q���!w���C"O&) �al@b G)u�P$z�"Ob��$,��N��Z�nS�\�D-t"Od�ć$!b��R�K4���"OL�����,M�"-
�h����"Op���Jߘ\7�k��ɴYZ@��"O@5Y�)�b�B [��*�j��"O��ʂ�ޞ[��pU�y�`:B"O�s�'�'��� �����@�"O<��t�\�0��\˕+L�
� �@�"Oj\*Wo��r��#@�?H�"O�5���`v>������`M���&"Oؘ��mǱS�$i�OD	Fn�v"O��ҮJ�2(5�.�)-"�Xe"O�ԑ��RA�JPx$��.��&"Ojar���q"C"��`0��b�"Ou�sF%���n�"5C��p"O��K���PzQ[Ƿ�N<x�
h�<y��.b�Z�y�,۶���S#�c�<R�O$R@DЀaM�ܰK���K�<��Ɔ�R��9:r�K�^�C�.�l�<��`��B>Y���M�6iTh�I�i�<䉖<@X�k�oPL�H�8��e�<�΅;_>&){筛�_x�`�K�d�<����E�ҐH�̈́89jUh6�
Y�<��S�&?�T@R.U����Cn�S�<	I��H��0! P�4�����e�<�-�0٣����ܳ���J�<�-�5>'0<���5xV���,m�<�B�]C���b-E�l�|ԓbC�<�D���ؚ�^V���HW�<1! �u$f����I&XB�#r��U�<���V$ @  �P   �	  >  �  R   �&  2/  t5  �;  B  TH  �N  �T  3[  ya  �g  �m  ?t  �z  ��   `� u�	����Zv)C�'ll\�0�Ez+�D:�Dl��F>O$���'h4�l��n�p�2���cZ��
J<�v'�l�6�H��́M ���n�SA��?�/��?��A�d=��pD͜�-��;`Z�"оI5HN/`z� �Pf��S�c.�#�uBի*����'4t� ᢇ�X�~�i����ε�fߗG�����-�OD����I�������$��۟p��ҟ�������S$Q�#�h�ч�$�!Ď����	� �Ly�4���O����D�D�Or�@�/�U��c �	�8=t�ca��O�ܣ"�<�������u�u�	�<���\#*�3aE��!��b2��.��p��yR�ϥX%��[��C� ��U(q�����>��~R��j��p�O(\�[�F@f
�V���܈T)���?Q���?���?����?i/�D�]�a��Ms6+��_�z9a�c\�oF�����%rٴb�6��>i��i5�f,�Mkr����?�#$՛*�򩂦I�kx��м-g���f��"�Mз%G%4V�8�C	X�t�(2HD�}�p6�IͦY�4�Z������'��	�n���04)��k�v/��ԛ��Z3�:�kRn�(A����� ����7$b�-�� �2z�\8�ʆ*+A\��O>����#%B�X��'�i���$G8џH�	ܟ\�|Z�
L2=V@��j��i���Ouy�)§n��)b���y�~(*P�I�dS-;���hOF�d�[��o�s����� ��5��#���{b��;�?�)O����O���5���1�E��8�^���OX���Q��xȦ��7<�n��*O��%�/M�t-u�9U#��D�H��<��G����k2�l]�	�5M�	韠-O�$����!p����"	Z9(T�'n2�'��O1�:�I">����nY�EL2Ijq�J5oJ��E{�O� 7m׹mҰ���C�G��Ԛ�H0ey�o�Z�zH�؊��O[^�5��W��13��%>2FUق"O$���dT�j���C
ҷ~�|A'"OΡ2hO��p��W�F�(����"O6$�sMJ�)�MjnRXDJI�R"O��s-S3��i�G+�0�aU"OD�z�gF�y� ��j+*��԰%�'���a���S��V�c��(Z��6��'���ȓ#�T�D�5Ȏ��ËE�E*�M�ȓ\�t��ħS�t��msUi�!����ȓ-�`�8�
�;;{z�BP䗂�P��ȓ>wEcfA	�8���B�������ȓDe������;��ԹY���'u�i��d��� �ۘJ݌}Q��(G`фȓ�H��Ž}���5�M�P]4|�ȓo|LJ�ǎq-��ɓ�d�r9�ȓ+Z�[vO�&@�`Ap���7���iRlЗM�t�
� 2JL�8Y�͇�7'#̘`�4��D۾#3��(�
��2����\��"R���Iϟ�ϧ]VY��H�UᲈB$�?��E,�|i��L�<y���p�d���0<���Q��}�7!ʹ����A`�A�䘚 z�����S�AR���%��$�Of-n�ϟ�Qb�V?9�� Y�|��YP)Qy��'��OQ>�I��B�X��$��e c� �N%��۟�D�MkӔ5Y����]f�qR��(#z�ؤ-Ҧ�$��:QH۳[�H��?��'[hJ�qV��L�Z�QLƷ��8��'���4/
z7�(i�_�b�\��'Hh��� J#��� %�nI��8�'�M��퇫|�M0�埂e���+�'�ZP #�!�(�xBĆ�[:�h�'%�z4l��Gjʩ5E�X��ײi��'�ޤ s�O���'��X�<
��[�=�<S�!V&Eؼ!�A)>0)b�K�/M�`2��+�f`�O������1"h�jcR�hؙTkF�j�s1f�6VB&I&A@i�jc>�5��Y��$�8� ��� Ȃ"����� �l� 6͒ByB-��?q�����?��c�`�`�V>xq�m81J�-\�)��u�O��Q�>Z@Bx�*ܘ v���'_��gӊ�oZ]�i>��SSyᛑ_�N�x�$� �X��f���x{��dӌ���H�a�a3�X"D-��ҥ(�IZja)sO�R��U"����|�$Y���ގ\�!�DU$r�`��o���cא^�Bv�'�LB�	�*.��%�e>޽R"I,~x!��C1DZ}bR �:~�"ꛢh�'ŀ74��	�7�o�j~ҥ�e�6�����_ ��)tD�?�.Od���O`�d��wJ�"�����J��z�� xC��t����l��~�X��'�� �Db3T;�aJ��3�y"�ΠZ{� a4�A^	VHH��0<��I��`@ش�?��Xl#���#�I�bm�y 0�����?���?���䧥�'i\�s�#�O�<�8%٢w��Q���q���K�
H� \F�fj�S��?�-O�͡��Ӧ�F��i��$Ƃ��(Q�� ��	OP��ɲwa�"<E�Tċ�"����˳(�͈�����W�QE�"|*��H�B���}�ڐYr���s���
�ڭ�I���S�O��"!��	�Z$0��'+$�b�'K|݋���5Ш��2� ,0|���A�OCn���i�1DȰ��Gʤ|�dā�i6�'S"����O9��' "T��04�ȥ@y��0��֊ysL��3Ʉ�����OR��p��Yg�F"��+=�,�rn��~��'N�3������*�6m6Z�"@�e��?"�D�ੁ ,4�%�"�ݮl��m�8�ć0dY���*�<a�h�h�eEO$`�.䃰�նd�T}��D#��?�u� �P	���ת� ��(�3�?Y�� R�	ey�X>��	zyB� 0F&�A���rl�R&�P�N!d��r�����O���<�+�F�D�(R�S�Ζ^X����?%�LRk<U����ɬb�z���L"p ��i�͖>�ٸ'�M��K�ǔ#���	x)�.ݚs'�@Ȣ�ښ&��xC��O��m���'��	�yE��:�`(\~��:v̆�R(��D6���O*��(c�$�%�ܟ%[Q�`�D<?� ��㢱<Q�l��'�ɿ$@{ش�?a�'�&�iB��3ߪxȐJ�7�0pHÓ!9DDxB*�B4��G,���}�r���0<AR	e�'��i�-ś|N���*����l-�4��7��F2�2HZ�o�e����d�t��c��� �RkjXc�K�2P��Ɋ�?��K� pBVdٱ��iҤ9���l�ɛr*v۴������O��1��RWx|�愗5%��=�W��O���E#_ ��O���%�S<Ф��+�l��FX�yPv��'��@c&�*9�rTQ��K�d�>��C�M� �(��a"��8p��X�g%?u��˟�ٴ��:�If>�	���?s�!(f�A�r��(�$<O~���O.�x���i�E75X�Mbr-�52p�E{"�'�����df>�؆L�@"MQ���?.5(��6�̦���Ay�K�3�t�'��'��F���!�H7ʨ+��12dH�O����J^TQ� $c�'7�����#j&fH�g��r������+�P��5�h�����h�DZ1�1Of��D.�9� ����$B�f�#�'R6m�O�i�D(�O�b>��?�7�I?WR����ʆ@�@������hO|�=q���&]���/L���Bv��-oX6<��?9�U�|�'��O��I y��G�	FC���]�>��U�u.P#�M���?)���D&�ɒ:E����Ƹ	�(@#Wii�e��$�^;���I+mNL��e��'C�1%���f6���J�nԼ᪇"Ii��l�˓ݨ�"C�� Iؽˀ��$z��3L����Ƀ�M����$�O.��c6�]6 V�����0n5x�iu&�ןF{2�'���V�x���1�P�pIH�2ԠN.\����ڪO@ʓT������i�5O���`��]7*)6|H'�'@����П@aDT$\�!KE�ƙ;v��JQ(��9�G��KJ|P�n��0<� /C�:R�Y�FϢ@:�L�T�i��)��.������RE�l��ej�uȤ��	<�M����?����]aW��F ��E�?a���?��?�J~Ҍy��;iK�㱇�/ݞ$*o���'�ў�+�?BG�	�hlpv�ƒn�X�/���$�<��D
?|�F���4�6m�O4��E��3���
T��!Z!	�O��D�ZCP<A��T���,��f�O��?�+�"\"u����&�R��"u�3�S~�I׼P��rA9Ŵ(g;ҧ"d�#�Qv��IĻ|u��'8��`�� ���C`Ӿ�d#�'H���c�#�R�����A+9�ԩ$���I៰D{�O3�<��AA�y�Z�t�$�d��D�OX l��ML>i����5>�a��L�yp��`�9�B)X�3��O��Q/��H��[���`�腝E[PB䉦ev� �
ή���;�.#@��B�7p�`�����N)���s,3Y�B�I�t:�Q`DGT�@Ӥ�kn�]$B�	�Wy.52W�$]���sI�4�C�I�w>]��>u��d��״˓MC)��*`���iW.�:s$���Q�0B��C�)� �8 f�܁$�~(���-<�E�B"O��7-@�L��Cg���!8� &"O���A�zx4P��#W0֋h�<�� Mz��Q�W���kQF�gx� �������@��+� J@	V��zk2D��pU��o�ƕ�e�xS�5�P�#T�`C@E]�P����>���9�"O��)�EߥVD&9X�ŉf#x4H�"O
��䉊hcry�g�	'����"Oh$�����=�,��*�|ݼ�!�I�e�ƣ~ʃ�ߟ|���b�-,A5JQ{���I�<����:%&^ՐrC�+� )��BA�<q7�
�'x�شř�1��̚��s�<a�� 5]���*	
@��r��p�<Y�FWd�|#P�аg3��A�.�W�<q H�{[*�١c1%:$b$��|CXH#<E��B�y�*lqU��w�������.�!���6Ő��Ua�*M��9�炘/f!�	�X �Y#�mƭ%'@��id!��3Eƨ� �Ƥ��2�䝈ib!�D�[f��3F���:y!u���j1!�D�R�2�,��q�(mpQ��j��	[�8��$��1H��L`�x!Cf%Z^�!�d	4�
���w{�A3���t!�$Y՛⋞	I������q!��ؗ7W��a�"��]b���m��N�!�D�.u��L�bꚭkTI�t+�$��}��R��~�C:�d$S^,qv �%�S��y�-O ~����b$�
:!|�2o�0�y�Η�I��q��	5�J�Z!M��y�� �Bhx�b�+/��`�O�#�y� �?9�z�aŎ�>$|���庐��'��`Q��'ڬ��B�C�S������G�F�Q?%�$*���h� �?F9*�b'5D�0� ��K�	!�+&t� BD2D��3�Q~��a��O�8��jT"2D��K�.�+�6$�l�&~ฐ`�=D���gl��R��x�֮7�@�M-D��#��\��mr��D7`���e)�O��12�)�'P����b*�/o�H$��
Na5�	�'����􂒵<u@�,T��d	��y∖�0d-R*_�_6�U��	���y�[�h���]�R��tS���=�y2	��Q2	��Պ �`��X �y���`�i�%��J��I[E+ˤ��I�9;�|2k]�8�@�9I0+%Dd3e��9�y���D���2H��� ���>�yr���Jy��`	���V�p�@S��y�@]�C^1+�MU�|�p�Q����y��yj�q��f��w�؍����,��>Y1+ S?��	L�Y0
��@�/ՒMl�!��'����@¹�Z�W.��L��	z�'�z�ڳGßK�X�	��Fb���
�'XI�� W9p6�0�c��ge<=#	�'�d(��FB:��@[�
�'�d���A�-r��Ha�g�=��i��D��f�Q?��Gg����u)� J.Bt��Rt�(D�L�1	�,/�x�2Eʉ�Yu�Xb"D�T��תX3�$�
�"�Z\2�4D����FЎ@A4���NY�CU�P'�6D�t{��R|�.uã��H��U��9D�`�򢔗Z��[aX�]<�l����O��R�)�Rn�8B�^�t������ "�'���׮�wV,ts�n͠d������� NР��!P�,�16Ɵ�w� �0"Ol�I� w/ء�P��Z���2�"O<ɫԋ&y�ƁHӣM�DSW"Ov����C+Ήc�ސmw6�7Y����a:�O2��.��p���+�!~S��*�"O�!���>���$Ĝ:8()��"O��'���<���C�\��@��"O��ːm�a%�5��֮qM`���"O���6�3s���d�&Gİ�$�'�:M(�'|Lۂ�ݥ@:n�
����M�c"O��PTbJ40t��a)�:����"O^��U!@ZL��F�:�,3�"O�9�Ŕ,mS���$؈<
�<:�"O��Ѩ �S�έ��DU�C�� �w"O�����Ɖ��C!�� ���I���~"SٴF����p�]t�t5:���c�<�P���e�xK���>��cmF�<�r&�v����A�0�2X��.w�<�Vg_UL:Y3E(����h��s�<i[�Y|L��,E	Az������m�<� ��,="r� ��Q�w�p��Q��0)��8�S�O�V<��Eޤ#�����A� H��a"O��* IY�ĄF��4��\"O)q��X� P�$�/*ي��2"O�Q#ë�I_@	r�o
�$����"O`)�d��r�� ad���؇"O���D�\�v�Ce*��^c�D�V� f�*�O�9��S�BШ��c(�`c"O21��y����#@K8��ep�"Ov���@:<�a1�]3�X�P"O(� ��)�Dkt�=��q��"O&�����P�	��%K��u���'@8�P�'��8�d�.+8L�BeVX0�T9�'�J�9n̠v���-y����	�'���ZB�4��
�ˎ�k�=1
�'Ҥ&�>[E �IM4v\��'��v-&^J�%�w�����)��'5L4"�.bZH�Zl�R�@Ȉ�Ĝ�lrQ?]B���B �GQ��$��$6D���5DC0Ie��U>��b)D� R����G�lE��L���(�&D�X�#��� =��
��I�ʗi%D��bւo��ٳ!�Tl0��E>D�\�%l�Qo
�x�V�1n0�p���OȤ��)�M٪yKS���a��W�@eXX2�'��er!��~������:؂�'~� �g�&5�(�Lތ�r�P�'��(�5gĜ@��=�t z
�q�'C���F� ���4�En[�@�'̕���R-k,�T�0��"xǾ-A*ORL��'	���V�C9��(��K�h`ʀ9	�'g0�� P�9*����cq�ɐ�'��Q��H�T�P�'��_:Z�'����Q�O\�@��i	1M{�	��'#��TmP�wJ�p��֑G��i��8Z���u=�����PA`��(L�o4pC��,D`��7	�����Βt�B䉗)"N�0#��n�6ʢ˺=�B�ɯh�A�ӏ��X���R�)
)
B䉇����(�����s�
-�C�ər��c(��_Ɣ"	T�Ab��=Q�I�M�O|�\�f�[�~	��抱yբ}H	�'Rdd�w �[��j��]t<�M��'GfD�tC��1��L	�N�T�\�s��� B@���ҦK�~��gFO�(�I5"O��I�'ֶI� Sq啍0غ8"O�C$"��f�!�ڳ0"4�S��'�|�����~��T�0���2Kb-BDɃ�aV�ȓ�*UD��T�d8�UA/��M��-"�`��|��l��çx��ȓx��Aaӆ���]xt˕,�$l������BB9X�X�	� ��,�\9aS�L/|�C���YP&��'B��
�	#Z`ʆ�ߠrT�� F(&��-���� �D�߾Z$ 	�J�/�6\�ȓ���!cM�"�x�d�M�.(��W5D��?�� h3�K����ȓ'�d�f�D\%��KF���Y̐���I&3n�	3 �*��c�-{�8���y�jB�ɱv7�#B��($7,qUg� O8B�ɼݺU17&���� �F̩@@*B�Ƀ��b�Y��5�޾+4C�G�XT�@'D�O�F�1����fB��=OZU� Aϼ$��qԉ׹M�V�=�� Lz�Ow~��u��	;�l+���|�	@�'��视OiqC���	2$\��'��D���߮U�h�s�=P"O H�&9+��`��	n�R��"O�`tj��^� Ts�Bл��a"OĽx ��5����KIq�����'m0�����M�0�	B�5�@�0M����vx\���DM�� Q�є �ȓaw6l+ӂՍb���%Ι�QM��ȓb8=x�j-^� "� W��Y��2��`Xb��j˲i�R'�&Y��Ɠ�6���M �_�8���_9Z����#�����'6 q�'���z������>��"ʲ�p�H�Ck\�3l�4#��i�'�FQӡ�նJ��|�r��
���s�'��hi�l��J�6(��Ł��d@�'��PY�l�E���1�Z���r�'� )��^�$`�7ό%	=.��
�'x<J�ëHε�'Ó ��9���
,�O�'�$D0�'�%7��s�,�m�$L������m�yB���e��fLͅ���Eu@�?z�gl�8���ȓ\Z���&��/����R�F�J�V��ȓ�
�����8`-�h��.W�B��M�ȓ:�v�2! L�"��[�5,�MP��(��h���� '���aH�&�>��qe���!�$�~����%I�~�d���c�2_u!�;H��A�$&�u�vxX� ߹\l!�R9|�����I�RUXp�_fP!�ɮ��0�iT
h�´2aد1!���v�0����*��U����v+B�X��p?���ـmWL�jCO�XV��!	�R�<�����rg����6kb������!�NpyOF%ld�UReJ\�~�!�D�n�R�H�'ڱ@0K5I �K�!�7 |J\��[-G�
���Kps�{�@O��W�4D��JΟB�E�da@
n��B�0%�X`v"H�po�p�A #3�^C�I4dL��	�2jl���J�X+�C�	G>�8�"�;Va�=' �2E��C�ɭ/��L
��M$���C���L#VB�I*�6��%�1��i� ��<⟜��%�S��3zy�iB'^�S��@P�L�8'	!��T4to��:t^A���F�b&!���' ���[E��rбF,�*C!�� �]8�5�D��G����Y�"O��0�.Y�BXxx�OK����"O\�+��[�،bvȁ�	d4�Q%Z�OT�}�Qk����ʞ�tGXB���#xf���/ṯ���L ȍ�`�,��ȓ&hh��bNzL���b�6�<��1�����;'J�xf	/��0��B����A.׾Q��h�L�[Ly��`NN�x��A�o9<��"�CH�)��7Xt���D)���RB����A2�/ԭ%�!�]4n� i	7> �X"FNǯ6!�d^)u|KY0'm������!�\h
�'�,�����<TA���C�f��	�'v`��兘{M��B��+�(,�ʓh�$1[j�'O�j� WM��\��5�ȓUoIs�k�#QҚ�� ��k4�x�ȓ8`6%;�c�*(�T���7�^u��ז�S`$Z�-~PU��`� �2�ȓE(��7��Q�H��: �>Մ�ۮ�P5��V �kI:_�b�'6�'�ɧ�$�	
�{F�I&�ŭ$ݚ��޵o�!�䗩_P� �H�_հ�;ť�%��O�6�8�Dү��'HPIu��>3Ĺµ!�#�� U�i��g�8��S`]��'@���'D�$Π#mN�3CA�drN��@�V���/GӦ���lB���I�<)2��znz�	�ȟk�\����Rm)0�ZT'&Y�YA��?������yr��.���O����O���!Y���ۄ�C;���mx�F��K�Ob�D�l���$t���*�?7����O��Aэڰ	U�� HN�2z���ڪM�Iҟ*�G������O����z�DB&A�	0��VY2P��	3%���	������O�p��O�扞RX��s��H��`	�Thv�v�KT�ã��	�[�,�Iğ�:t�9���?�'c/pp��ZY<����Ɛ�x����d���y��8�?���vK���O`�	E���s�¨�SX�Z�Z���՚�؝�剺8Ԍ��e��1 �O��X?\����l�ɾ|S�UY@gL$.dd)C�Kn^��ߴ)	� ��'N`�r��?A���?A�'Ӣ,�O���gDX�f�����b�'bɪ���iˆ4���'�	���)�>�e�<TxȠE��3m	+��yJX�!'��r7��@�q�π$�M����?+O.��O~˓���lH��I��D�
�����e� �w�i�X��	���)�O�˧�?I���*_&�"P@��d��  �[՛�Z����Wyr���U��2�N�'
jDC�	s�����3�yb��-w�4m�w��VR�Y��EM$��$;�Oh�a�O�6��PIC�z�6��f"O.!���8�������&A�X��"Ol$!E���,&vI��Bq�Ι�`"OЄ�@�x"�1�
��5��"O�y�4��H�l�v�F�&��$��"Oz��3손3gMrA��%�n9�"O���6��u�m1�`
-���@�"ON�`�H����73, d"O*��ei2�����S/M�b]�"O,򥃇D �l�r��r�����Ԯ15�@"dk��(���b�p4f���B#L�N���&Y�lTlի#�1@��;o;�82�˱N�~횢�wYb�N��#�i#�bV�^Ӯ����8�ٚ2�ޓ�\ �鑦x�};C̨Bp��I�@� \�&*`��0�`�.zH��/]�L}*�O���F�8WPV]�X)��	��{�<q��A���)�J�=��ԙ孟S�<��#v��؂3�Q�#�h�(��M�<!0*ə�tb��
*� 3�YJ�<�ƈ܇f�@��E��11�����|�<YA-�#k�L��&�peLU�Xp�ȓ���:I�X��Sw�N�(v�i��K�(�z�Ĝ+?|4*Ӫ�W����ȓ5�8���!�i5��q0�E�:�d��)|�I�ʋ�U!���G4�씆�4f�X�%�4�]�2���v��ȓk�\K����T4�L�0L�/�Hم�~�C`�4��s�H�!xI��S�? �X(F�ߘa��£R�~W��*�"O���@ P39fx�`\PV�Y�"O\aJ�b���>Y�2�Ӄw3�E��'�̪�`B�:��y�H������'ξ�����j��Ԧ
�wHY��'g�X:��G9Ihp����7jq(�@�'۲HFf4Kz6�)��ڤ
(�j�'�*p�FU/s�<�"(�#+Hle��'N��X�o�\|�"��</
���'�Lxi��U�w�~U����??({�'�,�L�8�x���u��-3�'�1z�$F;i H�HK3?�"(!�'�B�c��F�X|�(`���7���'�h��gЕ�&Mѣ�N� �'���B��d�s	A���
�'xi�!�Q����j�l�:f����'>���gn²&��m�LM�-��y	�'����-Ę<� �c )�9T{(��	�'�Z�ˠ�è]�.���f��Hjz��	�'��4"��K %<@S��ϚN���[�'nة �#G�8���H)H���'+j�Y� ֡_���R�o
�h����'�J|/L�\+&eE2*ZXq��	��y�#�*]NFq�1됣(����&���y��m1�d��A��JL��E�F,�yr����g�,
h<y6�χ�y��U��^��ࣈ� �$}#6���y"��e�Z��֮��,�jB	�2�y��c�L@!&�U�
 �)+RD� �y�!>�F��-����(q�I��yR�*><N��#Լ(t� 셏�y���i�Fd���)sP�{Èɀ�y��T�<c��D�ow@�3�H��y��т"[2�6��8KV(A#H
�y�"S�JL����Q ,��j��y"�
�<���9Tbu'έ�Q��y�FTA�����O�?l��]�1"ݼ�y�Fɺi�(�ƌ�jg���7�y�j̀}PĤ�"K�^uN�a�_��yb�J_c�d�T��	Y�l��ЁS$�yR�}�n����ݜXw���ׂ�ye̎e����s	�C�\�1�һ�y�Dܫ8%Ԑl�P/z�v&�y",��xT�����O�̄ v� +�y"�R#�l��e��Pmx١e�@��y@_��*�!�՟t��{����yB`W�L5d��ƇŪq,¨�pA��y�C7xX�i�fTi5�U8`�[�yb�C6]I�]�
�j����gI��yc�R7RhVaO�]�F�����y��ܚ�B�sk
�[�~��c�yZ���sm\z�.����.1�C�	j���� )�b��칱�͕
ݒC�ɽ}��zd�K(NQ����̑�&C�	&#r��'�C�'�2	
�@C�	�'X~ੵlE�wвu
$�7~8�B�I3tE.-��ϱ
L���C���B�!W�\�1I�?���S��	Wq�B�	5C���K0�1l��AF�U��nB�I�C첩!v�ׄ\��R���B�&��d��\59�j�#���.:�B䉒u `�'�S8ǘu�9�B�ɅW��{IL<h��B��X�B�*`�HZ�5f�"(j�͗|{�B�)� ���C�
��q� �΅�3"O�|��.��"��	A��H�p���'l�}{ J��Mg�\z��7����
�'P*��+��iؑnY�r!:�'�
uy��,�T ;d*�P@�
�'��*�J�[����bC؃L�Vu#	�'����P��2-�Ds"�I
sI�A��'���	p��!eЁ$Ob��Qq�'�2�3�8b�+�ONWa�@
�'u\�!�Nċ.�d9�r�J
�'��Z��]�R�# !�6�*5�	�'� AAP�_ X~��ƽ(>�Հ�'��1��ټV$dA��N�)�'�6�ȵ�Z�A��ȇ�!k�'�[����TM����B%�	�'�А�dA�S
@C�� �Թ�	�'q�Y{Wc_%�vXB�͑l���',�U*�f�'pl��� �`�5��'W0�9'B��1�aH�!��Qj~9�'^r�	��]�$���3�%ŧR��Й�'��(���e���;��جH{��H�'�ē��$T�U���;���
�'{�)���%�褈S`��/~�i�'>t31�^&��@#���'�vp�'r8%�Ҿa����ҋ�)p��`(�'��(b� .%<�����p�Μ
�'�A%�	� %ty����<w�p���'��XᥡŐ ���-M�|IX���'Ȃ��j0d��%�h�$Bqr��'O�y#�F��$��B��#���8�'�b!x���; �T3��{� }��'��9#��*߀�gD�p�
��'��"��9Vv�6,ˊa�>1i�'�,� B�W�("��B�D0S&�C�'��1��&x���S�#Jzi��'"
p�[�*�@�B��-Hxf4��'F��!扂�T �|22��);4db�'�Vu�Cʀ�DrY@��2U�����'���d)�H�<%y��NL���'?�X����;>d P��Jd
���'�`���c@�*��ղ"�G�D��h��' �
#��#A���aD�L#��Z	�'ߎ��g
r�p����>�x�	�'��-�Uj^F��	�)^aG� r�'q>�2teط���3[�}��'4���ʋO.��G�ښN�x((�'�Z��]�#�%�"��*;�u"�'t�h�B��6;(�j��/&����'���,"c��q'@�T�̼8�'	��W�ȗtHH�HG�Z�Jj�e�	�'���;��X�$^Ĝ)��E�1����'����VlD����GEʀ/�|�B�'�XW��Gh��*%��;�\���'^6�@H�����;F�d��'v��Z�� .������P�i�'��Ҕ^�4���R/��A�zԁ�'�&��g�.�c��ԠNf�1�';ɢ�k���z�	�aO�5F���'�`kB���y�v�ǘ�D\�'��6��4��AZ���m�:a)�'�~d�r���Z���w-�l�H���'�����Kv�p�o�8�����'��A��\�i���h���Zڑk�'��1	fǇ4W�txj�aBUKRй	��� ��A�9T� ��JG<Au��0"O2��FϘ;}tj��R�u�h�J�"O�9#�-,f:4��%ڨ#��t��"O��2�ʈ~�Z�{ 䒆P���"O���)p'�9zD"����R"O����X,O�Ψ����,{z���"OU�V�F�"����&-�&Y�"O������q%h("�ۅ�HY("O���r
O�/���!PkJ1�@��"O���(Y����ʃ�ek d� "Ob`�?Ϝu�bΓ!9�iʇ"O�����Q #&l@+!-�
{+N}:"O�t	��V�H%��!�)A�Xm#"O�!�n�2�n�@%*�1�0X�"O�}3S�����ac��.�y��q�<���!76H��kץ^�hdmKf�<a��߶@t�Q�
ß�l� E�i�<A$*ʢ$��y����2�T�k�`Bb�<��٦8��B���8�VQ��l�]�<a�[=<�RɈ���
�d�o�<�s��|�+��6^�!�I T�<Y��7�p�z'�I"3؂8�C��d�<�き�N=F���E_�N��H�OEb�<��.ȢX��0���2u���)U�<a#�ΆF�A��
S��$����H�<����z
��Ǫ����qfa�j�<9���-eG���4�
��`y���r�<!q'N��j�"$eO�(B���4	s�<�o�o�hj���2PGr�Q�%Wh�<Q$mK)�<�+�!ZN�У�HTc�<��*�{�nUh�n�
�z,�Eg�^�<A K ���{g���jXx����B�<��FE�='���	�\s�!PC�F�<����>u���0ץQ0`��pTd�@�<�'�_�2 
�)6���!�v�<��F��a�TQ�u�����1ۀm@~�<�tR�dn��L��`�JTs$nM{�<I�FS�2� ��ͭ{l�u���SK�<Y����X��d�ɧ'��4��`q�<��-����2�mrT�EL��'�d�[��ۑs`�:Ӣ�*Q@���'̼]p#��n���y��C�6��	�'M�Ȼ`�Y��q�����2aX�'�LI���L��1��)�����'�F�;�뙫9��+ "Кh� �Z�'�DAHfIә�@�J�iF�Y�bt{�'x"tb%�߁��X �E�S�p�
�'L��Z�(�
C'hdz���L�v��	�'=�A�EE���@���ML�	�'�09f�շ2�0 �M�{�|u�	�']JL�1j�e>��(r�}IY�L�}�<�o8Vݔi;�f�P���M{�<��F:Ru�$�4"�Jx� �y�<�ECؙ1�Y{b���MB4+��M�<�Ck
�q5�#g.�:F �*$MI�<����0%YTQb#� �foF�<9�`Ɯ$�2���IՐf�.�0"�[B�`W��)�&sf$H�eŭl�4&�@ł$X��ce 'U�����yr�V�n����JO|�	F�L�y�'N7�60�3%�M�zŲV����y�F^9|�^ �$��F@$��5�\��yBMG(#���'ޏv9�h���͸�y�]�������P��T�ڪ�y2�E�=��ݨ�b4T��y
� ,����]�5L<,3�#���k�"O��nǪ?��Q("�К�ґr�"O6��R��)}$ (w! a6"���"O9���]K7Ƙʥ��44��jG"O�<aI�:LT)kg�($"$��p"O5���
4��i�d��4�z�"Oܹ!��ƫAB������z����"O�tô���U�r���y8�xQ�"O|�cSC^�>B��+ �2|p��"O�]�`	��p2�X�pJ��_~Z�`5"O�M˱,� �a�NR23�]ғ"O�h1� �v+<)��MƝs
><�f"O�Tx��ʺj"��R�P�7 �}s�"O¹��H@�`+�)���:W,��c"O��!�e*����戉�-�8�T"O��2��+4x��Z �B�a�(E�"O�҅\�	�( �&I?{�rq�Q"OFl�� �!%�@�:��� �|��"O��#5���"P�B�� `O�0 "O�TI#�TG�leP�	:j��1a�"O4P��%2���9gjķa�Vt�D"O֍h&�S0
EX&�E��qf"O���p�I�*�E1R+���1z"O����>�:1����%���5"O��@f���Zo�9�"	܌C��
�"O^�A��W�RYk�o� �,�0G"Ot��=N��S�L�0-n�0Ip"O ���ZtxQ��
bH©[7"O�xa$ڲ'
&`���8�V�Pg"O��	C�^�\J�	3 �-��K�"O~A�*ٍ'����G٤ ��ѩ�"O͐��Z9K����S�0��"O2͋"�&t�|#��b��y!"OZ�a�<}�.�Y��VNbz'"O\T�VƜ�b�A'���p��"OƱ��e��B�f.�4��S"O�IءfZ!I�^p��E횥�"O�Uصw�$��̝�;��4ZC"O�+��0����2t�0�ha"O"yy�㜲��I�$��x�:�"O�8RÑ4s��8�M�0o�HkB"Op�����^.<���
��y�"Ov���M�1Xp� )p0��"OZ����-:�R���Y�Q�V��"O�Y�#�_r����п|��A!"O��BoRm6,��c���\ڒ*�"O&��g	5� A�h��]�.��5"O`!��̓7ϴ�J��q�
=��"O�슃��`��de��
��ua$"O����#��Ds�O�0���*4"O�*U��!��ʣ@�	`B�8C"OnTK��֪0p���!I�l�B"OI��D�F�x,���&�>ecs"OP�i�n� �Ҹ)B톹e8$:"O��cي'~�{�cͮ>3h�"OA���!Q$����I�T|H��"OVx``̾54Bp��E�3j�`�"O�az��"R��dĚNd8�u"O���)�8��k��ܝ�"O�m�f�\�� jej"z�rȰc"O�= JP�H�(S�1���R�"O�lۀAC73B8���;�r�;�"O���s/�q�,]K��$9��"O��#�#ǻe�9��^W�is"O� v�X��>Y�N4p3E7��dJ�"O:M*V흦x�� ��/��샰"O���$�@L)�/�"2z{�"O�l=1l@kW �H���s"O�l�t��eM�eXA"cx����"O:]Q�eˠgRR[Ǭ�L���{�"O�H��l�Dt�
ׁX��e��"O�xbB��`P�T�ã�,p�"Oz1 �f�����a()i���{�"Od18p��-gx5Z���o�1�u"O�9�7��	�0HA-A�MU���%"O�x˄&M�4�R���*�D��"O�EC@`�$@���F�m�v�+�"O���ʁ�}������2Ǥ�8�"O�lk߱r���f�]�c�DY#p"O `A5� H�k�l���%"O�P&*Ȏ/��2�)Q�^ �U!�"O��ӄk��\PňY*wq��{�"OF���J�]p��W�ѭqb|�K�"O�d���'�*@1��W*A�X�y4"O=�ѳ_�ZE#�Bĸg�Z� �"OT����35����!ڰq�|�� "Oq��H�d�r�+�@V*!���"Oz�tiJ+X��r�g	j����"O�$���<*T0峵�M�A�(�:$"O�U��GX7���z��lE��p�"O��4�J</�����87��tkS"OLUѡHdO<����Be&9�ȓ'�0\��� �r���n�ly��)X�XG)þ2*�����E�KH2��ȓAψp#�C�0�a�ac����|��Mx�b0��k�]!��n�ȓ1zx��J��a�a�&�
�/�Ԩ�ȓ",HC�;XrEH�L�D]���@pX �(��`?<�b�߃1�.Ї�TG\i����#��`D�x�Ňȓj�����G"O���I�+U�X����\\ �'��%�� ަ���s�+F%A	'�DE	�
���ȓ)=6L�d�+|l��F"�p��ȓI���c˟��}����;.�D��$+8����V�["�ۓ
2N�U��+c�nC��j��A�Ů��ٲ�'��1��<F�2!��O)�H��'��=X���<}��Ibp͙�FQ��
�'��$"gj�V����N�Ez�4��'j��	烇��q@�`�+I[ ���'?P�Q�=��¢�Q?I����'�@��2�,>�Ep��Q.~G�P��'��h���� uضʒ�$��'����@T[PH獇*29��P�'�0� -�(,@�t���
�Zo�ܸ�'9�;��_�XСׁSWGb� 
�'	��kE!�j<��f��x)�1��'��aC4�
��>)����p�H��'h�J��^�\�:8��HнC��x�'��:�D�yT�:�d�>?���
�'�tq8B _&��+0�X-�,��'���D����s�ݺ�,<I
�'S<5��4CT��2C�ٝ
��h�'L*��$�S�D����ŠQ#v\��'�(12BNP�8bB)�4,�<QWBDq�'zA�B�N/&�0r�lP�`� \p�'�l1	�~(�X7mŜ��C��� ���f#Y�_NJ�s�n�s*���"O��[�'���`x؅�Hv�^XY7"O�`ғ�зO��h�a$�+S
<��U"O�)ɤ�X e�~!3�!� ~�g"O���"䊞h��=�p�Э(gb"O\��D�"A҅��1d���"OЁQ�J�M ��Ŕ�	_F��"O�IbE��]�81BA�B���"Oҁ�"'�	z���2��.`2h<B�"O>{ �2]�t�a�(��"O�HPjf�|9���!fڼ��"O�H�ϚR�V�9@�Y��ћ�"O|�Q�E�Uc�i�
d���"O.��c�ܚ�(�U)۳wBD��"O�\�A��C���q�&0�ԝ�f"O0�Hp��%
��K���}����"O�ع�BAPeT����~�j�"O>]6gܯ,�51�^�	���:!"O���D��i�fh��X�d�1"O �Bס	�.5)щ���< r"O�S�i8��(�hV�v�5"O6q�4M\�{|f�PRN��"O�m`ej�3l��]�R/�*7��Ԫ�"O��W��#S�X�oP�/o�l��"O���GC,;���%ό!]`Ĕ�"O�q�D�,8�\+Q��"�,�0"O�L��-�%��5�l���y�"O�4�v�N0����l)uֈ��"O,H�Rl\%7�:9�g�L�s2P�[a"Oy���X(�`]��A�.��H�"O�p��.�75L�a���L.5�I��"OѢ��ʾ�~�q&�S=GȎ� �"O��"j6� 5�1hM/	3�}*"O̅rE#��g��H�q�
�j"O<@Q7F�U�����J	)�x�R�"O�$"&�G�up��I�(Ϝp�l�"O��V�Ϡxr1[0�-J��i�t�<)��V�z�t �T��#֖Pb���p�<)V!Q3x6��9kK�g>�(`�H�<1�țߊ9o'�`�:����u!�ނ%#f���`�=�th�r ��'!�$۰#��^]���N�o�E1�"Ot0��2C����Pm��0�� ��"O��
�'��4^���6mS�Ut���"O����E�~�	Ŧ�\�H�"O�H@��0L�Ωa$%ĠS����P"OZ�
W��WA��1k@'�\|�$"O$�Kcgy�YYu�ݟ2���;�"O�X�2c��L V�Y��X@�C"O���4�-(��'GN��d˵"O^��i��.��hե�)}��hڴ"Ofq1�		 ��$��bX�	���1"OjA�"�-���/�"��+0"O�<���C�C�%�b�ɽE~�J�"O���f-%�T`��Q�?L�9B�"Oq�gnW�hO��߬��""O�)�/�9�hkΛG~��"O쌰`�?8 ���n�43���q4"OԔAn��N�>���o�P�D,��"Ol�r��ޏ+�H�7NK$����"O�-����,l.�҇�8j� ����yPvx��kɌ5�``q��.D4�'�� R�Dթ6f���M+s�EA�'Քa0������S�o�:�`���'�RYa�R�3�����Н4+8P)��� ��y�N���B���1_�*�"O=!R� �t��%���L@, ���"O�C��7Q�̐U*��@�R��e"OF����%7��8�"��hl\y
"O��8#�,Ŭ�s�ےC�~�E"OH�y�ɦb�b���J�=2�JU9G"Op�d&Ւ8Df��D��8��E��"O(5{B
����l���/�}�"O��s��L�
�R�@6Ĕt؎�h�"O@�1%�������S7z�`��Q"O��"�+B�L���&��'� I��"O��s���~5V���#�?��P�7"O�w�@D��ЁC8z4,c�"O4T�#.U�k���ҵ�vF̀u"O�u��2xA�0�P�<2њ"O��rbQ"0L�[r�ȐU����e"O�iW� %0RP�d�(��� "ODԻs�5U� ���������"O�m�1C3v���a�:4�F"O�4BG�$��d�s��p�h(��"O� ���P��܀��Z�d��<��"O����6� s� �3?&�v"O������
M󨡢d���?)l��"O 8[���*]7��k���*�,;�"OBy��@�;�n��b⛰k3�С"O�LB��L	7*�[R�E�$�<�١"O4\z��\t�6�"��� ��"Or!;g&y����K�yypA�"Obx�"�3w�E;�J
lZ`�1�"O�Q
S�V�&!�t�@�&�ڹ �"O��8J�.yJXĚSgS#�=Y�"O�{�,^8�آЅ��P&�'"O�I�,�6M�ŀ�D��
���"O�FB��PO�;��C����F"O<�u�Z�x��	�m� lA��"O��RS�
�Y�&lr��ֽ	�@Y9S"O"�a��XZ R�j����"7"O�a���["YĈ��R�m ��"O��A�[ _�qc��+�D/�!��-[*�:�`�A�B����
�]k!�d��$,R�����bP���j_�Q!��
8|�q��Io������Z=6!�/U1�8�CK׳l皕�tgɥ!�UY��Z0v0�%�Iu!������z/ |+vFĲ&D�,�"O����#0Ť<SQE�~-\��V"O�PQ��^�Ƥ��O;.�2�"OI��cE-b���C�(�Q�2"O`\!F�{�`���B��7 �9�"O��;�N�:urm�(�X�Fp;"O�0 ւ��t$���Y�7ɴmQ`"Ov[�k�:hXpy�N[Ol�'"O�4*�O�)+5X$��*ց#�8�"O<q�+��|01�A	��1^q�D"On��5�Y�&*$�n�P�f�A�"O¤Q�ɾpQ$�ȦMԶ|��8T"O���d��QEʁ��M
hyڤ"O��fEO�m�|��`�Teb"��"O�\H�Y"^��11�M+2Q���"O�e
��B�Wm��Ռ�-A��"O態	
>��)��˙�V��\�q"OD�3N�t�����lH�c�"Ot$A`�ťScĀ*Q�Q/j{ C�"OԈp1(3l�.�0�&S�s��b""O� ܥR)�5}��٦��q���h@"O�u�V̌�9��u�#�V2i��I�C"O��6��Pin�!L�.�Z�'"Or�(r�8dG�U�r-�3���{�"O��a̝�a=n�(�&˕t<8P �"O.�z���*u�ܒm�(�(7��l�<Q�
̱qC�%�w��G�h��C�Ok�<�$	^�A��U�L��ԡ�Pr�<��#�(X�h��H���)�Fo�<1�#R9N�Q#����W� (�)�p�<)�E�	@��l��.�!Wm��Vȝn�<A��'R*�C�MI!%��A��f�<qЅ'�"�yC��b4 �^�<qB�i�Bt��*[=1t0#D_]�<Qg�6:|@]�$!�w$f����d�<q��0琥%U�c�D��o_�<Y�O�z��LB$K���d�D��W�<���/_��<#�[,=�m	��w�<yA��4��)�ٻu}(��3�{�<q�Θ�-�N����ޫC��� �p�<���ۤ5���Z4+N(E��]�'ELQ�<Is�Ȥq'f���JÛn�0X2�Þq�<��'��fV�U��MZ�Y�r̐��5T��� (D�P�0� J��Z��bc1D��˒@��q~���������L#D�`$�ÜPy(��ec�92� �%6D�$�Um����H;�!�71ZQ��O3D�D����)|��ЀI�J�����1D�� A/�%7R��c�j�W���	�H*D�t�4� -��
ȥv:45�g;D��ҩK&�P�D���\�h#�;D�h�ub�%�@��LV���R��8D�4�@
$q:�xjl�ex �Hvc+D�|ɠA6f@X#J�6Ĺц,D��r�A�1E;�4���Zw�� �>D�4��kZ�kS��R#OچVhҹ�À.D����l҄iIf�Iq�ęu�V4��-D��ЅO��"�`죰�&���dg)D��*âVSך�Xr"�yrTO)D��h�B!B�T�ꡎӈ	?>]���%D��q������2��.�Xh࣪%D�|F�I�.5���$��*B8���#D�4��c�+�"T�ҩ'9�� �i7D��C����M�^����G#�P#C2D���ց��S���j�$T0%bA@�B1D��*thݔo�\)�-�7I;8i(qi/D���t�*�PG!�?�8�ۂ�.D��z��M$]y���w� �B��-D��p���.M����=�G!)D��C�Ҁ1,d�i�AN= ���$!"D��#�ϵC� 87�&�P��!�=D�|��"��*��A��Ϩy`�x��:D��Ӓ���P#.
�[��[��9O6"=Y �S,

5!�$)TU����r�<Aa"M)B}�a��'ҍ�,A���LT�<���M�&6���Ѐ�\0R$SO�<���@{�>HY0�<ƪ�1Ꮑq�<��`Ԅd*�%�i�d�!"��b�<�4둴`��$�b�?��DĎX�<�B���fj��i�i��7b\�R�<igb�?P訋P��e1�,�R"P�<	ԣS�Dء%�ێ�VԨC�P�<A� 6G�"u���U�&Uؔ�@�<��C1
0�9PUÎ-=������u�<� l�c���e� 2`�40X�E"O�8p�
�&Q��	���
[�x$R�"ON������│C�v�u�0"OBq!Q�p����A��=!"O�@�C	�(7tq8�N�"t�"O��Х�7H�蒒��3(��s"O����.dh<<QĥG�	�M2d"O4H[���ԫ�A�
�@q"O(!�DO�3r�������P(�"O�� �C�I`���4���X�Jd"Ob�I'�\Ŋ�c�R���""O�x� )F�i�ᐍ�0�
d��"O���0F�Gh� u��'�p�"O�4 �gQW$%�
+I�����"O�)���|�Q����,�^�Q"O4!���9���#1��=,f�"O<����v쌘��f�Q^��v"O8����_hڽY��!zߠ���"O�}J��\H�t����E�~=*b*O�M�!cf���E�	�"P�	�'�z�g�*i���*DM̦m\x#	�'i��"�KLӨ�Ѓ�.v�D�#�'P�@r��T����à��3gA�'�X�ؐB\�!T ��V3^�����'\4�Idh�O�n{wM �V�e��'BJ�V��1Q���2gD�&�̰�	�'QT�3��C(݀��#���%!�UI
�'M�|j��I�d�`s�ƿ����
�'�\� �]+�B]��O#�*(��'���kA�_�?O@L葎��"���'�� j�B[�g�8\�V�N	(�֜�'�����e�#J��Qf�ͺ!yx���'�2X�,ܳ��0�%�ݕF���
�'.<�۷���<�f`h���1;�d�`�'K�A�v��,�l��Ǡ�8:�0c
�'�������I$Q*�P$�	�'׆@��DN�U֘�� Һ�a	�'�чŁ�>r�2�d024��'(����ף�E{$�D<n>��'�h���_���Q��� y+@���'!��)�"�t��(�fC6Dj����'�L� ����}m��xG��1>kXy�'O\�6��+o����W�3�q��'Af��A&r�����-�c�~0�'a<1"V(��4������X�`�	�'�b1�u��D�!�'+T��)�
�'��EQ� �TY�UM�2;�81��'P�I��2�KmN�/�6� �'<Hm��K���Ĉ{���o���H�'�<L!�㜀 ~�DN>kD�ܘ�''�����19��ϙ�U<(K�'���k��k:���#I0L_M��'�d�
���7�j86�\Ib�@X�'���Kd�A�oߵu�d9	�'ݒ�(���4Mv����gPoK�-	�'0�!�2L�Z�Z0PD���V8� !�'����o�ؐItFGQ	>�*�'�R<�PB��hC
�`�ҥHIh��'U � �k�:S{�J�Gя	�����'�| ���'�Yc	�uyj���'�:�#Ё��Bh��,Vh^�ѫ	�'�D(�ɜ8Z�p�*��ŕf�:�z	�'�rpB��91Ny9գÅ/��h��'�|=˗���8 .�it�HV��չ��� � �-ɍ $*Tb��!��@"O�(g(��f����91p�iR�"O�|P@bJ^�b��sK�;we��z�"O�\�c��E��5@�珮KG����"Oh���X8/�);"��=><x�A"Ojmң$�o����瞒7��0%"Ot�pĉ�!dv2�X�J�.TZW"Oe�I��S0,J�ǔ��r���"O�u�#)S���Ʀ+N	P"O�h9AD̩�qNɵZ"���f"O��Ԁ��#�Ȝ��P�Z@�"O&�Q�K�3b�����&��$˓"O�MۦL�A3���wj3�0c#"OHqv�B�H��
!�:8��"OPp@��V��=T�:�@ :!�Ra��3� _�`�XMA�& w�!�dģ;����p$ѠBR$+�O8�PyRnF;2�"� 'BB0��ѵ�yR�B%EdU*r��P-n�XSf��y���6�\H�W�լC2���3�^��y��.
A����D�b8IC�%�y��,5S�9�0j�n��=zF`��yA��&t����%de�5H�4�y�!"JebY&�X4a�Z��!�y� �\ E��n6.	���Ӡ�"�y2n�)]��8�ɕ.�z�Z�����y�ڳ[9b%Ib�D�(�x*��N�y�͙m7�L�T��"��X��Ԝ�y⇑�KnZ�Ps[��p
 ���y2 _��<��!@��0t	��y2�H=tK�Ö�����l͒�y���$���Cߛ���1�V��yr�Q�Ц�{C�Ýq)Px�@�<��A����ԁ��b�P}˂EPK�<iīM�{���*�%�?u㦔����Q�<��)WcB��
��z���Y�<�G���Q�,!r�	H=+��^j�<�L.1H��gd��y�֥C#Di�<1��(��y{5c����If�d�<a0F��d8�L��h�N���fG�<��K�5�y���!UȔ8�4ǅ@�<�3/�����(�|XHAC5r�<q��˙|<.��WND�~҄I��je�<�2��9;��)� ��kr��3�Q_�<Y�ǚ<i�L���R)\�����*�W�<���;� AP&6:֕Qק�y�<���]>����J� 0�D��R��j�<i@Oƾ4�nhi�^��H���h�<�ƈ%%���3qKK��-�R`Ae�<��`��`�xXb��&�(qf��I�<q*MTL�	�'��</h��FI�I�<��!T�J�#r��rA�$��m�<Q�fM��z�)��=u����Dg�<1F%�aRx�S��ʵx�Ċ�c�f�<˗�J�"����/qE¹Z��^�<yҀ�;v��8�$F�kn�ъ�$@�<��NةY���q���35��p�D�<qD儂
\��T����5q�M�u�<u����drqo3E�`AMs�<Q��<�Xm�v�ՑH�~1�s�<ɥ��zK���O��(�83mJr�<Q�IU(�( sD����R�4��y�<1�I�-XFzԀ���k9��b�x�<y �Z�L���A�L��f��b׀w�<� �	wG�H�
���;��	1"O��[�jX1QT̨�c��a��!2"O�0�MS+u����&�6Z�� 
�'.I��f��ahB�y�\���'Y�y��͐C�C'��l�Ё��'��$)���Z�ظ:�O�9_^���'q�H�B�`�V��SJW�l��'��I¢N�l����%V�U�F���'K.p	$Ĕ/2�Df��V���H�'Mf;$^��������l=��'$�M��#�s��26*�(
�E 
�'8pGJ�3�}b�����@
�'���!nޠ��c�^~�֘b	�'*��s�1a�:�ÂS� HTPr�'@�٠���8��%a���	t�1��'���Ģ�!]5��QDN��HS�'^��rb�3�V@[Q��)4����'��$3�͓%dPՙCiR�C+�j�'��Õ�/MФa�F�5��y�'A��1RnM@̪y�b��|���'3"\�0�I�!���0'A:y/�UI�'���b`�E�Zi `�6qB�9z�'�܅�!��(|���l5��9�'�Z����ڕ�㛒�b�#�!�Z�*b:t�4��_�N�1��H�!�D["ȤUZ�G���"9��)̄-a!�X�"�Ê�3�ܠgh�G@!�[�t:���%�1[��͉G�˗a$!�V:(�tab�M^���s�O�:+h!�l�Ai�%T��lA�oEYx!�DY�r��]at_���M�K�� ;�"O���iB%jz�!�"ȵm�4�J�"O���s�
F�b���3#h��"OX��@
'\���z��*\�C�"O�E�-�N�L��7�Y1V8�z"OQxan?+����`R�M�nPi"O�q���
Ә0Ӥ��h|l$��"O.�w��U��Pm�(]0=�"OԌB�*��?=��Q���1=���"O*M@���_f�����ԥw�ب�S"O�i�h��l�!�)�
r��E3"O�MW��nF�yT�T��Y�2"O2�	�I{0`<��գ1Ӟ�6"OR��bɃ"mm*pbpDݹ/h�y!"Od���Ǟ O�ލs�c��q�nLї"O��)��/ ���z�� ^���pV"O����|q|���`�5�|��"On��3��$��1��۩>��x�"O�t���0<���v�6"]���"O0���
F���[�.	RZ,�!�"O�]Z�nY/k���� �ų@$��"O���@��l�Th��K۵n "O%Q$�ŕz_d8@#
AX�B�"Od�7�Ԁn@XX�ʌ13����"O&��Rm��q��1Qr�?j�����"O�I�U"ŕHz��cb��N����@"O�
�n.uj�@��<>�$9��"OҀx�G�!9("���� "R1J�P�"O�MrC�$�ى��Z�J��T"O� �@'ʈ?HqY�߃0�"�P"O�lba�Һc�4�At�ɔ�H`#"O8usV�y��u�d"�"~X���,D��C��T?#3&$�CL�;�l��3/7D��bS��KB���S���SC�X�t�5D�� �%�M�$A��Б�K^�7�����"Ol$ 0��~!Fd�e	�F�Р�"Ob@qP�C�v�{�gF�~ݘ)!�' ��U��%��`�cm
"fEl\	�'+�h	���=r�����թ3[���'��E�� M�8 '�ŧ)?�4�	�'4��H�%Ӧ*���Ƨ��>���'nfɐ�G��G�T�f�B֐�
�'9����=,b�P���ݓ
�')����k�.[%� ֤�5�H;�'���"@y�����M�-�
�'j���g�Q�Ϊtc;H��	�'|���5݌YK�"^�9���'Ѡ�:e��w<E9��ͣ%��X��'��X7o�8M*vC؝� �`
�'U,Q�`�7��3���=��T��'��i@L�:Q6HDȓ˙
�l�'���b�Orv |s T7|�r�
�'������^�H�C��h`l�	�'�fi���
��`���M>0�3	�'����M���H�㓚,�lH�' �i��*�X%��h�#r���B�'���0W���f�H�p��=�08��'��!I���j9�ȣR�5.C� �'kJ�I�X1rQ�,!���3%�~�'����P�M�4`�bA��>q��'R|�kG�
,_&`@�	��,�Y
�'����NX�;�<y��Ά�D�~��
�'1�A���5p�Њ6�a	�'�ֵ
�N�xê�N .<tMK�'�F�9WHŢtҤ�SGA�5���y�'�����cI�]7���6o��y����'Q�	�(F)�ƌKq�q��x*�'v�9�H$!U0���Hk=���'Z����Z�s���� �+j�ʝ�'����"@�䴘��H�aD�y�
�'m⤑@bجz*�T	�˛�V����
�'�`���KY(���g]�I�^|(	�'l�|c@�	>��LJ1JC�)�����'�V�
�J
�"*��I0 Y��:L��'�rp�MˑH$��0c�)A�i�
�'?��r�K7�l�0�]�Vn-��'Et�"�J�I��Ipj]:_ެ�I
�'�p1�GʍL��*#DUl�=Y	�'�ʘ��@O�
c.u¢��Ȱj�'g��i�<ǚ�ue��]x�B�'���c�@/n����"R�
4�Q�'i��U��~2�FO��b��'$�y�qo�e����kQ9}|�@�'�  P��%^tz��"�s�$�'��X@�Kܟ&��-��L�zȈ���'���2���\0D]1b �"qҔy��'z��"��d� ��4O7�<q	�'��!V�C����3�5�F�X�'�����6朢Ԣ�.�n���'�.�@�^Ehy�T�Y�v9��'��Lj�U�'d� �� _p,�
�'�V<�v�׹/X���&�ĊT͔,[�'��4��^�@~X�s� Y�Pt��'�H��M�	�~d9���c�����'�l%��&��!Ѻ�.%` X��
�'R�$ V52�@!��Kl6Q��'=�e���$PƐ�$"CG����'j}�� ɼ1"1�v��<Q�%��� ��Τ,�d�1�®�y��"OD!�D�59��@�R�J 8��X�"O4�k)�8oK\��@\'�<Taw"OTը)����b0�ɸa�z9�S"O�u�E,˨G��f �	k������lCq��W����'l��T?����MTt;�f@�^i"�K���cG^����?��|#���%�[�rt�����\��D`>�^�6!B]�i���%�.��}pa�
�h��Y��	�W|�0 ���v`��`�2l�'�I�<Q��p�e�*�`�0в��O�oڗ�M����i�tکbb��H���DҦ+G6��`�S��?�,"��߸�r��@�M����I�M�ֲiʛ&*H�l����s=��	ׂ��~�c�I����'U�W>ų7��ПH�IȦi;q*Qo*Ձsh�h���5��6�j�X6���6���/V�nm޸��?ŕO��t��reJ�@�b<����G	(;�$M{A�iOZ����(��6��9S]"���U:�xd(rÂN����D�p�Y�2��T�@I1h��	�2�i�=���0��z� ��+��Ż�͈�bB�H�+˲#��������bX�p��ƑB�n�+�"J�l8v��ҁ8ʓW>�-w��O���ݭ�&*�:L �9�HA�6RQ�f�
�?�����< �P����?��?	�S?Qm$p]1C픀<��DQ���p�#d���v�� � *J>������:c�:qM$����dT����B�����̮8�d�fV�%j:��ˁq�$�ƞê��P�zy2��
z(����@*�B�(��Scr�ӿ�t��Φ��uZ?˓�?ɬOR�h1KD'����s�5bP�|�"O�0�ȗ�i�2�дc��5������L��MC �i1�'���OJ�I9mhH��(Ή`ʊȳ��S&�l��@�J]���I����� �%Nȟ���蟬�Bx``!�̀�[u聊��T/R{���i=���@P�/�Q�Q��)_��̓"�+:��	 f�H�Vļ����=�蔺S��V�d�kU���+�R��c�@3�qO��V�'��&JǗ}��5�7l��{-p�C<,��<%�<�ɀxD��?�;���b?6��H�l�.y�����y�@֯v~p)h煁 ��WC��~�%f�Zum�Ny���Hr6-�O��$�~�'�);q.�*'�H�Y���ӌ ,	.D���'���'ܐ�Q�FN��xK���b�F`2@k��|��D`'h���c#`i�CAc�'Y�q ��8$R8a�-�9�F� ����u�]�\�����<���&��E�<���$I"2�'>��,7m�!@���C�C ,n򍉷LNl&q��T�S���� �z��#%ѽZ�BT
<U�|"�sӰW�9�M3�i��W�,�R�Z+{�{��Q?�&\2h؛��'�bZ>�r���ݟ��I���CĮ��1(�1dmӚ#^�aT�L�8$����S�����U�|w��7h�?�O�����LmJ��XB�;�h��6LBQF�i����n�'D���X�$��}��8���*3�x��l�H���V��73��¦%[�����i#��(�+ۛ��~�d�D.�禭ء��;�v|���温��`?i��?�����d�Oc?���ȓ�"��D�^��lR��/ʓ*B�iO�'���Z�eJ��ME��Yd(�
H�<�K>�ۓEa8I�  @�?�   H  �  R  w  �*  �6   B  M  fV  /_  h  �p  \z  �  w�  ��  y�  ̡  �  P�  ��  �  .�  z�  ��  �  o�  ��  �  E�  ��  e�  �  3 � R � �& �. �6 �< <C !I  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,͓�hO?�zP'���|��6E%V�ၖN'D��At��j��KC !sx��rh8D�@+�-�65b��@��B��`8D��S�;���!%�*��u���6D���̒��;�mQ}\��Æ(�O�O8YGcĪ#�p� c�	S�Mi�"OBpX#T�~�LX�H�b���S�I���)�u�x� ��4����5�ĝ
�Q�L��	�#�6����jR��f��u��IXz�I�?E���c��Q��O@�5g�P���:�y�D��Ʉ	�&���B^6P��,�K����b����=��@�Z8
��`C���%�{؟,ϓ
��2��5�<�3Э�G���4�S�����a\����zQ�`C��?��O��~��c*Qkp�vH@:]�d�Hg.���x�G�+<]��ࢁ�#A�P���MCN<Y�'q��֑��	2*�*?J�����:e��[�?D����/�^�+F��)�xlcW� D�*��A�ߔEe,W�*��g D�+�O��|e
���;�
Aq�$>�ə;�Q��O5z�a&)��XX���S�z"�W"O�a�����>�^0�el��Ф��"O�0�+8Kܶ��A&�\��a"Oh��WQaWp ���I��Op����>	Vf�V}9�?.�Hq��j�l����>b"�)@>9��I�*��%z1^k��E{�N
<!~2�O�W\�e��H͸'�����D�
paN 1���N��P��J��~�)�g�? Z����R�r�X�
C�E�0��3�	G8��1* ����G/D"��%.}��'�ȑ7�P-S�5E\�R�
m�cM�y8���O�ĂA�[�nl��)�B,F�A��'q�O1�� O,9��Vj�!�X��"OB%�V�ɬ: ��(^#��5!��<��}����S���Ud�1��?b�XB��%E�~I���JD]�t: ���5axC�	3 �2����Lצ pT+E"L�pC≇����k�9
�*�ɰMڷ�V�P�'��8Z�Y������^S$��'f�CF�ѲaVʼ�ɍ�E��Y	�'{���`��lh����A&tc��ىy��)�Ӳ\���.�i[��x�A�ZќC�	� !$�@@��n��
��I�C�I:;tj�1��,{T�AxdC�I��j� �K��:�� �~DPC�	��tr�ǌ�.��˵�2G���#��:`� 4`��o�9҂ه8��B�ɢ��B��2'@�a��[�I?�b��F{J|"a%U�3�
1�%���iz	/�m�<Q@Ɂ=c�|�j#G�������Bm�<��c�$��)!�ʽ��er��]g�<9��S�-"a���}�
*�\H<�c&]�j����ǩ٣|9���A�u`�{��$��aL!�� ��\�O��ȅ�ٟ��O�����\�V����˫[!NA�p"O�Ѕ������J�C3�)�s��8]>?)�V�H|y�H8��7 ��n8��p<i�R�/^�ᰢ.лr��QHm}��i�M�?��E�*ctIf���u����F�Gj�<QA�
";�KЧ�0y{�M�P�d؞��=�R)��:v��S����T\<Ё��d<��-:$�*�o��mV\���;e�t0��N"�=rת�3#0�m��lk@�ȓS�<$� �S�?iN�bfe�.%�م�"�H���a���J�Y�F���ȓb5P*cd��8�9J 㓦&����	Q<1`ȉ��l�Y��@�I �yS��y�<iËǻ`,<�䂎 �v�	� Uy�<	���[�@f�@�(��� Fx�<i��>h�M�%K�}LV ;Fs�<	���$� @I��D��\�"!��h?Q����g'ZR�ꀂ2��E æI.\C�%54&�V�`&��B�%aNC�IR�d5�`̐'#�|ٱ�ퟑk�C�	�_߂��坙+� p�C1a��B�	!x������	x�8(Ӯ[�?���y���(5�:x(���a@�5bՂ)�O\��+,[�`�Ba@�o>�y2uJ��X�(��4�H����ɖ
.\�+5��f"]��W�u3���� QS��W�|��)�ȓ%��@�� 4\	ҝ���$r|-��I^~��� �����lUmc�/�:�y� �z�p�����pు�G�+�yR�}���bR{6�	�c׮�y�X�}p���ـDb���yB��,�$��FnZ7m:Rٓ����Px��i�0��7ϕhI�(C,Ʉ8��p/Oj��ĉ4^|2�xB�.R�4��GpF�y��
1����㊛�[]��Y��w�nB�	��`ɶD�-t�����$fpxC�(�p P�cD�NU�hy�$ŷ=erC��D�.��a�� G�`�b��L�#<1�S�? �D'�_��QA�Î�&��=��"O ���#-C�0�D��dvjt��"Oz���2x0E�eg�><j�m��"O�aJt#��#�,�1&?tx�e��"OVȫ�D_�W��)���;�p����'O�UGy��	��rɰiP%5"a�P��Α!@T��$6ʓ<l��P�E�0��옖�V�q��A�Ox�����~�ڶ"�(y"��
1Sb1ON��p��|�!Z�0hC�-��]��lB�0n�x��+D����ڡ9�>]b��&'��$3�g*�	jy"�韄��-F�J^<\YAfP�OY��"O8p��.�+�e��dS�>D�l�5"O�TP�]��cFC�+*(<I0�"O�h!�ǋ)5�@�IU��d��`ّ"O��K�F�Rq+�7L�@��`�+�yb���4���ڻcԌ���؇�y�B�>�TD�#��3���EB>�y"�T�G������< ��𕭓1�y�)J���c��פ��T%�?�y�%�br��
s�J�ڤ��į͟�y�&� ̬H��4:���g����CX�x2s'2??R�� a�+�}C!�)�Ox˓tٴ�	�a�fB��ТT�&�����/�^ cG�D�!�H�سގ�J��ka�Ij0d�v(��
�Ԅȓ[&5�Qmҷ<9X1kp���D0H���L�>L���ѐ@�.3�Eut�T�ȓC��I�@�daڠ���ɺ}E^�ȓ/:�8ʵ�q�K�b�b@�=D���� ����R�D�P�$)"�<D�( �
�
���BsNøY^p�`;D�� D��M�0X@�c0f8���:D�8�ǁU�IT*11Q�R�I�ؑ�R�8D�H��\1R�j�S)T�� ���6D�8A�LY1��98W��>���Ib*5D�d�"F_�rV����xE�-D��c�*F 4Wg���mʊ@h!��<��y�AT�FF0y�����,^!���=F��ir�I�jZ�Xc��۬F!��bڂ���D�4*QA�ɟ�!7!�d��y
�����"W�(�'	�:W4!��2d���lY�gYl�(f*Z� 0!��W�YN2��AB,O�P
3�΁F-!򤛋d��m�ċX+�p���F�J!��ʯd����t���F�Бg!�d�89o�!@؟���3@���!�$�1-���H�	Ԟf7r-��J�/K�!�Y����6O�=ov�0JɞI�!�$ҬP���KG�7rqA�bQ8)�!�Ċ	&I9;hѲ?8A[���o�!�d
4D�@9qt���:H���D&9�!��F2l���3�;0��*�,�)�!��&xp�ub��
4_h�@�,��!���L�z9�s�C�d�p�����!��D�F��e��ۮ}����H�:o�!�Jw�8 !�ڸӀ�Zd'O�T!�$Ӷp�T�����.5�4��Q:!�D�>E��AԿa��RQ���T$!���)�h9�(�!,�� D�G�rx!��7v�~�����)�`�i��B./;!�Y� ��%�WK.U�h�Y'I��b�!�ٷo��X�RnS<\�xP��(A!򤕡M�<��&��>]Z�Ş�<t!�H�Kٰ�!��2-tBa� �)D!�� �	��]�:h��
���� 0
d"O ��@�ˁ >��g	�*z���"O4��$�6�x��_k�J�"O(	b&�ɠI����u혽-f�5*�"O&\eJ��'3��-��i��m)��'��'c�'��'c��'�R�'�`IJ���K���¦��'a�B�;�Ħ���Ɵ��Iܟ|�������Ɵ���ܟl
��T�!u�pB�IO�M*ӡ	쟄�	ӟ(����I�����D��ߟ�r���'(��� �%����I�l�	ٟ(��㟔�IڟP�����+��wo�����zbv-�`ʍݟ��I⟔����H�	��l��П��IƟ(b �	*=4ޝ���Q':��ç�Y���I���	������I͟X��� �v$��i�8L��$$P?N�� �8�I�<����P��՟�����\�	񟜠�f�C��$d��6�m'E�ٟ�	��T��П���ܟ��IП4��ԟTh�"Á^�01g�A�]Dn�Xf�YǟD��؟L�Iܟ��	џ������I�4���]0P��J��\4G�@1��/��x�	�(�I�����������I�@��+ �a��@*X��T
��ȟD�IɟL�	䟔�	埸���|�	ʟ|J�� +:�"q�e��MV�A@�����I����I�p���(�	̟h�I�����Ʈ|�!���u�A��L���ş�I����I�T�� �M���?1�-��l�r�z҇�3E��@C4z��	ߟ�����d�䦩� 'N�2J� x֏�$e�0����#��lԛ6�4��D�O*Ѹ�hH� 
~A(�DݻckQ��O���M>C	�6"?њO��8���9��$��ᇉU��* �'T�Z��G���R�r��`Q�j�5���בK��7M��
�1OT�? ������50�ѣ臇�Xx�@-��?a���y�Y�b>�i���	̓'"A ���1�l��C=[�bH��y�J�O�л��4����4=?��`R��Hb��S��X�/��<aJ>��i�H�yB^�0�@a�D�?7����q�eU�OZX�'���'��>)���B��y�(�N4r<�k~2�'?�!V�S�ؘO?��	�X$����j` x;pkI�&�МP�*�}��my������$�I�\H���/,R�]
-�g��KצU�`*?��iY�O�	]=K����ٜqfF� �EwC��O���On��"iӬ��������,1�HѮe0FL�U�[u��4
�B������4�����O����OR�� y�>}Q�U��&�p���6���OǛ6�E\��䟐&?A�Iv��$@C�}Sba�0�G�z�=� _�8�	ܟ�'�b>A�䍞;������A砼+0n�~,R`��i(?qW��1�P�$Ґ�����L�$�"5�b�X�?L��(�O�u�X�D�O����O��4���Yh����#bcE�M�8�9�J��+Q Q!���1m�H`�H�O
�DG}�'�r�'�d����43�.1�a�H3c��\Ҧ��L��OBY���,�����t�w@(g�:���q�� ,%d����'��'���'?��'���j��9*������
2C7�`�b��M���?i#�ipf�C���v�O|�j$nP�ʪ�Z���B6�]��'���O��4�:���良��i�]��A:_n.��Vm� �,�a	C!-��ɍm��')�I�`�	����%#��:�m����`qB
z<,���P���'|7�^+/xF�D�O|�$�B��@�Š���E
�u���q$��q��D�Or��'&B�4�6�DЊ2��aA� ι����.o�`��r���9���ѯ�<���~����F?��M`��$��?��[4�7�\����?	���?��S�'�����IІ�??��RanW�|S��qA���\	��	�9�4��'���?Yq��4G��4�4t�i�v+���?��+���ܴ��$�l���O��I�6�  &�84��/�HDf�IJy��'j��'r�'�BQ>�I��@��Nͱ��Sv�Фz�LR��M+��)�?����?K~���qQ��w���[�F�-0�(\S�M
^��	���'�2�|��4޵[��	c�'=��p��_pd��&�(����'�N���!G矤���|�Q��''x�Aw�\���1���\��Ԇቷ�M{q\��?����?��ö<\��{�aѓbd�=*�A'��'�꓌?y����K�A� ��3t|i�m�0��'e�!OG�k2$Z��$�ߟZw�'�a3�fF*��(`�E�W�M�v%ΉLrR�'A��'g���'}��jPJ-k����`���'r'"�}ӐEiP��O�d�%��s�I!�j�b:�(Ӌ�p��dcc�x����D�I(E���o��<���F���֦�?i(r�սV�����@L\xs.�Ɵ ���j�����$�O��'6��'�v��d�t�nٵ�͜qt]3�[�|�۴���VE&�?i�����<f�� $!|�s#�ƨ}�J�����#�������	O�i>��Iş���A��"���1�ꅶG���C�P֤m+�/)?!���'����^����D������g�ښCv�9� mF˲�d�O���O�4���sD�(�evR�Z.r��x+e�K?5.�z��0Z���lӖ⟈ګO��O��Dڀ>�H���-�}
�Kߙ\N��[�ô
2�	�3���O^�'?M�=� �a���V	���0jJ;3=��R�6Oh���O
�D�O8���O�?u���u�^零����l���ǟ�����(�@����j�4��[�BiQ������6�M>	��?ͧo���� @�L~r+Z%-<��A���JW�P$��,�0I�%��p�d�|2S������Iǟ����Z�Ep�����9�a��ޟ0�IQy��nӶ`���O����O�'Ā��ICl�̑�4v4��'����?�����S�Ԯ+,��ԓc��	 ���$�Q�N�a��ź���O��Ա�?9�%=�DK�y�nh�5��5�󧉔i�����Od���O<��<a�i��12�/Bh�	�f��9QJ	+�e����'*�6*�	���D�O� �(�
ξ���N
>sV����O���շ"|ޠ�㖟@�4WP�d�~��L VA�}e�ۍpQh-I���<i-O��d�O���O����Ox�'{������S�� z�
�$���i�XL�A�'�B�'���y" ��n��szX�J��\l��(�.3$���OX�O1��C���.39�DT?tMF���F�Yu�,
E���D�Vm>Ĺ��U�O:��|��+�
��s�\� �7A�s1
�3��?A���?�-O4�o�R6���'
��PJ�K捎<Y}�POŵL��O~��'o��'�'_����	�A.`��D�2)���O^���);Wh7��E�ӭv����O	�4��%W|��桂1I��3�"Ỏ�s��KR�|a�G�0�0@�O��m r���	ǟ���4���y�!��6e><��oY�?�J��T���yR�'��':��sv�)��$X	�"X��O Xi�ֆ=��c��Eyf�Җ�|�S� �I؟����Iޟ�p�f��#�ɛ��tL� %$�[yB,k�`���g�O����O蓟��D̲��Y��O4W�\��W���`�PT�'���'ɧ�O�PaE�A�Q�:����
�b�h���
aU���O`�jFEH��?	�+:�$�<ђH�;Ad��&/I%�(��M׶�?)��?	��?ͧ���������K�ן!"h� �yuƕ!0a0̰��ӟ�y޴�䓢?�]������	9cZ�K��\ :��_�<�!�6��;���y�L���쟄�KJ~�������)m(�|xQF_�!���Γ�?a���?����?Y���O���qW�ۈ	��ؠ���r�2��'d��'4�6�_�(���Oz�mO�	�9�F��W��Sh(��%�Tc���	��t��0<嶥nZ�<���bs��gf�X��Ӂ�Vz��%�o��ud��ݾ�?YPd��<Q/O�������d�O��˗nS`�UjR�\0'��Q;P�P�x�Q�<1�i^H�O���'��$�w�f��`�0=H4�9 ��Q7�생'�΢>����?1H>�'�?����,��$�h�#x�H��)X�@DXׄ�k�"L�'��Ď	Οl��|r�[px=#2,Vq��J�&Mc�B�'�R�'=��TY�D�ܴ�6@�mD\�H��m��J�E���?���r�����b}��'2��Z�ƨrz�+aϚU����'�'��d�d1����O0ݸ����
K?�Bb�X$4���8���p���*��x�H�'r�'���'"�'�哟d��r)�s���ħI�/1�!�4Le(����?a����'�?���y�@ڷ>4ʉ�h[j8�H���/Z�B�'�ɧ�O��,�"�ɯ�y���D�$`C�%ۋ^8n@���yRJ� DH���I�M�'J�	Sy�T�(a0,	�G$$dDu�vm�0�0<�"�ih
�K�'�b�'TZ0�u��9_gV� B`�g|�<@s��FS}r�'�b�|B.��a	��{�B[�H%�a;r�G�����*��T6FY��X���P:�'��G�t_�!���:�t�S�SE0R�'�R�'�b�sޙ[��Y�2�ʵ$Idz���)�����ߴ^ ���?�V�i��'��w� �r�
�1�n'P�\y��Ț'�r�'`���(�"ݚ�O� J������ �T1����Cc�P;U�Ғ Y�L���yB_�`�	�?�I��Iǟ��"� �ul���	�s��Ej��H�R��N�z@�j��'�2�O��4�'��?�>����'`�5� C�v����?����|*���?�Fal��r��?��� ��ѡS�d(��4���ԾQ�V)��'��'�剃�A�Ui�ml���*'6��IП��	�d��3wA�ȕ'��6-׀���T"t ��I�ATY�t��
�P��
�I'������D�O
�4�f�JtD���"�[V	�_�,��gBv�7M|��ɩP������O7�e�'��T�w��٣V�V�/Iz�:���(Ytr�I�'D�IX<5��'���'���ԭQ1~1X��7S4X�T�!'�B�'D�j�IA�d�Ov�� ���%�蠱�݌	��r�*5&�E�p��L�	����ɟ�`Ɠצ�͓�?�A��s�� !���Щq`c�=�J�X�ʮ�x$������y�fW�\�x�u�I2c���a��ը�O|�o�H�p��I͟H��b�dm�~u�]9 dB`N
�&�����AC}"�'r�|ʟ�|*@
��<��5M
��|C�ȧ/�*�ҌZδ��|d��O~9�H>��@ 4l�}�"��.F�&Q�@�?���?���?�|:.Oʅn��)�l�ѐ��+K۠�dH
�~�$B��ܟ��	#�MCH>Q��[������F�% �D��W�ȱ�~P�a��P�	qN�D�QK$?�@�R����Sy
� ڸ#�F�*S��;7mG�?'��I21O���?I���?����?i���)B��T��d�g���Q�b�9}N<l�4<���I��`�	F�s�d����`EN'H!�b�ɮO�j������?�����S�'y]�ɲܴ�y2.�0(ن�#�B�+K�R�)��y�m1$F���?!/OJ��|��F��)���+@2��x�G�_�i��?���?a/O��nZ�{6@t������ɨX(D��Ĝ[�`�$�7Z.��?��Z�4��ğ�'�p�qi_?	"���F�vh�����=?qWo��oٮ5����|�'jئ��ϼ�?��cG8@�����`?&@HB�	��?����?���?)��$jѬt�/Γ$p��`jS�Z ���չe��BnӮ́@�O���ަ���uy���yG%��w�}KM�G�(��֯(�y"�'"b�'���G�i��$�O�Q�t�ޫ�:�.ߘM��Ԁ�C�"4�xg�Y�b�`�O2ʓ�?����?����?��b"�u
�N7C�08��յs]p�/Op$lڈ	����������?������		nJ�ʴ� s�0�:���QR\a�O����Ox�O��O�d�|aT�Ìp���I�	�&=Qt!	1tà�'���
Ԥ�O���|RF|̓���m�lE����<�FD�pKr���$�O
���O����=C��-[�f��L��tH/:14y&��+_��EG@���b��ī<1����������i�	���b[/K4h1(�oӉD�n��<���.�m�Â3��'\���wn��{��4}�KF��Sn�Z�'�r�'��'T��'G�%�BK��C��2�j�3�P�X�'�O|�D�O�xnLo��S̟��ܴ��\!*k��`M�"�@�$���H>!��?ͧg�&���Do~�A�;D�j$CR	��!�5GO�+30�e�Fs?������<����?!���?��P����/S��0���?i����ĦQ����۟��I� �O
 ce�۪7uJA��C6�>�c�O~��'`��'^ɧ���4E�����$;�d|X��P�%��M�Q�>F@26�5?�'%���L�;��l�Ǔ�c9�I� *B�	6�M� D��}p�J�>�ĩS�'�i�����?ё�i��O���'��Vi9j����ԗ$؊Ԛ5m����'��=��H-����xA�e
�~��,O�` �B
0z["Q���ާ)@���4O�ʓ��=�S�-j�9�
�d����1�"�&!�'S��'=�iOæ�ݯl(���a] _V����hj��I���$�b>]���ÎhP�I*OTd+n�"_�(̓%WP�ɱ�v,"��O�O˓�?�� D� �˻\���c4��LG� ���?��?!-OxTm��Z�܉�	����Q�r��E�'U��1
�73ء$�����$�O>�d0��~r�Q2̃i�n��E�F�H*�d�OHhAM�t\`�t�<1��c^p�$��?Č��6*F�y��-1�8d���L�?���?���?�����O��� �83vp� 1�Ϫ<Z�.�Oʡn"v�f���˟|ߴ���y�ۢ0&x�ۇlޏL���iq��!�yb�'���'�"�PV#�"���7,-�0��@a��H6�5
��√����e��O�T?O���|��'�?1���?��jD���F�=
�� ��>0mX.O mڡY�:��'�2�O�D��'��e	�0�+��
�rN�Xw�&���?i�����|���?�rM��^�"�2��H�mc�ƒ88����4���Y\��b���"t�J�˂H\�F�D��$�&\�����p�1�r�-���U��6��h��e$c61B��P�
U��<`I	����jYO���w��	�����֨!ZDU@��8��8
j�   	x��)YQ�����>�8@pa���D���!�@x���E*���1�b:��&3=1�����!ߔ �'�| �asSB5Bv1��Z#x@�(s���]�(��V�z��e"��<{��{���9q�"�R�Hv�Q@�"i���)j'�G/Ԥ���K�(v$�2�T'�M(O��D�<	��?)���P���O���Cg�� e҈ h��I�-�*���Of���O(�D�<Y$�ZtN����Cg���pK�y�f��,=�����ޥ�M������?��K�����{«�D�X)�fER�"f�q�m�9�M���?�-O������b���'tr�Oo�(�Y$6e�1c+,��e��0���O��DB",���'8h���&-�k��$C!ON:�m|y'H�7��O���O���a}ZcD)7��9v\��3%ޛ2?�x�ڴ�?9�H�"m:���׸O�0T��(V�܂�ǂo� �ܴ\��T�i���'�R�OWl�����~����f6�tZb,D!�LYn�����I�	o�'�?�t�ڬH�(�hP��&�Ω���Z��f�'	��'�����Ǳ>a(O2�䫟8��#�&
v���C��j��$�I/�Bb���IƟ$�ɏp���`N��-�|ՓDg��r2�y۴�?�1�ׯ��I]y��'ɧ5��6q(�葶ٸ9���+�%�#���];a�����<Y��?�����d��iP E��K4�p��X�_+⹰�T}�[����^����	LLĜ#��38=�ⷁ�LP*0��y�	�p�I��4�'��T9��`>};��ŉl�z��N���0Tfs��˓�?�L>���?���η�?���=S�D@��5[���0
�F���̟8��ʟ0�'
X���%�~B��S�����T�|�X�FD	��|h�i=��|��'<�&��qO�a��Z��ቄeք&t��y��i���'��I=$�2-pL|J����q�? De�F��^�>0��<XJl�%�i���֟������	d�s��01
��˛y�)�g�7E�\6M�<%-�F(��ɥ~����*������bE�B�t��I���TPp��~�^���O&�$�O ��O���u�ܴ|�R S�RN�`���
��DoڡR&���4�?���?��'hՉ��\c�0H����-\N9����D�A�4�?����?y����Ķ|z/���yfc��H�J��%��-h
v<@��������* /ˡ<�O��=��c�JXhf�)�A�K�2�"�)d���Og�OJ���*_�T<�c���j�$��T�i��cƒc��I���	/�	�W�>h��
 xa�y�i9T���9I<	�!o~��'�"�'���f�[(�(.T�PoGR�@PN����?���?-O��d�?	��۷B���P�ʄs���z�{���$�<����?����D�Fn�p�'r�L��w��yb$��*O�,vʑ�'^"�'z�'_�i>-��"xÌL{!�N�$dL�0� �Q[�O����Or���<���)�O�^�R�兺Ux lB��8W��[0n�:�d/�D�<ͧ�?�K?)C�G�6��(r)��U��X���~Ӑ�$�O"�:�̥�ד���'��\c����T�O�t�Q�Gɞ$��!��4���O��D�O����|�+Ok��\&\  ��6c�h�b!��A��I���bcf�۟����@�	�?���uG WU1 I*%+�?���$&˕�Mc����B�N���4l1 ��$-��p��?w���'�i֞I���' B�'�b�O�): ��S��ç�@���I��ʋ�I�Ɂ��#<�|��J�ޝ�C��xJ�{�ꇲX�n��%�i7�'L��؆qT�O�	�O���9�<�Ek�1 �p��[�B�J@mZ͟��	Wy� �~Γ�?I���?�p�Ά<� Q��\���\�`X5���'��(C��2�4����;��*MϰD�s���Z��"��� D���$���I\�Iȟ��'G����H��u��j����$[(�Z�(���h�?����~�ǂY�P��W�B � �Mk5��d~"�'�b�'��<sR��	�O��l���P `	���Z=�޴��$�O���?���?��C�<�$��n��Q�L8�� ���2���؟��	ҟ��'�h�肉�~b�n���_*w���(�+�W�ؠ��i��_����Ɵt�	�K�����`��<x1�&l]�`�JC㘥 @8m�����ILyL�T�맜?1���b��ǳ<��Zs�[���¥L6 <��ڟ���ן#�9�s���|��;�ȋ�[� �k^�7�imZQy̅ ^\\7m�O����O"��Tk}Zw4ޅ�bffm9(�*�2W�.9��4�?I��b؂�͓��$�O�>}��	�3Y��x�?pv���gd��4+�����ߟ��I�?Ey�O��P��l�1�U�B(����
�fS���ĳi���'�\���
�4�:��gG".��@`ɏd��k�i�"�'�K/b5����OL���y�Ҙ��S�,���CSj� g��6-�O��$R�S���'Bٟ�D�!�ʡ5����483R�qc�i<2͈*S	����D�O4ʓ�?������4�cZ�#F���'T`�'3��'��'x"S�H��<z:��3���*���ͅ c��!��O�ʓ�?�(O��D�O��dZ�RJ�pJs���/Lnp�eθ8>�5O<���O����OL��<AuO�{a�Rqvp%�1b{i�$JcLW�+[��^�\��^y��'3b�'ev5 ��5f�ڣjdXx�jN�-��
�%����$�O��$�O��T��ɩ�U?����jӊ`���%H/��1a��P���ݴ�?),O����Op���5��'ʅc����@X"2'A#j�(+�4�?����dE#�<�O���'���I	�]�S�Y�z�J`X��G�D��?����?���<�����?i�1��"}�4�����]�N��%�w�d�U���B�i���'�"�O�N�ӺÕ�Y�a�����@���K�Ŧ�i�n`�@�	��'#q�Pp9�-y�!�Q�f���ҲiFR��"Io�����O��������'��ɧn���+��mh�t�r/Q{@��ٴJvD���?a+O��?��I�"2�ъ��΁|XMR)B#L7Lts�4�?1���?�!�͉�'�B�'4�$ܸ��
��"n�e{[r��ډ}��'�R�'�¢U��,d�4A���ҩ�a�b6�OV�s0��X��?�*O�����A#�N��*|������ �ER� �p�ZşԔ'ar�'*BS����U�9dH�D�%��)�@
!
a\�K<y���?�L>q��?����y:�r�h�#
B�JC�V�Wt�������O �$�OT˓X�ڑ:R0��48���]3Jɡf��Mn��j1Q���I�(&���	퟈��|��� ��4�n��GE�2��BҼ��D�O����O�˓2l 4��t�= ��P�D'���V��e��7-�O��O���O�q)��(�l	�V���6�y�#���F�'��Q���#,����'�?��'��E��M@�$�)��K%�`{u�x��')rߺ�y|�ڟ��Z�H�8p
�D#��ƛ/Fl�1�iJ�I�1n�$��4C����S���D	�1���A����8Hg�'�&�'7r�!�y2�|��ɕ�wT �ؑ��7	� i3���3�����T6��ON�d�O�)FJ�tT� �C6#p&�!�4�L\I�p��i�R1�'��'����D�^=�P��L�ouz���F]"���l�̟��IΟ��PG�����?Y���~2��qr�k��F �B�׋�M;N>a�`\7ŉOxr�'<Rl܇J�p#�(�>�Tʝ*
�f7��O�$�%G��ҟX�	@�i��Z��_��ڤkC�[|�1hϳ>Yd�U:�?�+Op�D�O0��<��W/ n�B�d��D�:�*G�Y�`�������OғO��$t>ݚ�cS�?��p��1$��y��� �:{4�D�<���?�����䚑	�-ͧvW��\��g�ٗ
!�@'����w�	���	'�T��+�r�LZ�JѲ� Q5+��\��O���O��Ģ<�ƭ�!.��O�\p�EK4��ԣv�y�I��~���6���O��� j�l��>}"G�?CC4�{g�ڿ^G��2����MC���?�/O�i��Ba��\��;C�����6��j�+Z<M�0�I<1��?rƕ/�?�H>i�Or�qQqʗ6D���H��Yݤ1�ߴ��+�즽诟.������'$�h���t�&���S;�����4�?��8+~������ܸOeJ��!2pO܉ ���7����4;젡0�i��'sb�O��c���,�(�\�!�����Iڒn�:�MK�L�?L>ш���'6� �Gf8���_+T<2a���l�\���O���+HSƘ%��Se��ƪ5�B��ź���?W���p�4��'��8�d�O~�D����	p/���� Ab�t�t�Ц���		I��H<ͧ�(O~���CS�m��e3D�[�Cѐx��'/�ן4�	柸�Iʟ|���ڇ2e⍛���R�Η.X���Cr��O��D�O��O:�O�$�� 0
H�O���3q�RD�h��M|Ӹ�R��X������}y�KQo0��S�
�@��R#�8��2��޴듛?���?���A������x��h����Ufr�YC(��IП���ӟ@�I�� mڢ���O��r7��'`���D�+1�:4C�" ̦Y�	Q�	��\�'H�t�H<�6�<{��|9�,
V �#�ɦ���Py��'�v^>���ȟx�S=x�jHQ5�";�fQ��ɟ[t�p�K<�����U>W��]0cN��`%��{y��C��
\�67�<�qm�k���k�~��r���lc�4�rd��@᪡a%�{����&�O�, T�H 1A Ѱp�@����R�i�p) `Lh�^�d�O�����|�>iT�{F)af*+|@��b�6�a�'��R	�}qQۧ�I� aH���~ӄ��O�$��t�l�'�,�	Ο���In<x ��^:�2����S�P�j��>���y��?���?��!T x�v�� *e#�C��L� :�F�'Y\}I%$�$�Op�$$����q;%FɌ&��eZf��1sp"X��Q�\bP6�	�O��a�̐��*	 cn��J��!��F?!^���7�R36}+��U�WT, ��k/]�AX!>��=����:Ni�4F9�Ifx��G�\�9����ϣD��>Qs�׏~ĉۣ�݃g� �T.�sT�KP.�P�r8҄BZ���b�_��:�h��(G<�[@J�',T���+�|��X�� "�
����P�"�ʘ�s��,/��d8E�C�y�`����&#���.L�Y�zG�E�3:��8#�:A�&9V��K����pDDN�F-E�0�����M!�B�����"R��I۟��ɝ'��&	� 	%�W����T�[.��E��y�b=9�)?X�Ȣ<�	b�>�)�(�/b�vaF0G�<)`���7��i�ҵ8�y��2��Fy�����?�����Om0m+bG�8�� Pa�]�
hHx�'u�Ҏ��V�W P�$��%:Є�0>9s�x.�7	J�I�o�{1�g�˳�y��.����?.�*8IWb�O��OJ�P#��B]�C���~�Ӓ��=A��P�Y�H}va�O�h�矔	 ��8�tX�EH����[P�A�(=�<�L��6{���\�"~����t��5�6T�rl�i�1z%�YB�O�П��Iz~J~�N>)��'s/
[d�}U��;�ju�<!D�ǍG	����'/<�b��#<��)��Ά�6�ㆨ�f/����J��?A��y���)!#.�?����?��f��.�O���X�Z� ���U#tSʩ�$N�NL��Ŝ�����	�W��㉪vw��'�f�M╨m�ƴ �'��)���'�Y�Հ)O�\��@ާR�<0y��K/Fa���w�O0�B��'mr�IXyb+�'pV8��̗9�y+B�S��y��1G�ʜbN�wN���#)Q�r#=�O��I*y,�0޴W��ѫE�S���iҎ�<nI���?����?�H�$�?Q�����k͈|�H��Z.��tIӧ�<9�xj��<�R��B�!lO�q�aӑb2������/��XR$�R%HD���_]�]���I2����OHP��[(P)��)�*t,��`a"���OvZ@xD�N���U`]��!�d�	c���qJ�Py�=([����2O�%�'�剕J�p�K�O��d�|�4��p��k��Y�&<�f	I?�zY����?��f�Nd�h�O��(�T��>�O��Q�B���X�e2�Mߎ`� mC��-.�鋳M�~����}� ��5A^�exd�g���3�"��t剈M���O�?��ή_v��T�ʁf"a������	����
ۺ9(: {օJ�&ǎ���L�ID��Q�'�̆ �0�&F�z�z扅	i�d�O4���|�LA��?����?���h#m�P�ۓY��@4�bC���5@\��`�P��Vr�*�2b>�$J/v7��,m�`z���v�&%s��u�L�# D�WO"��S��?AA�
c�	 ��m�d����8C歀�4s�v̭<%?��S[yb�R�Z(�1gی�v��b���y2���j�{�U�i��\ �O�`Dz�i�>!Ǡ�aDh��@�Ha1:��sk�.�?��/��@����?����?q�@��n�O(�$�gI�R��T����ѭ��j�	$�.�0�N�?)��ИR*8�*g�R !�'
bx��C��|���'R�+��.h~�� �A�$��O��
�K��8�<s�J�ex��yq�O�ȁ��'�:6Mڦ�?Q�V?���ӗu;$$i�P�s��䚀�0D��*�c���`q�mL�>U�� �HOf��'7�I���"ݴ`t9y�g�+f=�1c�@�~���?���?Is���?����D���?Q��]�:x�c�H�O��ȐUmԚ�rQ��$f��T�2!k@��(� �c%.��Ɏ0|�D�O:ebMe�}�V�Ƭ X�7"O�Y�)��8�pl�A�n�5b"OVE�&��,�a@�'�r�h
�=O\�>����֛V�'rbX>�5f�Uz���S*�0������Y���I�0���(�f��	I�S�d�V��~��ŭN�|N�=�6Ü�(OB%�$�S3g>mzqe��MB$`�Vi�F�&�<Y�mR�@F��@�&vܔ�i��L�7��`�g!�<�yd\mLi���4XR]r���0>iU�x�@� 
��P��^�To����,�y���/_��7��Oz��|
`NL��?���?�a�%��4��N�#g�������p�������I�j� ����"�F-*S��",���AS`�Y����2La�);'�L�T�����lS�A�T�'�1O?��\�_[d���Q����-a�!���&v�K���`��qHmH�{��҈��?��(��d��軖�W2��(�����I1>qT�B *C؟���ΟT�I��u���y�HN?PH��FO�	{� ��E���~rbH+��>���|��i�3�M�,D�8J�Ɛo?����Ex�T�P�y�x���2�Ԓ�$��ԃ���O*����#A��q���+�����
%{!�d�4:���9`�	&D֌���бd�ȰDz��)΄d�4IoZ�{V����K�Q�LRR��p��Iڟ�������ph�ϟ��I�|j�N՟��ɓi��PY���fP�C��7L����%t�IR�Qfeȅ-�i�խm����D�V�B�'�0���mA����_3KE����'������A-2 ��;Cf� ��'X}�U�ſ��4ꆯ�\� K�'ڢc��h!6�M���?y(����>�{��`\D��$T���d�O��ć����,�|�f鄌~*,������`F�ūp)�s�'�܌���	�1��ғQs��l���0R�Q���O�}w�Kc�"�ǋS�P>�V�i�<�7�I�{����f�#Q~*���\�|sM<���؛yo^%�#��c���� 	A�<!%,48�IԟP�OA�Y��?���8��8�4M�/�c�IK~�,C� �|��y��D����`���C����e�'��s��"S n��.u�D��ܥ���fH�~��~�IQ��mY�gY=Ef�5�f�	�h�t�(Տ�֟D�IJ~J~�����$λq�x��EQ��ejs�X3Z$!�dX�X�L��B��h��Q(I8X/�����?a"�(�
g��q���x���`@⟐��T�~���؟,��ҟ(���u��'��ڹT��Ъ���/Ҿ�*��ء�~�b[���>�c�(�bݢv�U�����r?��mlx�P�g��)��%yN٢knN��v桟P�Ĭ�O���I>k�t� 6�،[�x`P6T9#�!�dH�\���\
x4 ��/�x�Gz���\�o��Pl*	�T8��@�FB����7N�������<ia�Z��	�|Z5�� ����mL�j�p�BH�U���ǂ��3Cx��B�B�ayrꉛ<^p�ăD"p�$��	yE#�J��!�=~����D��B��� 0�L�,Z����Lɑ\����*�O��E��'���I"nX�1!E��w∨�'�����z%��W�$�'����	�Ȥn�˟<��G��K��Z�N�;d�ТJ�"����0JQ"`�e�'��'�P��W�'�1O��h�"u
���'8�5c�
lת�<��+�L�O(�����'k�*�R�H.-6r�ى���,��u;��;GX$~���AiT<{fDB�r
�*���ڢH�૖�e����M{��
Ezjap�ٻ!��;KS�Xb��I�e�~��4�?�����$!S����O�����I�x�i�^9"H��QQH�8QN*5�9O�c��g�'����� ��[8���d78���R��&�(O?�ǫsM0 [��	R"�����F#p�*�d�O���3?�SF��?y�)R�3;x8	��ێF� +���<	���>Qg�ͭaV�i�aL�!rH��%
|�'|B#=�OS�ZT�ԐU,�x"��� B��'a��=
�\]	0�'iR�'��w�!��؟쁔�Q�?�܄s�F��	�ٳvl����'�0�O����(�?gd��E��+N�,�PU�Op��c�'�T%�a�����"gͥM��1��'X`�`���=�El�tPSFl�^2�$r�Pb�<)t�Ͽ&2�3`�Ճ\`Ը1Rn�"=���"|2T�ƳCV��%
�g�l4!f�	�"-�B*�7Y�'k�'L��{#�'��0������'S�c�$>�)��ة{��ƃ�p>1�jHFy��L�Z�������TI��0����p>���|��?����6q�$� �0<*C�	X��5���Q��-i�&��C�ɚ�n �IG �öBG)�����'T��ѧӤ��O˧>�j9b[�N1<���	d��P��H�3�?���?�fn��?Y�y*�
�ۣ8�����h#V��+��,%�¢BD�=
�����apU�hr�'�!c��h�0��FN�?͔	��!3��E�r"O����$�*�0�l ܠ����'|�Oz؂����A� �r%>�����?O��h ,����	�\�O��պ2�'���'բ<��k�me�l�ѤCZ�L@pP���B�T>#<ѵ�Z2�huq
�'��B&	?]�pU����O�C�ܢeȾy1�#�C�����L16���$:�)��LX&JT�F��P�ĵIi���L*D� Pd��i<��٠��\�*}�A(�P\����ĩ�"kB<G
ϻ@�Q��?���í��C���?���?	W���4��X{�A�s�@�v�L{��A�v�O $Rt�'z>R��L)s�A�$}�T��' $���)��E!r*��v2r'2�C�'ZW?�EA�����I�:L0�u+� #	���Ka�vB䉟ߐ�c�,X5�Rኰ*�-�`���SU�~��ش��ċcQ�������G!L� ��?y���?1##Z��?�������?Q��f���7D��Xd\@��������	����JL2���,���A2eܳQr����	�s�N���O��0�	՘l^e2�FBE����"O*5�F� �+��]��$�}+���"O����a�7L���#�����B7O8��>	&cL�N �V�'�_>��慕8u�| ��.�5XX��٠�f�X�����I.5��	z�S�tg�"f��`+�Eò}��a��(OH��4�S�H��`�-Κ=�D�pf�[�1.أ<!��]ϟ�D��e5#��tX$Mġ	�؀��͊��y�/W�BKl�#5c�8��[�m��0>Ǜx�ӗ;D`U���������F��y"J��S�6��Oz��|:p%ԁ�?)���?�a%I�	��S"='
��J���Lt���嘧��I9.tf5�Ŋ�cI��ǉU�*�X�۰�[j�����(n�]H&��;c��!S�/�r��'�1O?��ŵk&\��b���S�z�ף���!�ğ Q�NiseW4]�2� sHM'<*�T���?���/	�<�X=�q�� 0��Ȫ��Hퟀ��5J�<����쟤�	�����u���y��V�v�^*��
8�����~�n]���>�P�� 8��=h�0b3Ãc?92g�Wx�D��c��w�<ʶ����:g���� g�O��� ����*x��)p����
@�yҲ"Oֹ�'M�K^���pJ�5h	�)��Bd���Buh�B�ۦ����A>9�� �T���3���jg������ϟ��	�0����x�'���	��ܘW�M}�t$!u,S�|y��; c3�O|Y �X�x)㡃	t	��0��hjQ�`�0�O�	��'V�gH�"�D5�"��EF%�`��y�G]�L0+�~�>��!J��y2
���)��Ք|���`*�y!�I��L�I�4�?����	G�aF�ۦ+�&[�J�끎S�5>�I��O����Oy  ��ORc�ʧq��q0�� A�cK�8h��Dy�"ő��b<S�
�}�a D�hB��3T�<AEj�d;ڧ��ͩ��^��k螄}���c�2���H�(��e��"ļ7��X��	��ē^[�i8. ,C�Ƞ��S<���̓h�*;Ժih�'�哛_�P���ϟt�	Il�Y�P,߂*A@|
�.��W_0��6��ܟ(�<��O�@	�MުB�@�[�₳_�\5��l�,#<E��aM����I�iC��h�C2S,����?��y���'���R�Ɂ��Pu��.TX	�4��'���Iƙ3��:�HR�����Č@����U�8�T�s��>0v����ڀr���$�O68�T@J�V����O��d�Ot�;�?�;b���r5�!�I*T�4j'�O��3��'�Ԉ�-2�D��L�^�B��'fNI��J�p��� .6a�ee�=����>���o��l[�%!Y��h���j���b%D��)�Щ/��u*���.o|�1�(@'�HO>�Y����MaV4'Ԩs�>]yxY��f�;�?���?Q��+zh�K���?q�O>����?-<H�;5C\�A$�� �u����ɒ���r����c�8U�D�G��^�^��� aTr��O��Q�l��1PHu�	��Ɓ1�"O8ղ �G!b#���
F�v�	@"OI�N˩�H�;��z�N��;OJa�>�s��.RY���'��S>��@	Q�Rm���8�\Y�@(1c���˟ ���.�����[�S�$kC�"�.�I�L$w^�I4�V�(O�@`�S�HH���S [�"[��+�f�!Fo��<Y��H���E���	1Jj���ī�-`��R��yBς6�|�$�/��I�@�3�0>yB�x��ڝcj<*�M�"���v�T��y⦈,ۖ7�Ot��|������?���?o^&q�n��U�~���q��XX�8�3�ޘ���	4x]�P��Nz�v@r��M��@�%c|�����	��
\ј O���}Gl]3�N);��'�1O?���D�z�D\Ҩ��+'!�䒘SK�@:dهk4�B#��}�8	���?�� ��G��h
e�:xA2�����ɑA�g+Ο��	��\�I��u7�yG!͝j��u��D
����EU��~�J'��>y�B��F&�,�&�J�knN@�r�\f?	s��mx��ᥦ�2x��pC���~*���D岟��Ӈ�O����W�&��y��� "(���%"�0`!�D�<�5�OBZb=4�\�~|�uFz��iU;w�m�<w�B���̊,OJ6ay�aF+R�����$�	ҟ���*���L�I�|�W�?��qB��\�F}�)X1*Nw��� �~Uj���'�:� d�ɤ3TL�Qiʡ���)V��3=���jS��K4�*���T�(��p+�7��O�TB��'K�u�XBeR�5��*X�j$ў�D�`*WR��pqC�8<E�!)Q��y�(�2Et���F*_"/�&�[4Ɩ��y�h�>i.OP���K�Ȧ�����O��Ց2��) t�Y�b$A2����� )��'F"�ĕ$��T>�b�h��Im �p0�T$K56����)�:DG�D�˯^`����(S��l: .���(O����'	�>��6/�&h"`���Q�SM�ٱ�;D�ȁ�)�C(n�5"�&	k7�9�O��&�x�է\�?�eʇH +l->�Q3�{�x�rD&�M;��?),���#��O����O� �#}��@r��\9���u� Ym�$?�|Fx��.04~!���*���1�D y��Qc �)������fq{���:r%�AP0k� k
���u�S��?�td@���9Kw�@�(��%�
m�<� D��
�.��t���P1[��ɕ�HO�"�L�)E�Y�hULL
%��?kW����ݟ|+E'L�Y������0���D]w��wR(mI�@J��|0R����ԁ�'C�K�q�ą���\�`��r��o���Ug�p��	�Q��)y0��$\�X`��!1"�	�c6.��+|O���ܜ	�(� Ƨ�.�֙!C"Ol����+-��@B�ӜS���a�.Ye��������ڦ���ΐ�GMFБ�o�Y�`���\� �Iß����=������'z������l��$m%��ô�ʹ@�J���<�O��J�Q�`�"Č' 3z�!H����A�%�OL��'�\�~T��ϲ{b��[����y2I\�}lV1ɤFܗrC�d�ũ�-�y�
�n����/Xke�캖f��yc>���W�x��ߴ�?����	KtAdh��Hν��T�r.�`	�$�O���OB�P���Opb�ʧ`~��s��;B��5K�$�2T� Dy�c��蟄p3��Q��5:'iׄ+^�8z��I�%���0�'1�4Q��'�\A���ǋo�ɇ�5�X$8��լG�z�B7�˃PUX�����ē��,�U�
~^M�E�^RlϓG4�}a�i�B�'哹6X&��	͟|��<�
�K�ցd���%A��d�p���+��<��O�i�U	�pp�)X���kaH��]�n�8"<E���o�������'�A�cLGj���O.�?�y���'-����W$l:��p��.2�� �	�';�|	p��,,�*�.U�Cj��O�pEzʟ21:e%]��9�ѭE�Tz0���O����3��e�b��O�d�OX�����ӼCW)^,о��6)ܬ!�jђ����R�>AC ƷZ�Mb!���#D���g�'	<�01dZ i9:}��B�<c5��(B�ϒ#C�3�5+E�M�S�����d��Yu*�����.���sD�#=P��TT?����hO�˓D�Hj��	�J�C Wj�v��ȓV�mj)��Sm,���G�ve���B�)�/O�����Y2H�16*�ٰ�mH���ہ���T�IܟT�� �>q����Ḑ=�p��I�8�A냑EiH�wFŰ"v�i(6K2�Od��W��CC�5E�Z|듃�(]��,�Gc1�Oz����'�b�ٲ"Q0]�2N��jT�	�N��y2i]}�1�o^�x�.LJV��yb)��\�d��`)¹h���x���:�y�9�I$-|�u`޴�?������[ D�h�gi(��`����[~n��E$�O���O���&a�O�b�ʧ2� �R��M�+p� ���U-�Gy��ݤ��`P��C���"Î� WX�m@�	�h�D#ڧzn�����uԀkчܔ)W,!�� ����`9i�ʤ�`�&XQ�Y��	���+Մб �c�N�b��&|DM͓��L!V_���	\��ƗNR�'6Z*��T�-�48�! Ab��u��I�q�F_�z�cS��)#��O����N	5z� `V���'b��� X�J�B����Q��<h���ן"~���r�ȡ�V��p���eK�(*�'�ɟ�Sش��)����˓��P� ���g�H�w��2l�8�ȓN����A�MG����K�<A2�Dxҧ9�A&�I*{��XpP��gv"�Ac�-�.}�	͟pI��$]�������	ӟ�I]wNB�'�r���U s�K�B�pW�`��'��)j�+}y!�K�=F������!���~}6����?K�Pq���K0�|hg�V���I:BV�#|O0��5$�,n=L�r�捍j�h�"O��2a燖H�y���,CHt�Cj�R���������0�o�|y����'��`:����˟���П��	�u^��	ʟ��'CU��Iɟ�!Bi�VY����F�`|ԋ��.�O��Y��u�ڝ#��נ�4�j��+�On ���'��I-��7C�!ͼL��Q�y��$^�9�G�2M)܀H�K	�y��0?4`b"�H�J�Q� ��"�y��9�OTh�k�Jl6��C)%6�q��"O���$Bہ5P�tb���ߜ��u"O�X�#���l�gꂆTg�a##"O$u�"j�D��%�OjXu��"Ol\��o��z$�!��ț�jv��C"O�  Ը��		0\���v"^�j�r���"ObL����+C���BE�	E��d��"O0)�s�_�1r��Eώ�H�(��""O�e+ǩV`8��M����!"Oh�q�P� "�L�с ,�t`�W"Or� �%B��>�7� 7�����"O������^���;�.��ށJ�"O��`��E/D,������N��6"OzT�LM�0����했Q�`Y!"O�ը�g�,D��`��2s�R�ڠ"O��9�!DE (�����5y��Ҧ"OP%�Eڂ,� ���I�6{�Rle"O޵���;eu%��M�T�
)P"Orݹ�*�L�F���ꚢL�8��"O��XW�\

O�P��H�|��U"�"O�QB�Xp���H��/m@�9�"O��R��׻F�郱,�{��`�"O �ksJ�R�y��jܖd���;�"ON(�7N�.M�B*�h�)!aP5sE"OT��A�0B�x�%���w� ��"O<�Qʌ,>{TT�G�/q��!��"Obh J�|G���3^�2׮a@�"O0���`�:� �P�$ߞ��"OVxF�{.m:Չ7\&$�jE��?�M�LJ�Ū����pq�ݟk,\5T�8"
�F��x!�X�����<o��	�jR�|�=���`�H cg:u��4���q��]�Obtk6%F.c��\7I���B��|e�
	����eL�&�Ac���d�p��I:e�9,�nD��Jm2��g̓S8�A���!���R �L�9QV��3�C9�~R��"a�̋�Z�0(�i�K�{����@(�/�\�ͅza��� Z8Ib���'��]FyJ~�0":}��`	Ѡ���ё�_�I�����S�.�>-��*C��4��h��j�^�!vO�Q� Su�D���O	CǎͱD�=ml�R&�Z4X�j#?9rd�`�>�kg�YU��0Q����}�@��*M&	b��?d��8�B%�'Lt��X�[�L���?Hls������Ů����"��X���Ũ�q}L�5a�������̉�jG,�?�3�ɗ p��M�V��Ƞ!�>�D|	��<	'��(\{l��'~�@1�X�\��԰�)�37� {5Ȱs����a&\-K��3w�'�EyJ~����/�Mz�L�*H��H֊�=(���ɛ$BT@���'w���V�pY�CB�.lMK3��;}pa{ҍ]�)�ʓ"�xl�v+ˀ.�x���+ϪrÄ�aش��<)e�G�e���H�-R6}�1�?V]�ĳd�*4H���!i�P˓n��u?����+$ A���xp%���#?�3}�`�����ܰ�J2D��a��'�$I��C�/pcP�fɋ��T�C�LPy�S�����T� 3�(��TQ����,�
2
j�,X�D�<��nЏkM��%�P�6L�ʓ�0<�M2bB���Aϊ0A�e2�C�v~BᓾU�q�`��:-v�HEy�'v`V5 � �"T#�D=���E��=Q�C�S�d�T��N��H��dp��S�C6x24I5�l��Q�)Bk�\��P���C�!3SX4���ՠ�X9�+�t�k�~⟘!��R��BG A�k��:b����L{իƃX��1�Ne7�E�Z�bLITe�:45��<��@����� i@&Ef������.@�Ox�ɡ8��LCEI 
���Y�`��.[bVXi��Ьwj�캀`yi�T�$n���?y��8�S�3b���鶩���j���9]�b����*��F�7��`�)��?�b��:��E*��C�-�d�3�[Q���>I�̀��a����FǕD,�B�(�����*ܗZQ�����k	X}J�J�1hY�ᘛw�\A)giV�
BfM:�(��X�B��S����I*1V�D|r�_���x�lY1'�*p��(?Z��Q6
�>!�D�#}D���O��`l�s�����󤄁ZiX�R����0���X�B:+�JF|R#+ʰQ0�Yk�X�'��M�3��;/rl1emڝ'6XY&�ɔ}�~q��*�O��{���4gR8hZ���'H
V���Q"�ɓ��Ė|�R��QD�2iΞ%�����&��biT	4�!9��`܊� Үt���Ĳ���I@�%�$�DA?M�|�$�Y�6.nA��B����E{�O�~hzR�����)��w~� ��iɴ?�j�x�*'ԃR~�!�H��JQ
^H�'�J��]1C�����Ka*zĂ�K�T�0�fJD�ʁ'� L)�`*b��;a4�}�'89�2�Z4�e*]K4��2D��O�DhGy�C�r,Z5�a"M7���6L����d�@���tf </�hT���RU1O�*Ц��U�m�\�	�f������?iU=O� :pJ�]�E��G��~���࣬�$���&H���x��,~JQ�P
�$AG���[��2C����F�ֆK�E2�K_�%,1�'H�,�jl��=�O<��4�z��M�PL�\��'�	�Z�RD��^���$��p���Z��-+�B�I�f-B��m�")��c4RN�&4b�X�(�鼻pb��_��qQ+&q�ȵ��i��R96�1��9O.����V0rp�mԬ\����V� �I�3���qz ��\~�)���~)��H���J<�<�3��j�D��
˨��'zD���0T�e�Y����,�cT$�)��X�̆>+eH�� ���1�6&ЭuKl�V�4<O*���+F�[�)9AN��u���·���Qv��Sk��Y�gYe�'�Lp�	G]6N���� \=>Y���':l���M�A8�I,"�.�`ǉ�3g
歑�E|iL� ��"}"!ƫ^x�'N�Y�'�L�]�XpK�F�bT�,8�!4I�ޓO�-:�)	s�b>�${��(�����P�會|�y���u�bH�L>���>�L��ug�yc�#���?'렍�7oϦ�6�b���4I�
�q�*}�l�O\5�cl�q|�����Ć��d2�<�9�+��p;� pe�Ei�jAb[�����S�rI�S�'x��ҎE�)d(������x�TP� �OH�#�	�&��QI�;���*�q"�^�iE���IŘo���c�'��k�j�U��#�]�
�}!�Ɠ�P/.h�Eh�M6�d`�/�<�$A�e�4�ږ�=}�A2}�'�7�<\��g]�2	t軐���b��8�P�(�$M9WE��s���Ku�	S.�.=��d��H���%�p5Vߎv�d	�Ɔp�tSN�@�N���� H<�ڈ%?7���J��j%/�|@����{��I� �ُr���3	Ā�0<љw��@�FbȂ;�f���A+%(�u �Oݳ2W_�Z(C�HSd�bW��\��%��o_+6� +��I-'�p$Q���=-�O/���p��=3U�| 0�N#��(��'w�U����4{`}@��7y0�3'd��d��!��l��҆�!��<�슓u�Irj4}Z��*n�[�H��@ �6��k���P��	��yWxI�j�7R��+�(\���>I�ʗ�_���`M�V�@ AJJ�d,|�$��-�D���8��@�KV�b>93�\?8�����+ϕ�Z�MOL�2��O�����Z�	is�'�󎈆JP%�@dΉ  3�)�,53�I�T�O��J�	s2�P7���ΈO"���e��@��<Zv�C�{1[($?y��Dg�ɠ/��{4�U�f䤟�`!K�2s���Kd�H�; �ت%�621�(1���7	,�tt��]5,��U(�ꆋDF�U�D��G�Dʓ[��R!�3������gDU����/���D��F�8��+9e���r���2y�VQ[��`���<.���t�D5P.����4��6��\�F�9l�4���m�0q�����~
��O�P��J^6���r!#��Xj%��'5x-���+]A|�ғ�d���W��ؘ��f����WZ���u���1|�lYs�t|�2!�.\/:y�/߶ug��Bï�SRQ����^#">4p��D��9U�;po���v�!hP�ϫ.�7�Nb�>50D�@��ɽ1�<�Ԁ�p���!BDħ	NL���ï ��yBL�G}��F'^�u��˞�nM0q����U2aEM�ٱu��I�ހSW�^y��L�A'��9LYSǊĆ{�\1i�m�"Jb������<)ge� N�b����F,Hm�.��W�Y�0�IFLԍ��aR�z�V�0`�f����d��J���}B��F�e3��4 ^'?����֋�C�;����҃�#oneX2ˊ>��t�W�ϟ�S3*�H�	aKZt�6-����
(�"5�=��g�
���'��|��l�`�lM[�jV"(���ߧIJVQ
�Ɣ(f$��	Q,�?�Ϙ'�4��[�_��tl>z0
b�[�``���6,i�@�5!ޱJ��q��J��l��.�O��pH ظ��	�"*@��w<Y84�v-��s���$z�tH�~��)E#���ԋ8ɮ�ӗ��]-�Ź`e"�$Q/;Z�w��$Vz�#/�55z��>�'`�8:o �`kӊS���z�o�u�'����rG�b�Oq� .��|���b��@6�\]�/�/r`B�ɳ"�h
eQ���5_qџ�(�HD�+���R�GX��X` @�"D��v�ԟ��d�����p��� C���DHx�A��_�R�$������NE҄�7�O*���$Q�9�p�u�,6L���=O���'���f��.<]*���\>7����	D����Z6 H�l)�Β��0>Ao[4��ɚ�"��`�׮Tf�7Aߢ4����'�H6z�Ha�S���ȘIz�%z!ȣ��W��S �� X=Gx��'��D��DY��@2�S&!�~5B��0j���)d�:df�GTo:�bH�X�џx@'�̈́}3H�#РG�Af���H�'4"�M�3��:j�����c5��n��Y��%��ύ�鑤i7(��	H�L���*3�1_ B�	�i���o�>����'�$?���z���ˊhy�i��'�)���i�~����/�f��矴3ҜM�*��g �8�g��p=I$�'@���C匼;^����ֿ5:e:"�X��8w�	Y?�!���!蛬3W�����Ɵ���J�0S��1O���Z�NX�}�1O�X�FH�=6�e
7��+y;�x�����'��y�j�!^�5		�\ӊ�� J�g.���)� V��&�n �=:t�d�4���`E+)�x� ���'�CG���i\ yp��CHbiq�O�#&N;A�@,O���y&"OȠK ��m>�,ˁ�� ��-�ƃ�$H���iy0��`�e���C��O�-ɇ	��@K(,��'�\���N�6�	�G�k7f�����'͕[�^u(C�q�j�u�L1�"���P�JY�L���07H�`t��-�4�>����?U���1E�q�����k�n̓1����c�y���P��Y-}����Dp���4F~؜3�Z�i�l��W��jl�"�ݩq㬴�
�Ex�,؀+ɭU�<\��R�w��SXO�6�Itg�o�"ūRh���G�+�x�-Vź�gDm޽�G+Ŋ]?J�:���i����)*D���#11���Y63$Yz!�� ��1PwH ��e2E��7B��sQD�օLA�b�p?-2�.�Tn�$�ia`Ǉb|���D���ѣ]�l�V�Q04�2C��Ӣ#��e/��(�B�"�d�:,86�M�v2��V�I@�'�l ��6�$��%� �<ʍ��ΡX�| ��l�l%��-� H��=��� X���bf�t�@􈶆ʾ~N�p�p�Y�l���I1L����L�?�~-9@��*c���D�
�xD�9���ϢC���0��N�����D�3_~,o�~��_jl QE@Q�lU" AW�@]$C�I�d�1J�|�JӁ��o�`EJ2�3D�Չs�|�'i�ԋw��]Xz!�bf�q��L$D������Ől�B"�OJ42��(I$� �N^+x)X'N�	ܘ�Yb-<��d��$qan��lp����*�Q��(�FѲ*ڜ�� �C:R,H�P�%"�1V2�hN��jZ���$�S�H�R�-R�r��@�|d�rC��u��e�ܞK4`���H�
w�|b.�1:���R%눙e4�-ۇD�4��<��)�+2��[B�˒=�D�Kg&�z���<I�wHP�a��#d�� i%Ɍ*� E�	�'S�x��#�8M���2����7�7
�j@E��;#�.�M�'B(Q�ę?�]
�$e�c�A9P��'Ƅ�W�C��:zs�Pxt�9H�)�!��c�6��3�Gg��Q�L���B(9�b�?=DzB-��^���k1�N2."�ʁ�>�'(�#od����-N�ı&*�#���Y4@�!�$�8UN��L�;��mO��}������j��>Q�� f��Q �&G� :r����1D������=N�U%�c�Z]S�"d�����������vJ�%Ȏ��A�ޭ��i��Ά�y�#\2@��"��ZO� ���Ě ^�h��Ğ���։V.E7`����X��!��H��!�g�I�J���9I�!�d��
�ȹ��ˏWGDh+DI;A!�$�� ����
�;I�<�ႛ�"!��1>�.-)1Y�c���a%0!��ԞE���!�ݑ8L��bA��!�D�X_~�pB*ݮ^�4Q���O��!��c��a��KIE(Ea��d�B䉵H����X3��d�up�C�	r:�07*@�+p�I儏z�C�	�Z�l�٠�E:h|^�! ��5�B�Is4����D[r����5I�\B�ɾ�I��%H�p�N|�� �[�C��3]�I�D�K��S=]�B�ɐ��xb�i-�0�+���#rw�B��5ZN�m؃,�c���LJ
׆B�	�
�mp�Rf� MXc�ƍ5��C�-*PX]J��ٰD�ʬ� �~�TB�	��p,�BRc��-�c?B�ZC�	�D�PY�$� 8�A_(%�C��1.nb���lK$AC���p�ݍB&C�	) T�e"��DLơbc�<$C�+>�
2��~��U!�g�3A�$B�I����2Ɔ�kxE�va�mH.B�9�^�X��ZՅV�K׸B�IS���i���=L�6!ȄK�C�ɼSO��hri
�!�.�	���~[B�ɉ3؜-���C�l�%3��
B�I����s#U�ExܽX�g��>C�ɼ�0����u�������B�C��2�@łq�R�G���ڷ���C�)� �@��%R�d��G͞�@��,*%"O�\����(Ί����\: ��"O�%�!�[�1`�E���Չ8�h|��"O�P����_Fz��`�2���� "O�M��M�S�����D�[%� �"O��"�G'�<�B��6�r&"O��:@��"��<#b���F�9f"O8�е�R㮭Q��cw�i�"ON	7JXpt��o�6]��͓�"OJ�K����h�!D��"OTUS6I^P agg�)����"O$�+�R+*�) T	I?~�,8V"O�8 иIZ��uH3�����"O�I��@?t�)p'A�l��l�a"O\�b���C�b�JE��8p`�h"O��J"Ǵt�bϊ,#�n�S"O�a��	�wR��Ӵ�L=t�~�ڲ"O4�TK\�L-`a`�ϐ78}x���"O:`ӂ��uĸr&iM�Os�q�v"O qA�W�E����9C���}�ȓQ���z�2y?��)�O���D4���2����L0�r�Vc\5,��wx�E��ґC�P���02��!3v Ye`H-]FJ�/�5Q����� �hhB���H����]�|~�Y��J����!�	~�ja�$!*Q}�݄ȓc���I��Ԑj �8��"?�5�ȓH
]�Ĕ�J�t�kWK��)ü���v��\�f� 9,�e㧭����$��NL�p ��E�� 3o��{��}��S����fy�̇^E�Ш�i�3����֭5D��1aW/HO $ӔAô� �2�4D��y"Ė&C�`�5��M>y���.D�\���9�i;���y���ѣ�,D�Ҵ�R9I�P��@�Q�G�]��m,D���w��=*�5T(�?D�d��I&<OV#<����K��!����X�0��'=T����
�k��y*� M�8����6D�x�G�/ �*IkS�H���<j7�'D��������k�NpSP )D��J[ `��1�C_f�l�qDF%D��"�-�(w*�ci9N�48;�Ɓ��hO?�d�
~��CW:.�n��B��k�!�D�O��F�%��J�폠A,��`��iH<9P�C�|���68��Ո���a�<g�ZT��P��jK2^�F����]�<a���J��z��.�ܕ��@�\�>���Ex����B�oSV$�gl�X84ѡ���y"Ɇ�1����>I�Q�2���0=	O��h�'���Rv�ß�>��M�!,�Lԓ
�'Q�]���Ӳ>�p���L�*)�٩	�'��u˶��5#P�!{ .�(��)�ϓ�O��g�'������%���Q�G{��	F"q�j�'HP�bp|Q*�b�L�!�d��oز��p��+�v9a0�]�x�!�d�!�,(���h�����ǎ<����i$x�;�Cߟ1^<b�e�K��۔H/lO➜���:P�I�!������
*D�,{w�H4R��Pe�'&P!�#��^�����h�Z5Zu"�4A��`��%e��C��<<��ꈰ-eD0���rBB��V9�I� :�������%A�>ʓ�M3d�2|Op��`ႋȦQ���~!���'����&'��as�Zmz���v(�5t!��O� �1+T�'�b���
y��P���Ii�O��	��,
f|�M��. v�II>A��9�S�S����kW�Ov�{&*L�K�X�aP�#D�`0A&��Pؐx�+	*�H�iSL#��<���]xRre��� ���w�H�<	p����L�i�|�}�%_z�<��o���}@�)�	P�T!8��s�<y�Б'`���r'��+1K^m�<�Sl�cp� Z+�	NArQ�ri�e�<'�<XA��(�CΊ04t�S"J�5l�J�����V�6SE����P梄��y"�&ֲ��FB"z1�96(�/�y"�T,!�T��K�y�h��ˆ��yr����pC�#9r�0���E3}�"C��9�ژ�aDX�#�f���e�:F��d1�tY�����;P�8"�9df�ȓ*Ep\i� Ͽ+��%j�EW1dw����r?��
�4|A��a%O�Vx�t�ȓL��(t���^<��y`���w���<ߓ[Ī0H�Y��"
+D��i�ȓ����d�72��	  H�S�r��ȓFnd��*S�l�N�97%�>"�Pم�	0Px��ɾ|61���Z�\�G��Tc
l(��%_N�T��!T��C�Ikeh	goW
oPJ�H��V�h��B䉶�����X�fX`HyS�>.�B��;�А�%��w�13��[����LF�9Opd�%_�)��Y�n�^���s�"OP�R�(i��9�c̤������Oأ=E�Ԩ�<gc��a��1e6ph��hā�y2Jc��s��C�P��aZu4�y�a�HN���)Os^|"�ҭ�y��@,h$KDDȲE ��Btbۊ�y¦ϔa��e�8h=r�:5fҐ	!ў"~�B�ֵ8ԣC6�}��E��H��ȓ8OD4JS�Z0-��Ȧ%2���S�i#�������e�P"�X4��A"A!��04x�s3�Xפ�sP�K�\�!�DO�~\"��� �8d/>)���8��=E��'�Y{$�ݲFmJ̙�	�W���'/��4�G+}R�`��I�	���$'O�h@�i�.S�&<	�W5���I�"O~��S�>�� �g��{���#�"O"�ڰ#+$���
����E�"OL�KǺ}���3 eJ88��u�@"O,�A�Ì�A��1�B��|$Jp�"O�A�+C
$,��r�F�ȅ"OʁC��a[��� )��1[`"O��wdQ�!��L��(�0���"O����ùE�la���$#ո1A�"O\|�����[��A�K��5҃"OdM��G�B�$�I��J]R�:�"O"}*��Q�zD\h� oA/M=ΰ�W"O
�A�����P�2`	1]�%""O��í�<fh���rH~�"O�DY�,0J�,���΍j��("�"OX%"C�]�ݜٳ��Q� )FI�`"O�M2��F�S\Լ8wH��9�b�"O�tp�ΊX�A���\ P�"O"�r��R�'-�p�@(�x�s"Ou3�ȦM�@�q�L͹���"O�I���+��9�J�$"t�P��'z�$ғvҘ�p�<+��6_e!�$No�|9�'%_s�Vh(�j =O!�� ���Ƨ�m{��9!�V9!9���$"O!
&��'2���}�5�d/\O��bج�R\�F�@�VJ�b�"Oά��-9�.�qQg�BY��"O��Y��R�.\��'-�)`xnD�2�'��O��"�*]�u���u�Z�f:Q)�"O p��KU/&�`���+��=� "O@t���M]j�2`lL?&n]Z�'f���u��Gh̿hv�8�BD��-�"<iϓn~B�R䄏;���̓�}�P�ȓ>�0�㲦��[� A�Q6*7 �ȓD�p�@;��T�
1[�]���Hd8�)�Cfz[%��i���ȓTA��[ɢ ��x�����=��S4¼b2��.o��x���<L�����B�\���H��$�4�����51`�ȓO����F���H!*!�(f�dE|R�S�K`�W@�鸭�$��{��u��U�;�B�1'�fp[WD�.��H�ȓ2���S#i����b�A@�&m(���}��@��՞qw�SkR;	
X��ȓ�L���#H��0�C���o�0�ȓSy"�{��T�p۔�C*�fxE�ȓY���Z�)6O�:�$��3L�m��O�JP4MO�T8B�ha��Y\���t�~����ƞp`��5�P.r!<��\���$�:S�=p,ڭ!��,�ȓv��i��V�h�N���U+k�4m��C�"�ْ)B4����D'd �ȓQ[�y[%��z�j$�t���f�rѴ�������'ؗ&0�݆ȓ	Vд�T�	Kj�|��n�S0��ȓ$��!�ǂ�Z���C�.ՠ$ڊ]��g�ԙi��>	|I3R��8Βu�ȓ$R՚�`׺&�:HSq,�8��ȓFO�0�`��@ +��n"}��]���i@�X��.e�w�/�ԆȓP���W�X9JSTXW� A�
E���q
�@y�Ы'銝<h�ȓ^���g�H�f�ӂ�ƲJ�|��ȓ%U8�@.��9ᘕ��B�[i,���G"x��'���/]�}Pt�׉����ȓQ�Ib4�\�d��YP�M�1@�������9! 'ƛ1��	�KV,F����kN�����
�*d�6Ɨ<f��i��q�M�+Rp��Bf�K!K�<�ȓ��]j��2	qh��͕ e�\�ȓc���1)�G�Z$	 ���C�����D	�C�7;��a�H���,�ȓ[�T�i�NK�$��H���Zk@���N}�Ͳ��B�d@�Ŋ@�{R�0�ȓ[Z�� �L9T6� ���]*C�$i��Z�z8 R��2 �R�U����=�hؚ���� �n]4G�>a��I�����s��5{ՂM3ANP�ȓ �$�6&�6p4��UO�.Y��ȓQ��L�Q���S�$���cJ�7\[�ȓ3�����G��,�ac,�J��o]Ċ�!^�	�q�I�+^fE��'�hkŦH�+�*�1�dƳN|j������3�*��e�xU!�KN�<�&���f���eb	��x� �O��4IJ��ȓd�T�2���(�l2ӈ'$A�P��n�"t��m�`����d�E$SH8M��S�? ��Ģ�`J�0$�E?���"O��	E뀛e�N�*Qf�Y��-�"OLq�קu�L�VB�5��41�"Ojy�c-�.mҹ�#��u�l�p"O)�)U��H���"&f�"O-YR#����lP�I]�.Q��s"Or��T��.P�I���W�@d�"ObX�q��9 ߢLy��� <�U��"O�9 ���kf����i�/�ё"O�[%��8.�
u�. D��qP"O�)z�bzxHl�q�F�89��"OfCӋ�=�PAHfmN4B)�TR�'�z��#�ɮ6��h��iYx�qC	�'Xt��Kɽ�2����~9�<��'��Q�tK4}��)h���mo�� �'R��I�n�I�y�>g��� �'8��@�%��M�E�ʅv��y3
�'� ċS�"N������j�c�'V��Xt�;Zxd��!&	2'��K�'��R#N�C��IBQ-�6�N(��'l�x��i�����"UC���2�'7	��^(L��Ē���<�$(�'x�����pV0����/���'�f�F��u-Ysa��t/�И�'�>xx@ڀ$}P)� ʎ(q4�)�'&|��q��$E��YÅ�-d��(��'D�l�B�̫t�ȹ!�ھ��%A
�'4!b��}�d���.	g8k	�'���[�ˇCw8XBU��' �T�#S�L.�,��޵f�P���'�6����[8��Ihvh�%��'��`+ �?/��y��gAp��5q�'@8	�����//N]�y�|qQ�'v=������I�<o���'��aI�O�%��� �h��c����'��k ��h�0 k§J���x
�'�<������<z���1a��'�tѥ�ʀw+�=RPŕ�|qJtP�'��h	�#�U8\�7`K�w�Ъ�'I0:�e\�eqz}�g$пv�V�@�'����Dة Ȥ�膡L/{��i��'�v��6��%
y7蓷?��k�'!TI�t^���v.H1����'Jq���I�BX\Z�ܦ%��y�'6�'` g�l�aB��
����
�'����d�0�4�0�����h�'��l*ŏ�,�Z2�`�N�1�'o�T:�/��I,��рe�?���A
�'�raӖ$P��v��-ЂU
�'�.���h� O�� q��������	�'��9ru�[��b�"Um�3���	�'���`�d��~�� ��U�
�V���':�3�%�>��I7K�0	,`�'_ �+��+a0���)D�s�Q��'�D$��ZS�P[����jɒ�0�'|�M[�냋,��h�cύa��q��'�Θ������cD蟅R`��'��`�w)�6N�\k#(Q�V���'���`��� C
V<P[,�	�'A��*�d�N3�oܙW�ʵ(	�'5�5�gB-"c�eЄ�� �*MK�'=��1�*a��$��u \U��'-,�cgb̗{+yj4��u~-S�'��pC�]"%�Q��^$X�q,D�� �mK"�A�:jD��G��b�j@Ȥ"O���v���M�������C�4		�"O���B&3�ݨ@A��!KN���"O����(3޴a���8S+FM�"O�|2Ah��80��#NL�' ���"On8�&��-��� Ն��X� ��4"Ob�ȼ,A�(p�����"O�A"�
���գLJ����"O��#)a�@�T�Y�4����"O�Q�t�S�fX`�$M
]:� �W"O���,
M�D9ࠬS,�\�7"O}1"��*\$Z�B��I�Fl�1"O���R�,9�V90ؓ4��`"Ov��gg����d�6-Z���ٵ"O��H�f�aFę� �
-�:��1"O�1�E�S�& *S�t��(�"O��#6C̅P��
RMB�cyn1ce"O@�+U,�<�hA�G�̂ag�Y��"O��P,F�*�l�X�n��L�"��"O��"�v���5+�$,��A�"Oxxs�$����S={C�k�����y"�G�u省���������u�(D�yQ/<1�:a��"��+���f)D�06ּb����h۝l���锁+D���F�Zi�=�cX2<Ux��"(D�$P�f;z�A[�eT2v�f���%D��C�"P�S܍��G�7	m�1*Ol]�#L�6��p����_Lf�*�"O�P��d��Bq��Z�%EEF�izE"O����"��:e��H
�9*0Lt�%"OD�z%�Ȃ]i� :��F�>;+�"O2�Q�,�(x��� 25�!b"Oz�c��I�&ᐙ"f��	���pe"O,��⪔3-�`���e��V��Qq3"O$X@�g�
���Hs��v)N�:�"O­���&F�"7��a��$��"Oh$0�������@-W����"O���/H���`2`�3^M ���"O.���3jEᡮY3�� B"O����-��#�,k��,I^�ա$"O�Q�PC�@�R�O�:n� Ҧ"O)J�`�D�YzЍBG�����"O�ɲ�Q<0�($�sN�%+H���"O�t0��,�@ݪ@��
A.��S"OF Z�l���H�u�߬4�ͻ�"O| Ca� �{T!��j�B� R"O�����Q�t��2F�8 �w"O�Ճ�f��OO�݀��V�@ *�"O
y2���W�p��f�P;R9��"O�(�BK�_����Hň
$L���"O��sq�B�q�IX��̃`��"O�x�a�E�@�G���&�Qp"O0�+U,�Y�p��Ӌ璕s"O�I���Y*D�Fh �O9?N���"O,Ec���nz��c��9Y����"OI�V���N��aJ��:-��"Ov\ S�7n��Z#��"O;<dx"O�a�Z&ݚ�J"��#q��la"OF�����OW�����%�­
p"O�M �+��B��Z&�)�D"O晐�
z0�
��Ӿ.��ys"O:�(���Q��JuI_�0{6�!2"Ohu;�)��\�'�˱Sq
L`�"O(	Q��Ӗ�X`<(��"O� �i��C9r�a�`������"O�s��W���2����"O`�qa @�2�(�ڂ�7�d�"O$,@Տ�F[؜�F
Ŵi�:�)!"OX�i"�C'/% �Y£J@.�Y8c"O2�&	)��1�t�5���"O �P� ��d�B�#l��UX$"O4Ű�G(_.bDBϧQ�8e�@"O`}�a��0���U
P�V-�U��"O��Y��������c��<��"O^�:�-ΓTt���������B@"O$��AK�*:�T���M5���3�"O<9��Ă�q�r|YEy?�]1�"O���b��[��5Yg�?3!b,)�"OL��L�%�T���	��I�g"O�u��E'�t�
���1+x�"O�(���Q(F�a�w
�|��`"Oq�����H�ǻm���"O��a�߾{���� p��-� �'*!���w�N�������R��'���!�Ծ,C.h��b�k\Ľ9A�X�1�!�d�;q`1hUI�1?�D����+!�d=}�	C�ڳQ�����Z�3�!�$1M�T)��Dy҄D!IK�!�$\#G��ɨ��F+=�����ҽ!��H%3!��_�F��6�\�!��
��)� �ܨ��ݸ۔^!�$P�z��b�䗯'f�a��ܸu	!�V {n��kfT+v,���.�!�ՇY~��Ԉ�#]lz�鏵J�!�	8m/�� �_�$q��F���!��4aF������z�*�#�^s'!�$��XD�u���
Ӫ�z��ʹu	!�D܉TRn�"D�L2����$�!!�$ *9@��`cj��M{f��-!�!�$��X��)C��Y�ב�!��7K��c�LH�$=��C7���&!�D���<�A��F2�B�. �!�33���0o��f�U�A`ݱ
�!�D�<@�Z�`@)͑5 5`,�!��0YE<���Ճ2� @��x��'�ў�>�B��w�
���DQN�@P H�<i	�K���C�$7<v��S)	gl	��3OLA�M]�u�v4{�h2�ʭ����C� [3��
%-R����ȓkQ���p%�����Bú�I�JBf�<a�C���AA��!���B��
|�<��L�$$U�9��;+@�
d�m�<�Ӭס\�T�@C�����"�i�<q���5<~`�Nj�r�c/A�<�d�/�T�ِ�@=>d𤤃~�<��Y�6������΄��u%�E�<BAk�$�KÂK����2��J�<q��G<yՀ�B�	�E�Q��<�7��$|��4�ژ#mTQ���T�<�¡2B�e�#.�,�~i nR�<��h�*C %0�␧�4Rt&PM�<��L�1I>�#���
�p��E�]C�<Ѳ�J?Qui
ҋ�=�"����RC�<�3h��u��Q�SC;�UHS+�|�<��킓z�5��"ǊZ`�B�k�b�<�e�ȴ	�>�	W�P����A*8���{I����k��\�H!X�k]�;D\I��+���{�h>N�y�%W)O_6���S�? �x��V�v���X�E�<�J �&"O�=z��2s��z�D�-�P�2"O���!B�쌲 �I�W�ȅ�"OJd�+և z��u��b��W"O�ɲghМ*�p�6��YZܻC"O�̑�O�$:BH(���)`92�"O�`9s�T�%�r�P��{�|��"O�t�g�j�"d�A4��P�Q"O�d�sb�-n��,1b�D7���"O���jO	�6t��cM�Kx9jg�k�0�'�!(�ڐH�q*���1D�PZT�ˉ^�t1��$c�&LADe:D�|��F3rL�9���RHɁC�6D�4�3dX/^&��7�	r,BeB��5D��b�C�tlUq�N��m ���Ѣ!D�h��戩&Μ:�g/~�TcG�+D�<ЄO�,�i"U�ϒh��X2�+.��Z���,�:~mB�(��X���g@*D�h���{0��I�"��b�$D�qB�ʈcD!� .(���y��5D�P��
!��1��"�)���;E .D����oU�bv)ۓ�^fＵPV�*D���rd[�*:�\��3�{`'*D�C0/J���B� �;�Dp"�(��K���ӐWF��GEӝ ��HZi'W$B�	�n~.��eI=m�@SŢ�(!�.C�I��ܢ��ʸK�~��7���&aC�I�{ ���ulԢ/9��
��E >C��R�6�3�hȼ;GhIq�´d� C�I>(扁2/9f����'�q C�!	�iW��݊X��dȝ��C�	�nZ���w��L�ʅ9v4
��B�	�n���c4+�pyte�bA7X�|��db���dH�� �fCT(_%�� �$D�KčN�{�X�  �Ҭ~A!�F�>D�0�t�_�q� X�@0����7D�@qS@�s�Ar�	R0g�̕��N D�L0�Q9I�Q
��ko���3D���$�V�X:L�GG�#,8��W2D�kwY**fn�j�
��:a���%D�ܙqh�>'0����BJYLLK��"D�@���� O4���T�ItL"D��i��0�ص!t�R(�#�k3D�l�� 4Ѐ@&��_騜�M2D�Ԛfc ��@���>Rk�$C�B&D����b�&x�ei���7S��Y�$4��Sm�*���~ 3��J0�B�I`w@q���cZ,�CV+
�]ʠC�ɨ	�v��e���Rm�is��V&B�+l�Fͳ AA8��b���|B��&~F�� A�'jR=(�#òP'�C�	9'�>�0ń�^�(db˒��C��S����.XF@�9R���hC�	SӲ�3"��9����B��8C�I�S�PRE�X�V�h ;�V*�!�$�;c�>��J����k� wq!��spʌ��J���M0�/�7`U!���s���E䄍3�*��띝I�!��ͬ^T
�+��0 ���aQ��U�!��S&��т���Z6�����k�!�#'22�UL�� �TI>Y�!�$V�T��2"�@���]	V�O)p!�Atf-R���y�"y��	�LU!�d��c�(����{�(L@���HQ!�� (��GF_�"2J�{���0ID"OXp����G@r���6-�x�"O&-�B�E�J �O���lI�"Ov��tC\�P�W�U=P�n�8R"O�1[bf�gz2��wL�?����@"O°Ӕ	�+n���	 P�xU�"O��Dn>a2d��H�R"O�q@��c��$�#,�(�"OA( �&h����мR�"O�h�w���w4��hڜ_����� D� #ZN���I�m�`͜ Q�
?D���4b��tm^��u\�D+��/D����g��`�z�(�Y8Zb�ե.D�@�2a¾R
�a�G�X{�H���(D�@+�,G� 	,��ÊW3v�jB�B�	�.X�I�F[�A(@�@B�5^� B�ɜU��}�q�½|� �.�:I�C䉔j����P��+w�9�&�-q��C�)?�!2�m�\��+��\Z�C䉚�J���˒� aJ/hC�ɰJ<��2�IJ"򢨺s��15ijC�!Cj(9	$�DCc�8�Ԏ��|xRC��� �慬@�P8�$X�<C�I1n��MB�o�7h��i6O��|L,C�	
q��6��T 2�PJjC�I~�(��t@�F��(զ�\BC��+u(�|��BǢ=���is�\�:7�B�� �UH\%u⢘��G�}�LB�I�/�P�{�*�
 >$��#�>Iz�B�	�?W2�!Q<����#O:E��B�	�tZ�H���$�%�*9���"OF�*�D��[ܡ��C�65ƁX"O̤��F:Q��8 5G�)�H�W"O:Ya���r������(�r�)�"O���G�աM���ѳD�M���"O�R'�	�1Hi�gD׊�"a9b"O2D;��D��Di��2L�>��7"O��H�FY�6�`��
�Ah:�B�"O>�L���h��dց����"O��K��>.�T��Ɍ-h$+�"O�ᘁ脽w�Z��cl�)\�����"Oƴc��X�Sp��@�K�6���4"OV)�w�-t���k%
_"B�u�"O:���f�q0�y�s(�
w�>�2!"O���@�2$�(�Y �0�4"O��J.\ ���D����d"O�Z��	{�&�x桅�A��Ԓ�"O���F¡i��4iE�	o{@�I""O���g�6?�x����<^D�t"ONq�`F,2��L�Sl?4O`��"O�ajB(9-J�TC1B��A"O�ȉ'�K�H�򠇺i(���"O�P�$��b1��3���i���K�"O�%qF!�7A�p q�@V�E�%�"O��R�HK�m�<B5��^ϸ�t"O���7l���~�R�n�%����t"O8l:A��;���Ydڥ/��ɢ"OT]b�f@�U��J��PiƄtB0"O�<!aރ=;T}@P�[�j��$�"O������hCF�W�C0��X�"O�t�⍉!{ⶅs3e�5r,����"OLQ�n�;ҹS��U:gtA�"O���f��������C��Ej "O���C�,�@Kk����=16"O� ��I�"F�b��<��
O7E� ��"Or��⨟�2�8�JB��� |���"O�I9u�h,j�ڔkNH� "OLy���5v�L)Q��ښYQ�P�`"O�$�i�-K.tah>yI:���"O�}�	�a�,`�'��$5 ��"OxMa(��y8P#p��3k��t1�"O4����=WCT�[�Ǘ$��e��"O��;#��(4D���N�	�EQ"O�@r�L��`�#�e�SV,8s"O���-��Ou~��֓/#��C"OҘ*�斺6r��	#~<����"O8����ܔ{�Bc���~|���"OFX*��h������r"O�@󣋜;���	3�٨��C"O}� ���l9Վ��J�ZU�R"OX�'Oɖ:�X� ��M�u�j\z "O���Ð<~�	F�� �2�H�"O$�� ��7P��B�R���գC"OL1�f��)B�-�E�4*`�l*�"O���A�$�{rmI�c&dh�e"O�Ԓ��ߡ;m���,B�����"O��� 
T)D��L�����!"O �kR������[��Mr�"OH�Ф�Ά8�D E/
bB
��"OfA
Q�H���E0 =�ِ"O���X�~��� -֠2��"Ot��.�Vߘ�rf��6���u"O���3�Q2%�k����
��+�"Ov��㯀5<[�a�#B%kX�c`"OX����>3a�4h���"O��`aV&G�|!�LU/!��H"O:d�4��2W�d��- �4���"O�%��#A�d�ڠ�%L� ��Q"O���4�L:xL�ĊHJ�J|�"O.��Z�A(���jC=5���Ѐ"O0�����e6�JgDף����D"O�<چ[=D~у��F�]�|� "O�T2P���Vڊ�3�ɻYA⭒!"O���fG��u2p��w�͈]
8A�Q"O�yb�e$&@@�
��M+�"ON�ڷ���y>���(=g���+��'y��ĕ6�HT�$N�+[k���c
�x>!�dLR�T�skT�Z����F/�!���:��EA��D�!�vy(��^'!��U�x�\qFfP*[{Lq1��B�!��\2_���v�[��`.܏f�!�G�$բ`ҶM]�pv�M#7MݯM�!�d�5RUb:#˝�X]�CRI��!�D�,�z5y�n�)H�@c��b�!���`���j��m6�,�$�^�8�!��K�|�����Ct��3��!��0��5�6$G
=�f���-9 	!�$�����5�+k�؀(�n�"~�!�$ܪw^�赮޺H"���ggV�)�!�$ތ?t��o�?)?�U��4n��	v���@p�B�Lh\�X%E� ���c$d%D�d1�A��$M��a\�f|9��!D���AL��dP��pH�P@�Y�%l2D�@+n��.���ѡ�9&�9�.D���s��;��u06)�#S$�Wo+D���V
ÐG�0�@���0x~4�R@d&D����]�338�:a���Ku�03�D#D�� Dd�a���H���l�g	 D�� ��`U�M�⑘Ӊ1*x�9�"O�H�6�R�/�tH��H�t����p"O�	��c3Zc�G�3_w�8"O`�p5�L�k`��H7���3u���e"O�i��I�x�2���Y(Fc�XP"On\b�E
�!6�k�mC�&h��ӑ"ON)h�Zy�0��l���Vt�0"O�yDA� x�`��@-)��YU"O0T)�U�쮘��K�q�NPҐ"Od �a,P`�)Х���A�X̀�"O|);��9b���l߲���p�"O ��	An�B9x�5I����w"O����4W��8�����n�j�CP"Oz�9��Φ8@��X���U!�qY�"O����Վ- |�����8!����"Of�XR�@�v�
 	���;!d���'c���S)j��m� =�|,J�� ��a�ȓ9b�J"�H3]a��KչsȢ���g��]�E�	<���C�
�p�!��'O<�"��)F��Y�$�6f�"<	�'2�l� ���2P�2/�3g�J!
�'A��U�Z:���������
�'�X���K�{t2��ԢP%��p���&O�y����K��Yb	���%B"O�M���4y��x��}�Y�"OZ��3���- ��*��Mz�"O�is�<-@�`���3�r8{VS����I2�N��p��2qnؘ;��ڲ!��B�I�&�2�㉜�(�e��^�m��B�	�v�8��$���^�A�P4����O֒OT�}�k��p�#�Y����G�&�X��l���[�O�$�ȕ��I p�P������8wo�5�ݙ��HJ:���C���4鈉[��L��E
�j�:i�ȓ+j:9����:�Qz���,S�0��\��h��DµA��a��!z|<�怊�|�!�䃌=�m�'#�^u��G�_��!��[=n,�(oO��b�M�8	Z!�?2qft����8��c2�ʥs�!���@��8�ÞC~�SB�
t�!�$V�qDY	��68q:�Ń�{�!�}˨�@Uf��C]��Yǂ!)�R�)�ei��jw�Ϝ'���H '>8��'2>:����y
m0��FʒX�'������Ot�b��`Ņ�cV��'�r;	�z���G +{Y��'���P�d� �Ұ��C�#��Y�'1���W`�:{$	*s��q���
�':Ɣh��>Ms�h�G�
�eI4��
�'xH\�2\�Yf�-�W��&_�X0

�'|���KZY����
���Y��'�Z8�Р��	$,�)eb�� ���'A���`G�/���'��	1i�k�'$ 0ó�(y,����o�%�%h	�'5@,KM�'��^�+Ӣ����ɑ�y��4
��sF��![Z�m�K���y�-p)���u��Iఋ��y��@�zp���,�y��r jܬ�y$�n�>ś#��r^���7�^"�yr��246�;���!<���W%�9�Pyrdގ�8��H�-��8Yv�[�<�!ʚ��杛,
�*�jq���Br�<��}[��re]� �V���g�e�<��C�QHUpE
�Zz�]��LX�<� ��p�ӳ|\��*�B+[��"O��sR(?�d1H$Qq�!Y"O��yG醕21�H�Э�B�d��"O��Q� 
3 �1�+��<����"O������8`���l�����"OBz��W3ݖѲ��W^0�r�"O,���F�k����` SBL��"O����jD`~ܵpa�<}C�"O���  �KGP��4I��;Zt�'"O|A�# �%��a�TH�F=���d"O�Ś����-�uс��H*,�"O�A�a���L�N����L/b�=��"O�P����p��4PGhW�f�ԍxC"O�d�V|�����Cv��؃7"O<�q���GoL ��|�xtK�"O��x&6) h�۔aV"Or���"O�j��˦h��Y��@��ZkL��Q"Oti�b�	5=P0���)kM��C"O.L��z���s oG�>X9��"OPE��M�)��J5~��p�_���'P���P�2o*|;� �N$ܺ�'����JX'vv��R�]�|�H|J�'�lY���>zb(P��w7rI�'��@������>.��1	'����y��؉|�d��'BM�q-�t�6�Y��y��"��Ģb w�@%s��#�y2�'�\a�.O�\���r�c� �y�֧3A��	�.�7Tl����T!�y�I��[��k0Q�z��`aZ�yR��`'Z���F�y���  Č=�y�{�.��7q�� ��酊�y�m$����*�3h;��h����y�d��:�!`,��Y Z%qS���y��ߍ2�R�H�֚K�����?�y# '���R�%N1u:�x "��<�y����[��#5n��m(>�9��X��y2E9�"P�'O��i`(]�UF�$�y҅�=)ӊ}J�,�0?F9P���y��B [�@��]$���B���yR,��Kۦ�)�'F�D�Hh�J4�y�k�
c�N ��" h`v�{�n��y���,/�0(�vU�^"D͐�jѪ�y�挽�XѸ�^:�׀U>�y�Ύ�e�
A�����N�n���P��y�BCz��:zKx@�Ƈ�;�y���|0a��݈mTI��$�y�*�1|�N���{c(��м�yRØ�Q�\��+�+m��S�V�yRd�8� -��g�>p���dZ�y�@A�ivY��l����Q��,�y�"��sr��bd� �����7�yr�/D4��Gu��]҃j��yₖ�s�(�`�N�t����M�:�y�.�� �UFܡf�2�K�N2�yA��� +kD	AC�3j��	�'+����HX5u�2�AE[\��J	�'s�SE���:��p$ڃi�h��'nx�M�5o�p��sC&i�VX�'#�Ѳ��&0�eZ�" �/{��C�'��spᏨUK&5P5)޽&�`J�'��S`�\�f䤑��Av���'!к	�	5|�v��O
�!
�'��@�î�c���`�M�UG��	�'��r��L$�eI��}��2��� �L��$�>M����� d�ژ�U"O�E�&�I*��(l�N�X�"O�њ�B^�(�`u"�6`��#�"O"8�$J	DQ��O��<��"O� -� -��T�b�ݨn��{�"O耰�I�
'�X��G�ކ\�>��"OxH(%Q}��9{SB��JF�"OrB�f�X����dJ_�nԛ&"O ��#g��40�.Z9�b"O&��Ř)BqX����Y܌*�"O��wC#0f
\�pD��gn��� "O�����!+T����"Q�"_V5	�"O�t�3�Y�29.�����KW�x��"O>�S3!��ј��y?j��"OX��2j�������U:�c�"O�`@@D��ՂIa1��c"OZy���W;k��0 �(DE��"Oh1$��SB<[�a�Jt�S"ODX!$ֺ ����vk�+C ��#"O�d��,�RE�M��""O4qX�%�&B�P�"q��8
���t"O�ez1#\l�$��
ӌ�"O�(0�B�:-f�!�K0;X6 r�"O<l�P�fA�\Ah,E�1�G"O�0[�k��5F�yjg��Y�Ty�"O�`x��$������șc��X�<�P뀱/�� �(�:Q��P	���m�<Y�K];u�%jC��S���k����ȓR�J2����YV !S��I�3���'�a~r9D���"�bX����%\�y�`��0�Fd"3DH	0� ��.�y���̴��� �%_���eܕ�y����T\J��U�txV��0�ybg�O��<��&@��t�b���yҮ2JF"���]>"�`�Ȁ�,�yr�!o�A��)�l[���>�y��C* *[c��#R Eyo��y¨	��ڒc�7� L#W���y2#��l�@��٦0IB�	��׷�y��y��e��l�	vfD�s'�J�y��Z���P4%�?�.IY'$���yҢ��	Fxa���/��!��jX�yB%������<(µ�c�#�y �S��0 Џ�&;(� ���y� ��F]��Ib..�B*��y2&Y�I�H s�Wb�$H����y"+R:6A��Α�����疹�ybj�4w��j��^�yV�M�u#��y�H�,�jL���pzB���G��y��̂�e{�a��g�<k��ڟ�y�'E)c(�@:����[�h��5���y�^�-�����M7e��X��>�y�C�9&��Q�a�� ��S�y�J�� ��E���.Wr��v��%�y�& �U�B��޸����6hS�y&]��p(���>}j ���ь�hOl�=�'ne󣇊�;�$]�@D�h�2H��'�f�@0�"b־����/Z�H1��'���#eQ���%�%e�2nԘ�'�V$ �
�~@�e�7�d�
�'TR�QDB�#2X��GR�ሉ�ĩ<1��i�Z� �A���)~`աEO��P!�ƴ{��Is��2(Ǧ�+��_�j�!�7.������Pa��S��M#{>!�� �A���B7#7��ۧF�B�lb`"ONH3��=[�t�����p!�"O�D*�K�<[�����#2�Xˤ"O@h)0���sl6�ᗈ�=*��0���|�P����S:�L�� g�츙���I�VB�I�qUN�:�H�*�l{c��G B�	;c�<��G�/%=���3XC�I(j5�2 ڷ|��H�`�5X��C䉎7��eų3���$�;�8B�I!�.�P��J.C3��lUtB�I�K,���ս	G����ː+L�=)çy�PH7��#�.U��ǒ@d���&m�*�K�4&a3Ҧ�� ~�(	�'=Tp ���~�<��� �:I"�D��'Tdዤ�Q�3��x)�+T�D�X�'��Q�U)J�QP��Y
:Ր
�'��l���=N��LQI�}B���	�'`	z��)*�x�W�@�b�<M���$�<���)��2����F�j�tL�c�70�!��J9H�0���B/�28�P-L��!�R�c
�D ��֋1�ŉѓ2M!��= Xp��
ک��Hp��ؓ!!�d\�k�L���a�8�ܤ��^�Y0!��S�*X#��L�N�˄�FE!!�S�َ��6ᗣm��\3!X�ў�ᓻC��8;���A�L=����9�!�$��%s���b���0�w%T��y"� s�	a�'�]���vAH��y�P%!�Tո@��H�(�s+���y�AAW���#͡B𢁉�D �yb�Q��r��q��Ae��Q����y�ꅆeO ��	�>�	3�/ɣ��'���P�Od3�ɓ�a�T�'T4G'�0�	�'t��h�E�pd�E:�"юFF�<1��16��h���_���"�w�<i�!ܑ-�@
����u-��C Èv�<y)_ +�Pd��MS�b�ct�<!�B6>���)��FR*��!\q�<ѵB8b`0��GllN��Fϓh�<�%-�/����^�, ,�P@�z�<�OT�6 |D�Ç�%en����r�<��PT9���@�j\x��Dn�<�ҨͽBv,�%.ќT�t�����h�<� �G�9�B9� �-j��qQӄ�y�<�d$׃U��CF]a����r�<�"�۶�h�[�M|4]#�Yk�<y�'��K�5:��B�b�6��ф?D��f�=ÐڷIM�CCI0D��ط�1!|�����͟���	-D�$�H�2~��)����uMn=��*D��c��S�
��4^-���t�؅!��U?8d~��@�(F� �̀!�!���!x!z�lC�T9u늖R�!��T5I~|�3�%n#b4��k�Y�!�Č��.��$��1B��z�� S!�$L� َ ����I���ɘM�!�Ĉ%I�vxaրTl5PPЁ��(�!�$A<p�cI�z?�i����N�!�M:i��ؑ�n7r5���1!�DAX����QK͘(�@R���y!�đ�]%�	�g#�Z4�S!��QB!�>!��I� �D�9 �-�v���x�!򄐪z;z�ᤩi�� ��Z�J��
�'�(d�b��V��آA�/P	ޑ�	��� �i��q��EK�1-���C4"O�y�T��8�NXZG'K�0�@);�"O�<�6G!C��maqG�X�*0"OX���"���(����=�V+�"Ov�x�O�Z�,�"&��1[N2��"OV�@�I�Op$��J�&W6�Q3"O�I1�P?CF��f�I�ȷ"O�̱�l><0��%d�t$S�"O���![�b�q�$N>n��A"O�A��#�� KƎ]�Wj&��"Orl�ҥT"�y��lf��Q2"O�D�%h�f%����\,�҃"O"	��]���&X���hQ"O�u��N�-�6� 4���X�"O�9[��_�53��s��"w���#"Oj���d0]�1������T��"OT�f�	�p2vau��#6z�K"O|DД�ޠI��s�-#�w"O��Ru���}�4��#��o�1�"O����G(-x��q�R7wV��A"O�M�Uln �Z�f�,��1;"O@YV��J����Ee<np�q�"O��K�(�35�4��ÓPL�e�"O��Y�P�H$e��	��; N(8�"O�(��nD�ٞ4)�i��"	�`"OĨ��`�n���V E�֩١"O�q�p�ٽy�2q	��o�4Xc�"Op���L.Oj��ߢZ|X\b"O���4��� 1�e["~�Xؔ"O"�B ]1Z̸�Mۄ;a:�1�"O� $
�m����t�	\I��"OJ��sŎ�X��1Ic�U7\ˠ"O�)�Cש�Șh�ʞ0	
��ȓl_ Qhr,�Rp$�)��N���`��7V^��7f0��-�Іَ(`)��Y���K�+�`�v��Q�<���(r�"0!L�}��R!�Ur�<�Q��1������$��@��W�<�ր�4D�A�G(��=���E�Vg�<�"��9�2�$���ƹ0�j�x�<�V�S1R$%s���}���� "o�<�3e"����mߋT�B$�DƀF�<a@߶&�1���Q PKxp�u@�L�<��-	3V��D��������a�<)sD֨+�v�W�°!zR�S��W�<a�R4<�i��ȟ�4Lr��A�K�<qdP1:�\<�U@\���-�fHI�<q�M�s2����^>b�i�D�<�`%)v��1IG���%��́2��J�<)�@��b����P�C,D8ҧ�}�<��]���Ahm�94TJ��H{�<YW�^.K۞�ʐ�̻\�:�9�P`�<Q�HF�@���u��)���-D��c�t�X�; �X/B��m
�J1D����
?E04#s�X(Ǵ��5�<D�xㅙ�o�0$!�WD�<,�[HC�	� 4��p�"����**`�C�ɱJ?<m R��A���zb�*sxB�In���K l�~��i"�ɗ�K�B�I�(�	P�	��SY%R�T{�B䉟L>P�[����8�
#�F�NtB䉝j��{U��0���s��Q)��C��&mH\���Ҕa����,*�C��
5��Ē� $x�8�CJ���C�)� \�#q�ս�p�q2 ߵ&8>�c�"O�8��Ͱt�~e�q�ɓ|/ę��"Ory�����)�m����M�"O��!���g�,x�#�C\u�|�!"O��cnǆr���횔'h����"O����F�J�JT��Ýq��U"O�8�g+	�7J����xVh��"O, 1���Q1�Y���6a�$��"ON�Z�I,C�v9ӷ�Ɩn�
}cS"O�� ��U��Eh@E�\cL ��"O��`sL�V�ӥ�X�s�N�+�"OnLH�e�0�呣\����s"Ob�I�%�1	Z����ND̲�;"OD\X� ـz������5�pI��"O�%�@��,���d�U*y��QA�"O��Å��.D��Q�T��=J��g"O�R��`�Y���̸h(�2"O�ɻ�.ͳYۊ��隝^��T2�"OvP�TNJ2N��I�W�˓.���"O����۟��1�BJ�=F:��4"O���Q��1vL�t"���m.���"O$��ѪE�'�:8k1�A����"O2͘@*�"hغ���P6%�|��"Oxy��)A*��L�d��t%��i7*O໖XE`n����S� �'�Bݲ���}��@��*7�r��'��Q�Şh���[���.�d� �'�Ш�t��629�tC���,�D4��'J�ڴ��LEƐa��9��b�'�4�rc^��^�{Ӥ4�ޑ��'f����`E(d�.y�r��B�bD:�'�@���ㄯ��`P�ɀ�:��41�'������ɛ|�(-�P�͞1}*yp	�'Jh`{��
f̭)�E
�|s]	�'$��wi ./wz	��aY����'�N���eG*t�I(1�R=Ѥ���'y&4�V�F� ����O7>�9�'�����]�R�i"_��P�	�'mK�:h�.�J��'b�~u���I�<�sʂ-4�N�Sa�
*8J����ND�<��e��`��5��t���ZSD�B�<i!A?nN�� ��;��}� ��g�<5L�H�}i��L<(��
��^�<���
�i���#a9U��ɕD^�<QS��Q�Z0�	ǶWaj���Y�<a��I�u  ё��8Sܦ@!�R�<�#B��9��(϶K�B���'�J�<QQ-��>%�����jȚsp`��"ON���F����R��
���k�g�<Y�AU�$.X¡iV�;��@8��KE�<y��_�+^j�9C�vP�@�3gN�B�ɂl��;fi�<�ī���N�jB�	����a$�o�M���r�C䉦_�J��Dµ��E�ص?y�C�I5��� �D޽O��D,[/&/tC�8@؂S��;��萒nڇObC�ɖN2@9@�O<b#:Yrf��H
C�	��L� �l��U�"���_y�B�I�V)��&q<]3�FC�3?�B�!=��Т��V�8��W��n͚B�I�3G~D��a�	����$�N	�pB䉏J��-�����T��f�?+fB�I�D�����D�y����
dB�	44P<QqH�7l�+W��o�LB�)� ��a�f�	b(�c�V%v21`�"OVq�o'+��tc�JȬKX6@�"O@�e�%sq>m#6�OQq�p%"O��c��@8V���)��59$�q�"Of�:��[	y��g^�&�L;�"O�mj�'�C���BWg	:$�8�"O ���珪"Ğ
�G7 �8��#"O(u�'dˢ6�$�ul��U��u��"OH�੕!<��L�����Lr�"O � pkN)C~U9T��`�B0�'��x��V�8'`�?8��0+�'&�١��&#N�1���7`�:T�'����R\0v�e�_ S����'���S�5ZA���%Qɘ��
�'��X�W�UTN%��*Z,A��H:
�'_ �I`J�"v�ι�V�D�?ܚ��	�'���f[$'>V� wg� @�T�`	�'� �xf��9o�\�s�@87Ӿ���'����ʟFQ�i�����-����'���u�W��Jt�ݙ.��Dj
�'� ]D��E�f5��([D�H�	�'�\�Q0�êKTH�Po��O;Xu3	�'h�P��οf�Тđ�BH�(1�'�V*ʙ^qn�p�p���Z�'��cE�Ӫ(
�z�%�:��!:�'Ԭ��Q�N�p�B�D��t�'���Ə��1aq����p!��'���3�ŝ;��-1�I�24L$�'rla
�c˄w��8"́�*{|=2	�'
0xH'MXI��q���ύRxZ+
�'%.�)�˦�xB0�>O�(y
�'�8��E.i3��	e���{�r��	�':4�Jf �?�6���C�&�t�P	�'���Y�L/�6�`�%��MX@T��'�b�1'7M��R���;�L�	�'g�-H'B��"$+a�(��'��,j�ʒ�dG�HZ I<N����''XL:�OG�܅�
R��j�%��y���8'
$��G �M(�a��J��y�F��hx��G�L�	 '���y���>���`�L	19�(��ꔠ�y"��Y���@f�7C�*�نM�6�y�o]�~X��r�,Y�:�\��j˔�y�֋4���	5�=2x�U�?�yb$�)Uň�j̗�e7�(�T��,�yB�oEx��!ɹ#w�-���^� C�ɧ�pb`	_`m�vD�bh�C��|�;�)�(�lвFY ͒C�	���<37�L�_�<X3�ȑ+Ea�C�ɱ7 I:���@�$����m�C�IW�����Tv�:�{aF��rsvC�"i"� '�ʪh��3����V�OD���F�?M@�"��~F�0K&"O��k��bվTJ$�Z�'d��b"O⼩Pg�2���`�0���� �iA��䕹<O\��fe�CV�#P���H�!�d��μ�cg�8.6��	�-C'o�!�]4B-�@�х:-"�!��4�Q�lE{*��#�߮�ڦ��j�j"O�mx)��+��C���bߺ<�tj�X�����O��d�c�7`�>��慦�y�A 9\>b�k�"\m�M��-ؚ�yBGJ�#6�t�N��)]�	آ&�y��[,`\(a.F��:4Q�"��y
� ��1���<	b��/=;�qi�"O^H��F](%ԕ��Y@����|�'P��UM�c=2�0v��n��$�
�����:'g,����
r�z`�.�m`!�D�j��p�*�y�<{1m��A��'1ў�>�HW�G�0@�]xQ�{�j��S�0D��*4��'CP�X��^uA�}��!�	m���
A�_Z-SM�,$\��'�#��3�S���O~��&S�iʮ�@�� u�t�����7LO�)���y����b�؜o�,���Q?��	�Vł��2/i**���Hq!�DZT�dۣ�M�T�"��8`m�1��B�IDg[=NX4i a��>+��ȓ���S4 Qn������m\��'���T�]��5yu
��PEn���������c
@�K�[��ā�j���� ��{��)�i����B�/-#q��C�ဈSU�v�'E�O?7mӷN� �ቀ�Ft��qB!�D�o@���5.A:C
6�R�n�2]'�͓���hO�S
�Α�¾>x��A�4$9J��D��'���*��Z*>��%	:B�\Y:Ó�hO�����Fia�Jٝj`)E"O�0�akT� K�r��ܴ=G�`���PD{���ܚ���b��U�v�d��e�j azr�	q-<\��Kњ�p\d!��$-�AH�;J�h�24� �Id1O��D)�)�5>�2\ �� ?NF�sBE>[��B�ɴb�h�*C��TV�X�"�&])�b�PE{���-��jpl��� �X������y2�?%�.h�f���P����'O��y�k�1f����!1��������y�a�2��L��@ߣ%}���c�Y��y2��)���R�B��D���ް<���d�:�� 9��Ẁ�:�Ӧe�!�DL�ް�+@h�N�	T�K�g�!�D�<1����ɐ�>�H]R�.��!��mv(-�\I� &n�]#�v3�'{*̙s�üϾ�fB�$p�D�z�' 
� ��	�A� Q`a�(� �'�F��m���a�e�.
�d���r�)���	�>�@-̌UӲ h0ȗ�y)��N<I"��2T}N��V���y�#Ud���ӓk} C���N�bB�	#j�D���#��&�̺��4i;��I��y���)U��9!C]&IN�LZ��q�XG{ʟȓO*}�E��@A��!#W=5B��"O2R��߄�JLiĂQ�ܬ� `"O�pv#��"/T��a���>]��"O��j�(����
]��}
�"O�D������JT�����\?�%iT�'�OT,�@a �=԰AB��5 ��e"Oܔ�"O�7f����:R�t��P�����ا����f�-Y��9��h�N�A& �?��'���ص�Q!W�X��e� � �"�i�ָ'�F��v�Åt� ���J���y�'=j�u���
� ����W=�Bԓ��:�S�I��>9��4��* .�u'ݡC8�{����0���ۮ�2Ux��E�rB!��K=)�xu��K��ΰ���X�!���O���qΛ�4��Pz�/��u���iP�~�DX� ��c9TT��)ܑ�ybc˥+�����Փmd�`9�c
�M6jB�ɷj�8�#�M�A�x+��Z�(C�9U ���)�j�P�iЦ58FC���� <:C�T&2�2-��aR�kqn}�"O�����J��88�Wn�5^�y+��'����n7~f����uS�lJ D���b뒵#����Y���'>D�4�!/��$ǌ�Is�V?qSQ��:D�L�P�zv9��$U8����f7D�$��Nr�iʅ@3�vq���/D����[�?�������	bU�b&"D�l�Gi�(cBJ�#+G:I�Ne� f>D��
q�E!%�Qr1`��J��{G& D����T	N��
VAO�3z�h�(*�O���-g+�{���Sa"$�&dKA�lB�������)0����FO$%p�B�I ����t��=v��4�	&�RB��>� �״s���HE*��0-PB�ɼt��[UcF9Xo&�x� "%8B�I�K��I Z����ψ/gB�	�Ҁ�鱁ǻ���3ςc]�C�$��p#£!�t{��K�Xo�C䉉D���C�<=���Y!�ݬgtJB�	c>�u��d�Lꂕȓ��'�0B�	�"*�h��KQ�f�&�b7�B�I���02��<x��1���B�I19Np�)���^~6�ٳkE�b��B䉤1�9h솜-'4�c!j�VB�	x˴�Q�/����P�L� �$B�	�5y����-Mɬ�Z�
�0�TB��>w�� &�\,h���8���=D	H���4}�Ą+{D8���)T'I��Az1ˋ �y
i�bVсv��hʕ�ڨ��O��~Z�ǁ�%��GoP^��i�R�B�'��y��D
WW�ҤL-R^Ҹ	��@��~�xb���}�� N�t���n��j&a���x�炂i���sb��V���d���y"n�"��Ěw�ԧ

��2�P�y2�8��K�9D<�� Z���'A����%4��htoƈ�e�0|�tB≓,�HЀ�MbJ�ڶ�\%�{I>���'�$9c��=�ɑTh��FY�$0��y���	w��`s��Hh�L�3���yrƟ�%"$� ��!;���c;�0<���^3O&���l��D̦�Bff��!�)�����˄Q�^9x�%�1�!�O&j���E���m J��!�X8�4!��]��1t���9�!�D�1��8�G��w��u@p�R�&u!�$�+G�XH��*J�~�2i����:g!�E�ԅ�#��0�͌�e�\d	��x��7�S�'fړ&�%g����*�:��؇ȓ<�����X�����P%��P�ȓ0�l{2�˜]^����R	 �����{?���ɀk�d����":����ŝd�<�1)�#E<&��ၘ`/���Snl�'�?�!�aT��UóaH���HD2D���n+!�,\B��b�^xA`0D�|P�&;�� 8��C�:t bD.D�aHM:�����#��l�#�*D�𚣉Œ6��Y���u����3D���F�0gZ�1��
�9-�`ӵ�5D��J�@L�.PR�7��X�~D�á'D��Z�ć�:/n	k�̛�'gHLS�"D��5�۶�B��W�M�3A�� �$D����X�UtV����L ]�yrើfT$C�n�!�<�#��_=�y
� ��V��Bq�)e�A�L+h�"O@���`��1�bMs�A�Lrd���"OQh��m�t���eV�H��"O� vɇC�b1r��k��U��"OڍɤbJO]��*����5qS"O4;U(D^�rl�d��<{���""O�D�1��-8|���]�.MP|""O�x��@,�<A��Ǎ'-m�Eh"Oֹ���c�<ܰ!!Z^ج�S"OHr����#��س�-�y��׍"�24C�̉���k�#˾�y�K�1rn�3 �ɠǀ�	R�W��yr��w�ޕ`��
!��;lN��y�폘s\��"���ga�ar�)���y���4ʨ��g��n�ND�����y�kN/�T� VaڌiSX� ��ϸ�y��ǓMjƹ
v�
=i�ڬ�!���ybȘ��Y����q�j�2!m��yҫ�4�\Z���S��0C�΀�y����f���C��M��:7d�-�y�n�kr�h��@��@��d3$O��y�e�rNB\8�M�>{̌�Q`��yR�Y�$���E��<aӄ�J�!д��O�c�u�vI�׌[�X�*8�4O�0�pF��Ew�i_�$�%"O*�@�kX!l�H1�vo�2@T(�3"Or1+�iH�{��jc-�V�􉃲*O�`��Ҍ!ל�9�e�M�
���'O�=S�&�"&�)�e�9kJ�h�'B
d�hC�{��X+�O�b���')��	r]�jhe�4e��b�'�$yCR�6f�T�-!7L�C�{�<91�N0K��b �Ì�@=(�n�w�<�G�N�>e:*ciߊs�l���){�<��R�|�B�+&L�GcR�#1ƑJ�<Y'�
:Z��s���O�u�AG�S�<������"ue��^5ER�C�H�<��-��_� K dT�L���ȰB�R�<�@����~Q
���d����	J�<��F�g�ec$@�1Y��(��$_E�<9�lm�*��'LS�(m� :T�J�<9��A�8���V/�e_���#��\�<�� 
� �X�l�*)�����C䉅@h�ȗ/��`5���W+N@�C�%V�|y9��� ,	��
3AU�z�C��&cb�Z ���f��q�;eL�B�	�@���!��)r.����#�JdTC䉙��%�N4찃�Ǯe^�B䉩My�4�u��yF�Pp��B3R�B�	?:���'�1?���V��?L�B�	�m]d��M�9N��A�[��C�ɇo)�c��r�xҌZgC�B��6~���3F5K�P��X�"x>B�	������9� �Qf�W.[w�C�	�g��M�*�����;7�B�ɼ{�B��@k/d9�3V@\.^#�C�ɔ'�0��u���{4��k�t�C�	�{��|"%���e�1��ڟO��C�	�L�(ԀP����ese���"a^C䉋]:���aI8ņA��H) <�C�I
z�P�;@�]�wN �L]-b��B�I�
D���ǓrTp$3���V��B䉍5(� {���H�CJ�P��B�� �=�D$��Ov6�D�S^!�D��?�Uٳl�(#�~��$A�p6!�� �|���cbv9@�lZ%7��"Oz�����&�1�,�(˴<S6"Oޥ��}�:K���^��f"O���1V�i�-1fa�Q��yC"O:���58K٩�J�j0�=@E"O� ��,���29�!f�B2̉��"Ol�P6#H��㗥|�������y��0A~�Ӳ��$���=�y����E�Ai����$��e� �y"�C�,��Q�a�*�I!�߈�y"iX� �J4�,��j��`F�y��k��uHb��<��삅��y��.kCfٙ[�l=� )�V	��t��q�d��6�]kC���F�I�ȓDj 
��Ǽ+��X��?y�z��	�Fnz�ʆ7�]x�Lp��X�����h��0^ђd�
��#�%	6;O\G~�ʖ�Z���D]Q��B��pH��A�/��m
E�m��C�	�q�z�A�b���r���%J������	3nV�l�(��h���
��j��$�'�B����"O� �f\"F����P� ��ȉ@yR�V�+Ob��d�4W��5���X�iB�������~�&G�4�D1�QR=7Xi���)EG�����0�4�;Q�'d^0*wCC�s�������(.g�};���E"q=,XZI�>���� P��r�U�aE�e��F"O0ذ%m�*N� @�EÑ�p~,1��ORe���.����# �<E�t-@ �B9��L��<��o���yB+��(P�N� .}���V�v�9��`TE]jV���U�v��@Y�lH@1ɐ1��bF��If��$K	h��g�3F7F�򒬔;��R�N#z8!KTC4d�b�r��٩��O���[�T9dM
%�7љ0������\*��5C��?��'Cǚ���
w�"�z���? ��V"*��f�V�o��P�>�6yL�ɂ}�lL1���	u��j�+�"Na�˓R("����.��S�'�z�0b	6nI��Ӯ2�x�8�bL�$�h�'�9CȖ�w,���&|�d�!�%3.�h��S$��4D�?��&�˶��Ej�O~�(��0_���3�[�p��ؒԉ�&U����� �x�Cb�d��KW,T9
��4NO����W.^�D�x�C�9�?��g"�b��EK5�Sf۴���l���]T�C�	�E��pP�E�C�d4I ��7|\�I�0V�YČ��oR�c'%�	jV����!dS)hmQۃC��8<��I��☱$	]�V��Q`�D��r��L�w�֓L���C��'J�Qh�	I6~�`5�ቨf �ew��<8�,|DL�@�?�Ɖ\�!��<��M�O(AJىm�p��cHG�g����Q�.*����w�׎�x2㗓c/�U	K�R�LK�h���V$/I`��퉢�y�؊>mdE���L%A�$�q��/E���#J�!�Ă[��z�H�ZDeㅢ��:N(l�F0��� ������YJ~� �;�Ĝ�!.ꡣ�4|��i�KQ�B��9LGV�!t���jXa�KL���9t��@�L���	"v�xw@�T���3
�q����];V}ʊy�nѦB��J�㋸"^Ss���y�-��^��c�����Ai�0=��E�L�z�'��Z�X.��=[̙��pmc�'n����jUfQrE����/N]�1cK>����LX�9kçX�H�BPf�!5/XĂ2掔J|l��T�
pI&.� \m��$�ږL^�xe���	�,������L<!BL�UyTo�?d���:�cIKH<�ES+Nną
4�Z3z�j���iA0#8��D]�CǨ��D��0Y8!��cʘ:�.�}ay2�� ʌc��Py¦��82��hU&\{x�����y2k�<�̚%ʈ/N��x�@\��	�X��� :!Ub�'!�0IB�=j��*"t��-�SqX�&��k��@�j$\P����Z)���U���o�N����O4as���!����KhĠ�]�/���b���>�6qG{ҍR6f�Kǣl�'5�A0�&N ~�T�y�m�C��a�,6`�$�g%�O� �8����}C`��%}��t�$�'6�zAkZ5 �fT�O�d��l����o�\y`�5�tmy��Hd�!X"+\0�y�J�"�q�jLL������
���+2c*��è�'l)��O(����&���T�<��(��<r�R v�/[��}RB�.^�Pu���O��L�`�	.��&�H<jY^��{Rd��-�\c?�$`���B�Y�3�'��<,j(HG{��f��`*�E{�'P��5�G#���K^�]e���V-D��hA�̊M�LRB;r'Bx餮�O̼�P$J&@)x�3O�"~"#ID�w�~�)d4QP���b��y���=G�2�c4;̞�˱g�:��D�:��,C6��|�N�𤋄@���Soƹ	Z�uAP��}ba�R�\(�J x��U��!`����N5/1��G�U؟�j@!����I��K-u���N)ғwHT9��ᔁH�0C��:����/K�K^jFܘѮ��9�"OL�p�˜3xR ܃�
�q�ư�C�i�t�SV��xW�Y�dNٙ�"nZ`�Zt��޻;D0��Y=M3�B��R�0�Ja��\�|�Sc���h�H,9�*/D�	�e*W;1^�	�,�?�=� C�$8�Q`	3(��L�-�K8���rmK7S&0� P�L`28�e��
B���k��d���_Ta~��	?~qb� Mz@�d�O��Z�Fɛ#jкt� �,���|jT��$~�4yC�h"4��9�AS�<��.gǊ�F�_6��u�Tiψ���B��Yk�9#�]5J������9�6�4�XJj� A�]>k蚔�Q"O��RUS ~**�����~�����)Wg6	��B�@���nF��DF3��R9g��#��`@�¶A>���l�T�F�"t(�R�h¦}�5� � �z�"烏X�0D�W \<�}Bj��#1h���!���۳�0��'�����؍Q#00�띖
<�P���i�*ޜ���ֈn��p�!�d��t�Sf��>�00W�]T�Ƙ�M#?o )��A��w��9A�I-§%�4��D(.Y��S�h�@.�:*�B��e�a����>�3Jy��x��$�$�;QaA#<�r��Ǡ�d�I���d�+;�|���R�d0 [7�A�g0�z�Y	�Ƚ0 Q6��0�N[�bx�ґv�R����Ήw��{&�,�a}"�ߜAE9p��*
��0����'�~yH5��t��j�Ȁ�lPH0��S��6C��a�O�%� C-#	DB�@Xi��/�<Cn�	�LTq��I��Ĕ�+���F!�\Ia'����O�0��;0����=$�R4"����sUP0��i��y�!�P#t`QK�!GXPU��i�z$D�	R��$h�Q�AJ��Gy�'���S)��LӌA/�yC�JM���=��ám�P�1�!��x�Hᰴ�ӁY�Nh��n͖z���[��O.5�UkvX�4���=4G�͡�&U5%����R�9��:[�8{�C�{k�l�!�+iM@��U?񪒧Z,*���Bզ��@ӆIZ��*D�0!3��=1���I�`R.L�=(F�<i"�I� �� PMa���F�v$��%d�L\N,� �D�<��	 V`������#9 ��%�.��=�2)#�gy��0wN�iV��!�E���T��yҠ�.@B�e��4O�-�DNE��y"�ɝ	[
����?I�,�Ϗ-�yR��nRz��q�Wh��0Ν�y"b�4U����[�� ��y��G�6�8��M2[Gte!�К�y­48�(���/Y���8�#�%�y�oV0M�B���̈́SUdP���9�yR.�,7rdqj�Ο�Lߪ�ʑ����yBK���|:G-��N���ѡGZ��y"5xdn��#MaP e���yB�P|��e�`*Sa�#�yJR7��d鳡ז'�4 g#�+�y�!M)X9ܑyU��V����ά�y���;��S�k6�������y"�C���V�L�:5j���y2���'E4m9�	ư,�����!�y�#��-��?
��Yō��yL�>d��9C�1P����4�8�y
� ��Q��U|����f���{�"O��1 ��M
�x	��\�\�Q"O�p�c�z�\oIR0�ڀ �"O�9���9�� S��ڠiP"Ot����J)^jp��M�"��ԫ�"O*���B�'p� y&̈�k���g"O�b�]�
r�Qa�l�&G���0�"Ot�1R	�/y��jT����܀�"O��0��+A�F��jkc�x"O<���er*xk0c�vFd�1�"Od�X �Ұܚib��;;�ȶ"O���EeD 0��y(D��I��)�"O�@���H O��`p'k�+��Y""O�̙���L����wj���r�"OuZ�d�Z	��懘�n�p"OA)���w�x�0�fJ6;�	�"O�u���B5PIXU��8>V���"O8E@4�jdz`�V�J�V!~x(c"O��{�,��Y����@K�t/��"O�	�*N�k����4�J5J#�h��"Ot�k��"�P$��-G��P""O�%�g��4h��@"B�/!: ie"O�]�4fE=f*\&jy�(�"O|1x� ږ[z��[6�˶l��!"O*Aò��#*��E��[Yx{v"O�k�.�&d�x"&J�[�l옷"Ob�rJ�Y|h�c�
0�|��"O�P�ed�24����]�`wJpR "OX ����3|/,�� V<��d"O�ax%-�5gV@c�+�.|C<	[�"O����@�g������PPC"O�ё�n�=�܉�2��g�B%: "OL�S�P�c|�E����1a�p)m D���c��'k�H����&8%	�	#D�Dk���Fp��"oFH���?D�ܘs��G?�\�WLۉ�(��6�.D�@32fɏz���W`�,���#�(D��Zr,�K�8UA"C t�{��'D����
;u��Pp��/�2(�bM D��S���h�*}S@�=.��(S�:D�
��D�7w�� �˝�o=�R�6D�pj��K>*1ġar�̔OA*��N4D�,������H@�7�M�b�,�;��)D��V�ۘyJR�c5
I�z�Ƞk`'D�\H�.X4�T`��еk[�  �# D����S�iN���@(CB�]���!D�L ����P��"`Ûdkp=Q�B3D�T���DT^�"�.��#�p�ю1D�ě��LJ����.�k)ڄ�sg-D� 15�_0i>��'��Z��-D�h�h�,��ĩ2��/��`�S�+D�43Ƈ̒��U��y�ڝQ��%D����f�E����F2#ʆ�Y��$D�����nѾtp2�Y�Qr�C��"D���ʌ�X��0ťS�j��x3�c5D��:�k�/ �$|�fM7Xn��t 1D�D���/2O*�A	�p6d��&-D�x�� %9�(�"���N�����*D��%��"VZe� d*��B�+D���b�	=�� v-J�[�ޤ��<D��Y���:�0��f�W' ���h�o;D��Re~��l��	���誷J9D����ξ,J���P-%�jyB��%D�S�'�2�<PyI�D3v5��/D�� ��3�.H& ��I��f*&�((��"OX�&�D�7k�eP�d�C�.���"O���e�*M"��Sc�[V4X�v"O|�:d�L�D��scE��'��;�"O��$�\IA�RB�P&�`"O����Іm|X�'"N�e�J�cA"Oƴ���	9J�p;�Ò�6�1E"OLu��i�Jʞ0	H̴,��]�"O�i�����$�!0߄��0��"O�p"fH�[���F>O��(�"OZa)��^%C/�=��E	�d�@H��"O�Q�ՅwE$�j`��f���7"O���&�H2���.JC~�8�"O2�R���,	ܪ0#���KKz "O�Ѩ6�Mq��ႇ�Ơ����"O��4D��q	D�JA���2lIC"O֭s�)�1H�
VBF��tU �"O��bÅ��6A��!�T7d��"O@���@�Sc��� �3b�cg�'�D��e
� �HEs��=C����C� vȢ�Oʈ�EbC�?�4�*e�2})���,8�!�)W0i��O8�T��5\8��� L��N�Q�'�8�`Ѡgl���ϛ�~�82�'�|�c.}٨)�CV��}���^�K5L�+|(H�S%��h�<��ܪ4�x�:� �?W����M���剃&�L���LW4%��g���@�WjA�Cۼ)!��������&Aa`�m0�ԡ��hTi&z���Rb΀P3�j؟ ��io�A@tN_C��g�*��$����B��Q!L|rc@-И	�" �U~;q�Q�<Y6h��*F�Qj���2_>%+ee�N?!�m�c���R�(���Ӓd�d�y��*Sz��YU���7�B�	&-�I���H-f0"Urai��y��p�)O�Ѹԉ�xH��J?O�h��B��B$�墌�Re�}7f���zi�	��pq���?7��}��d�*Nv�ؓ�\9B&j�K�k[��Oze�$I��W��>�����(��	�l�@/�M��b4�.�Q�vf�fJ���̋%�f1�(S��_ ܉���O�U�5������l��4��@~⧗e�٪���*���!#!͝���4䮌3�,����/3��4�@ҧFhdPd� Z|�QX���&"�ɶCf%�e��g�axBeO8t@P�{1�P�&pv�#�$�&��O�	i��AC�����%��x�ӎ\(m�x�3@J֟P�:K�팈S����7��	t�'�es�M��w��XB��<a�E5,H�9�#�O	��A�2A�R`�����$K3p�YT��#F��牥�y"E(("�!v&��6��.�&tW��dҚam*���`�G�j@zO~�q����E�l1�[֠K����9��Z�{|�⧅�i=�G +��8LTt=t�1ԉ�zZ��Ɏ!�TMwC�A�ax���Fl�a�����^C�u��b���O��&O�t)�J�9Q0MQ ��+b���M���sk��t� �(���� I%*&ƢR�uS`U���<��b�O��m��n�4P)�9+���}��A�e�&�P��"D"�:�j[c�<��k�:��m2De_4��I:����\��D!+������m	䒟���M<a�董j���p�:M��Tz�E�T<i�hѢ�}�E��4��)vK�$'�v����Z���?��)Jr�؀/3W�֨�u�T8�,ٵ"��]�1O.�rU��a�����T�*uԕ!�"O|trwn47��!�g�.��e�3�'���ȓ�W�$�bXɓ�H֢c@��"]�yD!�D�T.E�s��>q=,!���޴B�'<(1��J޵Ca�$,Y�,����!�K%�LYd�E��y�	��s�ҸE��W?���Ǖ�r��<)��>��ⱟ�'�$i��GC Ūh)Ȕ�4��j�'خ0�+�.��@Y�CL_ܬ�d��x����̏Tx��8� �0dF���і��l8��6,O̘3O�+:y�(O���!/��N��d��蛰rI�0k�"O*L��t�йxQ�#7���A�>y�B
HrT��#�E��ř.���π �z�B��z���h���c,: YW�'������c'��4������i�
X�tP�!#����4�3�D��Ռ�ᐦ	3��9�c� �ў��i��`g4�y���E4y撉�푿L��x"��g�Y��n�d����WD%�Ã��{oUɓ��<K����ɲ=:XQ�W&є>��?��$/�!)~>�wY�x����`i$�[9P�dK�	�y�,V�/�`���H�g�|k������ s�1��Y7�@�O�9�SM��	��xzua�S�t���R�!A��}"i� D������G�����6�<�ٗ�Y9B�r�{�육} c?�d��e�v��;���1�K�.f~D{b�پj�-�2H�y�"��a��������G"�͇�U�����d@.n�6����=脤���I̲hk?�S�O�A����H���B�E��1�
�'����$\	#���s5�V7#L)I+O�`�.�X[ք8˓K��	�3\d��#�@�ZpRl��I-9-�HJ5oH�y��MQ��J�t%ȵI%,�
`r��IX1�cE
(צe�=8���D}�B?R�D�$
��s�-�P��Y&Ȍ��H_��yrʌ�\�ʜSG'P�Kl��疼�yBT �P�QM�?��ma ��y"Ȏ�G@���V)`��-{�ר�yh=?��U(�K
7hZ�)*	�yȇ�� y��ّU.@�d	��y���u���Pc /ؠ+D&K��y�惓8���T��^{��#S郆�yBoUs�B�Y�C�^���@9�y횤yԨ�� Ê�Q��\��@��yb��\٢Q�zW�@ya��'�?��m��p���C>y��
a��_�~�	p ĺOa{�߮9�H��OV͠��> �[���Ԉ�"Oz̢P�3d.����n��:�	22���y�
��Ö�~��� ����O�șy��C�m���o/~�(���'�*Yr�Rb`��V��-Y��x�r듓 �"U �'ɺ���+�>��R5�����ȧn� pPI޻s���A"O����A�/��Bւ�.!w���O�]����`H�f/b���:\�蕏@N�'��Y�AB��9����#_�-�דoi b�AIb�6�ć�A��9�g�![�!�r�B�C�:9+��_�6q���L��T�#�%}}(x�R�݁�p��=9�@�u4�H2���O,���A��t� x(��`X�0��-v`]�+�x>U��"O�<뱇ڵ>KLM(�@�4��#��L�q�E˓�'TSϏ2U,�4�2je�u�T� J�^l(�� 'h	�	آ�"D��v���C{E�!�'(tn4�V)C"nϬD�'�%0����Ť�bQ( Fz­�6�6��P���.,A1�F$��=��a�'-�؀�'.���1�'9�����!�$����۝YdU��}X�c�'3���i�%�jf��p��"�I���U0��O��A���i`��x���Rb�R^I����[�l`w"O�s.A�`7�S�~+Љ��|.ĩ��)��DD��pf��(g�K��Nc��8D���ʃ?ʐ`�@!LX�Kѩ�X�>➠���<Q��Q��0�`�g�����i�I�]�<�dH_TU�$J��/��9���T�<�2e=Py�ghƒF��Yq6@�U�<y�l�&=$T;���X�*�r�,_�<�2ß=5��`���I
B�D����l�<���C�8��3�߆0�rx����U�<�W͸W�PMB)U�j|QHP�	V�<A��Êa6
�)�\=���a_u�<y�^�@(b���Ν+.�V!l�<ɐgӝnr�ch�Q{����jGq�<��ᅁ=P|J`HO�	�&qQcIw�<ٕ)
�̵	���Y- �@ҫQZ�<�E'�)~���g!�۠\;d+R�<��(K6d]@˂aZ�i����#E�u�<If'ƥQȆ�`3�^,Z��C Gm�<� ��Dg8�����%f��1��"O6IҳC�%�h�j"��u�! R"Of��w��vڼq���1	��YC`"O�L@G��4'��=�7%��M	R�"O|l;��?'@X(DE�2K0��"O�8����#m�J@�ߜ<
$��@"Ojy*$��teD� ���Uz]AE"O@|"! I�!$1��k�j��В"Ob���H\
l������ߟ'�a9d"OP!01�@ 0�^1犓<�@:�"ON��5B��8 s��Q��!�"O܁#ǀ�"'�*V�=M� ɹ�"ObEI�'*"%��� �A����"Ot���"L���(q,�Rr��2�"O��*Gb�U�t���HyR\@Ɂ"O<���	�\EFd���^0Q_�驐"O�������0r��3'ZT U"O�P�⃑�VKL��*�^4 8�@"O�Ȣh�
^�`u(AH_�Z/4i2"O�ʴ���K�䜁�_�B�dC�"O�Ab�2.Q� SEҖ���e"O"Ժǅ�#خ�"t��9���`"OX8���Z��6i�n ��,�s"OHyK��-��q��Ѯ5�!�"O�(Y���y��6�_3���Z1"Oޅc�'L�~\�1�:�� ��"O� �R�/!L���`�O���P"OL��w ߡg�2�7aU&="2 "O
������CR��u��B����"Or���k����s )�!2�ق�"Oƅ������\�gOԣ\�F��s�I�Wݢ�pS♒,��
tK]+8{��	�x����V�����k&e'�n��~B���ē�>�s�e� ,+����n�����A�OD�I1x�OQ?��5�Ոx�@I�M�)�N]��f��@�G(�)?��6�ԑbnS�Y���gÓ�h�!��B���p�	+k*��e,��C�ў<��ӳ^W6l17�$(�,rnim���y�D!}�����N|!B���,$�cR헆��'%�#=�}�G�#b�ґ�<T|~�:�K8yH牡�yҷiF tO?a��O��'G�L	&�vۦĚe�z��E�vċ`�,�(:^���X5"vnϬ��4`��RĆ�Q�cy�S� �A�Ow�P6���r�����ia��4��'"�p8O�?�&��eqJ�aD@��,1 h�FhV��ēX�l�OQQ�,���0�C���Q��5?�q2O���;}Zw9��SU��	,�	c�Ds��u�s) �yB��0�N�9�4��)�)O(����
'Rc�P�B́AOT����88�VJ,}�����T�r(�0 %���l]�0��)�ynb-)ߴ��uY�O�Ԓ�vݥ��imq�Ɏ(��q2��q�F]𧶸��'��(��O�b>�yt!ÐE�p]���,CXJr��<�e�Ə�����X�(����]҂Tk���i Ԭ� �+�n5�5-5z�̙�'h�P��F�H��\�D�2�K���v�4U8p��K�¡@�=4��`7o�x��� 3��C���'������:�Z:���$�,�	�-�֕H��O�,"ҏ�+%��M�f�d�x���"�󤟄j�CF�� �0|�#�K�hAڴf�H~����K68s�vI[�H��Ȼ�ϴ4T@t��'?H���4Oר^�*q �
@�m����y�D�bD�CVXi�O�����dY`B'��o����
*���լM�O?7��8���X*���g�T�!�O5~��Z�͵?�I{6'ON�!�D�HI�A�c,i�胁9N�!�Ď�b�Ћ���/�t��1+ԘY�!��E�Tc��n5hu"���8oz!�䄓1�r`"wh�
��ؙ�	�8LK!�DW&�<8��E�q�D@Re�ޅS!��]1N yH⊘y~�ؙQJ�2!�� T�����}�2�B �J�)�����"Oȡ�ւ����dȚ�
�����"O�����W�W�R���J2-N���"O.ܳ5I�"x��\����#);rmZ�"O:��e���,k��R��wr��"O����؜z�pd���?S~,C�"OD�r��A�x���A-%MB��f�<�5�V
t�ذ�Ɲ���s��_`�<�T�«�؀�B̓+��A�[�<�!�S6l��䁥b1Hh�-�v�S�<a���;a������ ��5�5�L�<ٷ���W�~p��@�{�)R!��K�<���%nNh��`�<\�h5qw��q�<���Ƚ�b|a6#�:�.���E�p�<ѳƝ�2vds�fء����"-	t�<IL�1��a8�I�!BY��KT�<Y��
���̺�˻�<l��D�<�Q �#p|�:M��<`���@�<1R�Q�)���O�E�3�P@�<�3��6��P�t�DA��P��y�<	Fl�;BnY��@�#R4��E�x�<���w٠��w��`�8#p.�L�<�@Xz���Ir�2M�Ȣ#a�F�<YT�S�;�R�C�G�Z��`��ZH�<a$g@�]-J��!�81e%³��D�<Q�J�,-��B�F=W�\�f�G�<���w�(�N��?~L����m�<9��	0Ds��pQ�;r���Hg�j�<	�.	�L�6$
"iNU)e��f�<ɧ-�$0�K�B�%���`���{�<�cL��'L�#���lQ#2�L|�<��5W�DU��I(d�P�r�JT{�<yt�;�ڣ�#q��1�x�<�� &5�$����# ��2@w�<�@S�;��H"�EW8'�t��l�o�<Id�Q�s�@���m��+}�5q�iRq�<��)T:!��%ұ"V�2�ȓ:k�i�C�膰:��ޣN|�D���D݈'�(���S@аa��X! =��!�(I�( ŏ^�U��M��(�t BKщ*K��2>F�H��qg�ea���2b)���7:.�d�ȓlh,��w��*@�D���W3-�t�ȓa����&�Ч1�)�w���
Q�ȓ%�$��#웍L�LMдj��n'"ȇ�aP�s �W�^!��S���A����e�f�7�؁i��#c�ޛ{�j�ȓ`و�YC�:p��x&�Q�m�v��ȓ�V���,	�gA:�.��yR�[�t9�`82�Y2b�B��aJC��y"�'X�
��0-+T��8�F��y�dP�.�$Y�E`.�30���y�*D�z�&A�R�
�8���S`�/�y��Ȋh�<��O*��;u�M�y$�'!ij:�B�$�ސ�q#A��yb�����!��)�buKD�U*�y�Nѕ8�@�`�H4:V�8��F[�y������t�5��d0�(�#�yk�܈Հ��� �up#Y��y҅Ǵ
���ۡ�VA@����D]?�y��C �,�a��9`p:�����y�S�F��� c3�Z�S���y«RmH���� (�n��7���y����_����6w��CW	�y
� @܁��I�Xp$BMX
V��yH�"O��C��,�L��M���R�"OTY�G�˼j�N�#R� ��Z�� "OX�J�CP\r�Ђ0/X�"�~�;$"Orl�1&=yD5��i�"O䰂#b��n�@��MC.l����"O�����Pݎu�ѡߩX~��A�"O�9�f�B�%����]i���""O�p�d	��#��)Ss��&xZ�Xf"Of��0�U~~ �����O�6i��"O����Ǵ_g*`;��G�`dp�JW"O(���ܟ3�. ���>	V QX�"O��G���~p�̗iULĳ"O�9J�����d&��s��q"O&]�`.
�Z��T/�0Q[���"O�|�3l7O�!kUL�XA8�y�"O̕�����l�KU�j�18�"O�`�ҟiJ�C�i�18�P��"O�4��K�&%Zm(�n�Z��<a"O�2mI;���SG�,DF�,�"O"L"��N��	;��Tބ3�"OH�����T�T�i�/ϫ1y�M�"Ov�����Y� hU/�#{f(`s"O�{c Z�,�8�k������"O�91���--J����HB��"O=#����@.�6OɂJ��(�"O��@�^�b�����T�J�"O����ǂr`�RE�D�V-��"OH����Z+JY*'L�ty2@��"O�]�qi]�S.x哒�T/D`TAs�"O���	��u����.Y�`�"OVAQ�X'a����w�
�nQ���e"O��Jt�6nv��� �9�B-�e"O�`#�=2j�����K =vD���"Oh��'G$a0�I�3��/jN���"O��CS(�:PY@ $*i���W"O��8E	LB2U��)�#3c��he"O>͢ �۳-H�s��=ZO�}"�"On�b6$X?g��zW'�E���1"O�f��)h���PH`YQ"O����H͂}T��"��ʸ;c���"OLXY4�9q�(V��7Y~V�3"O�%h�&pĘɉ�B1(iV��'"O1�UcF��9[ӮJA*���p"O.e�����_d�!x���5��"O.��$�~�*�'n�98�7"Or��Tc_"k��a1�ҤC����"O��[!�
;w��(Zgb��Z
�RB"O�P���t�&ف�g=-��
7"O��vo^<V���z���|�}�"O�8���P�\ 2�L�ZP�"O�ayrl���<�J��[!	�aF"OF@���8\k�` �Σ�u�e"O���g�+0���Q�5x��S"O��9�e_��5I1�ڲp��}Ha"OpC��Q�~ȩҡ�.O�����"OШC��Z�d�hH	�c�*�>��6"Ozuz4g\-~��$XsI��@��"O�zu�D�k��x ��i�I�s"OvD�@��H�4�A�&?3��Ȣ"O��J�˙�[hy:4����R4"O�����Pv�J5*˿~�RY*�"O������=Nҕc%��5,�v���"OHd��n��ҩV�58�(�"O� ��AE�/S��b�ħw8J x�"OBSa�X0=�IK:`E\p�%"O�=*��Maci�⃄E�$$��"O�u#�k	W���8���\5C�"O���E���A��m@,0蒴��)��<�a�(r�a�LD(��U�b��|�<y��*怀���7K�1�HB�<ك�h��A v/*~���Ŧ\d�<���Qg���L�	������w�<a6��
^� �C�Q
�b�r�k�<	�Ɏ�,��	r��
iJ�!k�<�c@�4k�%�孁0��ت�J\h�<Qr�[&%�4u���ғq�Pt��&c�<1d�Ȑ6M�aLn�B����E[�<�%"ۼ �d�0҃@��ݢ�&OU�<��@�2~᮸@�f�"58g.Q�<Q�.^~�C��C=*�X`u�J�<�¤�3x[�92$�\����
���C�<��	�=m.�=Y#́"����&�f�<��nx[�L�rb�?$t8�	��NZ�<�� �@��3�	>uzzX�T�QJ�<Q��`����A(=���D�<I�O��Z���+7劖L��UQ"��[�<I�����훥s��s"Į*��B䉆V{�����M�(t����M`C�ɬa�4��MN�B|
g�O�u~B��<K��)��T
+�8�S�J�=q��C�	�;�p(��/YP��r�Ga�C�	d�b��h�f�"Ys�.
MjC�I��<Ӵ�!�`��{�6C�44��J�h�)H~]�w+��F�C�	kv5��Ȅ�X��1 ��!�$�I�ِ�M�-��x+B�C)�!��^$N��D������]�!��]�!�$1~�T0BH�-�����2>'!�$_�l�zDB����]��6��#�!�$V�*<�y!���.Cl��U��}�!��&y��lY����9�C�*W!�&A��h����'�5cԇ�( 3!�8aP^M���M�9���2g��<,!�D��f?�ղ苼�e��9�!�E�4�1�l5'T:��q���4�!��	?��غf��a���Q��^�c !��po����Ȏ%�2庱L�5@!��%�A	X'c� q��L�5$!��
���=x���!���K� }!�/"W2�Hs�Ĕ9�d�y�'�!Cq!�$@K��s�ϸ}9ƜC�F��]!�DK
\����DC�F/~U�#��kO!��G�T6��ծ~p}(��#4���<!�l�������Se��y2���
e���y���[��՝�yrk7+�r�k�oH,_V@��N;�y�C��F݄e;��@!{ht!YQ+J�yr�])p��]	E��d츐��"�y�K�4|2*�Ѓʆ�O���:�I��yB�=<����-v8��ر#��yO��}T\h�� 9spz�����)�y��;D�H�!ƨ0h�^m�E�ɧ�y��38�����g���k�9�y2@�; P  �P   >
  �  �  !  (  �0  �6  4=  �C  �I  �Q  X  B^  �d  �j  q  Qw  �}  ��   `� u�	����Zv)C�'ll\�0"Ez+�D:�Dl��b=O$���'h4�l-�fdre&ĳQ�-�I� f
|��aBHX���c�HdI���fh�Q
`C��?��O��?!@�K!.�YpNZ%([��ʿ#� �:gkE�"I6I`��٭l�s�	:�u���\��D�'�py��$�=t�tM�e-�[� uI'I�{+�ő@��O  J�(m�A@Mܦ�aG$Eן���៸��ΟH�bl�3v�Zd��� ���8`�����	e3�-#�4��$�O�+� �����r��3�R�E�؈!��9D�'(�O����O����O��i�+�Ou���'�d���w#_�I�p{��վ9Jԝ[��%�OZ��+@ �;%�2`�������'��듬O��2X�|iB�?�0�n٭4�Ft�UA#g��0�L�O����O����O��d�O(���|j�wI4)�0�� h�L��aZ+X|���?�cz��l�MK���?A��T�?���/�?����31�x���d"�����9#���a��Xܓ���;@��0f�E�8�|��U)\�Yҕ�ӎc��!��Ɉ\-�7-���]��4�b��h�4HF]�GRN����{�,}��k�z��3�i�n@kq�$/�(!a�
�>x��*ՅL7��u�Bir�Lm�MK��-���:�'�.G�1�Z�^���ځ�)�F�Rb�i�7���)�0�tI�$X�.��t2"&׶|Т,��(�)�R�*���/�����-ʊ�B�3/5�M�ѵi��6m
�O��dr�
D�2A챫��V3kQ�1V#J�\0�I���M�~���"Qަ鮫��(
�O�"ggf�sQ�0���'��OR���.�R7�p٧[�]�Tc��OR���Iҟdc4�۷�M#ʟбæ-�U��ŉP��	��'��	�x�	�|���>GQ���f�ʟsk ��ɶ<�X���J�k���T�οa\>��ቌe*t��.Z9{��3�GBß��h� �,�tӡ6�9�ro?Op)��'�B �<!BB�c�0���t���Q� Vӟ4�I��@�?�|*�'ئYX�뛬Fv��S�J�9��:���i>�
޴%�x��W��6�$�+�Z�An4t��	�?�ubء��'F�4o>@�x��d�ɂbT��P!.-0/!�d�<_:��0�&!7<U��c��!��R�~�L��e� ,$NT��B�d
!��3Z2"��Ѹs<��7ᜮ�!�$ֳ �4���F��Q<�8��Ғ=�!�ě̤���+X/�5�"�>�2�Ֆ�O?1CD���>�-qP���d�h�Ηd�<	���� դ\��a���d�<���6>����ߜI��8@&��c�<���5����̔0b�TI� +�[�<���I>=(\�[����H��V�<�@E����tcc#�'DK� ����Xy"bR2�p>���Ի9�P@ѭ#d���e�\�<!�%�*E/�T�TD�݈c�I`�<�-+�^0s���3/ҽ�\�<���sP�Rɇ�H�֭��oYY�<QWm\�A�( H[(������`x��p�l*�M��O,���cC)wDp�X��I#M��ʲ�'+���D���|���Lkȁo�?x2��`���赐�M7/�fE2�OL,�B�@Ó T��U-ֲMH��gDfӤD�>*�(�2��phnI�'C�Y�����"��'��7��OڈQ�C5)�T*cH��e�dJ�ƿ<	�����(�H�rh�|WD�b2cL�2�8����O��}��i[�I���Nڼ5�G��L�h�:Oq� �O ��u�A�E8����ٞ�Eh�M�9�� -a��v<��y4��� ���Ə۷ARlH��U�Й���N�~�\c1�5@+ ą���J�<u#@�pu�H�>��ȓRV:����Y�G�h��+�-5�	�ȓH�q 1��*е7cحf�=��4��O���C���?)���?q,O8@����'Z���tk;/,��@[4`Ű��@C�Oā��D�Os�˧�O�9IT-��-��ԏ�R$$v˞�p��p��K�u���Aՠ�n�1��eH�L��~����ٔ��ܭJ�Ő3��2L:��e�<I�.F����|�I�������e��	D�*.�īU�/}/|���I���'є	��C<M���WᄱYL<���?)c�i&66�4���	�<!�f��6���ii�٠���{<6����?1��?9��5�.�O���i>���:�(�O�\z�iېi�s=�C�ɞ'���SM�?�
��Ձk]��b�>��S��.��a�s�ƭQ���� Ȍ0���d�b����#����(�b]/5��X�e8D���'g^�8Q|�
� &�l�!+�d����&��{T�:�M��O����*aܞa06f&l�HX3��'��۟t��ӟ�R�d��T8R!� �?$�С�S�? N��M�'��k�&�|���6�'�l�XԮ�8�Xp��&�,�y��Y�8B���P+.�ͳ$`�0< J������Jo�Թ �ٯLBv���L7D��1��	�`�I�\��ߟ�&?9�<!H� aj��%��u�l�9c�m��,��^٘d*�@V��5 v��YC����By2��FDF7�O\��|"����?���U F�T���yǆ�۲.͹�?���W�Jܱ�����>�s��|S|��#Ŷ4�ʙ��/Ng~ң��O>1[���.V���p��!P��8�O=?	��֟h�I>E�C�7.���H�#)\e�����ym�Z��T	��P�^i�P�D%�O��%g���JT�N`6��1�X X�+�/�M;���?y�Y�n��I��?����?��yl�M�g�	t`��vOZ�1O�5�5�'������0M��8���L�	�R�8�y�EA��0=Q��� � h�	;FP�$��Hׇ��ET�<��e�g�c�F��SNK-r Ȅ���	�J���]��!��R���p�W�O,�ؽڭO�0Gz�O��'��M�� S�,�$�Q��n�,(j�/�*����r�'���'�R`s�m������ɿY������`\�axuN��1��܉5&T9 ��a!�!�d�(�$ރ/xb�
��[�PY���B�շ90�Yዶ *hm0�:0�a.ѻR�&����U�>]1�1�4U��O�d6/��=��OW�(ƢP@��CՌ��	A�	ϟ�&?e�<i�
�8�顡Gހ|8�p w'�gy��'�6��Oʓh�غA�i��'6�ah�^B��ơ!�����'�r��'l2�'�Bƃn���ʔ�>q�w��	��[�2�(��@%����zÓN��18T��9����`ہo����Q}�` ��۸���8P*W1�0<� ݟd�ɹ�M��x�b�R B͍S8ܱW	Q�x��u�)O~��=�i>��<Ʉ��'[X֨�H@3q$�Y H�Oy��'����?3�%�h�CT�R`�5y=�-�I^y>��7��O�?ͻi�+�A�/�b�)�*h�4���'c�ñU��'b��I��|eB���R�K�^�uh֤��a��q����s@������3�h�zp�$ϰ8mL����ҋ8�]ib���S��O��o����ON��2�J,�qH8�f|RG��y� �"��'���'����^��@rG�_�zb��5��j`�=A��@o��uy�>�Z�i�iXr����)�
+.�q��u�8�d�<	�-�:����?����ē%�Z9s@C�41�����>���~8�åzџ�Х[Ǹ�cu @�(�E0���dj��F��&�Mc`��?'��>c���R/�;4B���^ @w�)!4��Ob8n�ȟ��N�l�|�'��011��xU�@ �q�@ɇ�ўPE{B�'0�h�U)W$�X`���<�|0�@�'��g�>/O|��<�
W@��f
_vZ(�0�@�T���E+<b��'��'��	o�'B�Q�Pn	F\D��N�.B����Ϣ;ŤqI��N��`䜆7>LmБK���yK8'*�A��Д-�0p��'rLTZ G�y�P�.�l�v財�?!��~����'W�	ߟ��?!SFҏ���r��0�8C��H��?���d�O��&��8��efB��}����8�ʓ�? Z�8�'Z�� t�|�dn��a3F���XI0�]??Ғa��Oʓ�?A��?�k	8etL���ƭT�I��'f��C��-�ܰ�]�f4Z	Ó{�����d��h���#fG����o�P0�V�Z�6R�-�#���0<�����$�ڴ�?y��m`b!��4XV�2H�(>�rm����?I���?�����'��'��PӰi�t������>6�X�r�i>Q��"'T`�U$X)8���X6K�5����ByBL��06 ��f>el�ßd���+e�q�f���b0#��8�I� "`�2#�43����b�0�zfjo�%��LЗ3^qH].�q�'���82'mkZD�g
ȑ[��#}Z��<Ȳ�q��!�`�'`~�,�	�?��i�7��O�"|�7�ThhP�Q����u�qP�B\�۟���]����b�]���&O�-0�X1�,�hOt��Hᦩ�ߴ��R��D��e�,6��(}I� HC�'��=�G�4�Q��-Lx��u�(��t�D�rTC�	 9 $�Q+͹WX	SA��g�6C�ɟj��PЃ��ؐL��B�`3.C�I�<�h̳���'V���rm� �8C�ɪ/4p�A� �Tk�dh���
E8C䉿x�DJ�i�h��ұN�ʓ~�Zl��I�l6����F%XD$�:���%X�B�)� H�0Ո
���q����*6��"O諗��;P-N!�G�%.�ly��"OV܉���\}F�c.i��t"O(xZc��岬x�b�y��l�A�'A�K�'_�r���(A����QmB4_���'w���5��:m�J�P��!+��-��'��ջS�Z/b��Q��*��2�%��'3�͚4#�$��ū��C(��c�'@�`��m���Œ�! 9?,���'���� I���#ũ�*t�S��� K�Q?ap �>^�U)#��<S8��Մ*D��AR�T��:�gdS�@���;D��+㋘7R���qE�O&g���ئ�9D��#&�?e:�ۦK#1�0k��6D���"�] "ۊq���C/y�&U0T�5D�Ri��F���Kz:��X7M�O8T���)�qo�x��%GGLZ�R��#S�B�'�ⱉ��`���sa�a�tz�'�����@�Y�*hZQ��n�|	�'¼[���0eu���ڭI��A��'�.use�R�K�� ���>�-
�'d�r/�9 ~��F-1�
t�)O~"��'3�3���w����`Y]ux�'qfuh��J�k���ؠ�!@B|� �'��$CqH��O1rE1� ѮF��;�'��T�V�'"i���G�7@�$|��'n�Ħ��/&(�奜 O�\a�0P����p��qB�w����M��i�ȓ|v*1��� �fj�9��l>����:ā��s��8!3&�0�ȓJ��Z�k��^R,!�m�HU�ȓ\沥[���� ���Z�	Àޤ��ȓdR V	�w0�lKE*�,V�������~�a�ۯ\.�@SSJU `�:a[��q�<Q�Ꭴ	7hY�צ� ���oJm�<yV�\��@��"zz��Z�/�q�<i�N�719>�S�̐�1`j	 ��Oq�<��C��HO�!�W�,~-�A�bhp�<ဏ�=Ք�Pu�&�T���$���6�S�O���B�V�=�d�:t��\�8��"O���$O�x|ppv�̤d5�Y3"O"�K���qn���l��nLI�"O����@[�$���K
!��)��"O �h#��\z�h�
4��pY�"O|ܣ��U0;z0����B��@Y�:9�OR�� ��)�T�1'습%F�qg"Of�P����z�0�ǆ7<�*"OJpy�_����o���#�"Ork����>u��j1/��/!�ĕaoR��!ȁ�2�B|ӢΙ2|-�}R!F��~���(�,J�k"_�Z�ڡ����yㅼ��S�?�* ;�����y�Eu�D,���73��أS�@$�y��L{�K�Z43�^903�ӗ�y�J0_���U%Ր�ReO�y��:d�B<�R�������$�M��hO�]�r�S�#K�� C�l<z�0O�M� B�	ZyF��V�@,�juq��ѭ��ȓl�28��ڶh���-L�3Jl���L� -�p ������0����M�<�a+�
%(�
Sϖ�W��*���J�<�d��xc�YG��_��U����ڟ�q�)#�S�O�x<9�O��I~�ś5d�_��l��"O@)�݇Z7f�{�B�%'� 9`�"O� �C�ꀿ]��5��A�;�.�c"O��ZįL�=y��5���h�4�"OR����6yK���tH�H�^Y�"O��QW���m�*�3��))� �{TQ��P#!'�O�(�� ԿP3\�T��Q匬��'��a�e�)J��5	�	�i��D�'�x�2�Dٴ��8��#�+Q�z�b�'�,�* ��]�D���Q�R���'�p�8��;+Ҙ��&�7��[�H�T �4�"eP��=�0Y	N>{p���s#���W!h�����T�[C���ȓ.�(��w���+�|V��9�����_�����4yd��Jd̙Jj��ȓm��d�	�/���Xu�ŒN���R�،���3 6��2�G;L(@D{�n�ɨ�&@1#�P�R��U�p��8~%
F"O��7Jͧ%ELE񤠇.f��c�"O���V�\��p򀏇�`�����"O���4LKe��h3w��d�m
�"O���u��*5:c.�t�0B"O���S�Q��\�(kf�F�O�����)��؝x���2P+&I�x�	�'t\�b2*��qѕ�7G9H$8	�'�z}��mآ,��EQB���@����'�F�cG�/>�z�aV��3�0�I	�'F��)UI�-`��k�C4|�����'������i#<�	�����(OXp��'��T�ơ�.R�T�Q>ek�'� ��wIL��H�$[�/�t�	�'(��P�	/O�.8��M;I���'~<*E�^8 �^�r�1Xl����'���#�휾|r�aab@�8"���A�]d^Q�$��pt gI�T��ڒ��Ԇ�!�h臯�++c��K���!Z���Mo�m���*C����c�@!���sG"yZǯ�	W&&�0��N	I�0<�ȓ �Υ
��רa~��&&C�5����ȓb���4J;&����A>�rmD{BNG������ąO�5LX��#&��~��9 d"Ot����a`����]#k>��"O6�C2���;E���g�lD��qg"O$�ce���M�� d�̨�"O��t��E� ���I�d��˒"O����D�X�|��B�>e��Ta��'0��p����3��4�F�\�#Т<�.Y�� ��4�6��fDٱ](��N�_�����r�"�A�ʋ��CƖ).��ȓ.���rJ['��XBJTF�=�ȓ2PT G# �rZҬ��D	(Kd	��?+x�+�d��[g�]y�ؠ�L�')�`*�8:Zb5�/-*�p���Z���Q0pX�ЌL�"�"��q$D���4��z ���夂-��u
��EI�5�ȓ&89Rk�2R�.`�w��@�d}��(a�ᢒ"D�vNм����M�,؆��2]���2;�,hK�$eݨ����؋p�4C�/1�X��$F���b��#���C�	�K�*�{�0>P�S��d�"B��j� i\�DY� ��/�!z ���'������$
Ҷ�Wc�9w�^�b�'D ܃0�-�DTs���+u_@�ڍ��ȮQ?YA�ܮYs�d���.NKh$[��6D���&���|������.%2d�E� D�<3�e�w%p��0
-lz2Is�=D�� 2��ՈM�,\�]�"���{}�!A"O�రǍvY�� B�|z�b�"O���pn�:j$+Q̎!,o�!)�'����ӹE�v�Qe�T�]��"�K� ����ȓ�P�2�ʕ5z���b�?iU��ȓ):���q�Y 8s�A6�9oT<X�ȓO���b�PD��H�=8�L��ȓ@T�8���37hpI�'��Rʎ����b	
S��P�*E���V�p�'���P�y=�4�`��!
�����L��>܄ȓ�"y��B��B�stiP� ���ȓ ��|��*@'Y۪s�L�<9 �%�ȓ|Ph�	��ɀ.Ǫ=��d�G|A��lʮ;��5k�)�d ��GL08��I+8���I��,+%�~!ǀ��:Ҋ\246D�P��fI�+�,�G��$�v����4D���%O'`h|ڳ+�"��� �&D�LS�m8`���b���2X A��h0D��R��a�y%�\�g����"/D��C��#
|�0��- �A|��E.ړFn�D��̋k�D)�'RkP�1f\��y�#B�>���!&�D�h��T0��J	�yB$Z^�d���BI�yЏ��y҅�,U�0P���IL���ׇ���y�d�n�<u��A�
P&A1�&��yBf$r����ub4$:�Z����?�0dDD����ȑ��� �^�j���B��`8�_HB�ɼ:��z࢚�_&:�E8C�	�?�ty�	#`��YdB�	9-X����A�_c���֮�.6YB�	�xN�C�G*O�e 6oL�u�C�I(A�x\�ah�!<���S�-`� ���z�IÜ�̓@=N�H���O:"���OV�)M�jw*�#�/+K�-�D�ކ����K�l���O��dZ#]8��'�6;f�c�%����w�z��סL���	p����y�">y��d�z(�� Q�1��,j-��(:�K�c�i��ڋY��]"#�	�Dg2�d�O�c>��V�%.4�����_�����<�����(�!^�Gk�Y�H�3;����I���$�K��%��a�|%x�����Q6�Od`y��%�I�?�IC)���תH"�2�aTOX�FB�	�ڀ��',ԇ#�]Z5�T,x�2B�	1O5
H`di�9aN�]�פ��g��B��7T�h�oɪ{+�	��.�lC䉞@���K�ׅyh�U�©W�RC䉿_������E�~��"a�9  �����~���*(��A��7U"�!��fV�y2O��-������I�(y8����y2k����Q F�>�,�	u���y�f�.r�i�:�٠D���y�D��{�F}Ce��0W)�'!�y�ʔ,J��)"4��'3l�dVg��?Y��D]��x�3	�BX����H�C��Y�1D�h3D��?p��L{�oT_�T�Ƭ-D��2�R�0�f��g"�"doV�ɷ�*D���d+�QF����;V�Qa2�-D�X����`3J�Ʌ�3n���F(|O����>��%>.�\�PpFDW�H|�aA�D�<9�^�OR��r A�*#Z���|�<!$M�0[֒(�cJϋg\yђ�z�<`��64�JMQ�O�weنMv�<y��P�0���P���ޕ�ITk�<	 L2Q*��`�ݤJ�(�iBLj��I�vTDxJ?����	�f���J7P�k��32D��b��ܐa��N�Z��A��*D���&C�B���KVɠ3i�����4D�� �	R��1*r�U��C��<f���"O�e��S�9(�R�,V�N� k'"OL�F�Gd����KT�!�b4ZC)[��O֢}�&��y�n��O�B�����'4΀���6$t���8	��5��#�4�|ćȓ^��,�A��'!b=ئY�E��,�ȓl%
s��i��Ka��:V�H��gp�Eys �(n���3s	z���vf���΍�s�NL�TM��P�.��$"��D��R�Y��e���:�d�,t!��P�R�0@O�y��-P��28�!�$�>�.�Z��3(�dL�A`ΆT!�_M�L�〷B<4)��{����'�
e	���c	�Y�#+� A��B��d�f$�!l�_�	�a���ȓႧe2���o�=!#��'�R�'��
!H>��So�Q��H*?O�遟++̜�Dc4T��9����?��pQ`�	�c��l��,Ѣ^��'a����1���4�v�s�0q��1b���` r�'��'��iV�@��cb�5!ќ���"�'/2�'�b[>�Dx�*R�1���F�5g�@�صK����>!BT�$H 4�����i'�XIu��<q�YE���'?�O�Ҕ�`p��K�3���ӷ}�+��O�ax��ɜ��CP�ĵ$�>�@^O�HX��Ҳi��':�u$>Ms��*���1�٣Y%�<9Ъ\-�M��?F�9q�'X�S��?)���?q�'�:�b�A�J@��m�>����`U�*��&�'E�����'��P�r����u�o5�1fuF�I�k�fDjf�@;ž�AV'�O��F�d�
��ݺ���?Y�'�?�'K�uIS���u��#B[V�[q�Ws\,���O8
$�Ox�ɑ-
n�s��N���N�u���"� ��g��
7!�?y��Hߟt���pJ����OJ�I�O`��vʈ��D1X��R�dv<��oHП4���OR����}���h�$�e�?7��-��/�2a�'�J�d"��H	�:��l�<�q����D��>Ur�'�?a���҄� 0���8pv�Äo��t�|y�'a������?�׼�@��x�P��/�?Yoڈ ����k+8,�X�V�ƨQ���ը����Γnnt�I��;u�2���?Y7
Q�_c��!�柈�"��Ȃ�i��DqT:O�@ �'�r�O��1O ��;��`rR��B��@�Z�x���qӜ�xb#�O���?��S�g}R��v����&��/W�P�+A��y2�WV0cȟ�xp���@f� �M����?q/O,���O��$�O���{��Q#70�Qr�ƹ<@�8P�ݦ��ğT�Iӟ��	����ȟ��؟Lj�9���rk�7ot�	2�j	��M#,O��D�<�L~b/O0�iSOC�)N�p*$�U���S�,�ߦ}D{���i�6�r��^(�u�E�0f�����O�����g��C7M�I�$�P��<?!��O,^�TY�8�衐�KM�,&!�$R)RA��Q�� /Rxb,�3�\�!�DEp��8kpNZ���^�!�$N&_�"�%�>6�E��3�!�d�:#gތ�b��5�(�b�ۂ<�!�dT�xl���ۿH$Iqt�ҼJ�!�����%k��UeJ9j�!��P�tp�$��^؎�e��z�!�R�0�^�C��N�r��CB^'�OJ��B�$Ci���&	�o���h5&96|8��G*lf�1�:o����.Kd&�w���X1K�Ǎ�!�� ��<@{����	�xyq)w�����<Q�����a;��
@,R$:"�x�QDZ�d�8�����-5���� e�$1N���L3RSP%'����{�[f��huT5{#��hm!�䒸y����T�Vf:6�k�@\�Rf!�DZ�Cl k���3���.F- s!��+�f) ���?�p-d�!�<GJوd�
hhZ&IQ=q�!�$�Xd��
�(�e����gv!��b��jr-�w�n�W�	!�DC�n��pS�f�B��)�,�B�!��K?" >qHp̉�Ԛ�ѩ6%�!���p]D�h�E֙5���
�S5Aq!���+c���Q��Ǿ�`p*s�V�	U!��uZ�� ��.�P�r�#[!�č�z&�ųC"A�p������mQ!�� <4�e�]�(��C�� BAh�{A"Oz���2@D���7�f��"OP�B���#��%h���xi�- 7"O�ygݪ>݌$�MN����x�"O�ݚ�k8J|V�i���S=�4�"Ot�rD�Z��Ĩ�1b���2P"O�ec#�I��H�,{���E"OZWA�O$���ֆ�7UH����]�<�B�'5Y�A�g�7~���TG�p�<�w�ؑ7v2 �FU�f��heHj�<�䎎UB\�ᦉ�}C� �G_}�<�0 �)��,;ufX�`�!��$�a�<���q��: ԮU"�M�VC�D-(�pv�96�R���� ��B䉮��	�#ԳJN0��]�&�B���a��)�$݈j���g�.B�	(R��8���Q�̊1I�cg�C�ɜ<����`C�ǎ$����L��C��L���Dn�1��(BTF��C�I�R�����-�Iy~��dfѰ)y�C䉞f�(Z�"p�$��&�*7O�C�ɝg=��3%�K0o+$� ���G�vC�I�<xi��)i#����� �6C䉙��U�Í��Y��c���!�C�ɻkE|�S�?|�+0��-�C��#���S���4$JX)c��D0p��C�I�j֘@zL؀j���8B䉍v�z�΋B��dG޹MB�C䉠/�TyK�@ڀÊ�`��>kpB�I�ze+��)�|)`T�V�n�bB䉰~���[��L�@�N](Qc��V <B�;&�1��	��̈�mN(8B�X�l�1�M�qJdH!&4�!�L!=��p5�Ğ T�ٓ�QN�B�I1�����*����1'�)x��B�ɬRm���(�S�ԣU�R):��B�I�dЪ0��OŦL��C���1-�B�ɬ]�Ĝ��e]�b���hԂ͎eW�B�ɸ�d��G�6l�a�ǌ0s�C�I� H���&��9��=�V��T�<C䉡S�ޅ�e�_�2i����_�3�C䉋
HI�e/��.�tI�u�ސ3-�B䉉F��҇��.K��r�+�zB�I��uy��/m��-�sI;M*B�ɌPx��B�ٛ@4�q�d��#lB�	�3IJ��W��w،	a�*"�C�	QdӖ�F�^`�ͶC䉒R��}�rCέ!�Xu�N^p#�C�	�I�(r� � wF�x�n�q�~C�	�4ܚ	sG���PJ�1���$NC�	�;���b���/Ba�)�~�pC�I�/�|̋��S7�Ҕ"AE� W,B�I�#�q�+-ۜ�*���%4B�	�WjN�d�i�0�BŬ@6PB�ɽV%|A�q�C�G�3�,�6R��B�(%�j��pI���HBc[�qhB�	�DdT��g�@�o�ѠamU�?uC�a�Z)��%m��H�6!���B䉈^�fJ�/ֆZ�3K<r��B�ɊY!���sJY9C��RPBB�I:4��U�+Yd�
��E�HB�	�v�C���L,��b�B�4\C���Dk�3�(�G_���B�	eB����^��� h�e�zC�)� �I`&j�>O��@���0-��5�"Ol�P����d�ֆԹ,���"O��#�j��V�4x��>Z�vL��"O,�R�ע(en�贋����!V"O����*'�2UjE�:sr�B�"O9����Nxٻ�L&*p~���"O$���V�f�x#4��_��mQ%"O����x"�iܕΨa"O��i�dG�0�<�e)4)�-"�"O2����)pj�s��"[���"O(U#�*��[�0�ĻR�x�5"O
�A��P�l�A�$o�h���
g"O#'�)K7H�ʲ�Ţtin�p"OJ�t�L9�8D��53x�"O>�҅jZ�t5@XH3BL�'P���"O�%K&-�<r����_�
�l�x�"OVh#��ðN '��n��y�"O��;e �md�X��h���8G"O�ف�%�R�*�A���0O�8���"O�����2?���Tc'$�RRp"O` 6�],P�p s��L��q��"O�4�q�/(:� �!y�T+F"O��ѫ�7�ً�H�Q���f"O�1�/Ĩvq]�o4n�8�j�"O���T62���bS�'��]S"O��S'J%ʸ�H���C��Ń�"O��;C��1}8�����R��d�Pe"O x"lR�{��q'�E�QI���'"O�r��ǌ�ls��Y;�p!�"OZe� Q*g+�DJDH���4�8�'���'h�4c[x�0��Q<�)�'�Z��`��7H�P]hԠ��Ĩ�y�$O�~]��)@`�J΂L 3eC.�y2��=(Ĵ��W�XVG��f��y��Kx��͆?M���̈��yO@0As\��t�	)DL4Qc2���y��QU9s�JK�����6�y�>Kl�
��Jp2!�0O�'�yA3v�$���\ DB&	 ��y�e$X�ò�S�J�1�%��y�'�Xz���V"�,t��J�-���y����-'�a�B�M�ps6G��y�N?�b0a��zrZ5��N��y�#�=7p�,� �X�IB�|��Ͷ�yR+��8�����V	H�1����1�yB���!cJt�F�#J!l@��ٴ�yb�_|-<��$�E/�������'�y2��x5b�����BČ)RC�ɤ1��w#X@��� -`�ZB�	Z�P%#Sb�(*�%P�@C��B��? �D��ڟԶ�öH�0�B�	�F�X*�m�8
��1��+YLC�I-2B�붨�X���Ct���LB�ɞw�R��1��{Z�#�D@�8B�	B��@"�÷@����&@z��ć�|����]�R��e�*5�!�I/&�i�D�Un~	*�����!�$^؄i04�Z8b����.Ģ�!��H�a��
�J5TZԲqO�&0�!�� E���c�';C�a����V�!�D�!��� �.@zY��B�!����8d@@�Č���G�K�!�E�^t,0�8d�n3SFP��Pybk��XnBq��eɈ|��jB����y
� ������K�Vd P�C &�Ő�"O�8#��E4w�L�3/��6=Х"OqpF��+#����J�0"O��Z(��|�t �T��}�VT 6"O������Y	�y:W����qi2"O<P����YdٖC��mq���v"O6�Ivϓ4/�
���kʉ?�6*#D��I�F�;1>�!i�8YjT��t<D��b����S����'�u�c�/D�zթ�:t[6��nE�N�8%��.D����@ DyJ���v	�DL9D���L�|>T|��+�:�<f":D���JCx�p#���0���1@	:D���"�Q�l�������\I���E:D��rc&R�x�@d��i�*D����;D������8P�\q����U���zC�	�g�T��w��g�\�*&+D50׀B�I'J/����Ą�?�v��#]9O�HB�	>9,�9¬['3PŪ�i�	T�C䉼Tў1��h]�L�D��̙�j��C��`���E'Y�##��8�L����C��R?~�*����:�0u�㩈�=pC䉬{Y�|H�I��%�s�9qB�	�)9n=�kؽ��B�E܎;�TB䉿~�<	��i�' ��2��h�^C�	�+�vuc�kS&VMĄ�gn��&^C�I�V���B!tF	J�ə�<�6C��,(�l�G��U�p`��J�+LC�I�	�0dA��#%֤��A�<C�C��e���2.H�z��!�(�~C�	p���۔�[}� ����jC�	�cX����S�T����F�:�ZC�I�_Ll���ψP�Y�	��BC�	>}��53ϊs �d8p�"l=,C�I8��੓�yUL!iA�,5�C�?�`p"f�f�5SA���C�,a�,����~��uxdʟ�C�	��1�NK� ��F���C�I!Je�����(C����ͪrAnC�I4k���M;�x��G��*r(B�	#a�H�2ǇX�ܙ��H,B�	TD���#dB�dQ� ��a B�	�6��9�e��3��i�Xhy���?D�8�T�O�{Pt)��G�� �/2D���gQ2A�9H�O�<'�(���.D�4�Ǣ�r^`9�#ӥ6���ӱo,D�T� �9�j�#��T+R�5��b/D�h�肄wmBE�rO$X�tyq��'D��I'�3Vfr���7
�V�1��0D��; #ӌ|0�1��4	��0��/D�����kb6�g��<a℠��"D��꣤2�*���I_��=���?D�l[�dU�l!`"�
e��� v�=D��җ�C�.�M�G��4�&�A�E:D�X �'�#*}�zO�u� �zu�6D�TKf�l��lCR�(p1���c6D�����-g_F� ������qVl4��J6~8*4N�,��9�0n�e(D�Oʑ�dҽ	�Xh����o%~�9�"O����)ؓ^��8��@�'0X�(a"O�a��)&Z̕xӈƕMGd9	�"OKǘN�*}����&yQ�I*%�P��yr S�FQ�7���{ނ	��O	�y����%��\`�G��%��2�T��yBP#0���K�ɇ�q���ŨG*�y
� ��:��U��!�U,�Z�q�"O*x0���)&"-���3�F<��"OT�HSg�z�,����:��\��"O� ��1���0K�0�K�"O�ԩ&.ܼO�X�ʳ���.�5� "O��##bŞ����ᩝw�x��"O��x$d��|�J��$�Y�qR0��"O�ABPG�)ijQ�]Wp|��"O"Ѥ�l��}0�GNk�<۔"O4�)��O�:"�h�/R�#�Y�4"O�P�����h(8�֮���H)u"O���_}�h�RNCh�@30"O����Z9p<(QM�>P:*Cs"O`��\���z��X
�� "Orl�ēJ��	��Ѧ
4l��"O8X���9S(����+�D���"O��1!�k�������l����"O.͓�M�Ѝ�q�ܜ}c���W"Oj	���	�rd6L�郩V1Rً�"O��$@MC&iv��&y�y e"O��bv�3N$�)��%q=<���"O�����d���!p"Q��<���"O����ǔ1t��u��m�LE` "O�Ys�e_46b��U�Z+r��U`�"O��B6
I>�؀*b�%/��9�"Ov9PA�|�;�JUWV�H�"O���g#J��Z��&��R"O �q�N8����֏�/��"O�([�Gҳu�\��6��t�����"O��8W��8�<{W"Ī���X�"O��D��4p���W@S�R��"O����� �E�F��צ�P䀡Z3"OX���U������9�\�T"On8kk	�t���z��`�6I�"Oz���G��]�B�DP���S"O�xT�� $Z����$|A�"O\ⷩ�6
n��R �Xt�t�2"O�,
��P�~ m�
 ��Hc"OJ�	����Ia慫g�ޤ�t"O�p�b�����P�Ф��L�8a"O��8qj�C�쵛䙏VQ$M��"O��Ǣ]�+`�RT��T�"Ohm��@�j1���X5`���jT"O 1[�
�5ftPD�Ս.�޸s"O��0�6 5�  5ȋ82*`��'"O��c�
Dm+&�1l��R�"O�M����4��$L�,�N��"OY� '�Hh��d�)�R5!"O��q�\�B�v�V�%jQ�R"OR�8���D2���өK�{fhQP�"O����Rڤ�i�.VY��t"O&�
�m�	?u�D"� ��9�"O��֥��ǬA���Z�M,|��"O�t'ϴGڢ J���zo(��D"Ox�:���-^����ڳHg���"OpՐ5D�b�T�O'xIؑ��"O��BY�cz��u��5U�x���"OБH2FU*@�v�J�N�)|�5"O𬰡�6T �fK	6�B��@"O��ڥ%�g��(��G�N�)��"O�({7�CX"��; F	~yQ�"O��q�A:T�^���YL��"OP�bW�םGZ"!Apb	��$-�"O��4IEd��tb$Dܣ��l�u"O� 0���	Pr���t����"O�T���Ԭ]H����j�X�� ju"O�P��^/�|R'�T�g��5�u"Óa�-��K?nu�@'�3z��r"O��z��ܠ��9��e��!�G"O�����P�v�{���:Ԋ"O��+�o@�^�`ݒS�ߴ�B�t"O�Ux@�(Fu�ԡ�z�q "ON=Z�èLђ�� C��iXX�(1"O�d�楘O�P�7s�6(��'ԺxjbM�D�v]A�鏮S�$���'�\9�L],-�� O*I�\�b�'��d�9��A���.|�\qK�'0�Jǋ�q	D���ų<#����'f��`Den\pD�<Y�%��'�5�De�;�Ptd-H2�� ��'x��j� ��a�v<����)��x��'����i��ZoS�+��I�'�F<B"�]Z�dBOU�*���b�'�Le�a�ݑ	��-��Bӏ_�؅�'.��b�
�4�蕃s�T�E
伂�'����'[W�*`��>�l��'�tQ�q�G�d���C*S[�v�h�'vB	�����7*�˂�\�Z�b���'���I��P6OT|X���)w��s
�'����R�p1�5S2Fш+�ܙ��'M�8��nĽ&��s��
]�B��	�'����e_(6�ɓ��(T����i�&�(��*x�v����ۣ[!N�ȓ�n�I��ȪC�rA�t�����h�ȓ �~�)�KB('��I��;6����{bP�$nԶ`h�H�d����&�X����0=� I1Y�*}�c��0>Ǌ��AMTk��آ"�E'z���"+�-\D��W\{���(�xBKN�p.,�I���<h-rU��HO0��!/QW̥IA�D~�''/�\��A�	|@�ƌe� }�ȓ!� �1�L˃o�ZV��=���l�x&�h{�� K
9��O?7-��6Z��e�s
fiSe鄉E!��G�~�h�n�	�RmCg&�?^�|m�8}��0�H@�-h�e��h>#>q�BY()A�M��HJ�ʵ�Eu�P�P�hr��r�$�3���ڠ*���� dD� ��(3�L�Ͱ?��O�_H�����;F�]H�nW`��KI��pÏ<?�i���x��������*#x���3�#\��#"O��R�W�6�aQ"���6DFp��˙u�~�d�	6eҪhhGl�j<�>�I�;Zj$�el	���T�&%P�B�I9e{:��� �z�\��T܆a�*�Qڴva#VG��>ʁ�4�Nź���	d��pge�T&�Cw 0�����ڄ=h��>pHF��J�2?g��aW��, ��:�K-t(�w~����և�UlX���`֚!S*�p%�)�ɴJ�\Hb�J?V�V�cE#��7�?#�O�Dr��oS�
�����6D��`s�?8%�f�������.vw@���)A�*�&�Z�c�1�MG���w��1��F2N�����Q�b�Q`j4D����_����i� 	�4!��`�M��c�!_>� ��$r�l��Lb�o1*Eeڇg��9' _�=��{rNJ�3��D�'`J0+����E��55�Ĭ�$N�!gj`[��Y��YQ�'�d��V+�5B(pi�a@[�U����?I�Z�L�
s�F+P��4ːV�	]��N�{�m�0�֥3����^!�I7@�pD��f�
 \��4凒}��I�w�Q�"̈́i��7�s��k���B�\��w�U���"�+D���*ڎp�ƙӆ��/1����e���D?������3�IuB9����� ��6��4m�>��D���l
�� "��%����{6H��^��  �'��d1��(Z�l�uD�>C����½,�f��M[�81�����n�;&'Pmrb�d[X|�"O� T��E��>(o��0�cX �lQ�q�O�@{7E��^C"�O�>c�!�
$��)*COŁ'K�H�fl'D�̢��=f~"4���z��E�l"�$>u.���	,�L
˿kc$����4�B�I�H;X�q��&A|S��V$��B䉝�4p�-:C���AgGY�C���� QĜ�W�ڐkF�Fi��C�I?uʈ�ᕏ� ��xQmɰby�C�	B����b��l"P�;\�C�	 '��p6�F3�F�(6�9s�DB�Ɍ=):a2`�V��r�3N#�B�	��LX�E�)"&kS�B�Il�
�����
 W����&N^C�	�(ҍ�Tm�N��Ab�CC-��C�I�(���yw/��,C�	�$l�(%��C�I##l+wa�� ��e�'N��hB��+ʅ�e .��-Y!S��q�%D�̺p���̃dC'p�����!D��b�̷,:�ꞆD�pqj3%"D�`k�A�'gf��)�#^+Hq�pX� D�,����2��Zv�ߌN��)�'�/D��h��V���%^� Ji�!0D��"D.T�wU������-?D��@��{Р؆�M�bU��ʅF"D�܁s���p��g�=T)"�;D��۷&�P-�&��r$� �-D�Xj F�{c8�����p�%�%)D�(�,�F�ȥ�Q���V��-[�6D�(Aр��[���9p��/)D��a�@(|
��t
�	�4�1��!D���vO������(L��C�1D��s$
0�i)d�͵a�2���1D���Vl�|{�A*'�kd�	ӧ0D�t�cdʽ7�8E0dǊd����i$D� �Qg��_Y��c�`�qSf%�1 -D�p9/J3lր��)AkM>uB�a)D��t�" ��]�7�EZ��$$D�Bܸ97��c!L��T��B- D�(($�βs���qC�W�Q���`.D�H�wo�8?���5)�{G$<�1c.D�F�ӲHeܬ���
-�  ���&D�`��F��'�J�1 �Z�X�`'D����K�����эǀl�� �`�:D�0 T+�B5J����*���Y�'D��)u�]/U���7��nq#i%D�XP"l�65%t��5lʋA} ��
7D���E	S5qt�{�Ȗ�-��%�?D�0�ᆏ��
�K!���o�@զ=D�|���
b�|��ע\�  �B/7D�,�R� ��a��}�LG5D�D�Db�w$ (�C��04;p�B�/D�$�0��0����7?�J���#D�H!ei�7f�NP�bA�t�0�*Ţ;D�����	��\���X�/.�	�D)&D��+�*atL�Ŋ�%A��գ��!D��qw��%v���,D~�P� 4�4D��k`�ЫOo�cP��>�N��Q1D��	��R�N���!�H�m��S��>D����+u� sy��m��:D�\q��Q�.�z��K'��УA9D���V�P* ``t�S�Fql��׊&�I�v��jG'��8�"�S�ߪ�O��P��*T�2�P@�Ŵ�Ͳ�1D�t@�瘶?�p [��T1 ����$D�,8#�	�@RR�HBV?	Gi�R"D�� �XfM	#,�0��Y-O�<=��"O�3�-I��UJ�'���R�"O��墉�2%��I�� �?%@�f"O��ч�U$?]�Y��%���B�c"O�X(�o�5yض�1��;
��Y�P"O�����.N�z�0�A/x�D�"O�0�"P#M�y�! &_x�ه"O�+V�ԟh�Ȉ�CgN�\Vp�"O�Ha&� W�0!K6��0O��"�"O� �ϕ ��a�	�0�"O����̷(f�����\7���'c�!�կ!w��C+Ia����'��sV��0B`����f�Qq���'P�L�V&W9�.�Y��]�NZ �	�'��Y���S�-N>��L=u��U:	�'~�5:�%U�i�P�EG��#�.�	�'���KflW�*��s��̩`�R	�'n5��G��Ζ��28Q
�'U�А�eI�M�H�$k���V@�
�'Nhm�t��%L�Y�	Õg޴�	�'V���D&O=n>Az&�$U��	�'�F|��ϐ�P>(���J��H�ze1�'= �*վmbxS��_#EX�=�
�'����D��M/��8�(��K��+
�'j��b�$��r��8���*H
���'9:��DA�:h�ČE�X"�̆��� �w\�26�qx��F@���"���S� E�p�r�a<m0�ȓ0m�Չf��:L����͵�����m���C���F�Į`��y��.�x� ��hAz�@��'|�0��+����5�@A<ш��Jt��̅ȓ}S� c�[�HR�y w#������ȓMk	�N�*B�ݫ�U;�,	��I���B�K�.[tt�陎�D$��fZ�̠cJ[�Z��!KF�Z��ȓ�hdS(�&VU��2��<��W'z�0� W�z�B�_1|*��.��ۓ):�
�BQ�Q8A��D��+40`��#.~�ʂ K�X$C��Z��4�IV F$a��U2��C�	g(�U(�] uئ�����&itC�I�E�aH���'>o>t+�)�0�B�	�}���#���*m- `�`�4P��B�ɘjT���"kȁP��@�߂.�xB䉫f̊�RDL	F8�=R��B�W�FB�	/@*�e�?i%ܩJS��]]B�	%4z��+D���d�₨�~@B�	�09V՘a�N�X6Zu�U,�7|p�B�	�u�.��5��)uX��W
�w��B�	�jM*�1�n��>�]y�X�-��C�	��b<B$��;��uJr� ��C�ɕq���˒N=|���0�שM��C�)m����9nĎ��Q ԦR �B䉪j��-`�	�ĘaQ�m�-��B�I�?6�l�#��%\��rPI�U�B�ɧw�z�{��ut�r�%$0�B�	6^V�Qv�)[@!�� ��B�	(@Ǥ��jYO�@z@T&q|B�ɷ�n�CujT+C]�`��R5lRB�ɾ5ЬTF�W�M�(��2A�ZB�I|��|��k�? �؝��L�E�"B�zp�a�F�%.�Q3/͚/
B�	�+��(O�a.�5����B�)� "q��וi��A��a�W�U	�"O��ZQ䍨g2���æTY��H�'"OF����MI��	0 ��>D�q"O����]>rX\YI aÀw>8L�"O̼bfÂ�:�0c�G4G-j%"O\�;�JL�]�n�I��x��T�D"OF|�e���8�TCM�6;�6"O<=��Pql,��ЯR/3Ʃ8B"Ot�P2/^�[��"�݉;�j��"O�X��.�$=J��#[�
j���"O�ݫ�
��(W\����>G��4"O�H ��I�2-�M0,U�����"O�9(�l o��1f+Ea}P@��"Or����M{v�
J�\UҩC@"O"��w@�$s$�a�	�%<��"O�U��qh�ǩ	2.8R��"OƩ�Մ�7��q�s�Db��"O��Xe �?���#�'��WPF@J3"O�Ap��'��+�gT?F�F"O��ՌT�،A9 >|J3"O<9����?
�@�%B�m�t�A�"OV!2"@��G�jm[2K���(�2"O�L[e@�NY�U���̘$����"O	�,��r8!A�+��?��]HP"O�]X,�*<�a�K�
H��e"O����-|c�P"�Í7h�d��t"O��
��o�X���h�
O(z}z#"OR��3��#hJ�"Q'�	Ҷ"O2=��6
��4�F�.;�,���"O4]�n/��:P�ؓf\��w!	Y�<QDB�1?�d�C�>��}�E�HV�<a5�؋��� )� �H��P�<1��C;n�6��Q!A?u����sIe�<��i��@<Q�(��e=�T�
x�<�W`�/�hH�-�G��[J�J�<Y@�[�<��E�&�� EH�<����tk���R�Z bZt`���G�<i�O+Vu��`���9��"v��z�<�N52 �K�a�I, ��n\y�<�2 36]$LoS��`��$�_�<i#�ش3� �A����>�0��F�<����"\���3�e�0js>��� ZF�<�`
�!��AA �D�a�!:�_@�<1vHT����h�x�0��{�<����*��Ϗ� � S�n�f�!�dP�`c�L��#�=Uz��E�!�Ȉe�ޭHR�I�q�]b��΂k�!򤟄v(�����=<�E�Əv!�Ğ����z��ξU�Ph��ƸRq!�H%HH;e�׾b~�K����z�!�D1.�8��w!��-�� �/�!�D��[5�y�Ǘ�f�ԅX�FL8z7!�Dʔ>�h�tf��6� @	��-99ax��I=[������Ð%1�J�C䉼@�(���Дdy���c���C��.<2����G�b����]�B��9}�<�&�M$7�U��H��B�	Dadah"OϚ3��RT�Ƙ)׌C�I�T�	��-�kGv���YB�4��ГO��r���U��$C�����a2�ǖ<K����/�$��B�	:��{7�H�CA�,����w�C�I�o�� aa�Z�� a��6��C��>$�N-pB$$X`�M�3Z�B�)� z-2� T4"�
���%i��"O( �lՒ\0u
�aC�k���3�"O�`�D�J;(��i27 ӵnԠV"O�
!��Fpp�I�E3����"O��A�ۭ��!�cF|\��"O�E�g)�/g���s-ٓ{QȔ� "O+e��)U���&B(m�j�
�"O���b�G�@з�Q�5x`LC�"O�UV)сIB��E䖊x[�E"O����'ɟzA�񠷨[�DvRm#�"O��� ˁ�,�,QA�Y5J�4)�"O�h�q���m
ƕS� �0@b�"O��`�ό4.�����i�"O(E��K5/M����b!��A!"O�U�Ӏ�������N
�^!�"O���@*�.�B����3�,�Q "OļxC���Xut���Y�Nn�HW"O䐠T��P��1�%�!a[����"O���#�9d�>���$5X�u�"OP4�Ń@9����"<E���E"Obe�b��y��9Ц�VD`x�"OD��U�|C"4���9-1 D�"Ov��',�!i�I���	R"Rr�"O�y��H�kw�%r�A�6 ��@"O�� �ΆNG�x%ɘK`��"Ot�����$t�Y�W��%g�r-T"OZe���3�ȁ�!��0T,��q"O^��f�^�E�rqDC-/�|�1"O8��`� �m0���a��<���#"O�����u�Fq�t��J�����"O�m��}���$��8' Y�#k.D���I�<4��h�g׌L+
Yb"�-D��Q&�Y�)d�
�Ls3B���*D�����T�
X�~�H�rq;D��C��qr�֭�� �"�Т+.D��;���bF��Ʃ/A@�ȃ�?D�����%)׾9i�
������6!?D�lCĚ�Y��|Je*��
���<D���l�@nܩ��H�Fђ�I��&D����ĕ3s�9��$�o%P�3��#D�� ��Tުݠѧ]�<�	2$ D��[0L�6p$;���<6� �	B;D�i��3���b��`��)�l7D�l�!/k�v1z��H�45D�RU�6�$q�@��Zg�t�.D� ���Z&.��XRr�Q�6��,;�E&D�zZ�`�� 2 ~zA�ĮW�%!�&�P�tcϞ}j,h``� X�!�d�>z�%��̠.`�rb�Q�!��Ke���� I�s�ozs!�D�J��(���f�m���\
!�J~��v�
�no���#��Pybn/@p@�C�<��)�Ҥ�y�+�26>\{'ٳ,�a�UFM��yr�97]~q�D�u��dH%H�"�yb
�9Tt��X��B�9u5���y�N��hݣ�?-U�<KSc�yb�OR8E���*Z�x�"b��yB'O�%ݔ��b,Δnav��ǣ��yb*_.~%qh��H��7넿�y��R*$��˛es2�@�J=�y�˃�r.����DаR\������y���H9gL�4����r�H*�y�����/���Jw� �y
� 6L�d��jonH�L�![�,���"O��C��E�d�
�:$A�x�b�"Od!�!Z��E��ѥ7�l�#"O�q;���?Z�$4�d�0�
Q"O,|�t��,�][FcF3q��m�f"Od�أ�K8Y�����4Q����"O�(��'�H�b��g�e!��R�"Of9�6nT7�`Hd�_� :2�"O0�H Ō*Z-�QPg
�1w[(�"OLpB�ޤ{���F F�[K<��F"OęP@��O�б��o�3�n���"O����AR5*s��1`��:Z�}93"O�=Vk��S�
8��Z�����"Oj�賊�����Sݨ�"O�h���B�KLb�bD#LM4���"ONe�$GB0.�\BŢ�U�3�"O�0zU�����S@�^���a�"OB���b�].(-����F1\�J�"O�مg�Z�:��'-��=\��"O XQ�Ḑm���8A���W�P�*t"O�M�,]36u��q��Wp�����*O��z4���o�FA �L9{�i�'�ْǠ�^� :�ŗ�-�H
�'�:��o	�7����ƹ+� 3�'��j7$���`Z狊�q��=��'��(��'�3"q&L�nM7q�@�' �8 Q��"���&�b�@��'(��Aā&���E��'�����'A�y��-=��Q�X�J<��'��l0��ރ�������O
BL�'
d���۪G<�D�Þ�s���R�'9e��B1I4A���p�� �'�B<@�& ��90�aĀ���`�'V,(�jU�,��`S���|��'>m04�˗#����� ���'f�Hyu�9{N�2ŧy�< ��'_�9�n��(���խѢ]����'�\�x6�@�^���)J��ы�'��=��б.�S�#ܩ1c~���'t���GO�2b.lc �4*����	�'�"��,ev���薍Sx��:�'�>�$gu����GᎿ ��J
�'\yz��4�D�k�N�C)x�r	�'��$2P�	=������f`���'�aHg�
U�����o$�j�'/@��gJ8��(��
�"�V��'Yt�8ԡ4_"� �R7��4	
�'xL�#GH�;,���g��$u�X�
�'h��`�@1-zFe��!� _�<T�RS��]�Į�<�d��J�<a�'V4m�+�i;R,���G�<�7�7t�Ve!K�:��(��'D�<���/{@��	�%bpp�ӣ�|�<������6I�;>��P��
|�<Y�L�*Q��9Yq���^����h_�<Aw�w�V���߻T�.١� b�<)��
�,�5�ϴ�=��]�<�uG�d<\"eM2;x
D�WY�<	��I�?�u�t�1�x5(�R�<��)P':e�Ó��&�#�Y�<�0�rM��K ����!cs!l�<�W�.]�c��?
fl�4`�k�<��$�	uo�ͻ�I�]��i(2��j�<�s�l���r�e��Q�r	Г�Pj�<� ���1�%��8B�ΐQ�FXX�"O�Y򐇟�Lm���! 8AhF@��"OF�3�FҔt!�x�h܍ ���"O�qԪ	(�~9�!�K�D�6"O�HQrJ2O�p賂�D� s�ɰ�"O��S��7������$S�HS`"OP��N�1r�t���cVINDy�"O*ݱU�Q�?�h<x�ERAe[�"O�I�c
<$}DyyD%�&���3"O��BFӀQW��;S���0d�V"OJ��䏜5i�FHcGȀ�Ym���"O�P���9E�\��
\!Y0J��1"O�H`�c�9=\�I �H�=���:�"OʔpG�̘
���8�!��P�fD�"O�k���?[�l�da|��'"O�!j7O��&�P@Q0�e��ӆ"OB��V�Bhq@86�u��qZd"O���sł2�����,�
d�fa��"O�񺃆�W|�Ȃ!㚽p�"O��	�c��I5��_;h�>%p�"O�eb��E�6N��S�F��Ȕ�b"Ojx�@T���-�գ̤*ގ1ç"O���qHQ6	���OL3vpH�"Oh�����'ݲQNA |B.��W"O^��5�
7n� ����
!E %�"O�!�͑�:����r.K�d⦈""OF@1���)wF^��"�5|��=#u"O�	� N7Ť �(������"O�e@�(̼i�G[�N �"O,�D�M&�&y�����d��9�C"O�̙�'�'��Q�4*Z`��"O�
�g��k^�S� �	�ၱ"O���f�|��(`�̨/@:��0"O��F"O�=3�h)'�=k�"O����CVDԘC����8�`�aA"O"M�6�I�V��p��c��%�Ϭ�yb-ݚ/���Vi�5�2��Q.��ybKO<�ԡC�ɣ88>�Rm���y��
	[Ѝh6�J*3MlT3�dT��y늗 S��e�Z+y@�i��8�y�J��z�Aw��)۰yA#m���y#*~�U6�Y-N8�x�B��y�I�j�	�IL�>����-K<�y���d `�!��&X�x���ݠ�y����#�����լ��,X���0�y��<+$f��DĶr���Ʈ�yb!�H�TsG�N�,��G���y2aB/Ӗ���JD֘M��,�y��Q/Z�A�B�8�Je��K��yҋ�1 P�}0��}��j%���y�/3��xQ/.!�y�Q&X
�y��Y���A�k�l�P��%�y�A؋-g���D�^�j������y���o��a�#BH*��M�פ�(�yf�!z���U�Q�F�ضaA%�yB/ɥ4s<�k��I(	]f���B���y��	
���G� "U��#�yr�)VjB8�q��sQؽJԪ���y�/��^_�8qn	e����y��-Hit)�"���b����"���y�)
GCP��7菶F&�1;R�/�y2Ǆ,HL���"�=�p��am@"�yR��9��Uv ��u����y�Õ6\�RB�9 m��hЊ�y
� �i�ì�Q��<Aըϣ8�bT��"O��q��������%��y�"Ol��C���숡Mh��U�P"O�=1�c_"�����ձf�^=G"O�d�ԣ�'^n���ޥ_��U��"O�5ˤQ&_���A�y�ؤە"O"�CکT���֛j�F�;6"O�� �"]7KW��kϫ"���A"O�1А�H1O�ᐥ�!�A!Q"O�e�q�T.X���+�=#�x�3"Oֽ#q
����؃J�0(���"O����Ξ8J����!��=��X�"O4 �p�S���c�)6(J$"O�*d�H;�,9F)�`
|;V"O.|�Z)�2�84"�0���"O�ESF��(��ɹ�T!^�XZ�"O�b�d��"�=��MC�%wF�B�"OlXÏ�!bE�0o��;�"O����E.Z����`"�IR"�"F"O��)B�_��j�[� W0o��p�"O�,�%���4��01�֊oW��[T"Ot)��P�2ON��G�؆q"\2�"O�hjP�F wS�; ��8L�\���"OvQ��ϳp�8���_�q�nS�"Oڃ"�Oe��� �G\�$er�"O��˦�
�$��(qD�	�,B��"O��p�&I(Vi��8��МO�*��3"Oz�U	�Q�.���Ώ�P����"O��`��c��}����}����"O~t�w�H#!��T�%{LX�"OH�'�S y�j	���4C@6�k�"OXIy�mQ�pt�P�Feݨ&8��s"Oʼ;��u]�ńV40�Af"O��k�h����!�gQ`��"O� �R	�*#<�Y.8eJZ1�"O�Qm޹eF~��a�kW��`"O&����u�R����L�|"O�� �	%��ܣ�$0�L��U"O�5Od�i���\�-�t�a�"O츱u�v*H| ���/R��p"OT��+Uj�JՀ��6$�F`�@"OP��u��Qi�i�Eܐ����r"O� �� (l81�FN6R� F"OI��M��s:l���g3�[�"OTd+ �ȸM����`��V��PS"O�d�����x�O$s�3�"O���D;J�椒o��gV,��t"O�t��c
k���Q!l�u��"O~L�O�8;�0���-��K/��"O��!e�	09�{����j�J���"O�8�s��?N�`@4a�;w��x�"O�%P#f��^5b��CX�Sz�q��"O��ؑ�P>u�\���;B�R���"O�����O+t��� 6����!"O~,�w�40�tS�GS��n(�U"OR�XdA�	0ZH*� ��:�氬t�<1���S�p���?�t\#RɖY�<�b`�-"U�h�4.�z�$�ufBA�<�S�ǻ8��\[��[���Zĩ��<"R�-�VԊ��Dj�J�S�Mx�<�q�\�(}�Qo�-�N܂�����y<@� A�,�&��7��y"�Z�e�Mf�Ig�Ѕ��,˦�y���&oR�J#���^e��bI�y
� ���h�88�y	3ꊉ\�eS"Oha��W��H]bU����ɀ�"O��z���Po����S�<��u"O�Y&BG�bK�mR �
.}��T"Oz���H؎�(�U�0~�T���ޟ̘F#3-���'���^?��#e���
%��/>H�6�
�b�l����?��Ha| ���A� Ў�+����J���g�d>���mǩno�PC�Ƒ���x���%ғD@�M���P+*n���oE�O|�T����6Y\
�8%M�;gg�8�rF�.�Pa� �g�T㞠�P@�Ob=o��M������T򸀥�,Z,���ϏY�y��A�S��?I�L�M�X�t��w��bCM����	"�M3W�iț�	�08�
��[���`Jg&���~�G_�u�ʑ���'�2W>Ś6��ܟ|�	ʦݙŕ|z�U�d(߈Qr4k�H�Q�=�d�5s���ѳ�ɮd�P��?y�O��4�ƈ�1���	N��2/Ǵl$��9�M%�?n�0��I(VG�pщ�s�)��L����5��J�q�v,��hڀp�x���*��M�'��4��6�'Y?7��xn�pXRc�9n����5R?���O
��$�2U��f掽{�ؠѵ��r8Q�T:�4^d�6�|B�O���>�"T��Y?`�D���D�9����۟�B�,6�T)�I���	ퟀ���H7m�21	��A�-�TUZ�Bͪ|���b�&��p],�8X���m��?�c�IW���F�u/p|��ɔO"�i�ק�n xgÊ5G*�0ig$�~B��!#Vp����<q�$h�D�٤	]�wu�e�7�;w�oԙM��|��8q���I��'m\�s'g��?���O&�����'W$�����A��� bX�y<��qe@Ŧ�Yߴ�䓝��'��DR�/:��c�:M�^|ZՅ�=��i��aU0a0���O>�D�O�����O����O�I� �׿
qX<Ҵ�f��\�%��=����-ɦi�E�A�o�Z������$Z4�y5/M3%��Xe��/R�U��-���d��b�a�Z��R�۾Z�ryCwBۇ��'������M["
��=w��еf�:cʚ��B���%��O��DK��֝�|:"�Kt ��!�R4I��ț7&Kv�<	�$��1�&�ã�ιj��PC4�o?���i��6�<�b����'��_?9��(�	j���r5JX!)��sՠ�������?��_A��)S�D�X�vl;6�֖#GTQ�&fy>e���+BL��D�5��@1�2� ��P�0�Ѻ0���xRe�q�ht	CO�3��C@�2�SU�t<+�$Q6$�����{�h��?Y��i��O��桅�#p�L��f�1+m���� �]��.�)*�}baa r\ ��z�����
�p>��i^B6�l��hȠ�_(:{2d
g�,�����~b���7m�O��$�|J�-D��?���MK�R�#�A:�2d���Ꙉ4଱�Aƕ�1�*�:5���B�h�H�-�V�)|����N�:A��c�YŤ%YE�a�r5Zs���_�<��s��/�t=8�M٥5��ʊ���s�e�5*,��ٚafPhײ�t�~�D���'��6X��Io��MnN-I�� sFMFe���� ��v?��?�����O�c?kG�[	o�N�8E__d	�"�7ʓR��i��'h���FR=9V�M���ڲ)�2A���O>Iۓ,�1�  @�?    �    �  *  l!  �'  )   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic�'��}9�n�<Y'��{*�Q놏 $n��V(�u�<����8#¢][G�ÿr�(�@� �Lܓ^�XFDFQ?!�f���E8"	Q��ۚ3���B��#D����bڥa��a	��+s�����ѫJ��\"�v}R%_��7���t+�.�h�@f!����ƓCI���5�y������w
]+��
�p|�#�J/��{��
��n d
�!�'CX��y' � ���Gh_F�00�Da�H�Xx�3'��Z�A`�Ƣ81!�dK���I�$(7%"5p��"��JEh���+D�mK�+�i�Q>E���b����0&A�������;D��p�KSr@��5iA�f�`ɸV�.7к�3!T�h2��+�lc>c��8�Ԛ>:����C�a[�`��"��:��5w5�ZPJq TD_���0Xw�@3q���a�'����D4�Y0&HÕ>���V�6Yџ�bɈ M��q���eS�]Z��%��� �q��ZU9��&4��1㌐� &T��ʏ8&��	A1�<�T��b��!#�p��9!�k��?���	ڍ�%cIS�  �Ch�O�<���f8�˔A�3�:��u���jЊ�c�+���7MB'3�L~zf�|�I\�,T��&N�1ވ,��l���?�AL�T�l}
$�O�^<5��J�67����Ƈ B����C�(thq��'z�T�A�"|�NE�z���`��@�G���iU����'��^� � ��{g�L�;lh=�#呻g�
��84�b���V�ƘJ�Kɯmμ�#��6?1����[�x�C,���x�Q�"�x�OT2$���B%q��yC��*c���z�'�6�(�nV4a��y����U ��qgbC�ofDrF�i�XȎ?��Ϙ'�	�CE'#$�������H�'�V�F	k�.��E)ߋN(�#��S�?���ҭ��䌂]���#�M�z������t���j-lO�Tp׈^V�SC�Cb� :Ђӝy�Z�	6v���ȓw.di3���S�	����/
��>i�˛�/޸���$�'M�=`(��S�|���ۊ�,��ȓ���`B1� (J@f[Ne8U�Q�O6 A�O��Ȍ�Y��sKٲ<�\("�&�8�hf/#D�$"�iFe,4����xi&�[�{�6̊����&�����E%;��P��()�iC�g��{�ʉd�V�n�$9k��U�T�����6cnh�ȓPlH��@�u����l,��ȓY ��6�ּkےHed�i�p��ȓNX���M�ws�q˄k a	����z��e@Ec�
q�ܘв+��*IX<�ȓ.�(�Z��&>V9(�ˀ�<(�ȓUF�%1�OϜ&�iGeC�P��9�ȓ
8B�FG�8[�	���4e~���E��mcgW�U$�UJ�ɓ�SĶH�ȓ.���*�
����+���:0хȓW٬0F�W;��X4.V�6�T`��Pm*�#�Q�����>\��ͅȓ������<[B�ch�=0-d���s�t�{�n�mɤ�	�hN�Y|����Mx ��U3=�� �e�A�����
8@i�$�C�H5A���\�J9�ȓO�x�����*	�qc\�:��ф�Io2`����΀	��Px�ȓ_
v��l��rXhPѲ� I8vd�ȓ%��=2�Y"=o���ŉ�#!�p=�ȓ����!�"E>)�c�?;�ņ��L�p0';��"`h]�z%���[tȕ�U�W�T¾��@BJ�B݅ȓl{���J$t;tu����	����<����4�^�#%Ra�w�ƈ}A�\��n?���R2#�)�!@gM2U��;��*�"fc@M"�e�B)d��ȓ ���`��U%Nz�ً +6�m�ȓ4��\#'$��݉+Կ^�d%�ȓ�� ���C(d����d����(D��a�EI�J~8�3��|���3�`6D��1F�ŘW�������yT�q�UD/D�,"bB�GD���Z�k�}B$.D���TJ�BI(����Y(Q�̐;�+D�x)�ήeP��t���S{�Xb�M$D�H� dޜG�X�)G�O|D��Qa#D�0�F)5C�(���M	M��rs�"D����ȁ@��(��b�����{��+D��idN��+�ݨ�N48t�bDL*D�T0c珓C�HQ���cj6="�-D�P�Ӊ¸<9ܜJ�̝H0�Y%-+D���+��c�ĉr���K�U�a�;D�X`V��c,��P.��t�u��8D�4{B���>�0T+�����"xAq�&D�(PV�Y�h#��#B^&?�ܫ �%D�P0ր� _���z�a��>��<X��"D�H�+.`��H�%lk�4CpN D�����%||�Qu!ޜK�$��*D�1JQ�pm~:��7'���M5D��rh�6Z���
we۬t+2���>D�� ��{!��_��a!�#�+d�P!�V"Ov8��`.!^@K�G�*+��Բ�"O�y���3�̨2��a�$��3"Ot��D៭V{�I�'-L�T� ��"O�1��G�}����r�l"O�Ck̯	l�1���\Z�E��"O"�r���pj8�@!��!G�كe"O����vg*y+c�<C�$��"O�8 �f��.��UE\1r5$@��p.&��fS`X� j�GX�d��0��<���N��y���w��Ĳ�ʃ=�P];��O��y��A�$-"6d��7�� '�W9�y�gI�h��C��y,(TѦ� �y"�èz��4��� �i+Q
G��y"�8~p����D���?�yreJ7>g|��`�ɉr$���&� �yb��qi(Iz�I	�<9���;�y�ҏon>��)��w���rw��y��Dd��n׽u�� f���y2+�h����qDx��EE��y⭀Gb�Y"Nĺ�0�#5����yB"ɦ:��T�����d|%�$MW��y�AA*4��'�
�斐8ĴЄȓm�M �o�r@�pΔj�!����X�h��>��Ҧ,�J�X����p�C�и�ƭ��H�W+,��n�H���@�Q��U{�Q!���C�����P�#14�:�嗄-,.̅ȓ[�|pˢo�Ƹ��sV&@��C�9e���8v�ί<| ��6HQ�o��B�"M��q���s.	��"�B�	w��Ā�,H d����(O(E��B䉞_��� P2'���Y���B�I\$�CB-T$n���
�I�o�&B�ɯŔ5p0�G�RX�"cC�q��C�I�$��ܰ��*>䠙��`��C��E���p���"h��	�JP�}��C�Ɍ>��m� ����Ȩ��-У{��C䉇2��馬ɨ'ФkՊ�}�C�4T.�Hy�E	2�����3ӒC�I ]e�Q��`Җ* N�C��.-�C��������<Epbt�L�9�C�I�e�@��V���$�ġ��4D�vH�����B(�dB��S��!�.Dߢ�Yb��(Q°=��ߜS�!�B�Ff��*�F�����
3�!�0P�4�XscR�Rj���Ԉ) �!��"E�p#��mep1A��L?�!�D	�1�b�C���F�x��ͻ�!��d_��f��*��)�B�Wm!�DǙG�8���Y�?]�I�d���3>!��8g�� �ŋ:Vd��"�!��&`�zz�%̘H6@��ƅ�d�<�բ��	2�����[�'�`��0�]�<I� ��y#4T�G�R���:��b�<i�m��F��D�b��b��Z��w�<)��t�rU�Է9��QB�*�^�<�3�C�z��	4��=(�|uaԪ�Y�<���Q���8��M/%��
XR�<��
[
vx���w"֬n����M�P�<���1>�T�"S'\�!]�� -�L�<����GYI��BK��f�*�`�F�<YUʎ^a�p``�0eQ2�1�E�<�bZ�vg e�3l�4Y`��HYB�<� ��h�#˼~c��Ġ��)�l��r"O�!g~���" �3n�f�Q�"O�M���ϛ,�-��H,g�H��e"O���� w��-I�ak{��
�"O��)��9:�.ik5'_�AZ�qg"Of49b��X7j���'+P'X�`"O�;D�ޤ��!ADa
>�2���"Oč3�U��D�@"S�C�d4��"O���2b��2�����~@H"O2�`a蓲S���a5G0j�LP�"OD�"���պ�I��˦}:�(""OjT��
�����@�W"�̈�"O�AHba�63���A툢[|M�r"OQ�p#�UY�e�K�J
й*�"O�
�`��mbpiV��6G���1"O�����{'��l�
7X�&"O �ǲ���"���5��x����{�<��LW'E���*G#wE@e��D^�<����S{�D��.Ω4�2<Aq�V�<с�^=i8���,�~� ��GK�<�S*�������_$d���m�<��U�Ot�$9�G�&~MR�Ǚk�<�Ǣ����u�<hsjա��Ep�<��
�	���/Ѱg�)�7�m�<DD�\�3�V�I��� W��h�<A �A��H�& E��� d��h�<��08u|	��bـYo:]�%�AN�<�dNU5g�vD���U�2���$�J�<�4�F�e���0�9O�<|;vi�<�e����*�
� T<X }2�J�F�<��a�=^=D���EF��ph�C�UY�<a�I�s��0�'�R#u��b�E�R�<IP�R>h0��AE�j��P�j�<��/�8h��1�+�U�ĠH�d�<�4��:$�����]}c~!�`�{�<y�
^� �ѺWFr���x�<�n���!�MT*"q�Ar�<I�)��
D� tѨa���o�<�r��x�*pQ�I
��Ih�<Q��WX��9�<A�fձ@El�<�e�V7Cu�����	� �|`y&B�f�<��IӔDA�q`a�*& �'�e�<�� �i-ԑ��E�<����I�|�<��a �^�\{r�����K��N�<�&�Њh��Ay�KH�	m`�&��<!�bV�AWE+���/�H�aMy�<��%�"}T��(�)C�N C��Wy�<����sH�H�-�q~��D)�x�<�� �9G��M9@T�'�s�<1sծz{�$�QA��j��ܘ���E�<���B?�����8�^\3��K�<Q��R#]���w���Z�z�('H�C�<5n_�BAB�[FƼk-�s�N�g�<9f��/]+6�ؠIX�2�izw�k�<���
����{�P;U�:�p@��5�察=��C�JՂ �����Y���q�9 ����p�F�Dވ�ȓ%�lHQ҆� Q>ecVg�9 ��ȓY18e��N����+��L�<�0��ȓk�Ђw͝�0\���$^��hl�ȓb5QcD�]pp�"�F_�>I�Ԅȓ��a��4��]��P8U�@��XQ����\���K�no�!�ȓB������?z���F
�3X�A��S�? ���6���z�X;3 �,����"O�%�+��frv�1 _�� `�"OT0���>夘+`�� �����"OԨ��bޗ6��Qf-Ț*��Б�"O<t�l����ҩd����"Od�S�)^�E�J1��,�

�f��u"O�ڃ���0���!l*cb��T"ON	�/�7 ��I�!�;F��"O*X!��M C����O�;.�P�"O\ub�B��#�<W�QpvXK�"O�I1	�f1*�c���0� �g"O��($iT�o�R�q���#�H�"O�I��PAZ���t���n;� D"Ox���,P��`<(�����T��"O�e(�̎?V���AG�*<�=�"O�}�$�н=:�Tc�+Q
%m�0�"O^���`܋-*f�[�k��Z\	��"O@Q��һAd�1A(�85N`"O���5�Ί-;|��ǒ�4�"�#�"O�)�c��5c�|�D��h���d"O8<�����Ȗ�� �%"	2"OЌ��OG�˾1Ƞo�6l��)$"O(����ϵm�V�B $��h�H��"Odmӥ�?D�FV�ԄG� ���"O.�Bf�20)
�$E��h�"Ol3Ԇտal�I�"_�y� �r'"O�x�ң]�pg��˯&�xt[1"O����ӄ'x�$��EF3>\�U"O:�pr��p��I!��<N��M�`"O8�+K�xo�ɳ����*[&"O�8�pΓ�Z�q*�A݁��h�G"OV��V�ˆOPJ%���B�	!��"O��z�G^�A{�E�'Ƽ{��"O\0��	�F��L`R�R�.g"H�E"O��e�Q)ڔs&d9"bܭ��"Odd���LBW|����-f^
�Ac"Ot]����,��	��V�[C.���"OB�c���x��3����"O��V�!E������~����"OF]��E]�kJ�J�%Z���\� "O��
�f�nĜar���5fD[R"O��Y��� �̡@f�H�ZF���"O^�x��Զ��12�jƟ0;*4T"O|X[ �p|��!ꅺh:i '"O�	��i��#��hy
����s"OXS�,�1[Q�zgh�%��A�"OvY��IhT�U����u�"P��"O>���Q&RQ�
��
h�.Xٗ"Oj�"�Xn�2���;6|ap#"OJ��U-�9r�"��`�݄A7��F"O.dQ�K.Y[���@,ʪH��0"O�P'��&�Jg+E1)g
�В"Oq �7~j.�+R�_�vN��C"O�,I��)#9������`e,�xA"Oa��-X3�ȕ:�iM�iJpDc�"O��⒋Vh��Y���u�6{�"O�]SsH�eD�Y���ʹL�d�E"OF���G]�1�*,�eF��_> m�@"O� (b*�#<.Er�'1���g"O���F&l�W�Q�Qj�\	"O`��F�Ow!��`%0]�%"O���V�l ɂsC]�r(J��"O	*��Ԑ�hԍH� �xU"O$�1��2�n@�Ӡ߂	� ��"O� h���Ӏ1~�ڧj	%,��H�"O�d���V,*���B�A+D���"O<@S��H4W[�&0�q`�"O��ДI���꟝1���H�"Oj�s��(,��J�,V"]"O:xV$� �gI[�)� ���"O�ܹ�h�	`v��c�ԻCB�q��"O��S�B�pl�\�6��9��"O�]Z%�n)>Q*��Z���"O��A�H�Y(�#ō����˥"O���5	ޚ&�P6K�<�t�Җ"O�����V~.�X�q$G _�t��"Oҙ@��FR�|��]�%��ܳ�"O����	�  �P   >
  �  y  !  �(  g1  �7  �=  JD  �J  NR  �X  _  Ge  �k  �q  x  T~  b�   `� u�	����Zv)C�'ll\�0�Ez+�D:�DlӨl��>O$���'h4�l�^����Ο�0����S{Ȭe�2l�#K+����!cݑ�6E��?�:����?呀dYL�D��D ]���K�d�W�jEɂǓjU)ՠ(4�HDh�u��l)Q�'�?����V�rt	�[�9���股"�n�# �6R��$PC>���%	�}��6��m����O����O�����Xd�� ��B*)uz}�@AV9M�~��O�Di�(�O���?)�e�?����?auI�z�P��H�8r�GD
�?���p��v�'�"�'���N���'>�$�A�xs�+h�,a`P�K��4OV%+GjڶoՐ�+�*�& ��\�dDxR�O~�P(C���ҷ�y�+[��z�ϸ ���'�r�'PR�'+��'�����SS��;y&�H�g�XU�,��o��<i۴g]�Nr�VTl��q�4`_�li�i%>����'�n��2��טas��I�W�6�0�Q�DA�{bW?��$�ծ?3ĘrG��c��8����"I�<8�#C�se�r�k]��H�4cL�f�O��4�@�D�t�%ޮ8�}�ˑ�Q�2��vg��<<�7�`0̓'j�-Z��@���7X���ݩ~�F�n��M㑽i,�#�Ή�yM�鷭�S~m�U.F���Q�'��~�(6m�����4z+��S��
�}�Z����b���`��M������>�lC񫕈-'�QٵhM�;~���i�z7mɦSc�ةO�ބ{@D�D|���>�R�O�!k��T�d],rdP�ش ��M�'�S�p���K�N*CU>x2���'R��%��a�r!S�]l�u���'��O����O���#����O�t�7�D�4��8��V^:�������D�Oz��n>�hB��%5FV!�E���] �$�
+%�U�f�N��4.�n5�"O�ł0l־R#�E9t��f���Z�����OM�N��\��p]��'�ZP���?!�W����@�(t��1��f4�c�O,�d�Ob�b>M�^�~���3{�}��f��N��?a��4���n�7��k��?l4JTCjLCJ�K۴��',�s������5�T-����O�<p��j@�=D����R� �(L����QЁ��c;D�Bs�J�Xkv]sD.TH�!�u�;D��#��;*H}ؔ��3$��m!�7D��V �5O��8�7�� ��%�7�3D���Ԍ�7Vx�� �,���O���r�)�'V�Б4\>V����tM�5x�'{2��%�ː�r�8���:pn�)1�'ሤ�`���ܬ ��f<�ٛ�'~Ɓf��pA|A��\!3�|5��'c���e��F@���31�r�	�'5X,�8o�<Y��[�-2)OB���'�1c!U~�  ��O��C�'MLP�Y#^� ppc�R ����'&P�@CX�I�F�:��*�B}��'�
I0q�HD���Z�'����'Z.� ���F� 2u��(?��ϓUYp�{��i7��:�V�X�͊�G_���ׇ²}<��D�<����?��Ot�Ɋ����M�@�$)���2��pH�M4����D ͯ3�ax�`�n9(T�ý6��)�TN�}���6�*)�Ƌ\
s�0qa������	��Mk�x�9Ks�]��.���
�/`��,A(Op��2�)�'x��c�Ä�_��I��!���?����h�(l�`,�2�mz^�%Y"�Ԇ5kr�K�4��k���`�S��'����8l��y�Į'H��cr��(1�!��Y:i��R��y�
T��@ w�!�ē�\2y�F���x��ī^�!�D
솰��5�2Q��̎�,r!�dD5 �t`嬀�|���V�Oh!��A�=) \�G#i�`TP6�%�۵~����O��$�O�˓�z��I�:���B�ţZ�����Y4�$���,ؖ�֏���i'_M �+Ԧ�_��$e�˵&Z�T����R�Y��C�a��|S�a�Ļq�b���'���BաR��Z���*ܡ�^pɡ�蓮{,OmHE�'1���'8b���X|�nH#A��-��ă�H��y��(���͘��X
F�>��*�8����O~�l<�M�I>�'�R(O81�
n���+��N|
���\�Y��O��O��Hݺk���?��OQ�0�cA�2�ak� {�.M��'���xϓslL{c�Z9Y�Z\����)��d
�'dLKS	ެ#��L�8WnB����@�?��'#�h[�lT9.�T���$��'	���a��u?8ä�$��J>9S�i7�'�� f�t�x�����ī�W5<u�E��Ih���Zy�'O�'{�!��Y�x6*1	��_�F�� 6)�FO��Ʀ�hr��w'����'��Uk��@)2���y���?Ҟ��g�ǃ.�8Y0�#�0<��l��[�4�?���=��T���!es���£ڶu��4����?���?I���䧡�'�FY�P��#f2�Q��F�?�l0��)�a�^U��E�?lp�p���?A-O`������IßL�O�����'09�IĚ|���⥊>r�(5	��'�R!��:��T>�'��(�f��B��dp�d[�t�ܥ�Ob]���)�' �a���b,�!Rn��,
�'�Pr��>+ɧ��Mۃ��:NVl<XCfM�jw �0r"Oj�VK.t�������]Z�ٴ�	K}��9ғZZX�:��d ��XD�	����im��'�rE1��l#��'���'Gb5����#\5K32�k��=,���A��d
&�azb	
mn�����K'�4 %c�/Ә'���W��(r5��.B��SFT(1����M>�F����|�<�qA�(�$y���
��81]Z�<qb'		� x�H���i�CƬ���t�����|��:o,�`�K<^�䄱V ��>�H��X46�B�')�'g*����$�	ҟV֞ �B�uZ٢$KW�46@�RD�r���G�s��ݘU
�#>T�E��LQ<OG��VnUm�ȝ�0c� ����ĕm�h�8�(U�pH��(z\R��'$T7�En��?�����M�dو�(W�|�*-X���*t�R�|R�'��O�1O�c׏߼:�2i�wIg�h�]�x�	��M3��򄎴*�F�nZٟ��ɬ}m��W)D�δQ��H�2���I�����L؟�I���B�H4lxL`x�O��*v#����w3���B�j��/#O`q�I�� "4� ���7Lq�an�K�j�Pr�D�X{l`'`T�i����ǒkT��'C�7m�O~����]G�Z����8=>��VȨ<���������
�o$ ��B*
J�ƴ	SH�..�	�����k�S�-�Or�r��Q�G:��X�h�1ʬ͑�'d�ɶ.�,��4�?���?I�'9OIc�
����-�qo^�#��'��x���?����*h���|*����h���Ƅ ��5���3<�$D�'e��� Pɧ��Y:�Z�{����l�%�x��'��0�(�OF���O���6�'	�8c�GF�\H『S�B��%���D��b�eL�XH�i���JHT6.8�����X�'c���GLڢhˢ���ɀ�3� %��ljӌ���O��D��=�,�D�O��d�O���y�y��T�p�C$�'l�L�ɣ9,����7�3�-"`�`aV��A)D�'��J�4TDnc>c����D�������Z.�iJ���O���O����Oc>��?!�M��l�#g�	W`2��N�y��� 	6����g
=O�(!��~o�	��HO���Oʓ\�ԕ��oB�O(f����U,
�rH��\9���'�B�'��Ig�8]��x�f�=Fm�`4��
��Ā�SGL�8J�g+~���_5T�^��!���v�EH� <��zd聊-6>�Cd�':6)"&b�wr�a�Z�Ԥ"�#ͳ�?��6>�v�'�I؟��?ɓj�",�R��=����k҉�?����O���&扶ik��. |��� �n(˓�?i�T���'�ѐ�`i����r�L�LR�F=@���w������O��?����?�$䊙bi�0#�ԿY�RX��',���"��G��ס8 ���Ó>�ƥ��d]�
�a
��	b��#��*.&<�s
]�u�h�����0<a!�	ğ<�޴�?���(�\-�cb��ð�����. �~0C��?��?����'b��F��;�,�`�+���8��i>����Y)�Ұztʤc'O�����	qy���I*L6m.�	}>�lߟ\1tb��W�h�+��A81g�a������$=�:p�X�d��S����fM�&<�.�ZA`���?x  `�'�\T#7�1F���a-]���#}"�$?�t@��	\���VdO~b���?i�iF�6��O #|
QdM-h׌LKS�G�De6\��ZA�Iɟ���@����eҦn86�U�2?.%cΘ��hO��D�˦I�ڴ��a�֑`u��RS��@O�j@���)�6�Ў��(OD݋�F�,�<�	��Eq�P%��"O|�f���|N$h�*x�ڭ�"O����JV�G\la��@�<&q�Qc"OV9�%8&����@@�ZTX-8�"O��X�?�>�ق��  l�� �"O^mjL5)�e�$��!jQ((��P�X�a�-�OF�)���b3L�IQ�/7Z�p��"O� h��U@�Q>� ��� h�H�3"O�0+��K(-��Х��8��i��"O��P�gF/nO�Qf�)l�JT	�"O���*�X�L�;Rf@�@����'�>,��'3D��瑐<��HӃ.��#Ur}��'�́sfP�i�f��Н!����'��]��k�`�ฉ��+q���x�'��"�ǣ7P���EꒈW�:���'�.\+��3A*u{ Ȝ�w�`��',���`j�a�ج��˅* �ؕ�����4TQ?i�'%M�B��P�Tj��J�Gf���y�i��dn���Ӭ���D�S��	�yd�X���`%G-�by��#G&�y��¸8ƨ�i�ݥ�l1A��2�y�L�	o�9���عL�H飕���y��k�J��%L�@d0����?A!G�N�������2�$@��l�e�n�j�3�m,D�H��A�snL�3�o�F��d*D�z��Y�/�XZV�P�&vt���'D�0x��N*,�IenI�
�$�
�!D��x���&k-��w��Q`<�!sA+D��:@R�!#�Ɨ��M���<qc�w8�$��� &(��ao�1��n=D���1>n	��mS�k�`YxpH'D�lk�O�v��wM�Xޜ�1�'D�HH�%9=R�Y�&�3E#^C�!9D�����cR��#`F���B�f6�O��2��O2��	[2���c�[��U@�"OH$�s ωJ��y� �ŕ{�|�r�"O|�����-�0+�V6e�R�e"OZ����X�]�b��a�!~b4 ��'����",!�X�A�띙*h��)�'�`��nA�b+\<�v��D��e�'h�<k���@44��q��I�����փY�!���|�z��2bI��<	`�Iȥl�!�D�Wc,��tK)ߊ :rɖ$
�!�D��zl�"�J�f�Y3HQd!�䅡L�e�tʑ+-��!Y� �i!�d�#J|���!�Z�OC(J��v�2����O?�F*�P�Xq�Ȍ<G,�CӏA@�<aĦ��]���G���,�+��}�<����I~���	.�Ȃ@�x�<���ܼ|W����� ���k4�q�<�3MK�& J�3ƂH<���S���n�<饁�.5������g��k�g�hy���p>1�`ڌ8���a#��q��!�Rf�<�F��sn�J�7'%����i�<����CQT�Ǉ�2�2��	e�<�r�D<\?����$#鐽h��X^�<�1��c�9v���	�8�kS�Wx�<��%���b��kְ ��@5(���W#%D��x�
�t�p�hg���Йy4O6D�< �k]�H�� �DhݒM}���'3D�4{�-F�jq��ɱ(��4<���1D��
u�)3�&Q���c�R�H� *D� �s�]7Ȭ��+�'yc��贋=ړ	�aD�D��7'�(��#�V#�4�c�����y"KV��r��PE�e��a�Q� ��y�Iӈn�1p��T�N�^ܺ�)Ϯ�yBĖ�P��(�w�uJ0��qѪ�y�BL�3�ЙA�i�}XQj��y2��\�����6Y�����,�'�?1R'E����r�#q� :\��0#�%c<�-D���ĭI��A��#Z*� �8D�� T�� @�-�`X� dB�)8��"O�����ӻ1�p�c㋔V���"Oڸ�P��� �ĸ14�=b�L�F"Od�:�o �([qD�^�l���P���W�:�O���EA��zCҕb�L��c�^��s"OL�� 
I#B� �2� 5d0�ˑ"O������0N, P���`ﺀ�&"O�;Qe	[�x�$�/�f�c0"O��Q1 �O��H����(���Hc�'Ym��'�@�R#ѩ/�������蝲�'}.���@ڛf�	D�J���k
�'w�);B� `�>�Ҥ`�<5�M��'Y�Ѓe�[�~y�G獮%چTS�'�
H	q�L�!ئ.�'uˎ���'U��S���I�t,HUΌ<mG^*��D�*Q?S�E�{cF����R�dx�c-D���*L��T�F�C�l�[�,D�L@�
�p,�A2��@�`�{t`*D�@���$p<m 1�gZ4(�(D���"d�hb̄�w���k8�ZaK(D��S�#_"E���&�H�[�
�p��OةS�)�|���JʃT��B"�+3d�1	�'V�I`.��8I'���Ѓ�'	��z ���i(Wm���
�'��e��SED�������2��
�'��p��˕7+�`aā�b�,I�'�r�����8�HꆄJ�0���,O���'��=2 ���pa���P�Q��8�'�t�S��\�3n�Y ҨL�Zcj��'����C(�V)�r�l�Dʬi
�' ��E��0`���P@�'>2��a	�'_Zi����N��ȗFȵl%�ݢ��\ ��v#��zUϮ>�6L���zs<i�ȓ�*�c�B(�8�/Ӷ;��i��f�nH��-���>%�SI�-#���ȓ3��9��cSp���UE�14Z��ȓ0�\Y�iX�z�5���҈����&��ө�	e���K�C�LuV�G{a�����(D*�rt��"�V�7�B���"Oެ���.D�H ���,���ҵ"O�U#1	�A�ly��[[�@43�"ON�:�/�sɤ�� n�;d�8��B"OH8�U�(Pb�)A��X�0fl�"OZ����ܵ�c7哟(-�� s�'2� ���;o�d:u�S)r��(�Q��	LH���_쎼�땇P����/d�D�ȓ��5;�	H�b.�!�� RS����Q_|D�S�QJ�p�b0#N�)����{��� k��1�B6|�F�ȓm�,1�b���-0�%�',T�+X@=�'�H=�	�@S�`Xp`پ�pH�@m�' ���
�	�ʋ|	S�}����ȓUI����ρ2wfZ��!C�4��\��S�`�!V^�ZJ΍:�d�P]�ȅ�9�����۵}T<�H�&Ͻ.�����	QaV�I4 �~q���/O40b�B�%,E�B�ɭ|�f��uiV4V���"EūU�B�I� �p��E��;$����>	\LC�	<^�Tx�F	Aj ��+�E�C�	�O�faa_�d��=Yc
��sY�B�%O!>����ߓcV(����K���=i�&�w�O��H�g���;���ˇE��T���'�,�K�"�6'�p�!�ӱy,P�'�]cbM�!V�|y�Ώ j�<���� :t+ �n��Z��V<i�ݳ�"O�[m\�}RHx˰"ۋS�	�"Oz�:f̩7Z$	j�!\/�Uq��'�>a����	ePP$�ōJ r�����oNX�ȓ�z�`6,CE]$\p���j��хȓm>z5��J�4g�`��Y�"ͅ�H,�${U�İ0���[F��<'J���2�8�X�g�xx�� �9�jX�ȓZ�X�;C�J�(T˖�]�'����R����R8(�����/F6^u�хȓrEP;�!�6!��`�A���<N��ȓ:���:��G��:�,'[~���6�1����N ���#&j5 ���P5l�Е`З2cB��Q��;�х��8Dx��=���D��|x��􌂔0��B�	�2æȱb��ZUړ��z>�B�ɸ���P�M�	B$Ԩ�� �BC�I�\/U���߯x|X ��E�!)zC䉹p+D9�����n@걳`Ƀ�L&(B�	�+�r� o��Z,�	��/r��=�	UP�OD~����J?�(��ϹF�dt
�'z��3�	.R��C���1	���
�'�έ*wc�L������x4�
�'�ʽ#W�IB��`,E�l�]	�'�p-R��T�T<�2��=��UJ�'+F���D�"1P���%����#��*�Ex���gK6Me�ʲ^��P��>�C�I��]�"Iȅ?R�Ps@/Q2+��B�I�\Yd�Y�ǂ����L�kӘC�IFŞ��#�&�2|Уe�'cs�C�p/R{D�lh�f��y7tC�ɫ �����њq<@ApT���6�*h�	�Y@�I#GH]�z�]93$�����C�������>u\1 �LW)p:�h���D�	�f1t���ȟ0�I���E�1C!�a�#N�O���P����9`e��AĕC9��@�\�΄���K�:���O�)��#z�n���L��������#E�b�'�1����@�.{�Ȱ[�a�&@`4���Q���	F��ӱI�(9�l{6�	�j��!�O`�'ϰi;ԭrJ̹ᅓ�mG �4\��4�Oן���/L�h�O�N�f�O�rN��%��E���eF���c	��O��k���X�↨/YT��3��O��Q̧4̄��¤�wJ	)0f����Γ#Ҹ	4�P�1C�#҈T4�蟸���HP�n��D��"�t�Ay�8O
y���'b��������D���Y�#±~���ȓz���х Y�b�@��-%�Z�D{�M!�8905�֫ʤkh���o�!���*`��?��"�Ր�+C,�����?��%��n�O���a'�? ��EI�fMuA^與�݀$ hE
�	�!�h�� f�O���oB6I��Q�	ٝ�b�[������2K�?�NeX��ڳT�S-��'�]+4�(�1�G�0a�,�K�O�;2�'�2�I�<1Yk�k؃9Ӓ=(S�(fC�ɒ'�l[6*O�%���H�"/@B�$	O�����'1O��q'��Z��U��
@J�q��'�����ĵz`��$PK���
�=g�]�ȓ?�$iD`��*-6 �+�<a*L��v&,��M��d��(�"!���ȓ=�J��5aƚD���#ݤ&PXŅ�Q�ac�
F�-Ra�ZB��+6|ON�ꢚ>�q��SETE��a����5���_�<a��z�KN3�s SY�B�	*����A�3��O�U�TK
�'hd�9d��%C8�K�/Q���	�'���j����,��Ĉ��]��,2	�'��aWm���H��� '#J�Ј���O�'hB�QA��&x�@bȗ��`��ȓw��3օ�4����HK�q"�y�ȓ7^��ѡ��4�VձF�T=|��S�? 2܃�!ҪD�j�&��-h�PP�q"O)��?7xD��B�E�,�qE"O���5�,_88�H�jʹo�N�:�E%�OB�}�TB���%�J;���"D��O(j���L���B�Ǩ������`�dU��B!�x�"��{M0E��bŀ�С��e�N�r�o
.f���!�@G ^0�@�ȓ�T�a�ٻ3��QY��D?>���fp���(؛!V*]�VL�=%�u��7t|��DF���31"@2pĄ�"b��9=!�$�:746dț�h����j��C䉍�&��TC�-�9��OŖM'JB�m��e{ˀ�<����@�X'T�PB�	�4����b�$E>ݒ��R4]�?YW�D����'�R4��dC �����$*͖P�̓��'�j���'�B�'�t�J�/K10���?y�O��@�#i�N.��@����h!`���R�2�	Q�/�/���`fp�t�K�s	mzW�;\d�G����O�}�v�'yb�g���$|>M�Wǟ�O¹K��� C��.���O����z�']�|'C�96	 �y��?j�b��?i������i�_}2���r��q�J'�~$���V3j��'���'��ɟ4�IZ~����8Eq/�lG���R�L��0<y��X�z���H܎$�
���c�9/�Ov6�1�I���'d�(���I�D�����R��A�iyB@èX��d�w�B�'���';���t�m�L�]�V�z7�ڽt��-:b}���d�*[ �|����?7������5��^O�H�P�4KH�{v@���M�IҟL�����<�YwlB�'���'�$��a��0ē#�ҡ`�o�\F�'|-]���<O�8�۟�^w!�z�*$�c�/�x�6��BkЈ�I38�>���O�t�O��'(��OjB!�s���0,Z�qx��8�z� ���<R�'��y�@�'��w؟�^w6��=.��@Q�lX�ٲ�5H��7M`���M�O���_�~�Sٟ����?(W뙰*�I TnǭrH4Hȑ�G� �BϓD�t ��˟�
Xw�21O��0���46m�A�Hҥ��-!z�P�6���mj���O�扵oR�D�O�X�՟?���ɟ|�t�$<�x�"�k��A&nG�M��۵�yM�>�?���2���y¬������9����P�\����ps�6*H���Q2x�P����ܟb>�l��A�v��K��lz,n�� �ȓ��xf-D�"�����F�NalZڟ���y��'��'�^>�حR��)�J�U��d`�t�h6-�O>�D�O��$�Ot���OX���Ot�D@0%p�0*��p�H��v�LM���lRy��'��T�ByB�Q;O�bгA�F�V[&��3��g��)���2t,��l}��7F�0Fh (��d�>��|��q;�&]k�2u��Aa)xQ�ȓ4i:b@�]Ύ�uJS�H��C�s���`���U�V��0��|��C���؁{af�p���!0)ʣI�<B�I|r�; K�%O0{&���B�	�N���# R<|y��TI�C�I'4@���7Z��Ҵe�%SD.B��^ Fy%��(V��h�,),�B�	�&^R4:1mR�9t�q�� �8B�	�LL��!�B�dR��6J��;�b�t �� 8�<��*��ӌE�!�ح�|`cH"����j
�VJQ.ה?�$mQs	͘;��@��$5�Z��0���8|X0l�">����)؊������"^��!e��K�r�a4�?dA�`�*F��X���L�@*��y|�y��y�9(�y&S�m�0e� N�&r������"�y��ɏG�lY�D�BJ�r�nӜ�y���Px�a�(I� �S��Z��yBaW* ��R����A�H< �@�y���J�FP���D���c�n�?�y�䔴 |�jR�Ƨh:(M+��;�y���50�*��u�̳^즱k�I��y�.V��<��MG�X%��Ȓ,X�y��֖n[�-�ql��d%��A��6�yB��"	v���`��&�Tea�݇�y��6B��0���Bu��,�y� �F]�5+p��p�����yc�L��p�-M�44�J�#�y
� pHUcHY=L`��̆A����r"O�xЄ:��#3�	+e$U�t"O��q���,k����-F�9�V"O8Y��7<Z�z�g >����"O)���գT9��!��%n���"OX飑`û8�>�Q�l�u~HP��"O2[�d�@� �G� 8L,�Hg"O���F#�"{ ��n��k��lI�"O �h3F�vU��T�L�
7r	��"OP�0�X#+x،�.�$y3S"O^�H��T��i����-R��0"O��*b�ɹjz`=� ��X�PS�"O~(�d�_�_m�L�?Z����"OjQ��@U�����" )("O�z�hI�C0���n�^"�0�"O\�3�O!WCB5y%�w*� �"O^�A4CI+�4m�ʌ�{� ��"On�v�Z;B>PZ�&�7@|J�؀"O.��RC3D�<�/a�0�"O�"�n��[��HG�iV��"Od�����C�ޤ�gl �w�j�0"O隐$��f�P�*vjΟBIZ�[�"O�e+�)�5Ԇ�bs,�V<z\QB"OD�a�[� `��e�_�[� y�"O��`d��Q�0\�f�0y�"Ob�����c����7��zq�uiE"Ot���!�2�M�� �Mf���"O�����KOL����� �#S$��"O�	1��ҽy����O �����"O�bB�)ߎ=Ɇ�,U{�SB"O̅CEF#�:E�u�8bt@#"Of�
��L�A��I���W�\Xq��"OV` ��H�bZB��BR�KZu�"Oހ�偐�l��U��&��(9R��"O��`tBW�|͚D�$&��2d��5"O�iṙ�|i�x��EJ�9�� :�"O���N� ��}AE�w�@�+"O@|���.4x�&��{z 1s3"O4���gv9��)��lC3"OTй2�ͽdT^`:2_-	#D�7"O���bD.0|+��Fp�L�"O����cY$\a
y�ҋ�RX�Xy"Od�l�4�6�[�-�4f�-�6"Ob1� @ۣ8�*��'쏝>K:!�p"Ojغ�n��3��a!Q+N�qj*��a"O*x7.�6;�m����YZ�F"O�h$�Ӌ}� �@ǉ�NM܀0A"On��$��Y� ��ufD%8��a"Ov����ܜ^�^T���ĄDȜ�E"Oȕ"׈ �����Dk��Pw"O�i���%n����T¾p��"O��u��%J4�(*#�"`�BH�s"O\`��+��R��ɩc�<9 �"O��S��
�89 =��Ӈ&�tEҕ"O�,��B�Z���䞷E���B"O�x
�"�!���7��-4����"O�t7���L	2��3V-��"O&�Y��F�)n�E+aP�#�XA��"O�A�hp��3nC%(�0q��"O:E��CK���o��]K�"O�t��+[�R=I� �	��;2"O^�C���X>�4c%��_�VLb�"O����)�"F�%Q&
�V���z�"O@@F��:��qiZ����!"O� � q�aʨr�q�v�Q
��]��"Od���o_z ��j�O�����A�"O��	R��)�&@���G xxe�w"Ou���+�R�f����4�6"O.�B$7h$ 0��A,�z!˒"O:��**���#L�7<�,�!"O��rP��,6*�I&�Q����"O�X3�+܌/؎�����=J�peH�"O��0�Θ3"���u��+Q)�q"OR<p1��N��p�Q��3���)"O�܊����T�0���g���p�"O�����V�<�q���� ~�� "O��䀅�^��`'�^�z�bp"O��E�.wo4�p"K�jZ�1�7"O�Ly2ʙ�!pz�3i�98�1�""O�]���CdO �2��,2-~�ʂ"O�����O)W�V����Ԉ.����"O��r�* 4�޽X�#ε-zܨXu"Oj�� ,2bH8���#oq(�F"OP�k�#�Q��(�S�4)����"O@qA���\	|�K��(y���3"O�hb��E�(`�q**r^��e"O�jb�R=�D%XD
�
'gހ
�"O$�����Q!r�q�k��i3l��"O�q�`�Պ.Z:i2#J�3-rp�!"O�hb��|�ZykP�:��"O)XS�)l�XL�S	_�:��l�f"O��6�Ēc�F<C�:�xeH��y2/^*8J  ���MR�Rԡ5�y�"6���=r>Ԭ� �D��y"+�,@�mtA��j~��H��yB��4L�hT��5[�����U4�y�J%�&u����S���q�\8�y2* 2��=@�ɿ8
B(���yb �%y�T��O�aOX�۵�	��y�;�D�$ǅ�YIV�Q$허�y��T�nZ�-@4�7Y��S@���yr�̓8�)��O'�qR���
�y�C���N 11�Go� ����y���?�6С#V.?��)����yҫ�)gG��a�I� ��:�����y����:�0��ՆuG`�!��yb�`��e!�Z8PF!�����yB��b|@�r�D;0��S����yB�OALvMK��^{t����d�/�y�D��9@Z�[D��e�����X�y��:0�媍e`P#����y���*r2�+ժ�c�Z0�M�yB���x��E�Ҙ_Sj��l��yR�ȋ�bI!�`V�NƮp�V.���y(N�/���-I�MUQ&���y�㋵gH`���j �!KZ��� �!�y�Ǖ�B9@d��#ջ �2� �O-�yR#�e~YqLӛ������y��R-;��x��P���X�����y�k�:�XE;!�O�5���܏�y���&=��1��M<!��կ�yb�L�e�����`���@{�`��yR/Z<<�Xԛ�X&r�L@'oK��y��V�#4 ̹gnM�Wf���gŻ�y���v��U���JT��SW�G�y�Ad����d�Y�<B�\P'����y�!�I�u� ��	3��%�F���yb��m�� P�0|q ���+�y
� ��C���-��`�:@�U �"O���u�ېXc�t�4���n1Fi��"OZ�:1�#p ���m��|)|]�q"O���PCT/0�h�b�#�!����"O��aw����n|Z�A	9רe�!"O�x#�U�,V�-zB+�h� 1Q�"O�Q���E N�����Y�����"O���t�#r�ɒ�i��X��D��"Oh��m�aQ���gS� �1(�"OP�)�-P��ɂF�=c���"Oj�c��/�v	u�X�Ko�T��"OL0��(5.q���S�|�&�T"O,UJ��X�+�`�y���	L�EI�"O�r�!��5d���ʸ��Р'"O.���'a
˄e��w�0���"OZ����JE��	ȫ:��G�>D�P��ͣd#@L�e%I��J`�"D��S��G^@��!(F�[��}��F"D�;Ǌ�-}@���$[�)�B�:D��
��

Kd���oB�=@��2	:D�|ifj�*g3^}x��_Y�pق�;D���b��:�QR._%X���� O+D��Q"o��8���D끃tքq4e&D� �֊�z.d�K3�5\��b7D���F#�u��	��P�̘Qq!*D���E�`����82y��B��&D�X��UT��H4�^>�8!��%D�hӰLB�c��Yj����ktLY��%D�w�9���27�G"c@�Rw�"D�Pp%��V�p�x����z\(��%D�k��g�ι��� �t�h��7� D�� 4���L�*� ��ܕi���>D��Ӆ�^L\u(�	�Y�bD��.D�`7�ֳOa���6���9h".D��y�Ƈ�G�
Ղ!�[�!��H-D��R�<@\9�GaZ!��,D���0`ό����')��q
��),D�иSIY�1��z�WY��g%D�4#Ƥ��*�z�D�.w���P� "D�T�嚯)&�9���Q�8��i�t� D��i�$IQ�l����$
���iv :D��ibo͌@S�y!�&T�^�Xe�9D��B���`�j��6��:�~�sV�*D�\��%^#<��$(0��p�B`o3D��ٴJA�m�:�6�λ1����/D���J#�M��Ig����.D���I�rz�PL�sb:A��+D��S�o� T�����;x.A�3i4D��;��I���Sm��&a9��1D��ZF�Մ�f� l[H�d4D�\y�˃�tK�U��Kص�*dB�-D�İ��G�~H��'b�T�6(D��� ��cܖP�&��a+D�Q�0D�x8v`ӹz$,�!�]�g�Zq�<D�@xwM�E�Rqx��)�DI2Dn(D�D��� b��C�L|�j��v�$D����By�*`�J$ygLD�ӄ7f"�h����'���!�]3��O��aGV
�1���;V���d"O�'.΢/ef�h�F	��ybD"O 4�t�Hnd�f(��\�A"O�pzC܉G4@�J�E`(2��""O����h���#שK�\�r0"O��
��m�Q	�%1pX�"OXAa���r-�`��ܾEZ�@"O� Di��@�S� �í�.e(`��1"O���5�A��h1;wFTyF����"O�m(E�K!V�Ę��dI�E�f� "O�٢P�%p�I9������"O ��2��`i�N�H���"O�P�����a�VhC�?�f��"O�HiQ�>10�뷠�#��QA�"O�-�Uas���C��(.��4�g"O: :
�s��,#�B7-����g"O�,��-˾L�L��0C�����"O���a���QRU)���&b�2Xt"Ol��s �7/����ˁ�R4��"O̼iB�<�Ѕ�К`�2iXU"O8���.
��1Äe��)Y�"O�!�g��:] 2' 6���R"Oly�Q���'rT F^!Q:�""O����ݰD�z�I�OԶ3� [�"OJT`�)�=2�h�C�A*���#3"O��IG!B��|�W�KP�j5
"O|��R/?K�LK���g �1"OZ�r���5�tI��Z�T�N�B�"O�4�EB�=���ق���A�b�
W"O|�3am�5ln��bD�%�"Oz����F�,��ЦE�]�b�C"O��b>v�Q�T�0JW�"O���s�=�8�!/�'^M��c"OpY�B�B�l��ˀ(zGlu�""OA�k�.�pU��Jب���"O,5�#�@�#����4iʻ�J�Qb"O  9�#��J-�HZ0Q���r@"OЬ�RF�[��9�D ��� ""O\��E6#v8��n�r��5�"O(���*Y��.(�D�s6"O"�(��9�(m�eM��D��(��"O�<v昼U��K0�5k��)�"O2��vɐ�ɌՋ��ę~x`�9%"O�����D�bh5I��>�l+q"O3��L� �H�8��5�"O�X1@�c%�p�MH�$��#"Ov�c���&|�����5<��\t"O*��3C��>����Vb��-*�Mz�"O�e��ٟ,��(V���$��B"O���U�ێ+K����;�ej�"O2XР���:ԉ������Ps"O-Z��C�F������/�V�Y�"O�%��L�I�ˣ��Ze#�"O�K���>�ja��Z�*�,�(�"O�X���W�-��
4)�`���"O���⎆�{[T��I3	R��""O XS�d���l��Q
IArQ��"OR%�'�؂8�<�35"�1FA��A"O���2��ddH�C�X�~�@�j"O m �ϚxP�X���VƜ��B"O����H�-^Ei�C�4���Q"O�@Q�a�ҽ��c=hw �f"O��*U�&�"�s��,Q��#�"O4y"0&�!��� �+`�4�i6"Oڸ3�W)9�`J���cΦ�2"O� pmP�	B�ih�i��4��(�"O�$pt�X�b*�D P�{�
5�C"O�9�����lP���.I[e"O8�rw��9V�b)��H�;y0E p"O&A���O=0� ix�n�&h��'"O$t�e�q� �e.7"mV�Q$"O� �����QE`|uئ,	�zg�$�"OB\R#�(h�\�!��+0YP[�"O���wbV�q>(u����2�ib�"OP�*1��_.h�R�[(�0�"O4M`�A�:
�X��BV�|(���"O�	�w�ޜ|uR�2!��}p�Œ#"O���L��o2��;�EO*IX`�c"OX�"c�)�dL	�EA�N�Q��"OXܸ�JR]HX��+�^��0��"O�(24/�!S��ʋ�)��b!"O�tHR�.���IV�C� �^�%"O�����v'��4B�j"O�a��ңBģ��X�}�2Y;�"O�ݩ�f��,4��k��v̂�q"O���Y6P8�)�+��_f 8Cf"O�}�r-rȡ@���fY�	B�"O�T��`��)/H��H�{j��w"O~���K��y!-pR�I0"O�8{v":LuEp�nR:w����"O��ԉ�U�\�⦤Ktk��0P"O�Ѣ�ʀ��4�[aD;'N�@0"OH�{�h��j~N�/�f�U��*!�dU�fB64{�ڊN��e3�R�/�!򤏌H��I"` y����U"]3^�!�V��س� )�p���E>�!�Dӆ���@�%�
l$\�m��Y�!�D�1gV��S#КX[(&��
�"O6qT�%8�X��&��@���"�"O�K���2|��(�P(��e�� 5"OLƀK.���EI��!�h�#P"O`��6Q0�,�q�W�Z�tAB"O1�@0p��Tj�E@$�z��x��r
���D��/,5��*�cA U�@A��zGa~�NN�c�\�z�-S8Z�F�"�i�=^�)�omX2B≪p��L+UDD8Z(`�r�O?S�t"=٢KE�璉(&*!m�1�8�!+�{	hh�� D�`��7"O�t)�b6
�H���F�1#��i�� F�V!QI�����>E��4��ub�D F�j��Q�I4t����%��c�ʅ7|/fp�Ҍ<�Sv�i�Z����,.ӚP�cK������	:kd���,d�>h��&�)=a|�I�u�I����uE� ���;z@��
�*?v�QyO���D��uS��)d����t�@
]�O�J��G��d�&-HbH;Ñ~*e�N!2آ1�Gc�+4���]�<QĢ�+������װ:���o=�����d�j�z���S�yx��E��'�������[���@A�;���")D��[���:,@�Y�$/2�� �B��MST�(zK���	R�U��Q��8���� 	L[���T�E��BR">lO��������J�) �2 ���;� �9z�pR3+�9�hv�_�#�"����*�rHc��N>Jr�f�m�nc����J�ʨ=�%�śzy(� nh��S0\���d��%��@��O $�C�	>P�\	M�&1_����H�*S����`Q�i��Y���0�t�OA�:	gL�ps��g��t
Ȓ��>C�	7[��Ua��ֱ*(,r�%�._$p�ٴj,R�8�K����ეຓr�I%/I�a4�<j��@qn�A�����!TgV��Mo��;BĈ�?�`���[e}&�:%JϑcČY��'��`B�p5P�hF*� *��Q�#��4�Ō:aj�(ՄD:��'}_��9�.�94�h�jЍӘG�>C�� D�T�P�B��l�EУ�<k�V��d1t$�^�0n:��<��ȹp �EbK�4a�ȴ�$`�<Yw)�Ut�:��;��Q���֘5剪V��`B�����g��n��U�/Y����@��Q�t���	�a4�2u�~�#D�͡6�Y�*�=�� Q�O�PC�;}��s�#ւ�<Z3�� ]��p�_=<Ntc>9�?v�*���#�b��0��4D�� ��{0k\�EH�tB���g\�O�,@6�����O�>�AcL
�z �YI��32\�* ,D���E�0B��[���S�����l&���1'h��IҴ|����X&��8�FZ�%vC���U�r��$��x���Z�8B�I?�.�+�mȪ-���͙B8B�.P`���9(�H���
)��B�ɠ}���1V�|(>Brf��5�B�	�N{&�A�aܩv&*
�N�}q�C䉪t��%�$G�0yN2�"u \v�jC�	Z��R@�#l�J��L_
=��C�	G�����_�k2��"��.�C䉒���Aࠊ8ƥ�fƝSb�C�ɄS��]:���7-�-�D&�7StC�	������ߠV�v�#"�.T5pC�	�MF�ۣc�=NX�1��S�a8hC�u挽�mS�3,�iR'�bz�C�Ʉu�X�#4!�4e匠b�eƨ�VB�ɽQ�B�
r�W4/ڐ�{��()"�C�I	^��U��ቲU�N�ҥ�:��C䉪v��=��k�LQ`�AF��;��C�/$���� A03P$�I�$D���C�	�4vt<��g]6@0C� �4�C�	)V�ڵ|���"�Cy����'�Э{��K���Y��%�9����'~�A����/0�!��C������'=d 	�z��ң׵}��0�'��E���j�^�z�B�+|0����'�U0���`4`���>~Rb�!�';�)G��G���t
�wf6,j�'D����þIBX!�	��t}0�'��)AaL�4�|��(�/f�Ź	�'�.,)bJ{�rdB�C������'��t�BMO&H��@�䉼=k>9��'��`a$"�4�B3�L<+��y��'��Mq5�î1�L����  �n��	�'�����(Rf��w�SM���'�p�J��޲_p�0ǉD56#�=��'�b���
�V�>�[�i�'&�Dtb�'���� �x/�)9���]r]��'����h[?��,�QJ \	���'x�Ѱ��=�$�"p������
�'��݂��E�ZD�%{c�	
2h<�{	�'�9 -;����b�5tʠ��'����Ñ�2x�er�dO�F&d��'��dm	�}�.���f�=�
�'<���$J���3-N�G $���'|�G��2�x���u�	�'`bC��[��d8�,�B�n �
�'m�ɫ�L�z-����
p�"M�
�'x���LxXX��Q�m0 ���'�� S@� c���@�6�X
�'�v���jE�^�#j,]�<m��'.�&bC*
g��x���c�A3�'��J�aC��x`(�(�$mB"�'���)T%5H>������zK$)�	�'B�8�E)�1F�B��#mďh�ɠ�'�@1 ��n����tj�t(��'p��"�Nw��KT��+g��	��'�X�I�)���J$�6Hp;�'f���T��FoA���C�JC�Op�!U���D뺕�6�ًf��%�t�BgQ�΀���#~%�����#D�h��	�i:\%�0j��AP��k=D���n�b�T��tL��1H=D�� v��L�z�������B���;R"O"����P 20���	���[A"O��b#H�:����K�Xk��Q"O��X�.]*7�K�Z���O�<�yR��[��2�[�*��̔1n
C�I�2d�tcE�]mx���Ɖ$�.C�I6:��M:0	D�&@	Tm��	�B��		ؔ�*�K�5i��|�vіJ� C�I�^Kh��E�F��ƸR����b��B�Iq�pX�e�)C����pO�kX�C�I�!��4B�c�:`5p�M�' xB䉏2�RT�d���B�L]C�� bB�I�l? �[�Юj��Lе��s�VB�	�\�%��:\��H��/�C�	1>,)�4L��&e��Q7�2��C䉴=�:����S�"m��f�W!QPC�	�C��R�[5L����B��&�B��!@��[��H�bD�aj���_��B�ɔ&X���?u�����`�B�	�E�h��DC�%u�@�����B�I3v��Ѱ��9�Hxp��&	��B�ɊCN�=jF���9qF�� ��B�->���s#ʅB���O�K�`B�I.PĜ����J�n��j�k��_PB�eB(Q���W�lq"T��3XxC䉶�N�-M&i9H��M g\pC�	�#�L��ª�5?�:��!zt"B�	#3��l;��%����-�gg�C�Ii��P�dK^"�|k�k�3��C�ɴIC83����ztH�đ/f�lB��-4y��@M��0@P8�g�`B�	�=tY"���%B5�m�3�<��B�	78ɊI�R�/|̩�3&�]��B�ɪaN�8a�i�-��e�LǱY�C�I���ţ�b^�8��XS�H��C�I$:(���$B��T�����5BXB�I�&#N�0VN�n&"�GE��^C�ɻE�Zdt�S�W��y��y?&C��%Q�f�S�7Q�ꈩ�!_�W��B䉁<�$��B·s�����_�_��B�I�W��Б�	�3,!A\B�	�+6���ş�_�9`u�I J�B�I."��3@�q��K��ü4R�C�I3x⠭�w��)Q�p�EBB�S��B䉬4,x�)��ڛ_nL+4���C�gVR���"e��<I�蘘^��C䉤O�m"B�6^O�¦lհh��B䉰(� �	f�y�ѡe"�'EQbB�1V�Y%�����P�ȗ�9VpB�ɗ>�1�gƉC�VAk7�J)B�*F�<9�b��<�)���'�PC�.A�J+�R�Rw�`���ƙK>�C�I�}�hmފ)���+��� �~B�(#h�X8���R4* G��=D�B�ɻ��M`R똫2 �)h'���C� j�R%����;1|��RV �)e|�C�;SA��٠�	#9�h�	Ğ��B��PR�5b�i5�$��/B>Hb�B�	:f�е�P�h�@����,xK�B�ɤ&c���eJ	 g&�R�Y�B�I2{,���V�L�8}:=�1(�l�^C�	)l�1�a�6h��8���E���C�	�=N����ϐ*& �i%32C�Ɍ8�f*s���3��q@N��B�)� Z��6
�:=}�+��UR<��"O���B�:Z'v��"��2GL����"O,ݠ��ZP�R���[�J�:�"O���)�)i~�8�k	92Ȃ��`"O2��eR%������:��uv"O^�����z�r�"�+��G2y��"O.��!c�T�VA�I�' 4��g"O�@���Q��
�"'&����"OP��R���0�`Cóbx���"O�����W'6��U�DD�Ah�ra"O*U)F)P�'�p%��LZ�@*zU�2"OLH¬�.fr,�f�,	!̠�"O�8�Q��� ��E�F�T���"Op��$�͙ *>(�&{���)"O�P��гs|��d��|1�ô"O�����D�e����0��%)�a"O�i����(N�t]�7�]�q��m� "Ot�)�K�D{,�7�	xhtɒ"O�� !��C��2�B��&@<yГ"O��� �DJ�zbP�A#h!�"O�yiwEN�C�Pq[��(:��M��"O� �G�?��t��!��D}�6"O�,y�J�o	�y1aM���4z�"O^)%C8E��U�am�q��i��"OP��'����8	tB�!"O��ؠo٩Dy�́�?c��Z�"O�0x�od���X���(�
�;A!�D��>��1���\H��[�!�Dz	�vNB;U"�Ѡc)[�9�!�$�d�����v4=�u���D�!򄚄`|m� 3m�Z]�Wg�2j!�d���;!��'vbH�*'H/Xa!��F�/v�AB�x��(9w���H,!�Ě(L}Q #��uB�n��	!�DA##1�
b��B�:f�G!�$��gɠ��"+�b58���7�!���<J}b`��eҺ���)p�݇ȓ�0� �V�E�~ +ע�	�bɇ�`�*P!ϒ�5�tP�*NT�D������	�&|f�PTEA�q���hˮaO&]��=�vj�QGT�ȓu^��#�b� W �J��<cרM��V�c$���'�QZ4�	�}��_Đy��	p���r6�S�~�����s)jMzqCF�~�x�!*A$#�%�����lZ�w?ISN�&�RM��C���v���=�	�d�>i��E��5�`]��l:y:�����o�H��/�f8� ϓl�:��F�]}��`�ȓ
o��3B��uIF�@<yC���ȓ,d���Q	.r	�4!�l]�8Rą�M�ǁEGU�wO�)�L�;�X�<qEȔ>L�I�T�Az��2)WW�<�"����]Sr�Z'�f$!#Ej�<9� Y�W�H���Q�S���d	j�<A��<IْI:@�'*uB4��j�<�)�3'�9[��&����ׯ�b�<����mr�C�Q,x^p�����J�<y�抏!�!�b�+jDԙ�B@}�<��EU�NJj6(�&a�v}	��d�<q4�� ��YW)�ks��B�l_�<10�9V/��8'O�W
n�T�_�<q�I�j:8�I�OK�U*�`�5��[�<iW��7��!��%�}A�$X�<� $�Q	A.n�XDr�m��a"O�])�ś�hJ2��� "Db�	A"OtZ5l͛^�9�o֠c��X��"O6�Ї�IK�(@���C#��p"O
;��;<�B
VBh����"O���
�;^�b J*'e���"Oʔ�b��30�v	��d��RH|��F"O�%˶�ӏ a��'Rhy5"O���5@Lp��PG���Z�!���J�h!��ۻp�aQ�K�'r!�\��ra�B�4A���)�;!a!��Q�~ ���w�]��y)��D!�	�i���z�C��s���	�\:%;!�߮D��y�M�A�BXu����$��4��s�Ɵ�7l�d���yRŒ$F�� ��*P͠@�y���NM:xRbdө'eB����6�yr��	7�p+D(�:�ڸ��(���y���*#49B�K�2�5J��ӏ�y�)عV��"&`�HڦI�y��\_���5���.��6�״�y"$�=
�%8 %|8"��Kʤ�y�"� l�|	�.ݴy9x)X�%���yBۿV޵�`��n�b�K��y�B�M�hi��M� 7פ�O���y��0m�jy3��Ų)A �h�L��y��Л5�X��&
�4d�� ��y�Âg�بS��������"䃺�y���C!&�aP�LH*Lx�Ѡ�'�yb�=D�	���ʜR. �{-��y���px��Z�%�Q��X�5��"�y��1u�1W��4���10O�	�y�䟚mE�ܛ'*'2�^l �fU�y�G��yY��*�F� �t�H��J�y���1��1���*:�Q쀰�y�f��¤*�+V��(�s��<�yR�G#Oʮt�p��y��)Ӣį�yBh�-1(����<�d�Y���y�!J|�A�m�2��ʄ��yJVx@� ���*��Y5�	 �y�K����q�/�d]�d�8�y�&�*j
2� qN��s�Ԥ�y@^6mW~���ㆆw��@�d�yb��w���2
�r-K���y�� l��P`�'G3q�����ǎ2�yrJF;j��];@�kkʅ�`�1�y��V�U �Ģq�|��p�<�y"B��/`�3�EЀj�V@աV��y(D�{z�|�QK߀]�vͺ����y� 
�0�E�L�8r!��=�y^H^p����� $v � �T*�y�L=��RE��v�����yr(�&�=�7�KkL8Ѵ%^��y��
��H���K�av�ڄ�Ӈ�yB@F!K��%�L�U�S#�y�"�B���a H�j$0�*
��y�mP�|��ѳ H#98��CG�S��y2�!�
���@�+�\�&��+�yr�&,6(aګr�+v"��y��C���Kd�����yBӢ@Px��!_-�X�+�`^��y�#��E��-p���\ԄX�!�y�&A6~2t�&���ǭ�+�y��Y"E�4�J�	�	&��k�Y��y
� ��9��%N@��%H��P�su"O�$�p!X�
d+��x��"OL���/�43B(Rp�εL��)�q"O�b�%�PfZ� ��I&_���j�"O�yɂCԳT`b�sb����V"O^AT
V)�6�� Y�c��!��"O8�@�d�)�ޙ�ǠW�wz|J"O8@�3BۛsYj�뗏�kJ� 8�"Opq�2&T�r� �v�8q,�	p "OT�3�J�.�|-��lY�K��;6"O�j䆬a+(�CG��8��%ӆ"O8���ZD`򧈆�c��:`"O��@B� R�s�G����t"Ox@b��զ�Ȥa�l؋6)�E�U"O�'b�?�<(�b���k(B$K�"O(	(��ήMX��D%�-W!��YW"O�����	��!�!%�M� ��"O���ZL�F�ꑡ,u��Сp"O�Z6+��&d�4�`.�r��A�"O(P�Oma �g�.g�:P"O\��sf[�A�����Ton:Cu"O���qB�,(\2�2a�Q��a�"Ovd���X���yhf�S��"��S"O�ͫ�o�{��P��@^�@ىu"ORi�ӭI�0�-@r`�/-�Bq�7"O^ � 
6%I.�i��"&����"O�3�F�=a�B��H�T�>4��"Ox�9���rU4���Ș�Bo�	�#"O��6��m�]�%NO8lO���"Oh�zA��95��s�oںh5&��"O"�����g�� iq͕�lr��"Oy��J�m���6��.��y�"OX HA!�-@"6�:v�1tA�X5"OȌ���ԋ}�Np��/�x� c3"O��M2I	��H���H�1"O~�cQB׸@�!j�.�g>�zG"O� �ĕS����!���T�*d"O�%�A�??�����KZ����x"Oz}z��C�HQ8�R�KO�e�
�B"OFP�`�"z�`A���4��8�"O�i����=wBvH���^��$y�"O�i BA�$�4L2b䋪Swޜ#"O�L	e$F�}c����� �@�h(��"O�Y��*f�� 2R�7I���a"O<l`��?&������H�M�
8��"OJ|`W�)&Mrl�P���"O QHT�\�k���@c+�����y�"O��B��wʤ�q䇴�zh�S"O��QPj�~1"u���:�c�"O>LY��(a�l�����?���R�"O�PHp��>m?�ì �~z�4p"O�1����k�"-A�Adi��@�"O�a�(D* a � /gZtAC"O�]�q�^��i��]@<<��"O�@�6Þ�4f��#�*/
��U"O�`5�]�LfYȔ$^�qv�Y'"O�)�R!o�*��l6�=�"OfE�v���e�n`(�,)l��"O��)�/4)1L;c��j����"Ov�b�!��;>Z���W�vh�IP"OZ���՝w�p#e�&d��Ї"O�̀&J\~�#�';_wH1+�"O��B��
� �@p�����N� �@q"OԝyvD������� �;"O� �d���˾y�6$� ���Y���9�"O���E���e�V�4v҄�"O�,���H1aa ���I�BIB�(�"O:����V�d�(RO�����"O���BI[�R�B�I`Ϛ�*]H�:�"O����H5l�R损2U�� "Or����1ۊ�af�\�>*�� �"O�\;"��Nq=p4(H�Q!��0DB��4�fd���`@�^ !��A1��5��ǁO���� ��_�!��I (�~-�p���(�|4���M�!�$��c08!��[13mf)C�/Y�(�!��z ֬r��ͭi:;`K5S�!�D6I����J�"���:ro� �!�D\�h���  �x6\3��K�!�DQ�P��|��Ŏ-msr�Wd�
 &!�(*?�|�����*�,�[�Ԯ.!�K�v��M�'O4H��mS�Q�d�!�Ód�0��"��+J�E���C�K�!�D�sw���5��=��S�H���!�dA V0�#�G��0�$�t(�y�!�D�.3�-u�ָ;��-�'�T�!��6N��ё��b�
HHwT�u�!�D�;~I��C�d�6
�@(36  �+!��^�t��(ył͋�ĤPb�ӂN !���D�4����
�u�^����g!��ǭVL��1���7�(�4�Z:�!�Y=n�蒯�4Br��pb���!��MT�	�!��A(h�z��^�u�!��!Ia�Xs������9�B�� {!�d�jk椡de��M��  	U)
!��,,X�r��ŰE�0����_0?d!�$��~�P�hV��P����Ťc�!��]�xS�D1*=HB��d�!�$@3RW��3G�3o�D;��W.!��ıB�`�FZ��� �fʐ:�!���W�f�p1�K�_J$�+ �P�J!�䞯Y�(LҠ`�����$�ǽe�!�$�&*ǀra@�cn\��Q�X'g�!�D"J`���㥟3O���4hˮ5�!��W�h�W�����`+�!�8s��Iu�#0���Qa��C%!��
(3tF5�q���'��X�͔9!�DA�8��C�N.�@�Z���K!�)N�ZH�3/��9���>#�!��y��b��3X�4ٱ�L�%�!��|Ԁ�pgŦ;��� �H-�!�۷M<"�A0`@�"��� ��Py#�s�YT�Q�9�氡�
���y�F�o���b�?5�e.\<�y�fU�[h�i�k:~����%�y��ǅY.�1��>D�yj!,.�y2�-u>��%ߖSd^p��`Ŝ�yR�0�F])��ֵ��m:�m�"�y�G��hט�yv��H�x	G�L�y�&�Z1�q0�HO�-NZ�s����y+J���q򫆗"X�9��A��y2h+q�tid��=HUy#�c߽�y"�\<)�zs'�3�ċ6I �y"M8�xi�+A=+�N�(����y�l��N�2�ɆÆvā��D�yb�o��s���l����yl�=uL	rR�_���@����y�KK5-&�WY��y+�B ��y
� �4jc� �0���a�o��f`p(��"O>x`흒5_T	�'��fI�U"O���V���"�z)��̇a�9�"O2���C�"7µۅ㓗��Hi�"O�q����>&�����>%�����"O���t�վJ�T9�-��_���R"OT�`��VmA���bP�K�"On���ݯ1�άh& R�+���"O�K�҆a�.U�P!CT).a�G"O&�B��"��ٸ�i*�&���"O����E��a�p��#��(ό1c�"Ojy����&(��!(��_�<H�v"O��V�ҿ"P�Z�$C��"O��d]u>8��4\�.b|��F"OD�(��ʄ��+6f54RD��4"O1��Ğ�iW�M0��љ5FҠjA"Ot��6GM�:F�@�o��"O�u���!
�`�EE�*}��"O $XDH�\�T�aЄK�UF��"O��j���P���3�〼5�\�+�"Op�I�Cb)"�$�*t6"O*́����R�DQ�&+J�<l�"O�R���#e��q�Qr�eC"O�����$V�b܂S
O�D1D"O���ɚ+l��#�'0krzݡ�"O
�26�A�YÆ$�TC2#kb��"O�@T�
?+y>9Cu�I�`M�ljT"OHD�0 ץtO��S%Q`r!"O�0��C��`'T��ǥX�Ls�!3"O����ǶV��c'��ic�9��"Oly�0M�:8ƔF�KAlC�"O� ��M��Z�ذ�7m^Z<.�p"O���䎜�*֤����W��i�"ON<H�C��gxp��V	a'����"O�-�d2@ļ0�ē.���	�'��%��E(.0�2pZ�d	�'�P�D$��؛2�V!t�  �'��������/0<@ӑ�?rX���
�'?fH6H��Ԫ��etz�P
�' v�u���:�py��_�`+����'Y���ȝLd ��Ο Y�2�'� d�!̐�`b$
5��"p-�P��'bX-��y�~���灂f[�=i�'��Q�'D*{�h1Q��*$���',QI��*~z��y aֿ��$�
�'���l
���@'@AT0�KXg�<���#H��05K�Pt���4�}�<���
�u��j��5`)ҴC�I�C�<᢫D8`0L���-R����Q7K�@�<q0��n����� B+1^pA�pg��<yt�ɐb�x��⇨'��uD�S�<��l�����4O�>{��5{G�D�<T`���t,��$M9r�Z��!�ZK�<i6�J	<_���rE�5q�j�4G�L�<��2~4Й�
�g�"-���F�<!���~h��32KR��q�&�B�<�gV-��h��җ9�Ua�Bs�<�'��/�ܻӥ�}������C�<AЂ��o5�IC���,=mʍ�FGJ�<���gv�U�ŏѤp�B�Q��Q�<��C�:{�v���ˢaGF	�#�N�<i��?��$�% X���l�E�<�Ʉ#z-ά;�ǥ2z`�7.m�<1gH�I&>(�� �_9lܪ�jDg�<� �8�e�ȳ8���Ӄ�.+���g"O��Yӂ��_�:1��@4��"O��s���'{�+��է.�&l�1"O6�1Ą�P-��fI�D���#�"O���U�בh|:xK�]kX�Q��<+��X,%ٛ&�'f�TT?1b�$MR�	�՘w%�����H~H���?q���yҢI-r7���[uKDiR�	r>-��

�;x�@�lW�yŀ��u+ғZ7�df��5Ҹ�ӕI'Q��\�"�`7�`0�#ݦ"��L�g�"��#���GQ2㞘S��O�mڕ�M����Ɇ�F�rd�H�'�Ma�ʊ	r@l���k�S��?Q���DD��@veܿ(ra�`#RH��l�I#�M3g�iΛ��0)HV����N0v �&C�~�		�un����'�RR>mxCk��|��ߦa{�럈j��0��E4l���:Wc6_�&�u,K�HP��-A�A[���F-�?m�O������43t��5�j3�Å��l	�i�VTa �P��h�OS֙Qe(�2m�匊W��Ƥ�yAT2ȴ�BL: ����in"�R��MB�Ư`�R��/��i�B��I��pt��2$<r�b����	{X��(V��)C�qׯ�-J��y��0�h����~��Ob��x�	��lN�`��`C���S���p0����?���$e���?����?A��T���玲㭉n�+ԩ>�Z �q�P��X���BB:��S������nD�"<�E�J�a�h�yrd�>pA���̀�q�v�9eK�C�QJ'�����h�Or �P!�ҡ0��̕'6(չ��X8���DJ7&�H�e�O������OX}o0-���<q���d�~:6�kt
6/]\�����[!��:�P4�$��>�摹$�M?L��޴G��Ƒ|�O�tV��З��9����j_ 1��	�Ɲ�H�m�V��ߟ��̟���u2���ҟL�ɸ5-9P'��m��	��.#���АbD*]I `R2�UnLxC�lG�:G���c���&�h`��S�J���S���Y	��"Q�L����o�%u��떠�5�H��D��}�r�iC��SP#F�Or�KE�@��6��	��T�hHd�Ӻ�O�^}9�.ͳB+ʕ��I�NV@��'�(x1!*?� �����,{A��)�'�&7-���'��\J�is�j�d�O����)�C�T�(Rp�)�ّʮi��X�;���'��mӎ4�@u"��;pl��i��=�p��'U>�@��R 0�ه.��&XEz��00sF�X���1�"$J$È�uan$�[w�ܬ[d$^Ni��B��_�b��{�� q6qO�/t�$�O��&>Ul��6��P�-��`��u�F ��(ox�h������9���;���I��0`��M`�F�k����d�ަ��ݴ�M�C��(�P�����]f�ܩ���N?�GE��*W�v�'P>�3c�ڟ(��֦�`L-Z*:�ۑ��dQ�"p䐩	����%��UC=0)�Iۓ��?�O�$��0\`$c?x�b��t	5���S�iߊ�pDɑ7-�Ɓ�e��d������I�\}{R�~���RA7�;C H@�&\�|o| xR�i�����}��dw���)���%�;
�ޕqqċ�Ug�@�B����	ş�àT�'("��s�֕��-әx�4$s͗8tQ��R���M{K>i���bu� )i2�Q� ,	��;���t�`؞l[S�   �   r   Ĵ���	��Z�Rt���/ʜ�cd�<��k٥���qe�H�4��S66<q���\S�f�ث.�"� ��p3��yT��7%�7�T�E)�4Om��;��[yr�O�X��j1L�1dd&�x���+[�� ����,L�=/2}"6͍�N��$Q�샭Ub���

�z��I�xY�&Ԕ���(_�>PHP�N$Ap剁;��	)�d�%��f�	Z��1ɕ[؛&E�!�\Q��*m�yK0B�?�C�'���U�%I���� EHY����Đ7bxY��'����� ;:�8K�b�����Q ��2BaE!�ug[1��4�3̂�G�	�[% ���<J�b̊���<m.�fl�]��'��f���O�I@S����ny��� ��T��K� Pe��J%�����'�pYEx�Iз*�4���K�t\��{B�
�Tf�#<Y�*3Uk��^<����O�j���h���oӀ��O��A��D�Ÿ'3����2�I�@ph� �޴�N"<)�`,�f��!�K�#��Eva�
�Ƀ�h����>	g�%�3���{r5�� �4�2tb�,��On��'C��Ex�o�e��i:~�W"��[��b%�N��D`�(�w,�#<y�n�OR��S搿BE� �o�/:ty�"�ï�Op J<�4ϴ5�~��a�0j{�!�GD?��8�J{�OD	[7�'CX���'Y=�8�ٖ�EI�MQ�4s��X�'��P�h�OxM+GZ���K?�ǻ�H�� �8�j��$ʌ%k��:Ӌ$�I�Nr��I!�>yqeD�$��Q15�\�R���fi�G}�JV�'K^�Fx��N�$��4�vlI����C�5�y�'J/D d  �T3�p+s"ON�����O�8e� B�0 V"O�%R∛7I$XE�'cD"%�mS$"O��%f�Ud"=��]��{�"Oh��b�7xK�k�*?�<�"�"O� &�� �A�Ġ��/ժQ��p"O�LZuk��5^V`�&O��t��MҰ"O~���S����@�\�u��Ṥ"O�ٺ'hί|U����kɻN0�"O��X%�N�&{�(���Ƅm�t�+�"O���D,�? �$��V�Д=� |Q�"O��6� �&����R0u�#7"O.|�L���1C��F����"O2����#f� lʶ#����"O�q%=�q u#_����7"Ox��dG���ԛ`BA2z�d�9V*O�`�ň8W4���(>A��Y�'nrX�f;Z����Ç_�Ġ�8�'<�=���/H�ؑ��R2���'/�A���;>�m��BI�~�N(
�'���W+;cQ�����pv�a�	�'�6ܱW�)Q��DT�J�8
B���'9Y'͔�Y��dIv�%!��;�',6%�'� Lb��R��o[���'�P�1�B?<����M�t�\-��']�	�8�3���z\�*�'�D�1T��y8��!�Le�����'���;ԢO�Y��x���$���'�(�l� l��Y/6��a�'a���E!C��Hɹ�B�&(����'8�5� %�i�Е��"��L霑��'��q���$v����dۥ<t�� �'��XQ���4m<����$e�:�'~u��/܊#����ZD��'�Z�S�L����cէ�'�v,��'K��������15怖/�i��'�B��5���c�����K,l�`�'���Ѫ�.UG�[�j��~��k�'h\h8��G`�X�"�K�q����'��}"�ߢlx�$��ě�k~�(�'l-є�L$F�d����f��y	�'���IԌJnu�(iQ�ZY�4az�'^d�I��tk�P�%e��b�ij	�'1V�sNF l�xAvū,�H=y�'�4L�]Xp���T_V���2C���y���e��ݢ�XP����	���y���S�RA��JB.E�lI�����yBj�=_At��E�D;�u�L��y�J#dq4�@��Չ0�ݨ��ϑ�y��av�9�%�":0����
7�y��S��ı�)N��L��ƃ��ydQ� �,%��$S,��f[�х�3�&��A�W8wR�)���e�
Ѕ�!�v���3a�(�)�H(�ҭ���`�⤃�,j�`�e� 
�ୄ�?�x���6N-�	X��_�D׊0��Vtݒ�A]3>W�Q�P'֞Kp�q��`>���vo�
_Z��@ �F���@#�����G�D)����ȓZ��(��l·M�zeg�D0"���y��4�U��	V0���R�� =�����{BI�K֭?Q�M���鼙��1j�����w���񦆗T�H��6&0B�c^hJ51cΏz��H�ȓYv](��3w��!�'�;$��b�4��T���\V�%a䂭m}ę��4L�;B~�$10#�=Cڅ�ȓ �b�Y���4�Lв��
0��ȓ2ņ��qg
e��I(&�
3@�̄�S�? ���c�0X9`�a���T$� �"OP�K��
�L�$��K�8	��cp"OX���F3|'r<a���1,����"O*���b�'�fx�)����C"O&��L?/���2T�ή!>0��"OJ��O�6��x��a��Z\��"OܽR��%V�����B݈?�h��"O��k� چju���'
.,��"O�d�c�
tx���T7R&�M��"O��e$Wo�l��jݕ5����"O��h�/Q.8���'��Lx�iS"Oȕ�JM�~8����?"���"O��PG��A`'� �˲(k�"O� ��� k|�qI�S`�"R"O��d"��^��ͩ��7K>�0�"O�L	cۍ,�������l6� �"O�lҰ�'8|ٙ$e�9]5 �:�"O"t��f6l�q� �N�h�"O80@���e��ؼR	ȉ!�"O@8 �_lhx*�l��}��(��"O�eS�͙_60ѤS�w7Q�"O� R�A�h��:�C�b6���B"O�8!�j}����C66�T�[B"On��@�[o,�2����8p�"O�y)bJ�����э�57y�Չ�"OP�(��7Q�nuk �ݡ�&T �"O���pM��;t�S��х?����"OƝ�7��2�H���,�h@���?|Oft����,5�X�x�J˅̸���"O���3A��R��"���.a��z�"O�1�&D����C�ӵ)2X|1u"O�mh�I�.uoH(CH�	$Xt�"ON	��L��]�pHqt�M�T�UQ"O��+ ��,DFXX4 ��	��ݪ�"ONx��L	r�Z�/֪gJx�p"Oa���\�1*� ycDCQj����"O(��eI%��-����Z��X"O�8k����&���E�"�U�s"O�sF&�x�bA����u��%��"OD�X��0\�� �!�T�6�S"O`d۵�6I�$���A[;�ԩ�&"O�\R�i�w(@�� -It�m��"O�����v�H|JQ�I&ld%�R"O����n]���[���*�:�1P"O24@�H��2�T��h^��i�"O �zG�\Xh�r��=8�n�:&"O�y�#� +Z}[ul��6�u"O�1z�bW�X4�r��-���"O�u��
)Τ����4�.�"�"O$�22 �+Wx��	�1v�R)�"O^W�=bИ7��=J�F<kv)�\�<A�",NR��n_�����Z�<AR/N*R髢�k�|���T�<�!ިlI���Qf�9����P�<!�*�ҍ2A��P{h(��E�<IfXfˢ��Ofl�	�#�X�<3�s��|�uJ� RB(؃KQ�<��N�kw��@Ί	d��!�UP�<ٕ�D6k��8g�H�VÒ��F�<��#կ(*�1k����)� �[v�M�<�RA-�T�A$�//97j�}�<q4H��zJ�a�����@)�@�<����1}��ك�
ƭC�6�2���x�<qGJJ>m�Z�H�+����q�<� !,]7@j��"���x��"O~�S�HR?͐ur���rF���"OT02d�D�*JL�Qϕ�%"�Q"O�� 
�A�>���7����"O���F�:& �%��f�=��x3E"O�Pd�����Ӣ��#_q�Hj�"O��{��Q�@Қ����9KƄ��"O쌣�7bH����.�#m�A�r"O�}�D�)X,�����
'0����G"O�� P
Я5��X�J�lq���"O��yL�A;*�3p�4lM�c"O.ؚ#m�Es�TɦEӱ5S�1x�"O�� ��_��X8kt%��>�, �"O4��6��^�<�#1_�A���(�"O*�I�oJ&.|�YS4���@f"O���V��j� � s�(x"�ۤ"O^̩�hY�8���'��m:��"O���ČֆK��5�M�&b$k�"O��2G$�$YI�ʁ�,y�QF"O���"iR/��10��	]oh*S"O�ظ�
���H�2Z��Сu"O��� �O���ܻVdطW� ���"Ot)��"Cqu����nq��b"OfU��&�,
���u�7Rb�r�"Ol���Ȉ8�`Be����`�"O���aJ4t`5�#�	\�`	r�"O���kķ������̑^�6���"O:-���]!IW��8��L�^��"OV0
��?M"�	g��W��$A�"O �ʖn]�L�|���J��.qf;�"O:�I`kH;[l@i1�޶@^�p3�"O��R��F�f�P�d��:Ct��"O$�c��½xn��k���g)�X��"OXԘ���*�@�����r��0Q"O��`T�WnjU8T�X "hqr"Oȡ�@�ֹp���ےE@9�.��"O0��4J�;jY(ȳ��A���s"O4�b�ǔ)~a�11)D�U��a[�"O�%�@��Zh(��w��/N���w"O:iG�148��ӭZ�i����"O���q�� vMD;7C�	3NQ�"O�XKD��W
J��@�B7L���p"O��	T	[��	K�D�Mshd�w"Oh��C�#yJ�5ٗ�L�npܼ�E"O��'k�;(�̄�O��dA8}�"O��)kƢ.��!P�_ ;�T`�"OƩ1'��>c������d+!�Nk}�}��f���N���ݽ!�!�?��qo�@�>E���!,{!�d�1X2PL;��L���! �kδiP!�DС,�!�#g��7΄=�țp�!�dV0 �L�T
�Q� aF�O�a�!����z�����L�\�hS�9	�!�$�`�n-�trO�J ��Mx!��=r�:�j��UH�l�+Y4vr!�]�[�r�ޕw�Nѫ!Dԧ1^!�$N*W�bL��=|s��뇂�[S!��1��|��G+l�&AS���G!��p�hf�>*��D�Do\5F!�$�<LQ��*�>)����6���=�!�C�:���" ̑	#�\9�l��C�!�5^t��lX�N���J|!�D�~��Q�V&f�@P9�&�?�!�D��*k�
K�B$�4��E�0�m��S�? j)A1ۢM�(�93J)2D�Q�"O��8�J-�L��3&�(P#jx��"Ox*ŏ�k�tŨceGPz��"OB��E�DD���cC�R��P�"OV������/��\ �aP�0H�|
�"ObDp#f�3,^��CR 2��s�"O�� pʅE=�hC�(���`�G"O-���uL��9���QÌ��"O�)aW \�wΆx�D��<��P3t"O�H�6���RC\�����"OF�� �E}B8�B��7
z(A5"O�)�P��
oT^��Ĭ�H�"O�Aˣ+��^��@���
�سw"O�V�+o�Xci	���5xu(�K�<!wb, ,�![�o҂h�,ɣ���D�<���>I�����N�pR&�����<q�
���� ��6]�DQ��n{�<!��>������ꦝ�U��m�<����,6�*������<��l	`�<�a
�sf�}�g�H�pݲ����U�<�����0/4������o��S��G�<q5�I6��E�נ#d�)�7l�E�<�Ddڼ�8Bd
 YP��+�$�G�<���
.b�K��әO����!b�D�<	�N�I�s�*P�e�
u'�C�<�B�1y��U;��'Ѕ���}�<q��PIj����V�&C~m��Ha�<QѪ	����z�O�!q����CZ�<���+.���CƋàs��reB�^�<1�����q���, =H��M_�<a��#sN����pl�4��Ie�<�F`̱S��dΙ�z�(@dHBb�<��&S ��Ɇ��1.��pF_�<��r��x�7��a)���Z�<���
ay��P��,������j�<ɵŚ�E��!��qJ�:!l�j�<!")O�U���p�e�I��"��j�<a����� FOD��ǁ�c�<ɳe�)<��I	f��=�htJFe`�<Yf��5o���)4d͹[}*\�C��Z�<Q֢T�1�b H�o��=���3b�N�<�sD��j�85$C�H'��x��I�<Y��T��朹w��F{5s�NH�<�g��HH�m��ȡQ�`�ԢL�<��,��O�6�Ho[����H�`�<C؟n��h+d���$��i�\�<qQ�/wY�d�v˙4�W)N�<��P'B��X���ʘK�8��@�d�<1�gW G �
��ϕr�v����a�<����$b� �Į�T-ΥQ�FB_�<y�HN�2��0�#�65z5�u�[�<��K(��"D�˺�a�Y�<o�T�,�7,A,upY�
Y�<��ȟ-C�Biާs� Q��Q�<a&�-���7�#%��� XK�<!�,��-4�)���6��q(s�E�<�gQ>L[����a�9c]@��D�<)���I�0aFË7Zsn��ရX�<�R�q�:d��K�4{\d�t�DS�<�B�H����u�2L؍c��\M�<a�k���ʙ�ȣ���!1�_�<ɠo���0�Lx��qi�k�[�<y��Qm:d�� _�=܌�C�DT�<� 
�D~�d힦�	'��L�<� ���u�;h���	ޘq>B�!�"O���ďkN�I��M�Fנ�r"O�����X��Bg,B:8�Ȱؒ"O=@-�%mwN�� ΜF�\a�"O0=��H�vkx	x�`�tTf��`"O|ɺa�ׇ_��!���C9Ψ�"Oj$���M�/,`����1��JS"ODx���>x4���[���1"O,�!��!%���B4	�m���'HPɓ��_Kh. ��z����'��}�(B� D(��ƫJ�ADl�'Z��{������ɲzqD|!�'�^��0Aܒ��}W��oH�(�'+�����+�>Q��fZHA	�'
�����;/���6�ҴY{�i��'B$+$Kթ(t�9�Ea^}��8�	�'���џ@��}��΂�B8k	�'�����ׯ\����Ӛ}1�d�M>��O��a��\���.�:@��ȓ�>�k�c��jrܭ�2��YP��ȓ92|p�'��6p�<P���/$�܅ȓ��#  ��j	pU��*k[�̅ȓD/dlч�Ƿia�+�)j�х�U���C�M�Ly>P�B�O�\V��vlv�C6mK=l(8��-���Ʀ �GHH�$�3�a�"�"X��>�* h1�E��}�}�ZA��P@���A��c�V���C�a����=�����Tm�u2�����$b4@����y"j�/����&JF� �*�Pc���yeݭ-hd,B���(�Α��y��דa��Ê�S�L|����yR�W��n`A��7Z��jw��x��xӺ��׏-?q�Q�f�A� m�"Oܑ�U�C�d�*\ڐ$W�9@�8��'đ���@I$S7B�J��ŕ[i0i@�7D����@�/���b���� L4?��)�'X������+F�J0�l�s\���ȓ
tй�C��z]�m�MWJ�4�ȓt%n A��mb$�χ�"���:ъi9�'��Mf�G�
���ȓt	0��ACڰ�X̢Cʇ?M�$��<Q����(�<Ek܌��f �c>��ȓ/A��2���nXh�(���i�V�ȓ4�20�H�O.��(�j�/�q�ȓ`2�@2�-`�MhQ�P�m!�T�ȓ	A`<T/�5,��<���Ǡ31��ȓxfIE���p��B	� Y�0����Z�Jw)��T���PG2d���I�}�����.0s��Q.V.T`��<M\��B/^;Ԙq��e^&	%�ȓr�\��)Y�x=���� W�J��ȓ_� 1�nB ebyx�I�+s�m�ȓ�́ ��m@x�SuEJ
*Ϛ�
�'1����e�e�mڵH�4�]��'$T各N1Y(L �/� �8Z�'�fx��8��lD5.�P�'���
�-��N��{s�܋3_�;�'W�ݡP�S�adH�*��\�,�\B�'$<���FW6و�ӬW��p�k�'�ĉB0�J��r�����x�'��9���9o��]$�:cT<p�'�@����D1j����ׁ3����
�'�а%d�,xn������#n>}�
��� |���".��ԥ��D>:��S"O��IF-	�[�䈁�˞k,0d��"O(Ѡ΋(*D(��]�F�$�"O0\�tl�R���R���ar�"O��%�-CGv�a��RI��"O�p�&�'�<#R[�!��,�&"O��xga�fN�����o :4�&"O��q�"]�dd�ٚ�lL]���B"O��0`�ǹ{�\X�F��d��[�"O��Љ��7@d�B��,��x2 "Od5;B�y��}��ͩR��
"OxesQ�Ǖcj�Ыd� Md��!"O�@��(�*^��Ĉ�����trT"O�aD)���b�ڥ�(x��S"O�ȑ,�?g���!Ï7ZtIPU"OR�
6N��c0�#:<򭱲"O�y�bǗY��Uڅ�~-I`"OP�7��h����ˆ�6�ey�"Ox��� 7M�i�H���)�@"O>d��#u20�cD��/�$)i�"O^�J�bW�#�]�aՏ����"O����j�t��P  �}Ң��""O>�C�� aB-�$i�2D"�#'"O�Cl��$��i9 c͎���"O0Ѥ*��1�쐣���3\J K�"Od,�0�N�"�����OӶ%8�r"O�����756`+��6=Pq"O�q)��؝U�Ѐ۔O�3�b��$"O`ui���6���U���-�<e�t"O5jң۪f��c���8hֱ"Oh��&K�"��)�UN4���3"O���mM�
+@PA`�<i@�s"O���ȓOH���΁$>H���"O¬s�Z2Xy�͋��Q�� ��$"O\�r�
M�4��
Y{�ʀ1�"Ox���EȤgܖd3@ǈx����"O
�ha��Y���
[h��W"O8��'�A���X���w>^,SB"O~�)��˸F}>Lð@E�E8��Y3"O���B��^�x1�oV/hR�e��"O��B�(��j��Pbf�Z�v"O�i���:"u��*��_11�$4��"O���G�-d�p��d'̄�!P"O��ۃ��r`y�4MӰIf�ap"O�ҁJ'e�J�[�L82
ҷ�'`�`P.ZgB�@�Y8%�X`˷M��h�'1�����O���O���O>���O�5t���l�t�S�����P�F�� 9 &��䥀=F��;ËE<]�����y0Q���&V�D�:"L�%Jtp�ϋih JU��)��x���=�v�	�AK;m��Mc��@{�ɻm����J�[c-@�.=��ݜe�%������M�����D�%B����|⡁�	EX���-�N2���@G~�'cay��̣F�xT˗���b��h�q_�"���Żs��]n���`��4��`�q������O��w�D�ӂ��.]�Q��Ċ���K�)Q�����O���N�(=c�.O	<*Q�����#�t��ѳf�()����[�dZ$I�?��LQ剧!������5>��sw/�?���:鞈:���`�D�4:5x$�M����&��&��i�O�nZ��M�����ɍ,D��y[�A/K�t�X�E��MZ�hB�4��'�"}��=TĞ)#�H8�a�R-��A���T����ڴ�M���߇6��h8�e�Z�uX���O?�7�9$���'*T>�(Q��ğL�IƦ�ҩ�=D���q�ޜr�^C�� !�eJǪ�&B�� n��#��S!o�=~�4��)�R�ih��*tM�ՐT0�J�?�F�p��a������g����ᗸ#��F�.R��:��D7Z���5�#**Z����"a)ԑ�$h��MSUEKݟY�4�J�ğtF�ܴm�zсf�_6.�J�#���Y��?�)O����\�M3A��9�Ec�:8 q���dl��lu�l�T��cH �iW-_�N�����)-�.��O���O���D�O����OT٭��?�޴}��!Ї�� �� r���+\<Ր�OG�D��Hͳ�ʸ��%]�}����	�(��jJ>� R�j�@	>��!�%�T�^�����"(u	\59�HV7T�2�ە�U�"N�
q�R�uO2V����>��9#�o�Z�j���-�(@->�'���
��?�R�xR�'��T�ܻS��J*9��P�h���Ӧ废|�I͟h'��}"q��,r@����C�R�|�1�l.�7M��)'����?�'H�$9�� �N��Ԓ��@h��aG�͝l�P��'<�'��EߟN��'PR�Z,*1�7MF��8Ek`ʞ��@��,gnh�ui]�4jD��,�1�m���d�"��yS<%�@`��Zn$��`Fy8<h3a	�a:xȅJ[����c`p�O�����'8t@���ς2�X�V�_��0�p���l�6-�O���?	���?y��d恩qJ�{�#kb�ز�e�3�y��G'Zl\Iƃ�afȬ��ɞ��~�U85�6��<!�	Y����Iȟ��O�� 9���b����A��#;h��/��Y����O�����@���i�H�Y���E�A�#O�rԯ�(H|D�B@תhjr�bB�"g�+a�I%)I�ԃ��ۢR�rQ"! �;rDI�'�|y��*_���?X��@�$UX(��*;�$F�$l2D{�Z�l���O���O Q��!�/zT�K�¦��?q���O��I����u0��#ƃ$�y���'�46M���mZ�x���(���Gxz�rƊT��<�N>�}2��v <  �   d   Ĵ���	��Z�tI�/ʜ�cd�<��k٥���qe�H�4M��\70<����z@�v*ɾE P4%�M�R]M�Q� �6��Ϧy۴8��$ �Ibybl� \�!����V��XS%�,8@ɲ0�PK9�=a�#?t�7M�dn8,��W*¹
�c�.2���&�ʠ�"��RG�I�Us �j3͔;���<2Jڽ��%W� 9�P&�92���Ej�6*;�v�tTx��/0�H5�V%�?)�'�������%g� $�r���9F�(�fbSA}��{��c˧~f���'�(� >0�kÁ��<�cH�y�p�I֍�I���C�+UC?�� )�Ƹ��Dy�+�	�0����Xg7�	�q:\	j��W�8����J�6��#�ߢi�~�@���δ�O�y��?l�ڠ�ጔ\^8E˳��X�'���Dx��A}���	���ɲ G=r�`��+����ɱz��;��$�/��*�:Fu12�V�+��j�K�'�@�Exbb�2G@�`�+cx���13�� �}��LT�'�pd�'�ر�BD�]Y��H�!� Qhh�k(O�d������'/�� 7�,h5R���#@�u�N<�-�t�'��Fx��˟L@c�ýV���6���@ܙ��/>�I���쉂�xr���%�6�J@�=7"�-�~B��}�'�i%����'��U[���CK8eS�էRub����v�I4���	��iݩ��rD����y+pm���1-Ƹ��%S���'�\%FxҎST���n��N�(Sb�!H�AB�P8�Iv=�x�1�I>H�fak���0����)26ۘB�I?t� �  �a�U�<��	v��p���wv�T�B�U�<� ��RǭJ1I�13"%S�D�v�D"O�Y²΅�"�`��G���V���"OP�4d�+YȞx[�S@ڴ�@"O��"��U�@n��:�g��-Z��q"O��A.͒Z�b�X�ɠPR�|*g"OL�i��	�pcDM�H��¶"O�l��_��y{B�R-V=:���"OT%����d��`��@�Rȴ1�6"OD�j��>x�
mN�a��lZV"O�Y��?Nq@)����G�p�1"O��q�E	����m@�.�B(Z�J�ON�{`���M�O?�ɥ\�긻��מ6͈y�e�˶	 ]¥ã=:騀��k���#&�8h�6�>I���H��/��LL&�+��V�nJ1�g�i8����A�Rm��0f�n��T   �
  w    �!  �(  �1  �9  @  SF  qM  �U  �]  <d  ~j  �p  w  H}  ��  ǋ  Ď   `� u�	����Zv)C�'ll\�0"Ez+�'H�Dl�N��:O�1"�'"d7�R�)R�ĞH{b����L)<H�yi[i?zhЦ�� �7C~ݵo�?�ѧ�?1Hw

�mR{VA� t3hň4��IЌ�'�Z�*������.l�C&g����?��I+e�.}2���7X!���d&lŢB l"đ+��o��z�-�U�n�91�i:�M���'t�'d�'��$��	�$2$D�	`Ν���'�r���>/vMkR�T��;l����ȟ��ɰZG�8���+�
$�C� �~p��	۟��	⟸�I%���	�b3���`���CP�cf��*-�Y���7z����I�<	��*s�Ƥ��RE��{ƧBs}r�j?1ҡY56$�'d7p�ISK<"��|��oL� �P���ПT��ßp���$���ĔO����d����Z�"JPju�'�b$e�R8o�
�M��V��	�4��1`�i�DIyr�'�T�P5�E9]���X�^J�H�B	!ғJ	\��Ղ<�'ɊxC�jEt�x�؃-��@Z�|����t�T�K��W(]� 	ܴ�fC}���)�T��0�3CD|�ˆ"���H��-ݻzEF�g���e��#~��%�r�Ȥ?�L=��	E�P���zu[(�M[�ig�6�7.�<Hzq�ײ
��Bb�~aC�k��S�T���l�n��7-B�U(�4?�pX��J 72<�Kզ�.����fg�Q�Xy1���!�1���;�܁p��������i�7�Y����Q�ʥ*{n\�ٗ?�4�R�i���Q��ڊS����� �G�V�k��<Y�����X?�.z!K����������'j��Aҁ�`��t8�}t�uj��'��O8���O���4�Ŧ��O���2�A�{�� ���4)q�$*�����O���d>1	Vn�|C��0�IƇ���o�1@���Pb%_�~�� �!F2��M��I��
I�DE��5E��
���z��ե	N^lca(B�ByN,�'@#O&EpR�'ª�<5&�,�0!���'.m� *Nڟ���֟,�?�|
�'/P�-Y� ݌���+�7�a��#6��I��q �cq+�>p�E[��/:�7m�<��+�(t^�dNa[bY>a�����?�"h��Qo����.7V�حj���柼�	�F�����jy��'6�3}�(D�l�&���.��m�,�hѭ����/N�֑c�$%+P\�!q�5�'>ռy	f�T|(u�!�W�ƙ�'�V8���r?�f�1�S�?��'{NPh
5���K��,ɱ�
�R���I�� ��X~��
eN���%��f	� U��hO2��Fl}�Q�`�'��å�I&6��\`�J�9{�Ta�I�#�b9�?1�g�'W��X��U"nF��`!R�glp���'`h�u&�Lܮ�P��*X�`TR�'���I���?un�lA��Z�6��
�'��;�!Q�@��� G�~�%�	�'�D!���`�j�ёD��Li��x	�'+��z�bY�ep��`!�6|*�$�)Oh<j�'�"�b2�Q�0&N<9��!m%L��	�'Z�����<�x��i
�4>�I	�';2	K�(��jb�)�EK/7�"�K�'00\r�֜h���w�D�(���Z�'����f�|��l!`d����APϓo(��h�i<�w��h�o�9G��K�5��ˀ�'�2�����'���]"pĞ�1�i'V�����ߵJBπ�O�V���CO�!�&�xE�0O �C��<��/
2Bꈝ�d �?> ��ơ�A4���Kax"��7�?���p���'8��KǕ<<8�q$#F�4X� �S���ID�S�O���s�.B�t>|Q�Q9Mz��yBY��D��u��Qj�c�EԜbA,8X�2��WjD䦑&� �T77����?�'f�HP0�Z?�i;�L�
�.؂�'��<J���{�XA)��l����'lp��P�cJ��!Ə��d�:9��'����2�J�kz@�cV!�=M�B���'�X`�
�O_b[�^�y��T�
�'m�x9!J��~�<q��\�{a��AQ�i!�'�,� ��O7��'�\�� ��H?�( 1F�/!�>e;4���P�VH�ڴ�����9�ޙ��R>1�#D./��I2$�D�TŠ�	ǯ	�>�D��Ҽp���JE
��t�4ۈ�DH�G�����*L5����<����?\�h��4��	�w��$5��O����O��� 8oT4�:�P�/]���g&(<O���?�dA�rypV��"Ж����fy.z��mZy�i>U�Swy���
3vT�U�;vm�OC�q}��`��8O�b�'���'~�]��p���|��揆��dI֯�a�
�K,4|zmO����u[㔡˗Ė��fa@/
W�d��5�O�t��� �����<��ec�, C��1�O�9��,Ҽu����#��*��؀"O$���O E!+��F�	(���|REy�R�O�ⷆ���'�\��������K\:/� ����$�O.���O81�'��|��qR��ΐ&��)� �[��\�"H&tPT��("�z�B��'�R�pQ�G�iEօ�%�	�y⧛�x	���!�é</J�P4���0<Y�L՟tsٴ�?���z4���`�?hNȪ�̀;������?9���?����'��'t��sN��D.�lW��T�+�OD��	�wZ��KW.	6 ����ş�0Q����<���_{��f�'��P>8a)�џ�F�l�2�8e	 ��E�"'Yȟ��	p����	D�S�L��C���H��Ds�H-8<eh��#?�(�[����l��W�֌�`��7�dP�0���9#�Ob�$�"|���r�@� b�����R4-h�<�!� .7ͬh"���C7$���	�f�'G"�}j�L6^��)�K�	B�\DP�Ĝ
�M����?�Pv�U��Ş�?i��?���y��!b��)�uN�%�2DI�-Z&��'���h�nz�y%�L��� �����	@�f�G�L���S�YPa�RX�g�2�����d�,��d��xr��AK>٦dAşP�|�<�p!'aX�G/�;F5�\kaA�R�<G"C�=����g��4g[�lP�F͟��ɲ�HO�i:�$��r���**媢l�}�N��S��2�X�d�O����O`��;�?1���T�ýoG�PPՌV+m��sI�Wׂl˰��b�(��u�R���!bDգ<���V-^�p�+��:qr���JS�|�:a3�'�,�ڤ'����x����[�\�Z�E��?y��i��7m6�ɾ��O��*�/P�wR�u�5��م�y���Gy>�`B�I�/-l�5���P���qy���2��7m�O��d�?��!0Qk�"6�U��n_������O��g��O��p>=I���O�c��X��~Ȋ�1.�T�ށh�N-O�H"�	!$n�lXǯK�o�8T����<�j����;~[B�(��$�u�8;*�ʔ��U!�D�5)��4@ȚD-ZxCg�� e���O�$���=I����BQ�@��(��|b�Wt��6��O���|2����?�#����SU��n��z��]	�?��\�J9������Ot�g�Č���а��C+�)1Uo�)��	;����ңp=|a�F�O5U���W�x�z����֙'�t�O��B�'H6M�q��ڞO8ĵ�2." ���ᑪ��z���ϓ�?�����O�v�H��r@vm���O� ^ў�I�����<9�OǦ! ТKļ���֭��`Q�i�"�'��J9=�l� ��'R�'�r>��8�u��I�*TBtaS�t�c�逓~r���Nn�* �D�f��'A�ON�瘂_���
��M�,/f�#�	�2:9L��VN@�0i���⢛&�1�\x`a��d�����HV��d� *i�����O�IoZ<P5-͟��|�'�Ҁ˜:_p�Ё!Hl�� 5#T�I�ў�F{�'^�0�`�6�<찐oW�O�"��'�B#�>Y.O��'�?�-O�P� �4Ax�Z��_<1��§
Vv��d�O��d�O
�dº����?�����ܸ�� ���R��YP+�l*�BE
$@�2�]��@aq��'e�غ�Ŗ�=P��&j݅'�~�h�͔�;0���a۔H�>�9�h	t��9���D�5z��sv�C0V"�8��l�ܰYS�'�"�a�F�$�<����'���e��3/H��e��o�R�h��',ў���˟0�<a�l�
1�ȁ�`�,x��l���HAy�'M6M�O��u�h�`�i�B0O�	5�M	O�l�q`�7;�I���'���Ɵ@�I�����>([��uiB<p�"yΓ>�`���M�O��f-j��I�w�@��`Q>W���)��{�p�I)2��Icp
��l�N%QJ�54D��Z�S52 iӦ��O��k�X�P;2H�Ye����-�Oh�$�Ox���O~��Jc�$���)
�g�t{� C�J_"G����Oۻ����$��a�ʶ:�z��D�'x��!bJ\jٴ�?a����_7+����ܸh[ "͍|��إ�ĉR�����O���Tg�Mۺ�'��W>��O���a� ~��ҤP6-��hT�� �"���_z��B.I7Y]��"��8##q��L�bM��Q��k%�W�h*4Rԑ�0�׊�O�an��M������|!0�7���ҍ�e8�1rF�|�'"�?%B6IWMc�`��H.�h��:��"��`Ӫ�OH��7h���FU"b�W�yb廴@�O�����;���?�<EE[bʨ�{�ĝ'/�� I�^�<q�cŠ�ÅE�V;ҩ(�]�<�/�\���Q��`�a&EX�<)��
,����d�n�@\��GQ�<���G�tpJ�AP7v�%+��L�<Q���<���j�r��dJ~y2��p>1d�0pVBEP�h�5G�lH2�.�O�<� ��H��ϕ*5�\�J0-ځ��"Od�K�@��k �����\�E$����"O�)��$^�M7F!Q��Z�E!"OM�v �6\jH��A�`zN�F�'����'1�]�b	^4gY�ĸ��@|*���'���H�-�`e�dgI>v�Hc�'RZ�	��!�d|�t��A�^�I�'�tmQ��)[���2�]��'�`3��!x��Q�@J�:7j�{�'�d�rpn����y �Q�G���8����&NQ?�rwuH�mq@%C�O+�\C�8D��X��:~l�q ca$.cIQ7	4D�4���P�C�nA���O����餉4D���ra>�I@A.�7����3D��%Z%@	f���.m�^�;Ǫ<D������/@�2$W�<F�M��.�Or���)�'cFy��j֣+�8�UP^�f���'��I(o�!�4�T�V�QY2��	�'��1f��#C&��
�&ً{�Nг	�'��h�j.M�*Tصg�.m����'��.>�HC�HãVd�)��'� �S1a�4�!�Ĕ<E上(O.����'C����3'��1��@ 0��+	�'����՟j��i!�ǫra�ih	�'�ne�0��K�TQj3ŕ*q��Ac�'KA�0鋼���T�h� ��
�'��p���?t�&mR�%B�R2��;�-�H ��*m�L��^5��@�	�mF���8��C��J"����45"Be�ȓiN �Cɞ�C�,�AJ^� �Շ�x���I_�`�`
�ό�(8���ȓ]�5�p�U�]N���oT22�4��ȓC ��/U�*$�%��)vj�E{"�����x%�C� ����|5��"O�آ��ю+�EQ6�ěr���0"O	���`�&h���OB�p��"ON�TNG�_l��(��	e,�A"O���UNU�剢��,4�"O0��'�J8��
��k�$AYf�'��ɏ���&3�Y1G)נa
B��'P$��Ї�����.��tkԍ2E��(��E�ȓpL�$ c#�7����,�3Rb��sNyIA�_�B�dY���) �=��L���u�H��U�%Q�܆�;7�ec1#ˏ �`�@�	� vv��'�|�y
��j�ZG�� ����ӣ������ȓ�$�B�XXB�p��D�~
�x�ȓV�n3�ӎ?��&��x.�Ň�}˔QpF&��k��u��'A�]�Նȓ�� �E';Y�Ȳ��~z|8��I����	�-d�)�m�;��%:v�vB��?Z��)daYA��I8a�*I�dB��$�����^�Eg֡pT�^.^8B�I��ґ����1b�Zx��]�gԸC䉤	�rU �dO"0|�	�	��h$�C�ɻJj�K�e��N���X�D[�_�j�=QA�{�O&�E�1��jkr���	�1g�j�3�'��`'���2M�l����m"����'�b��*ؐ�>�aA�e1�U;�'5��V�y���ȥDZB�y��'�I u*QU����5U0 1r�'�>�R+lmHǪH�Mk�:����MFx��IY@��胄���20�ϫp��B�I2����J�;O_r)��� ~�B�)� � �Vb�9,$&
Z|��"OM��ͻ,i���djGk#�$9�"O���¥�;X��j�B(���"O8�
��C-Jh��`��kZ�H�Vj!�O��;�	)eF0� �
u�V��"O��2��L�V*&���^&3�lK�"O�03����U2��4�0�"Ox����WW�~	���΄(�Ry�R"O�Y��)¡L����"����2�U�'[�� �'��iҢ!��S���M!NO��y
�'<��Riְ)�K����E!]
�'p�`eǃ��H���tL� 	�'�HI��+9�P�čQ�br*���'��M����&%����a�4���'�������D_��H��O(�F�2��$ˉ�Q?}p,K�N$� �B�3biN�}!��S	}��P`Tl�$��RI�:{!�&\��UrD���8��rgGQ�%a!�]�H=�� �'ť�X`�`qN!�$V�\�{�b�3U�!C�dId?!򄍯W|<I�O_2rN��q��/	/,�O?=`��ɞ,L���&����@'͟w�<AR�ɿ���Q=I {�`�t�<QmH�7A�݋I�|�Nl��Ǌo�<�'� �1�j Sm�;|V�J�&c�<i&�S8�"�5z�(��B
]�<��a�]���A�neZ�����by2�آ�p>��yr��+7Κ)SG���u��T�<	�K0=_����'j/lI�u&�H�<Ag�	�-�2�LX�n�B�JD�<�A��8B����M�와��X�<�sgR����P�_�b
.��@hLWx�\�������1KJ�<�0�D%(��yC�(D�P!$h� %LU���ǻZ=�0!�j:D��3�@�j�h���C=BYp���&D�d���P/mN9*f*B�^R�8��#D��@w�r��e�\�^��7�D��y�Ѕ6�Ȥ�����T[7,��hO��˃��)*�= � W+pW�,˄����B�I6=��uMA���	3��>Di�B�Ɂ]����gꍛa#�eAP-�>�bB�;)��H�l�&Z<B�Z6l ZB��:p�2$񑨎�z�
3'@� ��C�ɁƪI0E@)J��tHZ�x��D/{��"~��Ń01Z��E���D��d[F�;�y�FDa��p�0�9��Xg�\-�yB�����!�.*�p�EID�y�Ȓ�R�N�s4���&���e���y�Ǟ.{�n��dG��x$;���y�R�F�p�������E|L)�.O"	��'�	c��8Gy谁��NDxU��'����Ջ}�4a��Ωd�	�')��[�/�>]�ژ9�䐴X��L��'�!�=s�0��ԉ��S�ܭ 	�'wV����!��
��XEӎT��:,p���N#�`�%�:�n�Yg	%�6�����ɨ� ,���9&HGh$h���Q���� L}=��So�?ɜA���>A)p��検�%�À��P��/N��#F9}�p<i3��71H��}�����_0.�FC�uIr�D{"�����ɒ7�Ѽ+��w��-N�(9*�"O�-�f	A?bQ��[���+�"O�`:��\�S6tk7�O�g�Y�"O� 0JvD��N�n�B��Y�:C^�!�"O�8c���u�~1���WR���w"O���E�/�hip�*���>Y�R�'������St�t���8)����|a���X��P)�+��v_^Րulݪe�Ն�^�~l��b�9<�m@�KD*;�e��Xo*ua ����L� l��e/ ��#��>X,���_^�}��n~�#��e���X��Y%v�j�'{h 0	�5N*T��@�`S&��`E#��5��d�4���Lʏj
�ҀkO�=iΔ��d��9v(1�M�2搕�ȓo*�����^
h�2=��ǩpv-�ȓ9h��Yр:w��iBB���B��� qx����c��U��G�0���`$D6NC�IV�tU Aʶ,�L��4xg�C��-���:ʒ�@�Ι@d�����C�*aJ�`��O� ��e'I�3|C�I�u;� ��nN�N��ՙc���{(TC�ɰbI�T2BH�:䈭J�z�B�=��C�m�O��(�6E1'�!��M�{d�z�'���ð�ۧO���e�p�L���'%�\�e�*%� �´Ȓ0tH�س�'
L=x��9c���SKY?nn�D��'�d�ð�;X���S3��`t�e9�'��ه�\b�����8z!���6�Fx��i_r���@��톀eÀ5g%<C䉍 ��A*���B�,� �܄w�C�	�bx�P� �w1j�[�"��C�	�P}�5����,+8��-�,C�I6;�Ĩ�C�S�k 4kt���:�*C�I�O�ę`��:_p<L�Q�UB\����v�dWT}Bm\$Hʈ��4vÈ������F+\�rܛ��\�rJ���ђ�?� ��=�?����?m��<�T]c��@&(�H�˜����)sB̏S(���d&H1e�v��'�NDEy�AL	gG|� ̠_��`"�aC�$+���V�-D%������ [�f�QadK��iGy����?a��i�b��\Mh�@?_b����
�6D��R�X��ɱP2�cp��x���Q������@{y򈃻�
���dO72��e1���6��'���*a�����E'!2���s��8Nd�ҠNI�!��\k�L�W+�J;�$�r�3�!�dU?r��emï4&�iGK� ]�!��M\��EĜi%0�Y�)�|�!�	P��ʒ�6 7��+�g��!�$ʠb�T�ۃ����l��]v�\�щ�"�g?�A� H��zAJ]�k��4�1e�h�<�4j�o�|�Cl�	 $Q��|�<i��@3�f,ZVG��k�pp��IQ|�<)�^�T���ÊƵwE�'�w�<	ҧ��o�4q�J�ri�-�x�<���٢q
P�$��H'�����%�O
�`���@������~&�qD"O)(�bΓM��dj0�/_���"O����%Fa\��tË�`6��S�"O� �!�%��%��*-�L+�"O����ʏ9H$^��U��4v�*��'ʤ��L��c��@>=*�0_� k3�0D�� ��$��H%�Ĉ �T�"`!D�@bV��
�ر�v�����B%!D�(��ȺI`Tۥl\�rVq�(#D� ��b�/A���
�h\�,�Z�;g@"D��[1�	; %�3�T'0�@�?�əl�"<��0��� Tx!YRk�,��"O����Y��]Jq�E61���z�"O,��g���`9!J�f��G~���"O� 5��ɭyҴ�B�EW�J��p"O���ǝ=?�z`�PoS+iH�w"OeӠf�s �QA��"3���b�I���O΢}��0�0Z�CA��]S��ۨM�@��ȓ_��&>KP�� �3tZ�ȓv�1��	C2:8NEy�^�`h�T��o\%ar�W "U�7F�(pHx��ȓAT8<RA�Аv<F�ڰEX�E�͇�jS��Qȉs�$�W�֜�\����azb����䥒&
_4��Yʧ��n;!�D�eB
����J�/xd]p�Z�l!!��@���A 7H�H�ݵM�!���<�&�� IٛZ�d��`��x�!��I~���tiɻA醱1�
˱E�џ<�Wc�'�M��?	�O&���"���^G��L�����?!�ɀ��?!���?9���?�y�O5"��
��{�樱@id�E"��D�?)yV)�D��q���k�|�
F)� m�D� #�(m#��Om�'^���y��Z�a�χ��3� ÷ ����"O:dq`LD�n������X�,����|��i>	I/O��3T'�:l'D3��U(N����X���	���&�������'�z�$'t�ҕ�G���!�"�y��$P\�O��hH%��2z�B��%GË0Ø�?Q&�L�8��?m2�j@�=z����lh�Rp+�h9?!��O@t#�>��y�,ө+֐C�Y1&(�2�Öo�2M Q��D�N�tAC�3}��9��d�q"�*�& q:��� ōS�>ɀ�O��}Γ5��!B�Z�C�Z�{���.g'�!�!�`��M�Ĉ�j����S�,��D�U��E+z!r ٙRX�$��XZ�0/��D�Te�<~$�d1��L1 ��њ���/%L2����	��I26�~�'�>6m�:(B�bCZ<<���I񯞹#D�	l��'��#��̌z`��*%N&�ЉC�Ê
)#�D����S��'�lK�Ov�����GÀ�Q.R1?����BaY�ʓI������?I`5ҧl�����%����S��8A���	:����:��$"�9O�5z%�OX�����]����kYh���Z��'�l��I(T3����6A�]"+��M��B�	G|�D�%X.$N�{��Uwp6M�O��D�<����?�*O�����۱D�h���O@�6�s0.�˦y�	[yB�'�\�'�?A+���ر��4��.�Vx6
�9�V�lqy��'5�	u��Ly2�؁v�QĄ�_$�1a#��l.>B�	6X���0�#u<���Oϝ3B�	���Ň�j�g��PB�ɯ}�d��̇v%䰣� �H��B�I�:�2<�2��C�(ZF�E6U�C�Ipfp� ��01N�8$�[��B�2u����%�6�Ƹ�τ�k�C�	�eL!so�X�ޕ��ʗ��!�$"U3 a)����̪��%�!�DV�_H�T�5�5����ظb&#<��K�?d���D�$��L�REb�S!RO�y�A$��yR�ш��xq	��;"t�� �
���'*H�B�E+`"#eܧs���H�'�! H�=�\����(P�d �������bOI�d�V����Hzk��؂-���|d���2&8f��t���'�Z9[�ID�P� �K�^ G��!z�"G#}�d�!��]�i����->ZD �Z���J�B
u�LQ;d�9K����ŋ��X�B�/24S��
�U�q2@A�?!�-Kv�zv��7qɧ��~:HB0�\a��F�M�����@�	bR� )	6�Bř�D��[p��D
b��0Ps�Oք�����S�Y�F�`O<�7&����4-��6�'���Q07�& �j���6-Fu����O���dܙje2(�CQ(n�,eH�O�\�xR1�u-��j�_-	�����:c>89�#K�6e��'<�B?u��]i��'r��'~BK��"�8��M�=�L��]0�䠃�ޒ#�`ؓ)!S K���1����'�rY(�"�
Cb�����|@8��ڜ{) 9W����P7囌۾�Y�DBV�D�^K:��0�,TS��&0����F�R$��Ѻi��6-�O.|�Q��Oq���Ц���S��IGQe�"a"����x2�F�T(>M �.�
4#6`X�O͵���HOBʧ���HN�$e(���^̔{4N՘�����Ț!�<�	����H;[wO��'$P8���c+���=@��M<�4@��ܔ���a2�ט`R��$M�? h���юq���vAY,��U�
��i!6��PcRU���gr�AD|b!Ё�^�+5��![*���%`%3��H���?���i��V����S�+�.`0��w6��ǧ<�x���hO����O�Od؁e�<*Jtic�5*/��L�]y��')V7-�O�A[��	��i$��i���%�S*�-��L��!K6�j�O���$Μ���OD�dI�gD���<ݴR[^-(� j�2���.�t�剏7�ֵ�R%ˠ"2�yƬ�8��'�!֬,��.]
�P�˓@�a�I �M�b�O� z��$�X�b�ٮ[����>�Ѱ=qBˇ�NU��yѮ��o�sЭ�'���'��Ia��� ��n���B �EU�����KsVU��'�剛'^��QU՟��d�O��i� �:7�\�gM\H��R�7dRm�c�ͻC6���̟��q`���
g�U9W!�p9�S��^?���D]�5Ⱥ�1��Ξ<�rq�c%��ͅU�E��wZ�S�5�'-�B� w`	�,\1�k�2Cj�$�D�b��O���7�'�M#a�˽R���If	�S�H�R�T	T!�H�}X9�&��1�4��ܚw�x'$�p�vx��\�a�x
D�\�W�	��Hg�8���O���]�8��X���O����O���wMhM�t�{��4����؃�F[-XEJ�䪓�{'�`@�B&/Mjc>i�O зj-#:�y����*&"��Y�pZ�*�+k�Co��e$I���T )?I�h�03��x���6K��|'��D�◟����O�"�|��Yit�1����Ujd�ȓz5��'*�����Ǎw���O�Dz�O��_��cu�%�
�U	ޔK!p�ɥfL<X�Z�X���?����?��!����O���>)rr�{>�-끭GP[z���ϵ�����W�����6�'��@���i>�Ra۷IH��`�6X�i��W<#V݆�ɗe���Ғ��U�e��g��6^��2��O��m��M{��;=R�z�G�`���-�	[��C��
� ���6\�\0!�/4���˯O�b����5�pi��:ڲ���8j>��]�lG{��	�\�l���O�Z��P��V��ذ>ץ�!0:�B�4K{�)�V́u�<����P��Z�mޖLI�Ty��o�<�B腟$���f
&ފ���#@�<�/V%F����C��''SbtSm|�<a�P-�@��3Jz��L�r��L�<�QC��	|xݫ�HR�h�>�
pKK�<A2��=n扒'-��Pwz�����`�<ɂ���(X�/Yy&��UhC_�<9�ڦ^2����E�&llH�H�Y�<ْ�ҥ!�m�x��}�OR�<a��B�o�|,a���e���tFX�<QW��$${���%���>9�`(CdW�<��I�#CEf��3�Ґ[t9P4�RP�<t��������j�j�;"g�H�<�G�ʔ���V]��ђ�k�B�<)Abݣ/w81B�.��6�P<�CYY�<��^Dy1�B�Gd`�����S�<�gMħ=�ʄ�T���u������F�<�q(�&9�A	�?^��%�SNB�<q�ّ]Ʈ�ŇշEs4�I�g�<�����'�C4?�<y�'�b�<� ���U�T2v%�.	N��d�U�<�V��O<���D�q�.����R�<�7DR�YX���HV!(�~����XM�<��`�
lB��sŃ�G�|��hJ�<)� _icF�zg�oO��h''�G�<Qd����0���u㎕q@ "D��7�B(i}�XH��	M�L�a�-D��:�Ӿ\/BCw�2�<��D&.D�t�3I�\%%G2�.��p�'D�ls���oV���Ŏ�(� �D1D�PI���M~�1�rɽ2���cS�0D��(�E�A;�������P�I.D��[�J���lx����RF�@ rO,D�����0�d@(�(�5M��4p�A/D�� ��+R��,�1�U.Mh)D"O>(7bA�5\��@d�+"\��h&"O质I�;�`��1
�Vۑ"O�e�%���p!r�֣e~(U#T"O�@ۀ��%a�B��g�/dD1�"O�i�c� Si,ŁG振!dx��"O�u#���y��1��/�-y��,�"OLLI�I�f�H�7��oq0x�"O�h��>5t�2$/��^�B�"O���M�$��� Q  "X>��f"O
t��c�W&�[�/�< ��� "O�y+K,-����0�1|#f r�"O&���L3S�s�� <
h��E"O�T���0�$�#���4t��8�Q"O�
��=>���ҏ�����3�"OFt#�� {���n����"Ot�P���16 1Ь �Tp�])V"O�2$�;m���P�
�`�q��"O�z"*5:Iʍs���
9_�!0�"O�:t��B�NH�2�
�JB�1�v"O�Y��̝"�jY�8Y)a"O�s�YS��,8e�c�Z�"O -�S퍥��p�F��,H�0��"O(����K���pj�hh��0"O����l0vw�u3 ˅�8��3�"O$�1w*F��|����r�X���"O�L�WVE�$	5��X�"O=���^�>�4�A��g�Z��"O����E�D]B���޲c�(�"O�h��R%K����߽_<�d�`"O�p��o�`$�b�N�s8�C"Ol04F߽�Q3�C��Z �4[a"O��W=�Z���lј	-��#d"ORY��m](v�XI[e�] ;%���"O�I e� p�N�s�i7D�I�"O.9����� h�����w"Od����(� ��Fጢ*�<QȠ"Oμ�h�8`�jw�������"O����K;UV��Y�����	�"OL�rfo��3đ[�Nov��"OrqS��~DF	Z��dT���"O���꜍#�:HW"N:p2"�"O��yA�K�r��+� �^��6"O��v�Z&TKH� ҆'h�tY�"O0�H��ܔ\��<3�jؼ
�蝙�"ONl(��ބA��{7ꄈV�xMW"O�P������䑖HH�90s"Ou���I�8�.Z4`���D���"Od�sE?��⴯��z]<{*O�}h�K�w|X\gL�&�Vy
�'��8��
X�}Ɗ�1S�	G�	`
�'�RH2�o�%8u���>��8 �'n lx��w�j�HޭM����'"8X���ϹY�ڹ`���4UD���'3؈���B�h�l�+!�U��]��'��p��\,+ę�_�;�RM8�'�A7/�W����셤.2~���'��@�I�cO~%Jʀ�/?�P��'�^�SeI<����4a��Y_�̀�'	^)I� [-��TDE�
QQ4!��'_]�� �(@���9��&3�X�I�'���Hp�P����p�S���t�
�'!��I�m2JH!���$
:���'d������u�^��HڜLȖ\���� �����BE��j���>e�J��"O�x��� ����7i��H�B"O� 撲#w   ζBuf���"O���Бx���Z�� fj���"O���aH��M"��{7fKVb�X�"Of���O1��䥄�nR&\�"O�mz���EUx�!P놗?klLS"Oxhh�ʒ4G�� �a
�]u�Y	�"O�
W,�l���HO�mTr"#"Ovɉ��p�"l�S�#sRCw"O�镦���t�Ei�7 �����'O���GO��f¸[d�½Rw�}�
�'���G*��?M� �f�!xDy�'��xsF�"A(8J�C�z�h�	�'\P#�ǝ
��%#�*~�:|�
�'a}[ F�#jtB@�ī�uȄ�0	�'�xAC�*�Oz��A1�ɐ��P��'jayg�+t(��� ��Fav��	�'�����j�����87<�T	�'7�����;vi�I����$(m Չ�'3��@4���͙v �
"�ri�"O��T�V�\J�d�G�}�ku��u�<	�!V��Ν�q5^OyK�r�<��̆MM,S ňiZ���$	q�<�4Ȅrf�����Z."��J7Ml�<!�;a2�M��' ��`\l�<�4jٯAF|�&.��w��]WMOj�<1e-�:~�����fL�S��A�<�e�
��=�͇*U"�p�`�a�<qs��(��<s��\�%"K�U�B�	�e�T)zÄ��R��q�w��|vxB�I�2Na�u�
�@�<�,��EC  $D�\�c�Z�Rv�B��"�x�;��$D��J",��C|�JS��	�( ��N7D�`��BN�=��mk1iS(,�ʔ�9D��0@�I�V��Ш��,e����8D�0 G60�p�1�N:���tj8D�T��ީ@I��CU�g��$i1D�����!wQ5��=S)|���9D��С�N.q��H$�;FN�s�"D�$S!�̣5����u̞[(2�D?D����Fb6l|�"��tj�%ȗ!D����ܻ vB�G��m��}p�:D��HF��.x�l,z�)\20w��8#N7D�����d�X�(�:xm�K)D�����s�,9Ra��
Yd�!C�,D��
�`� 4�L�&���]^Jc@�+D�\�O�hM��Yẹ(�\�G(D��ɇ�*�Дr`Ǌ�|KT�3j&D��C5		ev�z1e��kQ ��d�#D�DY�����6J�6�"X���?D�D�Tc��PV��3�OQ~ZP�e?D���A�؝x�!{Q$Bj�.�91G>D�h0�H��6f���Z��s��B�<q�܏�0���@�(T� ���C{�<Ag��#�H�@$M;er��a�	u�<�c�ߌ)�����6K�>x�!��m�<ѧ���Ra�E�3�:�"�`�<�	�}3��HBG�2��T�%��a�<��*���Y�G�K�2?�`��/Iu�<�#��:`�:�)�E?A�N�X��s�<Q _6O���ã�7� U�s$�C�<��C�,T^t�0�J�VzI�� E|�<Y�9���*�;-Ȱ"F~�<� �Z2'J7]��
�`�()��D��"O�(��E�g+�Q��[�"Ȱ��%"O.���i�@؈DI��#I��R"O*�	����8�# N� {x��E"OFA�$΀"
�
\���F�m�4H�"O�dˤ�Ϗbk���ݣ[���"O�%�A$I�=�Q�Qd͂An`ۃ"O�	��l�&�Z``%%�X�C�"O4���ך-�p8!�y��1e"O���b�$TjP��F�\ �"O�aWcӵW�+W��5R�<�i�"O��sЊ��i�k�Ab	×"O<�
�#D?~�J%+'��
����"Ov����7O�D�T�R5[�t�c�"O^I7iܢ<�Th {�W�c�!��/��p���-KSZ�i�n!�$��!bfn�BP̸��ƅ�O^!�D��09��0�B�lR�@�V!򤎊\R񂳀��]���Iᮋ�(C!�%�����I;wlrZDM�'w�!�$�=�ՙ�F)bwl�JT�B;t!�$��2�������ZY|s4�:-;!�dȩ>4J���ǋ/<Vi£a�
3!�N>5=�u��լ-��@ �2$!�~`<T	1h�mY���iT"�!�.qf��f%�W�T��HV�w�!��(�!Ct+Ӊ,A��#�f�e�!�dD#��I�'��/!N =��C�g�!�Ӑl���-�2.@�FFS�].!�dSr��|	��׬@�Ȁ��d!�D܀Q��z�:w��tpC�D�C!�$�U �pkT��ӊ=ʳ�L�E!��J#v[lq�Q �Y�`(Y��ސd�z�i&8
���5 ���Xm(�		�#"J����G�g(�1��X�<�T��0&�Z�@��2D�����o�<���[}X0ҭ@~��A6h�R�<y0*�B�ڑ7@jO�iɱ�!T��$#��W�̐B�,�N,j��5�"D��Ŕ�-�<d�#!ӣ�B ��)!D����I��:�,��DR"L�zU�s, D��u(ԅ*V��s�*-��l�W:D��ՠ�<^��Q�f�!F�x�K+D��h�dB�MNP�#iƣWb0Pk�	.D�|�V
�
�:��郐Z��Egc*D��y��� Z@H��-#�d�P�g,D��+C&��F�bXk��%%.��P�+D�$���-U�f)YT�ņ+���Cf*D�$��
�E�L0�"�B�4�Z��=D�d����:m�>�qȏ.�	�ҁ!D��#��Q����c	Q*IF��ir�-D�0 g��,Y�8Q���Ӭ)hʤ�$*D��p�*#����<,��%[&+D�$8�!B�2t�Y{��%j�&\J�"*ړI�m���Z��:F�r鹖�m���G�<�Ĉ� �s,`���BC��y2J۶<������d�Dd��%��?ɡNA
�j�@tJL&hR�7N��#}ʣ��2�D�����#&��"��C��y��ۯ�`�q㥑{dtiD��)]8���Φ5��e���41�_>���Bh9D��` �B�<�R�r6�Q&��>q4�Y6UĦ�B��D˦ 0�'$j��0a���f8��I�h�"�,qC��'/�-@P9+H5�C+���!N>�G#�1�?�f�!���� �\���h���җ~Z�Ո�h	=*�jwa�O�!�(w%�s��P%&5[��CGv
�pW��*g�Uc HQ�%���sb��8�M��l�Tˁ����C���u�����SC�r<��K���xIHէX2�L�9�BW?�0]{����4�
T#c�̊k���
ۥWxHJѯH%���� ���tn�4qq8H� H�z���'S���$��0� ��c*2N���"��	�B:^�vc_;ٸ���=R�0)���.Jwv���+��Y��������M�H�� �O6X;�-�,M"�C`��*k7�q��e��s"��-Zd��D�.n�r�v�J�P��� B��y��[}s  9K�?yb<D�K+<[�d�3�s�4��%�� >����S]3�Ik>= @�[�y$2R����M��A��-��(���0?Y�@Nן��4�V�,�����
�m�t���I��,�$��W��1�H߯HؔY�0�F�l!����N��]\��@w�Q�m��	�����O�Hҵ�{���{mK<�:90��+)z�-Z��D, q�ճ ��"����hղ%��Q-+ �a��I8�и���ºx^4ih����d���	�*P�	��A�� ����II`eU� o����X�B���(5� �2A�N�n%J���ŝ��!��B�A#v,�7��]ca�n�x�K$�"G�iq�+�v>�����$˧4WX��˼{`N��l�e8vLY;o�2�j�_b�<���e|���'�F��j�� ���Z�K�8�B�c&��F* �  ���%����Z	�PQ��S��ڹ ��M7��<��C�]ڸ"�]]@.��2+Λ1;���)?6a�Ю+�b��g�y`z���'0�a��4l,Td���d&�ēM"2�*cI�8`��&=vli�".��RV����a���ًyX���7����R"O����+K�e���m��b�P͠�Lh8��[T�o���+��<z���/#�T$�Y��.\|`���cٹu�,��.oY���@F(���2z��+��аRd\��`�ʁ\��)n�"e�T���:X�Q8��O�*�`���^�-�3�\�	��(���7�'�z�I��ߴ�?���~���pT�":��]Y%Ń6~42ăc��]�)�q�Յu�h�E�'|<ܚGᗐ"	Kf㔄x�p*�O�e�AH['$��ܴr<�ܛE埀,]�	Jd眔XZzpo��°�a�Ҡ%�ܔBA�:i���#"O|�	�I�k�~��*�v�lg�g�8�u��?���b�m!������IE�Qlf��d��sq��0K���s��L� �� �O�qu�͡�1���P0@�kĩ��6���y��T�e��k�@���g(�q�2�"O>�{�j%S�O��!G�B2X����^����0"O�:��LqzMAG�M�c�y҅�|B�]�#/�Oq�.�#@�Y@���k���|����"Or�І-̠@	���7i�ƽ*1"OP�qu��Y6-JblYU���R"O���r/NT�&��#��g���pa"OH��c�l��@��kϴJ�ܽ�"Ort�	@�N�;�ޠ���@"O�$��E�b���!���3��̂"O\E���0g��	�bדM,��Z�"O��M.kܺ� �G�`uR9��"O��p+�$g��e����2��<�"O���&؋
�Xbf���2�n�1"O��a���"m�S@��)Puj4"O,���Q����'E;`i��ȥ"O�$�r(�EW(Z$hP"OB�YB؁4kF-�������g"O�Ac�o��6�*�p�� ���"O�0A���>`�4�r3��=Y@�9�"O����"� b&�Yb񪖂�T���"OTA��H�F�*�YGCD�t�����"OZT��R2G���
'��W B-z�"O��s�R�>�d�`���%���y�\�.a�ӈع&͜(x��'�y���'�:7/��_-P�횄�y�)�'j�V����߸U��a�g�ȏ�y�AT�q��s#�T�P��!d��y���)�������\��
$L˩�yb!ؑ)��ݨb
�P��5���,�y�̴^�"E�բ�Vf�R�%$�y§RT*pA��*U��{`��&�y���83;���(P�\�aK0�y��^ j��3��KO��p�Ɠ5�y2�ÅT���ӄ�
F�숓���3�yr%�D�piCF
�z�H�[�����y
� Đ�!�T�e�ŋu�*T�̸*�"O���D�}�f��R�v��0��"Oث��T��.�(��!?�1�"O� �ꍺ@W�1��.78�ܖ��y�N�-.�)BA��n�´���[?�y2��XaH!�&K����*�劎��O��G1ʧ:�n����	x �X�+Ӎ^|���J�|�  e��c�%����L� ��U�A:��S�O�̣S��z��ə�ΥF3���'���+#��*L&D"7J:?O�@��O�M�@f�4��݃Ǔ:����V���i�N� HR9;F8����2�v�.	��PEIg���d�+a�<���L�@ՔՆ��Zʨ���9_,����o܊p`�Gx�
154�SIK2>X��3���1�)���$=N)����y��M�M��(@��E�~I^��T�1K�u� ǜ"/\���՘E`6�s����%R�utH�Pq�=@��5��b5D��bk �T��ݑ�Z*�}b䖡j��I1'�=0������V�n����kՊ���J_�1��8��+ե#�h��Ĝ39?R\8f���+U��8"z��y��
 c�(Ҭ©3�2 ��'���!��6_�<xr��ӓ}�r8ш}�l��\�4m�B�38[|����Y���e7����
���ר�8E8��ȓosDt���!K� �b���*�8�2OT��^� Vk����H��9ϓs����j����$�V �1�ȓ5P�b�`�k,��� -6 �EY�ilm`u�%uŢ���uw %�M#lpHsm�%.��|�FIA$D���I�/Q((�����"F��4�K�[��ܐ�mmcrI��ǉӺ��C�-�0?)4hX?|���U@�2Ax��׋�r�$a��`����!}���GCD!	K�o:³�J�d�m
`eH0 \���-�Y�<�Ɇ.U�Pb�\)����3Al�PU-5a��ʚ�h̛����<q2E�6Ö]��ي!�DE�a�V�<Y�/�0C��@p3��)A�Ҩ��UyR1��$w���,P�n����ԨO�mX��)d5�Z�N�`��$�'j$�"�I2�lZ�ȉ���	�lT
:�LKf�Ѷ6A�Y�%'̼�p?�&*�)WY��ǅM3H�&��"* P�t��$�	���Í](�Ob����l�q��9��'v�4<��'^��Y�)�?
��� CKr�~���'q�P�Qd90���S��}� ��6i!���w
әU�8$��e�t�<���[�U�q'�V1F�Y9��]���D�"�T�v
U���3��	xa���t�B)�Tٙ��^R���I�L�	Ǎ)�$� ��8��L���(%�p��O(�.t�T[u�ʛ�lP;�/�]Q���sb[�������4�>9V����1o�������y�)�6��qe�ݲ#$&0m���y���,9F�|��)Q��	;�DN���T� ��>�!�$rᵎ�;n=�(�"U,�΀�xR�U�v��zBF.�����m��w�j�W!��y���#N=a���C>\���M��yb֟'��P����~�
q���\0�yRCi��}��ω	$6�����y��=Z��Q�`HFu(��V
(�yRG P�攸W��j��`e��y2�ϏGH����Ĭh�d�4�º�y��]�7�!a�����f��yb˯[��P��`zi��r�U�y�Ɂb��c�P�y�xh�%����y$�2tִMKpKZl1���y�NQ3�,E��&^c L���ʍ�yB��4�6A�,����s/8�yҤ��.�fH���T	0�2��R��y�I�`��T�#�� s�d�'���yB�]�R�� �K~�R�jdÓ$�y
��*�d)�0#�'ֿ�>��ȓ�����Q�Y�[`�F�$&	��:��j��I ��NX�8��S�? �@�ӭ+�ʗi�$ol1�"O"��gc>X���*��
o��{"O�<�"���E��q(*1��"O΁��NL�R�:�zBH)��a��"O5c�hۂ�,����T�d�D��2"O�4�a�:X��E+q�I�
Ԥ݋&"Of�R�f�`FV��Ff�2V϶("F"O�JBƍ1U��[V��j譋%"O�@v)мC�|��% �_V�(�"Oֈra�+JX��(D!Zg��4"Oz �d�x�����K/z�)�F"OL���O%n�� �K��ON�Ă�"O$�� �5k����-ǳXݢXJ"On� /Ξ��!S��N�`�T�r�"O�ܐ�jͥa̸��t��b��YY�"O��Hc]�Tk��
Uͬ! ���"O��X�@0�L�Z`L�&5���w"O��ա0���B1�^�y$��r�'1*�R	R)��ձs-���s
�'РT(qf:w,�T9c�J���0	�'����W���K:5;�ڴK�4(�'CJ���S%9P$���� U�0t��'X���j�*�,���K�R��'�D�a�X&/�>�A���	r���
�'Ga��3d�d0Z�f�eT$��'ULq��7me��zb`���\5��'(�آt�������%��1=F��	�'�%'�>R/�]k�̗g�$A��(΂�CF)˦:�S���(04��ȓl�8�a5�B 24ܐ#hY���ȓl(���u��U�<�N�%h����,���Z�����b� Sen���^��H��U�X���d@3�a�ȓJ�^=�%�0t��넶aB�����ec# U�]暭��K۝Q n�ȓ}a<��vl�6�(�1݁V#��ȓt4\� D|Ȁ}Rǚ�e����	"@�TŰ$mQ�\�Ry�r�h�p�����,����+�
`�!�۱�  �)*8}��ڴ�S�@�!�DR�T5d�3���c���@�
��!�D�\���I��4N���d�U�@�!�ā�U#�H�`Ԓ�n ���0�PyҠN�-��Y� �R�/�.h�-P�y2�*	�̈"k� (?�UA7����y��C'����u�ßx���N��y��G�2���nC���H�/C!�yR#:s�(�� 3NAae�D��y���6�h���i2�6�`� ��y�	-�Lј�G�N�r�]2�yc^�{���b/[M,�q �R6�y¢�=\���f���25�ͽ�yB�@-M���s)Y�f�ػD���y�(�S*��)3
���1;t��y'\6 �� P��^�-��г�� ��ybK{�$�0�o�*v�L���Q�y���"V�.P i
,i�~���炠�y"���g�6�������׊��y�J��WgfUh�C�E��%菭�y���<|�F�{Cb���Pm�Yp��'�b����R�t��@��! ]�Xa	�'�X2t,V�~�,�2� �����'a����
3��������x�'�t4���E�D�J��բT�b����'���5�#����i�
V�d!z��� nP"�`�=��8��A6���""O�H2� ;O���A��6R��hU"O�)�#�Q�/�܌S�I�'��1"O���	A��x�(,Y�{�"O܈jB�@]iJ����W�P��"O.U�Q'ė�Pȃ�eZ�=hM�"O�\��C �T)�O�X�2"O��yr�X����(G�eX��"O��ՈW�, ��E��@U��� "Ojxy�g���igB(WY�l�3"O@���(i�Tp��`H
#N����"OZ���#��#rdU�7o�	?��c"O����S�b=�<:�Ύ<1�0��"O`=�U�
,��x��H-.�1��"OL����=We����h��K�ɉ�"OT�3ԇM�'��ZS���(�,�(4"Ob5tF�N�"����],e�VLcu"O}q�č�C.x�tـu����"O�����N/v��D+�)�YC�"Oj��):%,%	���d�>@�"O,]
2 6�XaVE�z�d̐�"O�P����`��yQ���N��h�0"OIpp�S#Bҍ:��R�V��c�"O4ݨ�g��I!4�Q������3r"O�fn��M���Br��@Ie"O����ʚd�t�PgW�N�V���"O(��ч�]r�d����]2t;"Oل���[d���~�<��0"OxQ��¢aVmI�IM%h��U�t"O������e熸�'�[]�>�2�"OD�1�G�*zľ��g猇��B�"O �ؓ�W�n�*�	6F�+B
���"O8J�	3��!�E�*a)4�:"O�]X�Ʃ57���C�>��T9"O��#�lArX�AÇ%PG���"O*I��.�7�����'ځg4��"O�0Z&��6]�vh��FY�R�6�u"O�y�Dh�!X�q��_�"���[�"O(��N�jC�x�D�N����"O�	��l�xO@,R�B��޽6"O�U��HD�%�%a ��2I��S"Ot�Ókx�����*v�`��"O�ܱ3@Lb8!*�)+�6��"O`H8l
x=3�_?o�� ��"O�J`eѝ�F�a�˯q���˄"Ov�8F�M4 "x��%.S�t�p�@"OB��2�R���uC�M/c���'"OP�@��N.$5JE��e��J����"O:c'�Nw;���b
.v�e� "O��XaA� wzV���
5��+7"Ot�G�G�VŊ�,�!�1h�"O
$��gY%cn�mb��=Ji�"O��1���&�x��@�W�h8��p�"Ov��;<��'N�^!(�4"O�� F��q��pրր�ju�"O\�D�N�	��B��Ӗ7�J��"O��*��&W���rh�,X^0��"Op�*@m�TF��(��MO&���"O�)Zd�ޫ;#R� �>Yڤ�"Oޙ� �َ�,|`���BS��9"OT��H�%�$Yz�IP'b=^��"O�ԙ1C5I���I�
� d"On-�3��F���ʑ�،�yS"Oⴃ`K]!l�����M^�a��!�� M�����X^8c�,�-T��"O��xF�)S1��J�&�c�ʼRW"O�����(Y����O�8.�hB"O��rb�=L��qa���n*8�	�"Or���i
7`��k�<]**�Q"O�dqO6x|$X�
�' ��yY�"O`d ��(L�d����A�nm0�"O��Rc�G4!=��� �ػ�<��R"O
\�$O�3�X$cP��e����"O�qX6��I@�`����A��"O���AlA(I�6�P7���:�zH[�"O�x+%,�!_縙��쎌\er�"OB�{��B�B��D�n�0IZ��*�"O�Q�WBЯs� ���D�&�Pݲ�"Oj]	#�\�u�\�z��


��A��'s:sw�^�~!r�IG�>%6���'9t� 䘜V�H���O��9�'�z�X��$ �N�rV� �[����'�"-k��iij4#�D�_�d��'��щ��w|���Ej�X^�5�'�h���ВV��Q ���5g���'tR ��ҖQ#�eyE��'�laR
�'ߒd"ߜ4�.}�TOK����	�'C<Q�ϛ�
r4��#)�	�B	�'Tj��P�Xވb�	�X����';��3̝�JI���u@��Vf���'���C��C l�.m� ŋ�`�D1K�'��8b�I+o���Ǫ�Y�-h�y��'WF	J��d��c�@7N��$Z�'�J��C@�%*z]��Ȑ>��8�'\Lx��d�(nέ��Z<�\؈�'D��Q��K��\�S��,~��'�2��r�͉	�:��JM'ȸq��'kR�SqK��Z��$�
���'��r�7�����lۓ�ܕR�'Lx�8�.J|l���EZ�[�r(��'���E_ r��J��*LVx��'�^�H��}R>�����"Ot���w�V4�C�M{�t	�"ODm��H�6U��ȸ��4`�db�"ON��0/P'�^�y��]57r\d�W"On�Q��:r��Kv��9Bm����"O�`�tB�Q{V1��U�a\�u0!"O�)�t� T�,���OJ�I�"O��;$ )a�ΙǠ¹s&����"O�}��j�y�"ɳ��:*#�P#"O@q�,�p	���o�S�ڤ3!�dAV�!�CC�P"Rua�h6!�����C��Șn8E�3�j!�d�fKfq����K��DIcĕ�NV!�R=T�P����TEؘ��C�V��!��5N���A��8����J!�䃮#0��+Dᐌ,B�2gL�"v�!�d�:Z��m1�'ܸe0Rl���ȉW�!�$W����F0(0��S�D;�!�dC�H�ތy'\�Z!��i% �/z!���,}=&��2#�,g��:5BU)h!��c�v�:c�=8K�D`��/�!�D�>�Hq�&��=������tc!�d�Jl:-�?9�H��E�!�ݝm�r�9@n�
dkfE�����z�!���ܘj`J�fn��&b	�Fv!��O�⩸A��p}:��Ί�7�!�4V������#1�X�i͌�d_!�� ��*&G�Tԋg*ۦ$fƄ�w"O$lBs�%�<M)2T3!]p$�c"O�0��!7S�U���5%�p��"O�t�pѢ)˔d�E$P	P>��Ӵ"O���������R��[�k�d"R"O���.ZhB��F)B'f��I�"O�9�� �*� ��(鬹31"Oj!��*�9	���a�4m��]*U"O*��cf\.{j�����0:�����"O:�Ȗ�:=:^�:���+��""O�|Xc�W�d�#OY/_��˅"O"(�0�� +?4���ŗjo���"Ol��T�=׈l�m/R��i��"O|�եY�TN�I3a� �܌;�"O EZ��ɦ.䆤I��Z�����"O~8�A@T�Xll� |֬��"O��9��FE�:�"���^!�"OF��"�?<�e"��I��[a"O�Q�!F�����T��ֽq�!�$
#h �S��Է3B*@����!�D�'z��p�d|+�	Тc�!��/o��s�.E54|��dbW(1�!��<�P��f�Q�=I�d�Ǡ�W�!�T���ёW�Ĕ+,��Æ��<�!��+C�~5�w혭5'��Q�W+/!���XXxp�!F���#�NU!��
��x��援�� (��#MP!��ũ(�h�ŕ��4��ڒ;!�ʉ=@����+-� ]!k�wJ!�d�!1P3�C�R����׃C�!����$R#+߈�E��*�--�!��	�3��[�n��	�8���>H!�D��~�[� �Se�ܚG��@D!��E���i%O�d|lI#�G';6!��C�j��$�9Z`�����l!�DRhs`H���T-_�	����Z�!�D�L����À�"2Z}��'�!�X�)~5��$�m�C�=!�!�^�
��%�0C�`�ӫE+!�$U#$(��hI�l[z}�c��d�!��
�(<ۗ�ZP ��Cd��?�!�3iq���f�]O4$��Bǳz!��_6x� �Pt�Z�8M:�D�[a!�$�3PT�Cׇ��}@���-ܐ�!��[�v9�c�K�7�b�.�bK!�mt�fD�-?�nU����
7>!�O�=袅�+�^��d��F!�ʡ\?@�c��<W��U�E㍘X�!��@�.�ɰv��;��]��Q�<!�ەR�"�Rc��Q�ݸD��5!�Č�l���Q$K8pp�2�#�4s!�$��;s��[7�ȍc����	- !�$�� x
�!ͧIV��H��Dc!�DQ*w�
ث�߄9M�ѯ� �!�����P�Jŏ?;N�
B�׭]�!�WP�R���"D��D��-�!��,-?,�!OE�%���k�C��~�!��R��M��՝c#:,�6�G�d�!�$�+�M��-�@�~|��×J:!�1��!���K9D�N5ء��#2!��G�\�rDs�dȈ�a��G@	]!�$_�(� ���:�z�����a!���7�t �� AwB@r��S�'!�䆴!P@�#�^9,a�6K�s:!�� ��Hv�A��\)��ͻ2���d"O�����93���v��Q�0��"O$��ф�>p&�a��o眄K"O��c1��
�d� 2��C�LNm�<Y���57OB1�eBлꞌF��Q�<s�
�a�HdbH9&���v��L�<��o�I����tgҲ.}z�H�L�<�d��#Q:��f�ȱ"��<b�+Bm�<�#�Ҡ(�(���%P�c�THs�<�f�S�b���+<���*l�<�gf�3�Rd�P!�H�ZQ����g�<)�a+
���ї D����Y�<	�h[�{�.�xU�:u�N�
���~�<�tO^�#I�@�$g9&�N��Ĭ�@�<���S;tx�A�;X����G�{�<���L?VȜ��,�(h��LB�<�Fil[��RARs���I I�<�q��-$��	����U����OPn�<	Daթ���D�#&�D��qN	j�<4����e�^�dy�	O}�<���@+1�p�c��%�%0^�C�	�Z�ۥ�ś+���B��^�B�	�\��A�Яt�`+q Ǘ>iB�-�N}��N�y��@���H�/
B�-Pd��6i��M{�] �`F���C�	I�ԉY��.'|^(�%�ɰ0�C�ɝc�� ����`�@���B�,C�	�kC(d	�=>衁�;)�B�I9��v�։*>|����u��B����e��%�G�*1p�,C�C�I�RX���%��I]�x�KQ:9,�C�I�Q�p� @�(O���#;4�C�ɀ^��lI�DR�q�1j��F�~�vC�	b@����I�&����OXܬC䉺|M&���d��yl�i��Tg�B�	�A@�uC��E����`�Z�B�ɂm�V��/@��Ҽ����RB�I�:��Z�+ ���$h�q2B�ɄE�N]�D�ˍU{�@�[��<C�I=!�6pJ�&��f��uXC�X�6:C�I�5($��FAl~�(R���h@nB�Ɏ\�0p�P�vv ! �W6i�C��6\N�8��	(d�x�[�6D�H��̋Iy���VɌ_v��Q�l"D���"E�d)�	�C�%1y�!p D�����L {��%�Gև ��S�*D�,M�<�~1����t�����h*D� ��酪t1��ᘓS
�����&D�̰���|3�EyEĘ�M8� �T�/D�(񨗺�<�!CIگ\�̀�ƌ,D�\���ؗR��A�ٞ���Z�)D�H
�B�u��VJY��l+�h&D�0;��T/	p|��sBX�wb�|�1	&D�lE5��\��A:_w�Œ%/1D�1PM۰u��x��S
h��`�+D�P���Re�	;���6/�~��#)D�l[fƙ��z�Q�̙VMt�s�(D�x15�ڠkېd��&�� ��`{��'D��*ō�.d����J�|�n;tj3D����K���Ш�K�\.�Ғ-2D��@Ť��AV��H\bg�Q���,D����m`�0'��T��E@�0D� �]� ܔM��/544���,D�\��d�PO
��a�+t~"|[��*D�� �xY���5U�Ɖ�!mJR ��"O<�r���C�h<�Ì�&(�ii�"O����Y6��$8���1}��"O��j��*��M�b�FxQ.LK"OTt
�h̪l�Pl	7oĲQ#n0aA"O<@(3퇟T�"q�7�"�"O�����$����ī�����"O8|��%\0e7^�Q�@�:-��D@c"O�pZa�%
�
4S�nɓi�m�"O���2��IL��V�<h�z�	�"O*Y�'�<fd,�`�"&2�>=*�"O� @7�G2fh��ٗ"O��R�`�	�\��a�$.g��{�"O�2E(�� �)���<Z-PE"O��eL�� �Ju�����"OI�2gH�3~Q���W�A
"Oju���|��Y�a	�Pd�4"O,�pd��|r��ځ��ݠ�)��|��'�:����N84;�`�65�&�
�'0d��t�X=`�b��A�)%���B�'}:��b`]Mo4a���!&�
�Z�'-������x�P/G�h�H�
�'Q4Ep���$�h�p	�VnЈ�'0�|+0扫2:�|�W�/&��=r�'U�}��Q�?Ђm �%-����'zܐ*�jB>�|���[4?,�	�'E��B��OYd���`֤5`)	�'��� #D����%H&�<{��)��M�jx�͊�3c��qBn���!�$گ+��g
@P8Cw"@�D�!�X�v���,Ni��D'�4F�!���>&,`y��е��\�S
G�%�!�dۖ,� y)5E��*�Z �3*�.>X!�TȦe�p#G 
�a94��{���G+D�0�Q���~�q���v9.��P�(O #=�U�W5\'"LQ�g�K]���E�w�<q�B�92X�|C��(�,�I
�r~B�.�S�O��@q��)]��;���4(:h2	�'A�P�ɽ��́���#/��9P	�'Kh $��
� ���'��5;�'�ce����Q�l](�F�Y�'�5�aU��Th0'�Y�e젢�'�NL�"�C�)�O�_�����|�<Qpe=Ϛ�1#k�>UKH�4��^�<9H_	�n�z��O�64(|�\�<鴂_A�fm�o5uK4�;�EW�<� hX�rZ=P��TQB��Q�g��B�ɚ0W$X�ba�����K���s�B䉍H80`d�=a�d��(�>��C�ɥ ^]�6���f8��Q�9�\B�I���=��J��^�<����ܮ�B�ɫ80���<��r�oϢ1	XB�	�a9���>q��r@M'[4B�ɕxk�,���Sd*�t�MGb]6B�	;A<�iTđT�~$��#Z
�"B�I�b��m9㈐8AD���NB*X�FC�ɫ
c2T���9Up�!ՄD�.C�I�Ю�B
�R�(���{yC�I�E���]�+���vO���B�	$��yjr.�y]�\hb�S�}��B�I((�`��!�,6Gx4�TGR�P�pB��l����ICiâqЧ��U��C�I"��<��Č6�����+X�b�B�I�+l����JE���� ���� >����[.}�m�%�62�`�"O���|
r�x���j-B4Q�"O� #Vi�
bf�̈�D#i|tx�"ODD8���e{�$Y�Uz@�3"Om�!��/J��7AH��vE	�"OL�#���8f|��r�����W"O���/�`���A��I�v�J�"O��IS:ڨM  �O�[t��;�"O��;�,X�����a�~��24"OB0j��-@�4h�Jt~�l�s"O��ť��=P�����36|�;�"O,5)1#�<Q\M��"<%x��I�"O�u��G�Y^�4!���Z"O�M�S#^o�!�D�кd�j�R6"O���W�O�/zp�a7㊆d��YБ"O��z%��!�x@O�?�D���"O�9Ҁ�I4ݩ�@ùà0��"O:x���Q�c�����N��m�"OP��C��.v� ƃ30��͈�"O��Y�P�>�Jq��B4V���	�"ODpAtŎ7d��b-	U�!٣"O���b�9=TM�����}�"O���^(�T�'�րc7Ե��"O��c@�ئu��Q�� ",xYRV"O怺�͚f�ΰ�q�G�')͓�"O2i���>;���%���rp*x��"O����I]� R Uk�*_bNp�"O(у�S�]W$����Cp|$!�"O2�ru�1
"��(F`�1?
�84"O�i0�H��Q�Z� �L�
�-�"Ofm�R�@]/��!kJ����"O�@s�_�(h�0#�ċ~�DPS�"O�i�mB$y~Hqw�Z�z�V��A"O:�[��W�<
�苏]��MJ�"ODE��m���N��� ��"O*]�RÜ%>��\��b!�~]H�"O�\pp^������ƅ[��MP�"O�l�㊷s�S��N����s�"O�����;s阐�%�?�Xc5"O�����?^t<veM!=�Px�2"O.HCV�_,_���P��OZ~��s"O����`R�������Dd�U��"O�X�g٧��-��lZ�Hm��"O&�*B��2dC�Z�ǋMZ8���"O xŊ��n�-���T By����'�b��8Ca�b����F.�u�r!ʯUi\q�9/��$�O���Oa:���O��$�O^Acc�r��i�a_�T�ԕagJ�)p���Bgo�uZe*� C��s4m��C�Q��/�e¹+wa�:���
�� R^���݉k��#Ӥ���
��#%�9�MɅ� c�9���^�
 f�,�ȸP6�ɪH5���հ�M����$ӼR����]�|��fƇt���Y��ٽo5 E2f�`�'aayR�N�r>�c���f�T�T�ܪ4e����6Iܘ�lɟ!��r�`L��u��'�"�S���;bR��U΅�f���	0%\u(����'�2�'BX�����O�MۦɅ�v�<$�!Bk���@/#�T�s�F9E1|@���@�h�<i��J63��i�r�1sT���&�v��|s!	�< ul�h��,2�֕�B�әM��+Sg���L�1����MC�i��V?i Q0S��ِ�±!�\���e����DY��?��$�"z�x��r�t��Lk O�H8����4_盦�i��$� ��@L+^%c.T8�U��sQ���M+��?�+���8PI�Or�dӖ5(c�A5+m�x�mӒu�a��e�t�В��P5ߦ�P�֭^~�Q��A�R�O��Ա����CE�(��Ȼp����T�iM��GCP�Yo�u�a�.�Ms$!�p|� oL6|w����A�V����C� ^+p"�Aґ�˦��c�O��o���M�������L�:�fU��M��V���b�D��~�'��mX�p���+@�9C �����01��/��M+Ӹi��'��S-��q8��F"_
5��HAT$�����?��P�*~�@���?9���?ه����r�|�k�Ny�����=��X���$%�,�q�j�YJ�[���u�|��S�P�F�іg)�� ����U�c3�P!�H�����C -��1�'#C��X  �ºc|��$.�@s�C0���z�Ƭ��%Ҵe�LA��5*�'������?1�x��'<"U�DJ�G�j-�1ѳA��y@�!R鵟|�Iܟ�'��}*�*Ǳ)?Xj$�|��A�ժ��7�ɦ	%���?��'�8i1a*Ʊ�`�Z�BG�$HX�s�H.;,Y���'l��'[Bϛ���'�d���bu�b���n��1*�W�H~B=�A��2.T����bں}#��X8,���dZ1\�!h�l����S��I�='����K�7-��nZ�2_H4�p �2������#�@�OŢ��'�D��A�.��i�w}\ܓ����>)�7��Or˓�?!��?������������^�{Ș�ygi���yr,-A��k��^n���Ǝ��~"eC)A��7�<Q�N"������O�B���ɒI�U����P)�)s���d�Oz�$؝=��TO3&�	�B��Ri�S���D��0��EH)�D��a�Ș=�t;��#H�t���D!=��	�rCƘ4Ul�+ԉ�g&H��O��R���>�b�`B�8l$��j�@�O�alZ��MS����i�:e-��8��Q�vl�$�bSdˆ]Sߴ��'��#}��Z�٪1�U>>��Lar�1����d���ߴ�M;5���6��&�_�;�~�
�Jq�'��' �O"i��  �   d   Ĵ���	��Z�tI�/ʜ�cd�<��k٥���qe�H�4M��\70<����z@�v*ɾE P4%�M�R]M�Q� �6��Ϧy۴8��$ �Ibybl� \�!����V��XS%�,8@ɲ0�PK9�=a�#?t�7M�dn8,��W*¹
�c�.2���&�ʠ�"��RG�I�Us �j3͔;���<2Jڽ��%W� 9�P&�92���Ej�6*;�v�tTx��/0�H5�V%�?)�'�������%g� $�r���9F�(�fbSA}��{��c˧~f���'�(� >0�kÁ��<�cH�y�p�I֍�I���C�+UC?�� )�Ƹ��Dy�+�	�0����Xg7�	�q:\	j��W�8����J�6��#�ߢi�~�@���δ�O�y��?l�ڠ�ጔ\^8E˳��X�'���Dx��A}���	���ɲ G=r�`��+����ɱz��;��$�/��*�:Fu12�V�+��j�K�'�@�Exbb�2G@�`�+cx���13�� �}��LT�'�pd�'�ر�BD�]Y��H�!� Qhh�k(O�d������'/�� 7�,h5R���#@�u�N<�-�t�'��Fx��˟L@c�ýV���6���@ܙ��/>�I���쉂�xr���%�6�J@�=7"�-�~B��}�'�i%����'��U[���CK8eS�էRub����v�I4���	��iݩ��rD����y+pm���1-Ƹ��%S���'�\%FxҎST���n��N�(Sb�!H�AB�P8�Iv=�x�1�I>H�fak���0����)26ۘB�I?t� �  �7j<C���Ci8,|�)h�E&}r{�'.��=1UI�jR�IJ�!v�V�"2��ʦ݊�ቮ[N�dхĉ� �����I4]q��P��8
$b�TS�I�j��I�5�A� ��܅0�cL�*��� |�#<�`0�	�O�TaAFS���bK�#���t�Ɉ`�X��'�bh	w�N�[�:}X�G��>(ybHJW�'��&�t1�f՗,�<�1�� <dXm�������	(S'�'�����h��OB l,����b���xy��Z@?!�l]?��	��� \w��H�A�
h��'i w�)����;�O���H��b#��KF���Q�6�tD͢>�� �4�"<���5D�ThF�H�_2���A�<)@�� 2  ����C���q�.D�l�#�    �	       m!  �'  .  >3   Ĵ���	����Zv)���P���>��'���qe���OT|#�j�9]ֈ���
�*U��r"O1�4ŋ�/^LPi���0HEfIqJ�O_�����+�\#��i�,IP4�4>z�Qv��:\m6�1�I�Sg�-e��4MD`ri�i�rA���o�B���I�^p8���O�f�Q櫁�d��k�}�"�Xu��s���*_V0d�2#ښ!=���$�89�]ەNL&M^q�&GD���	��	ßభ�:������q�de�1a�v���l\y�)ߍO��q�2�'ˆV:)4��a%t(ՙ�oR.�:m�QE\[08q�ۜ���'F�Ƞ� 	Z���"�����Z���񖂍�)Ŗo�ğ8�A�ڟйܴ)��<����~��W�1���IhV4�vM"�ɳ�y�O�qmV� iT'ޜ�2� �M��qsV���FyL�O�}(W�+C3��C���`;��yռ�����?����?�`��`�d�O��%�z8�[��>Ղԣ�0�� �i�-M����S�߶x=�b����O��k�Fd�|�{!��TB h�@��0k�-;%���@�B Go�bs�3b�jz1h!��B3b��-A$C�6b_� Þ�%�Z6m�æ���yR�')�O��W/X\���It��P�� Y�0B�	�3I��	f�m��)զ؁��(��	zy"���B��7��OB�d�?���/ם^<�4�� >����r�}�6!	��O|�d�Oj�f��P���!mK�w�l�m��F�:%�I�@��:tP�X2�m�'��x�Ah�`t��2/� T~����I`Ս]9N���)	BTH̥ ��	�s��D�OJ�o�꟨��$ �Q+��9s"��p�n� �v����9�i>uGyF?)���r�]1/���
q��M���?y�ʟ�x�'5�p�D�Ɋ�R�bĨ�Y�pYg(�>A�	J9B����'��'��D+G:Yb�'t�� �C�cQ��S�L��-��mj��)a���O���?A/��O2��`��n2x���ؗn��y���'�"4yed�-{�Z��E�ѝ=��?��S,ڕ1#�9���7P����ȅ�H3��OZqo9��T>�Ss�t勳[:��SQ�T�,�����ww����I؟H�}�qjSu��J�r��)3��W��?QZ� �'S�> ������8/:�@����<:-�Ȓڴ�?)�?4p[�����?i���?q��}u�n�O@�F�T�MRRp:s��2L��Ѓ�ڈ^�����3�&���F-�`	��(OD�ٷAԭSv����X2x��`Ps��J|��%XsP��d+	�6�3�]Ĥ�wȌtC� s��~�t�'i�y��?����'�	׫x���q䫎 F܂�����l[!�Ē�tYP �3�Da�hPGm�+7Q�f�4��|���������a�	%Y��`���=D���Rcɒq����O����O�����?����į��DN�ĺ'o�-/��\�����~�P��6�׍Yv���@�Oqxȣ��(�yцh�S��T�y�u%�iK41���D�O� ɤJ۞l"�T��]�p��`"���Od��%�)g�%±fUL�bZ��Ʀ�G{��ɅS\�8q��:zA慹'��m��C�Ix��ztB%/��B�s������'��3��p��J�D�?�Zŀ�F��P���� [�XHvCo�B���H�O��d�ON���	��hI�A�A-h�ԟ�R@C@=_�����A��S�ؙA�ɕZ��`qS-��'4���d��� B��Bi�
���<@�Ņ�hO�=�@�'n�6M�@�'="�	p��'h�9g�ھ0����'�R�'��%ӵ�>R ��+�It���
�Dm�ɟlS&a��iD�k���i�eϥp�j�lc�\B"G�;���V�G�	Ӱ�GzB���=ת�K5B���HjaE*�y��U�֝��A�|-�Tۅד�yBRb9S�B%&��vgͦ�yr#ψ`:���wH@�T�Е�yR�'�	�n�P��)�(��y�b�#�L1v	T">+�e˵ᒱ�y���B)IGa�h4B��	�y"/(5�bh
��O�C�K4E��y2FZ{FhKB([�;��� �"�y"Ƙ�V�B���fP`�H��Tb@�yrI�0�ޕ�JݘNF¨xdh���y"��<B�E��b		^�T ��]"�yb�D<%쾕I�m�:���MC
�Py��8j"�z�F�-*�`��u�<���c�����0b�n�8�]N�<�Ь	$���:�a�&s�h�j�F�<� ��j�H切�0�6Y`�ďC�<ɤo��w5��0�ߵ/Ң𳤘_�<Y�*���9J�À�x�`��B\@�<� �\0#�/dhlh �>SgE��-�3p��C$�Ζ&b��2w�i?>#|J]�<�$�V1��%��L�@�X4
��1D�
rI�14H R���k#$yӮ�2�f�)� ��ɆP-$*�	�]�H�Ђ#Z�̹�"a�qm,�����J�\d��ၨ���cGΎ� ��P ��\)J���x�-�lh�� U؟P�󃅯3�y�Mۼ5�m���3�ɬ?"m���5��;Q��'�47��d�L*Q���ABG(a  UŧJ�y�AE�Q�&��T�]%#�@y�D�BG\�tWi
�o�\T1t���M���?�sS���?Q��O\m�.A'����cYv%��'�v$��Ŷa�l� �7V"U�΂�L�� !�i  �ĮK�j�RYQ�M���Q���H '��%��&�;m����Ì�O�Q�����X gh�$��.�+M�j�	�Ǆ�o�s�
��Ri��0P�X�2�
S-X��@Y+�BS@؟��" ���с�ޟmW���Ic�@��(�~������B#y��i�	L8
@r��W���s���o�� n�p7*[L.�Uq�a D��@�
ߡF�@�h�"��=��<����pkFܸv�2y��f�����O$@�j�*��}-�=��O��Z�)P
Q�&q�6|����'��HP��9���7_��s�ütL�	���ɾ68 xr�����J�`��z��j��7��Onh�@Y�@wP�l\�O8=��$ՇBrK��@J2��
�� ��|+��0,w�����1��BnC�@�S�4>���-(�O(L�#�!@.�=����+�@�����2 �U�':���g�H�PP�"�Oc�ܔz�����6m�Q�4��& "!�'�R7-��:5++D�0@u���������w"#t�@C6��/X�Pm���������x��&t�4u�3B�>�ǅ_1-� ��ȷr���2�]\8�0���� 6��p�SdȽO�~��@dD�g���z ��*)��� �G�/��zĮ��'����o�]�'+F�q֫إz@�1[�B�}R���d?'=�\�l
�5�tpY�#�^k��pT���Î0�Q�J+gC\�h�MPkU��Y3� �O��v-\��#�BRa�<O���q�^q�n�"�(�`�L�t=|�h!�]�S�X�*q[t,Q�Tk�I�4x>B�Ix���׫Oz\t�>`�3"����׫N�hA�Y	pc�S�ft��.i��1*�O���P��M�f��q
B
�4ب��')4٪�M^�N%R�`�\^"ؑH3O2g뾽��*ͺAVJ��'���p$r���+(�R�F~� ��n�L����1H�@uUhЄ�HO&MQ��\�?�w��cຈ+6l�$%Ltj�F�ސ�ʝ"G[PL�wA��vX�t���'�V�J ���iɒ��w"��{W�� cU�D�|X���'gȸu��!�ִK"ğ�I����t��w`�`Ĭ�W���Ö�u M��'�:D�c��
k
��rvDCC�K\F Y����1J9��(ݴH(��� 0+��2D-�����T�H�G�]�q��](�a�.��!��'�O�q{�9�$�mywF��� � "tR`�V�w��6��8����"��tSb�^�W�J`���dSZ̩�e�]?*M䘒�Lӷ/#�h��mԆ^4�Q���G(y-I�p��rDL����#!�d֎z��,�� &T�~4F
�7�V'�%�`�|���i��a���v���
tdU5&��y��'�8�afO݉~]�p�o��\�2r�O��1�/|O\u�ELI�#3��r���)�0��"O���e@�c�@�W�`��"O挻�&M)C�8�!ᇟ<)U�ā"O�,�ǂº6���� �%d���y"��nP��m��.z��������yr�B�d��Q���+!��aѡ쑓�yB`��L�L���,L�e}z%	���yRd��H�ѩ�,<�`����y��_W�X��ƀח���eCG:Y�!�M�[x� gΈ)5W*Җ�@�H�!�d�xLʑ����Lg�@[��� [�!�D�>@�Qp#�U�d��*��!��8��H��V ���f���{�!�$�<��q N�_��A�L�v�!��S%o�S�G��0� *�hS��!��e{
D���Z�S���BC/�!��2t����Vl�m�J���қ6!��L=�T�E!�f��@'� r"!�䔌9�ȴau(Snڠ���T�A!�ǚ<V�P��ˎ.fL���'R#Mh!����\�U��)QM�x�u��G]!�� j�8eX�*9�l�p��$#V.��&"OV�$J�$YU�<�q��4y�P�"O��7��aN���X�j�c0"O��bg�0�p��l?#պ���"O��e`��y�F\+eͮb6vy3S"O�	s�d��ԉ?+"d��"Oz�����]�u�%k�7���آ"O Tb��E�t�`r6*ע	�>��"O�eC�ɒ�z�r�Jw��'REA�"O����&�'y�@K�HԡW&B��"O�q:�mЇI��%P"�Ëf& ���"O%��f
�!�H���>'
)�"O8�ъ=��`DKJ;E�q�"OV :���a���'�}��"O�u:≚6�ލɅ�p�(� 6"OR���_�rqCFћ'Ot@@""O���VjTw����n�
 A���"O��c�� n($|��\�BxQ]6��O*�}�>d�,�UGI�Rx�m1�J�{��t�ȓ{ �Zp,Z��i�Ui�]hL(�EG����'�Ja��f&�Q���[4CA�ד3����@����VANb�l�J[�)�"�%�B�I�#��Q�C
J����*���O�����
Zy�u9Fd�J�O���� o
Ta"�2dEr�	�'�Eâ�#I(�9�鏁\Ӣ0S�BAp��<��j�O��1%���� �D"��T�Ln2�;��߇/�����P�;�J)� �O�P7:����L U н����KR��	q�'�{�²�O���a�p�@�����U��D*�[��Աf���b�C]�2�m���[�y?�B�I9(3�!y����g<b< �-؝Q|�Ox�zD&K�{���(mdo<9F�dg����Rf�H*%�B�0�:�y�.�tg��*Z� �qĉ��mBqHsnQ� ��a�?h��L~�y&�����3F���HY�pR%L��?! .��B���a�@��Y�@�9�.Ep��Y]F> ��J� ��w�'��,u��0��|z�Iul2�b��$ĽB��݀��=�԰ˠ��~�B��CcK����T�ވ���Y1=)L��� 8&� ��yS���h�:
V9�'��L[�R�j(9Z��	pIs�t��WcLI��"��Jt��3�D<��O�
�
���x�����l����� ���`����"jӐl�F+�?��~8�'X�� 7�P�+?�`�	�4���M؀��A;mQ���'�Q�W�,eu��yo��-O9�Dz�B�g�y"�N�p����êb��•L'��Oz��3c[�O+�|�w��r��נ�/a�T�r@�v	R��4��.�TB�ɄlM�1卑����ـ|
�9���a+
�A������ |&�0D��@�h�l�2�uۘM����/�y�$�J�@����:h���S�A�a�P�JX���)���|�<�0��<T�H�ɰ[P:Y��OW�<�D#C^,��Tj��J�����ȃ֦�a`��%4J��P��v���k���AvfM�daI)lOέ§��l�`!�Ӽi�(��q�I�`mjAhe��W�T z�'��-�$A߃_ �A &�e[�{�A��,��f	�h���G@�Z0��H?��u"O���Br�q!�S�dp�d��o8��"�xr�<�g}��ەk���Q�L�c��H�rݮ�y��S�a�.x³�D=3�D����:4B�|{N��d�=yd	�ŎV�V)­q%�-o;�{�*�:Q��I
�)� 62Q�h�4�C�	�;����Ŋ�܁��լ?�$C䉯#�H��ea.	��Hsa�<S/$C�I�- ��7�F�vw�䐶��,i�B�	3��d�Ɔ:K�T���T$)�B�I�6Jvɑ��Iw�d��7|�B�IX�>�B�1@p�3���Ii�B�ɤjD�(�g�:T'&�ޜ.�B�)� �q�s�QO"Ց��^�7 �p�"O`�Bc�U	rʈ�ABg��Qe6i1�"O�s�(�N<ԡF(׶!���+p"O�*�`�	.�����(J>�Bݳ�"O�m�Q��%T� �&� ?�(��"O�\1��%Lx����b38�lR"O�]�f���l��#LU�*M�P"OLē��}#�܀`L\HܺB"O><B�Bч����!@�+kB0!"O�pC�C�,�4�ɑ/�'�<�r%"O�L�b�Q�$� A1daP�R���"Op�0C��M����(3���"O�l��Q�eI��2eG���0"O�*Ó,9!���c�;_B©�p"O �"��43���D'�z����"O:��5�E�j�ti���ӑ$�zh��"O�
��T�Y�|�Rs^M�.�:�"Oʰ�G���ږ��8j� P9�"Ol�0��F�.e���	��qP�"Oq`�FRo�<i6)�?��y�6"Ob��3I�������;����LW�q �[|z  �1O��܆ȓ7�� !'Q#M*�Hu�^
#�I��G3��tn�%"���sSf��1�<�ȓF��i��g�~Ũ��{���ȓ�ެ���Ů2i>�KV�ٚń�]:���-a�x��`DV�pp�� h�h�A�-6��#�h@�S�]���A�U9�rY�7�("��ȓ4�>=I�kI"�dx4	+xǶd��D �أ3�G)y6 0@PO�I����cf���!蓉,�ΐ	s�׭``L���h�8���W�:��R#�^�R�؆ȓn�hؐ��o �Ś�EM�dl�(�ȓ}  �P6C�?���&��#
�6a��ӢP&ݣGR:�iҦV�^� �ȓ?���0�G[�/�����z�숆ȓ<p���5eH:/w�Ys�̉� ��ĆȓC�\H$�0#�r}���/����ȓ�F��aFE�OP��ecʲ3)�@�ȓFo0!�WmFm�x�2L4E~5��wz���#O��0 .[�{�܅�sUB�b�T}"�GJ(2
��g���c`�U�LsƝ�	�N�t���9L�dI��wU
�P���	;�2�ȓ
K�����z������� ���tz�)�%[�W�>E�En�_�Q�ȓ[9��eM��rH v�Ƨ;����ZU@x��dy~-�%�	GHN��'�X���l�<Q��8Cp��
`�tb��ě6=�,EH"�@�(06��aDP�!�Ĕ+ZV��ĭQ�b��Т��Ԛ_}!�	�M�:��$���!����L�e!�$�>����'�I�RQz殈�U%!�DQ� �	�0Jn��y�-ն!�N=�8���6����uk�(N�!��Դ��i8F,֞%��ꃠ�y�!�D�d`)�'�O�$!B\�P�!�A�2�4ړ�	�|1�4��W3!��ƛL�>�tK�&6�*xB*ė%G!�Ċb�8���S�tySW��&-!��*�BQ��/B�qۥ��(!���ՠ��!�Mcr�!�p���4!�ٻ^Y���L�4d�0,V�g�!�L�pLh&J
ZQ������P�!�� �(s�.B蠕��a�lT�!"O�Di!BR�0w��hB➂sT0�1"O*5�F�ژB!VHӔ�F�|fnMb "O��	����@<hs�W LW��J�"On𒖯��hԖ{4aT�s��PV"O�,��cV7
�+�J�<x�<��"OV���. �pp��j@j.+\T��6"O�8F�j��0+!#�8	�& �&"OB���^h�\�â�HV"O��XC$�7�eyE� x���ib"O���ID*@�n��bͧj���"O�����	��� ��D��qI�"O\��a�!il�Y���=�:���"O��2TMJ�|3n�h��ݨ��g"O���G��k��-�ciZ%��tK�"O��C2�ڗqa��)WSʐ��"O4��"�u�f�V�Ѡ)�vӒ"O�`� �c�2��)UXwDɣU"O��ȑ��G����Ygr�#a"O�\�C���Z�� H @|��.�!�DRt?bM#aJ,1��Lx��M�!�$�
t�<K"�S5f�9�FE�?�!�DU�~��r���+8�� ���#=2!��<1�n�P�ŶP�c�E4_7!�D������Z'����!\�!���J��a�fLJ|�>�1U���!�D��f>(�&�� ���q�!���pH�"#���#ӿyO�ȓ%E�`��oJ�����\�[����@���
�lG�g�q[�-W�`z�E�ȓ �Ax�%�Bb};ƧU94_>��ȓnM��jC�2,�ITG�~Zhl�ȓM{�=�PӉ<2���S�1v�ȓl'Xh�U��_�z��ӌ�D�и��J�呥D>b.h;��W=T��̅ȓi̍���I�$�4c�ʷ�B剭9HK	; 2<��M&�Z�f"O"�/�L�Ul x��'@�l�C�Ɂt_8C�l'^زa!1O«FٚC�ɉP��Ѩ��u�!*���f/JC�	98�U{�mU�x�n9rg�+�C��2H�Đ����:V9��%ч��B�I>W(t����f�$��f� �B�	�d�.0��1?^i��
�K4B�	\�^4��)[*e�J!R��(;�C�IV�Bǀ-i3>���NEY�B�nj�A�ʻ#\�x"� �TC䉅iT��%�<� ��r��yNC��\Qn�{�K:E��\����N�B�Ɂ �����\�0�|�g�^�u޸B�	�>�*�h+'�`�B�_�^��B�ɹ��9��h�>f�P�b%k\�&��C�I1<��e���Z�Ia�rE		�HB��,j��uZ��^�?�Ԣ�"�eFB�I5?cD��)U!"*�<�9�nB�I8tJ��ʖ�U�C�T�җe��
�BB�ɗ,�(��E;l.􂄂�j�B�	�^`��!���L��B,?T�C�I"l�bA��m�����QBD�]��C䉱�6�����V#�ZcK]k��B�ɌrZ�P8�@���u�$��|B�		'���i�L��e�`9�vi�(��C�	�w#)�P�:հV	Ç^KB�(��f\r���$�.��C�)� �<�'��!8��9ňA5��#f"OF��pC��4G�M:���f�Y�4"O���P��5|Pܩ�AP�s�� �"OdP�#�Q;Sr$ŨS-WR�@#�"OD�C�����[#��X��mK�"O0�5DF7�Z�r��	�(�����"O~�`"��1L���˧Z9�D��"O@L�F$�61F�Шg�-#<P�b"OV��Q�3����속Q"��'"O��9���SX� !.Z����"O�='��Xe �̋<~h8e"O�E1�)�*f�IR)��~V�D�"O�Z@�\�sx<���fB��s�"O��A��6*��qg��8e9�PXd"O��&��q���1W.Ʊ4z�`�"OfdXC��x<I��=gr���"O���֬ў3��H�2g�W�D�"O��[��+�JU�0'�8E�P� "O�m�RJ�h�!�Խin�j�"O�x:E�:;��sV�ޕk�]��"Ol��ѿn7�@z$��.s���"O&��b��Y�%�T�A�@M*�b"O4�v(Խ#��(�d��?�e"OZ4:�#7!��2-Lip�"O�� �Q$f��T�_�/,F�0��'��'�t�Hg�LP��}�E+L�9~}��'g�}��d�'���	��ʉ�f]��'�l\��L�aZX�QC����	�'��Q�Iy��Kb�Յ;�=#	�'��=(���)����!�_�GJ��'T�͛�dR7W$�<�D�W�;H�'������?C(	��b� ^#���'�H��ѨA��eP��& ~U`�'
����K�x��QMނh���*
�'��=��΋J��F��n����	�'���jց�#S�EaU��t���$��%�OXq:��N vY���E� \����P"O�t���Œ_��h��=F��"O������NHl8+qC��tL^4��"OT�K��G3g�����U�d�F"Oz���]?�P�r��(a�m���	�HO�6p>�H�`�7F8�|�çM%?#�B�I0LQ��JGeS�d��JB.��I��6�%�S��M��AK�a�t�[U�Z�)�����N�<�c�M��Ie�ĩ�"���	K?�F�'��|8��H*N1!�1��9	�'kx0��K>,(�!p�ń-à��ʓ+��� A�9���1f[�QLP��ȓl�"xq��(M$d�P��C�B��X�ȓmw�!`��"���5��5=�,ԆȓE��x�% ���$x��*�-�&��ȓM����$�U��hk7@6	�h�ȓc��=�cH�-Xt$Hm(�ȓ\�`�P�M��pċ�Ӿ��l��/\>�s�0M����e�ws� ��%��1��]�İ��
P)9:Έ�ȓ`�V=:b!�w�Tm:ǐ!nC@���y+j��0⏂z=�8jX�0��5�ȓ�>\�7���&�i�Ɲ�t�@\�ȓ9��B�n�P72����	*��݅���m*'E��2��@S �,�Ԥ��a'6E1wG�=1�E����(\F���74��3�K�1(� }j�F�"J��ȓo����AV|W�Z�d�U52\��S�? �!ʂ�̉;��,SwaA Aj.q�"O(y
��Dg����v	�!5"O�H��Ԭd�iq�"Q��a0"O�=�L!q��`���P�$�0���"O���DV���H`�����;�"O|�!UcZL;ƌ�%#ݝa���"O81kEV:�x�AtAˤ=�x�"�"O�!e�ϝX�$*4�_�f�&�1�"OJ��5苖)�x,9`-�"x��QJ�"O2�b�HC���F �#h����"O���3h۸H���R�J�>R<xv"Op�sq�>J�Z|	��Q#9Q�И@"O>1�J6!�M�4g�K3T�K�"O��(%A�0+�Z�����||ʅ"O씪��T+ M�9r��q�,
�"O��0��^�h#�F�!��"OZY+�Z�	>4Q&�O�a"��"OhAW+P�b�М2iT4e����t"O��d��%2��R���r�	�"OU�҉8!;|qIWgS����"Ol\�g/�"r���+sd�	0Q�"O^�٣b]3~�=!�C�LV��d"Oz,��O�d_&x�(��bKz1�"Ob��rj�8�%D��+�"Oz��4ჍP��A�᪃.,�6��%"ONĂ���k4���O
y�6d�r"Ox���ⓝT���#_=��!��"O6t(2��\萕��	�+!�~��"O��r�)4���i��ޑ_)��2"Orm���KB�U�Q��	B�A��"O����-#�j�z�@�"?2({e"OE!E)�*%�ȍ�յxZE��"O����#4�X32�Ěv]�ɉG"O(b�нJ�rt�r�&O6�*U"O�:�@�U�`���L�=d�T@�"O�܁��Y**�����N3�Ĩ�"O��s%�#������0(Z��D"O<��b+G�VEb���}p�m��"O��K!BJ��$xR��C�E�0"O�Q$�]-Mz����� #�8q �"O�	'H�bL�r�P�n�j�"Ov%h��-�-��o:��6�3D��3!K�3.�^��t��B���d�3D��:ևM�(I8R�ɺa�� ��=D���4�݀��U��+}��h�!:D��
`C\�A�1����=CSg7D�DI�Ւ�م�}�ʹR��0D�p�� A/~�R]A��;_��5�0�*D�p�bj ���y�e�D�y��8��$'D��"�d�;����#GΦ�ʣ($D�@zVM�eR�t3@4u�u� A"D�T Ԃ�)^~t��K�8�Ni5�2D�H���;u���1�
�*=xC�F%D��   �   j   Ĵ���	��Z�tI�.ʜ�cd�<��k٥���qe�H�4M��\70<i���:G�&�����0E�5��y��cA�6-Ħ�q�4x��$"�	}yr��2�p�Y`f�lٖ�&�H�܋'왭e�a�=��,)�=`6�ĺ)Π9Q�$�x��)xׯ;w<�ɋI�q�ǩ�{���(�8YvN �q�	 ��U	"�$q�Pa�� �`����[$��͔9,�%�	�Q��`�d�?q��'�0�%ڱ��E�*ߓU���p/�EdUI��A�����d	*3�i��! @9OT��U.
e,�ɏ]�����b�&�FŉrP�G����d�����Au���t�nY�t�P(H����OF�����BTƕ+u�ҸuG=kՀY�[H�a"@\�Ƹ'0�Gxrk7�YP"F�]�CF�p�p��	�*���a�Z��h�����ڔ�290�x;�6}B&V�'C�X�=�SDZ��`�W�\&0��bb���b�ቮ^���%dV����!�c�(��Z	L�Bc����A(��NFM8�%=o��*E�)v� �'�B"<�d!���2,<��-F�+U�"���*>"4(ቻ��s'�'즥���Gb:}���HW|I��y��y�'�~�'�xa�ժ�r�ϼ@�(@T� <�~���k�'��M$��s�'���Be�1]�X$��*�/F���C�+h�ɄU��	��i�M��Kp�dņ�I�ɠfQ���s�O���'��Fx�
b�DN� n<�2�� C6��d,�I�@��`���I��0���E�W)��a���	dQlC��5>�� �  �&4D��ic�OZ&�g�{K���"�3D��2�g�*�~|���'�Xyw�.D�|Hb�	;_��dy3c��W�@��4,D���n�����[	T�9`���ybO�5V�y L�1&��;T+�(�y�B�2�`�F�_�.H� �#�y� C7)��q'�\�(ke���y�l´uB�5I����X�H�HMJ�y�MZ�E%R�RþP���¦R��J�'������=�\I"�iĞ���Y�'�|�T�K&��I�Q�� ���Z
�'�N�E� �� [�@�H��)	�'��C��W�l,��瑄\�����'U�5A���o�C�F]�i�8py
�'j"��`��%:p(Yǋކw��$��'H:)��ω?��j6���i�4��'ðĠ��M�F�Q�Ի�    �	     (  �!  �'  .  W3   Ĵ���	����Zv)���P���>��'���qe���OT|#�j�9]ֈ���
�*U��r"O1�4ŋ�/^LPi���0HEfIqJ�O_�����+�\#��i�,IP4�4>z�Qv��:\m6�1�I�Sg�-e��4MD`ri�i�rA���o�B���I�^p8���O�f�Q櫁�d��k�}�"�Xu��s���*_V0d�2#ښ!=���$�89�]ەNL&M^q�&GD���	��	ßభ�:������q�de�1a�v���l\y�)ߍO��q�2�'ˆV:)4��a%t(ՙ�oR.�:m�QE\[08q�ۜ���'F�Ƞ� 	Z���"�����Z���񖂍�)Ŗo�ğ8�A�ڟйܴ)��<����~��W�1���IhV4�vM"�ɳ�y�O�qmV� iT'ޜ�2� �M��qsV���FyL�O�}(W�+C3��C���`;��yռ�����?����?�`��`�d�O��%�z8�[��>Ղԣ�0�� �i�-M����S�߶x=�b����O��k�Fd�|�{!��TB h�@��0k�-;%���@�B Go�bs�3b�jz1h!��B3b��-A$C�6b_� Þ�%�Z6m�æ���yR�')�O��W/X\���It��P�� Y�0B�	�3I��	f�m��)զ؁��(��	zy"���B��7��OB�d�?���/ם^<�4�� >����r�}�6!	��O|�d�Oj�f��P���!mK�w�l�m��F�:%�I�@��:tP�X2�m�'��x�Ah�`t��2/� T~����I`Ս]9N���)	BTH̥ ��	�s��D�OJ�o�꟨��$ �Q+��9s"��p�n� �v����9�i>uGyF?)���r�]1/���
q��M���?y�ʟ�x�'5�p�D�Ɋ�R�bĨ�Y�pYg(�>A�	J9B����'��'��D+G:Yb�'t�� �C�cQ��S�L��-��mj��)a���O���?A/��O2��`��n2x���ؗn��y���'�"4yed�-{�Z��E�ѝ=��?��S,ڕ1#�9���7P����ȅ�H3��OZqo9��T>�Ss�t勳[:��SQ�T�,�����ww����I؟H�}�qjSu��J�r��)3��W��?QZ� �'S�> ������8/:�@����<:-�Ȓڴ�?)�?4p[�����?i���?q��}u�n�O@�F�T�MRRp:s��2L��Ѓ�ڈ^�����3�&���F-�`	��(OD�ٷAԭSv����X2x��`Ps��J|��%XsP��d+	�6�3�]Ĥ�wȌtC� s��~�t�'i�y��?����'�	׫x���q䫎 F܂�����l[!�Ē�tYP �3�Da�hPGm�+7Q�f�4��|���������a�	%Y��`���=D���Rcɒq����O����O�����?����į��DN�ĺ'o�-/��\�����~�P��6�׍Yv���@�Oqxȣ��(�yцh�S��T�y�u%�iK41���D�O� ɤJ۞l"�T��]�p��`"���Od��%�)g�%±fUL�bZ��Ʀ�G{��ɅS\�8q��:zA慹'��m��C�Ix��ztB%/��B�s������'��3��p��J�D�?�Zŀ�F��P���� [�XHvCo�B���H�O��d�ON���	��hI�A�A-h�ԟ�R@C@=_�����A��S�ؙA�ɕZ��`qS-��'4���d��� B��Bi�
���<@�Ņ�hO�=�@�'n�6M�@�'="�	p��'h�9g�ھ0����'�R�'��%ӵ�>R ��+�It���
�Dm�ɟlS&a��iD�k���i�eϥp�j�lc�\B"G�;���V�G�	Ӱ�GzB���=ת�K5B���HjaE*�y��U�֝��A�|-�Tۅד�yBRb9S�B%&��vgͦ�yr#ψ`:���wH@�T�Е�yR�'�	�n�P��)�(��y�b�#�L1v	T">+�e˵ᒱ�y���B)IGa�h4B��	�y"/(5�bh
��O�C�K4E��y2FZ{FhKB([�;��� �"�y"Ƙ�V�B���fP`�H��Tb@�yrI�0�ޕ�JݘNF¨xdh���y"��<B�E��b		^�T ��]"�yb�D<%쾕I�m�:���MC
�Py��8j"�z�F�-*�`��u�<���c�����0b�n�8�]N�<�Ь	$���:�a�&s�h�j�F�<� ��j�H切�0�6Y`�ďC�<ɤo��w5��0�ߵ/Ң𳤘_�<Y�*���9J�À�x�`��B\@�<� �\0#�/dhlh �>SgE��-�3p��C$�Ζ&b��2w�i?>#|J]�<�$�V1��%��L�@�X4
��1D�
rI�14H R���k#$yӮ�2�f�)� ��ɆP-$*�	�]�H�Ђ#Z�̹�"a�qm,�����J�\d��ၨ���cGΎ� ��P ��\)J���x�-�lh�� U؟P�󃅯3�y�Mۼ5�m���3�ɬ?"m���5��;Q��'�47��d�L*Q���ABG(a  UŧJ�y�AE�Q�&��T�]%#�@y�D�BG\�tWi
�o�\T1t���M���?�sS���?Q��O\m�.A'����cYv%��'�v$��Ŷa�l� �7V"U�΂�L�� !�i  �ĮK�j�RYQ�M���Q���H '��%��&�;m����Ì�O�Q�����X gh�$��.�+M�j�	�Ǆ�o�s�
��Ri��0P�X�2�
S-X��@Y+�BS@؟��" ���с�ޟmW���Ic�@��(�~������B#y��i�	L8
@r��W���s���o�� n�p7*[L.�Uq�a D��@�
ߡF�@�h�"��=��<����pkFܸv�2y��f�����O$@�j�*��}-�=��O��Z�)P
Q�&q�6|����'��HP��9���7_��s�ütL�	���ɾ68 xr�����J�`��z��j��7��Onh�@Y�@wP�l\�O8=��$ՇBrK��@J2��
�� ��|+��0,w�����1��BnC�@�S�4>���-(�O(L�#�!@.�=����+�@�����2 �U�':���g�H�PP�"�Oc�ܔz�����6m�Q�4��& "!�'�R7-��:5++D�0@u���������w"#t�@C6��/X�Pm���������x��&t�4u�3B�>�ǅ_1-� ��ȷr���2�]\8�0���� 6��p�SdȽO�~��@dD�g���z ��*)��� �G�/��zĮ��'����o�]�'+F�q֫إz@�1[�B�}R���d?'=�\�l
�5�tpY�#�^k��pT���Î0�Q�J+gC\�h�MPkU��Y3� �O��v-\��#�BRa�<O���q�^q�n�"�(�`�L�t=|�h!�]�S�X�*q[t,Q�Tk�I�4x>B�Ix���׫Oz\t�>`�3"����׫N�hA�Y	pc�S�ft��.i��1*�O���P��M�f��q
B
�4ب��')4٪�M^�N%R�`�\^"ؑH3O2g뾽��*ͺAVJ��'���p$r���+(�R�F~� ��n�L����1H�@uUhЄ�HO&MQ��\�?�w��cຈ+6l�$%Ltj�F�ސ�ʝ"G[PL�wA��vX�t���'�V�J ���iɒ��w"��{W�� cU�D�|X���'gȸu��!�ִK"ğ�I����t��w`�`Ĭ�W���Ö�u M��'�:D�c��
k
��rvDCC�K\F Y����1J9��(ݴH(��� 0+��2D-�����T�H�G�]�q��](�a�.��!��'�O�q{�9�$�mywF��� � "tR`�V�w��6��8����"��tSb�^�W�J`���dSZ̩�e�]?*M䘒�Lӷ/#�h��mԆ^4�Q���G(y-I�p��rDL����#!�d֎z��,�� &T�~4F
�7�V'�%�`�|���i��a���v���
tdU5&��y��'�8�afO݉~]�p�o��\�2r�O��1�/|O\u�ELI�#3��r���)�0��"O���e@�c�@�W�`��"O挻�&M)C�8�!ᇟ<)U�ā"O�,�ǂº6���� �%d���y"��nP��m��.z��������yr�B�d��Q���+!��aѡ쑓�yB`��L�L���,L�e}z%	���yRd��H�ѩ�,<�`����y��_W�X��ƀח���eCG:Y�!�M�[x� gΈ)5W*Җ�@�H�!�d�xLʑ����Lg�@[��� [�!�D�>@�Qp#�U�d��*��!��8��H��V ���f���{�!�$�<��q N�_��A�L�v�!��S%o�S�G��0� *�hS��!��e{
D���Z�S���BC/�!��2t����Vl�m�J���қ6!��L=�T�E!�f��@'� r"!�䔌9�ȴau(Snڠ���T�A!�ǚ<V�P��ˎ.fL���'R#Mh!����\�U��)QM�x�u��G]!�� j�8eX�*9�l�p��$#V.��&"OV�$J�$YU�<�q��4y�P�"O��7��aN���X�j�c0"O��bg�0�p��l?#պ���"O��e`��y�F\+eͮb6vy3S"O�	s�d��ԉ?+"d��"Oz�����]�u�%k�7���آ"O Tb��E�t�`r6*ע	�>��"O�eC�ɒ�z�r�Jw��'REA�"O����&�'y�@K�HԡW&B��"O�q:�mЇI��%P"�Ëf& ���"O%��f
�!�H���>'
)�"O8�ъ=��`DKJ;E�q�"OV :���a���'�}��"O�u:≚6�ލɅ�p�(� 6"OR���_�rqCFћ'Ot@@"��.H�$���J#s�Yi4�G�uaN�25M�@�!�$��pD��Q���N/��z4
�J9	Cl�|�	�
�Q>�4���",S90�F� sAN�hͅ�Ax�H�Z�j�v-F�o������DH�dcԥH���&�U��\5���B$'�H����>\O�)��Y�"���'�Hh��VW�	)��&`�$��'�����j�x7�E���Ex��+N�$��e$D�]�S45WT�G��q�p=0CdP��� _�y�g�������mI�k~�x��닝�F�h��Z��$��=��;��L>၎�ͮ@��+�26r~�`�Da<ᅆ�6���8"'� {�1�dpԴ���c�r��o1ɶ��������G B��<)&��J�ax�-M� ��@�Y�pi�T@�o�'��4����D-��{I*Pj�'�քsaI�f�6�E��r)�V�<ic�0�:}"�
"kօqiY�����KjZ5 *�
#JԵ�PQ�v"O�9&"���i��#�tmV �w�α#����%���{<�MB�n0<��O�1O���f�=Qy�$�,����!�'r����|{���v,
+c�����9�q³/��,G��0"*1����D�Y��ؤq:� ���Y�k�џx��j�0������'�`�2J��kǀ��+��zA�M	rGX�pϦ�
�'�2*R�W���ݲ %ִg�Tm�,O2 s��S��P�m��L�U����Of���CӔ��C�-Y�k� �'��0��H������ĉ-s�<u�� :䰛5�_˦9�aƋ�n��OT��O"�)gÂ�C���ڐ�To�YS��'�"�+cˍ�J���Y0E�6i�:b�
K5�	�@b_�E�i�%�����D�,,���&�� TI �&PџX�sdD+,dQ�&
@A�A�&��b�ltX��}�xyC@�E9x����b}�Q��JV	h�S$	�8,:���',Ѫ�@�1�t͑C�j1�Q����
LH�Pg M'>�f �/��(�!��N�q�&�*�c\�Q�M�b�<+p��g�b���1/�T?����y�-����};#��t�I�#@Ƹ�y��ő;w�|I�.�)3��[����M;v�^�o�֤:aN�p=� ƄOO��PA�:FҨ�Ӧ_]؞�zG�X:U����7I|��)E�I�r�8�ض��u�dE;"OR�"R&<��	2&́Z7p c��P�[��3�j1F�>�	@$�3$�TڧME(�,da�l1D����	N�3�@.�<�\sB!ºX�8�1�Rd���^�*���F&�8�xI�q�Z��!��Y�#Ü��D�Q���"�GR:�:6ę������	�3�,���O=�%���Mz:���JJ���_�v|{F�Êr��T9�CCbp��O�P��p���S��e�e�٫l:�����╂D�-XU~ز�a��`�ȓy?�DSFܖZ�Z�*X�p���N�$�[�&ژ ,���)��q��@� �U��?0�x| �㏡^��!�ȓ�bE�k��LQ0g��*���ȓr��0�GB&58�¬��%��S�? cT'�J��X�'C��E#"OR�j�CY&rp|�6����B� �"O���RmK�L�\����'M9�8z�"Obء%`�}��ga��pQ�"O�����09���!swu�"O�yy���JЈ�;D*L=	L�w"O�A���o%�H��+߅l(ԣ�"OJi���m�hd�>�}S�"O4���I�(�DL8�O�.Фݳ@"O8h��N]�0$�16`��|�PU"O|�Ā 7"�iKD�Ć+�Ny�'"O� ��<Y��}aqc�+L�⭩�"O�BǠ�h��1Z��ˈY$:�i1"O}��%�Պt� �,}f�YB"Obe��1\�,)�l��n�⨰"O��jg�R�IZ%���8�f��"O�٨�E Ȝ}y��zR���"O(�@�6b�д���pR�y"O�i�j�X|bF`ե@�0�y@"O`�&��/P&��SM��(m*A��"O�ERí��N��p�0f��N^����"Oڡ���6���'��7d�q"OA�'JI�ڌ��Z�<+<�y�"O�0j���I�vP��,t�,p�"OpZ�%��SW9!�_�JdVyA�"OpYFG�7jhN�j��		8~��B�"O��&FY�,<�qY5��53���0�"O�t�ġ��H̬U:t�W(�r	+�"O L�jA1s�ţa�(�΍��"OV�؅!\�HN08�CQ����V"O�Ăs��r��2 	���891"On����2;� y��K�>[��g"O(	B�K!a�fi���#j�Tx0"O2 J&l���֐�DO7yc`��"O�|���,X'�TX��+.���"O��S&��k�6��0ߝq(�� "Opx���V"'jM��O}"����"O2Ac����#l�P�֥}���8�"O4L����A�b��6a 8�*���"O0`C�U~�]2 ��4���""O��S�蜉&�J��4	ɷa�V�e"OZDH��E�3SިC�*�t� I(�"O�A�pE��w�&�b$I�3����"O���ݾG:��[�iF"z�n�xT"O� ��A�F���� �Fq��"O���F:��Tա8_��!"OR$���ťx����d�:���"O��a��d���z ����1�"O|�1FP�_b�zģG�g`�9�U��[��3>}R<A�ő~j�!�.�Ph��������Y#n(�D�ȓ.��&ۍR�����_+�)�ȓy�� �Wi
dmy�l��A�p�ȓr����Z�GA��Xb�û!ÊՆȓ>u��H�B5=���p�\�;N���0�Mb����[n�P�L�8B�N ��5�бQ@m��c��eAR�¬�ȓ:�F i��[�r���ڒ ӿQ��`�ȓ;jHiB �\>S��pRfl_�@�z8��vR`��W:��ꦪ�11��9��j� !d#P꽙��ԫ��Ԇ�OyP]���B�U\l)x�ʋ�7�t��ȓcN�Ae'#h�Xͣ�ߝ7��X��U�<8��ĸ1�б�琴5����ȓ^=��g��:>vUIv:):���S�? �y0�l�
l\}��d�����"O�$��#�_�D�X� ��o��C "O���d�>A�4��L���Ⴃ"O��X��Ȓ����MWy��I�"O��c`BF�/�6�C�,N�B��(7"Of�[(��\�����T3�ă�"O�01�J�����S���"Oq@�51�sAL��+x��"O�Ȓ!qi������O�֐�p"OV�B��#dr���Q<[���A�"O���Ӌ*o��Z��A-Ra�h0"O����K^�s@���?'w#A"O��IڣD5"踖BR)=ϒ��D"O�| ���ZO ��V'_Pĩ�7"O$��ɉ!bJʐ��ŝM^`�*c"O�u�掅$VŐ��F��ʅ"O�hp����y{�������u**da�"O�1����(t��5���\|�"ODC�*P>�~I2"��K��E:"OʤQ� �c׈XY�j޲'���kT"O\!h�J]L6]J�)�#w��)9�"O�|3�*�c��"�">/m���"Op}�bi\���UƠ�i�"O��K'���C��6m�@�"O&��s��@$��c&�ٖ�`JQ"O8+$���YHv(�!����ؓ"Oތ�F/U2@�J��tcϗ~$Mk�"Oظ	�]����b�Ѐ;J��3F"O(a��M��yv�_�2g��b�"O���7g�69��d���ԝTdp�+ "O��J�D�K(���CkT_E�$�P"ODQɣ��-3��{
��
�5�"O�!���A�zQT������?�\�0"O��w�_�?.<m���\Td�b"O~��C�D�"�����^��B�b"Oz]���kFb����$9��4"O�s�'5x@a󂥘�s+&�"&"O��(����D�T��dB،n�4�%"O,)�vaOHZ���CB��:� �"O0ĩE̓�I���c�=j� (Bg"O�T�6#ެz�4��L�9�|�J6"O�eC��4 ]���+w���3"O�1��D�-�$��5`?[Ui�"O8��-G�r}cs-�$��"OJ�f
� �L�(�ՠ�8�(T"O"�h� �n�NT*���/��,�P"O$�3 U(6S�Ar�Ė,��1 "O�@Y��Z0j�\�X�$g��0�"OĔ���M�%&bY��ڧfZ�!�"O��X���.u(,@� #K�a:b"O�E�`4T=XP8�?.*�q�"O�XY0�ӦaДr�Ò�JT�W"O�Q#ahS/(RzXb�E��TYF"O���˃:��`�`Btcb"O
}A�� n�ܰ��ʃ�.���"Ov)�5 BO�5�R ;t�P"O�J5ɞ�'����.ٜ8k��x"O��J�� +����.u8��c"O�9k �2N�Պ�a�RW��F"O�5P��P�MZT����N4�Qp"O�:�(%'t% �@����"Oʍ{@�L�
 }*@�J&f���"O"xP���Io����ϞL��y�"O�pp�92��Y��Ǿ�
��V"O� ��"��/r#�Q`6���d�@�KQ"O��{�ϔ|%J媧�P�ymei�"OȅK����S���Klj��"O�u���B{W�DP���4l:t@�"O$���&G�b�y���`��"R"O�Th��\�`��|s�b��1Z=ر"O��T�)�TŨ�[,d�Q�"O�+'��]�!�Se�0����"O�d����r��]�f
�?Ld�a"O�X8���"Z�V	S����0�"Of!��*;�1t�Q�z�,9��"O�d:��
6�y���ϳJ�����"O`�2uN	�&k�j�	��9zs"O�\k�b��"��� ���!"Oxt�EI9z�6��؎2��u*S"O��X1g�i�r��4a�0}QS"O��I�+@�c|�mX�� vvT�@"O���WF3F|��n	�p(	�"O�M���D ���V��bSpu�c"OvH�AЗyX�;�c�2���"OjHxg�&�� %��n.��3C"O~	��K¨g�1%M�1X K�"O��aN�8�dp���#.4�"O��D�&i���+rD�=e+h�S&"O*�'�;��j���(T2NQؗ�'��'�4u ��H�(<ja���~p	�'zB8�pjA��A�g�Q�$p�'�b]�Wc��4ѷ��PIf8[�':.�f@��H�V�;�d �HL��B�ay�惊kv^�+�a$'h�ȓl���ro:B�|�c���;$�D0�ȓD�P�����dj�Q��b��M�x��^5z��F+)k�tY��k��20� ��=S^]�qމFԋUa%�H��ȓyT(�!V�&w�̋��#�xć�@�4�bU$L?�����n�����x��'�6yG��[��\�VӌKQ:�h	�'�,h�gȣU%��Q���mF�$��'�t$�7�Ԥs�*9(���e��$��'wtay�I9w8��.�HA�'���/Ң:9ƌr����-�B����Dq����C�8�����6[J� D�3 �!�d�*]������X�\��@��6�)��=����N�8��_S��"#�!D�t����`�ġsa�a���#�����ziΜy�&�;z^�@h !^;{�
m��r�  x��>�^�`a��#9���ʓ}��(IEI
���5P4&��q�|B�ɍW �腵U��9
H�.D�zB��!q�D�g(�$~��Uk7G¿`�:C��<����RG�,�R�Q&6'K�B�VM���
)j&
�0-�8$rC䉘XFZ\y�c[�C�:e(޼g���ȓ�<�b�ȷ?(�1� �Tt���G�t|ai>�1:��W�+-�<�ȓ�hʰb�m�R�������5��?T�zrk 2���ƍ�=)�]�ȓ$&��a I^-t"��w#>\��r���Sn[(zxq�b�TK�V���F��<��ɉ*:V!Ѳ�Cc)�@����%K6d�/����vͅl�29�ȓ5��c� GTU�Ŏ��]��9��Z��Ed
ITU#f�ȓ��$9q�Q�_o���I2���S�? ����)D�H����<��s�"O�HVAǼΆ$b�	�<I*���"O�	G�M�TՆ�(=��:f"O��8B��$/w6\P�D�=~9�$"O�+�8nW����bտ"p�Q"On���-��W�q1Q��4��q�b"O�� *���qe�6��Q"O�X[@����ic� l��M@R"O��"�j�=IA�2eͺn�.�XT"O��ؒg�P<i� Cѐu���G"O��!�ʆ	E�HJ�!��U�`�6"ON�0D�&��9`���~��U�#"O�8���M:y�6�g`��n<3�"O��P�K�ͰL��/\�?19a"O���F��-_��P0�7hj9*"O|�+��$^UL!�D�Q53��H�"O����Z�$+LıW�][���"O�P� 7B:a��/ V��(r�"O$��a�n�8a�����Kn����"O�� %n�W��������m��"O�,ɢj���=IE��˪��S"O�(���©r2�e�]a�"O��ٵ��>�t�����.)�8�*!"O�� LB! �B�;�E�Q�R�"ON@���;YB\��b� V�h��r"O4�0m�ZK��hT��w�����"O�h���{��� �*˴-Nh��p"O�-�O�(��@��.l���v"O�,yCN�V@�H�g���9ΨQ�"O���&�֐��y��fC#�t��"O�J2%5�.� Pe[,�� "OHD9�B�(;H��ƭW���8:�"OV�h$IO?|�Ĕ��Jڸ^��t $"O�5��W/ET���(]R4m[$"O�a��Ԕ&�V�XW��A:nmA&"O�T�-��C�US�`Ϋ<����"O�Ű�*�a�����קF|A��"O�����
�(r�V�3��(w"Obx��J�O�81���~7��[E"Ox�S1G��J��Ƀh�l|��"Oh@�bZ�x���̏h]�9cd"O�\��kĥ~��WkC6`�pق"O�sE�"'?�%�f�ˉe%����"Oĭp�霝A��-����6 "Od�9�H�0:�,�H��k�<�!�d�uTD�j�坊�[r��a%!򄓖J���:ɶ)Dk��+ !�ئ5��*$58�Ƚ���	m�!�dJ q��uZ��_�t� }8w��Q!�$�6Ǩ�1�&����|P��ϫqC!��A>�2U�b [	o�F z.ڭ�!�(D�Rt��a����S�80!��>A.� u'��.�v9�яR06,!�dU�Hg h  �   n   Ĵ���	��Z�Zv�J�(ʜ�cd�<������qe�H�4��S66<��ʄxG�f�َ%� �8�MαmF���򄒻�7����۴ub��=�	Xy�dݰ|N6��#f�%~rN �E^+Wa�:��]9ap	�=���3�l�&6�	o6MhP ��=�r	���G1���Æ��C읏8A�		9�[�H�y�If������`kP��%m�<&���ťR�Y��MN-c�0E��$S��Lj%˱?�I�'�X�06*S�!RHHh�A'$-�$��O1��2r��By��G�FO,�0Fk�O��ϓ&}�|�E���y"�ƭR�#���;>+�!2A �"�~"h0�N����	��I6�ꄹ���5Jv�g\�a�DW��۶O����K&�\�b�H�iu�;�X[�h�a�͊c%���Ϗ�[��y ����O�����^����
^n��U�
�~L>;B�!L��'�f#<Y�D �I�h<ٓ"�� �`i�g�߹�6M���O\���D��
a&%�1 e���RD�ڈ\J`�s����O�!�O���T�	+`�p&��X�����^�����I=vO�O`�E2�.ɰ �I~�U��6�O��;��DI0�?yC�\==���RRHKS�TkDP̓zS#<�T�5��O 4P���\_�A��뛳-�d8�Oʭ�H<��-Z�MK�G��H5�d c�S-pi�ԚG��ßp{�u��
��S��?�2�>���~��d �j/�X��O�UL,�q�d�?�OJ H�x˵˞9���5���*	��μ>ѱ`9}:�#<9���;9�+��ʴw�e)Eȑw�<�qN� 2  ��*�Of��e@�&+�1sN�9U��)��'�� 3w^�yվ�+�h�O�U�#�(-���v�C"�H��"O��S�Vu�tx�e������P�|b���NA��Tm�xun�}�6��_z�{��ѥw|B��@m�J�<�p��D䘲�
�� *V��X*KzIpI�	;.�6M�*W�BI��L>)�f��.6
1tDD����E(<I���5r�Qf�M1(xY�A$���X'O�<�V�������z
� ������9�q%3��I��'�@�b��Q�ka��]
&`�l�҆"M�$:��N�{��������yB�3hv�!s�o����0�����*_Rp3�i�C�y`�$�>EQ-`�D��ț�Iq(9�!?D��QPїo�6�s    �    �    c!  �'  �(   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic�'�C�\���E۠_����p���T�?D��x��=X�`�JTԖ�Q��7�	�e��)�A�Ur�O� 9s�jƅQsp�r�W�U���'z�ٲ�	D�LT��R�m�Eg8S�O�;@e�@]���D1�g~��:FFF5�0��8Pe���׳�y�d�(�R�+���:�P�ѡ͙&�&��E%U���y�7�'��0q���`Pp8WÎ�� �a�A��r2��=/��@��?#� "��71
J�ভ�/c�1@p"Obt��������)W!T��2�x�C���Y�mJ�.8<9��S�5�E�G��*u6���@�%2ǂC�I�ut�1�)�]Z�<�bӥl�YC/_8c2`ڡ�ڃ>�6\�2�1�3��ոkT>�y���	UKD �2�B����d�j�Ը�6nO*�t�Yˣ )Z���C�;*c���EG�%a�=��>��x�!V�U�7�
dJ��+O¹3Z��Ǣλ�2�����A�J��Px�%8rcX�l}v$��.4���C�P�^�XNP�]�����8?���0;:��k	��(��C��O	 ���.�1gb@3L�X���'�RP�+E �ީbF"L�=�LS`&�!9Ruv�
&$��ڷ&�ŘO��', l"bb�Z�(��S�sZ��	�'� m ��>A�l����$t�d@"'�-@0��0���xܬL@�E�!d��y��{$}��5����f����0<�$��5|�; sU<%{��]�? ��1�
�������R�C9�K�J94���r�2'�ތa�d�8]bl�3�5} �v���Bo�1Ў�@�l�{�O�
ycuȓ6��MB�N�F��y��'�](� �(�`�eH*Ġ	��Iϥ2�P�����]P���F� ���G��Q�Y�MY&� ���0w��̆ȓ0��	�LĚ/�Px*B�Պz�����`KD�����b�^����(U�S���4rHoK1#�a{b�Q.)��l+bLB��P;��)Yd�,;UB�8g)�i �k?D���xH�Ix�e	N����1�	=d}B ˓�J��>)2�k\��8`�#�Q����=D�D�!�),��5�a� _���On�"��v�JC~2�	~���D�-I��mO�x
��c�[.eS!�G�CK.ph�"Z�!vd͠b��\�v`�%N-^EI0�'�h��� ��5#�!�?:�k	�M���-OrqR��J<���:D�/?0����"Oq�"�K��P(� �<Q.�1�"Oґ�⛭n��I�4_�0�"O��h�� 7IEftc�O�@iZ@P�"Ouk�>_�D����1oڜ�"O���e�1YvVD��/#X�Aؕ"O�(����(���.P�3�0�R"O�@B
n����E�Z<3vJ���"O����?
�.��3^�\����"O,tc�,�<TI�qNT"��&�+D�t7&%2�x���`d<��H*D�p�qB_)G}�)�.^UHl�*��=D���c��(��(�``�)u/,���$>D����&6WB`���s�Rx`�.D�4@��E 9�z���N�0��1"'D���̭� � 2��B��@�$D��B Z�#�L�`pmV���I�%!$D��a�Ć ��G,	���ԣ D�dk�l̊W �:���7r��ū�d-D�u�M�T��a@�	<��A6�(D�  ��<ܩyr/=�L\��*(D��+$��hY,\��l�y�લ-,D����m������*�$9�.D����B�:�
�D?�d��a"D�(``�:c�]7���:�i3#�<D�,1c�0U��#�dA�[*vLAG�-D�Jt��|��8 �Dw�( s �,D�h�.%Z��E��i ]0Ѝ�Ţ?D��cfNV/%ֈ@��' �Z�r׃?D��ĸ-&� 4	�%"

���<D�$��΍/dZD#vf.� ip?D���T�˩r�~��Y4 bj-ЗJ7D�����;l�x�%� �\�K��*D��kP��qr�ʄ�Jo$�q7	=D�8QqD���A
%I�6xq��R6m0D�x�g 
u��zC�Ӂ�0��:D�Ԁt'ǉ���qc$"�H�#�8D�tju왉N�҅�'ˎm�H�7B9D���c-�f�`���9�"���%D�4rC��(�O��.^P��(D�,�AJ�=T����n&���E6D����l+>��z�Y/����&D�̉�޼4%��zT�T�P�x|�#D��G��e�@�{�JS�=�<��%d D��!�Ȓ�Ix�@��'R�J����3D��Cp͎��0��&��F�@�3A'D�� +��:&d;�%]
=���R��*D�� �>4���=Xc�Y�/7D��j�)I���9Q-�@Rp���!D�0`�K0?،����[��\�,D�� �A��#�Z�j���ڝy��Q�V"O��P��\�RM|4��2 ��W"O �aa�9]�̰!t��"BFV�xw"O``�"�L�I�$uAg
Q��v�"Oޜ�b�])!�����菸�0��"O6�vAD�!��M��I�+e&���"O�x�Q��o<K�)\�W!��"Ole.�
-ሑ�a�F�	�|�R�"O*1�q��Ci��z)�1�8�	Š�9��!8�xX�dKE\*Rd��e��(\L$P�!D�HQ5�
�~��Bd&@9P=D�����9H�PU�c�]&?�i��B<D�D��A�%Ю\���M�em:D�8�rg�
E���e3�Ѱ5�7D��J�,W�y��P��QZ� D���)�=CL��OT�VQJWi?D�X�P��0$�j���l5r��@(0D��s ��%`1��6�-H�xQ�/D�|�FnF/T8)��i�f�Y�#2D�t���`h" �Wf\.FQ��0D�$�ua?<��Qs�.ڜh Nݻ��9D��SG�'��"�+S`�n����7D����D.xs~qP��P�T��$�! 0D�8���U<0^�����>k�Pix�1D�P���A�,�{��H�9��D<D��35��T����wI�o���Z�=D��A�[15κ]����(l9���$�?D�d"r O� ��3��"c��H��<D�� Sü`e �Y�H �hv�����8D�T�B�.���J�I�'N�{�3D��80#N1'�4�����P5��%2D����[�$n@�ᠡͮny��I��<D���Ƣ۲0�e�̚-�`�+RN8D���w�U�������S�&i���2D�t����PdY�*ǋv:�١�*D�8��'��e� �@���#�a0�2D��R�E3iTN,ڥ�H�fl���(+D�����s�%ZWnL�L��&�>D����+Rq�p���]$�r3  D�4c���1�x��g�Z��(cf�(D��#��V*g���B�be��J��%D�x+!@]�lM�i����n�C�.D�l"%&�{�t:e��)G�8%�c,D�t 
�!/�p�󩇳I�
�s��=D����� '�h�	��қHF&�a��;D�����W�?���fc3��'��q�<i�#H�f�6����s�����gYR�<)F.E@��v�.{�L����C�<���C+"9bS	ީ%���h�h�<y��@��Reh�V�q��H�<�fmI%^����JT-W�1Ӌ��<���N�Z�f�ޖZk%R��B�<�O�Ab���b�a^�9Td�e�<��N
�@P앂�ŕ*q8���Eh�<���Y�  �|�OXw�^��c�<��I&gd0�BbeB�k�Hڀ�Sz�<�&�KI��5rmծR\XD3i[j�<��LG� �-ba��-<@�Z�$R�<�2_�}Fq�JS=qU� ���J�<q�(��4���`�#���:�AE�<y�i9	��< �Oߣj ���ь�~�<�!B�gG�]{��!=A�9j��Ty�<Q���>6sD��eMĞ~ d9A�s�<�SK
>0�2�C BN�..����#�l�<� >���.;Xp�f\��Z ""Op����ɠc욜���38��p�"O������\��) kD:	��"O@`
!�O�|-��ٰ� ��s�"O@P@%/I����r��,v�Xu�q"OH��QM�XֶȒ��+%%�u�"O� �q�)��Y E�;
����"O�4c�D�{r�����$9�"O�8s%Ҏ7u ��-�|l�6"OPP�JT6&d�)� ��f�����"O�BU���4�捐��H��x��"O��M
�ZO�-p1��<p�����"O�mL�i�n����<]v�XQ"O%�g�%k�	��\?Zp��"O�����P�}�x���сL��r�"O�<�W�?tтqÈ�x��%�"O���`NΦ)�T�E%E=��ɐ"OdM��ٖ"
 ���?^���D"O� ��v�|=K�ذm�.���"O��� ��������ױ-�|��@"OԵ0�Q�+��@c�]5�����"O40��킠.� +#KQ�l��@� "O0Ar��1��A�䩈�"��Pb"O L�S!ˁ�dc����Z�"OH�z%	׬P�ĹB���azG"O��!%�	�\�f����KR�Z�"O���0BD S��x!�
�FLU"Oa��1]����#�m!,�8�"O*���D��e�dⅡ1#h!�!"O��Q@��!�d: @J)g�T��"O`�i%���u$�%�i�j�"Ou�����8R�2i8��"O�iVȁ1���Ҏ �Ln�m�0"O(����>&`�g�C� xb�"O��BO
z!ҽi���Pm�P�p"OiK�lXV�`i��h�Qxt��"O0$� ��\� G�n�af"O��ѡ�SgC
��Q�M$Yx]k�"O�|E	3~D�f�ͳ2>J�C�"Oa��fB#ז����h��	�"O�`�u��_x��x�����A"O��{�CS�~b��B

�(�FPe"O��Y��W�6��b%��o�$T�$"O�iH���K��-�j��q"OF���T�| ��!��h��R�"Ol1����j�}Z���R�j1
0"O<Ԫ�+[��`KDj�ٰ���"O|��
S�R�~����_�jqK"O�Ȫ�L��p8�X��,�8�R���"O<`A�'ð���`2F���"O�$�ٯ���!R�]=���"O�x�@��5�JM��I�O/�,�@"O���v'ģ~��G;	�X}��"O
�g҃0~X(ö�yIf]��"O-p��w:�x4G� B!���"Op书KŅ�Q0V�?d���P�"O�a
Ul�Px�����j�8�9S"ON�1�3 Z�}9�hR4Tp��y�"O���T��$9A��-�,@�"O�5`ㄹ-�q�2�� f2�ۄ"Of�ZP��
O��ëƱp�����"O �2��L��% M~�"H�"O��1'៰DY6�n kâ�"O@1 �B
��v��v�(X�X�Q�"O� *EX3B��H��}�w����"�"O���,ҹ;,a˲I�>�h}c�"O&d�7-X#9�mYa�Ҳ-_]�U"O���@�ؤiݖ͉W��"_ �!�"O�;N+r�(���	ƞjAn��r"Ov4���.C��Y:��҈1����"O�ܪt���fQ�]	Ř<|�Q�e"OH��4gI]�~e���416e�U"Ot��A��1g�|��vO��Hl��"O�8����N�eR��M"�p�У"O6P���B8�<�'�*l�^p��"O�hR��N�7��l�u̗�^��t�s"OD�Z���}�z!Z�M�=fv�Ȫ"OZX�F�[�&5��
��D1����"O`�Cu���B$@𲗊K Ojh�³"O�A9ݞ.:D��0jʋz�Lh�"O�X1���L󦴙`C�-(�,{D"O�� �+�M��ܓ�A�';�
`""O<\� CP/�p�"��3?�5�"O�,Z�U ����ܭ&��p�T"OD�ȏ��p��ga��~��m��"O�0��화�����8�jq$"O�u:gD\6 ;�@�U#��2�����"O�<!!�	=�Fa;EɃ�ؘ��"O:"�(٥����J�+�٪�"OPC&R/�ĉ��ł%}r���&"O~jai�3�HI��٤uU�i�1"O>!Ȓ ]#0s�h���2Sp �g"O�|@�� \lH1�t$�e��F"O�P��(׮cYZ���,��_��"O>�Ke���@�٥�	2eH8��T"O���A�xz��q��D�G���"O��3��Q/6��!sƭ��=���v"O���ťl`�t����A��Y�@"O�p�Hϋ%"���vH��"O�$o�ٶ��¤K�}� ��"O إ!G��Eq�C� ��h�"O��*p틎+�ԱH׃	�F�,�b"O�ER�n�R�S�?Zӄa�"O�s���>殡#Ǉ���Mjr"Oԥ�$��)jƃU==x�"O�Ő�E5j�R͓�䗜/�ȸd"O�hA�bv��UAQ�-.�E��"OEz��Zg`mi�j�34?ZP�V"O<�����Vu�ӊ�e/jeB"O�h��ǅ(dH�1Xg	V*E�|��"O�({g�٥s�9�'c	o�V]33"O�3�	U���=�A�-�h�3"O�(Q�#��L���+e�
�5����"O�U�� �ZW���'���nԘ�"O���`Y�4��H�,V1��K�"O(|����pA�$�� olS�"O�p�7+ GW��2�)ϰjaԔ��"OVpCFc��N����1L�Q@"O��O�C��'εKݐ�i"O>�$M�4*Jy��2o$>�Z�"O$�hS��Lh`���I�6h��jR"O�i���N�,�Z��!�N�7"O��k�IO7���+Y{�IR�"O���wK��k� �l_:.@C"Onp���%f����6K\5r6l�"OX\��N�1Vᚁ��&��P6"O����C�<	I��׷d�t�'"O0�РhE�5\:�G�rq�};�"O� �M�dKڜl��9����-{Q�1��"O���e�>`��+��23���"OZ@��^FԸk�g3���U"Ox����;�n�[U�g�@�P"O�H��� ��M�W��%a�5�"O��jY�1@�e`��O�1A���"O�A)�
��p{�͔x0�:7"Ol8�Z���� ��u�@�"O~�G�8IS���J�\
ViS"O,���"��~I	Ā#�8]2"O| �Lk��b4CSA��(�"O��ؗ�F-0~ c!�>���{w"O�Ç$�#n��(��@Z�UJ�	jF"O��!��  �   p   Ĵ���	��Z�JwIJ(ʜ�cd�<��k٥���qe�H�4��S66<���EO�f b����Ɗ_)2$���Ϙ^86�����I"�y��D�<!ĊɠH�hp"� Y&:�`�<W�0��D�c�㞤IR�ɼ4��˒*W6�����;qz� �m�=���V�(�`[���D:vVuR���d��(4�ġ��$F�ar�L&[�B!�!a���M[T�Ĕ0�����(�Sߟڝ�aa�!RЁg�\}���G�bU	4����e�cc�!�O�p\9��u~��o�|�R!8����q%�,r^R(�u �!0�m�R�O2� ��<�y��]��3�gÉG�
��Ł~}b�+S���ӨU�j�Qv"�&Gdh��g��>�rq�=IG�8�<��Gj��נ-	4���,h����c
��[�S�x���س.H#!Z)28 SPa!}��K�'-���=Aw����4]�Q�G�VX�v����b�	"Y��\@ԤWDxF�b��f�lyh��� Z*b�|j�ቌO�I1`,��E+_F��6��2X��˓i��#<�0M*�I6���ņ�h��k��7GD♀�����r��'�2���)L/���ˎ�ZH1�y2�NV�'��$&�4�rĕ�N����k ��5�V������I1C�'*v���cbpiTh_�@��Ct�r@�m��Ss��y��YR��'�8�-O뮼�h�_c��Ya�%�8wJ�ko߄|��y���]>�O�3H�(�4� �D8z��cn�!�nt��&�>9�8�;Ǆ#<���L�]�M���;J#� 1B�d�<��h�= 2  �"���oH�w�L�R�SC6Y�ȓS-$�K�ʈ�x�P<�3 \ �"���f�`T(�� tX����"�h=����k��EAd)E�m#"퍟D8���!̪d��<Ԯ�btGA�Mآ�ȓ!���Pe&���f/¬	�"h�ȓz��iҡI[���Y�͒#e�Դ���R��ī=;VX��oWH�@l�ȓ.�|i�2o��R���a�&97�хȓq��з	7_�u9;Et���'���wnƕ����V1B@�ȓc�8Eǘ�<N�� �$ձ\�~8��L)�I��)�f4�ɐ��*|l��ȓf<�mԤH
da�p�j�t�&)��� S�LEB��'�8�L �-�
4���� %J��X�'�\��¦�v�:ɬ�'q�Hs�.�4���[e"��H�(���� ,�� y*zX �"O� \m2�-�5��\�Aˍp��Ȼ �U��,�a3*H���)��<��*�?`�����W �6��l�E�<!�͊6 �t�� ��.��)�����<yC�M�Dy�­=\O�����9�
�`vm�y��	��'�����O;3�ra�E YjN��'�K�f�^0��y�"@�lQXt���T���`�!�4�O8��f℃\Ӭ����)�3d��c
�w��Hq! ҠZ!��77L��r�8k3�I� �*X <@�C՚*�`��N�"~Γ^
T�
�W/7:��yqJ�i�Q��9������Ϙ ThY�p t��I�y|��i�'B��$��F����
�J��ez���a|��
#Ḑ�e�ӣD�d��k�d�5	�F2p�a��'׮���AQ�W��-��������䟁?��u������(�8PI�Z7 �h g�]�>m(q9"O2h*B�\�^��m0F��7o�@Г& �Ĺ�uH^���)��<�Q O/OK���8*����\p�<�B�Sx}� ��]l��t����l?�3`E�-��h�e���G�EU��� Wb����	��"1��'��r��>FP"��'��P�<��'�l���%�	N��Cw�I*���'��mV�B8'����JJ?���S	�'�d�"J�"h���8V癈Bh��'�~(�����<�P�됞w+bɲ���^;�>9(��W����S��0d�]�oK�!�$��P_x�T]�d��!�n2p�]��A'O���hQF�S�R('��O����6Kv��(.�~��7"OD�8�P��%��x H���@@��9�s��Y[JT�'�T/{��I�^�Ԉ��;M�� "pD�8l�
��d��E��9�m (���Q�F��"O��`c��)c�Ԥ�sB�`���'�ea��JSB���AMGG�ȓ�}��2 ���K�e��( D���79�O��b3�_��$�k��D�2Vz͙	�'�L�
�͂0Jz�p��@�(^��ao�+�<(�$癀�A�����7
�,�I.�\�șw��К���P+Rh�Ј5q�X	�']�L��;�7��i�����!ʗK3N�p§<D'�u��-L�T�d��'~2�k$�ݗ��	=l���Sႆ$"�KfD��4�4��d��9s2���}��!�L�$S� �i��%����T�\�1Кt ��H��B�J�K�I��q
�'�M��`\��� .� |���B�y2N��~�����7h�4��h�-��wȏ)7�e��[�I�a�$O��CBڇ#�Y��'/���P!�z�b���J*�0R��Έ�T�'O~�ҙ�AB�#-�����|�l���j�(� z�w����5F�h}� �G�ۡ�i	�'����Ռɍc��X"w�Y~��e����Q�0��H&t��e��j�_x��H�,�a��pz�
�y��M��O$��%HBaJ��׌Ϝp�D�	�v�<1��]�\;rAS�B���%C�+'H1I£�.C���b�ه^4�͂"�$>��bĬ�+S֔u��	�;�6|b�˔1n"ɚ�����RjȘل+וO
�eKpi��L�r���J�nu������� �ѱH�y[c���N��AcJ�sH��'�� c�؏wZ"�&#���s��06Z�� w�D�@mօA"�9��(+EtP:�Ɲ% �䑛wo�U�A�'X-(���V0$�~�K��5j�}���C; ��q�РxP`1R�M�^�$�c�A�@�1��E�"6����O�r�(Ѿ,��'��)��Y*6�����[�:��э��d��2s�O�iC�hj�DV+pB |{
V�t��4��2;�:æ��6v�b˓>���`,;,O��[��LUߊ=9!�E,����V�t���W��+�nK�#��1��ն`LL�>i��'�M^�0���i��(D���Ñ\��	1��t�M;�-�H7�������s'N5 �l����c7�>���I�F*B+�? ��K�*P<�3$]�|���H!� "ZM ��UJ�<T����w�^	W 4�����X���۰<�D(�2zz���g��n#s!�J8����j��x�2h�L�A)8���@-?���`5B��7�е� �"O�5�6
Ͻr��m �B��$� �Ap��S�I��h n��Py�#}�k `t ��������
B�<	D �8i��xK�i��;��ġíѡE���v+w��b�����H���G3�Y$F;Yy!��H���j ��n'���f�F�W��	���,���Vb)|Oi�DꄖVy�\��3a[�j�'n�2�ٕ �V)��i����NS�R�~dpG�(�6��	��� "�zv!���Ԉ"�O�rU41����)�Tҷ�Ա�h"}���0@|��70x�y�@Q�<A�jTXP@�`��3$g�`ƬZ7�RE��EU�dC�I�k4Q>˓��8;��8�����[�&����ȓS0R|����l�F�rQ�R� K^�l��u�rm[�T+n����O�]C�:�d��qmH�y�{r�֝۞T��g��������TO �ք�`l��+D���
W>Z�^-qg7p&��@�+�I$V�Y��蔯~��>E�	��}��KH8RP@d"�L)D�����P�����K�_&n Q4-�;}_�"����	N��~Bi�)H�M�1�[�nɚ�dņ�y�k��(JDO�Y�X�"P%ƍ�ybI�#F�=���'eĂ��-
�� Ϗq��x�?L�9��q�$��P7Qф0�W-�7=� 9��-D��p3̝���,��/[� ̼s'�&D�$����r��8�X?�)��"D��:�,�
1�����?zٔ@
C�>D��Hǝ3^μa�`�fN�ɛd�>D��h4(W�s�� �Q�Jt����+D����$f|��f!M:L�6'D�l� �$kVӃ��.��ܙ���� I��eta|Riؕx30q	AK D<�u.�0>)�`�.A�xa��L\�{��4S)����ۢR�\Ʉȓ=�B��� zg^9�4���`�|������	�g�O6�#i�|�ӌ�i�:���k���y ���G$!B]B�nSL��3+-i��5��Q�FĮ8Ѷ���=�Ъ�ZL��~�� �u�+@�؊��U�U��K$U�.�H�㉒V�R�3s,�Uܶ�sPJ�<�h̀6m3~`p�A�V�W��X�!�'��`#��`���I�$�N1�
�+���@�+���W$��W ��V.��+0^�' \i��8|�B=K�N۔Q~�H��^= �7��!��]G0-��&R�}��ɂP�ڠ(ƴt�DҁXa6��G��-@����X@:%��O�"�+���M7g�q�r�U(:� �  �J�5�az�j�A�X̓^j��h�DηE/���d�Q�0�~iI�״SC�|;��N
�`�ח�?)uϵF+����!����'���t�է,��"�h�Z���L>)��CX������@RU�2'ت�2ԐթK���	�'��<��Q���l� j��G6�?��l��$4q�FI�G��y2�9��xV��j�Yv�J�T&%Ё�ì�1U�L�1�H��b�'2b���<���iÌ  �tR�R�z�rP��	\�2K��j6$C�ɽT�.� �GD�wdA:\XK��ζi~<����dB������r��d�V!��? Pp��z?1Ǉ��=�9X$�O�(�x2�݆Y�=�`"$,O^�0��S��<kܴ
i��T\- 	� �0��K����^}��ѳx	,e��Oqy��W
A����Lr�I�0a*W������5�8Od=ڥK��`e8�4E���˷��G�b��� M 'X�]�I�(��H��1��dQ��K�:�Gr���
�FY����آ;� |�b�A�\Y��E�Ơ���K�O����N�R3d$���S�|�Hَ\N@ �vb����?�Px���o�2�90��4��"�+1hn��iқ���.�,��f�n�>�) �n�D��|�n�7\�
��Q�R0[�4XE%FjX� �c�$c�
�y�Z���
Z*:���.�-��)��Dl�^Q{�4q�ص�M�"~nڮ/,� {Ce	,���@�
x�O��!���z���	Wed #�UNJ��#KY'��I�l��lj��\X��y���K��ģ���en�(X�ě6k-���=a�u�'UN�u���?K�`c�Θ	9�<���9D\�%��'�MԋόO�����,L��C����h�~����]�tY�� E�%n��!�CA"�!��ŗd�`T!wj�( �sR�A$D�!����`�pP�
�����NS!�#�ڝ��I�O�
�����%!� w�y�$�.Oٔ"t�)P!�dӃZZBa*QkRC����c X�m	!���+z1�(I&r��d�q�@�K!�$�φ�H$h�03�� ��34�!���~�0��6.ǁj��\��n�>}�!��
Y�XXcCY�f���@�^�!��O5��e��H��S�Ʌ�e�!��Q�Pd�O� t�,�!�� �P�c�P4"i�Տ�mX	�"O�%8�mR�#���0D�٣[�T�4"O����BOS$�q@!4��"Ot���B�*�3R��K�Q��"O<�����H?��� ��Z"O���K�#b��S`�C�p�L*"O,}ᔯ�N"&���Y0X�hٵ"O6���(��:�c7cP�P�XP�"O` r�F�M��2�m��~��4"O�i�ӌY4̖�a6>�%lO��y��ا[�����Je��f�A��y҉&0���0�(�NW�����'�yBL�=�f��̩~e���b$*�yr'S�I�v�C ��8`�ĝ��y҇G-"B�D�E� v��yF����y��{��er��}b���(:�y�Cԛ3ʘ����t�i;�H�y�䞁,<���˜�\�*�:!�R"�yB	�t���Q�"��U�>i�`���y�%�u	<k�њ������D��y2�/'N�,rC Ս�&��Rh ��y��I6O��2���3}�e:3���y���7ܮ%���
5��(٢ �:�yҀ�j^��CP� ����=�y��`��aϾ�����&5D�p���70��d�68��-3@l5D�hj�藇:�%�Y�^��c7E<D�p�bF��\v���f�U3��L=D�L{b,ښ,h�
�'F}�)ju�=D�8f�66t�k� �[�4�91F;D���2��y�ұ� �U>4��#6D�Ъv]�K��Spd_�jt�27D�D�2�Ջ@(�1�?�ѐV�3D�x�1)�h�EJ�C�	��a�#:D�����6W��+"ݍi����%<D��3�IǢK1�\8�iO/� ��(9D���ᄝ�nM�A� �>�ꠘB�4D�ԋ�^W�����	Z����S�2D�3�N
h�N��`�K?v����2E3D�8��4�>���"ǖ{r-
�#1D��(��&Tg��9��ѿ7��(��.D����dE�xAK��6�zܠa*D��!!��DX�X3���8�T�r��5D�8sB�'A�$T�C�^�^sD3D�����ɣP��l�q��.���Z��1D�أ�hK�WX.3��D=D�� 	T�"D���a�v���y��^?Q��QBn5D��	�Kфej����Oe����$D���M�\�x`�R�(�j)�c#D�h����nn���e�!^��1Po2D�Tf�alHU{��+*.=��3D��I��3s(�ّ�E;7P	��.D���𤘋+	Rܱ�dB�y4F����.D�$1��Þ*��ذ��/�:��d�1D��{w@�C���� 1T�e!�5D��qnO�e��&� �Xc�'D���N�9Ʊ�P�S�<^�`���0D��١�.�R���]�~zu�WC*D�8����&OC�i�O۪|i@�o+D��x6��	"Q<�i���6�HA��c&D��&$%=T��Y����0��Q�3D���A�G�7k���*
2����!2D�`�І�F��XЂi_+���ڤ�'D��h��߅>����%�ڷ-{�)׏(D�� �I�F�"�S�]�xK�0��'��)@ �$*CI�&g�H�@��������rd"D�h[5鍽{�ޔ1f��<Fl�\���"�K� |sei=�H�(���n1(��q���$�ʅ��"O��� 6��Irp��H����oذ}g|Y����)��<�qN�xd-��/� w;��T�Mx�<��%A0��k5\6����U�<q���)���a�%3\O����#ˬE����F<�)�C�'�,���X/�L����fA�A�*W ~e 		�	� �y����:ij�l�6l4� ��OM�@����&�(��Ă$	B
d�^�13��0A��S�"OY��� ��!�f��()��Z�Qf��`�H_#��)��<� ��1��E�$�~5"(��G�<iW�^�x�<��w���e�����`��<�g,CzXr�`&J=\Op�z���i�C�?	X��q��' �U�r���!�� �C��"�����m0Bԓq-��y"BʒY�H
�k��b}�q����Oꤢ�� /����$Xk�@iU�4#2p�R �Y�!�X	�����L$T���ψ1(����Ѐ��*ږ��L�"~�|�����U P�j,$�@�ye�]�ȓ_Q��X3�ʀH��L˲(H2f�h�ITP7��Ű=�`���&����!ȝd���
ҥFX���5��	B�E&,���L1hQ��,�$�y��؟z3�]����3�����ą�y��,ݔ���'Q9#,��C��y"fɨQb�:ƂAA���p�dѥ�y�Nʊ��6�M6.P�@�K� �yԀ)��MΫ_�`�Wƌ�y�EM��J�ΑLHμ���A���'Iʴ���R�S�'9
�*�̜<?6�H�HD~�Є�"�R�ʔjR.��cA����FQ�o�m�ɱ�LE��Oq)�%ά0���Ɖp�IjdO�t�&B�ry�s�,�6d�!�#�Jg,���_���>�0@'6Z����i�NR��rA��wX����RM����R�h�Ԣ�=E 49�a�0u�i%�-D���ǤK
��[�	ξW!�PL*�S~!� "�Aؕ�M��B4�c?����t|�9Q�B�#x0X(��+D��dM>Q����F���~�᥎I���+۾Bjn諁H�[�vb?%�Odhk�a�0c��x�5
'd�HO^tЖ�&]�򙛣LA0m�SÁ�n�tQ���߸8�P q��<0l��I�� �ʀ�ߒW�(|`j�"F!��D�>&�lm�� ��D�J$1c��$/�=��"�Pn���Ԑ� |��\s<�󌅠>�f�34��k�(T	�%8�\ ��-����Y�L��:U�ܴ��D���%8t�	���%	��n_�T�t��-�S�r��B��!�D߄V��;�lK�(ؽȥ��/��!y�� �θ��`�	YTX���o��% � e^@U9�NE/,�^p��O�������y�<H�E�-�H��I[wZ�)��]�r�hR�̣i&t��Ռ�iq2��$�'3r��C��^����v��	aO�eb�'�;1)���2/����:�i��Ǻ:R��.8L��M���h��ǉ``�(��ďi߈i��.�|�h�o^��ZQ��N�-e�bL�a`֩
�ꥨ�'St: ����UA���d����V������^eo��za�W{Sv@�O=��]Y�F��|���w�N�x@Ư~a&މ|"�=���h�@�@$F�d�b}	�'�Y�]�և��QKz�+��gv��eˑE�I�fr���%�1��S�~����e
/���[q��*=�џ(��"�/��aҖ/�2|�������@cœj�>�����$�h5���|��]$�l1��I3+������<r:0�E囚g�\˓C��`L�j`��#u��j�|#}�K�P��u`�"^-vl41y�<q�H^4{H�r�)R=Fp�	��E���yy�G�)6�"�sTg_�)Xȭ'?�ԛb��)zc$���lڨ�`c�)7�Ћ")�kh�IW�#3��U��ʝ��=��!Vv� $S�e��P97#Q�F���	Y@��ݰ�O.OA���fw�3cF��y2�g>�3ǓQ�F���A	��y/�q�^u$_*1Ķ�X7-Y8��'�n��6l|�G��됇@��8�Ԧ�4,�Y)6��5�y���-b���y�m�.[�`�V+H�+B�B6l�����:PQ>�S�? 4i���2u�Y���S(~��M��"OHI넀�) <)��,P8.�>4�4L|�R	� ��ă�|��qArخ��r�z�"ܷ.q�C��c�X]�� ւA4���	��y�ꝌG�P���/?k@�ywa���'"����N�P�t$��Ӿɪ񙗨�f`�8P �I�C�I-+�.���O+Q�paF�5N��͊m�X����*O:�K��Y�TA5b¨]�s�Eܹ[� ��!/D�Ќ׀TZ]A���1�lӘ�2��@(,$��J!�'���5S!`Z@ڥ�9$���
ߓ\_T�S��^-(�
6�M�cOZl+f�4t	���� X�Be!�d�t[�����P�S��[ i�O�m; aL(�R����0�`�F�uY�2��2o!�ċ�ٰ��jVH��C뙉'�̋��J�b��OL�}��9�xd��M�હ���,�� ��$B�䓼r��K�F�MB��ϓ|B6����>��=�B�CJ��yI���N%fmb���C8����Ʌ�F�d]��Z���n�=Є�G��,2�!��=w�A��@��!Su�ǅj�!����ad�@�G�T��b���!�Ę�}`^��ŝ�D�{G�~�!��L�cU8a��O㪬�T@D��!�""�I2bo�7٪L�m��\�!�F!L|ꅩJT�i�aPSU#|�!�DN�!].@V������Y�K�>X����VP�0��\��@Ӗ]3�0�$stم�0o�*����̟��gJl��%냯K�l���Ǐ,D�P��/����$q�M���4��O q)`�ϒ�~�eϡR����G��A�O�B�QG�j�)�)��n<Q��"OHi�dI�0�$0�%gG�e0��7�O�@i@sJ�Yw~�Q�'Q��Pb��h��Sq�{�+
�TXђ�,ON�����`�*z��05	�`�E�5,�M
pj�aB�$	 �&�?I�Y��N�)v�/lO~ęU�(d�#��	/s��a[��r@��\�����ȍ=���0�����)�Ŏ^3j���[wb����s�,"�
4v(h�'۸��@k��`pC��P6z\6AX��
�.���F�U]}��eaנ��+C�|J��y[8Yp�w?ęz�^!6F)ф�v�p�(ӓ��`R�*f���A�U1~�~m�b�Q;��QwkI(�q��ו)n��î�p�����'{�nu�Bf�
>���<a�c��98������i���Aov�h���/Q��P���N;O�!�֌@
�Q3���*Bl]���J27زP�s�^+-`M���x��8K���$?��]�
�8�hy5�?ZA�b%��pf�8�S��M��ȂX�<Q N�Gx��r�����
R��h�g/>k��,<�y��E��CL^�1�
O�%��HD�RV� J��J:�L� o�m�T�J��ȠO��{A��#���ʖ�ĬQT���z?�o��A(~K��M��8:�F8��l��F.,O��IԨ��v6��48�]�ʲ�����[��0�$k�K�S!�K�I��= Q�Mcy2�E�+�8�� �a�~����V03�@���oFwVO���e	�<����4k��=�e,��R�:�q��t��}q��n��
���S5Z�j�@��S�\��e���I$�'^:h*��A� \t��#�Kuh�� �B'`i��@�z=�ԉ4�W��h�0�ӼYa�ѻjP�6��m��_��ć1�A�fAV5���u�B-v�ب�E�$b4Pc|��b@g�z[I+���V4��'���S�*�t�@SN��*]3u.�9@Z���:-I�Jܶ��V=9l �$�Kc���!!M1Λf�G�	��� Hg�ӧ������o#�#d�����R�@������z����0|J��ǺC�l����}�̭+���^}r���7����4.Qx����S�}��9"�)��;�M0��P�{�qO$�p��@	���S���\J�@�{� %��i�`�B�	't�`	T���qKʘbC����">)��N-�ȣ|T�<(��S&/��?hpP�,RP�<����7 ���)��w������E�<�e1)�2�+�$S�R�١�%�}�<�a��F��KvC�K2�a2��}�<��JC����j��MG�%��a�b�<���Y�FE6��dɚP�P�
Z�<��k�$��$C�ޛ0��@e�P�<��8y��@�<��UX�+Q�<� �10W�'%jl����ш,Z�`�"O�"�S2�|�2�S�6� �i�"Oޠ���n0��a�T/��Aiu"O�����ОMU�-�BgM �X	�C"O���nV�>�y�#HA�,��"OpP��İ*:�X��S�1�65!!"O�#AF�1vq��"�����"O��J�DL�ð��ʆ��I��"O�\Ba���B`Bn �?�luӴ*Od�Kg�[��=���27�8�	�'��]�df�/;Y �*F�%�"��	�'�EG�D�i����/,l��@�'Ǟ)Q�(���L��ō"e�f�#
�'mx /�fz.��@�>^�0�p�'�
�p/4
��p�G\!y>�8	�'��i��W�� ��g���49ڽ��'0f�	.$r)L��e>Y����'�(���fϨ��i�Dȣ;���'��ar@Z�,� ���5ː`��'�t�����]�T(�A�.[w�Mp	�'��,	��R-Zwba1�W_����'�j%0�ƈ�3R@� O�W����'à����/�8�d�E)�)��'u�x��"ε��*P
M�:"��'m$�Z�Yuj�R��F�2�6���'����cH�,���fX2%$ٺ�'�6T37Jͦi4"Թ��(:f�'�~-���$(�F��$C U�&���':a[�$��n���\ �����'�~i�e�֓M���1허)����'��k��>E|�a�`���_�4��'@ �*�͂c��tBӥ֟C]��a�'����`��7���z��;�8I�'�L�鷈:w�ā��$֪S���
�'4���V�^<�%� �I3��˲#)i:��Ë�1-����|Oȝҁ@�Up,M����<u?�]��e'
�y�헰+�����������L���fɊ�ohy��,�D5��ȓ<�p0C7HY�{@�T�Hr@�ȓP��%��^� ���F�e����M�����G3V%�-�"NQ��b|�ȓ*T�ƭP���ӧ�	����<�ÇGI���O���J�)V�@Er�Dd��
&��'�`7��؍�'���B^w� �3?�')�d�$�4J�f<���V\���kFA��E�,OrE���O=L��W%]�,(�hT�g�B1B��T�|T�	U���(1��	�fǓ0��	�M�d�8 ���@}rh�6i@!�֡@���	Ll�OE�Ub�H��%v�u��h^B�HSd�V���Rr�7��%���O�?�yPƋ4%�А�œN�	�1Ad�L[�@I�A\8�'���	ׂl}@��"l�,xԜY�)�ZQr)��'�,Ô���Mx^Ԃ
ç)�R��G��jѨw,S�R�x��Ż�~B�=c�P����+����O� J��p��cyp%%�����8=|E�X^M%�����۞r��d9�����d��K�UD��!7(�<a�kFy��IZ�a�J����w
L����تΦ����,��	�'�8<'?-8I~�6#�20eb� �q�$�6"
�h2И�0#�V�m�;a"��}n:�+	�{Q��B���=�4��/O�V������������|xX���S�{��@�b�*wU�  BF� @�h���OV��'@�2S�W�?����j�|_�<еJ�xg(%�@K}"��.U[��3S	I%���Z �\ �+ZGjX 5l�	C�D�$�����x�f�E�~�>q(7���>sPF]JY�@��`��S�p�^3�ݠ��Tb�ѩ��\:�!�$-]��J�O 7.5ry@p��
%�!��/1�X��AӑL��(c�'�;e�!� 
g"�9��L�S�Z���O�i�!�d�>.(*yJR(�8φ(K#��2!�� ��S0��?iT���J��p��E��"O�)pE�ڸ��q
���7����"O��!���o�T�ZB���8k"O>�`%o��%���($���mrX��"O�I��ŨN�@"q��M���ɐ"O�h��K��P���	��=A���"O�;��Έ@r�� ���0/2F"O�%�`����	�b�:"W�c�!�ٳBl⸒7/��>i�	�v�ͧN�!�_�S��`��-4hf��nE	2�!��4d!�Հ�m���P�L�!�FY�<=�;U6����"�!���I#���'��I�pxQ�B�[�!�P�R��A{U@V�H�P�����&&�!�dUz�>�o"Z�&H� ��!�DX%=��b��&Z܈c�.Sk�!��-_$*w[�byI��"!�=~�,���@e>NEZ$��'p!�^�@�Z�0��L����-z!��2�`�"�F�SH�!#g�<r!��3WO��j���a>��B#&�:gp!��w`�t%R=r{7JB-S!�*W�|{���-�T���F!�%)�����_�m{�@�fA�$)!���{���;rT$d ����>Yj!򤌆@�T�3b����E���]K!��[�R��!S o�w���(r��y�!��-?���J>|���T%�?F�!�d�.���g#R�tx�U	��aK!�D��_a(��ԁ̏P�ĹQ)B�#F!�כ[� �k��(��	1����m�!�D����4#P ��0Z� T�A"[�!�W�y��q����O�@�	㉈�!�L:o�.Q�q��6�D9� ND �!��0-PZ���ʅ
����Т�!�ĕ�GjLfB�Ut��qɅ�!�$=xޑ�a�: �r��6)���!�d�&@E��
Ԣ�F*h��P탄b�!�D�>|�t��$�Ux��<�!�d�F������'���ǂ���!�$)3��c��-Y4Re)G�N�/�!�]%o����ʰ*w6h`�R�y�!�$�?����ӛjZl}��`	J�!��͒Lŋ�̃{���@" ��8.!��LJV�P�b*��e��rr�̇%!�DÁZBJݲ�	�r���3��|�!�o���`$Z�t�0#� �!��4E@0�#���4#�aD�!�
'��4��([c`��+VN�a!򄛙R�&�3&�8nC�11�lS6rP!��VG;Pp��M�P*Z}��J1%�!��Ǟx	�B�3��*�jѵF�!�D[>Y��ģ���0FըQ��O�!�dNcs�HA`��� ���*�!�d %-���1&a  �0�RW��*U�!�Z�4�& ��LSX���g�<q�!�d:9<�5q��4v��y��Z?\�!�č��b{�M��	�R��фW%�!���}P� �`߇�4M(���G!򄀃=F$`%FP�d�8����ZIV!�A��� Ʈw�y �\%SS!�$������-�-a��7L����R�5�r�!mڹ�lI��y��֬P��D�!��}ɦ�9&ڗ�y
� �D�g�ʁgF` ���!j.�#�"O����Z�<M��$�UW��Y�"O�a����"'K� �C�<o6pI��"Of8{�C�>�j&�<`%pE�7"Oj��b�Ēx{�HE�]�5�Ekc"O�)���\&0�@8����2�`"Oz���ߋ�2��v��	� �r"O:����
)��|Z�#	Q�ؘU"O��q��#ҭ��E%Җh�2"O,���/�`����#�+)$ʬ�C"O���D� �TK���d`p�"O�)sW)��Z��#\K�l�"Oʴ�P�&�>�I��k�`���"OΉ+��ԇX���X�^]�~@BW"O��D�ϯU�����KW3v�� ¡"O����n7����٢#��	b&"Or`z _�
�xE�s��r��a"O���&-L���A��_1R%09"Ob<�'gq�0&j�1��I��"O5�$�B�E]�e*ѹK�}��"O&�xD
N�0i5d�xS��i�"Op�P"i_�1��0��P�'<L�5"OJ��t�V�H�� �%[��§"O�|ђi�"rHhׇ��pҐX�"Oа��C�$���ǔ$��u�0"O<���gÈP����2&�-�x�W"O����
�HO�Ar��W
)��iB"O*���ܧ|X��{��Ü)�X��"O��R%́�#��cg-��#�V�iD"O��qv��B�Ѻ�픛"�d�S"O
d�d&�6��X�M�d.�qW"O5rc�7>l5!���Ѵ(�"OH Z� ˕)��`+2%��[�t�"O��`��8��ph�a�z�Q
d"O������(���OR����"O*��uAH8^�~9��d	�\�R�"ON�"(�;��	t)�._�,5�"Oެ���3�j��'y�.�C3"O|��n�r~���`��;m`Z�@�"OB�+pD�>ڌh9�k^�r�z�""OD�[�N�7'��y��a�t�"O��*���k���U�/b	I6"OȰ!�f�,J�COQ_���V"ONI�S�ޟSs ����g��%"O8���K�{�������|�� �"O0TZ��H�sm����K����"O�%���()���F� 9�(d	P"Or(���f��]��Z�7�P�q"ON`��c�d�YC�k���*V"O]���H$"#j$��l�E�z"O8���ӎ{���I!0�d�a1"O�l�kȗcGb����kYr�qC"O֥�U"���Ait�X?�ũ�"O��{��ѯ2�@,	��̵P�0�"O�;���a�U�� ԛ=A� A@"O$XV�v�� 7�1|���	�"O�`�ǟvg�t�U �V��e1�"O������4C�,��(Ȱ	5�u��"O���#�X�{�����@�&y�D��"Oy#畑 ���'�D� \{ "O.Q�C�Q3
�� �wE�]1֕��"O�9 D_�"����]5x����"On\�g���p�L��N
��"O�FI
�phQ���
Ҥ��4"O� l!pa��	�d ����/��9�"O>�"�[:J�0�"��s��A�"Ox 4
�:|��1uDFb"O8�1�˞I���&��d�)�"O�n�*��Dh3I�����OժD�!��Ƞ@:ݙ�l�j���0��!��Je4���J55�Bu��D�!�ć�?Qr,�g��*�	`d�!�D��V�@кA��"*�j��D�!�dD���1,�!�F��UÁ�_�!�{G��6AN�/^Xj�!�H�!����@�Bd"\�f)`���4�!��V�j��M��-��`p�E/�!�$�L�Pq��C���=;�D�F�!�d��Y� ���
-'��I���P'Oޡ�d�$5�
�p��:}J�`Z�A��y��� i��S��O�]k��i Lӊ�y�Cݽ|#�K�,C�H�ɛ��V0�y(C�nhct䔤R�tH!d��)�y��]1�̀a�ڟ���
����y�%����9�ԥu����D �yb��r�ŋ�'o(D�5��-�y"'S���p�sJ|H���d7�yB�NFP��e�)<m��(�	�yRlZ�r�B6E���!�ϵ��4��'���@eD�1=�A+&Ɛ+lX���'�4��̗�xO޸be'�	r���'�^�J�V�9�rk�/�+�:Uq�'���QmѢG] �td�3
z��'�*B�@"�@�3JC%����'w���fȀP2<�B�+U��(�r�'t�����W�������Y��)q
�'^u;fE�9}�0�K"A�����'��	�n�?w����B��<C,�J�'����a�Т�F�5����'3���@�1��`"6��,&e4p��'��ԁ�Ɍh U��X3�Xx1�'ǾMA&���S�X!*����h
�'֌����+U8Ȑ�tO(u \0
�'�����.Km�D0�	^<t�X�	�'Bh%7��w�pT��9 �D��'p"����X&���#]&Q�;	�':�`E��q�<P6��C�
�
�'Ѹu`Qfխ	e�l��4�\�	�'a�})΄1l��A���W���\�	�'ox9��j�T|ma�\�_���'�x,���	
 W���b�� Pm��'J���e杹��,bả�f��i�'$�����6^����C&'���R�'{�E�biB�{�0��#���P�
�'�B\��c�%#� ujG�H4���@
�'�Ι*�@Z+L%�D!��-#�JiB	�'�xe����b�~l��-ƍ!�P��'"����L�e�h��2l�
eI�':Z��aش"*���e��j	�'l�idA�O���A�0$�i��'��4�P�	��+�F�#@*�@�'�D���Kj�^�"��Dh5��a�'JhH����L�Re[W⑴p����'Lb�"�	qF�]����#��Gy�<aw�'\��UrU'\-p���AFPt�<� ]�L��@��E���m�<�4��0�6i��[0ޘ��#�	f�<�2�����dE��)Nq��hM�<�+w�   �   �  ,  �  �  ,*  u1  	8  "?  eE  �K  �Q  /X  r^  �d  k  _q  �w  ~  W�  ��  ې  �  c�  ��  �  '�  ��  /�  ��  [�  �  J�  ��  A�  ��  ��  ��   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C�>����鞿6�!d��x�^��I��~�!��
�l����v���:�9a��:uZ!�L�,Ƞ�#g��UԀ�e��t�!��v.qc�ʁA�P{U�C-h�!�DD�x>B��cG;c�lK�,��"�ayR�	� Q2���F��u�t��� �/��C�I�Ld֘8����D��T�U�#�fO��=�~bh(e������M?��m���Tg�<� �������T�����R�g��dR"O���ѣi�A	�͖<|l��"O�ȁ�N��SO��µ'�#{u�L�"Oҕ�sGY�>u�0@�'B>]ԕ�b�'I�O 5j����)ɲV�л�"O"}��J]�P#JLa�׊R�Q�֓|��S���O��Ḡ/��l"�88�n�:!�D�	�'X���P��u�҅� D�l7�<��'{���6f-虡4��	.�<�R�'L�Q8�C d� ��욯zA��'a�l�3�F!C����4},0|ϓ�O�4 6g�'���z�h�!�P�R�"O�$Kue��Vrl��MΈӲX�S"O�!X$�ZD��z%��B����C"O:0���b�V�a@���VĪH��I8�\��׆pT����Y)i3	=D�$�&���;�#!a��9��H7D�|��BP���x� 脖~g�T�#5D�H��
�Kh��Fo�Z�s#�'D��)F�^��$H�/ǐ'��(#D�8�\�.V>���bYO�9�4m%D��3"�Pq�f�2P.p���(B��$K
~%x�b1Fb�la�CN�.��C䉮T��[#A�$I����(��AC�C��H�XtN)qH�!!��A��C�IHh,����s�6C K�R�jB�	����#塕��Z����}�B�ɥ~�� 2
?<�[�"��nZ�B�I)&�ĝ[uj	�%��a��;�hC�	�f�-� ���=��d�E۸a� B��;}�܉�e�1(��1��ġ=JB�I�!�\3�oԾ�p��C2h�C�	FxXz�g��dp�Հ	c�C䉇>�6���a9yVa�W�vdlC�	�!2,ҧ�?U�*�����5�0C� XwZp''�q�1c̀�ThfB�I(wM��+����k�I�@�ӽ	LB䉆���F^�=*Q�@GB�	�4�ܵ�!�� (Yv	`s��7�B�	?s�r��d����hj��I(8�C�	�g��d,�(M>�h�h��q��C�	�TTx�5��<�� ��&��C䉿[.� �� �a�P��/ԌV�tC�	3F�!wFY�b �'NV��C�	>=F�m�FǵxZ8U�ց�	tLC�ɦ:�p�n[�u�ҴY�!ӣd�BC�+;���U&�<b��T�@�����C�	<+A����Ǜ �R�I�.ݻs�C䉂Ԫc��T/T.nL���ܴS�B�	->�N�9�N��T]@xËZ�a��B�I�E�Ĭ1� ̮j��� A��'�B�I8[�2�r ͫ���TP�]`tB�$�0C$�!O�偷ƛpuNB��]EdP�o�4'��m
D�ُ9.2B�4$�t(*d�8X�}cRd�+DB䉷L�T���k�2n�i�CE�[SB�ISQji��6��{@��/'�C�	�sϴ�;u
�?�X�:b
��~/�C�I�F!*t��N�:�0�h�-	NzB��<�C��3}"%���CW@B��&`H�ܸ�Ζ)��p��+� .fC�	'�n�x�$t���2�I8�^C䉟2�F�@�╧Nt��q�ŪXtB�I15D�"� 0h},�H���yA�B�)� ��aF�H=�`z�aN�'b��v*O��xc���2�~�0����}��'���� 0����
Wl��*
�'��ԁH>pxcG�o�����'\za�2mF�3��H��ˀ%o�����?)��?����?���?���?Q�=�q���-xpB�ѧ�B�j��9��?i���?���?9��?a���?i�vD�U����;�Pĥ��?P����?A���?���?���?���?q��S�x�+��� &�h	���#OVlI���?���?���?���?���?��j�$X�գ���l�o�d����?a���?���?����?A���?��(b���[tu��+�B�h�J�2��?���?����?���?����?a�I$>�K�m�����Bl����?��?	��?���?i��?��,�lyGm�1��x����n��,���?��?���?���?����?��g�x˷EǂP�C���'�
�C��?����?I���?���?���?�7ⴹW)>��
A�������?	��?����?i��?����?��s��A�N &)*�n_�a ��0��?��?1���?I���?����?a����*��)[�|��� ��r�J��?Y��?���?���?y���?Q�z�(��P��
^CB�ve��A�Z)[��?	���?1��?)��?�c�iC��'�:�i�ƩQ+x��r-dԙt��<A�����0�4)�f����s�P�p��&�:�S�C{~��nӘ��s����9��S�Z�A�u�_�ƚ-��՟�R�(����'Z�	P�?�����uc2&MD+0�ѯs�du�����Of��h�d�Uk�19�A�v�R�q�2�a�����#1!#��L�'Ad��w1���G�[	7��%�ECN��xM9�'$�?O��S�')����4�yR���B�@T@��)T����pM��y�9O�����ў�ş�%�dȌ��#QV5���%`�L�'�'67��-�1O�0�vg��k��Lץ
�ؑ��/�����d�O���u���'|��Gw��Ȃu B�}{�O4�DK�1
>	���I.�?��H�O\�p�n߲iM�:Q�F�Bc�m ��<Y(O���s���$ޑ6��$ѳMyE��uOv�`�ٴX�t-�'f�7-+�i>�ꖉ Q2�8��Q�'�a���o� ��ß@�	�ED�n�q~�=�,��&c�<hJ��~KL,�&ş)���#�|V����p��џ�	џ�Rp�N
W,
��IV�LH*3��oy�u�mIB��Ot���O̓��d^��%D�8Gr��i���Hb�Ʃ<����M��'L�>���O�;5($s �� �h��MM�Kx�S� �>��@jhy`�ьO�ؖ'c(`�C� ��,��D�	H��'/��'�����S��ݴ`� 	�@F��	�/􁻂�D3`.d	�Z�����g}r�i� 	l��tK#�^�p� �G7Y~���D�Uo��m�^~�닥�ܠ��w�'ojk�3=� !e��!'2<)�+�T���O����O���O��$9��b�.Iy�$:?F ���>/�(���՟���9�M�$)Y���dNߦ�'����M��d�di6�ώBb�(CUFN:�ēM���Fu��	]YD�6�7?!g����(� 
����s���?�Jx�$��E�F�$������4���$�OX�$R)�e�5ᛧaU�l�FnUd�$�O�˓Z>��.M�\��'erZ>�05#�+$�����LDA�=�l)?�_���4 ��v
&�?]SGKE!F�:�tB��@¸��4u T0h�I3���|��`�ONd9L>9����IF��Q.2�Ψg�ކ�?a���?����?�|"*O�$o��Zm�U��h�r����L_!h��I�������I��Mc��B�<�4w���E픧��=9� S{$��sǿi��7mC0H+�7�??Ae힧����3��[�j�x���,Ү��qe\
�y�P�L��ܟ���˟(����ܕOΰ5���m��eg��$��XXmq�(x��-�O��d�O����dD٦睈B]�a���q#~-�
ӈh%ډ�	��
O<�|z��0�Ms�'�ص 7���NcHLp���A#��؟'��)�4Ǆş�$�|rW��S��k���FTn��"��6%�Rw�\�������	hy2�{�T�*�OF���O��.���P�C��Ii�r�Э8�����D�O�7��]�'e�:D�P�1R���i�d�	ǟ$#����2U#B|~��O2P��	�x���0'��(e�(ј	h4&ז�"�' �'E�����"�!�3����^�qo6`x3�C���4.G~�S.OBl�l�Ӽ#����Is�y	V�A<e�L��E�]�<���?��i0�a�ia�$�O���WJ���!*�v'z���n�4���2#�F�RUp�O���|����?����?����>4��D�5����LN2,.� )O�o��+�m��ȟ���X�Sȟ��G/�-?�н�d��Y�b�*�(C����I妹��4Sg�����O���H�3U8�UY�� Q�YggI*Ly EY��d�*\�n����*h��Of�(2��2�K�4�X�d��蚘���?	���?���|�+OzUm�
INL�ɺ/?� IRa�8:x(�cC+��H��	6�M#�2$�>��?׵i�\��R�*1ՎQ�G�N��Q3#7��:O`�d>Bf�Z��Vb�	�?��=� vmS��A%1TCV:l5t0s�4O���O6�D�O$���OZ�?ᘡ�.n�Ȉ�ɇ8�Z�#"��Ny��'_F6��+5�)�Or nW�	&P(vă����j�*@M<	���?�'hҰaش��d(<	��E�ϢiR�|
��G{J�#�C*�?�&�,�d�<ͧ�?a��?�U�O�"ߘ8{V�5i���Y�	�?!����������ٟ��I�� �Oh�I���.�J�*��6�&��Oܘ�'R�i��O�S'Y��YA`�<1B,�!!���t�Dy�eo�()ں�s�:?ͧZP��DH���bd��q!�M��1��ɮ�	���?i��?y�Ş��d�ͦ5q���$u��j���v_����+^5A�X��'��7�>�	���pӄ�b��;L��6ʍ[=���EOH��P�4*;r�4��$��X;~���'��5��]�5ɂC�5{��W"���Iuy��'�R�'���'��[>uP�Ɠ�e���QBOϫ�j���gۀ�M�Q�?a���?�H~j�v}��w�"𠱩�
,��(�EC�g�ԵSv�b�v�l��<ɪO1�0�1�}��ɡv�j����W�Jq�偄�qUd�	�js~q��'6H�&�����')n���J�X�����V.TEK��'��'m�Q��"�4h`Bs��?���'�N BT�O9z�*q��@V���i�B&�>Au�i��7�WC�ɤi��9:R�II!b��2
F���*�#ϟ�t�D�|�c��O�D��0��#�d@(5�pBvI�(]�
�c��?1��?���h���$Λ<�f��S�[�8s�Ao҉H���Ϧ�P�B��D��:�Mk��w�t�d��3[˸p�WlI��`�'F�6m�צ5�4}��`�ܴ��Y L�6 ��z�v-c���m��!�@�~���cB7�Ľ<ͧ�?a���?9��?���1]lM)eeA�S3���r�U���dW��M"q�ןX�	ڟ�&?�I2de<��4�E_@�y���إ
��IY.O~�Dr�>]$���[�Ş_4�ځ��o�(M�wӄ#��!���\����B��f�	cy�
�nH����K$t��Y@��f���'zR�'��OL�ɪ�?AE����@g�ż'�� Y��'g�@H  ϟ�a�4��'����?���fk�QθZ�K[vhrYyA-V�2�h��iH��e�X����O�q�d�N�& S�b�ײ�0�����Z>��O&�d�O����OP�d1��R�L0B��7�^	���->t2��'$�ix������?�j�4��7����N�.6�6�`F���\0�x��'��O �Ҥ�i��I	T�{��&L&�`��ǌo�� �p�ؿvn2"Lf�	y�Ob�'�Ɍ�J�4�A()8[P�ԗ���')�ɮ�M{����?A��?9-���(��Ģ|.��S�D�	���8ѐ���/Ot�$g�\$&�ʧ�"�c�X�n-�HA��:G�2�#��D�$�N���"}~�OT��I#z(�'���3V��VT�[r�ϊsjV��V�'sR�'�����O��	��M�1%KmȾ� #Z/��
�!��zF���.OT�l�`��/�Iݟ�w��	[��ٛ!ǆ�}�\E
\🸠�43�pڴ����H��Ÿ����+Z>�$��2�r�U�1�D�	my2�'���'���'��X>�WDF3Ӕ$��,%s@]A����MK����?���?�K~�F!��w�h9c�[	T�V��W!�_wZ����'�2)%��)��+��6k�� ���M�p�!�'аC��б�$r�����#|B�H]�\y�O��Dؼ�p���f��سQ�Y�4��'���'3剸�M���I��?���?�sd��l<dK�C��L�2`C�����'��ꓬ?I��H��'V�Hq*��Z�,ʳ��)+:(	(�O4�ٖ��(J P:`�IN��?`��OF)x$$�3���Ԥ�<�l�`&��O����O*�D�O6�}:��4&Te*��4k�t��0FS!{GR�(��K��f�ɸB�'�J6m3�i޵����u;����$þ���i�j��������;ش�R1޴����(oȤ�'|�8��6?��H���9$i��*v�7���<ͧ�?���?���?���=|&�u�aE�L��%9uFY����Ӧ�1
	�,�	���'?牝T�d-��!V1b(�3���>�P�S�O:�mZ1�M��x��t���k�$	׆��l?�0Y%ˀ��T�aH����Q0�����!"ؒO��.Ɋpk�@��#J�����|���H���?����?��|�/O�oq@v|�I�E
j�!�J�� �VA��ɺ�M3���>����?���i'H����?U�zh!π�(�S2aWd������lA�S!������ld�Beǡ�썣+��H�B4Ot���Op���O�d�O��?���E�`�8����U�3
d��b�Gϟl�I�d�ٴfy ��'�?��i[�'&黳��-������
�i2O�W웦�q��\|6�+?q�ȆD�ШB���3#7�#�윀r���H�O�9;J>�-O��O��d�OĽ `�����)��� ��E�g��OJ�ĩ<�'�i���<��柠�Oz��(�	�H�Ĥ� d�zX��O���'k|6MS��i�S��du�|B�I�Z��"�F6Q��	V'uSB�RS_!��4�P����ָ'?2�h��M�8�h�A�.x��	�'�^Dt�/ƺڂ� ?tI�	�S�~�-Дh"q�A��Q=�P
�e��5<��@�쟃�С��B�ncn���@NR�iX@���HvgĐd<��6错;� Q3�O�R�\� ��e��oP�yh�͹pT<"�̟E�V�Q�'��0��̛���4/���H�B ��A!"��*��Ap�,�8���f��[���,o��kf"O��g�F8�(0_XeX��S���pT&I�c��'v��f�7��ݫd�L�y �E8F�F��q�Ȳ ��k�� ��D�F�[�|��`�`�����N"r��4���Ŭ<a>�F��e�A�!��F|-�FDN&aI?:<z8H!E�bXlaH���-H(5*��.$���%"�K$�� �c�O\uP��� >�6q"D�K�9C6�9Å�O��d�O�,�@:Jy�nW���y[�IG��������X��#E�k���Jg��)�(O�<s��*�� �	�Y�"+$�r���T<E ���9P��a�'Ot�'r�D����?�O~����t�z�c^���´c�:��$K�����?E��'��	�-��`8��`��,�>`����'�'�����
Roâ:�&����O���D��P䊦o�m�R Y`+'4!��թ	<��!�1Bz<�ꡨǽ4!�C&��A��;W Q�pHߋz�!�$�2��|�Df��| ��J�AH�Z�!�d9�Z=K���bg��%��br!�$g��e��m�� L�9�4BƃXh!�$Y�f�T-�5���B�XZt�@�y�!��i���`1�Q�T��
C���,y!�T�{V��%/���P]PP��H!�D�7Ul�@���h����Lև!!�䕘6��B��Q�چс�AJ�r�!��4 Vl�$J(P�x;6�)=�!�ě�a�H�8P�%�9��$�x?!�d�/&�b�F���l��S7@�!��+ێ�(�NA�+"*Q�� �2r�!�d�Q��"U#H�a:(PoZ:9!�$D6~=�UJE�N% Q��՟;!�6NS*���	� �'�n�!�$T�r�p�ra@A���u�<&!�DQ�.o
��'�Z#'���׉�2�!��� �@��A
B9��-Q��|�!�$D<��y	d"F�b�^1"�m՘x�!򤃪q54����YXX��l��r!�ĝ�[�6��GBY��{�K b!�DZ%�X��_�8�x@�%��uK!���*N����(����cӶ28!�"z��Lyˎ��jd��O�_L!��?-h�D� [5G���V!�䃠��(z�SN
}S�f)R!�ď�{��S�'߳7J���Q�T M!�&>�$����
n*�U��O[d!��s�<�)��?t�l�ir��RL!�){z���n�;u�>��Z~�!�$M�17[Q��E��yұ�л�!��g�A��{��I�V�z 衇ȓL��air�O�E���Ƃ�4`�괆ȓJ=�!�*w�x)�JB�d��"O��bR!JZ��݁B%��g}t�KT"Ov����&��)���)���z�"Oh�wM�0�p!��u���(r"OL!	R@>R��a��f١��R�"OvL�7K�e0�����ߘXՊ�s�"O��%� =hV��U�nӪ�2�"O�}x���ј�cW�W�N�V��$"OR�ă��3`ٰ��W�N]�a"O�Ps��ϻT
�#
6`��m�V"O:ԃ0-� &���cJ���[�"Obm��a������#��BGJ�k4!�D��N;��h���)eF��b�>!�d�#"^ �B�B�B �͠���EG!�l���k��W�H̢I�'d�>?!�D��Ji`��Q\�,�QB�?.�!��C7'�8.)v`m�7IM6 ������ i!C$µu�p�n�30���"O��A�a[�F,,l�-C&�nyx"OB�0d��2HL�x3���eې�"O&M f�G0
8���.I�bl�q"O�xcGE�X$A��+�|�"O�ѣ�FG����Q�N-SC�q�"O�B"��@=�H!W#�+vEp"O~���X61���g_�"l��T"O�8I2�й_Z ���'˥����"O��Zu�h�挠��� LN-J"O:��чѧD�9�4i�#7�t��g"O>��C	}_26'Y�<%R�94"O��B��������ܪR��A�"OL���"�=p',ac�Ϗw.c�"O��!��8M�H��/#����"OR,ٗ�qIr��:E~0U��"O�+��"���bg�'5{�LJ�"O����n�S��qq�JE�MD��T"O��
'� 
�Xx)C%'�UI�"O�p���*3`�9Վ��.�Pl��"OD8���܇pI�`9�&��T��*�"O��Y�,���N��e/�g"O�yg"�/v�$�H�#]�*,d��"O|��p�Z�1!i�R��A>�y�"O(	榓�]3&�+rb82�"O��sVk� j�M��K^�K�j��u"O��!��r'��:3Ii����"O���Ǘz�A��s�^(�"O����o"*469 G�HXŪ��C"Oĭj�DI+!����'+�=�S"O���0��zڂ�Y��Y`�y"O�!���>^��)UD�_\]P�"Ob]��HV�+�\y�RC�]�։)"O
�fE$ }B�Ŧe���"�"O���5�V�?�,����Xئ�	 "O��2��������#��9��"O$)ht+�0Vs!���'=���A"OVy@oϦb$ ����A���"O�E�N�`� BfݿK�zE �"OP�A�'8Z�����	�$;PLB�"Oބ2��ԌPW�p8������"O��� �]�%�X�* (V!�@��D"OLb׹�V�ز@��*_�P��t�<A%���}{�ms����"i�4�]G�<9�/�2q���K_=b)x �fQo�<1�4a����ڒ!|�4��Q�<�LT�P,h�!bU�P�:�[��q�<	�	.XP�S��ňb�y�"��q�<a��ݒr�&)X��
�d��f�[l�<�I�7 :fa�k�8���ʑA�<���6N��Q�g��V}�`�+�{}�Rx��	���)a��FF�_�����%8�O������<�N�LѤ0�&mj+1�o�<qS�D�;	�-�DI�D@h(0�KZC�'�rHi�0�k�uc2�1*=
��� �2���O�����G��d$}�ek�.����N�i��O?�ɝDB%�� I(�:X�R�2"�JC�r�($K����
�2#/�0J�$��I�D;�@��$��#��lx��b�ߣRt�Ň�&v<�p���A	��$�\4 ���O���b�(@)*�!�92A�Ѹ'�J�D>�Hr�'IH��'��Ip�/Y!*��E��Oƃ��<ȶC �@=��D\��yr˔;1l`5��D�zH���jS�W7L��&�ņR/>�ZmE#)�M-F��é��9�����S�? ���Q��
/3j80�(�7 rg�i�JX�mV-ǰ>���(�$ً��:O���x�@K؞�Q�aǵR/p ��$��z����Dd~)b����w/v���S����c
�(�b��iH8EDx�	׃H&�����T�9�lyU �4;Sn�b��E�T!�䄑(�� ���L�H��+�l�N��b�/ �' �>���8�pv��~��(�c��*Z�zB�ɜ+~J���Ϩ]�]�Q��(BP6�_�`zZ��R�lCP`\2H�8���I@��%q�$?lO"1K ��d���~h}�1��0��q����7�^��ȓ�$�s��JzX)� -2B���?�AN�Z��H��I֜4�ԑ7'Z�M��L!�Cě�!�d�%/ND�,�$�l��C������թH��b�"~nZ��ҴB6��a�
	+�n�vC�	��`��=%^� ��j�L�@��+��'��xb��U6W�B�`��IM��u1�D\�d0OD���64����*5���r"O�-��/�;l�����!4�)��	�dm���):>@\�a�܄0��IBᏑOb!���u�<�&��?A���z��׬]�����p�=E��4�p�C�\H�I:��N:;�&��s/�x�ph	�K�E�G@]�#�U�'��[D!��=�0�ӗ:=zr�- ;���c�JX������u��6m�p�\��E.k~X��K��^�!��,&I<tXf뚾H��@�d�Iq��H�Ee�D��>���!��Rq�TKc��D�e�*D�<�U�76���ӵ�!.l�`a��tӪ���
LK�S��MKCE�4cBᲖ�l��)Q�Cg�<��Ы-�E #�^�^	�`�g�WN}r$(a6���d��U2QТM�8X@=z���)~4a}��3<��I.���e�Q� ����G;6B�<3ꜰ0&EG	:�i{�Oq�"=�!L�)�?�"�D�.@1C[�t֒��<D��I��J�5�<��Z�G�8T�C�d�4\����w�S��Ms�F	����B�_.Q�Xm���[�<I���-Sr��{ �. ��f�Uy2��p>yA�\�V<��KթH'9bA`D�PN�<iDh�c���#��L0lJ�UN�<A�nX�����*	(�}���J�<yG���'Lx�D�E|�lp@�_E�<�5bz����!b��{�����[�<����m�V)*hj(�S��S�<�Qn��6����'ԦN��Kf��L�<y�Ē�7��r�*�96�飰��l�<�`�ƨ!��I�愜��A�Ġi�<Ap���/�:���J\��xp��l�<�ҦȂ[F����	-[<�ي1̇e�<��f�l͚l8c���j¦?�B�	�nw���#�Y4U�2aCj�i��B�I3&�I$,
�-P���_�`&�C��8c2R��E��x���T!�C��0,-��ȿ4i�ZV�Y0`zC�Aih�@�G��BU���=@C�ɑ*`(�j>>Lr��?��B�I� p���+9�d�x�N�a�B�I��h�;��E<� ��&L��Y�6C�ɷ������( �I�C�	*n͸���e�	^&3C䉁?�b�r�o<!���� 7)לC�	�Yޚy�FK3e�l�h��`��B�I�i8��W�5=���;��B�I�U��Y�v�?A���HԤ��L�\B��`���JgIka4�Ǒ_!X"/$D��� �ϠVbR�gL@%Yܼ���/D��  ��nR5W$V�b��b.Љ��"O���a17U4 �0́�S%�	��"OPi��jY�W�<�d,�?~ZI�Q"O�`�-Ϟ �R��g+�5�@��"Ob4z�,I�U��4
�)Z�3@"OXM�1��X%Z��6� K�l�s�"O��ƒ3>�
���a��I�:��'"Ov$ ��2j���f(s���R�"O��Y�,ʙ�
,1�%�YkX�F"O ��'/̀���CϩR~i�#"O�Yڄ�ޘ\&�\Ygτ' ��sP"O&ܰ�
5Y]\��c"0�&@J*O�S������sV�1�`S�'��񩠄�3�1U���K��XJ�'A��0�*W<@� ���ِ@ 4�
�'ۆ�RO�1`����OH;᎘r
�'BYʴ���V������I,8�ƝS�'�^գr�[�k��Ea��ڢ&@��'�ڙ�D�2<���ϳ~2�!��'����F֟N�,�AY���K�'�R�!B��YD�k�i8~�V�C�'5�y���΂2��ᓢ�Vs1z���'[zDZ*��z49��4l��@P�'چ��g�#+VX�q�[�d����'m
�A�#�~Y�P��,1��`�'W���OA�J|h"��<�x��'͒�R�f 6'Yb��`Ç ���'%��IEOQ������V&��'Ȣ��g �4b8�	�	��}Q<���'8�����'�� J� ��@��X�'#�]s���|��Q�eEm�X=k�'�h̹!a�ڎ�C$�� TT�':���ʃ��,z�i�)i&���'�8��w	�>lܴ�C���̴��'�P\�e-JBg&�h�]:!����
�'�z%�S-S�H����s�ܸ
�'�2�Fn��'�&9�v� .�ab�'-�)S�N�Q�;A��-l�έ��'-´Ҷ�N.@�q`#�ؘ\��\3�'�q+���S�9+��T"?3\���'+n��iNb����8��(C�')�xpi_H�\�h�JP�/a ec�'
,� gV3A{&����(�$�Q�'5���˖8�vDQe�-ml��Y�'�8���"L�``Q�
�����'��2&�Y�2��{B�]�;p��'o���@�6!iQ����*���y	�'���b�# ,M�I0�����I	�'4Zy�AOP*L!z�C��N+9æ��'<�:6�TE u�&��
i�	�':�(g�B! ���R)�]!Ԣ	�'�"I����첢k�,�F���'ў��f�46A�[�&���j
�'A�8*gC�Vݦu
�ψ4#�<z
�',)��	(%)�(���t�9�	�'��XC��O�>	zU�O�X�`S�'$��23H�x��q�����v�����'�xY �#�+�"itO�$�@	��'V�]3�EE���������'���{��& �������"�A:�'�v�9r�
c`�0K����;�' p�AAǌM$��06G�=Z�'����`�pE��b�ŋ�'���	�'$e˓�S�i��%*�iZ���}���� I�F��&v�"�R�P#
�[�"Oj��nC��X�Q-D,u6Mp�"O��V�&���;����"O��R�l�b� ���#h����P"OԚTm�)=�@��bQ������"OP\��&�	]������L�$�D"OV="u��BRx��qC� �����"O ���aֵ���K!�Y�?��Ԛ�"O�@� �ʍRQ��yCAʎ�ĸ�"O�5Xp��_���Q͕�K��ՙ2"O�8��&ڋ��	P���cܤ`��"OJ���gUHD��p��Ы}��X��"O\���])X��-��c�F*a$"O����7
NLm* �_�/�(p1�"O:�!�'vH���l�(V,�4"O,���ۈ	5�pr�˅Mv,��B"O6�K�ʚ20[�l�-ɚG^�l:"O
@1�LD
J��h�U�R�ոd"O�9B��O��KӬ�&8Jص"O�=���L6D�B�"�N5����"Oܘ�@ ��P�N�"F�S"O�l�0N�"��9����I�1��"O$�s�@9jEBT�@�r!^���"OD�r%(T!Cv`u��hs����"O���H�r���P&�V1'�fi�&"O�a�Q��!zZLD��ǈ�A߾��"O|$��K8=�d���۔a���"O�	�#F�h׋�iqL��G"O���piX�R2�I�kÂ>il�0�"O$)Iq���!�/�CGt�JV"O�%#ծM�mBdXc��Qb����"OFk��N�WP� I`�/O�̊�"O��;p'�r�0(ʣ�
 ?@�p�"O��@L�"Q2�[�14��p"O�;3L��(�����:@�y�!"O(x�b��!%��l��0�y�r"O@�5圐i�<���L�;:VFA�P"O"��Sn��`((m	;<h, �"O���af�g�Эj��J�Y"l�"�"O�hT�\10Ą�ɂ��+#"O�l��0W$I�E��P2�"O��t��@�R�3���(��J"O���jLo-������74�,C�"OF(�UGaJX�!Ƣ�C�]r"O��YR�F6�
�i��B(�fd��"OB���cT4(��e9��9æ�w"O�Y.�1%��b"%D�N�Ľv"O���Ǝe�����CM'��H;P"O�i@��Ff��$BɳC�����"ON��ો�V��a2���T�Bh@�"Ot؄��W�yC������"OB�[�d�0 ;�92 �D�g�%��"O�2ri�I��i���oؔ�""O�i
�_��+��@� �|�jW"O
�{&�P1����V��
�0��"O�M	6#�*�N`0��2;�,�!"OtQ�Z/�6����
�Ŗ� �"O&�`1"��.i�gh6�fe) "ON��e�F'U�.�7�¨B��P�6"O������X͊5
C*Řw�40xP"Om9��+�Ui0�_�R�8��s"Of9SV(���-�!� |�"O��*d���P����qm�r��s"O�����4Pz,�r�oΌ��"O� �H���[�^��R�ΎF�!3W"O��Ѧ�;&�
�ٳ�(�����"O�́���P�����b�$�i4"OZd  ���&�9�����F"O��Z5t� ��۵62���"O~���'�uN�� Ê2M0�)�t�'��D��(��h�$ �O�r�=�ȓ;�$	aTd�V�4�PR�6��	��y�Z!�ܬ#R��R��?4"�}�ȓA�ָ-9 a���]�H����aJ4D��u%;\E:��CA]��-c�*O A�T���X�n���n�{���D"O��#6A�JNԥ�$`	�Iѐ��r"O��@���1��(q"�;V'��ا"Oj�:" �>e"͐�A�u
� ��"O�l�r#ʴ<�L1b�<_�	�"Oh	�I:6<f-i㠎�;��u�"O�-�T�Oo�i�f�Y����S"O|ܢ�ˌ5�~��u�ژf�e""O
pA���T�p ���6"O�����K�AA���dR�0g"O�����.���#�N]��r0�W"OFU���&�~�K�B�~Э��"O`T� �B�q �C�CK�"O�T+3)��|�U"M8[��-Y�"ON����.EcDq�
B��d��"O�0儋�R�TÁe�p�ޭS�"O� ;���f�$� ���c���X�"O$H�C��A��U�BM��/N�T�"OJ91$ܤ	��X�ۿD8�x�"O4P9'k�G�������MJN�`"O�IiFg�;D��d�`G�}��"O��@��Ne�%"ǡU
M�*D�Q"O����B����a�����w"O��" = L�Kp/E20��"OVԓ�I�|P�=�)_�Q��"O����Ίd�� TB
:fni�"Oֵ����@�^̸g�@��h"O���CBT�M� �����"O�!�MX-P�fPr�^]�k�"O���D-2rc�V��T��"O��k\/���
�k �5Kd"O��a$��>ܡ���%T��"O�q��b�b�nm�w�[B�4��"ODmQ
������� Q
�I�"Oڬ��@V.`���
T�9�I�@"O��9��\[&@��R�T�D"O^�y�]�+@��A�;Y�0�B"O($�#շqæt���܇��y��"O2aԩ9� 8��BÑ �~���"O���a��Da:�h�n~���D"OxB2��!@������"nl,y�"O� ��n'A|&�BP��P_\�rS"O��>y�bG_>S"��"O*@q"I�l3���#��?I�#"O���R���`��	�m�F��"O��	��̑�nА�핳M5*$�"O����ڦR@m��˕Y n��"O8��`I/M����*��jT@$"O�1�E��d	�
4�J,W�H�+3"Op�P�ˬ�ܘh&��&>�(��"OP�Zq	�Sb;�抣e6&�U"On��g�K�j�BE�P��7��J"O&��螂(�J@/���p���"O� �s���v�F��4�i�<�cD"O�I�$�!0��Q�#G݄}�&�#"OQP#֑��y;�^��:�h"O��[���d}Ԕ��>,$��5"OB):_2L�!��_!:>�0i�]��yr�4͈U����(�l�w�Z?�y��@ld��0拷�쩓VjP�y`����Ҽo��정��$3��	�ȓ"B���R�%"�H���L���ȓ,{r`�3����t`X��_8��ȓ��@cA� �X�w��;�l��ȓdx]p%�C�uH 8�I�b�х� ߆0;AGQ�t�:t҂*R�B����5Z'AV�&d����K7Ji�ȓ˰!�IW��l�Qj7�^Ɇ�b�D�l�!((�֤\
��ȓc��U@�G�t����T�$���m�(!��$C �L��%��(�9�ȓ.�T������`)������ȓ��S�gU9��H�&��[�x�ȓ6̨�cង���Q7-�k}4���POZW�6)F ���F)xp"O���D)BtH��aID�� �q�"O����k�Z	��u)�#j稬82"OR�y�F%S����t� ���"O��p�=c1���ǈ�^����"O޼��-*�� ҡ���\���"OZ���ָU�^�� �ȟ(��͊�"O䰊$j@.K� �ׅ�$�|��"OD�Dm��U��d�#�0�w"O\�`'L��{H�Y�գ�?�Q�"On�Q��؂Y$<�h���;:mA�"Oq�3����}��- �"O~�	@����Lb G�*e~l��3"O���rd�D �{@�P�� P"O*A��OȥoX:�"Q3���C�"O�J�r�X�2�O�����"O$$c��_9>T@��:��4��"O�=��qk������ 8/L�Z"OF��Q�.~�6�!WԌ9(ܼ:a"O&%!����|M"lJD�ۦ$P�T"OjĩE$.A���ظL��|�@"OT|��9MR�b"c��E=L�+�"O�H�񮓯6��H��E;̹B"O�@1�ޚ(��9@,�S'N5��"O���e�9F�ܤS�JX"^�ٻa*O�Y1T	�Kba
���}��y)	�'w�Tѣ�D?8]ڭ�S��<�ޑ��'f"�Ig/њtb-1$E�np\m�
�'&��s ��#w(�f�S�_���	�'d���cԋA��j60T7	C	�'.�C֕B٢������FrB		�'����.�2�r�dK.>���Q�'����6Nͮw�x���S%v��2�'b �����)A��a�NIG�)��'ly�%�ͅs줼S�n�	b�8�'����*)����+�$K	z@��'���H�+�.��8 TI��B6!q�'��@�+<7\��-%A(,E{�'���q�œ?BG����8����'���#��ݵ{�H=+p�X�B���x�'���@�u)���@΃DJ�q�'�j�!C�yG�a[�셞B�ȩ��'���@�ɢL�QcQ\B���S��� �E�$D�yj`�Bc��(xx��{T"OX��a��=3>�)��R!No(��"O@�x��2������MW�@��"O��[�Cѡ}@Uk�$n>T�"O�l@�O��P�����vak "OH��V�c,�c��h��y�"O�CP��c��4�;#���`�"OD���R9"nB��w떈Y|:8�&"O�b�������Z` x�e"O�a2���Y�T�CҨ�!ET��3"O����\����-h1��b�"O�d��	�.�dd�m�
�*p"O�`����tۤ-&�C
�����"O�}���8<pAx ��F�D�6"O440��]3C� GD��3�|�5"O�����DIP��`��d"O��YW��l�a�T�.�xYې"O�����T	�e�3��&\Tlp¥"O4��ꃪn��@�B�F����"O�-�r�W�4������K	1^��z�"O|(�fm��V�6AW�0%4�%"O�R3������!ǰxӈE�c"O������
�z�ՠ�&�F�#"Oj�bs� U�x��o�~��x��"O,�"���>@�$����� ~~e+"O�9�^:(�b�Va3zY��#�"Ob 3eτ�	� a�t�<K$(qQ"O���p K7Z��H�5C��2DT"O��� �E�_R���X6{���X4"OP�+�j]3X*
�`��3��4��"Oh�i]�M���WFP�q�d��"O��B*�)�\�H�l�hH�"O��fhϮ*>,p� <am�5p�"OʱӅ�V'i��J�O�_V�T �"O����2Z|�K � �[�@ �""O2�SƬ�I��`��O�O����7"OfL�UB�%Q�:@1�b@�+����s"O�	*�MVj�q��׋j�޴�@"O�=�e� b��1���_����"O�=��,�%�
�C͂�_��1c"Ot�@`�H���Dk�
�Y""O!12��{����I�y�8��"Or�b�F'uK��qۓh s4��ȓk�����7x���9dN�r
&$�ȓ@)��pm�;���%�г.;~��ȓjhm9�HU�D��Ap�/T��8��ȓr<���ä��F��Y�`e�zهȓ/0��sa�Ia�Qn;ꅇ�&4��(7&M@�	qe�M2*$ҽ��|��}�G��&�z)���O�*��ȓ����9-�)�RŖ=E�r�ȓi�J����o�й�A� �g$��ȓ<$��b��3?`ģ���2#EDՄȓN�B�[��+"��}SU�׬��ȓCe�[G�:]]6�9�_�c\|����BcO�>etT9j���!UVh��#3UA�#�63^<4�H��ȓj��<��@7/8��i��Zk�����a����1LB�m�#$��-f�`������2���`k�9����Ĥ��z"���.а*u���AB������W�L�z�MĆ\ڂ))�-P<Gt��ȓ�����Ȝ�7D�u���� ��@rL3�O	�)�,����Z�D����S�? �4�El^%��1�5�K�
���e"Ojt�7A�3W�<��!�;z�Ѳ"OJ��'B\��i11*�2K��"&"O6�k(^��lC�iY�wH��y��E�D���K�V�"�1D�·�y2N_�B�L(�í[G�,ȓ�'�yR�0�p���DU.	|d&A���yR���P�z�z&�S"}�r�b堆�y".�v��Hۧ�ֺa�]sD@G]�<�al2�ꈚ���.)�]ҥ�}�<�h̰/A��/��p׊��W��a�<���U��h�G�	�t���5��t�<�j�=~J\,�A�Ğ�j4�Wlp�<�d瞽"��#R�v`���p�<�Uf�.>0�B�6^܉�NS�<)`L���z`�Γ[(L�+�Q�<a��	��lɷ%�n0���`NO�<y3�M�i��h塌����eEO�<!�Ay��8���?M�;a!s�<!S!eȆ3���2u�EH�<q#�'LCT�PSU�|�l9��N@�<�VO��ZTȄc�~8Șb��u�<�E�j�����z��0t��t�<᳉S�W��D���]�B=���m�<PB�']Vii�eƉ)�d��c�<Q%1Z����^�t�����A	E�<�w� )�x�	���`*�H�d��e�<�&S2��8ɐkK��4hRi^�<��@��N�t�Cϖ�f4(A�$S�<yeK�Jn6e�o��a�N5��*�t�<�sg�=c�`�'��c�=a�o�<�%�3y�*-�Dτ�6����#��l�<��-C�>Q�JX�n��]�3 �s�<�ӌ�#�P� ��I�tlj�kHU�<a�Ӽp�ذ+��@�1�萫Ӂ�M�<A���O���DD^�v���e�o�<��i%~.�`�ǋ�4{bPk���g�<�v�G8ze:�b���h_^�(�_I�<I���8Z!�ѤX�`+n8xdF�<�P�Q��2����M/��1��-VI�<�nƌ&����큈G� @�Z}�<�7���`9��ˡfQ0+ʰS%B�{�<�1o�D�U�s���P9�9{�k�v�<A�I��8hZh�$��X̮���)WX�<1RK��l���Z2�K�̈���Q�<�⋕{����U��c�:9���U�<y҄�=th�!j�fW��F�`4D�O�<�W�P$b$ք^����aV�^I�<�7�G�*�<0a)�)pnY�BO�D�<��I�6j8t��3J�2�����@�<�3�Bj�zͲ����*M��Dh�~�<)6�" �V��"-ON�!�À|�<YSN�>�V��	ؐ`5>�q�kSz�<��(X�Kyl��ve�"�F�+��vx���'LD+1B���a2U��i��d%O���u�~R�"�ܞ����"O ���A[>��X`�DK�{�La��"O�A7C��}�D���D	U�� ��"Ol��� o|����B�R�|T@�"OВ���3ZJ�h���7x�x��"O&��m��c&Nb�� �"O� 8��� (j�|Ç䒽pC�d(�"O�P)�l\��J��7ߠf���8S"O�,���!���a��3 �LI�"O� ��*w`з,�Ā:�D}�
���"O����Nɼl�������E��S0"O��b OԿ4���a��܆&��9��"O��p� �w[�`��fҼS��=��"O����I��$	h%�랖D~���%"O|�X� ΰZ�� �C
jN؂7"O�9�
S=k����d*�Ch�|P�"On�y���3B�P�Hu��}(��"O~���)œx�.q[�	E�m�"OY8��	,J��PfߋX�e��"O�u��H�(��a�ܳ��("O(�!�&�6�3$�0i�؀��"O����$\���t���;�"O8�ã�+|�L�*���g�2�
�"O@a�vHc|�dC3��|�h�S "O���6![�g삡�$�&���"O���'D_� �WD0A!��z�"OD8�1�Q�!,�TB�$<�L��"O,��^�K��L8�&O�B�09"O~i0D�"�ZX�ͬ%��$�w"Oj�R�k_�
]y��X�U��0�"O��R��9x�t���mI!I���U"ONA[%iEo��t����F�0e�t"O��4��uD��	8*�Ќ+�"O8xp�G�^��uږ�\#�*�J�"O�<kQ�ǒ&����A.^����"O��@4�Z41F��p@R P ]� "O�0J�$��f*T�ϓ.Cab�S"Oz�P��� wΪ��mΝ����"O����ʰ;2�ē��I�߼�1�"O
0��D�5��������c0`��"O���g�dNԴ	0��F'D|�"O��C'��su"�B�Ȑ>E�}���D(LO�YQ#@�	R`���OL�~��pI2"O����\3$I�yXh�f"O>�86��L��xKfΔ�_Z ��"O��p��||<���9iC~�S�"O4��I��"$��l�>O*��� "O21�P(8�rt�LҰ5z�A"O��A"�Y�T��@ ��-qX@Qw"O����홻%�Α)�(�̄$#"O�	� � �BZ�g��d%
�"O�Y�
�8b`XR�o����!��"Oꉺ���BC:IN���uH��|�!�$���`u����={B�h:���!��ğ��q�.T".�=��'_vz�y��'�1O��p�� /�U�5�?pQ���"O,�**��l# �85�I�(J�k'"O�d�D�m7p�����O=D�)g"ODLi��ЗA��UJ�8_�ԡ �"O􈈆!�@�V�����y��"O�LS��J]b���f�lp��I�"O�Jq	�.i�r�`��n=�I矰�	çrwR�Z�!�i[���G"Ht�ȓ]T���\�"�T%#�E]�^h��*�~%��H1DD�q�Ӌ���ȓ?���TJ(
�.�Ag��+�ʐ�ȓI&���C+|���x�$ɉ�p��ȓC@`R��}�"�
 �̯J`��ȓIW��7�LY-��{SL�@�0��NNl�j��2G��	q!I �t��Wԍ���?ٴ4`�%��!��ȓt��k�cUv���OU0�z���}oj�"�拍��S��Lc/Ć�S�? l��5�\?�!J`HYgܽ�"O>% �b|���  IN��"O.���п7҄�SL[8 />�q&"Ox%A�#κ'e�]��N.X&�m�"O0GD�.�t}hւ,X�+�"O< �s�W)�جw��k`b��'"Ou2�o[�\�D)�gU
\U�� "O�Hx�ϋ!V�N�B2G^�{��v"O� R�c��{��P��&U4��"OƝ٠"U,I@ �PB1n+���s"O�����	/6�;�B	_"|��"O��U��,�	إ��9�T�0"O`�S �Bs8���DJA(�"O�e���B�m��|��@�y�n��w"O:�����
.����!J�ē5"O�TA���$�|�*BׄAН�"O��ub�R0�};�@C'�b��"Ov`"�,C�h���@���Je��T"O�<If���%0$X,W�`�)�"O�y{�/�Nr��A<y��t��"OTH���=�l�ʦ8���z`"O�����%�Z� >9ҒU�g"O>�Z�Ǝ�W��@���:�B�2B"O�q�5�[
~�l�o��a�i�"O�P�ii�J��-�t��I��"O2�b��]t��X���M�W"O�6�P�k���z� � h�~���"O�d(	??aDٳ�P>Y�>a��"O��X���(�lh��،s����"O&�vI`; ���"ĥy>�m�"O\����[��<��!ޮN/0��%"Ot�4�/}t�z�� W�HI�4"Ota�s@͔=R�	Ǭ˨#�$�j�"O:�q�횋P�E�ԋO�S5V���"O�t�����Q8�%`*O b���"O��kM��0���2S��0la�|��"O�9J	޷T�
���ac�i��"O
��e��G�ةq���2va\T�"O�Lx�N%t�D0#�֚"�(�"O�,�C�0����b�,I���"O<�āU�A'0�:Adçy�`��p"O2�aɂ�^��[f۷NYf�i�"OȰ��$O�<ĔAS���-��u�g"O�,�B�)�2R#�.��hiw"O�������)�7�U5-��Å\�T�IK�S�O��\@� dB��qgX@+.%`�'���`��оRi�8Х,�=�2uK�'6�=b Nؒh�E��O@��;�'C��bBN�T����\i�'����,�Z����#M��6ܢ�'5����A�.7ɰycE h�|8�'�RAGӏނ	�2�ŚtQ��Z/O@��)�)ʧ�B���ΧYT�\���]1�\��`�L�¢
*(�)��#!�\����Ar&K>C�f0Ɂ��8a��ȓ2�(9w�D3mvI�]�UxL��ȓ7��X�e�.����3O�J�d��ȓ 醨��))}�� b�#4�ȓ|d
2�ġ:L\d�t#�$t��a�����1Vz�@ �I�g;�|�� ���j����Z�.�#���)���0��I�5C�T�S���i�l���.�X@�򇉅n�N��e��%je"T��\����:�� ��"byj%��S�? �y0��]�N���Y��3jq����"O��p��p��pJTA)k@����"Oa�	[�L����t�� \949`'"O%�C21Ը�Ue�8s���"O昀� �i�`h���!H
�"O��i6!)ekL�F�Ն)��
�"O$}�512��C�X�x�"O0	g�<~n���`������'o^��Rl	�<�݈��Z�ER$�'Ђ�Z2�� %��T���U';Ҭ|�
�'�t�ä���P@^�9�
��g�2�:�'�6�P��W������oM�S���'5j\: '�6[\��q@�$��Q
�'8��*EC�#��ps�,��t�U0
�'d�esv#�R*
�1/��a����	�'� 0�	�<Q��a�0h:	{
�'Gb��U����|%i�	ۦg�e�	�'X��+X�jy)��C�k���G��`�<�q&��|�d��̄/ar��w�`�<��0��@��,EK�q��I�Y�<&B��6EtM:3��#u�X}�֭�O�<ɗ��8V��BL��}*ZQ �g�<I4˕�>�`� V�V9�eA�^�<�e-td�(�7��^R~$��+b�<!�9�J���R/k����/�u�<q�gȣg��Z��7��{�TG�<!$M� )J��7�LZ8�q�Jh�<Y��m���郞��u��m�< dY
.���՛v��"���`�<���T�k��xVd�C=h�z���[�<Q5�
6-~B�&����dB5�DP�<	�L���p���_@��r'&
u�<Y"O��'�p��ǖ@�䙥��i�<q���VQ��C!7�v�Y�UJ�<��U�j��J���b�(؋#@I�<���P]�ڔ*��ܲEQh\e�Nx��'?,�(A0�P����L�t��	�'�:(!�*1�^]���L�3 ^H*�'d��j�%�	-�d��p �~���'� ����\�ntc��_6�L�
�'�@�!�d��	�4�i'�F8.�F���'t��%�A!~�J�f*�= >��	�'{���,Y�?�P��2m����t�	���'q�}��-U�{�Z� �jQ��:	�'e<	����%>��������'���R�ѺH�r٣R���߂���'$�+���"K���pO�#un`��'��쁣��
K�2Q����!V����'p�y��B�3d�-��%�* "�xi�'�%Y'h�(@���kR����бr����F&L���qf˚M@l�b	�I�!�d�>w/.�㔦J�tD6�"�d�L�!�@e�Y���8�1��
�g�!�d�Q �%������g�&_[!�$[�9t���_8i�V	��b� 1!�qt�4:TW�U}^�
�AG,# !�<, Q%@�@l�����F�]k!�A!��	�a��wX�m$ �`!�d�SH��3�o�)BFpcc�݌Q!�d0g�QX��@�E�Y��o�?H�!�$�#"�2�ISbB�u�,8�h�%T�!�W�A/�=��مg�j��:&�!�i�jYZ�D�� ����B5�!��Օwa6��2�C�V�z䇔�5�!�� �᳗b��5ߒ0!��	�HQb�"O�-�C��;J^Y��	�6uԴ��|��'`az2݋v,�(j`L#S)p��"`��yr�Q�:���H���`�1�F���ybg�L��Q`��]��0�@�yB�."q�[��A-���k�i��y�ᗃz�%D��y��Q�:�y�ʂ8621��J�=qo�)������OT"~b2���K���"e�,v7LP8RC�K���0=�di�:Pڈ	�"פO�HX�g�G�<q���^4�� ��"���P�B�<�!I�P�8���5x����z�<����r�`�u�H�H�@Tq�<�M˕R1�9C�냒QK��v�R�<q�,:(l�h� �3��0p��IJ��?�	�'6��ɰ��B 56\�^�VA�u�ȓ��h)�EX�k���k��H:l����Q��ab&g�HR<�9@@�l{PU��z�P��J�W�8��c�<@�z���J%`������(����|���ȓA2ĉQ�>&�pR��2�:9��a̓2�B��n��^`�Y�Bl��s���G"�S

��4�֛�Nu��!0ԨC��4A��bG<k?}S��Ò;��C�Ʉ����hU�`�1�6�O��JB��<U���Zf#��)JDK E��
�FB�I�zx�} ��(5v�hn	�c�0B�ɸP�$i���@4A@�j3�\W�ȣ?q��)Zݶ5`��� xr��v&�"�ў\��	�h��@��"��e��Y��H�C�I �ιc�E�K&�� �K7 TLC�I/�␙EH 7L��U�E,N91 C�I8g�ʀ�+n8�%JᏜ�C��2A����w+��G<��iwꎲL$C�I <>�� ��ɿ]R��gE�����d*�)wHh #(��#�8}�"���4B��H !&�����4#�@'��F{���G��U�
e�DBG�������yr��L%��j�W�y�t`���ybAA�.���9C,6�x���OX7�y"�@0\$4������&FB�Q��y�&@j������JG�$B��S��yRf]�l��j��F�@# 9䎏��y�)F-(E�Wh�9d�RC˝0�y2��m`�i��s��1�@ŜpI!����Х2��P�V�����I1!�Ğ0L���A��޼>��qR��#00!��&:b�Kdș�l�8,r�&ײ*!���]U�u���� 
u2L���; q!򤟦j�F)�4k	�+c��g#I�:�!��P�pi�a!�*U^�ab�*�!�DǑP��(qb��o:������~x!�$ԭA�R�z���@1��ի�rh!�D
�\�D�!��*�Ä�
]!�d��aͨ9�����F�I�Ĥ�(p!�d�=�vթ��d' ���eD!�D��=���#���rg�}�g�!�$�'s�ࠃ-H8v�%���!�
*&�4��k��a�@�;!�$#p��0hС,w\���b�5�!�$؈��D[R)��|S��^!�D�^FҥJ�Ê*"T��.� .�!�$X�t�L���iǷR"dU��ݖ{!��DRm �h��jb�\R�� t�!�� F��eG�]��+r�P�BߺQ1�|r�)��;9C|eb����}Ė1B�N�=Pq�B䉡;L~�Kw�Ʌ$����&U�b�rC䉍>�4ɑ�b�h�A�D�h8>C�.6ta@�8W(��2.TD�JB䉳OW0a��O۩b�I��b��H}�C䉬,�%���_ݞ��Ev�C�	�
�n��%#%W��sD����B�	�>�~ɓT���,����H*B�	;��4��1QɢȰaKD�2�bC�	�@|d8b���M�dI� ��B�I���Ű��@�i�((�%!��_HC��> ��`c`�v�(|��e�?@�dC�Ɉ>2|�A���-W�8S��G,Z C�	�1W�0$퍫]]D�d�<;hC�I�_��8UK'Z9\!�w쑝Q��B䉒,M:����O�Y-D�d�B��� ɝ���E(�p�!�"O ܓ2��,Nɮ�	�f���Ca"O������6�L�#��o�ʵ�T"O�:� L�s���9Ab��v�"O`���e(Ǣ ���Y�#%���"O*�����p<x Y���!��`"O��CM�R�.mbBBW~826"O�Up�(��
1 ų�(zYj�٧"O��!��q������qQ��'"O�#��J(lb�j�)?=x@"Oj��GhO����J�wN�Y�"O�d ���+��ݪ���vM��h3"O�%hf���5�6D��M_�>���Kf"O�YKV�-4�Z|a@ύ(%���`#"O�Z�Æ5�pq �����L��y�N�&n��hs�Y�5@00���!�yR%o�U����.��h�Ȕ��yb F���P�X/Q�*�RC���yR�O�ѣߵ7m���n	�?��ȓj�l�۶�?z��}k&ÒGP��ȓ�|��$��5V�I��N�P-�܅ȓ7�*��(�i��튑˓3+¸��ȓsن8��׆G����E΃-�<5�ȓ�|�)�#�R�"!д�]�f�4��ȓ4��3�-�B�}1�ȜHVDH���t���A],�$=c�ѠS�Ņȓ#��Y���I�NRTc����fQN-�ȓ^�b�	�lQ%<�"��p��E�d�ȓE ��
��XP'V�q2� 9x5�����l_&=a�t�ӱn�0ͅȓn{����C��$C�
!���ȓ�T{�瑒2�l��.60\�ȓjt|�gP5
�����pS�p�ȓ)��P����]3�@nRY�ȓ��@���;J�0;#��/hB��ȓ4ƜeK����/�4��Ƣڭf}!�d�20:�k�F�[����E��/!�B�kq"5*����(�@yZ�KM�!򄈱�$�JP�ݯhu�al�	!�d�9mԖ;oO��eHG*	16�!���.-�m�L�$& ��)_�*�!���=,qn�����{|��G�ڟi!�$ܫ,u8�:b�Ѿ���P"�,-!�ǌ�
I�7��<|�4��Вtm!�,:�*qm٧/�|��ʞc!�ɇ;�ҕ+"� B�8Hҩ�<a!��(V�BŨS��X��C��!�� �Ũ�kɚ+b���6�Ӡ8M<MYW"O@-�Eh��GKv9�rG�2נ���"O��i�A�~H�po�����U"O�	���U�� [�+��<��#"OJ���B�x���j�
v�,a3"O�@�D@؎h��p��RchP�@�"O��w�Eb�xDk�K��;^raH�"O9�S��TՖus�HB�~'�u;s"O��kpH�(<8�ၰ�]�I!�I�&"O8-�嬅d_&I"�e��8���Q"O�,[%	� �!�V���H�x�"ON�c�	�vt�aI�0F�p�4"Or�#v�ӸVa�h��4-��P"O��ÀFO7j�qJa��C"`��6"O�\��I�5�~�� H#C�d �"OD5)�(C#a�J�Z�'��{IV1a"O(Y�Ƣ�5b"�e(� `���"OZ�SKX�Z�L�a��Wۖ"O��Վ��!.�"v��=~��Y#"O���G���X*w�3n7\��T"O��B���72h�]��)��J��k"O��ӲSt�&	��(
�cb"O �Y����L�"I�3�^�S�d�QQ"OBM�Ph���)r�ֳ%-|�P$"O���Q��r0Ec��� �|@"O��p�o�!F��Q��["d��"O��sda��%5~�`U,iV��z�"O:	�Ɗ�8�dI�#f����("O
�	���PW
�2a�2��$"OH�J��
3����hI7O����"O�m��LtP�Q�Ι�Ol,�&"O*@� *��@��y��5�"O&�#���u��Y��?�:��"OސZ�I�8=�ԐR1S�c��I�"OJ-r�䇓HV��S�(����[�"OL9�J	�<���sG�$�0x�"OV�@�d��4p�#���hն��D"OPq֬B�G
��T��I-�	Y�"OF�"� �5r�b���fܬӷ"OĴ+$F�f�*B�T�M��z�"OzyX�遛b��+u�����"O�T{�O� ����G1Wt0�"OzH(`�'xl)��_�n>��#"Od��!�3�0�� g��u*��[S"OhI"� #D�p91���h�1ZW"On���V�r�d��hȝ(�vT�"O�]�4��X�,���fٝ~�Dܘ�"O��y��ٿ#.t|ʧˊ;*T:�:"OL�C��,�LT�mְgO��"O��4d���M��,Ǻ2O\Y��"O����W ,D��
C�s���+�"O� ��,DE\d���JT����"O���dE� p ��V��3r5��'U����H�\"8�W焊G.�"�'��;զ� qu.��Z�j�6a��']�E�#�I�h�<qc�� ?\M��'�v�wr��[�a�-B��e��'�V�)�咇�L�iT8<*�Ը�'$f�A򨃤y׬EA��1-��L��'H*�k�j�2Cl8�ʐl��+����'����P N!�00�*Y�[	�'!��8��
/`��2�� :M���'匕�. ����-"R.��"O¨r�'8b@�y��Ǒ
o)�e"O�  �8���a��m�fm��&Er���"O����e�z���8>jZR"O�P��k��t��cf׉G�x��"O$ �g,E5/N���E� ax�"O�Ay"�B�gߞ�sd��RE�@A"O����J��<�h�JtC0JC�Hk "O�T�`E�S�4�b��S>H3a"O�}�� T�D��騐����M���"D��C�`2K������`���3D��ƏZ��H���G�����*3D��4AŏJ�"P�H��K
�Qx4�2D�����/�
Q������B��/D�|����P��e�Z-@g��h �/D��e.ڵh��LcF�� G�4i�f�-D�(y�OZ8<�zq�U#�$��1D���� 12�\�k�`Q(���e,D�$���8z���a�S
����(D���l�|3fK��l[�Hj��!D�����R^¶���%> �����#D���qkA�ل�C�(M1�$����7D�@�#�8q��,
7��:M�����/9D� �5���]���pǆah��9�j7D������%"�̹7�Q]xHqAIb�<�C��4KO����	ژh��嘥�IX�<�dK��d,��tǜQT�MТ�K�<��"Q�l��8fbN�{ɂ��cŖI�<Ag��������ܾ!O�aA1dC�<��fJ9����*��I� !@�A�<���3�xx���]��]� ��t�<��KM�=n	(��X4�셁D��m�<���A?p���8�������`�FA�<��)N�V�nY( ��;H�`Q	�A|�<��סFDv��@!�Y�||q�)t�<���#$WH�PԎZ7w"�9�t��m�<�1d��[z��33��3 ��1��Z_�<i"�Ȗx�bݢ�hX�'>� ��^�<	4N�n.���[�0�3��Z�<y�[58�p0��_�:��SG�Z�<釉*k��ɓH��8\AYcG�X�<1�@~,ze{�Q�Dw �j5�X�<���ԪNS�0� ��&,��i*p�RQ�<���9Ąl��`	";2���b�<���-�*ɂ��8�(��Da�<���V:v�N"���\���`�r�<Q��U�=@!�R/�G1T<��cIo�<�SfX1_�t��$�!��aE-Hl�<yA��2"�h]�Sh���ܙз�A�<A($E�JT�6���9>�Ҩ�t�<9�!�0Ĭ���}%�蔌Ae�<p$�(taPo�WR�YHԯ�c�<q�j��?]d�!@��8�#��Ut�<QuCM/xn�:����B׸ZrBنȓ4A�¯T�$E��Gɝ���ц�=�����m����F�%*��݇�i��A��HE����b�j}��S�������HT�֖�<�ȓ�X}ÄK�.��V�ۑ ����ȓa�B���i	�z��ro��\&���ȓ��\@�ΐK��岷�P����ȓ@�~-��%P��Ja�R%�"���J+ � �\�6��cI 3x ń�L����L�#�&� ֹb�&�ȓm���Q(�7y��<�Ңa!2kKG�<!���ް���ܸa�rQ
��<� L�3��\�N�6�0���
@�*���"O�\	��T!'wv=�6�S�-甬��"O���T<B���$I;ֲ��"O�qQ����.�4 �Ï�K�=C"O��S a]�`}�QJ������"O�}�qg��H��t�#m^5k�F�Q"Oh�86C+%B��*BϳYE<0��"O`hHa�F+M��G��� >rX"O��y�,rI�.�'6,�B�"OPu��G&��{�C����"O�8R��< ���C /��&�T�`""O��JtL�QJ���sC�i�B��"O���F!DV��1)�!A3i��
�"O\�`5䔉S��d�b��A�t�Z"O`D�s�  �<�#Qg*��"O�}���C�OϞ���AF
\T�aP�"O�:iƲi��˳.[�L��\Z�"O,����
U_�di D,�άZ0"O41{7��=h��\�v��+M�����"O����'ބX*:l�R@7nLMB�"O���P�#"�pCD.O�@�az�"Ok�*�T ���,�(`� �"O�0S�쀑*���l�)!��3F"O@}:�����(�j�"�X��"OZ�{n
'?�D��3�:���z"On��T�X�M��<�2�H*�ZA� "O\T(&��OA��îP�sr��8""O��	P�Ln"J\���> ~�L�!"O��j�WfT4 �/�Cw���"O��	h�d�d��\q@��"Ov�{�l��б��o´e"O���)X�G,d��&�ΟCC�i	�"O� :RO�@_,q�Ǌ)d#*�Ї"Ojh��Ę��M�G�;��ӕ"O��r��l6��@O,�� �"O
LP��e�<D@��O�I:6�"O45Ѕ,g�	�1@\! ��� "O�@yU&
=�H�6	C%-�ŉ�"O�P�M�8 (�k��L�G����yB 	�{��k&n�>i�ⳇ���yL:Q�V�X�M)`�@����8�y��\+%�\���]A�q9Gj΍�y�/���>4`#.�V�����n�'�y�aĘx�����B�K^b}���y�MG<l��ٺ����7 ���ì�yB.S�"`~m�2�A�'^h(B��y�c�Jp �V�ܣ@�)�w`Q�y�˓X�|�`*i囶D\�y2+����`kC�HfB(�	?�y�cͷSF���$B�\�������y"hZs��86G�4Qh�$(6��y���2%1ܵYV��Q��p���y�D�PY��1q�F:r0���ǋ ��yr��pv�`�G�ΘcH�j���y�n�+����_�	�V�CF�Ȱ�y��4y\!��/�t 􀸶�ِ�y��V!+,���M(�j�UHO��yR�2�ޙ����M��0(O��yr�ɥn0�2 �ģ%6 �CJ�y�I��P�yO��V�@�P��y�ؖ6�je����V�V�IQ��?�yr�S%{�x���Fz̈��C��8�y"F'F<�d��	ۛx��+�Ɛ��yBoW��ָj ��s��Њ��[��y
� �9A���lm(�"R�75�V"O���b�
\�e!���/2���"O P�2��3������y0 ��D"O�J��U>/N���2,T��c"OB0"|P�8�I�$�����"O.�#%L9y쑢�a�x�� p�"O"u�"	�W��qb�5f���""O �Y)P</�\���}`U�B"OT�p$Ӯ$T���Hp]�I�7"OB�2U(�/3	t�1g(��L�j"OĄp�GN%���7�˟i�(�"O�dQ�\�D�P$8���&DX�0"ON`���ȈR�l%���q��� "Oੁ���%'���jg-��z~�s"O�{Ť�.+bR���KN	�\�
�"O���`�ܠ���{Ɗ��z�|�;g"O��C��;a���ĩT��8�"O��ZNV�IE�u�%�{{4�@"O����!��K���7@Y�0��"Ot��gM���9cK�J����"Or�#��V$��8;q�V�}��0�"O��&�Ӫ}5��@C����"O�qɢ+��f��t��*x�Q�"O:ɚ��W*o&�!8!�Nr^� "O&��1���&�����4�>��"Ot�A���BA"�3�6A�P�"O�嫓A�[�������s�T�a!"O�$v`P�Fm�`.������"ONi��j˧y�Vŉ0(�Q��p�"OҔ�1?hd��'H�&v�>��"Oր�F��Z�z�S�蝰0���C�"O�)���eu��*��|�bT"O^��1�[>Z�X���*P���Ec`"O�`���JL�� 8n��L a"O�<�F���F���j�3�(�!"O���AG^�Wc�ˡIǊ6�h	�2"O&AP��
.mP�9 k^�t�5��"O�%�����[;~490����z-�g"O��cqA�p$�8'`�=,����P"O��`�T�=~~�#�nWC�DP�"Ox"�Ƴ&�RkI� ��U�7"O|H��	�	:�t�8SJ<~|yb�"O�p��4,Y(,@�	���is�"O^��6�I-�b��k�}��	� "ObyQ-S2�$M�$
S,���0"OD����u�Р 	� Y����"O�@Q�NݮQ�ҡ��D�B��<�"O$��ڸ|}�Y	Ą�	c�p
�"Ovc�Z�l~�	w�E�Z��"O��fa׺n\��P� 
4O�a��"Ob!K�����\4�y$y��"O>��W�(6P-0�ȊA#x�f"O��z5O��[�����Q�D+S"O��b��w�y1�/� �@���"OH� э~��Y�Go�?^@���"O�!Aō�O↼��]�r��"O"{��&�`���];(7�՘�"O�A�@��s�j� �_A�yj�"O���򥗦#��Q�DH�[2�]+�"OΨ`A��!%��1BÒ�*x��5"O�!���#J�	�C�
����"OV)FL�0��8CU���V^�:�"O8�Yp-߰� ���r��P�"O�-�T�:���m��b����5"O� �HqQ(�9k0�qZ��	:�i�"O0���MW�t>�JCM�c��MXV"O�T�b��(7>�k1�,	�h���"Oҵ��ӅFO�(
�㕋\�} "OjD�r���h7��եL�"�@u�a"O"i�'(�6ڪ��n[3qў���"OV}sv��;Nn�ڱ��:�0�{ "O�,�iب%\�x �g�?,���"OD��iG�$`kw��W�PH�E"O�9�B�^�&!A�A�n�Ka"O�� �@C�$���o�RO��"O�i����0Ce����hs�h�+2"O2��(R�~�Aᐭ�7ۜ`h�"O�A�� �Q��{b���(��"OT:�ё'���b�k�;y�0��"OP	D�Gˎ�h7J��pLu��"Oz��fI�B�L����Q �}��"O�I���c�� �bIV�:�Y�"O>\[Q��`�~1�*G�V��tڤ"O���҉DN��3�*K`aZ	��"O4ub��ǡH&�E�C�ܿ(�
y�"O.��5/ ,:��S�³T�|�zU"O�ɲ �T�]��K3Q��"O,� ���BG�:UdM��㛝M�!��Q�e�)��2<r����!����,bqgI�V"�9�UA@�)�!�@�z�����."�<�QV�\�fF!�"sr0	WE�e��A���&,!򤜎T�,$k��#LlZM�$D�h!�DTi�ɻҨ-u0t@�c	�o!�d���F%�G�!~�(p-�u�!�:��I㋚�$��ݘ
�!��A6x4,�td��tm����2U�!�DK(\1���1�����	J�!�ė*U 	��ᕗ^Ķ8���e�!�D�&�2- '�C�0f%��i��=�!�$��UL!Pc�{�|��)���PyR(�2hX�Ls���oVZt[b��y�K�-Ҥ8���� ^����� ��yҌ�/KW��Ӂ�#Y1Q�R���yBۭ�jԙ1#���^yyb����y�o�(x�F�TjW0��bsB�y	�=P���&��7b�R�U>�y�BϏ3�>Գ��.�@�����3�y��G�^�����J�z1�ᐅ�y�N0
0ir�Q�t�0�
�����y¥A-G_�e�Ǔ�@jU"����yR���Mn]�蕊����m�y�	�n�nDj��T�xϪt�&����y�D,K n0��_��iㅅ���C�ɳ;6+o]J"����=М��'����,��;Q(pk0���a<�-��'~�y���[= ( R�l�V9�
�'V�=J�a���5c�
QǬ8��'��i���0�����J�n{�'�:��@4I�5�ț1�3
�'�̜ia ʔa�j�3%A>�L83	�'�� �/3����`K?Nꈫ�'�j�b�ǚ�a"� ���=X���
�'X��j�>��P)�$��|h����'� �çh(}�|���ʿ��9�'��X�Gc�"<� �@Ջ,%@��6�\,0��
v{R�{WFMx�t���A�S.Ze������
9Tԅ�S�? ��� P03�V�Y�ʥ~ȢD"O�]Y�>Cf�="ֆ�,��9q"O�U�d�'4Z����W��aI�"O~�fiH�A�����?4V$�aG"O|qiT��~l�Y�D��)@v�&"O�(�F�2*��lY���
GL
��*O�Е��h�\�2!�����
�' t�Ϙ�Bb�R�G���{�'�F5���TG+���Wn�D��EH�'@h�ȝ2�}�PKM�oԎu��'�㍐�j���V���a�L@�'t��S���0�^/X�ੇ�=�z܉A��_�� 9�)̓\8���ȓe�ĳ��ݑl�<J7�&k}� ��H��} Ǭ�?+�.4HS��1$���JO�(ɥE�a���a! �B�)��{�kƎ��@��F(��v� �ȓ:7I�D)?Ρ�lV�3���N���9�+� +�6\ G�
ݜ���7}���O	�AA,�Ud!��@$��H��|�ׯ�*���`�ް�B�É�h-@�={��ȓz�� ��2N��ȓ4�K�7,�i�ȓ'>�X��&�.��P�7�(I�ȓ/�,�:6ףg���#w,ӈD��H��#;�8�V�ɲA�sá�WFE�ȓ$���FB��>~l�ȓ%�RE�wk��t����@&ي4 F�ȓ#\ �#/T�� ��ʚ�=�޸��M��Sv�- #���Eك&�0��ȓ2�b����]�Hf@�k�ޣ:'t-��TT��2���@�"mN�ϪلȓdN��'e�6)D��B`��n�<�ȓV�Py2�@%њ��Z�&X�ȓV���H䀅'��⡦Bv�&��ȓ@&��e�
�E��D�ԅ�i�b̈́ȓ���[��U�vפy+D��a��M��wܱ����	x�����	�lhD-�ȓ6��zRh�i&P�
)���ȓ����ȉ�>�d�'AZ�!��l�ȓq������7�PAx�aF �q�ȓo���qM�4i`�mȥU�VT�ȓs�FH�ŬC�[��҃�|�p��PU�U����%�ԉ�K�(�ȓ{EN��Bo�%����b�ԅ<�@�ȓ?��p��/�aB
09!� �:����z^e���pNl�(G�P�V��ȓq�0 #Տע4�����]�@���$����
�$�3�mQ�6�����7,.�P gC�:� � �f	�Wo���:Z�x;�� "
�@1@��ދJ��I��t��a%�{�8 `�/e���ȓK��1����>�\ccL�S����,�Ry����9j\�����[X�L��x����#��<1ؔ�#B�ftZy��g6��glD�&�����iiL��ȓL��-��I$;�2��ӧ�1H�8<�ȓ8��,�&m]9Y��{7鋖Tr�<�ȓ�|#��=R~�!��̝'��)��&x��&kϛ�n	i���7��ņ�jb(W�q��_`���ȓD�\�����	KO��	�J��XXY�ȓ|A�X�&
(	r�
DK�+TH��g���c��d���"�)NC�)� H�Cdin���ʇ@ƚa"���"OxM�E&Z���ŠL y�]�"O�|�7��.z�`�`�C���"O�4� \�s��Rn���"O�M���źdp*����>/YĒ"O(L@�o%r*TYc��.K��j"O���w)w� �	��ݕvWʬS�"O��	��6z�Ljn,(3Rp��"O��4�_0}yJ�X�M�]�"Op��ԨV�7�6 ��
���K�"Oxx���ʤ��"C�<d��d�v"O�XS� /;r��t�RHan�b�"O��0�zD@����8b�����"Oha�7ʀr��Q��c�5�Ї"O��3p)�	>��V��	v6�2A"O�y豍ƓEk"���HT�kKr<k"O
��玨~Z2&� K,�%�"O:\ZB��	={$��"&�D� "O̫�Gk1P���n�"1l��'"Ov� Í�}2���  y�^��"O
E�I\�p�|�R�"�2p��"O�0�@D���u�P�z|B�"Od�����#���`�\�
���1"O������%ML���-�f�D�0"O�����\�f`C�e
�Ph}3v"O��a�!�5[�$5�%���d�K"O���E�B�\8:�8�ҮO�!��� �zQT�V�mN�ř��%$�!��6i�5`%ɔ*Lڑ�"��M!�dC-!6h`�2�*���nĊP�!�$Y�5�x���VϜ|㴇��^$!���(<"���`�8
�E��G�T!�H*o�j� Ì^�;��<��Ǖ�b!�7O�h��bV��zi�A�p"!�D��]�p!�H����$�s!�d�#=��;EF��U�8�p��K8	!��?%J�ɷ&��tg���虄n�!򤁯7-��!c�X���>�!�D�hC��#���4 �y/Z�(�!�$�	��k���s�t�I�!򄍧.0�Ei�A�cj�� ��^�!�$�2]��C�MV2HR��s�σ1�!�� �aN"��$GW?�퓐CE��!�dI�H��!��ܣqB�I�#�g�!򤅧\��тӮ0W��%¡��+8�!�dMH&�2'�
�Z2U� L�n~!��֋	xt�b�C�ww��(p�$2w!�dC����PWIi�X� �H�,w!�$I�"�z�x�	 R�X-�al!���Ȥl��#����'[H!�䝬=��q�m72�P�0�O��x-!�$��j3���B�� B��j�<��N��k�ŉ�f�:��.���ȓu�������r1��+~�*�ȓ%[.C��(�D�"� *-�`���th8�J�˘�f:�*��@?9C���A��=+�F�9ڎ���7T�B5��@�R�����Vd$�+pV����dUf0���9�0L����N�ܥ��-�d�t�ӇWv��ۤ@X��2-�� �@@�gI�L�J�I*�LV��ȓ ~J��R7U^�9䞼����a�L1�`�-���r�ݠe�\��
��j �øG���j�"^��Ȇ�S�? �=���� w��\��:��(�"Ol� ��;gj��#Oэ�&�P�"O�"UA���r�C��|���"OPD���� 6)2���U�4�A2�"OD��@/]"<�"��6�ˏ1 �ʴ"OH�yA�L�$��f#��B2 !�"Ol96(}�2���#M�� 
�"OZqɠeF�9��[�,ܪ#�jK�"O��d����h7&^9!U�
�"O��"���ifB������K`�rS"O2�$K^'1����}B^��"O���G&@=����±)b !�"Oz�
r��x<��q��f	l`��"O�bk@�^�na����,*��9�#"O��ؑ��d)�B����t��f"Of��5�Y��`���#*yXa���?D�h�@A�$*�h�3i�.-� K*D�\���5�p'ҝ)�6��'�&D��R��EN=���c�ì�(��!D� �Ѕ�g���BGhB5����!�>D��:gA�OLT�DdV�U���
P�;D� ��	�&gP�C�O<B�\M���9D��Z�/�ѸT;� �<�~�h@�8D�:��ߣP�^�q"��*v�p��G<D� ��IC�s��$("����<���$D��+�AE� t��(ǥh��z�f8D��s���S���s�:Fx�p�#<D����L�S5AH�o��&����9D�<2'$�D��D�����b%D��i2�H^%���G� �ɤ���7D�H3R����V ��L� px]�0�4D�ء�ر�6m�#I�>f9�w�0D�P��G k 0�	F������;D�����y]�ah�1V���$.D���Ȃ�Nd:|��aA>�d[!� D���C�� k�@q�dA�ckhQ$T��r@�Ymmh�9�-Q��8�a�"O�]��m�C�*�@&�E<�0���"O�<�o�&L�B�KS%˹8c,��'�(]"�b�-V��a#�P'iL �����!����-�4>htER�H !�!�D�3/�DC��|G0A26#�1�!��V�^&Д[�͟mMLu �i�){!�G�����z$vx�&�H�!�1 ɡbә�4��!�DK0~9N��A�ث6-��A����!�D��
,+wl�,SPa����9�!���k�"urF�	�L	�d��6*!��XlN�SQ!c�h(i��W!��6庵�d!F�p�^�z��Y,d�!�dS
��[rW<���H�H�+�!�䚥N�z�'$?G|$�A�Q�!�D�?C��C�,Ɲ!�����a��!�d�-#:����-(ʮd��C�:+�!��$An�ȃ [1{�����Q/Za!��W�/B00n m����!nİv�!����=D*�"��7(�����!���z��9yu���������5�!�$FzN�M2q�I.W4%y�ϑ�
L!�ė-'�.)����AD!��	�'�����ԬM"�p�"a��R �3�'�����"v��e�"k�U5����'pԁG:=���AG�ZM$�ϓ<��ag�V��D&y���$	�e'��Q
�qs!�d�?0�����=s�ء�j_�1��'x�\���?	`��� ¤��.�b��tp�f�{�2�Yr"Oڸ�j�((4�
��t��SPbͺ)�B�,�(�9�`$�3��ۗ{2QU�?MH��A��T�E�!���y��2�PR�x�yeÉ�A|Z�:˚� �5�XX��(")�4�HX��G!F��ط�(�l�ttᥓ�A]�)��jb7Ÿ;��@�0�2. }x�!p�<9Dh4`h`����`�sy�ᙇwPh�#'���i\
���(���sM�x��9�!��8yg�`X�kA801�EC��(u� ���
���3#޵Wq
�:�Y>�<�Q���ű@��+��Lkc�UHX����F�0F�ɓ	�6�]%
֣�x�Z�I[���0[@y9E�Vc8�:F��� �n{��!��Q�$�q`P�3|4��Q`D*it�=�Q ����ƅ�m�}��K�+�aҴ�y�X��z5:Ƨ�
���!3���I�"`{T�	1	Q=Lxu r�l��ygA�h�(y��צ�~Ma�.�yb�Fo���*�e�}����BX+�|���kX*AP��W��2$��Z��o���Fy�D_P��\k K�pǾM9ҀS���=GL�'.�7$��U�:A����v2Z��Р�bt���]ݮMr ��a8�	�g��ed���tn�uK�����;�I�Rq�U{�F�����3	�j��0;5G�?�°"�m�:I��ƑP�qҮ<D�4J ��p���I�MK!>�ٳAi\����bg�C֪(��iѾ��-j ������@ߙHY䵰"�=4$Q�4�w�<!�.Ҫ�q�#j׉(���g�֮$�6����P>�h�����-{�r�"�Nҫ|��<YքR-xh y&��z�Z�*���i��L�QC�������M�P|+��c@��'�Q�]�p���4U�"\s���:�p>��	7�8�RM��-:2�ã�b�ũaϐ�H��6	U�o�"X�a��I�qQV0I���6y�W���!�$�1\���C�e�,�p�E�H��<�%�^�SU|��2�M�qU�U��0��O�*��;�Z�����8����ɞ:
8D�ȓ|���Y��Cf�\�RaB:q�,1�7)I��* �)�.0�K��ӡ|���aP�"ʓj� qK��ͥYIH�yb��9b+�!���j�|��.��c���JTMA0m~�����<C�(h��
f� �vN�-ւ!��"\X���6nA:�I����	�=�h��K�<�r�F�v�m3� N���謟FAY�R$���@g�6#���D"Opzt�})�!�0+O8�a��v�|  �'��)��D�0@�P�J'§�V��MXa�c�#d�n�(p���6L^C��-�h=�#$��$�nM��4��l�R��=E�s�5-�֘`n�ٺ���N�.:V����#'	P��ӟ��{� ��wj2�9�M�,9��D.� !=�A��@��.A��c��,A�	
�� l ���(��Aѩǒ8Kh	Ex2�-#�hɑ"����Xgh�����ah��oOЄ�B"OH��&j�>���Q��V�{OF�T��)m�2��͍���S��?tR�5�Y[G�\�VM���Kv�<�R��98�N� �EXr��f�p�<9�*ÈJ��X��A��\1AM�q�<3�ސ[�����QQ�t�E�n�<��k=\��)�i�?�`��RC�o�<IM]���yqh���e�A%�d�<��+7~��W&�*8���Dz�<y�	;m��*%a��e�E��`�v�<i����j��+V�!xvB�P��]l�<��Y$n�: a2M�"X��U�� �D�<1ǌ�'ǘ��T	�=��9�	_A�<A�L��:�F�R��W��ܼ�F�B�<S�ױt!��0r ��4�L��M�{�<�Ģ��d�!�Αei>�C7/JL�<�CG�*F1��޽r�4"� O�<q���6eFua����%˕@�l�<��\5?���WI���T[���T�<9�+��d�0�`ې'��H����<9@�ǈg�(�b�ě�88E  ��m�<ѵ$��t�)�:F��DX#��j�<	3���Nu���7�B0MZ ��De�<	�f��$���� �,.�n��i�D�<� �LsE��L����_$~E�T�"O�(Bp�ߡ}��;uF�"x>��HT"O�,)����r�`[�f;7��@��"OS�%�7임 �ޯ*����"O�ڲ�!H�<٧ٕ(�� !�"O.�f�A`�
A��#�R��Pq"Ol�b��9:�c����SV��"OB���N�3�hX�!\�.F����"O�Yє�P�_r�Y:�[�i� �"O�EZeH�3~� U²�4@G��92"O�@��·W���B��A����"Op�ۢ͑(`�,U��ѓ\���"O4|�r��$?,�1׫�3d����"Od�I2j��c�RA�F�D���U�G"OT$��
k皔 @�PZ�0Y��"OLU��ɉ1�$�YBW.(`ڒ"O2�[G�܁`�H�(�s���e"Onњ���b�CF�ߠ��D�U"O�U�����ؚE�<1����"O�$3�ț����yb�5�mk@"O�P�ԯ�'���!�G��d4�@� "O2,���8�}k�� �"��"O�Rab�,C"���1�
��F"OX��Ī$:>D��d�=gPI��"O|l�w���Lu�����ˉqH��;�"O���M�:5�Z�{� Y8O�ܰR"O������>Yu����τ�s4d��"O��yc�A�[(1*M��f?��T"OԠ��9K����퐮z� "O�<��"]3\�j�P5LK.�IY�"ORLr�Z��Y��k�#1^`���"Oh���"3hȹ�)!p>zź "O,Mkp��.%�V��F9Ctp��"OJ�R� �v�����G�ok��3"Oƅ�.7DQ���Z=�0xg"O ����?10�V�J�L"�["O�t ���[�$���&חV���"O�TYюW2*h6YJL[��"O~���Ht����#*�=	�:��F��'w٪�ڍ�	�Kd�)c	;D��1�HٲJ!�d�=j�����˵ l*p��ԁ24@ѻ��I?��gl�|�'�$!Ă�V�`˅EA]3���'@tB�eV�X_��4�I:W���b2j�E\n5��刡LA����	�`���!�9yYDT�%�խZ���d�*r񺜀D� *Y��ۖ L�.�![��P�4���0�l��*���!��ېI$
���F��f�'�$�G��	<"ђG��3t4�F��)Pu��h�+��nO<�Ò��1�yBh�X�vq�F*��t��1�&�U�x��8�厗�n�t�CG���i6P����L>��n�Mc��i�%�v5D"�(<i��n�|P��B�p�9g���Sa���&��pҘ�`T·�q%���G1�������!,�!��Φ/�axR�ߦ<� �(�mX�z~$])��a� �`�T��h���� �̵!�Orh6Ι	\͜-JT眄wU¬�Ɲ�<C�N8澨9��H��!���s���xAAaKG�]0��IH�~x`݆ȓu�HCu@Ŋ-�b�&�Qq�A:7K�7R@�ಯ֟[k��(�G�f�'��.Gf���EW$B\F5y���KV��.Dn���*݌?�n1�`�S�6���X�����C� =(5QC	��<���(D�`��ƥC�u`tp�Bs�$�F�6*��kC#��w*��ʳ'��w�u�%�]�
�ڡ��-��\�Ɠi�0�#f�\��%���R4cS���'���cDMZ�m;D!�m^]dΜ ���L�`��� ������	4�!�$�T���x��`�
t��(q�dG�Q��!��0LƠXLC1�ĒO�`��iP�l(��u�$=�0
O4]�$"��v��9�J'�%��^�8
�c�N���0=� �PB0��=`��ls ��6��@���'���
�A9��T�sF-����4�Aa!�;{V\[�H�I�<��g��&�h�Rp�7
-$��M�ɃoR\v%[�}����$^m�Ojd�d攈c���6L:f�����'�(9�Ĩ	��`��Mv�6*ҒEJ�b������ � ���ē� ��슰(�@�"^sBh�Ɠ�*y��	��.u���ՐEi�y���R�yԒ0
щ��
�Z��䒠pL��/�I%z3v�zr�z�#�	�Y����<�g+R�X��<AR� ~HiR!��Z�<� 
:>��T ���,��g@J��@�c!�v��d�!(�B\8��^�y��.�>�I�)Cy�~5`��ѻ_y���ȓw�@��"{���×0*k\ ��_��c�"�$h�"��%l��<�ȓR5B�+�)n�+-"n�`�Q�"O��rA�I&��óLs˜u:&"O�ѡ��՗r�`Q豮[�w����"O����D�?C�Z�;6�]<��m�T"O(��q�Uk8�R%�
2����"O�)�'f��lF��&*B�*�,1�d"O2p� �(�X��P���w�1�P"O��%�47�`1C�,B
M
2,��"O�tt�2T����A��q�	
v"O �Y&k�<������&h�Q"O�)3a�)Q6`	aC/�zeb=��"O4%����302�{�,�#zEΉ�q"OdS�l�s$r)c녂G���kG"O�p�����*zpu�j�8st��[ "O�}Y7Q��R��d�Ot֥�W"O�̓���o0~e�`�!P�D���"Or�C�ʁ)M��l�� ��p�Cp"O�q1�
�z᎜c�H� dy�xr"O��8hB�о����/fb��"O�a��SC�F�pǫۏXfN<��"Oΰ��a�;%���bQD���� ��"O����C�h�:T+vĞ�[�z%�V"O��r�N�0��X�	Q�a��8�F"O,��r`�#k����ȗ~���f"O�u�VC�;pF���7a^}��"O 9���t�Q��V	)g�ċ�"O2|�2%�Z�8k�)��at����"O�EPT�D�MZ�И�'6P�{�"O*�s#�V�O�u��ѯd����"O�,Z�M�:\�,p�Z8iT^Lq "Oԉ�c�����r�.��N_Z4��"OvuZq� wƴ�'��%ʐF"O��!ਛ/n6\X��ſP �q�"O�]�Q �4	N�� �M�[���4"O|�
GEU�lf�8�ϳy |T"O���I�W���J�&ů\QFy
A"Oh���zҥ�g�[=*�b�"OP)CD�B�iu�\�a/y*�$��"O�cg���>���J�oT
P��"O���P�Φ0��уM�7
�4��"O JN҉�6�Q��D��.�"O^�8�V�Z( @8t��ag���g"Of�7`�*�`�)���W���4*O6����ܱv���
�V�s��1�'e���C�	���cϝ	�f�S�'E��1A`ʐy;Z��1fye����'�Lِ�cwJ��PPѱ$���z�'�81j��p��m G�A;���'��cƊ	#JR�0:'@";�$�H�'|~�DI*%R2��fG?�h4I	��� R�Jt*R�|.DT0&�,)c!y7"O�)�k��v=5��C�?ri�t��'<=��׿��	%I�.IC1�O	6xձ��� C�I=7 ��R_"�8M42[�O@�ib��jg�t��Ef*�0�g��p�y�o��g?�B䉺�Tͩ�)�?H<|9� iU�(}��Cq.U\~�a�+W�T�}&��W(��'���"�1g�h`��+����Ø+}N�H4�>H�Z��a&y�h����GE���K��Eʂ]$t�վ��b�&�w�@Ah"�Ō��]�J�q
g��V���o�J�E���W�<Av��8sD�!�w��*��d�Jgy����dL���"�>,�����	�;|:%q�Ƃ+H4�`�C�f�!�����[d���o=�с��D�I�t=apAڸD��p����{�Z��]>�<aa-��u��Y��)V�8;�Xh�KsX�H��D�5d(�y���G@�F!�g̍.k��s#,-X�`xxU�|��`��	� F���+�e���p�.֊YJ�<١%T�&J�ۥ�c���(T�����O��	�@�&�����6VX���'���w��9\���-�8ĩ(��x�ց[���1%vd�q�I��E��w�rd[G�hW����Z[(�B�'��lĄP��* ��/��u�h�BI��A �#I��R˟4���o�'�Fi��#Z@���j\�t_TX��n��Y
W%D�n�PE�+�!l����@a��q��i��d��%j��^�I���P����&�]�Ipu�fb�f���D�l3�v�c���8^�:܂��51�l�SSY�@�C�^�(�V�%\}�PC�I$	��`��b�K�耺t�F !<U�`om�"A�F&S{^a¢���.Y���4�sޅb0�U�Z�b����u�j�#'=D��hB�+�G�4���$LV�a[^�8ⴍ�t#�/�J�z�cF&G���0��J8 �Kt�X%�@����5���d�9,Wfܢ���6 H6��t���c��y��̒�{�Թ�L7nH��Cv��5Y�$!��I"c�(��F�Q��q�%W�DB㞰����'�-���j?L�j�L�)���0�O*��R�Y�8Ć��k�?T��yC�'�8�"4��mA�XId�<P�zlƩҪDL ��$�B��kE���a�0��~��x���T��sƞ��vg��F�D�b �,D���-̸v�]����(0��A%i�t���;'�i��\Ӳ��Q�����9r�Q���'�~<�
f�XC��b�7\O�	A�%r�����D�thVH� g�iؤ�8��^)d�,�AFĦy��-�K8���q�_�jQr!���U�Sjmke�#�	(����`�f��}�����dȨ�k�t�]�E����ȋ���@a�
�yҬǙZ��BF��Fw.`['*5p�t���.��`͸5P'��v�:M;���k���-�!��
$qiJ��nD�M�!��G�E-D��3�%Ji�A#A+E�3�v�S���<�@L����5�Z����D|�EA�JZ�#%AC�Q���rPEX���=	U͟/S�����AKx�Y�͔.J�x�t���WZ���	�N��	a@v@;��Qfѣ�I�+id�#<i�;.ƈ��F�Sy�O��Q��{�>4��f�!FX�];�'��!q҄٩dH"���Y'7�F��qO]&O��Z�Rz�)�矼
��%�����_�q��\��$D��+��<,��9GK�h�
ݛQ�"D�P!���s�v��@�eF�89�� D����&Ǽ_v@��n"tMR)� ?D�\#�FݏB,�u�p�q$}�cd?D���E��:�\-�fC�S���ڷI1D�xB�ٰJ�=�[��40��L�!�$�PMz�Q�Lϔg�MjA����!�dJ�Oc�)(e�ǝ	�����x�!�dӪ}G
8�D�=*Y>ݐ���*De!򄏛[ǆ�p����x@���&�#?a!�$2�	����7DT��(�84U!򄜫YP�@! 6�������:G!�ĝ3��Q�m��<����-�I!�$<vpƱ�5J�7)R}�흽P�!�YGB�뵁9?�@�\%�!�H�Bx�A��� f���oB��!�^X�u
�@�N�>՛�?V�!�� H�8#�Ϩ.�������H��"O<�YS���@6`�2��<���"OHU�A��_`��,*	�}S!"O��#L*RL����!��n���[u"O�YA.��U���ˁ,전�"Ovyc��ppSS�I49��"O�x�/�t:�h��%/�Y��"O�AbU��eD��
Ts��,e"O�)�V��/)�(b�j�3��J'"O�aCP�2�2H1		��!S"O��0�ǻ�P(r�h3�a�R"O�3 (D�/,
9�ѧ�M��@JB"Ore���L�D0 -8�������"O0DR�����|�*�G��w����"O�����$��xYW&A�T����"O&)�e��x���%�����"O���ូ�Q�O��g�d�q"O�<�P.�DX��J!a����"O4��B��}*8y-ȈD�����"O��FYp���B�M�)
@}Y�"O�i3��$+,PP�6&�p�\}��"O�u�b�ށBl��)��J�
��!�"Oz(c�_�}P�Z�gU�_StJ�"OĘ8@��T$��D��@���*W"O>�s�cI�1R��PD�rQ�X�"O��P*8&�,��Gʞ		@�qA4"O����ZTX��2G*���"O�T8ң��/�QF���]�D"O�,)��		~Z�$SV�F��rA��"Oĉ�J��^��c��X�A�p�&"OR��R�!Z���Ыk� �I�"O��"�ŽT�^�:dM�/r�6(ʒ"O�	bu�R��J�.N_UR�h5"O���Vc#����l��s312"O\m#�L�6m|<(ؔs#f r��>D���,�w�	j�&Gu� ��"�:D�X �/���Ƭ8��?
y��ɶ�?D�8� ��#~[1�2>K���(D�䛃�[�^(��y�R�F�����) D�9d*��/,���BM/~HD��s�;D� �a�Z�H��5���)L�f�2�9D�xa`��b��[@\5B|<i��:D��ۖ�nz�8	d�� i.H؋b?D��I�eĜi� [��W!FdLB�N/D��b�ؽL�V��'l�lE*D����.F��Za!�d��F�z��&D�hI� I�6�J�k�*L�
�����$D�x�����T���3rf̂,D��3EߏN����K�B���� D�$�A��2-��zW���8��<D�xs1 鶴�5&ݝD�
����6D�4ĂT�-�-�]��0��8B�	�z��L�k:@�J e۶)FB�I���p�W�eB� x�W�$:B�s��$q&���8�p@��9SB�	�H�vE�C �Q`�����Q&C�I�� I�bذ�d�b`f��C�	1ne�zs�é�����`�=�B�I�q�D�1l�96eHAk��A�O܀C䉩��L3S͜L�N5�C��m�~C��f��LD��~���&�6QMjC�zZT
�3M%���o��bgvC䉟s��3�-^3k�U�@�	/~W�C�/?L�H�c:&�X�с�8�<C�)� ���T´C�uC�m̊��l�C"Op��3�;v�;Cl�{��љ�"O��Bu�ҏ_o� �,�p���S�"O�]��MތH/tS�!n�x"O�����,
�Y;7l�a/�ę1"O��hW��(F��Cu���[!"O\���C.v�I�'*<���"O��#�P����"�$6.�2�"OI'$D�z�x�x5!D�h����"O8k�@<DZ�$����<k�"Oz�J��;|C��r��{G�!"O~)	��F9k��|���SJՋ�"O<)��G���6a����aZJ	Y�"O��B2�;1�A�a��"���
�"O��{`@�)�\��/iwԜ��"OVؚ�+�b# %P� ���2"O :D�4K�tض���9kBi��"O��jo�������4m\2�ڇ"O,ܰ`Ʌ��89�����9ؔ�"O!���?^�ҁr�(�Z��<3"O`@�C��6}�l��B"5���@"OF���2 ���K"�A�!���j�"O��ѱ*�+g(8��oB��� �P"O�}��͈���bcy�"O�0ʷ�3�:�b,	#(_\�HA"O@-y!O	a�)4="D�[�"O4X���}�RHt��'�]ʢ"O������Lɘ��ۋ�I��"O��Y�A�|�*�8D�� #��Mb�"O�\:U��+��m��'�(�� 4"O�]����`�ҥt�ɉ�X��4"O^�Kd`�,��m!0e�F�V���"O��"񥆉|��,P��FPt�xA"O��' �:�Zm��E%29���"O��A!IQ�����4]-r90"O��V��'�\����w0�{"OVɋb�-���c*�j�$*�"Oh9�Ř>*�����
�z�����"O�ZÐS����rE~�\��"OL�y��Q
��ue ]�`�D"O��4͵EO��aD
 0��k�"O&�$R1=t.��֗S5��� "O$Y�a��6xA���1<�
�"O�E9���$(�9�nO$_>.<h�"O��8g���M����a*ļGJ���"O�E���Lrb�8��U;D� Y��"O�x6�ҜX��a㗢��� �2O2���ٵy&$��1���$�1 ��ɫ*ϒ����,@�X�$�V�f0B�I�.�BMjs�_&?�����('3ZB�o�n�x��=*}�����L�h�C�	��� o\��Z-)��Ȗ����(?q��U�~}�5��M��`�<1ԌˊX��-q��UQ�H�1U�
w�<�a�¢��@` "�k���S&)�l�<�*j.g�=�.Ԫ��_e�<ɶ疼KpxH2'UM�ܐ��J\�<�rُNHcƝ=S$pZ�bRX�<�g,֢?%v���G WE�	��nJj�<���7h�� ��DP��	d��b�<rDث��E�2�r�,^j���E{�G(�����"	�2��x����u��<q�����'v���yU�C�2LP<����&WQ��9�V�4I��ا(��$A�أx�}z��Z��76O�9�'
1��?y�>0nԐK: ���E��E�f^��D	�����?� ���Ԉ;?.�Ivcէm���Z���H�'
v��i�'`��p�A�&��Ua�.��Oڹ��i>��\�`y��S�/ت�����!pz��%�P{7��o�S�.PX�g�ݺ>��S���'�%�'���a���ӟcԘ����! �x|S`�ٿZ�>����(O?1�WDϺd�	�	��ł�"ac�<��?3mZ��kMe�2]
4*^�<Ys�  ���'eV
K��,jEq�<�%[�M̆���d��#u�� ��v�<Q�O q���A(��(�6��G�u�<��d��*��=�t�zA�^p�<U�K�N�0��q�5JӁ�v�<���%(�p�ڇ�w�p�³#�r�<A�čA�Mh/	s$��+��s�<�0�\�P�2��@�߂��!BIW�<�� Й-�0�c��,+5�CQ�<�AI b��e�,j�x��&h�<�r�S��Hf
�*�T�#ĬNb�<�p�O��t���n�"t�ƽ����C�<!4�TPj�!]:�����=T��J�M׊GP�[��(1`��,D�$��h�4���CF�0_?��;�+D����n�?U��P�a��t)�	��(D�v�i�ê���j,�+^Rܘ��'c�0�����8�ʹ匊+j��x��'�\	/Cd'���Tˉ8_(rt��'[D��@�1~t��3����2��'��Ĳ7�ù^�003��%Py�i��'z`a�� ����oV�xXҁ"O�Q��R��m2���e{�"O~���
Ւg|��f�OV�8m��"O��{�jP%H���S�|x�0`b"O��"��t[r:�o#O�\"OT��c�޼G�D����G��};"O<� "Q�Ԁb�G�K��9��"OF,KՇU>�\tq��2\{�"O�Dį��@�y�i�6)�NܢT"O�3�Z�i�D�V��D�aW"Oz��S�L� �q�����p<�"O*Ⱥg�?}�x�Zu%VT�\y�"Ox�Z �I3"\���� ,:̪w"O�$U*.�:�c�@�#m���@Ot�<���4\ܦ�S��R �e �iF�<�0�<QLxPc��X���t�C�<i���q4�rD�O�S$BY��|�<���W|�qhEF�	(�\��NJp�<��-�8vA\�����f3�4��YV�<IuaN��{&b�*�n!s��\h�<���:H
fLЙ�4���Ίm�<��@'NO�E�D
H<�!�:�	���S?�b��v�C�!�d�;�Ԑ˄HG�a�Tat(��=�!�d�)U:,hF���p����>�!���f�p}�$+̀{�d�<D�!��;�p��C�� n��i�cܓn!�1y�J�" ��J�����4x!���+�ΐˑiBS����T�'
!�B�=^�yжK��+�>i	��I�X!���(}���#T�2]*6�1a͌!�σ.2 ��ߒy���cj<'!���x5f�s�)^�+׊ZD�C�{�!�$�|O
͡P#�M�E���	>�!���
�3qO��e���1%�ՐF�!�� �,��l�0���!"�M�!�� �4�se˥H�N�s�)��aQ*��"O�ɘg�ωS��E�O�{1Δ�@"O<4BfIE!g��0���DЀ#�"ObT8��Mӄ�x��>�@��"O~��@��Jy����(��+�"O�ܱP�GC�0��0[ɪ1�"O.��"i�&E��ð�>�.�k�"O@з��&/6��j��LĲ�"OX�C�jB
8��i�>��9;@"O�ҥ�%HcV�۰g��i�DQ "O��`Q��6Yd��(��[�B�Q�"O�lySǅ\��j����\���p7"O&��`�M:����83��ɉr"O¬�0�)[�X��W �F"F1��"O̙��A�"_ܲ��ɪ��/E�yrN)
Ll�����	�~�� ��yG�L<b��d�BVI�`������y�
ڀe�$Qum+c�<ēE%Ԍ�y�X"�YG�C-^Ȇ�B%O*�y«��l���b%l�;f���8 +@�ybM�2<�LAbq�-
^�,��
�y�i�d���r�9|�´3G`�?�yr�7|���8�h�KB�K:�4�ȓ_nq�1�ѷ	N$萦�+O���ȓh0�"�����['Z�9[�̈́�~s��b��!�r,a$EB�2�:Ʉ�,,x2V
����i����%�0نȓ �%8�mX*���V�R�5����!!g	7~u�����ޒ
��-��{��T�&̂��ʔ�We�)-�l���$�.y�p�֨Czm�f)�r�L��t�RI !��+;�4�F��ni�݆�7V�m�"��Q�F��e�%���|g�� 瞹+�A�SI��j �i�ȓ?�*	A%r�lx�Ğ�_v�����s�K�����E���i�`���-��1 !��R��72)h͇ȓP�Ј��ŕpf�u�i�	hE���(yy�B��WQ�|�'���8�ȓj�"�Y��XZ�P�(�*n깄�~�*����	�y���TBD<XSd�ȓ*q^��m��h!<0�&��k���ȓ���1���{��)��ί>M(X�ȓf��" Z�h�b�[�wX���G����׋E�7���$Ҽ~�怇ȓx\t�h`-��7P$�s6"\"h��@�.��b��	=�|�U&�5��}�ȓ7b� �I��T}��	WKP�r�J�����QCːx8�6�3A��9��b�� ϞY�at���捅ȓyŎX�s�R�q�X�x��A�5����^�bd�d�@ ��bBi��<�F���elv��S,�gꌨ*��� �Ą�a7�$
���T�,l�րB�4���qr|˂̀[w��!����y�ȓ	>ژ:�I�es���.�(Y���ȓ_nD���M�8�%�P�ը�2�����cGGD�J�, �Rl�ka*M�ȓNX�z��߁	_$��jӔR�\���0���g�TE�4��c%��sC��ȓ_=4�RDwfe��KW+E���ȓVs�T[��?/����R/T��0��G�r�J�
aĐe��@�7rp��;��Y!	�01�A���S4de��S�? ���O�>+�TMc��	3LY"O~��#cP�Qy�tP�h�
N4Y2�"OJY���N� ��8�i@�dhm�"O�e#�AYN	��&ޮh슑�#"O0�a�k4m�~�c(ҳ
s�}��"O,2��D1,a3L�:;�Q� "O�u�L�� D��e�"Qƭ��"Oޭ[��/�>�D��RW
̊A"OX| f��&q�8r�M|<\�P�"Ol%�r�-%�uʢ�!4-"�z"O��pʍ1m��M�D�A � C"Oބ�IJ�,a��Cm޲|z��"O>�+�(Ē_d���'LJFRF49g"O�8�FJ�{A���*�<1�=�u*O<e�#���KO�M���f���
�'=�Q��#�o���D�r�ؕK�'*|H���M�5vјU!�>�&P��'��%� �!z$t�����G��k�'��G��%�����a��P_�eq�'�����	Ю6u�� ���I�H�0�'���Bl�=���1� ҕx^��z�'njQ�#�!=�TE�F(H�;�xd�	�'�0�ڲ R�,\�+#��?3���A�'��[�l�;ޔt钣%1�XZ�'}d=q�OT(+l.������(Bd���'H60���̅
�;�!V7%:&���'�jh�C���&<0Hpd��(��k�'&F�;�Ζ�5������$���#�'8
0��j�c�m��5p����'�,	#���d
d}8��ye�a��'�ӄA �"G>���mϚ{��IB�' �����C��V8��d	@�G[@�<�&�t����7P��A��x�<�b������(�i��8��ae/F~�<a�fG�`Ɇʧ��
7�N��ZA�<ԅ:S�6}��A�npj���g�s�<A�o1p�u�0
8�l$au�Pl�<��N1Rm켁`!�%V�p��	B�<Yq�D�06U�a)N�q�v�#*ST�<�E
�
A�]hP�L+"pP���P�<��ŋW���	��I�x���+�g�q�<7b�'Z���he H��b��Øm�<9ԅ��K�\T�F�ucd�`��!�yI.~�8�I�G_
���
��y"�,7Cz���^?B� tH�hܒ�y��7C�\����F�"ȑ�V��y�%SA.���J2Bi� � �D��y��b�)��CR�:����ǆ2�y��D+v�^���AL;�ptYrb��y���	�@ب��S�d��ac�B�y"	��j�Bd�T�^�`J�J񫑈�yRf�.j�1F�G�j2 ��֪�y"Ɏ�=�e���K%��M�u���y�fD=���S�H*O˒���I��y��$����hKS��� �0�y���[����$Ets�ّ����yR/�=��Ҥ�O.W2�4�_��yRf�D�n}��K�op �	��y�j�)5�n��FJa8��K�AR��y�Ȁ/I<�0eŔ�{�`��P�y����f1� ��M�k�hI��ˋ�y�oA'!>������dq��T�
��yR��zGJ�B��n��1����yb�?%�R �7.������y
� ���ЂE�'�X�+�.;��2"O0z'�T�[��U�K���6�"�"O�dxV��	�^A��*ɡe��I�"O�A�VgV�m��u��	�$DB$� "O�=��E�#���
--�\ �T"O���biQ4j��-�t� V�z�1�"Oaa�bU*�RP;6�� ��٦"O��X��ǆe=@
�k�=� P��"O�I��6l� A�0�
, �JQ�"O
a�� �Z����g�'g� AI�"OĀ�f:M�T-3�
�[�\�"O�����Ǫ?��^�D���4"O��x�
   ��   �  C  �  �  t*  6  �A  5M  �X  ec  �n  �y  ��  �  ߙ  s�  Ũ  j�  ��  ��  H�  ��  ��  D�  ��  �  d�  ��  '�  ��  - s � /  �" �) E4 �< C �K xT ([ la �g �k  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+a��6 \��	�<4�d5h��'�B�'���'	�'/�'�B�'��I2w��5Kk����e��U�D܃��'�b�'A��'���'}��'��'�>��5�\ h4tIR �>���'l��'��'���'2�'���'b�Iz�k�fVЂG�[�x.(���'���'/2�'��'"�'"�'�^�qs�S%V��c߁Lb>ıf�'��'@r�'���' ��'h��'J����b���@�3MTV<q�'�B�'�'���'���'^��'��`�$�͡9Ql�#[�=�"���?i��?����?!��?9���?A���?P�Σ9<�x�
�&�+K[�Jъ���O<���O��D�O����O���O��DLw�eȴ���ŢW�2(�'��O0��O���O"���O�d�O&���O,���ƏX���K�8�n͊���OP�$�O��D�O����O����Oz���OL,���0�"&�:3�f�j���O����OD���O����O����Or���Oؕ����JT�
�G�Oݨ��Ԣ�OT��OF�$�O���O����O����OH�0t�ʰ[O�XbQd|�^4�G��OP�d�O@�D�O����O���Lئ��iީ�ć/TF�U�ՁN�:�Z�34�ڂ����O��S�g~�i�"���]�j߈��'�M�Z֢��-�&����@�?i+OR�T������I�h$�c����9����O���CAp������f�Z�Oz��1!�+:� #D�5(�����y2�'��D�O�@誐b_�w��u#�$�Z�b�HbӢdS��:�����-%�d2���v����
��;���I���ϓ���)_�+�7�k�t�f��4�<�x�iF�}v�YEw�x�G�r��u�����'�|9�`�ۄ5p�2�fP�J{Tq��'��	[�ɯ�Mˣ��A̓^�n�f&\5�@@��${n�9��S�D�	��t����O�"Ip��1]j�*�iل��I؟��E�P�	40b>��U�'50P�	�Z5<����� �<����M$Q$Ė'��	П"~�3�(e���Ζ,S=P��!GR�<�G�i�8���O���?�i>�8��D.=���s C�d�~���a�����I9)	��n�k~�6����S�)�H��Ě	o&��f7V|hM���|�V�����l�Iן �Iǟ��G�[�u�h@j0��X
P2�
Ey��g�Xy�@��<Y���O&�wцf(0�` �C,�u�W]��{�4;�>�4�J�i柒%�D�^-1�}@D�U�O��a�թN�n���@�+�OL�t����Vnl���N<�tT��ҵ��5�>i$���3�^]`F� �	Ɵ��ӟ�Wy�j���Z1��OZYh�D�4E`U���6��%Ka5O���0��Oyboh��8oګ�M����y1��r��W.r�$ڸ,��`3۴�y2��, ���}�J`���'F��/H�p��n�Pn�L9��ރ(�����(P��y��'�b�'�R�'Wr��Tn�f4@nR�C��h����<N���O>�ڦU
��Giy��'.�'c���"F%K�Qx��]�f�p�(��}�\�m��?9S��ܦ��?	3$^&��a"J�:�4!^�}�p���+�OP��+O��oVy�O��'a� ��J��wAZ:ݖu����x\��'B�Ʉ�McV*%�?���?	*����7-�_
�U,��} ����<�' \7�Kܦ��I<�O~��VhC>��y�OWi����獤m�d\
�*���d�ۺ#4C�O��/O��)b�0�� �K?;(P�HEl�<8����O��$�O6��<9`�iV�츑�j��,���Sc�	Ide��I����?9)O,hnZ�E/\�rs掕�ZL�f��?$��R�4Km�ǎ���F>O��V�w�� �'^m������F>ێ13iʌv��L�ٴ���O�D�Oz���O��D�|b�[�+�&@�Ҡ[0	^B�)���"��`
�([2�'�����'/�w��H��θZ/�a���N�,�t	��'҂=��iE�6a��0�nҙH>�⦖�D�و�n����&��uxӜp�)O�DnTy�O�cԚ6�,��Fe�1T�<c�
�Yf"�'b�'��:�Mk�Q*��D�Ozp�l��]�@Y2�z�6���&�Ity��'��g,��@�|�ѡ�EH�8:,Q�`cO�m<��O��C��N^�ՊV���!^w�^a�ɶZMW. �1�T��eo�M�@܎K���'�r�'7�X>i��&��u��ʱ �>����%-^�
?�̠��29�V+�
^������?ͻx`u��A�:Fj���G
�$?H���M�r�i.�6�;J*|7�r���I<Ht��O�:�2�l��3�虧��)pZ"l)��iy�G~�J��|���?���?���R��:��� Q�,���(h��}�+O�%n(DI�'kB�iΠ;������7ަxіi
#@r�;�6�kӢ,$����?-��,��3SG�J�h�.�U��^
Θ�3���fĝ9Rg�^y�z���mf�:���^1N��䩏�=��)���?Y���?a��|�,O���RL���*7bH��d�-�� ��mN�yN���O����'´i,6���EMP)�/�[?LQpM�u�9Op�$�)"�8���')����u����  d�'*���p���>J���7O��$�O�D�O4���O��?�:�h��eG�0��k~����FM런�	ɟ� ߴ�j�ͧ�?9���aB���!D*m�y�ğ�p�
�!N>y�i��7��Otxq�@y���ɵv��b�ȞB#����AKG��<{�;}*���"K<�M�K<�BW���	����̟X ��4f�&�8�G�X���HßP�INy�a�j�#��Ox�$�O�ʧZ��ە��h��ɳ��	
�a�'�����o�)�CV�8a���%AK 9>����� ?�u⣫��� ���f��hA4�|"�%G��QAM�S����!�,R*��'�"�'���[���4iyR|� �A�#�������Ƭ RwJ����d�Oj��'�B�@�,nQ��#f_��;���-?,�'0f���i��O �""����w��HZ��Z������&���c���'M��'��'���'����-�V�ނY\8�{�̛�y�` ش!sJ�{���?i����'�?a�ӼcB�Q�!�.��G�ɠ(�8Ӵ��&F��'�ɧZ���:Ҁ��MӜ'�B��V�1,�"�G�a�� ��'.lea��PF�|RQ���I��l[��L$:M���`H�9w�|�Jv���Y$k������gy��h�]�ea�}y��'5`x냈�<=�BҤ�^S\�B�$�<A�i����?�d�#��5@�e�@�`�Wu���O*`2���g�T��o�<��'D/���?�?9Q)N�p�9tI�:��i:��$�?i��?1��?���	�O^�"+	R�i���)3d�9���O�yn�g��H�I쟔�Ir�Ӽ�1�T
M����i���!X�K�<�2�i�6��w�F��fOs�@��� �Q+�T�4�(H�jX����i=��C�,����$�O���O �$�O��K�K(R�i"ܦXj���QKO�^���\��v(TZ~��'�����{.v3�k�.Zb �k�!�˓�?����|���?�dI�A~:��.��R�d���*_��3�46��	�=�PѢG�O~�Ob����9�*�Y� ��0nDA@XD���?	��?���|2.ODonp�`�I����hD��&S�}Y�c�b9�I����?�)O>���O�n@>�6Y����"�f]�#�W	i��L�f�g�����*�+|<�	�<	�����GŢ|�ԙ�E�3g��(�v���<����?��?����?����A$l'��k!a�p���Ȋ9!�ǟ���4W�Z�O�b�|��P� Of	vB�x�����$&l�'32�'q��b���7O��D͡T� �@I���4k"�Ϳ��A�DI0�?) �*��<�'�?����?�'F�"M�"p@�͝37�%���F'�?i���������I���	ş@���?�e� > q�Qt��(��+3?Q,O~�d�O��O�I�OF�HF��0�t�IR�C+,D����Ld���5��!����?a���'IXy$���勆Z��K����%��"�N�ߟt�	������b>�'>6ˎЙd�H���I�k�HX����O����O���'D(7�	��"L+@Æ%��-Q��]"Mv�Xm��M�T.$�M��'-R!Z#/��S�L����Be!�-H�Q"DhǍíY���IWy�'��'Db�'	_>��B������G)�i	��y5H�M#c���?���?)K~����?ͻfD�	��Gz�\��ɀ�>K�jQ�iaV��"�4�������0���C`3O��h�C�-k�2���[�*��-��:O���� �?�
6��<���?�W���5�L��cㅓ_U؅���W��?���?9����d�����hyB�'��4����]n����fHu�j�bg�Ĩ<yQ�i.��$(�䉽L��y����!�2�3e��7LT�ɘ��J�!o��$?ib2�'��9��:&��<���O(E���+��ם�D�������ퟬ��h�O�b+��K7�)���K$^o�`1ȚJ�rF�Oi��V����[�Ӽ�7j� G�PEK-L�Z�B���<q��?��|�T8�ڴ�y��'�Z�Ф��?��)v�ؖ�G�X;^���x	 N>�)O��O���O��$�O¤J6�� q�9{E
�<U�=�'�<�ĿiT��#G�'.B�'��O/�&�:v�b4I��,O
�'��,!��	��M{t�i�|O�)���I�([��*DB�& ��1M��e�=��(�G���MP�5c��'�Z&�$�'����vd�� ����t��4;�\h��'Zr�'�����$W��c�4��x���Āk���>��p:�#�b��B��?��������Ϧ�����Ms��M�S���W!�8l&H�ѫ^o�2S�4�y�'(z��s���?��[������I21��uh҅Ȳn60���qJh���IƟ\�	��Iß(��䦉�I?��B)k��B�MC��?����?)4�it�(b�O���'��'x�zB�R�Yk��O]2GɚL���7�$}Ӡ9m��?�u�\�̓�?��k�m�HJU�"y�abTf�aX`|:VN�O��hH>.O�d�O����Ov��3��/5�vq 4g�4]X�! �O��Ĳ<a4�i�6��t�'��'��5w[����IC5�L���X(����d�O���+��O���,' ��1����q���!
��P bȔ�x(\Rc_�L��Qy�I�o�	23� ]ѓD�5P
��H�o�;���	ß��	ҟ��)��Ey�j��8������̹�Ν�1��4�eA�/�~���O^��(�Iyy"Hn�H`��#�8�Zɻ�m�M�M*vRƦ�4&hl)�ݴ�yB�'���{D+�?ER�O� �%2�J�[|�+�M �O*B� �4O�ʓ�?1��?q��?!����IT�5���*c�F�8|�w�)/?�MmZ)�`���ǟp�	j�Sǟt�i��跀r�V� ��]G|����J=�M�W�i�<O���Z���=Þ6�{���J�7l"�@��$,Vb]P&�{� xs/�5��%�E�Jy�O=�D	����Hd!3X7����фR��'��'`�I��M#��P��?��?E
��P�q�\%+=�3�S���'�������T�	�O��}��hʼ)�u�������	�|+��a.�Y갈/?����V�$��?�'\m��X���"��PN���?Q��?���?1��I�Ol�K1�I� :n]�g�\1& (�����O"<lڅ%����ş��IE�Ӽ#��	�EI$�:y�P���<����?�'��<�ش�����y�@�?�ñ
ֿ����٪&�L��Dh�i�kyr�'���'�b�'��{x���G�8�� VM�	���(�M#�gM��?����?�O~��Mz[%B�kL����.N.ب�.O,���O>�O���O
����k� ��A�b���c �~Yڰ�v�Z!�'��YV�RF?	N>�-Ob,�#��N�4��w(եS��5���OJ���O*�d�O�<iV�i� �W�'�ܨ3�D��.p�sO�,ln�+r�'r���<���?�;Q��Q�i
< ��e '��Q�<Ȑ�fU:�M˛'+�+����'�����B��.f:�@"E�@��x��߷`>��O"��O����O��d.�S�`��P�A���]�"�-Ay��Iڟ��ɲ�Mc����|Z���?yN>!HҢYӺ\b���.Q��0b)�7��'ݦ6������+��-��?)!(�"Xdܝg��y��V�	��a�O��qN>�(O�	�O��D�O��j�B��n͹4�ű
�1���O
�$�<ɢ�i�"�Ba�'�r�'�17YxAb���>�P��M�z������y�4L�i�C$���(������,<-&�4������4��e��%��Ob��G�]88���+D�X:�l�T��O�d�O
�D�O1�fʓ4��&��=��0
��q@X"c��r���1Q���	M����D�O�� 3�ŀ3B��#���>[Af��v��O<�D�/w��6y�<�Ɋ7���O���\����"ϭA0��Ec2�� ����O����O,���OL��|z�cQ"c� @���S_2}�6� �[�fɖ(�R�'����'�w���)�K^4{a�d�clz�����?������|R���?q��X��M�'����6D�=E�pɊ���S����'Ad�R�+�ퟔ0��|�[�����u�p�L�P�о�F�[�Bǟ �����ry�az�4�YD��O��$�O�q"��a��3n�S}h�`/;��y��'lr�|RZ�9y��tGXsw��(Qm��y�'i�17�� /o&���O���=�?!e��O~e�g��w��D�O�q[�ѳ�	�O��D�O����O�}���c�"0�p��u���Ea����b�&�&��B���'��4��Ъ�O�s�^q�f��{.2˅9O�1lڑ�M�b�i_�iG�ii���O&�`�P1����<��R����.��������`�>�O���|����?���?�?Xҹkq	ҙy�K�D!{u��)OVAoZ6k��I̟���}��̟�𓢁�TP�J�M�&c��U*a��zy�ia�toZ����|r�'���.Z-�2���%Zʀ[�@V.ic��3�j�}~�A�\����I{B�'��	�'rt3�Ͷbl�G�S+/��	�	�,�I֟��i>��'�7�ܸ\�N��a����<3�ђ��A���*���O(�0��W~��'��V�dӢ���̺!Vh��̎�qt*����]���7u���	Q��!!��OB����&�MH���+*LD���g��9��?���?!��?���O�fu*���7�5�v�C[���5�'���'Z6-�8�˓�?yH>�6��%(M\����1iY&��f�n��'2�6M�۟�I����7�)?�6���#� �z�g�f da�n�)Q������O��#L>�*O
���O����OAS@��_6�S��͓|��ԃaa�O
���<�q�i��h��'3b�'m�S�F��G	�R�����/Q�F���$Ϧ5�����S�$�P%�9IF*�%uZ6�)$�Q�u�%ڕ_�d#Q���jXbi�V�	���zQ��>C�����M��M������I˟��)�[yB%e�v,Sa��9>�����Yd^��]W&���O���4��ky�lӖUq$��#�Dpi��@����3�M��M�i��YCs�i��d�O��{�mG��A�<!��N�
g(��V���H[�a)�E��<�(O �$�O��d�O����O��'&�12�L�AC�<Ab�L�}(@�B�i> d+�'Mr�'��y�y$V�M��53��Wt��}�+ʳ'�2�'�ɧ���'��G}q�f<O���^���1�N�n�X���]�y�
s;���	�o��'>�i>��I�x>\��ҋ�K������4xH�,�	������'��6-^e����O���Q?!d� ϛe�*ԡu�P-\�4�'���'�'S��[��� >�M������1�'5�LXP�xl�io6ʓ���#��H��%B�8|+��'ʱ  mTc�������I�����n��ywg�Z�� �2���l��h�'(~B�lӦp���<������yK֩��xrl�.]��0۵Bҕ�y��'2�'��#�i���?��EbRU� �����X�sG'e}~���#!���<A���?���?����?��(%Ԧ����%x@�������Φ��'ߟL��П�B�ჩw��ܺ�%L#6�P�N����O�4�4���D�O2xz'iP-��%`!NJ�(2ɛr)H�6m�ay�I^��JI������v洜���� �E9c��

��$�O
���O��4��ʓCc���̖\b��	7�`���ӣv��8R�E����'��O�˓h�V�e�^�n�62�&0ҡo׵jx�XK��L/,�RwFҦ��'�T܊7���?��}��;h8���ESJ�
��ȭy�� ��?���?Q���?Y����O���b�Yp!b��
�?~�,}�w�'���'�d7m��(��	�O���>���12Px����'�&��o�@�8$��8ܴqR�&�O=��2�i�d�O0��Z�J��0Z�!��D�k^/&͐���pp�O���|
���?���@���w
S�q��CVbR� ����?�/O2�l�ɂL�������O6�`8��8pA�%�& �� x�O�)]�f�O~O�I�&YB4�X�,m�c䁺�J�c.�% �\a0p-ʦ=ώʓ���!�O�<sH>�p�A�j���S3 �1���	�?���?���?�|Z(O�m�7$T&1���&q��(�)�:\�$\*GLҟd�	��?Q(O�o�+���m��.�L�U��-�|��4P��v���$ۛf0O��P�+k���'U��˓��uy���Y�`m�u�]7�-̓����O��D�O����O�$�|rDB�8$�Q��BݙP�6U(��[<k��/Ä
sR�'n���t�'��w���秞;0�y����,�&8R}Ӽ���v�i>����?ݠ�b�ڦ9ϓ)F��е�T�OHM�ҥܧ6�|��_�Z4�`�O�}"I>1,OJ���O��:!�ԢteX���`ۜH�|�����O�$�O���<ٖ�i��x��'aB�'�X�SuXPy�P1%?=�hq���<����?�O>�ƣ�B��Y�a�Z��t���<i��~z�i����M;WY����)U>���O4���䍝<!ԍJ�H(�­�A��Of���O2���O��}������[v햃"��q��D5Xs(YA��J��k�3�"�'�2�4�rmz��x��#W�,��;O����O<��\��6`�0��+,���O�	R'��{���@Eܸ~�����|U��������IP�	��ęC��~.� K�N�m4����m�Ly�ioӦA3��Ob�$�O��?9Y���)u��7,�x��թ��ay��'�b�|�O_�'�4�P��9�	�f�U%p���΀�c���)�<񠶜�;��Op�O���l|�DaO0z~Xݱ���6h�\����?1��?��|
-Ot!m��(eB8�ɿO��(����✣$.u��	�P�?1(O��O����W��(����DH���M]�$
@��h�J�Iٟ��!��:���%?��'ҿ3%�����2�͐����S�<!���?���?����?Y���M҈�`�ޭ�FHG�P-d�"�'�r(b��`�l�<a����7x�գ�HH2������a���ZK>���?I��g��P�4�y2�'m���K -��X�*��4��^3�:�T�'"�&�����d�'QR�'�
��¡\�LƎ9R�lQ�\����q�'%]��.&<>mq���O����O��'#t�� 'ôE�0�2����a ?	*O����OȓO�ӿ<�z�)I��cu�0yњm��������8��>?�'j��ν����L3#Θ�����h�������?����?��S�'�����z�A3CE-�Ɛ�k��hA�[;IT8�'b�ĸ<i���,p�v��?#�J0�7(��b����?��mҬ�M+�O����OJ=�L?uq��>~�RP�d��D�"�p���':��'I"�'��'P�ӻbb�0��Ʌ2��%S�&�9V��ݺߴO��8���?Q�����<a�Ӽ[4�E�T��D��mQ�i�O��?I�����|2��?AQ��M˚'',L�SƊwx���#0�~ �'g�8� ��؟��|2V��ğ�b���:6⅒�K��>����g�����������	ny��h�&8�7�Or��Oي-A�R8�%L6@�`����O�O�T;���q��l'�@:5ゅR�b���Z8��dx"c����q�=����'+ ���&��OB@��%}�DҐN�6K"T�Z���xc@�����?��?)���h�����i�0��Ґd��U�.S̘�������wP��l�I��?ͻM��h0���w�dezXH@+�Ň�<1��i/�7�ڦ��DCҦM�'� �ƣK�?�� L(3'��X��R'����'�i>U����|�	ٟd���Y��+���"82M�th�L�'��6m�d�����O�����$ʧ�?Q��O�u�ؙ1��B�x�V�k�Y+��d�O&7�P��p����`�{f�@\�x3��*Akq��,��j�HXQT���\�l@$�'��u%�`�'4�a2c�� �J�(� �&�n�h��'I"�'�����U�,�ش
�0���?y��R�$]�r�0+Ĉ<M�]���?��U���ݴlO�Vgo� `�E.C�1	N��p�H�a#���E �!��7p���ɉ~ʸd���Oi���;2J>=����G��6��9��̓�?���?q��?a���OG���΄	8�~�񀍛n��\X@�'�R�'Q�6-k��|:��?�J>�سOJ����]θS"��C�'[�7MIȦ�S*�8nZ~~b ��� Ν���U+N�+�?�ޑ�V�9�?P�$�Ŀ<ͧ�?����?q 5Pkf���o�5�pt�A���?����?�HٔER��A5�?i-���oz>���XJ���a��^;Je��i$?a-O�Xo�6�MR�x�O��Ď��:d�(2��
�z�c�IG��E��	bi��X�O���и�?Y�h:���;�L9���z�:a�*��u����O&��OP��)�<i��i T��U�W�P�l���V�@Ddx3��P.Xa�	۟�?1-O�n�	'�xD���A�\9���/6�
Yiڴz���\�K�V>O����K̲��'cl�˓AUrEZG��&9�-�"��U�t�͓��D�Op�d�O��D�O��d�|
� ��R�����.P��-�l:�VA���B�'(B��d�'��w���E�'eVL�El����hc�&p�(y�	I�i>����?u"�Φ��=}�e��^M4Q��a�.e�0�S& ���OH�
J>!-O��$�O �kB�E�
vؽ�r��qF"H
��Ox�d�Ox��<!s�i���'U��'�JeA�퀮:�tq٣�z�y����<�G�i�r��9�A�S��d�ER
>�am�.e�d�Ol� � >�����<���5�']�%�ɝk��x��a!��E�Q� V���	��������IZ��y�g�/�H�=X� a١@ضv"�r�plC��O���O���]�[_��pC�� �Jqa�D�sJ:�ӟ �	П�9���ɦ�͓����=sH�ITKe<���� B�.��3�:$�֓O$��?q���?���?�������ی�:�Rt��k�t`�(O��n��=z2L�Iş|�IA��ş�P&�%J8��;�+�H��Tx��xy��'(b�|�O&2�'*���e\� Q����	�C�d�VlCSj��,�<%E�dF�	T�ryrA�\�6��#-Z��*��5N�*F^��'�R�'��O��I��M�u�\#�?�G��}�jP��g]=��A�r��3�?����'�����o<�M�r �+/��iz��Z+j�Yzw��:pj ܴ�yr�'�.�[焀�?���O�����ڠ�'��4D*&�z��,�7<O���O����O����O�?�P2-��j��cł�S�D]`��	͟�����ȩܴQ14ͧ�?Q���$¸�&ų�,uqd�*��E�x��jӨ9nz>�������Q�'M�)t��Gz���F�6!��\0�=�t���,l�'>�i>��Iݟ���r�ZFA���M��ؙd�ӟ��Ily�"|Ӟ�ʂ�Ol���O��'n%$<j�)a�����D���'�	��M�B�i	FO����~A��#��4s��pc��W�1��j�:R��Q��	����?�Ё�'|I&��sQD�(H����M�] �ږ�W����	՟L�I�b>�'�86M�&U��Q�Iɐ�dYð���	��� ��O��d�O���'nN6V�PLࡳ�V�)��8#շ2���l�5�M�@���M˝'�O]3@�Q�S���A3�V@P�� :|҅EA(	 �ĥ<A��?���?��?1-�Z)�f��eA�]�Vg�0*���5��;u	�����	�����x�D�';�w�� ��A%7[Dt��'A�K�ڸ���'h��|�O]"�'��e9f�iU�dd-ч`F�8B��c��4h��Jr���'u�'<�	ݟx��g�� U!	Qʒ ���۵ll���ğ��I�$�'J,7m�KHr���O��$[ =��p1A78i#�L�2?M�� �'(��'��'ɚ|"w��:��
�t;�v�x���,�PT�R�R�1	,O
��Õ�~��'��:��'v����p������'rR�'��'��>��'R|�yÌ�+��hʒ�Y�v������Mӥ��?���?��w�x<��#F&�j��3K R���'d6��ͦa�ڴm!��ڴ�y��'G�$���J�?���4uƀ�wM0Bf1��Hׂg�'F�IƟ�I���I����	�1InHA�K�Ie�����c�.��'dB7���H�D�O���&�9O��xWɝ�
��A`f�p*��[)�<��i���d=�4������ y�/� *nt�sj]�r�΄�@"OW�
�x2�<�	2`B��(����䎟`���C�G�i��%��B!@���$�O����O��4�~ʓJ{��
�GsRN
c�Pb4H�={�b��J��o�2�'��O�˓F3��O�6��ER8񻶥��8�˓��8�Tx�%$oӤ�@X�i�P��miJ~B��C������;&���� �N<���?����?����?����O�f�HB,�$Z��)�Տ�?�놘������rߴcB�-Oh��4�d��
��q�B����- ��9%���O$���O���Q#+�7�i�T��=�~$ʄ�|?�M��k'Nij2���~|S�4�I̟x��ܟ���.�*��,ऊ��d��������ILy��aӖmЃ��Od�$�O��'x|��ʖ#Q�Hk�ՙ$)[)L���'[�	�����N��B�i�9�x��(�(y�Z�����'��ya��	�L�ꇧ�<���m#N�D��7>h0)6��k7��q������?���?9�S�'���æ�
eB@�{k� �5���3�ܗzT�������}�����Orux����;xu�!�F�4�Sҭ�O��$Aib7�l����fq�O�剂D#��g�Ut�`d�Յ@	~��`y��']��'���'�rS>�8"M\��^q�#��|�=	�)՚�M�2)���?���?��'���O
�4���HqB
�<��p3v��Y�8�2JͦI��4;މ��4�Oi�$h�8>���2O� P�C��U�7;H �Ed]4]9��3OR����ǀ�?���1���<ͧ�?�`%˗/o ��"�S�I�h��ŋ���?���?�����Iצ���E��t�	Ο�Z�&�m6\*�H�
���ql�������:ݴ�'�h}B���'�ҍ{��ÙaaN��'��)�WR����Ě���Y��0�r��ytu�b�B6 P�
�$D����O��D�Ot��"ڧ�?����Rp؀�1�]���Sf���?�'�is܅B�'K"�'�"�|�w�t�ZR���"��Hz�kżo�ј'u6MԦ�JٴM�X��4�yB�'�R��`���?�Z��q:G�S�|�����?��'��i>]��ߟ���ܟ �I�`�4��T��Pd,�vL/9x�'�&7- F�|��?����'�4��<p �>�jY����u�������_�i>m��͟��B�w@���!�(p�����=8�b`z�$.?GG=sq�H�������:��eA�HJ�^�Zqȗ7AA����O��D�O�4������j�7 �b�!UӸu
ek�g�>q�h���'��O���?	�Ӽ۴���p!����S�p*��1�N&I��bش�y��'|"a�DI�m�.O������=��h�!�T�T�T.J�Z��:O����O ���O��D�O��?M�sE��pߔ��@
6H�<�������	Ο ݴ�d��.O���O8�Ұ�@�i(�	�mG! ��yI>	��?����ܹ��4�y؟l��F=�t���E^R�|��"Ҏi`@��]�uyb�'7��'�B�Rl仄��_7���2ȌC��'���6�M;��Ɉ�?i��?),��<bGl�1�j��
��6TZQ�����'-2�'xɧ���'����nH�m����HBU}�Y�ꏳm)�0���iw���*�Ǳ�<&��ڲ'� r�~�xǃ���&3UES� ��̟D�I�b>]�'��6m	vV�c ���:D2��U�P�V�6eu��O���O�H�'[67��9)����@ḙx:mz%A*E�X�oZ��M�]��M[�O��*DE-�*M?��ƪ_��T9�&XB������i���'|�'���'��'��S1F��XU�Fx���2�B��
�vt�ݴ*٨���?������<��Ӽ[����,���J�|���MR�Uk����OO1��<j�`���	H�H,�6�F*��	�Dn�}<��ɓo{n`�"�'��T$�p�'�'8 	b�gƔKH`S�&0|��b�'\R�'��W�ش&�&�9��?��b-�y�6&�gB�,	n�2kP 1�⚟��IП�'�,�vJ�4�y���;XV@�Z&��O��3p��i8�l�m�<���"���d�6�y��+\fH�5��)�n`��O
3�?����?����?���	�O6D0QD%f!^=i��ӄq׆��B�OΘn�4q]0m�I�D��X�ӼK�K��'��p��aZ|9 �_�<y��i��7��ئ�
�D�ƦM��?I0��g�����z��]� c^�8V,Ց4��b:p��M>�,Oz���Oj�D�O ���OJ(��-Yu��ӄ%%�D��i�<I0�i��Q�'aR�'[��yrcY.!4�˅)�&&"l����?:��	Ɵ���N�i>!��ɟ��"�c�.��dO�핖�ߢcS��� �"��dA�mǊdA�AL�O�ʓY�v�Y1-��	{�u*��6jf(����?���?���|�)O\��	�/�b�$A���qR��5��M�b V���OP���'��'�ă�+i�Xٕ�ʗ;
&�9c�_H�����i2�D�O�X��kˇ�ⲛ������u�e
��B��`����)v�$���(�I�L�I˟��
Yn`,�׀�h��i%HL�c�����ß��	��M��|j��?I>	���ufz���')��<qq�Z ���?Y��?IgV��M��'��i�����:E�X/R�4�A2BT�n.l���/���'�ؔ'���'�b�'A���V�2ZȬ��� F�l��5�'X�Q�D#ܴ-�΍���?9�����	�5�	Ռ$���4�A�~N��ey��'��|�O��ĭ6l��C�.@*� ĆP�KN�k�J�f��O6�I�0�?Iҭ!�D�.}�-���>yJK���i���$�O���O���)�<���i���7'ܰu� ax��%x��dz�o�?ywr�'{b�$�<��m���6B��d���iAa���J�@���?㥅��Mۛ'����c���SXya��[F.9���5����K��y2T�������	ߟP��埠�OrY�Wc�Fj�D ���v��� �eqӂ�z���O���O����O��W�[���a���.N|YA�!
]����O<�O��O|�$NQ�B7�z��!�ͤ|��sR/��3sT�@�H�@�HP�'��-���<I���?���C*��IjDӇ~��,�Z����?q���?!*O`�o�v
[��џ\�I��xyA�P�3���3��;����W�Ik~��'eB�xr!�>�\w�U9keF����X.�y��'�Z���$R>�����U����J��+�şԓ��I���x��	5-������H��ߟ��Iϟ�F�d�'si���M�jd�0����S(W�Jx��k�� ���O�$�O ��ݴ~ L�Y�hӳB��B7@��	!�M��i��7-ǎHYP6�u���	(u� ����OLp6l��zŊ��FLE�5!r�S�IEy��'b��'S2�'	�"�(+�8�qD�n�Us���4g���M�c�Ȼ���O�����Ę>f��ԉ��G�bq)a�� �ʓRb���OO1���yP� �|[`D����a!ǌ'�
y3�7���1� m˴��O<�M>�,Ǫ:��(n���b�*F��+M�OL�D�Or���O�<	��O\rE��⵱��8v�����I�(-k���?y��Q�������FL�a�/[�^ ����<V�.� F�˦��'�X�D�G�O~���'���
2�U<XЄ��r�S�g�VP��?)��?���?�����O���ѨEL�'��X*ld�'#R�''7͋�c�$��?I>I�l�P��#2��IP�h�mM���?���|� ��5�M+�O뮓y��W�9��yh2��?r�,���#�~|�_���I�x�I�P��b�].�pnC�v ��P��ݟh��Wy�kӮ9�#��O����Or�'tx��� _�U��`VoKP�l��'a�	� ��`�)�C�'r�c	٠N�2(rs�І:t�!�����MSP]��Ӄ/���3���>l;2 y�!~ݡ ��$^4���O���O���<�i<���A�q�X`i].p��a{��I�?b�'PB�D�<A�iBޙ��O�3���9v�,=����$�}��n�{�N]�1k>?���HT��)7�
�f>��%��o!>]P�J��y�S��������	ȟ<�Iϟ�O�vTR���0����D�_o��(a�L,3R#�<!����'�?)�Ӽ����-G �  _1&�Ω��扔o���$c�@$�b>� H��4O��I�O�.��5%�m #���O���]����f�'�%�ԗ����'A��J�:\���*J<E L����'��'��V��{ݴ.�|Ё��?9�8��MJ�/������H�/��H��RY����4k���/��0B�舢����Q3��G�T�8���OZ��1��,tJQك����ӄd^Oʟ���g��8gO�5"��bT���<��ݟ��I��4G���'����|D�s�	�:ɐ}�q�'l7��?U��ʓ�?���w7����	)H���j�|�^ 1�'MB�'�R���<4��'M�j�|�\��+r�� mB8�"�A*Cy)@����|"Z��S�@�I�� �Iןܒ5�$
xL�@��%T��Y���Bdy��e�|؉F��O,���O2���$�*f�,QRh�*,�N 10Dֵ��ʓ�?9����|���?���Ǯ�8Dk���$hZ�J�@�f\���w�V~���ݺl�	,��'�剽j��XB�"z��q��DG,�����ئ	�E����#-�:#�,M@���khK�˟��IE�����O����OF���5�p����K<U��*rj�A�JX�1��J�����	.����^Y9qL�v�R��G#�#7���"�9O����P�8aB!G�)2{�Z��,�����O6�$���F�6�������{'Xn����GA��^v ��I>����?ͧ~1��K�y~Zw��MƄ�2u��𘢨^x��X:5iU�`N��.���<��"E��e԰���E����sB���O�@o����Y����IH�/ �2�n���ٺ<5
I�+���D�<����?QO>�O[����ڒ"�V�i��6B8�h���KkT��K���i>�YU�O��OD���DN?�  ��[�Ld��[O�\m�3^��%ؖ��(��5���Ȋs�2�8!�_ß����?!(O��3l�.
s�ä7��}����2^����ONU���+��i�=�AR[�*O��ȇ'�'z����0��6Jq�t5Ox���=)��V)3��Ѥ�%�
D����f�ӋC2��'�2�I�O�J�.A~$c��P�/�VY�"��J*���O�O1�
aC�ЀJ���#���R#@V~��C��/g���5�q�'1�'�	Ly�'$	�-Z��D*$�Z�C��,�0<�R�ix�K�'�2�'b�|��H�]��);�LA0F��<I���?�L>0n�2}��1�d$J�,,)S��I~RɆ=H��y���WJ�O��q���?��Ǝ{���Ԫ�na����M�<q�*�6P(J!Ơ��9�ȊWG���?�i3.�Zv�'�B�'��O󮇶q��w�C�\�@J��
�v��O��d�O�d�b�ƶq"�iݝؕ��{R������'*{䬵�ǎ������D$��j�8 JGL}���6Ʌ�f�H{e���q�4o�"����?����O�"�Xu	V�IF
�A��<(�R����t$�b>q�QA�.sJ��Db_<y�2
�-+ttN��2��ky(�|��������� �V���S�3L���Q+la|Rif��� �O,�#,׊e4�H�$Hߌ!����O��� �	ly"�'Fr�'R$�v�,q���!)T!lny��\�w�J�Z�O܂����ě���w�hX�+��i$&�����_��Pc�'��b�
J����� \�
(��_����'bgo������?�	\�l��4p3/��F�@�	c_� s�%� �Iş�S�.E��b�*5?��t|V�㒎�8�X�W@��0F�ʒ.8�~B�|BR��?Y%L�
u �@ �a�`l��;&�v�'��6mKs*��D�O��$�|Z��? j�բ�M�aDP\�רSi~�[�@���%��g�? ~i��G�xS@�g	��S� |�E���l}�M0��E�qP��|B'����'��ۂ
�b�(��G'��.&2��,:��J�4k'�)s�E��Y������}�֕3���2�?���?�b]���	n/����A�,��a5�_	#@���	ߟt��	�V���Ӻ������V�L"B�� ��T�S�@6s�5�"x��'L��'�2�'��'���H������D���H!&Y
$���4QO������?���䧖?�Ӽ�c�M�q5p�����6����ri�	j�6��OO1�6��/��5��DļzD��2��n�0,���3_��*ހ���V���O�˓�?1��s�8��e�?�T�*�ҧe@]c���?����?)/O��mZ
%:@�������$�D])���� �Q�c ���?�.O.�o��?H<���^!+�T��2n�=�)�%E~�eܤ="D��$*��N}�O>N��I�N4��7).M��T85B��H�95B�'��'���ߟ@��b��,���ǑT}4�x@P�|ش8������?�����y7CK�6@�RWDQ�l�������y�'%B�'�:��bK
����us`ɲ?qJ�o����AV���X����$Mu��yB�'Tr�'���'�Ң��6���p%+��o��n�$剺�M���?���?�M~���AK2���Õ5�����g��X�&�H*O��$�Od�O1�er��
���jVL�El!��#ߣ��5�`�<���_�y�v�IZ�}y⎙�rl�l:xjH��O��0>r�i�����'�T�2
V3R�X�͸"�	�d�'b���<	��?���bF5S����LtW ��ܱpfX�����'6|���bzJ~�;'n� )@�>g�y	$(����X���?i���	H�@&|h�`鰥��Cr%�	��@����MS��n�4�' �'x�o[�:��@j/fጔ�D�|B�'��O��:��C����F)T<	#P�S�E��F�̄��d�F��X�	sy"��P9{�X���ȃph~��b)O>�Rش;~T�B��?�������!wԚA�B��-f����Ǘ�Z�	my��'��|ʟ~��u�T61�
�r!�_7=�P9��9jG$(@�H�+[l��|°@���'�;6fT�[VPH�/H�g�N81�":�t�ߴ<7������j�XXk_�K����?���?�"T�$�	�Uq�A��� ��9�G��O4��Iٟ`�bI{�Ӻ3V�A���$P����J��i`���I��}�q-w��'s��'w"�'Mb�'��SZ�R�2��Qy�w>1�4�P�����?A����<q�Ӽ��h�2�� ��b?�yy��V��?!���Ş!�d�����<!����F���ᠠ��R�uY��N�<yiC �P����4���d��,:�H V�dx��c$�B�����O��$�Ovʓ#1�䉠<���'g"Ô~��@�D:g�pj�¾N&�O���?y����'���5�WQ{$	,�bI�'��x#FB��ڌ�$��̟����'O�ћ5C��6i��`U�I2�rh t�'j�'�2�'�>)�	=n*L��: ��K�"��e����I"�M��i� ����O��݀%@�Ix`&F���j��A)���P��Ο�r	%@�����&�埔H���-π���8q�<�a�H_�����4�&��OR���O���A�l��2i�T�:��GȀ-�ʓMd�Vl�*Br�'r���'�6A�ѦC�E��h�k�qKx���W����ǟ<%�b>q�M�'j�2w�N.��q��-V�Z���x�/?��KQ�m��D�����Ĩ�L��CE��E��`�7�����O����O2�4��ʓr�D�f&R�6��ÒMצu{ڵ
���y�'��O6˓�?Q���?Qp�G�7�D�� =eu�SPh��>SZ�C�
v~���ql��W�'���h�;A���P����h}+c���<��?����?)���?���4��$2`�0�����'N �0��E�`�r�'�"At��ĳl�<����{��)b��3PǓ�o0\�*�|�럠�i>�3�U�u.�z^���j�T�@���L Y�ڜaD�'T��DU�����4�����O���F
G�xd`��׵ ��c�JD���D�O��=o�6�^�Gx�'�BR>	�RM��&`B�p�D�4J��t,#?Q/ON�D�Ot�O��8@3�"�6��<G!�M�B�4Ǝ�2�,��,=?�'td��dX:��ڮ\��,^�=J��ҥd_�x�^ܸ��?���?a�Ş��	�������|�i3RW�6�lp
��U$�%�'���$�<��0�r�K��@�X�Z��!o�X���?�I����8�'�vQ�5cB�?U���%Є�߅&dtȻ�Kќ"WN�Z�Iҙ{$,�Ǆ�e�<��2d���LMAՏ2L$h�wI֒>o>L�pJדo^P�A[�K��7�:i���@m�sp�Ed���?c�A��e\��S�bI�a�y;��#��mڞ%�`��
_^7^��C�xp��`�3��E �b�D%l��F������0Z	J.Y �@�d0 ��˳Ut!I�\�c���OJ�N�:���^�ۆa�5j��d�%nҥyH$�	��Y�w,����HV�-zG��*\I	&��).�Y(+d�8Q1�Y�*�ٴ�?���?��� ?�O�����V˄C�[&4�,b�b��M@��9�S�OE"�)� �[N�R����ǜjvlyd�i��'��-G�On���O��	w��0d�ǁV�ؔ��űk�c��	�f4�	�,�	ȟpgL�(���`�c��\�:�Oʗ�M�F��RW�xZ�Mc������B�++�	�� ��wj�-:�}}ҦQ ��'��'�]�hp6)�Z���%OC�ZUؒ ^�'� ��H<����?YN>�(O���G_*Q�hU!r�[�V*ʙ���]1O����O����<�v�ТB7��%H[L�.t�� !�-�Jܫ2R�L�	�H$�H�'�����Ob�lC=%��<Y� �Is�%�sQ�\���I\y"��'c�D)���}�9����<`��\��iC�����~�FyB�Ѕ��')2�YE$�-<0�V�0 ��l��4�?����򤅳>�&>�I�?]YA�3<��iy!�٨P�(`G����Ms.OD˓x������4��F��c������
)M��pA�ݻ�M�.O&�/_˦qK��@�d�b��'<�93`�*z�k&C�� la�4��БO�b?���+Z�&��p �OEv0$9QIs�`5�Kݦ���ݟD�	�?A�K<��L�����5�Q2G�p���1�i\��ˋ��Ɵ�rf�P+9p@%�����!��3���M���?��� 2=��$�O��ɤZL�bR&�!�8���N�2c�����0��H�I�4Y�`�
%�w6���X0+�MK�UPJ9s�x��'*�|Zcr�eB��+j���f� ���D�O����O�ʓX"\yj �۴a_N	�Ē9I�����ߧb3�'�2�'��'��U�dPr�*D��H�N`Б�>���?�����Ā-2` ��';� �����=E��Us����{�H�mZAyr�'-�'�b�'c�U�7�O�]��Z�ma�١ĢQ�A�NY��T��������}y�I�;|^�'�?���.or���`_,H� �N�	+��V�'{�'WB�'>�BF���D�a��ŕs��;&k������'pb^�t(Ď8��I�O�����Tt�O؏�*�6(���4c��N�	蟈���#���?i�O���AU�*����&iZ*^�F�!ش���˿5���n�ݟ���џ|��)����b0�C�Q �@��CO
,��p�i~��')��b�'i�'�q��E[C�N03TX�Qϓ�� G�i�=jBf����O��d����'%�j�� r�PӞ��@�,xX(�)�4q�Xq���䓘�OJbh"���`��pPTpf�UnI|6�O��$�Ol8��-PO}rV����h?���S�G�v-��D&,>Dp�˃G�4�H`�<��?���OY��C��6���Ox1�lK�i~⯛�}6������O*�Ok�R�4 8q(D��`�6�h���!W6 �Iky��'�2�'��I�d�����2)�SlZ/s`��IH���<����?�T�y�EAO%?�n!�Po7�Ҡj���?1(O �D�O���<C�^.y��I�) (�C�G�l�xx*D�6���S�`��i�	ޟd�	�!H���	�|D�)�)`�SBW"nm�蚬O,���Ol�d�<1w"� 	���@�D��.jj=�S�-}YE��/ �Ms��䓀?y�>�`��{B��0N�t���hV

�5"UdΜ�M���?A)O��TK�g���'�2�O�8�Kd��<abX�I���,����G.��O<��Ӓo������?x�(竔fఅ+4ޟ]F6�m�Ry�J�2)]�6�Y�t�'��T�/?���}�.��a�5R�~qRu�Ҧѕ'�' ������v��k��{��L*jYڨ�ß��MA$I0#L�f�'k��'���)�4��\�Ʃyk�D@��I3h!�r��Цmp@�Mܟ��IAyb���']�:�B��v�.��xC�F�&^6M�Ol�$�O�R��K�i>e��{?Q�U$4K�8���],�,}�P� ͦ��I]y�卻;�h��<y��?I�V�0؁�Q?T.�x5�R�=[>�(6�i:��XG O���O��O뮅�K�ڬR��3r� �d����I�ۚ1��R�����'
r�=��`��!u( %�F7�M�3Z���	�x�?����?Y�DȨJ>�b�B��H��q�e���P�RaSU̓�?�*O �$M� �@��v��k�@�w�|��c�ӧnK66��O2�D1�	Ɵ,�ɛ9���"�x�tTq�J��@DH1cã	*��9��x��'-�ȟ�[u J���'5N�����^Ɋ�`BC�d�&�B�|⟠��ϟ��`bȲ:{lOj���\("9*dQ���}��X�T�i�W���	-�P��O�2�'��\cİ#d!@(�*Q�d�)bJ<	���?	�T{���<�O��ʈ�E�"�I��<{�z�S�O�$��u����O2�$�Ob�ɸ<��,NUh&�Ӝ���;���c�t�l��x�I ��d�c$�)�S�I/ ��UAL���%�X6�7��U�j�m�����	����S���|r�O>3x�H5O��4Ь��6� |~�v���"�'���J�3?�3�W��8�Х@���B�x���'��'FTH_���-�@����ʘhr����i̓1/x�a6���'tb�'��W,�$ ��	�("LaQ�lӎ�d8y��-%���ޟ�'��0+S�xX�Q0�ڂHv�ya���$�<v�J�d(���O�ʓ�?i�� *����Y�2�t�dG��<<�C%Fƚ��D�Oh�$=�I͟����-��-Q�c��A��}��ʆ=Y8���*�c� ��yy��'&z��؟�@ ���R�]/�����i��'�O@�d�O搨cADݛ���~CHI��B�����A�<�듉?a���?/O�4�@�L~�ӊ~ov��ׄ��K�YK��K}����4�?IH>�-O�]�FM�OB�OԅQ�,�9�<�xѬ߲I�@b޴�?Y����$ܗ(�%%>)�I�?�؏(���g�|j9���Z�fOʓge:a ����'��� -E���!���=�Q�B-�?�M�-O��#E�Fצ�������y�'��*0~�,�QCƟ;x����ߴ��<`������Z�s�µ3a_�<����Y;����1�i�8p%�'��'=2�O#�)3A�4R�rp�`�O$A�iy%��i�����d��	��y��I�O0��#[5hdT҄��+�^�!��妝�����ɟQ{2���OT��?��'����J�GR���E�?0~l ��4��|��	�S�d�'�r�':��bG.�-Ag�z��+ON��$Ov����Ƴ �&��'��՟ �'�Zc��|�b�ă`�B�ۓ�
=�<���O�	{����������	���'�*1H2��55(��tML/;��b!ڼ$������O���?1���?���G��+�F����(a�r�R�kq�,�'��'��\�H* $�����O��&�>�2� :wnԪ�A�M�*O��Ĵ<����?��EK��͓-M��)q���Q�D��,��$�:̐��i'2�'"b�'��I�*0 �s������*t"�1�����Pzra ,
��|lܟ��'��'q��y�'�&n�x�bEi����4{�
@0���'�bQ��@�	����O��dퟘ�3&L �C�<�΋)zp`xj�ώ@}��'_�'�����'�U���';:�Q�@8=� 5r��(�@Xn�@y�II��67M�O���O��I	f}Zw�>m#��2Pwx���Z�I !��4�?Y��<��'��	a�'i�x���Dޭt0��̘���oZ-�p��4�?q���?)�'R���qyBhܾ0"��@j�{��9��eE}�ٴd~��͓�䓇�Of�$�pa�$0eG��1� ��<�P6�O��$�O �ɖ�J}bW����B?��@F�L�H�b�J2��L�ӊ�¦��	^y����yʟ����OX�dF0�T���"K3p+���1L�x�o��dHō���<������OkL�"�(��*\v�`)�r�Iq����r���	֟���̟L����d�':n��l+�(�i`��29�T �$�E#2p���d�OBʓ�?���?��v:!����l8�e3"��,��̓�?����?����?A.O:8cb V�|���i04��h�~X�Y"bE�ݕ'j�S���IƟ��I�\�H�I����KuO�^a)�B2��۴�?I���?1����r�`��O�".�(^Ȅ����,z�p�(�b��`�f7-�Or��?���?i��<yI� 2  ��|U۷�/]� �֣w�`�d�O4ʓ��@'_?E�I�����x]�1:c'��q�L��EL�!�8D��O����O�D�u��Imy"ٟj	��ڌ*�.!vg��,a���ѹi��I3X|$۴�?���?��'<a�i�M ��>it8�4��c��ع',p�b��OJ���>O��d�O(�(��A E���H�L�?}@7�byA�Me�J��O����D��'��I�@x��7�"s~���ք2�ɫܴV��������O���޲d��Y�f!T�rQj�R5�Ih>.7-�O:��Of �e}bQ�H�Iu?Q$ʟ�fj���@���6aRBA�ݦ���͟���&&�)����?���B��@�i�#U{B����it�;�i���z�p���d�Oj˓�?��1�%�h�4\D�P�jܕE��'
䭐�'���'���'1�s��rR�L�Yk`M���I%��AH���,��d��O:˓�?Q(O8�$�O���П�L����	v�t� �\5�4QW:O ��?���?�,O�I�����|R7J�#���0�HJ���SG�UԦ	�'&�\��	ԟ���)���I!z.l���I�'^@��CW���iZ��ٴ�?9��?�����՞_�.��O�B�K�k��z��];�3S7M�OX˓�?����?I�I�<�H�d���n��m�W�Mp��uCl�X���O(ʓ.��8DV?}�Iş��ӟ3���:�	� ��2�[0a��کO����O��đ�=l���'UB�F$5��Qq��)d�-m�Py�nR��N7�O����Ot��i}Zw�f�f(ӇL��`Ӱ*T�s=�b�4�?���P��'���vܧZ�B,�P��]��4��a�z� �l
F� �ڴ�?Y���?��'T��`y�a	)X2r�1�TL���;wF�c&�6�	X,�;�$&��ǟ��qIԼE��8�BN ��{��Y��MS��?��](�9�V���'���O���'ƽe�İ�
`��8��iW�\�0�o���?���?�����da���J��.�p5@�U����'NL���M�>-O^��<��s�g�$ ����q�����I<���cy��'��'��ɬTq�a V)2,	h�+���2'����h�����<i�����O����O��	 e�6f&�H�͊�8N%�!��"^�d�<	��?y���������|���"$�M(� �oX~H�#�ŦU�' �R�P�I����I�#�F�g/:i���_;Wl�(��� 7�\l��Iߟ��Ky�LE6��맓?�q�? (��@�H,��(�Kİ3�PX0�ixrR��������	E*���[���B95ľ��7�Bf�D����!,c�7-�O��D�<�e��܉O�b�OԾ+��.�J]H���?g���#�6�$�O���+{���$6�d�?�s�n�f�Rq��k�v���wӬ���Y���i�p�'�?��'G��	?ZT���`ߜo��$`'��<�`7m�O�dƧ.O��?��6��l��I�`ι��P�ń�#l�7�.H��mZ�4�	ڟx�Ӌ�ē�?�'�ьg�6�3'�P+D?@@��+��T%��O׍_���|����O�雄B�
?� �CT*�`Yvf@��%��㟌�	�E���3�}��'����Vь��w��������{ܴ��GlN������d�Ol��Okl�$%�D�d��z1�1�ƒu����'#8���@&��O����<Y��Òlݢd|f:b���1�b���e}��%}�BS���	ȟ��IMy2#�q<��B�X #x�s�&�[ (����3�I؟`&���	؟�H���N;��+r�ݮm��Ģ��^�;��zyB�'�b�'��I?s�u��O`�pSէ�;��8Á���Ia��ҫO����On�O����OX,�2O��R��C=B���(�n
�XqlX}��'g��'�前e��jI|�P�#`�d�o'�а!��&A��'��'L�'��#�'�C�& d��*-2�vg�<I�.<nZП��	fy��4\����$� �U��]YN�!�%	�Y2��ĀD�	ҟ���rurx��h�IkZTNY���x*S�<HFD#����-�'Pd�H�Hzӎ��Od�Ow��C�y���Mu�D�Zb��..��l����	�E��O��OF�>AY�$�QO,�kQ�M#��2��}�:͘2�W�A��Ɵ��I�?��}�$�2D\	�`ς6;m�d)��Ф��7m�j�-�D#����p�G�N9f���^��b������o�͟��I֟���EA5���?Y��~�@$A�Ȫgհ^�n���e� �M�L>!�&I5@D�O���'�I��b�b&�����<�sˬm�7��O����BNW쓝?K>�13�s�@��@�X����n,��'>Z	K��'��	��H�Iϟ �'Ezʐ�;&� %��**��
�3GH
OV�=ړ�~Ҍ�5Wn����"c/�}�d-Y��MS���D�O��d�O�ʓ[�<!K�>���2���z�|KAm�/�*� P���	Z�'i��Ο<@�F�A�f	��N��Z=� �Ċ��d�O��$�OT���O� � �|z��� ɪ�	�D��)d�[�>ښ9�5�it��|��'u剞#|O��`to�MsF���A�c�`��ļi�"�'q�I,!�R��O|����t�

b w����ш�kX>p�6��
l->��sӂD�!+� T�`� �*h���Ar�i9��'2$AE�'a��'�R�O��i���q�.q���`�IyQ*2%n���D�<��g�n��ħ��B�퐫;� ���H�	GV�l�{I��i�4�?i��?�'A���QylW�zf��ٵ�F� 1�GȊ/+mF6MA,[��$ ��,��՟����3����SeO!�Ф`�H,�M���?!��4�ڭC�P���'��O�V�S&vv�E����S�dc�i���']�,�yʟ���OV�DX�
�0�� ��;��q�j�,o6�mZ�|C��(��D�<����d�OkL�wL]
5�Ƒ nR�8&
D�^\�	B#��	����ǟd���'`��Ʌ$e��8a��
8ji�pNձ[fZ�����O���?A���?	��M�x�F���":H�PB����T�'G2�'.2�'�剞!C�L�O� ���A�Ϣ�i!�?��ٴ��d�O���?���?�dF�n}R�C/%^��C2M��X�&(���M����?1��?y(O��5�M�D�5�j��sP D�������D�K�M����O��D�O�[�5O*���#u R]`x��Ó�esjh��"k� �$�Oxʓ� �z'Q?���ܟ��Ӆ�N����+J�x�x��L9gȮd��O^�d�O��Dί2@�|�����8>}���&�թq�:X�T��M/Oz���aE妥�I����I�?M��O뎜V}�1sv)Ӷo�Ĉ0�[a���'�AJ�y��'���'�q�j�V�,�n4�bˇ��`5N�զq�7��)�M���?����J}�U����.Ё]��0�$M�j��4��Mӑ���<���� ���p�U��cz]�Gg��v�"�{VN�M��?��Z�m��R�\�'�2�OH��T<����d�³j\�{�i�r�'�Α�yʟ@���O�䚻�ɣeػB;0��b͖� ll��EN���d�<����D�Ok�S%;1�h)T�F�x�����C�K���'a�'�b�'7��'��Y>�BG�.T�x	�G��Kj�2A�� ����ן����L�	n���H�0t�a�w�[�#�m�T���o�FDl��3���?A���?�.O���n��|�',�"�� )!=f�(7B[}��'`�'��O�p��S?�3MժM�hѓtBN8phF���>y��?����?��3mH*)����*:5~$IT,�z,��@*Z��o�ן�$�P��Wy����ē-��1w O�����c�?Jy@Y2Q�N���'��>�	����nɸ2��t c✶R`zB�I(3z�|�G��^��X�pd�!{�&����~�-�ukM6V�Q���-?c�I�ҷN����!�(S�v(Rr�*� �}��	��_�|����P�x�I3*�:#�8�fL�$IaF
ڙ>�:����kҬ�!c�|��m	�(�07Ĭ)��(JT�d:E�ؽP dbc��s�D���B8o>�-����:T@���O�O`���O��$�κk�دZg�ePʐ4��[@b_�qY�݃f �J0�$ �n��,�T�1�ӗ��/
άPUӹ�<�� ��(�dD����e��%B鏰B &���L"��7}��X�'�6�h�N%D�X<�HZ�#�X���'��I5!Gz�4�أ=�e.J�kZ����$H>!bL��DI�<�f�0t"�����I��E0g��B~� ,�S��_��f(�^�|�b@��>\l)&bB�?=  
���������I��Yw�2�'��:��+#��	@,���ug	5r����,ܡ"=th��W؞�BCU�a,��F��ܳp*D�!���k�#�}�ycۓ|�p�P0D%u������w�QTϜ����IM�'3�O���b��Tste@�Bi����"Od�"���"իf�E��@�ZF�$�p}�R�����4��$�O�l�6œ���-q��ϯ5�R�awg�O���i��$�O��2����C@�%Ѱh�'��9��-ݻf݈���Q�C��KǓ\�r�ZQ�w������OХ��1Jl00��G+c`&1ZG�'�(���?	-O�%�q"��?K*-�h�g4�8��&|O��[eΚ!P ��@� �~ H�Ov!l�Z�٠�ː�lG�p*��� � ��Ky¨^0q 듆?9/�6u�	�O&��2��'��j���-!�j�e�O��d�9AY`cqh�H�O�M�D&����0���� B�-0�J��uV*c"��0
�)��IдR�n�Y�Ic0�	�h��q�љ>��`�ڟ\�	l�O���6u-��'�[��ՙ��ِ�yB��	t�Q���Y���0g��0<��IT�6�R�lV�%5d%R�ʞI6\lA�OL��O�*�%W��T��O����O�*  8���8G�f���/D�ar�0�!�L�eFT�I[��Hj%�#�3����4��=�W�	�;�+%)�=`�TK����H�@���,e� }� ��|r���#"ph:%�
�8R������h���O�)$�6��bЉ�L��ps5��?�Ņ�o�H\��l]���)3�6T�F��'�"=�O���-b(���Q���������DU��X�7+� <�}��؟���џ��]w���'P�7����%@Ʈ����l�
o;<HѮ3m"�x[ҎBX�0iǓ[�jApa��Y�T��Peݑ\�z� �	�;7��;<
�`R#3O(�"닻M#����)hs�|��bZ�
�r�z�xXl�T���|��P�4-�^P�#�~�e�3"O^�:1���-,43g
ֳ]z�P���ID}"T�0�&nт�M���?�F��>����N��BnR��?����nxZ���?��mx��7)�Nu�a�_��?ap��"@�$��hL�J�����!�u8������ȱ�T�NT�ڬ���Y�W�l��1���l����_�;�l���a�B�'	�7��O�iP��V��)���F|�q	��<����������E��^�PS���cm*����/�S�O��6ߖ<�0�s�T�q6���^	!�`��,��hOn��qH˒B@��#� �G�\��"O.�HE�$ -��r�Ƴj`�!J�"OH��LO/0�e�EŰLj��v"O��%�����ƕR� 9
�O��y���svUJ`���� 9���yR��]���B�@Bu��F��y�J�<xC6�!���n�L����ʠ�yrK��3(b���d��a��-�SjT��y�K�\�b��F�Ш]P�,)׮�y2��-������Y�y�CB�yRŗ�� ��F�^S����ˌ�y�)W�w��)d��]!�8a6HN9�yB�։2���L�����&�yo�<]�,�À'V0A��:�@��y¤ݡY� m��+ծp&����y�F!�2ԣ�� �bb��ra��y2�h%0�u��	���&L�y�[8��4��s��M����y�$�8.�J���j�X����d��y�P��NT� ��!@\Y�s_�y��߿V���)�K�9q���@�1�yR�/f�}��#��DS�������y
� �}X��>9"�mPt1B��"ORr έD��"�e�iÈ��"O�� fEI���h�Ӄg�؜��"O�Q�BD�D���)a�	x��\K`"OP(Z���_��I�%%�"O.H��(�(MA��!�Ά-Ѣ��T"O"	��MC�J�,EZ����B�E�D�!�I�V�X��Uk��8�1� 8Z�!�$O�.� ���j̡Z�]Sg�F��!��J*��A�P�L7F�"*ө*�!��-'D9
`�W6(��G9<�!�d�o�@Db���>�E��E��!��BY��D��- ;W�%R#�-�!�D�~3����ĝ��(-(C��(�!�DNp��|�5��o�՛r�Rs!��G���U�c�P12�TU���
d�!��#z �'L��$F���$B�&�!��/o�8-b D��v�(�m���!�dA�W�V�&R	F�:�G͇�M�!��Y�R��Ӑi�d���
�f�!�M֐T7 L�~������Y!�܌ie��Pà)Tp5b	@��!��C�9�L� ��_H֙`c�K+V!���|&��6'�91��b�6�!�D�(�"aZ�)\0T3���5o�!�-���#��F�<Wn�M�!��=��&�D/�ɂ���2!��aa�칆l��8 C���kr!��P�-1Ġp�GO�$�걠ц�sq!��1�6����8�&����݉]P!�d[/;u|d���@�TPf岂G�p)!�dI/4�:H����gDrH��ڪ�!��űIK��iF�֣\�\e����8�!�ه<����@N�+&�8��;7�!��5ef�y꣌�%r��]���&L�!�HU�̒2����(�a��!����QMT�g���sk!�נ{!h����S^@�&���N!�$��E���4l��~>�H��R�:!�䈟k�("3]2">ը� �&~!�$F9{�y���L�6�<���o!�TaD��T3�á�
���'~�3�C!�꜒0���I��'�lj�L5G;��J �{l�܋�'KJ����������B=zu����'��Y`�@��<��;�g3q�����'���9�:r�@���/e��1��'����!��6h!�`H�Y��e+�'K*Yy �ȋY�<���D����
�'�$�2��4�����9*el)�'m=8�Ϛ�Pm`=��@Q�xL��mX�O�c�pE��'����F�ӓd1���4�w �E �'/TL[���O
=���uH>R��1P*p�1�O*չՉ|+��C�F��^�p���'cH��c}�ǥ=-��QBg�!,�&{��
�y"�ETӜ5���N�a �4�<��'��A�gF%�'O�h��E�9fចp�"�$M\���x�8����˰,�li�ͅJI"���9W�EEx��IK��$ē���^�1�%��!�$[�q xꠦ��Vb��c��2��e��hۓ �,�(��*-\�Ia���Ѳx��I�(�`oZ�?�� �J?�r83B��D�:C�5h�� j'��bg���!i_�udxö*�r.�d����I��?��;_T�p ���))6E#!_��S�? ~�ZW�.x*4��:�Jb��F�q���	������_y�7M�8��S�4`I?Wt���M��>��Lh�Y��0=�&�Q�mn6,��<��fImD���X�2�xH�E�ӄ��pLծn�ui#]��'��'Q~A�&�	�,��9z��]/X��+�y�\-P��k������yZw��ɠ�e-D����
t�+~��`uC�/u�@Y��'�T�ǉu/���'�1���c6`Oxy��Oġ�G�	V"�T��A`٬j�n��q�!�`Z�T��% J��y&h�t��<�`� ɇC$�I�&�6ol���	�#�yRMʮ4�m����h��?�aS���S&H@�`��+	 ����a1LO0`��ǔ�Vp�08O8�����}�3��f144�KL(@��7#ɧ�?iKS����'����J:c!l����ՀPs���yB�ԂT{�0���(����dK8'��Ub*��hm�eN�^Ͷ�q�EF�En��:���f��xc
�2yP$��
#\�p���e҂3�PQk$?u��f*�U2- 1�s���{e��I����U�-܈][��<^ONC�	�N�� #뇌���i��3�>����0&�n������F��p;��
�.uN`��iv�|R��G<9hyu���b4�p�a��V*%5�(����yB�B?'��3�ئӐ-r��F�4��0t�ЌU�lm�n��J��|�fV%�psgnކF=I��V*��'5,	 �W(=evub��iFR�J]���F�v�P'�W}��)���5k��fk��|���I���MRd�)y��D9V���:&��!�с|���H�i��L����$�&LXm�coư=�� �ȓN�������?�s4��R7�$�#�`e$n) u��y89F�tO_�㐜z����T3� �QO_��yI��Pb|h�p�X�^����EL�)<4�!Η�H���D�����L���2�4�im큆>�^�p��94����M��)ڢ�ȝ��1B&�(h���	�۔��hFX��`S����!*Zy;P䇛=��q��?�O�1��MW+<X�6��9&���:��ċ��P��8��'X�L�Ҧ�?%�bI�0����';�A�""��b���T$�Kx�;	�'���a���6���kT�H~�"�q�'ˢ��b��	Z�U��C�%\�4�
�'a2����-ؼ�G˫le�@
�'L��ŕ3"!� ��k	�]�`(�'#���E�$-��ة�d�c�����'jY)�+��f�	�2�.k�-��'�����Ⱦq��uC)i�B*�'z\��Q떧3�J���f�fT�
�'�XrD�\*6=^1��+�i�^�	�'�JT�&
xv�pdIU�^>Q	�''��:��).�����R���Y	�'��PN�|�$�V�^�Li�Y+	�'���Bs�S!�i�h��J+��	�'��%0rN�zI�U⟖u�H��'U$}�Chr�1�F��gI����'�l��ɋ@N�D�RƆUwp�'EN$2%+�O�(�4蒁6X�U�ė�27��Q�'���P�&��P�RD�(d��1�i�M8�ّ��2D��{��ߦt���['}FJ���e3�[W&�;@�H�A��8f���KàF�t��B�I�������&tK�y���@3G^ƴ�����O?���ahJ����r��$��	��hA!��;�@!�Dʮ3|FP8���#��	+!Zf����0#hj��G�Nc��sU=Z�!�� 65"5p��4]�����^�I�!�N:1�Uч�pY�I)ѡԤ�!�d�3����2.X-TJ��3!�46��ɺdM�"<E���]!jfD����� |dH(��>�yrOC?Y�.L
p�O�ּ}���@���ެ]��O�����V9'���k�%/�Ɯ���K����$�@�:���Ȧ�C<8����pA�{�<�Cϊ�Cn�i�Zԡű!�������#3�$"|z���4�|ȡ�4{�d0���m�<	�i� ��Ū�_�Jtق �ey"c���OQ>� ly;��*�����YOZ,;s"O���E��A�,�Ӎ��?~|P��|R���7az�hՋvRU$m1 UaF�Q��p>�ԅBժ	u��{�}��%�iGL9yG�]4�C�I�\��J�4r�sT�׹aRh�<Y��G�X�"~� �02d��(����&jF��eTJ�<��/�l��R�ʹ^��kp�a��"�Wm�S��?�%��9�t�r;��U�b'B�<�0n¡-0r@�7> �uA���s?���.p���$§H��h��Č�"�K�Aj��|/T=�)ϓy���sAM d%�ms���'4�ȓ
ݲD�1 ^?�B�zp��-p�Fy� ֪բdG�������뀌ײX4U�D���yr.Ѓ �D+��J�ZƢ���:{����J������« nƜ=�s�W1Iݤ���j͒�yB�!�|����C�P$s���~b�Ե,�\<��	�]F�P᭖#BH��� �G�"���@��eΓl���ǯ��~%)v��ZB*p��[Jف��3C�$Y�kӶ-�Tt��YL ��P��1�4���N�LUd�ȓ[��˂BBU�>�L��<�DA�ȓHV��SF����Y�� s�݄ȓ��]#�g�gIh��C�1.`�x����s� Q�%�&���ᅄl��y��98�0��@�t�ʩڦ�\�L�ȓ#܄��儹�q�5�D�[a8L���I�� �+@.@�j��8 ��`�ȓ�"0��'�����5}�(�ȓRbXp ��<�.l��L̴a��ȓ@��$�+|V
���C�3N0�ȓj� ���G�%9:	�3�O�M��d�ȓY}|�P����|>���N�3�&��C���l�K���#��= <���ȓ]8D[2�Z�tr�A����#*>���K��	�`��	�֕J���PxBU�ȓx,��@I�[.8�ɋ��݇�Cv�h���F����'5�ه�E�Ƹ �#l�5��W-)W��ȓ*�DC6n�&���BÁ�%�fY�ȓa�����j����*e��`J��ȓI�L��"�1
7�@�a'�>W&%�ȓB@@y˂���Mݲ8���ݞ!bd����`HG��:kK�2#iG�i�vчȓ6s�(˧Ύ����D�k�d���T�lQ`�O�t�܁-U�-+`L��G2\cK�7( �iC)-�@�ȓG��c�\:il.���)��|ODA�ȓ2�v8�(�,���H����=  \��%��4iA�˅z���� � ���n��� b� ���&��o�,��ȓsR� ��R�IxRkg�/b�����'�:lɳ��ژr�(W'\����ȓ6�P���E� 0q�@օHO��ȓW�Kw�L�K7� ��@��)�ȓ9��@
��ܾ1�z�c�������:q�N% gjOBx�e�Z\�<9�H]�!HQH��Q�2 z	H]�<1�%�<W�ȬS���4�̭�a�Xn�<)E�Ɂ&��j��,*
�[���r�<�4��0c��ͧ ˖��7h�T�<iDL_�O�Y��c�Z�*�Az�<��'9g��� �<�A���s�<�qn�#e������(��Dȵ�]C�<A%��Oލq����o
rqR!�i�<� @�Q���.���v�9v-Ѐ��"O����^�#@�������!�m�u"O����
�L*�� o�w����"Op(�Fd�������Q�Ru~��'"O䘻$C��Y�vdh4��
S�b�"O��CY	.����4���Ʉ"O�<j�h@&X�)�0�D9{�H�'"OH	�%H@�ji�t��b���D�@"Oj���')V�
d�aM���ȱ"O�- Eɐ�Q� 9)��b�����"O�$��D@9D<������)� ���"O&lj�͞)�L}"��˘?��T��"O�����Ð4$J�;0�O�B��XU�$?\OHy�C/� eۆDr��f�
!�a"Oȣ�ѝy�����Q{�.uz�"O�p��$�X-J�F��Q�,\�@"O�0������1!�
|���"Od(�@S(5|2����MZi�h�5"O��ч/�@��͗,-����"O���'��M�� ��e[��>D���㊋�jWx� T�+(���CS�;D����	�N����!�E�[�1��9D����U�6��d��#A#�y 0�9D�As��XY"�K�\^���B�9D���LD�p��y"��/#����f7D�����ѷR���pdTb��3D�
Ʈ�oϴ����51�^��/D�|�7nL�r�`4c�V�A�,Br�,D��bC#ۮ2�)!2+'.y ����*D���$+h:�9FkΒa�#�(D�`�g�����p�ނ'I�tCu�)D�@iV��Тsi?3��ܢ"�;D��V&I�@l�#�*S��py�&>D��j䗸v��鷈�60@��@9�$8�Olu���^�1�Y�jC�~Q�"O�\���+yPL�Z�IԤP$��q�"OFu22�1�&�2q�ϫ\���6"O6�8p���d�,x�3�]P�"O�m�W��1:��r����%�$"O X� '��ͥ
�em�b�g��yBh�	FBuPad��p��y�,Ǉw�*!�C�L9.�\�A�T��yb�@,T�m31�.l�L�1&��y�n�-��T���H�!��@�i��yCP�y�2�1��
q{�Qek
>�y�o����c]@���K	��y�痴`:��S��+1OPQ�A�^��yb.m�i;��)�Z�ja�Ϯ�y�l�'�w��x��iD&M��yBE�*d#�<�0eĘ�n�����:�y��	 i�:�K�@^�3��Yy��ԇ�y"�ڱ�b����#78蹧��*�y���@ab��2�Y�X�%�Q����y��U3	 e�%Ōg����ֲ�y",m[���$@�&/��!���y��E��y�d/ۨP;�D�p'ݍ�y���S�4�����9u���pKА�y� Ȋ%(����*��DC "��yBɘ;mݸ ��)�V�<P��*ѳ�y�+��L-Yd�\Cr��YC�#�y�)X�@B ����׏nF�h���y"EW�0����.�\�t�p҈H����)�S�OX��ڐ�L�9G�h�#�Q�n����'{��A$ͫ"�)���e;�<���� �y��,��P��K�%2��"Oġ��[�F�(�1�L9�A�E"O��0&�KChLKV�QZ�k%"O�4��;?W ��f����Q"Oh���LQ�	$츅����ܝ�W"O�L��e	N����r`H�WD�գ$"OԽ�����if�<*7��k�"Oz�z��F)9�������91b���"O����`��Gx���-�,Y�&� "O.2�S8A��p ��"D��ԚQ"O6!�W��b&$sR�= d��"Oe����{p��z�C��6&
��W"O��&-�\p�A �9!)6̸�"O�,�(�_/�4��$�Wt��"O��&l��|��)�w�����"O�Y���7Op�f��0�D��e"O� %e�j}~��GJ?�peS�"O|i����>� ���F��P�c��'��d�Ď)@Ӂ1� ����K�A�!�DI>be�El��t�p�qŸ@�!�d�%�l�y�
H�0ܴ��� �!�D�W�媠%����$�� !�!��R���23�C�tj���/� ^�!�䐌[v��0g/�8H�чJ�~�!�������C���=HΩ[Ѭ�3V!�Dׄ0-ĩ
���D�e3lĉ`F!������(ʋ\� E9f)LH<!�W�&<�}k���'[q:D��h	!R!��0��p��~R�옧�7B�!��-Yf~%;dnT�i�h� D���!��!5;�Q0���|�d�2���"�!�D̡����OߵY{���p�F5�!��M^�,)�"Y� {��E��a�!�؏��YK׃��]q���J��W�!�\�o ��e
fp �,A�}�!���m?nȋ��L��r�u��[�!�İ|1 -�`K\�o�F�{ga��
+!���r��a�pcU�C�R�u��M!�Dĵ-�Qv�.H״�P����k!���`T����q�d���K;7!򄃾hcҍ��S�Nl!T��%"!��'�	Y�锪q�Vey�L^�d	!�dϰBK�=9Հ��N�X�L�<`!��U�%����H�B��i8�e�.Y@!�dY� ^�Ps�ҝI�Ё"u$�*R!򤄭!&�8`!�1�R}r��v�!�d5��0���T��Ar&���&!�$�#O35�Т�3�(U�LH�!�d�5�DѰiʸM�JA�sc�`�!�Ȫ���ڐ�G!N��%�����!�p�߅{��!��F�pI��"O������z��遗u>�I+�"O��:@ ��.�^�`��X�N8�"O2�+FHS�JbۼTٜ�в"O8lAg����y3D'M5k� �r�"OH	k%	0��V�^�z@1;�"On�#c��	���2Ck�	�l�["O<9ɱf�6�[�O� ��P�e"O$=���Ϯ5j2��⭌�B��B"O�\�����_��)��KT(O&J��G"O�l�	� 	aa�L�7~�*W"O��*��e(�S'
A�g�P�5"O�|�T�c�� 3L	p���C1"OD�� �R�@%2��'��AK��"O� $h�栃�x@ƨ�-a_���"O��{�K� ۠AY �&`F1at"OJ����!j�6��E�MVB��"O��� ��<߲�isa�xTRę�'<.����?J#��G(Q!��
�'����a�	$gr�v�Z ?���
�'�h�D�Ҩ=<`��4%�����D*����rɄ� ���1�^�&fJ�`"O�Ep�˯*�6\��N�
8e
2#"O������N�����F��Y��Ȼ�"O��)��	-qh�񵈎�q:yI`"O�LRsĂ�������9�<�P"Ov�V/^G��y���**XH��Z�ԇ��(%�f�s���&/h�[U&%$B�� |j�`�B�4^���!NI��C�I/�| �"tL� ���
��	TX���7�3	�$| W�"c���2H6D�dㄮ����U���yE�5��� D�4����3<�(��� �=n�r��!�?D�yF× *+�0�d���h5�$=D�PB��Ѽ�I�ē�n�r����9D��A�ڳ7�`�����h���!2D�x�k�������͠bjh� �$D��'U0)fmb0#�74�-�U�7D�����F"H�K\�+�8�F��X!�&x\JC�O#sh°����&�!�d��L��5�҇0L`�Q�N�/{�!�Z�>w�m�0�Y�a�BT�VG�1n�!�Ė4OM�hs�Nō��`�C��
y�!�d^o$|��j�}%"����N9�!���B�L�-
�hhi��Ù$5�!�d�ah��g(�6,2Eص)X��!�S�;�*�eM�.���.(x�!� $a����}D����nΌN{!�$G?S���`�#��l �d�ݟCf!����
݁�(��2�D�3�E�AW!�$�o*���W-��$׀u����,uN!��Si3�E��������%im!�.Vز�٥�=Ѽ�Q��� n!�$̓�,�BB\:C_����,3<�!� �K�V����BR^n�HW�ۣ!�!�� }��k�HƁ'A�4ꃍڔ3�!�3"~Y�aǕ�.��L��Ǝ5k�!�dԧ'+h@��J�g��%�6d�2V!�dV?e����ُr�];��Q�>!�D�A��Ӕ�E,b��C�4[O!�Dц6�L2`��v]��Еʙ�1!�Th���p
�oOԈ�T��1$�!�(Z���׊�mL��8���]�!��ߣ`��[Ti��HH\1�-�:d�!�� n~p����C�r�J���&ɟ
�!�D(V���+�F3��0Ia@���!��4Wʽ�E@Y�"�h�Ⅿ�!��3A�$�8�fӥT�X���P�f�!�WF<ٕ�Ҹb�ES�5B�!�ě�5��ɣ#$ޖX�@��d�!��ւc���*��Y���8t�0�!�DZ,J��h�C��`�`#,�!��6�Ptg���-ҖB�P�!�$F��`�l��@���u(�G1!��ww�X􌝶2�E#��?!�$�$� �WJ0i��f� =`!�֋k {�K�Y�@x�oR!��C���M�Sd(7G���L�{P!�� ��8g�##��8�0JL�N��)3C"O�%���I�i̞=!�n��j8�r�"O�&f	�j�}�g֠hK���"O
�G^3I��Y㇂Mb�c"O���q�ʞD��"@⋉AXt�d"Oh� ��J:> � B��aE���"O�irpܛt��h��[����c"O6Y���C�$�b6�@ �B�"O��P���'h���m_� b�"O��2�X�V$S��m �Ap�"O�p!e��4D�aB��/���ʰ"OQ�v�IQ�q�W�ڹ8��}BG"O�R��*Zz(ś7掣&�v �"O�a���I {�"�c���b�¹�f"O8�ˁ�N:Y�0�,�lD�"O���"�
'�hŨ͖+)v(�e"O�UJ�5A��mK�&�%Y�n��%"O�)�����8���r����"O8E�h�"+6ܤ*��U	A����Q"O҄@���K��mr�#O,e�Ht"O�ݙ7��DH�2a�W�0bC"O~�h�W.Byy�,Լu8��ˑ"O��ǯǕ:x5K�,պy��X0"O� �m��(``9i���;y
��"OB�:S��������L�yz�"O0����,��Q	��K�4D���!"O*M�SC.OQ���E��>J?�`�"O��Ȥ�SJ��S�_<�Д"O��H&E�6�-��G�H�b�1"O�D�%lC�>Ӗy*G�-)��Y�P"O��N�����hP3|��w"O�h�� AS�H��F� 9��|j�"O}�Y5�hq�S��Q�v�(S"O��q�f�7��h�$742�,p�"OԱVC��L.�B�G.!����"Ov]��ʀy����A�t��8�6"OP)��`P�r����.ޖO�P��"O���t�Œ&�r=���B2oߺ\B�"O�A2��
u�.`�ϖD#*(�v"O��*�f�Y&�9P�R�W:�q��"Ov\CR���׶�aR���?�PQ�B"O����#lvD�T�Tqkl X�"Oj5f�'=���������`P�"O\Ғ�ҸjH��:��w~��"O�(�$'�;i�E�@�D9Xh�8�"O�T
jV�^�P���J��U"O�r�B� ��ك.S_��T�F"O<p�$�$��sC��P�.I'"OJ%�!���K�B7D�l�I�"OqQ�`Ə)?R	*�n��X�"O��G�!kN�rd
1'��)@g"O&0����ay慚eB �L����E"O�Q���+��ɹ�!�#ug��$"OĘ���3(H ]�@�M��"O��+�A֓6���;#�]$Y�f���"O��A�6`E{7���t�p"Of�F�^�W�����H[(7̼�d"O�t� d��v�"�t���"OT�3�Ҍi�����0 �E�2"Oj3sc��o���+�Mҳx
B�R�"Otr��
-[�b ����7"Z�pq"Oİ���A/!�r ���+�Q�"O�I�M��pe�Ή0d:��"O�f�R0�6Aaf�D,_n�q�"O� Ā�c���fvl�(�CCU8)z�"O�`���810d�9��O�D!ۂ"O& uC��y����B�U�@P"O��H�k�
H�d����j@J�i"O 	��O��C���Z�/�u ��xd"Od�P�M$~Vl���/��"��)u"O���m�+E�Ei���<`�ܐ0"O�]����0f�,�����s����"O���TKKp�)�J�"��MCf"O��Wd�l�,�QaJP/:�"i��"Oҩ�C��qr���Wi�4r{�Y�6"O�Y��.�;
�EP$ɓ6i�@+D"O ��S-G�:�zG�ɽb U)0"O����P�V��aT�פT^8��B"O�آ�`�.c�f�{R�B�|Y�XU"OD�!��9�M8W�3I�M�C"O*�@Q%��=jPK�UٜT9�"On�(!`X8����:�D��G"O�`*�CUT��ToAI�؋�"O:�Cb��r5�h��D�!�L�I�"OJ���E�*-�D�2ƅ�i50�E"O�� U�^�=�hh��HXI12"O�����8�P��T��W���1"O9��@ل9�4T0�͔):ݠT�"O��H��őd�V\��Z������"Or���]3�;�H+<�8���"O��J��ٽE���;P�M�1��蘷"O�܊#��M�ꀙ��O���9s�"O-�rƚ$zhP}Cd/�S�T�P�"On=�DBJ1O�4	J&�ۑWt���f"O��c�%�'OL!	Pj,�����"O����Z�u���$����V��y�'�C�RG�
9�D"����y�'��xi���N1$X���Q�=�y��I't�$��ND�f����é�y�D�:���	���'�p�1�I�-�y���Q��4�$)��J �yR�ָa�d��#� y�0�$���yB�U;6О)
Pa���2����y]
@Hҙ��&@3������yB��%x�H������1e��V�M��y"ĝ1R:�� �� �[K^���c�3�y���o F��я��Tʐ�vL��yr�63F��-^�N�@�b!��y�+ϔS:���b �Qy&��.X��y�/�4�0ԑ����C�ܝ�`
�,�yb�]�Lл��=d� �k�FՒ�yRJ{���p�h���� �Q�'�@�f���<_�ي�� {���'6��ZFgD�*�d�[�*ׄF���'�X��$��2S�b a��a�ƈ2�' &�rge�Kξ%����6Y����'-P��Ӈf�� �х7�T��'�A���c�5�!n�GǸ���'�P��%���!��Íii
���'V*h���[;��3`�Ab>U�'h��D!�71��qpwnǑpy P��'�	"CZ�tw��_Jf�
�'꼽�q#���1�a��V��0H)O���?�����J�$�Љ�%��!��O����ޑib���U��<6�!�$�{�Tۂ��
&M|�b��#0�!��q���%��>�ږ$�<�!�J&�cBA4@�zc�4/��p��� ��̇	D��C����"O
�4/��+�x����=R<��wX���Ij��ქ�:�bAh�b��v����wh�<���0>�b�ύ2����^^FQ�Aq�<ٰ��?b��D�p�N�v�fԺ��m�<	�h��~�0-�Q�<a�P
�l�Q�<Y3⋉Ôh(�JĹf5� ��Uy��'�H�����U�-��cYQ�)�	�'@4���W	��*�'��,�x[I>���6��51�"��'E �� ���-Y���0?Y!�^� ����J�9�p%ٔ�C�<1�c�!2��M[�N��
��$i�C�ɟYZ�I��Z�X��Xg���a1�C��ٲxy��^�dT�e��GߍT�B��0?����M-tCg��#"XDu{��	Hx����m�Qa��W菼bѼJ6�����!��9���0 -`� R�j����jd���R�ؔUZ��E�m��e�ȓz�(
F*�)��q7b٘McHX��gh�$2ScՌ�D���E�YN�H��P�I��ޚUtU��f�X�ȓm���ХD����6�M&O���Iq̓`����ᯒ�,8y "�
�&�@Y����i�HU<%(H(f�d��l�ȓ�
�Y�HS<oAX1� .G����Cn�\���]2&s�0��X�Cv̈́��r�S��d$�`�& ]���[�r�bK�j�*t����1Q����<�6DT�8�`�DK�7ʸ�ȓ5�,��"J�D
�]��ISOu�Ņ�=�~�@Po	��ܘ
��ҿ,ި��_x),j�2�̋�쎵��\V�<�F@�s����c2��EQ�<��G95�j ��Sq�;���A�<���KV�ԕb4��[��s�<	cĨD�IV��$�ԙ�r�<Q���(;,T	Fˆ�.��!�G@i�<�b$W=nV�#��M8)F
E\�<�FͅG����N��E�FBc�<ѠeI�i��`+l͛YWR<�$LV�<t��,b��s`h�T����T��k�<ID&�'S��A8bgã7(��$��d�<a�oוD�`��ω�H���#C_H�<�P���2�ab�̕uFh���TT�'rџT�A�"$Q��#-͌
͊ѹ�!@V�<���;eP����:dqւ�R�<�q�
�C���K���f�x�A0��Z�<ɔ*� ���2r �\�yi�Y�<����AM��x1�؈Cψ�;s��E�<Y�A��|�i�:��@\X�<��(@�e٦�1�+˔���[lh<i�i�)6z-���G�&=pD].�?��'���8�bUqT�pc%H8�aI�'�<�ٕ��I�U�BN� ��q0	�'�
GS$n�p�Xr�J�"D)�'�N��A��_��#�A���T8
�'��U��CR&7?x�)��Q*�)On�=E���&5y��h�{�pU����y�ꞈ}m(H��dT�l��C#�9�yr�I�o��ڕ��$`�NݙR��(�y2d��^��x���T�A�J�	�����y҈׋^ffђ��:9D�3֌��yRC�(/�R"4��R�Ce�G��y�L0�� A�>Jl�m���y
� ���*C�D0�)��pm��u"Om�)ϙ�$MAF���SYxI�$"O��36�S�gf8���e�2}��"O�	ya�!a}�aj��n��h(@"O$���!K�	JR �D��9�"O���� ���`�&�I��"OT@� +�SOQ� �e�z=���Ih>�I�|��S�S�/�>,�.:D���Џ��X=`��HV74:,Kc�9D���C��2"=�0�R-B	:����,D���v�X�fE{vIQ�Ez���b%D�|�2Ƌ�O�~e[1@ě�Dyd &D��kEB�%%�ɢ��C�J�����y®DsC�ȉ!�1l��@Tl٭��'�ў�O�T�;����*���!p���nn�
�'�.@��P2����WlE%a�zT�I>���0=��fR3A,QB����5����p�<��M��.E��{6�G�C/�����s�<	q'C�W7`A9�ʉ�J~ޤ��O�v�<�5��mr�I��ӹd��5��@�M�<)M�/>2��p�'�%��L���	L�<y�>��B2�&F��B�o\\��̓lB2wo d��}C��(uO��%���I6��}q1D�P),�`�Ò�uW�B�l#Zxn�3�՛㭌�W}HB�I�.>tX�u��,����^{6^C�I'~`�PS��Lt�Q��>;�C�I%tM�y�&�I
Ӥ=#�`��C:B�ɛxh��C�Èp_��q�YvV�C�ɦD7��y�`��I��nv�4�'a~B#�9 ���-P��P�{#F�1�ycS>Y�X�6J$�V��nP��y�EP<Bi�$�2D���Ѐ��\b�C��kt�lr'l�&��:3�	x8�C�	-	�BH�%oV9P���i�+�~�TC�XL��ԨO�y�~qH��^�W1C�	�\x�!hU4V�aU���^<�B�I_Cb) ���#�F5�-^l��B�	�h�b�;���+l>2���\^��C�ɏU�r�aᚆ^�\���-Z�C�	�
.���t�\!	,�yS!v��C�	�rM��y3�ƙ�0���'ޫDF���O<�>u�A�#څmG �x���?�B��ȓZJ����Q�c@������q�܇ȓ,�*!x�H��4Ȃ��)�EK<D���3O̟�XY�@�(X�ٳ�8D�4���є?��l1E%�r�D�"�7D�dT.�  �Z�B���-!���i��6D�l�#H�_�80�)I03�Z1 $�7|ONb���ǝ���@p@�'�X�3%)D�d��ǔ'Y�"d�uJ�	2t:��(D���̞�p �K�E�'=� t:��#D���6ğեD]�jqv�Y��/�!��ƶZ=�z��ǒ+S�P�! +H�!���B��Y���q��=�c.�;8�����ꅞ$N��S�ލ�`�-D�|Ӧ]�c\E1�^=EY��� ,D��e�A`��Cq��_��$j'&5D��s��!h@����)\�=qΠ��=D�pb��ݔt��L��pc �;D�ԊS�Q;����2B�d\L庳�5D��1f�M(v
9j�i}���m7D�$ɓ��7P���iu#�$��2D���B� lD>pI�.��!���0D�� ��2�c޻U:�I��P8`.Ԃ"O��$�A�d[���U�^�&"O@�� 7�Rx	�۟R��I��"OpL����Vܴ�8�@�^��k�"O���+�i�`�P�ͬ���"OvԃH�c�6��̘v�vDf"O`�rc�V;��ā���tU���"O����C�v��yp ��'na:�;E"O��a�Q5���Y�#_֩2�"O���c 2;!$�͖CE��b3"O^U#6��u�N�˰��uC���'"O.�+PoJ��b�6��!���"OHc�
X���딊ֿtj��"O�4{�nY�n��T���� hBZ���"O*��aK]R�<t�p�	,N��pD"Oz�)"��r�r��E��V��Y+%"Oꤋc!�1C���儹����"Ox,Hc떅[��-���^K�Y��"O"ZÎ¨\hL�2�$E�f\� G"O���d��]|�y
w&I#vm��@"O�%�a(ξH�I���y�S�\����~$�t��3�ik�+F�8B�	$��e�Ĵ?� �b��=8�&B䉗��UYF�.)	��I�� |ZC�I(\	"-���ۮn\��琷vJC䉬y`�@Ӭ���d<)cD�	S��B�I�sV�P�����Pj���B�Ig��C����Z1Ie$_�t��'eџ8�<�6L�
<� "��6�싒D�N�<����m����[�$#d��k�v�<�f��: Xp��2/��A��*t�<����jz�q�@��-8o$@S�v�<a�G!����,�T��n�p�<�p#A??T`�Ǫ@�`IS'o�oh<����`z��U�@A�q`�(�?�ϓߘ'�:1�.кRQ�TA��
_"T���'�����"�^�h7&�ak�,��'��Km�7k�Ld���)i�j
�'(0#�)Τ T0���;u|z�h
�'$T9��c�i��5�G����h�	�'/�@D��eR�'*����K�'�����Ն>�6�QG�	�4��		�'����r��?\V�t!g�A2|����'q��AW�)�24�6�ҳe!�Ǳ�U�I�u0�X��G��|L!���*R>�����	4���UG|O!�Đ$ٔY�iU�Z��,��gƠ2!��3j0��G���\0�TrD�
$gN!���{L���}��A9�)C�[����;�g?!�@p�ЂD�I���#�ry"�'| p{Tҙ"p\��ڔ;�L��'Q��E&��6�>�ص$(/�.D�r��N�a��Բ�"�.� ��N0D�d��E־mt���q�ǹ4R|���M<D��'5t�k��?pU>�҅A'D�L�A]��̽�#�D�W@N<�vK ړ�0<��)&}�Y(�lE�@��@�G�<�����X���s��FO�H@��<����>�x0)��� �
̃G�}�<��5U t����8�TX{��^A�<!��5T����E���@�C�<���ϪIR��ߌP,��q�B�<!bJ��X=f�2f�1Y_"�2'i�U�<��ύ2<D�2��Ѱ<e����WG�<� �Q���N�
�5�5��S� ��C"O)Yǭђ7��)q�iȒa�p��"O^	�E�!>���)�;Pzc�"O�U��f��%Ub�� �B4H<��*#"Oh(��4)_`��/O3�A��"O&Yb�g�Nl\�慜k*=�"O��`ҀںWۈ��׮տ!�F����&LO�T�"�Hn�
��i(JQ�"OBi!�,[�`�@�"ѡZ�z902"O��1Cf�yB���F d ̭�s"O>,Q��.F!��O�s�,z�"Ob��s����`$.\�ʾ���"O��x
��V�2m�7�Pe��'$�UMXX�+�>\)T��T�~!�D�"p@W�ށ�M��ᅰ4d!򤛫�\ڰ�	4�`��L5!�$[4�(u��
L=p�*�����9x1!�d%9$����5a�� ��*
1!����0%�:C��h���!�!�	Y�x%yU���w�T�)Ь @�}���l×K�C��D�QA�%
��i�$D��{'jV
)��G��7u�n�8�� D��#FX�$��}�"'ĉ`���	6` D��;7@�9XF|�H'Ė���%�`�=�O�˓Y`��'�]3W!���d� b�����'���3f�ۨZ��� o���꬀�'��,��	(
�8hqu���\J\R
�'�x��� _lG͸L����y�h�?�Z�yCO�G\Bp�����yr)��}򾐫�H�BO��&%���y��Z��˄�E�0ۆ��k���?9��
#`��E�Ʃ'�"\�G�%#;j�H�'b^${�L��E{$��K��Y�Ř'U���3Z�~�T!������'��;�M��0w ��+ئo��p�',D!А�N�0m���B�j����
�'*N0��
� 2�E����hR�'W�$*EP7��E�C�hW^��'�$f/X�j�$Ż6�)[�85Y�'n`X�fI�H�>�����Z��	�'m@=:tmو'Eb�$�8TO8�
�'�����%K���ҡ�C�G���9
�'U�Kf/֑v����gaȲB�P�
�'�B�z�m#0� �WD�'��M;�'j��i$
Z�*��H���	 �⵫�'0D�@ �݄r����i��@F�H���)����+Z�0���G�X��Ä۔�y��/>���s؃�~�)�)���y�-
��RD#�ʇ�j��ˀ �yBk��*���咾�(��F��y���>f�����#�O�������y��N8%x���M��w[^�j��9�y�'Ŝ&�p�
6t��U%n�������2���Д��#^ `�\���8[�"O`���!��kRm��x�P!HT"ON��@$�����LS)u�t �"O���E ��_�9S1.��@U�p9"O�݁gꀰp�DM �lб1�2 �F"Oެ
2`#a�9�+O(�� ��"O���@j��	��R"O�a;E*��cMd�I2	�%��a�"O�Y���H9<6XY�R�ם*z�w"Ol[CCF�WIj�������&M�"O칲"�<#ɀ1���e��%�"O� ���w�ɜC6 �����8?f��P�"O��K���0_?8L[�$H�z�EhD"O>�:�O-4\����%f���S"O�X2p���0�\��bZ*{�hyڅ"O
���E\��Fyj�c�?l.8j�	@�O���d\��+	�j(`��I%�y��Z�P ����u�`��$Y4�y�K� �L���"�0n�6̀2�F��y�aVQ��b�Č �q�X��=q�yBȐ�9k�4+%k݋*����kY��yZU��\��E��j:�=KP���'Q�C�	,v�bD��.�by���B���C��/,5�G��&sth�E��IyC�IE[(m��)ܾY/���� �e��B�Iml���LD�#�|)�d��<&C�!�"%z�	XaN(����3�B�I+]~�0p%菇C1����I�R�B�	+L�����+��YH�̌�S��C�I�ZlJqp���ش�ٷ�	�)��C�	�)=:e@��:�B���
��C�{���b�>�L��	�LB�ɆR���=x]�c���"�B�	�
7z�[�/F�\�Z��#�� B�	�iB��AM��wώ�u  #s�C䉅o��0!�Fڢ�!��߭���=!�'1�D�C�Ȧ^'�(��L�5ʹ���	0��E^`��&��+���ȓRL����A"Ylqu*�?kl��[b���k^��0���"�옅ȓ3U~A�3�۷��![�]x0�ȓ�hi���ּ_�9�ϫ\��̈́�EB P� O�z�ș�C��X�Nl�ȓ_����U��3:x����^R�I��@�"�u��;�ð䚢�f���~=4�Ĩ���z"N�NךT��`���l&�2(� �ΓK`@�ȓ3��8 s#��	�8XN�4k��l��	p~��Ս:�jq"#ҙ1�b�E(]!�y��o�N)��$���a�Ug���yr�^3k�B$��J�gW�mR�'���y�#0�0�ŏ� ]�^d��㉿�y��t��� �3]�^L�&k���y�ٳc�����i*Z|j��­�y���oh�Q�+PT  b�(��>��OXX3􁆏6њ$�r�ĳ6�H�[�"O ���֠ �X�
K�78z\ٗ"O
��s�� Ea�X'�џr=y��"O �f@�a��Cb�K�� "Od�`��7NM�� F�*G�8�"O��W;0Fճd ڂ]7n��"O,\��'S,�M*w�M���5Q!"Of\���(�|��FΟ$X��uy4"O�M)U,��Np����Q=l���+�"Oh�Y�NH>Ed�R�%(A�αʅ"O ڗ` #D�����G�8�k�"O(m�W�X�,�I�)(��i3�"O\y����Y���a"�.)v��S3"O:Ē�J�k[�U�TBK�@ź<h"O�5y���'�`��sO�� "O0=S�Kܣ{4*<��@َ~n�E��"O:tx�j��|uR���d��}��"O�}+6�#=*$C�eX�B�N�xg"O��8���h�-P珴"�00��"O4Ĉ�</���U�3�H��u"O� �p�6j�v!d��E�6@��"O�P�b�A�=+�B��@-j&_���'�ў�O�8ؓm��P��2.ѡDs�'� "�.�"q6�[��Z+!��D�	�'������� �, ���<b!6��',��1B'L4t�,�d�]�(8+���xr�A&;�΄cB��P�.��v��?�y�P�X6J`����t�,�#�5�y��P4T�){�/8il�X;Q�,�yR#W�]��D��Z�fIT����$�y��-aI�떍�p9�%��yBϟ|�\����O0L4xY�-L��'�ў�O��9�a�t|�m��+F���*�'ɂ��q��$��	�n�&m��dK
�'8������1��x��Jg�|p���"�B�*A���U����s�KǪ$(z���&p��Se�9x�(��ܝQ�P�ȓu����-!d�!��⃖?�B̅�I��(b� r A�#ώd��u�ȓ�鋀(�+�R=Yc�X��h%��3��\id
.i��`2�� (�t���	mEb�m��T]��05O�� Q,��	|�'��H�K:^�$R���!�
�'���X�g-]�h1��-N��<�Z
�'��yh&苙R�<��/�� �@Q
�'$l����K̹�3b�1q���
�'ND�[r�S�!R�=HSdL1gL�J�'�PD�a[!���Ҋ��R�Q�'�6щEK]�|��Ro۪ �Y��'`*����C�"`6����AsD�����D.�Sܧ/���$�G�Vk�1#B��8p4d��b�V����̘�l��H�K�2)��%�z5�T���gEƍ�$i�5�R5�ȓ���鶄@/��Q��䞵1�����H�B�v]1��Eyg��e�l�ȓ!Z�pV� �o��E�Qd��L��,G{�_��G�Db�9$��py�A��`4b	����?����0?� d7n�$\	�K�3 ���k�Αg�<�'�i�:Tj2A7 ���SGF`�<��c�3v��5x4���AA�=�"�A�<	Ō��5/�5;@ �p9��B�+�r�<�VN��!#�!���i�8�E q�<�^�c�!����p��`�2�rx�Fx�퍓#v�œ��;t�Ys�h�/�hO���D�>Iti�,	U�4ա3I1Li!�D�Oqf��� �4OkB\��Ĭ<�!�DlBh��ç���"}�a�L	!H!�$�'5ops��ĸ?�(m��ȷH�!�d�7TCTi;�Hֹ<�� ��b�!�����ÁTEFH���ƷU��{����V��`�
�!K;�<p��R�t�!��Q�H�ZE�*3-�(��#`!�$�3_�:��W H�%U5��Җ"O܀��m��-�=yt*����踶"O���,+�ܘ�s/��!�"��"Oƙ���ˤiQ1�J�<�Xf"Oڝ�T!8h�,P� E�N�|�ہ"O<@�J<>j|����k�p���"O �e�pS�i7jծf�614"O��� ��
�RxH�Ϯ=�Y��"O�(D�c&�����&,��c�"O���%�4��YԉS��.	��"On�+�MV6�̜���O)q�b�X0"O�X3�f�rTF�1J�s�h��"O� ���ܨ
�f)��{�P���|��)�S�
��:�C��0q�ΙB�C�1k�ܽ��Sp-pI�*M�\�C�I�M(���D�sH���>�B�	�c�$-�U�]�Tm����E
�
^^B�ɜ�P���cN8Pl��qI,��B�	
p6Vhc��D�s��t���B�c�1���
�_V\ Ql��cަB䉣V*X(�"/1RP��mѼ"�B䉯;��Id��zIJ�c��S)pp��D9?q��W�Y�9
 j�*g�!#�K�<QU*h�"٩
̤C1�F�<ٖ���2�R� �ϥXL�|"�$�A�<��F�g�x���Ǩ����d�@�<ل)�\��ACb���~!��������h�S�O��q5`\=Zj8��qDSj�j1[�"OZY���W�6.����صA�>�X �'�ў"~�aɹ)��!��E�!���{�+��y�ͬ~�dq��g�*y��6�y�m��^j\������J�`��Ĩ�y2�Adr�*#�?�hQ��
�y�$�YX-P7/��n�V���.�hO6�Ot��?Q��@�z0�j�@Wdӎ�6�^���x"nU3d He�N %���Λ�����?�	�HΓ+`�Yk��
��	"�+��nz`������w���
�D��aG3�؁��O�d��DȾ7c��i��8�Td�ȓ\ڀ�$�T�ᡩI�cU��t����5Tِ�������=�Ɠ2�0 ӣ��z��0;RA�!T|��'bt�R��� ���H���]>Ș��d#LO,�hՋO���JU�X28�v0�"OBD�6Czb�*��B$U�ҭie"O��!ъ]�<vx{�OC"kݢĸp"Of5��k��?�ͫ�Ol�BȀ "O���"�].1��A[��M9&(
�'��$��>���y���{l���߰�!�d^)h�h!R%CJ;����lR�f��O���D� Xxk��� F�@�C�Ժ1�!�D,I)�FM�<U� �Ir� �!�A?� �����j=�!Z �!��" ��x`�%u��Q��5Gz!�D�tX�r3��VY�-��OQ�Ti!򤇽k(L�#�E?YZ���\K!�A�\�Q�T��s���؃88!��x����E�R��-���f!�D�&��|�T�.��e� C�M!�d�]��ԡʁ�T�$�а�;�!�d��R|P���\�H0[!&�!�Ĝ+P�t�3A�#rx��â�\�B�!�$�}��$K�p�R@�ٞ��{"��y��'᝼v(����h�9Y�!��Z�|Zs�׋H�����@$=�!��5M�x�+ ��\��9UO� �!�3
�VA��/V�n�H���<�!��N;����2MFx������P,i!�d_��Е�'��2�h08�.��K!��7H6L���R�h��G/B�}"���"2�2�4X��F�|����#D�ԫ2��]��`k�:"3�bq� D���G�%l/���u��7��q
pD9D�,�u�����E�?Bz� �7D�hcE�
s��țA��o�Qj��8D�P�G��9|�%G�_/q�|��5D�� %1�C�?^�����0�a�"O�M $&�O��p�@D�,y� )X�"O8�8Vɏ�K�<L��Ʋ��,"O���w�X
>�t�`����CV"Ot(�a]�8�v�;ÀW�x���3�"O̴�����>x��;�c"O�Q"VFĢ�d	C �s4��z�"O��S���U;��@�J��<��'1Oz�:��μq�mĄ߷��t��"O ��g��I�L՚#հf�"�zv"O���P%T����ş/u���p"O���4��/+�d '.%N�~L�Q"O\MmT�'L}����1�J"O��+�r��a����!)��e"O�<��EE�|�^�j��έ(j��Af�')�	�%܂!��tl 9�� ��a��C�I��d �`)�u�!h4�>i~C�ɨ\ء�3� X�i Wv�C�I�0�4<�Ό�Y��TC�	 NY�C�	�d��S (���i�8nB�ɘS͢���J�81���(VC�	2RHHXG%ܞFY(�I֠Z
c�����O��ɱH$�Ek�Ǒ�"�`xH�N3|���<A�O�=���Sg�d��d� PH�W"O��z�	�NzJx�GJ5]7VT#�"O�e9�;!x�Q�f(˦�&,�V"O��2��ЃXp�Pe�D�ish$��"O�\ȡ�	�r4aE�ٙ$|�P(�"Od��6�-b.�p)�/�2�H� 5�'O���$�t���k�
�Y3����'ga~��p{2C<fC��2��(, �A+O���� <Jd&�Z�l�1/�� [��?EM!򤈑J/>4�f�.h�P��c�  +!�Ү����f�.hY�1��Bk!�E�4��D�YL��2�$NFR!�3�L����R �����*^<ў�E����>�2���uҸ8j$.,%B�'�a~l��}��#���xJ�У�OR��?����0?���.6a��ƞL�}����<Q7C,7���\�$�na����<y"i͇\Z2X�FG5F@�a�&�g�<���[�g�MX�n�8�H "�_h<�� w��7�C&�)�WmV���Ov��6�'ި-MA�Dc!�8h��`���O����/?�c��8O�qS7 9E8��Q@�����s��${��
��4��49x�@��p���`�7M�p�ꕀL�o��X�ȓ?ݴU*�%*{5P�Z%a�?B�:%��H|��؅"U&Xd�9�N>I���ȓ!���z!�4e�U�d��!72���g�'��	uybk��;�N��/v�Z4�s��)�Py���3m�1��N:3yse���y��V;8��hpg��^.ɺ�L��y2��=T�l}�p#�1]D~�*�y�@Ԫ�D][�E�[R���%�y�l�8o�pB�
�'$�!P`�A��>��O��2���Pw`�*FD��y`�'1O�%
�i��-�q"�	�.�H���"O�٩�H�G7�<��< K楑#"O�Ii�#�0���8R��7D �[�"OY�3N��l:��q��i=�))"O��2&"~X��JG�A�^6�!�q"O�IH!��<7�xf�_9E�h���'�1O�KԣK3z����5hY '"O� l���Q��ƝZ!K�q��s��'(��O|6�����ˁ@�h*t�X�!�DE�)��!E�&؄��G:1�!�DC:w�񂗫Y�\�b��֍@�!�ē�h�#v�?m�,
b�	�!�<��� h��lR�+����R�!�	 �@��-h��/�+S�!�DV�<�l���ѝ+����& T�Q�!�D�.7@� )�!v�<3G��>�!��.N�={G�OA��Af�ɱe�!�d4���k�o��"&�)Y��V�!��R� ����x�K0�_4zw!�ӰN�г���/��&YD\!��ޗ,����D,*v��RAI!���y���� ��.�G��+�Մ�h���B����#�`؍l�  �"OP� ʰX��TP%�E�j41;#"OH�"��ڂ����qʕ g$t�F"O<E;iR��d� �&��fft��"O�ݻ7Ȝ�2)(A�ɣkJl�`"O*`��B˄[����4e�G�h�6"OfTK�e��*x$�j�F<!B�&"O�'O�sZ�A�'2�A"O�e#��Z�x�i*F�@$���0"O��`�D0}H��c�Ԕ�f"O�d�KD!Y��05�~��"OT�w��=
�؉(�e�$6��h�"Ox�鴌X
a��d�r$�I���Y"O"E���ހVOJ�7"R �@�"O�E�^�@TB#��6Y�1D"O�e��&�+�ء����kC�䠂"Oj�����|b��R	ÌW �k�"O�Rf����Es�U	q@����"Oa��G̗u%��
�ER%$H~h��"O̤Y��D+_�����L��y�p"O�u��yG����- ���;�"O~� �	%i▙�� �<_׮�� "O�P�î�1y��L��N,z�Q"O�X�6l�`��nS'�9��"Ov	r�
�
:M�ic��	xh&"O((�ǅѩpjd���@�0�
a�D"Ox�ð	�}�
-�A��0�ѣ�"O$�P�~I �����`��'"O�(�r�
�,����:G>�a�"O�)�G�,]��h*��_9(�
�"O+EW|j�13L9�,�P3�X�<�ǩ;H�>�H!�28D��7�VT�<i`ӿܜ!�mpږ8����h�<��g�T0�ɶ⛲C9�q`�f�<�ڞ7�@�H��2R�4<At��z�<1�"Ns,P�f�*@>�@��w�<a�n��;�A�Dڀu����$��s�<Ѷ��|3@�X֭?Nb^|��Zh�<�G��w����&�0�t�2��c�<�P��7e�` 8@��=<����Rc�<!�d��B���雂���p�`�<1���?���r�Q�<��'�[�<93�F�@I:��o�l!���W�<��JP����QR��%}\�xɞO�<��߶���(V� <$u� ��G�<!7�V x�4`�w��v�Fy`��^�<a�n�/4Z��;��R�����d�<I��O:��s�MD`�����`�<6F�JS���5쎆9ۜ]���U�<� T�׫�
]a�m+�ϐV-��"O�TP���o�uS��$-�R�"ON5veЕM�ѫ�%�,���6"O E)(͊9��	A�EX2��1"OX��	]2�����N�j��*@"O6��#�K0%�0�F�2����"O���DD� �ީ����8��1C�"O<�:�'
�����ꏅn�2��5"O���b�:*]8�8��:���A"O�q�fX�K��<�.ͳB	*�+�"O������>�����1'�!*�"O���f��hՐ 1�\4�= �"O������&� \#��ٕ~�ܥ�"ON�����6��@� k�u��JU"OhN�Ҵz��[�3��pԨX1o�!�d����<Rv�[�j/���A�%#l!�;�ҀS'��QK����"�G!��W��H�V	�O=�\R��/6!�D����PgLP��$ 0����M,!�dL(%>΁ل� 3%�4�!�/@&R+!�d�>�+�S�jH�/��h!�;p�j��ү]!_�j� %C!��ZJ��4�%��/\$3T�N�!�$� ����B*` >MK��!\!���9S2ԍY�)_	J渽Sb��'!T!�$��7��S�(��n�&�`e��@S!�d� ��I�I��~���c�n(3!򄊴@ iH���.�����j!�$E*,�|Iy�	�bFּ�T!�.~b!�x��CE�$@1��5f�}�!�D�9�j&�R*f ؀����$�!��Wc<\��ɖ~����ٝq!�´O����,co$1hNo!�d�77p�!�6Y�F�[6`�%Hi!��+����%v�	7 2.\!�D��c���b�N#+�\��N��2�!�D������'yNe��� 
�!�D ���B���Qt�H�A�C�!��B/I
6QZ�٘|_dĠ����'��aVIӉP Z�r��C�<]��'��ʔF�)�(�pș	/�ո
�'G2�g�<=K���@��(ʁ�	�'��̹��ڊN��y ��LV0�'
�� ��L�.���i�N	B��8K�'��h"��9s�T�����	Ii =��'�H��ѯH
�b�`�,�E?\0��'���C�+��mR`�M7@�I�	�'��Å�L	1�8�f ̰=�L�	�'II2�ƞ���J4<�l ��'��ݨ��%��MRv�,6���'O��B@�<
�:<�D�H�'�8-��'pl=���K�;��d����&X(|��'�X����C�
]�t���P�O��`�'�R���JW�G�}a��?�y�'b�u@s#�2-�X1�C�E���l��'���B��<�Ή8smَ9L H�'T���O�����y xl#�'�v=J�ۏP�qs��$o���	�'5�0 �b:w0��q��=k�&yb�'���¦�[M�,�C�3 ��
�'�鳳���Be��j�^�"�&,�
�'�&���?&��E���.h	�'�6�9p���мI��n�B���'����)osXu�ak��Ep��� 9
��͐Uj�:��8q�y8"O��B�gERH(�	@�h�>�"O4XR����D�Ȇ��1I�JE@s"O�)�� ^��uطGC+�<U��"O��`P�=^�8ܩQ`4�$��"O�hA��1
���' �"��H0%"O��� ɂv��]y���N����"OB�i7"���.|J�nP/|Д�r#"O��XafE�oi2]@��çmTL�2w"O�YXT���ڵ{���+d�p�"O��I�J�g<��ނR��IC�"O�T����1��`A�iK$E����"OT�h�DT�W�Z/����"O����S�1��ѡ�DV��rV"O��t͋1{��A�e�Vfu��"O��p&��-�B� 5/�	��B"O�2�G�6�vi�`�9Ztt"Oh%(�ł���m���ꤛ�"OfP6�4o{F���F�6�8�1"O�=a`�<���:p&��z9�U"O:� #���ݮ	k�D���d��"O4q��KK�C��e0��ѵ,5"P"O�A�$*;>���ݳxt���"O���1,ۃ��Yy�"�sh�б"OTT�D�L�D���+��ʧ"_��ʡ"O��%E�$�|e� ުxwY{�"O��9Ҁ֛:�8X��"U�0{c"OJQk�G�!x`��f	Vh@�d��"O|�:�kÑ<��Ty�j����x�"O2��$/�*G(����"{ʝq�"O�P �oU���԰R�߸2B���6"Of�����7A���ʱw:>ɠ�"O ;�fF>M�d{`a'gE�(��"Ox��a��%F�� K�VE�%��"O����k�6V�2l{����d�b�A"O����+B��\#����u��p�����6=O�c�"|z�N/�L�#�c>N	�hx5W�<�'鎱/Lx�Q@�1a �2���<��}R�'-�S�B�(�}�X�{R"��'a�h��D_��i2Ve�}jnВ�C͚&0�B���/���e�J<S��P�AAU��������>�Lǣo�X0�s�"t��BIDS�<a��}��M?N�&i�sF�H��I���O�0iA5�R4m꾘���K}Cx5��'�Π���
0(���Xc�/og�i0�{b�'�� 	�h���@p�۔Y��������Z�V���� �[5��׋E�O!򄗺5Uf���bOP4m����W/ў �ᓀ	&2-�G��1	�(��SKՙ2x8B䉿NP��eN�t�BlC�@��N���3�	�Pf x��)�(<�R��{RC�I?��Y("Ey��Z�!Sy�c���'��>�I,=4L�ŏ�-e������?A��B�Ru�fJ �I�Ν��C�I"Bܻ6�4�Z��T�P[�C�I!PV u)�030���E�2a5�C�	}�\�9��a�1�*�8<��B��j�"��ГC��x�A�Q>&�RC�	�D�T�3 ��Z��9�.�\b4C�ɿ	͸��d��+Sl�[�Z*V�B�I�,����(_�"(�$a׈��B�I2P$�!�,S�2�aP�f�7�B�	7�X��#�ȻJ"N9��aȔp�B䉯(4$l�Eǁ�Y?���D��k��B�)� hG��zN�DT5�"���"O ���(��ܽjF��+&����T"OFزQn�L|��@�(2���8�"O �Z�?<�R�k���*
���"O����1*���;2+5�%��"OШ���>]��I+���(H���U"O\Y�-�DX��zB���nP�f"O���t�U��%����=�t���y��M	-�h��K��x��e֊�y�/<x��q�-t�V��*��C�I8ahz�j�ȟ%� �`^?�)C�)��<I�i��_�`�7�?%�T�;��^k�<1�E�Ԇ��2C�d�u��Xi�<�u��٢񭜘08��*F}�<�a�XOl�}f/���Ab!c�Q�<���'+<T�f�_8��7 Hf�'jў�' �::p�G�=N�eR㍞�m�꤆�h�2���jD7yC(
�����b�ȓ-�E+��!m���(��݆ȓ�l�����TZ�y� �i���"���H�h�XWdI��I8����~yrb�u�P̐�lT�)�f�����y���2W�ҥ��@ʆ���S懔�y̑�+�HIc�M	p\P�3�y�@�$@�����/��f��,���y�JHQ(����!*Rب�����p>���5?�G�]�yR4R�H�B�b�gǏI�<a�͛YǪhch��e�ABp��{�'Nў�'7�FB�W	Y�بxk�*�:(�ȓzԤ%آ��/����L(X�t��'�Ii��~�\Ni:�QEi�3B@��D� ɨO�#��E�{ָ�""��{Rݱ`��`}BJ>�O$��A�^XVmc�eր'g�P�O��=�'��'��jMD�Ā咢�ÃCUj4��'0���(�*w�m���ڇ5�(0�O>�'c�d2��|�p,¸:�X���B����,A���x�<I� �=��|q@Ǟ�\0�ß(�?����O\��e/��-SrL9��K;����P�'=�O�[ƪ	-e��J�h�+��ȹq��ēM2��S��yB	�	�N���=����Q%�y���_�h�
�gΙE>�Ӆ�Ƅ�?ُ{��'��j�&VP	7C�Mݒ�zL<9���	Pc�'�&� �g\�Z�QP�	C<�N���'a�ݱ�C]�;AJhH���>��H<��'�1OJ�?�g��1�pD�&W+~A걋0c3D�Dzg��q��UJ�*�<F���2D�8�q������W�G�yu���/lOl�	�j*Pd��%�&��V�|�Z�Pse�,��O��d�<�t!��g��`�
c�P%��O���}�ٟąJEEI�%�|��5#�,oj\�x�"O|�*N�.!B��Άbg�k��i!qOl�)�I~nZ�b x3�iȈe���4�J���B�I�GY.��	�"y x�$c�s����ɟ��?E���Y  h�h�'�C�<��+��y� ��bi0Ix��ѐ_�3�l���'/�{��(y�>;�	Ơ��y2�'S.h8U�Ϊ�9��F �r�tm�c�8)w�	z�"}I�˙=h����V�+lO���E��5$�p��D��QT�%��s�"ڧTs��)2'ʸ`���ªS�G����;���ɷ�I�S��@���J9'����'�ў"|J�HU�1���A%$N�(djM��%Rr�<!����e�j=�b�L��:)kJZ�<Ad枆o䒐�F��	b��0�GS�<� B�a��	������H8�::�"Ob!k��Y ���[��1`���O:��֕a�	yW(��_��p�3�L�-la��'/1O�3�s�<�٢�}>|�ȄV�L�	J��~����!<Պu�� �T��2C��m L��;�p?��o\:>�%���HT(�Ta�*�b?�����'ᑞt���7u��e���F4v1~�jw .�O�I��O�!Hs�'�5�c�3�Bp���1�S��y�0��y&퐮j��bP˖��(O.y��%$�'�@�r@��Vg���bb�d�4�����J�gT�tu�8#L>@\�e��}�v1)"�Z�2sbH�m�M�±:�����E��)�2V-�y�>i�������Fy�:��;9B,�E厰�y�ݳ%����X�0f��פ�HO@��d];=H.�I Ԁ�t�7�R�!��L=��ϓ:$�n�X��X�hh!��W�&�PDceo�"c�ʙ��C-A9Q��D{*��y�U�~B����
1��(Ҥ 4��4�Oʵ:��D�^�Y�7L3?����'�p��H���	;@����g�<���!��}o�B�	�p��X-�g�Czx��Ȕ'ў< Doҝ\�P�Q�Onz�@� 	{�<a��� &5���/�+b�S�y}�|�<�g}�Q�0�مݧ{E$D�po���yb�DIn�"�&{�݂ �K���IZX�(�򆆕��0��V*�r@�*D����nV����&ΦL� ���*)D�|��cF�$����@��&j�i#��)D����5]f��ф�<rIPH(T4D���$E��J�@�����wz$��ׁ3D����nW�(u��Q �ԡ�UF�.}!�d�O�0���ͩ��L�A�T�(|�&(>4��1ׯV j�2�x���UA�	��'*LO�⟠J�GI4�QQ*�U�Z�3d�'D���UG�IE��UΏ+%����e'D���2�f�#��%1+���6�%D�01(R)k!�����Ą)ق�A��1D����J,E�n=K�쁐�>�xC�.D���΁�<��R�$UQg�-D����J·b頑X����y��.,D���p���r>%�գ�5�^��Wh+D�@��Y<(�y�*Rb�0��>D�xؐ�§|52hzG�G��@s1B1D��05#G$F���b�(Z�V�8;e�#D�p��F5k������ �z$��)=D��R�a�24���#��/SF
�"E:D��J��A�X���й(�����4D�x��kԵ���p��a�l�Bԧ&D��πw�@hY"�r60q¬&D�$� �	��<Փ�m[�N &��S
1D��{1���SQ��)C+�"h�u.-D�$���$OJڰ8S�@[�}���)D��ZT���(j�@ڒ���w tB�'D����	X;#��8�ơ�`��A�0�9D�J��M>P���i���A+�]�d�*D�T1�n$7���J�dP�{B��"N6D��H3D2rH��gM� ;�t�XR�2D�x�geZ��*9*%F�5�N�1�m1D��ڒ�ߚ!�l����v��X�/D��Rw#؍ ;z���'$قp��*.D���$-FD*A"�Dl��u�P�-D�����.L.��y��W=��A��J!D��Ӡ-x�AH!#�hd4�0f;D�� �@�bԐ=�b�.t�d��"Ox�C�ˤHZ�1A�_7���;c"O���A�Q5R[�T7
�$]hp�!�"O�M*6�ܰ7�|Y�gȎ%Sj=��"O�`	��)7v�{�ǫC�|""O��l_�
�h#GU%U�JѺE󤔦R�T�µ��F����/�
1}1O�p�d:��C�FW��-i1"O��bW4A�p ���)�"q+�"OΙb̂H��H�"FH1o_5Ha"O�`C"Mu�)��K=2)a�"Oܡ��W�- ���C�c&��ۧ"O���iK
zM��1/�u*��""O&����ݣR��Xpu)��p�Y�V"O��؀μ�)��ًh�=
C"On����;4j%�Fߍk����"O��y� @G:$��%1�Th��"O�0��R(sl)���E!g���R"O<�3�� t�@��7+J�3�� �"O:X��3C�,���L�]�,IQ�"O$�ɠڜP�@�X��/f�5� "O��X!n����Y��1���"O��2�o[�"��q�DnP9����"O�d�k_�}Hq-٬#�x G"OJ}���\j�]���	�i�2"O���&m�w�D��B�C�^,n��"O]B�2`��6��q��{�"O�a��"÷U҈D�B�ӿ6�$Yj�"O6=���`c�Y殃�XQ���"O�-9��{c���,&-�� �"O,32MZ>K �Ę��֢~��C"O�9@��J1��P�eʗ?��Q�"O.ͣ���>�x�ȔɃ��A�v"O��K�R�@��˥�S���CV"O:��(X�kaB�'�����"O�I�(�2Uh��x��ɫ<��@#���sJr⟒������^@[�л""G@J�� "O��	!h�����H[5�≮��͜��'l@h�𙟔��A<ua�Ya�dρp�h=�'$:D�0�S��_��q�!��8?x���d�3<�(y�u�'@b6�<�}���/Ehn���h��7}����N�,�re��1��y�6�I��yri[�6٢&ұ߀����͘'܎���JU�Ş.]�5`5�^=`�T�S���y�8,�ȓ(������[���IS?dS�d���*�2+B<#|�'!6(J&\$��l����p\<E��'W��B�G^)�H���	u$t�s�-���ΑL�ِ5��
�`�:��!o�|��6n:�	.]O������!^� 9㖃�̚B䉋1��x��ڳ=6�xkf�R1�l"<�q�U�fL�~�!�p��3Э�E:v���΂v�<���ۚq(��͠N�^ Ч�E�(X��I�B0�)��<�DˌY<ĵ�a/+/��ĄH@�<�2"|VT�aE\�.�ֹ����<�%�cV���A���p놭��`��c�b�.�a|⦘1�~y�+����/X'J[�呀Z����ȓgp�䘑��4U�p�aw��XEx�nГ(��E�Ą7lb��{����( �J�%��y�C��1����n�U�qa��-<��9sN8�)�矔頡[ 8���Z K�1i�8�Zr�(D��s4���^�`����?(7�{��)D��;!�F=Y�&<z M E��b� %D�X�!�֞T^2�{5CY3����%D����F��!�6X#ƅ��y��z2K=D�4�Diº+��y0�הLgR��1�&D�� ~%1��ܛn��jE�t����"O���K��LY�� �j�;P�N�t"O60"Ue_�.�;�ʛ9��%��"O<mR
�Gf����Ǧb��M�S"O$�)5�[����)'G�Z��:p"O�xu��7�a{�ɚ�[ܤ}��dG-o�:u�q�3�MR�R�
f�P��E.ez��ȓa��0���4:}FI9�o��)	�0�@F1���'R�I��x�3��y��y�L<t�X����.4�t#���7_J�Ȫ��L-#(�3Pm#�`���M�y�І�Irf���v�Ԋ\���g�Ym ���ԋ_���ǄXi$扣;Ԇ���T A���	$B䉱sO@pp3iU>A9��c�(S�H�>�O��[$�R�N�&0�D$��(&D�"y̧
��		ӈ��t�~�g�E97hЇȓk����@��d49CK�:��9����|)
ܕ'��k��,=�⽤��������#��_�|��Pȋ'Z~�ԚwO`�`'�T�|@C6��%?��\��Ft�ZuA.F�f���	'h7|�Ö*�	p2�=�����*�C`����l21�H.�yb�@���Db���,�D_	��ИF)(9t�����M�t��0hNk�(��^�_=���䗴L�"0��`@��J%�K�j��'A��zU!�i�r]��8O,!Fd��<��O��N��e �f¦JJ�XԩG�co4Ѓ4M:4�x3��m8����.O�OR`���ٶ!�J@Ȗ3O�\�d��OS�YsB�o<������d��<�~)Ae�07;�(Q���q�p(4"Oʽqč��	�����B���A�@��B�h�����SY��)�	�&ʹa������g�$	/l�10B�5'�5�uI�3 
!���Od֥�*�Ex08b���$Z�<���d�F�4G�!R��X�Ů O��2���|�43��D�*ЌA��'� 4A��L�y3LސT�|!���
pzq���k�
8"E�;��D�(�P��F��P�Jg���&E@�+"CS��u�a��7^���a2q��,P�ߑ@45����y�by˂�'��x �^r~��N<U��q��iX[Ќ؏1��#'X�2������1ɂ�X��t�>�vN�����+�BlR�L�yp��$y���;E�?�6/M��J��	a6X TlP�f��=آD�+Q��x� D��q�'��% �T4����GW=O��Cf�����'���Ot�0j��X�$i�.�w�a&���TI,`:ۜ��9��
,!φB��  4���Vᛋ��tl�07T$�5h�n��I�޴I؈�Rd�ǈa�!�Q͕5
�Z�����
+�v�Ku��0
�~b��#�p=ytl2��x�����^���ۇ�ʊ�F<�g��<u�����-�>|���P��DB�g�Q������,S�iÇR9���>��!���y��J/uf�'?a�jB���|�r��+h{c�ǒ1
"�P�6)��@�2���5Ux(��	��ˤ�R�V����D�\w*�5�r��eo����ɹMn&�@��,M<�gR�-�� ��UȞ2�F!��RH<I�`��J� ��5F��7N�5^RX:񍔎3NHs�푑}�DEÅ��$�N� �A�D��W�����
9B�$�Y��ΰ7ϔM:v�V���<����cj�!�$LL�N1�iq�̽C��ۓ�¥/a`xi�@�6= ��;O�?�*T�"���D�cM�A���X�B��-���C	�L�H�"̩f� ��I"Hh8�p�D�/̀Z��P�A��9�D��FؔO$��W�A#��(�E�r����h���-�<Rb�97h
x�'�Q9'�PByb��.;ݘ��3�Ϳw�����(8r^$��s��=�����9�V�s�':ؖ���L=t����Hպ�y'@��0�D�6x(��O@���''��K�O@�O���1[�	��0#�cVv����Ƃ��u� )��V7fYQ���d$�'�P�ȥ�-=mn��'�D�re%`�8 �b�74b���թTRqO����=)�U�p�
�'v����^>T�He��_۪}��n�<~���Ơ^��˓>����g�yH"?Yq���<&v�KtBއ&��X���æ�	0�E�r�J��p$�m��pbWuT��H<���A
Yi�K�E=bɖ����çi����\;gZ��+Ów0Q�d��<�C!H-t�(Z�◛{��xPAM_;������)t��wJ���̧��#��'qh4[�
Jl82DʴS
@,�R*	#Q?�x�dT����rdJ9r:p!*��ȇy(J�S��-A� ���W#P��l���>'�.E�Z��d{�Ř_�R���!J�=6����'��X!%C�!qx`�'��ٟx�%�Y&O��
'�Ԑ;��<aB&�5\��'ut59b��B�g�"l˖��SD�8� 	j�@�J���O"z��Q�I��1�L9�'mΘ9�F�M.%k:iZ#)�:N?���2E �k8��j��3�Ol5(g�E7O��A+�/�lj|�C�Op#V|�L>I�ߟ�m$��2x�FqC�O�4����O�k�.�iYP�[0"OV����$�: 
�"�	_z�3�'�@��� "-� 0喉3����π �L��n˾V`�t�U��Na�)�C"Oh�j@�"v�T$�*qiH����V�U�ްp�M:�3��	.�2�*��ӺJ�.I�e�S�>}qO��"�i����r9ȧI��Bޮ�X��(jU�S�H02�:��MJ�0?q����b�؆�^9Un��ià%�DHH>�$�a�Cķ.����`�>Q@��D����@��-V`�h�b�bh<�)�-9�c
e��)� G�3���rOYQ9� Y6	2 r��>iK#W�EW��1�T�2s&�8��*<O����ձ7{*�(�OlM��W��h9�%�����C"O5@����^9�D\�5#~<:��|b���0/fjԪ�C�OI�I�3�ͣS�-�gO�����'�TQ���Y�REr��A�
�hd9�ɔ�Yɚ�'.͘���>��
E
����:����e�ah<Y�K�S�J]`D��	b��5�ći���YEnՇD���lڹg����1=Oʥ�(P���'���pRD_l�29��c	�:y����m�>�E#�9}�6m߹K��i�e� |�%9�
�[P��z�fO�4_46�O�&"\AP+*LO�h�&LA43�0�0ቀ�S2z��Q�|����P5t��dΖm�P#���2ǺB�p�Lπj.D�'�����,J,��B�I̂D����m ��@}~��l���#�@U�H
�X�h��9.�-٦J=���Π<:�>f��D�A)��,��Xem��n<!�$��9Kl�2U	#&�`�  ��,�5��d(T��Z��Vܲ)�!ك8Ih�"E�O�j�O��F�ۈc��q�ꐓ_ʮ1��'���نӖc�h�l�90� А K�&~�.]AF�'�ذcÉ��
�0��$П>L��F&O
�ہ�I2NFџ8q#$�:1TL P.G/%� )iTGOl4k�lT"���2���;��p	�'�>�3�[�c�ڄ�� �)]����(O��Z��Sq�x��Nc��c�a��\l�K�~��ѳc������"OZ����4R���ao1h1��ӱ�U:o��dC�	ܽ�f�fC>^�~2��&�����h��Uz�!]�J�"H8�K5�O&D��ՀOHTM��LI�+�����ٓHbH�����N̐лb�9,���D�ox��b�P����&[9.�6���D4�'��]��
Y�� ��i�2����T1+S
}*"mF=dQ���\)���x�g�gh<���Pf���E�;����b��ڳ�C.E��7g��(�R URb�~��zĄ����8��,�>FL�ȓb~������/�n��'���ӒY�Z+�(�"�G�N���]���U���=Y���ZȀx �.�"r�&�� I�kX�@�'a�Q$�݂p`ȦVqJ%���U�j���'�2E�B��46h L�� H:O�di���ݤ4&�"=!q��1>T)`�g�'!�pXx��A5A���� Z�w��؇�qx��ᦏ�k��aZ7J�3[tv��I(h�0�����w��S�O���� �wI�8�/�.�P��t"OpQ򠔾*] ���n�,��=Y�^�p�tΖ;2�t��'\��+@k�ސ�`��O�V2����RVP˂��l��a��J>�V�B'��-��'ʼTI&��klF��G�| ����˕e��x���I�wذ0�t@��(CA��t�!򄀤L�AZ�IX�>3	iզܾ)w!��R���cV3G�Yk�ݷk!�$�jU���7��
\��Bg�"+!�=P.}��Y*��i R���,!��4��8�ݽl#<(�q-��'!��G:1�=���Ȃo�Eku��6Z!���%Bv�hr&�+��̒GD���!�����X��A�fF#r�!�.x��MMU�d�"]��!��0:��*׋��>�V��#H� �!�ĉ�P�,k�7*m5�a�0�!��=��P��#_��ebQZ�!�ӕS�X8�1�i�1Igj�C�!�]e�� ���'<���oəcb!�dE�#�z�R r�(��|�!�$ۋT���6aӯ!���u ʖ�!�Ǔ �2Pi"%[�L`p��j��!��YX�40gڔE}(S�'��!�� �u�L�9�\������x��!"O��BS9 M�L��%U�.� 4 �"O��yu�(6��se�P�.��}�f"OD-��-şd�,%A�#f�<4"O���  Y[���S�ю�= A"OH��� +)�V��&���z��ȑ"O����+&T�P�3�3i�R���"O�@kT�M!Qu�� ���"�HhG"Oh���$[:o��#J�9o��"Orp ��Q�Ytv�Ĳj}�T�C"O���&@3nhKP��;W@a�"Ovih��ߧm�jh����J4Ӓ"Ois�ܺ&����l�,i�`��"Oz�&Ǌc&͈f�	��	�"O͡"�ݳ[[`�!biϪm��a"O�䣧�K�b�^��0�4��`E"O������G�!-Mp��"Oҕ��)�=*�][HFZ�'"O��q�M�셺�k
�~&a��"OČ��:�e�U�� ��lK�"O��z���	/~ �*C�Sd9b�"O��hvO\PUH�?/z �"O��j���4z}T��ƚ6/Xó"O~�[5FX�(�g倔��M��"OX�R/�0k3�x`#�e�T;�"O��������q��>d��%"O<�0�-�ꝁ�OZ/W�i��"O؈�3J���r�홺I���$"O�9�G],L�N�y��,$>���"OT�%�Wݰ :�eZ�\�&��V"O��w�Z�����FXX��!"O�9;�D�@;�|���UM�i��"O�����<~ ��#�;	F�d�"O���DM��8ˀ�c+"N�K�"O@T��Aq���2D�9$.��! "OҰ�V��=��YE��%,� ��"O�
���hQ
�BcȓS
���"O
��֡�3HG���B�@��^�"O&u�排
�8u�-�,��jG"O����	x���Z
�x�tC"O��"c��|��`\�U<�U���N1�y��E:b5��WD��p��<�y��S'����é@�j��l���y�kC�/-^�J�&�deV�M��y��׿`��e(ăٞY�^�3+��y�JS�R�P���F�a.���f��y�*Ư<�R�55,`�hb��y�*@���("�-�>w��l���yR�[:9��
>3G�(��藊�y�J�3Y�35H��]�v�����-�y"!7�0 ��EX�Q��	Ȑ`���y-�tQ��T!�/8 t�
���y�@*g�$d!�)�2>E�=�2@�9�y�+�;�P5A��,�$�+%!��yBa��gH�Y�d�/� }x���ygZ�$��Pi�3<�fh��b��yb+��{���9E�.7s�|H��B��y살-^2���'�6s;�0V�Y��y���?a��qs ʄ�$�Q�H]�yҭZ�Cܵ�3g�A�E���y"���0�h<C ��\-j�d́��yb�O�q���K�I�.&������y�*�L���r�C�2!C ��y҆�:4J���e�0x�~@���+�y
� �1�E[�@.����7r���"Oʨ��#'|�qQe�&b[����"O��b� ��D�CA��"O�q��Δ/�j�á#(Y>\` v"O` ০A�>�V=q���~�I��"OP��ЀJ/^����ਃ3UcP��"O6$��D�>��`��!ƹ\\���1"O<<� A �4%�Ic����)�1�
�'�Ѳ��$b-����B �x�<�	�'*F�&�Z�(���H��Ps�����{Bh�Id��A!�ӗQ����l�_��X�,]�ִB�5����6oW��x�ƚ��L+A���>��8 E��O�y3&@"rb�P����qs5O�qS)ΨF26�hC��w��iZ �X�5��RT�	4֚��D˙F�2ꇄx�(�q �]�e��yj�|�<�!��ܩg�󄝬P�Td���Y,"�0q���ÁT�!�9�,�g.��uԈ@�,��'��iBA�*�Č�1����H�w��&@�]#`�ۢJ;C䉳6U�`BsO F��##��ŉ�7�P�a�^,���L���H7َQ#�/ڞ+ú����-4�@���7`R�	ZgƄ3_��(�S@�{TLc�嘣paF0��	�1�� Gύ�lM.-�#j˒p�b�󄍑oE:��*ʐs�f�	�~�2+��~��H�Z4nB�I$��%AB�"y8�KF"E�j\�O:�c&=iR\���?�H�,��$D��.@`��
�+JՇ�5��L蒊��Mڰ}H��}�0(xcH��,���'�zqx���`���Z���b�b��ǜX!��_<]Jؘ�M̏Uz��$I��3���������,�B�j�:?���.��!�`B�I%M����-^*`jx�pg���FB�ɬM�(:�C�%[$�{�mY��HB�	!��[�j�s�z�B��V�L�pB�	.Px�|C`i�At��`�`4{�`C�/ ���C�.XPˀ��� �jC�I�\��T�N|�G���p�"C�I.S�虐tAA�)�5���:-8&C�I�.��&��/\�rcWdX,,C�������ׅe�H)�UΖ�R�"B��lF ȂJF�,�Qc�_�C�ɐCV�؇h�b�"\Uk;��B�	�������9U�l���)�4��B�ɓ���S&0F~PRdO,�C�I@��ӡ�[�?�>��Ѣ^�zdn�?Q�o���O�JtL� j�j�KS�H�xC��	�gųG�� ��'�@1�3n˦p���Mw��pR�O4��ϋ�4j��'�|"�ߗLl�OȒȹ� ��Zh�s�	�c�ޤc�'V�=����#SL`J��USzm`�^�zk�e*�ħfxAX%�wa�I���t��]�	��l�b�[��`%oϰF����72�jQ�ʞc� 1 тom~��V��>��QZ�B�F4��f_y2��4lW�Z���Z�'�LP{�a/��� �9)��JN�|��дq3^\��,Xi�*|8�D<�Ӳa!�:�I�9��ْ�D�m��P�������'�-`ѬX���tk``Q3g4J��a� Ǟ����� 1S���;�r�Lر��\S0`Q2��� g�˂��
�:H �
f �B�1�4	��M�_���QFKi������ث�J��n�$���.=n�ɪ�~��Rě�A�����ʥI؄w�|0��#�8CU���dקbƱ�al��}qg('G7�p�B�cм���N�yӜ@B�C���39��e#�����O�{�hK�H��� ����ĸ@��>IQ�"��An
?f�u`i�"��'/�%r�,ټ4`���Sb�6�h��Pɜ�c#�/�ORlzR�c}m���'	r>�h�c�% )�!{�g��x]dp�@璍C2���ax㟀3g"�9CV|x�݌^���
��&��#��6;?8���H�--�`��D*ָZ�}����x���.�h���ֹ[�X\��r��,��)����6ck����)�oIay-Ʒ6�j[�MRۖ`�I�s6��Y��S�FĮ�Y�o��{B��'C<}��_C��,�}&�xE���{Xh���6oH	� �8�$6mB�pk6R<�| #� �Pʰ�0_�y)�*�	,F��d,�
�j-(��'9�@�5a�i��U���pL`��CO�]"l$�d��O>T�O�ms
��' �b�c�.>Iv�����P�'�lj�bS�[=$��&"�)��6/2-��#� _f��������d�'B�,]� �\�6�0���ip$�C�ɐh���ƈ�����Iõ��-�fi+}��o2��}&�XC��	0��m�v��"؍�I<�	���`�4�S|�a��x1|$bg8[1��ya��%��Y��'� d¶�K�S�qHԔ�PU2��B'm��'�TE�� M��,��B���':�)����0N`%X�fܩ��']B1��;;�YP6���� �Q'�$4����er\���`Hp�S�'U��i�& Hɹŧ�=`c�$��$&X��e�<ba��&:p�{&��(2�`	c�L\�bB䉎D���S�<�N���o�.wo�OJ��d��-qe�X��i��2K�!q�!Ï4��c'_%_�!��M�+F�0c�뗟J�|�ڦ�5��t�ĉs���h8��?�'R�5�ϣb�~-�"�ҲDs�x�'�<��F��Ϝ�`1�FPp⒊ �\f!��,Y��M{�h�
O^P�!E��-������Yp!�C�nό�x��F�.��y"ÝjŘ�8� ��k�C /����,V�>mBu8'�K�(�2+������)� ԇ�I&u���tg�2$��`P���:�O �H0%�9�0mzPG��Nq84{b���Tؕ� O�'p�� q��\�t�TL�$��qA Mh<�� (������o�d��6��Yx��ڴ�|��B-��Q�&�; ��,3Zp9��[>m�@o`��Pb������oJ��2��@ D��@�kӇ�D1!S�`%Np;� �5�8ix �7r��9�b�e��H�+S��F�I�[��)I(�#�o�8$��2F牀�������C0�i��&[��8��Ò�x�f%�0Un}���M�72��� �Kx�����*x���/XZ�`�:��")R���J׾]E�hA!L�l)��b�׹':�cPG�Q�z�#a��lġ��D�������\��I���Y���yD`92$'�z�b���{dr �����˛"��)�jD�<�MJ��@��y2��Q�p�Ҩ�?c��"K�a��)1M�-'���Fجa�)1N?��G�"�$�dȐ�p��O5�T�ys�(�a~bA��Xr4k��ӸP+��׈D��#v̇�$\0��B�}�x��	N0`��y�O���$*�苵M�V��嫊�hO&�;G&�$3�@%�BMs����5�H�|��p(�EX1`�<�A2�#B����- ;��x��n���tOԼ1�����+�?��h��H�P�+3Ϯ�����J�F�i��f�� �N��1"4��m�����yr��gd�	��j�(-���`�*���yR&�k�l���lZ�u���?UCE#5�Ɋ@?�%�&o�>;�0�&"Z�G�L��dD�T�hT#%;x�Y�)_���1�F�j��A
�'�8�-�|"(���kT�\L�s������u�f��	��O3���(x�� ��Ւ`Ď4��'�bD� "��)���6�V%grlE���$>	�1"
�hwhӧ��&�9�Y4�0�Ň)n��m-D�Y�I�J���#��|NI��<�2��	I^��?,O�]8�Ú�*\�Aˊ�)��'u�HBL=��L��1�q  �G*/�,��O�є�I�#|�P�]x��ご)Q�����ɝ"}>9[`���N�RdӢ蜋hl���k>D��,܊�cV(V�<�I�(h�C�I*�¹� `I4|f�� ���,�C�5��t�WI�("��%� ��1ɄC�I1߰��C+�$����c닉a<�C�1m�&���+_�,,F�9��5�(C�I�-���2�_��BJ'��=p�ZB�	�N���FO�X�>�����B�7D�|��F߅w!@��p��7<�����8D����Yd�6�)�d^<�����4D�|���*Z���٤`\9x�B�k1D��'`U�a��r!�F�	E�@�D�%D��X��݈S�m��m�� 9�Z�f"D����ވ9"8h��	O�*�rc�,D���6�d��I�'�=�|�c�+D�� XM#G@Ө$�,��1	L�	��Z�"O{'�[?*%��H�(]�0��,�#"O�D�P��e^-���+f�RT؅"Or%��֮2�r�BV�O�Jfd�t"O�!:�� �,S���D�AB��y�"Ov�X�A؞H�r�,H =�R �""Oͣ�lM,Z��Z#�Ν3�<�g"ON���b�$v���z�!�;=b|"O���˂9����J�	E)>H�A"O���'"�a��(i��`�h1"O��ꓫ¬T�"��'h�:@��2q"O����>���+(�aN���"O��C�) �P�2S�g_=AX�+�"O�X��D]�!H�@�-ʨ%|��I��+"s��1��H�mG��`�buQ��yb��>�Jpq��-a�8Kc����y�F��A�N82r%�R�P4r�kގ�y�Οwqp�4ED���A���y�'��18��Z=�H�Q(�
�y�Q�}z4�Ra�S�_�j�1I�6�y���5i�z���cڠX�����yҍU4H#&��ˌ( ��U�]��y�풄Z������h�L�1�m[ �y��8#`���a1���s��3�yBe� �४e�ք[�� JӅ����m��(��Y���_�x]�4��5�J,/QȮ�Iҏˈ������T�=Z�+����?����tf[p�)~����,�^�Ue�M9$D!٘([2L�&�>�R(V21P�`�Vm&��bp!��I���ʔ�ݒ4Uf؁�P�H�F�&\씠�J>E�����[��QdD�)�n�q�Nʹ�?��/��5AD��J>E�tk��ӒoV=#9n0Y�b�)ڴ��ۂ�'�0LQp���A��;�!QF�i	�'�����E�]����1J�%N���3	�'���ip�J��z���ZEm�3	�'�,�F���i�z�H�q
}	�'B�KB ��(g�k5KK�={�D��'۪�SGbƻkd�8 �H:I`�;
�'S �lS&�nBċ�b��s��9�S��@
&5y@�¨&�`�$��y�b@=U�2��Q�	�4=lU�C�
�yǐ�'Զђ��0'�E�U��yf��}A�0Ag$/Sl=���S��yrA�4���Bc�M3>��ș"(��y�e*�*t0Q�O�B��l�����y2��xpAq��.7<�����ņ�y�R�4��h�E�@�A�g��ybD�j�$�pu+�2}�L!�B�^>�ybn�1(�x-�D/�	w�>M���yr
K�QxM�@,w�lpX �ݭ�y"�1�N����o���S2�y"�9�� �A�t��yr��%PL)�p�ͼZ����'�y�+�F<�X��%���,�;�L�%�y�Í+\T��e�	~0���@",�y��i5�ܒ��4{pV ��%�y�c�l���&��$:�AM��y"��+���`��n�n���&��y�-Y-uI �!��B�V��wcM��y�fV�xoz<�J�+a������y�(�F2Vpy&F�?Y�  ���W<�y�G�nh|M2�+ٳcW�i�1蟨�y��VF�*�ALT;L�X5�d	S)�y"���]��aj"̛IH[t�)�y"Kԝ5U��1C->X�`�;'�'�yB-�-7BJ�т��8T����F�Ï�y
� 11$#ȇ'V�	���P��6ነ"O�ʔ	�#0������ M�jغF"O�����V�(R�b�\��-��"OT��7Ǝ�kBLLG�(�t"O���t����@2��qz���E"OVLX�.�*3�N9�!���Hn�8`1"O���T	Y.z���!&O�=[�Q+R"O�K�aW�.�^"�@�$r�HF"O,SsmS�@Y9H�/؉9q�\(�"O�Yq`%�,M���*0)�Wm��"O𥰒��,r\�`�g�0if���"O�	c0��&z����D�NAZ���"O�m���ިn�Ѡ�ɪ%��X�"O�E�0��s�N��A)0s"OX�t+G�o��0�@Q�@)�q"O�x8��g��H�/�2*ڐ��s"O�9�C��70� Is~3^t�"O�a
�5{ Ф4���"�"O�l���/_�H᪀�d�|Q�"OTuj�A@HD�J�"��f�����"O����[�3)��B:����"O�Mk�f��_)`�0�/��2�`"O���6/�: ����*zp\�"O�A����,	"�Ćr`���'"O��@񢀽`��mG.�<D"O�����c4H���@�}�"O�u��$�)[��܁V��na�"O������,B�F��2��	�ŉW"O����(�75"�
���Q�`"OLQ�-F�s�d, �#�#Z�5�s"Od��G�H�_���ᜦuW*uS""O(Ţ�H�/Y�r��a@J�H�q"O@�E�0^�j8�C/�*.��"Ob=�sd�i`́BAS�sN���"O��%��gkXdC�/3V]�0�T"O!�⍍:�Nm�f�/|Q$)k�"O^PI΍:.|��!��S9W�썂"O�� Џ�\s%OH�h���#"O�]b�ث �Jm���ʎ+��L@�"O���ѡW H��Q���(%`1"Oh�.���|��4!�Q"O��CIK�x���XW�T����"O��!smOD�H�w�1
�2�X�"O�Q�剈�5�NI�P�G�{`Td9�"OTH����,J�у"�7N� A�V"Ovݣ�'�<Ԇ@�� K�&Mӄ"O"fĶK�|ՉCo�-1��T��"O�{���e3eNL�V�J�Z5"OX�	�a��qӈȉ���%s��V"O:��a��&SDfT�̈́�ec�� U"O�i[�]R��`�4�X�)����W"O��1��k�����DZ?a��ec�"OXԃ���F�d�xP#� �Q�"OL!��jT�4=xc���v�$��"OҔ�Q�����I�.�y��@�"O�m��jZ$���[*7�cS"O�=�%�#=u����oS��y�"O�$@��C�d�܅󔯎+r�^�ӄ"O�`�tɠ�	�f����3"O��KW��j�(B�.���HR"O��1jWW�}R/Y���A"O� ���p�̢
�i�
� �"O��&��Z3�81fͥW�Z��'"O2��2'U\.�#�уŨ<�"O� $X��$ D�T��C@��a� j�"O��it�T"X<ш@�	1>�f<��"O�"f�H�6�|����+Q���6"O�|k���x�~���$	2|Hz�"O4�� �P�Z���p"Ԩ`���"O��3��JU�*A��	o���"O�9G/�rr	t+�&djƥ��"Od����[�T\XUE(��(W~��w"OH��n�x��*8��:�"O����NT���&�F7�R"O�ݫP�������W�/�ȺW"OU㗉Ⱥq�=�`�;>x��"O�e@���"ͺB凖�f��"`"O��Q8���J�D�u�dD��"Or�{Ǡ#ɞ�`2�#(���""O@���/�b�P�,�`�r���"O^�Q׈�67����@4F��1�"O,����-P�ի�i	�zp����"O
л�(Y ݠK��FX�� "O�i�w�;Q��p	�H:��E"Od0��c�7���v�#<�lٖ"OZ��Ń-��$��G��Ji�EH�"OR����߹@�N=���<j��M{t"O���分)���Ja��2��5J�"OlYX��K��ҜA6c�$�*�i�"Oz�
�O�CM($�&T	�h�P"O��"��m�ШC@gЩWY��:�"O H�ˌ-9L�J�@�,P��C%"OL�;Cř��qH�b�8CL�);a"O��@v�>z�*�ң��702���"O�y�P�:2�f!zg�Hb�����"O�$BW�˶�̉���5�ʤ�u"O���B']z\䃵		uJnPr�"O�����Ҽ�rmH0�� +�;D"OT�c��ll2�[V��8r�a�"O�0:bo͔w�(��ݐZU !"OFu��-s<V��+[NU6ͲB"OV�Ġ�h��T�	�;���1"O!�p�$�����%3���"Oʘ���/��8���1#QI��"O��wЀ3�P�2�I)n���0"O�*�eD�W4�����5A22�j�"O�I����C5��C�߮7%����"O8Ls��.�"}��)C�?��u2"O�b �F�!8�rW�[)KB51�"Ox!�2H�)�|P���e74h!�"OPɘ� ϩJ4�$��(J<QtJ�"O�24���P�(1��ߖ~ Xa�"O�`a��� P��$�·�C~XF"OP���,�}42�u��6��"%"O,�qkǱ.(�"�e͝/Ң"O���a'��UP0�Zr�Ib^��"O��MS�V,BT�/X�L��"O�0r�_���jqÜ�5��=�&"O�V���Pe��Z+_�b�z2"O^�"���P��K�o��zـp"O���eC��PEb�Ha%ݽJ�b\�"O\5��I�v��b�Î�[]��y�"O���� I�6�扠���	p���"O(��Y3 h�C�FU�k��("Ory����'w�0:����a��"O�l��b1	z�ya"hJ�N�Be�"O��t��A�ȓ��D�Nq�"O�e�u#�\�-҅搊|[8%�"O� X�I�!f�#fO�֠¥"O@A3�d�#s��]��k��5��"O�0��.�lآ�r��")�.<�&"O��7�J�e��(���J�X��"O,�I3���=����w@�.��
e"O��UK�S�@�X�OG�v�90"O��˰Ɓ�%�:�O��i��= �"O��3B�W::��܋c@�7��J4"OD���@V�s[�Z�O !y٘�$�y2m5��D���qҭ���/�y©I
 w�v#�� ~�!�d�A�y���"K<M��{��	2���7�y��7;��8 Fa�v��I��B�y�a)E�Z9:�ˮ@���+!OQ��yb�ёqn��V��=Ij �p:�y���Lnq�bHH|��D�����yb��nb>H��"I�z[4̹��[�y�D�j��  u��&j������y򇜫����7��K��y�.ٌ�y�I�M�b��˓-D@�z����y"K�2:~��Z�b�6d0�+�I�yr�Y�r���K�ϔ]�R�H�^�y�FZ�6����ǴJ�^ tIT+�y���$eD☀7AѓGɌ$��K4�yrj�F�j�a�-B�����煵�yBD	*�F$c��<%�����y§��B�^z�d?S?mak���y�g�*N��ŠڗLhġ��D��yb)A�|E�[��5<u84�EC=�y�K �DRX��`B8ۀ��1��y��ibji�# �,:����ᗗ�y�Nj�U��@�!+�HP��Z��y2.̑�b���%ë1F���ż�y"�B�l/�\0R/֎R(`�ȀȐ�yr��?^��q%b�N��y��Ν�y�*�'&�h4"�ʰE�PX�a�#�y��"�R8�A1":uhfh�2�yi �	�bS�h.�F����y���"k�nE�"nç4<l�B��þ�y�N:sHS��҈4��t2�;�y����j�^� ��;3�}P��^��y2$+"j�m��Ɏ�/aD� ��U �y�G �JL:�*�+
�;�.�y�-�p @  ���?y��RP��l�@&,�%�a�����Ɵ��	43.b� �	����I�T�*,A�@ u!�tڀ�@)�v�S�4�?�D�Ě:����'w�S�(As`��?�Dq�5$C�Oy�(� �Y9�M���FV��<����?y�����@�C�F�#d�I�,��P�cJ�!K m�i�|��՟D�I�0�'V�' uSʇ�D>�<s1FF�!v���.ٳ��'[��'��؟p��KxrcD7������/�Je�*妩��՟��Im���?� G&{k�<oڌ5�t8��b���x�s$���듃?Q�����O -��|Z��J:�U��+E��+b>�b��Mכ&�'+�Of�D�'Cc�uוxb"��`���׻.6ͺ�'ڐ�Ms����D�Oj|�a�|2���?i�'u���&MP$��h�foR6w� �(����OpC��G�>�1O�3� � �e�n�2O��[|⡘$Q�,�I85`���I⟴�	�d��yZw���.��,���h������O��d՞��#����aR���WG�~�|HW�LԛFD�Y�2�'���'���]���Ɵ����۰g�P�iC� fNp��˙�Ms���D�V�<E���'��8�`λ'N�����g1� "%~�.���O��$A�i���|���?��'�.�W�"L��|�Wf�4H,� �-�I++z�E�N|����?y�'�-*"e_)I��;f��?N|���4�?i������O���O��0s���7T�P偕�x�Iۑ��>�YB���R�!?���?�/O0�䔫!L����R�Mw"���KܷlZ��Ф�<����?I����'hb x�|�8���(�U�GD�o(��%$�1��D�ON�D�<I�66Dys�O7h,	��m3(ڀ	���Y`���9�	����Ip���?1%�Ԯ8p�-o�� Cҝi����,�����?����O2�)!��|"�'xD��פB��1��)��sJ��
�4�?��'l~�P4o���K��TC�+ Sh�$"�J!8_�Xm�ӟĔ'WR�1@e��֟@�I�?ѩ�o�!� �I�O�6���D�S���'�"�@�zxx�y��J���/�̈!#���=n� �"V�|��8M��P��۟���՟��SQyZw� U��Ԩ+��)����|1s�OD�DR�Y����O!2������G-�J����W"Z�6 Pc��'���'+�$W��S�(�wN��uq��p�Y�d�\!�����M�gfΏ\���<E��'N���7@ �Pp2��#�P�6�g��x�����O��2RM�<�'�?Q��~�յ{��I�R�4YG����2B�"<�����'^�OB1H0m�85���G+!�v QR�i"
æ���П �����=Y���	bV,�Hq� k�b��g"�z�ɔ)���?y�����O�����O
C�@�p��6�
T��Rt;���?1���?��b�OZ�90j^�o�d}@�L q��PP��i��0��O��D�O�˓�?Q�cG���T.����ՙG	� H^�e�R��M���?����'crĒ�O�`hp޴+���VȈ#-�u��#���'j"�'K��ҟx�  }��'B�iY��.�`U�0�"X�f�c���D7�Iޟ�擆	?�O�0f.>Q�A�13W��h1Եiy�T���I�R�	�O3r�'��4%L%-$��i�;:��9쉟WJc� �	�*�>Hk�(�~��H�c��y���k�"$�e�a}�'����'��T�\��FyZw�\��¿V�4ܳ��.1(�p�O��d��\���r���	0%�&�Q-V[���T� ���c0<B�'�"�'��Q��П���͋��P���B���[��Mk3HьU��m�<E���'^^hɇ��H9�D6�C5�~� !�n�D��O��$U*0!F��|���?��'����:��a���T�:8�a���'&V$��C2���O�d��|u��]s��d�C�/LbG"f��d�:�N˓�?1��?��{2��7�*��A�` L��aղ��C'C��������	Ο0�'��,Ϸx�� 8���?�zt��ƙ]O�0�g]� �	쟸��q���?Ã�(�r�z��.&$�0!��T�=���r�ÈS~��'W�^�4�	�����'&2�	%̋!�bm@`ɕ-M��l���p�	����?���<o2E0�lV�A�3��N�� c�^�0���>���?Y,O��ă!i#bʧ�?ׅ��d��¦�ֵ}�4����N���'��O>�����d)s�x�C� ,ϮL;� ��xE:��`� �Mc����$�O)C�b�|2-O��I����&�Z�$y��Y,. �>a�jXp���Me�S�$���`'�Q�q,W=Ȇ$�hɋ����O���$��O���<�������8ժ^0S:��XDB�)R���p`[���I�~��m9P";�)�S�IH�!7�=*�Ȅ�n�;2`7�7����O��$�O�i�<ͧ�?9C"ɑ`�V�+t�	!�z�a�튔F��Bz�Ś�y��)�O0�BT,�V�`{���x�,A�p�ᦍ�I�`���dEL������'��O�]-�T��s�X����fx@�y��X�E��R���O����I\1 �%\�.�x������b7��O��3��<����?9�ĸ'w�5����,�1"֡3�噬O�LybaWoN��蟠�I}y��'�@�z&ۺ2}榔-U��[BE;g���ٟ�I埌�?��Q�������;y���%Lѕ2VL�������'J��'w���4sEGD����
�ذAǈ�'���p������	ٟ��	T��?��;�In3�Is�;(��yGΞ����?Q���D�O^|��|����<�Ԃ3+PFm4B���ـ��i�b���O �D��~��'Y���D!�X:�<���M7fbJ۴�?A+O���@�xp�'�?���J�i�b?��r͛ �S�/Y>�O���Ϗ4t k��T?H0��+�Z�ga<����>��~$���?Q���?�������(a@l�
�u�o֞0�"(��R���ɓD��x��6�)���Gh�{��!��a(1��07T6�Q�P���Ot���O��)�<ͧ�?	A��!n�ԫ�E�j��aV�T?��&��s�>L�y��i�O�5� �� ��>p��s-%|if�i9R�'}b�-��i>���ɟ�v���:,Jn�1t#T�k�>Q�P��/���$>������I�Qs�=���Vq�%e�^4�L��4�?��n�*R��	Fy�'��IƟ֘�s���q��;z���S��TV�p��q��?A������?i)O����M���a�啻%\��� D't�D,�'��IПĔ'�2�'@�T�)i���cD,w+��A�ʩuTT�r�'N��'tPa�p�';�T�r�������B���[p�X��ؑ�M�)O �D�<���?	��u���4����	Y�`��=��+��?�p}�irr 	���'_�bb`ѭ���d�7j�٫�,�Y��J�-@�*�(o�(�' ��'�R)���y2P>7��^K [�ą� ����6�Y�����':T�0З�S��	�O����Z-9"K֐��A!�)b�:͚�B�a}2�'��'�F�)�'��s�D��a�6}2v�Y��X����6�m�fy�癁w�7m�O$���OZ��b}Zw}�5���_�4e^`q��;Jx���4�?a�r�H����$K��m�}��&�c�`\Q�i�,q�`���):�M���?����pU�4�'I��C��|����e'<����nӮ�t4O��D�<y����'쉳�\��(*0�����ͭB��&�'"�'*�����>q(O��ĭ�t�G,�tz@ �6���m�b�i�oӀ�Ob�3�8O��� ��˟ˠ���ر�ӯ�(��9��I��M��> V�$U���'2Y���i����hȹm�`����)���Zz��!�FyB�'$��'�I/2��F��(^Vظ�jwU@��F���ħ<�������O
��O�M���ǅ�`Y'��#��P"��S���O^�$�O(���O�ʓU�4���;�|���NG��I#�/0�дi�����0�'���'�c�����W�{�љ��,v���Vf[�9W����I�ȕ'�r�E��~��{bT�7�٥�N����B76�8i�&�i��Q���	��\�I[���Z��4z�f�ۦy�AW�C�Tbڴ�?�����QQ��O���'��4�Ȧn���Jץ��"���kZ���?��?�]K��|:B������q���j�Q�ά�SS!�Ms(O��Sf�ަ	������I�?�ɫO�N)��©F���I�f��]r���'Wi���y�K�~���O���l�.�>L&
��tX�4N>ir�i�r�'B�O����򤊸l���Y&�>=X�˳@�
���m�R4~�۟�I&C&����'mV�q�_*O-��MI�qP�A�i&b�'�2+�##����D�O��ɇ<��tK�J
N����%��6c�7-�OP�/���S�D�'�'��#&蝁A9�󫚝zd�eV@}��d�7}�X�'�ʟP�'Zc�>��f��Cgܤ�S@�g�$0�O쨋w7O����O
���Op�D�<�C^�Ztԉ�E� 9��VD�irW�\�'��U�X�I��0�Ic�u� Bs���J�L�&��)p(|�4���X�E�˟H�	Sy���"�擲"Њͱ B͓1)�av*�f�0��?A���䓐?I��+����iŲ�a�Eo�j)[�""}$���X�l��柀��Oyb�r]�pI|�a%�V �3�lы2o������ro���'��'���'����A�'��K���ѡ!�%+��L��p�.�D�O��9��4�a��4�':�4��8�z�(3揑<X�B�e@�l�Oz�D�O���A�OȒO���97�R���L..<�rI?�r6��<�� ���/�~�����%���1S#� /=l���f�
%��A�`�h���O��ХE�OF�O��>)�#�Ȕ^��՛��_�~'е ����o�����ğ��$��'V�p+�Ǝ�f=s	R�y�i��y��qp��O,�O��?1�	�0��Ӡ��F����H�Ꮈ�ݴ�?����?)Rē��'�B�'�X�Jΐ۱�ʶHI4�#�[i��|���3��.���O����=jH䓑nA�/A$$��읉t�oZɟ�s�:��'��_���i�E)��!�DaEںP�C3M�>g*��?�(O^��O>�$�<I�Ɂ(�P��,��,� �Yu�݌�@���x��'z"�|��'{"�Џ0sl�xE'�{{����\�f�c �'w�Iϟ���ҟؕ'��� 1v>����.(Xj�ђ��.\K�M)� �>���?�J>����?�&���?󩃼mJŢ���q��#���+���ܟ$��џX�'���[��'mƽ�N�o�u`�D�S���D�iy�|��'x2�R% b�>	�ې;�<d۱�<� ɡ������Ο�'�"�y(���OD�	ِX:0r��U%��+�oN�"���%�\��ܟ��``b��&��'8��1����eQ��[RD���mty�& "̀6��[��'#�Dc(?���M2�5���3,�4IEm�֦��I��0Jr�Aڟ%���}z��Ǭ����hV%ۤ)a1��Цm+��^��M����?!�����x�O
f���S�a �*A��&�L$�`�s�x!1M�Oj�d�O�uF��':q�΀��
�I�M�</-$���pӪ��O���W�/Rn&����эU'y�ħ=�bY�Ʌ,"u�֙|��/Q{������O��D�	L|>r��J�ہ� +��m�ǟ`
��T���|ʎ���#A !�#%�#��`5`êb�6�'�"���'��	� ��ʟ\�'Rh� �Es�cH1��
׬N�;�F4#8�'b��韰�P��=����gnۃw%��� �.yƴ���}y"�'�b�'���'Pp�۟ ���!7\�9�c�ة!�(c1�i��	şd$���Iş���$�4�6-\�]�f��1�2\�2]�pj+�������	ß\�'W��Z%�~��[�R���ܫ$P�(&�>b����V�i��'��O%ڠ��ڠ��@�ЦZ7�uHDhX%JQ�f�'qB�'�R�H A5�Sly��O'��6l�VR>y����Fk�̲l&��O���47�x0�"�T?��gA��@ �	�
l�\��w���d�O�Q�M�O����<��'�?�����
��b��$���t�XT���Y�	̟�� �45?b�b?]��95`	��ɸ0����"ii�j���R���	�x�I�?u1�O˧n�$��k�& ��(�H\�]�G�i*(7�D򟂒O���/e^J8!�oˀ\�h�ڑ��=����O����OH�h�<�*���䡟�Z7�L�:�c"��8M��١h���'�:L�Q�:�i�O���O����k��=u
4)c��-*�H��@��ʦ�I�,3n�'�T�'�?�L>�.D]�lt�ʜ�
`�',9v�	�"	�Aг������4�Icy"-/y�́P���./Zœ0����禼>����?a���?��Ț�?m��30�O7k�DU�P(�+f$rY�A�|��'��'�b�'���kf�'e�� �W*�ZP�d�/�����x��˓�?�I>���?iB��!@9�mmZ�U��90W��I
�2����%�l˓���M�Xx4:çKT��w�[����!���c*���ȓBN)��NL�#��{Q.��Z����JcV��v� �*&��"/����w�e���ǉ��t.6�RC�M�G��"AA؎V���C`ƋK��ؤ�^%$x\]�6o�#:�L�
@�{�0���Fאb�L� ˑg�X�&��$*���7"Tp�y��%^>ap��F^<�@2!Z%Oh�d�Ab�
��Ⅾ:��f�O����O��9TBS#qC�HCd�"�>�80mKtQ�c4\�$	45)q+ΐ�dH�O�1��gG1'n�ݐ脩d]`��¦<wy֨�q�W)�"��3)��k��ɭR��pn
2V.����9a����%����c�IP���䙓��	�X��'��+����FX� @	d��<)@0�ȓ[n��P�E�U��Y�Ě�k�Fx�"=�S���#��9�
�vQ9QNנ��'��1�U��"�'��'�v���H���g�ԑ��h	o�^$@���R��PB��C�4���g) �P���?�=ٓ�S�Iy�0��(_?}��-��
^�B��.u��=J�@i�g�'��qKҁB<X���xf�E�t�0K�'��B��?Y����<�Q�	''��zg�/v�����	�Z�<1���
��`�[*l�D���㙓|������$�< �o�J����"5XX�/G�uY~����t�	ğ4{���Ο��I�|�1�	)@�>T���Y5g�"m�@ł�V����,�VT�z�_���<a&�K1/8|K��7�$YWIv�7��>)�t����-?N0��	�)����O�@�'xcB��D��"��`�7ړ��O� y�Ȥi�0���$ V͙�"O<4�� <5 h1��޺�Y�9O�=�'�I�55��s�4�?������8�
|�7�ԙ���;-c,H��-�O��D�OP��!�z������S0~���|*h{~MK3͂(~�� �W�'b�CnCC~mb ����9)dN�ﰴq��-��i��݀K���C!\R�'�%��Z��gl�"�D�|�$�KW���C��ͷF��02��?1���9O�iP�ۉ&�ڵ҂K�8Ln����'�O�\��G�kf���)����K�6O�rv�Φ���⟰�O$�D�'�b�'HT����g?����l��F:����XJ"�xd5�T>��|�IS*�M�vA:9���gƍ�BV$��dP�X��D�J>E���x���õꂵ+".(� ��	�rԋ�	��?����?������Ҋ]�{�UP NK  ���Pҡ��y�'��}���9k_"�b�Ǽ0�d)�/��O�Dz�^>��B�$�i  �x�����ß��K/��������Iݟ��	'�u��'4҈�v	r`�B(�b]������~�f�u������ɝcFB���	>v����ʐ>$���ńpw��I��&H���K�@<���ˁl�꤂q�N�N�ָ���ƃ$��Ռ;w��mӪ9l�V��a�S,,�楙q#ŀHRj��`h��izC䉥u�H��� �|H��3V������Ē}�Q��6��'�M� ���	:���� �Sn��Ā��?���?��t��8���?)�O=6x9�,�>�͙4��.��(��ҍ'�6��(X�~��X���'�����UIӰ|y�"Ğ3?$�#N�oTDB�.ֆK�$H EB�	������dJ�AiR�'����E,K�b��ѹ1� ��'K�O�}Γ3k�sʟ����K�ŕ?tTQ�ȓ�$KgC�<X��ӤK�>�L�����qy#U�N�7��O@��|RgOF��+f��89��[���	F�5@���?���=�`}�c������ �|Z����HA�@̕=�}�S�	6y |J$ڧD}li�B�n��a��c�<#�R�Dyr�Չ�?ɋ��@�s����Ƨ �h�0�g�13�!�!_
���:��('۔�a|��;�R���X�ģ	�M�xDJ��T��H�p�TnΟ���k�T�ؘE0"�'��
�	G� ��R��7�4��w��+`��Hi���'�ia��M9H1LqK5ͭ~"���;*����@��:���GEеUTn���9/c���Ŏ�I#��փ���>��'��tم��<M\���,�Cϐ|�Ai�O���"?�[��?��Ժ3P�Eʢ(˕'�^H�3#��<y����>1w��tF��;GH�z jR��A�'��#=ͧ�?�Cއx���:��Јn�@�Q�&@&�?���J	�\i���?I���?)��j���Hy������M:AfQ]d�ré�����*�"�4yaE��p<��b��*��sD�ɦ�\JaY]?!R�?@o��fg^
t��x����B:�j�#��Z#�� `�: *�Ð�Fx��'n����O��arX{�/L��YA>���ȓr7$� f�``$$
R�N'O7V�Ҁ��}�$[��P�o\:�M��	�6�xep�f�3[����#Ā��?q��?1���������?��O�Jh��O����ƚ�}^�� �Ɨ�Z&E�EXY v�ٖ`��0<I o�7$�:t3���('*��@N�d\�����$Pl
=ˢރDjP��	�-&���֦���E�/���`�,��D�"$��M˻�M���/3��<A�He�t�a��"���#��HP�<����?tH��Q�i>|�cr���<���i0[�(Q����M����?�*���#$�K�>Iq�%�p،�2�±9���D�O�����$*�|�&�7n`��eם$���ٷ�r�'(���ӳ8���d/��k슁H��)0�T�<!�N���IF�S�pƧ>sx���0%W4ef��T������?E��'�`|���%|�5�[g�R1��^#�'��d�gڤ(�A5�������'!^���{�����OF�'0�R�����?���p(��ڤ)R��t��u_�1!
�o6��'�>{h��Ȧ�'���?	dl@�t�)!BldQx|ˑ�_�@�� y��U	�:5�E�",U"%G���r ���\��qyg.4F�|�1��?yC�i���'(�O���',�A�D䠱��U� *sF�ֲJ"�'a�}b�S(�4��'�Q=K��U�uŒ��OP�Ezr��>I�MF[�ji�f
K#CؼY�BNݗ��xB�=9�d�)D�i���펛�yb��2r����Ψ`&�� "+͡�y�l9BvyB��U^���E*�yr��W�Z���@�	
򭨑��y��m���d�C' �N�pj'�y��*����F(�0Dڄ� @��yB�� 	�)b�k��R�t�1"���y�#T8a�� #P�4N��b�
&�yb�ϠW�̪F&��x��T�G��?�ybjS�\gj�5.��l�֠���ʄ�yb��fR��3�	�f���+���y��?g4��A"O�Y/���K��yB�_�#-dtZ��@�Q�l��bO��yb��.8e$U)���V�D��"K��y�g�]�.����	\0)���yr��8�&8�'J�$�s���y��@t�D+���%r/<��1���yBbM,i�Ldǎ�9l�Ұ
���y2G'w�,8�F�_k�8�P��y2 �g�*�BrbH�h�RYć���y��>��S �[8]��ICc)��y��F^R���*�9`>����@�y�a��.,F�p��6\\ޱar��4�y"��]��Xs��T1V�ٱ�o�ybh�
�R��2�$ Įţ����yr�	�w	�m]1
*P '�y2�1H���x�cB��,S'�ͱ�yb�%ź	h��M" gF��D���y� @l��#��w�� ��y�J�#J%���Vn"�9��>�y
� ��[S�ݴe�psj�g�\ls"ON�P�ʚ�
)n,����\�$�A�"OZB�[ E���	�K�fc "O�0��,��z�N8p��A�t��"Ofa�h"�������#�,� F�>QGAW+kǦX(��`�"~�#����1)��Ց�l�Q�*G�,���Ol�S�"W�?����r^K��x��˚8z�@�.M�mc��H�C�s�<��U�8l2�»d�T�2K|*�eĥ7I��長u��JE�H:l�(��#��HAP,�℈�4�����z2�Љղ�O�KGo�E�H [֌_D�60��%.&F�RP��xCrb#n���`dj��� ZԈWd�60$�����״"�Ʊ1��X3�(@D��?+oQ�L��$�-���<Aʐ*��'�"����6�>���A��D!��!�>n� iq�*y�h�5F$�|B63轢9�AB2V0��v�=����8
F�7B����фQ��IG�e�e^���eI𮼢!"ضn���ɨZ.PAф��)^��L�Zw��x�7��+�4��v�>��IC���S.܃}94M8g
���3�c	��?ٓO˴n`�%>�y�/��-���"�[�T�(E�'�[Qyjm􂓷N�\#��C�9����Ɩ �8x���UP�'��e�O)A�ltKGO�c�Z`�ۯ?H`�Qb�^�4�xb6*�Ev�ܸG9a��T
�K�"#�ɏ�`�Sv��p�8j���0�ƨ�V
"o��IF}���&ؠIeb��e�!�p�'�ּ�@dN�*�!�ς�l)4��`݉M����%j0jx<Y��jq���Dl^�]�� �O��睭I���AJ�p��PХ�ơt;|�T!|��G��#)���3���h�F-A���^��]�`K�:��a�Dk��<�E��7�����A
<�Ub�jP8�mc|�'��!�<[J��;�c�h���Z�� ������'�ƨ�����ħ;G��)]-s�j<�P�U��y �T,�(��(C4$!Z�-��G�~�C�ʜ".	2EA���Y�5��S��	Ued(zZ��$(0����(�区�<��I�B#�'r�=����)��u9g!�8Yr(����	�1�<�6�,���#�Z,ml�%�K>�?A#b^�*�]Y��;y�*%y�-Ou�.���{�F�?嫂NԜ@纀д�Vc����cKְ�=�L�H�ˎ�!��8y��D7P��ϐ�l�rʆ�g��iI�c�n����1�6�����#���=���1�uw��-_^�a�1.ʆ3��>�<qvRc�H���.>��1�o�#� Ton�y3��/z�L��̩?� �y�DR\���Qc�!Wszx9A��8;�@5"���Y�p1���S$H���I�NvX�Z�A#>s0-�'�x��4�`���EZ��o�%�b��?Eb�� �T6ݸ�lA9,���Xq�_ư=)��U����1n�b�� �A~�0�֩��|����(֙q9�]y�,�e�O ��O,Z��XI!s��;1��bs�͏ɘ(� �	3e� ��F7�u��P�_����L8!%��W�R�P��P=B�T�#�Ĕ3�~���o������቟~vŉ���n�9[�a�,M8���shG�(��
����Ѐ뺟�����AkL	�K�F^r�23��yYph�΄ 1<�~�a�-g�&���l�}@�jA"�&���p�'; ��"D+R��1�O���杻��X+����E�
|s�&U�*"��䋳v)zU��ͯ?̾�[�� �~�|Dk3��s�$U���K�Ez�!g�H�O���"҇��(�&�%?����\�d��1ۑ�N3�aإ	*ʓ�����L�$�0ٕ�^R��`��?�˅Hv7�z"읬+���!!�4����gB��x�jZ]���g�'�
�ZG,݄0o����B0{I�y�JX�H
����5D����ְYҸ�+Qm�yü�h��
Z�n�!�ۚRU����"_�qK��'=�n�r�f	�Uo (���D��ʓe V��O8�q+�+vK�wF@��͉70�*�k�ḿ2�2���'�.���%��a��QfC*9<����ҭ��ɦ�y`%��O��S5$J�w
�$9Щ�h%�I���V6D���'㠔z�/7'�Y��O�<�"ŕ�8۶�	���!<	C� �m�\�͓ �n iʃd�����O���Ȟ���Q"ak.j�����$�@��oW\���~�g?��# �~��e�B�b�̅#�NE����C�L��~R��P���a�(F0s=<�s�ȴ5��	�S���T߱bS�Γ?��,��l����](�B�9rY��@�C���S��:�\*���PU���@%`�\��"��"��	�e	E�K
Ur�E`�I�Ou��/D�M��x�t��!�E
Z++4\��$�1o�; �HAia��\qB9e �u{��}�Iz�+��^��������G,���?ёH>i��L4S�h8���k�q��X~R#@��-᠍/q풕�bB
-'5�g}Z9n���#��r���㉖1&��Qc��\x��z�⛋66b&jÐ0x& a��ߎ'���jg+1 "6	�o0&��ֽ<��py2�؈k,��HT�=�y8�՜1
�CC�'���J`%֠N�� Kޣy��0�g�+�b�h�<a�ˈyh��K:�<���|��w�R�����HӖ�뱆�'�0<��֮r�Va�2LO�q�.����ۂ�����b�@ƿ�<�p���y� �d|u=��W�d��:̔���W%hy&�'��(�/��X�mR��ۣ4�t"T�O���� %�$a��
SL	6(�I�uH��7� ���O�J���� b8q�@�5H��qHyT*���-�1s9���ŪYG�C�b9s�P�u�H�	X19�:��T5��Y��!Cx�|���p�h�O�X��	�q�p�s��J0Э�!Ǘ.V��HPw��x	c�A�~��h��܁��P9o�,�K>*�.1,���.Cet*6lY�$H9��PdȒ�y�-�%7����᠝�M��� E:Y�E1�`�S&ph�`�I�~��<"�G@4�f`9a
�O���'��ܩ�J�_X��J�ƿ{L��0�ڽz-��N��p��g�ŭ���WB�%�y��D�] <e�BFm&�\���A4�B�M O<Kw��Ș�M�5I����.��v�0�(��PDX�M�"l�O��$��#8�D�ƻ�` T��'/4N W͡,N  sÓQy�u
ؘ*�ds��@ ���Ow��$qB���pr�ăV�U�;�t�0�f^0c�:K��^(�^�G/�hOv�bW�N35���0��Ī-WP�%��̓ebQ�ۮ��CƎl*�k�N�>].�1��e5t��4S%@qCKF�094�(��7���2Q
T1w4dE���+b�TmҕB�o"���!L�o*.� RF��d���(;L�T�&��	&mDL��O�A���U��.?q/�*�.f��e�����4�!�$1���[��܃Laq����QC~�D�q6�X��T}r�6`��e�ѠB&�����߈��D��pN�]#�H�d�%��*TiLax��
��%�� &!�Ia&LUg\FI��*\�7$ �����C�m
Gm��K'�D;�
A�;&�[5�'���H����fn��͔�FB����O�e1�-�E�	���WI�Փ��\G�����MC�n��.Ġh(���i���xBaJ
F��\J�@�Ow�Q��-u���"��م$ U��G���D���鞜sj��!6�<Ս��n�`Id��lS�c�O<��X�h�QD �02��T��K��C��y��A����L�$�+p��	`D���'��K����wˎܘ7�ƽ� ��ÓL�����מ���"�_$��[H� 6�̥z����&�{A��U�`�L�K�|C�aR���<YA�3��0F�T2ig�$��XA~b���$Zލ�*ƓF����e.K��y"�ܺd�r)�'B�(д;�F�ʄ�Χl�<�ȓ�jM�5-��VJhѢ��M,�N]����&S��j�
��Ń2�Շ���<�6���S3�ܶ��ԉ� ��m`L�$%\c<Q7�̖?7������q�D��dfH�q�0D��M�.��sú�9�):Oڭ��+D%D���N� :D<�@��j�'vX (�2��cf�Q'r��A�u�����8D��!Y2��eZ�>� [6���y'H�D�;#�+x����v���D
p��(V����`�|�<�����n�`���CD�a���x�t,vS!�"�����Vq��O虚5�^lh0Q�B�ۃ`��A�����tÂ�O�<:��5��O�:mQ7��?Fhh*`�4�y&��65h�a����b��M�3��pԧy�K�R
8�RA��]8���)ڼ��~9�P�B�=%n�$?qHg�C�9-��N�B�P�LK1��`˧J�Vz���$/eJ���"�<*�c���O��zc"�/���ŷ'&H�NɈs�RA�'G\�h/���L˧x��sŪ��y�ݳN6YU�εv�*Uhe��$��	�+m"T���X�	.��y�a2�O�T8`CO?.aĩ�rfƚp�r�����>�ԣ�F�8*o�$�E�X=�%��tj�P{7k]"��L��5q�X!(m��Ze̓�J���Gi���{"�yӐ4�VNΈN,8� ��	�4G���'IbpȒO�$z�h�Kg�:Nh�C=O��o�2t0Z���%7�����W���ݴ;}0w�}�$�g�40Z�穠|��iw:�D��U���CE%{��rs�Si8�<���ݟ�pA�*v����dg]F�l��F(+S�D� S�Hv�cPŗ�(���
�HO2�c7�yH1��C��7�RE�0�D�;)"M�i�ihq��̶a�Mr��ԬW� r��;���&cr0Q�W=O��	�S�l0"%;Uԭ S�x��Z }X$ B�#�0�I ���t��҃Mt�剄���}�  w+�Q�����?�R"��f ��C IցEa����J\�E��Ծ2� �8� �sP���Ƀ6M��sCK�!�x�%��7E*<j��y�ρ��\ JЁ�����?���U�󮏳%�� �d�C�;�Ȅ1%�O)�9Y�Ny� ΄~ͤU�� ��Ń�
D��U@���x�M�5	C+��B�f]%$��Q��6Z� �����<8�
��y����|�&M�.s�p8�&����'p9�"��4c�	z��9O�VJUh^��@�Ɗ���B4k�D��f%�H	���(VZ����Z<Fi ��Hq�dޘpe���� P3>���J�lΫ6��SZ*�ʓy/�ɬ�<�R(Azl��0d�i*�o=���N1w�dTK���M����3�:�+⦌�*�@�RǓ3��`̓�9�T� �!�*HL�8:�a�KV�	�t+ 0��P>�����^�N+$@G�S)�H���㏹n��D��%\� �F�f� ����~�c��WJ�i�`+�,1@I�u�F|$󤬞�H6�Ē!n�y)���h��!Ēxm�y*���'��x(���$|�i���O�YPA��Z�j�ㆀ;��[��Ɋ>S,�$G��D4�uK�}���4"�X�p�o��t*�I�j@J'
>��Y�B���'�$ݹ��Kv
8�O"~�Jc��;Avt�ï�&�����i��x#��_����,ˡ9��xRf�/D�N�*@aL>kVI
��oeV�@ �����"i�d `��Rޟx�3�)� �P*v�]V�``�Y)r6DA��FEH<q���_h�ix�CЛj@�Y8��V�<i� nC�\+BD�0�nq��A�M�<�5'��v�Y�#(T�CVf=3GM�d�<�ao
}ۘ��r�Z/\f�`��h�D�<�BA�4hJ�����4<ۦ����}�<񓮇� �ʔJE��}�H@�Qo�<9�;]����p�9�pU���e�<���C��Yxq�Θf�}���j�<�r�Z�>���W<xz���� �g�<��@��Mh�C׫�5-�h���`�<�q�ˉ8�0���5BxH�!q^�<�g傗K�Lz��޲so��I5(X�<Y���(jc�pp����=��9�5�PU�<�R�v�y@֥%+�XI�O�<��	]���F`)%�tb��c�<ٖ�ˀA��y��[�v�V}���Ew�<��	
1�^��Q�J���0�
�s�<i�2a��ꗁӇZ�$�!s�<�� �
r�� ���Q��,�Q�Ap�<�&�u�l�!+��Zx=I!�Xk�<�A(��p?�A���H�� �Ae�<�&k��j����P�oA\�R�^�<9�I�(_�l�:d$�&;�
�ŝ]�<���&x��	�Pg�gk$BT	Xq�<y%cO?&U�ժ��x�Ybab�j�<qu�+��I��ޅ|��5�\e�<���Ӄ_���e��"eq���b�<q�S6!��	K�¿�qn`�<9�.ȞV�$�
>�����_�<�n܀ZJ8:ak�.z��MI �UZ�<��lT�c����Y�]Kz	Q�A�n�<A��7[���Ă.7�t	�'��P�<�g�Q�'N|�2UGS�2$T��d�R�<��B�>�㤩�&0��)j&,L�<)%�/#B��'o֢2T�Q��F�<Qgj�S=�����ŊEv�ق�B�<���\�:���2WjUA�j_�<$j�zk�@���\�MjHI�� b�<�g&��H�D�<Z���Ї�`�<q"Ś/f�E(�.V��X܈do\t�<�/��}Ψ�´ǎ<LN��Xp$�I�<�qɎIRz�C���8���0��H�<QS ���!�D �,����E�<�R�%&���҆�%h+���g��B�<� Ӭ��VK� z�nq�(�h�<i�B͟S�LUz4j��BXۗMj�<�!-ӻ:f��� A�����f�<��脾s,�He�ɧ-���vl�e�<A�Ί�C� h0��$�J�w�F�<���1uF��6�ߝm3�H1�o�w�<q!"���܍�tiqkxP�CH��<��AM](���J�S���Tdt�<�3%PPpF�{šDؖ&)���s�<���֍�������p�T��,�r�<��El�����><�]���p�<��v�b7��� ��q�
y4PC�I�dڈ�p�/	/Q�ܝQvd�>$�C�ɛ"�J�Yc��5{��9в��6!��G>p�l	��H�P��@ku��
e�!�ě�a�ȫ�@�/*��`3�ZT�!�d=TX�uh��pd��k��!��'KF�C�ʒ�yf��*-Ɔ��ȓq�T��Cm�YJt\��`�U*����S�? ��$i0�83�i��w��p�F"OT�A�K�9s&��+���Y�"ON �C�ϰ8, ܈�+���1�"O���'��t��|𒥌%�J�1`"O&���D!y:^a)%/�0�����"O2L㑁��7F�|��P2R*f�B"O$��٩7W��A���B�^���"Opy�`��g/�A�կY���A"On�h媃.w�T��D��rc��"Ob!�7@�^^T���i��x�8TA�"O��s!�"}Fұh�i�3��`"O�$���'`�ȵcb��_���r"Oڬ␇ַ0s�\c����z��8��"O����X�m�Mq��]�ت�"O0��)�:<M���(�b�s"O� 룍��(ơ�㉈�N`i�$"O�$���A�lV�akW���a:��'*Oh�;�`'�j�{B���,���'�����L�d���Ҷ	�|Q`�'O��"�*6ɪ]����:��
�'^n���1i6.\�@C8t��c
�'t�ݸ5˗9f�Y�f�C�*b0
�'5���S�UrB�Bu+����	�'���ZW)M��e�O/�2r	�'��8R"וk�V|�t�_V�r�':�k�@m��	�J-wbQ�"O����9I}hPegP6_N|`�"O�a���ևH���kί^X� "O���"���8���ӊ�)*�J���|��)DҠ'��]q"	��	B��C�Iu���X�.K�/R���4`
��C䉾:9<��셤e�XD	TC�;P�C�I?_���;�i�/qyp[E�s�\C��+u�~�)V�L'l��5�Gi�"'��C��,R�بS�69���s��H��C��/��5�9Zgd����د~�VC�I��n��f/K�2�NYH��'G�B�I;q�b鋔oWf��TI�� *�B�	�&>|�S@�*\����5��a��Oj�=�}Ҵ�[%`&np��O
@��*XY�<ّ��Wx�Ӭ��_;�(h���U�<��lHN�Z�H�:T8�SWF�T�<Q1O.c����K:O:�k��TO�<Q��*��<��!"&�$"��N�<�k%-��+�MΤ*���1�  F�<QS�[�k������+t���AlTB�<	�ȖcH�t��o�f6,��1(\F�<i��A�����'J�}.L�<�����=�G�*-Wza�㋟E�<��pB i�䥃D��AQ�SW�<)�,[�x�F|{r@�."�2@F�T�<�7i�G��a��O�&2	�r#M�<YcX�>N��+U#fT�eR�FH<��ǵGs�[p��?o8��U��1!�L�M��!
�g��d�E��O5@d!�S>�ʔ��:=�`�b�#C!�d�0`j(����$<��V�H!��
?j��C�i�!�h���*ռn6!�R4`�r��g���m�6%�S$��J�!�$���[�,� ��T*�c�U�!�D�������L��}�U��7!�dS50BН����_��	3�E3!�$����rb"�8*��dp%"�
�!򄘺eq�a�������[3 �!�� >�����Bp��E�#0zH"�"OԘ;�+՛:����ӫV0XJP�
�"OD������4�;��C�sܖ��"O��vN�5�J\��nل���� "O�5oV!}=Ɲ�r.�4��Y�g�'h�I;v
� 7�<j���#��:`B��,M��yz�'G2�΍��K8NG�C�I2����4�E>i�e9��_c B�I�A4Up�j�=]~�z�ğ�`����0?9��X�S��av	ʩ�^p��eTL�<YM��7ft9jw�Dp�eTJ�<v�̲:E�(
q+C�$k�n�IV���O8�y�Ȍ{�	�0�4Y���{
�'Ⲙ9�T"NQ.z�K�.|j��
�'��$�Egݱ@Uha�a(��	=���	�'�����B�jK�}\hE+�'v��W�u�@�0%��?oа����'T��rI�	O�f,)�Fޘmg��8�'Nj�c�j�(��8 ��b�:� �'z�̳�c��n]ҹ ��a��i�'j�"�U�~7�X���[x���'�|���
�5�r�H���i��]��'�JH�2AWA��y�@��b�����'�@]��ݑh�8���(���tp��'�R���b�0Ext�*���?6Q���'L��bD�Ih� Dj�5- ��'$�I8Gh��<S��u⋛b�r��'���/��'����ϽB�d��'D&i
�n�3��(b�߶&�VM�
�'�Zț���3[�Pɑ�I�%�����'ou�j�&+D�g���p"K\�<��Ǎ�40��"S�لL��eȂC�s�<�S�U!5�B�9!��FW�� �G[�<a���P���	%(U�<���QS�<Y�@��	5���%�RB{�<���!{��b�C�s��ʵ��b�<�R��|Lҝ�5L
# >�@�ZZ�<��!��Y���N a�%���m�<�Ӌ�W���#�@S�����-�j�<�4-��2�����-1��ȳS!�P�d3�O9��"�(6T2a(��-}� U�'Z�]�-���#�
ND�m)� � 5!�ē�=K�8�$G IԊ=����2.!�D�V��I�0M�d�z��ac�,#!���TL�Z�"H�\Y�X9����?!�� "�L��t��AG�i�훗M�!򄛬��-;IE�8�X�+R���S0!򄈖@�� �EK���0h�q�Z?H!�r���\���5��-�����'4�|[��F=0�+��F��08��'sF���'J�l�)�E�)EHP���'�~Eړ�F2�6���F� A!`L��'�`{t��yE�pS�bY:)��H�'�b�ɗl��G�
p�s�Zs�:��
�'�ވK5b_�A�^��u,�,i�2	��'bd�
 h�'�+��ēe�0K
�'������20n!�c��+~���	�'�N0�t&J)=t���B��:����'�88U
9t�xc恧8.v\��'�����	CZ1��M1NA+�'��Y����+�>E2ଡ଼�[�|�����X�L�, �f�P�Pe�k�!�!�dK�*�D��iɇk������:���Gy"�@r��5\{@�:�) .�6)��"D�� p��`�|��B���!:��z�"O��D#\�m�X�����F�(���"Ov�����}DtE�%�  *<"Ds�"O�A�'˧J�,@,�Y��!RT"O*A��e�,HF��k�dѐ�"OH<{�F�S=`\B�e�o�u2�"O�Q�t��#g�}��.��p��"O�냇P& O�<2$��< fy1"O�y@`L/������F&0��"O�A��GY�^c�A�\=(���"O��ի�.L[��a��*5S���F"O�l����'v"VxӇb��"(�"O�AC%ԇu,�t�O[m32��"O�\�pE��&�(��D�{H�M� "O�\��MWse��ѐn* �"O�T��jY�P2<|�m��	$�S�"O^���G�K>v��3��K��1�p"O�!��H�;V=pˁ�Z�2�[�"O|�i֢�7ٜe�����֔��"O�%#R �L� ��"/�%q���"O.���J�-Z�h���4Ih��"O�<a�N���36m[S	Α2�"Oֽ)�'##�D�{��S�O:�qE"OtYv(�5e�\�'oL�b�\��"O�8Q٤z1�s5�'4j�t"O~�H�Μ�s��@��U�4"O~U�2�ʜ;�^q�����^��#"Oj̠�Yr�0b�)ڎ��"O.��w��m��)��N!�ZuA�"Oht�-�\��9ڴ��%�>hا"Ot��3
�2�C0N�:���C"O:U��MO>�1`�BB/#�8���"O �5�Š#��CL	�f�N�9�"O|xp���HuS���r�.���"O,ar�$4C��a����i��WT�<�#c�-3�Aۦ`T#zrH�7�e�<Y����m騙�u����B�&��y�a��3��l�@�_B4�9�$H$�y�e��vŮ	�R� �0]�  t���yBjo}�5��lK�q�Ty�E���ybd��Z�|��HC���h�뇓�yRj�W��Q1)�4?��qy�H�9�y��E �J�h�L�ijФ�S�y�Ø�8�n4��q������K��yB'ܥ{p�Y�Ѡ��a~�!F��&�yr��*.*�"��	�X��9��
��y�D�_�T	�ҬMX�F18��y�j���slΈhZU�B�%�yb�DWv̛ %W�k2��)����yҮH�Z��l���.1��y�bB'�ybnK��]�3nݒ/��T٦	ѩ�yb�@~�<�'H� ?@y�Ȓ�y��R?J��HC��ܬ8�6�rt���y�WQ��()��5M�9A���,�y2�@.��8+�+�8B�`��3�=�y��0Zp�����q`�%�����yr*�X�~ ���Z�4H��`ܓ�y� _�p0P! D��]q�逹�y�ȝKp^My�ǅHpf)�g�Z�y�P;x��:#��9����I���y"��v+�%�DHþGό=��\��yO�G���ed@������4�yrm��a��[6�:6¾$����y��(y����'��SU����y
� ֘ڗ�М�`�ش� �(��"O�T�$�����u�S�^�hI�"O`(��B߉X��Mv�B �p���"OF����#�"Z	0H A��_�<q�ٗ1c�1 ��IPD�2���`�<�B$�,��HXd��;Rt2`o�c�<�ƮX" p��̧	*�)��b�<��拖#����9 �\`@�L]�<�'a��R�`@�[7CN��
S�<����W3��Qr�0SgH��TO�<a�gԂ3��@��#��A2# 	M�<ё'�L�|D�B�
f\H@���`�<a�M�zU��R���gYq�<!��F>:"�i���(
jT��/�n�<�bFG]=��/�0b<����T�<Ѷ��I��b���cw�8k�o�U�<��蔖x�L#Ɔ Hj"���)�l�<	Ă@
&�9;��ٌ1Ƹ�ϟr�<���UM���K����`]�J�k�<�� YH"���ٽ�(Y�Zi�<y��1E"�viG�����c�f�<�4K�c|�-#��՚g�hH�4c�<Aq��Ii� 2��>l�ډ�pE�[�<駤H)Hp8ySi�#UV�-�Ԇ�r�<ɲ�3\�����cW(k�b�[p��e�<�V�P�
rD��E�,>3���CLF�<1i �
���qъ�+7xۄ'Jg�<���� ��M1O�>�鵬�X�<Q�Ӎ`�|"�mʃ;2Rm�DB@`�<	bMO?6�J�P�ƿgg:�rgj�Z�<Ap����(Lb��6g4�%��~�<��#ݚSj�Q�rJK�pr$��1�P{�<!�S�X\~��C�K��P(z�̂N�<A���AF�H�abZ r@�^q�<1�*��l-�!��	CO����[n�<)�jP�P����Y��Ѝف��A�<���
<��0�w�ʜ �$@}�<��A�:h��9ՋY�U�\�$B|�<����� �D�B�^�J0��F�Py���%Xu8�:Fe�q|^ur�e��y�d��u�h��,ӉS�n%#��y��L5!�f��G�I��x	�GA5�yb؈��v��"u�� �ˏ,�y���7h9d�ȼmO@�1!���y(5pZ1����OLC#GV��y�A
���,i3F�`��Bo���y"���O�FL��K!Pqؑ��y�gH��b��a(���9�"#�&�y�HJc?0���]�qzHQ�\��yR�Ƌ4���9GO������ߪ�y��X�}4p$�j�0k&�#�o���y�C+֩q���%/~�MIs����y�
W�k(����ϯu9�i2�oʽ�y!F]z6a7��6 :�C(��ybd�:x�tJ�kP#*P9�����y��#AL�±-
�w�8��`D�y�b��e�,�*1�6f���K1�R��y��ݚn�Xw�>Z��(��yB'�-G�$�c����8
���y�J] F�l�#���
Cݜ$0��K��y2EH24�"�0��Q�H)8da���yB�&X;���5'��V$����T�yb�Pl��,9�kXLH&�y���yrK��o�pʒ��SѲ�v�_�y
� �*�,��"G6��G��Oł��`"O*����X����
\cZPW"O�9iEա*
�M	Q����x�<�耹(~ ���HQ'u�^I!�B~�<9�,R�6� g�U�d�P@�Ey�<Y!� 7a`A�3 ��h{6�%�^�<qf�ܻrz��O4U��ɷ"G@�<�ႌ�
�E` ݅d~�U�[{�<���H�y�b���<2�<��r�<�_/Z���A��'�y!n�B�<�՟[��<� \�����|�<�V��/> ا�ݷ[�8hdJDA�<9�f[	Ha��L������C�y�<'-G�C�ּ��-$B����}�<q5Α#�D�3�m�.r�lȐ��_�<�r��_�Z�c!��2�.@T��Y�<I���I�B��q䈿gM[��Y�<Y�cD0#,E�@J=7�.�r���}�<Q.о'���Ea�1�*�*3�T@�<�w�,x�|Ҕ��#8~4��|�<���480R��	�}�����y�<I7jG3 cnEC@��4��Z���s�<�"nY:L�ƨ��L��|l#��q�<1*�9H��MP����b��_n�<�Ϛ�S!�}j7n��?}��z�+�j�<���ǁO�PEY�H0$���uA�^�<Y���\4�Y3 �3I�Ƙy��F�<Y㩕y�,�	�ǅ\�"��@�<��=vzٺ����&� ��A�	w�<	������p��U撨�F��u�<��F��ѨMK���0y\i0�̈́l�<�f(�2�(,y�Q!s����%[l�<��2Pe�Q�­\���� f�<IaMP�r�n���B����(Kf�K�<QEJA�;������ܢKA"f�l�<���>vŊ��Q4 ϴ�b7�p�<��i�N�&��`BJ%v���E�c�<q��X�P��
�Ȅ3�,���o�^�<�ů����&BO�Z�4h'K�X�<ɲ���Nu�H�e�L�H�#2!T}�<QS&C.�&J5��Y����S�<A��a2$�d�IlH8�D�[�<y�@cI�<��>�d�1��JX�<�ѡÒw��=$L�\ t�qC�[W�<٥'ΕF�$0	�GM
D�IJfG�T�<����ߎ��d���l'D�4O�P�<	�Ɂm'H��"�
�h4z�
f�<�w��cZx��L�gcܨ�V�R_�<�P�Ӱ=���X���<|���uU]�<�1-��%%��уh˶LV�rj[U�<��K��5I�؄��9,�a"$i�H�<��%ݼs���H�,��hኍ"���E�<�G�O�"?�[�Ȅ�)��܁ao��<���� �>��\�ac[e�<��a��*�x�fػC4�% �_�<�t�K�>����ܲ��0�Š]�<�v@7:����'&!X؝�g[p�<�B@;�p�cn��$���䇝k�<W}, e�F�	�C0�Ph�<1Do�(Ì���U�3�!xE��m�<�� ;Q5,|㯊�>�~U�!MMR�<IP�	/6�м�1nPR�*�� ÑJ�<A�N�R��a0M�A��(ΗB�<	C�
�U�T#F��Ӷ��U�<�  ��ަ�l����+�V0Cf"O �gg\�b�<��`�%'8��p"O���%kE&1Y��WÇ����!�"OD�@�틃>m:��#�w��\��"O�y�Ɗ�n���!"�}��13"Ox���A���MZbA��qx��R�"OV��b<7$�H!" ���a��"O����H�� !��U�J��"O�(�����,TT ޠ4w2��6"O0��#�Ǭ'��}xu�Wk��"O4�*�[�
�x��M\1Qa0F"O:ujc����U����B^����"O��ٷ��n�0�`�ݭ>��1�c"O6�jU)W(�X���G�<8���hp"O�9�ăD-tl�4g�~|Ψ�Q"Ol�ydo��M�He
�#�����"OxWI�:�H�!�r�(��"O9(��^� a����6n*�8"O���hQzOف,V��r7"OL�;ŏPf�)X��V3I0���g"ON�9��Dz�����A͝��c"O��e�&3>��°�4!	����"O�)gK� d
�,C��3���Q"ObD0��1fz^�J�o��h��"O�Mrr��&C�Z�;��w�@�"�"O��a���Te���7�*#�@��`"Ov�;��G�6���p5.����"O���0�`��B�ML�"Oj8�rj�4z*�YA�bP�^�����"Oh��6�A3 �a��%RU�=� "O���@�vrfMȱb��3�l�4"O��%',���7!��W^�홐"O2���+c�2=R���{ft�"Ob����2W�� � DƘ��"O�q��◇K�y
�o��;�V�j�"OҨ�"��*j@�Ԋ�F=\|���t"O�l�d�ߐb �i0o�ǮLQD"O�YQ�
�u �+�p�l3�"O��1�O^l�y��_4��!�T"OF�H�k�*�25�,�@u�s"O"\A��-��,z�&��:�yb8Ǝd �GN��Ҁ$^�yҁP�Fa�I�)A�q����P��yB�M�Z
�*�+H�"�
����yb��fv.@s�
U�>���G/G5�yRCK�A�:��S�
#o�4];��ȓwa���r��Z����`�ѳ&��Ň�5\��_�6�$��Z�� �ȓsc��Yw�^�K��X�ǉ5!�
4�ȓ������=F �t(�� HF��ȓG��DI$֫\�tXw(ݓ�0�ȓ%��ꕄ�U�VP��U�z`bć�b80<�0�>bu��[���D����ȓ	yTQ��E��]�!ÕW�|��j9Td�V#�.I�{�����݆ȓ^<���ъ:�*mJ$�"rxe��bpT�t�UJM�d�;j��I�ȓv�4]�e��w^�D��7$�l)�ȓgnH�� N�xl
E��N^*U�����9�k
G��U$�|Rل�3}Z5�T"��g*�#C��w�b@�ȓF�@�C�ÍX�~pc���1n�݄�A ��%%޷-�|h�䣟�2 Ԅȓ�`1�6O�4zt�!�ǧER����S�? "dy��Ѐs�v� ˗$! ;�"O�T��'��h��)��2$PPr"OT��W��(N�,�lB�0�
 "OZI��(+b���+����K*0��"O��Qe�ˉ�����Q+j^��"O�ۖ���$�0�!ي:jR4��"O�5���W+d\����rR�:d"OfT�$���%<d\A��P�]�"Of��!^W���C(ك
Q�8�`"O��u.(����F�EV�1�"O��۱�LI�Ā���]�8>�T��"O D���Ҟ ��eQ�IO14@x�"O�m`G�Z%G�� ��73�UY�"O�!nFWsvd���8J02Q�C"O��:��ݽ6�^� �mD=&}�2"O��C��0�d0��JZ0j�5��"O ���	�19���@�гR>�b�"ON���'��2����H�)
!�dS
V�B=�����L�d�$t�!�P�c	�|�h���$K���!򤞷?a���)6�Nyz�J��!�$H>4Z����	6.d0D��!�D^��� ��J^;6��%�J/!�dX,=� M1�NU&( M���7 !�$�("���R	�b)�����|!��<p�H3����d<�5�5	�!�$�35�v=��B����h��.#*!�#��ŦT�~A��h�>�V�t"O͓���;#n�DQs-��Q��"O�0�R��+��B���%d�B�!�"O|)���Z"���qǔN��TBe"O�A��B���ʌ�� �~�bI�"O����h�G{�i�W�Д]��H$"OU�p٠W �Yb �"o�r�:�"O,IH���:�8am�!X��`3t"O|�
���>x��<)���a@^YZ&"O�r�Dɓ�>51��܀��05"O,�P��z�\��,��0]\�CP"OШ�n�9��3n�1&�R��"Of\zhE0d0��&��:8�8��"O�[�"I5Xċe���A0����"O΅�U�N����χ~*X9��"O���woC*r�6Ɗ,7�D��"OTe:����Z$� ;׈ʉ	�A��"O�R&�އ.� �a(��#(���"O�A��	\D��%s�	�w
�š2"O,���J�<��@�O�pũV"O��L*T��)��H�N���t"O��:�,�Q�l%� 쏛qVĔ��"O��2G+��[�H1�3kS�D@n�J�"Or�(E�12`5qvJ�X3�t� "O�\뵉Z_���I#{���a"O�9��)P��abj�2 ��s�"O�׏֪s`Jh�t.ė �X�Y�"O�4v�?,�p��e�$�P�i*O"��5j�%!�(
",�Yz�'#��9d���% �F˖�$I�'Ͱ�@��в'�
=  L�Hm��'e�\�0��]�j
� ɬ�z
�'� ���eѬ|��YSC%M!���	�'������rv��A���9%�@�'I@�nϓ!� `�R��.��h�'8�ш��3C ��6�U�x}
!��'JjH�t-�1b�iW����� h$r -I4'�(
�産*��}��"O����W<ws�	:�ŕ�V��"Oj�{Q�؄}�Z@�;[h����"O�|��Y'zm�է^MHF=s�"O*��
�}���s��I��y��"O�5�E�)�<��F,�� ��8�"Ot�� o( i���(l�E{�"OJ�b��ע3�Ɛ(�%[c����"O���MT$���C% p鎸qP"O�$:���e��A3�܈*���"O�9I�R.R��F�gu��9�"O��p��)rǠ����\M�XR"O����I,%��+��`e�=��"O�Y3�C�,�(5���9Z��"Ov�{�Q�R�:�k�"�*�
=@�"O��8�"P�,�(oO��]>H�B"Om[�Ò�i��@ փ8�m�D"O�a��
m��y�W���3�^��d"O�0s`f�R��XZ�ٙ �8(kp"O���Lɒ&�ɉ�L'��H"O���_	U��A�e�E=A9�"O����+>�MH`�&V,x�t"O�1�W��ND����ɩ�@T�v"O
��j��vόX���.��\��y�Dz�x	I�Dk�p�T�-�y���:}h$����?ؒP0#��yB�=v<&��6��/ٸ48b#�yr�ŋ=� y	B��/��걩
?�y2��K��;��߳f�J�Pv%R�y")��f�D e�z����y�B�Z�PԱ4o�-RQ��+���y"�)Du��%������jH��y�� Q�:9�3FU*Lϸq)u��y���H��(_�3�����y2č�>�j�_Z\ȴ�"ː�y�GUj�*%��E_�M1���d��yRI$S�2�!�؍O�nE�6��PyBΛ���PF�	vRR�a'�\�<�gH�e��݋��%�B<���|�<�"o��s��D�
'qt>y���o�<9�ٗCW�1��T!K�
=CT��O�<�T�Gf�GEՠ���V��_�<!��F���������B�l�Y�<y��?Ǝ���u�abei�R�<���V;:X�4*�i�*@�sD�<'燝U�����1frFp�r	@�<iW$�
2����#�J�z`:�(}�<�aLN�e�HE���D &�ER�fWu�<J�L����FB�.�0B�o�<�$�íf�*�r�ºA�����@Hi�<���[�$n�q����y�T���]f�<���*7�E��f��n�p�b�&�`�<9")�$	<0`I�ςtP���l�Z�<��F�3<��Is��=T��y�m�V�<	p��K�$%��
()	0�pE�R�<�`eM�!���2�%+��-�D�M�<���qd�u�&A�)6�IJ ��n�<E�^�H��}�,@%Si����Mr�<�q�$Q4f}x�)� Ɋ| GGr�<�G�ծ�Lcu�@ ��Ԁ�y�<��A(��3%
^Tg����+�|�<Qd�{]�(��G��y���@d�<	b�ؙh�kP�@� A�S�]�<q! /O�HPK!�,�qQJ]�<� �����D
Xe�s��tLҼ��"O��馆4E��0�1�P�b��i��"Ox���D(�l��ڭL���� "O��ȡ���	I�P��b��3��*�"O��B���9� ����M��]��"Ot�8�^�	��j�J�i�ĉ�"OҌul�l{ pM��*�jMh�"O((�EjV%D� Q �F;_�dqt"OVXd$�t���{��;��Q�d"OJ�0��6Q�X�d�w�ެ�C"O��&fۦW��h*��4|�|�[�"O��& �1�F�k2��#0�2�"O�X��Θ-�0��A��x\A�"O��i����XW��3�aD�B��Yʴ"Obu�WB��L���q�t��"OV��0��'"F��q�6Xl��Ku"O>�PB(�A�0�`b$g.bU�"OHuSBD3%�L:sޒ�Ś�"Oڜ�u-�?jc~(����`6-2D�0�2
�u��M��"֥W� A&i.D�h!ʳ.� ���oI4w_&��&�1D�dp啑>�4��r�9@	�P��$0D��V��aղ�3ׄI"�|Ċg�,D���q�H����UH�1�8-s#=D����
5
�:R&��Y'���:D���ul@%b�z��4�j�e
7D�|:�c����3M,�$ �2D���*m����.Qخ���/D��W��z���ZՃ�_�`	�G�.D�L�1g�2Vx�3a׻7r>�h$�'D��a�ؑ8�N�JpmV+����D'D� ��K�,A��|J%�S�x�>i9T�$D��BS+j�
Ur��R)[���j&�!D�`#�L�|�����>����!D�,(T`ڰ;�yW�Ut,���=D����I�es*��Vm 1�0��P�1D��ȗ�K)����C�v����q�-D�H���2�,���M�pڕ3w"*D�@���!C>��ƸD��MR!-$D�P�FAW����c�"�Vf����N,D�p���*]4)2��?mi|��L*D�����p�r��" R�M�*XB� ;D�H�@���xvN�B�Eʍ$��D�p�9D��T@Ɩu�l!�ƴ!�hyf�7D��x�
#*�q(�,_]VxiE6D��AC�	�lR��d �4t��4D�Lz�`���x���)D�2�p@)1D�4:�K,��h�e,.H{N�v@$D�dJp�W6r���p҇1�r��)"D�����E3!q�e��C�d�:@!��?D�@���2�Nt�5��X�R%)�j<D�Rs�
=/��l���,c����5D�,ɂ����5Y��9F24�k��1D�0�eG�0~�,���
8�Vt��+D�D�6�Ѿ�1�Q��6~cnx+&�.D�8	#��J�򱳦��Gފ���E7D�ذ��ȳ`��t@�Ҙ<@Z89��)D��rר�E���o�7fDP�06�#D��zDh��:E�a@�0
��I��6D��Rw�^�P����2)W�.+�M�5�6D�, ��#<�I[%l_47�\� ��*D�����,Dx��ް=��xjB�'D�<��/�50ݨ��F��,�����`&D� ���?,<H!�*~�ܪ��)D�� `��
;P��ꔌ�#M��r"O���q�%G����2K�76�Zd"OB T&��Qf�9���=z*�X��"OV�G�N��N$Y���2��s"O�QYӊՏ��@B�[-?�|�@5"O��I%�(<�0p���
CT�)�"O���eY�r������	�"3h@�#"O��	��&P01� �X��)b"O�h�/,\`�Aք@|�YC"O: ��E,W���0$�K�$��"O8�"�H22��irEY�W\��3"O����\�b.�U1"��"3����z�![�eHs�`��ôk�Y�ȓlV
9��U8g�V�1j95SH�� 4�l��*�$|���hf��*-ܜ@��XHx���P�P,��FX�ȓ8I�����M�x�Tx��H��W\<���,�r n2xI0��۲B%�]�ȓ!�,����؀v|�P�r���z�4ͅ�&���?���Wŝ�I����ȓ8�X�p QgdlC�@�$|@:��Cz	B��ζK�Ή���D���ȓ��})����2A{�݂2"����4�tsd��XU����3]���ȓ�p�i1+H;�0��  D`z��ȓ,ѤX3w!,eªQi�d�6R�h��̨Q�s��PoF��M�;F���8k��j�D,��X8d�NX�lE�ȓ	��1ѧ��o��Y���� ���ȓi@��Ĥ�D����#	�PS���� er�p���ͺIXpG٩u�RC剓Ci �ir��&n�M����J'�B��;U`xmY��e�Z�!S�Z�B�	t x$���;q��)�d.ϯX��B�Ʌr>6��	� �P���K�&ׄB�	�Z����Ġ�4��%I�Jx�B�	�]��kt�s!���*�~���%D���V	[�>�*���iP9y�B��".D��(6�؟y�]���3n���O,D�D(�� 6c� I�f�!����D+D���sH!J~ 4MK,v��ѠB)D�P�ᅂu�H�"�G�\�NZ$�;D�@�V�����1q�b.eu0��5�9D�|��B,-b69("��.,Y�07�5D��2��Pu�*�B�G�{���go&D�� 5
Y�I4��5W���0D�)�ɍ6�$�0����X�@�j)D��R�O850K$�L�ʶy(c�(D�T(�
�z��΄�z����Ш&D��)��%l��� �_�Ԑ���"D�(��O�:34hRr�T�����6D���`/�g�L��r�H۵�9D���U�J�V:��C�W�3)��0B�;D��!��eD����т48�	1�:D��� ��I8"�SĎ4:9��R�9D�,� ���zb���4�߀%��Yj4
4D�����Ps���9*��#p�8�T�-D�$�E(��iW��B�O�\G��cF�,D�tY!LVm���\+�:�sV�%D�p�`Uh���q�l��z���׫?D�x�b�5�|0�E0��U0%�<D�X�aR4��rs�lv�!3�#=D��2EHI)p�
P)�`Ď}�f�2Sj9D���RM�s���Y�(F�e�Z2@�2D�� *鰵��+���`B�<(�Ȩ�"O��S��F1C�e×3&�"#"O�`�4o�3B���I�.P�&�D!#"O. 9Q�K ��ͳp�ϡQ��{�"OZ��&�H�6�4��k��[
�P�G"O"� �3r`80�)L�6H!"O����\�w� 4�v�ƙO�1��"O�@��)Ҽ|�W�כ2�b"O��{�#8�>�c�i_y�|�Z�"O Qbf3���U	K�'�@�R"O��ɇc�0��=����{Ղ�X�"O��F��a�޽�Fg^!�Ђ"O�yY!��6Q�^�AF�*	��)�"Op�S���=v��mR�>I$|T�6"O�$;���P��):Qwh8@"O���%J�3��X�B��au�8ȅ"Oj�Y㇈�2D��i��R	��e*�"O�y���ѣ#�=r�?? ��"O�"�d�Z��d T0J�8��"Or� 1W ���8
�j�"O8��H�5Q~�pA�����k�"O��#�}ʥ��M�=,���u"O�(Ⰵ�)
���� O;�-
s"Or�֪�8�8�R��m	w"O�`��"ڿ�XQ��&�
�X�"O6}�w �;��κ<?�$��"O
�"��?\	�VŃ�C\�X#"O�M0�i_�1~�qR&%�v�R�"O�@C�F�M�M�"%�<mP�D8�"O��&_\H���T��H�"Oµ�FLЇ"x i@���*<��"O|�����4T?�� �+KcQ"O~Y�G�[-t��e��Ն5���g"O.�0�Ր]��Q�Ї�.e�d(�&"O�-�4-�n|�l*�	-B� 4e"OD��	���� ���P�r�[�"Oݑ� ��(,�ʐ"@�h�T8�b"O�pᥣ�6�HQڣ��}���F"O������b�
�[`̐v�Ш��"Oȥ`aK�������1?��"O
q����6E���y�C��x�F�R"Od�S"Jb�V��CT?����R"O�4I�1N�85B�b��mh�i�G"O��3A^�Z�LP���^�aT���@"O��bP�2`�Q��G�!;ju��"O��f�ha����f֧	�Qh"O��#��Z�.5zƧ�5|^ d��"O�la��D65����B�7LDy�"OF��k��diA�Ģ9�u@"O.؃�MV�N*ء�	<$���"O����E�0Y�~�p��O�/&У"O�a)�A�)|д2�Q\ȼ	�C"O�M1�j�6Y��L�+5��I{5"O,IZ0hȧHN�����1!��۳"O�U��	l��a+�� Z�r�s0"O��ŤN�'��1�U�>��QP�"O\� ���ݨ��X�g�8�$"O�(��׋�jh���S�f��`�"O$���+t� �G$f�l�S"O�q�ț#�f�2`"�$.h(li"O�9!d k�Xs W0!�����"O&4{���o�n�qT��0g~�P�"O��eǁ�4�P���g|ĭ��"O8caD�?F��T�5��5M�� 7"O� *��&j��`��T��M�=M��A�g"O�вs�X0h$���L�;Ό9�7"O�����}��8�cl�����"OV}�`C�b��Ċ�đ�o���z"O"!��.�/&���h��ڠ(�+��O�<9��ʬ�Iق�Ȼ+�����G�<��B�;w��ъ$슻j��}	V��]�<9U��(5V R��:4����E��\�<a���# p�3���Q(��Z�<��DL4��%`Įn�jyഀ�K�<)��r��4���̤O�	�FƋF�<)����hlI�$/C�z����Þ\�<��n(k�TI��(S�q\bEX��Gp�<y �Oc����$M�6�Y ��h�<��Ѷ �:h�gD�p~P�5��N�<qGf�<g F�A�X�:�`�X��L�<�`�� K��aDc�<( ��G�<	��A�mHa;�癣d��p@���C�<	4�@�Kh��D��~\��F�S�<�b��
�HаQMpu�牌L�<	2�^�'E8����)�ư��`�H�<i�'�A�v8�F�;���k�n{�<�E,��4���$&��%5, �"�y�<2�ȄQ-�bE`U�L�,��E�_]�<aSj��5�d�Ł�i]>�uG�q�<1'��� ��U��`1ፂB�<�p�_�K�BQ[֠�e�9��FG�<��B�%]Zd��C©D�ޅ �`�A�<Y3��p�����.[�MJ �,_��C�I���hSj\O�x����0.8�C�	5��J ��-pfY���7.�B�	2!��]:R�^��$��d�)2f�C�ɴy�v����%I���!)�7i!dC�	B+J���Ɣn�@�1�a-&C�I8"PaP.�#.X��$
=*�^B�	�j��1�"bڶjW���ʄR�XB䉯��U����X����]�DB�	��@���Br�((5O�,��C��*_�n�R��`� �����[ZB� gf2T@WKΐ[��T8�́�.�dC��9U�"��0#¼z���MA�h�C�3K��\��q�>���ޞ�$C�=�j�#��*�E���v~ZB�I������BRY����.dC*B䉰:�����O�U��х����.B��+�H�zs!а3.�5���)��C�	�$b�]����(\��袩��y_�C�ɛo����H�uv�s�@�++�.C�I�k.��0"�٤fw��c�靨/�B�.SiB��Ϸv�Ф��h<CA�B䉧!#� 8f�<IE��(���'E�B�	 ��@̀8w���T�R��B�	����'�K F �����jǚB��'<���Н,�0���IҾ'r�B�	�[��V���`u�1�΄lGVB�	3	|%����7P\�0C��<H�.B�I�j.�8g�-<�f5+ǌ#:��C�	Ur��c�2A@>q�'J�v�C�I+G�}�,��y�2٢�(]��C�ɾo�p��AK?X�0튅,�&"[ B�I5]�yТ��Q����! 'k�B�ɰZ'�� 
��d�xx1,R {�bB�I;�\1��	�M����am-K�>B�	�Ь�Bg��/l]��@w&ڗbw
B�)� �%hDL�20�l-�p�Y�*�R:1"Ox��6���D&]1�� �j	HE"O�q4���H��L��*R�3�(i�A"O2u�O"�drJ��]�22�"OfUy
�+4G�M��&�&HȆ��"O�t��j		+� Pa%Y*��͋"O�iq�!C�L,�rPE�
��R�"Or �'�^�<-KW%�2� S�"O�eYpi:��[F��^�څa�"O�l���� ;�uz��"Od=��B�oږ`r�
D#:WH��yr�^7$��iĕO��Ġ�eȬ�yR���Is�� � _�U��͖�y�ᅥP3>ТE�E�(%�-���V��yrT,�X�����7/DĀ�k�y��0.�@D��R&/N��$�$�y��D��"Qk�
�0��@jU%Q�y�K��h�z#	�'\���������y�k�2,�`�@:�l9x4Ş��y���e�T�∬q�x��>�y���7:2ht�ԥ�%e( �2��.D�da��Y6e�H� �I aE�9�R'D��)B�ǧX�F	KF,�,�h�PE�!D�P����MN@���ʄ5g�����F<D� �C�h�H����Q�
V�6D���#+�~��T��Č�j�1��4D��T�ȝe�j��A�Sc*�;t�3D���G�^_zd2�)]"X6�S�5D��!!��(_P��9x�y*�4D�4I��	8>̅�rm�~���J0D��K�#*�~�@���"�~x�%,D��*��r�~xp蝭$�F�O?D�(�c�N>T��gG��a�$��4�=D�ܢ`	KdAP�fC�3�Nd� �6D�<p��O�!���u�@�;��)�6D�tӴ�5~ĻF�Ea~b"+3D����;d.�ʃ\�l܀�"2D���B��7%\�xt�5*-!��*D�t
�K&	Ά%)B��9��H
��5D��9�a�'<ڐA�װP �AzF�(D��� Ϙ��|��b԰;��Q��4D�l���.Z�(0� �,$E�}�'2D��#�*ǽf�v���O��Z�K��:D�ȃe�(�	�L�n�4{�*#D�4*�➀B�J�c ��pa�U#!D��R!�D<}ך	�׏�� �DY�p
;D��:�k�1�D��d�X9�Py��4D��vH��D����X/Y�����3D��B�jĶ(,��GדJ��	���0D��閭� {�0	*�$<��$�,D�؃3��(�(q"D���I�l��&h%D�\��)V�`,9�@N$P�B2�8D�kFe��'�䉲�Qa`W�!�d4O�"g�U�Oe\(jV%�|�!�$�k���ؗI��X>��ʤ%!�D&'h� *W�4ѧE�;!��,���ۗ�/>�4x�DdV�i�!��mF��Ҏ�so��{עB�*�!��D�tY"V*��F�D���5�!򄐐
�v` ��),$$�D�8&�!�4)q�`2�ۗ� #�,�,W�!��w'���	��8y�]�!���N��QB�$�L0��߫v�!�d�;H��5	{L��@�.}Q!�� � �aK� ~�˶����b"O�����/1�EA0\�* @�"O0h��]�$�ʣ�VYd�Y�"O9��@�`�<���lF��Q"Ođ�&�ձ)� �J�'X$/���U"Ovq��E���a��C����x3"Oj,����B.꼺��ԏM��D �"O�(B4�Gܖ\!ϙ��p�ٱ"O�eK%��>1`��-��c*�2�"O4H���W'
�&��e�΃pp�Y�"Ox�r+�bn��GG�7�Fx	�"Ov$O��@Q�8��G �ܱ�`"O�"���c
0���J<�2"OƔ�Ʃ_�J}�#BZ�*�ً�"O�c7K�������ٗ^��1��"O0|�$��;���
%��VЮpha"O��qU'��Y�L�E�F�M��80"O�d���/6�����:6�*�� "O���п:��X��"�/8��P��"O�� ��^�d�	�̍_ ���"OQr���0���Ə(u��	�v"Oz��P�EJ�u�p�	VWPi��"O�bF�LP6��O���-B�"Or����$��tC�F�Z�)R"O1����<h���"�Q�A�PB�"O�l���(m�h���^9���C�"O��I&�����$2�߽��X9�"Ol!�U*$�@�aռ4�.��"O
|#j=<� JC��I��ɧ"O����%�)Q̸Qr� ;sU��QR"O|U�gͺC<\Y�dO�p���@""O��y�"��-`��x�G�3;(�(�"O���3�¼���I���(RC4H�'"O M g��3>3�b�.ٷ�.�k#"O���  R�E��<�G�Y'8�^�%"OhL����]� -�q��2�|�"O�����w�h��#ޒk�,�(T"O^���;=rc�1���c�"Oԣc�yI��S� ���P��՚�y�
W�D�|b�狞t�T,s�BJ'�y�E(2� ����t9x0u�X��y��
D:ܜ�
Qh���4�<�y�˒�v8Yʷ��Vy�1z�c��y2F�yjX#@��cȖ	��L��y��U��*��-λr�(ɘbO	�y�늴AJ��b����	S͌��y�C96H��e��2zP:�92O�y�����A�r��%	�y7@֬�ya�
�]� _�G�4&h��yr��8s�.�	���CF<�(�,��y� �� g�-�R��<!
}@�mA'�yB�U�o�P�@!�0��h��C�
�yr��3x���� 3-����t�W��y��	�$/r�2!h�+2����V��y���:v�� �`��$��i�����y�o����C ��:!@kd�ԑ�yB,�,�x�teH�zn�S���yB�9�ZA���:��Urc�%�y��<�ލI�F�S���Р�"�y��T�M�ir eJ/���G����y2�\�{�.M���ǰ
~�Ё�	�y,5�F�aլ?z h�I�C�y��EC�N	y�c���E�ЀƑ�y�&Ȣp�X��S�[�*,Y���y
� �ѫ#�5A��
���.`Eh�"ǪA����3B�(#-]k�Y��"Oh�����u��H%���!Ӯp81"O*��b��쵠��J�P�"Oތ�7�7fP��̉6�\�!q"O���`�µP��Aq���-/N�Y@"OE��ʷM���ˑ�G�8��E
7"Oإ��Bܮt��(#�ޑ�"O�x)�IJ;ș�a���8�5"O�D{��pJ��a�*O��,+1"OT��"ƕ�`f�t��b@#*M��"O��Vf6B��-
d�.���"O��QsiY�xخd0�d��T�ڃ"O�Ś`Ɔ�9�aJu��8@ `�"O���f�ݛ�#P�&��(�"O�2E�M�4�d� �OW(d"O�,����k�(�K���H��H&"O|=��-ه[��Ap���z�>`�"Oܔ�$��bmtiG	ɸ�M`u"O���W�J�Ѹ �Ùa�Ʌ"OT �B�>���(L�)��Y�"O\dv�Q�<&�b�_v�X+w"O$����rϜ���gY�.��W"O���(�C�p´$�8-����G"O|�r�#�3s�鱀$�%r���S�"O��ͥ;.$�K��P<w�Z�#�"O���@�$D���!�J�U��3"O�t+dG��� ����EtDj�"O�T�P��`Dj�0�$x���q�"O�h:�(�1o�.p!f*�#D��$�w"O.����73널��OȻ�F��q"OXmxE�Z!oO��³�9�lyҖ"Oʤ�$k��e#���!zf���"O���4�.J�� �c��<M�T�"O�D9t�ʪ:d�!��("�Z6"O�11ǎI�ix�p.��a� �"O2���O�8d�
���rpx�"O@M�&���{�D9�,��$��pH6"O�x+'�ɵrQ�@B�D6N�D	A�"O�ykW���n��R�S(zƾ|��"O�M��#u�����,w�<Q"O�p��'��-�9*���"�"O0�1AÚ��i�* 3-@��r"O�D*W&��!
�	@ɝ�pw��ۅ"O�(�6�IXdY�g��\��!"OA[$ ٘��ԣ��N�E�h4h5"O�i�F����3w*�s�h(3�"O�����E�<�E����L��*"Oҩs��� S� z��I��z b"O֝k�,]�H�����,�7�PЉ"OވЕ�!t8�)���ȗK����"OX��`K�i���r��y��t�"O�|"�C<'0�<�d�V<Q�Ne�"O`q�r�
 ���q��@��B"O��r�cԚ
J���\�4b]�"O�5+�,F�<����hS�H��"O�����.FR�I� �o�ޕ��"O��3�i�d����@n�C�2 2�"O꓃M��R���E���"O��YG 	
;�`{楝�Z�0"O���P�m:DX�7P��  S"O��B��Q�'CB>g�@�s"O��H"��	{R@#@TF��"Op��ѠʭZ[�툥/O���H�"O� X��@����$���/0,�	�V"O�p�UG�!y���6�Xh"Ot-��]�%��Q��
�u\���"O��8�c��?J��)D��*��1�$"Ot��b�_�x��@B��A�a "O*�Y�K	��,a�T�3�U(�"Ox�� #9!����{Vnm��"OX;�*gрj,�F`dZ2"OĉHB뇔$SjI�H�O�����"O��b��RY�*�5E��/�LY�"Op�"���d���p3�T2�nȚC"OT�R���e�*D"���(*�*E"O�'$�w���C(W켌"6"Oz��r����@bT�Y�b�A�"O�����CQ��h�)D��1�"OlLy�AܷfV�(37!�<B�"x��"Ol��0
U�u��O]a�0���"O���R���B��1� ƃ]�N�"O��i�-2�� �m��<1��"O������&nɌ`����-k�XE	�"O��9�KI�"dġ�)��A�9b"O@rPh����!�ʥDuF��"Oz�i��]�3�,����ԐOw��0 "O*����ѬP|����!eؐ�V"O6���K[%Kvt�Fn��z|�k0"O��9EΕ�,xpal[���q"O�Y�s���0��8�FB˭	��r"O��H�� $:�H�(U�Eq.�)"�"O����d��P� ��1,3( zQ���s���	�[>�ɢ��'��)�q�J�-�O�<
 ��8! �P �&���"Od���5z����s�)��9rO��d�l�C� �"{&�P�KT�,�!� 4z8T`��5 Y�vҫ	�8݆�U�ʽJ�T������M�މ�ȓa�P�&"^�I(��Ă�Ŗ�ȓ�@��@����B���-1���'��5�$���~$���_���a������	�Z�X#K(6 j�	Cnŵt��B�	%ST�sУÈJiXA�֪H~C䉢* Qr)N2�B�����29��(*	�',H-�QhY�ž���$Յ{�eX
�'��!�l׼Q�p���O�0r�ΐc	�'�p�ӈ�%Ai,mY0� �5]a	�'f�Ye.�q ��w$�"v�I��'n�P�ug�2)�]FM�u���C�'b���=m��6_��p���O2˓�~��$F�T�y�d��ԁA#9����3�ɩ�y�o�?+�ܭ��U4s���N]>��'��' >ի��5�=K��1a��� *LOH�'L�$�O�:�B�� �qw^$i��84��܄㉼XN
�X��A�ZIڴbi͢yW2�>���Iب`���X Kэ^RZИF�+!�䝤-�nd;�I5q���1%�<6��$.}��>%>O ��&������f��9G���'1�	7f���2��&���P�����6mw�y	�������>r(�ug��{�����@�S��`��W��|�DcF�%w����*� �Q�t��P�ȷSl`+��������d��x1���Ҕ=�����!�$O�|3����&β���R�!�d��O.��B���ɂ��y!�R�e@��x�&��z��J��<j!�d�+g=���%�K��5qg��"gi!�� ��e�H�{r1�a�9!d4�"O�qAC���7*���Wc7��Y�"OF�!��H�q�a���0I4��"O�HP��P�g���7��@A2� �"O\a@�c�cD9s���zEh��"O�qh�nI��,�y�ދy9\Zw"O ��!B�*�����/v�@"O^(�w�$k��ě�i�J��1O
�=E��cæN � :�&_3K��SѪ���y,N�,1Ԭ1ը^�+.NuA ���yJ��S��!��E���H�g��>�<���D�1Att����&J��1�f���Kb!�ߦ2�>�CZ9��Y ��_��|��i����gG��s~0 �%C�V!X��I��X�Iܟ,�E^	1z&����ӥ#���s� '����{B�)�	g����CI5���k4c�7>�!�d���#�I0�֝�"G-R�!򤖨7E -�D��(�LDsfB.N�!�سa�bu�*�.�ZQOU�!��_X�� ���{�"t�B��\�!�@1 ��S��E�;�@��O�$;G!��	3�R���EƝ�ԉ���TB�I����;LO���C�S�z��lح8�PiV"Or��Dœ���-��-E�"�R3"O �C^	�(�ċK�M�� K�D����Ӛq������8^�["�ݰ4�>B䉴j��!*��l+�МV�B�I rtI��N����r!�J:��c��D{J|JG��q	2�*b��#H@i1rc8�~��'�FM�0+�u	�l�b��$����'	 	J҈ϗ5��UkR�Jjbz�'Wb&O�qY2)����&T���͋�֘'$r�$!��B(]0��#I�1$L��K#�!���{'��cc�0w�qz��΃�!��R]������hj U���˓X�!�������Cmצ\|ZE2E�ݝLC�J�����7te�1D�B��vB�ɡ'� � �H��_-?�:B�	�B;$��!�@�p�ȄB��G�H?b�d���`����UCN8V�8��Eۚx��C�I=uB%8��|l�d��V<ܪC�I3i@�E�Ւx�v�F� h��C�k>쨨Dd_#|yv0�ᑲ9�C䉀 �H2��L�x!R��M�)�ƨ�`�)��<їd��p4���#��xSh�	�H�y�<Y�N<�ht"ga�P�AB�s~��'N]��?-�̭�ҀѪOJ4I�'��,+eA��Jd�P�)��X\�	�'�ṭ�U�V���;AΘ~�f̫듸�=>=Z4�N$$�2(("+�%�C�ɩob|h[�)E(a� t�&E>�|C�	9Fv���L<U�q�V��C�>������B�==Pp{���?gZ؄F{���ʓ�~"�'�v�hN�iNp�@Ϟ]�Ε�rO�ubr��uy�!��j��,���
���;�S�Iٖ/�8����fn�-JъE�a~�^�(��B5W!L��� xO�� �1ғ�p<�!�ۺ.�|<q�ʙB���6	�U�<����*Q�I��ᙙ (UCW�B˦Yz�,�(�����3NcX���
�46�����'��)F��-3J��#j_�YŮX`�	5$�T�uCC�2�j�T/ǔb��¤�.�R�R�񄇓��@bE�O�})q�lɊ0j!��]�Bk0q��
�9�^��Q+"p!�� �`� 3k҄��G_�����"O�|P׋٫B����c%\'io��;'"O���)9r�#��D5?n��{�Z����T�'�Xq2Ԍ5*��$��18h���'T�l;�d]�`f��ZE�W&.^�y�O��=E�TnM�G+t��$[��0�!����'�~ ���������Y�O�3S���+B���y��Or�"~b�(R�	ì)K�m���!0t�WG�<�d���8���an��;���F��<�ϓ� �p�U�^���*йNO����	�<��(y̜#F�ӥ'�r�BT鐰��x"�־f�q�B@�BtBkt͍���On���iԘ	��С�cI�N��Qy��ܟT�1Oh�=�O����A���A�*?�j��E^��!��b� t9���^�m�C&��2�!��"L˞|�#��5wP��Ґ���(�� Y�8*7�1o$���W(��il��'���iy|�^��C"�:}����Dk�);�L,D�L�m�7pexE�E��>t+��)D�ܚw爢 %���!i24d;%�3D��Y�JL;g�uhq�ug|�F��<��5�ڤi����4i!�;Nz���s�'�����H
�j��As�#�����'/v`��*+Ql���e/����'�����G����D�)d��'h���E��6�ͪW@ۆ%@�š�"O���fμn]fq�Aώ1P�d��"O�ԙ���D����2-c$1J�"O��H"���WY�/]�:sz ��"O��*E�<g{��I��ӿnm�b%"Op�Ǜ�XP��u��2rT�@��"OB�hMU
����J˕e_(U��"O��³�
�c��,xf(R�Ub3�"OF-�H:h�8)�@�L?8Ha�"O��ŏʰ#�dŚ�B��1�,��3"O� +�c:]�� 5]�"��\��"O(<i4�F��f@��@�V�<pc"O�ZA�-`��d*IfSjԺE"O,����5�L!W���Z8 �!�d�D0t�Y�D�hp���W<)�!�[�q(R��C��'Hc����#C�!��w�p��)I�7��I� _�w�!��_4n�l� `\�p��Tk��c�!��ٓ0n���焠K���D�7*�!�D�g�(�F �"6i4��gfܶP!�$Jx@t�� O5\b@���J�!k!�$ tm����(^� �<1q��?Oj!�䇴G'�u�$LR�i�B*a�Cy!�D�
�pLR���@�$�+��ξdv!���7Cr��Zv�R�#���8���8Y!�$^�+��1�F��e�`1��"�:�!��j��𡋊�Sj�`3q'C�>7!�$��(���M�m?H�2Q�Q0{ !�Εs).5��&F�I&�J�k_�q�!��͚1V��_�};�h;��1D�!�D�iȼ$�)ׅ$
��QkE%F�!�ִ ��d�򏋫V�nP�֧ø!�!�U�6�ŠCY)_�u�'�%�!�B=�Zm!χ�O������fy!�DB�#�0��qI�>�������J^!��0� ��]�	�s��AE!��L�\d�hj���X�Dd��.�fP�X��H%Qa~2��
�ׇ,���z�E��y��Da����CN�&�֌Z�� �y
� �m�fjԻ[�H�6i֒3�*�z�"O�E2%,H,z�d�x�q�F���"O �4Ԣ{������V)�.e�"O�kBi[Kh���.[>W^� �7"Onq�D	5�`�0s̀<P6�M�"OZ��b�.v1�� ��E�j��3�"O
����Y�?�\̓U�vVL%Y#"O�[��%ԦγmLF}�Ԉ0D������<�#� �r��a/D�D�e%Ә*��p��ř��y �%1D�����f�D�w�V�>ﶉ��.D��+�a1:�!�"�U�X�U�6N-D�D�o�7hp��Ff�
\ق)ؔ�+T�H:��\X_ư��m�x��Q��"O���+�ТB؜�B�[�"O�ȈQ&�����ЛIW��B"O��R���|C^��տY@.}1�"O��9'�&o~ BtfߛGjl��"Olu@R
�V���(������V��^��y#�'	��zCh�ZN5X��D)`�bq��@��6�D��	�F�rv�ә=��b7%Q?�Rlp��ˡ��	����O���)g�;(���'�蝈������Yg/W����"��~�L��gbʐF"T�Ū?��$�a	��^It╠\�"�J�����`@oՐE&�	h�'/�D��	E�e�h�)&��	�qF{҉K$�>yZa�*i���;f��ɄB�x�ʗcجXc���k\�B$d��}8�Dإ_��� ��L>1���;�J!PR��!	�pQRP[���h�c�O��Da,N�@s��(�\�XWAQ%G�P,����:=,�P��	'u2�� z�����Yb�ȁ�	�w��Ș��4�t	c1WܔDPw)L��y#h�|±M�v����!@�4�n);�Q���"6\�z$
�jR*R-lO����)I��!��@�.�h(pG[�	�t�t��K���A��� {��p� &J��%�$i1h���Ol�D�>�TBO"'��u�P1j�L��`�P;!�2-bR��A�	; �81"���_>5��hս��+bHS�?���A��v�1���b�Rx��%��o�iР Gߟ49�Ʌ�oQH�ӄp�)��Ǔb��e|� ��e��n{bK�%0��Y�ǌ�zV�4�񡇳#��% �CYa{�,������0iŌ����q����0�B�)�S�b��-�<�t2A�ï���D�bH���$Iż5�*Ih���}����cS�&�N��/��T-��o]J9"y��)��mD �l�//�8Y� �F� A�����Y����B��e?�N*sJ�w���49��i�:XS6Y`l��	!�pGH�[��`���^1̀�����s�t����ʔ_�1���(�0'�G���TϘ�eGBLсJ�?.��$���F�(|��)�����ҩ�Ry҅�&7Sp�zS'@b�@��$XdhR��OPv�F��)�Ш������%�oN��b! �XS���,Pt �DK��1B`�4���w�p$�E�2wք�ۇ�¸I|�ثQnBW&+�->x4�����z4�e�2vԀ�ӗ��Ky�̃��C�`T�5)Ȓ�2) �1SpHu���F�[��Qp��%~9s��ն[�l�dɑ�*p�bV1Rq哴6�`4R�kL;o�$%�5�Q�6h`y3Ǣv�ʠ��k ]= 3f55�n(n�v�t}"4�¢ l�Ъ��݌JD�)�"��e�V�����;L����ٳ. �
��x�acՌKE�s�Hh��D�Q;>5,֎�|����2 y�F/�3o&|� x�0$@�4m����"���L�wk3#i��I2l't�x�˗�L\6�U�A!+�Ji;%߁.f5�%8R`�'�T��D�K�Z�9�H�-WМe�' ��d�a��1tF��T�U�"��p�e��
& ;��^NHFQy��J5\\x�1�C�rK��$��ֺ�bM�O| �p֋M&��dC�L�@CSE/�Ms���%1�`���Țmc�L�u!P-�Pzɇ�?����KX�:aaH�0�ʐ�ei�0=)�X%G59�k���]�R��B\T]jx�SA�����U2;"�%u�����T�QNc��Qd��85Т/ |i�d�GsT: � -�8��G�Hh��	��@$  �����~
U�d*"o"v�yqE��R�p�	�6��=�B�OVQjp߂U�� 3J�b��O��8s��lH����>���`���`:p\h�`U� �.����[� |�:�#G�d
B�1�
B?���X Ǜ#e6f|8@���tl��
���W�<_y8�k���L�z��0���&b9�A� ͜�!����I_)�P2 L�!�8P뷏]�4�*fĔ Ŕ�92+ô~�ҝ+��Q/gKV�Y���$�"`�Ϝ�:�z�'A�̓D�֔�8	���+f���1D&�>A�)�wrR%�'� 0
�Q��+��R���0ׇ�2fu�4B# �榱��E
��Ի��&Afi��!�{�F���h˾��Pr� �6\ �-���iуZ�vu�'v��P��XH^(uKC*�+jxx�A�@[�ɜ=�4%S�2�R�¶�W�r��a,X�LT<Y�j�)mvd�)W�ۍ1��ec���"~�V�j�-F�L׌�)K>a�m� MԊ�9c);ғK۶%�����T���2sC_6*���4Ȍ�+���*39�u��k�+I���P�HV����^�,�����荂,�|� k���Ũ��� ��q!IF����E~��<1�q�N	L8,p��M��Z솔2AU�D?^�KY&�u&��qCN���j��+Ƶp�Đ XaH�"G�(
�<8B<�\<
 �PbL��Pb�g���(˵�߇T�0ii�	C$��ǲ]��] �%]f�Fm�C��u:����&N\�qHF씧8A Xx' �	��y�nѭN�ı�&�4i�0���) ��M��)T:s���Ɇm�3<	u("Z�P�s7��hтiS!��Q��%��)�V�4�0�R��ޑ& �E�!�� >�j�"����c;�DU�Ҏ��	��9*��\�"?���nՄ-�:���J]�#���)�c̼ �TIВ>�!�D�U���b |I��Z �'K��zp�5��أ�D�0/��2�a�3x0�EK�?�N���	�-�&aj1._�B��7�(�2">	��ڥN(��/Z�F���X(~�6�b-����!*�&E�^
�R�j��[�����O��������Or���A�v�b��@'-8^� �'A���ԫ|<e���ǹ8bpA1��N9N��|���)������@'u�$HZ�G9?:��'��A��n��Ϙ'8�5a�̑xm���Ø�,m#փ�5����J-Cz4��!j����A<��1�i�tHK�"��yqB���+�����Pg`C;E��G�D�>��{B�yq�IA�n���t�L$�Bq(���W�
� `�6"�*|y�T� 
�Uq��P���2[��3�u��X�ZH(�(�.R�W���E1��On-��B�L=N��#�U��Qq����Du�K�S�"��cI#0���1��P似E
��8��$:�n?1�eE�Q�D��Q����	�I�����G�>�t��N'��D��:T�	0�|}.ٻ$� &B�H�qC[<ܑGǓ?ND" �% ��I��F�?Y�8�5_���I��'mP���Eȡ_i��:Ȝ� ���̚��$Q<\01V�"y����m_.\�eJ��f�������ٲ��إS9V$�̣z���XA�^�]�����8(68A��t�~�@�ܺ*j:$���C�0=�SΝ1��X���BN�Yr"I��M��Np��xd$\� -�L�H�{���(WI��AH��];0n����0�]B���3H�;Wjl�熊��'hd�3���	� ���Idb\(9����	Z!B�zr�Ũ4N�0F��.A~�J-�N�r��_�e;JȲ��cR�����M�������h/�l"ٴ����*�ViI!��,^F��̌6M��FA�D@/ZHl=�o��8��*0jTK�.3��ܣG�I
LG��!����/�r�cQ"$���Ȅ�YA*8��G</t%)"/ڈHO��L>!2oZ�IL����fL/v�ů� H�j�t���f����Z�T�Z0����N��� �M,q�9CE��I�z)��a�)c�([����Or0�M�2#�m���W�b���D'����ɯa�aE	�D4�uh6���L�x�*&��p��EA�'c�*١Qb�
��4m���&�T��83H��aT�"���S�*�N�뮎��x8%�H�p�\�Rդ_�mnB��d/�X�rl���dӘ��m	1�����V�I�t���
	>2�Иx3�_^?�G��-QE���#ޖ �<�����(AGXXz��ȻX2�EYp	�ڄ2$d�����C�*MpB�T����4B^�?hQ�
�5е ~qR�P����%ȕ ���M��n�E12!a0��Q#c�9{�2�ґD�!���;e(@�R��&�!#f6M�tn\�V���4|a�t$'*�ĝ��*0?��hA�Œ�w�L��!��!@���M$Ru��C�����m�������T
%G	�S����A��"tѠ�ͧT~��k�-M�
�-!���+D
�ig�
&6���������}�b�0?	�CÚ$)N����#6��d�d���s7.�!��Ը+nVWi,d�b�L%5D��bݖ0�\q�f"W�+i�\Js�K�[.�AY�Եi-�&�'1N�0���|�(������a���#j����k�2"�yp�J� ���J?�	��ә��A´�N#k����S�i=.h�v���dU��a����wa4��Ї�38EF��ቘ4=3|AwƓ���'c���@(Op��`���§�!��@`#�5tnDy �f��/{@�h2ឌ;|+O��H�䂼|<�v���N�7a��n$������h3B<��lD�{�xR��p���`�G�JŢR*H1|Xup�Ñ9��88q�U�/�� ���4H<�۴! �µeU `〉 ��%yRMY@���@" s=j�ґ�Ĩ��u ��6E�a�!�F�n�c�UA��d�\8"� �/@��۳��HA
p1K^  �2��8=<<٤����`�?���CLH%�'�>L�qߠG�@ �</3��p���O�%�䏶p쳲C^��,d�Yvyx"�ڀ��t��@6��r��9e��׈VgzT:���*���F��j3r�`e�ǥB�����	(��@�e����-肇^\��ի�"ۊ"T|0�(r�Y��X�+��P�eF0��	�g~���Ҁ">��� �¤�.Ų %G�e��|2������I�lX��Ӭ��xx�#�-[�7m�����88ʸQ�GG�Ш9Q��O�o]����%|q�kqm4h��8"������ҔF�|-R�٫0ܬ�0B��oܓnTb	'&�l��$Jd+�U�J���EG�qbv�i�Ӕ(V�ِ���F�:�ATF[�w�<A�r%�XUit��O��a�O�҈��b��,2����;tBR�~6d�����	�@��M:�Oƍǖ�s"�=G�-,01���`�
�9�-�!v�֝ɺ�u�H ���8T��78Lu%YЀ$)��M�AR�����R��@�U��|2t�ʘ
22X05k���!ci�KϺ���n�Y�"P4����D�ʣ)^�-ѶN@�5'�9CI������ؓo�yS�1�襉�gT�d�wT�Th��ۚk}�xů֡|�p��E�Bٶ����!�	!l��X�� T0��m��IߛT��d)`FҊx�Zy�-�$O��)��� b(���ʔ6��}�ԩ_�Q��XA���~�&��A898�����e����a�b��#��D{r�&gG�tc�&'n��Ĉ�ܞ1� d@�U�QL(���+R=Fl��Ysȃ#�L�iE�SN�0�3d�~�Vʏ+#��|�ٟ�*�A���8YP�R=$�����P�IS8(��d�Z�T`ܺ1,qh��@e�+I9�!�'|`����ø+X�p �ō)�|a��[-t&��R�XАr�m������/J*(�"���m���!� ���`F9 G �8���gOS/T0�qQ��uh�[��	�|�&զ��0��G��u�Kן2=���U�_�GXu�@冏K�n�a	^�����Yx���KV�hO2d ���o��U����%z�X�Ă�g����7-��a`�F�BF8pXF�l��]���݅ r�a�R��ۆy��_�<�V/�!��"�&C6�d#>9�D�E�䙨CDS�S!��P�Զ�x�8E惈K~���Ό|TMa��Vl"��$[�����O�D�Rc!��?���h7F�?��YC��ܓՖ�����n;��CG�|��A�o9��k�ܴn�1�0m�>�p�&[�<q�FN"�=X�(�2����B�c���yRoрQ��� �.�,�H��Ξ!�)HՈ3ɸ���胏g���m�-	����C�x��ؠ�O�E����� ϩ;��W��	���,�.�Q��}�������F�⥉2���D��LзCB9gͼ!�g��ul�oZ��b``g�5A�� {g.L�w���� ��� t�q!�I�dCZX��m�P��}RA�[�����I�9Ԓ�x,ݧ~�u)O�|k�c����b3� .���)v�P�6���4E����X��O�b�b<H�#G3Ƞe�UHT�-�0vͅ��Mj4�L�@���a�1�X��a�$@���c$� >J�=�Q=��yrtO�<@��t�2�V��1�AU.s�@�5 T%�'#O���� �� �8�P�#pdԃH�6������!��t���GcB8t�������ysT���.�#{=4�;��xa駇*�(<���C;q���ࠖ{v^���N��y8��ۄCp�$��+%'����Đ5ڪa����L�V�Z��:DaP�M�HPʄ�D)!+�͠��1ӸA�j�Z�1�%�=6�)X�K�/��͛e�͑2ZV��1�� A����"*��[�b�Ġr�?_���w�ȾW�P!Q�������ޏyG��{��#u �k���(������I=P�H	2��?����x�� �Rɚ?ҙ�vJ�3���0/����p󤍰.��ɋ���
o��]�࣏=�����-�K���P�J��n��E��К ΋�1���`���|��q����<+��U�V��G�OjM�W�!/i,�<�`;r���P&��ɚ
����C��+@�?���pd��xF�P�1,ȇclT��3��@n��lܵ7������ײk��L�57�V`��R{x%(OQ>�ᰲ�(z�E�kK�y�#űN�D01� sRxݺ��Y�c5L<�����t(	B��,iN�%1vC�2H�n��g�ƅ{����j=hZA�A�]BpqN��
\)��"���'����J1g��R��S5��IXtaJ.T���|J��nځ@��
%�R��4��/���(��r�IH�{Ϯ!��*B+"��ePᬐ���'(�
uRd��q0�ԆSM����y�y���	�1���@1.Xn s���Lq�CZ�)�8�F3E?xE��^0*�V� Ë�HR�|�iؼ�y2�1��)��E����7n�1(�R���IW�\A`�?x��%���D.Jl`���z �GD�j���PĂ$�O:��֠�-t�7���s�4������i
�t�0G�;w�$�����l �$��F	pp.�cW����.�Rf6����Z�ko�}0*��3�a~���X��j��׸-dD9J���/�I�G�Q�`��b�աc�Ȱ�.Z|pu�@�V:)lH-b�L .�����Ă�oïE(\���` ?���@4�X�y�5(�:��8�cG;X�Χ-�`��B�2�F��!�8PV���ƍ<%�pa�(E��Se`T꺋���-m�$��%�Z' !8@*��������-+�4!HAS�_z�I ��6�4����8ˀ�Įk�M�፝�Q0,3��/\h��BJQ��e	�\Ip��D���fPy�ő�,�D�h?)��*.�hL�E)�/'0PyJ���W9�����F]��]�eP�9�f�VN���©ŀ���D mϪs��C�� �Dْ���z�+�%�0�����+M�q`/.u�&mY�oC����>����	[�oV�c��{��l�?q,U?XF�ݺF�9��сf8-�R���H�{FI�1w9`�4W��qÛt�>�zf�?�=a��@�o����ǉ�l�Ғ�J���t��{�OCy���q�%ǂcW��"e�0�j9�e�,` &%N��p?iR�؃������]'n�I(�._�'~����@�.w� H�)[�S�VX!��ǥ8�`R� 7[��B�I8�H�����o�y1b��=����*(�`p���!b�ի駈�Hq��/S/7@(�bP��<I�%*3D�T���qߐ`�G�ڵJ]>Q�auy�a�%h� a�倆���	�)lrXH� W��@I��G�h������z��ѱ�Xs�,���85(�g�N:9�(��'��a+�NϠk4l��s�����ƭaD<9���įݨp����n!�*���@��y��W�N�x�Ț:r=�D��� �yB$P�u�^����it���N�6�yB��b����%
oAHt�N��y�K���TzǬ;e�b��e���y��0�P�$ΐ	YI�MA�Ζ�y�%{bV��R��&̪̔&��y2���TV�i�&��*�WJ˳�y"߰fU��_[�8Ƭ�
�y�=+E�]0�߬[D���	��y/޿Q��(���J�m��D��y��M7|���JA�FI��#v/6�y�E�E=��3.J�6v�B6�Q��y���;r�=@+�|�8�
 /�5�yREI��̰9�ʏ?g�8ݒ��3�yR�::�T�"��*^����$ �ye���6*��Ie8y�D����y�`�-(&t����A��)����;�yBfQ!1q�KƭD�q�>���@��y�B&EV�a&�S��#�K�y���A؀�p%�-C}
�ȇ.W��y�I�L��$8,@)<h���E��y*�4]a�t�wl�X�^� ����yBr��ѧO\Դ�6�y
� P�3�7kZ4�z��U1$zP���"O�8G��2tc�9`��� ^h��"O:�3�<zn$A��+aKb���"O�Uà\���YД/��Z>^i)t"O	s�gҡ� �"VLܥ3?|q�"O���KD1z��;�L
;Ij�S"O�}���-mV�sa-��x���e"OZ�X�쟶W�j�6�ڪ.�"��U"O��˷C��H[��G%ؘ�e�"O�G���'�\]2"�ŰoA�<x3"O��`�ҒvIR�+�Jܑ?���"O�Œ�J�����ɄS�p���"OF-��DW(O��� iP#ir:�T"OX͋�S�@4�
b	ٽK��#P"O$�[VA��`�:Q"\�(�ԤB�"O96�ʁr�V�7��g͢�xw"O�q�%fd��� ����v]�U��"O0���R�;�������w���j"O�B�n�m��c}��D��"O��#�Փ,�hL�"�weT��"OȲ�h,w<���K]���P�"O<�� ��O.f�Y�m�N}�%Ҷ"OP�x��	8h$��0��;ή(����f�j
ç�j13CZ�^��c���h��	A��326�����\�؅ǘ�	�N�cڟp��`9����>�fY�O��E�EJ������'�J1Js��,)�[5�[,`�� Y�%I�|;�h�6:LhT]!!�0-��W-xJd3@�D@�K�mz���'�6�Ilܧ)t�z'�R�WB��c]�	[p�D{�"� ��ţ$bՑl���pG�].�)U�.HB�
q�НjX	K(\y+��0!5��D(Q�@@z��L>���X K�	�2g(3a+�9�6�ؠJ��b�)0f�䐡g o^�F���X! W�y����0����j�C~FA1噥o3\�0���p��Q���(L��W����B�Ȕp�* ��rӂ��Q��,0�X瓁)J��`�m����*C�U؟t�_dM���q#F�!�݁k.�O��#��=�ؗW�&B\� M� 9SZ]��-;!b]B�BE'����T\2,���▤+����8R�'K)�(��6+/pl��ރL�R,+a&Q�s�n�OP$1�Q	w�zE�rFK��	�*3e�i�)9^�K�*䰴��'.IܬZ1�D?v�z�D��*'�Q�B4�\�[ǎG+簰�J�4  \|ě6˖7[%�b��ANpHb�F?l�~Y��/�^$9d@�E���ug��$J���P�پ%�t���@�e�_���S2`�
&�P�<:�ω��'h��	�������cb�`궎��U��1��)�)X60Y`�oWc�O�|%�v�i�����7^����L$�QГ P���@�vbP��o"��i�´���އ8��@e�=(�4p��EE��a�kF5]�.���k5teVyt�i�p|�eB�.�&\SG�D���Z.E�M�5oT![2��`H� �#ª �Y�V5�E������+ �v��WnM<8ڇH��mɆ�
�I�����w�M\.�1���ڗ�,YSv�H�}̨�Ebق�u�1,��a����7'�Y%��q���&}���pQ���<5.TyA��]�`��E(ɗg:��S�T�L}�W�[��`I�Ú�5,PqQ�\�j���i�p�@��8�\5a1��@�6�1�mN�Qaك���^�Cdm�7��p�=�D��:B�2��O>dJ7��W#�,(q��/pJ�*�c�'v6H�[ebJ n(�R�$ޡ38xrGCd݉�R ������M� ���KR.��1W�!��C-����%> ��5�]�0����P��C*��J.t�h`ѢH;wW�`)C���&'T:1�A�8�F��#%˖3�R���$�0���8]�DQ��D�?Q*i1:�H��c��6�ƥ�0Lˢp�*�Y�M�>��a���ɤ0"��<��%�t"08��(�:
mP|��|y�%����ZbՈ^_�9H�H�P,�#��̯$�T��]$�9 �,�0G�i�H��Zwd	��{.-S�ʌ�(﮴��X3�M�7�i�X�QFE��(S+���<J�L�dY�})��0'�t8ð!a�N%xS��7/�Ɣ��aЍQ���I')� 2�.U���ͻ�0uIq�� (��+��GD=Tq�F�d���F��Gh�h��YѲ��ӟ��Q��~���f��/��If)B>L݈����l��e�rېd�(�K�쁾J�V�1㉆�c�����r����?�dC�0R�b`"T��f�3?)D���g��Zg�����E������q\�b���.-"t TH��y\�(qGE+s	���R�F����agĈyH�j���>�m���ܣU.�������Y�È���5��I:D`���ϡ@{����F��s�t��'�?	�iJ�皯_k��׬�;{L<���k�%v�тU&ټu�`���$S=����,��H&���`Ȍ���H��	Ez-�YxK焳b���[�M wݒ �ش,]V<6 �֑��A
3�rE�b�d
�i�Q`��-��8Mty�釁so�\�b�4��t"G#<����"�����jL��M{���QD�k B�^5F�1s�ŌCr6`��87(��U#T�5�\�P���Bh��PŃ�DJ��5�N�4�2�OH����/5�6I#���V�@Wp؁�'�=��	���z9�rh,��	C�8���W�D_`ġ��7��q�B�k�5O�@A��:@ ��O#(=Jl@��K��p=�㨊�� �©ՕC
�$�ХZ@L�)���F@aAT�Ͳ_�]���3�"EX��TG�0��e��CK�='�� �HqQ�N�E��	�S�ܞod�I���6|��`�G�!D���1�70߮�Q��J�`�%ÂnѢz �*�.�����9�H�.�9�w��+ 늄ȡ�'ޞ�x�ޡ.��9�*ݧ
;���4M�T��7�J����!3�1Q����B_*89C��:Np:S�[�Nhg��c�i!�䃀m��۳"O@5��!i�4��K�U�-��oԣi�P
�f,i���%Y3Z�D=�����!k�$��J�]�1��?�,qЊQ�4{�����;S>qqW�'R:}Q����I�Al�$^�-�G��Ỉ*��ǂL��	�E�t����<>Ȇ��NR�H[b#>)���L�-��gY�A�0)�,#����I"m�
Ȓ�G�W����ͅ�?���L���7��� �PjP�����~{3�C;c����>�~��ī �Cd`��4.h���W�˘OX4���7F�c_�3�r�+��c�䆾Wdb��g����l�@���KhHٲ�E������:X�~ex�,+Z�}I�����*X�7�5�`%�h[�$vls��^?GDȨs(3S���``B'|Op9+�h[�	��D�7/�'ZK�����L�_B����ȵ��d��$ܾN��̓�E�(
��P���;�/*1����)���9*%J��`�L/}"��E��ईhb�77q�����iB����E�)9�Ex��M�6������,_\���t��p"C�Y��T���'�&�Cņ�z�P�ҟ����#m�����>�$��V�y�O�K=�!����"2��$ZwHN�3����#_ [�bO q�,�7*��CJl4ң*�e�z @!�|�����#?�,P�놂 �$�'*=ғ2*<�$d>5OBh�U&H���z3!1KI�3C���\j�#�H+0 ,�t�Q�7JHh�%&	� ���C1 *�xJ�`�*��	y��@+YI��XbB% ����'�T8	!œ	C�<�g�[�bR�F�ůdC6�p���uݨ-P�f�klL�
��C�D�,�#M���{! ���M[ڴE�&�0!�:y�2dj��1;,�`�d#�$�1:(�h�'����wjB%@3J(ۃa�0B,�X�(	�^,4F���3��5r�2J9Z&��J4�:�Xtg�W�d�����*��- �)R�n7M�)`+-Ѵወ  B�d@�m|����i�0h)�D��$��QMNU�L02r�IN�bb�����q�,;	p��&h�~F��G��7�n���A׿m�t �w�Dzn�m����~��N>���v�Ib�X{�q1�D�n4�M�-��#�Bm�E'\�>X��F�^݂�9�o_s�YP��8o?�eQA�"�@E*g�6-1��lì��9��B��tL�r@ѳ��� L�<8�e��d��q�e��6&>^��NC�9����m���X@v�P=ii��oڼ;Z�I��B��L���:zz(��#�Z�((뮂2��e�Ξ�J�� ���A9gxU����k�6B 3Z4�
g�n�� ��+'
(�E �*v8���o��mQ���(WBmKP����x�d�@� �
�P���yA(�6]Fr�q�� *QI�V  =(ő&ˉ5���	�FwAMK�=̀���,2j5+'��м�s�L要���.a�����'s8�a�ʐ�[c2�rfHO�]"eɕE6��E��	�/18h�ՂД_\�ioZ�)��(Q���N�R�⛟dI��K�	�|�x�E(�9�A#L��� ��-S��x�2ϐ�m�	��d�)
h��J5�+�5���X�L���@FˬQ��`�2o*d��� ��2oM��ۢ�I��j�@	��I�?d*EL��ֽ36�sSz,�s��SĠ��b9������ʍ�
`����&J�=����lK�>�J+b��#�OȤ��D�?O �p�+^`�����l����,���r� Q���~Cx��ɬZ�0� a��Wp���$�m���ݴ"`�sr-�=$h �j�C�j��M �Y; �t�î"3h��Ξv����]�Ȩ���{�	�B��ŀ����!bg���.�,�y��َL���i1�Y#s�8��k�C��F�)Xpŗ�8�$9#�$��e]����`�/&�t@��	�O(HA�E+O���q�"�X��Ŏ>+��H�T�_�juh�b_�n��ē �H�˵�ֆu/��-SzHAA�Q*w�����<�8��Ӓf9��:G�S^�lMEC5#<R�!�dP���%0���3Q�G�$�|(2LƔD"RyX�R��{J�m��1�5���1� [�E�A���L�@%XuH�'R	��C�j����DP$+9��1C�K�W���Cw�\�r�I��c	6�8(�.]=p��IgK&.2��aӀ� U����s�Y�#ٱ<W�XSf��Z�H7�V�c�=�刄0g�P��`ʹq�n�2�V/���A
 ��r�C�ޢ-P��*k
|q� �8*8$����V.��fA��A>���b����+%���|��J�o��Qn�4�O�}8��)�d�?�Z)jP	H"N�𰕠��8����!�	҈8��j��_���K�91�؀�#M���5�Ϙ<����q#I���*8Ƣh� `�J�8����Շ7�f��q��C~��� f�K��pdI��(�*��G�\a�h���S���0��;-��Yqv� �:1h��:����g�j�˟ԉ��]_٪0�u��x����7NCȝ� EG/]YȜJ�i��Xؖ�H81����
�U�d�p)M�l������\���)�����B��#'V5]Â��Ɇ%>�dL�/<whE�U�On@�q`�CÎ�5\���#�i�$�DS�/�bd5%^:��V�Y�*�����T$Eҥ#Y�h ���ϓ�.��$A��_9��f Y�8��2I6r.j�	���)T.fq. �Z��7q*f�1�'�(W)hmڴ��F�u��$�uξ�KQ)G(��c����ӈ����I��l���Ѻ!�I��m��;�4�1IG���K��5Ӗȸ7S?��-��:��uA�,ـ:��1�Lʳ>��e�s��W�']<�`�"|��R��7z�8�`�AЩ\��a%��;U��+�aC��%��Q���k�%ܾg$�'Pw��§m��+����L;������[��	 r)X%Gj�'�0"�!N5J0����JM_��%@�i!A`����ze�y"Ý�e��PiĆ�P������";ʹFI��El��%��=������OP�:�-�*b����-�ta���Pb���'o 6��]�B�]\�(uF
x�|0�.�ri���� ��W�-V���a�(9zj�Z�l�W�RHS4N��[���s/@�`�EHķC�Ҁ��ŉ��hOL$����L��D�RM�#��=h�$��-g����)�|�	2��1AF0�r�8O��L���&���'0:����+Ϋd�I���9�j��Q�[X��Rf�I#H|���DG�,w4bt�qK\�$��%A3��SꙈ��G�l���bIߐ5s�8{%���>``4��)�~���Y��F�q�#7J��	�tg��-�Dy�$ɺ((Z��c�r�()^��5�3Hr,\����E���B	^8z�	%�� "I����e}"uP0�W`;�����(�6�V�rI8��Z-*Q�+�d~(m���f0�����RŦ����%tN��X3�\�qt����S��@z���4���S�AF�l�H� �(M$wF����]8rt��ƎD�T��4*���7��P�����h`�Ł��uF��Ɯ��AЏJq� ���[e�O
=��ȉ*�2���dC�J� �a������B̟,!텋^h��ψ	����*VPh�OZdi�C��%x��3�ӻ1@��oݕ?i�Yx "�+��'�(00�+UZ�ЭI�N�|��i3O�j
4����[�$4�&_��8ٰ��Ӽ58���j��i��r>ᛰ !X�"4����7�,Ř֠ܞ+�i����murըE&�#�剘��ɉգ�l�LK� E\z�m�78�f�j����i��t)� S�y �2�4\r��X�y�/�w8IQlB�`U6��%� U�
i��0�>HZ�e�Z6�G�v�p��Q�
L�Iw��p�n�2��_`��Dېv�tTg�/p�f���E�#D�Q��ǔt�|�rG�˰>�܀W�&��S6LE:x���+A�y&�pB�>a�@��K�?���<!'˱;�Ԝ+RJ+2>��  N�r��Ke�̺ ��Y�"����;��^�T��K��^,="��� =q�����:'�^���i�*x����.ڕW�n͑��D?[���׍1�	?Z���w퐌O�i�I��L ^�E闝a0~,� ȃ6R�"�RF�/&�r�6C��*\K�M�)%b>�J��`1r ��H4W�>�Jƣ���ǘ�a�l�qM!�2���ʭ�~Bˍ3o�pGIY8Zp!���2|�д	��P�s��e��e��;���Go,j<�q��S*�p4�Cf�5{������f�4�:0�;gY��(��9��kQ}�!���YS8I�j�0>� ]����#@���еe��1���SKP�~��!*�*Ɏ]Y.-!c:�l퐒�@��H c6a&~"�V���m�J�8t�5�s�� $F�/Xd��	3=�<���G�$��EC�R�W�d)�'=�8i�i�.�J%i�8�*���eǟ&���I����@j³y��9���E�E�̭#�ß��$��k%A��b��� ��-�̽7(���5�0XN;0ƿ���j�A��  ��D�Xz��n-u�HI��=h�M��"��+*PKء�2�I$h/�(�qÆ7��=Z�(¿n�A���O),D(��"�(� fصL{rDӸ`�8;�̖�O��E��;��?I���8.�j�լE�]^��·� M$��/��_�P��Ee�/x1��r��+�z%��̅>XV��gc���P� �p�r9ځ�Q�0^���MB���c��A.��b�B�0j���!�$j.]�E���*T(�#�c��{"��FҴ\d��¥C�5`���aSH*�'��Mٴ�8�����O;pQ����Y�+���J��A 4����	�.K�)bN�`�4oFVb�u8u�L�Om �dIH�t�1�晅Ulܐ��>)�Dǁ��TX�Kc7\�:��B?1w&B�]��8�a�W|HJ?I)6ů�pP䆂Z��X��W7+$�e�+?�Ɖ�� �mz��D��p��}��m�7m���a�D=0�,g�O��<ej@O�5
�ҵR&a��sQȤ�c�F$��H�;&�u� �S�`�r�S(>����bD���Gԓ+�� ����� ���WyJ%��*I�:�5��NM�1���q�甒)���}ΓQ	&xU�T�z��xEg��4\�GB��-Rj콊g�U]�S-)���0�ڗf����G	�d0�����i"TӲ,U=���wF{£U�VXޤY�<$	�y�Ԩ��I�yJ��"�ԟ��X �T��ޝ�%,�(+r@ r�vcđ�7V�[ʼ��'�O$� �M��b�P�C��(�d0�퉮H6�t�o�3�툇��4� h�#)T���3w-�y�*��/.�0P�, �f�C�,�?�¢��<j���18���)�/i�yJ� ڀtAʥIGŅ
(@:(*�'���b���
j�a�FNߔ���C�X��J�	[�VXT�GO1Fx��A�x�D�P����e8VX�gi\�p?7�Q���%���-%j�� W9p������N��C��${��,�aj�9Bz�Z�	��6MF�?	�h�,��b?�r�.\����J�9Y���3�4T����D�D�֔�[�}ބ��"O$p�,t9�`7�	X$��"O��"��ʙ��!G�eM��A�"O���f'���!BE��A"��"O���ҧZ�h��l���!6
�C�"O��RS,O�&8Q����*DQR"O��Q&�[�Ew�����3$ �!�'�����)3>A��IK(2X��'�����+�;p^8���A�n�,@�'2 ]₋�D�@B��Ρ�2i��'��������@eH^&	�>��'�u顧G�ZE��6�di�'�~�q��<e㞙s�NΥ C�|��'Y�-��&Q�+�>��ҋw[ q��'��,���ūGr=p��A�78� r�'_ �(�E[�`��ds���\��I��'�N�2��Q2	�N�� ���`�|2�'�	rs �����H�ilPQ��'�v�iB�a��9#�׼_/��R��� F٠u�X7�X(����@1"OE���,�nak�E��q~�#�"O�h�!R�
~��PVc�PP�8�"O�y�Phέv+�呀25M��"O�����Ux������6P{"O5�����X�T�L�z��p�g� �Q�1�ɵID�@��؍�~r��,�A����nJa�0!K�0��7�!�d�,����	6L����R��$ ��Q󏍎#SO\	Z��_��M�ᓸr�C,M!
�<e��S����4�*8���f�pOQ>%�l�]@<�ḟ�G��"(�䘏�(O���Xd'�����B�֤ۆMq�\��`����h�q�|�-8Ց �A�{<�R�e
��M���E':����Sⓔ�e�;b�R���C�C�lM8���=�z}�I
�����+{���ç ���[W��,B4��D֕@fH�"I>�y2d�Jb�Ij>["? �䐤&�:��8��S��b�Ik��C9>���$>���ǘoox�rD��gN`�`'cX0�~���G��?q�$��v3�х�Ӫ\���!M�q�w�EE������j?:��Z�y\YK1�ؕ�`��_��m1��(�����=?�r$Y�/Q* �%C/��41�X#Z3J�;�� ,�5r��OՒA⟹o��h���}��LR�0�\)��Գ#�ȩ�%C:Z�&Q#�UBXH93�'3���Z�[>Y���c�0c㖰^�d,��ڥ-8�J317l�uk�"OI���	�[��[��7%Mh%�L��L���9��J;u�x[¤�����۟Q�֝8�*��a+ <(��s��,@.��'�T"�'/���	��1.��겠@��z�3N�5/��~2G�H�)�'O��I E�`t�I�*��=2�	�~�+�V�i�@��Sp��X"ŉ�
���|��A��i�:�A6?��'e~Z`�FF<mpD�@+�%R]��n�t���'�Jq���O_��gE(8������S�F뼥�免q~���'\����7��ɴN�ڴ0�'LK�3�����O��ض�Y��M3s�J���>�"#��eVT��V2l~� BoS�ovHl��f�R\Q`�˹vӦ�8�ď#@�X���Є�S؊H�ve�pO\Q_B<�ȓL]� `Ջ�::�h,8�J�x�b���:U>P��o��|��ȡ�u��@�ȓ5 ��ׂ��+N�ԃ���K���� ���iV�γe���!V-׸����ȓu
�L���$Dr�@�a�R�"I�܇ȓ�ܬ��/�'\��\*��7wj8��/@)�vG�R\�8��l�1������a$��3rx�v.D>����ȓr��;s��0]:�D�7��zdt���Zb�tۄ�ʺK(Ke�,ZlC�dQpͪc�EP�d������s"O��!K�f���J����f�1�"O�$�٪KԔ�Q���#�Jh��"OtآE��	�dtX�ζSyl�"Oh�P�׀@���y�+U�~�+�"O�=�P�ۄqK�m#�ݿ[���D"O|��uA� ɮ�9`�4.���$"O�t�҂R6Q���eة
�9#7"O4��΅�.Z��B
�M""O`A+���o>,1IDa�Q���W"On\p��)(L,4��	��1���"O<Y0�.#RX��j)Ht ���"O����M�T�B%Ѕ/��*��|#�"O0�`�	I���c:)�	�>Xspm���0d�ղTy�|JG��e��-��MJX���s�ǨE��q�,^�yb��.=�RyKb�^9+�$��K+�y��J=w.8����%J,@ڰ"ŏ�y�F�;-�n�ʐ'�M$�e�Z�yr�J`H�@���|��bý�yb��20���Llk��P5�	��y��O$���2Kb$����3�y
� ��iT�D@�럨=���"OzXCda�.aƔ8d)�Ezl�@"OV��wE�����È�am��"O�#���>��k�슩+E��s1"O���m��2�n��s�K�!�p"O�ࢱDMQ�����AK�1���z�"O�q�+؏X�V Җ&L!`�2lJw"O�0�sOaq��q�0rBE�"O�����Q��ځ�#�|f�ɕ"Oz�W��'#����*;I �s�"O�p�"f�~	�i�uյJVl��"Oqp2�7akj��I��m�x�c�"O�ib�$)bK�2�B�Q�0�`�"O���<� Ā�w��H0"O
�Б!��O��(�r�$%� �!�"OJQ����#���@���1�R�R�"O*#� �W�D +�C�|���2"OFI� 9^�x5Ʉ�	veN��1"O��`ͅwz�١ǚ�,[�0"OF囔�0���С�_�I<�0D"O�uؐ �%`�V�#���!'N�!"O��$��(���s�H18t�CU"O2��$��Xe�L����*!R�k�"O`��ٞ��mc%�^���"Oh���I�(4b"�fU�L�R�"Oʭ��&�eBT����h=40y�"O��!�'���A�#%����"Of���K��҄�WE.�8��"O��J�e^�@���7�.���!"O ��i�X�A�$�	\��z�"OZ��B��C�xH�bDT�X�@�X�"O��K�2H��PgË52{���t"O�`����*GuL�H�+�zy��"O�Z�N��D��(GH�xi�L� "O�)���ŧ`��`�eL>yU��{W"O��+D�u��R#���#�UkC"O5���M�~,�� �O�x R�"Od�R��l�*��#��}��d"O�@C`k§'�I�桀��r۴"O�THe`Ј,1������C�T�[�"ObT�@˞-,gR�x���Di�"OL�`b+��2�MZ'c�-^�B��C"O�tm=VD��L�	���"O����q�l�@K�:H�p(;�"Ob��J٘
�J%5,���R"O|�[��m�$����Z�"Y"O�9�	�G"8�֦\���"O�Q	g�A*e<����2�vu0"Oک���ʸP��uA���N����"O�)c"G�l���a�=xu�X�"O�,8rM�����%��D��"O!T��0D{0\�%G{�N�15"OT����Љ�6�K����J�"O(�jn�!��y��IڒQX#"Ox�n
Xi���AbZŚ�Ip"O���M��c_fTi��J�R���j�"O0<	�L��:��M��i��e�lLx"Ov�B�@�#�A!����T� "O���E�܃>6���	�� s"On)�B�p�<�
�(Ђ���"O|�9��8H�H&�4� ���"O� ߫�(%$G�_�d�B���N!�J))Һ`����"�&�"�OE�[7!�Dɻ��c�"��VÕN�j!!�� ���E��;��0��]�D��I��"OnD�O�0t�|����ؘ(#"Ov|*��[(��\Ñ�+�n��"O9H�n�B�Н�և
,A(�!�"O�ɪ��I���;ֆ̔5,ȑ�R"O,\1Wȅ�~�4x)uEޯq�IG"O~ #�
�yhИZ�.äU��I�ȓf�� 5��J~�S&��VTH���Yޮ(kp��iG01i��LU: ��:�v����.4ː��bc�*)�ʀ��|�)��O�R5PdQQ��#Ofe��:��P���h�1���!K[���ȓjϲY%�A�g�$� �,$� i�ȓ8cJ���Hҟ�j`Eᆔ?��`��}�Z�e��W�u��ᛑ+�%��5z����I^�2T��#��M�Fۆ�ȓ{�<i@eX,p؀�)b)�G|����c�L���e�o�e�"��?wxp�ȓ�����S�=g��l�P��H:"O*)�!ɉ2h���+O2�p���"O�JQ�)�k��-��i�5"Ofu[@��.T~e���m��x�2"OdMKC-B�P��1�Č�*S�h��"O��c� �a�l�3�Οp#l�Z�"O(l��͆,-�P�ڑ�\�\4#S"O���dJ����ST��`�(��"OvMP���2=�
,ȥ̅c���"O2]��gڽ~%X��(�+*��R"O�a�"�	�U�w�eN-��"O�%(��J�e��<�̍C]N�{�"ON(i�����p��K�!�0��"O�Ը�f��(R4b�
�;]��:w"O��K�K9�h�P�H.��|��"OFt ��ZRJ������*�<4"�"Ovi:QD
�3�ܴ)�CЯȠ�Y�"Ot}��^;�P�Iu�<T��|K�"O��LX*��E��I�e�l}P�"O�-���0s*�J��4y�<xY"O����/�M ��	v��F� �XU"O�w�OO���YQ���:�h�"O�kUoєrN�K'�Dg�]�"On���?�*ɀ�i��ShK�<Y��WK���@!5� I��KC�<Y1��>�r\e��a� 9�fD~�<iGZ?6W���U��h��k��y�<�AeB�:M�sb�=l<�c�x�<�ShG��B�$X�;Aw�<)����/��eB��΃����Tp�<y۝s��̊ zG�Xa��B�<AE䎂k�e�fCQ�����&�B�<S�A�U�$Ҧ��HzHz��w�<ylE39��)w钵�	RS��I�<&��8R'�x1U�bD�ia�H�<���Z�8���b�%� <^�Y�BA�Y�<�%"���r�Ȣf\�{�(L��G�Q�<q7HP�FI�p3UMO�K���d�<YqM�	�^Lkj�'Z�xK'�x�<�fNR�O#����)��Et�$C0��r�<��+k@�H���O�:kؙ ��Zl�<A�,��W����.��B�`��j�<aF��4>�PRecĚvμ��ц]c�<A�-v8d���\=��ș%�Pk�<)�N[�m�،	"�W�]�&��a-f�<9EI�%gP(�ɍ��yD+�J�<� ~��d�E�y+7�ȟ=T��x�"Ox�Z ��1�n(#S�MR@�"O�9�3D��#��@`�i
��K""O�m���պq�Z�
�mȗ}�i��"O$��UP�[� d9R'��-�|yH�"Ol�s�*ٚ~���f�!�i�4"O�����X�Q�I�$
�"O�<p�n��pni"1jG�O��]�@"Ol0�ǀ+&��=0b�T��ed���y"��F8(4�3��59�,u����y
_
t�@���8�� :a*Ź�y2&��]���b� y㤄�sE�y2➂m8e�X7`!C��
�y��ƽ��`�D�	"b��	c��yb��$��Yô��l��!Ó�� �y�I�=G�H�c��^��̀����y"J��'��(�fآ\V�<B���y�j�0a4�uJB�}z4iQ�̱�y�7j��\� ��w��������y�ǎp2h�`�#P"r"5�¡N��y"	U8�Ra녓6R�l�r,��y�o[=L;¬y�$YZ�pܡ�bX��y�
�4LD<�C��5Y���cn�H�<I���!�"H9�.�y+>iz�	^w�<���W�T�C���%5`�e�J�<yF�O�W��� ��"A?0)�0BAC�<�Γ�=N�!�2�B�؋FlIE�<��D��t��eGK�t9iP��v�<���D�_)���%K�b����)�s�<y&*� m�!�D�Y8�rYs�<y��U�0g�|��x���R�G�y�<��_�N\�T�%BS�{��(�!B�r�<�IL9W��D[����B��f�<aG�É?�N�w얺psjy���_�<�P�
�B�J����ó�����]�<Q�`   ��     �  d  �  �+  �6  nB  �M  �W  `  l  �v  �|  .�  ��    �  G�  ��  ˨  �  U�  ��  ��  8�  {�  ��   �  ��  ��  �  ��  � � �  �/ l9 @ \F �L �M  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|`I!'G#\���%�T��'ItcbꀀK<�k��̥:O��'������Ǝ8�ݓ���"J�S�'y`=c �d���	%�BPiV��o�<)E�I�M��c�Q'��I���k�<Yb�`��s4��/~�����M�e�<Կ��رD�E�?�t�Жgd�<��j�aZ����Aّ'�F�r�b�<��"���e�ďfe��ѣ
�[�<Y �{�<Ԑ�[�0�Rѳ6aE|�<�ǆȕP�,x��H�o���ۀj|�<��\��!G	��lhP�qI}�<�cێ�,����ޣ��@�#��x��G�<��Fъ��u��Z�JQK�%v.1���� ׋� ^:�Bэ]lr"�&���I�-4��Bbʴ9[��g.A�$&��$@?�vĥn9zt�&D��v�����Z�<�5��@e�
I
p%j�a�L�'�Q?y[��Ph�d:�
�Z�bg/D�$2��q�HÄG��R����I�r�����䕘!��8r@�P�Fi�	� ��!��̲��u*4%#\l􁦪��,�du����	�j�����
���k�h�7EB���˃���.*����u$ML�BQ���C���C�I
|����d�2�y�e#Q�B�	�� R��g� �t��B��1�s�Ee� "<E��'�����?l�i�|����y2�6�Şw}��̞�� `�d�ǁ���a����dE�D��p�i^�;>��S��%+�|�L3}2jN,m��+�lRu��iT�y���>�����Q�g�عQ� ��Mˌ��%��|ph�9IV��1�!�;qu��UA؞X$�>�XR��V�ԎPԜa�g��:]&���d(8a�МA��řcYx�h�G��%ڧ\�ƠB�!3]��`��G�44��^�Ȅ�-J�S�d�Ӱ%�'
<�'Bў��$��Fa�,ʕ0�i�9j.!�$�!i�;��@�f�I�Iſ+� �牰D�-�Dk�;�Q���c�C�	;<�4Qd �
����'�4��'��Bm_�K;�HاA�H5���|�����Hȸ-&�tbr�Žp#��v�/�yb(Ͱ6��9�L��o�(��^��~�!�S�Oaƙ�gh�[8|`c��e��e�'% �;?ʡ��� J���
�'��s0i�3y�Bd˖��Vy~9�	�'�F��A�^_8@�D_�M}F��'����7�[�Y��:C��JF���'�*ex��N�d�B��9;� b�''��SѪԮ4	�#"K��7cL�8�'����d �el�0J�g#����'�HS��Q��*�р�	����'a�|@0l�9�0�p�A|�`<��'/x2���93�]���:%���`�'W��P��҈4�����)뎨2�'R2K����y(J�0�D�Z"m��'�~���j�$)ԡIg�0����G��O����^�E�� �9rdx05$?��{rɚ��I�m#��Q��Lm��$*Ǹu��ʉyr�'q�x��H��t��ѯ���r�H0ND$��=�3U����"��M�霂���.�69���ȓAR�L��/�B��ǭ��-����=���?Q��Ӟ6 ʝ)��^�%x"T�&��~�<Y���7?=f` ���4~D|9qM{�<����J�Fa@o�`Ѡ�sS�Q�<�[y|�d[� r:���`n�EB�`�'F�|�ڮe��)҅��F��b�O���	^���O(���b�>�bI����O��p�	�'eF�Js��#y��L�Ǆ�U�
yK�}�x�鉷4��9{�ɐkL����N4Z�rB�IlZ6�+l�	<�ؽ���Pdֵ����'] �cV�`����jG�%��9�'jX-���_�"�ba던�Da	�'�bY��R&��l�� ���$��˓�(O��5,��N�R$�7/T�j�~�J#"O�BS�]9af�K��G�Y;b�s���=lO�A��ydVEk��ה:0��"Oȑd<$�X���$Υ|����"O���t.R9ǎM�1���S
nj`"O�:AJ���,������eh�ha�"O\�!��שn=Ҍ��$�	'�<Y
�"O��#@E�U��C��W�9���"O�؀�J��}:5��k
:�P��"O�D�G@فE5ZA�Cj`D����7O���df��	Y0i؀}�~��)I�5,�,���'���ɉi����AE\���z�&I����5�I�|9������?& �S &�T|�B�	���0p#� ��� �<}��B�I�Jz��5B�% dY��T�A�6�F������ ��A��ƛRTV�BpH�>���6"OL�ke�I�Z t�A��V)(��2dU�p���h��Q#w��
T�� s!�F�H�ZC�I,A:� Iv�CQ��2�iħX+`B�8P��(��_�!�l�s�H�3
R>B�I�T=dX�!��N�ZAz���._B�	,$��rVk[	l��-q-�)
B�I�e|Lru���Z%��� $��>r�C�	0����ThW]jP��-B�6Z��#��c%O�>�ȉ0�F.`�����4�O��$�QԅƪuJ�AK����>���0ƈ3D���� 	F��AƂ�5�a �M2扃5���?�|b���b�c��$��iIGhd�<�0�� T�4+	I����a�`�'O�yB	Q�$�� ��>;L@�cc/_1�y��%&�&aYF.đ-�E �Ј�y�C���v�Pg:��P�7J<�y�n 'Ǻӑ%�0�؍qbC��y�ώ?~�Pt,(t������	�?����v\8���,�H�Pu��!i|���ȓ@��-Ӥ@+n�P�Sd݃B�v,	��O�����!3��q9�(��D���fcҖ^����)"?��,�;�2%��۷�����(�f�<���H��z�eZ�j�
1I�<��l����v����¡К3^lm��	�!n��M{�O��e�k�!�"��"bN؜�"O$Iǣ�W�$�����w���S��D�O��s�{����P=j��1���{�|x{V�D˟̄U24�K4�ҔT�X��CDP�(��:g(I�&�ݱ*�������>�rԇ�,�*I�K�J��f�3��!�ȓ%�M�adT/J�������n4�ȓ�Jt�0o�zB]��j�b���^=�P������[Ôpc���ȓSܐ�bɇ,�����ODN�ȓ&��MJ�� m=j�%)F@�م� �]Y�Fѫp'T�C��J�[@�ȓ?�,�B&@�����1FTl��b3�Y��N��z�	d�.n�B�ȓ9����[��䪧(Ų!xPl�ȓI�@��Q�(]�r�I�Z<��O6�dұk������@�]�(��׈��H $��<1ѧԗk����n�hU�ݢh"69YŨ�<�\�ȓ[�p�Q��L�r��a��_p&ȇȓq_Mb�o˗%�@$�+�# �����<_p�+3
�h�F@�3$����@ua���7���9�'A.S�\�ȓ:����<%�.��P)��(����|��6�Ѯ#���ޠg��=�ȓ-�E�� '��ߓ4�� �ȓ"cr�@�0!{�	�fΈ�
@�T�ȓu+�,J�$��P	�)+vN6Utz��0܅�P/ٮr�\��v!�h��x�ȓ^��`�$5)x,�N8�f�ȓz� 8��O�]1l�RT"�39���ȓ{/������-��$~(�ȓi<ش!ĭ�_<"c/ק!а�ȓi�Y�&T�w�^��n�%4P��ȓ*�f�K�JB�$
��R�ĩ�ȓx?�W� ❩3 �.��\��`�Y Th.���)˯vD�ȓM��R��+�:v�Փ"6E�ȓz #U�$ut�A��7-�4q��S�? ���*E��t��Ś���(&"O�"&H�8��U��e)���u"OnQ�A��r<x�D+^�@:8�W"O�h��&Y���k��N+/���"Ob�p����U ro[�[Ά�[��'��'��'��'&R�'�R�'Ӡ���J<OT���ʗ/p�4���'���'t��'�"�'A"�'�"�'�4�Q*J�$BLc񧆈aR��!��'�"�'HR�'��'42�' b�'���D��'�� �1�u�3�'��'���'���'���'���'h�v��k��<"#��>2\�E�$�'���'���'vB�'R�'E��'�Dm٣��"D*����Y�r<�f�'���'���'>r�'���'��'&����
���`}�&�ȐF.Jp��'/��'���'e�'1��'��'"�����5`�P� �R�F�RC�'Z��'{B�'>��'ub�'�r�'@����k5c@�A�*�-5������'���'�r�'e��'or�'���'��)�ը���e��Ȓ?'�=�F�'�B�'�2�'#B�'7��'���'_dQWhV gg�0S�M��˂�'���'%��'��'Q��'"�'���AЂ��t��!�,�W�'{��'�B�'���'���'+��'u�� coK==�vlz���f�R�*s�'���'��'���'R�a�����O�Ձ��	{����rrgjm(*O��D�<�|�'*7�Z�-	�&z����g�8�Y8W��D9�4�����'�	�"�� 5_OՒ8S�	|���'��U;f�i��I�|��OO�A�&�ۧ�U=��d�aM�?�6i�<�����D?ڧ��;"n��d��PE�,T�+�i����y��i�ʦ��4uu�i�����Kt)۱��
}gJM���Γ���I�k�\6Mm����&���@Ad�p�t��q�q�PΓE�Hx�����'���`��\�#�l%@��Y�F>rU�'��	n�$�M� HKZ�2�i�Ǭ�?�B �B��}*�2�>��M����y�R���V��ctK�����0�GH>?A��Ǩ�I�PO̧ƪ��P��?�gM�i�J���ì��q{�D�+OP��?E��'l�����R�\$�U�g���Dl�c�'�D7��7C��ɽ�M���O몬��.�j��m)'N��-�'���'�R+�>�f���ϧb���"�#e�ɴj�:"��
�.��^�z�%������'��'�r�' ��;����"�cg&�"{T�i�Q��3�44�ݳ*O�d7���O8"�)�f��dAb
1VH�U���D}B�kӠo�1���|�'�ZT��CY|١��C�~0��/�J�9ї%$��ҿp*<y���t�Oʓh��مϋ�!�x�b�H���񉒎M�����?aPB�9S?�-ၩ�3H�0�5�?���i9�OV��''�6�_��50�4���Y'� wh� �gjފ�^��Ğ
�M��'�b�Ӝ *$������?�\c��|;��� y�ڈ�Ai���`ј']b�'�"�'�B�'��OKra�	�
����G4�l�-�Q��'��nӀ�2:����O��O=*R�O?'�ে�8�8�i����O�xlڶ�M��'L�xݴ�yb�'�͸����w0Z|�F�b�uq��øG��z'�E�m�rP���i����?����?yCP? ��K�/G&⌈uI�!�?����?���_�ၣ?�?1��?��i(�TM�q״��I�o �f�)�yr�T.��|·6O���b�0m�;m���|���U� ���Mdld"��,PVX؈Tɞ�4F�TP�U~��O@���+��'�d��\K��u8��V�ʩ��'�B�'�����O�剠�M{� �c}�M*GB�9T;�U�ڄ?`+��?���i��OH��'��6�� /���DY)l�`�#���+T�l��M5c��M��'���$�@]��&<D�	Y<P��q	�2oN��$"�,���	oy��'4"�'�B�'��R>1ZuK����T,�2-��$zSˎ1�M�$�Ӛ�?y���?QL~r�	���w	
M`��G#T�� fJ�0�h�,p���l���|Z�������M�;g��M1RL�(6�����$S�u���'��r�
�O�[M>y*OT�$�O��21f�W0��T	̙t�-#�D�O(�D�O����<�i�1�T�'�b�'g���vHژ2ȠD��r*�2�'��'��֛&�`Ӡ}'���A�'Y:k������Rmz���ɠFi*5�A6+�8��'������T� �'� �W�݀g)�����T��j�'�D�eZ�Fa���� š�O<�oZ�\1<%�I,j޴���y'�U2j�r�@�ؚ[R�j�ѿ�y2�w�o��MWo��Mۘ'D�A��W����5j`�p�5�Q.p���O�T�
@�ג|�Y�����d�	�l�Iş�Jpm=Z�FM��aW$����@k{y��|�xz���O����O�ʧ�?A��)���#��yJA�ͅ.���殮�ش��9�I矼����+��p�Mb�F�2�)х����R��x!�	�u�u���'�B�%�d�'�h��6�I�>���;e�PVd�4#�N��FL޸b��߱2�A"ᦂ�E�h���FbBJj����(�O��l�M�i��a!Q�{�|����0��A3�(XYr��3OR���=F�Y��3�0˓�bU���  %!��G8*mhl�cd�4sn�J8OzB��6#��8�5��i:�i���O�3�|ʓ�?�Բi��M�ΟJme�	�ƅ��Q�vx�Tb����I<�#�i��7-��Pq��g�������$\IZ��Q+J�/N\��,�z����4�'��0&���'���'4B�'\`�[#��#���Ѡ# b�����'��^��
ߴ_^Z����?�����	A9L[���6�ۤ.l�YiӤձK��������	�4x����O�� X�� �.@���1�����I�$��ӓ傓?P���?Y �'P�@$�8 F�C�Έ��'X�l��m��EA��Iǟ��	ן�����	yyB�f��Yk�����;�뚙+��2�n��d��$�O��0�d�O�˓e����9.Bܣޝ[�f������qv�6�Ȧ����QΓ e�q! "�|���	�?�S�o�H8�nO�(�f�QH�d�7-Y�����O��d�O\�d�O��D�|��p��$�%U%���)Dd�@��igL����'gB�'��Of2!q��J�0<p�[dҎ}-~ 
DU�M:`to��M���x���Đ/�V?O��	�g�Pn���5A��[!D�v3O&	AĦި�?I]��'�����T�	=_'�1��Q�l��UA�fDll��'���'qrS��[�4g����+Ov�$�*Q�qFo�'V��Q�T+<?\��ЩOm�*�MF�xB�ց�H��dK�c�J�j��y��'�� 6F�
� �QU�<�S�>b�Fşp���_mQт��[�d�"�K'DϟL�I�<���D���'~�U�C�W:�pj��8��'7T6��<<oD�$�O�n�ϟ�&��(msh)�^��*�#T�P�X�:�M�@�i��6m]<rհ7mo�d��*3F�#��Omh�S4�L,5� \8�F�QE
�!Jl�Cy��ѬxÛ�:�͈-�B�� B��j9,����<�� ɉ�r�%�A��gn 9��=D��&�MsöiD�O�����IǬk��-����~4���A �73�t�#�ԢNR˓[xĨ��o�ֱ��&�	Δ�qR#J5 ����k���Fݜd?:���G�����*�2e@���6"@�BeP�1O�G�Z���ІPW�K��H)�|0�T,�(ކx�3ɉ�jÀD���Y�,�9�O��3���r�-K��M;�_�:�����QîY�a�;�J��\q��PR2 �q�u:�̍��tx��M./(<�,R�	���Z�ʊ��\0��E����C˂�/����aK4�,0)q��D9`��#N4*���J�S�x�T�Տ5&�Ā�eO'ސ�(b� v\���E�	?Y��kڴ	E�Ю�pg�����|�B�JC�M�	ş�&�H�Iş���!�>Q$�
;M�(h(d>)���]o}"�'���'��I�$o mM|����(p�q תډT��P�q��2G���'��Z�<�IğLq�� ��8��ݙS�2^2��B+�'k�ߴ�?1���DΠE�>�%>u���?�؏k�V|s���i����/	�7�<A���?����ş�?Y��ae���4A�US��K'&	��u��_,�E�i�P�'�?1��%��� �nU�4�3���e�B7��O��DZ27p��|���&� � �߽�&�	I�bX�=��ArӀ9�����I֟`�	�?!�L<ͧ,�>]���R�KK�`�S86Ҵp���igt]�gY����ş@�3�	ϟ����ng�*�Xڱc�]3�p�۴�?���?�,�Z}����'�b�[*T����S"	�]\@�j�!����?������<���?a��U�X �뙎`h� ��SY��s��i�2.���6O�I�O��Ĵ<	��Ka�x��ꖓ=	����CUt��6�'���x�y��'�R�'R�:ߢ��4چ4�>��&[�wT�����?9��?�(OV���O���w��M�yy���q���!NT2^1O����O��<b��8%�󉁀[7fT�#��$z�
3c�-!���ݟ$��؟�'v��'6������)�/�B|����k�i �\���I�d�Iyyr��/w��i���4��%��E@)S%v��l����	q�Fyb����O&,ҲHG�*�pu��,ك`�Q�ݴ�?�����ܲ5�d%>-���?�أ
��T���
�8S��D-p7�<���?A��^�'�?y��e���4	F����Z�����&yӼ˓O���i=�맢?9�'eR�I�W�S��;��p�F��6m�OP�N,�S���ē@0�PϘ:�@ L��N+�1m��Xz�I�4�?Y���?��'Gꉧ�4��!�Izm-W~����,E�6]&@L���?9����<q���Ω�tʜ�X?JMP���eȚ���?���?���T鉧�$�'*��Ԯfޒ1�BȘ37P��.����?���&��a�<����?��'��eX�`ҹO�8�Y�M H^q��O�Y��<���?1����'Ɔ����|h���m�z:���Ob�����d���\��ty��')tDk�lQ�k>N�e���Q��̛
#���ן��	�8�?	���z�@�����-C�K�t$,ixi��d�'���'�I��#j�s���qTJɠ6i�(1P5��ܦ���蟨�	a���?���$�x	nڊvW��Y2�ŦgΠ�1F\����?a������O�y�,�|���)�j��B¢G_�4���@P�d9�p�iW����O�$:s. �|��'��[$K�{�tu����$�
�۴�?i)O��$ڦ$���'�?����ڷ�E$3��%��3�����Ί�D�>���x����c�M�S�Ĵ<�@���t�4Ś����'I��T3)���'���'+�$X��=� �)@5� ���eŘ+
�ڑB�Q� �	6Բ�!a+�)�n�v]���D�J۔L{�j�$��7M�%5��d�ON�$�O��i�<�'�?���P[�]��n9D�����+1՛��ڕo�&وy����O�mq���'-��*��H	:r	h�o������|yd�5|��i>�	ȟ���m�t�Pn�& ��ip�O_$�`Y a󤓟rꞤ'>U�I����rȠ����R���r�H�dIo����8##�ty��'�B�'�qO0L3�m�,�2��F�Od0�]���NY�j�,��?�����$�O�db���	"4�2�k�$���d��.<����?��?1�R�'e���DG�\2PZ�d�v@5�R,ֻY���OX�$�O,��?�f.W��d�߃)����HM!S�:�X�KD!�M3���?!����'����!z�d�4ZFP9Cĩܱf��Q��Ԛ	9,��'���'��I꟔�	�B���'��- ��{6����&N�yBv���nm�R��$�	꟔*�ǝ%G�O*����M����%���B�tb���'��	��\ j�w���'�r�O�zͰиKB��SEȠ*�v���*�	ly���O��isLY���U8-> �LC%ZZ�	ޟ�[�B@ڟ`������	�?ᕧu7ɺr���f��*�̹p�"���ķ<�#�y��ħO<Xc��=Db�1�J �7���l��'����I��,��ݟH��Yy�O2���~���P%^��=ð�E�Nv,�Ox�Ex����'�~,+P�V��L!c����� �s���D�O|������|���?	�'7L�3˂=66�A�4�Ӄ,+�	<Hp(L|Z��?A�'Θ��#+n;�a��cHI��@��O@�0�/�<����?	����'��0k@0z�D�!K�>��	�O�!i�M�&��������Vy2�'L*�K�D��?q� )s�����)�J*]������4�?q�r��hc�Ϥ�@��D%/�M���
I)A�'qr�'��Iҟx��JLR"�J>+�
��p�GGp�tZ e��u����p�	[���?A�L�.tj�lZ,δ�A��Mk����đ.J��?)���d�O"���I�|:�'!�a���EԖ�Y��C�?�~<�ܴ�?1�B�'�N �W�V1��]c�p+u�O��0C��B�~ H�m�ߟ(�'���91E�ӟD���?Q᦮A�b�J�e�̶a�*�!����'u�IV6�t4ъy���$*eT�Fb���˟�X�Z�
'Y�0��+���������	�X��{yZw����"��+t�ur+��ҫO*�]Iz��;��i��^�B��b����0QFFS�����Zd�'�R�'��TW����D����_,��[!C�j�z1�����M`O�� Ԛ��<E�d�'�~�P�*�X�P�����l_��7�h���$�O����#y���|���?��'�n`@�K\�� T�pæ9�ɱ8��8I|����?9�'�U ���J�I26o�)Y$� ܴ�?�X��,OH���O��d2�I�&
-��C�&�d@F�@&\��;�ti7��M~��'B�Z�P���>��P��N�<��8q���s�T�Є�Nqyr�'J��'��O����zp��1C�"Ԩ���ᎷG^�8�aF�l��	֟d�I]yR�'�LHk�ҟN���Nh^��5! q�T�t�i�B�'�"���O�u$b2,C����>+	8�sS�z|�h��#���D�O���<���:�0��)���d�z� �x��7!\8(��y&	mZ؟��?�bR>�W��Q�If�����;1���`� 0j6M�OF��?q6'K���	�<��';���	K�,�,C�K>B������O���Wˁ�S�1O��9�`aS%WC�����f��3���?I@Ö��?���?����B)O�n�*zb.q�5��
��	;�~��	�,�G�� j>c�b?IkU�� <���"D�dIV-��{Ӵ���O���O�D矨��|��-�|)"F���Bua�1C�����i2����M������$��QH���G�P⺑Y�\7_,,oݟ��	��@٤�EEy�O��'����-oT�k5Ø$/L2��F��<OD��<ɦ.8C��Oq��'���"H�I�'�U�Tb��2F�"g��	����'��'q��D�&:�ۢ��N�|�R�N[���I�> ��l*?���?�)O����W��˰���#v�<�		��ȵ��(�<����?)����'�bL�6}楪j�/�� ògX
��j ������O �ĺ<���U��X�OpI@�hE���ۂ�#"���2޴�?!���?�"�',ht�%ǣ�M��Q�	�>��GNό)�� ҃�l}�'(�Z�0�ɓ���O=R(�}()r��ȭ&$luG�@�%*<7m�O����I��lK"�#�d0�4�@�ǉQ����,T蛶�'V��ޟp�*�L���'~B�O"�1y�����-h��޼7�F� ��<�I韤HC,5T��c��']�����43�l�*���U���'�2�?���'K��'��t[���$w�����}����$/Ui8��?���ڮV��<�~���R�}��u��՟
��p�sN���q@�
�M;���?����Q�t�'�� �Zؼ6%ޗe���Aר�5�6��]����Z����櫛�A.&�bՁoL|���i���'@rL�oɒ�����O��)� <��de�2yR�B�J
眑��i�2_��B��v��?	��?�dŎ�uP��g��?245)԰>6�f�'#�u�c��>�+O����<���[AB#hc��J�1M@���Q}bKG��yr�'2�'��'&剶��2��,M��؀@�ܙ۾lI���yk�����O�ʓ�?����?A���5<m�a�Fx�ڴ�$Y�-&��<����?����dRL8ʹ̧q�:���Q\6z���~�L�lZay��'|�	����ޟđa~���Ƃt��hC1
�@n�p�T��MK���?9��?�,O�t��`���'ҽ���W6fV�����c8J92�t�����<���?��bJl�' �$�K���f��2ZF9�gH�F6���'�rQ� O�4����O�����T,�!Ck�F�u��H��X*��t}"�'�"�'��c�Oh˓�����b|X���/'w�y�C���Mk.Ol�1σȦ=�I�\���?��O��I�@K��3S�:
����C����'gB���y2P����Dܧ~��ըW���+���l��A�m� �h��޴�?���?��'���ny�F.Yʲ�A#*�1
�.8�W��]w~6͑�-�=�$9��ӟ���Ǘ'��
�9&�+���M{��?9��`�vS� �'I��O0���MV7faL�Z'O�1��-+ķiq�'l�ڟ��I�O��$�O�|S��.�D�u�W6X��]�b�ۦ���<!���4�?���?��*���R?Ʌ�J1s��qڱo	/"a	c�UR}r�V��y��'���'3��'��9x�J �0BD=Zº���b,���.��ı<Q������O4�d}�X�`$2�Pxrj	�t2R��#Ρ&i��<i��?����򄘆"02�'^�J�ɆjȳI�Bu���2#�,<mZky�'4�	��I���Lt��⣮�e>P��ģ�r��Ie�V�M����?����?a+O:�A��y�t��5�cM�o��g(4k�Z u��=�M����D�O��$�ON���9O
�'j���t!�d�#v
��C֌�r۴�?)���ǖO�`�O�r�'��Tj�((YnȲ����#�i8P�h��?���?��D�<�O>	�Oz��h`	�I!�qaV��9f���4��Z>:^��m����Iҟ�� ���� 0���'���tB�
j^�E�A�i�2�'�`Tə'3�'�q��P놀�"|8�2��sn�l�T�iTz�Pt�b�����O ���~T�'��I9L@HhۣZ�4`@p0-2X�޴Rfb�ϓ�?.O&�?��Iͦa��	3��mX�ED����i���'j�e��d�>1+Or���`0Sힰ�H�[D��i}��s~Ӯ��<)�O�<�O-�'�B�ޢq-����?8��-�u��,,�7��O�us��x}�Q�0��My��5��~��,�#ƅ�g�eP��?����#h���O����O����O>ʓ/�V|���L��l̘ n�"j2}hM��#�	Fy��'T�IƟ�I��[�h�,�H�Q�	e~�GM�h���?���?�����$��k�I�'�\$tI�C���ܿ&|l�Iy��'���ɟ,��۟ a#Ag���?%_�e�@$O	$iݒ���/y|6��OF���Op��<QńN�@��ğ�� �����)#H�!��M�K�N��?a/O~��O �$��* �d'}/��m48�����!X�5ӽ�f�'�R^�x@
�����O����Lm�pe�->@�M	�,Ա+��V
�g��I��Iڟ ;��a�'�0��.f���+�'I��J���aZ�o�Ly��U'^6-�Ot��O��K}Zw �U
A�ٳU�"	�U/X(eV���4�?q��WԂd�V��s��}j�-;cr�=Yc��-i����gB���wl��M{���?�����T�@�'�ؙ��a?.���@�i ���$1sld���
67O<�O>�?��I�YE�-��KV4VP��)�7�8�4�?���?y��o�Ity��'��D��U5 ء�&

�i�IF���'��I���)j���?��U58�A�$Ej4��a!�<+T�P��i3���0�*���d�O�˓�?�1�J�iV�O?4�15��6��ml�ޟP"��m��I��p�I��L�IayRIK}��j�^-A�X�"�K�9�`��±>�(O��d�<����?a�P���A�¦�4"�"�SI��c����<Y��?��?�����@�@�5ͧ!��� �Y�[�Fkd
�b�%��IP���	�:��	xb���B�5f�P��8���OX���ON�d�<I3jŒt��O��@R!T$fu�`�7a�nl{@�~�H��&���OJ�D�L�O�=rv��v.Va��כ�i�W�i�R�'��ɏ.�� J|.�M��'oGh�@f�e��K��}`q
�x��'�B�Z	���|ڟ��,�.Tc�I�!��)6�i��I*+�drش}�֟$�S�����$��X3�Hl���^�a{�iI��'y�H��'J�'�q��uBM�K��Q!闆Qkеˇ�i�8�[CB}���D�O���䟸�'����j��2�K��`,�q(M�%��)�4F�������I�<y�z�<�QwHWa�p�Dn�&�:���i���'���@)vb�0�	N?������	1 ISPE�q�T!f��<����?��� #�`�K3|c�m�HR��ŵih��.bO��$�O�Okl��0,lY�e�Ճ}��k���"S�	P�'����П��	KyAY�ܓ��ݰ/����@mO�6�:����!�����%�T�����p� �Mq��N�&�PQYtkSm"�:��H�<a*O����O,���,�2���|�a�T`�@ ㊊D��ѡ�F}��'5�|��'4R
�yR��>�Zq�Y9$���+%��q,ꓠ?���?I(On�H��[�St|��j싈C�0=:*�
߆l ش�?�I>���?��߹�?!K���qaJkLXj�ኩ3p ؁Q�a�R�D�O2ʓ1�n�����'s�t`�?f#����BQ�p�tjp	�3Q��O����O�L$��a��HkS.4�#�ɪ���5L�:�M�*O�<�@�Qӭ������ ��'mzIV&�;�Ν�A�X@{��ش�?��S�N������O����B��:w[��31���>�P�b�4�Ԕ�Ҿi�2�'���O��O�Cx,����=����G�q��oZ�:g2����l�����䜑f���g�=��/i� �ӗ({Ӯ��O���B�6���O��'�?A�'k���0�܇��b�)	����%��#;
b�0��ß@��#R(nBQ:V�g�V�I�Kٴ�?�S�٪��dXJ��'��'K�<z�H��(9���R�8M�$�`�C�>᥌�%�:��'���'k�X�ؒP��,�[u��g�j	��K!� ��O����O
�d�O��4���-0�xl�iA�j���a��{.4�&���I֟d�����	�%�� �I.0�X��
zp`
5�+>�"d�޴�?����?�M>���?Q�cS&�LoZ5���9��x�!�NH"Z��?����?��?I���?��?1p`��E��	+��H[��8���H����'��'���'��x���ēx\�	�#��}@��.!,Vx��x���O�˓5��1&V?��I˟L���0d4��h����D���0qݴ��'��������k���W�� ��zk4�r�ɯ(����'B�S���'�"�'���]��-x�&�6��L�풐\�$��7��Od�dDn7,}d��ɘn�^	�悅�:���Q�ĶC���%U�a��'1��'����'0�O�,Y�'�U�fp@���-M3�X�r�Ql�qw1O>q�	$V1���c�F8a8�(�$-	 ���4�?���?�oȴ~��O������
�I�]�LU(�,�D]�p�/�ɤwǌb���	��I�&���tn�	tL^I��e��ش�?��g�+щ'$r�'9ɧ5�+��&Y�����`����Ьͷ���D�H1O����OB�$�<��́�BG���h�:JUp8�v�.[ ���C�x��'��|��'��&9�*��C$��.��q�GRg^��q�yb�'B�'E��'A�)x�՟��B�,�E��hwC�7����Ƴi���'�җ|��'�R��$��D5NG��;�U9+�Aj�mF�^�I=O�2͉�
UJ�0C�e��K���b��b�b	��t<�fPS,!�Ͼk)�D�tiڱy�
ي��� ;����JІ٣&��Z��0�qg��T�9
D�:d�T��[��{/}R�̈��!��*�μX�ءrg�ŗ>��S$iӿ|� *�1A*r,IS�;K��kw�Ūt�h���g:A�y��e�a��&k@8:cn����::HX���]��`r�d	�4/���Ȃ;,��'xb���Xff{/F)(����e͊��@]�&a����\끍�<�O�1��Z�K�&�q�ʐ!2�@`m�%t�4q�'j��'�*�p�%�<E��9!�0���L�s�(@-ژ�#b	��?�U�iB��?�G���B�VEJí��sڎ��5�M.,�}ϓ�?!�kl�hj�l��f���R��*̡ExҌ=��|��P�T�Rf	R),p ٪MH���?q�cJ�j�Z���?���?9p��4�d�Obe�3�H�K�<iEk2[��Ѓ�������ދa�����ɀ�x_����8X�-I�^i�$�
)U��I���z�)���%iX)�Ac�?�=A��K�1�����#Xr���/f?qE�N��	K�'*�ɱ=/,M��G"j,I��g˖|v&C�I�Q�LݑTg��W�Zpjf��3����?��'�9 �kd��x��Az�.,�s([���Tg�Oz��O�$�4u����O���:/0U0P��YR$!4�3
�z9�fb��e���	t�欆�	�:�<�r�Sd��X�1��/D���g�1w�t�б���)�T ��ɰv�4���O0YK��'t����@�"��y��#5���O�!�5υ5pء�"�F�"�8�Y�"O��dka��i�D�E`i�1O��'w�m�~9�OV���|zC��_��Q�@�	"��`�U�g�Ƒr��?!���U0��!`ʜ0��ƍ%�*����B��e6E"��N�U��)���u.Ri�A��-��Cv'��U��E0��Qr(�fՔTf~ИPb��x�,�Z��)$�2�D�O�?���e���"e��*��ayzI��@w����g�$]�q �%�� S�S	�n��$�g�I���;��7G/�[d%�.!�I�M�Pms�O,�$�|�[=�?!���?���\�	�&�=!��d�U�>0qf��&�(G	��:���kB*��c>�DHh[`T��ֵB@Z4��U�D��"��Ⱦ�*� �8vj�ZE�ċ[/�"|��0�Q�)F*46t�&�Y}�1#n�l��[~J~�J>�W�+O�)p��L�|�G)T�� �؂ӫ
0�;@D�1r�I��HO��@̂�`#�H3�P���`���N���ßD��@�0����ş�I🀺_w�r�'��<I��f��03��ӻ9�1R�'(���@�:��i�b�=O6�Q�/*�n�� �űB^����O���-(AB���d�\8�\zu�Yk���h����o�b|y4���DD�O�d-ړ��DٛWuh�Av�B�o*�d��U�#P!��B�&���j�����ЙFzʟ�ʓ(p���i�����+�+:�bU�۠s���i0�'���'�2g��r�'�)�;C�7��O��g)�%L��� �'8�����'>FdI�U� C�	Z�)f8��W�ޝD�0Py�"�O-�p�'4R6��k�}Cq�
Y�`4�f�@��lZ���'����?Iْ�E�JJ�	qn���}8��+D�p`��,s����VW$հTEv�;�O����)�f�i#��'�d���1Q��+ˌ�3V�	����Wd�ޟT�	ៀ�	̈́M*bx�<�O=�2
IC@���4^/MD�6�I�����8�'&��Br�]#0ƴ0Bp�D=5QGyB���?Qd�i��7-�O@�'k�����L��r�Q���8i�d��������$�>q�ar����#u�]�' �a|B5�dT�!HZ�Rag
�Z$�C���1�d��|5��m�@��c����4-�r�'�B� �D�� Rq4���m��&��,i�bb��g�';P����D�:�Dȩ4�1X�r�s�c��k���"~�I�L��9jЅ�dN:ܹe�%�Fф,�Ɵ���W~�'����@$'� P�YN|ڴ�	�yr�'"�}���0k�r7�Քu����׾�OEzʟЀ*���f�N1���8`u��,�Od��]�y��1$��O����O���C�����?a�N�v�t�V�X/%]���1�T?�qa��r�����ɝ~�fZPhӨ}��2�^�97���u��mCe�.|O�i�˂�����c<�2���O ��J�O���O�Y�l�	ky�c	:=y����`��Ph�Q81����y"�E�|�E� �P��qZ0B�Q͠#=Y��J>�?A*O�,�N�˺�AcErx�!)ak�/bv����X$�?Y��?��z�bD���?A�O4���,�%Q�6��D{����F�mS�p��d��p>�����k:~,��40IT��Å>@�n=�ND�I�l��I��<��Ҧ����M�9���JG�Z�R ��S�K��M�����$�O~��'|�>�Q�NV�0T;Ǡ��d�ȓR�]8$��WLu�pJ�k���%��Igy�Sp�7��O��d�|���/,�#�JD�
���F��%f������?���bW���@��&ul�2�M�u>\R�W?c	 ���1�q��EN*=�$ʓN��bP.9%�$�Sr��q=��s����Ol��Hܷ	LY)G�	r4����ߦ�޴�?-�8�jg��=0���ǘ�S,��4�O��"~�S��8�E.��������/->4��I��ēz�� ��Fۿf�\選y����'Q(|�d�+<b�'�"�O�0�b�'/R�'6M�DcO�xq:��c�Z������]0����:C�@�C��ق�^_�����>��X���W�r���J�ݬW���c@�lo<�P���-f�ih^2�&ܘV��A�pIӶX>��
I�����l�\$�i�>�l���I)�S��?9��J�e��Ё4W�?נ��7j�]�<I�!%Q|p���l�$-�'!�b�' �#=�'�?���3�L=��#��p`Ze��͑!�?9��:wuHiK�?���?)��ta��O����	o:X��F�7j��%2��8|h��t���=lO\5��I�G�(VV�=v�� ��O<��ѩL9z����@���&=?�5��f�|H����?q`n���Ӧ��t�'tRT�t�WD�<nB��pǮnt��d/&D�,9�	��q���a�_�9�<�(�� -�HO��'������oګX�B�Cq"��z��!�4�#� ��	���	���� �����|�R�im�T��4^��ĉSw��Ci��? p��ɴ$��l��Φ�I�S��ZH���-ŵY��)6�O�5��'��6���~�]��j˻6�5�s�c�*l���<�'r��?�{��AưaR�߃-�P��*.D��agkNm9� �@h.��(���k��+�Opʓs&h�FR���	A��g�^�LxQ�E]�ɂP�L*d����'���'L��`M3m:T����4Q.�T>��5�ZT�h��
�	S��ӣ�1�����"Vpa ����3S(9B���?Q�AMKh ά��Z$����!`+���I��M����R�X�v��s��	1/S�]F��O����/2�<����<�l4Afx	a|�L6�� nX�U@��Pǐ���H ��n�P�>Ot�!1̦�Iğ��O��<s��'Tr�'�!#��2�R��3kLin<S�C����"ط�� ���3hF��'�ϿSC�V�s�:H�1��u�PH1��15״�ZԨG�/���R��#�J�/B�:�rX*���fV"EO`Pq6�ד$Jpl�bF ��?��O����O�8` �<D�ų���?]L,t��:Ot�$3�O���\)������O<0lж��9�HOʧkRD���GŐ���ڏt���2���?���+RN� ��?����?�ƻ�����O�p�@�WN+|���
������O����GvN%	f�']�L*�+�^2Ҙ����9��3�'�F=� A�~L�ϓ\b�J&��04��;W�ʷ<4�`���a�����et�V�f��Y�@�I_y�� ��� ���"}���Hӌ�y�nΟakT\�`�/K<�B�*�#=�/��O�.;6��@�O�\V�8[��І!򄜡g�~�K�
�� �F�hS*s	�
�'u �� *@ +2�Q��1��=�	�'���۳��)* 5�͚w�ba"
�'�x��D�� ̔e�@�Сk��a�'�0���Ц&_j���$@�ykP��'��LAh�#<���X�o���'�z�:�EzN~����)e�$��'�>x"�AU��HdN0ML����'�H�Xti�V�-Z3��/=)�|��'�|�¢@�J�dP��@��1c}K�'M��r��s����s|��	�'l8%��d�\������B-zȸS�'��pU���Lͤ��`�
w��"�'�N`7b��~y���8�X���'�� �Q��D��T+��`2�'�tY1��,D� D�6fȠp�X��'$^�W˄*th�$�g�X9Ԏ9��'7�)��tb�g����	�'At��`�Ћu'���SkZ�x0�'#�����fÊ���M/NGP�2�'��	���G- T��B�ބH�>a��'��l��aG+Z��ǢPG�T�
�'K�aE]�0Z��%�=Et0��
�'$쌢�H�j�ܙ�D��&��R
�']~��&μKZ:��&%�t��Y��'�d���F�P�qv	W�Y	*u��'�� ��Ը��$A5�T�{6:�:�'������ "�q e/�ׂٳ�'7P�H6 xp y��\�|��e��'�J��Qa�;�T�S痖��<!�'�b*҃\�Z���PwD�R  ���'t�m!W�X�s�Ե�f�K��x�'܄(�¶tE�a�f�� 9��(��'$R9�U�_M2Hآ�D>1 �	X	�'��)� ŔB>���ҹe@�d���R�RM+��?`�ɧ�S�3K�!+20��y�U��_�Ҹ+�H�}؂Us�O�x�Q�H;f\E�7��K��06"�,
d�dXedT����gϜ�(}fq�?)��C�azX��JG
p�5E�m����J�%ւ9P�+V�i�l��:X$.űGo���0����6�N��A�B<;tf�X�l��0JB��:~J��"�O�(���Vk>?��M�*�X8hg������P�_�<����rVj�a�'>����7����d�j�8"�ȇȓH��sE��;���B�/ϸ<���L*�a�@�$Th͓~�q)�z�%��jG���; �%��a�tEP�fުB�!���O�V�i�B	�?/.U���@�Oפ�n;O���s�S�^����E�Y�F�+gJ�{�>�\Ѳd�EP'�A++[�ĪE�.O��B#$�e�JX�&,G~��I6��4X~�� i[&/�٘v���m�a�@�J�d���*|Ov-J6��֕�#C/v�\�����)�O� ��}�viA�=QG�ƘV�t�ɵk�6���:O���@�φ�JOx�hZ�=��B�	�WHxkČÜU�<��v�`��Qx��wÄӾ9,ű��d����|���A*�ͻ\�2��+��B��(v��	�0Y��,�gt@����$G��d�Y�+�V�✡�i��;���qGם1����;��P���|2����F�6��K�H�ؘț�� BT��"�n����=��%��-T%ΨO�q�2H�!�.Ӈ�K"]Rt�`�ȇH��=�Ν"=��1򷍟FԞ]�@�̑jb�(з��O�xc@�ɅL���"��~ʟ�i�o�"OFu;�hĖv;a0㕟��r���mmv!�d�m������؊*���Vf���i>RA|+��ês�6�ڤ�ݥIF�!їb�<�8�b���~���O�a ��3T���0�
9Dw�ۂ�&��<A1�Z*ø��i6��	$~r�9V �P���ZÅ�.>?��ɹ#�2B��q������	\�rع�jJ�?���!��-`;�8Z�)}�K=@vms��4��@U��צ)"�K�y4dT��(ܠU��M���b.Q���CKV�x�XA�Ʉi����OTrphF��F��M02-]$�"<a�2��ĠP�O�L�'����@-W�B�V)G1m�|�2�AF�"Z���a*x$�
v�SQ*��=�Ә*}��O�w�h����Q$.�(��{��;�'"�d\�J>��/͛4~��I�x�D �!�p(Q	�/�䜡��	�����Re�c��=���h��6(<�y�#�Yt>��I�vojL�F��5xb�dC#��>NC��ˤi�F�%B��H�D�`�%<}2B4�S��@�t�"7-W�lF�xP��=S,���*zNrɊ���AE���7�B�>���w�*�[Ն��:´��@1�0�E�$���y��ߨ2�,��:�?��'�JvV���
SͺU+Di�6v3���6f	O~R�¨-lfE��e�2^?b�I���'/p:�O�C\�����Җ�y��y��6���ɳ�?9�G�ܦ����¶��>�c,Q�km�m�dY8NmڼP �=zF�͓h����H>����V�'V� ��)#?��b��
<6pD+�'�z�0v��R ���dWT8�L �c֠�|��%�64��i��$�f�eŗ;������@�l˺+�I_������\kd�)��R=����w�se�SI�|l1V�x��B�x2j�D���ɳe�<P*��~�˖7RG����CT�C�<�b�X=A�򼲢*G=�0<1��@���5����%�ׁ<T �#�مx~l�sF�Ɣ@x)�>j�}�g�x��*@��5�ǟ�6NH٦OL�NM�r�r���9IB���>A�h]7l󒅐���@���CN��%gN|��+X�d9�}#�I-j�Z	�;��I���"�Р�%O<���.����m)�P���2V�i5�����mB�%*�FJx"/O��y�$ث-f@��&ƋQ���2�A̛\˂��aX0�ʈ	M��;A\"���M�q/�I$1��OԜ�	�+�睔j��(��ҧn�����H�.m���B��-�V%�y�.P1c$ˋ羉15���Q�йo�
&剹Y$<���!���3��ժ3_ę�A�>�������� �ҳ7{H�ٔ Y{�'m�<�uM�b�2	����>R�6$BҦƣ{׾9Ce��)�`�#�0n��;5�����'�� �r��N[X�\�B�^�9�T��1?��9��,:?q����#��q��I��h]��'�A?�e��S��*�H%��x��%S��Xp�W"�y���7o#.�@l[;��<BtŒ�?N}�2��I6��1O��������,���w����ႌ �Xz>��N��!�D](@b��kgk�d�ru1CL��]TT�"
�<����vP�|�<!0*��--�aE���lm�=�b	3#M��J:���Ҏʣl��1E�DlL�i~F�"W䕟.��B ��x���z�k�2�����ާ�Qn�grN8V��yU���$�\�Pe�is"#��0�S-�82�i�G2�(y���Y2�f���gb�&d�֙� *X�T�:Q��$A�Hс/s��0�Ƅb�Q+��1���
�>A"�R)H�d�H���,pȘHaF�SDb���B@��@������O0�/%nn@��n�?Fy�A/\��O�)����݂0��?������ic�C�C&h��D�גJ��87gƈf�:`��8+d�,�"�H����kg�S@�'�h �G�6+>�$�Ϟ�Gr0�����<8@�fK]tq��8 ���yB�k��%�ǎ����������9��(u�R)��ȂF<(�Aդ��7���Qq�'���@��W>>��S�B}"iX ��/�yb�y�~�cP/��A`x�C��w~���U�)&�2I�wm���c�Ej,Cs�+u��-q�c�X�!So��r�^�;d�=/^�%��jҏx��m� BI��f����S"9���E�܆(`��o޼$��b¯8t�l�JY�GHf�C��Z,���A�J�J�u�L�'5�� �\��|�.ɗV��-ʟ'�P�)�2����#N�{�,ZB%ږe��˓x)Z��	�(ۖD��\�i���?i��	�/�YR����T[U�ԆZ�1�V�q�01u�O��LlΓo��XP�	�U�U���AA�o)f�tb�@�"\X�a��� 4t��pg�_&�)��	�_`�S���!8��:3#�0/`�P��{�<�g��7;�(��Ư�(���O^��觿kc� -�������v���x�	�x�����	HH֔s�	��==;�ġA�֤3�A�Gޘ��Pc��P�.��xbH��)��o��=���T�Z���h��M��ݒ���8�!��	D�b�I"��s \��/�O�"�ɛ`zp��IL:R �<٣�
k�Dy1�5�7"���Ӈ�Ґ %��>MՐ��<�Ѕ��Ew�"��U��xƭY�N��)�G�0�a@O�'\�D̓�� �
�8���ߕq`ǟ�&�l�BF�%.sJ1ө]9G��8k���$��P�6���Ҧ,��4|p�+�z�������!pv�]�E��<���;]\=B�o�w?��k2 !4�@�m�^�1��aۇI`��	J-��<��i˧h��I�Jo�? �}�ARF�ԁ8r�:�v���΅E��D�cW�I��:i�B�?Y�GaW?j`�]ZP���Y�9"�E�OR�}�� ���@�t	�/-��3�(�&3��D� �T�d�6iM�@�-����C����06�a�R�6;R2��EI]D�(���i�<Yn�UV�s�)J�X6���aV�[�i�W��r��Р%sʹZ��9�>����$�T؅*��]Fd�S��S� ��pH&�^� b���L>�?YUcV2R��TM,mKf�NɆ�f$!��݁UD�вl.za�m�'�?�O|�	�0�׎ �l],3YD kA/%�8��#d�.Y@�yB'EF8���w XiR���Wp-��'�;dZm���o��sq�'�ҽ!D��}HIu��Sp,������$�&	�e&ЙL��hЦ�O ��ɂL��\�s<�a�|�d�O$f�*La�g�%Ia�-N>
&�E ��6R�fyp�,<P��E��_�|��A>=�L� �LQ�15pD��7+����7�D- JWW�aأ}b�'(��HcÁ�G	~4(��&|D�a��J�t��y�V�6��LP�O>�џ �F�3&�,h��ޤF8�����)T�0a����?��Lh��P�8�>�u?�Oa���h�bO��pH�Q����"KC�(�K��	/G�xB�M�.��$&m޹��̓\$������=Y @8V���m^<�A�O���	ґ"]�L�f�,^�ISF�.���D28�Z�J�j��%@^ұOp��ϕJ���Tbу�(���'�d"+ ���gS�D�p��'�)��� V��8^ $��;^8���I�<ɡI�so�\rC�':��8R��\��2�n���|��u ��F���OU�N�{��a�9Se���Q�źc�A��6��4M@���?A�-ީD���0R�ޅ8b�U��-G[�,2�l+r�R<q^*�⒫p���S��SP��B�gźl6]�`��0~t��m$��xrE��6K�d���i��e��J<r����3q�k��R��~B?O��i�hH�="˓b zʟ. ���� i��hъL�n�`)�h����'��4�e)ҕB�H��T	v1�82��~b#��>Už|b�t,��p"�"v���Q�OXU��D�+��T��1��B�'��9J�j����,6��ʅ`�#~`��P�I5<� �Ú���]3��I����O�'�_�	-Q&� ����*�p���o{��(e��yA�8�ÓU[N�S�A?!�.͈��ԙ5��yZ��DE��Q��îL�\���O��'J:}ڑa��7c��rV:� 2nL�r��}R�JJ�}"�$T����� �y� �Z���3�U�y.�YAg������i/��q��
xc�A
���b>���`F�2�����=[r�a��0۱O�%�"�Ք]m�����KPld���=�4�de�z�/O� �"���عQ.� ]�ώ��*m>�x�'_�`"�$���-L�Y��_�f�rȂ��ՁcI�U�չ��t*�%��^b>Uj�Zs�C�'�����B6�� 7i��R~8Ey���?Z��aQ��Q-2v���I�L���KD�(Ց�`�+:�d�@��`�C?����V� {����}��&V &H<`�	[�ѹ2��`��IA�Y������=2t�I���j��9˅�P��$Ɋ{��H��$Ο��O���M�CNí%�>%ZeW�M�M���V��Op�p��M7�]��`Y��6�	0'���8<|��h`+�
.�m�CS��;}"/��J��i��ȣ�ۊ[�}@ 3D@9z0�k�	Z�Y X�4 ��sS��4���e�gy�O�xQa��v��L���Ƹj�<��5��d�=D��T	��,O�見Ic`l�F�R�>�"(��$^�n:��0�+�.��U��gyI�>	����Xyn��V��R��l�����P���@�&���dO���;B�εYd�S�K�	¼!�2.^?!7�0��cT�)��i��-� Ew>�p�$��H��%"O�U���Z�$,9Y���S��%�p"O�8p�
ʂ6�� �SBO+.�f@�""OE�!�� +Dc���5mѠw"Oh�Q!KF�D��f�[WH1��"OX]���G�9��Y��.��&[r��"O�0��O�l��P4K��+M̠��"O~0#&���(��P�Xl-��"O�X'ͮ/�(�ZT��:t�6"O<<����Q� � e�G�"d(؁�"O��#���Y�L�r&��tcnq�""O�� *B��9��I]�/_8P�"O�`�ӣ��<����H_�EI�� �"O�xfgH=8ْ�		��H�K?D����"�3�8��j�\隭�/?D��A!O8f�V8�H	�zf*��A�'D��y`*	�7s��K�����D��	'D�8�G�
��Ͳ�`�#��A
ǌ&D��P�߰6W.��.]7f��)p�%D���F�^K�@��Y<rP@��	#D��
p����t��!�J�Xp��&D�� ���jO�gbHUr!�H.(�dj�"O%R�ñkz�U1'n܉
��	W"O�	P��F&�p �$¨�W"O��V ��bj򅑲���2�"OPQ"6�W�������#�� �p"O���w*��R=
4`A�A�$�x�"O"��bc�`a�P�X�(p�"O,ss�
m�@}StA�'i�A�"Oxt�3�]C���T�ܦ9M�	�U"O�4P�0'����R�խ#�Hp��"O�ԫ�,�3U����Ǟ�&Z�l3�"O6�t��$s�0��fNV�^�b&"ORX����'��j�A��Jm)�"O�*d��8��Z���L}� �&"Oa�B����!j��Mo(�`�"Oveq�iԴ��M���S&L�2�"OgÆ�ِ��F$ c4"O�D��ĒY-�iSR�V0i'J(B"O $�)j2ZQ� �ȕ
���""O���0�%[5n���!,zd�J"Ob�s���S�v��4Ć/8�V�'"O�����,̰m��"�t�� Z�"OȜⶬI8C0Q�����2��u�g"Ot=˓�ϖ6�hi �fɓ	��L��"O��R��NZ\,CF:�t(2�"ObyѲ��q(��坒*�PY�"OJ1$�^�\��q�B�xup��"OxA�p�=!��5q'�&>f`x��"O�LiRǌ@���*rDU1oj�ds�"O0С�̃k�ܓ��.�ٸ�"O49��L>��jĨE6@�mɢ"OPme�3 $�k���!�<��"O�����A��tH��z�Is"Oqjc��(KU�,�t�·m�z�3"O��9��ܻjD�
�Ϳ$�D�F"O 0	`D�:*���&h���ޕ�"O
��b�:y��#'�_�����"O��!��X9")�B��,B��"Oz��VK�#iN��W�A@@�"Ov�����%>�U	"F�k��Y��"O.!���Y�cˬ!�r�߻!p	�2"O��{@cH�`���Q�@I�:fH,05"Od�`%
:�C�O��P��"OT;�Ę�l��D�c�U�p	R"O�����,PD"v��#�U�"OT� ̙X��=`a^w�p�"Ox-�����;}n�@��C�UZ�"OD1��R m��h��R�   "O����D
aN�E2vf�l�M"O�����$ô�J#H�1O����"Oh����7�X� b'_�)�浺�"Ob�c��?$Lh;���P(��1�"O�,[�'�4�fQ��%Miv�Z�"O��P���@��qK!cӋ �E�Q"O�,#�I[��e��b( ,���"O�����>d#B(��gQ/�Y��"O�t�GI�,e\3e�s�x�x�"O ��T!nI���)y�@�J%"O"AZ.��Hp> c�����` ��"O�h�(�,Z4b��'��-���`"O�Pà*�Z,J��ch�#X�>iX�"O�d	TT�I="5T�k�R��u"ONY @C�(ȱ'� [���q�"O�eH@��a�`9�2��.'�$�aR"O� �xy厉1nBڵ3f���Z��bD"O�ux"dԥO�hub'��7S���f"O����	фL3\)�6��*�f�h�"O�q�e�e'��v�	-�u"OT�j�)[:f����ѡH:\���K�"OH�s���!��-�+K�H؁�"O�DA�.�B���J݊:��*"O0$�W*��j�Y���'u&ժ�"O�����S�G�\��X9I��"O�XsQ�!w8�#c)�
Ֆ��"O�5�M�a���d�@5�v�	l��!%EҶL8DI�d��?O���5�3$���DI���� E7=��L��B�,�yƳ1�=Q�C�2KL�c�Y8�yR
� �
d��P+�&h��$Ø�yBk�e��*j��q�lt�H�9�'�ўb>�h��E}�\�R #(� ��#�;D���QI+�ycC��?R��T�k9D�8c�-�I7\��%EЩU4�ԉ�k8D�x�6ˇ����r��)=�"#��4D��PF�$_����F�F��Ĥ2D��X��K�W3��	s�H2WM
���/�Iq���u� ��@l�&��*g�MI�|��9�~�8EX�b��)�ƀ֖l+�P��Q��y�@�F���s!��2&�}�ȓ7�vdp6K��|RU��j��o�"%�ȓM��Up���:���N�>@X��%:�0��Qa~�p�\�"�J؅�U��b��S2L��&@��f�ȓ�ttȕc��1pVusb�Ǆbꔩ���g}���0��Y��F<hx�`"Ucύ�y�G��-6��ҳ	I�/?X�:�) ���'��$�����<��E<v\��R�]�}����"O�Tؗ`�=D�S�v�@�8�"�S��y��j_f�Z���jD��"���yK_�g�TI!�Խ{�(�����y�"ڂh��9Jq�F�nn���aMA��?i�'\��r�3e�����5��' <�(r��y0��l�ij���'Y����CA8W��+0�˥�pɲ
�'�.lb�� b�53b���!��k	�'V�\Bs��8V,F�r��vl4��'��,hD��[�~0@1�>n�Z,{�'�z��$ȍ
0X�pl7>�+�'��]yT�*�@�
q.6ꮙ�
�'�" ��K�ipa�(�OP�B�'�h܋f#��Q�:�i�j^S����	�'�������.s9T��mD�NV����'1d�ąJ WP�x6� �xH�0��y�iڄ1���s#��-�������'��{�B� jY����"�fl�B%	�y�/[�3�L��\��8��Ɨ�y�ꆄ8��و��©[�����Җ�y��@M� �ьX�"<�d��y��)�j����,�l�w/Ǆ�yRjBr��e剴�|��8�y2�L�.PT�j��]�k���GC"�y�e���ju���R���I
*�y"I�"�I2�υ.¬�&^��y��&f�����o�|P�h�=�y��![$*q #��j��Հw���y	S'9^��{�H.y/�MK���yO�V�ƍ�1�Z�]�Љ�!�
�y��N��`�!0�@�!ﰼ0��
7�y
� �ZDg��LyF��F�pE��"O�U���qx�sD��-�$̚�"O h�!��kn�`0c�?U.>Qӑ"O��*F�M���T�� <A!ca"O��c��(������C7�Jh�"O�D��& 9���!��A����"O�cAl×��xd	�� ����"OzT�!
Y ����ũC���"O@�!�\�j�"(��n:b��hy4*O�eې�B?��v�K� ��O������l
ve�2�J�<���sh��!�O8 �H�Y�|�; ,��6w��"O9+5�&a4�z�	�Pԁe"OB����X�1UPT�B�H�o�n]�'"O��/[9z{�u
3/L�^U�*O�3c��Z,�F��'ڼd��'6�H#���$W���ɡ�ɱ�:U�'z|"� �D߾њf(_i,\��'b���k�#Uʘ(� �^�P��0�'�,ɡS�T�t\a�E ��ڽ��'_}�Ƨ�@���N���)��'��� 'C��h֣�/K����'Z�cGK9��jt� ���"�'�"y��U&|���0��"�'U�Th߈9�8K���<�2"OnIs�7)�����Q������q�O��]�G��D8���l�:R� !��'���8�iX�~w��P����A��'W
�(v�Gb���Ƽ��'\:� AK�-)���aՉE2=��'�y��ũ�2Ai�6Ob~��'��Qz�/O;jMBѪ�JƝ2�����'�Ɲ0��u��p�Ů�/$��Y��'��m�aӞ�>��N=#)B� �'�b�bȐ�i`D�IG.nlɪ�'���ru���>��ŒƧ\�j�x�9�'�ڵcD�x܄�IQ�a$�Y�Op4Z�C�*3~h�#0K�! ��}z4�d.\O����;����!��"g"O���M�9d}!�L.,�xa�%"O(el�m@*����O7!朱q"Oj0�4�G�l��R�m(�॑|b�)�Ӝ=$��q���7���'�4	�B�	u��4J�葃h.\��&@�Z+�C�	��rL�� �`k*Yhpd�� �C�?&�p�����0b�����-rC�I�aH������5g�\`3��3�\C�əvmXD����4*��8�$�Q
^��C�	'C�`x�G�g��M�2Ώh�C��2RB������+6L"���J��B�	�51FA��P	>��P��E98�B�2Qj ����H���RT���B�	���	� G/�y2��V�V�fB䉫L���rɇ>FѲ�)�J|F^B�	�6K�)�W��D~��Ga :Q��B�I8��x�2��\$P�����x�B�	�E��-P���J� ���P�B9�B����A���ҟrʶ �Em�5��C�,/�Ȱc�+m��XR�^�9|�C�	�-����çP!��0��� BB�I$/D��5K�(j�✩��B�	<<(6��d��.8u.�![#Ay�B�	<@���:BHа>r�{��b��B䉰&Fh���`���J\�:+�B�)� x��ƫ�%�ڑ	 唗AՎ�ے"O����&?�R��'�A[�q�G"O.��E�ڧYm���°a[jaH"O����8vN���M�u5�<��"O�!�A�%}2��JQ/1н��"O���腯M�d���	� ��"O0 x��C�i�Q��M��@���0�"O�e���;��i`�N�Bܠ�##"O����N1!�ִh4@	!�6X
�"O�q�pcȫ6�h����.�X[C"O��������ꆏ�z׮ȳs"O���䁍F\H8�H�!�
�+W"O\���CO��*��ȯX���P"OD<*�mB!Ͼ5�P��#�8|��"OL��m�o�Ԥ˵�� cǢ�*�"O�E���.D�L�  "��,`1"OҘ�/̑A��YK�Z�e>A�g"O<Zr�	? "<Z���>^��zb"O�T� &�.ː���6Or�C"Or���#>_"���)Ȁ�B93"O����s��asÕ26��=�D"O�ѳ@�ϔ/~40
q#ƮBFT�+�"O��YO�]����0-��	:�D�!"O�K��e3�X��w3����"Oj�����Z�cƮU�$!���p"Oph!"K�d��������֜²"O�
G�)|!�Ƒ�F,��"O0U� ,���dP��!@��P�"O*Hi�L�[�r��p��b��B�"O��	!)�5}?��b�J�"/��x�A"O�ܓ�A[31Y�B"I�Va�E"O�0���M�=s�U���(�"O����
+��Ѡ�̈��"P"O�@����4�h�[�O�B��u"O
��M(_/Xp���(X"O���ꙊxӾ)�#�;=�l�rW"O\�#U�ā�j�)�H9C�C'"O�t�b�?H,�JVkI	9��m�"O`h�e�w��@٥K[7Tnv�S"O��1uIP1-�h'M*alt�hs"O�M����I�\���޿W.�x�"O���ӗ)�)?��Xq'ۦwG!���i��BL���*@���/[�!��E��-"��X1�,x��Fp!�D�+�\9�̳5����6lO�V!���#�nвP,�-�B��3j^,�!�ڜ.H�XbF�|m���S�F�W�!�D�Hذч� C�p9���đy�!�Ă�EA�D3�cW�w�8�t��g�!��+J��4��;QDr���nЙa!�,��0⬛#d��0�pT!��G���TY�˴U^*�H��a!�Dª���#�ė�iPx)�5Ξ�GT!�$�	*����N]�AA��3�͇$X!�D_:װ9��)��j��b����8�!�$�L��l��kG���H슂
4!�D��ߦp���8f�l�%�"t"!�W�
^Nm�蟩o�pM�kց!!�$C�����P+P'WK:T:B >j\!�D��9�6����"d��W��7>!�$އ6R�%���(<X���+�1>!�D��A�۪�PF_��k�ϸ
'!�$�_i�� W��x(x���D�-!�$<	�<�iG/�g�tQba��!�� ���V�ق"J��3������T"OX�je��jr�رpGݨ$؂���'t.QK��8$켉����M�]��'
f���$m�s�C�:	�X��'n(X��K- �vD�s�ȏ �*�d�<��")F�z=P���j>ms��N�<1�M��L����u�O�L)�� e�<���X5��Z�[
e+����@Z�<�D�3g
԰��_�Fm���O[�<Qt�2UP�@R���%t�A�`�M�<�w�oO���Q�I[TMB2hAD�<��͓�'�I���� ��S�W}�<�G��+fD�xvn±P��x��j	b�<!$i�
i�I�#�x砐�@��C��5*n���ՏoT���d��E*C�I"U"�|P��\�T�j`�1�ŁB��B�ɬh�8�
'�&"�r�r�O�$#"B�	2�.���J ��j����+u�<B�X��������)�T!��C�qj|C��<���b����`t��(mx$C�ɦ_|��C��P-3�4L�W��O��B�I"<�q;U
>�RHSIU
Kk�B�� b ����c�6\I�ťr?�B��;zd]��	W.���Dxq�B�I��|����YL���M�?�rB�	:w����@��N�(���j-\B䉥}��j�O$�"'
Q �,B�>'s�L��$x0D$�[ �B��=v�*�q�`�:[(� w�Y�q�C�O������(r�d ��\��B�I> �XA(��&1�;�m l��B�IXk(4��ۦ<�mj��Ԛ@�nB�9?O�$�b��`�NQ�.H�m�B�I:Ov=�� >���7��=tǀB��0N*y�/�eM���"� 2�vB��"d��!��
�tQ�b��f?$B�	�p��5`Ə�\��*��K�u �C䉩:����=���@�Յw�C�	���<��EF8{����0$S>w�C�I�	�5)q.ה3L�:6�Զ��B��6}�j��fI�٪�Q��2T�C�	���1rbG�N�v-r!��?LC�C��2ri��s�����*���.�pC䉆v1fa�h^(Y�<=Å&�u�<C�I���4���DO�.���H�	q%C�I�Mt"X����Y���!���B�	3\��Dh�	�m�5�ad Y��B�I�v8p�"�(
=&/X�C�
;��B�iif��\/�)y'��5���R"Oإ�u�6�bQj�F�OPn-y"O�$����+Rvx����!��y��"O�D��	B�|�.H�NL�w�,�"O��Q��
j`�� 4Lt�W"O���*2?�)Sc��V��t��"O:�` ��+C��8w*��R�"O@C���*VTXi�C�����KA�<�G���S�D13�Klh���@S�<�K'[�<|�v���^`N���#KM�<!@�[o/r�u�=4�R9�˅G�<��.E�$�F;�%Ϡi�x�)�B�<i��Z�Ct�� ��]��u���@�<1��=~a\�ڐg
-xV�a�k{�<qu�L6m>��P)] `��M�<Ĥ����wLW��(+1��O�<� ~]Y@N����P��C��P
"O��s��0�(Г'H��k�|YB"O�"�#�>*���Fl��SA"O��A��Ƃ��%�����R"OA" FU"
.�1dɍ�?��i�B"O��;���R�$�+SIQ�5�\pc@"O\0�A,V��|��h�1eE���"O@t�C���&��V�Z�r�"O����h�� i �жٚFў�p�"Ol]��� �Fe���Q*��p"O �3DtZL��B��K�4 "O 	;vχm��\��'W�(�H�"O�Ir�4]�Iu�ށ%Ƶ� "O����6~���ȵ�P������"O2X���P�;�vA!�M�>�\y "OZxAbaJ/��y�U�&��i�"O\��"<N����b�?AGv�b�"O�1��@��z��A`��@.��"Or�f�d`z��d.�>F��5"OjH0WI�+�j�┬��w!�e;�"O�E9R�ǆe�(!B�yf�s�"O�8�ƢA�Nрeȡp�*���"O���L�*�X��C�B�]��c`"O�<�M����l`G�� ���!�"Oj��d咜*�2t;C��6�(�v"O��fA���0�	��ŕ�6���"O�\[���:b|�`��L�!%��L��"O.���Β�P����E=s(8�"ON pÄ1E-*�Eɱ_�B���"O<�
����T+u�+��H�"O��#�XO��)I�̥>�
4`F"O\���j5`�2���#�o�P�"Oˤ��MT���"�3���� "O©�bᝆ/ �b�׻�dXQ!"O�" #Ļ>hR�f�
"�(D�r"O�`HÍ�0o�~��Q��*߼5!�"O��C0/S�w���ڔn�v��"O�s2K��y��l���A�A>�D�R"O��C�54���q��"$,fQ�Q"O|�����?��(D��T ��"O�@9֌>a��U��IP�hŀ"Oj���/Y�����RX��`"OVU�e	S-p��;�愗6'��"OJh�n�#tP�KP�O�8X�3�"OX�ѫ��e�� G�ebN�yB"O�yg��%Y��US�&P�Z�
=��"O�m#�bBn~y:��κ`�ԉr"O����#�t��Q��*�:G�x���"O*�a�űa��c�gH���#�"O�lxe�;�p����07�mC"O�|Y��#ӰI�Qe��\J���"O����:'PFhRFٟH�X��2"O���E�u��aJ�C�1`p� u"O�#�E�+�h�V�ӃQ2�X�"Op�s d�q��ӣ��	��y"O��8THC;E�J)Cd,H�M��6"O��p�a��H�q��� ��"O6��슨q�0	�h+O����"OHi�A�0Q�ĭ`a�V)xT#!"O�y�fH�>qt��x�G҇�|� "OtIR�@�2���ɱ%��X)�q"O��R�ѹ]f���� �"O�還��<��#֡Z7����"O���5D�1Qe�&.0��W"O� B�
��[�b����ղn�+�"OJ�35��&M���S B�g��p6"O
� �B['R�E�b�
�OU>�0	�'�0��%/�� h@P�3Z( ��'�DHb��4j�8@�g��a 	�'c<-P�UD�����+B S��Y:�'B���!�)a>� ��3C	p��'�*(�e��T
LӳE҉z4���'B�a*��G<M�u�W�9H6Y��'��u�ͫp)��Y'my[p�z�'�$·��>C��1���+ *��8�'��1H�m��5�|��Vo�7�a��'�hi����� �RY[��@5e`��A�'����Ge^�i&�)pHǤ+�}
�'������E�M!�T�e���+5v��	�'z�k����~覨0$��vI*�'M��[��%QKl;3O&$�<�
�'�=Zai�	 pB�I����(�
�'��@�J4]�~\�a��ݦ��	�'4�\0Q	,q�4�KQ��=t���'*2$�d aU�*�H8����'��T	˖�4]�uÉe��I��'���Q'�
�`W
���ȟa�dՊ�')" 6o	�gO�<As�J;Rb��'��Y�R_�0�(������'���š¡���r �n̨K�'$�tIt-ȟ+~P��-B.^/0��'�t%�0LJ*D�8�hV�J����'+�]q0B	�Z��D�(<J�X��'p<
���1�1����D-Ɯ�'J����k�`�^�?��a �'9r���T&bP�V��6�z}��'�(�aG��N}��9���7N
�8�'o��&��E���+�mϥ2'����'K�<�%I��e��{�C�.���'l��Y��:o�٫c�\��	�'OZd+"�<M`�ۗ�TE���'Y,a��J�4q�x*7IN&�~��'|��Q���9W�>�{���..����'٢�����V�E �
�8	�P 
�'�t	�I\"&��qG?p6��	�'d��^�~5�� *<����p�<q�Р�R�fM��*Ӯ�0-5D����E���h��t��3��q*�#2D��k-�O=��	 %Ρ,4��V�/D�0�H�^�M����!>�Z��1D�@��g�#t犱B�	KL��'�3D�d���Ԣ�i#&M�OF� ��2D�D���$ܜ��l	-��b��1D�`���~x(�����/U����@f1D��Q7 ��8 ���X����2�-D����M�����pV�p�D3��*D��ⰋD�S�  	���؜"�I%D�R�A�b���MНd�=�w�5D�Ȁb�F$Q�,�$H�>04��C��/D�H��(��I��u3&��x�4�+"D�\�FOK�7<�aN'��x ��<D���f�S(Ᾱ���
=��P�>D�T�U,S3_��A��2��%iю=D��:D�Ӝ$��@%Aț�e��b8D�P/�L(�%c��>%�l ��٠"fC�	���T"���d�$Q����TC��
�\���f�-��l4�Вwp�C䉏=�h�2(I��0��Z�&��C�)� @�Ȃ) ɐт��	�4`�0p�"O$�%C	 ��}�P�G���)R"O|������@�h#���N��""O�t�dG�aOb������ɣ"O�0S�N�c��hr�M5@��Cg"Od}ʐM*o��$is�T0ԅi�"O��7H3�T�:�jq����"Ot���(=�����T�\� y�A"O�l2e�a0摢�GМ/�ꌂ�"O"��)JA���QU斪%�驤"O��k#9k,t�eЅd9�Mx"Or��	�.m�q�����m8�١"O�ZA-6������N#�q1g"O�	IF �
Q��	"M� �d��"OVfD���#1kA;rB�3�"OX�d�$R�]ұ� H��"O�J�B	�l04��'�/AK�	�"O8
� 2;�a�ŭ��6Ke�"O�����+�d:E-Ц}��]�#"O��!&�ۇzX�y�,�
��"O��`ЦS(B�AbeÄ�H�c�"O��	��v�Ve��cÑLƦ�"O�h!�!�X�%�B������"O8��4h�)�<Ի@ѻ3��"O���C�����A"a �h�9�"OJ�8�Sak"L��ƴk�|͋"Ob%�.�\�����0x�ɛT"O��yPᕓ ��)�Q/J���S�"O��5�߹n�.	yt��9��9Ce"O�BDL�%�
����R�vN����"O�����>x�"k=$�
�"O�t�"�Hݞ�2�J�, (HHPE"O~u��@A0*ڔS�邥cu�ك"O���֤9�^�)G��?���S�"O�cv%�}���ӷf��ё�"Oa�wm/0�z!�-2��a��"O� b�lۻDֽ��%
�P�p�q"Or詵(N+-@��Ǥ�7�f��"O^Ё�K�<~���%2)�Z�"O�1ҡ�\&0̼�[�d����x�"O�ejU���\�fՁ1F=�(lhS"O�p�@�X�lp���b��`�  ��"Ov �@:^$l Ă�(0�$��"O:hX�	
�\؞t{�G+|ؐ0�e"O��S5i��x� ;%�
�V��l��"O��P�J�)�|����ۍ-�%a"O.pX@�#�pܘ��B�<ʤ)�"O@2"+�a��@��K�_��Ѻ�"O�����ᆹ4a�p�<!6"O�Jኋ��:yң%�'S�<�
�"O�D��<�c��D�gPذZ�"O��آ�Z7v(��"�d$��"O���a��#m���#a^�l�bg"O:԰3�w=&��.��
�޾�ybI�y#����K�?Ǥ��6��$�yB)�;4~�ň�hU�/�B�4�y�	�����ᇶp(�i[0���yBmO7<�t
!
�z��x7����y�������h�����)��yr��"K���V��B����4�y��L�?��IhT�0�E�u�އ�yB�ڛ���%ÁiW�x��1�y��C+�ZEQ��_c ������yB�Swyl���#�P� ]�%d�y
� p�V�v�5�	H���"O�+F�p喝Zק�V{>d2"O��"ō����H0�O�2oy0m0�"OTH�E��:f�1���K�5�Q"O(�9��14<D,A����y�n�sW"O����@�:u�B��ѩj�}X�"OZ�$']	,��q0ᗽ_r����"O�e�V�� E�b@^�7"O ��%^;q>�(FFGb�E(�"O����fWoX�\�w*X�"ΑpV"O��1��t�>01��P#(p�a�"O��{�d��+6��$E���"O�-�#5V�<Lcĩ
�Q�zM�"O0�EB֤	f�@9GH~�$4A�"O&H{��C�PO\|*�GH3�
���"O�a(�Þ�x�&�&�o���"O��S�Ťd��`$�R4�|Ȕ"OJ��F��y�&lcգM
*1p$ c"O,c4�PdH��fE˵l�N��1"O��pb.R��=a�dT8T��8�U"O@a���^D:eAm�(1I`"OR�(��dQ���A�����yr�M�@�F|��gۅ&]�؀���y"��)I���H��C� ���� ��/�y���]�P�&G�� �����ybe�����p-�x$JЎҴp!�d*�HAPD$d�0����:S!� �n,�"爤���r���B"O������,����(��nu�u"O<���T�Qzn��,T�e����"O\���ÍM�0L#���=�t 2"O�()�)��I��1ԇ\5S�"OD�A2+J�7��S�N�p�T"O�0�F�={lX��@�+���r"Op��еK|��j�EǺi 
�y�"O����<D��⢊�F�LE�"O��{th�E����A���X"On$�r��43��d#��9"�M�V"O��g�С��4�7n���<2`"OV�z������R��R�(fiB�"O�u��)OZ�ĥa��4NU�yӁ"O�hX Er��I*��@�G�>q٣"O^�i4c̄V�xȻ�J 2t���"O���$ئCi�M�D�\���"Ob�p!��;נI8�*�4�i�D"Oh�9V+_�'��{�D�"+�f�	"O���5�;,5�0��T�@�E"O��Z���2E��j�:4�ʕ(C"OF���m�,)�4�tj4�Ä"OF���(R�i@��a��E2d"OF(�B׮8 K"O'jhC&%"�y�� 
-n��6��=p�Ҵ1f�Q�y���W�0��i�#l���"�E8�yRDگe��H�k�^9L�)�[�y�)ǧo���p��?��A7���y�X0}�x}�䏙�K�(@��y2�
�U"8��� H+`�2u�V�y��%W0E@WE�P����?�y�hI,?��j��\����4�yb+t� Eq�B�>O$4��LV?�y���A��AthG�|���+DB���yB���$�>I��]7},���c��y!��F7�E���q��Tjc�]��y�������"�A�W�F¥��y
� �90���"�9DjH�
K0�)�"O̜�%hJ?����5^8�3"Oh��L��΂\��\�ri�F"O\�S�!X�3�rx����*�<���"O�����4%�}�wh��Q�\�"O�aH�N�Ԡ�A�DV%�h	d"O�A(�C)`6r]iʓ!J�I%"O^ ���) ��4dhŹ`�C"ONp[��=fV�l�'�����&"O�!�I* 5�+q%�<R�h9�"Ox�r� F�,� ���N'N��P"O�,xp`�XD�ۂ�Gn�x�Yg"O&<��Y�<�v��R�������"O�M"�b�צ�"��mHX��"O����-
e�P[��/; 	yu"Oj,X�����t���c 0lp[E"O �Q��)��zAB��{�5%"O�ez�L�u疽3d_8��4B�"O�H��ᔍ�8[�b�fu�h6"O�JBG�1��\��
K�ib��B�"O�%��	�rB�{��޹@��(y�"OXB��߿#WXT�6�c��Y�"O�ib��MgN��#�AHv�:`"O�qUG���db��
pV� �"Oв� �BtA'��Â�C�G!��!s1�͏m���" 
֒�!�Յx�\�*�G)hb�yʰ��<[�!�D��E�h��C�Ui`�xa��p�!�� �84癹r^Pp��ED�0k!��Ax�t� ��B�ƌS�C�
�!�d�?Frʑ��N�	4�j�ۀ-m!�¦1�%A�o�'>���AE�Wi!�d�.3�(���[c,��S���F�!���t*B���%N~�|���V�h�!�$Wd�lQv�U�v,,Q�É�!�E:�n:W�Mb�x�u�30�!�6P�dX6�)><`̪�A�,M�!���;�Ph�E�֕G�����<m�!�$A����"���k��R�L�C�	�.rb�x�iZ.N �Bb�K>T^�B�	.h��Ԣk�"yf����mH�
��B�	84�&C&��,�n��kȕ,Z|C�I�Fkv	BWI��z�:)�F�ŧ|&B�ɕh�N�CG��0,��RiC$�C�I"��e��T�60�S̈́6���IP����l����[{r(�b�iS�`���A�5D��P�#w�xx�f�Q9Iʠ1` 5D��"�b&P�h��O�(Qb����3D�йF�!i\�t���L�HNLy�*O@��Ej�Iuҕ{U��)�] "O���V��$~���B�,`Z��"O�I��@$�0m��D�x0ؼ�q"O��0MR;&��݊��={M�D�3"OvL��O݋AE\E2A�<v�P�"b"O2\���À_���SkX��|� "Ont"�kS'�ʽ�r/G�t�ȹ`v"O���ǀD��Zh���T��E��"Onlb�(Y�6�A��؀n��"O؈���?I>��2�ds���"O�pяY/ZF�����O���1"O|�� ��tt��#!ΝM�4�"O�!� �,Q���JG�^>p��Pp"OZ5p�@�OE����"�:�	"O����2H�&����[7"�4Q¤"O� ���F-M�8��I�8v�y�%"O@
�gL'������D�n[�l�"O�I�/��A�Z�Y,i���r�"Op��28�3��|�nX�p"O�u� �G	νY!�T�M�rHSP"O^A�V�˘u0zY��,��rY�@n"O�}�"hɃfsv�{�!C�#�<��w"Oh��� ȉ(a�R���"s.܅k�O� *F(��\q�s�+]BL�J��O*B��=>����_�Cx����,�B�ɸNo�X�$�E�@v(Rơ��|��B�I�}� �W(-j0�$�ƈRcpB�	�c�����%s孲W�9c\�	�'��C&HB� �$�ևD�T~�-��'F����N>d�\h�փ�Y��!�'a��� ��=97�� ��^��~�S�'�D�� G[�gEL}�e+�$J����'�X�C�+�7k�Z}�u��;yO��;�'���17�.~6^�,�u�:�2
�'�N����S>���F�-q΢t�'W�x� (}k��Z&fb� ��'�ũ�ȃ���<1e���a�<��'���*&F�3<\ �k�W�Q
�'6N��g^�l�/�N���b�'`���#O�;Wh�����B!:zf<�
�'�F4R1�.�d��r��7m�x:
�'&m�$��J��P�G�S�&�H(k
�'&!+�.�������vux	�'Ͷ����׎{��Ѹ7�X�t����'�E���[�$BǁJ1I��!��'�6(�7�<��VIG�1�'�������2�͊a���2�'����\R��M�'��']�l��'����V�A�`��x·�"	L��	�'�"d
3ȃ�;KP�bW5DX s	�'B��VE $Fռ����@	z��l��'WA
�\ 3�f��#;`M܈@D"O(�ȗ,
�|@d-��$@*�w"O葲����L���bɢO>�C5"ONH��C�;��� $ζ#.8h"O<]�n�
?���v�U��̘�"O�At�X�k�4h ��)-�n��7"O���O�2FA�䓷��%{t�"O�)�R
�/d��Tj��es�uzG�' ��ȟ�G{J?�[�nV�q3�(Y1"�C����&b=D�<��hW�A7�|x��3*{D}Ba�5D��u<�vea,�/2���5D�T��*���1f#4aU6�c�'D�ظG�H>w�"���♼y���ǀ0D���bh�>(2�4:�eE�8�H�@"-D�(���LO�r��b-*�zh�	 D��ڢJJ/�ra�~���f��y���*'��L�t���jK�1����y�f�/%��U����Pi 1��F��y��D���A��M�>�pt��y���7%P�iц��Bw�r���y�,o�����ڨ7�"hH$�y�$S�s��X�-�pY�����yb�.�UQfe�3!��a��`���y�阚Q�f}#��� �舳��W��y"d�p�%흗z>i0`
��yB��?)zƕ`�b��6�p{F��y�
Z�����	Yt.)�._��y"-�NH I�Pā�'E"l�%���y
� �Qf�	�]����2�HIr "O�}ȱ��"~���XWE��Sڌ�҇"O����Y]{�Ր���;����"O���%ѭ����F�׊h�h�w"Oԍ���I� ������Af@�R "O �@��*��F/@	;j���"O2���f�Ѳ�o��_�պ""O�t��[��d��c� 6P�h"O���O�B�X�bD�F'$P���|��i>h�ʍ֟�&ě$c���AVb��z+��ʅm�s�<�瀼/fn�[��!�.�z�+�n�<��!Z=)����1N�"EE@J`)�s�<���*�p0���I'��F�o�<��m�.7��Q�G%һT�hiD�e�<�q���\Ҭ��n:}��q�A{�<�)ұx��"V�E6��hƬ�x��~���O���3q�SX�plC���U�Z�'�$�(	"���%�Y:����'2�{�`�%}�j�J�L�9�
�'��ysE�Y(���cD
�DBЀ��'16��w%��A�#Iwh�Bf	r�<QǪC�Z�@�M�5n��s/[S�<��,6;H���Ԇ[�\���F]I�<Q'�Ėb*�!�F�G��B�m�<q7K���Բ��τ���a��e�<��Y�[M�`RbF�:�qᨆd�<�3GQj��a;ѭS�"iY�E�<!�+�+����	
�����W�<�Ө[�2�:Hs�c�k0��Pŋ}�<���D�I����塈�i���iK}�<a�i�~�T���#� x�T`�Rn�<A�厄ka��ZF)J�LȖu
B�l�<��
,&]8hCĥZ��ȹ�s�a�<�rN��BK�)��	��$N�p�u�ȓg#�qAD�;���{�iR�x-�U��#�!�V��DE�y;������$Z2���� ��c��χT^� �ȓb�%��ꔣVB|cd��* "��ȓ:  K�:*�jDcD�%+���ȓ~�X�a`��� { ꀍV��T�ȓ8B��a���#��-����S��E�ȓY�B� ��FjJ��ǃ�/�:=�ȓX
�("c��&�n(���ٺi�V�ȓ,r�ѳ�EP���!_9K��!�ȓ=�*�;��������4�� �ȓjM`@�S�N�c�e�\�!�ȓ7��5R���<��ĭ�-n*~U��D��.�=��$�G�V,RT.ф�utp���N�;��A���! !�$B x?ƴR��w6����'?!�'Iei�Ҁo2}4#U5!�Իh�@�b@À�t�1��f3!�L�S��s�$�Y&�E�-!�DLW�m�E��� ����&Z0�!�$B�~�p�(ą��2?H#e$��H�!�Ȟ<�Lٲm�7�*5�7c�5g�!�҉>���B�mF���:�B���Py2�U�H���Ǌ�=�:T�!��y"Ń�Ī#��2vD��QR��y����J���ra�s�БV�J��yH��3�Ƽ����y)�8!�
�yb,E8<�X,�ŭ�bF����y�j�>
����	š##�]������yR�Ġ""��&C�
R:�@h4�N��y
� �D��� ?|�+��Ӑg�z���"O~��AW	\M���"X��Ř"O�yW�@-p��E�G��h3�"O\h  �6eW>X���V[���"OlY��
�"�e�_(*C��$"Of�A�]�i���K�3?l���"O�)��Bˍ+Ƹ�0��	2<-��"O��ce
(�;�D��%�U�1"Ox�B�р[]�È)c����"O	p�H��$�p莾-�b$k�"Od�cA��# :�1V�
h��	"OF��C��%*=3�e������@"O�ա� �x]��DKi�xY�"O��8r��)|��r�̗2�Pc"Oz��LA�D"v⛤�P`�"Op�����Q1��b�@L9�(�CG"O�D02�ߨm�N�`��Czv8r"O���s)��A�ub�:��,Z5"O:@@;����� <kf���"OT�:��H'~6����iS?f�@��"O$�3���:�.tS��q~�(��"O�E��!�I�M0ˑ�'��mS�"O�;�Ȏ(>�A���=��ɺ"O�,6A�����S��M,ֈ-��"Oy����(vg"��س.`l;�"O�e�Ι*3�<0�	�!\���"O��`��B6b.b}�ӈ�z�\�ѐ"O쑁�	>2op�h�ᗅ5��#"O�0iWB�d�!3O�Xq�r"ON�J4�ێ@����!�G g�4"OHp"�Z"���K��ɿO���i"O�L!bBJ>~���Uΐ�j���
�"O�xr���^t�h��O4]�c"O�ɲ���=�����጗5xf�yE"OFD�R1J��`?�9�%"O6"�L�=e�(3m�%> �ۅ"O��)K�)r<cu��$*��"O6q�F�!��,��3pH�"O��Est(��L�
���"O�q�C����J K�H��;�"Od���A9q��@����;�>��"O�;s�1z��(�ЊJVXJ�"O�Ƀ�N]m�j��V�[*�
G"O��z!��<<�-ST#T���f"O&���hʴ
v�������C"O$��&��%*Ȃ ��l��]�f���"O	��m²Ll�*Є����"O���e�͏f���TI���L�R"O^��!��!&���$�#��		�"ONac�g�$u�˵K�h���"O��@�Ǝv���#祓I L�s"O^�P�N]�\�͓sE=(.�uxg"O���`+��7E^��E�X8����"O6hP�$~��� �z�V�y�"O
yam�N���$_�\s���"O���� ��L����E�d\x0��"O�hrOGq�}��-[*^?f��"O��AE ++����clN�?L�b"O,)���B�x�@�%�[4��"O~IHf�ÝpR����7%x
2"Oj��5�6;��ӂ��<$�م"OXu�-��`��iB����+�)��"O�X{�%��3!Z���gD^����"O�LCE� 4�;�F�T{���S�? �a�A��F]�y3�&A��a6"O6�0%˕5+@ȓ���(4!�!W"OvE�C�3��l*��˂I	�d�"O|[�"�=.�&�Z�[$	�L��"Oj�V��2!� �飦�%v���"OD
�J�#��\�����%�q"Ov��3"�(q�]`�S��4"OrذRM�U�ΝR�H��@^9�"Of�{A����xq���A�B=Rj!�S�3�X(���J�Ydf܍iU!��O2N����)���)Vf-S-!�D�N�L��G��f�{e��0!�ğ�6�l�2�&<��<��j�>^|!��K	0B�bA��q����<)N!��%	�ի����z#�eh��M<!��T)
/|�Ps�J$
P@�5��V(!�$<YxyK�Ub��yFf�.1!��4n*�:����Jh����߬
!�$�d�puA��P!����ĢE�!��X6ez��-��(Y�C/�@!򤐉4����W�f�s��ӺH!�
�D�H��6I������л�!�K����ڱ��8��E�cόr!�$�x��h:a R�c�f����	�+!��B"CIt�{ED�$�����m(l�!��ܥq��i�RJ
k���JVl->�!��]e"�S�T7g��-�w�ۭ4�!�d[�s��QA#F����]q�I�!��2D��0rD@ �<�F����DP!�So-�QuH�"i0�!D�?!��K%�Q�,J�{p�K D��%�!�7g_��{w�T>f�s�b�	�!��8loޖ
03�r`"ˊ|9���'5�Q[c��>N�܁@��|f� ��'y��6n�[5���H�r�t] �'?��Ҷ$�-�jT���X�r��PJ�'�P�I� 
�䬐����x5��'[�X�1i�g7���̈́M�L��'��m��卶n�
 � d�
@ʂ�`�'/�4P5&�aDy����4�>� �';.\ ��9`>�9���ٵ.��I�'�.0z�������fS�W� qs�'��&"/HŰ�$P�8�
��'���n$V�0�Ι8A/����'/����n�(d͜�RJ�";�Rp
�'�μsT�%��0�a�Η`?ܸ��'ytYv&׌3��I)A(�k�|��'��q���+M��x�p�4y��1�'���R�-P3T���I��L�n;�,��'J-)���
�]𷃍k�1�'Q�=*$��xnU���j�+6D����/F�H�����m�Xq"8D�`�j6P�b�IC�L�Q2pM#D��c)ϡ6	���M��@Y��� D�l8�hO�bo�pH�33
���&?D���҅B
��8�S�H2_�P�A)(D�ģ��ͣj��\��.E,ss4ġ&D�8gHP"<��hR���3D���0D��j%�״z��=S�[-4����J.D����C<k4D���ivP[�k D���-�i�&�·�٘R�l�#4�"D�XI#GJRN.�yw�����a�a�>D��r�kCT|ذ�ˬ@;�5���7D��*V��p�8ApB��2���!D�� ��� o�6l�䘣�G	},��"O�L
2�ػ�l��H�&�\�W"O�LZS�[�k0�\	6�A�,i!�"OX�6��R�^�va�"+$dab"O&��狒!.��qQ�� 	�,�pt"O�]�'��F7D�j��3(�(���"O
��R�3�4���1l��x0$"OP���B�P�,����2]O|C2"O��#
�&}�$�S�6֠Uzw"O<M�Q�p��Z�#Y�x&��"O܅��f�u���jrW�r��dZC"O�8z�/��gt���C�@6��uA"OBSi9%�Ȅ"�<9}Jt��"O��
0�߈������@�"O��BF�V�M�h􇇗^���*O.͘ e��� r�`d��'��X�ǚ�c$��k�F��i�L�
�'ص�ؤ_�nӥ�U�fp��	�'9X-`�E%&:t��%ռ`�J�"�'��D��+Յ]�R�����9&	LyQ�'� 	���-q��}����	g
�0�' �� �MQ9(bn<{$蒺+��R�'��Zf�H�v�͚��\&m��,B�'�d|;�0|:ܨ�S�R<1�L�
�'�N,[A��-P^���F7H,��'��b�<��83�"�t��')�UR Ǖ�v�^������Q�'��q�qR�tR�t�=�J�h	�'�t�`��
|2��R����0�j�'�@u���p���ݠy66 ��'R����R* �&�q��'�
�z��Q�;����4�޹�'A\��G%#��+q�Ȝ
h�S�'[d��A(Y�C����q��8��
�'��x��3N��}�F⎜hƩ�'m ��Pl%u�#V�\-Tyq��'ߖͣj�}�X���M�6<5�ɲ�'���(�(�'#�6@��ߴGN�,{�'8U��h�<�7�h}(�r�'Ő|j�-ʙ3� ��閝����'S�����[+X�DԺAMI2�=�
�'�|��w�[+V��䂵s@Ȉ
�'��*���8;br���/wP���'�,��tL�4��!�l�l���		�'������+4��#P���'h��F���ta�B\i�	�'}�P�-S�8�� ��DF��8�'�L��,�*'�8�hpB�IK�$��'c�4B��όD�!! ���t���'GLL�G#��P�1ǉی
0�i�'6
D�t��A�V͠U�3Vup���'��t��#Ҍ�0q��ѩK����'�Ν� e
�wR$���EWc�-Y�'�pMajD�:��Bh�7nR���'�)'�:h���s��&,����'��y�Á�?��d��Y��q�'�HV��l�	��D��=�D���*D��H��
(����H��[~��GG+D�0��ǌ[�\�1dE��)��j<D�|���@&R3DQ��b�n�zV)/D�,`2fޕ/c�h���]�|+6%%�,D�X�Ɖd�*|�@�+9���!�I/D�t�v�R���w�X,,9|�hq#/D����[A��z��:c�zQ���8D�� ���q1G�p�a��#�ȹ��"O�k�j�-O�LIf�è�����"O>�r��a�a �(�+eR֔��"O���E&\�V&LzA��Ok��&"O
�JuQ�z�����l8l8"O����Q������ ~ �I!"O��7�+S�<q3��R:8/�6"O��R��(�Z8�C	�U-R�I'"O�'Fw>� ���CrH"OJy��f�\z��RS�_Ȱ8�"O�M�婔�"!8�qЙf"O�h��+e]~�rGo]� #�l�S"O��m��\U�;��̯y0!*"O&��F���$-|��(j�"OJd���x50��*�7��uR�"O��r��@��TR�HF%0�2���"O��s�oo�R���)���9""O����D�� HI* ���yS"O �7$^K.�,P����"��(y"O��� )@�|~���WC.|H�"Ot���V"c_"��oܡ:,ti�"Ox����	/>�*8C����/�4�P"O�����U�9 �`&��#/�Lj"O�uH��(�VPY���>)��U�"O���͖p���R�6�8��D"OH2Fo99�䅻7k�.�jl�7"O�M�#�4�TX�'�X3$5f݋�"Od������9,xp�
-���#"OB$�M�>>�Z	��``dt}�"O~  �V�b��m٣Ҿ��d�c"O�Yǎ+� ���L�GgH�"O���j�)��|RG/S(g�v��s"Oz���9�J����FD��#"OZ�k�:Uy�h��n�9*-���P"O~�@�`�^�x�P��0�ѹ�"O|�!D��M�~i�3�o���XW"Otl�5�A�]��}��ϛ�u���7"O�Mjw��k`XD!ʮug`@�`"Ot�kĹA�d����Jq����"O*`)!�M�f�:P��?��%A1"O�����t��Q9�9����"O�l("c˒~J����U�?��U�$"OF!�g�U3Tc��C��L�`�"O�Q;����~Y���Y��D�"O�0ё��/x�Lu�T T�l�BQkr"O^!�I^>w=�-�V�Qz;\!`U"OH���Q3AV�U�%�U�n0����"O�9�õ�Dq	��א.f�S"O�x��-�U�y G^1�l]��'�.䩵+@�C�dhd-"�ڹ3�'jҝ�@g�w6,�D�ܓ�|ɹ�'�v�3���0�Đ�ΐ�h��R�'�6��Ή�d)l0#��dl ��'��c�.8v��!�=_]�h�'e�Y��K�C���XB
c�.���'��@r
ُ@�-bV�B�S�h��'����󧊿3��Bu�M��A��B�<	@l�%3 ��(�L��b��0�D�@�<)bQ'�$�x����;��E���Yd�<��.�	D��q �����ċ�f�<Y��D�#E  *���ogL�6/Em�<qF瞈�|l����ZO�AF��q�<���{���c@dΝ]4��ûw�<�&K�.�D$;#՘BS�9A�L�<� �	��g�=hvҁ�
�`*�U�R"O�pp�M�6����S��bL�"O$P1�����Ç��3�,BB"O��K��>q�e�Ԁ#%CN��0"O�$�X� ��}��@@k��i�'"ONYP��OR��q!a]7�h]�2"Oz��6 6���+dKS�L�Ll�D"O� b5`�!rmƘ�j[�bU�9��D0��)�'S�X)���]C���4���ȓqO��ѧ@S�-�<��L�@@X��%�tec*�`6�d�[y*Z}��v��5�o��`4��+q�S:b��=�ȓI2�\34�B�c�DI��f�x+�y�ȓHQ�����A򈆄���ȓ,+ �6%H�Pb�[�������ȓ]:T� g�0�L
e�#*��ȓ����hR~F$��]�
����Y�.ay��"{� �B�9,`Ї��G�'�L��fP�a D��i��a(�'n��k�w���Fh�2����O�x$Ў"��)1�P������"Oz�Q,�+w�(]0��V��@!��D#|O��KD��8�ȓ���f�08���]x��k@�4�ڨ����.,PD�*D��@��+�Vj\*/PI-$���$0?�-ٖ(��IǪ^�oX�(*V�c��E{bM���c�
�� i!qKW��y�b$4�e��(�tyP���y®���̐�or� <�J�-��'0�	r�O��ɩLE',80!V��l'���fh֣�yB!�l,� �k�9x�,P�@���y��)��-����h�eJ�
o��<I�,D�	�!�OFq���Ŋk�����%���f��L*�`�3]:iSe���B��H��&6�O��j��)# !	�.B���bhU�$O�L�� ��ؘp ш(��dH#*��G�* �OV�Dz�Oo�Ie&�'�S{�h[�'�?D6�͓��	p���q�=2@A$"�U@d�9SO-�I: �Z��$�!��8�`+àR����@� ���$�_�x��W� �J�n}كl �ഊ��9}��Y��4�0Ǖ�P �����<���Ĝ�O`�q*C1dsbd��� 2�$``"O$e؀���M����0`���Ւx�BLl��(��5�$MP�F��F�p�0`�"O�)p��1:�M	�G�vU2���"O
�ta߆���jd��6�,���"O��a���4�l�� �e��AQ�'3b�=���(OX!8��E�Z�%#���0XF���u�'��c���< ��@�@�!��Y�"	�'7!�dN#"Լ�֠��N��x��	�����D�De�.Z"�O�vmA�-�y��.,O���"ۗwJ^L���@3��=xr"Oze�bf�{(�=0��Ԟ80�*OЅJ�+_5���k���=���	�'�rLY��Y�&���oOe�	�'`QG.S 3{�$��ÖV�F���'8�11�����h��Ğ��ı�'��p@��a�"M)�J�7���I�'J�žp��@�a��'� )�ķiLfu����-�q�'1��5�����q�J� OA����B�)�4��D��"�(~6u2De�#�y�cH�M��D�O�o����b �)�ybaͳ[�U0�kQ 1[d�qL,�Mcu+�0�?	/O��G��t�? d�J*P<  ��Z�=?| "Oh20h]#
l�;&��*#�d��"O�M`�ᐤV�	�R�ޓu��T[�"O$b��J�T��@�Ǉ�@�����hO���3W|С9��Y�Eab�`GF�=5�!�$�`�Y�P��|h�/�=H?!���:��e �F�,��4�g�;�!��-_�$ �č-BL��%��!��5H,t(S���[��Ay�mS+y���⟠Җ�D1ʓ������Z�g.6�!��Z&��ȓ��ɧ.B��jLiV��{�̕Ex��)B��N�V��hB�W0��Ls�+�X�<RB�4_X ���=�( [�N�<Q�n�"&��!��O%2�f�ga�'�?��b哶*��ȶ��6����m�ԇ�	�oSdU���VL��� �P�T6�C�In�z� �>n�ǮN�x�DC�	:@�@XZӇ�*)@� "��oV~��{}Ҙx�Y�4$��ݖ������H�$aj�b�[�C�	�s�3���MqLɣ6�η\����`؟ܸ�eA%=sK[zv"e�3�H>OBџ�D����4e���w��7- �f�h�J	�'�}�m�b3"�F�"�X�O�z-O�ҧH�M��˧uD��3f @�"O��Z��̞P\�@䄓�{3��3��B���I�9��wFط[���vOұ;!�D3<lD@6m��l�P�(O��=E����V}pp��7�0Q3%���y�BǇ!�TU���-?��������y��|2�'�*� q�#�^����U0<|  ���Mh�d�ju�!��h�HH�T�w�!��	=��+���$Ep(Te��֒>Y��<%>c��ْ�2S�U��"�|��s�>D���b@5D��H�+\�H;�,B��<ɏ��&u�V����ٛpv��H̟8�nC�I8�djs.� (k��!ň"AL7-[���?Y��8P4n@�GIѕE��X�5��c�'C�'�r��|�D ,5
���m7 ��yD�b�<�s�
(�t9ⶌ�1�V(zU��_؞`�=��b˶>H*�X@�z�����/�[�<1�i�p�@�x��� (��`a	W�<��!
�HA�9���P�P܂L #�M�<Y�� d��,��-D	5bJ(�"MVJ�	]8� ȅ����.XHFj����9A��#D��͖C�
D��
��o�����!D���h�D��`��A����r�s����0�)��]y4I�d2Vu+��@�N��"��1D���&��C4��#��Y0kkp,���+D�8�7�ؼl�
��2�C&�TH�2�+�OԒO�D�"�����r�Źd~��E���b�'U�����7:p�c�&��x�h(I����	"w��9be�Q�_�T�h�l �v��C�	������
?���Y4�\���O�˓��S����Bӎz���@�ېc:����u�0���7J�D���
[�b���h��t��)�tK��#�Ǝxhj)FzR�' ��j2�\�+�>�2C�\�߲�YCO�x:7��;Jεz��*���:1"OF�r�HϦV1�;�ޛeN�\�O��Y\H<��bˁ�:,,T�B�Id����'���� �GBG�$aP� EGD|r`"O�ܪ�[�VQ��5 D�a��"O�p��n�Q��p���aJF Q �D,���$�	+�`��Z�g�i�c�ƛ&&!�� Ԙ���C�찹�&W��]���	ix���2�E�7hy��(@3i���B;D�|�e�շ%��M����qM��Z�3D��Ӄ�V�2!F�Z��R0����0D�Hs$gԑqzLj ��Y\�Ha�.D�h��-��U4h4fL7	������/D��J�ܘ$b���J�rT�R�a;D�pi���p��yꁇ��./\(���5D�8مl� t�@��&��i����&D��`܍f�]k�b�8O���SE(D��3s��J���f��rz9{Џ:D��v�Xot��&� (�PpRa&D��AT�r�J��&N��ZMyB@9D�l
QC�r_D��p�ͨ�V5���5D��D�*�Z�����8�$݉�#0D�h	�K�!|bحh#��.�$Aj�I8D�Dɂ���8t�U��&=HB�/5D�xc�e�v�Z�Чf�$)���+4�4D�H�R��h����%&�R21D��0e*-+n�K���/�R+�O+D��)��P�~eʧ���1֐����'D���uP�:�t�w�	/FŲ�s�e*D���aI��a��(0%�L�ؔ�=D��£@�8�&d�5eF~�Y��n<D�\sWNQ�Qæ���C�:XZu�R�;D�#��ȼg����ݞJ�\b�o:D�H�ˎ�S���@GK�\f�聃�"D���f�4sp���[�Zkʐ�%�?D�|!��#%v6����Y�<��H���>D�4�GD�L�����
�Բ��8D��DB�v�BM���6�����;D��Ȣ�ճ7|��DÚ'/�*�3$ ;D�X�2�QG�q[0ᗈmW��g7D��	'nT7��8(�J֢v��� ��3D�)��)��$6`�6��@���<D���QFG�ZN� ���F�U�7D���ӥ�@�����MX>�8�0�"9D�����!�r�h��
4  �"�+D��ʧb��U#�eK���[..D�L�%��&��A
�IK�erB'�O,=AQ���f�@$`�X�&L�u�-��:�"O��E��?b�#"G��h�s0"O�	rPF��	��Pb�_�i�z�"Ox��F���DJ�@K>t�^b"O�1a�ѥW�j0C��J��J�"O� v���,=�n۹E���Y#"O���U��AbЬ�͆���]�!"O�����@13,^i����j�"O��#IV�� $��x���2�"O��1i	-%��P`������"O�Z�	םkA���Dھ.�0��"O� xG��F*� BdO�k���9E"O�=!g��-+�\H�t$ �o��c"Oꌠ���F ����h�^� B"O�e�b��}c�P���"�\X�"O��vOs� � R@�<��uj�"O�p�r N�(�e�&$þ AʝkS"O�	�c��e�F�Q�ؕDMnśD"O��#IS�;�( t�ԩ
q�0"O�U�Gʚ;�Ĳ���	�@��R"O�Y��I� f�Hj�b������"O����d	=���0E���%-���|cz���%+���,���C�V�O��U��8	hB�əe�\�ƪ8��al��vR,���̪��0H��A��S�? &����@�4ja,ъP��� �'�,�U��%B��L���G?mY �/�
I��xJ|����4��ZR�H�b��x��7
�<Y�ǀ������ �1��$�Ɂ�\�zEy��5nxz�7E�?�!�D����Η�T���H���Q9��O�U�l�E�E�<�)��0�6���|o�H�ěv����`>D�(F'�����!��U�P���߁cu�e	AI��|6�`I}���3�ur��sY9L����@L6zS ����b�X(��4O�h�W�j���I�/Z)8��RU�ǵrm�xТ�
|ܶ�� ݮ�p?� �Q;+&�|/i�܄s'�acB��{��'�͸�M̌�	�
�۲���d�!�<j7٥Dd�8�iC'g�v;����y�C
>mV!{�`E=f���_7r>���S&T1  D�#���+K��y#���5y�^�c�NE�珻����	%�~�Y�mлn��ڣ�.�	�A�^��q�)P�U|z��#�n�2 .����F�+H)@��(O���a�ߒT��I	ՉD�v��fh#?�aP�̇-oǪi��S�4�"	�%�_�C�z��V�:����A�t��֌��-M6�Z�M�X��bt�F�k�X����A���� H��mk�aψ6���?�:=�M�%	���\Iɒ�R�dx:!,/���{aU��8�zEJG&1��r�ٽHaJ��ӭV�nh*џ���I�n9A閌Yی� Bg�#3���H�K�nnA`���0|�Ǝ�.\���
W8��y�*	m���(�"+���PE�IR���̧\��XQ3��9�I�l���"���Q3�؀��Z5*���ŗ�.����e�Ȓс̯+�Zl.�+�1���a��=z����F�K�?����'�Ħ+���Hn�m6�l���>x5Dp��+�U����V����/_�<��+rr�@`��dJJXK�aU7���Y0I�$4
��p�$5��$�?�� pv#��ހ}p�� uw\�c�̓c?���BƐ'�l�d��A{�����,A(`Q�l
C������O��2�b����D�_tz�u7H��B4\���3EPn�am���p1���7*;����E��l�.�d�#æf�����y��E�<�@HD'�0_O�	AT�F��X6�G���sF��;'���@��|�#Av�r!W��<-束%������:tnF�;����*���	+�r��ջe�<)��{>�ʠh�8qb\�CL�*���Bx������7���H�7M���\݊Q�ؚ|�a(�I�?>�(O��������"@��V�=��*!���<]ܙ�� G�up��ci!�$ǐp~���)��h7��r� �C,Ru6��#��7R�"ػr��z��ݻf�(8�nYEH}yb�ڴ �������� b���!�&ryvT�QhB4�<��fh��DyGƷ�0c�i���������HJ�j\;��cbK�C���yg�@w�
isBď�&�,��l^�r��Ig(��?E��';��c3��`J��2�K��ʔa�ãI?2[*}`�dX�P��H#a�%>:��ScB��Z%��6��A�w�4@%f�>Qc�83�� Kfl��'9�*#Ę�M hrU̓N* (҃Bj��2����y��(��4�؜Y�c�f��G(�g8x���̛6��Q��`���6f4[��^ C4���3(4p�s!�³#��#� ��'��(�c�:!z��CF?�<k����&<�%�SeߚpePk��̷M.�Y�%Z�O\�!fE1�����K��`H:���D���R<�3�>sɲlkSυ�+
`D�9�X�S'lJ43�J`�A��D���<p̴h���s�B-��g��0qJr�HF.�ϟ��B.؜p���>E���+<���QΔ, �u����-*�r#ɹ�T�" �Y1�lx �O=���.���Y�ec��~��ϭ7�npQEF�t}��2a�A-��ɮ#��)u����%��^D���X�k�F��2�&���b�S��I�v���*��}@lޚ&�	p	Y��Oh�r�ǹ(��ہk�Wn���D+3hma1C��O4�q���Z�,�Z��V�?`p�DI̟zH�!���/a{����V%��ܑ�d�B���j�U��I������0��/uINU)�ۓAz�0�q�[;t�n��+�}c(O;rAW ̼�Q ]�9cL�i��[�Va�C"��J�<Q�/0z�� �۝}c���rS�,<����!���'�Ȋ-y��Q��C�y�<���ڟyj����gI��?qF�V
D���r���|F�H�˂Z���c��<�Z��a�1~�B��'�K�~utE�@A��l��öh�{�L��gVFP��N�h����*Qў��K����T� kA:�� �C(�Ɏ;�� ��/��裁m�����c��<\�0�R�J�<�V���[�Q��!��
5r񤹚�JD)*�������s&AUn纝���U�����	�`L��[8[�z+��ظ�����h묵�+F2U��;VzР�O�*�@�b�WK�مȓ�h$�O�iv�`�N�u��|�@J�;�e��Ǎ���HW
��b8��/Єo`� q-��q��H鐺i�\����N�j�2���<TH82���j�����V��5<P@ 2�~�dK�U���Q�](R@#���v�����~Aq�Áo��	1��pϮ�S���f�&,���&$���	4=�&��q�K>aWRH���ߞ?�vL�3H�F��FE*���n��8�2��$��e_Np�2�=�bd��HS7`ʐ����&�L��g�<&.@kvlX	���x���FK"����ށ�!f��_}� 9䎎8]�L��`�΁q��=�LE����ŎL�8P�I�#]~��(�u����AH�"iC�+O-th�w���(`Rx�1,7]XN�OPp�q���^_@MȤ�7y��ѣB���\i�Ņ��O/p�^�*�i��W��e('ϒ�UcF�R�'�Xa��u��y�ɐ�b�"�Y�N�T��iw���}oZ�J��A�rK�D��i�5��
t���*�)��d	$)�4^�-y@�FI��M�B�F��}�e@�	rذ�Z)�F���# �|*�$k�W8]Y$���E;5x��"�e	h��EÊ*�V�Gy�.'+�0�F�_�X��B��:3�b�M!�v��5j��z5	'��(��#%d�
��P���xp�I
0R�xaA��	>ށ��⚈Wo�	�V�N6�Ո��		:ҡ�G��Rc�9���O��� v�������P�ORF��t�D,����$z�IJR�>E�Oڰ Q�NSr��7I"t{�`b��
sv��s�IK�3���$����!�H<ɇ�PNJ	+�a�y�&]�����y��$�T1`��g�Z��8ajܴI}���S�ρ��YXQ�i$N��&i�|r`�a �R8"إ���9k����g�� .��=լ�p�e]�P)BU���w�����-ۍ0P�:��!RO�l3_�����ǚ-� 8@*�(&o��t/i�f`E]�pњ�X��ͅ4#�%	U#]�mY�-� ��D`ےQ7�%D}�E�L��i�GG	�Β�k�6.�H���&{q�0J�̩<�¥&r���i"H�3$�6�[�yT�l�4�ʜ�.���K3�p�Ƒ
/�ay�K^�e0t�&��R�q����� �:4���cA���XK���A΃�G��͈�N�2�������;�"�Jĭ��[��
^D����.C�A�xq�7��~�����(K�p�nOV9Ss�QR���Z��-�R�C��3xM!�Ο,B����/;��q�f,�G����� M��F��M���(O��pMNK���!��6m�j��<� g��h��&(�|��"�X�!f� ���L���)�L��p��e��8�
$-�l��RM�8	X�!Q*�1r���D�(���PQ��)CwJ�D^lٱ�	^x�,de��mS
�~.0 q��CRP����7r� �هC�`q6q(�O�Y[j��?��BQZ���D%Hb����C���m;�&�k��D�����W��5+Sc$-$�a 38CE�"�tA��G"�
�.�
2�F�P2�F��?�!OX 0許sK�� �z,E�F���9i���-M:h�'�ֆK|�!�$c"�%?�x�Q�ȡ}߀E)��>h�0P��l�'�8�M��J,�'�ϏXr�Q[.hJTm	�y21':D����.�p��ܟ�qO|]y+ҺmW����OP�4��D�W�v�.����� �IS�̄!�~Y�;H�M���þB~��#a�<]R��*Ǟ�O���i��4|ST���.A�fx�I�4��d?�M�'e��	�0��I�c��}�E,��28��)e�*'���b�L���)�B��ðl�6�V	��ؘ:��UKu6o��j@a�LF5
��S���,h��,�p=��"�63	^�����l���M]�OTDX�s��"w��aV�
����4�At*)��ď76�!���~�����#-N�ҺoD�Y(tE��q�@��g��P��}�'Q�.��&DS�G��$���>H3R�P���{*]D�L�04�t�U�'���@�B���0Ó�J0P�H�iH�x �Dݽ`dTq�� g ,�Ѓ8���h�n���	H?�����΅`�����p�jᧄ#:�^min=g���kǭvZ��h���3殜�r�~�*���;K�Ls0�ɯ/�Ā�.K�3u,���ʀ5Ē��2O����X��úI� DS`,�-+�ШCq�1p"��T���91�Y��$B�`K��
�ѓ��.�x��D�4Gcn�xʏ6^�c�abNx+��Ѫ� ��8Gn�(�@D�Dd~�0�Mˌ7^�$A��g�.	o�6�qq��h9�]�t ��ha|�%>����b�T k�C��t � �r^���E0v>7m�",nҐ��m,�Pf�F X��Bע��i���O Lqe^7~IZ�
0�U�"%��	$%=L Є��?k���� ��Vm�DH'��!ƁӇih�)aLV�Q�(=X�.��d$I�F���|�K/ C�V�q!D�'�J̐�/�}u⨋� ק���+`̄�Z�e����9Nf]����8�^��Oڅ~}�����z���S���_��A�i�Dp@5��
HE��8c�؆T��MX$�'�X�
x��䣓#��2�2@@ѩ@�v��ā��?>Z�3���hbߴ9���Ǉk�M� 2��k�i ����lN967�i'�'q̥�ả�W�ށ��X�q��#\�
l�v�C�I�,�ŇݑTQ8�����k� ��$A]t�5����_�x����O҆�6v�|�d�K� Bp��@�Y%�O�9��L�h�l�j`���H��z��N����.� f�j�)v��p�t�c J�@�>16M��dM�AKLF�?�TK�+`��lh�	b"�x��O�?�����玆WIJ�`�"
�<�`Ż��ݾ*t�H(�䔈`'�X�3�V=9����(!��ՙ�!^�L�{&	G�2�sg��*��ڤ�'~�0 ��� j��D�$$��S&�Ac�
�N!�f��OB��#%�3t� X ��"m��p��dʹW.�y�w�d��*��f�V|�t�P�(`
�Cof<���H�8�-�2f�q�%۶c�7*�L�hŁ)l�!Jg�Ѳm9�H��+ċu�B4�R�� r��#�5.�F�P�Oƭ#B�!5L�I��愝���.q�qO����e�waJ|�&ɳJ�ʼ�Ө�
Pd��Ƅ�,�BU9w��)X����o��jn`��B*U�w�.���̌4�-��&6�/�V	Y�!�D���	�#�r�ɳ	W�!��
=pl�lzbh��9�d)r��X�%�H�3�F�& �f��c���$ʘ�Sf�����}���Ĭ6�v���׼d�Q��������B�J�,ZyR��l���k5�A��s�+�y�`����8P0�0���V��8J�獗i�Ґ[e���
�� Cu�!�y�nȯ��͚@N��.VB�g!�I��a���q딕@�N(ҧv@t��CC�;��!��B�QyM�g�ڿ<9B=(��� �ig��|ܠ���#U6��yq
Tse��-����g�	i�!%�X�=�X�k!�W�|�����'�����\	]���M4���r����
�΅�_���"b
��Y����K	����qED��𠕯	/5,��H/�RN ��*����'2�"����~�"H�7Vx��-Y2Z^L�'h�*$�Ay#%�%}ь��d>�*�HQ3_l�'-�VF`駈]>k̩x��+"�$ꗽ.�����܋ٴL�=i3NE�hS�tq! �'U��y�ׇ߇7��s@��">�+�	�%~��1��P����π3u�ڗ�����_�Tѭ�e� ��\��0���^�D����"U�\ 1� �aD�\��O���	��r9{B��X�~Uh��ѫj+��h ��?��K��|��B���ii����m�p�W��+T�N���&A�G ��f�x�����Uja ���$Ëe�d��47��&*V�:�Z��ɗ�,w���A��b�f��*�o�`���ǈ]%+�U�BD����>L���`E��#�2	��X!�~�K���6��$2�O�z��mI���8`2<<*
 '�>��y"JJ�$�*#����M欙���1	n��'�ͲV�`�W�����	s Wz��$c)@�O����!Iۺ����!3�Fq Y�WXJ�s���	����Q 7��1!%�վu^�c�49ue�<qT�QS1@^+K[X��YW�4�"C"�p�Hel��AI�(PI�!�ݱ4��
'�, qD<��Ч��Ke`� ZB�� x4pvcì_�%�Gn��6�eʖ^��� ��>vrh%�q-�7v8,�1AW�	��k7������>��<!q�_�c��x׍��n#L�ѳ+�I�r�`�r�\���D>��09A�ߩb��H�mT�m&D��ûie�������� '�
'N�P�&O(Ҏ��) (~�(�pŉ g��U�|"�E�F���e˵��t�M�.�Zs�*VL�l�`��$��rA �#1mX�:e��4��l�=9��C��2���k{@@ǥV�X�M�,Q�p(��gD�wTA�ˀ����jGkzBhEхT� Xᭀ/T�`���&�A�~M�5�P	��#N�9KdL%9T�7�IRJ��eɖ�FԂF�⨃�nS#)���C`�WԾ��G	�/jϘ� ��>�`ae��8�t�l�*�ם8QLq�B.����$$�R=��o��.X�x�DD�/�v�'\����H�g]X钴Dҫc��ApaE
k���h.�$�!�'Z|xT�C-�Aiu� y�Y����B7����W4&#}��wZ�h�4
�j���P���R�H�o�D�`�d�T���zu7�� �U0V��eF�{��,M3�ă7�ܥ^z��BF��v�8��d�=z��I��Gn>#>����Dj���"���
�0�2��&
���@ߤL`����:��y�H¯F
y���H6bH �-ǜWx\�1��P(Y��LxPCFs�p���`а�\&�� P��Վ�������%b[�������5B�3@��D-�)c��t���Az�V�cv�Ǿ��OL+���	���?��%U�w�r���{m�u���ޣ�yB+9���� �K�C$��MY!��/69������)�'\N�ѷ-[#l��5j�QBć�798PK�O�+TB4
�)Ӭ$���=ф)֒Y����$#B��	�	N(><����8�!�
I|��2�=ut%�q�=z�!�ď�>��a��M�#���;��֐�!�Һj��թd��Y�*��W�A�3�!�$H�'/�P��NԊ/��VT-R����ȓr��e�A�D�D�V�� n�21�츆�oN��R���NND�:�G�2ߒ��ȓ$�(5��F��U�,Hwg֧| ��ȓX�P5��b]<hMP�S�8SD݄�=�����U�U�r�ӵ��-�����Ԡ�>@u e3�Я "쁄ȓ/%0�h#�F�!��Ĳri�*8���I��"d,B%K���FǕ�P�*p�ȓ!fn�0��0�4�0�W����H�|��cX.'�<�H&�_������>US��K�\����R�K����H�=�$l�)���`F�M�U3��ȓ0L�'�>A���W�D�T�2��ȓAF�QCi[�v(������ņ�[4p8Q�ڈH�xh� !Q.�:��ȓ�*T8�͌�H�4X�!� b-��5o�8ӫ�X�]�U�51&H��	�|���=C�L�pGΔ	bڠ�ȓs��8��'��`�Z"�DI�]�ȓ��}C�ܼ| N`����E���ȓnF �J��,9�LP QGR�p�����v�J��ʄ�y����p� ��TW���5�b��2v�/K�R�@�"O�lc�[�H�MҥOE�J�̼�`"O�)�d��$I�ҙ�a�٭8`z�U"O���fEC�$E:A-E:>�4!�w"O��vG�rD���J�*R���f"OZ1 G+ZaJ�K��C(?X�+7"O�%�A�,��X+Gg"7U��b1"O�Y�V�.;@^ ��f�02�Jdɤ"OV���lC]e��1��X�u�,�q"O���bCD?_$�p�WJ��C��(��"Ox��fʞ�.;b)�V�Y!*���"O�m�$�ƖK�6XZ1H�"���!�"O�� ��J!A�&�qŇA-=�� ��"OŠ�щs�h���e?[�b��"O�)hSl;K�9a�a�[�<��G"O4��R�"ǼL�Bϗ�>��"O@�!AfB�d�n���,k�jl{7"O����JC6J�^�ǁ�9�E�""O� P��nGP'|��2��_�6�D"O���#'T�%�� ��dXs�O=�Bm	�!���O�>(E�
$C�����Ě7;�(��3D�xfK�h�����x����<Y2�Wp�U��0<i������e^�8��I�ƕpX����ͪc(����,z0p,k��2
Lb��Ų�'M@�!���H[��`g&�B�ȍ�	]IJ��m[�K]��@G!��_�-�$��H� � ��C�4S�!�䊕c�� ��	������UA�'��P!�k�!<�y	`
]�Z�9�)�矨KX����ӂ�n���q*z|!��2�V�҅�P�h�8�K�@��1)J�-_mUY�����`0�<���b�@�-%�m�C�@Vci)�e1��2�B���+3����hՉ �����Ȁ�.�m�f/�/���2Ŏ(+��
��v�Xhw��8�ddb�bZ}�V��ɅwŌ���.�&(�����]�, � N�w9���@Et�da�#=C @t���g�~�;T���!�]�d�ޭ���L�Р��`�>h��Yaf�\�I�d��(��rTj�4���S�.�8j�ʒP���	�l���X��@�zz֡:#�XM�㞘�rl	�f����{�i�{�҉`��5b�(�٧�Q��������M�f�S�;�`�cBuɺd����"<	S��j�����\�J�Q�'A$F�����Z�N+ȓO���c Z�J#��Q �$}PRt-�=8�հ$�F�Sw��iT&Ɨn(BMx$��.C�~D%��[��� [�-�V��H?y���w.|h������AL�'	z0 Qٸ
g�����t2�˄�ފ����B|��8��y��F2��)a�N�U|t5�t�M��~�		s����k��!l���ӌi�"�I�I��A�K2dȈf`�+0E�d�t�@�9Nܙt#f>�:��I4M�4��aH6fĈv��-2Lh�a��E05��>GJ�z���$�1h	>, ~�-xn-��?I��ˁ~���e h.}k��ͺOO��e���"N��F�g�ڠۤd�![�&tIpb�m"}c���:LH��%N�qf�51<��ӂB�d���P��z(8dBc�.-\	�)O���	6������ow>T"G�����(/7Wݲ�r����6i`��ɥA<`c�m�����̓�'ʘ���6T٠�"QmТ�&qH�<O��7p��A@6;��aKN�&K8��30' �NP��虴`�d��4x�@��� mu�Ο�nM�IF���W�N�`������PnZ� 5�Œ	�.���'���$��\�65���V�ND�; @�kmXM�\�z�� �	��7ӎрt
�� Mbh�p]�|z#͘I�D��D�� �%C�� 92��!�R�ȿ����g�R��	oZ�GW.���?V+���JU;dl�cTU������(P抅���n �Y�՝/�@Dj���5J���ٶ`�X�5K���& �`H��ҩD%�`H����h h�s�E�V|�����ąu�6�E��9�J�P��_jy�CT�Q_�Xs�#Ԝ{�n�*a��'޺y7R@���Z��y)��M�Uq乫��&( >I�(��Q}�@hu�;���x$r��T�?�]��mÇĘ!L��Q��^47"^��A!7xA�1�D�����A�)��<�â	0뀴�Co�;A�-[��M"=+� !�	8;�"�+$��3$�0��'芨����G����1dmΨ��C7O���B�a�\?yCƍ�o�Y��ǖP�b�P��'�	\�<��E��o�����iR0!��oZ�9A�@m�1�*ejf��2|�tؓ�J g�Q�O6X���Iɤ9��A�5���Y�,~&㔣޼��Éy�Þ=�
����#-��Q�B'�2K5�����dz�b^�4A�GB�z�<�0���C(���o3��ŃE�Z,�+ߧ)�J�>��R���Z幱�1R�Ҽ�A�?,�"#��Tw4s�N�(~Kʕt��hdj��9��2��y��ѻЮ�$��|ƒ�b�@N��?!!�jKt��G9}���D&Y, q��W�k^�b��T<G�PQ�!�#�`��^�j��U>C�J��&�t��v��FP�+��Of�0��
_	�Sf�*\��YRw�>��LT�c�֝V���$�U�K�A��n��d�&��@ HK����<�"f,ӏ�4��K�|�u�C���j~�bC�� �p:	ށdv�㞘�4o 38ˊAhs#י�d, V��M�8�c,��324]�c ӊc����P밬�p-R;:�(�ؔ�˅�J
xJ����\)Ҏ��M��Xค�g���e֡j�	/�M�7k�
�Bq�M9R"���wp�5�����] �E"b���'O��H6�N�Yu��W�fԩ)5��c��̉e'�d"����UO��`F��\����&
l��A��'VqY�H�p;�)�AΝ�)�	�@ð���݀��ʠ]5�eq�� ��B��K)-�����Z�L(��.�,A����r逝Y<�I��D��`)~M�GJv�L�+�K�8�1OH���=�ެS6�5r��)7�?��x�s)�:f$��c�N^Vq����_$a���2f�>3���IU'
IX������Rs٨c��A��hQ%썎z���C�Ǒ9��YD(Q�����ɟ<T|��Ӏ�E��lAumޥ" �'.��x#���d��H %+&D�""#��w��Yed

i�¸B'�@#%<X�wlћU@�����+u^*rÔ�r��1�$�j�̘���M� �4?�ii@��]� 9ksЅ�jA����D�х�36Q�0[?1�U�,@�����Z��р���0xPY���v�0�2b��<=@G�':a�q9���$[R��A`��HOB�{ƨڠ3Dfxc��3�!��A9g��	2cF�7��=�0!� _V�#f(Z�0@p\##�0�5�%E�c��d �.��h	LQ��q��!�b
�v�V��Ơ�u�'��ya�F�9^��ka%�sㆀ�0��Vڴ�%ѰZ�x���`$Q��Y %�ů�_��4D.��)#K�b��=�p�ܑ1�TX �^.5@�ZAG�]��y9Ę|RE_��WŢ"���g��^�a�ץj[=B!8,D��U�]���T�a�P&!p���d�^�����/O��Uj2�ƛ,F��J�=��@�Q�"b��r�� ��S��Pm��x�#VQ�0�0*]?e�&�%<8r�!�oB���cрДl��l�S�V�S�<� Jܽ8���-t���3bB�6�dX��n^�'�=!"�t�@N�q	4�Ȇ�5�l
�XEi�l��Tb "�~1��(�S��i����"I*�5H�V���x�	ڴh�1����Ob	�0hA�T�&��ND1H���J� o�^mi7�R�2�N�t(=�I���
 `�i�FA	�Ɠ�4℁k���[&��u̘���T(Q�����%�/XÀ)SQm�� ̎�U8�E�X���th�Y�Ĭ�0%h��~�^�CG+Z�0}����x��5i�I$�����o	r�|i��G��L!J��1��СC�<X�L�C�,_'�m��4;j��gkX)<�t���kĹIv��!��{����>X�D�I7� ��c*38TA�!��1�eè<<���Xs�@1��`#Z2���
��64|	���8��.�"pt�x&��� 
�2�Q�W+�;���Ч��J��1#��>��YҘ���KF����͕-���YP�ɘn�t,��_��bֆ �#i��⑤G?:f���R�����ݱ�`H��&�Kd,�r�ӧİ<��	͏9��tpUJ��I�Ε[f \"0�0DP̒<=w<��!nͼy�)��BB�8�3��ȋ��#1�*|(��'q6����?~�B�))j�P�BزF}�X��D�d��'��d���Z����s����@L,��.�������Q(`@t�zx���L�sd��V@]�MS��,w����	�x���PH_���J'ϙX̓�T#��'2����r�F=  K77�fIB�ʂ$:<�rǪ� �D���%7�� XB��q�H!��~)V��ਚ
R�F4��+°7�h��Ǣ�	���x�NE�n�$��I/��Ę� �%3
6Y��f�$I���Ɍ	6���$�J3�����Yȇ�F� ��,�M������`��\�v3��Ueσ/�ɐ�.AN��Ժ�gaA��qj ��12�Դ��ݱy�m� �ŷO�T$;�N�*�	�G���^@�4�а�`�O0a���ڥR"��i�.QPf]��_��Q�0�I�} qO*|��D�?Ld�Ғ�Ì�f���8NV�`d��*�4s���Y�����%,RL8��@j���'�L!Ѡ�*�����<D,qO�d�R �}SdI�&l>=he�6/ �p���6F��h���S�Wu�`�� Yf<8��Q�"�l�����ݼc�G?�A�z�Y��Y�e����C�4�9dʇU�MJ��/O����LP-o200���B��_�|��a�=�@��{�NYx�����C��0O^(�h��� �3]�8� ��U�M7��:��
�8��a������0��˞������rH�e�a��S���!�iT�8�v�H�k3<p6ʑ? ��G��n����wzL�m_�R�\��fb.XƖɱ	�XĒũ�灅--&��ǨS�U�Ɛ�CʰW�\Y!�Ӊy�*
��9?7�Kաɔ%4���� Q�ʄ�cJ0V�Da�'"^���"��4d���>~���{��$^���E{��O��W�=hl�1���9e \[P@�h\���1d>�cfA�D�@�ƴs��9&ႁ:b|G|�"�`�n��c+��fV�� ͖�!)�iN�:��TQ!T��vJ�]a�j��+͖cB��pm�##.�EXV*R�z�TlYlM2)�4�8��)�6�7�ŗ4��}�ô'b�0ȡe��4�� j�# `+��K�_�m��mS���Tab5$j�����(ɋ�*�7�yg�ۋs�Y�$̎�Zd���OQ�0>�kL|��(`d�D�~$t�v��ڥ� �kXrt���h$���A���c�ʍ)�Z����*\�c�a��>ޤȀB�'^��C��ęH9��`�N:���Ey(
(V��5��M3��R��O�������[�WA<Y��.��T/ ��hVL�I_쑣!l�	&�1J���N$����y�'���%�	{8LX��F@��~��Y���WcŦod���M�w�ؐumшx0Xt�&恘	�j4i.H\��e���!WNU�e#��ܰ��C(�4�^�	R�'V!q�C�-]B�lSU��?PMȢ�Б7&���D��P���!U-^ ش\�����J@z ��05��X`R�V<(� �b&i�l��c�'y�tSLV�%s6AT�(dv|Uc�&x�^)3�M� �BVg��uQ�e�ɔ�Ԋp��*a}fa���{�X=0�RGA�hT$H��� �������O^}Ѣ�π!ڰd�g�'H��ˁ�T�+
�8`bM\�O�ꅐ��BELt!*��4I����M:�DD֣v�pm�4@ݎI���zƯ�m�|T�6�ȝ1,T���@�f� �v��'lٞ�Y�B�:i��:�O�o�rt�7'@�dP����(Z^؈�\�haj`yv%�?����	*V��Isf
�` ��+2� ���i�c�K�m>��rIR�|�¤�6��X��c�$�L�5���Y�U~�@�� �$Gw���3�'�����	~n� �*z�~����A�Opt<2�`�d��G��	���A	,A�^�ˇ��Y��CQ���dr��(*�%��Ÿ_b�\'� �I$F(�� �&/�@9�@gȷq9���$Ӻ\�e����!İ�&��\�����9x^Z�Z�A��l?6���M �.*�G}��.:��5���+�c���C!��
�?��q!��ua���đ>���q��*� [��	N�
_�qx��,��A`��@�q1�!�L���BiJ�"�,O�y�ԁZVmʔ�&Z�-����YM��&�+*c���2IH��U�d�Rk���F�/��,Kq>�j�!a�W�ƜQ�Ɣ��ͪ�S��
C�APmy������-9!�}�͝C����h^� ��[̄�gs��9KJ!x��C���`�F\B��E��8�Gȟ��
�f�O���O�n���q��gr�,3�L������r��%��f�+�����^��@��^�?a���w�΋R�z�al\2a��
�ɖ8倠`�놞U���k�^���K�pEZ��E�j��|��#�̏OW��ʂL�nׄ���')�Ԩ�e�./M���M�{^@�!2��ٚ�MjЎՠ�'$%����E>oJPq��m=����ߧ6P�;�D�u~➘PS�@>5>\��/��4�8���	5ߌ� � �8N:,���O�Y5̚�I�5b9�#!\������@�x֜VZ X��0�?=<l���"+�ti��̾�qq�͔�qb|�KE*�>�-K�j���{3��(VHq߄ݲ,�&�Y������0I\HBb�C���!%�I�^��*�D@�%'�p T���SӐh�%O�(sLx�"�G���q�M$X����`�ఒ��­ F����i���@W��)=�&�Pd��/���k��r���� !	�D)��4Y�v���生�� B�ǥ�	+�h����W���K|_v���!K� \�1�Kأ=�V �GH̓<�\<�E"P����F�$_�
�dԷr�^r���+;m�A�U ^�gEXA[�� U����s�Z&]��P����Ԥ9�
Q�C�D'8��`CWwo�M��<,D`���$�>*TD�C��3�`�YǦ��<�U�7J�<�%��&Œ��:�0�c��J2L��`S�
{Ҹ���?R��!aD��>�Ҡ:�:�K�h�ݒux����%I:�j�F��%�8qRIձ?���`�l�*�	�A�!�V-#`��~B�Գ:K�uO81�W��]�0XT����\gD� z?L�`E��F��ّ0��tL0%�'cX�<p$�i�L��֎[[�M`�"��Fd^!�,��o�����A$LDT�D��?	�VȲ�M�A���*��QEb�'�/l�ąQ�se�0� ~��͐rfA�EV��GQ�Fh�=��Hʆ!:hA�@M J쑭�`����FP�X� xS��za��Y�j�c5��I6�x,�7fg����F	U�LȒMV8x�
��$�ܙK���;�]�)�v��7-����'��A+��qb&��t�`�U/_�4=��y��uL���EN�;��YS��v��@�˨[������u���&&�-�rʖy���D'e�09pF��0`|`��U$["��I/`�����ȶEY�����R$���B���-���'8#�$�e�d�p���!@�x���#Xa�q��3��	*4�W��H�V�	'��)��E�?OR1q���xڴ��;p��(#���yӱ����q��
�"S��Ph Ӎ�9rȓ-a/0��q�A:�Ȁ�L!�6�3�(�S��J�}�p�I��DБ��{?A�o�h��h�&�"��'����-L�,�3�*wZ����$k-N��q���2�D<a�%<lO�=I�	$f �;5�*|<QSd�`Xe��;Q���jH>��;P���b����EW�O� 8�0���mK�8���4F��ڼ9�#`��fF�V��`	[4��r҉L�;��8��&o*���ø7/⠒j�0��і'�ڴ��*�(|2��OQ>��p�^dW(,��ĨC��}Q�B2D�+�M� 	,h҆�l|Yp�1�ɀ6�(���'�!��8l	�qҠd��^���
�'�����O p���0�^U����'(*���E��K�-��LA8O����'�xt�c�׏ (���Ǒl�z �
�'Ja1��8>k.]ؖ���ۢ�X
�'ivQxc-��̛`FV�n0�	�'��Jr��i¨˹LZ�L7�yR�^a���;���|Ұ�Y��yRh��^�r�6+
\7t�!�-в�y�I��B�b�@�Q/�)�@EF��y�*��+�)��M0E]��)�e���y2�
�O�T��u��0���l¶�y���6k`���0:����y"ͅ�L���d�P�-�j�����ȓ��m���Ʌ肤i�D°:_���:���!'T�&4h)�N*)z�8��s�� �ǜ��#���WH�����){����}B�����'p��`�ȓq�X��C��<��C�ov���s�����F�71#��s�Iğ�4���o�N� �e+p��#���{����=\�	���ԜL�]�Ð~K@�ȓ#{6�ʑ�M�:>@�C�g�����0H�<��	� (h����덄zN�u�ȓk�H�a'd�<f��N�!�>���	P�a۵��8��m�Hw�NY�׍�������`��ĵ �O��@��#���'P�����Ab8F���[�`{ �P��ʦ��h�C�x#�O����6��o�8�P1��;x�n��LI�����T�+�r��<�a�4�sը�z�GD1bC��A�X�xt9G�
+7�'�a����`����3�I�Y�V���_� ���v�>1�4�O�O�j�	w%�7|�4Y���c����J<�0�?�S�'j�j���K�J�R�wl*{�'c�PFy��iHj�*H���l&L�3CK�k.�VE��ȟ,ȡp�O)I�2��.�L��x���
�����3}��!� �I�`��˒[����}�p��%�D0���<�(��9Za��.Њ
�Z���٪�Ƅ�|� ���k�X�P��-:lqO��V�[f�+���vE�=+I��un�=`Ĺ� ���oV��S�O4�� �(�P8����M��0EQS�I�B�0Y	���d���s��i%��ٷ��(�>�`�#Iy�eX��p��m��,t ��/��O�'%ɢ5,MxP�m ���Y�}" �`~a���+� [��R�5����&��S�1��6OR�Z�.2�g�? �	��FS7w>BT�T�u�*��O���'m�O�Su�8]��ie�
3�$��(�/�����OV��M<E�D�D��xV.٢/W�TH��B7�y��A�$nha�4�S1M����b��$w���D7^2:O�<�4�zc�b>M�"#A�u�|1���!/��"R�5?id+d��p�y��)�:0���a���6r#ʹs�mT�7���Mޟh+'��S.O2�I�h1#0�L�ƙ�B$V�����˓�y
çzĬ���C��F�C1B2DC��W�O?� ��$��?]�d͟��)�?�DǮi����� �x��1{��0�!�D�3e>z�YЯѧx���I�/M�!�$�!p��!,������!�ɮ��0����I�n!�(�i!򄎫A
��9'�T������$!��إpM��"�/ ��B�"|!�F3>\^�i���#F�0yTC\,�!�$س"<�+�Kܕ̦xR�L	�0�!�$��r9R,x��ܪ&� �b�m�8q�!��zfr�b�G�<A��x0lV�!�dZJ,���.���%ք/!�dW�eQ��+��e ������Z�!��FF�vC�;[��Ac�3mx!�D������2�"S�ӵ�D�-�!�D�-��Ԓ-@2j����K�mQ!�d̏+�Δ���D�o�Fia�n�-OO!�ޮp�ȉ�̉=��d� MK�Q!�$ �	S���f!!�F�Wf�Qz!�D	�k5�S�Ԃi~@i�U�ͫq!�$H7!a�<�AŞ�L�Q�nU<xc!��9�\*@���qP���A�!�ĉ%,��d$M�	���6<�!�O�H6��A�/J�L6C�σ=~h!�d��O�bL��!�n�K�v��t��'w�5�AL�zxt�'gB���	�'��r�ƦQ3V�Ń;k��)��'�q�pJ�}/y�3d��l�$��'($����	�i|>)���ٶMd�U��'�lP���b$�(n�BF���'�1� �+TѸ�� h��|���'��H�s�C�df*�@��^��t��
�'C��� �H�EJrG'U� n�)�
�'N|RF(��~���F���'�ֱ�'��,�Q
)}H�V�Uht���
�'Rt���K�H�H�Ћ[~�Q��'
����Y,J���ӌ� N2����'�`�'�#x��9:�+% b��	�'�LI#uLR'e��L��)�%���	�'�"����8�V�&S$���:�'��KW7W,`,���u�]"�'�ȴ��GIBjVG��PV�Y��'�0D����$ JH���GܜIB�'��m�#bZ	s̺A�t��(�f�+�'�v�0��>[P�9��#:��)�'��U{Q�X�~0��;��ݰHn\P��'H�(�`�@�Q]\��lV(@ZR���'���s�H�8��92�O�8*ϒl��'��(��î\�P8#@d҆�"����U�MO�k�L�G�Y70����?D�h; Šw�a�6�(L,T$>D���TʛV�j9�T�՛=�,�Vd=D�h���H�$� )֕-,����d/D���'��I6F�;T!�e&-p�n/D����E�,�a@�(_�TP$��% D�����ߦe����e�;ܕ��?D�� �2N��0���FO�����>D�� ��c7C2=^2����g���
�"O�UyrC�qx8!��F^��e��"O49"�$����OW�x��"O��2#��!`��ဘ�Hy��9�"Om��̘&d?L����w$���"O��Sc�
9��@ӧ���S�"O0�b$��J��a�V���5p� ��"O����?Ttss��&8謀6"O��r4� �d�$Ч���M�I��"OJD�գyL~4�v'��.:" @�"O����,[V"���ĎD^�S"O�P[7�S�cR �g�<x��T"O2����׸x��Z3U$���"O*��# 5P`( ㍐3�=��"Ob�H7J_�WDx���@k�H�<Ap�ܢ\��YA2`
kP�xI�&D�<��A�_��O�L��$N_y�<avAC�cEĐ���W>7��4 �ŏq�<�s�Y4�6A��eV�]�EqB��n�<�F@CS�̡�ViՁf�bYYuiKr�<��*ǣ,ь��̏�3vx���o�<�����wo���4kM��}b���l�<�ŉS)~!Pʶ��\��8�Ch�s�<��aѥo����D��:�,=�w��x�<eeW�Q�t���Ju�"M O�h�<�Eb~VՑ�� PF x@"KY�<��bHm�~���һ�HtH� �N�<	 @L�Bf�X"���
T\�æ�C�<ƤH
h��H��l̄N)p��!D��PG@4r6�\�U��F�~��@!D�tQR +c�����^�D4c � D���u/��$�S�	�r$�:�4D����È,�JD2cʅ'�I��-D��#�K�8^R��k�IǇ���2�G(D�����@u�*$�Qr�%�e$D�d �f� ^�10�aQ,g~n�	Y�!�ۘD�T��#K�OF��g�M!!��ā
�|�����|O������3!�d�c�1�����iH��XU �RF!�DJ����0�C[��9��.��^A!�!>�.Es�eƱ![��@�mJ�q�!��� DH���˔AO�r���!�ݱD�V��'DQ��Y�Lĵ�!��]*NI��5/�̢��5=�!�ē5hZP�4O���faވ�!�dϋ)Ը�77�I"�#P!��=z����BL�3V��R��!�D �X���J��!5~�b2�)Ai!�d�y~�e�A
N��q���ʿV�!�$X�_>�8��F�����T.�!�D	"j��Po@�B����f��!�ąaK>1&� g^�:D�#�!�č7-��]{0��R\�5h����!�dC��&�y�����%�)���!�D�;SD!����c��8���B{�!��;r�����&��k����A>N!����K�7vP3Waֽ:E!��,U���s���0r�&^�O2!��-\�|z���0{�r��Ug�� *!��5z�P��A2~�R<�0@)P!��@�CE���EN�	I�(�j1m�B!�d�J���3i��\�Y1,M�G!�d�t�v(p篎�uݸ�r��&,�!�A�7A��f� ���ȗG !��  ��fo�^UH���\j'"Oк�c��Sܤ�s)A��4܀�"O"\�BBד^�bQZ�h	�\ך�i�"O\��dMD8����H3o�xQ!"O�)�hHu,�"�Ƚf�$%2S"O����H�v��bÅ"g�x�r�"O�< e��c@�P�Ď�t����d"O��b'�&Q
�ԃ�oӘ6�0p"O�<Z�iY]��ه���h'�L��"Oxd�B%ϩ@���B�'%��c�"O<S7�<�"=C��E�r�,4q"O �����"_���*pb-1��y�"O8Z'IS{6�!��x�J�s�"Oހ �!�h��xs�/ǬǾ���"O�Ti4��X���4P�x%�7"O0��U$B
X�� &Ώ}0P��b"OzDU� �cxP���u"�(�"O�1 $S� �M���S�`Az"O��W�ܻh��ҋ׵H�H�"O��q�C;�~-����$t�Z(�"O�L�r�ˌ\?Ld�C釈����v"O�l{FV$k ���͉�T��	��"O�4��AD�0쨡�4������B"OZ� E�8H�@�Ѫ�W�HEa7"Oh��# �/�V���jCU�}aq"O�D�5c^[r
|�Jˊv��@�"OxI�w�P2{�б@���cV9��"O�4C�L�m>h�X㧟%&W���d"O�����C�eTXx�G�(��y�p"O�����X�?��)�t��1O�J���x����*���P�1I����ȓeDf]SB-^e�d���q'^H�ȓX�Ґ�VF�%y�z���E�'v���HJ���e�G��,�D�_�~B���^\cf��x`�A��%Cr��ȓV7tH1��YL�ZY��%@��-�ȓ"��!�D�T�4j��J&MR =�B�ȓ:��q�e�u`mJ�/��o��5�:�+e���*����D}+tm����3���]�>} 3�N��4��>b~��e�ٱ)�P�����M�`D�ȓx�f���lsP��cž@�0���|�@��V�ߊZi�j���D�xĆ�w(��5Lׇ;���k�f٩38^ �ȓKJH��`��ʦ䚗m��-2��ȓ
�+��
�. I�!��z�"O湛T��/0��-z��,7���"O��h�.��e��][�hM>�Qse"O4��!H��n3Z4��f�� ��Չt"O�2���kf���dR;M�d�У"O�}�KM�!�D��۫`����"O���PIW*J��I�hȳ9l����"O ��f�	�����/e�a+�"OVyK���9�ܵ�B�Km�~�H"O6��/
�,\L���E0'�`5�6"OMS�DV)�ʸ[goF�*�xhr�"O6��XB4L��H�tᐌ�(N#�yB�2zR="�肄#��uz�L�9�y�L��E2VKޥ0�� {���2�yh�WĪL����2,*�sBK �y�h��h���B�</`&<���!�ykW�.U��L& �F��5F�%�yr�6���B
�h�<�r)��y!�C� ��(X��C�ɵ�y
� ��Wk_!�
ҊR�:�� #"O*0˶�ơ,=ZIJ3J�A. �"O�@
�Ǹ*6��a$dZ.U��;�"O�)��9!���2hT�8dPV"O�|���F��Jh𑧀#2�0��"OV�i�i�(W�%�D�ׇB�@Q"OƵC���"$��|� �?���7"OQ�Q�Ӛ)��Uz���7���J�"On����ӊ,��a3A�	 }�,P�"O���d�T�IgH=�sD�(׼���"O�!����`s"��#�X(Y	�"O�r�.F:d�
L1�\2SW����"O^L�wL�t�x0�T}R�Q"OR�   ��   )  �  ?  �  �*  �6  �A  �I  ]U  sa  �g  n  bt  �z  �  *�  m�  ��  ��  7�  z�  ��   �  C�  ��  ��  V�  �  ��  ��  ��  3�  �
 � �$ m, �2 �8 i<  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��Y�1/l	aCڷUClM��%ɘ��n8UZ�&]�KR�P��,%T��<A����!Ez��F��\���i�L�/Bl!�S�t�3�a[��~��	9"O��"��IvH�	��EL6j�"�"O�aY���VAv,84jٟ.��"Or�{��+Q���A	L}>q�e����D,��ʆJ��t(T��43 �B%�!��/@��*e��-�tF�Q���hO񟶙��$ڸj7�7�B�Z�X�,D�|�7�g�Z���\� �~���|\�S����M�o�|P�L�"��uȨ�Z�'�L �r�ϓR�<H��Q/_��e���$*<O249��G�/{@ыR�%2��Se�'F�,���s��P5�!�s��5E~���b��ex���*x��ᐦO��HO�����`h%���a���
T�V"O��X"�@57�R�6#�^vʸ��"O0d�7@ 4i�8![���Z[�݊�"OaZ��R�,�"�;��T�xD�9X�"O�#�EMd@R�+F
]�� *��'Z�̈́	�dlqi۹&�ͻ���z���$=�����"	t1�.r��'�a}�c'
�ǓE�T�8c��Ұ<)W�>�O�����mF���& q��I!���F{���(aDQ�p�"Ǵ���-�2�1O��̓�4@�2�3�  ��B�G�ecʜ�R�.���"Od���/Ƽ2�K�Ȗ6nƲ��3�O�=E�TV*�\�b�Z,�T�k �N��y�J�v 
8��&�b��,��y2�
/B�R�x�k��1����jD���>��O~l��M�Vk��8ċ�4$��1�"O����B�)G�"8ȡ*�8U(Aӵ"O�l�E+Y�U>�48�Jӡ/�����"O�-r@�C�\ ����$z�t�R1"O�����'6��]?Y��R"O��³C�&���	¨|����"O^�{��G�
�d{�"hh *O�M�5g¤%�-ۃʗ1)}2�H�'��Xp-�� �\t��m�kJ���'ڴ���"F�<�b��$����'Hٲt�S#����!�
k�ܒ�8.*�6ڰJ獀�6vP9I4e�'@���m�|yZC�%x]��N�����Dz��~���IX�Չ��^k0NXǎUd�<���F'W1�%I O��՛"�Ҧ?�"=E��D��I���5yb �`%U;S�؝��B�z;�Hņc�6�����d�,T�'_a~���T_���+��X�<�j��L��?a����8������(c��BS�9+q�|��]fI�����ht4tZ$
v�X0�'�a~���[K� �	��C����᠂��y�A �f�\�iS�n�*����y��K"��0ՙj2�䫓bR��hO%��)��8�4={�I	
kƞ�v`[:*�!��·|&�!B��� "�� �ռ7�!�J�`�����<�R����t�!�A�_�t,��-�'!��;���|�!�dӗg"%pEhތ�2���jȓ�!�ɲDEz���$��o�ӉĔ=r��x�㉳	xR���7`�bAj�O��
��dh����i˹2s
��)���&#D�`X0�Db�����ᗘm-z�j��?D���"*��Ae̍�C׺r�0�鱤(D�\E�Ґ +��)i����㤟�D{���H%��1� @Yh&�A� =!�$^�yUVxi�V9eǒ�Sr/ފ6�Ѱ>�a!�[}���U����k��A����'g���r�Np��d�{�l�X�'���:�/��{()q�R�v����v��E{�'99�\B���T�]h� ��z}
���9�TPh��/f��PL.s?6ɒ��9$�t[D��
K�,���(�X�Т�#LO\�@�"J�O	<�PSe$*^���a5D���Q$_%&|غ�)�5.�;�G4D�d�Ǝ�D�Ea��k�d�)�O1D���$ޠ�����H<P8�H�ƭ<�$�:�S�O8*���~'L6��*��i�"O�$�LUaa�q�ƦN8eLy��$^�<Y�~�R�� �-I��{Ώ�"`���	J�	l�@b�j%N�

��n@�8#�'k��4	ҏu8Ԥ�TCֶ6�L��˓�(O��#�1d�����BS`!1"O��@���.�HU�1GR�eEޙ��>��)>�S�'~|mc��ǃ>@>m1��@�]Td�ȓs�\��Eő�2��Ɇ���̇ȓDz�8`�Z�(�8=���B7�0�ȓw�.��!�U$��Z4E�}DD܄�`�0��2Þ0�쉁ōT�(�ȓ' @����	$Vd�T��	�v���S�? B!(d�ʑ�xǁ��W<�D�xb(/���%��1��[&H�8a�"N>4�F���i?�p�ҒR7�m`�
VUԵ�EK�<���+���p.C[qK+���D_�Q��7�eq���H�)�ȓR@Q0���*���� 6D���ȓN��U�@�ƈu[Q1��ο"�:%��@��Ϟ�D�fq�(�or�ȓL 0�	AS�8�DI�F~��ȓ;����g�ӱM��0�i��;�m��}�|��GMQ5
�-X���&T�(��n�Z��@U�]d=���д��\�ȓ_��e���΅S��!��.'n�@��	c}���.A	��0�!P���z@
��M����s���C��5!�m���	 h	�"OjiBCN��l��B�]�!�f�)�R�̅�	,��"�j
�>Q�P�����~V2B�IKO�
�F^�%v��%ƅ�>SDB�ɞ|��D�g���d`�h��+B�I6
P�S5�(��!h���\��B��ӟ��'L��$(J���-܅+/��P /*ʓǰ<�� �Tx@�1c�D�+ƭk�'g�I�h��h��Ͷ	F�B���(�MD"O�}��%�, ���U����{I�<I����b׌ѓ�"ڰatz��[��C�	5�]I ��D��=� ��;�V�=yÓR����G��<��M�`,(�����?7E	2(�V�ì{��=��Y�<�A�We��}�֪��5��=(�ZT�<aWob��r�LN�3����FS�<yfɝ7�*�:��Ͷt �h$Rt�<���؜9�Q��	�5��9b)�o�<1A+U�����F��!шP��j�n�<�U!�2���boӱuH�]a׭	g�<��n�9���I��-����/_�<		�7.�����f5�dx# Yv�<�w�
�������*� 8G�o�<I�i	#�Y�^�,R(YQ�"�E�<�t��!Dk��X%����t����y�<Y3&H|�6p��i�D�0@��r�<QT	�Z��r��+�0%!!Ak�<��&G�k����� ��'�	h�<i��$`�zH��b"x6�Qc�k�<�a�]T�t�tMU4R0�a��Ap�<��E�&F�����
8`���u�<i�I҅D�����e�!21,�Q5��n�<�GN<����F��_��#��a�<a�c�(��q)��\1JM�Qx��^^�<�E�|����挭.�&�P�Ht�<9�%9\����$G���q�p�<�r��1��u����R5�ea�<Q�щh���Z%K��2��MD-TZ�<)F��~��Tc�#�m	�}��V�<�W
�w^콂 ���d́'EIN�<i��ع"zB��@�cs�:��H�<�WMӟk`"-�S��j��
�Z�<�V��(gDT��@�=u�B}��b�W�<��΢<˜�����`2Q��}�<13埦ZN`��N/D޸�p�O{�<闇_�F��,�o�vG��R��B�<��2u��8#�E�_K���"E�D�<�Wʄ���-I�ਂ�&G�(B��1"&~H'\�W9��!���QBC�!Kz�$��,L��,!'d˰ �C�)� �����E\�k!��$SH�"OtM��imƴ"@N7 OV��v"O�٪��`�;r�[93�@�"Oܔ
5#ԙg���W%O/\��@"O� �tl@�~r XפM>$�$���'�2�'r��'2��'KB�'6�'�@�A�E(uYT�+���(22 �!�'�B�'���'pB�'�'8"�'�H�"�Ȃ�V ղp	�A�\�r��'���'���'��'	r���isB�	ߌ5j���F����o����O���OJ��O�$�O��$�O^����Oq	aP㚂��!CcA��$���O����O��D�O���O��$�O�d�s-J(�w ߲���+	"��D�O��$�O>���O$�D�O���O�dJi�\q2P��)������{�V���O����O����OD��O��D�OB���<~�ܻ��� iԙ� �7���O,���Ol�$�O���O����O��m�Z�[K\"� � ��8dZ����Or�$�O���O��D�O����O��_�Q��8l��5�i���@�����O����O���O����O����O��d_��8���M8�����'ɘ�d�O��d�OD�d�OL�D�O����O�����܉��U</b��k�;8����Ob��O����O��D�O��D�O���0+��e8��
 ��s'�A�����MK���?Q��?���?�׿i���'Z����Cʗp�~S���;�K����������$[��qA�	1 0
�Ěs?='D0Y�-)?�E�i��O�9O�D߇o�V��� �a��8Rt# -t���O^)ا
o�����Td���O�"�cӬؘ~τ55��7*�mc�y"�'+�	s�O�6L3��4'g���'��+xI��N`� �#��>��1�MϻI���u��<O�ܸ�Jt� ����?Y�'��)擽0y��o��<iΈ�R��U�p&įN����A��<I�'f@��hO��O�i�FU3�
�a��ȱ+$��#�;OV���XԛV�۞ט'��=�R��;QɁ���<0����	f}R�'�;O4�9�$��D�25pyp�	�	��d�' �h�>00]����H���X�4�'H�� R)��T745a�Kڒw�x�T�ؔ'���9O�Yʓg��9���[�DU a�:�Ӗ<O0-o1%������4�L�:ńL�v�^��d�;���#=OH���O��dÀk�b7�1?Q�O���eF޴�D��:	%�Ā$C�2ah���CC�r�l곤C�}&�|�F��T$4K�+ĭ$R�9�A�8u@�8+�@D8t2��镤��*#������d3(����D�d=�x���%u�����-@Z$��� �a:�
"ݓy	ZI��i��hf+��S����U�b��{DТ;����V)&sŹ�OK�y\,}��ݥ9�E�sDV����14�f�����jj4�� ��}���H�OVriK�O>bb
ȸ�,���$���^2�TCg%��Q���YqJ�[n��d��
�h����O�s��@22�	OgTu1ì�'2<�Rg@�|���'g�'��`8?)�+��x��uyw�F�g4��2!V٦a�	��ԅ�����	ßH���?����]�D�G�zT��ڒ�b����u�i����jӊ���Ox�D��fQ%���,
1e�����F���	��� 1�4%Q�4v�(�z*O�d�O���d�O�H���U")�J�����.Ly�I��ܦ)�	�X���(!�՚K<ͧ�?���E��}s��U�n�E:��N�����V�p�I�@"�?�I� ���<i�
����K��5�$�r���MK��uz����x�O�ғ|Zwi����� b�&���A΁M ��O�A���O,���O�R)�i ɝ-}^���M�_�P�ڀ쐚r1�'���'��U����֟H�Sk��7�.�h�6���'J�\66c�p���(��ay�"��YDt�S* �����H��p�G��>n��?	��?�)O
��O���'P?�Ȏ$:jSFإ)VX��u�>���?a���d��e+'>�C阌;Q���ȇVֆ�i$���M���?�(O�D�ON=��I�"';DI�0��;@ubw����f�',�Q�h�$G�)�ħ�?��� A�kn��Y�+]U<*��q
ئm�'�B�'x[��Iꟛd�l]��G�(�b""� �M)O�D�P��Ӧ��������*1�'��ՠ�+�/:�&I�m� ��4�?Y�j\��(O�S�?Oҭ�4E�0(�jj��Z9β��P�i�hf�w��$�O(������&��ӭ)�ƌI�lԀq�B�$�ǡ�<���40��=(O�$�O����On$���q`)Q��$="�0Xq \���I�h�	�# PN<ͧ�?Q��~����K�7I�	C4")\�zl(2\�L���|���.�����ğl�����R*�� �G?4`���4�?AsB%�����'
�_�H�#��6h�ف/�]�r@�Mk��r۠�<!���?Q�����~x��a�PA��c�ٌen��!\W���������'�r�'*\ !���4*���\0�r��Ø'q��'�����K��Y`Z��~>�P%-���l�{ҫ@��	� ��I���?Y��#}>��l�2��܁�`��,ˎ���f�+K���?�������OB���E�|�'a�M1��F�FƊu@U� �ډC�4�?ɋ2�'p:a3%�ējI¹y'��+E�r�	G�lZ����'��($���ڟ,�I�?�s3��V�V���*�A�K²��'�� ]/s�X��y��� @ePլLU�5�F瓈媜h"V�����x�F���՟��I�H�[yZw(�p���}!�yX���i3V��O��Q� 5��`F�����n� ɘDh�W.^f�O%Uۛ��,� ��?Q��?�����4�V�d�y�F$3���'-,��7i�0[s�o��� �Sj:�)�'�?ɐ�	2R�m �@�9���ŇT7����'B�'�&E��W��ܟ���[?9£%�f�[dF�K�feV
WL1O�}���k�S��0�IV?�p��#�
u�c��H�ĉU�@�]�If�\�'��',r��K>dӸ�/��V�)�!��*��ɥF۲�K�.?9���?q/O��� 9_69R�/�'B�\���!�&p��8�E�<9���?Q���'�E 8c*��ZC�\�e949�U@H5O�<�qT���d�O����<���.�@}�O����cד��,�ՠ)�I��4�?a��?����'�>�֦��M�%�S�A�����Σ~��Ԯ�}}�'R�\�|�ɽQJԕO�©	v�)ygl�?!��i���n7��O��|�I�h�x#�H"��%��%��)z�!ZT,F�6��F�'��⟨�S��G���'�"�O©���N�uƌ�+�AF8f��I0�&2�I�����#��E(b��'	�0l0��˓�1��f�.l��'_���62�'���?��:���P�LiNQ+���Z�b�>���X��Hm�S�'HVP}�c�$G"�A��)s��m�G���� �'��D]�����r)%E���¢C�!��lS��M�p "��5�<E���'�ݲ`��Y��@J�H�GN��bb�l���O�䑝zx��|z��?a�'���{�#O�_�d�� *֡��R%d7,U�O�'i��ُ;��bf�� 1.��� ƔJQ�6�'N-4W�p��ݟ���Xܓ'���5j*�J1)�+&��Q&�h��E(?��?Q+O��ė�:�)�j� ~r��J�D�D���<���?����'���S�c6�Z��t,�V�L�*j������d�O*���<�:�$���O�ͨtN�l=��	�
�}\����4�?���?����'���h���M[��b&dc�*ݚT�,�S�Qi}r�'�T�p��.�\��O�BaGA�<��QG΁=Ԙ�;�i�)S� 7��O��0��gl����;�$�/^J���r��;o�6�m����f�'d��П(�B�Wo�t]��+%�Be����G�zi˓�H�^E�d`�}��'�85e�1՘��)�.C,RQIaĔ`\�i��
���	ʟi���՟���㟬���?��u7b���y`�K�(Z��B�IC(����ON��s�ʭ1�1O��XUr�F�*s�m�R`#E�U���СU�2�'e��' ��\��ʟ�Y#
�I>�D�"`Ԙ������M��Hh}��<E���' &��G��2w@-)��6y�v��OzӜ���O8�D�z����|����?��'�8@[�BZ�ge�QYB@�	7��I�e<��5,=�1�M|����?��'꾹�1n\�	R��Q��I��HS�O"�;���<Q���?�����'Srȣ��ޯk�<l�@i�i��x�O��:V�D�5l�	�����Yy��'��(�!��]��Q� �BE��)���#��������?Y��K�ˊ�������A�DDh#��`@4�W& ?���?Y.O��$�����5a�*�I֢Q�%�X����=�*6-�O\�$�O\� �I�9�TP��g��)k����ّ&J��r�0e��P���	埌�'���ɥ;���$J7�I<F( �L�sH��!�U��M����'1��ЗL+0�jM<YU`N8y�j'ǚ'�HQ�S�����NyR�'Jx# W>}�����Әp�L�9�Ŕ'hn���b�~��}��'�$�S�������	��!��zۮA���T-��	��Q *�ҟp��Ɵ���?m��u�L�4.���fIԴeXD�z������O�I�V��;�1O��F�[��.PRF��6+B��0鰴i^�ӕ�'���'B�O��i>q�I)x����"�|ik���~	05��4/�)9�+NP�S�O�r��W=p;���7߆���;V6��Oj��Ob��p�<�'�?����~�bR��]��l�$|�ܠ��F.o��b�Р�)����'�?���~R��5c0\	��H�} I
G����M��=o:-O����O6�6�I�cr��K�
�Y4�2o�N���#�p�0U�In~��'t�^�����UW�ZRJ+6I=˷��(��c&��eyb�'���'��O���s3l(���mv�����Z<K�豪E&Y�1N�	����Ify�'@�cVߟ�1ݹ�E����h9�����M{��?Y���'��$�t���ܴ��m� �8�Q�l�o���'���'��I����T@�`���'�6�����)Y���SG�U�A!�~�p��:�IΟD�d�آOĪO��oB.o2�zE�ï8A��鲾i��V����6�~i�O�R�'��,8~{]+ed��&�r,��H$"��b�|��$�8��B+�~j��L42�s��H��`�"��G}����9PJ��'��'���U��ݖS�5R��Dh ��%�t�<��?�ħ֠#�]�<�~*�홨}	Bd۲&�>2`���˦�j��ğ4�	ğ��I�?�����'�D�R��U3x�<9yB�ݖzC��{Fdӎ0�$�@�X�1O>1��+׀ �8��%x� l!��M�$X�=�&�iz��'b�(Y'g��i>��	��h�H},I�b�q+�@3� �9nq<a��F0扬(�@�0H|R���?���K�dd8��2&.�u�	\Nh�z�iF��,N:�����ORʓ�?�1]A%���x�ā�Qcֵ=/�5�'&uZ�'���'2��'�[��0�L�N��3���R'�$"�k��Ȅ�O�ʓ�?�-O���O��D,)���x!�\h�Ԃt� x :��<O��D�O��y���O&��<Q����:$�iO�G�"�2U�L�Yh�'M�Ni�FX����GyR�'���'�l���'�Y
U'����,�f�l���A3�`����&Z$d��O$˓(�֕ppY?i���` ����Ņ�Ш���۝dTn�8ݴ�?�)O����O �D�z��|nZq�aQ'�������	�>Hy
6M�O��d�<!�̅L����|��?��F莚Z�PH�m���U��L�TyR�'B�'L���'�s�@��8�q#Ji$ y��k"�oZgy�l ,��6M�O*�$j��I]}Zw7�=k]T�c�MҊ=.��'���9��ꟸ��A`�X����,�R"2����А�iF"�X �*I�7m�5ӂ�mZ������<�S���$�<Ѷ�K�XH�ɖ8Z���(���6D�1�y��'���N���?Y���!x��x�&-J�0rt%K V
�&�'��5O  D%�>y/O��䨟T�T��8y7�t��D�IT��"�'���7Gf��?i��?!G��	^�+��;Q\|R(ں\�61OHp���>�-O��$�<���+wo�$v*���F�	�`A[%�Uj}���yb[�H��ȟ��my�(F���bmU�E��uB
�F31n�>�-O���<���?Y��N)��3��?y�ޝP�	�-'��r��<����?	���?y���d˱n�tΧqW*�Wɖ?X(�W�۰���m�gy��'����$�	ӟ�j���~�iH9JZ>�y�M$���2`�U[}b�''b�'���p����N�DH�w���`�sմ�v�ݱ"3��n�����'�2�'��J��y�^>7M�DXaRU$U=.\�9�g돮r��&�'��U��RW� �����O���0	 ���!�Z�C��8E
5ʥ\}��'FB�'��Қ'$��9Fj���-��lHVM��g{��@
Q���m�[y�Bտ�V6m�O��d~��)J}Zw�PU!��j�� 䇹�X���4�?��K�
E�}��s���}�$�G�>����˩<��M����h`:�M���?�����pX��'�q�1�j�襹��*9%��Z$�s�й�8OH���OZ�� ���?-�m�8A�9�$���k�&�����M���?Y�'P��FX�8�']�O�h�IG-!p`㊟���AָiJ�U��y�/l���?���?a�iJ3s�Q:B��3pG�H�Ʉ�t��v>O&�p���>	/OL�d�<����ˎ(�L�����!��@�1)b}�d��yR�'["�'R�'t�	�mgJ��)�?[��Ċ�#�<u|<D���Ĕ��D�<����d�O��$�Oހ d�˪�F�'��	0rJ���:2��d�O��K�^�6��OT�E{t}��>�Ҕ�r,�*�m��ረ�V�"^�<�����$�8�����σ՟L9�lɑ,�n�H4���`-z�������O����O�ʓxw��cF��D$�0��\r"�[Z����4a�6��On�Op���O����j�Oz�'�8��c�D�t�6H��*���sߴ�?	����$A��&>Y�I�?M�E���);4i!1N�a�1�4�ē�?���l�Z��������H'r�Xj�\�t`�PZ>�M�,O�,�#ZǦ�b��$���Rx�'�XLJ͒"(�4�!1�S��,���4�?Y�upd1������O4h(�Y�yYZ���\fp2ݴgی=�i���'���OZ�c�x(!��$ܥFY
l^�Rd׳i��5nڡHT�-�I`��d���?�����T��� �%k�H��a铍R뛦�'�"�'��`��=���O�����|ёM�>�,8��? �x�fӸ�O�pg�M�S۟����`�I�YsvU[��_">P씙��/�M����&������O���?�1@h��,ʂI.���ᯋ{��'P捺��'^�	��	ɟ|�'V2�qD��)��8�B�*H����G�VO^�$�O��O\��O�p��;�6 HG�S�T"�a�����l��<���?q�����6k��qͧHa��SJ�P�}4�@5�:��'���'�'���'�Z����'c��k$Kс>J�;�,R�X����J�>a��?Y����D�4L�@H&>�RT�16�DM
V�J�;�� zR&Y=�M+����?!�/�z�������&��闍9~�{�J�to6�Oz��<�')Lx��O���O݊7�@qE ��B�\*i�2E �$�O��� ���(�T?���%Q`�!Aj��K��h�pӒ˓I��Y*c�i�맪?��Nu�	��ܺr�#?��Yb்*+�67��O���[,���0��0�'/Բ��@�+
d@Y���	�W$�7-	��EnZПl�Iɟ������|��&SǮ��@L�%A����U$O��?��Aʛ�?9���?1��)�O2��FҜ=�|��bH$:���f�����ҟ�I�q�L�N<�'��I,I�ؼ�c�Ű�x1�ǀ7�t7�:�I��&>��	��T��8612�%�(�lx�ħX�� h��4�?����[����t�ɀD�p�m2��y�@D�%�l7M�O.0���Obʓ�?9��?�)OV�� 4XsA�>)� �xb�D:�Ig��5cw�'���I꟰���˄l�,�ۤ���TH��A�3'�6��ly��'���'��'�,���'B���^sU� �^H�����rӊ�$�O0�+��O2��E�&��Ǹi�j��׏c�hX`׎�&z��AZ�O`���O�$�<���\�������D5����I�uvZ�B槉�M����?��������O"Tu� X>2�6��U��9\7�\��4�?���?9�k����?Q���?���&���Z�'iPAb7��LD�D�x��'����\$\�0�y�����!	BD���gܝnF����'��-;��'=��'���Q��X'xn������4 <Es4&� 7��Ox�d���8ك���U�*�`(3t
A`�T�2�J�o��ŅesH7-�O����O��i�i}"U>��kT�"MriqDm �f�n�	��ݻ�M�Ď����'���|b�'�$���N+"O.��V��T��y"i���D�O���F��f���O��'�?�'.������;��d �k�>.˔�&�I�d7�AK|����?q��v�t�z�/�9C��]aR����m���i�b��*+^��'��꧳?qJ>q��_6�<	�'h�ay��n�/F�|z"5��8�I����py�hH���"�?}���jA�V��쉤Ǩ>���?���?	�����o�.�A@�<E��$�V�:hvX�t�|"�'R��'R�'\���֟��3�?f,��&�Ȍ���1"�ir��'�r�|��'�R1����4i���r��>uڦ��#�"V��9�'�.�R逩.����O(Ω{��m�`���:8t���'�����,U+.6D�e�
�1��p�'�Xyh��h^���&��Q�ұ������j�$[�KA�{���f۾�����D�����cd���lY�Jܢ�B�J�1�����ǼR�NEʇ���&����3���W<"|KtiR�|�d�C)F3�HD0׭��R�ʁ2�nǚz�Rd
O��@����m���2%�^E����O���;d� U	"�V�,~�a�h �I ��:�*��r�]h�������$:9 ��'ۘϿ+gb��"�b%\���y�fԡrv����ϧa�PT��oĝ@	F�3\fV\���2Cf�,/�G�M�<3�l�2$ $3�l�rҬ�$5TҘ�C�'q�����x�O����Y+�"�����-/t�"O���D���Y�$�\�֝ۡ�	�HO��@�����,Yͪ	[4��b'�i�I͟��s��NNa�Iʟx�	�[Xw���'G����&I���p��:h��,��b�O�3��g 딍�
����č!-Yl�PrH� �>m���#9t�9�#C� i���?�=Y�)c�@�pƾd^ք�u�K?a5JUɟ���c�'�剣'�tXF@�.��9S�%C�rdB�	#K�Y�#�#l�q��+ )-�^�I���?ŕ'�(��b�:9!�"��o��ᰱ�S�C*q�Ѣ�O����O��6e-8��O��Stf��"�@
"g(u���0��
ܱ/Zj�!?=@|����%y���Ó&-0����
0����É�;]���x4�5��	�P���O6����Y.S�
	��.�	���5E%ړ��O���:,V��RD�V�z����"O\� F��h�v�b�fو��6O2��'��I�ndDPݴ�?a���ن��9��� jVr�:��.Z�ˆ)�O2�$�O���E٣|� ���O8\?ne��|:Р��W��H�D�Bo}����J�'3ni��Ϋk��h�W/Xޠ��V�cl,ꓪS�z+|�ᬓ���5V(�B�'� )���)�֌y�N�D�|2с�%s�Xದ��L�${錳�?q���9O�`9���5R��Sꞯ/�`�p1�'�OT<����C��Ĺe���� D:OМ�4O
ܦ��ǟ��O!� 1��'3��'�Hpd��9�2��S�OU4Y�.�v$`�k��/�T>E�|�	$�V ��UIU�pkq���=�R�P,��,�U�O>E��pr|�Q��=cEF��� u�6�7�Ǚ�?a���?Y�����'wJ�X�m_�B�B�� �y��'��}�*�-,�� 5n�sbT�1�	<�OX�Fz"T>	�'	v�8%���']�T���Ȍß��	L᨝�`@�ʟ��	џ`�ɥ�ug�'5r�V!T�$I{��MC��9sK��~,V�* ��j�"J�m��x��	�4и�R�Ҳ�Dx�aɦ{�~��k�H]�t�O��Ybu�'k�Ua�*F1ug&`� �Z<���'6��3�Z՛�-l��� ��f`��LQ�>��D�2��0 )�"Oni볥ֶ۰�`Ҁ� �fII�'�����M't�~mo�OF\D{6��+�lĈB�G�d��I�������E�ϟ����|��Ό�&5$A�g�L,/Ҽ̂RIV�"Mc0cܔL6�|�q�E���<�%�zZ���r��1"��&@X�)
�[!�X����5V`�Ѧ^d�'�&D+��?	�e��v�5Q��;@��5hՒ�?ɏR�s����
*��:�X�&�����$D�|�e恢D2��m�z(2mh�x��)�O$�)��T�s�iLB�'&�R�8 B�j�#m�f��'�Q�JEd�� �����П��0
 ���<�π "�"8�q㛴|zl�v剫V[����(ڧu�P���=4{
M�"/�LC�<FyB�ˣ�?q��)����[��Ջ2�����Ty!��0(D���vÍjwԝS���ZTa|R#���13=���H]�d� D� S�Q�$*$�±oş��	G�$�W`R�'Fb#ʇ><j��OB9f~d�)�b׳&&&��p%��%��s�XY��"��~���;xU��'Zt�`Q��Ǽ\�t؀waN4h�����b�|Hz&-ɗO;�>�n^�s�,	�$�C+Z~@tMO�x$�(���O�$$?��d��?9�ع3����ߘ�)� ��<y���>i���/�V�H���:+1�`�w�@D�'	�"=�'�?�ER�	@����H'.�� ��C��?���r>�c����?����?��*���ܟ�A�6M6�(�DЫkؚ؉�｟$[C�I�6Ѱ�R��ί�p<q��4�Nu���#��8��Zp?��LN;5�F���BUW��x�E��X�Aj�e�6�*���	]r�]�2�'�����O���l%�(��a����+�����ȓ4U��p�*I���/��j	�YR��d�|�*O��ɂ�զaX���:c�>� �T�?c�%#�Vş���ƟD�I�g+he�	���' FYu�ҝV��ع%��xH=�$R<�~�H4�k?��8�F�Z����lK�?�����`�C�Ig!�U%�A�Äݕ%��b��D`X����&�үd��"�lÈN�*����Ֆ-^L#aJ�Q�?�C�s��U���D��4N���)��f0D�ta��ҹ,5�Ɍ�hp�6jn�`��4�?�+O�r��)�Iԟ�O�|ܰQ�P	]������Œ�d��O0���'��	��y��T>�`#�4_�r, Ҽ@���z�H:�v�D���&�F�Z�K�z~�"7N�0�Q��S��OX��(���O�\(7�O�
� &ߧ\A �TD�O��"~�8�4T�)F��mq5A�-n���I�ēUDZl������k��Շ{�4�r�Y0�i��'��Ӓv�܁���,��#(��Iї�ưu��+f#��(��}P�N鴐Zf�!P��遾��I8��O޼C�˿S㾕���˔|� � �/>�vd:�(W�<�Z�Ȇ�?�Q?��Hb�����U���ck�,׎L)���O��m�X�IS��T�IҟS��%�z,��.R�BM�JL�@��Yx��� L@�����0����*}�Ǫ(���|C�O^ls�"��@�W�Y2y~�u��b74��92톊ܦ6�P���9f`WP�<���2:}8A��R|dq�q�<�%%�,�������B�BIg�<yd��-L�z����(_V����O�<�խ4O<0	TO��x�]I�<a�MH  ��A�˖J��+�� T���d�[נY�TD�?�ȵ�si6D�<24��{Ah���� 'G+NO��y�ƈ{�p1��Z�dfp �Va��y���k;̩���Y�r]�%�B�yR�J:nN���A#]:�xţB��y�NN�w��$�ÒV&ne��i��'�n���͘ %x�\��5C{zq[�',���kz�*5HR�V�<{DhP�'|��K4��Z�k73��R�'�d(����L��!餤�22?%��'�N�����޺���-��3��u��'&� �E�ۡa\�,�JN7+b����'�Ji���
��jx�)�#h*�I�'�Yfm�'3 x��@�=JYVl1�';:�C$�P�h\��X%'O�G��h�'d� (%�ԛD����50���'hN��E*BvT��$�;���'e�A��X�2�6piPÎ�[l�[�'��e���M�x��t+�� 
�I	�']x� 
Ӊ,BJ���?y�h���'S"ՠ�]�D��!�'%�r��'��q�tb7:ώ��q�ֺ԰��']J��W;}�QD(6bD��c�'�BY�uD����0��5+b�5���� .u"g ���P{v�5
=�;3"O�{�M��z�ys�7
,��"O\�$�-;�"=I�m?'d�[�"O��;6���v��s", )�lV"O
T������X������4 ՞>����gX32-�U����<�
p���&R�}:�8R�̱�|� Z����@ 7*�c&�ȇ�ē��1�@���Z ӕh�ȴy��nt�PH�=I6�sƈ\{�S+$��m���O�z�a.K~�tc�!��)%�����P�9����/Z6�bؚV�ɩy�
�G}Ƒ>k`�DefM�"�L�7k�k���^4�V�(��3���ri\� �dbE����5k/�@W����Tj�f4����'V�
�s���
*eFl"�XJ�|aӦ�O�QkB�E0Cq��ABaA<#�(��q�	�f$^1O�<d��16��k�S�4�r�]ґ���Qa�;3�R/r8"���/?yqjV�:,`e����+�2p����nj@�ۻZ;�Q�@���C�`ϓ|���5
�	����,y�1��*gz�B2}�GG$䅹'�ԪW�&u)1N�"�t�rBNF���cJ�r+��N|Z��״
mF	Y�Ş<vb��F/;L h��g��zb���%ǚ.|b�� ���9Fha�#.�*�O����.X��Q3��'�z�.��`@��<�6�R5��G:����%& ��샧e��; ���<A��<|R��;勄!H�4(+�@�:dl �c���O��"G��f´�J�O�6B�6�Dߔ_	�T(��^��
����L�( "i�����$���̓� �P �����ɼ;3`
V(��3#ƚ�W�v}��DH~bJ�Co�����p��Mb��	*�5��c��@;�c��(�dْ�'3&!Y���w1v�&Egݩ��,¬	��p��Ml���;������<~�Pq���Œo��0���աh:��K�-�`���':n����K�J�'��K�d\�0C\!�:ષ�^�{��a�C�5L��t��:�脹����o��x�o��7��C�.��| Hۄ����&zQeSh�X��$�dC/�ug�x�)�!Ej��kb�R��.��GBD}R��A|��#p$]�l/y��',tL��O1 �R,� �A:8
�3�{�(&\�qO4I�'0�X��a���:���n�+�65� ��?��U��li6(Y �����@��Xg��zI������Y�^��I�ܥ�SÏ=Gz2 ��{�ώ}��nǫ;c0�q����j�'����e2��!6ləx+ڜ����N@�X"�'C������9�	�՟��<���w��P'��N����(E�;h�(r���!5�N0���L`R��䂖O+�3��۵*�D8���'�.i��
X �M�R�(3�O�>�S��9+ ��"��]�.e�l	!�CZ؞�	ѭ��m�$ט=0�2���L��
"Ȕ�)��mH ����	�<h��'���H���`�O$ C�����=9�,"7��*��$B�(I��'�FPyv�I&���O�ظX �P1����]�rcv�J���k?�uE��OnZ���Gz���$�F���U��z��1��DQ<:�r��dL��̡�c��H�ġ�O���ɋ.[��j��'3!�0�G�dϐ��-���p?����D���� Tgp X��Qn�ȑ��(��8��*Dzӧ��O���2!�M1��4+�=�$A�8a|��Ij�Ń�h��4`*��\���I!l��{utK �R���� 9w����O�����{����F�#�h� p�U`�Hܑ]�X����I�;�F�!�`�8@��Tb�@̱X��@���\�y�`ȐJ^��8���:\��`�����˪#?�3�Q�*1Q��:���1D�ĊK��p�<1@�Ԫ4�qq�3��g~�(�����Z4a�hR(�P�$B��u����}b�f:m�Ϡ,�0����
/[FhAc��æ.��Ik<l�'�d����?ͻWnI� ���j�buR�-�i/r��/ZQ�t��3:�Hx@��8;�>i�6�U���1��|���'n�rbH�:I��O<Y�H��6�*XX'��1|�.�����u�di�4F�x��s�����?E��@Ip��%'�(!�Q�X	��	�D��Zv
��P��g�')��� ,)�%Q`�lj<(��OR)I6��|Y�yR�-5���$`��б-�tJ�)N�p�[�y9�fD��p?�g,~,P��b
S��0�ɏ�N�f��,OLDJ&��.:�?Kn��������$�����7�޽  ��m���wO�%��.�,����FI�L���A�n�*B���NP���0F-��OT��?Q�Q��J�QI�.�8�q(C� O*��B-��$��P���B�fՃҮ����K�5{M�0~"���O�=*v(�>���O��(*���1x�*a"��'��´�0���Z�J$��a]?b��;�B$P����	�0�;A@pF��fʕZD��&��[ff�Wx��!��2Y:~�#��� ~�`L	�e�<�P-���BX��sִ0ږ׽<��`y��U�v��΅�AvP�:C.\��j/��?I�#\S&� 1��*Vq�HKgD��a��2a*2��1A���n� o�����\!"7J�LTH�is'��;0y��	��&A��J]���D���-.���N�Ge|�J��+`���0��<yP�W�t� � �C�Ax���n�1��T.ш<�$�A��'?��L�U�h�"-uȬ�������/�$x(��7����1l
�k������H?Q��e���� H9��,w��adk�Rβ!����eF��0��]=6�$�Y�H8��7���i�'N� ��0�,|ZQ�M�2-�DH�E4�H�O,}XU�D�S��3�b�q���*�)�X�xu�
3#��X��,.��0$�U��1q4j�5���O��V��q��qYR'�#A*R��՘>ᶬ^�T� S�a��'&j���8�@T4=
,j�Hvf�݉�mE$�굑g��� f�bcNʽZVE�d�N;9�����v�`��W�Y��3�j`���b����ě��<G��`@�ˍ,2uAS��g�b>mJp�޺Zq�$3���W��E���F��lJtÎ}�N-�W�V|�ڨ0�jG1��ɐ���0y�z����}��P�*?*�'UFP슥E]z����K�I�K0,�YW��J�p�H0.L�!��ɸf�Dʟ\���1!��%�%�ׁ$Z��bᖤ5�l0S2�[��`�Q0i]z(�tC�:0��(��%0�V)\���� K� Ic�֓v�%�'��i���gm&I�"�+����h�4d���8Vf�`$B7-95H�$�N*�L��DԮs("�Q��P!1�a~�F�X<X��fa�;�|I �� ���a^,ZQ���*F�4��ŀ|ٓ0-����I`pb4�t흵�ƙ��̆vj��:$O���p�L�X@x s��Hp�$�W�-��tȅ�4ϐA�'7�L�p�R`�<�;[��8T�O8���Ը-����nX�?�<�A�'$�l��� 6C��#��(*M�4! [�"���àI �:�Ύ�]�a�&��.-�ӊo�y�c��v����D�%8`\��f���$��`�����&C2v��u��Q��*0����4Ji�l`֥ݳB���F-qL�u��'UZ@�R�ʔ)���{��L\*�Jѭ&h��M���Y�W�ܴ��Oq��x�+�C�8����Xh�xo��h�VH�,E�!���2�=�r?|��S�֓[�f9�Eر,/ P�q�O��H3�Q�lB�d{��[>H�+G�|"@jp����39��� ����X-.��8;*��@Ex�����
��((�G�΅g&���W,H�K.p��$��;��]zb*;<O(uєA��a�@�h��;jm�3���:�(��3\�8��n2��5$i��yC��7�`扬V�(]�Fo00Ĕ�2NM�B�B�	�f�����"-6ܐ����n:,�x�Ι���!�		H9�0�&�O�s�0�"�c�Ճ4�C�#�bqE���<o!�ԁ0�Ӿ58"lۆ(��H%)'�?-��#ôi���I��h�t�'t��UI O;*��Pg�=+����I'�
� x�ՁM�~�x�`� ��?��"u�N�� �� i�ܡ��i 0�(�� )ܠ��a� ��c�V����E j��9�ZJ~A��@��i�w��T  �quT>c�Pʄ�� "w���E,M�Ԑ r�&1�	2.�%��A��ѓ��H����'�$oƆGD��:�K\8>\1�DJ���U����?F�oܓ�xb>�R.O3=Z�*#��6�B�q�,%`�5ѧ�K�r���c'"�<7HQ��#i�qr� n�0��
�69^O\  �C�b������G�r�̧.U��U���W3 ��S��8p�V�9��HX{1�}�����?i& ��{c������Y�"�9j�����䜱MD2,��	bQ�β3Fr�]5 ���[��^���Ê���'���p'�5;�45k�����>A��^	��qr��L${a†V&�U�p-�#_��S��0姚�+	��fh�N����O��5hݘN�p�
�ڤI���+�7O֌�p '�Ɉ�M�� F�t�l�0a��B���1�+Jz��)���j{)X�G�/JL1O(Z�O��p<������'!G�-_h��0CNQ}� w�b4�r�ǛL��5���=L(�#)W���I�)��B�"�i�Y�TIP��  X�j�S� aS��`;��{��z��!(j!,4K2ˈ�����s�>P2��S�|z���&rS�Ic�]�N���4lB����X2)��6��֯8�s�l���S-�<J���@L�tKS^�|�pU"͡@���<�!�/���� �LOܙ����<V���unKB����ɍ�(�X��gm�<i�Ǻϓxޖ����0 P�?�B,TL�0嫄:%}r� �̦����_&|�R��_�B�����IC>II�Y(!|Q� Z�):K�a��Γ����%�6Y�:@��&!��	ܢ(Y��
�wH9��!��k���f��5_����S8�����5.V|Tx���ß��@��4y+e�=r����@ 2�2��(\�R���d�� w�H�@����ˆ�Q"�y��4�"S�
�5U��lyס�6ؘ'7�m{ө����JW�9OP��%��j�dȁ�ˊD����\�:@��K���	)G8�t�ҥ�.}�bX� RC�䚐-z, 񃬊�G����L�3߮ۦ�2H��r�}��<����	�=ᑆMe�S	�v��ɪ���4
�9J%F�MC��O5Rq�B	Gi���Ǔ6��1k���I�J�cTE�G"��k7��v��I5)����V>����D��v C�A�Rb4�k�H���8c�1�H�� ��b]ve��t�7.�c�ā����x��AW1=c��[5�K<h��T��
/�y'�;D��#V�Щ\�F�m����'jF �e��GB��A���O-�ˉ�>(" �Q�Ƅ_aA��	���LW?T����uk�O���P������D~� H�y��a�8�䚸]���'���;.��w����O�V�9��Hf^��-I)M�X����i������ux�$+��+[Y�x��G�g�nX�0a�
/�6ТoY�d|Ex��5�&��bjq��I�ٟ�y�3�)� ~� �)�#'���E�AT�����mH<1�1��u ��@�T)�Û�y�cS<+��`�#O]a��0�!�(�yB��4)�� �b�:\��kW$֮�y�C��'\�\ԡ�ce~�sQNE��y-�<?���M�EMd�pֈC��y"�6�DA�n�DV�դœ�y�e�;f��i�V�.g7� ���P��y�'X3;/�![cU�fW��B�B�<�agD�^��	$o�IQL	Y�u�<�ԀR�'<$lQ1c�-RR�I�p�<Q�Ii�p���+<@ u�7��`�<�����y��nH����0 ]s�<��F�+�����~�>����<T�P��eK�w1���HG�`o�L�� D��r焮�B\�c�6"ߎ@��;D��C�N�(Hֵ;d��1#�r�F#D��i~m}
����^=\,�e�!D�� �ӺI������$�:L�� D�L*U�1
�J��O�`<z�vN>D��!��G�z8򯃶Ail�{�f0D������7`"T)�h�=�p��p�/D�āFʟq���E�YX�#WO;D����!�"L(X�t����`0��O:D�$ˑa��~v
�Q	[��1Wi7D�@�HٳA��L�A�2&�zq�T�/D���ŀװ���@1@��0��+D���#)I}Q�Pr�D�  ��ɶo*D����˻ }�a�r�]1��)i�*D��"�� g{��$�!޼�1`A;D��JD���k-p���B*}g�4sO9D��ke�G�E�.,�c�M���B�e8D��0!@�-a�����ބG��Pwo6D�X�t��;^P�uc�`����3D������S=&e"'χ�*|]P6�.D�P���8N� $	�=�Ti�Uf"D�H
4�^#mK@\E��2x�B��e"D�J��ۺ$bRp��D*0�E0�"D��0�ϣ���Y��_����?D��dG�'6M�V 0(�%���>D��k��E��liP`d^�/��e�"k7D��2$��,�RȚek��s�j�B��3D��j���FX���gJ�L&^�A�1D��o�<(vV������P�n�C�<yGK,NT�J�G�#�4��� �}�<aE� =��� ��^�����^z�<�n�>�����⍠��*�s�<q�i�ZBV)�A�j!#^y�<ɵ�U!Zx}��U�]�����_�<i%��w<f�s��%s����]�<a�a�O�fՂCV��HE��`�<�w)	_2�5�.�\���Я^�<9���p�(8�e/؈]���!��r�<�g�/Y"t�9����d�7n�v�<t�U�%�z�� �q��@c��s�<�"OE1+$x��Ŕ+�bų�h�<)�G)��8�b�Zx>����c�<QH���=[�S�XJ�e�	�y�<4�	��<Xq��ѵp.�e��s�<	���œ�*3^ v��EV�<Y#쒅[t�e0~hTTC��Bl�<�B�F�G����V*.�����L�_�<�� H�	l(4s���֌���^�<�"��i$m#�C�(f�dA�Y�<� ��$d
;Z@ك�R4
UD��"O��!���Yf]�c,�;G�Y�"Oz�ۢ�����,֓G|�3"O�륬ۄ��e�RK��.�b"O>(����E���� �ә	���a"O��a�b�3ъ`���˽K�V�@"O.}2�ቚa�^�Z�A]nN܁"O�=�	޿{f�a@�~�8��"Oz]���Z�*	l[1(UW�ཻd"O���H� �pT`07cs�u�%"Op�c"�"3 ��2��#u��"O�<����-Dj��#Lǿ4t�k�"O�C
�~�pLJ����?� `��"O�i�Hր2�
�7+��g�8���"O�Ȳ��P1y��M��ꎞ�<���"O��BGx4`�G7w��$�"OJ���V5pX:��fJ7���a�"O��N�40��!��a�,ˡ"O�D��r�����%&{��t"Oj`x-�S�b�[��B�,]̘��"O�hU�=ok��HgN� ��,�"O��C&
MGA��K�Lk�r�xc"O��k!�۱x�i���EQL!1�"O�Y����r�H�6FO��01&"O�M3GМ���{t�F�)�*��@O8�%aB�-��Lj�`Ǉ*}JIH�f5D�Hct��'�p�֪ʦ[j*�J�L7D�p�%C�&q�( �&��Z��T��5D��� LB�i� 9�d��u �S�� ��5�Sܧ
+2pi�o�P2��3�K93��u��
�0�{��z��@B"ܷ$%^ ��H&�ha��ږ��TP�ʐ(U�֥�ȓ^�:@�����,0��`"Te���ȓpU�*��9`����/K)	�ڜ��8w$�`)V4ʚ�RAb�9 �ȓ|�V��1�կeRĄzr�����ȓL$~��A	�$����cO�W����Mr���d_2$���NʄPn2��ȓtv$vE�
y��8�ҷ��y%��E{����P�~Ix��E	��e�J%#�B��y���l�"@��N�ꬁ����y�戙hy$Y����V�YPK�y���>u,� G��(�.��g��y�(P>T�|��d`[%):(m��yb��1sRu�T	6�޸Y����y��v���F�+
��݊ ���y"H�;�6 �!�3�ީ�w/P��yB�]�!�d��H['qE��H��y2�'p!�`���� &c�����#�yb,�'3~���l�8���[P�Dk�<i�R.��|C�]�?Q�=K�mDt�<iUE3{f|ݣD��U��jq�o�<��c��o��!j� |N�{cpH<��	���a��y��W$�< !��2�PTȱ��\�*���[�!�d4�
�A� �Y�̈�"�!򤗠k�L�[��~L�
f�	�=á��Y/.�J�@����C��؅�yB�*��i@雜U�v�r�e��y��J"f(��ZCFΓ]0<T����y�,�7C�L@E
�Z� Z�D��y��q�dc�%�&M[!D ��y"�S�%<�Y�t�ڔn�}A񨂅�yr/Q�`pug�$�
B������ Hxq0�7�e���.I�F#u"OƐ� ��q2�G75ڌ�2�"O����^�o�,��IV"�f��"O I�D�5�J�N�����'"O�����I��z$� -�N�F��!�'���-{���#5NZ�XT ۅ��?�TC��?1��P��NFr8Ȣ�8H��C�ɡ4���7��{�0Ȇ���B�	�P�n��Pg�4��m[� ��q���0?1�(Y�~�:l�長{�8+3�E�<a$�:4~��я5L� t�d�f�<I��{�|,�W�Ȱ&F�y��`��m���O4�<��E���A䈷!ؼe��'���:6� L�ll8�,�p���i�'ND��W��=~��d!�&L�`4��c�'���2q�S�,x��ͣP>�M�
�'9��ro@�&4��L�K<�ۓɸ'0ܰ��T1o�����J���K�'_|%�Ҡ����I�r'�7JH�Q�'/v���H�E�<�Z���,L��	�'�j	�"*��p��ҥM_�9n,�z�'���!�.��Q�|���э1x҈�'`\�:b��}ښ ����>�P���'�>C��U)z�0�:�'@�dS�m��'���v� �+H��c�E�]��k�';���d@E�o�8�cO�ln��K�'�
1iK> @'�^#f#�c�'�xX�g(=v���C>Z���j�'��Y���G�8�nH�K�u��'s��k��.X֖͙T�Ůp5����'ct�C����3�0��AbS�h�Nuh�'���h�V�H�L�eB����'���Cb'�4=>�(�o8�B��'���X�L�a�\e��Ó�iFP@�'ab���N�7�,�
A��"x �'=6�Z门ep@�p���%j�%3�'=�ؒs���M2�R��%	�t��'#�\�W��+��!3�նI�:���'��X�Sg�X�,�Yr��A*�P�'T�Mɡ�и\Je�a!�>�Ĺ�K�|���=XH�S�#'�����D;����f�`��c_ <�p����~N��8�$D�,��	D9!~���e��)r:�k�� D�PZ�`O=;vxk�`Y�!�J�S�=D���F�0<��q�i�-ll
]��:D��Q(�c�X(�cjW�p�.�ڒ�3D�pE�F�C����!�(���2D�\S��-4��8s,S&\3�9��.D���`�Z�'����D�� �ه*+D��+�O�hT��;4	Ζ}��h��)D��J���6�`�r$i<a��%3b'D���ю���S挤Sx�iKc*O�AX%���t_@´�Z�,�=K�"O �b��(@�L8vˎ�!$"Ota!��O���#t��!ńp9"OH�$I	�O��|�7�9j��
�"O��z��O�VŃ�E��8���i�"Of���+͕sHܼ�R�0n �{�"O@���@ݦO�<\r�c��F4Z���"O��;���/Բ�����0 "��P"OZ p��I:m����6���I�Tٱ��'���$#v9��K��vǐ���D�/UTB�ɵR#�!(�A�D��q�G.u�N\ˎ�*�g?�CMJ��)���%y$ܐ`��SM�<� �\` /�CbH̐�'T!,Dx�"O�U[�&�h"���H�-s%n��w"O0yѮ��[w�Ȧ	��-�"O�H���C8E��bq�K�p:X���"OH�� '�=d�Ld��4D����"O�I`��/��c���6H�.��V"Oz4�D���#t��;|v%�"Oͺ��A��ԓw�%f���!"O��%A
�ib*ŽAlX���"O4��w��@$��[�H̠Z\|�V"O(�{Fh�0�N�kW@W��Т"O��&��9t���0 ��V;`t�"OJ��coܞ���X�o$����"Oi@���""Q i��nCV�#"O�@��aIg��M.�$3A"ORh�툎a�*\QaK�^(ʑB�"O�t�!��:2j�m�&�7l�Jѹg"Ob��'�
�=> ��o�D���2�"O����O�D��hI��ܨ0I�B"O`�Cbk���%�g�E&VՒ�"O�� Vω�zh-PQ�݅ b�A�"O���E%@g\��B��I�hm�"OB������UJ֊J�l��"O(�I�z{��J
�4�2!�0"OJỲ��;;
mQ��Y2d��x"O �f��<�D]��Nz�f�0!"O�uI�[�:$@�!�)ψ.�L�i6"OE�����&��P��1W�t
#"O��S-K�/�)9�%;�"�ۡ"O�ً�Ο�R���5� �M0BD�"O���ڞA_��)P�\�.��)�"O^�b���~
��c��Êj0��G"O"35Ā:,��ꌐ?�}��"O�݈�E�7y�@ I�
 �y[�H�"O��E,C+Z���#I�M�Xi�"O�����(&A��xBry�R"OL��U�W۲������(�����"O���w�#X�8��$�X��u"O*љ���O��ЋԺ�,��$"O�#Q&��NUc���i��K "O�i+����4��JS�̱�BU"�"O��`��%*�����@�B�x<�"O���� (�(����[�i�0%�"ObL��IQ�J�I�g��4n^� "O�Q#,�%GtaB��=�b �"O.�Ae�Ib�^m��D�~�cb"O��$�T����V�G�wނq�"O�����7H"�RSU'O%ZX:A"O�Ld�S&h�	�t��y{<��"O��2�]���	R��
3x���"O$���Ɂ�;%�Ac�ZBb����"Oޙ�M>y
� ���:��G"OHi�&!C�}N�]P��J�;�`X��"Ohu�A펕mT��C䆹Q,�\��"O� [�\X-���3���&�S�"Op�ꇎ�mƈ4zqg�1/�43W"O�q�C��D�>�K2�B*7�.��"OtԠ�΄!,D��[7�"O�ݱ���"�-K��^�2�J�j�"O@�:�f͌�@���5}i`0�"O�P���ϲu1��o�6X2x��"O `#�$�����[�D��(Ir!P�"O0Z�،ـ ��	�p0�b"O��A�{G���E6%'�I��"O� `�Hq��Z:)с\;���"O�ڎ[i���� �4)#��0T"O����^�
4���iuN��"O��vbـD�Ă�Ζ�Un\�@"O�l¥hG|vV+�nT�LŮl%"OpB���ԺI� �O�p�R�"O�M����|�=��Ĕ��`��"O�*5�Ɗ8r�e�ήu�fI �"O�iP��<d}���d��43�"O��S!Y�ܡ��,ީ�r�*@"On���\�L4�`�l�/9�ָ5"O��!�o��+����}"l|J�"O�
b��x��}9&k��"���"O�*׉j3��"i�6漃�"O�H�a��E�|1Ag���#�"Oz	�kTo{�
�&��(����*O��s�DJ
F�@���:` 	�'������!��dI�	��h"���'�����M�F�~�8t�^7�X�
�'V�k��9H̹�f�3Y�"��
�'n��ə=�"� J�M�F]
�'`R����i{�a@�/�|����	�'�l�y�H�:�-4z�i�
�'n��2t�-a�HuG���x�H��
�'�89wh��X
��Pf��3q�|�	�' ��W�}�D�B	��[�l�Z
�'��4r�_{�Fm!�N
&x��	�'Ҏ�Iu���^30�Rq �1 ��d@�'\-� ��)څx����NuP<H�'�$PiӉ�?7����$bR2Gr�,�
�'��T���_�'�( �c�K�M�*<�	�'���Qw��9����	Iv)�'�X���X� @���P�k
�'�B�Q�M؇s��]����N���	�'� ظPk��u4J��A�� `���'d��#C�s�����NEP�r�'��P�鈏{������I1��'���cu���s4�ZQk���6U+�'������� EZ&�#���
�'�aSA&�y"�:V� >���'� � 4T�\�Nݘ!�y��I*u��<���Z[y��H)�y�I�/rBޝ��	C�O�4�!�+@7�y����lyys��xX����@��y��q�",�CݻZu��K��y�o]�[IT�T#\	~��Ie�R��yrJ�*R�ʌ���H���q���yb�Q��v����ݑ~��@Á�
�yB�2(��
�$�=`7�X�a����y�
��4��QT��E:��z���6�y� �o��i �ȳ;��"C���y��Z�]��p���+_�������y2��uR0Y`�bU>
���$J��Py"�]��ܑ����)6���x���X�<�f$��3����B$PK`�H��HW�<���6]��ձuOT�~��,�l�R�<���*U��Ic�ᑗFߪ�0�)H�<i5�^:y�*u��f@���|� M^h�<�B�O6 i�r�ND;fl�i�l�\�<`A�V�`��.X/F{����GTY�<�+B�r�%�fݴ@Q���X�<I ��]�2u�0a��{�Ah�̒~�<�p��=��\JG���\2��[�.�t�<�QC�~1\paю0
�m����s�<� \���L�$m��3�߄O��8t"O��(ӳ���v��?�Z�"O.ố�!/ܜ�v�ԝRG�=!W"O��B�(��{c��(h)��g"Op8��5�
��̚�04rACu"O:�Sjy	�\��@~5�uH�"O��1�!�D��0��o��y2�Q�E"Ol��*N0(�r�@M��"z�(�g"OP�5O������G�Cb�9�v"OFA`�OZ�*�� r)0cAtQ�P"OR�BA�?B��"��*ŮY(�"Ozm����jH.\RgN�q���"ON�qA7h*�jS ���P�S"O|��7bD:R-�����(��qD"O�a(BK���2g�F8	.TJ�"O����	PQ6���e@2�� �"O^e�"Ƒ�!�2�G$]�n���"O*9A���Tu�IsF�J�\�݈�"OT)A���s��Ԙ"P�p
�,�""ODTq���6z!�r��.[���#"O6�آ�H�5>M�q/I5��h"O(̩f�
�s�x6L��.��&"O���œ>uQ^����p��5�"O0 � ���xŘ�<��[#"O��ȅ�W�9�@�҉��7���h�"O�xˢ���j{0�9I��P ��;�'���p�%�%d�A��Fε|Kh(�'��-	+�0a�|��6��+)$D�x	�'d蝨3�غY��!7g;)�:�@	�'�l�`����'N]���D��'ڄP�G�ˍ��	z'I1�mp�'�R�0��C'\LI��!p~���'$�UB��V�%�lQ�I�:fz���'�~�k�J�T�j5yaI	]��;
�'�$D�A�ɒX� ��W�zeP	�'_�=;T��!�|����Z T�(I	�'Yz� @��9�v�,����'���P1e�[�ݱ�hנ"����'��V[\$� u�.�k�'L�Pԁϧ=�% ��f��3�'E�D�Iެ�:̱��g�@�c�'6
x6��-f��IU�ѥX�`q�'���I	3����k��Y@�}��'6�X�����R�k A	�R�2��'��Mʂ�����5��$��)p	�'O $c�ğ�[2n�Q��I��p��'��3��I�u�jG�� HM�mI�'B��u�B��DJ���i�|h��'��MY4���$d�H�(��e��!��'���3e+y?�����2K:AZ�':�]�P���r&N1{�nۥ5M�J�'�U;��n�����͛&�ޠ:�'��� @���C"��;	�'�h����L�y�E�&H�
8�Y�'v�}�6�	�}'2�0F��d�ҵ��'i��!!�ˉVR�eC��R%Lt���'�,|�da�z�hxG��M߶9Y�'NU;��#4d��8Wj[/tK2�'>\pI6F�k������	p�4 �'�8�Z�l�qb� �(ҖURH��'��= ��
e���&�������'e\�
Q'$ ��ᝧ�h���'P�0���W�l����Iԩ y��#�'i�a��D���-P	�{���S��� ��8�m��?Ϛ��H��d���"O���gHyX|���T� �"O\�pD��)�%�f�q��M�U"O@��ZސTzr늏���"O���aߐ��|����
o��Q�"Ovx��C\�rH ��W��-}�Y"OJ%����m�hT��뛘d�  T"Ol�@ -Q�081�I�8���!q"O��9��;�Z�����640�e"Oֈ@�@�^�¤r�C�6��!"O�
u���a�����
&�lИ"O^�y���9�@�'%����"OF�#�`���݂��H�h}Q�"O��k���:��g�]�`��b"O�D��#_�H��\�����_�V�z�"O�4*
/� Qe�1@`�2s"O@!��g/#X	�N�2�0{�"O0�+� �X�FA�����\��a"O����cW*>{�e	 *߇"�|9S�"O<��6M�,bϮ� �D�p�:��"OT\{��=/�,�sl�"9x��R�"O����Ťw\��2à'h�J@��"O��PD���;L�S�_)gK� 0#"OƀA� E" 0����#��Y-�9��"O4�I��@�zZ���^�աC"Ob�Gᓲ;���� d�ޭ�q"O��ƞ⾜������"O�q�-X�+�0H�'i�&.��l�"O��`eK�w�*�+��Ǫ0Bq(�"O.u����DF,�ЅΥ8&��9&"O޸CS�E�&f�A��[*׃B�<����X �XRG�fdT��q�E�<9���aj>\D>A	N)�#�}�<���4m(�`� 	8.A�DЖC}�<)d���O��1c �\�pnڨ����q�<9�j�:*�i�+�m��E�iVS�<)¦�k��i�˜���L[�YJ�<!3����<a�,]#BNɲe@�<��D#0�$�#	:ySP���a�y�<�1WOF��R-!'@��Q��^�<��*̽P�q@��+kT:A��b�F�<awkZ8�-h6�/�^]�l�i�<y"A��O�|%qu#��@OPi�<�G᎜�=RQ�ȊgtDcE�Xg�<YP:	la��μ\->�fe `�<���ڿ=��I'ݰn�&= ��B�<)"���B`B��K�1� ����f�<9�៭k{�U���	H�؛�hi�<) ��#F`t��i���Z)�!�$�e����
�".��C�L�#�!�$1\q�p �d�#�5{Q.5v�!��Љ|�#�ы^H��vKd !��H��၅���x�%�r�!��3��M�2`=�0���!��Z�`�J��F�D%��+�f�M	!�d�4~�T�Gn��n�b�$�/�!�M�u$��A��+��	���
�!�d�$�*�"��,"�p25a5p�!򤓗c����H�3rhx �	;7�!��&q2P��k�h��2�>h�!򤆊8�~�8V�h~����J%b�!�D��a|����X.p�����M�!�䐴[�6iӱG�_�����C�!�d��e������ɻ(� �5d�oz!�� *�s'�I���r�;G;%"OT��0N��4��)�kP�,#��B"O�a`�N�E��9�s��
h��%�w"Oz��CM��ZG�5i�D��q"OheS�a�h�;��ѝO����3"O&��vL]�S���]���	�'�Lt�Ucɫ�͠�⃶�$�
�'0}X�l_'�<A� KI=39�A[�'��IƪW�yh�:�.ڲ-"�'k�H�3NS�3j�Ip��',>l�'X��٠��As�xZ���/%�:I)�'���G�>(�pK�O�T���'Wxdf�@�ÆJ�
v��'��5���"/��h��X���x��'w�͂���&*y�|A�BN���x�'�
i�8cƤ�4$�x�X�#�'S�|+$B۷e~�@C#Dv�"���' ҝ�n�$0ļ���
VbWf���'Z����*B�6iF)a���^t\�z�'G81r��;F�z8���'�x9��'�>� �(C�V���Q���3�a��'����5��L�FaZ�-����
�'�V�Xc�m�l��g����
�'� �b�5DG�O��ʴ��'�Qaw�:�0�R6-Y�B�ص{�'C�Ic���N(D�RT��5K�he�
�'猹b"M�Z�mZ�a�Ffjx��'��X���|��xbA�%;��q��'a>l3#,��t6j������8�|��'�&b%��$0N ��J>G'p
�'�us Lʌ3�t�2 [�,����	�'�ZpHS��H�Dp'��/�,�

�'������[�(�+��� �Nt	�'�f	y&�O>mi�	R!O�-�0�	�'U^�X�8��$֦�#�A	�'Ƙsc�	�v_r��e/y^<y�'��dK�cц�ps�m�4j	�'b�-mD�Iv���sd�%R��2	�'E��[w��)��ᗍчl\���'�$]�Ώ,4�6�aP���٩�'^� :�IP�R�\H�V/J�o���`�' �K@��'���q�^{�P�9
�'�6pr��'����9l�%�	�',4 )3!C�*�8WM�1uK�1��'�P�8�f�6+��$�3kŞfTH��'y&HZb#�]80��i*coL�i�'�.���ŕy+h�0���.Vj��'� �9E���vԑ�"h,�>�:�'P�}�"�Q3������x��!
�'����)Rn��1�IQ�> p�'�8��j@'VYM�%�/	�r���'��QxW�\�4��aq�̞o�hy�'x�x��lU�p�r%���E�/�#�'&�(��5۬h�%F�)m��T��'"�l�� �=�J P\�$!�'���U�I���5#'���
�'�2�{�MCb�e Ux]+	�'
�s�	�6r�2�4� �⥋�'���C�R="�^%���U^�	�'L���J/s�nY�#dD����'�>X�s��j:`�#�&/(�� �
�'��A�(Θi�4I��_ L,H���'�lXxV�N�_~��+�QI���	�'�rp�$IH`�����!B�TM�	��� �x���[@Ru���0�N�`�"Ov�Ң� �q���C/�>����"OZ��#Jw�� �(�/�X郓"On�×'ʪz�V�b��LmPAp&"OV%z�M��:�T��P+����"ON:C~I a䉛)-���"O�吅$�;]APؘ�'�����"OL�cbC�g.��K���'P����"O�0�n�}ԞЉ�m�c��|�"Or��S����$���M�<��9�v"O��(�[�|Pɢ��u��!8�"O�P���G
�,��*�<��@"O���5�V�(���jU{���3�"O<��"ȉ_��D�f A j6���"O��p֪?9�}0U��<,c���g"O���C퉩�,R�LN5f܍�5"O�d�&�ΗG^h�FKByv���"O8�1$�xu����t�7"O0�k��V�lPd((/q�hcU"O���آ ">A���>���� "O>���$ؕ��YfgÞY�*5s"O�4��K�:�c�"q-�Pi�"O"�6�Qrv�b�g�(s�Ҕ"O���faR1��(1AY�!�6�8g"O�Y3Dk٤4jl<"��)R�t� "O���S�C8�4�1$NyL58�"O�Q�R�ٯ�S��v�<K�"O��)'���4�	��9L�th��"O�]�!�Ej��EH�|}��"OfѤӭ��q`��wPh0�"O����T:�|���m^�Si.m�S"O4�E��x����̋�_J�0"OX�RU��(C�jg+�;G��4"O����Nå!����f��t.�j5"O&X�O��eM>	PqC�=jT�%"OpU�c��;�����>%2j�"OD ��E2ZU`C"܋ �a��"O�<Hӭ�$t |�[ ���ȸ�"OB�Q@(O��0�H��O5�QA�"O�����G�{�]@�K�!0e"O�t#A��}�Vh��h�%$�*��"Ob[ ��?"� ��%*F!*C�M۴"O�9	tc�\&-yg��6Ӯ@r�"O��	�eݸG�0�c�H%c�8�"O�X�\��� Pa��+�>Y�R"O>]��*�:ԩ���G�4����q"O�FжJ"�	7����"O�h�"KH(�<����r�&q�7"O�$:a�4�H���@+`��Ac"O(ɩ�U��ݳ�
�?��Ԣ'"O`�j��NvL8�bI.�L���"O���c����Ua�� �����"OB��ć�vN�A�R8x� ��"O0DR�ҤM-X<�3�	�/$�{w"O0�@�摴8׬�� �]�,��d"O�:Q��N
Q*�_�yjv"O4�*�H�)0����:_��L�"O�9B6�;B@5��rV��4"OĜضIU }�2�3�pm�%�"OJ��D�
bP�)�K޼5S�U�b"OvŻV��8�
�	�݆q2j�SB"Od����ʤA..�*G�`%�()�"OzA(B���0̲К$@[�(vpR�"Or|��b��B0��*q�Om���"O� \�C��k���:cQ�7iD9��"O��A�E�
�)�o�l���"OPQY��ǵQvμ�c$��b���"O`!��uI4��6�.H�:�"O�h����Z7��w�ņ~��̈"O�0#"��G�n��W�-\�h�"O\d����!{>nQ`İ�"�(+�!�Mm�r��� x�^�����M�!�C�rʼX2�
2?Դ@��"r!�ċ@܄�p5oI$g5T2�%��Q�!�$�JZh�㶧[.(}P#��3�!����\:��S�ŚH����7.�!�$_$dj�Y�OW)i@����\��!�$OW�x|9eb}��i��3�!��!��h���D^�Kp�
%�!�Ď���d�U�܄fMyҥ�!�D2*p�aH�@?W84y��ݪV&!�d�4���Pb�q:�!��ٱi{!��dNX}�Eb�(IRPcw��
!򤕫j�KVE��a
2,���&!�$;Ԝr�k��T�Q��Z0Q�!�\�25���Jha����P�!�P�*~-Bv�O�}S�\ QK��w`!��X�Rq�N�`2PY��Q�9!�$/NPl��W�K�^��03c]�wu!�DǷ/���d,�O�"����/m!�$�e��u!3I��K�rL:e�T�d!򤂎#�QCׂC#�Vѩ� �`!�d�+h;�B$�Ԣ����v`�@�!�Y9*A�Ң��=�^A��)�!�[$3�n�JG&%&��,�a̅3�!��Wd�(�%��\��m��T�[�!�$ѽO��=���٣a�@ēb+̋B�!�B4#_:���/0�����K�{p!��@���� w�+�5F���jc!�Z���m�8��A�o�!��'Z����ŝ(H���%�K1g�!��r��iZ&�[=Y�~���
;�!�D��.:�p� �ՌL3�KU�@�!�]"�0��[�R�f<��L��C�!�$Cy@�drD�N�H����,��>z!�&lg�b�@��r��P��j�$ie!���9n���1�ď^��i�Dɑ�o�!�DA.*��0ϔ`P(��55�!�=�}�+�u4����1�!���-f�6lq��	�\-J=���Ɂ$B!�d"��i��H��NF��cf�*2�!��.����,
 .Y�Ñ�M�+�!��]�&�`E�RuK���C�B=�!�'
�t�ĤaG$�����!��܉_�ޑP�-^2߈����T�u}!�d̼rڰ�h�Viـ�Q'Ȫ_W!�d�?5 "!��ˈB��@���ch!�$��J�h�`@��[�R1����/@4!�'��}"�	z����2��^�<�cF-�B	���l�����X\�<�ԭZ�=`1�/�8Fln!��U�<�D�f4𥳥�7_9��/�S�<�˂H�J�pG�����D�P�<�'XL�����PK|�RV�R�<��3[�qz�&]�E꓎�F�<�r��;/hIȦD D�pY�qnC�<飧�9B��"+�#�����N]v�<1�,O�jXp�̉-D�=5a�n�<� Dc3L�b���Sv��!�E"O.���I�+��[ԭ��"��"Oqct��$.fH�Xc�ۡ�xE�"OR�[�d��j���sĥ�
F���%"O���A��	4�4�dS�,��y��"O�4�f���@Aμ!ЩZ&!~ڸ�b"O	za�2$�r��Ǎ
���C�"ORqJS��(���T��c���""O��a��s�R���/8��-��"O(i9�fӯ	4(�0E$�$ �N�A�"O�d�Ң�1b�r8���6,���"O��&���fo:�s
��P�4��T"O����gIO:^�z����a����"O �C�_�Oy���$�[�*8`H
 "O��c�j�ł6	^0/3���"O֤ F�(&װH���m-p �"O����eP�K	��ӄ^�z��D�B"O���wC��tMXyid��Bf��[R"O�J��K��$��E�lc�dqW"O�Q�f��KZhh���0c�iPc"OX�cWgܩ<�{e�F}����`"O2��2JQ�	�
D�PH,C�r���"OE�O�N�0�*P�T��̻"Oޔ����!�fR(9	�a*�����y��Oexȇ��-4�N��O���yb̯g��-� U��A)"�R;�y"�4�l�7*T6�~`)����y�CA�D�c��(���տ�yB�X���X���"K������y��K��iX�́Dz�X�AK��yB@ �v%yV	 �:2Ir�";�y�lͬ_Ϭ9#AŁ�0v�,{p�@��y���=���넭!>�F��L��yB���u�����AP
4-t4��,φ�y2N�7u;n-q�c��+.��!�F���yB�D�K˰Mڃ@�*%`�qcH��y�c�-()�b�9�2�A��y��O�V��X�A��	��22l�<�y҆@�<P�bH �A���ξ�y�ȑ�Q�L�KQh�3�ҹQN3�y��ڙ%&Q�q�Z�)`@�&튤�y���1��eGͭ�5I��
�y��Y�H+����P�.�8تgk���y�i�',.j��V��R>Ap���y� �D�E�D(*�0�	@��y��X9��I5/��?�@�C��:�y���g�����
�L��H���Py���v�9����*� ��I�<I���KA���7�/P���A��<�B�
A0��J�|Dk���~�<Q5�ۧ>� �X6ˎ�]���&�Sz�<���K�jZ��iƌ��%�EHx�<Y��1eZъ��ސ|Oؼ�0�q�<������(`���N!���T�<�닔~v����I)�Pq�j�<�$-W9#�P`�A
G���ҋPc�<9q&�:Jd�cQ�_pC(D����b�<�d�M`�8� +A��*��'�^�<q��h?�Hc.��IW���3FR�<�w�Fi��mq6�[�*�:ّ6�z�<y�^�Y�-(2� �qDg�w�<�'Ԋs$6�r3D[�:�ʤ�e��w�<�敞TXJe�g퀵c�.@I�<a#��~B%P@�5�0��\]�<� ��A��$��Ԫ���'�����"OF�� 훍b�z�����C9�y�p"O�<�Î�2c�L��C��M
<8V"O�$��mӋF5�P t$Q ['JE�"Ol�aD&ʵjL)㣢t��1c"O���b�8Dr�HB�kʹS�"i�F"O :�@��&�x�U�L{̤s�"Oޘ��*�vA��Dп
0��4"O�1�`�M�jq�	0�<��"OH ����V]	�@,W�H��"Oި���T�q�R-"@&C><�
y��"ON��@܇ �p�dEY�"��9K�"O�M����/�H�X���{t�Rq"O��ʂ��-l�|�0Š�$,�Fp*�"OLM3'� ��8�/�<~�բF"O�����5m$n�2D�jrPQ�"O��1�G0e�`�D�1>S�T9�"OPe���Z<E�Y����!L|�b3"O�IUR�!�K�+@0�-�"OF�*v��8O7��;@�A�yOx��"O�;$EZN	<�㓫�=v�P�"O��T'�H���[aʘ'>�Ij'"Op��!���q�@#�3h� �"O��b"#7y��!���3,<�"O�(�LD@�2d̒�f�q+�"O�#Gӯ
N�u&��l�t8ذ"O8Z��Y�6A�;���f
yd"OvP��ńr�pE:2h�+Z�&("O�QJ��Ov�$����T;$�Z<٣"O��kW�,C0��7'HW�8;!"Op�EG�=�nA���Ԅn'P��"O���6�3
���ط��}����"O�(Q@aU:-i(�Qֶ5�:�%"O��b[7h��"�Ɖv`��(@"Oшs���ز���PQ���"O,Yy�ㄔ��ܢl�5-�x"O��c�nC=�$��s,٣1B��)A"O���C�We�0��*��W)n��"OL���� 1(Ȥ�A% Y�pj LJ�"O�œE!!$Nё6�QaG���E"Oh�"e�G4	?z���M~]�"O�-XԊ	�)�D���W�1ʰ"ORE�V�خG]���!K�����V"O�Ÿ�bѐH� 	 *��o���S�"O
a� ǦU�$���Pd��#"OFm;gi��)�%��Ѩ]�ĵ
""O�@'���D������"�"Od��5�d�P��.�`���"Oz�y�i��SQ���R_*`)�Y��"O�}9�\�j��#��}x�Z"O��4�̆�~��)ԔY���"O�Qم!�
�� (�<�2,�"O�I!n��:��89ņ
�v��"O^��eр8P&m���3C
���"O�y2E�I1E�KP�ע6<(S"O�U�Ү�Gh���E� G2�8��"Oʵ#��Gn���/R�f)\Y3"O�r7mI�;W$xH�'N�|��Cb"O�Y	A �s�e�C��	���3S"O���7�}|�y����̑y�"O�9�r�%7qR� �DÎ��@�v"O����8XY
��%��U�}�"O���`�˂*bؕKԤY2H(�;�"O�@ۑg
�= P\�I_�Z#�\�"O� ��B7*�,@z�������4y1"OȚf�B1!Ǹ�����a �e�"O�{%˒"�M��sW�[6"O$4��F���ɰ��_�`9�V"O�ؤB��N�\����@�o D�+s"OXqZ�,~�:�ja,E�d�YP"O�\���T���GaS,0l��Y�"O�� BH�;>e%!A,$�!��"OpY[��r:����Ņ<wr�i�"O4�C�++c�� ��-�u�$��"O�$@��O>h�>��"LTxs�"O<�&�	��K+�*b$@"OЙ!DE��q��e�s�=r\(#R"OL0�S�N2md�s,ai~�`"O2�!t��5)��R���yW��KD"Op�Ԡ�M��`�M�F�a�"O��)��}���F܌HR2���yRLS #j� r��G�@�J������y�͎���yz©�� P� �Ѡ�y"#
�0�.}�t�#�r�
����y��Z? ��Ui�d�$1w��d�D��yB���(�pM�cg�/p&�*��X��y�_,4Q�HG����#(!�y�?6||ztW���h�c�%�yB�Zz�&�A@R�o!,�Ї ��y��T7N��ܸ%�>S:f�;��P��yC7f\�h�ˉ� j00�eH��y��U�3�P�RDf��!���y�>Z[R��7�Z�I�l�@���yr�I'y
:|!A\�I,�shE�y"@�4!|�D0���Fl)��]�y��ҕrN�	t T9M�Dz.�:�yB�ۼd\� �c%��
�mpKқ�yB�,P����˗Y���%*���yb��(9�&(����K^�h�uo��yB��$�� �r JT&R�!D�G��yR�P)n�b��R���F��yb�B-��`CƴAczp�&��y��I:+�`2�%[�H�� ��
��yr @�6���k(LC�ԡf�J�y�ĲF��$y�#�����z�� ^�<�v�@�. �a��uB"�P�<��ՙETd����!�)��)P�<1 ��F�	�@�8�����K�<�7l�:{|$y*AK�HY�u��E�<���.y���IV,�C��J �}�<Q��,y8��!ߣL^��*f D�<U!ɽB��aC�ҚNST�B���[�<�gƘ�O]/,lh��R�~�$�ȓ&���c�L�&5�Lq����꜅��|��H`�Ĺ�t����[3W�(X�ȓ�2�j� �D1� �A,o%��VDJRg�&���`�#ߥ/�湄ȓC6lܪ�푸(_8���B#up@e��&\���q �5�� �AJ��ln����k�L\�VFW9FZ�U�6���n�耆ȓO�
�*�m(�L ����*�<��ȓ;{R-:�M�]4�0��H�,��ȓQ`x����|޼����g]ȑ�ȓL
�2�+ͷ /P����O)#�I�ȓ5�V���(2�Ρ0'$^C]H\��,H�1��B��vܙ���-K ��ȓ.ȩ�b�X�H1p�J֖/Y�9��Ig4q���T�nLR�K�B۔9�� ��S�? ���'`�4Ri&���A��Bf"O��S��ք	��1�n��(�"O�i�nI$	a�d{�A M�"902"O��(��L3c�X�a�N�VL�Xh�"O^<	��N�Y �%:�L��Y<P�A�"O�t1��Nت|����,c'�x�7"O�-���D�d�Ҥ���m���;�"O����W&_���0K[�o���1G"O�,zL^�J�F93P�)7Bi�"O�h�'d�1|�TR7	�T�� E"O�q2� �J�y�hG�v���@"O�ِ��;H���K���\�F��"O����e߯pne�d�O�z��L�"O�\"g
�Br242E�w��5z!�ݿCI:���+
m7��Zc�ŝ
�!�$����B�4N� q{�c�!�D�V!U�o�4 w4�{�"G&}
!�-2����w�ә]dq� đ�V�!�$Z"!T�Sg�gJ����m��C#!��#ӠՊQ�_$� rLX�\0!�$&
x �x��AF`<҂J�bA!�dJ�j@�8� �HtL�=���Dv�!�DԳ &\͠7hH�q74��C�Sg�!�Ā��(� ��X'4#�q��$(�!��K�����M�'D��1�VƆ�E�!�Ā�l ��Z�J۝9�\��3!�D/&��҂��2,���	�c�oW!��R	! ���Ռޥ@�1WLW�-F!�d��_����J�O��*P2VB!�d�61|����3��R2#�Q>!�DZ���@ U�+������^�!�D�46Dt��B9��yk�� �!�䇥K���G-0	�tI㫊�P�!��tD��-i�<�c�Om2!�w´㤎N��*�*v!�d
�;r�<i��G���3��T9d!���?�Խ�bj̄��ۢM�(p,!�ɺo"@� �	���0AC#P0`!���:O|,�����5U��9�Vh�\�!�~�sD��?���uA[�5�!�d 3�^���08��/���!��L#-��%:2�R;	(>)�l9:�!�D߃z�J���bK)Lj��sd���!�D�"��� t", �\ɳc�mP!�d~H��AI�<��p�)��J!�D�9i�wEٔ����2a/!�$�
h��I	���Q�04��֢C�!�Ē1*�*0k A�!�d�$g�<l%!���%8� H
f$�+�!�BH�!�dKm�`�+��7`��%2���[�!�	���W��"U�$q
1GD 	�!�D'C�u�#.w�����}�!�dQ��8�AO�z�6�)w�&5�!���lD2�ç��ab�0Af!�$�ޥ���3�J�o�3ޞ�Y�'�&!�,�:��"!2�p�
�'x$1�ᮕ>>#d�PFW�D� p;
�'G�2��Ų��y@nԱg��[�'B����ǲM����7G�h���x�'�V(�eK��l'6aӦfV�NbhA��'y�����-Z(�P��Ţ=m�Q��'��{P瑮y'jQ��鏸2�Z�x�'��a��Ǟ�K���f�+2��(1�'/dM
�P�a����/��R
��� �5�/�$�,�s��Y	ZZ�Y��"O�0x�'
;?T� ���4�L�5"OtA����QumӏK��F"OD���ȭV��bl��O`PA��"O�	3� ղ��釛mo8�"O�Lb�g�:X��A1
�643T��F"O�⑫F�J���ah�/�젒"O�!��&
xJ��@�{%�D("O�˔�<���PsF��
�:7"O�,�&�,h�A��
�ͺp�b"O<u�'�5��1P���r��4��"OT�%�8Kl)�ÁW� ��8�d"O ,a]"$���A���j7"O��ȡи�`���(���c"O�)4F�0D�����)Q�L��A"O�Dy1.]40�~�)A+ �R���"O����΍!k�ػ`�� d� "O�p!d� $��P�\�;Y���""O`a�SJ��Tc��bHFY�"O�Ijp��lh���T>V��%��"Oh�^	�4R2�Ë ހ 	S�<y6�Ae8� 9��x�h����y�<)���k�t�� �مPM�lҠv�<�B@�6���&�RY�Z���@Z�<9V�-1SFIa�&��{-��QcE�X�<�S�6���g��U��}q��T�<i���7M�61��A�� ���BM�<��D4�x`��1���Pg�<��`�i���_�`�/I@�<���t<`�� ��E�r�����y�<	1�17����B�傄�s�<�4B\��>��x�̝��P��pC�;1�VɁ&N�����kK1�JC䉹G<�
�昏'�@{��˯M�C�	�[��\#�Pj��C�l��v[�B�	#F<,���@(S�����G\ �B�I
>�)EeW.=�`��ˇ��B�I���A����I��t��L��C䉂~#<�J�a��I���f����C�I!d&Phc�2�p;�ܿP��C�	�Q#8���e�\V��Hr�=f�C�	23% I� �:G�����X��C�I�v����f�4^�	07��j.�C��#�0����JcN� �B�$�B�	�ke�� F&�lv)����v��B��6m+�\�Ƈ^�,y: �q)dC�	�E�!���ѱA����Z9>��C�I0^��3���:���C���"s|C�	$](и"'Y�5.X�a��O,[P C�.�\m0�#� ?t�BuIےZ�(B䉨)�H4�s��
F$a8燕)1&B�I�8]�� �̌��8*Q�֑N�\C䉺B���)���l༰��Q.3u`B䉰Jk��3�A�(W;r��d9?�B�I7jd�[��Ȟe@Q���m��B�	�de�\C�h ��dŘA��Q��B䉴Pޔ�#gė�0A�����(hzB�I�HdV@af)��4�,�9��ڷo>>B�IZ>�1�I�eU]���X.�jB�I&�48rP��z��<��׭<ȊB�	�-�4x�4��X���r2��a�tB䉬*�IH�K@�Q�℩�R�'VXB�ɰ�6�ӗ"�7��dK�N5!�DB�I�q&�`�"FT�?v��Y��D3(�ZB�)� Э[�j* ����(�dA�T"O�ш�b0�q�Уԑ5��i[�"OƘ��ΌA�j@R	�٠а"O�<q6,�����R�H�E����"O��h"�+;��1��
!�l��t"O����ۜ$����4c���3`"ON�`A]�[W0�!X_������b�<	�O�*F�8@a�5��ڳ'�f�<%œ�{	�UA���=^�Ų��\n�<I4EJ�}�9ѣOA���j§Ph�<Qt��vf����ō~��M��d�<��O\*4_h�Yr/���<aĘX�<��,�< ���ȼ��&F�P�<1FOW=|��Ԩ�'��/�Z��)�K�<Q�)�-�����V-�N�z1�O�<	��[_��U�%�M�Ȉ%�J�<A��;=WD!�unZ'�B�d�^l�<yC�@�NLr��!���pĉ�i�<��Cyʎ�Q�� @���8kJ`�<�Հ��l��,�l q�������R�<!V�;|Ɔ��C�tU�y�U�R�<��Ⱥ!�h�`��W3+���2��s�<���b��!���zxB����p�<��IR���N�<+N�K	�R�<�G��SP���$H�u#��S�!Ht�<�2O����F��
~n^)�f�q�<I@�]e�Q"FZ��U�Aj�d�<����,.�V��%We4�ҁ3D� ��
0~��Q����ö�-D�l�௔s I��)Y+4CF}c�6D��j�@
<�H�r�� ��S�C5D�PQ6���^m�C�oV-v���Z��5D��9ANG�X|�+���� O�X��,3D�T�������B	ݮDKWd2D��
׋�`mR���8��ʖC/D��YDъF�d@y��K�`9�1��d,D�d�h�";L(`�%�O�r18�>D��s��L�(`@T��˔z�&�2�!D������`�:̀ࣔ�W���5#D�tiw,��RS�!�n�&#���K D����ǉ1������Qi��B 0D��¤��@;Xʇ�O�9s���#D�D�I҄"�ʥ�uQ�f����H!D�  ?�vU����p��,a�(!D��wgԜ��; A[�I�F}�I3T�D�0*C�Y(��.$'6z�"O��R��"�����
F
M:"O�\�gKT�i��?U#�|!"O`HtfƏU(���0��%<.x���';챙f�J
$jp�fL��@�h�'PJ��WB1Ld�e�J$ ����'!�Z����hp�1+�{^���'��(S`i��
S�`��m���*	�'�`�{�#� ��A��N�k!����'R��BbAA0\(���e9(}��'� 3�Y'!
��V��
\��ē�'�9SPE�:����H�6$/(e��'�05'��k.Ԓ�o�_ބ��'i\�8��)pB�n%��A��'[dg�T�� ��'!��`�'�P*��R���4�`��6z�9�
�']\x� �B�՚P1ao�YzV�{
�'F���cb^�Vc�+�O�O
8�	�'
�K%o�828L�WeF�v����	��� [4� $�5�s��1"�c�"Or���ə"X��e�c-S75�d�1�"O�����y������c�p��"OF�K�d�4��ɘ�D�V�h��G"O�CI ,�4r�Cնd}��r1"Ot�)���MJG�Q:0n���"O�a[��9oR�;1a�3O��S"O�Pp���	ĄX����WG�DB%"OƩ;�b������=%�
�z&"O� 0���x~��	��=_�:�2"O��s���j2r�bA$)|
A��"O��Cc'�BeT�!3LɾI	؜y�"OHH2&�~���sWKO2�����"OlX��F�
�HH�QJN�v�by��"OF����/!x��g���&ЩA"O�r��4B�:�F	|l�ͳ1"Ol�����qV��Vlm��"O�4[�A��^�lȨ�Î�"jn��"O葂�R�&7ؼ!���N,�sU"O��ʑ�l���	���2L��=G"O�#�E�p , {�U�^zR�˶"OHy��l�8Ƈ�`C�<�Q"O�@�%R�[�hU��G6�q"O������=V� Ug��)[���"O<)SPb�gtm�2g�X��g"O
7�;J��KGWr�H��%"Oh�Y���>/���Bv�@�K�~Tx@"O���A�!L�qU䑊{����"O�M2e'�<�R=��e��� 3%��|���	�C�x�d �8[<;u
)���)�O ����6	���:feG4@�6�Qp"O���P �&fA��Ë�x{�O^��HMo~�  &�tܒL0�'*Z!�D՛<֎1Z���#=ZȲ����/�@��ȓa�� ���V&��8�G�!�~���7 t*1�H�w�r�$� G-�l�ȓ�4��e�T1�hYWO��<,�8��~�AN�R��a�SjԉRSh���	�Gz�	�bײ���+G̜�A�  }��B�ɚGg��A���.�H6�%,P�B��-��c�j,�Vl��@��lP	�'P"��!KØ=� L�b�9#�'R�qRDE,f�y��K�Y���
�'���j�Κ�g^L����S{�u��'����W3H�#2o�P����'������2
�*�@<JLP�'���;m>��÷FUv���O˓�~��ƟLF�4`���[@(^Ě�S����yb���
F�`�q�ǷO�9�S!���'M�'7>9�B*�#E�J��d��{��I
�,LO �'t�d�f��x��.�h�@;T�>I������0�0�8�g�O�5J��Y :أ>i���է+9���6'М2�.���H><�!�$��a=2 �6� 
m�DM&�J�v��+}��>%>O���!�xİX�P�,:�Y��'I�I�^�q��ǃ4Rv�A�mW�c�T7ms�X��>9�$q�%�T���ֆ7k�Ї�	M��\n(p2��}nu�4%��:t�����rFH�.�� �so�(�$��������󤋵.	0�B��nT��oP�=�!�$βq��@��͇�h�aV$?U!�$�8��"5�#a�T�#ω��!��=`t4���E��uڌ�oY�I9!��H�q�Dц�΀��բϝ<}!�� �l�'a�#O��1��Ӡ=�l=j`"O"l���G�:0� ���	H�>-Kv"OQ9���h�����*Tuب��"Ovh[���H��Ƙ�g�`"Oڅq��Cz�^�8PF�$:X�e� "O��§ �����fW�K�H	;�"O>�q�2<X�0�Bc�?nԮ�S"O$�*�-$�꒢֐(���>O��=E��o��C��	������7�y� ͪy������ƀy�&�ɦ���yr�;fc��+��Y �"��F�C3��<q��9^P2���^<R@��(��D�!�P@pت"/!,��pDݐjV!��9HbPBB��#�%0�O�ay2�'.��'��-�e��� �eK�:��)������G{J~�H�%*�N9��%��<jDl���U�<iVC��9�r��#NS�n2(�4oUP�<�G&��%��dr��� �ʍ�f��J�<�ACX2X�0U�D<xB��H�<i���F�@P�DN��,pR*�O�<�p� �}K�a���;��-��fI�<1f�4V`x"���qlb��V�TAy�>I�~S�@�r��3��K3`�7�8ȇȓ,�8yK`�j��D���4DVЅȓ|��X1�ּ+��Iץ�����>��'^a��!F�E�����X$;j���h���y�Ӳ.�"{�퉾f��	6bW4�yR`��oQ��Ŝ0^���d͚���'�ў�����}��:UO('�4Ī�b�� ��ɩΐ�C�V1��)!F#P��$B�	�vFh����>Gܹ���XO��C�������_���9D�E�JݚgN-�I��4�?�N~u^3����G5PE�D�Z�<��O�"��)-�k(��Ӥ��R�<!@M�R�@i1�@7DU�i�� CP�<�g*�� �L5r �F��B]K@[��xr��N[�I*���X00IB���
	�'���Xq/�"�Pɠ�אLj&hC�'�Mۗ��?m�y��ͣ�ź�y2�'�Raؑ��Qb����?W���'�r	bJ��A.����I�`,B�'����p!�m�d��`�D�$la�'<��wA �UWȴ��N@�\q��'���� ���������QS/WPg��<E��'�"��wd9/���w�9S<R�'yj�"��P�:eI�-R��y�O6��$�.0�y�Эf��=5Ě�w�!�D�&0Z�G��(4�x�#�H<!��8Y�f�PA^g�RM�F �I�a}��>�5f�Uu��9 0`PE���x�<��J�{�|�sd�4v���A���y�<A��&\0c�j��K�l�ԧ�t�<�uѮ	�U�fa>R�$�G`׭�hO�gy"�O��$�/�$�
�I�d��*1#ʽ��C�	0q>�%{ՂJqar��FR"p�HG{J|�(H	Ul4q��%�a�`��B$�O˓t�NU�׹GU� ��)Q6v Ez��'B��5�ѨM'������H��
�'X:HpE&�.7�^��dJTNdP�4(����%~^>т�	BV�D��|*!��6"OL���g�s�6�JlH�h01��qމh@Y,��c�Y/@�D!DxR*^`8�tI��;$��e��|E���1E D���f�S51¼=�bkk�)���3D��  �*E�np�	�H �U�BP*""O�P㫝}5�9	����$���"O�2�-ʻ_:¤�7� Jèe�dY���A��o�'O��a��/{�z�ВPTR@y:	�'�ؕ�V���F�xmq�(8I^� ��O
�=E�tI?��0!��	0N���Т��'k�`V����A2���V���K�<���cџ�yR�O��"~Z,�2��#O\�9s�yi� ^z�<Y�@BR��Y������hO���<��nX�A�X' �Bh|�������<9�;������Z�pLxtf�;��x�_�"G��%_V���I�+��O2 h��IGh�BՊ�*� W��APLP�p�1O~�=�O��$�=�$�E �'�>)P�l�9�!�d�$<��� �"�`y:`I��l�!��@�]�T軂#ި �����(�<�!��+x�;�L�{���WW&:��IEy�\��$��'�� ��χ���y�� ?�E��'S�T�2MF�+�����R+L����';��3"�@���5����݌pi�'%|�q��]� \����|P|��-O���Xm�4ب�X1w%�T��@�%�ay��	�L>�sF�%,�@,��J# �C�0M	��H"/�SZ���@� w=�B䉸[���E�({Ȕ���mK�T�tC�ɂ9���D\��v�P,˴�B�	3�t�
�@��$n�h��Ό .B䉀~��a���F�S�Jp��c��L�B�u������yx�VnХ*~�B�I[]HԘ1mɏm�R�!6���aoTB�	..Ez聵%� G�õ�%�8B�I&`؝
p�K���A���hB�	45�*,�qoB� ������`Y�C��U�xK*�=88�[r	̻1�|C��#3d�r�`]�p��Ș���}�,B�	�G�Zy#�
�
3 �754C�Ibw~��
*��6��]�@B��'g��=R1Mȅq�:9�DU$M6B�I�56=Xk��U��*uh�0D�4B�	rN���1e�4�B�c�*̛7�C�4v��<Ѡ'�'[<���/�~�C�I�AL-�R��38%#˂9�C�IC0�����,7L8��`�f/�B�	�-zL���!�R�Aa�L�jC�	�H��६�D=N��'��s�B��������[H��(��B�Ɉ������oa�P��M��fтB�5�jL���©$��#�`�34�C�	�<��xHV)�<~�@�P�*:B�I=Ptp���ظ`��<z'��}�XC�	�q8s-֋$3@�0��H�o�VC�ɪ6�ʥ���S#f���A ǅ\oHC�	.Z4@s��!���K�!�C�	�i��B��>���[����.�B�II���R��N�nmp���f�B�Iiؚ��Ed9N�R���D+:�B�ɲrNN�";�(��t�6wbC�	,<�� ���شU���� �B�	<Y�*��䂗�@��Q�(�0w�B䉦s��Y f���\����J�B�	�Z.�� �{�h
E#��t�8B��y��jnO$�lHb5히;!��釫�)a�����L���,�=�,�Q0f�?|���
�'�0u�v4�ě�@��s�\ �
��� ��1MX�h,�IFW�Z�fy9�"O��3uoҤzwb0��.��	�p)�F"O�4�	R�\�dpj�䍉*^LZd"OP���aS�)��+e�D4h�$!�"O&��T�ɴW�⥲b"�r}l�!�"O޵�P�@8�Ԙ� ­6N��S�"O�h����9u� ��OF�/NN�i�"O~���↼5��,2�5]BTH�"O����js!R��el6+�0
�"OR�2&�`�j�a���$��II"Oҡ��L��{�����˪:�H)�"O���C��=�Z�����&Q�J�sB"O<8ac��lX��e
f1z�"O*��
��xv��1H��%z�"OLi�"��n|���c%�A�b}��"On���,�j}:��re��l#PH+b"O�p��h�QL&l;GAˎ|�e�2"On���֍S�s�n	���Ahw"Ovx�t���*�iڄ�X�%�"8h7���c���'9܌�z��O��(���L1?�Tm��툭Fs$��	�sG2H@��+�@Q��+`�l Gd���I;W>��OgZ@5�B6Q�X��'�����7J�6��N�o�҉��t�.ճ�X?��B��V9':�ʷ��;a������O�ff9�s�ê~�p�;&JL?��Iܧ&閝K� ڍ\���1����E{��:d�,�F�ע@!v��)g@�IԽ2�IF�g���v�/u�J�ˀ�S�P���5B�v����L>�� Լ,���:B��: �=
WN˦���%�\�J\�7���C�کZQk���(����L4v8a[����胈#��d��46<X���9��,�t���wҭ�䏙�Ryˣi� M�&\b ��I�����v��	��1g"ӼacJ}`dM�Oy��l�8���W�]j٢��'�p�	���ąѱl	�ip��	
H4����'�J\���Yab���Ø:|pv����l�I�L2���O?1�0�h-�В�%�w�:��g�:qT؂ƒ|r��vD��fBO/=TFMGR�|� ��1�O�Q���2�����k����dA�Kw$�8��'����Ȼ���炍3�����@��:k�حۀ/�m.>���nă1�|�������z|�v�
o�Xx��ֻi���?��;u��Q鞟\s l� -J�b�Z�!��c��ɑ����
ը� Fɕ1��d֞ @'?�[!Ϝ�^�D	'Oŧ<Ht3QC�;���z��Ζu�NH���5>>#|�b�&p*��$
�,$ 4��z^���F�I��ؒ�O�}ȳO)'3<�$>7m�>��� bS��K��!�d���
�F����=q��ű��+�����*	��+7�[�(�|���?i� ^�Nʘ@�w.�"yp�r��= �|���2�W�T����2'S�S�	����+v��y��+=���#�
�2�� ԯ	�����<��T��LA����� ��=�� ���K&6��(ďZ��?���I�F��ƨ���Q�O[U͜�T�ԉn��\���6h��u	u�H K�@����O��U�6��WȖ�4��9E����5)ѴB�x��r�w툄k�)X� e��ǉ-/�i1�.�8�?���зD�l��BB�T�D�-^^xq4b�����5C"�x���eWD&��2��Z=��x"
֬]Y��H7P"|%�kƲ@Fɂ�+�4߅�j�5�\�i��!p#׶\i@���^����f^�<fM��y�G�<{��ص��H \7��q�(�
�b;{�YC�s`� aw�B,%%���7�I$@8�&�s� ���Z�y�yф�(7��h'��kp� p��٣[�%那�sZ�ܢ&W�\8�$K�9?�I��뛟 ��;v(ք�~b��P`�@�w��^YY$J�#��y��M�x���8���aI��k.�Pc�t�7I���xu�d �R2�9*A��8p�*FL@Ȧ�3w���J�Y
�g��YϚ)0Ac��2D@&u�,=�c�@�g����]�z���a��^�d�K�b.'���'��8^h �U�F?D,���jA
~���FX�|�b��%���"lF�e�N��C!bح\!H���.R�ࠐ��;,��5��j
\�R�����#���,_&F ����m��DK ?�y�QV(�f�� �Q��?��#ܖ�r]��LG	�3?��,G���R�٧9�0��?5P��,��,��mʃ�����U�/�J��"�&?�4�#���;?F��l�*,����"��wC�B�ɗb<Qbٙz#b�KwD�a����,ЋO���8��ȓX���C���F�0�o�
l� -h�h�6QD�adA@��f���ˑ�c��)�%�C�X�Gi�0V(��ڠ���-��1�
;H̼��ǃ����-S�UJ�:��z%C��	}�����&b�z��S��+P=��Ɛ 8>�H��kݼC,����}`9�C���K4�ۂ* �/O6����	l�d8�T?Kd?@c>8q���"t��1eC��C��]�t������z8�D
�Ck,!���>L�a�3gE) fGs���s�ʊ�8��P�0��J��>��`�P�HO��EI8C� ���ѣ ���v�A�\Q���JQ<,�b�H jSl�%��F�
���oѡ%��$���4XY��#Dd@"n��9���p-j�o<HF)���XԔ�����z �ij��	�Mǐe!$aR����hQ�ҥ^"����B �z�kΎ� I��B(H͂Et�����X�xbڨ��T�矜Oj9���ؤ�HO.k���Fh���cO�$����&̒�1�@M��@�'#,|�0�HL��,�x��ӛ	�m�bG�!�ΰ�1���<as�n|����AN�K"�]֦mʁ @�+���� {M����Φ��Ri@�����$�;-o�h�����/��6	���8I,���S�? h䒱��<ULLp���:*�0$���ƮJ^�S��A�옄�2-�l삑�<TIPHѮ�8.� 8�8�����V">Dl��A"�~��C�'�x����1oH�5�Q�@Wqzy�s�Ҹ+�.�������I�D�|�p�-��c�����m�([u�">!�h��K���6Tu��E��3���2&�|OH���OX]�1�a�S`�I4��rs��i>n���H!�Y$Sv�#�eG�:��
`�$ŀ�c�-8T!�l߷l�t��l��O>����5KZpABb���qS�� @��D(Z0�-�����X��LRUQ2n9�]`d�[�ة�+��W`1�փZF08|�u���#Z�G2:6��8�ri�7B�98�Z%�w��\՘%�A��'|&���c�5|O�t�'B���t�d%M��w
�;$��k�ͦ#OxH����/z�ޡ; �;��`�DG��ިv����Pٺ�@�/wJ�c��Y�?ດ��I�x��1h�@�c]�
�4P���(�ZQZGC��1�1r�(�E�,I���U�v0xS�i��e�h�J�'�,��1��H�1{۟ظK�>]4a���$��ۤY����ӟ4�Y$�_$HeH��#eԝ+� �!�.�A�a��9W�|�%�^�=Ӯh"�#��wmL5�e�_����
& ?|�0w�աET�t�5�>ғV�4M����^��E3b�7D�hY8��&n����k[�$��A;ԩT�>]�V+�=\��E�5A�vaX�mR&AG�}Xt�_ ���p���eEI�^A/�8��'��0b��C�z����RU�Q���V/:��꧈j�zq�E���z��CA�/}����n�Ӻs6)�5�M��4|�!	��G.B(�1c���4\�<AaJ(���4]�8Ei�'�x�b� sPy�k� ��a!OƍV
�l��>��0�Вcwf� �I'iJ,,�B��(i�`�(%�i�"�`@�C>n�5�N���V��0*pY����`>�}H����.��4J������;f$d�p��mN���j�!�r��f�7"zq��A��(�(
�,ϐM��ܴ$~\h�#���Ѣ�٦;J�y#b��E��$�|+B�F�D���ƭ8[3������-w#bM��Pi���˥��i���r'bVR���-�;_=���N�r+veh��k�,t�ď�.b���ʃMyQ�CJ�*]��AVp��ׇ)��Y��%-cIQ�IO")xe�2ɟ&�Q���,*J�8��"?7� h} ��U�ɟ�b\�Ć�I�%�vg�?�u���<p8�Ah�v�i��"ǆ����ӀB�AԾi�V�� �֣�YZ��@�k���B�l	"�h��`STn��l �Z��h��U&K4�T��m�(5H�a`Z,]g�TKq�?H��:q�i�P���͔n!���G)�D�.�"	|���Źkȡ�&�x��@�9-�\�oں����4Ü�8M�XE��u�4�c��M?��:7ʐ7@�͡�6����e���w|�$IS$YܦŐ��p�B(���%h��1.�r��L)B0}� χ8� ("�䚵>�^���R��b����!3O�M�s�Q<}� �G�
�:*�$�6;�R�0��5��K�n�#�\�A#�"�H�[�E>V��4"𙟔���Kx���9ԠR)3/rh����"� �W�\�y�����샹HR��0���X��4��I��l�(����ɍ������{�𕊦�OT��p`*P?^���	�cZ��*ģ�����["p�j5#n��d#�DX6��j{h�*E�3(Dn9�A�bJb��FG�/�MkfE��Z�����!yJ&t*Q�ɵz` �KN8�7����x�7A ���
�Z�:�]��H6-� E:\�ɕ=&E���҉a�!4��4K�R�3�$���2�Pf�>��$I�BqJ񌚣u�ҙ���l��}�0��?�*�ag���x["��H��� g�.p�r�T&
%��=!qf��1��D�5'�Gn�x:�aP1(þi���2�H�L�	�"�)oʅ����?%�U U:�6��7g� \$�5Y�N#'h�u��A)r%�Ep/O�F�+��B����0W1a�EW�4�ʣ�}#��C��g]z=i�ϙ#9p|��g�߯�j��7��1�+O��P�ᆛ�T�+����k��c�EK�'~��Aʔ�ո��戚05^�� raG��D��j>{åK
!X��6�S�V��lX�R�9z���n�05q�iJU�*!��� ��p<��E7%^�P��� 9y�C<VhcrAD�'n)����t�@�����������<�)X?�9�c�L<�����FE�N��䃞k�z�
׍sv�!��땯L�je�>La�#�۳�PݚpD�"P�@�ۑ ��=p�9��K�	E�8"�딼Fi�'���b��/3��3�P�NE�*���'�&tyEH�� �r�� �U�d� ��
�V��p����HB"�!J�pE[��z(�@�Ǎ�$0V�D/��$ɐן&���{��!�GB���uG(@?v��\�T��=KD02#���M���I�����I	Cj��� ��{�ZY���:1��H$&��u��>d��ōO����7���
��0���k�Z����ڈ|��H�4:l��;����w�2�� ��'�4H�m��V38%(��;���P �B��0�#ӃR����H���2@�'V1<)0��ށ:�����C:��Q�}P�E�W��Y��lk��3@��g�ٕ{28�EhQ 0���{�� ���H�I"'������_�3a�<"�"ҁ�f�" �� �<a��{2 � %��!�_ �C��9:�HS�'Oꄈ�g�nM`0 c��W�:�X��.ړ:%.ЉĚ�����!L�t�� �L,X�R�qJ	��PN������Ȕ;���  O@����D�ڡu�
��Tj�2R����΍VK�p��L���O�x�Ӭ6��x�e���X(�4?��aa��?�J�ů;V,y�c�3G�t0�`�+1�F�����5=��(s���	�ʜ��+����f�X!Z1U�d6�h%��gP0a̸�E�1^y�adV�Or�H�&̚l^��H�aT�Ix9��'0�&ªM2��"���2Y�zqV Y�1Ut\��1\V$���Ɠa�yJ��&X<ys%D0\�n4E{'	i���K�(Κ�De��GK�
~���o�=1���1���'ys�,�@��n���c�h��VM��W?m���$�A�Ē�
Ť���F���e���Д��O�PJ5|�.� �`�;OT���K=z�����_,�h�A�m��!��㆛�j9�%�4u�S$7��kȯs��� N6S�l��C��+"�X'�ݗ�"q'��P�]�(e�m8'��: bӈs�Y��8O`��1���~͑sB��C��9��2_\a��֞=*@�t�ٓм�QEԄ�z��BՋF�����0T�F�l6R��e�}ƠA���=�4����{^P��,�66j�1cр��>(���sv͚:�hT��4k�@A �/	B�0`b�ƒX�>��޴n+���A�F�� �2����!���E ���G`X�2��4��=;c>���#
x	�mS��"�����=.1���wP����O�	��i�r�? �DZ�"��)�$�Y+"敳�Í'$vY��Arܓ�*�����r�J5����i6	8�HU�R��s��m�Xi �P�E��a��*��v���8���k�!Вm�X0!����^�5F��4��uY���c����Ô0��$�?�A2��ӌWȆ��EL�}X�7m��N�x���ٰ4�(�Y 
=lgƕ�H��i�^��EQ	���Ff�8/�`���*�"76P`!ՠ>i`̝�2(�,k�T :��E�S���7o
��Ø5[�����-�z4#��2�I��
��E�4�!Hǂ1d�J�Y7_���SD��/�hh@^�B.f��	��I\P�g
�I�"F}��պ�!�9{2�`! ޅC-`b��xq��G?�QV(��q�F����fPe��`��u'�N��� �U6}5�aR�v�^��t��e�#ۧa��u�G�]3֢@���>>�Gk]5zc�%{A�Dݵ{f�+�K�N|b٫ @u��A�g�͑w
^- �KK�L�p�îm@�a� հ���Do��6��F�wXk��ʞN�`�0�O��Cd.�3�%���D�:L`�e�s?y�	'/.���J�e؆j��ś��l�`��.��j����w9DD�#�3<�ұ�CwJ��i�_9�1������T�$�)0�t�S�O��p�@ ��R)B
?1���#C,E{�Yx�a�4�"���ɉV5&�r��Z�ZQ��<9��H��KF�ҟ+��)�JE P.<��,��e(�'�T`b���ʘ�yr�٫I�:|��D���(���P�z�%ƶ@�P��^��
Ӧi��E��P�
X�j�Ox$H6j�%�!C���4x�A�D��e���X��L�C�1*V��� m�X���Lt�e�5�����`c��� ,�����^�<�#a�ʹ@4��[@�۩8�dE���a�la�a��V/��!D��y"�Ɛ�J�q�`��c�h�SW*��A�����"���%5]P!�P-��T�IH�E)t]�IJ�%5�O�A� oY�&���c�F�|I��ە	���K��9?F�I�L��u��ؼ"�����K�H;��49A�.�f��2b�<( =Ss�'���	��Hv*�ȅ���q���� � �y��ͨ"�F�k���xt#@O�VzԬb"�8��a�П���
��@�C q�:�0"oAbj#>QA Bz\X��YC�!���|��Ϙ)H��1FK�Lih����}����t�e�L�$כo�@!���O��y�B�^w��+�e�(_S x�s�O�����_�*+T٢bA[�Bf��O_@��E�5?����#�zM��%`'��ࢋ]�TI �p?!��R��`hb�ʄ@a�H ��
�(Q��sU "ӆB�t�T�x��C
b?.<i���3o*�P�e�Y`��](��8��� Ԝ3"
!�OF)���]��.�A0�Z4L
&T�@D��K ��1-&�m�t�6N4�2�D ?�$�Y�:�s������*�4���ۿ^��h3��<��=����O�o�x�d�ݐ� �RLĢ/v��
q�1�Mҁ�C_�� 4�O<_)��3ړ`RB���	�j�.%S�H��9���O^YZ�Bъ۸����֝[J�!ò�\�>!Jva݆��@��=
�u�%O�e�~B�\:s����B=S�I��hOp��.��)I&��0O���'6k|)�.�c�88��*�ŭ2D�\���N�2Bxl*3���Q� �b���O��1c$G'1T��2�lЯ�~���Nwf�����jdj܂"��$P��C�I�\]`T���6wv�C�,f�a�'w�����F�'��18ϟ�PK@K��!�l�R�ðUhT��w�7�O���uM��()��bF&�%gx�%�A$��W�`�ۯ�x��E�M���^���]��V4��OLQ�
'��OX�	3S)�Y�^��v�@�D���P�'�D����r�\��U�a� � �'�(|��hP�4gB�,��	��I1�'~��#�=\�@%�di���'�C�,�1|ΐl���݋f���'"�XCK��dCd$�K�X\��'hV89����Z)q�9�t�'����G^�S�!s��� |"�j�'?nl#���?=�Ț�$y�H���'� �УF�K����!DؑD{�(Q�'j��8qM�ۚ����i�̙�
�'�R�����}Hd`yL�d�d�	�'ɌU�b��s������^Ȕla�'� �[��٨t���
 %��M�*`��'�KG � `|����ٌ
g���'�
M�%�ޞ-֚M���O� j|(:�'rD�f�5����b�����'�f*6f؍TΘ:�
G5h� p��'PNl�cl��j��)�I٩?��mk�'}�� �a����MR0�XpB�'w��ȕၼ}ގ�t��;*	`���'��\Q�G!o�ԩ�th�m	�'�Z�"� �@iy&��ynR�a�'��LG��ˮ�B�,��e���� ��ԥ# j�q�aK]����"O<`A&���S~�%;�Ƒu����"OLu�c�uE�@�$��&ꈭ"O�����ܱ���)�1�t"O���`�%Dlf�:�d��M��%��"O��0��W4ڡZ�b:�I��"O��Bc�و��D���&�0e�w"O8u
V�=~,�(SG Q0�\4Ip"O��9���_Z)r��T�$�i�"Od�'jA�'�<����!8�N�"O��h�O��R*i C�\�X����7"OxS!k]8W~��c�B'z���"O(����5l8|Hg�*�z�!�"O���!�#DN���r�K�4�x��"O"\y#�Q3I��X$O٭$�<�bC"O�h��ޫ8p��C휭s�x<�u"O<k�.�1P<���įs��p��"O���¢PJ�L���·�(�( �"O�����V3/Ԅ4{g�S'����"Ov�{u�5�;�L�E�mp�"O���-�(-�\X[�-��4�@p�"O���h�;���[��L�B��� �"Odm%$,B~��I�Kԕ~�$�A���
?g��$��'��� �)�\�� �b���>��1��A�Є��	IR����5<C����Ȗ.����dE����-^$ �O���Rl�%D�<|�'g���}"���v,O�I��ܢ��4�l�)�j�5�,��!��F���@�
($�Duqn�+}y���˪�jrϔ6��	cܧ&*�auƒ�	��Y���ūVu�D{�	�)F^�����uQ (J�*��A �)�����`�
!s0�� *K�Y@̵���]��D_�Q]x�:��L>�[1ǔD�R�X����Ԩ^���X�
S �p"Q�r�
�o�<BXG�D��0R^��c'I[�b���4ŏ0:΄��<r���/�\����kp|��Z�A��5J���� ̚f���XK��#��� ���S-jvp�%�>G��5"p����(�$�D~n=�a΄7��H�!�O�|r&��<){��,7ָs'��P�q��������s�ѡ�坵.r�	��`/:�+QQ�'\x8�cw��@IS3��#��=ғO��� �9����'Q��pi��K�`x�I�N�\5�b�7*��-W������͔z"R���-�b=�8�^=�'�6*��J����^�|�����H��IY`�N�>5��h���/���IY����S��O�'�uOׅ7��S%E�V�<`ɗ��Wmducˏ9SY�!a�.C~,��`�V�`ѷ�;��'p�1�&����̴�+�	�
�ig���n�
h8A��z�d��A��[�O����i��-Z#�
'
\!��~'��0�J�0�Ċ)Y�d��MP�s�`)���4ML-;`Ѡ<H%i!�F�b�R�fHH�a�)�� ��~�(v3k��hH�iQ#:Z1���`�P�S�I���l��(��c�9]���$M�G�v�1 NҽQ>�	�p�%��gA�O�R٘T+�%w"U;G��?�A �P�w>�%��3�p=�� �z� g�]��4�Q�Z��I g�t4���H��r)���ߍ���Cv΁�Bg�	3�a�f��H�ܘxć�/~t ��[a����O��Cwʉ�RGF�0�u��ƚ����s��6j�
�䅋\Z�0q��bn7	�B�H��E-�䡊u����?���T� #H�r�
_h�$�
�g�d sW���z!6 �c߰e���Qm�3u�� �B�u8�KF	�d�j��)������xɌU�B���iA�T��� 'E	�z2�\�xI�f$���?A����#9�A��&��9O��PgEG�_��%Y�.�.W��@���"}�uAn�=J��b�H}�j0�7�����.��P�L��"|�a)��J��:�
�2qpq�,\$�(e� ��#@�^s�ֆ3��˓K��R,�[�,gg��K�(ȗ'q��:��/4a���I��6�r�gJ(d���RF^?�`dQp..Rv��:6(ڬ5e��べ�����-��9�GB�1U	���1hG�x��x��t�J�(�r<��6P�-�z��	`�dIc�m��k@+"�X����S>8P�:�ģ �i�Oҥ-�"ɣ #T�F�F8 !͒`�*I��'1D�Z�O��A�o�?�℣<]�q��v;&p:d��O�8a@�-�)#C�@�ъT�
*y��B��r38LZ�+�B@ߥ_b�o�M�~��"�M$/��i�U����?لlW�-��l��M�$^`�3?��$_a���EƎ�~;��Q�?y���u"�Xl���GcѸ{T᳇IK�P!Z�еf��{3���}���Y�bĈXc��Q��B�RF��B�z �I�'aR:H`�O8��p���e�e�p�3����&A��s��=���Zq�8���
k�\j��\��J���G1	�����
&v���p�O�AhDn�\�h�r��5�U)���C�'m 7F�,qX�E���s͸<�����M3Ư��m�T��2a�BR�k �^f��e��T�,V	R$��>r�1�' �`xu�х�ı�O��RP�� �u3K#vѪhS�4P	�Ḣ��6Hm|�:d.��n":C��,H�u��F��B�}���R�mr�>�� Y�p�>�)�B9�٤q�8�1�Y���O���P��OȔ9r��E�t(������(q�4�#cV�q���+��Ѝ҄MϘ-2Afs%� ��4PCg�����EC��R'�p ���u�^Pד6J�+@!\"Qh]�!��5j�A2b_�����-�݌I�&[�%'�勡oJ,R�~uȡ-�7o�yB�~�)� "���^�2��ebYQ��p��5)@@@�Oʆ��
�,F(o{�I�BAĆB�:��կ��h��#��L�xÏ���*�/R�}����4<O:��p�� �� HGKȞ+���׵i*��rdT�|-��T�>��x�Ł�(BR���V�<TF)�CϋY,�J�F��"I�."��a�(D��c+�D�����G�2��i)G�;���Z��/\�v�zS�ޔqvh�CkL+D����eJG�6��Iw�f��@a.�_���	amģN��*�`#�O�2��Ï����^{���'��>W�D�W�À/h����O \�ZbA�})h�����M���G|�I@�_N&<��ōx��I1w���e�E%D�ԉ�m��A��@!q�^�8�r!�)���Y�Q�aI��:����dQ ����J���д'��0�$,P�.Ѩ�ݝqr1��$;3�ܾi=�xh�-Ԉ_jVLؕ	�2��	��Ҡ��K3�3�I��j����*rL���iȡ	a\`��
�		ฉrG�.{���@f%��/y��n��/4T�bҬS=?�F$����)6�9Qw@Ȓ$�0��.b��(Y��S�R!b�4=��и���u�J0˴cR%�T�#i�(g�$bO�2N? �yA�<��Ԭ;:�����O�N�G"�yj����џp(0�߈8�鑴�w~dl���1���Se��3m�0�G�$z�[�
ɸT$,=�&�â��i�G���~B�6R�+����=��P%�1(B�ABs��:��[.�	S��s�T�NXy��e�<qe�� ;�^����ŗ��$fn�[+DmJ3I��[Oƽz1#ʪk�N܈�b�Oa����)9���V��Z*D#=��O�&T�8*bi(E����'g��lEu�$�L�*�ˎ{}di��'V�2	2��F���������fABs��O&X`�'$jht	 hͻ1ky��BE7]paz���6����ƛ� ��T��M}Ш�q�ڍyk���a
��O�:Y�T'�8>�ɠ�ƚ��쭻H�<�۴�M��ft��Pǖ�"��PQDȯ<��O�T	q�/�ybg� }xiA�J��"1Cڐ
{�y��l^�*�x�p�ϽA�ȉ0�%
��m��nK$��#�	ܦ��T�xӤ��b	Ç=�5�'�0�.6��5oL�(r�a��FD�]Wiδwj�P�ִi�0�U�I�m�4���̛mӂ|94�V���󶮓m�°�F͈/Cކ9JD(X��qa�)s��:-�wB�����I�0)��
�Gֈ-jO>��G��FՀY	�`JJ2�؉�$D4L� }��U�7����Ȟ}BRx�D,R�=X}ys�KM:���wD��M�0U��AT6�xa����`�tc0�C
X����R`"�K6��	�+�B(��.b
HixQkP�bXFX�R�ăw����fB�&a:@���JF�nڗs�B�����k��C��
P�JYqwm�L-�n��Bq���B�9RT�A��&D��R���K�$H4RV�x�ڌ���r>v�ڄ�ǣE����)	h.N�H7��l?���KdP(i�!�)`��)���"0�t������2X�ћ�J	b@2H��
�&�Y!yTN	���K��I%5knp����S��{�ឞX��p�FN�d�+u.^�����Im���Iԯ���c'��<?�h��ƌ5N�i�b��/X�i+���}�<�#��U�%(��m�2l��q��Q�}|�ڣ��(@�N_���(%�@	 �����Kp���BU���!X��V:�|1�]�s)@}1O[�Ft5�ӏ֣.y�={W����=h�Ė�lYf!�#�ؖ{�u#�ՐbaJ�����<`��!�ʀ"C�
/Cs�0��ϝ7kjt�"�ͫ4֪��Ī/�^`�,�4l��x�TM�mZ��R��{˼}_�P�ĭ��hH����埮Y���ȤI�^�̓�H��5�è�~���O�)[q�� +�[�(�걬�?Y���ҵ[��\䛅����t���)Zr�G�\(����⍾3*� �@G�,�HͲ�!��s#
0}�������ፎ��O;Z Ա�-O,@�C��	J��� ΋�W,�d(���:���� ��<嶐Ubd(L�K�hY1*��	�.L��gV�5W�A-_PR
D	�v˥E�s�І�ɨ*싅�V�[�}i�Q1���0%-H,>c�)#��s�9#QKۍRԎ��SFa���2.�e"jeӑJ�^p��#怩�q�ܖ&�đ�A�X����+f�'�~�����;+@. ٳe2��="Wϖ�J-Լ��cM�&K���|%�P�VGw2Ұi2ᐱu
0�BΗn~�0W�'�����~"�t��W��bed��*�J�/�=~�r� `MĨWC�q�˓,����.���H�*�6�8�z�O��|P��UN��9���+X^��y���"o�N��Iߘ7�ԥ��%Ȝ��-�f�T�>��x��Ɠr�f��WC��5t��3H�hYf$�.:z8��H���8��`���Fs�h��W�K2f��C8O��		 <���48V��BE��p>I����N�V���� JBωڶ�����1��qI�
�#'-䰘q͊�Kb��)3�����8b�B�Ҥ��T�I3��i��y.ꈀU �/DZE'.I2.@&����.�I!��K1�ĭ$`arj�:tC�YI�a��qT�` D!`D �P���)�����U�WD
F$���Г��'Z����?Ad�`�q��
g�Aٔ��$p�4������f�~��X��@v�l��c��Rߔ��i�	 O�PW��0<�S�h�i�;D�nu%ƒmf`�5�8m��{tkV6Rf&}���F����&q#��|ڦ �_���a���Wo@�(��0d���5&����	�)w� �1b�A@j�k3�]/�±
wO���� T�V>4%��� )��r���\J|H`D䕼VĈ�*�������$�DBP�S%l-�����?�Ɉ{�����/�+�������'�PT0�f
�w����1阽CPu��1n�9��Y+������"�PhXc��~��ߋu����!��6?i�s2Ê/W��`WJۛ�hO~�Q%������R�Էy"ґ@�����"mGl��t���F G@�#�����W�I/B��0H�~��е&��A*�ҟ�@ �םmj�� �{����P��z���R��Hl�����V�d�O�.�I�'�~�$�A��pu��Qt��`mVdC@Pd���S�D�
�Gݒ���`��F*���T�>�����%�2fߓ,��a"��q�N��)�0/j�!�k�#�`�i�Ś��-�����s�
4>y �.b ���*��ي�!�  �D����~2�R��.~d!@�픘�hO��Y��Z�0��OŤ[�}@�d���Q����E%^�Q0d$p�h���ŉ#)�@hnx�4�G�M�z��Vn�dx��⃘�RHbP���i�r#>9�l� uVrk0�I�k�,��уZ��*��9s��R�ǒ+���eJ����S��-)j�OTf� ��9Iz� ��I�z�d䱃
ǲ2��<C�%\�X�@yf�|�ܽY�PQ6��9�v �O�1!T����A��<��� �����܈
�Ä�@w�}R�oY�i�X��`�̫9@�1dG�'"��f�T�	�֐J �E�F|�YB/�ɦE���*CՄ��F��<(v�]�"YB�
4��0)%`8�Q��f��Y:�%T+@ݐ4۲�G � 6�&%UXi�����* =!5�:������[��E��&#�T� � ���X����Q+�O������2��U���ٓ<)��X��">�`Bs�֟ �#��Re�)�#n�"���N
l;@���Oj�E�Vo�Hٴ�x�ˌ3|R��;�n�>�������'~lҦņ_a�����\3Dw�d���ȕ��c��Ƶc��IFbN$c�T�q
��wcph���؛c-� ��h>��f4b��!��ρ#o�H�Q�ʮ}&z�÷#�uz>	JD�� ��I�����(ɖ��+ދZ���l��?�jacYz]d�SA�#���zTNA�O��U�3Qiݎ*�o*D� l��
�9�Q��m  �εjD��M��A�c��k؄7�>8�Լ�G(&b�	�GM�mΊ�ۣx��}��P!O� ��X�>���h��g���$��iƘ�Co	�n�buq�-�/Gx���#G�0����
֗��j��	y6f�Y���o�dy�<Q[����
��)�2�HQ��Ja"�s!�L�Ύ��(�	�F����=�d*�LX�/�(�8�ͅ�Lj0�K1�쟌���W�6�eY�F4r&�s	�<
�j�)Îٗ7�nb��9�.�3�xpK�B�"7���z��
�F�Ze���>�p(p��!K�hp$����n �$�tO
G�Vi� h�;�l(�j��<���F��D���Z�Y�t��U��~���oѢ�zt��-Eu���c��Q$��f,C�f�z4�ϼ>���` �{c
p0� ˕B�F��B��	@�'�@�H4͔.z"0M��(���WƅC�`\0�%Y/y�`X�ᬚ<vhJ0x�#Y���g釧ˢ�[�愃@�j\��Y�}�vl.�yGm��jA%��SwZ2@�2��]��̧O�l�L�Q�1��$�S�����ML�{�8(�@�
Tj�p��I1[����'L�>Y�f�5�M��ˍ�}� =HF �Pm�`�6T��S��L=u��9k4��*��DSB�o���[�$��B!ۿb������ߙm@������[�� `�:D0 #�\F1����1EM�*֬=�]�U`Ւ{ڊ[���q����Po]�HxTgCK%J����Ɲ�Qdw<�t�t��r������KrHQ��
�M�b�P7�	�;�4�ҮB��+P!�&a▴�@؟��FPݥ�$���@����xxShůGN(I�A��p���`�2�L�T�����7ON��.L$+�P������<q�ǳi�a~҃��ri0q�%�2'��C� �d���LX�|YH s"i@>#^�Cπe��E�#��k��ĉe��	��l�^�	S0�!�.gQV���N<�-��A� i$�⵬
�[ڍ�'l� �1�	�
�Bl��	І;���f	Pq���`iE�O�A���@���dG�(*�B0g[�/�(x�a�$���ւ;��8!E�	U,��"��"���h�A%tk��)�XPƀ��q���G���"-�����	�L\J��:$Tb$�0H�/�л���e?�2C�C��iq5�^t.:�!��/;�](�o�V��]G��u���T�X�R!��Iط�����=�&9����VS�I��KZ�~sv���(I�[��[e�68����g�+M�����k;WQ��>�2_%B�Z�J�*�t��m�<Y�?�+و*2�����#��P�h[ީ����d8(x�F�[A��޴��I ,��
��T��(�?�=9��V��F����%:餅��c�U;Jv�M�{�O��ꁊ��P����Ǌ�n'��@��#����$�m	�3��7�p?��H*�! �U/	T@��I[��Ōʪ#�D�s Ъ\��v���ڔnHش��E 0z�07"O�1c�Z�u�t����+ZD��;��'���x� ��]~V��u��{?E��Ur[8-{�gϨ}`����U�Zz!�d�}���rI ��O�-mT˓'E�5)d��>�����Oz����� )�@�ꆶ_������'��=񵢞7y[�}��Ԃr�|�2�a���^9���G<��L�o�`$4(ب)�$�
���a�'s�Œ�@�`�'3p�lp��N-+�
�~�=��aVtCBތFg*�rq��_*(5�ȓ��!���AU� 5I��(�t�ȓ50�]�w!�D��c�J�IU��ȓ-l�q�RӵcpF���+���
��ȓo ��k�m��ȷ�+�VU�ȓF�L��A#�5z��)x���s��,�ʓyp,J0�����{W�;	)�B�I�Ba"�ش��3rYw�ݒ)�B��R��=���R�[Un��V�\��$G{��U���v��É�y�!�d�u�Iq�W72��%�c���!��Ǥ#PĶ��I_uV�H���?�!�A�JP*A�Yw�)ࡈF!�!�)n����u�@�Hb�� �J�w�!��G�r�E��8P�.�3�Z�z�!�dǞu�>�C���np����	�!�䇆I9ve[�ԅ#�ʜ��nõ�!�DV�dc0:�"@ _���c����\r!�Ău����g��?ᜑ!@�R�:!�� �!���ջo�(���'�<5���;�"O��K5f؟h�^%	�fƑm��!�"OX�!�A�{qX�ct�["T�fu+0"O$���ہ0���0�N֚��"O.�u��0��d��p���"O�X�#�G:m5��P�hJ�s*F�b�N�;}`����	�%���3�B���~�䁿i��0��4(��r���$J6�?��E8:7���� z�$]��.QaT볣OF�O���G�M��k�JY#$���d CgS���Hfvt��!lӠOQ>�KV"ȚeEP�#E�j4]Z"�,�d���(O��B�r�
�*�9�ք�S��ij�W��P�韞McҞ|�&c^�"���)U�z�ť^*�M�C��Z%��l�S�=T_�u����z�' ,��QґA� [i.��I/���A��Xh�'Va���CoY�v�f*��:��j���y�O�!r��m>1��c��j��t:t��h� ��Hӟ���I'CF�I�`��$>	2 �9wS8�JVʟM&@�0�ĂQ��{'�C/�?�t"�3{B(�����]2�+Z�&�pĊD�@?�5�a���c�ܴ��J�G�J�c?�l��&  �bt��(	�A!��q�&?�@�`�@��%�"�`� х�9�؍������0���OR�1�N�<V託���}bVAKMѺq�'��]�$yt,	�f����[�|�؝'Ɛd��&X>1d�ةcx������8ibZ�U�@7��2��N�O�M��� uxR���	(_��9��O�_�f=-�J�t�I�_��1��_�d9	��A���i��K2n�F����H�X����v�K~��~b�+�z01��y���a��
:ʼ�Q�S����'u�}%��|R�, +�B��T��*y�P�m���:�'�T�#��֝5#>�1֌ �{�VyY���#p�Έ�w�C�c�
6͘�/���0|B��Ѣe��xP�����q�e�Ħ9R��W~"��=a��ΑA#�l1�b����j|���'�,Z�iq���)�%A$		���@��T��1��d /�J��4I1�; �S<D~� q���9��ܐ$ �<e���H�t�<� ��'2���lѱ#28R /NY�<9&�=Nne�FFF1?�9����S�<��섶���R�n*6��C���W�<	u���n��d&�*/���v�]j�<AT�[�,�z�)1�, ����Ac�<a�N?9�<xb�\.+�i���D�<QЇ�2Z�qb�B�( mjL۴)�i�<1�U�y�NԘ�Eݠvx��7�Aj�<����&f8���c��q��u�h�<���1���.X.{g��Sa[H�<���L� ���@^fњG�@�<��K����6n�Ⴊ��9�!���D�~HP ��m�9�f�Q�!�ضB:Z�hr��ag�1!s�O�v�!��Կ.� �0&��\��3ƣ��OO!��w�� �kE >n��A�ݻ\!�Ę�i��ڔA_�p#Ե�� �	r0!�֛zݘ�R�LB�Q��B��ќR�!���^0��Q[�}���ʁ/*�!�D�Ukl2F��	� ���ϓ)!�DH"OH��H�냀�	cT6!�X�0q���L�-|p�q�b�"D!�͘D�~!AeɊXe��;�!�S�!��	t|2谐�G:j���hv.��'�!�߸.�t0s��;~���(sM�<'�!�͔DФu� B5��xIe,�7P!�W�%�X�`�J�Z��1 CL_7`!�d��X�e�-���k��0K!��)J�>H�a��^$�*�i_�A�!�d���!s5o�h�S����!��6!��z�e�saZ��ǧ?H�!�d�/�,="���C\xS7�Իo�!�DEq��X�&�Q'jL��` �l�!��� S�6x�)bHVH��P��!�� �@
!e �(��ㆵi3���v"O�|{ׁ]  ��!Yp@@9,�s"O�Ѓ6�a�L!�/��_��]�7"O�Y:��7^�&�iP.F'v� HJ�"O�[�C�<:|ِP͎�&�R��"O����P�Ph*7DW�Y��Ir�1D�xq����__:u
`�SI��k�-D���f�*H�VI��S�=�EKj+D� zb$X�m���(����Dt\=I�-+D����݊k4� ��Vx�`m#G�6D�
wc�E��"�eՋv��DB��5D�8� ��gs�3C�*U=P���)D����j�"?�`� p	3+�*�"Vj'D�dA�&ݩ><P[ .U��!�U+%D����E�tG6xR�z���dn0D���1%O"*]�؛���3�)���1D���E � :�(un��d�$��g@.D�Tz� �0R�2��U��LA�+)D�,�q�S��+\�ZL$�hC��X�<�w�P�`��@�c	���k�Z�<��&F ;�`��N~�<=�Qe�K�<���&88
�������#n�R�<qG��4"�"S���Nd���c�<�6K��4)�D�����=�L���Rd�<1$B�&耉��Ԫg.`,B�N�^�<���.�9bKmX�=S!�A�<1�b >J<��"�_p��rD˗}�<1���>P�t倥���8����q�<�͘�D\mHA-	\ptrW�@g�<) ���M��d	��G��` Aa�<�_�(�|���P���\1�%Rt�<�$�_!Q0#�D	�&NzD�	e�<q�^�Pn4�
���^�a��b�<)��ߠ)2��C
��v�8T��G�<1��Ƭ
������1(�^8�r�FF�<�r��/4��T@�.'
.v!����~�<�����i�S�s���aa�|�<y���!l����Lb5�`BLa�<	b��:�h��/
9?��)�d�XR�<��@� |�b$�,�E��d����P�<�qC��9�^��̒)"'���RE�<� X&��i� �j+� HD�^V�<aEE[	�a`��{ضQ�G�WT�<��d�4>�4@�jE7Ҷ�g�
F�<	b��`���t������b(h�<iW�E��D�"�"ӊ�� �d�<�G��l�d�i�N͈M�0Eg�^�<A�d��lZ�D� ��xA��,^�<i5iߎ]������6k"H��D~�<a��
*yN���2]�0%��N�O�<A�K{�\ԉ�͝$��YꑈAw�<�4O�)Lt�ɺu�,y�x���J�t�<��� KMٿX�J��FFk�<��K��4���!ֻ�60���Je�<��V����P��X�|T�'�_�<�G��4���x \� �SU�<��ǂr;�阣���=�]y�%�R�<�����9�1��+N[����bO�<I�A9S������R��`���f�<�R�N, {=3�f���unk�<�tFѦ8�ĳa��F�����~�<�W�n/�̰���/�ll	#�\Q�<Y��"m���f#I_G
|�e�T�<i#��&f��s/��(�0u3�`EO�<� \���⟉d�
�J���P�0I�"O�5���rO2=0U
ݓk���h"Oq���L[����?#��!�&*O ��E#�+���i#B��H���'HC����p	 �ꓳ�v�h�'U��ZW�A`�.Y�b�R�yH���'���b!��,JڑI�d��H�T��'� xcd.� $�Vuh��3t� �'��Q��έ7����*x ]�'W�h� ��� \7A�8>FH
�'�b��CD[줵����fUB
�'ҒXx㣘�;r3 i�3{���'�9��A�5�h�2柵q���h�'t�s��O&G�zm����#S����'o�������)��Pv�M�T8��'+b!�)KC��ҵL�I���'�@�cB�� [�J�zh�Fs�P��'xT�����	��RtIK�0A䘇�n�&<F��:skh��tO�,*[~��#IX�!"�y���fR�5a�ȓI��#�|��q�T��� \V`�ȓ8C<d��R?+ L��Ţf�$]���~y�vd@8�ȁ�	� G�:��ȓG54�uD	0�t03�x���ȓ�Ȑ;͔v>�lPF��9d���X���	�D��_n^�+�bN1
� ����t@�4��FLb��P��8M�bчȓx�� K��΍U ����/�1<��%�ȓ9zL(r��tztm�nB� �̈́ȓvG�E�r!�]f
�3f���"�n���q>�J��Z�p��5[�Ҫ,v"�ȓD�ң :e5<��wj'Q�`���P�"0�
֗:�.h�.̉,�a�ȓ�����N��T�t�  Cڅ ]��ȓ5'�"��?��jd�ê�p��ȓlU�C��_�@p���3��.h��e ��`6.��Q!�;�iÍn: �ȓ\㔼�	y��,q�5&�Z���5�uZA��?����f�0cr����qQrpYW	�*3ڼ�8��˫[��ȓ�^�h�]�z�d����&'_����,_L8�V�
v��I����W����>|T� �����h�O����̆ȓ|�F�{e(F�Y���9���A�\��ȓ.L�=�wJ^�ZБtLR�G�z��Ί4�l��6�w��?4�����fL���j�!\�堊�y	�e�ȓ[/��`�#wBФ8VKˎ*n�0��bޚ\P��;{���;�hǠ��b��=
  �	�0L��C0�%�ȓU�yAo���[w�Y>hʈ�ȓx��!��_v�1�'�"9T��CE�u1� J��P�umK�;�hІ� ���Vd��Ɣ*�jׁm�v`�ȓe�e��H̶R��]�O�T�ȓ��0"&�^�bo�}���R�-�l��%o�YA��{���[f�\�>�ƕ��|��܁_���H��-�0\䝆�&�:���E��=
�kC�
�A�%�ȓ:�������	���Q�􆘄ȓ4�%� FS�r ��_b@�\��-$�4�s`T�Z�b ����`���}�FI��#��r��9�UN�2����{�4���¾!`|x�&�2-��S�? ��bWk�8ע������UqA"OV��瞪;vDYrfˋj�lrc"O�� ���7d���T�)`��"OJ,꓇_�n	T�cGő5EE�Ĩ�"OV]ReW�?޶��RD*>A�@��"O��9����Ë�U�n�� "OF���OUs�d"ƢŤ-�j<{�"Of�㑅]98�����!D� X"O�eҁd�"E�8ɂd�@�Xx@"O�]"E߬c�$�Q䁍���"O�T�B�|��c��;�b�+�"OF�#��J�D������H-D���1"O���J�T!(�cƩ�	P��� "O�%ڑ�דg�y#�?^e� y!"O��S����d��� �NG����"O�qB7����@y�1,F?FP�`"O�QK��#;r����k�4�0h"O�aV�ŭz=fk1��<��W"O^8A���*)sV��s M�+�@�"OHZN��D�&�������6"Ot(V�O�]a�йE��2��@K�"Op��F�+d���� dY�'�����"O&�KC�X�X���ŅnoX�S"O���T���@X*��2���{�'c�Ȫ#�Cp��DꋴCb
���'b��!B�.C'�� �l�GTr,��'^�)�-ėyU�i��\�Ff�c�'Nu�$t3���F=�-��'��2�hB�ct�CP
:9�,`�'��4 �-FT������ni�'������p�	3�����q�'��%Iq�V뼔)�j�O�(�'�T	���>��1A\9�fX:�(2D���0�E�BDݡ�Ғ�b|q&D��p�B׿��9��N��U3Q�"D�S��   ��   O    r  n  +  a6  \A  �J  �S  Q\  h  Kr  �x    k�  ��  �  5�  w�  ��  ��  I�  ��  н  3�  v�  ��  ��  ��  T�  ��  ��  ��   �	 b _ Z  �& �, `.  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,͓�hO?�zP'���|��6E%V�ၖN'D��At��j��KC !sx��rh8D�@+�-�65b��@��B��`8D��S�;���!%�*��u���6򓑨�E�3#νw;@R$��Kv��U�'މ'<�m��.[&�9�BM�3�ڴ��'@�X1/�U��yk�H�+Y�8仈��?�S�T�ݚ���t��e/��� �(O��d��%۰��w��
K����d�ҢB�䛿�X⟢}�wi٪M,�Ad`�,M�<Xq��N�<I-�� �J��	f[p�Ё.D/����#�HOP��x0��0*��`�2准N��A�!8�O��hG��:�޽`�y�fC�<f���?��� �S��H�eB��B�2Q��!̟C��0E���3W\��"j^.ܤ�r�S���ĉ�t�f\:%m�8/���J�#��xb�Ob�>7M1?�cɓ�%��H��k�a���ç �\�<�2��*�L��(� �&�cg(^�<q��(4`�l\���`�e�Rx��Gx��
	N�`
a��j� ��5ㆳ��'^(�EyJ?�ІI͂X*q{ C�5,2@���'D�p���;a�h��A�&3d�ͩ3G2D����iZ27R�1��e�'����.D��(W�Ϩ��A!���(A4�IqE���`��	b}��K�kD��i��̠:�D���eգ�p=ٴ��C�:a�T�\*͂��D�CB����	�'��rF�U���j@	�[$�� �{��']�O�Oe�A��M�G�&��ӳ����'�ў�}� �0�FF'����k��W�L!��O~c�h�㉄�\���@��}2u#����k���'�a}Re�"~"��@K�J��A�W$bU����ɾ���m::MbGh �Szn�c�S�azR�D[�ux�%DYT zQBgeQ;aY!�d�>@��xt�[<0�a�I�u�����'����`F�;֢	*��E�ՂA,D���O\6���n��e��,rgJ?D��!#C��f\ک0��0JR�l��2$��SF�]"'�ZE��Y��)3cݨ�yↈ%O�BIzv�[J����ع�y�[�V�P1K�*B�%��5�&OO��y2m��p������]6 ����Eo��'+ўb>ّ0���%.E��)69MR��I6D����#�
T�^Mj��H��&���2D�p��(k�d�ree	�� 0� 3D�܈SB�#5s�#��G1sư�ٗ�2D�x,���Xf�p|�����I>����+�Yվ� 	��b�� oI*��B��+w��9�P.(�4��&p��b� E{J|:���J�i��!��/�r��W�<��]�V�L*SLU�.^-�T�S�<��E�E�̝
�B�/YY��()M�<�Ơ#q'~Pv˨V��H��
OH<���֑.�*ԀR�\U#&��S��%��{R��Y2�[g�R:�}j��	�>a{b�'(��R�k��'w[(�kÎ;) 2`���\1�cg] _�	@���3J/��G}�ŕj�O�� ���Y��A,^o�`k��d?O�4��O ,�ظO�"Z��h�u^��F{Zw5�O̔��"R�.((Ԩݭ4�93�"O�y�+�_���Z��ع"�!4T������9��xFz���7�����m� T����?��D֏&˖�G	ؐЮM�TNON�<qwo�;8T���l�O��ts��G�<a�y$��!U��#L��רM��y"�ށ)�J��K���W�Q��yBF��v��TIU)�1I_ ��!�3�?I	�'p����I�;��1�H^�d�L�+ÓJ���35�4#�SJ J(y�'O6D�8S�&O��d�$R� 	];��3?��)§8�����֫=eH��� Qf��|��&0&	#c�!j|�`��M��VV���hO�>�� &��A�D(%�"�i$"D��$�I�^�F����5�`<hu <D� �1���;�(��
Æjv���q�:D��	�j��o �H�� ��'`:4��l-D���@�7َ��4�ʒ��x�Nl�p��ɋ3����N�(W{� ��K"X���Dv�"o �A�D�[��F2F���[+yh<�c,A0 =���"���.��d�D�<Y�a%�!�ËYzպtZ7�Bx�<1��I<i�i�7@�����qx�|�'�\̀dW�E�����(�¸��'���C�]7`�r@�$�s��̓�'N�H�j�0
�fd)�kxTh��'u�s@M�4q�z���=n���'"LQh��/@�$�*ci	N y��'���)W��L�jS����W����D#�O,$��k�61��!����5@D0qr�'��D�E!�?`����%Ќ7.j�&#*D��Kr�&t��m�6!س�Z ���-D��F釋r-�XY����t�9t�%D�8R]jD�6h�@N� �	�$�0��)� 2����A ��)$)2+ �H�"O\3�ɕ�v��eqVH���;�"O���*I�N�,pڐHX�~� d�@"O���h@� w8��&�'���s�"O
	X�o�9�H����ڤ��'��Dy��)_�a�R��R��/&��a� ,,OТ<yu��2t�pie�J2+9�D�"�	X�<�O|(�G�T�]�<����LSGv�r��d`�<�>ͧO.�	�\qh-�G��~�@�a�6�j���'Ԝ��N6p���'�Ÿ}���{�\�4G{�'Y>\�ǫ�;�>p���6�@݇�#n�t��O;�A�$ь�6��=9�4�O�O��iQw�ό2���t.��4�I�'�����5Z�F�RD��4>!�PY��-O�9 !��i���)c�74a×"O�E��dƄ`��4¦�=r�ڴ*�"O�}p�ю#R�0E��i�J���"O�$��^�p��!�Ժq"H���"O�h��ЩNZ���a�/�֭�R"O�41W��)A���� �?b���z�"Ov8)��V(<M����F�!x��P��>	�$��	�׸>%|���R��p)��	Xy"m�.��ܚ��afN�z�$��y�Ǘ`
��ۂ��UK��˄K[��yr�	.��v�F�S�
YiA�2D�dC�������6��d�(�a�$D�DS���3?^lm�E-]TƐ,C@$D�,��/IVy��Kچ��3��"D���f�P+o���eM��o��<�%;D�l��[�+��A �S>��S�+#D��h׬'�J܀pi,IE����5D��0�F��A	�ϰ���7�2D�@a$̒�(Q��`�*��f����h,D�hg#�ʞ��G��N��k��*D��4Lܢ@̢-25��Eeʸ�s�&D��7-�9]䠸q'CX& �0�DA%D��૆#a�RD	���>]�V@y!"D�`����<x�ajw�W�8-�p�m>D��1��N�x��v�փ;7ꔱ(;D�d:��ڮCU�AB㇖g��<�Ҡ9D�(�UJ�1 Hp���3��#� 9D�l��'ȤP�~�!a�S�q!����9D���ϰW��()V�����r�8D��q�ŀ8���bm�	�*��c�*D�y֪��@�Y�a�I!5�2Qivf'D��P�c�|���Z&R�N�/%D���Ʀ
�@:����@�1Mbd%yF*Op���݁�8 ��]���0��"O�I��ī.�>-ȗ!��6�$YK�"O�� �O�,G ��U�]���K�"OFaa˚+"�
V�[zte��*O$�ʢ���Z���L��I�A�'vtH�AU0U��Th�� 5,cl���'�-�t�%o�~�@Q.�l���'�J��h!1N�Y���!N��S�'R�kW�̣n��(Z��O#}eJEp�'M<ƕ�B��ƛ�E���'� %u�%}"i`�Z<�"t�	�'΀� QHU8�U�4�8�	�'��TBЋA$D�
QJ$E� (�����'l=
��?N��\
$g�'�nԓ�'���Q��X-�:�`@-\��R�'n��� �1Q:���C�-n$59�'#�-C$J0_�d��2�_��d
��� �Xʆ�D�L�"-�D�q��,��? \�
�'I-0$!!ATvńȓOHX��F���n��X����Fώ��"@@���	��`K�=Ilv���c�nY��� v>�X&�Q�@����ןt�I�0�I�h�Iϟ��	ԟ���{��` ��
4xJi!VK�s����ǟ��	֟����� �	ǟ��I��	��>�s��� f�8ԀP����I�����۟�����������ӟ�	5Yg<�k�FE��r ����+�d �I쟰���<��۟��	ӟ��ߟ�	�6�!��;((�2������<�IʟD�	�������������Iǟ��Ɂ&Ⱦ|��X6{=���B��<~����ҟ��I�	��������I�����:V<���A�tV�2�J�1�F���П��	�����џl�Iʟ ��şX���	�F 3B
�1t�8�Q�|�%�	�X������	����I蟬������ɱ,:�SD��U?(yr�,_!������X�	�4��ӟ���������d���i����#AqB^��^�f�����$�	Ɵ��	�����ПT�	ݟ��	;0ӈ�8g�[ht̤��$�*鸩����������I����ܟ|�	ҟ��	+�TԚ��+�`�Aq��|�����$�Iٟ$���������������	�����*�#H����4��iʑ�����IßL������I̟$��4�?)��<$d,K�@�-�t�(�E�T��i�UR�L�	Wy���O$�m,keH���A�(R�B��7���|��f�$?I�i9�O�9O��d�0K�~����>6\�P�L�=9��D�O���wGt�����ԡ�(�O[l��F���9��r�*�=6��y�y��'�IA�O�(' |�d���_�.���1Phh���8�D6�S��M�;J��LY����"�h�ئ&>I\^أ���?��'h�)�S�pR}l��<��b��RJ̩���#c���5
Q�<I�'<�D�/�hO��O���Fhŗ�8��G�k���(U5OTʓ���FD���'Č�a�5�@���H̘J~*hjR��NJ}��'��9OV�Ũ
T,�}��ͨ`�.��<�'�bR�>��1��d+ן�1g�'$$~�ؤ�3�Ig.��2k��i%�ly"�����dT"�V��p�����F�5H��Sʦ��Q�7?Q�i��O�	�� ���'/�h����+��D�O��O��I7�m�*������ �k�mV*�.	x�@�0��`j5����4���D�O^���O�$N;'�A �R%ԕ;�\<�L�Sg�&�R��B�'�r���'�n}��(\V�%����)��yj�o�>�ݦi��d�)�Ӟ=����Q p j��!��U�|�<�"���S�O�y�N>�+ODP
pj�D褥�2fA'h�.Hz��'=�7���L��k}� U�A�e躁�!+΢����XϦ�?iP�t�I�����J���֩ߟJN5�ȕ%N�rplA~�4WX��ӭ69�O� G;&ȴyV�O�DT���,˓�y��'���'�r�'���Ƀ7|��P*�bt�	`��1"q4���O�Ҧ]a.�i��'|�yB�߆�x �rC��1|Zp:�|r�'��O��a�������<<���
Y�U�ѪG9IPT������V�&��\�������O
���O|�Ĉ,{ �����r���2K�-f�.5G��O�����=��'	�O}W�����i�D�0kӀ��j�y��'b
듥?)��O�2'3�z)�`��AnݔBA����L�:��=x�U� �Ӥ2t��D�	 |x^��f�SI� <�4&V#q�\�I���I���)r��?��Ė���@��"2%ɗ�]�Y��8Rk�/�<�'[(7m�O|��?�0[�����y,����*���`��a�t�Iԟ�
q�Tڦ���?!-V~�i��$S�t�.�`⌢a��r�#W�Ģ<����?A���?���?Y.�:H6i�"٨I�&O�kL��n֦MH������	��D$?�I��Mϻf)���&T:l-��:p���j��?AI>�|�uG�8u��Qϓ-X�xW�''ux�l��o֤��w�pB��O��N>	*O�S.pTEҕ[,(�1�r��[�F�����E������	���� ��e��'�qڂ|�v�C����ş���R�	�n�B,[�GM2|�T��snB~`��e����Z�ԈL~��I�O��R�|ٰ�P��>u��p�(R����?���?����h���ĞR���%�{~X��#d#Q6���ݦ%y���ky�OlӺ���E��]��,˷�����l��t�f��ş|�Iݟ<��f��E�*�:��Mj����L���_�R6��TE�v�<ة���
������D*�MK@kL��jB�ʍS���M��D@�?q���?���D.O�r��8�V�ǵ�k��9t���?i���S�'_����K�?P_�����8��0�M��^�옴��W{�$4��<�𠝠B0�XC��D	q���u�S7�?����?I��?�'���_�QZ���ş�*���&9�r(�f
]A���bhW�|r�4��'����?��Ӽ3��.�Bb`��>P��m���0E+|t�b.{~b���a����ӪBD�O�� : ��]�8A�N�oX&%��:O.�D�OF�d�O����O�?e�+0��H[�zCfMZ�C��X�����ݴY�l�,O��o�n�c8���!��,���s��H6�$���	����K���jP�&?�a�D�j� C*��Tn�����E'Y���1�/�O�YCM>9,O���O��$�O�� Ƅ�LU�!9%� �j5�7G�OD�ķ<t�i�hj�'���'�哚(ϫ��*P���R�:xbE*�O&��'��'rɧ��,0�tt�@�	���Q#�&ѯ?q���2	�)kn�Z��	S��~�� 87��
� �zZ.�(V�L!�v��	����	ןx�)��CyRCgӊː�B��P��*\1q�*��q�ѭ#�(�r�����]q}��'�l��߀k�č��\�{�j��a�O@�D�y?�1������0nW;1��ԟ~��� ��1�A� �l�Q����<))O��OZ��O����O>�'�Ƅ8QOѡ6B p�tiI�.��` �i�Q3�V�D�	L�S�P9���;#��7&�H����w	��jތ�?a���S�'��M��j��<Y�'m���E'X
d�Ѧ���<نa�>X,�מ����4�B�DN�|�&xr��Z�3�������I��$�OZ���O0ʓԛ�/ȔU���'D��]�\D^Aq׮ �N�ks%=r�'�R*�>!���?9L>)7}����D�7��`pA���<���4J��S�
�j-O���ø�?y��O%0��
5��k�n�ia�\:�"Od���ծF7�,˄�_,}F� ����O4�oZ6�r��	ܟ�2�4���yGd�C` LY��؃W��iF����y�'H��'[&���i��ɂ" ��a�ޟ,! �= �Z&J�S�J�a5
)�d�<I��?!��?���?I���Z�h�Y��_�=�t���9���-"D�X��t�I�(%?�I�UÔ�H��اIy��u�Ԕx��1��O����O��O1�t��� �$$��{�#��j�j�!i����9Ҕ�ЪQA��a-���s�	Syr�
?O�^,�΁7Ƕ�����0>��i�z}�$�'DTcWB�	&Ď��el��7b����' �6�8�I
����O��D�O�t�v����y����d2:A
��5b3H7�<?�)�8����s���-`�^�Ҕ:�d2 9jՓ�s���	�|�	��p�Iџ�&?���n���B�ys��$=�p��oI��)�<^���O!m��"��'��6��OZʓ	5�UJ�*� B6�Xe.�d���<Y��?��X.2q0�4�y��'j�4��[����ѢI�k{���^�x8�I*d�'��IY��.�EzRfE�W������hlHGxr.h�b�i�O0�d�O��'l���P�g�
�����Jm����'���?����S��_�yv�Ö��
p��aA�e݆S������֔Bq*�H$[�據[T�"�~��)(��\��J��pI�P�L-!����<��ɟd�)��]yIc��U0�-��!4i{PF�.�p�R�Lؤʓb���ćW}��'���Kߖ�xQ�"ˤ]�"^����	�5+́�2I:?���͋t��)3�4c�Id �Mtu�ȱE�:�y"P����ԟ���̟ ��џȔO���юB�^��a��DX"4`�D�pӪ�«�O����Op����d�ɦ�]�N����G&;����!����H��?�L>�|�6 �; `͓Oظ%��}��Y�Od�H�C��y�	n�`Q[CI�(N�T��NU�\_f%�E��?(�$i�O�U���taX���O��Wy�=��䑆z$�Wלe����g#�:�M鵄ZX6��Dy"��
,�
 �`�1M�� �ţD����˵~�<����W��R��G	�K7MP/ V���Дo����*z��#�Ȼ.�:�T�Z9Q|d��n*d�hlJ1)ܢ�@E���4F�>��6
š��}Z׍Q/}$��˷�ǥ	�x�RE)�]� -Q�r�R:@b�d� A���6��q�Ĩ��<<\9�!-v����OU�tBA&n���Ȣ1�Ĳm�Φ-�	|y��'���'WB�ZsT>�cu�UРZ����k]��7�Ҧu�	��'f��#��~����?q�'e���S�I]�B�
���֛H��ʄ�xR�'2"ˎ�E��O4�&,/δ���I�i��|�b�*Ɣ7ͥ<agL�'kP�&�'*��'D��a�>�1x~��1�	a|y�ք�6EO��n����I�(�:X�?����ɏ3x�#�-�>%�P&��+�M;��F�����'-��'�����>A)O��%藊zr�x��M]ql�A%����	�u�ߟ&�������7�(��B]��4k���Y���'U��'E���G�>�*O������D�q����q�wl���	|��Oi���x�������蟔)���;q���F�6%�hS%(��M{��W�Z���V�Ĕ'.��|ZcU��#T��K�X��a	7D҅H�O`|�$�O��$�O�˓`	�q��I�3A.l�"��h~���[7N_��Ny��'��'���'*����͞�Jzv��'�ߛBhQ�T��9�BQ���I��IEy#G
Kv�-aT���(�_����f@:~l7��<������?���,H��'���3'OǕ}���C�}�d@ȯO���O��$�<�c��V��Sş�3�!�A�`x���&^���`ߛ�Ms�����?y�||F�"����	_T����!Vt$��߽|�"7��O���<��!�/^��ԟ����?�A�	�&��QݱJ�K.�%���ݟ��ẘ���d��^�j�!�
�p��Ӆ��MK-O��Z�KHߦ�������T�姀 $Ii`�ƇwW��c$�	#pI6��A�i��'���'���$�|n�:�=�U�H�!,�i���:Q�B6m�	-�m@����L����|���ŗ]��b`J���L�@	ǝ���'}��'�R�L��y��'U� �T�؀sF��۳�"L �	�n�X���O����
 ��%��S՟��Ic�(���_�`���cWI��!�&3�4�?A����Y��V>Q��M�C*U"S�&Ip��Y+]*Dڰ�M���ɠ8^=�'w�'��'�AH�Ç�ʈ�hM�:!1��%I�1Ox�$�<��7]�HIV
Y�[�vqr(U�}��K�����O��=�	�����j�>l�A�	@��IցQ��ȹm8R����?!���?�*O(��R�A�|�'Ɨ&4�|�[2��8+�补�Z}��'m2�',�	�ORI�|��9����R���˴�ڠ.-���?����?a)O촲A�KU���vb�J@U�Q�\`��V-c�	ڴ�?�J>*O���O0�O��[��4LN���ɐ�_�2��4�?�����$,��&>��I�?ט��^�i3��p���阯 �@6M�<���?q���?�L~��CU`+[����J�1[+ԝ�æ��'�ڌS��tӨ1�O���O�N�S�0�I���*b���y�Fؼ �@nZƟ��	�����ɭ<.�����F�����냱*�^����8�M{𮛟�?���?q����(O��F0F!#֦�%� �#b���4���#�O�����)�'sĄ��T��_c6؁���!a,P�f�i�R�'<"E@�*��)�H�(	գ�B|:��e�� 1�ZIF-�O�4'>�������	�j�`�BA�"[6� �C"��,�ܴ�?�Vˁ&a���4�'��S��BA�����9+D-�4ߦ�M)O���<	���?�����dǬ�N��U�8c��ixU`G�"t�҃��|�IΟ�	S�	NyZwA(8"j�&E�1p�\��Ԃڴ�?�M>I������OzAW��?}��Cְ �:�B��n�(��j�H��O����	qy����M��N�� Șb�9 ^���ZL}��'B�'��	� .�:����d��T��N�a&�t�� Gw���l�؟d�'8��'cr)��y��>�v��&Bʰ�g��#9�4�S�����	����'%�}2D-�~
���?��'��x���rB<\0�K�&Aᰠ)�Z����ɟ�	�L�X�	����'����4+>�quB�FVd�������vU�(�o��M����?y��r�[��7e��E��	R�R �pd��B'�6�O2��A�{��DT��'�q��|��#�I��0s!�΍E��TI�icD!1�ct����O��d퟊��'�剂�HC�*��dxd��Ei�>�b$�ܴ5��̓��$�O��?��� e�����ެ-(� ��ċ�"�(#ܴ�?����?Q��M���ly��'!�Ā�4>QSC
ʌWvy*��B�����'k�	�Z}��)���?q�OJb�X�r�Ǟ���{B �9{u���'�����>�/O��$�<����5	�2�4�p�ǘ�uE�R#Z��50�	ݟ�Iܟ���Z��'��hK�1}�N�X�H�����0��%d����D�O��?����?�E��-�\p�P/��;c�@Ã�٧%9����?����?���?�(O�m�i��|����tBH�dK"����ԎZǦՕ':T�������I"0��牝���Cb�0�-���J�`z�� ش�?���?����Dڝ>�F��O>"I#�$;P.�.A猬Hv���4]�7-�O���?���?IG���<�/OB= ��� ~����!���R���������'�R��t�~���?�������dT�6P�\s�]��<8�Z���I؟���%wQ���'?�DP�r�@<f����� Z)t�L�n�Hy�ċ�L7��OV���O2��Pi}Zw��I(,��j��U�Ks(`s�4�?��Ԩ�ϓ�?!(OF�>iQ���v�ht���8(�X!�&g��x��ͦI�I������?ᣩO��!p�*� �7���cW�w�2��im8���'c�^��b� 
�{��0~�r!� �s�h��p�i�B�'�rX>�H�����O��	�-�t�U
+#&�slӱG�D6��O˓W����S�d�'�b�'��k��*_ ^ �6J�`�0uGb���ٶD$�,�I(%���&�����P+JD񭏧0+*�M�ĸ�<���?9����V�H�b�+߈CQr�f*H&S��ࠏ�j��?i.Op��O��df$|�C� 	Sg�H��k_�;�օP�b�O��?���?)(O���co��|�a��}8��]>�n��c*�B}��'�b�|��'�B�_�~�dH�Y}6T)A#�?s �6)˷(��ꓘ?a��?A-O80ɷ`A�S�a<�7�6c8���9�-�ߴ�?�K>Q��?�"+�<	J��R�[*nCX\���֩=�N�BB�oӊ�D�O�ʓ|j�q�Н���'��T�[�O.�!3F��p�P�V%��2b�xb�'�"�O��>=����e�"Ll��5;�6M�<	3���6ʪ~����g��P��Z�,H��B�*���bW�mӢ���O�$o�D"�D%�S���5�u�ЦZ�D�3̛ R�6M��%�Bn�����՟(�S��ē�?Y�N�6w4<�i��i��sƬW;)��V�_��yB�|����O������	p-�@��JԾj~z!��馩��ן��I�89:�}��'��� ��%���X�29X5	��%��ٛ�i��'Q,��$�/��O��D�Oh�xW���K$%B�ZF`]&*�ڦ�	Iئ�3M<1���?�O>��2�d�Я*gMMBdJ��O�D��'��%s��'���������'�l�9���69&��Vnc|�̙ԁ@
d�O����O�O����OX���_����&TP@�Qo܀��d�<��?�����@
4� �'n�����A2�X����}2�$����e�I럈�'w}��ɣ?���&��/Ԇ�҂oǱ;M�ۨO0���O���<����+Y�O��y��A� 7F���GB�[����}����*�$�O������J��<}P$>� @M�6wU��0� ϟ�Mk���?�.O��,�$>��	�?�%�*O��*�],�i;2���ē�?���c��[������EG�J���L,�q���\�Mc*O�,�O�Ϧ�Ю�V�d�4��'Wj ��Q���P�� ;r��4�?���>��i������O��\�#�L!q�^T����kc
"�4T���y�i���'��O��c�D��Z t>̈2һP�xP6!��MK����?QO>���'4�IJqIQ7!��bԊ��ujΔp�d�l���OX�DF�4��>���~�b�n?��y��\@l,�چό�M�K>�T�Җ5�O\��'t��Y#�Ӌ�,)�Όp���K�$6M�OJ�q7�
Y�i>�Gy��rM����Q������?Y(O����O��D�<A�'�1C��U���O�(9����T�*s3�x��'dў��hHXu!REZ�7�,e��H�4x5��o�埔�'K��'�B�'�"�K�����uB|��6�R�<�Z����Dݛ��'���'A�'��Q�!�t������;>��1"�,�l)At]�����X�IbyB�V�F,��b5��Ĝ��S��I�$�X�j1G��	ٟ4�?qf�O�'d(<(r�b��&Z؄����!$�o���X�I۟����$1Pp������I�����Epm[ x�J��ќ8>ܱ�M<����d�����!Dc6$э�z�&ZEFW�)�N��?s&���?���?��������d�J�hrh�S��)sաQ�M�����Fqr����e+F�Ә�b*k02y�f�iе�5z�����O��$���L'�\�	,[s��`-ƫ �:�UnB�d�����?Q�,��p���������J��`��&�'��'� 䊓C7�	�����q>��ǪGE�Q��EA�>��Ն������x��g"$,Xl�!͑�#enѺF��Mc��Y%�=2E�x��'�R�|Zcy�0kd���w�.p	S�_M
@��O�쒦�$�O,���O��"��(&��A�T!��"����J����'-��'-�',��'�BH�QAؑ4%�$[�AĘh�F@rt�L+��']��cׁ,�2�HCӮ;iv��'��b4�	�ݔ<f�0e�!2�:Q�ɲ	)�щ!��~<��@��>:gp:�%��O.�5hʢx1\� "8��ǮUX�*
n�C���X�a9��G�/��\a�a�;z��0(ի�*}�(���_���B&Ԯ2ݜ���'2�9P%����]��J�<$ |K��П{H
՛Ђ�=�L��2��{�ʌȴ�� �]A��V/��y�/΍B١�ҙaK�MS��M����G��� t,��h�!�	?(�|}�e��+oY�����Ρ�D���ϟ�rdCԢi����SKM���)j�E��?�Oc$۴�J�,��v�Ե%ݶ�H�̲`�[�\kd�
��@�R�
��eǋ#����M?��W P&,$���¯�p|Q�!}2ə��?i��h������0�p��%�5S,4a*b��,!�D� X�r5�t͟	2d�8�GaxbD>�74�q�%nU� {�<��C�?�D{C[�X��䟬�����T���ID��ޟ��=,�J� 楎�GG�U�7EȲS��e�W?��(6D![��>�3��ם$��4�H��FĹS_�[q�EH#�Ř��$���d���L>	�/�' ��E�a�]�4Shq`����?��O������d�I#s�:A�� ֽ5�d���w�C�	�{�0�sc���I����!���P� l���'��D�/4���$�T>
��}k���E#
<���,2j���O����O���;�?i�����B(�8�P�*N�aS�H(��(hw���?�Nm��2lO.��6�]��*؃ 'g�ŋ���*z��
pl��.����!T�8�E��3��+���L�-HD�O.�d,ړ��'9�e��C	9kV%3!��x3z�K�'xT�䍀!�1�'�� ��y�ȥ>!(O��v�k}"�'��3�ju-b�{G ��tW4����'�R�ńwr�'��i�O���y��?R&�-��2��#ElQ�G��d�T9���	%r��}C����C���'�lx�E�ߝM4���a
�'c{XU�
�|t6M�	�$�'"jmS��&+v}�d�[�Љ�y��'��H�mT�U�`m8u�TV�>���'^z7-fJ-��B�8�\�Z!+8i��<�5@
+`�Iꟼ�O������G\6�t��c�~a k%͂�i�b�'-6DA��ݪF����	_}*���'2u�W�Z(.$��K�Ʉ�B,X��O�zbI�02S@�z�π 6����	O�$4{G����LsQ�>QƎ���h�IJ�O�I;+iڵ�#燵�)��[�y���#�X31�����/�0<�鉾�L*�D��(������Y���ҭOT���O�p9�DM�����O ���O�n�3)`&�j�i�3�H�.� v4��@������c�t�XA'�3��'���7�ݘO��`�
M���ٲ�_, ]��=y�!�W��|"�y����0��dL�!���m��7Mwy�!�?�'����DL`p�9�nD}*��"���yRT=��Q$�� Mi��	��D��'E*���D�*�$S��k3�q�$ۢ����`��i
���O��D�OF �;�?�������h�|ՈQ�˿E������?!(L�E+ڔ�l4r(Ô�0=��G/GҺq��KQ�HU�d�i�W$�Xs�kX�����CCk�����2cG���V�G�b<��F$kW��D�x�4��'�b?���'..���l����pk�E,D��8�K�}�R�ېBҳNh�d�0�	����<aaO��c�&�'B+_{~\Đ�ɦH��"d`�����'����4�'�:��x�D�'��'�*Y�cN�y5l�3�
9}���>E�?٥.��scFd��\�:@=�%�m8��9���O(�Of�`�A�9�4a�'�Z+M�I��"O�t)d�J%J ��K��׳i>a�O�n�?"�~���N�9+F8���yX>b�t2O�*�M���?�.��y���O������"�R4�7!�T��#��O��$��Mz�D1�|�'�@p@�D/Vq\4)P�C�a~"��O���&8�S�'-f���u#��)}>)�"�W����>}�g�"�?��y����$Ĩ�����L_yc�,W��y�ћ�F���=Hܢ�Y�
X��0<���ɗdT�	0H�#t��PΗ�6�BxA�4�?9��?ф�U�?I֩����?��?ͻ7�%�ӎ��M����0NгW_Z�q�yB�ݨ��<����q��ڡd#D���Cց�_ܓz&���I� W*}�##�]��e`�b�T�<!%����L>1��A<�1qcLVZ�HE�R�<�A��&>�L��"��`8���E~Ҫ!�S�O���`�fӖ%��	00<�PԠ��L4�Z��'R�'��Fsݑ��ǟ�'1o&E�tk�%BH�����;��ǫ_m<����n�p�)���7���k��J�q��!��m�pH*�!��v�� i�$,�<� n�埌��	 +�zQ���6n~̠sPI��LX�B�I�*�XՄϰit����11�db��}r� �,�7��O\�� K��	hqn�*�Z�B�
�34�$�O�1e��O��D>���ON�O����I�68̽�'�����&�'�P�b�X!�d�8�-A7G�ʨ ���-�p<�a���$&����5�X8r�78�e��h5D��[D"�/��|`t � 'J�1�>�H�۴>�8L!�ϏPѮ-)L�/p3nM�<�`蓮p2�f�'�Y>�d�ݟ�auF��)i�H�Łˍ@��T�KUߟ��� xs`L�	e�S��O���G�K�,��D�h����>a��EP���O^�-�B#M=d���b(D��9��ɳ=_��:�)���M�"$������X`��ʽ4<B�	��h%�'���H؂��S���F������B�'�.u@�K��(�1��h߬L���̲>q��?�0�)E��!����?Q���?�; @��˜9�F�FJL�4@Rb�E&y�I��Nk��xa@�U?��|b%U56�Pia�&�4�Z�22W�N9��+�,.�l�e4xQ����|r��9Y6�t�w�D�w�p��H�)�"����W�O�i�O��P�t!Łp|K&)�JdQs-D� ��F#h�H8��MѦP����`*?���)
-O�Q��Z3<�P��@]]��}j�A@:2�1yd-�O����O$������?1�O��x�wąB����&�ط ־�c� ʛ�x�ɞdc��c5 @�d�)���eS��k�'d��[B�͉+tS�	A/3�2����¢�?�
�@�����cH@�Hb@͆ �@Ņ�k4�0���4=�����P�y%��<Y`�K�4��'���"Y�.�2fE�D<�m��8"�'#D�S��'�R6��i���I&���Q"��ē���i�zTYu$[�x�*<
�Z,�p<qc#�Z�����
�X�dʣ@���I� ��R]�*R�-b���C<R�'z�)� b� P
h��snÌT��X����O����(��A��&p�P��M͡q�!�AצIDEF$y���c�Z�z'��� oo� �'q���Q�c�2�d�OB�'j����A��]h��&*�쉩�+G��TA���?!�/���?y�y*����[��$��GG���`x�aH-<��'n������)�� ��4�S=!/j$80�;;�yF^���H�S�'TG�Ի�I>TZT��0���ȓ6�dn��~�<�׷x�l��	��HO��ť��0(����r^��p+N����П��I${���hC�Ο<����i���,�*G�d�3f�^	,Tt8��@̓5���$�O~D��Ll�<PQ�eɚt�qO.,I	�	W~�hG�e��� �֪�������ҭUm����?��9��G��"����l��y��'�D��p�����ɂ"� Z���OʸDzʟVʓA�|��ԇ��a����*0�̥J4��\��	���?����?�ķ����O��)4^\"Cɢȴ��s�A�`�c)�@[�a�`FС���y�4�Y�i�a��B�	b��'�E�ʝ��ӣA�����h�O����J�8�
�`B�AvTԈ'HȹC}!�D�66@r��ղSU�Ȃ��z1OM�>y��^�B���Ο@1�I�.�84��.˹"�ބsd΋ş��I�y���I���ͧ����'��R��ώs�R��VMW:H��Q)M�:H���#�p<�У'��h���I2P�����k;00h�Ԧ~S|���&@� W���D�|?A������d�0%��(K�_��x�6�V�X]1O����dA~�9��_�H��Y@�D(W!��j�DK.8��з�z��[�\9�ĵ<D���o����'�b[>9�$�՟X��bʻj��Ā�!�kҠ(aT$�Ɵ<�I	o��uK�R�S��O�y�f��3C$t[��ȠW�����>��!I�w���?�
���o:���f�
0��� "}���<�?����䧔�'?]�SU�IZֹS��(q�<1����<���J���F`W��`��$+]}� ȏ�Ø��X�5�N*4�*1r� �V�:��'��'IXiyG��ND"�'����y瀈�O�����gٍ|��U:�_-z`D��6+S$y6\Y�D�^�v$m���i�~�dC�fߨ��$d���7Ā@��j�)����K�N�����y'��f�D
%��})�(D%Yx4CR�E(���*?Q��Hß�q�'^��i��)�|���ĩ$��0�'���Apˈ�����q��f�����O�Dzʟ˓S�n�+Q���"4�Eo�06z�)
A�,>�v�p���?����?!A�����O��Ӕ5�$��`�@�>m0 ��O��t@�
O`��$�U���q�F� 4Ҩ�r`f��PxR���xZmR+N�	td��4B�*pJ����?�H>������~�e��4�M'k��-PЊ�N�F�<�ਜ਼
(:��3Z-&�!��|̓%��IIyb�PZI�7-�O��ّ@�ʽ�$2D����W,����OR ����O�$}>�aV��O��O��p�kz4�W���3�TW	q8��e�-�I!�X���g��2R�(ԺN���G�1��|���t�l���
�	��yr�N�>�b0��sK�#`N���x�q�H�ZbZO7��	���$��(w��E�*���'�bV>y��^꟰q�IW�PR�(4#ڊT:D�[؟��I�c\|I�f�:�hapԭZ��?�O哋!�VtPE���]�So�D$��'u���ES3����2��Xv�>���S�9�86	�mJ*@dk$}�?Y��i�l#}"�'CAB����F�J��`9橛b����'�v���	�Ԥ�E�6b����������ķA\26�����:~��F�'i��';be���@��B�'x��'��#,��Y[�߷[�t���'�4�<��~x��ST��&2����&j�t����1�ɛb����_(c��IP'*T�J��D���w��c���D�Oq��'K�a�1JJ6z*f�0w*�Z�ȸ�'^Z"&נz�����-�i0�O@�Ez���Ƽm����"�Ch�Ia�A�&e�D� J:B-
���O�lZ؟ ����a>U�Sm��rҔ�"�J9=C��2A�Hu��2�O��+��0
��(!U� \l��0\lE���(�h#t�('� ܰ�m�ş��IΟ���ay��')�O� F��� ^?UN��4]�Y��@�"O�S�D�	3�i�F�i��AAA�~}W��[��ÿ�Ms���? �Bj�9�����`��q��鞵�?!��9jt�R���?�OSH������B(<�y����P�$�Kv#�PH���	�-���H�ViB��tE�����A�K,Ot��U�'n�'�z��A$� �N-
G䀖��Y
�':az��[�9���6���>��	�'��6-�{�������#
��Th��)�1O�I��E�	�I�� �OH�4�'"�ܚ�b�#9���`X�P����'ObI��mi�T>�O����c�'=�L+�jٶ7]F��OF���)��3 �`�����U�8mvB���&�'��q������O�:�Zg����=��o�SRF�'�6���E�~�����I��<��HiÓё�� ��3��� b�P�h8#�,D��!���_�z�8cՈx��S�0D���"�[���Qoئ�rUz<D���%6-o m��LL �J��-;D�겎M�[�\�#U�y� LӇ#$D�tٴ�R�#�)S�Q�U@���#D�4#׍ȻA.ni(�@�4 �����L D�\"g�ř6l�����ƠL�-(�G>D��Y�gG0��$B@_�l�����0D��*��v$�3r�^�.��� w�/D������O��Ix�5Kn�kWJ,D��K@a�"c}~��V�9)jD*�d)D���A���|3"�8I�b�xi'D�`C�G݌[GL�i�HU�
�L|�t%D�0����	u�J�ؐ���f�H��M(D��rk�&��yp�Z�h�@��&D�tTB�rGء@ę�IR~���#D��
�.k��u���$�|$�a
!D�p"�l�$:φ��Ud��!l�t�c�?D�$3���4L�H�
�b�l�8q�>D�Dy'��#�X�^���awm2D�\����A�*�W!��'"�iR�*D��'ͩuŞ��ӈ�l�ֈ2��%D�H����z���2�ْ@�h�*)D���v �0i��B⍖�1�Rjr�'D��+5�sĞ�@V5&="a0�8D��5�K�L���=3߮�P�6D�T�R�ĪTe����Q��@Y��6D�0��f��)��	��ʑ�@98	�c-4��A���#������'���$�<m�:�B��Z�D�00�I��<��C$[�D8E�#ct|��,�\�'Pz�����E��B��rx�!9�O$,XP
f�������?�W��W.�:<8�Ņ�#y�i ��OmDr��§ӣ3�\i8��'�B�8�!�I�z���B�(>��� ���%�)�'y`�}B"�µE��%����f}4ݐN�d�ax�'�-LTp4����	�3��|�Q��в;6N�I��?}�`GA�'��%q�G�Q�0LkG�
�"~��9�FǗl��q�P�$�,\$U�4�j,����@;]���<�TD��N#,���H?r��!ȡ@�v�'Z6S`��(K?0=և�:�r)�'�B�x�H�/���3�28�P���'ԮG
Ġ��9}3\!���O����OW���+��NbDɜj���y�^=��h���h�rAO�g��E}��eh�a�Ft��iZ�a� #!���6�(O�>�kT���`V��	%U������zHb�1!L�8���4�J1�r_ɼ�B�L>X۴%�D�V�N80�F��@=��=�ÆܪcfB���-a�������'��T[F��G<� �DE�w����I� 	���{J�|8a�ڥJ�\�3��*<O�}:e�ʅ
9\�1���0Hhd�ՠ­(���ȇ�"k: ��ɭ>�3Vtl[�	���2�hT�Ft�'�BY��/� u��#�ʒ��<T)��D��j�����O����{���*GnR�b'�*O��I0A��3X��p��OT���|�9K0C'	� ���U�$ք�6/��D�tp�� �	/�\tiD��օ�2'e�=�iX�:
`�VF�V Ś4a2��!eN�*��B�]�* ����P����2mH(����O�;2T��q b�ɱm*?q��ȴ(b��īK�*1�Ą�Wy"����'��$�/�i`��;LĦ� ���R)1���i�I�o���q#�I	o�1���v��Ba:w�ax���N�����)Z�O� " g����I��?@�6)+�����G6�>��JqΕ}j��R�+�:A/����@�Tg�}�Hc�7��UE:�`9Lp���13*ISQ��@��� �?��?��?q���>��������ѐ���	��b���'��`��dD��Sm�K�`,¢��E�8c�h#�O�����F�=�,ԁ� �O��'@���gAy���ip,V�9�^�9�'Zɹ��FGbԛW��C������%���k@��<�l�S��*�SV��F�h���F!11>���(O��Ҁ1�pm���ӑ$�:p�%
)��'\h��G�������R��=���ȆG�:�bh�C�/;R���'�p�Ey���)޼��?��,H��;n
L�3G��y��]���ޢ\a����O�
M�7O��S��&l��!
�����`&��Y�$ߥ��	�O��Ez� Ҟy�zIإ
)Y�8��D��'�����EQ�}s���C62-���?�I��9RP��X0:@�"�̃f�����*���D|�4nB�=jңX,D��[��7�Xi�� P�
sFX�1���8W����Qìp焴��w-�O�h�cL8Z�)����:?-�(2��H���'
L! Va�]`h�x���v�C�b��d�[�A*V�V+"F��1� ֹȖp��0�I/$�8��?���$`R B�W	6T$�*�$�=��M "�4�z�b���7M;�'�xaÖ条g켪���$J�� U�,���u��˟L��Rkoy����a�\ m���f� �Dy��K�Q���~��+�>Q����_�iB@h�0�[�m�F�~р���O�)�@���l>x� ��u����aM]ش`d��w�dӺ�O�Q7v�X�� Ns$Mj���`�ʍ�P.�$e�*�
�D�ğ��̈Le�IP2��@�뮉��hO��c�Γ!��
ާ^�>���|�2O>��$� z��=�!�1O�����އd��D2`��b��X�f���|J�?LO,U��w�- ��̽:�L�ޞv%�KƎ�"0��ݩ������k�2ݟ02����`i�m�X7�<B���iĆ����Q���q��1D��]i��
p�~�ᇮZ
�>A�`˵&�0���׬Q�~騡��џh���V$M�+E�&Ww��+$��?�A9S�mpI>��O�!�S@�;fn4]�R�O���k�(>m~���Ȏ�Z��N#��D{j0���hO��"2P�[����/˸2qx�{�V�l�ɽ(����q�:9?����7�s����p,�+My���g�0X�0��P�ϛMG��А�?O`���"S��svƄ-Պ r, uΤ	���,g�`M�V��!bGb��2q��p�����d�R`�E�'o�?n��5eˌB7�����	pC"�3�Q���aN���ä��<O
ꡯ�RU�@�m�Q��� �^z�Z���JT��
U���C�9{�����ꈳY�Ь�Q�ig��j����cNf4@�jV�X��D�YPb���v���=�ܐSu�қi�%�թ�O���O8�I��C)pS����'��y��ٍzF� S@&�=�̤h������� 6����?QD.�}e̥j_�M#c�QcG@�!E͆�3�J:�F!�� ��<yc�_��y���3��5��nX"s�jћBa�5��'�(���u�TT%?��XH`�NA�:H]�P�R���Dz"��+�$�y�(\=d�Q*��Z	���!p�:����@.�$�+�!X0+n æ�HNe�OVݤO�U���� ����mA�iU�O?��17,Ҥ'�*6��mh<����0uf�D��LM%���� S4A�$!��Y�Z�%�Ĥ�O0D�O��IB�Y"�����'�d��w��] �-`�@ v��r�AV�=w����C�����t{,�a�'�I��.ծW��AA1�>&���K��Q=~kR�D|�b�h���X��q,3Go�Y dJJ�к �1`0�DZ�VP�!ʱ`�2�>���� ��a���#]�u�Uf]o�'=b!�'�$q���X7!�n�[�'K:T#&�?D|���]�=H	���S"�>���A�e~bS>��$��MoB��EB�?e�&��U�<���5pp4⢋�O�i[���#lL`�In:(d��>��n~bE�8H�P;U��N�|�s0h=�?�����갪���G&ѡdM�l*S�%�	@'>�ˡ$G7x]µ+�è��a pꃞ\�ru�'#f����x�M	]�F���W2@��ñV��yK�玧@x�1�+S t�8iA玗4��y�����ywo
�	��m�p
��r�f�y�A�9C����4��6� �j3�i>�;c��6\�V���O�ӄ�vA����NwB	i�cT�x�8DD��B��ɈPy�P�j�&�����!����u+
�=g��c�P[��aX��x~_?A&��7���w�\^�E8�>q`2�<s�ԋF�r�d���I�4-���'�?�7OY�(� �MҠl���)��3hP��pN�8<v< �	�B��0���#���g��,%��g�;�L�t��Y��B���vF�x��,�p�!�� 4�H kc,��{L�p�	��M�|ڱ�۰"�$�S׈��t�Z5�a$�'"�)FAR5X(H��'i�q���T���b˕�F	
`���^:gj�}BA!��?i������R>Sl���?)É��g2�qYt��Qk���,A<)ǁ��C�0�MP�VӶ��h�M�
8���zQb���uk1e� ]�\� ��?�J�-'E~ٰUj҇j��=a�3O�9+�Ö�>U����Gp$ؒ� �(����E�e�SOƓR?��ҕ�'o��)UlI&xud=+�L��)�*��O�I� �gް �ˏ7[�h	�A�>aEF�?/6h����I�d����;��Y� ��BI�w¥7�@)x�hѫ6C	����u/L:1�
���I�1),�j�B��$���B/�Lc�$���R1oJ���&_ �D��|2��O�<I��胪f�dJ�	)H���'<H�U�B�~� �ފZ�(�a��is�6m�?t�������J��{��?7��b;�T��mSN������P��t����'
q�GWo�pŎ�igL�MA<0�k��vMjAS�|?	�葡[T�iVb>��.�F��R��%��nޡ�9� ٦}����'�"�q�PR��|�Ɇ=e��)qH�����#�T�d��m�o=x	0��O:N��BaA���=�'Y�)��Xp'դ7��h�W��x̓w �i��<␤�V�ܠE�RL��M����D��!�� +2��	<-~C���CD�:��Z�nHK�䕉>��M�dM�O���eN��T�^���#̤
V$�I�fh'?�8���Fw@����[�xaDؕ,�����&V?��x��	g
��t�:���:.� `S�8]n�AS�-N���i vU�`����|F|҈A!hJP棑7���@���~RJ�_4�S�:[�(�� I��s��2�Lßl�p�J:+��P�яP�g�<���ٶOw������ڰ>��N!�x�"[�C�\��z5��O�ĉ4l��<��^U*x�&K\��:���gV�#�\�VF_++K܉��'n�퉐�?|� ��DL������h�j۴#َ�)�ЈB�ҙ��
�����RP�*`'����D��,� �X�B-7 .QSL��4�<��d  Y+2A��Ѕ@�
�P����� ��j�\|�8���I�
�"4	Чhö����'��q� �P |�24��9��d#D~��Ѭ�*e�E�Ӆ/��G�a�HԢB�=�\�na���0������K�^�a ��v<m�ƣݸ8u\� ���][(<cC��/�ڌ�W�%�O�a3����s���`�J�A�a�)�G,��M3$m�P���L�O�x&>��w���^(�Pƌ��,�
f��p?9G��vİPb�DIu�8�0fhR�Sv� �ԭ%6DQE��CƦe:g�x���L�p�0�����"8)�O�3f%�dō,E�`���<aǈ��`�%Wr�(��F[#��4�V�J$ry4�#7�7o|Pxr�>1Cf�//^,�����YJP�@&�F��8�.���	Đ�pcCG%`��ئO��aƇ�* r4�ĵ`0<0�&��[�l� $O3��\
�0eY��2�ժV��@���C�R��	Q�-�1\�h��'�l�إ�H�����v�#��޼=�L�������C��"��֬�̩�>�ݚI��Q	�"��-B��.t�*C�ɦd��c���n�@Ys�Ťu-`z`�B+|��<���A�����	kZ%��(�>sVu",RzC��+��Z)q���&�-O�-���ݕ+%� f�v��	�`C��0n��v��'�A1uJG�?	G�,7| ! 4't�bK�N�'j�m�����vNp��Y&�ȂI����)F2L�Kݔ7�1sЦ�)��� L������U�D��$�ڊr�@�{w/��o*p[��'	�T4��V����Mʜdz��^�s*(c��;O\�� �Xd�'����2�ҭ��Hx��`��T�PQG
O�I��m�_|��:%͚;�ڬ���
Tf�Dx���X?�AqZ�u���[c�5�~b^�KPd8���D�m������а<1�a΋���8).�2uC��.�{C,�Tn����O4�+���wD��C�� �0q�I �l���ı% �W���	&��䓂RGf���ON%7f&��PP#b�bDj�M_	�` u�S-jX��f!V�F]���� 9,��qSq��N�- ��*���,X�I#�)��Q�����V0|���`f�)N.�C�Ɋ9�,��1i_()h�S�*�����=I�O�ر��'o`*V��'>mª�����
�'�tP6M$b��p����l\��6,I'%S�A���=!�@	�͆�;ϖTS��M1���Ė�{O�c��;���o읣�$��%~0h�7D�8س�/d�lQE��:>�6+9D��"r)�ɨvET5�6�F�7D�$a��M�t�(R���8 �,�A(D��Pd�����̲:��aB�8D�(Ю��mG�Hsu(�:�٠�,D�@;�N3��\�'A�!��{� 8D�x�1%Q�&@�4+2Z�+���jm5D�L
փI��(��K̪D���c�3D�|YC̾Kw輹C��R궱�7D�8Ctkz,���
.�@	�� 6D�L#6V�P����2V5*�`�#2D�t���<'�α`""��dm�%qGh0D�� �i(�Ŏ@�r��2����8��"O.���Bĳ]|�pJE�I߶�"O��ge�:}�����4SĜ5�"O�x�Wf�5tx c
��_TNC�"O^�9tLr�I��nɍuk�B"O=z�l� O�@�,Q~���Y�"O��qd#���(M(���$p��uZ�"OB ��
��b�u��	�(���"Ob��^�i��b�ׁ%ʥ��"O�а���ְ���A�a8� �"O��愝&lnxa�́>��� "O��H�(%�q:$�]&9��7"O�Há�^-	��H��ݺc�.��"O~�2�ŚeV�0�� �v�j�"O�˧CW�za�Q� �͒�%D�T��#V���9q!���HF*DH�j(D��c��	�"9��、='p �B�!D�tv���&X���-_���c4D�Ȳ��[o�>��6�D�y���E�1D����"t�壵急VE �w:D�܂KצB� �Ġُh=���c�:D��1@���;��h��X�u^H�둨9D�hSe�N�O �T��DW�*�y���7D���tL�{�:��)��	��"D��	��Nl�����X*�Ua�L#D����)�SH"�b��ޡ�n�q6`!D���C#�U��,
��� d~�� # D���ՠ@+�̹K"��	�P�( �>D�d�W�I�F	`H�A�"<PH$R�f!D�<�AW
FX]��eS�xkx8c�<D��Q��Ţ.	b�����4	߂%�Qe%D�t�fd�[��ɚdȐ>��p�$D�(�D�G�I�>�ɁkN&��U�� $D� XA)�R*$��GA�(+�0�@� D�08Sf��?]v�br��$���!�
#D�4+��_2 
����:y����=D��b�'ډ~N��CVm� v|d���:D�8���0�]J�]�3�c�!���+")�u�Ѭ�Je*АE`:�!��SC����#�Q���z�.P��!�$@�i�5yo�w� �$L_6�!�$N�Z�*@ �� ����$�{�!���l����.V��uhp�>Y�!�d7SԞ@3%S<�d���&
>:"!�M�i�eی?D�%Rˑb�!�Em�e����	*���Ū� !�OQ��׃� �=zI��V!��:,��<0ƪ�-�� ��;ء��@1��#H
5� ��1JL/l(^B�	�JYJ�k�հ"�Ha��K�*B�I'��@ජ�/}VdS�e�n��C�?k��d.�<$&:�CĎ�U��C�IF�����A���)��C�	��Ė�A�FIHE�ϋI�p
�"OI3F�^2G9La�� x�p�e�'�ў"~"�Ӕ�8V�� hY�G ttB�Ia�>�𱄐b��k���-igf��$h�9q���U��`����g�yҌ�8_WB ��C�%w'δY�@��yr��1�aO���TEO��Px��i�$51�P�H<���r�]�a�.���'4"Mba�A�F>�)�*Y�,�:��2�S���J�Fl ��.���,�����)�y���K��cC'EA����"��P���π ���e���i�X8��A�X�$�a�"O��Ʃ_�c� �d�H���ב|R�'��}���ٳp]:���%Z�@,i��'kN�h��ܸv�e�v
ȳI�ڜ'yў"~*pEZ7�F� �dQ.)����N�<�Fԓ)�@:p�Q�Q�%����s�<�AH�0JJ�s�)\�L���R�HF{��i�#Ŋ}��i)H�.I��m�C�$s�F�2��H+�5�7�Ԙ�C�I�)�V�7�ܝR��D��:�8C�	�OZF��ǭ� 7�2p9%�@4xL2C�	�Z�"L��-	�\B
�9�+��I�0��hO�>U�%�"@��0;���d�T$#d�3D�Z�޺4� �͜�Gd<��2o1��6�O�q)��ÍE����� ?~`bh{0"O~勔MM�{: ����ގ,W�q��'E��X怅)@(�/�ًu�L�y�!�dܵg��k�eХ/�����+g!����ykq/D�jsc�;wR�F{ʟ0Y:��ա'�.���៛V��"O$�R/��$k�D-'���8Z�<���'��9i��׼O�dkF냩Vt�����$\�%�h���ű)'~���D�/&!��=v��@��+q
i�$$�8G!�%B,�;�E�8
<�.	��U`�'��|XB���)#E	�E��>Tp�'����#�l� �[�`M����'ȼ�S0��l���1�" �zX�B�'5��tה*%~ŉ�SHX��'�5"bٿ+�+�usTUk�'+$R�B6NNȀ�,�>|l�	�'�J	��V2� ��-�j(B
�'�y�E*ˢPl�!�J<� ��'5r\�@��2Kezy�P$P#����'��	�jM/Q��Q��3�6Ѐ�'{H��Z7�.��S  =(
މ��'vt�`TMNX�t� ئT6�H��'f��1�(�P4���R�U:�������OOe��M�b!R�M%�H��gh�Т�-h��UB6�T-r7�,�ȓuxPb�/��!F��+iݖ`��hC�P+�R"���פb�>F{��'�a�E��v�����R;/���2�'�����*S�#��%YUI�"W�Uq�'(.lkV�T�`��]���!u*�Qx���'J�(#!X�F_Z��c	��*kh�	�'\�q�جE+^iqs���)���')���ƿ{�34bPB�6)C≝F8���a��d�z��j�n٠B�	? �~)XV枎K�N���PS�B�I�C��Bd� T@�FR$V�C�I8tĨd�׋M:]��)ϓ��B䉀/�}�A"��	��*��B�	:fjyHw���/��$�a˚s�P#?�����T���pF��+T≡�2�!���,'[�H��ː�N;�0�p�O 	�!�#(�ؤ�s��'9X:��	0K!�d�O��� ���R�|0:�)�H���[��'`ў �q��/I�$4ʱ.M$za�2&�OP�	�$��cr�I*\���yU�@ bB䉝@�45���*2 �Fcɛxd.B�4C����tg@�o��&��'�C�_@�,�T/�9X���w�NX&�C�?*LD]�Vxx`�K�\��B�)� :h��/� j8&�s��',N&�+E"O e	q@̂Q���	��y9Tq�B"O.�Q�ʝ
M&DNH {e"O�@�Pc	�(�M�'jStE�D"O�d���2w,P(h�ڵ|�:(��"OU���+8��jv�T�u@\� �"O���Ǫ�9bq���2�4 $Z�"O��Ƃ)(�a�B+�� ��rR"OhY1� B6���k��,@��"O��2t[6?T6���U��k�"OP��u�J/Yv��$�Q6�&�8�"O8) 7��*E_�� �q�T��"OXe)Rhޟ>V���L>B�ȼ��"O�[R	���%�Ǝ[Ep�uk�'
2Hɠ�5f�$��3c�)B�8��'�T%��[g���b�ʞ'�d���'uf8�b�V�I2��Z���좍}��)�)<5��m`e�ʹ71��bW#]1�!�$6�\���j\�t��A�Uc���!� �G0"E�rl~�yC��ŝ3�a}��>�Uē�>xF��+��ET�]�Ga	b�<yG�l<\�S)B��H��VJH�<sg^�.����1�ér?P�A��Sk�<!��ʰFXus���+&Y6�AD�R?����S�dR>���됷J/�(a��޶o�fB��+N���srJ5 <��AE^�(B�	�XH<�	���P�(a�ri�iT�C�	, ��4�T
ɾh���"q"��#��C�-�����c��c;�5�C�0K�jB�	�H�ểW&6H�5��DR�.>$C�����+�&�3y�jek �Q.p�B���@a1F%�24c(M�B�O�8!�B�I�<���I &��TՀ����B�I�i�,!�D�i	,U�g*�1{��C�ɿ6�����R�*��#��o�!�Đ����˰nVdӰY��ˋ�����	�T~�u�2+]"92T�&۳z
6B�	�~H�J�	M.x�VP��ډvhC�ɓ"�j�����bxhd��r'�C�I�nI��x2�^�-�L��F#w�C�ɛ���0tkW9���H`����C�8sJP��U@rFv�Aa��!� B�	�j�.�`�Ȧqe��ŝ���C�	����B�� )����[�O[�C�I!,D>tV�E+
�n�����C�I4�2p2%��9 9B�c̽��C�ɶ0�1	�	ȝ=k�HvA�� C��J%�#��7:�A�����i5 C䉪bVNh�#��c��M۰�ߏZ��B�I�&4ѣ���)z�h��S� :�B�	�h^h#R2&q2e� H\p�C�I�lZ@�҆�qD��׫� J��C�	�IYz��-�(�LӅ㗳FX�B�	#�����jJ ll���-��+��B�	%h&��(��̋#��E�c�V3=$2B�	�PҎ��i�fε��ּme&B�	��>���,�P�|}ؕb o"B�I���)c��*�N��b��V;B�ɜi�0�� l�:�`��^VC�q�8H���:hY���,F�B��*uV�1I��.b���+�Ç��C�I�&I*xP�ҏu^찰&f'��C�ɌK �qR��6B�̨�g�^�JψC�	"D:���be�5!��8�C�9M�B�)� JD��O�={&��u��X,*���"O��+��ϣ	m�!a��FrF۔"O�e8Ĉ[4��eJ���*>g���"O��!-C7D@ �+�t0�"O�� B��mQ����
�} ��"O� ��m�TY��2�+�!0\�a5"O�R�mڔ\' ����R���@�"OV�!�~�0܀P!�#�L�ba"Oj5HRh��+�TԐDʋ����S`"O����6%fQ�I�5M}l�"OV�(��j����D�!e˦x�1"OB�㥇����2h�J����"O� !�-�� ,^̀��x!����Nx!򄂾�t1aG�#g��gZ�j!�D=����R�:STy�E	�5h!���N�p!ё��V�F��31Ns!��N���gζD�Z��M�p!�N���i�jMG��l�B�A�}g!�A;PƠd1�O�K��A%	^�UI!�dP�5�\���e�r�ZH�Q#!�QR`y9g刪xp�<�#ǾU!�d�'*Ɏ(��.l�@$r�(5�!�Dء8G$iy�0 ��=�ԋ_9A�!�ُ��LK��!x?
 #�M�z!�d#(_�⢎�9.�ԩ���	%ij!��̣E�rq䕮?���� �@D�!�[�f9�|*�=8OLa�tKZ�"�!�-&���g�#D�a�$kJW!��%}�����X(r�(�ů"�!�d�s{���h����1fȚQ�!�J,�����1&2�����f!�oMl�1A-�1����#A�q=!�> g8P�H
�n˦(�A�^"[!�$֥5����'Hb��(�6A��H!�X{6��a¤߿Lú������!����&�)��0�Z���!R�H�!�$��������c�TiT�IE�!�$�9�l�J'Ø�]�\0�'.�!�$�"4na2�g *`��<�!�D@>>�p3���
�����7�!�D �{3`��	\��E�H��&�!��S�5?�y�@�W�hq�$��w�!�$W�HŞ�"�&	 Q� �@��ƌQ�!�Dϵ��#n}@m��,G� C�ɑcXhl�s��'Ob0*�b�z�B��<Wl�`�����ar0<��	A�w��C�I�w��a'ܗ5BzT��z�C�ɺDP�1i!�7:�X�3hE ]��B�I�6��H#���8�k!��86~~B�ɒI^�c��[6�aa�DIh�C�Ik���ҁ /$��y��G!w�B�ɏ'e��ZSg�g?�q`"�.Q(�B䉑k�R�r��ʕ��E�2)A�ɆB�A
�`��N@�� �o]<�hB�	�<l�x��e��)z�CAV&#�B�I 4�ָ8���j�ڒ���;�B�ɳw��$��/;0!�Q����C�ɥ2`h� �
=*];gH׳4��C�	�T���5�]�<�cB��9/�B�	y�Tl��	�r�q���B�ɼp��2��9��(s�
4h�B䉬1����˅�y�����E�j�B䉗V�4�p�Hm�4�ؓ��'WZ�B�8+��{$���&P�˙�
�B�)� ���$h�p�RQ���a�
)�"O��G�O�
���gՂ�"�	&"O� ҀגO~�T:dG�<-�dQ��"O:y�d���؋r%�r�N�$"O��J�N�?��<��*	�^k�,�r"O�,y��ä�$e
��\�؄��"O^�cb�I�k��q5(K�"��J�"O ,��$ͻ?z����Us��� �"O\Qq!c
d{4X�e�� #BX#�"O�E��iA
w��X/�\y��u�!�D*Z���&ְY<h�	'�Z�!��/#�N�E��+)7|�A��N�kf!���*5�r.�"%V����M'J!��4e�Ш���X�R	p�ڲ�w/!�d�a� �a�)-rX��
�E{!�I1>um �M��A�ZeQ��Q
H]!�DH�6c�J��u�P�ϼJJ!�^<N��IxU�K�P��@�#D?!�$�9Z�\�I�b���L��`�?E!�Dߵ[~@JE�1(8�җ!�$�7\��`(��ϸT������'�!���d|���)�)WJ
�#���!t�!�$�mY�\h��Q�I%đQ'�އ$�!�D�d�z]Ip����Q�8j�!�D�6J�hܲM<*e#Vd�!���$B�����L�bqڌr���!��O�#����dA:Lk@��'W=t�!�d��X�����ā�)S4��6N��!�ě>v��-��Z��Ҵ,3H_!��ӑ���z�$�>Zp�&� $�!�D��w�"II%哷 �����$/�!�dI�Lvԁ# Ȃ�T���#g�@ �!�V9Qn����k�I!�g!�D�	l����Ȅ=Va\[cB�`!�$�7w�~0�P���y#�mX�o�!��[�[�t�˧�H3
����m�Q�!�Dϗ"���q�&ӹ0�PJ�/a~!��ʨw[d��IO�mޔ���
�rj!��|��<��ΏP0�f�G�^/!�D��A��o·-�Xԑ�*̳Gq!�䓣n�L����8o�
9%+=Xo!�M=��e���7QH1�D�ʂ9k!��ԍ-��`sG8'b$ӫ�a!�� a�Z�s��^���ܱVkŰ)�!�̪k��X$�.�� [�*l�!��%;R���F̶1����@j!򄊮@�m���½g�"��t#�jE!�$͕���WM�j�r��٨@!��)K	NEz�E�`:|r0�58!��`46Ļ�c�=dY~,&Ač)!�D7]y҄�0 Qf!�@��!��]�+B8h��#����(��g�!�R�~�=�b W:��i����-H�!���Z�.��3I�4��I�֠�=�!���T�0`)F����xA���v�!�DG�VBֵ97`EA�b�Rf�, !�ٻ[L2�ȉ�b �����ٴ>!�$ �e������92~���A�m�!�D81���/W#FL4r���	P�!�d�5'�J��劰;�����K�7&V!���5�ms��]�C��|����Py��g~��r0��m^d��aϔ��y#ַ	�3�nU)`̦a�񀇣�y"�$CB�EPr���VW��[A��y
� 0�F�G;E�s	ѨT-�y"O���Q̒�1)
=ks"�5����"O�iP�M��F|h`��FL�7�!؂"Op�؆,�d�9�N�aH�}��"O�	9�mK?w��㔃	 aH,��"O��i�Ǒ��-�!\0��t"OF���O=9������R;(���5"O�+T"( �t�	�)��'��Yg"O����̓t4ftx'	��K��T��"OPt[��}`�YrAgN(_��x��"Oty�V��<�����*_�`��"OL�AG
��D���F!�Υ��"O�H�X��ӸhH"���-�!5!���Yx�q c�-&����H���V-�v�p&�A<����M��ybٿPv��H�哹dq�,a���9�y�P�k",�P��/d���&��y�в^�T���$��T?�����#�y�ID?T`~���g� 6k$�17&��y��U"�����5�� �Lޝ�yR�[�24Ș9FI�-�����㎛�y�Q�hl��M�$�0�r�f2�y���*S��k�Q���Ԫ�&۾�y�1��ȩQ��bBl���[�y�MV�k� X���B 6 ��U�W:�yR��{�2p�d��*�ܼ�$!	8�y��\��3%���S��E����+�y�kY4F!�q:MD�Z������6�y�L�%n�zȳ�D*��		�T��y��(Z�^�	�-U%AEz�� �D&�y��IV��$�$˶"��3����y �E��4���� g���
���yb�]�>���2fVl=�́��0�yRB +�x˱�)h��$�C��y��S7{������c�	ek�;�yHUTQ�p�.Z�)��E��y2�[�*�d��W-O}4@qe�y2fJmު���#��5G�bR�M��yb�0J���G�"*m�������y��ݯ(��P1�ߖ%:R 1@;�y���9��š�C��G1���Ѕ��yBfR����k]�*�(|ۧQ��y�o��Hcj�*b��(r���D.�y�����$�"�>I ��8�C�I�f=���'�u���U�JC�I'��!��29���o�x"\B�I���E�^j���H��G���0e>D��g��6&*6�`w�K��x�1�1D��˲ȯ5��]�g��C�� p3a5D�1�C=v��`	����2�D2D��#Ŀo�XQq�/E+0�D"¨1D�hڇ�H?1�����϶[��Q���0D����� S�𝢖 @�=,�:B�I'?�*�RC�$1讕S��ڙ[#�C�ɫS�9Ŏ!Y�PUB��^(#WdC�	>9B�Ӈa�0"��`/T�8C䉗;F�d1"j��.�M�2��2/@C�	.a:8`��ݘJ��P�0 �D�x��0?FH�K����  ���ū��]m�<�wfF|���� !�U�qg��j�<q�C!�-�re�}h��WL�<Y'�U$2I�(�V��GJTE�<�t�ƯC�n�5��P3vy���C�<م"�y�B��#G�j��y��Z}�<� ��5d�r�x0
�*i�L�@"ONmx3J_�mN�)���/����"O��"�n��E8xd{�0-��U#D"O�dN�D5�X�v�F�Ov����"OP�H�;c0݁�-�*a�O<�y���fy�̸%�C�YX���Z"�y�EƬw�����m,��Y oQ,�yB��
XY��6@����c=�yB�U�T"8�����< "�@�!�yOՋ���!!�A<���a��S��y�bH�;
���$7G�m��yR�WuD�	Üw>�i���y2�K�g�1`5�9XcX���ޫ�yrg�!	ۼT�2��IjF�I�C��y��@��$ZRh�42A���/=�y��[#�i�s/D%+ ���%L�y�o�))��|:7$@3&j�T�ŀ���y"�RJ�T�S��$�ZM���"�y2�C?R��i�ꏣ劑x���y'̉#����D*A�~;^=K��Z=�yBA 
ryα�fU�o�9������y���?VMc��
k����"ض�yb��T�����O,X-����$��Py�Dݤn|��pD X�+y���RU�<	���:��d�'�,Hc�e\�<��I�<E`���")�95�B�NS�<i�����
C٣���ц�W�<9�K���L��u'^%KJHr2K�T�<Y��X�Qyg�ܞ�L�	�Ex�<@�P�)���P)�<�y�&��<�%�
�9j� �"VL��Nq�<�a"Jj4��cI	�-�s��e�<afa�	7��y:eeI8~�s�dx�<���˖*�jt����OE�0�b^_�<��/�,Z"��S��{��P�g�Z�<@^�j�Hp �B�$t��N�K�<��eə-�BpJ4�&dfzЛ�"K�<I2U�v:�1���N��@�H�<���ֈc� �ae��7��P��k�<�d�E �0�;�4j��<!���c�<Y�^���54g(��c�<��fA��0���H�c(�:R��t�<��A^�x�
�{#)�
*I�]RC.�l�<�����!k���"CI�$��q�<��j��U����T�� LZ�X���l�<A����yl�Qs#�<A$UX���i�<��i�K�D]ȳ���=[�ݫ`�i�<Yg��;/���(P�
?M���3�(}�<�6o��R��#T�����C��]�<Q4k$^�ᓁ��F��؀INA�<a�Jعp&(q��^1v�N�`amd�<�5��)jߦ�0D���'�`� ��YZ�<�������,��ǔզ-��a�<�`���ɫgE̚QH }���^�<��%��=�SFeΏAB.�G�R�<am�>Rb��������i�n�D�<��^�>����v.TA�HA�<�$AZ�9�<��= _�yAF�}�<1u���:`�+�� ��1�S��z�<I����\��CK�P��,����x�<�ޔWRm����s6ڭI��?�y�B��B�f�A3n�	hۦ9��-�yT�S�~�b��bcb��1���y��l�\ rf�O�S��Hb��?�y
� ���$U�
%.���ڍ[.�Q�T"O�h���]!%t���	ҹ?8>�i�"OČ��0�EI0�Ч"O�`���CL���nV>0��p"O�@��˳&L�$[�Ku�P���"O�[��>5.J�"�H�O`¤/!�d�k`Rђ�!��͹�eQw!��ViV␒TI �|��Sc�X�!��G�@��KG.+2���� �!�䂅M��h�׌�6b>j�h�M=7�!�dG�)��yʥ��~�X���J�!�^�o/�ٳC"ֶ%�M�0���!��߷3�)��G�5"����i3(�!��7T��y6K�6�FpGf^�xn!�¿-޴����)�`<3�g�J�!�� 9lvD���lۼ�zЀ�0"�!��J6AJ&���
����E�#�!�ܓ���㍲;<+)�Ꝇ�Y���y���7S��E��t_^�ȓy�|�E��>]5ި) $T�V�ȓNFPAFO:a�Lɷd�fI6u��4��l�5	ʖ!��� ր%�ȓo1L8҆�,Go�7����y�
�'����P( �������.�(���'Pa9���o�~TI�$�3-R�h�' 5r�+��}���(��	�'�d���넥P��P/��ٔ���'# �J�[���+A�d<K�'%V�3�-F7}��-�&W�Q2q��'x4y�	�=��K���W/4�'y�,Z&Y�z���c[�WCJe	�'����v��Ÿ4�җM�U��"O~=҂�ݳG'R�A�&�&P7���r"O��)g�ۥg�	�V旺3)�a[�"O�A
q���9~PႆC��#7"Oty�d�Hg�M	q���Y)�"Ov�
gϓs@�3�5;(�a"O9��B]�� #5i\	�:�a�"O  �ˍb����ITX�"0�!"O`Iˁ"5-��]X]���@I�l�<�0 S�1u�|�7�чG��R�H a�<)G���߆�����-�P̲7hD�<�#I�x��s�"�[���j�A�<#g�d�D�R ���[��@��jD�<��a�0%O@M Q""|9bvnB�<A����{O��jƚ5��ip��S�<��2m�"�Q�X�|ji�2��M�<ǋ�m.�4�#O��E�%p�G�<�CXw&��#2/ˡ:���D�@�<�\伤# ���l�s"�z�<� �T�<��1d��|�Pc��s�<A4�7�A��B�*������f�<�DI�1^\��O)	��E2�Db�<)RK��6�Xi��Թ;ʄ��׋�S�<!�'ݺo�.��G���p3�pId�S�<!�$ߗ.�d����0g|]��`�M�<��"՝	���Jâ-�.y룏�R�<yPⅆ"mdL�!�ȧC���X���Z�<a�N�T��E#Sˋ&!�|�w�X�<Qw�ʇ���h��=b��
0b�[�<i?��]�gjҩM���	 �X�<���"jNqS`���<q1��{�<�ѡwS�P��sajTQv�x�<i%�=��I���.)XH�&�D~�<� ���ff~�TE�d��=�� J�"O�dZ��א9�} ���M{Rț@"ORT(��OR4dX��lΗ`o4���"O��q#o�9V�e���/$i�@+"O����gV����2�ͣ+7t��G"O���ݶU�l`G�:H��Kt"OV�bF�S�Rhb�����jd쫢"O�P��$��L� U���"O��YBԼv�f�6�0d!rT�A"O��H�/וe̌ B��&{JY��"O� ��ޮF������I1}�,��"O��+�f��`�HX�޶Z˾��"OȊS�3N$8�㬘:q�P|�"O��kEF�2ּ<�k�=���T"O1�c��J�d�u+EiqLdv"Olp�J����x��,[_x�
""O8O]%7GFd!6��! �,��"O���"��
G��F�h� �"OJ%�D(��f�&�H  P��"O�[�4	�D�X��IZ��}[�"Ov�Dɇe�����R�?� �[G"O�=�Q	$l�f�bF2����@"Op���C_�ՎL�e��}��H "Od��4��� �c�,�}b"Od�x�"׾�ֈ#
x���CB"OX̹d�!4e��H�#2I�6Q:!"O��[�]�X[��hF�ҪP����""O�+��)nV�c��2n
P���"O*e��f*N"���#��-��z�"O`MqF_�X����J�8њ,�A"O��T�J�P��:%J�-(�L�ҥ"O $��F�=w��I�FÒ�f�ZŃB"O~�`q��
��� �3gR0 &"Ol
�l�z�p��M�X#�*�*O�H �Ni�PR�
��qh	�'#��sg�3�2��pG[�<e2��'i�����ɲiL��
�NС6JF�3�'l����*�X���*���p
�'�v� Sb	4N4(�x�A1%%��'\�Dɰb�)�nu�YØ�	�'Ć[����,��*_1���{�'͸5��y��ժDf<
��
�'<�g�/�K�8z!@�a�f�<��C�H�9fCO2Q,.�3vDn�<�C�Q�t�B(X1=���9C�
l�<I�ҺH�s��V/N��I����R�<�Q��D���,nqw��I�<�I��W�:���)�~t��8抐l�<�2 O���!���H|�hM�$�_O�<���!n��-��ʀFj=H�IO�<A4j�6L+��
:t�8�e�J�<�gN߅I ��*�X q�`p '��L�<�!�Z`��A�Q"�|5`��F�<��)1+�T���3.V4\Xs*�~�<�	S;[�3o��\���x�<q��3��	��++0^�2-y�<y@F�;$ʤk�� ��X!T�Gw�<q��-S�
M!,���(��
h�<y��$H�	����jL�� 'e�<�ȏ6-�̠�f�Ҫp_8���`�<Q�*nb�q
��% #�t ���Q�<y2@ϙҼ�J�(;͠�6�_J�<A���>D��-�9_��b�}�<���*�8���c-8j�U��D�<� �9�J��(�K�h�J��q�"O��i�O�n�����Q	��q"O�=���.���EU����`"O<���n9�&)�*��U���+e"O�D)# �0+7BL3t'Ɯ`3�!a�"On����W�$�4�T��z�5�!"O�i�`%�aN����'���a"OJ�A�6]���3dĹ5�BA�"O��󈚡���q%��R��h�"O$E"�g�4�D�Dg�
IUnY!��'������G�w�.��3ϊv�(�B!8D���$�ݳ7"��`:qz|�ʔ,7D����OnYk��8�T���8D��(�(�w\�x곁��)���-2D�8���!BY�e��D��=I�1D�X҃��)`�$A�$�‵0��9D�ܹ�*Y�
�I�I ��n%�p�"D�,IW�� J�L��g�@�p�+D���bMeբb�$ɟ&��6h-D����e��D���m�.���j��-D���c �I�~L���Ůhf̐2�.D��*�O�?\��  6h����0D�)�B��gb6����ϕ���"k*D���I�3Z�0�c�F�?Kbz��j'D����ϙ0�L�	W�ȱ~ �=���#D�$C6mȍZ�8�ZT4|��?D�d������[�J)o��BE<D�d��M�S��0��A�6�Bp,9D���!�\%:vY+��s!�ݹ~�xC�%#�Z�q��	:����<=:C�ɢR���g+E�8 @�8e��f��B�1x�$a.IB89�b�xٞB�	]H���O�o�` �*N�5B6B��6���2ec��l�PD��ڱx��B��I,Lu��F;?8*�p�%�?�B��k�N��$g�=oiD6fѮ4VB�	��q�w�>'m��C!~�XB�	�:pT����F
Df��R��$RLB�I�&�|���R�|��W��&{�B䉛 3�x���_�M�T�a�	�\��B�ɥBT����52�8(�DS�|��B䉘VpP\�ӒAГ�U	"4�B��=Y�t�"�N-s��i���T�D�B��+:�<���A�&�^���-ѡ�d�9WQl@���$,&d�2&;M5�y�
-�lqK���'0�����Ԛ
�B䉽"�)�*f%H��g��X�nB�ɒ<�T4o�&C����g'04B��>\���A��:
 , B�0L�^C�Y98��Dm�@ۡ Ѯ&�C�ɪ2ҠܘU��9`�έb�̋^vC�	�TӚY)@�Kf{���w�L(@*B�I�N��̫t����!�4ΈD��D�O J#�6���p�d;L ,�Q�4D�|av(��`.Hxp�Ćq�4Ġ��?D�t�1/1r�(�I��ǺgCZ���>D�,Kt!BJX��*@B�e!�Y�c�<D�p�ři�`��� ����CS/;D���"R4CF ��w(Y�_�>��eH:D�|Ys�>B�`�"A�Y ���$4�(zA�{�EI�E_S��H�ek�B�<� �DN��n��J���3j�W�<���1k��1#��p�"H���J�<���V؀�(���s�`\�DSD�<� �A�C�܁R�41��&F�`��"Ov���b�-|�n�QRF�MV���"O|�)�h�	9W����O�N� �(�"O `HU�W�̢�0�DK�M��� �"O�1z�j�#w'�-�$iW�5�e"O②�������Ǥ@�xځ"O�AHtN\AlP�x��n�,�r"Oz1��cj%��R�l�Z�"O��"BeLw�����\	[ɘ�q�"O:1Ǯ@�>���A�D��θ "O�4�E�A�1��C�f�hHk4"Oȓ�ǒ�R�>�`"�70�J\��"O�Aqd@%n>��"A�J��ju"O�L�R��"<�v)!gO�j>`6"O�Ń��=5�p��@��4o\2d��"O81`DE��""l:UkESx�&"OHIR��6o�Ȇ������`"O0�ᣌ�d��5��X�����"Oޥ�6�^�Q0"��j��~�°"O�p ��X�W�L����|�`�k�"O`19�c��4
 ����7!��C�"O`���D�=Q�d�L�����"OAR3�K�j\��`C #\�yBa%W��h0��Ww�p�*�kD��y"�Őo;��i�.�5$hR	[�Џ�y��H�Nl�!
�+9�� K��y���4C'~���,	��z��[��yR�p�r�C)�du��ER>}I>�*	�'v|Aҷ%G:��'�G6bxH�1�'��m�b�J5Q"��g�F�`f�Lj�'�R@g�p �����ф)d��k
�'A^t�!����b���ux�Ű	�'[5@��
�]%Z��Q扲>�l���'>�t@��ݿX9ЄK!�66*�	�'��@�B���4`!B��T$-��t	�'� �10�T��#rl�(.�my�'�|u���)�>!���+�!�
�'�] F �,w��D��+��G�B��'��`�!�8��⇄�5P(���'�H�����?Q�0��i�>�p��'��ۆ�H�A��2lڞ݄���'kf���>]{�����B�~�zq`	�'�T����gKެ��T�r�t��'` qir�:-���d�q څY�';���1KƞlV�����1q��	�'����b�c��8��K<���'/T�2S����9@��۝.�� ��'�����[����3�\:"�>��'�p�p§�EMfpÍ���՚�'N�5j$N��صs-G��^���'���F�F9'�fȈdmƖN�Ij�'�T�P&�U�,�ZʓH��8�
�'#�E��d�N�s��D�R��
�'
��持G�(��FjH���̰
�'��HO[�|+��ƂD(P����	�'=<LhVb���@�Y��ֵ^�L�	�'� �īX8fr�*&d��[y�8�	�'�&�b$J#V�Q(�'Q�ZJh;�'�
����H�J��%JI�W9`h�
�'�P��f��g=�����C�=n�qc�'��X�S�ۧF# !%��5&��	�'~�\���*<s�9�T&�ZT4��']�0���?`�M���	(Ω	�'T��p
L.e8�x1a�P(|���� \��$�=pvH����$!����v"O.�+�$D�F��*�2,.5�q"O��80,�:��� H?<d�RE"O�!qL��uU���q�֜L�����"O��A�C�=��XQ^d���c�"O�݈���E�h��Y5z�ు"O<� EE�]���R�I)m�+�"O$��P
͑e�A��P�C�a��"O�PapĒ1.��;P� `U�,�"O$RTE�>�<�a�L�GC�\K�"O&����ar�D����	&(��(�"O���F@+2V�{l�v��C"O��!�I����D�K�C�ur%"O<	���$)q��R��V�|:f"OD0x7f��lx��DFЮl��ȹ"O�aYƢ�"?��,y�ߛ��p�v"Ob� ���3��Ya�CX��6$��"O��S��JhEء�Q�er�"O�l�3��S���Q ���Km��3""O
<2�"ʏV�`]����^-��"O�}�6M��$��D���nY�Q��"O�ݘ���S��9�5�YQdxѤ"O%0�i�c>d��
�
pc��pQ"O����I�,�|�U��U����"OLPR&�7�����" �%Z�"O��3-B&&������*-)"O�"�^@b�����*#�Ƞ�d"O��Sף�*�����/�2QZ6"O�0&�B���,	�DE.��`��"O�4B�J�8	/b�;�$KEņ$�"Or�'��%��<�DM�N��Q"O��(�Ň�f傦�L3W����"O�=p ��\6T�ô�?�Ԙ	�"O����$G n��C�A�+8����"O~��EG�"$Ȱ�K5c�ޘ��"O�,Cpa��o�:țV��nD��"O��S̉5r�T��Ƌ-}�;R"ORu�v�J�d���Fd�.}�1�"O��1ר�?K}X5;�$�>'`��"O��@ԈA-$NLI��I�ް�3"O)��Sd5$ ��E����i�D"O��:�V�7C0�)!�J�p]Â"O�*���E=0�xP��3� �y�"O��k�ǎM��DoV�R���h�"Oj�����b� �����ɠ"Ohݫ�j�-�� �.J�ge 4h�"O��8�*�(���:��8To��2"O����)^�
RF�ƍ*���"O�a��`�'J"|�K�a�T��@��"OzL#�eO�IE�t�� ��h5R0"Ozty�řEt$t �����a"O�}� Δ��B���.ب�����"O^h����JG�1���;�N��3"Or@
�O�<p�޵%˂A���P�"O�s�JR�U+�����i���"b"O^�����'\����J��@�"OB\�%�;��l�DU+��=H0"Oڵ�5��h��qd��{���E"O��i��&+�2��ƀ�"e�A	#"OP�K�aQ� }��@O_ 8�"O�쒁)��Ws��2f�Ur��`s"O:���H�	�dтn�2}�<H@"O�
���kp���B^�e�D��A"O�CᏛ'N��SF �da��"O� L IA�g�(�(!FZ������"O�L�!�>3(����eK�1�Ԁ�"O�Q�1�ʏE�ll�'ע7u昁�"O�R%�K�"������,a�Z "O�1#���
�
��QFߙRI���"O4�����-��@Hp��;�&�"OΤ aѢ:͊什�A� ��QX�"O搉��¡6��<s�,�p}*Ux�"O�U��L	�?j ���ڹ�`�6"O�� S�k��HKf�(a�肣"O�\���
T��(!�
T��� �b"O�I�wFJ�u%�@bA�(
��;�"O�m��h�7Ah���"��%G�
��q"O�]���Vo����FV f�2�Ѵ"O��Z��?u��x�bO�c��	��"O�M�fB��������&E���'��'��)�3}��O�jz�hE㏸�Փdf��y�y���*HV�lsS� �F���Q�'i�I���3(BY*c�E�U���`�'IR���G"o�Ʊ��-@ L����
�'=�|�ҍ�1Ch�YJ�Du�
�'X�`�r�(+�x��f!�5{|\��'�l�����-<#��ic��w#(d)-O�˓�0=!��DuC�ѫ����:�� Pe�]�<��	-Hy��� �R����P�<q� c�F�0��	:�ZP	�F�<)ѩW�ys�e�GME�7�� d�A�<���(��C�@��e��C���<�` �xR���[�i�X��d�V�<�e��>?�X��.I���E���V��p=y�'��H�F��w$��Ժ�a�4D�l�!�v�PQ��)�kf��6�1D�����Cl�Z�I�:Oj4ղ1;D��p )�("�t���W v�\"U�9D���S�H����	r����Om�<)P�E:vD��$��nj��υ]�<y`%ӲBhX�i��_S®6�N��?qJ>	/O1��R4j��F�4�B�k&LݛI~9�ȓPj4q� �χ> xA �Ř'�.ńȓ�F�j��ں3{�К�ƁP~ ؇�nU�t���Oޮ̢s��1ymF@�ȓBr��9VfΜ*��yé�~? $�ȓIN5"!��.��01�R�<$��ȓ�VLK���j݆��芏8��e�?�ӓ:��}1$*&ހ��GA.�$U��abL����7"�Q���^ԁ��Co�Dc�ùz��9��͇6X�D���8;�]X�K�8R�H.C0K���ȓi�A��G8��4j�H�5b���ȓL��8�@�mֈ�p�(M}�܇�*A^m�U"Y��t��1h��?��Q%���'�ax��q����'"�"~\8Y4O���y"�K�4�����A=,��]hԦ��y���Y�ɰw�N�����E�y�P.(�=#a�K::4�Ҕ�H��y�J.ZAn̈P��n�x�P�	��y��8$��y�e�U76���2�y��7z��S6�߱z%�xҗ���y��^H��Ew�*����/�yr�
,"4����EN6�b�d�3�y���'ZRyB�ǆ+�.U�&폏�yr��3�D�੍�#kƄ�"��3�yR���c�����)��S��y����E�,�Z���'��Ųa,O��y
� ls'��Eh6ؐ�Aԫ	����3"Od�9��E"`�0�Ѣ��D��"O�陖/�"LY����ϛ�V��ѵ"O4�ҧ�Bx�p�A��25w>��"O4�A�� Hn�P���d����*O�|�vυ(X3��S�n51�T��	�'� 9w�L6A��d�6N�(����'��qf�*B��L"6��$_���'�J�1ש��'���#���b`���'t�{�  `�r4�gʍ�n��x�'�Ĺ�
ٵoB����̂���'���2��Ҁ,6��#r E3�`��	�'U�P($c@�AJ�Ժ��U�{���'���JV�Ѝe#쬒 )YkpE
�'�6yy�D�N��+`�E�}q��
�'��}	Ө@�?*�"�` �� �
�'$@%z��V��X�s�'��iA
�'f�)�_���$��e�<&���	�'�0�F�[�%b�X�͎6�Bej�'�*M��L�^A��9��R $0,Б�'�qf�G���WC�.���'�(H�CŰ
6*��6OȆ}M�M�'��XBp�Z�&`j��2�&v�����'�$�q/�f!�¤A:_�,qk�'���#�[- -�6e �S TX��'d�i���ʔ;��s�DAԠ��',e�k� �S�l�j�:���'5���`D�/j�$Lː�Q�d���b�'��Q�M�6t��A{%��0^^��p�'.ZL���>"�N���~9�
�'��e�e�\U%X�:���8���'���S�W7 ,�ȲEV/34ݓ�'"t]j1V/8	���D)ո��1�'~z}0K&_� ���&���p�'�*���e��L�^�����k#��
�'�Fa1�KGz\t�Q�E�\�,UH
�'`` �*�\Z𪗒y����'���"*|��PbeP���y�C�'M��tatjةx�(q"@[;�y���O7B���!�&d�K���&�y�-��md��+��u���X �G��yB�<H)��'mh3ز��A��y���0�(x��/(=�h�t�T�y��D� Ȝ���ǁ�Cp�뀆H��y@$T�J=�q��/?��hC�̨�y�#� ��`q� '8�T�rW�U��y��_�� yEA��(��yxV��y�F:N��xs��/<���Fm��y�)�-~Ȯ\�Ba� "9�)�e_�y��O�(�`��+1�5Qi��y2ɘ��j9���
�8��QG��y�?�B9��̓.a\��P���y�;.ܱ���D
{ڤ1�I �yR�H/} ��B�ˋs�����,"�y��-����g�f} 'f��yb��h81`�ő��T�!��y�l�d�X�惇�X�j�x�@�yR
݅Ki6�s��
�I�^�Sь�y`�<4u����j!v1	$gT6�y�n[��&D��/.l��tT �*�yF�Q%@��qkbT�*�J�y�iA
j�(PYD�/H��s�S��y2Â�Q؞��h�}z��ڰ�y"�ۊ:N��� �f�6L
��y
� J�땪/v��t�Փ1=�6"OPx*�#�0OR��v�0V�0 "O�!%�	��N����� $�l:"O��Ҧ�w�~���g�/7���F"O�7L�$R�C�B|��""O�MW��.4ʕ�f�öGf�͉R"O�-`D�G:�����lZ�cT�"OFr�aȞqK��Ic��2Q"��2"Ofm���U�Wbf(�ǯ_-Q�a("O�m����mբUB�.ՙ0� pc"O>��ue˔u�½kw#,_�t"O��vO�dz�S��H� D�d"O]�ݥv2�%b� �6Ry�V"Ot١� 0��1�!k��X@�"OB�( ���(�0�D�(oۘ��W"OX�C��#��y�'��/gR��"O��Pq���%(�Pe���Z�U94"O,�B��)-^x0��ЖSl�]��"O�9�.����2�FO4w")��"O��ǔ,d1����� w6�%"O(x���1KHݐ�N��A|@�[�"O4�+��-:��g�V�7[:���"O��Ѓ��*��h`W������"O���3���
�h��,��w��-�a"OP�:BW�C���(BFǆ "te��"OĨa�eғ5|�����T�D��I"ON��'�E>Q}|��A�	j^�!�"Op,�QǛ4|�-
��݊Dn�T{�"O�A��9~&<̘�.=[�j13&"O�=	����Z�"1�V�N1ȶ"O�0sm��f��Y��߲x~V\"O��`�IG,&\ �Y$lJ�vtTHe"O���+�%\ a�L�:+Z��c"O�Tz����yX"�R�A�%�U(�"O4���Ƴ}�8єJ\>d��=2�"O|��E*E�	���bp�^���"Ol1���(8�Af�� �|��"O���F&v�Q�� >�\}85"ONE��Z)E���Į��t���"OjS�A_u�)��cU�`
ԣR"O��Ys�żN�"A[8HM�p�"O��cuh+Jb`)B�P�<�$��"O����`D�+����nϺls��*�"O�mbs��Y4�x��Y�'[�ۑ"Ox��#IΪb�2�c�!J���P"O�ث�/4$ӄc���#�JA3"O���&�?"\��7��v�t=�'"OV�`F�h����!�ء�.�D"OV\0p��	~e���� ��$3v"O>0�0�гV˺�#�"���D5��"O ����"%������b�Mb�"O���$�ɒLd����:<�5 �"O��33��2�qb�ʕ�E�<�Q�"OJ��$��qpx�RDQ�Z�9"$"O����DX�"@��It"O0�Cq�Q�$H�!T֒�d��y"cN*`�8�� >�4ȖL��yB�C�{3P�e���2������^��yڌm���@G%�"^ RC˘�!�_=o��iƪ��^� �RHZ�U�!����b�:���y>@Y�΅�!�DQ�����*uZ�]"�����!�d��fn�+�l��uK�	ZE��2!򤝘G�\4rC��RB�u/�zN!�� ���֗_Ʀ���D�e�RTx�"O�]�h�(l2�D��+ɸА�"OJ�%C�7����s�D,���"O]�%�%-ߘ*@�F��f %D�hӤ#�!z���k�oۄ%;+��!D����c�6I��NZ3d�x-[VB?D��dA�>i��#��+5���>D��$�
Rdj�ɣO�*�Q:Ï>D� �&nA)-�.X�F�J����Ջ D�P�Dӡj.�����Sﺠ*� D�q NW1%���CN�i3�X��B>D�(��)����Pr� �#Rr"�җ*>D���	�I΂#��F�,�ˢ�=D� @�h�԰a� ��*�$�qe<D�$BU�θn�le6*�;-�gJ7D��Ue�r�-��n�c5a��f)D�1K���4�ŠW+�ʕq��9D�4�w��J U�1U��M�j9D�(���� j��@N�b/l���A7D�P���
�`�!�"m�!�*7D���E-��Ś}��뢼���5D���ӰxPb��CVc�Ջ�*Ot���A_S��m�,Ԫ���"O��v
9@��`YsM�\�����"O��� ׄ�
�B&�/��љ�"O4j�o�(�hͫ"_3k�)��"O�a"����h��\7\0 )�"OX�;���	�$Äቸ	r@Z3"O�Z@T�l6��[�����&�ybӝ(�������q��Xw����yrf� R�M���	�b�ALB��y"��&���٤��_�:U饍�(�yR&���]Q�^G�ׯ�y�J�n���C�W(Q�+ˈ|&C�	�O��ѱ�_�PD��ǅ'[��B�I�8�*������9�<=z�"��F��B�I�m�r��"gY%$`Łň�B��B�ɰ_��Q�E�
 �zBI�%'�C�*f\��c�đZ��hj�DTm�B�	�a��eQ䓔r�мR�h�<E��C�	&C%���䂈2���T�
,��B�	^�ەȇ�`�,��
0j�B�I�nF���	;A��b'�7��B�I�BT�@Pjش�� G�ˡ�DŦ3e������-�Rص,�{H!�$ ��p���� ��Ȓ�6T7!�D

�`hV��8���j��I�!�d��L��u9U.O3G�*�oMj!�D,Ow�sU��:m�ݳ��Ãt,!��ݽh��dz"M�E���P�Z�!���2wf�<S�:Y2<U3bbڇ%!�d�"��QAգ� &>�����mH!��L��p�`3~9��	V�[0!�\;f�\�
���(ΐ�ըO�y�!�d�<j�xsHS(!��S�Z:I�!�d��m��yw=�脠b��!�̷xθi���ҎY��HA�H#!��Z�p5$�� �I�A�V�{#S4p)!�d	[*
�ǼFo��5n]J�!�d7�"-�7���3Qe;n�Z!��Z.���h�GџMY(	�#� -!�d�4Ť��3��Jt%1�j�!�Ĝ8mv�S��'@&�:� U�A!���5[��<;���'%d|2�TD�!�� r)S���?)IR��n�=ܰ���"O��G�L��t{��.4�P���"O���b�B7�DK�`��j����"O�IT�R�H��a�ک�F"OJU������ԉ����
Z&8Tڧ"Od��#�<_N��@ĈQ�&�!�	[�O�fc����#x���DE�'��8��'�\��g�8(�]��X�2��'�~8��ė=�3��S"G�������*�' ��Q�.	kv����H
I#xX�ȓ:��Y� �Qd�r�b
P�)���ढEE�Th��Ĉ>Ivt�ȓG��4
5� �la�8�8"#��=�
����ĀU9v��Ǯ۲%��p��M� 'W�V$zt�[�Z���BFq�<Q���$t�I���w�|�4�Pp�<YT��`�5���J�w�@��d��w�<AV�$kW�	�K�������Xw�<�0mF �*��S#ցITBG�Rv�<	4h�-SP*8ؔF�N�y�c�p���<R�[8����G
?�aI)�b�<QSH�=F];u��&y$
T��U���O�4y��:>^���\���.�y��ǔA��,R�`�2�R`ŗ,��d-�O��f�U>��l	S%J7|�i��'��	l����t��>�F��k_�"�lC�ɲ[�,,�h��t�p�ȃ�,b�<����:����2q4-��$'HJRh'��*�`B�I�v04-�P+��E�n��C�=,)Bb�$��p<Y��4aζ��֪��W�l\�'��x�'>�?QQ�b�4���P���|-�� �l>D�H+G��1��ʴ��e�$���E=LO���&�D�����S�z�� �釀~��^��H���K2䛂�Ez�$b�����	a�Oㄕ�Lk�>�!ꇳ>$Z��H<1
ߓs@$0*#���,�H�+J�\r�Yưi(�𤖝3�F�Cc�.��D+��K�Q���(�|�S宔�:�N!r���"`������2\O4@��+X�G{Eʑd��6��<�C�i�Fy���i��,"��D�p�\)��&[zJ�4P$�)��<�  W�un�rEŖ:.6,iS��b�<����%c�� �+_�{զ�<�	�]����%��f�����ǟ�n�����hO?��r&Z�T��dr*J�e���+D�p�bd�I|Yd�T�wv�H�K>?����=�7��&�8�h!��((�P�+w"^w�<��\	�Z����S�3㨸��v~��'���� c��QҲh�O*�	�'�X`⍄=딁��K@�|����'<"L�cLL2�P,����
L�Z	�'ݞ�K�!?���c��3:�5B�'O�H["��6:~!*�ć�,>q�ߴ�hO?7�W:+�D�3HA�~��ӬNW!��#:H����L8�b����]7\!�D�]�^M��oW
@���؇+B�%&� D�H#97�pS.�/v,��`O��yrF��t��x��+K��c"��y
�?�$ s���Q3����,��y�K_)Q���	�E%���˴J#�䓾0>a�#F.S��:�+��z������`�<ɓfːG޸�c�ؿk�ұ���Be�<��h�t�"� 7n~e6��"�F��E{"NT��M�iA�D�ivL�V/!���Ms�|8Ci�.L̹ ̛�,���hO>� ^����TSpR �q��;l���c�"O���s'ź^���� �O<\�Y�"O$-�u@F�y6���$�+�lHC0"On)�� �,[��RB"��c$�m�"O�9p#%Smfm�� ܱK!�=��O�=E�D��.6�vM�K��	9�MkP% ��y*�}��<�d,�/| �S�Æ�y��iό��=�����'��X��I�d
�"E5^�nT��"O`�a'��5�Z<�#��:.Q�e\��D{��I�;#�8E�5ĚO�Tju����!��
n|q�b�C�����FLÞk��'���$͘
vt�1��:d<�+��?��h��(�@����A�l)�ˠ&�jhKt"O�t�RD���h鐨�P���������E��ȁ��
�G1;@�q�"^�y2��(��S�"Ҕg�b��s�"��OT#J�Ȇ5�F�dK p�,�`�Br�<р͟K-4\��L��,�'"AC�<�!HT58��$��3Q>�Bl�{�'4ў�p����A���͠ ��6�E��H��Y��
ޒKCĭȰ�@�K����S����,h ң��k^��	���-Ğ���j3D�p+�KԹ�p)���j��� �;D�,��lX����Ȕ3f4(pZ`�7D���u`���P5������B#D�B���?y��K%�J�M2���'D�t��h�1A)�=���bPHS��$D�L
��<�t�6o�!f��=� #D�<�֫����s3��9{�Y���<D� �X��}h%"�*��GE�<0�O �=%>�yS
L���!�NO�,( f�9D� ����Q��#��ҊFe`H+��#D����ƫe���z�$��d���3*#D���B	�_�0��e*ɤd��P+�!D���'�K�)�����	�#^��3� D�8���8`2�D
=PZ�Y��&=D���` ֙oɜ��R�
1^�y�n:D�� %,�;T?Ν ͽY,y�V�5D�������,���A2Y41�w�1D�d��.�%��GA?�8��*D� 2�_�E\�3��^17=��:gh*D�i��Ĥ)�He�[/�|�-#D�л��W��B��!W�%��AR��,D�`ae�Z�->J ��aڇ�r���
*D�4����8��q&*�
�\E�7E)D�H0"��r?�� D�+Ft�t�3D�<AwjIr�+��@ʤ�$���hO��hm���]T|q*��D�kZq��"O�a(�� n�-鳡�E0��c�IG�'
�I�4h�+�G׀w\�1@c#��C�ɡ\��Ђ��K/�E�7M3��N<�/O��=ͧC�Y��bH�����j�t� 4�ȓVe�lt(
,44�sF������ȓ�����"\^�h����J�����I e���$KZ���'��U�(�6)��k�NB�ɰ4�$�4��%����?+�#=��|<��݆.�vj�O�X+R�ee�JN!�$�d}��Q ��F��g��r��O�=�� q��!TM
��DD6]�`#�"O||"��� fѰ�n��*t���+�S��y����V^�	�g i8�J��yO�@�xlj��*����iF�yr�͐
(�k4u�x�(�+�yRow<:Q�*_g�LDkB�@&�y
� ��)E�3|bL��C��++�\�Q"O̱�h��W|쵭/
�A@��y�<	�D* �Ta�P呠2  u�w}¬7�O2]krŜ�n;L�2gɣA�`1�U"OPq0҈��fh�3���"O&0ȕ!ܔ �A�)$g�,����4�S�S�����LI1tx�f��Q�,C�d;�0`��K���I�4��2M�=Q�V����O1)�ส�!ڂ3�h�ȓY�X�WD.V������rĥ�'�&�c%_!��C~�ԡ	�'�(I�2,L�@��1���
ļ�	�'u�s�O�%����W={͸a��'�x�!����(�H-"+7�t��'�t�Dkʨb�u�u�����
�'>�P��3g�<�����9^rpR
�'x���H��v�M@n�C4"��'(�9���iv(!���¡;P��c�'��!ĈPZ��O��~˶���'YʈX���}Uށ�w���s'��R�'zm�*�{m�� ��p���:�'�$�a �14�}��do��'`�Yc��ǲ!(��3��|� ���'�N�����9DQ^h6���hvb�'��-@�!��N�R<(�����'�4	@A�����A���<t�]��'���Z���8ږ�Z���s�tMh�'�m�B�TYE����тqll���'�%���ì#��tRB�5p�H�j�'X�@��d�+ ����%ѕdYAy�'�J�a��_+{�M���κ��'5 �;1gLX�4��cK�=𲱉�'�xyYӎ�:�F��V�k`-�
�'�n:EG�|��tb!,7�x
�'x�����<pN�9��C�{�f���' �R��Zp u24��:c=|y�'P|Ap�k�t=.��#��-�'(N����n?2�����
LVe��'�B-Ç��f�������00�'J:���
�}� 2T�`�'��]�Q�vD����	$�K�'誵ʗR��4���6HE��qN�({&n�Y苰"T�ӓQ����M�'6���[CKQs���N�^13'�@) ]{C�ݕ}}���Rf�)�K�-���z�*�_�.��g���QE	E�i8�O�����ȓl���؅Ԩ j�pG�q�1�ȓj�����L!ޔ�P�D�D���8�#��5l� �S�m��P��b&�}�T��&��xrc���p�P�ȓ|	�)��`R�F'2�qDȑ�[t���6�qoB& ���3	גfa���ȓk�j�B4E��[d�(��
�$�$��ȓ<�@Ph�`JS����-��D��d�\�zPdߗ����2�ϬM|1��W�Μ�����Sŀ)^ӢЅ�s�z<ra�2Me�%��g�Q�i���fśs �I9���C%(�HM��o9�4c�m��<���B��,y�u��DF����0<�`ѱ�������xM���=� �'Ö��vB��:k�,�2s��3Q�L�s�R
7��B�-'��Y�H�6B]� Qd$Q�C䉷��P;�C���M:��Q�Q��C�)� ��17��v�0Qrn���4"O��`�24�b����P�1"O��)�/:!ȁH��_�"�x��"On��r�U�(W��UH	d)>���"O�\4��N�P%���
66�k�"O��)��9P6����049�"OpI��ʑ�%ٔ}�F��*�Z8�f"O��O 7%��89��;F����"OJ��A���g�a�����h���w"O(T�A�IDl�oB� ֪���"O��#��_�V���I$.��]���K$"O��HG���&����P;�ȅy�"O��Q�C
�e&za��Fl��0�V"O�x����+��iA!��N >�a"OбC$�@*(vys��C����([��P�䋯4��1�On�ȓ� �r��:�p�i�g� �H��ȓ}��Xxf��V�,�QE�̂0fơ��\I�@h��meLhq7fO|���
B*�rf(Eز�A#DY&X���ȓDV���~U���g�8L����\��kȕ�p���7s�y�ȓhY�t���7E��kg�L�a����ȓg�PhB�N �&8����9��h��\�:�!J�*!F��J������CiKSh��mؾeuu��r}^)CrT�$��p����4=b���*���q��O�Ψ+F���ȓhb�H#�H<j��,�9��Y������7�͎;C�1�7�]WW��ȓ"py�^�A�e�T&P�z�`І�}:���"�;� ��V�ӪB\�ȓH�%��V�R�`=���%5d���!�)8�g҆;�� H٪N����?Q��>~@
�[���'YPL����n�as�@�z�!�B�|�xR��	q�,���F#q�" �w �&GZ�'�#}�'���2B��V(���D�BWvQ�'RfɢD�«5��ɰr�U�5�Ѐs%E�HB �bS��)X���5i��P!�F']P����j��z�@�64Uiရ�֛VÜ7O�X{�cȲH���B��y"��L�����=BN� I`�
���'U�8���o�b|���ӓ
dB�����38���j\W��C�IV`jA���N6�z3k%%=� �&ח|wN��,O����Y��i2(�
[��؁F��@qƥ�Ǭ*D��ru�ȋ;Ć�	�N
�1IN�{�X	Rb�'�Â>lOXb�,�D
�DBH�8�h(���'��C�"�f�CU�i0��k�Β� l��"$S7>��� �҇R��d�G��g��C��㑡z���rnP�ڸ'�zQ	Gȇ�=�*g�:
i��i��O&B����a�E/i�N���F��7*�'�J#}�'d�<��$Skd���א]��"K��Q"��>�&�)��	ՔQ�'����/���z,c�3U�́��j] ����AG��0>�����b�P��!�Ah�4tG@�ޟ8�JŨ���q���@P�y"I�l� \Z'�P�|*�,�n�ij�����dBQ�GV�<�H�'z��@�&@6��t�dc�
�Xe���ui2���H:^��`�g���yW��!ΐqxs�ۆp_d a3J*�y2�@�g��4�r�Z�q,����j\8	y8	&�-}�5*�B�O���f������E�A`��y��A�eO����\�N�{Ҥ\�����A�Ҧ���m٭X���`P$CQ��tc�oޫ[ܘ��N��@6���ݨ�P)��������%Ը��O��"���W?��B��(4��	��J�r��ӿ5>�p��8�zH���˟nLB�	�,$�mj4��y6x��冗4����ߥ@�fm���X^d`q�0.&��?�ϻ%Ҷ�E�ӥ8�����Y�<����9)B�	�,��Տ�8P�u  iY�"`X� p̓]����?1	"�%�-�
��q�P0e'xa���6f�E��I]p[&�%,��� �%k5,�#Z��"��~�T���'��)��nX����ڴ6ِؒ%(?V}8g�,�复�U�O5�h����s����ɩ����C�EP"O�=��O�,n-b�s���4g��i������������O쥉7	��w1L��'l]XL@��"O�0qO� d���fIQ"�5�=Obf�츧������]0t!���$���Zg"O����ϗW�TD�N�Y0t�0V��CQeӻ<bń�	<[݀���bQ,X�Y"��G�?�����Uy`��n�EČZ�=���jË�l�����''b��U�K<P�āiu���b�Z��գ9V�zV����O���O4):�ܓեL�,K�%��'����VEO��D���
;&'�A�۴Pդ��#���Pӧ���k4@���A��[|�\2�@z=�����Z~�T:�O��3'�ݱt�B����$v(�x�U��f�6Q��<�c�'�&��3`�j<���'�??�����y�g��=����a���ނ�ݏ]N�Q�E%8|(pC�Ыn�U酆�
��x�ƌL�X8��W�H������fd��4�%}�K ���1i	d'��'(��,��$��{
�3R'� AK�B�Ir
:��T��	$r���PI�7[�:� ǀ��O�d�Xb�����I2����.�s�L9HFQ�Jl��-�c<x
��'n��e��f6p�'�n���л7��ă�'I�>-*O��C�*�&��dƛE4��i2��1X����S��\R�,�t�+5��m��V5!�$FE4^��Շk���t �$UZ��$"Oʡ$�&u���c.��CA�9A#}�2�3}2�A�8��t�>E(ع�d�)\jx����34��@b@
�l�0 U��(�a�(& �HA���a}�ù4�dq�S�H,8-�1-÷��<�s ��K+65�mC7�y��� E�F���i�?<����f�lC�	D$�Eb���T9�d@�*m��1֕|�D��(h����ʢ� 5D�����-0x�h�(��-<-0�+U9�y��L�\�Nd�K�<��bN?|���JD��Pd��M(����L<Q$��.D3l����7(j��q��\xH<��Бy�ah�Ë���@GAR����%�0�p��9�p=�C�7E���5�̤D+�59FRW8����-0���V��,KXr� �M�J�֡k�+˵5�X��DeF9!!��ݢ1H�0H�p�I��φ��`������
�!leZaàY7#|�Mk�th+�'�7`A��q�\�<�'��!B@���)Ǫ?"���C��y	5rtU~�t��#A�	;Ľ�|�K>1��a��(�C'ӡB(r}�s	}<9 b�@"�=��H�n�L��^v���ƨ�!�
|8d���\/�d���{x��[�"?���mF�>��QKU�7�v��+�k5��D��M�;[�\�РnE�pZ6p#!l�+g`�ē�FْP��D�Y_�D��jZ��Ț�세c��I�T���%EW.a+�!e�[�+J�QC���ǱR��X�56�"���x!�$�2I�����˛n����)�Vmj��m�(���ٶ�!	���:e�~r��u�	c��*��;d�|��"��_Ê���ױ!�qs󠓶;���b�`T�Xqr҂��2*M�c�,pR����&,�y����k��h؃�؞{�1��N���O���ˏ�;����߁$�`�Ii{�Ç��P�ǎ�x&*pɒG!$�8 q��#2��iXAe��z.��(���ٕ- �K�O"BK�x���[�<��~��L�
ݪ�l�k�T)ȑa�J�<��$]��x���� 4:��hB�U���$|1ё�A�6��ܤ�z��c!�d4�Ȑ�X�,nNt�4g�!5�~B�ȌzĐ��R#R`|� CX�c=��y�F�^�"-u&�
3C�UA�^UjaybB��t3XAI��tF栣�H�,�O�bWc�g|Jhi7�N�(���r��@,wY��� ��odnDbw�/�la��9$�,�EH�r�ʬ��ߛ@F8 �G��>Qt��.r��*�=����dջAc^��~2�d�SKt���DK`b��EkUg�<Y��R'. =��͇ "⌘rfDG%$�(y����)�p"�)fGp\&?2�x�J���Z$�0��	WD��G���y"*�?Z���-��*��`AVH
��?-H ��m�(��pQF�'�$aKR ��o�ژzAG���T\��DQ	V� iC��T�YU�P�C?ym���a���y
� X)"P�c��zӠ[+��0�`"O�ٰA��T�X�HQ7<9#�"O��Sf�+�D����{�!@"O@�ѷ	U��ؤG�&Ci����"Oi������E�Z*q��"O�yB2B�WG"�;ҏ�#dP<��"OpRǫ ��)2��?�"�"O:���޹>36����ǳ|s����"OƠ�P��Jzpx�TfX��ٰ�"O�}���];B�q0b�rn(���"O���&�\�Q[���ЈC�"9%��"OB(4]nZ�BD��r� `�"O���Ğy�%1��A�<�B5"O�T1��#[*z-���}�mhg"O�Yu �?ID�7L٭qh0aS"O����喃.�tH�CkιP��*�"O�(s��4�ʴ9��x���g�J�<�T@j���em,jL@�#ɏD�<��R�K06tYBL�M�4嫢BX]�<�#)	�.mU�@�z	�]�VDF[�<a�#Y1:O4���&F�e��Hs4�T�<����va�ŪG�M
K%�ٕ@�N�<��]�ZTt���R ���0�C�<�cN��qz���_Zv���O�}�<q�A8TJN��\<a�Z`z%m�t�<Ѱ��[m����>&@�BFx�<YR�ٳs�QR4�&�"$���A�<�6��L]�M��+��;d�=����~�<��of���ўo��A-Z% L!�D_��N���N�C,ess- �!�D�+|�q� S��#D�Tl!򄌲 E 4��.{	>��pB}C!��j.Z�I#*� �.����3�!��X6v�h�)L�)��Y�d`�	U�!�D�6t��� م�G�6�!��ű0��;a&

����,�x�!�$]5l�ȕ�$�_�v T�᥋TLV!�H	8��Ӈ)��@��t� K,{S!�Ј4( �q��;ژ�X ��h�!�$ױy},McuK�9;���G���%�!��� t2��q��dϰ(�����-!��zB@�q�
y�1�P�#2.!��BNH<T/,W"4ӑFϯ�!�$�w��4���0M��q"�L�A!�DP` 40�	ÚO��p�@T�|�!��( ��p��%O�RL$�1�!��_�Q*͒��ԙn<ĳ�lXV�!�Dԕs�8��e�\�}r���"!֫q�!�Ě4\�X�ŭW+sP��"C��<!�H�@�r,2��lT�lQ?(!��ǭr-¸�6/�8s�}� �T)Q!��!o�U
��]�9t�ST�k\!򤛁".�bզ-xzq��N0A�!��7r�@���9l�v����k`!�Ą*^���*^��IR����a9!�D�(h����S>4�����f��v!�ď"9u���eϓ�{�a�7OΙiy!�ʉL���d&թEk��3a*x!��'}x�S��	S�m)V�L"k!��a��s@B�d�8(HӍ�0!!�D>9��l{1��{�d��˷e/!򤚣�������+ngv���(!�d�$�`!��_�������p!򄆞:��Aa�*K�a��T����)�!�� i@����bڎ�c���5W�X�"OJ�$�ӒB	\}�'B�*	�	!�"OJ|zǦE
/�9AbE�`:)��"Ob�e� ��$�獈�a�"OА0�^5p,�`c��12�V1r3"O���T����Pl�֮D*�"O�l���<�v����!_`"@�r"O��u��#i��U1�S&m[D�"O��p�m�Z�Er�[� 3����"O���sm�,�  L� ���"OXi�@I�i=n������)s�"O�
��n]���,ܜ;Mҭ�"O�0֨I�*qL��᫉ 0���R"O(��s��3kb�SVLޞs˞u�3"Oh�1e��1��ɴ.��x���c�"O����ŭ:,��LɉT3 P��"O�����Ԍ~pZp�'jBl4X��F"O��0�. -0n�H�`@Ts�\%��"O�d�%I�f����1QR�s�"Ol)P7�փۊĘaK�*��豀"O�� ���5��бl��G
P� T"O.%Ѧ��xu�j9p�6��"O\�X�/��5�М*�
U�����"O.���#Ú�c�H�<HT�9��"O��[����U��G	������"OPT�h2]\�5�R�� .��u�w"O�p�'�-cH�1e�>0��8�&"O���RI@�jst�P%���$��"O^�����q��Q�&\9�
��`"O��������hU���*=:�"O���%WrQ����?���R"OR�K8ER���Oj��E�B"ON �M��bapE�R8'�1�`"O9��&V1}��ʓ*_	̩��"Ox4��D{
�%�u��jmHe��"O�	A�G<V��ʄ`L4�\�1"O�)K�C3
�X��R�|�"OY�%��J�2�q%N�>r���Q��ޜU=�(�Fk:�a�"�t�#[���CJ�]u���ȓhE��PE��!mش败�8P������W�V(J��3��Y��
��V/n�d��-$ݸ�#��)D�4󖫉{D��6�t��q˥`F�o������8ju:(C�ƀ�b e
=o�X����t�N���	���Iy�l�W"XoZ�]���#�g�F}-�p
T?�C�	zSt��rAQ�S�Ȉ�c�νF�z�Й1�_ I1���ңMU�O�D@��#$.�Q�V��`�	�'7L|��;�-��_����C	��`��<qW�'�gy�L�)�r`�,���akǽ�y���sB�6�q�C!'U�8EסE3iO�шA'!lOL����� ���b��1(��F�' (�؄#��D�	ѿi�����k���ۀB�$"� ��reG�d���f���KV�H9���jp���'EZ!��O�(�� 3��Ӕ1 ���Ra���Цx��\1S�ވ|�'��"}�'޵�E�Tq� `쓗ꊿTL�hP�bVPM�Q�O�4�}���
�UO��ɏFSr40f���1����A�_\�`�ǂ`at 3��1�O��{VO�Fnx1���� �'�p	{D�"��@��[f/w�x����� 41��ѥdήh��ϐJ�V��T"Op`��JOQ!��z��]>1Rx	�FG�	��X!E"���;Sņ�&gd|���imޭ�\K+�8q��?[f�[��-D�l[�¬3`�Yx�he"�oR��Ń�z0��0bC[�?u���C�'{��G��1N�p�hQ��^ܑ�Y��8�mD�J~7�3z�I��F��m��q�3��+� ��Ǚ7a0t��'��",��p�C+o�;��Qq�`vJ����G/\��5U�pA�@����i��15Bˑ3��t����
�y
� �\�Ҏ7���`�&�$6GƉ���)� p!KΟLr#�\:یH����{�혅m@ ���YTޙC���%"7D����	�1vޝ���_&^AN���aY:���0�\�8�u�'��I�	2~Q��I�*��8��<�@�Cb^����+|O�`D�+���A�4=)��S�Ŀ
x@�AF�*_�8���<�H����'���Ԡ�?+u��ِ��O�H���d�)s�\��!�'S4Kf��t̓s��h�P�ȓA��5�����Rƙ#��΋1�q*ܓh�.�=E���!�����|������[ */�D�ȓg.�R��mͬ�a�gQ5�Z�ϓ wZ5���*�)�<�@�4��/��1r)�贅ȓ^ ��HF�9_+�e2h��;�<�'�x��ƭȡaz���2+�\Z� �gU|��'�%��>��^�II�Y{s���v��1$�x�H}0-��r4B㉧k״�pC/G�(��� Y�P�4"=��ӷnPD��a�7�S�}��$ۥlX�'����e���C�P�E�� �0a���b�5*�7M�0+� �q��S���)�禅�lԇA���,
�Mg���� 8\O�9��-S���̥]`���b^_7�y�S;|�������q�
�"��y��O:{��p牿�6�;���$՘'�2�� �%T[q��	y��)+v�%p�Lۜ7`�a)��%��Jǌ��xr�'.�I!�+�S�n���\�6piʂ�=}��W�*n��d�9*�v�'W�条U8	�$ϿP�
8C��K��B㉇x�YW�J�!�q��QPi�t�ǁ�7w�pN���I;n��q�v�<�s�������ɳG ȋ2NI�G�'��㇠Ɉ5DA�'��lpt�_�0��:g(��()�)O� fHܠ^FH��On
���U��&[��)s��'/��'��y�"�$*����~�։� ?;�)��Ҽ(6Hq�%�����K�b�^�<����Fs\혗 �-,�t���mQ�Y�d4A�>��A[�����ɮ�<9k��d*n��5 1xT�B�I�O�XDc����iBt%K�[\H۔��63��)zP�'�N��T�X�_�P��SbF�ClMH�_�Z��#��2An�:�Q!"�'4$�Y7j���ȓ6�H`t͘5����U-IV��<�u�D�}L^�`��I�9���{a�%
f�QI�(P�!�6Z����
eWF<�c�"\�L`�E�$���(��ɵ�൒��qǸ��KR/�$C�I%w*F$yu���)��d��U�yn�B�ɑ@��4�q�<NX������v|�B�I?n���e���d=�P���&<r�B�	&	 �haF&_(u3�r��4��B䉳'0|pz&k�ь�B�n�#jw�B�	f��p� ȫIYZɰ�۳s>jB�Il���w�-h8����,)�BB��;���p�!��q��Q�[rnB�I�u���R)I��| ��	R
@�?��
٤%w.b?�"$0 	��Ď�Id4�:T0�!�D�P��y��I-Wݢ1��R���-I`�r�VM�)ҧ�f�QO�^�yi���a��Ȅ�NBD�+�$Xl�i���F��T��XC �zc̋�W�-��*�Ԇ�W̓n��a��Q�h��`�eY�l^����	h9��'�ɔD2���L�5_!���L�Y��Ti3O6Q�E"��J����䆈0:H��qBRGz<"�)C�#�Q�� ��U�+0yX��'�6 	�F�3?4`	!�0b$���m����CVH<a&
�*F8ac�^;]��=�/s?!��[u���ꇯ�O�!#�&���!��D�<1@a��G�~ æ�Z �yҮ����&
� ���pjچ�?A��K8m��
b��	������RF&�%��Q�
7*4�a�Ad�H��/�O����/şS|�|�GY�PE�uA�Ж5ܔ�Bg�6�?D��E� �-,Ol��H[.ZnU���W�
Q�@ؐ�	?`����!$m2EȅUt�C�W�eS`h� f�`�p�r����Y���p��@��*�#Ohz �'�ڐ�-T��D��|�8��)���O��� �C�=�F��fhK" �b\��'�U�F��`�,|i�KNEFQ!��i& $8F/B�d���qD���'f��O� ��he�&n�tC0��1�]�P@�ȓ:p"ɥ@��<�HÁ�%�'���Q�����y�K�%,���r�n�$$]XĊ�p?	�"X.t����f���n^v��e1j��pc0D� ��S5�2��F�J�$�{��1D��ŭ��B�n A �H�.�8Ċp	/D�ȹ7!\$��a�gㆥ�����h9D��۠-L.y����	܄��3D��"�ڍ=DT4���� ��3�)$D��P$��9&ʝ�Fj�)jpn&D�ȁE+�e���EyH��#e�2D��"�
�5�vKƍ��GȰ����7D���PbI�^��|�s�;,`d/>D���t���J[r�@.Mf@	C:D���'��w�|�2��@�Q2��7 9D���FbBA� ��۔>� �2�d6D�r0� 	(D�{A�/o�8�:T�2D���0bI�b� 8���$��-Y1�/D����Ձ!�`js���y�D%��7D����b	# �iv����#P��yB߽o�A��h�8�c`��y2�Ͱ�v�����ݢ�F\��y���]�|��! Aj�t{��J��y��<C��B�-˟Dݘ`�휨�ybm&�P�Fʀ�1g��`�@�3�y���{�p0�q��!����W���y�J��β$C ��t��'�0�y�c��b����A�RT��CN�%�y«�7tn"��@�[6����Gȿ�y��7Q��#��h��vh˒�y��^��N��&�3�)�E�(�y�F�X�d]�A��k��3N� �y
�S�v�(�JW��Rd�f�Ѧ�y�*�x!���ɒ�L�8��.�yr+P!!��M��H=mLp���yr��(J�`�	W�2pڊU�f�2�y"i�&ߨ���(����= �@K	�yRX;��-0tmo�D���*L��y�(��gP$\���W�2��\��'ٞ�y*� �6��E��F햙��g?�yR�1��ᬚ96�X�sWA��y�D�U/.m�+�*����N4�yoR�n�Y�l�	EFO�e�X�R�' �����іI�������3
�'�ZD�R&�9{%�9���ׇznX���'�
Þ�J�x\)�.��{Z"�:�' ���܃&`��).E�t�L���'��I����/"D8qF9��5��'�,I�@%���F�*;s�4q�'$�ya��Q8F�0�5I�"ff`��"qT�4��V�����SB��	/A��y���*� ����U
N�:T|EFx����1i���x�f��Y]�5��H�H�!�䆲y�^��ɘH6�,��d��g/��%�S�O^`�se�@�b�@��1$d���'�0<�!uf�P��eD5C�>!��IÉ��9�5�*^������L&D�4��O�ӧ���L�閱(Q���.�-R1Ξ���A������ݻćٸ*��`EW8>=#Ճ��e���#�'Pv����O�)�\�"}���J�xI�˝�?�l��7ʂ/atܨ�O���v����?ӧ�)�)Y�lU%���=P\ �O�&s����<��߶�y2��m�OA���B�N6~e��0c�ߥp��`�Ĺ<�2���y��:�g?�����N��	�V(�;��(�O�t~�p���=�O�剱舘b�k�jEq��$;���ɩ�D7�3�)�'�a��h:.k2!8�X 2K0$�qkQ���뢖x�O���G�� �x{0C�xȄ� ���:omԉ�����0/�p}�f݈M@a��@���4��'Ǡ/ۜpp��!A�=�Z�x���Ó,�&>	֧�i�����֭lcJ$:Să�gy�듿~���3��E��'�{�Γ�>%S��"�3�'�>�����%	�t�h��9!�/^�J*�ĉBj������D��R��񢴂(����0|���ޡ3F$�
tɈ%;��lх�A-_j�2sd2?Ѳ+��0|��i1;Vi0�KA�q�4ܑb심K���CՆ�M�%.�;S�y�ç3�b] &cC�`N�u�'I�$f�h�2�	���M���;N�&͘�LP���Tl�F�Oܤu��OE�Y8�-K%�$3W�9��m�~�V`��c�2TC�E:cߓ�~��I�Sm,	p�P�\q��re�K��v��# �O�?�("K[�>��m���K�A��ݠ���"���Dכ��	V�,[�{%"��9�!��0� x{�Z,=B��3o��#�!�dM71���&Mn&u�G-�'|�!�$��q6�l�!g�2v<�L�1I�:�!��:����"P"4A�
S�O|!�p%�yG([4p����f�-_!�$M
-�������B�U
b�}��"O`]����a�L��3LE��W"O���L٤_�.m!�+A
[2� B�"O��A��n�.AYGJ�8dya��"Oȝ��ξl�<`:S�J�>i��cf"O쀨f�0D��`i���iM6��"O̥bC�M5��	e<5R"(T"O���&˂Pbia�x)*-�"O��3��=Tnd����Zj�Pkg"O �"��F�^ł�@�lK����"Oj�Q�$ѐw�(�8�"�iK���"O�ȵ/�4C3���a�'	=fh�"OlF�=N8�a��ю|~��"OZ�+q�Z�)�&,�2_d�9V"Ox�ÑÍ�j�Bc��4{:J�kF"O:刁ɘ;8,���*�8.Xd�g"Oѣ��^�fq�p��	^]HM��"OE��9�T��&�Z�unD �"O�KRB�$w�jh���ڴS�|��c"OZ�K����{�8�'�,%�ػ�"O��
��l!�s�עt8�p"OP����͉&��rR�Ξl� ��"ORHñ�߷JŨ�5Ér�&@�$"O�9�`Ӫ�ʁ�s���q1�"OԽ�f���L��QQ0�� Rč��"O�Q*�%pJ����� �BP"O@�j��M�r��i�.V�%v��"O��q�a  2�vĊ`�M�2SPm� "O��BCQ��8�V@]�&�*�г"O:���A�/��
wE�{vظ�"O�-8��[�[�����hR� a ]��"O6�Y�f��B�@�;BN�\�p�G"OPk����b��
��%�"O�چ�U�*�����&��=�R"O�Ȋ����^N�18u�V'M��`"O��K�oK����Z!c�'Z���"O����� O��bV�U�E"Od�r�x�����L�I��l�c"O�L�t�߀`�Āh���p� l�E"Od��Q��V&PCB�?��X�e"O�z��:I�l�C�J�UAV�zv"O�4��+I�;��ĥ��u>b43"O��1�O�{Ylu���U?`��"O��rI�h��Y��A�K7��:�"On��*����;K�	eSP\��"O��˞�jO��T)	"
;�ɂU"O ��d�"qrNH�C��-�H��e"O� `D���R�A)�A���Y�"OLMːN��qARɠ"� �9]耹�"O�l��	�7mRp�u�Y�GD�5��"OBE���6�����'8B��iv"O��K���G��Q�3HJ�C�%�S"ON�ò�>P����D'O'l��["O~�@�DI�E4�GC�@��4Y&"O~�D�Ρ:`Ѐ	��R��h��"OЁ�҄Yz�%���J�]C�$�G"O�� W��]0+��0+��b"O��z� ݫ%(��4�_4\N�B"O&	���J����C皭�!�"O�a��T�Vt�G��$�x��"O5[�h��65�u�� :T�
�"OP��pj6�\qA��ȸT���q"O�	�:�X�*V�F�U�����"O���#��(+g0���F���ģ"O�l2F�+H�(9" \?��t"O���vD-��Ts���)�d�C�"O6�!�@���FDg4���"Oz�#���υ�A��ɓ��'O!�Y�D�����H��H�s����!�H r����Ո1����c �;=�!���3\K��[�Eot��(�
"!��B��q2�Ot�l�3�eS�!�$�$/J.ͩ���/�N���%	!��.mL��b���E�Ā�4�!�[&]��I��o�;I�z���.ہ?�!��F� �gkC�laf���,ݰ�!򄂑o����'�F�d'�Q��K�*_k!�$_�w- �׫|�>�[�j	�^�!�U"Zw.����߭b��!:���&�!�d�)��P�B��e��L�]�!�$V�
+j�a�|4�D�'K�!��>F�r8��֟/o�%!s�S�p�!��(:&X�SE@%[���$Ι1�!�$' CԡgulN0���?L�!��Q"��"W'fQ�4q"JBK�!���������j9P��U�	�cs!�d�%�&h��#�o)p�
�B�6!�Z>J��uc���/=�ȫŌ��R1!��X�� ǥ	*��a�X0.!�ďM� yZ���Z-�SeѾ*!�D�GP��x��W�O�(Uy�dX�g�!�D��Q����j�=�Zz�i��	�!���$7~��'�/:�=K�E^6n�!��w8��GJ�L
m�EF��!�ڭh*R�#�ǊZ�P��
�!��*D4z��A�C+��c�\�Z�!�䖬_���6�ؾ`�nUAw��n!�$B��� Jve��w>R8��
;!�i�2���D��8'8�C��4!��Kg���P�Hq)���C�<�Pyr�-�{�.���x���]:�y���#,&��t�sj_)���'q(��&�^h���BfA.e�u��'��-�5JϚ��EЕ�a :���'y�,s&)
�r� ����ӌ���'*�#&Oȉb� �JӢ��D����'������P�l�0����N�Q!�'�tC����4#pBwy��z�'TƤ��"	�+~�����l}�ժ�'^��C2��U�)�ի�6?�e��'�h��iW+'&VyXT�F겸���� �`x����$-�=	��1�p"O�D���H��T���~b��""O@���ψ�S�% we��mk�|�"O��竑'���Z�@�
�$`�0"O��	p%ى�xzuC
�SS*���"O�(�V�L:xS�q5�A66�p"OD�ca���J���Eoɺ2RՓ$"O��e@V�g>`놏!nC>�a"O�j��Y�8��XNK*(8"��2"O�maem޽|vP@쎳'��D"Ob�"�A�`��z��֐�"O�E��:WJ1��	ݮA@"OH(�� A_����� ���3"O^!Ja<_�Ly��HH�l�(a�B"O~��gQ�漹�̗(�
���"OƔySj��m��:�	!�n��5"O 肂��g\A��^	�δ��"O �J�%��x{*RDS:	��'"O�E��c�	R��8k��Ƣ�4M(�"O�Aɷ�e5�5�u ·.���Z�"O��� �R?��Iwo�m�*��"O��H!�ݷ_�XK���
��5"Oz��4L�:J�D�C�M�<4&|0۴"O�Mcŋ�4cѾYG� (_�$iU"O0��J�Ex�� !L�x .剗"O.��v�K�>o>y��T�� ��"O�5D�5Y�b]qJGw�H��u"O��0���0DDK���e5~��"Of�C��  �&�kD�ʒ (���r"O6�R-�8j�d�;���r�"O�d겉�sJ4���R kK�\�"O�Ik��&?��ȳV��q���#"Od5Z�*C>J�����7E`P5�B"OPC�`q���BFA@���"O��K�N�_�,FS-U�"O� BQ�B�,ct��E��##"�!�"O��gB�2�2	����;#4���"O٣���,�4��FØ�v���{�'fX0PTmcY�}�Q� �g����'@����J�A�P��9-F
�ʓnHpV(�Wp�p&�94zԅȓw�Ղ3���h�Sp�X�(�t�ȓ	������}�ҹ��j��.�R �ȓ{z�Y+@���[�J
���W����ȓ��Ѹe��*AϚ)��o�A�� �ȓ~�a��:+�TE���L�0��X����'G�=1*�s�LW	#o(pa4D�x�7"�!Ҟ#�Δ�V� D���,D� rEH/`��]�5%Ѡt�mk#*D��!.-Ʃ��&�8�v\�p'&D��hש|�r$��,�o�yرe)D���e���/X*�4�I�l���c�%D���C+��Q3.!�6჏WA��(a�$D��R��ϰ)�,41B�α�p��$D����
�2Ek�Xi#l�7'H�L<D�@��pm�tS7��!;tY�A�4D�T���Ϡ_&�Q�
�%x�AhT�2D���Dd�
�=S`-J�D����3D�@)�"h=��%Up�4Bu�;D�(2�e2m��F&��5K�,D��J%�G�[��JFe�6�
}z�-*D��"�D�2�dY
Y�e�0a<D�t@ K�b��#�Hؓvx�z�<D�<����
�"�"�=FL���,-D�� 6��f��0���˲i׊��5"O�L��G�>zܪU��.Α#i0��U"O���A�,<��dR7q2�h�"O$���+K%>�[��g����@"O�$���Ġ-��QrA�f�J�x5"O�-x'ܺ,�PI��gD44yd���"O`)�LG�1�&�as��ah�U�2"Orm� ��8
~�0Zá��[�"OF�i���8$��IRAO(TP���"O"dĦ	�|��/�"<-��"O���e@�!>^�X-�"8�A"f"O�L� ��!eln�"Gl�k �X�#"O����g�3��`�u��=�*��P"O�!(����]P���T 9L�0�"O���cH>w+͌K)8��d@O�<A�   ���9;��)ࡇsªD�g"Oz0���x�� �w�T����b"O�(���K=S�ę�0���8�B[�"O�`#� @(?b������o��0�"O`L:R�m�5J 6�Ƅ�a��t�!�dڧ[q|u���E/ �!��_!%�!�D�	0�J2 ;��٠'�Or!�թ��:���Ҽ2�R|�	�'x��xǈ�1^.EK$��t��	�'� "�щ"ш(�Ԉz��8��'L�y���0���F$T#� �'F��Qd��)F�+�%Gz���'��8��\�8�4MK||��'� �f�ٴr�X��sLۨC:@M��'�VD� �ɇ5���3��5Ū���'�tEA�ڳ9�$+��J03�K�'Xx���;?
���flQ�/i|I)�'� aJ" ��z�����/�|0��'�4 ����Nq���/��\�
�'V�J���~\����oASGNU��'m%X�*Ǔ@�؀�(�:D|xz�'�ij�j��#?������9Rʕ��'�>�yC�׳+My.��9/�'���X6�_�X. =@2C�14.X	�'�~�c֨�(룇ݘPY�� D��2��O2���� ƙn(xȕ�?D���	/g̨[��ǖ��9���;D��#�B�O�t\s�1s��9yb.D�� ��:���-,`1�' Z�x���"O^D�� R�|+B�)"&֐#��Ԑ"O��8�c�>�4U94n��c~ �"Oj`����������K2_y�s"O2L�FfϡS�Ru��	�bxPP�a"O�X��*�n����.W��T�"O���'��a�Q�0��Fk��R�"O,ţ�!�$"���rD ��KhL��"O�uq��k�Dh�aT1Q�ʷ"OJ(��Ɂd�p PD�NP:�� '"O�`����?fEl�!f���O
���D"O^p���D2fP�qłBܬP�"O�h�a�7v�V);V�����Yw"Oܼ����/C�Vhi"IW�e��p5"O^ś�L�"�+$H�B1��"O�8'D��ڀ3T�R	l���s"O��͕^����+,];:U""O=�'�1i��+�ӨO�<!9�"O0�2pω�}o��j��^�yf���"O�	�CfZ3t��	�.�8G�蝒�"O��ǅc����X�ߪ���"O¹��eMd��vI�f��l'"O��vg�%N����ȓ� �!�W"OtQZQB�]-x��1�N�of0r�"OZ���c�
y
��^�9qȝh�"ONd���*5Q���I.2`P��"O"A؁�ʙu�����h�`���"O|A����4Mq�\�e舄:drh��"O
��p�F�]�hiT�TR�
p"Of��#	 �t�!#e��{;��["Od����X�_d�!�u�� "��I�"OD�၊�H�İa͖"��Xs&"O���H+��d��E�.0�S"O��at��!��X;Q��4^�J�s"O�T�7v���x����""OV�r�.ܯ"p�����.����D"O�ęA��9"���w)�v�� c"Of� �(c~D�P��-D
�u�G"Oӳ�ŢJ:( ˱,U L2��"O*qpfF<I۲��,:]p%"O��� �>�9��.	��&"O~��GA��~B,K�i
� W ��"O ��u Kv�B*���+17�c�"O���S��i�@8
����a4F���"O.9����>���5՘	8-��"OD�:�e��P�@k�G)4�"2"O�m�q�ߴhbZQ���=g#��J"Od�q�L�-��xpq��x�t�"O��5.� ZJ��J�m�XyT"O���A�9}�9��
	82�؂"O|)kFf�$M�(�n�- z�|!����hҧ��	.���ۦǂ�Or!��ѹ���ad�*o晁�Kr!���|�dM1Fm}k�� �*��z�!���KZ�B@H�5���b�*A
f5!�Ěr��](���u�$�Rw��yJ!�Ē�ZE���.wv�=J�+G�9!�$-V�Re��N�X�H1�.)�!�$Z>k���v���"'�ܛc�!�*b�j���
RI,� �A4!��p�����I1Z\�f�Ч/S!���N��$�`������@��C�'�!��N�w�����!T��ĺ��v!�Cd�k�
A�G�J�a�Ϣ�!�� �H��p�h�[��yd"O"�x���-{�0JGaRpxR���"O�S��T�zt�(��v�L��"O4Y@�D�^D�s`���,���"O�|@Q	 
  �ȓ7:
`�CC�x������^��ą�0���Y�H��=�L8�Ǘ/�d��ȓF3�8
��g���J#ْX���ȓ���઀�f�@�Ā��W�Ƙ�ȓ?+�<Q2,ܡMv�M�5�� |>��ȓ=�&q 򨉺݀%㣋޻�4ɇȓbπ1���]ސ�҃�H�Pćȓ	� ��M�4w���k'�9B^��ȓ>��L�e��fB�6`dq�5�ȓ�(�:UAֲ.���2�<V��ȓi�Q����~�p����r� �ȓ5%��� �Q�4[& �2�J���>����Ci��VM���AO_���X�ȓQ}.D��G�c\�2#��Bx���ȓX/��/5C�$���UO�dh�ģ&D�����Ɔ6W�<�dB��$��2�)D��т�_)d��7�6)el{��&D�����)&��٢B)<,8"U�%D���"�X,)�((���-)���#�"D���#k���1;�@H�x�l1�f D�L)��.}��j�E
&l$UHԫ=D�Ce!#.Z�#���ɑ�I:D���GK�f� ��S�]�4l��	�,D�(��i��[e$a��o`��`�5,+D�TA�J_R���"�\�6����b)D��*V��i�d`I��Y���D�܆�yR]� ~�ӀK�Q�^D�F���y2����8���^�Q�ڕ�B��y�5'F4�(��=����D�
�yb��%(��Q*P�/�>�qCL��y2-�3�Z�����'�B��%�_��yrj�9Q��0G*ϼÄ�j�㏋�y��
f�Ҩbp�ջsHL򃏘��y�(�(y+րp�e-*�h�
� �y"E 8�Tb�ռo��m�
�
�yrAJ�+vX����a-
1�E��y��#�����d�Wd��ť�y��*(�8:6C
9E�h�$��y���\-���ԈX�'����@W��yR��� N�����\����z/ �yB��B��<��cJ'M@��q�
��y���Y�����>U��t��;�ybj��N��q���ĔG�"x(`& ��yb��0��pk�A8>H�y���&�y��-H� 9Q�n�C�q eC��y�=A�������j�X� ��ybD �mJd�H��Y�W���a@D*�y
� ���Ѥʀ
�q3E�	{�{�"O^��N�?vGt�Sa'4}D\�W"ObUyV�@�RKv��Vȑ�
$�)2"OLr�'�9��̋���z���0&"Od��O�jf�BO�+lJ�"O�Qbd�������.b�2%"OΨ�WNO>*'�,T�9v�����"O��3��D8� ��$.	q0�B�"Ol��ǀ43�e�4c0H �"O��B�^2d�U��\�f�~�X4"O8�
�G��Z���T�U�T`8q"O�`�Ѫ�V����e+B�{eйY�"O� ��d��)Ĝ��3醍W+�5�U"O�P� �[�xI�d�˧,*��ذ"O�1(�d�B T�x#�Q�R!�YF"OK���Wy ܣg�)336(Ҧ"Ou�bi��:�D�M.���"O\�t&�X{�� ��5+^��Q"O��	B, J���,g,8�'"O*�`�eG�J��}�d�,�d�C�"O��s�iR#,`X�ZF�Is����'"O�來�TOB��
I�Ѭ��g!�],v���������̍Q�!�@1>qM��I�[����FjO�q0!�M?;���{�O<q�T�	��!�M�X H��ԉ�0f�ƀ!6��*�!��ݚv�@�p���%�zAaԦ��<�!�dĄ�����Jw-�� ��éx!���2�:et��&H�ԡD��1�!��X2��o^)L�,hH��2!�J� �x�Z�5Ѐ)iG�1'!�DB�}�H�� Ƈ4�pU{͛
!�D�ch�k� Y�S��{0�/�!�Ā�	g$���g�.��-��Q#!�$)=R,aP�-̀P������!���1���r���l�HiQ���!�$��R��%y�ʍ,-���*Gk�>$�!�dA;�2�QS���l9У�M�z�!�d�	��Q�c�8݈�P'�Q��!򄐌6���'eT5'2t��혜^�!�$Z�/��9�G��ZsReӑm֑F0!�B��\���蚦)Z�d��ŕ&3!�d��%���)a !��U��Ŏ2J!�d�A�<YK��-�f�fG��T�!�	 ^�0#B[��9"5$�/|X!�䙊B�f1��j��]}%�fA�I!�F. �@0cT v�у�A�[/!��N�r�A b�i�8��l݆-!�d�(xu�׮Ov���-X�!�J�?��]*��\�r�gT!Ux!�$Բ|���`�=w�<,(�e�*�!���Tꆍ�TC��n��� e=\!򤘿G�ŋ��_�VK�x� o��O!�_6���ꄊ��U:���c.F�
�!򄏫"1�B!�/r�<=��,��4X!� H�P��Ah�pn���K�&nW!�D�@ 怪�wXhZFT]k!��	K��1Qwaȫp�� B�67N!���Msp�S6U�����*~�!�ĉ�H_��`c��%�N%�R��=4�!���Tl�y`�B�}�.a��}!��#�@�����x��lh���B`!��S:QWba�����McU�=hK!�"`��[��7X�HA�W��'>!�� ܭ1��Z#AV@@
�9C$��g"O.x��̓/;A�
�HA>y,,p�"O���� jI���ӜV]��"O�D��cS'8d4����ݻ53��D"O(!�O�7-�C�C'y+\�ْ"O*��
XM��M���X8p�#�"O�}�%�FLiv �w�;���"OV%�B��	QA+#���{&mP"Ov ��ִp p�M6'�会7"O��sff�jP�����1c��"O����P�>w����-��Jh�!�"OF���֦+߬��7��1 9ry8�"OZ���I�t�.Ua�,ʵs�4��0"O����䛍G0\����/@.F�#�"O�Ɋ��X.Tb�}��e�X�x� F"OX��Ċ�t|n�Q��%)ϮY7�'Oў ��h��eF�CQ�N;\Lv�h�J4D���K��<�H!B�R��DI[G	1D��*0 +{Ԇ�{�%Oi��y�@*D�<Qk;(�<��%�5����B/-��p<y iKv4M���K!y�80�&\W�<YF�=��pA�	�c>X@�V��H�<�q��j��C٣����+[`�<Y�������!֣O���G/u�<�U�R���+	�qC��¤�Rw�<A�Ί+
�$%��̄�8qZ��t�<��[�����zn>�+��u�<��F!%�Ҍ�w�M�D`����y�<97c�$�2�ja�;Ev��CI�|�<�b�G�rM �� b.�ⵘe��z�<Q��1^>V����Z�VC`�8�Ɣ]�<a�k�U��y�>=D�S��	B�'7ў�'Wʖ���%8��ˡ
�<o|���ȓC�>�S��X.4l񄅻T~Э��;���y�I�<��ā�.iŅ�Ic�%5�(�%G�-{��3�I�(3��E��R�1��޸�l��b�I�L>���ȓ0V��ړNH�e�����W0>	��-�0��ΎQjK�lZ�/	(��'������" Q�x{�͂��\��L����LQ� ��m���5:�X��ȓ�&m�nSQ:N���AB�i���ȓa@ب ���}�V�1�U5.��A��($0�C��ͤ_�Da���d$���j�r�82��|�4tp&ӣb����8"Ds���u�)�(������&��8A+�.q�b���͚N�lM�ȓi|�y��^���"`і:"��ȓ����KJ'_j��p����5���u�������'tЄ�M����$�ڸ	�^1-��5@�g�1����q�����M��W/�)o�q��z��"E�T.]��G�(�
�ȓq*�eH͏7xD�s�� ^Q��ȓ[�8Mi"�3){��SV�;C<���+�����8tr�	�clO˂#�[��hO1��Q��o4pur��ŤN��� �"OT�A���l6*���h�,��a"O6M3�kޢ]�*� 1G��X\�"O$�p�(k�"�¤�8���!p"OB�T�ح�క�+�P�	R"O�(�#n�1;�T��Jݛ>�6���"Ob�i"m�8��s�E�p"O��#S7\� �L!�6I)�"O� 8Y�6�Űh�֌r�%W)4�¶"O�e�"U&������^1;�$��"O�0"�,���x��M� b�P�S$"O&yBU'�/eP�8�˛�M}<5s�"Oti�̐	vs�\�d��/�x��"O�%s�Z?u�&�qedˁ5��Q�"O�b�^�MÏ�X���"Oz�t�LG�@e ��]�(+��2@"O*QK�h�_���;� Ӽ)&�q"OR���7 �]�ab�1dh\�"O@� N��.����M�,8�"On��B�37\���#�<{����"O��
Um]�j���!�����Br"O�h�l���6K�T;�!��"On�K��^ 9��� 4��/���0"OzW��5!3j�	���1#\�3"O&͚ �P=$�%i�mL�Hڭy�"O��0D��- ����	��ȁ"OFĹ���rK�LP@K��f�u "O��xPK�+X�F�T�C10�5�"O ԫ�>lԩA�̎Kv	
�"O��ȁٓ&�j0�b��
#; =��"O�}��%�)���)��O� x�@�"O��%�W�D����$��(�	���'o����� �Q�|8�A�!��U(�B�I$O�B	�B�z���HwFɢlJ�B�ɸd<i �f��C���jQM�1�B�	�D��m�,�p�{�%��?TlB�	�UT���Fe	%+��A��[&�6B�I�RSh�{ׁ�5P���S兜�6Q:B�	1V���gЕ2x"�!Y�j��B�	<)m��%I�6vp<�3d�+Z4�B�ɬ?�j�KC� �ib�15nC�	>Ұh�e#/5�t���>4~LC�	h�NňF�>���K��+�DC�	7L���f H�Kc�HȄ-�;pC�	�	�|�*�6E�|@�a�p�B�1]|h)w�B�*��!
�5BʰB�ɪYg� �7�pm����S����`��<����fur�E�?\ub��ȓ1z�}�Vl
=	# ��!L8h&�-�ȓ`��-�C��	%��L�t�M)5�Q�ȓd ����Y�b�j
02�Y�ȓf��Չ3n��fB����	��e�0��ȓz����)H.* ΍!S�W�i�����رj�#��>���Q5CT�ȓh1"	h�I�b' �&�ڳ%N�U�ȓfn�p!�H�r���(Wb �cL����D{��Œ!�]iD2/-�-����He	BN���Q'�ij���ȓXiN���T/z�ltS�φ�R�~��ȓE~x �K�B<x�� �W>n͸����|�Gׁ9M��j��C�`Lh�ȓO��ŲGL�*p�r�J�b Q�	������'�Ę>$��RB��G`P��� �"�@�%%@ܜ�p�H�~����ȓ58Ƹ��\�1�ƭr�&�Q���&�P�i�ibH�:��G/��I�ȓ���k�(��I�~ȡv��T���ȓB����P2�>����f_�͇ȓZ��J2#N3T4p���ͩ6�D�ȓ��h0�̛2]R*�c[�k�Є��d4�`-�0 {~i�� .1]��$cr����H=c)b��D.�m0܇�S�? *��.�Y�	��`'\�Z���"O���B�:h
,k���@D��"O*��`�\(#��j&o��@��"O&�:c��2qb5� @6�t�"OH�  L���D*GÞ/N$�5��"O
50��ʑt ���, �M��� "O�={��ZCb�Dr�,��H�̕P"O Ii��"a����Y�nDyW"OV<! ��R��樌	�&��"O��c�̀ �4T����0W����"O����`�5 � !lH�)�JQyG�8D� ��3iE���$��[:E9��5D���G��3u}��Pw��3>X.Ma5D�Hc��A�8/��q
֊Xg��4D��[�KM#I4\II�ԫ`#�e�EH0D�`���L:��0#���+G`	:�-D�l�1o޺6s����Ϙ�&�||���)D��A�&�9|�{��C&';DXpR�<D���$�"����R��<d&2T"9D��U�UđbǊ\V�U��$7D� ;s�>V���q��m�g�5D����Ҕs7�x���X+|-���3D��RE��AB�Dsa�	3H�,�W�=D�P�$���ty"���F(N��� D6D��B-�:%��P��ŽkrҴʧ7D�p郇�$@6P�5�4����+7D����j��ִ��ر^��9ӠH"D�``�"��-�r�y�$��H��-�-D�dB�/�3�6�kH*df���C>D�X���5B�p$�!F�~���=D����eɐH�]�B��Rv��<D�Գ�@�e**q bb����Q�b:D�$ ���@���+����y�Z�Z �"D�09"kԢFC�T�wg�'�\�꣮5D��a+�&x�4������[0���M4D�4ca�P�L��,c񁅚S�K2�6D���S-�'�N�����"o��\:Bn!D�$���[v��P6J%{UҰ�S�=D�
��X�E0�sD�]�`�ڶ&D��"e�J�ME�Z�-֏o�b�p��"D���f̌Z��Q�s���T�@��!D��/	?�0Q@s�\<UD�$?D��A	U<��ds�-�aVB���n*D�(��c���t�7��;]6�³c5D�����P ?��E 3��8�hI�K D���D�&R�<�f��?Y)B�[��>D�8�1i�-s�(Q�wǫyw���?D�L�"�շ~|e{���,�
�H��<D��h��0T�x�G A( ��t@�'9D�,���g�V(�f�C�W�>4iC�!D�$��/��hPR���Tn,�`I2D��*��G�-����kug:D�l3�G�O���Q�[�0Z�8�%4D�d0�b��w�9�*Ү��V#3D�l{Ԯ� E5�BC�L�4�S�I%D��1��L=��xRw�۱y�N-[��-D���$%,_�j��G{9TTr �6D���(^�;�Ƞ��ڨo�2�@�c6D��c�_�O��s)�3&���F,3D���dҭJ/PQj51Tu�
4�$D��+�̖M� !�A��'��8�.$D�X�i�<����"G^�:j�\��#0D�8x���^�h�ia*iܤ<��!D�"ҏדo&��! ܕ	�b��wf+D�� h�5�Вjqd���ζP"B*�"Ov,q��@�{�Q�d���>,y� "O��#R��Hl��FJ'$�A�"O�Y8�+Sprxhٳ��V�%V"O��{b�V^�
و�g�Ic8�"O����9Ii�A�FT�%xx���"O�|�̗�#�n}�҅M3)eD@" "Ob�Q�D�4W�0x���]^^���"Of9M2��A��/�n�V6n?D� ��GD�I��B�O$�u�� =D�Ш�W8S����̓'3`��':D�8#E`��d�k�'�W�AQ��+D�P���ߎa/P�S��;�@���6D�t[�̔��Y�F��"Uܱ0��8D������TZ���D�?3��u�q�:D��hC���D���F�K�;�Tc��>D��زDzB�#��G,rN�A��<D����(q�H[�BF�����ń:D���/C�}?��0�B�pD,E.4D�sQ�*V�x}p��߲<m�ab"4D��Z&��$Qmx���/V���%�3D�@)�M�8��=�B�%:�vX���6D�0��)��N$���.�3^�`��b4D����.}�d1@�%�"�k��1D�Tѥ`�:?0�Fj>X�V��3D�<�h\���\k�
A9vk`A��A/D�B!I�a������s	�.L!�dV��"�!'�\afH ;!��C$=f- ��۩ D�6g�}�!��9J�`s� �6R'\Ȣ0÷m�!��;f���`l�\PŪޔ"�!�$�	l*�q�,� "�H��e	J�K�!����� �)*-^�iI�!�Ĕ�5*$���zh�ѓJ��!�C�L(Ӭ-/J��r���H !���hb���w�
�p�����i�!�æI���+5h �2��s�����!�$�4Z�l�)�i�� <#!�T�l`ZB��g2΁��@�!�D]8G�3i�:M~��"��3q�!�+	b���C?eV9��OJ�!�䍑T�kA��a"�����E�!�$��(k�PY."���.9�!����ꕁVh:t�b�֣�8B�!�$A� �h���3#�ģ�%� Vl!�E&/�H�&̤0�<��$�V�RO!�d�7w8��$hJ�A��YB�զ2!򄟋(���!f�IY���p�O62�!�$4RG����G��j�xv�٧[M!���Z�nICF�S Xr�b�5:�!�Ĉ�7c�Jv-ܘ����R!��n�X���:�p�v͡o!��]�T�T�P&K�I��D�o!�$[y͂�����c�V�Kq��R�!���[?����,�~�v
�k�5&�!�d	=B���bƊz�n�#���H�!�DU�LmT��"iU1B�^�)��ͷ) !��$?�ޡӓJFh��G»V�!�DK��]8��э	n�Jc��7!�ձ[Mz}ڷC�(V�h�7�7D!�$πCZ����Q�>R�]Iv�##2!�dQU2 P0j	</A����
"!�9k=�e
A�]�-H�R�.��Y !�DN�,�`Ycmޠ|�M*�#�1T!�� v����?X��+ʘ-v�$"O��ڐ���U�.��#+��:����"O|�
����~���&)�1#�~`�4"Ov-��#��
�*��D��½#�"OҬ�E-
#K�� �T�-�~
�"Ol�ӧ�m@"Q�a$������"O�]@���$��J��T(�D�Z#"O@����T8:h���Н�.�a"OT��WF�6M|���b�$����"O|%���[��0����ݮB�:��q"OP񩖇'c&��G��5t�@9b"OD�!u���)e4��O�PIyw"O$�3��!w�z���*�V䩠"OR�0�Ɲ�tU�=Ф#�dA	5"O\��}Kd�BQ�	:�<��"O�4��D�O\�Õ��.���C"O��cIV�����`B�p�Ҭ� "OT�&��gnT�@̑?�b�"O��Z�@0�F��RV"�bT�<1���#d���n��]�yCǙg�<a�`�r��@�t��s3�M1���e�<����f=x�J'!��-Li#�M�<a��V�p�X�qC"�G�\DIb��E�<)�a��
�p� AL0�XW�<Q��C0 0 �A�u��QeE�S�<A��A�S���`@�ϋ�r��N�<1�M7-�>�y�&C�~gHaj�h�d�<Yl�0=D �W��8�L�@�΋a�<Q'B�i��=�2�+<�r%N�f�<�&��>@mR�#�&]��i� �h�<�a""���EE!<�u�"B�k�<� ��Z8qf�ğJ~,��!�b�<Q����b������@C&�[�<Y���s,.)�#�_�<`̥A��q�<U�I�O{|YR�C'g��U�n�<�%�7�\�B�!¤y�����)Gh�<��fO�W��!���)h
��7��e�<��
3=��s͉�F�ၧ��L�<��o�8
1h�p Ļs[�0S��P�<��d�?Y�|�P������L�<�fCQ��3��9)����f�D�<��kA%T+��c�lۏFr ���~�<�` ;|�iȀ+ր���R�|�<����e9����GQ�:(�pb��u�<��40 ���*X�Q��X�䭇u�<ѥ�� 0H�1�T�6��|a�o�<����n��Qц�UWr@	�˜m�<!���X��
��|0��HR�<� M{)��|	@��ao)#�~B�I�1:�@�N�5���e#A%&�bB�I�?��X@��@�_��C�ɧ|��I���onX�ZE�BE�C䉌2G2 �wNH�,T��N��&4`C�	,G�uk�"c04��BIP�6ÄB��/ R�փr��U�fL?j~\B�	���C։@�d$��Js�,	�"B�I��&4ۂe=Qx���AQ�T��C�	S�4p0V狔]j��)PNLM�C�Is�B|0�(Q,"3�̑Sk d���?��?����$$@F�ϬR�M�D(�
�y��.�j�'A�O3䨨n�6�yrm�U�②�d�/�B��v!��y�6 h�yj5%��R�+&����y2�N"X�f��E)�\��Z�0�y
� ԝ��&��@��f�˳i�8���"O`yaDE�^�p��7�^�j=�t�A�ILyR���X)��g��$�PbC�Ke!��O0o' Y8U�I� � �*g�ǀ~T!�dS	���Њ�<!�8Q��GC!��	�[ލ��ϖ�h�����,'!��#���¬N�\ϲp1'KX�!�dX+dA�xb��Q�y�d��jP�r!��Ӗ8.Xy�ri^�*�"���FAQџ$������|�B6�T�{P����D:pM�P�<i�C� ��I��M���Ź���J�<i# ��W��Dr���B���S3�G�<IP�I�4�:���ƃ�4����ĨJo�<	RF�2�6@+��D�0�;Ьu�<�SJ�6t�����c0�	��@�m�<B�+ .p���ܢI�2��b��l�<���R8���Is�US4jEs��'T��
Ս΍kf���1A8s#`٫U2D��+U�}R.ðj���8k�J0D�|�e��4�j��^�q��Q��/D�p���u�ƨ�p	��YC�]��/D����-j����4�וhx)�4�,D��q�[U4$:��Ŷh�4*D�6��B��k���V�X�b��NL�<a�DRCR�ڲ��9u�x�9 ��D�<�Rg�<�:x9��R�����VE��<94C�x��
'Hҽ+�D���V^��%k1D����h����G�#iI�=�D%D��yg�Q9\�.(@��ً��-)�A"D��� �@)�J ؿ
���*Q�!D� :���{X@��A%���A�	-D�h�j�q�����D��l�8�)D��rV���~����kK�hsׄ�<�+O����#��)�A��&��c$.��q�!�ĉ�FA��㳧��#�0��G�#�!�dѾ>�FaʳxhXl�#��wt!�ڿOzRd�!�(� TsD��
b!�D�>\4a�����A�f�ZsU!�D�o¼�K �C��!�~H!�r{F�!����h�d�ʸk!������rr�ʑԐЄ.l_!�d�[�I� �L�Ftb�ퟋ,�!��Dm@��! ,	�*"Ԡ����W�!��X�ıb�R"	���p/F�E�!�4c`�(�jӬ	��xQ�ěOg!�d��a&�!ye���^b���.�.D�!�D\���[�I�|��bpm�)|D!�䐿f�@�0��)��(�k�|�!�� S�z(���WkUd24EܒQ!���r���(+7�r��Tj�$C!���	A���ED�<��3t�)!�$ľA�\�A��R nJ5Q�Iў,��I,9lK�.�0u�0�TJ�3�B��e��p`0zībkK�,���'�S�OR�e���+phf�R�[�	>4�+#"O�2���*fm�I�G,lPJ�"Ov����{����P B�]`��"O�P�������J0"�&��"O�,��fX	Fl�h��"9�L4k�"O���ʓy��V��-����d�|�)�G�"Q1��"e���Af)@6���?�S�O���S�Ɔ�|���:�c�
)�F��1"O��pa����`���Eu����q"OB]�PC�*L�u��)\#��Q�"O� �!�(=��(S�^��<M9�"O"	��Ɏ�Vk�d�C�Y�)OL�X$�|��'���>����0HI$��d%��{ c�<	w���p��y��H0z��M�c
�4��|��|��D��
´;��+�H�b�m�<2�!��5��d�(�����pOF�s�!�ϱei�D�c�Aw{`4�$�"!�d��� gM�Ye��"��L
�!�$E�������� D��!���'�|����3WW"I�U,�8���Ȳ�4�vC�	*Q#*�˃̒����z��U:���d�C7�"~��bC�����'����k9�܄ȓET�ຄ�,^$��B��Tk�E�ȓw��C
ٿuo0e���%�Vd�ȓ1�0��e�U �Ar*̞W����ȓv�2��W`C�ΜMQ�l��l7:��?����~b�%[9(��j��
�`�`���YB���hO�'
8�9�DA�.q�HU��'o�6�[wl����<E��'�0i
�(��?��=[0B�\�b10�'�Xܳѥ|��GH4M�>���'�yxЯ��n�"�����?�4P��'sDt�Q�ݘ8���C�31�t��
�'�l�@��ؙ@e���@	��W��1���hO?!Cg��b���4`}��5�h�<	c˂�Mhek�ծ=((�BT!�⟐F{��ɚ;;���2
F�M!lUcD��)FB�I�'^fܒ�%E�c����C� t$B�	�?/���m��P;�]�Sn����C� S&��\ %K���C řS�^B��dM�$�Y��a�jX�˚���;?y&%�rh=33��K6t��ey�<y&I
<��qӁo��e���&�Q��`E{��)�h(i9u�P�n���jX�4�|C��-$)E�R�)���� .�.x�C�I=!��q��/͗ Z�M��C�7��x�a�<$��Y�GB���C�I�E���w'�*ފ�CIڔrӲ����O��ɮ;���y7*
����B���0�zC�Ɇp (��Yn8�@�V��.,�T��/�S�O��Ic#I�tډrCL����v"OL����Ӓa��u�4��+H�:�;�"O0�Pr�M2d�,�R�� 8DV*e"O���q��)F=�HDn�$��W�'���"G��$��J?T��w!�?qbHC��<	��z`n�T��`��-�#�nC�&�*���ؐk�h|�Q��1˞��Oj��{�'�v x�@�YI��Aqc�g+�'�f�؄��7Y�dq�	��� ��',5��D��4aES{.�L��'2�0�ԂXH�AP\�o� y�'���+�g#$�\ P�,P`��8��OP� f@D��Y'��r��"OL�:�e�]&V�Q��&x���#�')ў"~����)
0d��L4Z�đ��P��y��H�>��£OB-Pm��9t���y�)+G���c��	<I&��/I��y�A4�z���K�lp@���K֕�yBd�F�ڒ�!e�����%�y
��Nm,���X3gG&!q&B7�y�hC�<~�c��\��BA��y�A�|��ԤV�\� :���yBd@�Xc�|(�B�Lx� q�ė��y��?>X,�`K�G���U�Z(�y�h��
hIрǭG�"\p�I[��y
� h�c�"�.��)���c�J�{%�	\�'8�hCF��v��:��
�`�+V�'�ў"~"��W'7��k��O�y*ѳÜ��y��>.�	��_ o�
�R�H��y��=C��z��e��X���y��ٟV�^l����[ P�1
��y�cܐyҔ `���L4$��)_ �y"i�'.��(�"U�w�|!!M���O,��?a���T�UB�P�������$P����yR-�V}H%Q�ʊV�|�nS(�yb�
�7��iy�D��N�\17`�<�yBHݲ4��5��,G��5	4�Q�yRUd(P9RӤP�:;@�s&��y���?.T�i��o�<1�M��g �y���38�]��#4y��t0�����O���.§4�d����L�s:��d�א8%聇ȓ���� b��MU����&��v�z��*�.�D�Y,��f.��[�TD�ȓi�A@$å��8ۅ5"��1�ȓJ� i1�@@�~S�bƯ'^�����@�ۍ7j�D&^"�6��ȓK%��q��T(Rٺ�@,�,�F{2�'W?��/�3¨H���:@s֙x�N4D� �Ao�5!���4R�Sg��2f�,D���D,��A�������A�%D��j���8Ch��z�$0D�� 2'�h�TԢ�,R�1%���7�8D����δ;g��� #���8U.8D�,��	J�~�z��O��v� �<D�X��ȬTDZjpKLI�J4���:D�p:��Q�]0�PA�--$��ah9D� @�nÅu�bXɞ�3�ꝑ�<D�@��E]�IX�0��m��bd��b	:T�02fF��4��cQ*u��`�W"O0X Џ��"J�:C�
��-C�"OP|ۀ担q�N����J�n��Tc "O~-+�^��p RT�U�]u*�d"O���j��|j0��/8y���"O��À�M�E���FN���F�y�"O:5�W�g~�5���ϙZ��YA�"O��0��5�~��2Iމ;�%��"O�8�` ȡ^^��g�"���2"O��J�gV�oh�:UȂ|�@��"O�C����M�ȍ�1�S�K��l+�"ODi�D�0�"��䝩5�x���"O����>l��*��C�Dn��hF"O`���F"^�A���3GLL���"O&��j�V���[����d�0@"O���%&9^�F䡤oM�[�d��"O�<�hu*,m*g�A�4��"Ob����F1	}�H��Q�&���k"O^��C�����H)f��E�x��F"O��c��#�LxP�NRV����f"ON�@3ژ1�H�$�;z��r"O�%b��3D�M�#/�N�����"O~�)�+8(Ҩ#�.��'���6��Y�ȳ��i��}�����nPS�+�D�O^��� "Y]D��ކ4��3d"l'!�Ĝ�JT��|����#�
e!�	V�T�3�N {^X���aW�%�!�$�0?/hC���z8|� ��
4�!��лz�|�Q�똨%&��z�V�1W!�;c�nd �Fk�8�"\;�!�$%�Ԥ�v�4A��ҁNC������Iz��� ^�J��E#p5f��$��2ȂuYW"O� ���;��a���W,���	g"O0�+�5-�B����MB�X%�"O�z�
S6�hL`�Iʜ�Di"�"O���f26z��5N�%TD��"O
��F��5f��r�,_Op�"O�Y q��+X�5,���	H%	E�m��Q�H�S��I�{a~@� ܋K��� �ϝY@�C䉋A8���СZdJ`�4�K�1/�C�I A������3��١'ʕ�(C�ɹScT(����!p�!ܕX�FB�	��H	��ϙ/�ڹH! �6tB䉺b��2'd��<h�xP��;:$:B�	�L$re��G9�,l�c��	v��C�#Q_����L2Yn4؁@iԉ�jC�I�_�F̱�J�����w(Q"�dC�	�k�&H��FS�	[ȉ��,	��4C�I�Gz҉���Wy����"!(�C�� Ӗ��W�V.|�k��Z�Y1�B�I*����`D� f�6K�%c��B�&3�J��2�ۓ-��@�ǓNFB��o�ٛ!�	9L���d�+Q�C�	����G"A� ���ƍ�Da�C�I/���!"-ҋ[��*��L�Q��C�("*�����	��8à�
�uaxC�I!<Š�R���b�\��cE��pC�IVT�(���hGv��򤈡z�t��>��|���
�jw�u`��]lGƙ e��8�!�� y��y
Q�Z Q8��wc�8H!�dџW��Y���%wN��RGiM+!�Dч�Hy�$���K2.�)�I��!�U/0�3��_�z��Xy��R�!��ؠ|��Ĉ��;�l��%��<�!�dEP�!�E�$A��vH0�џ�IO�O�B4!��Q�N����A�D��'�Ĥd
�Q���Q�:	�
���{�J����`K�+��u�!�d�&<�&���d\>V��ѤjαXD!�J������\�EE~Ux@i�N!��ؘ�����M�f��E�ah
��!�D����f��%7i�Y�ӆ��'aa|�
9¶�ӄ��`B���y"��(̜� A"�����2�ۗ�y�Dޛ"�0�Kd��b�D�B�Y��yn�8�����j��T��\�y�����#�9ic�k�cF��yr��$e�-iv�(u&za,��y®��\��5!�2jʪ���g���'aў�Ov�
� �1-Ju*��ڤG����'�d]�
^��J��S2"A��	�'��ӷ'�
�a`�#t}��'n��Q�M4$H�����	�z���'��=PP��(p��3�k�#�<��'R�l��L?~씋&
ӡd�V��	�'e"ećX@���EW)Y�X�A���?����������K�� 0V
ŀ�K��һ B��m��$�*F�7i@�f�.�C�ɨ+�0l�sD���	H�Ş�k�C�IT� E����8Rj��OپC�3	Y����C��	�̀	dٮC�	{E�m1 "�̨�d�W�B�	�3�ni��� ~�t��A	����E{�O��d��TT�(A��f*��B^	_3�)�'*
&�
���-h�@��Y�\��LX	��� >h�4E�"6���ffI�II"Ox���bE�E����Dȴl��њ"O޴�ƣ�(4�zfe�(��=�"O�I9�Ja�b�"A.��.���"ODW�h|H���Xj�����P�I���OC�� ��aqD�%@_)K����,O �D1��p�'� �c=&�(e���ݴI�$��'�n䢥��WHTh�"l��Cs|L!�'	ɘ3��uVH��ʞ�?���3
�'�nѐ��C+|���e��>hZ� 
�'��ӧ��� -���5�K�2>�h��'(Y�h�jؠ& (�̂��D*�`�I��B;� ���R����'�ў"~r��Ϳ4�v����(Cff$x��yRH�j"��Y�`K:wz<P�Î�?���S5X�|��͓~}fe�Q�Y�^�B���a�8ѸrG�) zN(�D-�J��ȓ&z̅ I��S���(w�U<z1L���F0��Pq��F���S��R7Zj^��Io�IVy���G�(&�p��+[��E2�n�(��C�ɸ9��UK@�ΏU��Y�a��e�B�ɖ
W��dd���	aFA]�wp�B�g�(�rC�ɒA�H�h�ۏ ǸB��5JN��¤�V  m����^#�B�Iie�)*��Nh�TiiA�A4��B�I(#�����!M��y��ԏh�|ʓ��$��)w����MA38$e*a�"�R��A%D� ��S�(���1�dةF" D��kp�Z-_�T̛v#�"�h��ad?�Il����	 Pp��#i�2Eֆ��adV�LvB�I�fH<�g㍊)����a��#�dB�I�M�����K^d�Ԏ��38B�Iuʘ�zv�0*�L�/�:C�I3_zpuHs��wmn�ɉ23�B�ɝGw��rE-�fi���H
��B�	�K�IH3Ɛ��P=.")����?	����S�O ���rAX��Jq�RaNd��'��*@��#�R0/�=X�&�P�'zv@� �R���'E%A�*m �'��	GI��V��9�3���8���)�t�������'�59��x����䓺0>�5��	
��\)s��V��v�<�`G3F𱒇� {����b��y���hO�'��,!̟F@n\��VD�ȓb]�qG(F.8�az�J���LɆȓ��d�3*D�����e�)Br<�ȓ,�Z���)�*�
q����1:�2��?Y���?	��IL�c�
Ա���� �sp�,(V!��4	�!�e�߹&�j�al�  Q!��(W�[ԉ�(z&a`5���Iğ��IS�)ʧl[���%Z$&{p�Q� �N����c�� �S�NUjM���X5:D�ȓʖ)k2Ϙ�EP$iQI��y��1�ȓ8��"�G6�j����(�G{B�O��1��i;I���Ë�f�ՂM>y���?�t���?�b�ձ��Os��H��<J�Ju���Z�B�H
�'�0:4�
>z�mX���.>�^I�'Nv$2�I��ܽ��� "=e>�I�'����8\�Z8�J�9#&��'<�ɣW���kN��# ��>'�zY@�'�&���́	�dç�ėLR�9�'Q�aÐ�@�C����W+�t���S�<dExb�'���xp`ۀm���#Aٚ�y��G�}�(i�6,o��\�@���y
� �0+��L�s�� Q�^�~�|�c"O8Mj�'�i����C�09��i��"OR%��m��T�f�h�m�"V<:02"O�tу�'���C�TY��T�'�'�O^��!?�);���ᢘ?{@f�E��P�<1f��6N���J�	�:Zl3���h�<a�$ό�@�!L�cDݺ��{�<i��X�lRX��	��z�e�\�<Ѱ�{�0ZB�f���u
FX�<�QÕ�=��PL�|�9p��V�<a@�K0�ҴB��Jz�(]` �V���hO�R^&�a5�$�Q�cLn��x�ȓH.���J��U�F8�-�Zo���	_~B됪W�J�R3`ʴY�h(�t�^��yrf� h��[��Y�"��GE��y�'ՠjƔ�Q䜛W�� a�)�y�[�M��9��P\"�fٵ�y2�ΫN��@2��[M6�kl߅�yRn��3U�T�'S�E�ȹ@5%C5�y�N�5gs CI�P�h��DGۆ�yrd�2ڢ�(�ʜBt�X�êT�y�Hٍyr���@ϻ?�Q�")��yB�лz��Q��F�<�t	{�$���y2IK#M�A�#M!6��U�a�X5�yҬ�df�#�
)3��	X��y�Ƃ�v:���ֳ1�$�Q��*�yҢѨR����������B��.�yBL��z�2�A���a��oE��y��L�!>9Ġ�*>�Q����y��έ%��S�I9N�QF虑�y⢅)Gtz9��#�4�ڴ���yR�؀EX���%ɕ@r�����y�!ߓU�ܠ���t���aumM��y��)P��Cr��>���t�P��y��[w�D��46�&�s����䓒hOq�n5��0��)�F�i`���p"O�)��"��\q�n��r��"O��j�b��QrT�Ĉ�"O��1��E��Z踄J�?��p�"O��(��\8"�Ĕ�E�PN���B�"O���a�R�`  	f���_ƶ�QU"O$eB0�F�q��oS�f����&���O
��&�Q]~G�FS�D�F�Z��	 	9#��Q���5aC9A����K���Q*		N���b��o^9�Ɠg3�"Q��6om�c�oT�KҮ0�'���v�K����Β�<5J���'\�ppU# X(�Aē�/�ȹC(O�$/�O,��M�
�z�j�G&EL5�5"OZ�r&�O�����:5t�"O�(9��_5�
]k��?Q�=z�"O��� ܕ0���񁯄4D��iy�"OJ���h�
^$��R��U�:�(��'R�|��اdע �� �4��9sdF>D���&V� ��ȡ�G<<	����I!D��� �_�p�p��--�n�H��,D�l0�
3R�`�ǫ�s�`��4�,D�X!'��7;��A��=U���H�*D���'�ْ�ĵ2Q�Z�	,%��(D�p�!j�$�NE	ŮĴj�V�{u"�<�I>���O��k��i ����ƙ40�tB""O��Z���U��\r#��z���1"O@����L��
Ɓ�AR�3"O�`��C�&!n�� �;H����"O� D�`��W*ty�$��&]��ku"O�4iVhJ�*�z�#��̑VV6��"O�\``E��U8D�B:!Gd��a�'��|"�)q�ƿQY�]����6�x�B�5D�����i�z���D .e�f��$�1D����  �Uӳ�\��N�K��/��B�����c�n�SS���.�}+VD1�C��	f� �@/θ!wzy��Mr�tC�I�A���� �.ٞ���+L;H�~B��xON�x�n�[ll���G,:B�%BĺI���Ww7ZD��K��+А�	H<�'$�k�P�h�b���|k����<AQ����g����#��� �q�`��J֦㟔�	>!sU�'qd����~{�~-���5D����@�� �۔k�`���!D��
���Uy���]�\�2�C��;D� �����]�$X��nێ5޼ᨦ�8D�8:#�X����*""M~ VPS��O���8�O~Xg��O_�	#R��*o&����'!��$.�Р��˹C� ���aéL���r��`b1�+:AL�͏�_ɬԅȓ5�@��h�8���i��z���m��c�9�Lиb�\F��E�ȓf��Tҵkɐ����ǗU�Ṙ�Yq�\Q&���
A�,y�$`�'�a~�n��`M�H�NLي%HS4�y2A�M�89Q��w��52���
���hOq���x�6�
i��	8�����"O �0ǃ�����P̏ ^f��A�"O6��cË29��"�=6=5j!"O2	;���>d'�KP��o?�MZ�"O�<����\�HФ
� Cx�3"O��)�G	$M�V�P$�ۮ%�n�(�"O$� ᄆ-x����f��X���q"O����c�#��41�U�]P$"O�e�� (-��8cJ�1U��c"O�i!b���}�w� w�,�"O ��a�4��	�#(R!Mn��w"O@� �� �Bݨ@�ӌ9 �(�"OZ��d�8=��J�>a"0PB�"Ot�hN
`D x$�_$%��d��"On��r��!4���dH�e�1;�"O6� teπT� ��Ħ��D��"O�̙¢�:����H�'Ά�{�"O�:�@U�+Ɣ��N�&g��1	D"OX`���4+Cv�k0�_��΅�w"O�tk�N�>e�*�Fѽ��c�_� ��g�S�O.-��	�z��Ր@�+���'����:"�ڹP�ˠym2�C�'�,,ɲ&Q�����A3�,("OJ��Qn�6L�P-�ƯӚ$L�)��"O��� V-%v�Ń%�I�FMd��"ON-�S��R#Z�(wMĂC�(�;�"O�=���(���ap,�v��FV�xG{��酴^��H���G���B��~T!��A%-u�y .���0y@`�S!�d�?BZP�) B:z��$��[�!�N!p�؅�� ÄZR�W��1N�!��>mܪD�%N��$Y�)@W�!�݊J��E��)�;o�:�'+֕k�!���K��E�ʹ
�XسhY?c�!��HZ{�Y �p��uS�4u�!�$-/�u�aϙ8���IW���S!�D��*ފ8p ���ꨲri��%�!�� �c�Αg��t�Eg�8%
]0e"O��Y��7ZT3G��2��Z "O
!�*Әg���Ae�U� � �"O�,�"J�iX�	@ �N�B�b�ʰ"O��0d�#F��l�s���fc ��$"O�D�AE؀F�81#Q�\pd�0"O(��"�X��tR"��r��	�""O�5��E	=�ޡ�� ��y�6,"OhQK�%����G�*��A"O(<0���Д�T�I�N�p�{�"O��{�瓥%� Ba�F���"O�H2�ȊdP #�.�=)^�D	�"O�2b`
YL��! ؒW�"Or w�Фw��I�P�Z�l���"O����ѕ?�|�ޒ"�u��"O�a �"A+Qתm�UHT�
�P`yA"Ob{ǚ�-�f�RF M�.� V"O��@��4b�Rb��}�$��"O�0�Zi͆�r�A�=��G"O��4�l����L~q
�"O�qB��f@�:%�=#X*d��"O���pc��2B��Ʌ�V3#U���Q"O� 
�gO#� ��ᐚR8�U�"Ol�Itg�e���J��/l�U�"O�ei�Âg�<�5莝����"O��9׀�`�,��጖�pw�(��"O�,��l�6IY�I{Em��|�c�"O�X�h[�M����l_� ��A�"O�!��9R�\|�6ҹc�j�z&"O�Y;���CrE��
�"�B"O�$�f�5g� 9xK<jp�)p�"O��*&k��a��U@qj�o~�-�p"OĀB%O�.FP����!z�%x�"OP�XP
�O��QE�\֞�S4"O� Iw��:*}pXk�N�+a:H�@"O*)9���Y����`�Q�l��C�"OTM�R�
����v(U0n�x�h
�'������*�LLq�6Nq�
�'?�E��Q�l� `�*Cz8(!�'C�A�
�!	���0�W�@�fi2
�'o\�+GBU#R1 ���`�	�'*`��EʣLf���GF�t��'a.@�똚�R�B��T79��Uz�'���	�/�*%�%��$578`�'�R�
��9 � ��C1R1�' \y�G��0C���*�T�Y	�'�d���%�Cp��Z�F�+´l��'3<����D)W����V6X��qx�'Vt���b�$2|S�#ҞI.�h�'�pᠴ�ʌ���[whG�P�e��'clh��`	�I�q��?W�z���'�Ԭ�&怫t�@0�ը�?z����'�
�a�S&�5�HO�k�\���' ���7H��uޤ �,�h�(���'����.�Fȱ:�� *h�=��',xA;�ϥ}�j���SR&	�yIS,�HrQ@j�};�k
<�yr�Ċ�d�+h��f��HX��ȅ�y�a�6�2�j����h���tGܼ�yF�N�J��W��]�� ��NZ��y"e��A��툱c���i%�Ü�y29�ر��`^Wx�sSeٛ�y�N�h�f���AI&#����R�S?�yX�;�s��L
���
r�*�y
� �h)c�W�"
�y��Pn$�e�!"OpĢ�B�nc� Wcm ��&"O捩F$K�`��P�mO�0R,�Z�"O�!���V�V�:u��_��x�"O��	�&g8Hx�3.�	e|2� "O���c�<��1�l�-n�F"OVB�a 0&���1Vl�r���"O�/��[��s���df����!D�Ԁ�M.7W0�qbD��oj� �=D���G�.SXY�1A�O�����!=D�p���>_�(��u���w։���/D��K L��2)��-P�D,D��0u`_(#^a�a�KV���rr'D�ܻf�N�`R�QC@�ǒA��y�&D�r'ew֥[�ؑIp�sB�$D� �IYjoJi�����V�@�g>D�l����v�$dQ��B��
�7D���Ҏ��g��ٹ�L�*�@��ŋ D�(�@j�8�1��B)hTF���<D��H�d��d mJ���-#̥B�:D�D[�F,M�L��N^���	�:D��J�W?H.*���o�SY�6�4D� �t�	 mq1C\�)u�4D��c!ξa͆Dy�@ 0�A9Ѡ'D��c�o�x�2���
Q��$�g�:D��p��]l��j֫S"r �H�6D�p����F�X�	c��O[*��4�2D�,Pa���<`�g.�0��|��%D�(��tFΌ�꘬b�T��-D�h�%�ۺV�ɐ�B�Ls�|��	.D�H�n�-|��+%�Q�'f��2P')D��
pȀB���ۓK
 *�����%D�0� ��5yl���e	�8B�a�!D�Ț0+��XP��
v/�(a6~\s�N>D�$Y�O�*Z*��bt$1M�����<D�4�\�#*!⒩���z�"M D� S��t�:���/aO,���3D��u��<�{�,�5
�m�C1D�HY�'�, ���+�̍�.C,�.;D��	G�b�r�bŊ]�
�@�7D�Ġ���L��=�0`ɔ�YZ�!D�@�U��>A>%��-_� =��<D�P�f$P:Z&Jȹv��Z(�Pd�<D� �b�<4�I� �	����g�/D�|���d{HA9��0��0"�I1T��If��yn����ˇ�k7!�4"OhEBs�6F��㇊�-Mh���"O�0i�#�9+/İJ���	Y9*X��"O"��-~��ڢ�߳Z4��w"O�!8W�E!�zq����7�x�%"O�YG#�1wh�2S��1� �"O����
2"������"!Ҁ"O<< qKZ�JT"wV;E�Đc�"O0LhO*6H��2���;\d[�"O�� l�4T��b�CBSG���"O$=��d�YgX�cĉN����yb�>M����sfD��<Yچc� �y��k��}C�A�y�80ƧC��y�ܓg��sՌ�-��0�բ��yr+	���LS�rh�%���y�F�Kl~���膗k
$���ᚶ�yr+T�3��웄�NZ.�Ce!ߍ�y��1!`D0�� \�6��TrQh���y��7f(8�k�� �X��f�]!�y
� 4u��%D�^�$���IY7���"OhYrh�%M�&9��̎���"O"q)Îԁpl3Qf$��k6"Op����/b�0|���&"� 1"O�d`�f��o�*�H6Mܫ9� ""O�9�"b�-z�Ġ-Ʊopv09"Op��.�;a�<����54T�y��"On�s��
}�N�a�ٟG�e0�"O�T�D�،OV`BQ&Øb=����"O�H6�ѣ�M�7eL3}04"O�\9��62kg�Cev�[q"Ob�&#&:��!e�<Z{^��S"O��`�i� �6Ku��k��B#"OfD��E3!$��d!ւa�.t�S"O*K.��;L\`@�C߆�y"O��3caF�gqR<xP@�r����q"OMxT�5_,�M)`	о{�"1�g"O�5� �"N.d`�F�W昐;�"O4�@��~���s�%��9"O��HE�-`!���	k�>�3�'�Pl�p$��:���ч<u�l{�'$�жcR�\ AKW�dI�	�'u�İa���V�H�p�j�}f�*	�'��4KlXazu�ǅj٠|��'䲌`𥗥  �뤈��dq���
�'�ʰ�4��+	 r��dH�c�@@	�'d��sf�| ������_6����'�	��`ۆF�`@��Q%�z���'�Y��b�-,��@fE�4#Α��'ښ	��Ā$����G�&�y��'|��QjH Kz�ɷdB)S�e��'�>��V*HA�������0�=j�'Ҳ"���.(zK7@������'V6ra���豙����U
L��'tv+���}�HE���R�	q����'%�2E@ѧeW�tF�{[^aP	�'�u0���7�U��O�8s��t��'��a���g��avi7q���'�p����4@���z`*	�'�=W% �5��2ix(��!D�: b8p�i��!���a;D���Ƌ_����bI$���)9D�0�C�ߍ#�ڬIe G6d>��[e8D���R�.���G��D�5���5D���NxI�#�,!
�@aa@?D� s��R8T��@�RE(qi�i�C?D��8Q*A"#YhaI��";uxhɷ�)D��Y7���8b�Q3�m�\@>���&D�tKU�!")H�pB���4�g�"D��sv�M�1����5�@�`�٨��5D�ȓvĜ���b��K�l̾)C��2D��s�I�{
^ �,��Z=V�ra�/D��B M�j�zl!��@��hP�2D�������4�F�O��h��*2�O<}�O��S����K���gj��~��̋A�2D�|�5lF�K%���?g F�2D����G�d�8�'቙H� E��O>D�T��'�+u�aX��=@�(Z�#>D��	'kN�e�� �&E�j�d?D�l�Ƣ&\�
���G�Q�XX*��9D�p�̏�/�$Hjbf"k\��M7D�pҕM�.��@#b#���j�0��*D���Bg׷sfN`�p�P�te.��T�(D���Vh�1g���mK�a|ހ�si%D�� `��#Źd�� 	���rM$S�3O����]�Ԍ�ĂW�#�蹱#dS�n>!�$�2�ji����;$�ݳDҡ�v����X�r���efF��@�o,��hO���+���ڂe�m�a8���y�x">��I@�<SܙB@�%����n 1!�ǘRG��r��۽Q�����)!�dЎ
dȜ�whU:Ǻ)����F��O����5b�B���w�ΰ�f�2��7�O��#�)O1�*�R�����}�"O�X
cj��o4���eȯV��	��'��D�t�>Q�4��z����I�tn��*��DRn��yrI�o��q�+�@^�鲤)L	�0=y���W:5fHhAgKٶj�bĬԮ�(Oi�� ڹ�voW���p��hV�vn�%��E{��T!�
B�$z�߄���KU��y�`�!��Ѻ%��ީ9����'?az����T�؉�W!6�^���'J��p>i�>q1B�5��Pj\��i RƎßLΓ�~r�'b?��O�N4+�
�>��f%Yۦq;��ɧ#ĢZ�#��!U�	%��W��{��n�<��!CI�$�����&dS�ٕX!��Ey��)�OvXrf�ɞvW4���E��9��Q2U�@��	p�p1�W��;r���y���Ysh�	�a~2	�G�t1��p�a������>���<��d�Hx��Q.��YGXix��	D}��'�icfg�N�[�,�R�1�'A¸# ��6�p,Yf�J!H���'��M3�ǵ5�d���H�@-v�.ON�=Ys�Ę�.�@w�7��]�QmR73��	a���;��DC��	���/��q�%�7�r�L+5�O�`崽��)!����(6D��y��;=�HHS�+ {b���#�uӈ��m̓e�Q?!���ȍ"L|�ad̚Ίɑ`O>D�(2S&7� sSO?dXEԥ<D�ܸT皣J�fM��K�4%8�$:D�h��Ȇ�n�P�[��	n���o7D�pRb`�Tl��@#�C؅Af5D�,�pFۿ-Z���hHH̚%C5�1D���a�
�/�R �¢�(4d=��;D��pb�W�%���|rdX4�%D�h8��$��
��Q��H�T�#D� Y �"3,�i)�`�' �@g�5�O�II�F��T!r֪}	1��+?"�B��HM&E��Z�[,@�F��0��B��)�L�K"K�*�@� 蕭-E���$�/U���<ad*J!h,�"q(�{��}�؞D!�Q�`jqJ�G�e��I� ƀq'!�P�/R� ��i	*�d��c�!�D��7�VL����a�B��S�HD���D��,T#Ԧm`G�H�\�����!10!����B��E26.���P����9+!�#0�@ԲLG\8��C�ߗp!�$׳xsT��Ś� u\h��b��P!�$��x����C�)6���8���)�OpHP�{�����&�Qwo�1IGh�!BL�:ǒC�Ʉ2X�ar�B�&V<���g�mfC�Iڟ���G�F6er�AE�Z(��
��2D���1�]�/�
[d�C�X��;f`%D��ȡlB+'@�5b��η��d"��"D�4��ߋT%�T�G?V�N�6͟jy��)�'I?���!ʗ�8��T�����K�jчȓ'�
pH7�� ,��@���Z~��� D1A2�]�%<z`#���BD��'2��z�S�π ��[��a��䭟7M�R�"�i���o8�Djs�Ϧsf��Y�'6h1�2�(}�)�ӫU`P�A 2^p���һߖC�	%m.t�f�\��z�#�Q5#%���&������?8|���Av���(lO�Lyb�'oX�%K����!Y0����	�'4Xt	�B������2fp{�'L"�I�`l8��,B>UX�bO&�y2/�W�B�*��F�Ѭ��1c���=��y�X?x�`L��BK&I���!��N��y�L�{
C�	J�"�qAk܌���;��&�'a���0�ǉv���`��Q�;�L�ȓQ���!��6h�L؄�Ѽw��<Fz�g2O^���'�#[��8ũ̻b �%J�በD��Ix����Hȕ@g��P��A9E�p��"O P�G�B�enp`��^0X�QA��'f1O�PL��6�Xc��W$V�bհR"O���Q�D�a�����F����W��;��)�'M��2�C���([�"�M�rl�ēR�J�P���
� a��Y�"�8��>I�`+�OH�wj��p���C�ɋB0H��"Ov�eH���R�P��V����xb�'B�0rA�I�{g�"&48��x{�'�h$�7�
��>U�� �(��p)�'�LEӕ���8LXǈL�I"ы}��)񩇘N����kFƄ�ZAMA�2�!�d�;w��5`#"��`�0E���["=�!�$�O���Eɐ�̚Ē�K�ay��'[qO8��4��%W�A��툐A��ȥ"O��a�FгA�9�r�P-N^��"O��� �ϟ2�����q�.���"O�����,� ���3>B�0:���3�(O�c>�j�&�
�� ��%X8H�����$?�S�S�k�u�s�W@� ��b�tB�	n���bR0Ն�q�C�;�^��d�<a��+W4Aq�JE"(��+�W|!�E:6)r�҇a�'o�PH�-�/o!�c ��x���;��S�?$o��XF�d�K:SR�ܘm��4 P���D/�S�Of�!@֏�y��0�S	�2#�TT	�'�hI1*�7k��p�+p�h�'G`�A�#�3Z1�8��%?����B�)��<�hT9�, "t���Z��&F����'�a}�J4x�4ȗ(��~8
YzBJ�y�� &~�XƦ�eGɹt� :��?A�'����G�Q�m1&�_a��
��'�>E0�iq]��c'#�2;[�����5���2��3�޾4$p
	�T�(Їȓt�<Q�G%O��!1@� �d�dH�ȓ4O,|&��6q�z̐��&*M�)��x�.���.�� 2̤���l�D�������9��m�2J�ݚl��{���*'��L���bko�D�ȓA莌H�郭iR6H*w�g���ȓn��4[�L��,.�`Z���[R���ȓC��@[��ˣU�|˕�A
xt���'4���AC�h�8DB��d��B��a�r'�8lET�qҭ�i��Y��
L�)�B�Y=!A���[T���W���؁Ŏ�D�ũ�FA�u���ȓ]�*�䚔Jæ$z���c�V]�ȓ}c��G���Ň�7)���"O�U�G�(I��!�\x����ʡ�y���*$�����)�g,Ξ�y
� ^l���TPґ�jL�+L���@"O��� D�<:N�TKR��j,ne)�"Oz����5�̨��T�(�T��"O���`�Qܰ�Yu��n�ف&"O2ܺ�O���
V��?R+x3f"Oh�k5σ�:H�|���˖u�v�9G"O�-�f#��5������K��� �"O��ң�k��2�"�f��EJ�"O����G�\�&�BV�N��j�@�"O�a� % ���E�3m��3֔p�"O���Uj4sy�L�k��'��"OJ=� Z���ēd���3j`���"Olt��%�@�iႦʂ h��2""O�P����8 vdR��R�n3h !*O������p#�רc6x�"�':�!��Z%o�VT ��<
�:���'����&�&I��� 3��i��'����B	�{�y���ܒ^~���'۰a0VKD�j�
 ����L���q�'���ZTk7$5|4@Ņ�6TR0��'����$G]��9�U�^�'�>4�'X���cf�\�2Tݞ	����'oL��K]#�D��&C���)�&�2��	j��U<k=9�$�Ш@��=�d��h �92͆ȓUD��F(J1=��u�f��E?�؆�2��|pCV�J��0J�^�V�r��,���杸>ݪŉUD�8XNv��ȓ\���6�ǄBN ��m��r|��ȓe�TY��~Pec�*DZXx��tq� Y1�T�W��b�*�0���\�x�҄O�
z?��z�̉�X6� �ȓ<Xข1��0��7C!.�椆�k�(�I�BF(m	����5���ȓo�T`Icm C7�0��]�5�>d��2d�H���!��`a�JM�M�"���H1�̀���#��I��ވL�d�ȓZ�s(�U�Y���" �P���;%�� 2�U�|0�a����񢕄ȓo��% ֨M��� ��bZ�a���ȓJ[L ��(�$q�(Y3�^�*��m�ȓ0�x�J֣�a����t�>`����Z�>�;b��6�N�bd���p ��ȓYU>)��U�04;T�ҲQQ���9,����|B��.\v:W#\O��e ��\���
��T
�o �db�,�)T=��ȓ�Ni� )�,YP����?^�'�����׎>X��1��f�O�(͈B�v���A���z�0���'LԥA!�Io�t{Q@�1O�6А���v�с��O�q��!�u�g�	�?TU�I�Yf�l� z�B�������\�`7+J	v���`�/c�$��Et�����r�p5�T��:���F��U9b�?��h�9,��h+P�O5nX����|�)�g�2d�<�J��2?��pF�0D��� A�+(*�1����	����f��DYq�Q��&l�w��7z�l�pE���(��4J�h�Q ��ހ@Uzd�u"O&e:��I�&A!qL �%o �"���$u�� ��Q�4r�Q)W�&a2ׯ�&I9�{�C�3�����9(�(��'�0��<����)�$��G�1=�${��@'n,q�h!RhZ|��U�X�"Q�y�"0��Eg��Lj"왑A�3C�T��.�3�*<�@)Q=�I�7*U9HN�)�#�6dl�rE����9KN�=kA�k������J�z܊��Yy�'���&Ko�O8�ч���vu�CM��B���)�a�,��Pk;�MY�n^�g,����J���!r��ϻ"Z䘉��\�HM�F�I�;�%NYʽᐞ>!����u'f#]��V�,^���ŉ.�bB���1K!f=�ℍ
W�䰢��"U�9�t����'��\�� �*���ř0 N�d��4Z����5�0N�(8��.Gb D1�I? ,B��
�S�(�C�5�F�Aʓj�0X%�Q�g3`��<��Oƈ*E�ĨL]�=
� �ǀ ��ys̏5Xu��+5�[c������P)��5��Q`-^�2h����ϖu�PT�����)[wR&<�%K:®����E%K���[%BP�ʓ�$�f/���]�!�t�_��B�'�԰��N� .�T<ZF�V2')�0¨�o�5��jĠdp+�&���S/�����D�߹X1���d#��.,�@J��5��õ#�<L0��I�U�tM�'n9Y2���D�Yy��9~�����wN��X���-#, �Z�o�U��L1wDڎ!3\�Z"��/`�xE(MsE��0bc�/''��'�޴x�g�;x���R�$E<`\��4r���ǭ�%MtTJ�S�����?5� ��iP�Q��33����;D班UQ\�2Ǭ�^����Gr��J��q���еX����s�4X����]Opz�:�lI�}{�t;a�f�����-VԐ	�ƭ<y�f]�2��L�6g�h_�c�����Y,SҘ�O��<5#�i��k�GW�/O����΁T;\ ��a�'yv�D���Xݴ�>��JK��ͼ� �մ㨰����?��8Ѣ�I�	}He�A.��)�S�M�*ւ�� ���矙$R���A�*kǒPاE�Hh����M[��R���l�~]^`��FJ�Kٲ�K���
��t�EĔMa����]��ល7l8	��&ݕHD�ܙ�̂ �#�#(g�}�N:�<� ���3f.=�"��OK���Ӭ�"�3&R�>Y�`AM�
|Ҝ��b޹Rxc�#�����`̻*���'_:` ���5�~�����T�0 �RA��{�'�*GԌQ7 ��dE9Vx�����sj}�ǠA�RC��#gY	/MĨ�@֖{ t ���&�r&O�"�&)�6H�m��	�@�Q�m�	ݒ��C�%P���X��$�˧s��T{��T3���(�l�0b��@��1sZ�qc�މ��%6k�w��HK����|:��_1f�����aB�B�P8�����) �(��0i]�'.8�ß�"���:�H"�S�}�Fi4AFH��9"�ě#1֐0���уI�`%��B��bN�-B��H����1]#�zFdڠ7ۆ�7�x��t?D��Ò�p���I�z2��i���:=$U*���B����M+`�N�|Q�R+2�v�sF+p��RA��FD������!Q�P��GY.�(d;Ԅ�*Y�8b�`+��X�X�>��'}��W�;rEP�C$L�'161
m�	x����:E�,lj�C��uڬ�����tHF��� <,R�mJ�z�� �;4Lqa'�ǝO8���I�EܓI�����"��<z2��g�>C�@�<�&)F � !�@����s/�a�:B͇�J�l@!>�*i�0��Y���ہ%Ev 
��P��̩��'r���7ǎl@t�B�"͡5E�e�#��6GJ�)����/�4�D�>o�D3Ԥ0oGz�P��"3N���8�P�h��p�C��<y���F�2�B ]��
�;L,��G�]h�6�P��46�4��6g$N����>V��`[jR)i�h�t��K�������mv���DA�sV2L�2A��D�O�my�eB�(� � ��h{���A�p^ d��-@����FD"�U��J��tF�����Y�BB�	�vT ��ω3�|� �q$��G�+������9� ��M;�D4l��A5"�l�;XȬ�P�I��e��4!e��?�i���
qܺ��mG�;L�a勇Wo�����g��Z�#D [�D 5�/��AHo"0X(�K�Sf���J<i'+/"�Ic�H�}u�(�����'�b���d�o�Y""Ofd=�.׊Z� ���@ՙv̡Aaˌ�d�.��Ы*N��@���p`��2,O�3��u!��˦"�����Oa���U�GȬD��	W��8֭O��@�T�
�(��� E�g�����XT�(�܇R����R
�*�E}�e�c|�u8����^�(���Z�,i��_���+E"շ,$����4��=*1. 8V(RE��B��3�^#��%"��'<��XJk�����#4.��S`�"�t�|Cv��6�E|	꼻�˻".*��'D��~>��`˺'%:ĺ�&RVÆ�㡌��8�x�dm��j$�!��	>�(��!�%KѦ�� &��Tƈȳ,�.�ēp�ݻ'N�V��,��S6�!�-�<y�2�JU
��>�4	A���p�͋WN+R�� �㋓�0�%i'͑�$�����R�V�f��c�˓�KMZsf���鞩O����E�
�(O����/ǑYth0�2�
�3h�c���M+X{%P�/�����1&nԍۤ �4P1��H5f��'���h@�@T��s�FFQ@d�5��%6�ƐB��N�'�����GBYPD����'2�֌r���>�4�� ��y0p���6�8���'R�] 8\�w�Bk�m;a���Hp4��Š�z>d�K���2���G�+\����H»w:����LM�:��ӂ�i8YP�Nv��y��tP䰫��Іr�` q7��q�(���8|=A�T���S�9+��1��A�Ms(tHq@X�5�b���2*�L�dG� ��{co�x�I�"�꽋��X�=V�0K���G��q��_9��	�#��UZ��	d�M�&�����)ز?_�5��@�����.{����j�"vQ�U���r����Z�����\�J"=)g�΋T��a�So���t #��R���;���F���	ǳT�P*\�Ul(�@�Ę�r0oZ��F����A�DL�(SC��t ��Y��O �9"B5'`4#=��;Y��1$�
 ��(s�!4��{�U1 �x�rl	?+{,��F�X��B=C2L�( ����炩i
�}kphT3%�p�2�,�=-p8��& �6��$̏�.�Fm1·�3}�1q�3:y��%�)n*��x��� C81��NUС���]4o�8[bd�<)W��Pg��Ӵ)�3'ln8�N�_��x�L�!3b��E���OЈO��Zv�MK����k�����ʨc,� i�ߝ_3�A���>"���"�b̐O�����Xm���[��
)c(���gl�f�f�PF�W�L>8!���y�X�y��'�lX2���GLW�&6&x���*������PpjaybCB.v|��iʛg5�qg� 4&|m�yX<EIc��O���r���5�D��zŉ�ӅO�D0@��DQ�7�J����[..�D�3�F�
K�q���pc���+
�'�|�t �HT\ȡ�8��l��bL�O�$����dكkK�!�p�OI��zp���v	h��٬>�d3�'f����Wی����L5v��Z F��zH��-=�Lc�.�.b8�q��1?i�M��+݋|�Zl[Q�S�F*�&ܥm���ꄴ�0�y��ɗ���"����H�3�ӈ*��MI ɚ)�����$:54��,ߕ���B�
���\�c�
-��a����.��Y�I����� �'|/�i�@* ?�a{��Ż,@]�tC�I�&���dU�Y�0�� ��M>�}�4�ӹ[IX��eHS�p<���c�N��fK)�SdZ��� ���gD'37�Д�	�h:H�������X��}$b� h ��A����+�AA�,���c�F�5�|�2 �ő0wϺ�6HK�;2���7�C_{��k>�ئ� ����� �n��<��$�\@�R�Q� ���O�^�I�'��d�:.�
4v�X9�!3��Yq*D�a�ҭXS'L�cdm(��X��F,FN�?])��J�HeP=�� �	d��"��
6����D�>�c%f��L���Q�P邙#|�f�ŚIU�P
#Os=�IZ<xL�q���
���ć
�2��ѫ�
�zRn��Y���V(��	�l��t)!a�kJ	��E�� {�t�΍�Aˆ���R"+�'I�o��h��Ӧ(����N�<:�h�qNK���x�i
0�U��ޓe�ް �ߌKX8��I6p?�	!֭�����d�ýX˄H��^g�ʜh�I�NP6��5L�6r�"�
�*��f��*��1N�Q��Xpb�e�)K�	�� N��8r]%��ik��!\���!N�Bq��j�5 ? )�EGɲ*=�d(U��yC���#Yu�'�V���B�8K9�l
e�S�/����H�X�T
@�Wb5K'�]qx@�B�)ƔN�
t��%�uҁ���1ᤘh6�6B��Trs�A4C��"�.�c��Ms�
̤5D����&_�Lpf��%4��E@اG�t1RE�Bj�5�㏫^�QT�A�#R�x(�f�� ?�� ��F�@I�e3k�:U�Q���b�vɻD�3�E�'�M����P4�}�tƍC�lܫrnѫR�Dk��7Jb��0���=)����%6P0�Y����F�z���NЩ�E��*!� �3���!jĹ�bő�p�
̇�	�=1 � �n\�-�~��� _�Gԉ�A
� OnA�� YxT���Z�-rD�i��ٱ�F�O3����ꑡJ`a�v�^�	YiT�ʒbB 4�	jw���.��k (Stn[�P�eÀ+�UTLxh ���C���@E�7�ƌ:0A4^�Q�G�o3�Qwg��!!C�ܗ{��U�V�߅��<a@%\;s���Ϊd������ Y؁k� ͌_b�����	8H6�"�E�u���uFO�`�����R�Qʽt�C�*�(����[�Z�88�r�ϯ��?DÈ#w>���gMYB���)�-c�TIR�B}֬�e���:�"�M�#v:�0�\K��HQ�/f�DQz⧂7 &	K�LY�v�X�`mݨ/����	�g�8�{Tb�1m�RYIDl���Mx3��qutY	�*�ZDZM��z�$g�D�*����H4�i8C&�spzyY�"�9~"iA� S�&\���a�R�G��'O�Py�ߧF��sW�%) 
@jW�
�p1�Ej$�	9u)�`� ��I��� D�� ����/�1("U�t�Y�Bqb�2l=\O�{���+^D�	��!f�\��^;4M̉���#��="j"q��3D /TR�aB��#c�^2����c�Թ&^@!���R&.5�!��~�'���!U��W�O��yKc&�&���"vf�[��
�(�52k�1qB�	�eg]��,�!P�zas���$����f�_��,ReHW�6c��)��Q�-M����[K�@R�dIR�y��$j�ҧ��P$j����$�%Q@��yu��+n@ʈs�.[,`p�H@J
�N����V��s���`�W���\VHEk�&9�(O�5k���9O�: piJ�B^`m�:OΕ�D� �� 9�e&?��;Fb��K�($p�I�GTrq�S�ݲb&����08DH��x����X����V���G��L�q�7�C�����g�-R��U3p�� Wٺ�A�)ΟG�P��$�@�?J�
�"���)��KyܫáA�Uܴ�"��A�D��t��?>r��6fg��l"<Zne��( ��'T��Ki��83AX`�dg�����BFnI�t�j�$�al���P�պb�μ��.ǩuK��b&�����;`�ޔ�dΆ�sA��λ 6���FR=�¥!����c�e*0C�j0��g��Z6�o�����?�@�"߳:�,1�aG^N��ts�CS11���07�ܐVF�DJ4r2"-cCkȎp[�!�dK��XW�34���$����L��P��d$	�#���!��8|�T e`݃NJ�pRA��F��wL�V��$��!���d9~�@m24	�3���i�tXL�rf�N�Fφ�rY`��i�;.�|�P�� �W��mۣ��1"mz�s�Q8l�=W����0BUҠI���E������9ch03t���u
�mH�,N9]�%�&G�B&Q3��̘��8
�bY�4��UzCB0�� 5��u*��Ѷu�ܬa��
#1-�ps�$5 Y;��wm:A3Q��'= *�/7$z8�)w��6F�}ړa���\t[�grd.U;$�%9<����yw ��{/<EU��f�(�����(�H�Gb�VaR��=.t��� �$x)4I�O��a�F o8ɛܒ��P��B'){h���f�?N���IQ�ը�?��&�Hb<ͻ�n��D����P�yo�'�H�14MP�uO�9��nW�}V�4B&�ŜG�qS'䚱N�d��7�	�g�@�4-4sF���NW�z[�<Jh��G��%g$�_����
6v6X�uʝvJ����K	=0�|KW�!�		<4�`�� 'Y��H�fՔB��r�  �0�2�
F�_kPY��\.sdSC���g*��զ�@��z����2�*�J��ÌZa@E1t��7Nd�8ӵA޷g�N�����I��D@��A%��Qb��/�!;Պ�c�`b0oۧX�F5�ȲP^l��I%�p�����m�� Sq�$E2�|RM�8\�P��PB����"�O(,����9�R�\9O������'%P,t��k3+!��=}�uJR%B%��Ò�]�L��'>�ϻLr�q��Z_�^&>&�H�)�=�.� Ȓ/-�4}�"ދq�Fd�S���>����S��ēM���M�H�L �W�N�,9q��a��y ���ʄ�yq�lۢ���|���M-J�F0�7�N6-;e� ��61N�Y���1M�Xl�օ��b0^1(�ㅚ�T=����4o[�D;��D��i�f�z`fG�5�6Hj�C
Hl�X���|��q)gå2v��q d��gZ�(��Ä'3_�3qkO�PǶ�ǁR�L����3��4R�;�Z�h��pÌ��[�_����46Z���۹m��P��K�x�؁oD�����L ?��X*�<�W�71��b")�z���/k�O>��J*�h���I>M��y�{�D����{p)Q,XE�ԧ�1^�D�ڣj�ZN�[1g��j~.�%*�+<��eo��y)� �f��|b�սy����E�Z�93�)�Vţ���X�^h��'�AE��O�0�O�6+�b8ʵ�W-X�,�b�B�`h�B�]�|ц� 憊'I(��'F�k�:7�И��D�t�>������J
!'a^�`����]!��=�`IF?*��s�~�  c`�\̈��e�"u����T"O�  �X�dG%PѤ�@�oK�fq�PkD�I5F&�P���(:JU� �*m��� ��ˉl�.B�ɚ*v�0l��&�u��KU��tB䉈?ph�p����Y~N}����7'�`B��.524����+&��+�*�	!
�C�əI#n�"CE�$���P�L�C�	�,/� �,�2*�,r�l��:<FB�I.��Ũ�M��Q�����K�yBB�I�M$Ԥ�G��26�Q3�ˈx �B�	x ٣M� ���U��L'*B�,��h�l�
�0A��H>Y�B��%#ê�YG���Kn�K"S
�C�.l�ؓ�A�ђ<r׫�7[�C��2��)��!r@�[1��n �C�I��2 ��Kn쐒�'łB�	��y��LW�:�L�D�ȟ-7�C�	�Cr�!bw�l�$hb�H� mSbC�I5/����	g)�hH#�$�.B��8<�(�,��:Z��i���q�B䉌j�n�3�Z�n"�1��P\��C�?��ĹU�Q�g�h�� �Ca�C��X���ª��c�^I��L��C�	�ḫ�PN̂	uDBQ�Q�"�C�<
��y���*2��3/�B�	o*%��eͿv��xak�/qRC�	�d�PHy�M���#+��B�	�p�!�B�W��KeG�<��C䉽����!"�;Zz<��̂�i�tC䉻	Q�1�7M	((} �5A�2xۼC���ЗCP�n�:��r� 'b�B䉜"��a��*@Etbu��c�xB䉧!Fu���	*![��ѱ��>�DB�I�:���0"��a1��I®�!
.B�	"n(x��Y+��#D��zd�B�	8���r�ߢ�|�x$üe�C䉜`q�̀�a9�.��4%�2BC�I�7����"A"NJ�[7�
&(�B�	�iG4y�t�0,�^�Ҩ�,��B�I4V�=�Q�
�ewʀQjĥ_�TC�ɲ*��cT
��K��b�C�� �B�l7~+&@��xln�[֯ndB�I7qF�,ɳڌ
��"g��K�C�I�<j��d��<Hį-5l�C�ɺ`Z�K�G���5���	 '
�C䉣a���	�n���#�mNB�I�sA(�vΙ!;G��5@V*^��C�ɦV���XC�Ҕf�N5ӆ"�(ƸC�I dXz ,_ �\=���F&Jΰ��$C(Vͺx����>Aa�[̸豒 	$#j��1IUO�<YDH�(� �A�G�#��)���8�O)��/A�C| 2�a4��Е�bG�L�@���������ȓ 4.�A�L�!G�rm�R��r���#C��6�z�'�ܙ�4�>�3��H�X�c`�B(AN�]�vm�<���d�$z�,P0�cL&J�x ᨏ�[D����l��P>�x�DO��������?��H,�?z���jCnD�x�B	�7a�l���ǩ	&�yſi#̘Bģ�)@DWG%}�T$��'��\�W����ř�A��"�p�Or��cc��sO�%���h�ˏ�i�	O������� L48��c�K!�d�V�LE"r+>#b1����w%.) ɕ�&���0֣k�,i �bS V�HM*b;�1O����c��E�B]��ˆ�xxF�'�FU��F6zl�^tXs!P����Q� ÞDyFn��0Q��]^5�'�t1�%.�2C����e���RE�L<Y���j"f��)�&��Is�US�2��Bרl���r��P�!�@���e�	��RR�X]�Q�p�e��3!�?�
j�I��xs�ՆWd��aM�,S�|@�$
	�12TM ��]3�p�Z��GĦ�'Wf���f�� \�S)Ct4�[��r���k��Ŏ:�4Ygc�p�$#���]�7W"\iSk�8bx�5"�fU�m\X(���7�V�;��أBk\m���D�4P2|)�kT9a|��c1i� v��-�Jmqp��Ea�$��S3�JY��.}H'd	���GZXyv�QP̅%>/�D��ؘ{��<�&�&-�L��&m�����h�n��m�>�ț�s���ZP	.���0Q��U`��Uh�:^��u8�l0?9#P��ܺ�)���0��c�Ѱq�R�� �١$����e^L4��H&�@�:��C�w��K��Sy��:w�U;0oXId ����w��-ʂ\�z~���n��l��u����)P�������M���FJ_I��=Ң%�~ZힷQ��T��^= ��A8a��92fe1y��uCQ�U��3v�X��?�7@�_?�%Ɂ�`��=2.Oz�0���)"�Q��A��{�	!�� *{t�j�X�F���g���x���G+$��e�Q!D�{y��+ )||�D��v~�r�҈][� j��f7FB7��)R�2��%%�!T��˓Z�B��$B�*�F�26'��M`	�%C�^���L}�"�Z�mR���Q*䏕o������-f�(y�!�$C�Z7�C?�lm�eL�'	18u�d��@�b�������1�'R�p�Q"XE @L:���&��ϧ!�M��E���)��ݲ|ـe�G���cG��� ���KQ-
�\��y�Z<uw�(��ݾכ�aK�|����I��]B�xh�H�.[�@�c�0+���I ��R��I�o4-�B�;�3?�c��b$��0A��rr�T47�N=� ҟB6��N)$�NU[�K�j6�A����E��R*O4��D�C˾�9 �NW�Qb��҃7PL�al�����Y5I0�DJ��	���'0�>8ce�Dƴ��aŋ>]z��V�"�-��S����be+��`��k�>h��ɕx8��:���8�qc!���|���6���P��4X��UC�>?a�*m��m�VNH?
�.�x�F3ޙ��o���@h�s����V.�Jr ��"����;�O� 4�E5	.�߈�f�w��u}����Բhf}#��G~�WG߃O�R#0��7 +v0�t�2ovUC02�`���.I�h�T �ՅGmv�I�=�(��O,4r��̫����D�<���Â8b���UD/i��A�=?+��c�F��YN0��&��8'��"[�o�Ԉ��xRg��m�|��w%P�7�^�,K�@��7 �7H;DٓR�]�۸'��]d�L/R6�0���CЁ��>&�	�I�{˔l�D
�h.ȨP!�S�vÆ4�l�K���<�7,�H���Ƣ�>)����r}�1�V�B~2��G��hy�mF�X فt��U��\"f`�5Y�v�����J`��yE
̧f`Y��o۠^T�oY�1a����,\��4�ç1/2Q�3o�%AҰu��lٲ+�yI3��?�nmj��Z5̌��Ж7%"M�/���}��̙�(�Yͻ[�
�xf�̠Q���H���C4�����f]�c�� �<����[4��Rq�B�A8.�mp2i�	^�r���	�dp(f�^"�h�����)f���r�D�����өE-Q��z�i��*/Xj�ə�*�:bF*`�ܙ	�@�6H��It��**�bh���\�T`D�7�۝@�Ҥ�B�'��ћt�Dj�x��)b3�z�'�Ԁ�1�Ǎ2�Z�b��ڢr����̻Ld�8��E+g:�JG�޽H�NdB�1T�"D!@h�$�O��Òm�#��<pW��:r��=(�&�`�΁pJ�<���G	(C��oB�a�nH�$,�p�i�5��Q7,)p`YU�^=Fu��)�O>H�𤐂��ɀ�

�mtn��҂�,n�8�YÝ+�����G�(#䪖jә!;���"
�ns`أr�n�ɜ;D=���@_sf$ �R�|�#>���G�C��(�3�O� �J@J���?�b�J��֮ND��q��\�ց� ��P|Ŋ��	1A���U�]	
cay�Ϛ�!�a�|�Z9��Ƙ�y�!X�r�,��T�	�n�v�[��BG��y�@� ��f��ը!A
r��x#��Y�t��@)�)³_P�>)w�7#��=Z����S� <�A�
s�P�r ����A�vn͏^�nD�D�խ����]�j������ƕM�L����:��U��NL[�xl��+u�+M�?��`��RrZT!����� �V��˒j�놝���_ Zr�he9������X+l0�,��GX/b�|��h�$�����-�2K}��bv��<I���2�ɈKր�d��`�l�D��\�I�p �bt1:+]y3"���arP��,D$�	��B�7%<�#!��s(�Z���3? Qq3BS���E�'�3/�$!*$��kl�`{�D�Fs��b��FK<��vFO�s�F8`��D�Gw��MR��X�O@��(4��dmd`aO
�'��h �(ЌB�n$qֆF7���0"�IF��ȱ18���G�N˂j�=+�zӑm�W: ���K�'9���l�?/�j(�m�S2�#���:�|퐕!J�lm�K��F+��BV���[���f3R|��i�"K.e|��U�J8oj�c�ڙD.��j�Z� �q$J)n��
!Sْ�n_0�M�Q�
�m��Z�Lқ42��[��
�O������+�8�9�c?cg�4�A�@GТ"��a�%:��V=Ga�AD�ʠpu�@�Y�X����L?��M!dn�! ��'�l��ϓ��tJ�˻/�N �FK�~�*��@��$2\����LE m�L�wϒ8�ljJ9*�\�֡
�<�ЮY>��e�H��)8��ɑ��� `�[ӊ<�D�=�c� �P�	�s�����!�&	�0E
#M�䝈��~�u��J�$7�^��d/_�+���A��e�曫���s�#�?�,P��;3�ޘ���-�d�;�A$�!�h��n�`b��8$WP?�5���[�H�� C=t�:Y�S�߈a�h�$ ��6X�3���%8B���AT��`Å<p�.u��Ğ�e�b�	�O7��{��X�U�8�H�Cٸ��٘�i�|s3*�%js�׿��Cw�V32���F���-�-Otyc@��]��agEv"�aq.��4���v&x�����BaC@1�9�h��P!5�t��癷@x�� �N�c�=*��>@{�MCD�N
4�6�Q 5�`�S$g�5Gv��P�N��H��Ź��4� Ŝ���9@�a��zUZ����9H+	3@B y+%�ڭH���Ã�;�v�A��RC���I
70���m��GM;%�z�,MqFƖ9~Ҹ ��
6�����' �GD�q���,w�ўX�A�40`�Y ��n��1B�$<�,#�Gu¤�R`�XMP1�!�!f�|Pa�[���y�����I�wĴ��k�H˂H�m>U�v�@;s�v��[H!��(J<L[T��9q?t��e��i�����4a Ё3�Ǟ_N1��(>IQ@|{6 ]�"����A��[L(`GJ�S�.���O(���%�|��p�B�#��#>� �)A�yvJ��"BT�`�2ԓ�2m���''
*#D�8�B?\z1Æ)��zrN��b�
b�"�ӵ��O����f�u��G��3^i
��^kmN�Aۓ ���s#m��]��$���U*�5�H�Vڬ0�0�O*I�H�c�a��[!�(y��ʳ	T���ܴ|��'�"\�s,�n�HM���H!��	hfڡ��O��2M� �pkG �i��V�[4LjNx��Q_��3��#��A�ܴO]�!��T�#��"��I۴��'.���u�
� }�)Bz>�jaD�8�\fA�?G21�#8���{�pJT�ưҘO|�tRtG2V%ܜ`D%��P�e����$L�FI:!�B3DRRl�1���	,.A�d
T$1*<SE�?a���d�b.�[�O'�����g�M�ҥ16�>)����ݘf:��F&���m�"6�"�s̀-
���Y���0r1�l�p��Dj*ղ��ڜ'o�GC�zb(	����d�PH4ˑ)�8M�ŠpJ��ҵ�O* ���ФA�&A�dT@�g]&y��b�)�N�q��Ƅ_)D�BDɞ:~��}j�
M -�ēQ��ي��G5{Bޭ��ѣB<�+6��{lz\���]�=�j$�N0dH�����5xG΅�3� G6�Ę,zh(��W� ���I*��{��'�2H�X�A��,��p��)���ã�Ⱦb$�9��0x�IJ�H98R�ػ���v�~!Ч�%���Ӄe�?j6�iO>�f ��^=ll�d�L�T^2�"7
Q`��Z���Dh�n�D��� F�(���顪�Q�T	R䭁���2D�4����X9p��c�@�@�>i�l�v���'Yz%�p���l���.B�r|��3�֐�����+�6(��9Qn	��	^�|7�\�2���'�.&rp�1��=t6��フ[�hx 'e'�Ot|�Qg�2(*��w���TT��SX�K� �b�+{!��` �*9���
��3++�����P@���K�M�����1.@�Q�c��R��2
�')�ax"�ͫ�`�0@b�W�*i��k���*�pfd
q ��!Q�5I< s�bN:�x��/�
��p�>�H6R�r(�<�|�"_�+Dܐ�㨜%Œ�s��X:�����M�A7F�2s�N�+�ɘUw�����ph*=7C^��*��V����4��]A�`&l[�$E�:�LZhq�%�;<O4!��ꑫ^
%�F#�DQ����R�n���@��h9��!%]?H�$	�vJ�(T��#ۛB\���ĬSj��Be$��vU�80� ]%9O�*6�:�O�jdKF��{����V�T`�t@�6'cuɤ��w�LI�ŖN@Ts�fPJJ��g̀�R�@L�� �4#ee���(4X�q��ֱe��%r��y�axҪ�"��	#wo)2��k�-�w�]Cb74y��`UNH�Yk�A��' �|SSg�P�H�%F��~~�A{w�mX�И' "�c�_%l�~ɋ�JI't�	N��W�U;"�^Ȑ���ap\����-}�D�SB��8�hz�G�2��%�R	$���c���p����/�zU�񈉯�p=�7��uNd��SM�|%t0
�)�"{4$<j��*9B�t��BF!&��$�����pDv��y.` ����y2k��zݤ���B�,}x�����v�ўp+$�޷)�>������"�Ѕ/��)���D[�g���ӻI"n��,ʀ��-�Ve�ywv����?K¶<P�ߑh]�e�WG�|��5a�FK�:2AU�ޫm?pq��H��'i���3}�����C�P�⡚fC��y���Z1�ܶf�r�i \#oN8���G)�U#��t�)�f�R(�j�2�!�c�Q��e��/����V�1,����)��<	�eR��`p��J�[���(����VV29a�G�'"�����
t��C��H,v̳���?DE���M�=��TbF������	��Uء�NE��``�P�KC�U�QW	 \P��e� � u�d�^d�h�ĝZl�LYMHK�yȁ��%T^��U�� �e��%w|zD�D��?C����.���̉$�O����	ҿ?0��Ճ=�Tm�#	k�4�;A9�B	�s(Ն>7ޕ�ƨ�>:<��ӈT�;�JY��c�m���3�r�H�ӽiuڤ��(��(�1	��A�.��'͊�M�4;�jh�OoT�9�K��fy����G[�J:����f� ������4z���d�)d�-!�(4&d#ڞO1�ͩ&��'R��S��=�hP���5��{e��8��������j��>dZ����-M=�n 0(M# <��Kv�_�=��b��K�gH*q��/�@�V�#��ϫc���;��{�ޑ����}�X "g�^"btN��=ak,M+�F��;�>��4O�?�D�3vF7%c̸�̂;H���s�E<bj(yK2��>�,���X!;�F�+��vypB �0i�[���$�֜ˌy2��0'�¬��+�>"�����1G s���8M�*��)3L�u���:��`���]�ְjs���n�h���m5�j4�O�+6I�a�v�>��x��gޑ+�D_�Q9�:s�|��E81@�Q����&�.�+OǮi*F�k�ߒR�ӹx=rE#�b�'�h b�딚M;̬��(�U��8EgǡP�F�ᤣ�Oޕu��	Uy`4Z5��H1ތ����y��Zg�����?l.�l�h�یP����Z�ɳfB�l�z���-Xc��a%��k$�d��V�َX��A�P���R�F 8������0���E�=+�t0�)�j^t��yihYd�Iî
<X���d�/Y"�L��=-@��+c���!L��ʵ�:|ɨ��˘<1���3���,^ ���wl���C��	�%K��;�BC�~������D1C�pW��X�X>��k7BB7}������5^˒-�5#�:q.2�)#���l㖕2É/lU2Ȣ M�0�\��0�>Њ�eB��X�I��̶h圙2�ɂ/mT0̲0�����wD�I��*ע��ga@pCJ�y�`L&�6�j!͚�{�p�DE��%>	̻<U,�p���� d�; ��܃ÅS(N�e��Q)D�K�N�<T(�@��~��P�xAN0�����yi���"GP��ÀGIQ����i�& b4%J�|zuL ��Jĉ�.��FR���`�ș2���*k|	��C�$xp��h�/�_��i�2Ɩ�x:L@���d	I��x���߸��dyAȄ��d!vc�D���!���^�ypHΔf?
�X�Z��p���@u�(��G#T��ĸ���
WF����ДUEB|�HZ�M�%z����,qh�T)��G�m{"a[Ր&�Av�2`�u[� ���T)��<I��n�8�%Ėj��	Z�LXd�O��X�'�I��@�"aю0 p-h�{�G��Hg�>�nDF���7Lϖ ����ap�%��!Co��A�0�MKLN8%�4�>�O�d���4&q��äUk�Y��'l6\SB��<M��Z��(���G�? ���)�n��3$�(Uf��g%9q�0%yq�ֺ?B���$غx{�qBR�hOb�eR:D0�/9LM@!HSm��#��z�aD=<$����kJ�AXT���&�>��=���m���Ad�|-(q,B��yc��Q/y#~�1"O؍C�(״aA(-�Q�Ɓ`d�c�	�:t܅K��z��r-Ҍ8*�|#�B�=`�C�ɟQ��I��X&��凒<X��C�If���S��W*���uÑ7}�C䉩x��a�)͛;��x;�g	
�C�D��0a�]@zd�`�D8&��B�4!k��y�*�--��#A��U��B�ɊQ�TP7��+-���E.��wN�C�I<k;�����V8L�@A��	3�6B�V��;ei�.ņ��$���=�C�	U������J�d��|T���'|�B�I
���3�)S�}ٸ����(o�LB��5ZF��q�M#}�TP��"�<F��B��2�f�_'|��P'/ֲV��B�ɰM�n�#�/SK���O�1K�jB�	&[�Z��u�٥.o�h:�Jؐ
όB�I�8�e1�OO@I���򮝹j?�B�]o�2�d���5�T#A�~B䉆J8�1�\�H�p�Z��
C�I�F� �b��1�R��GB�^^XC�I
kT"����ór�b�K����C�I�.���b���-�xX�G§\��B�ɾz���cab��^�EJs�W`pRB�ɒ0�t��S0����#0�VB�ɢ]D��w�	K�!�HN�`B���ܤ����FiР+� FhB�I�}J�# j�ؼ���#.�^��W����Ha�gb�>���ŚzD� 'U�(Q@D*˧[MR�r���8�tZ-Ol1A1��0|�R�!�@DZFBJ�%B�! ��R(M��I�)��!��&K�Q?��K�Y]�jɄ�0��!��n�T���H'��q�,�l�)�'F��ak6��"s'4�)E �:�6ec�	]6fRh):gb3���:�~2��߈R~���THg]���˗�SY�'ϸH��s���h�e���h�K��y-�EO6�$��Nľ�b>��!N�X�$QJ��u\���7}�ȵH����y��^�JZ��s@%�!z�ȩ�Ҡ��<i���ȓ!Tf�j�VF	������d��g_���d��2�-"�M�e4�݇�J^�a"hL�bU�C�[^�(�ȓ=�8q�e��i��i�7/��;��U��`XP��cNƏ&}�-� �Z5(
�Ԇȓ設S ���.4a�-E����ȓ5�F��+�:��q&�Χ?�\�ȓD톄0�G�p�sF)F!q"����1��Ɉ�ɘ�Y�лi�8�x��E��ˢ-N;P/p)�e��=^6��ȓyN���D"�2:�dA���=x�h���g�L��ՅN'��5���*�1�ȓrXz� �A�J-@i`�*_�,`��_�");���Nئ\����:�8X�ȓI��:R�F�P<�䋑��#k��ąȓ^6%	M�?a�%��A��)��cd����ۃQ�@X���Y9�2��ȓn��K%���
����(*x�ȓY.\��$R�%y��ʀ���xPb��
ޝ
��}kj�
}�I��{�M��K�JL�R����Z���v�%��.�81B4��J̤oY�D�ȓg;z��� 7f&�J�I���Ї�s�����L�s�����W��݄�Ll`;E	�-�����Wb�U��S�? 6��f�5W�Z�{� Z+4(4ؙ "ODq����24�-t�W�K���H�"O�(��_�&��X0�´`����q"Op�K����P����a�����"O��(���k�8`�� h����@"O����2��q�f�ȝ)����"O2�K�G�D�9���έJs<P""O�|R#�ܬO�F-�.8e\m�3"O"���$��B��4���"O�� W�m�6 pn
�TЂ�"OP�2��>0�|�d _o}2Uɐ"O
zDХBi�� ő�4c��"O-#2�'e�Z8���	�yct��"O�q��AW�cU�� �o@PKV�С"OҠ3h��'�`���$]�d/܀��"O��J���&�h�s䂌x�X#3"O@�u�� [@I����>��U��"O�suoL���$�橗g��yU"O�s7aA�Z'R�A4K��3���p"O4]�.�/w�+I��7n�10�"OR�3F��1&IP�b��@�[WY�w"O��Q���0W�qpG�^"!���b�"OT�q�@ԙf�0�kkZ��"O,+P�ڝS 
��4-%&6]Q"O\�2�Q5H�P�Q"x0�"O�԰��G�R#.��fL�_ܪ��"O��B@-K�/���q��'3��9"O�A��J7O>.�Z��J=��u+V"O }0⥙2<cd<���Wm�diu"O%�fZ�K5P�t�̍b�����"O$�@�B0[R4�q��/h�>��"O��BU�дkY�@�E�ٙ8Ҹ$!�"O.���dՒIj��a
�D"O��vF��.�1�c%tq�$:0"ONĲ�	�L"���b�1J7�h�"O��ۑB)�ژr�a�( ,`�"O = ��D�!9p��d���8R͐R"O�y
 n�2&�{��X�f�qAS"Or(�$ѪY��`1A"��z!�M��"O��X�ț�M�\�$�
/lh"O4�s!I+	:��!�AH�0��{�"O�$(��_ >��݊�S'�X�r%"ONY�d�&c���k��oF�2�"O�8��)�1t�\x�5%H�M^�W"O�ք(��rǦT�`!0k%"Ov�S%�p�M���4#h��"O$���^�)���P�A��"O}{��m�z���ؾv�P5	7"O
���E9j���&�) n�p"O �s�Qd�f��P$D	�	!"O�]Sv�9�������-Ԑ�Y�"OD���VM V��q�C4�n�I4"O-0DIF�n�����=,���{�"O"����0	0v'<@�Hr"O4{e���t��=bW���@��j�"On0�PLθ!٤�X�'�/zr�+"OP�@�ؠ"f��TH�Z��"O�p8#�ٛ3�  ��o"�`I2B"O�9��vC&�{��E
#��ٚ "O�Lq����M��`���9|�[�"O�Z��?Jx���O�����`�h�{��N#G�����E��
�H��my����1z������$%�Ć�|�*�p�	��,t��f�]q" ��S�? ���<}&59���1�xHi�"Oz!��ܤK�v���m�?�B$�V"OXu��b���b�+R�U_�q1d"O��Xb)סr��pza��
vE\@��"O,� (T>u$t�A�bI��9"O(�� H�m�P=0�A�946d3�"O6y۳�G�}�@����v(�D��"O���@�d���Kb��#��"O�d�����<P�pvK�D��2"Oh�h��\:/���W�?�}��"Ot����:7t����B /ٸ��"O�ݪ!������*� k@͙@"OH�YR�:"_��5ώ�G
�4#"O:�#@�=�H��0�C)g�eXG"O�@��*m�]c��(��H�"O�d@��������dB������"O�����8�xH�'�E�JK���"O�!"�m�4LS�4�wl��"G�4Kb"O謁s&H�?]"���76J��T"O����Q)Y�Rhk���G2���F"OT�˧,ӴX�� #�X q0��K&"O\X�*�A%�X9��!l�y2"OZi�j�!&���kЄP�^�t&"O�I��N��d�S$Ӽk���"O���A�?_�2H#��ػ�*�2�"OD�3�I���Y���-_pr<��"O"и��éQv�E�E�Ik$a1"OphY�G_�w�J�+��� Xr��h�"O��k2�8��laS�""^�aI"O�㑈�""B��豊 YBRmS�"O�����	]`�E��,�"OR�X��b>~	;��C=Ny�ar"O��$�Na���� �  !T�]��"O4�1$M�޼x�a�-V:	�G"OH��u�Ue�^�8Fc^�L�ʦ"O0(����4(sD��8>;T��"O2��q"�'�����f��7�$�"O���6l.@��1�$�1/ -Qq"OyX�.ޓq��t�P�G�	zI��"OJ,�g�.%��QV
�%�"Oh;��ɳ]���F�Q�0�0�"O�(����s�8��� }�d9�"OPD��mX�c ���ƈ?�v���"Oz��j�%0���*�����%"OVSDؿrP<e:�Z%q�"O֐!4m�9Y��xb&bK"�.��"ON��go+T�4�6`����&"O��J̞n��`��!�06�~!�"O��AP&�ua3��,%�V"O"�p7�@���΃4q�p���"O6�j�GT1tĨ7�+D���p"Oht��M9T<n�XW�8{]d�"O���"��R��U�D0Z>�D"O6���g��]bZMr�"؅EG�i�"O~�VJ�����ͪJՄ��"O�� ����@�9Ҁūe���!"O�Zb�Y�~�8�CF�����v"OxA�5�ϦM�`�W[?~�
s"Ol]���=qJ�I���p��q�"OTU��сr��5�e�,|�8s"O~h�փ��s������N$�R"ONl{҃��}Q�N���1��"O���4+M0y� M�O�{ꄁ"On�H3bå_�@5�Fg�&�zI�s"O� ���a T>�(]F�F-Lg�DЂ"O�mucR�N3���dD�3ZL@"OR��.ӑ,���B��/�Nt��"O0���,@ ���k<��	V"OZ��T]�2(J1�°I��b�"Ot���N�I]̠�"��/��4P"O�Ya�䝡%�p+���
Ni�YQ"O��T�I#@�q2�6dd�)F"O]0%*̑A�9�aE�B��8(2"O.�{5�Z��T��fĠY�4�:g"O�|1�jv�[�&^�P��u+s"O&��E
��'"��`��&_���r"O��k&'BO�v�$���e"O*�h �R�E��q��!%��,U"O�5��Ϛ3�VL�� d�����"O�囒�Fv�@Sj����"O���4bٺ1��@_'��B"O�H��Ppy�`bC&2�ڠ-�y� �d��š��م!�s�n�r�'}�+ƎS����5�̠�(��'�ȸ)'%��Z�����M��i��,#�'��9� �&Sະ{�N4a��Q{�'�"yǥ	2����C�\����']]����V�����%� V���R�'�� ���ѲQ�� �C�:~���'۸x'��<�L�ccE�/Jn���'���!m�v���N�(��s�'��U�(��FpVE�R�Ѷv*N �
�'Qb�9��|t�"�ى���
�'��D3��Üxld�u┨d:Z�S�'t(8W��2ڴ$�3rN,��'զ�G��KgBd;/�!*�pA �'^�ؕOE[5���cܭ!�ؕ��'(DB��[c�hZfB�/M�<`��'�ʝ"�̋�E(j���P�����'�@$�!L�!&4���w��3	��2�':���$��?(zL������R�'AH
 ӤMS �9f$��|���'�zF��lt�0�Ą��t�����'Ɋ�C��1'Q�9�D��l]6e�'�4�s���=~J�C��$HZ�'~(�)s��%ErP[c���`��c�'x2�Q� �"�I�O�<[�����'p�Pd�5-�T��u#�(M��U!�'�$eكK�} ���᧐�p�u��'�"�J�)�WˎU��D��HX��'ְ���n�/2�.��"�W>/���'9l�S�@���)U�Ђ�L���'~�P�R��\uڥ�Ɖ��6�@�'���B�dI0s���;w䙽�(��'������B*D���E+O��q��'��0����<�����Aiz�"�'贡�H�j�����8&�$�	�'J21��]�.e� �s�W�.0��	�'>��J�A�Ug䀊 	Љ �>���'�{ע�z���;�O�nY��'jv`HSI������`�T���'iph���Ք5B68s׍��U��89�'f���Eߍ @0�Ɔ��9��Y�'�� ��Ǭ\��p���ҐG�:Y
�'��i�  ���   �  �  �  '  j*  �5  0A  �L  "X  hc  �m  6t  '  ��  ֍  2�  t�  ��  ��  t�  �  T�  ��  �  V�  ��  ��  )�  l�  ��  ��  =�  �  �	 F : ]! ^)  1 n7 �= �C �D  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr�	p>!��L�>P^�x�#\`yq�~�tD{���O(dG6â�ߘ<����F�N�B6��~�'.>I��]�(��d_�R>`��	&D��3$l��� ��'y��T"`/"�	�|az�H?X̴Y��ǘ^�B| �e �x�@�?	hlHG �*&���ɵ@�<A&��H�'�T)r��u����`��/T�i�'�S�č��F�P�+ 8x20��ĺ�y��Y8#N�P��1�P	�BL��'�)�s�Y�1~"AۇlX<�XAL<��8h�B��.z��s��N�@�}�'fvM$��E�d^� jSG�>l%��ρY7H03�,D�������b�]S�lZ�r�̹�'i��1�	��~=Xc@ѯMb����ėL��Մ��?�Ox��W���`�~�p�B��>eBV��H�Yw�^�]�*�x� �nN}��/!D�����^����b��WL����O�B���J�l�٧�QM�H�R�ϘB)&��$:��«z��u;!L��;-�Eaș!��5z�y���6G!���.Q��G{*��\�Ǭʓ��-W��S�ə�"O^���.ONA+F��6[� j���%|O0`� �B�v�ڍq�ڂ�x��i�ўʧ`.Z��y��V�k����=y����&j$�y���^9la��&^r�8Ql����)�O�yA�B��6-�Kd�+�j���yrj�8tE�Q���T�*�2����y� G�g�j)"q� �O>&ݚg��,�yb�D�#ˌa�E��^02}RgN���'|z#=%?�j�a�/>o��rw���b��}�S� D�DjF��$o�`t
�H��,�n��1�>��p<�R�� ��x�h�&RI�$��`�<)Ǡ]�S���C�g]wh(x�ԟ4*	�)�d�p篆%%Æa��*`��H��Es��:u��n+���ᑧ y���A�^89�`�<�0��%kwL1��9MV���&̟f��CƸǬ5�ȓ��q:��Ϭc����U�� ���԰�&]/+�d<sF��4�.��ȓ׀)��[�A���Ȕ!d�(U���Ҡ؄�P��3�ǶnO�B�I�'F!�6�@��$ZB*�!Q��B��7s���$�p��� !+ց?��B�IWL����C��sT� q� Եa�B�	�23���BK�8Uzuq1�S���C�)� j��Q/�9�1u�M�I��Xq4"O�����	_��K�	��7���"O��L kމ����-u��Z`�'A�p�<iڒA�Z��N@W���H�n�<�`kÌf(����B�"�j`�"��<Q왻Z���z�䛫b(h9`�@�v�<��4W�̅RQiQ2Ć�k��Ui�<yW!R#b�H%B�̟�`�.��M�<!@�s��@�B���$����L�<A�}��D���^F?�5�p�RK�<�3��-6�&�i&+��
��XGjAD�<��F�a�<:�B!|��aE��i�<��c]!ؼ,��&�06�ݱ��i�<10m���(C�I��8�	w/{�<�3n�'�$={a��;�\��3�	B�<a���zsҥ��F]5g��(i���v�<����~9zBd��W�.��!�o�<�擰a���N?W�t�e��f�<!4)��%9g��7iC���W�Z^�<Q7�'+�𛅏�6?:P��V�<Qt�t�T<Jb��Xd,�3"�k�<��a�?pY��Ht
�*T���Kt�Q�<Yv�H6�\xa P**�Hh#�n@T�<1�
ס�ΡS���)
ֆ�I�!�z�<AE���)4�1χ(U���p$_z�<iա@6��$�9V$0�q"�r�<Qt�]%L�4�2RF�]�jq�M�m�<�Se��\gX0���r�T$�6��p�<ɓ蝟Wp��2T�a��F�<ٖgE��(
@\��2G\�<ī�}ߖ�I�E�l�`�[PK�}�<�%��{�\t� ��>D��� w�<�c!H�Kھ|&�Up�!B�q%�C��CWx� �i���-���
�B�Lu�u�4�R�i��#Q.p�zB䉾^5k�)�T�p1�3L��>^B�	�U��a���=n(��3��i&B䉺k�����Īsx`y%o�'x��B䉦*I�ӁRZt��rD�<U5�B�I�Y�ș��#|�(
�� l�hB�	'���+ρ!AVy�N9}rhB�I5���۳Vm*�b�E~�B�I����U'Ѐh�^��-�B��_�Di:rcʸs�6DY�+T�O�C�ɩNQ$|2g��E��P�a�im�B�ɭQq����S�)���sE�9SzB�*�ع#́����;��â�NB�	&��
nLo��LXg�I2^B�	;����#�����e�KO�B�;i����55�R�Sd���xB�I�E+`�A��Z��h�'��C�I�q�Ґ����/~�Da#֬��0�rC�I-�H�(�ѾSJ�ҤJɂ$XrC�I	���w@�4�>0�BL�\�TC�ɚ@�B�� �� 1�I�K�)� B��T�@-�4OW?;7�ơCI�C䉄Bq�Abe"P�'&�	���	=fC�	3/&)9��]� (���Q�G�B�I;p�i�OӤ-�&��c��q�
C�I�4(��];y`�M`�/�8�B�I�o���3 �X�-"��G��C䉷s.`�B�S٦	9TΎ�8\B�Ie�θbu��:P0��'F7u�ZB䉃>Tb�"�ɏ%�P�āc6B�)� |��V'�4�H�P��-]�(U��"O^�3���h2j5�F��o�6hp"OL,�2��9<ct�AބM��A	�"O${)�+3�y��*��U�D8�"OJy���C�H�쨰1�
U��-��'���'�B�'��'���'���'�~�����|���ZW��tZ �'�R�'�R�'���'���'���'�jp�5*��I�x!�b�7<��'���'��'��'���'=B�'�xt �j	Amtp��@ИS8���'���'[��'��'3��'|��'���Eb֖_�x�b��ڠ-�b-Y�'[r�'TR�'���'��'���'UZ��)���pi�f�0,���'���'��'���'���'��'�\���A�SJ
hbB��,l��U�#�']��'�"�'���'b�'�2�'(�����{�f��D�;��'��'I��'��'���' ��'1�����^�p�l-X���}�Ty��'�"�' R�'fB�'y��'���'����F��
�1RN͏@�"+3�'pr�'���'TR�'2�'���'~&Y������ֿ�K"d'�'�b�'��'��'���'-��Y2c@6����P�y��tkS;5��'�b�'�"�'Z��'���'?�<�\-qD�ѕoSb�"&M3<W"�'���'��'���'�`6M�O,�J+"�I�F�]��9��L�I�*��'��T�b>�z����5H2�9+0�˩g%���R���J����O|0oy��|Γ�?)�&�$�<!ⱉíURȕ��Җ�?���{j���4��$j>a������<�N�IV၆"r-Q��F�.]�b�(�	ry��	p���w$̳+OH�����(3�@`�4^�,��<)��4�k��Ƒ:�.����®���Pg�ҡQh����O��I}���!�0��V<O� Y���>�<�2�%��B�� �5O��I��?!T@:��|J�{%> ��G(ƅZ3ƐC������D-����z!4扨-yx���'�[�p�h@�H�x�̍�?q�_����ޟ����D�2�T��#�	+!gZ���a��O^���!H����O9�?��g�O��È�^�	�#(��@t�pç�<Y,Ov��s����I�.|RL�<N��tb"Er���ݴGc(��'�b7�.�i>]�w�3iy��$jݵ=�����~�8�����	$vv�]o�D~�<�"!���_ۤ0 ��ʍ%.�aXW� O��8���'�T!��'6�i>��ǟ�����\�	�<�B�IԿ	����&З;��A�'�~6�F����$�OR�d�|���?9�B�,��òm,-h��VD�7M-�	Ɵ���w�i>��	��\8vƛ(J,p8�g�.�@���9��oZe~b�W5,"�h���?!6*��<	)O��*��{_�i�I��O�����O���O����O��D�<���i�V���'��鱓*	�{�N��':���kq�'��6�<���OD%�'�r�'�2�����f�:�f��Cd�_؉�B�i��O��M���s����߹K�S>�y��ʷYA�q���t�t�I����ԟ��ğ����Ń6A�䄃�eH�P݈I�UF��?9���?��i� ���_�,�ڴ��56��b�*ԴZ�I���0
w��AK>���?ͧ�(�ߴ������g$W�o��i��#g�1X$挞sD|�	�����O����O���^�L-��3��-t���� �O�V�1#E�l5�ʓN��ƈ@:��T�'���O�'��E��0��H	�hqDq@1	J�y��'��ꓙ?���OUR�Q#'�i2B��B���2�0Z�L�pFS#]���?1	f�'�t��I�4�	YW�MkoP#J="yx��m���h�	ßL�i>����8�'<7-.����	O�lu�EZ�{=���H�<����?),O��d�<)�Z�@��V"R� (��jW�N�����?�ԩ���M��'�����M���d	zo`��%śg.(�䭆KD�Ķ<��?Q���?���?a)��="#CU���D����\�T�C��I3��ߟ4��ɟ'?�I��Mϻd��ԩC�7v��Yxc�3[U<�J���?!O>�|*6Γ<�M��'o$�j4	E���(�pFV�tb-ڝ'�P�Q.�ӟ��P�|^��Sܟd8�nȉ@K����,ִ�,ږ�ß���ݟ4�	fyҠu���+�O8���O:d1�׿��Qb���	]��y*Ç"�������O����@���x����FBњ#l;?�4 �f���7瘝��'d��D��?1fO\�$�^���B��\H�c���?����?!��?َ�Ix>1C�
��7��}0��4C)V�J@+�O�n�}S�����<�4���y7d 7|-R��6oL�S���E�ɺ�y��'��'H��豰iU�i���	�?YÇK���HS�Ř|<��&�C��'x�	����I��t�I˟T��;4.X���']�:� W�ʳ":�'�,7���BT��$�O����b���<�'hԔ3<�"����Gla@�-��	�|�?�'�?���$z�M�m��U:FP�2�[�)M�Q���Dڜ�/O�4�dL��?Y6O�ON� !?O��M�R��m�4ga�x�3Naj����?���?���9q�=K*O<o�-y�d�S��� /N<'��}�B�eQ����M�O>���3��ן��	ߟ�!C%�L�� ]<>��� �e�	�el��<	�� ��JS�*��' �t��� ���g�#<Q(L3���=z�s8O|�D�O �d�O���O`�?Q�䬉�{D^Qk�f�8�R�9�䟤�I��|C�4���'�?y&�i��']�H����=?T:�	p�N�HR�|r�'��OQ��c�i��i�!�GI�!,⍹$@q������I�K�'��d����l���P]��07.ZU��uq��@�	ȟD�'C�7uD���O"���|27Cz5�8������@&&�T~¯�>A��?�O>�O�b�I�ˈ06�LRr�G5�İr�)�D~��p�@���4��89��I�L�Oz=����>���C�J�?P8��@��Ol�$�O����O1��˓D��v��m��QҦ���Ti����"�F��y�F�'���y�T⟐	�O���\��FTۥ�X�q�U��(��n��$�O�5�4�q�F�Ӻ�%����(�<ᷥK�
ͫ��A�]� ��FM�<�)Ot���O����O����O��'V�t�d��"�=�p��M�"ೡ�i��X;f�'b�'�Enzީ�uMS%'��Tcϯz��ɀ"�ڟT�	b�)�Ӣv_~�m�<�'��+cW�� d� N�ջD%�<9ve�
A>��P=�䓉�4���$��.���H�zc aQ������D�O����O���E.Q6:��8�I����8R� ؗ���K*�����	"��=�?�T����ߟ�$��x�g^1K�*���Y�r,"'�>)3�&VǞY F�x̧RƖ�D�8�?�!�����q%d��r�KlϦy���� ������D�O9ǂ�U95�5�;���2���\}�`uӦ�Yq��Od�DMƦ5�?�;���qJ��B�ͱVϗ ����?)��?q��1�M{�O��S���1�*"fҋX���P���8�$��f��)�$�O,��|���?	��?!�6�� 2� I��ƈS��6�\�*O~(n�Fmj���֟4�	@��.A>�a�c�����"�@́��80�T�d�	i��|����?)4�X�{ծG��>W���SFC 1pz|0UM����O�����k���O�ʓN�^8D!�, >��H��1p��?����?����|�.O*�n��u�d�I�y��@TM�z��9��J�7d���ܟD��sy��',��ӟ��iޡ��)"��5ȱ@��E����Yf@�B�iM��O����������<��'��R'pdF�&��|0t9���<	���?)���?����?�����V�P�pta˴V#t	��%�T�2�'2�r�$���:����զ]$������0��U9���f��7�4�	����'ߜ�e�iY����z����t~D�s�g���կ&���V�oy����#�Fpr��_2�ܭ�-N�u����4\�$(:��?���i[�=J0z�C�@Ж$���:��� ���O6��$��?A9��
?p������+N�a���#����0a�3\6�����Jş�h��|rE��-B��`B�%H��4đ�)��'oR�'Y���[��1۴?�N����3;R�Â�W.O��!��N�?���'�����
n}r�'Q�is+��t��ܸV�ŧP�,��'�ҏ;Y`�Ɛ��ʣ'�12�T�~
eY�zl�S�Y� ������<�/Od���O�$�O��d�Ot˧��X)��N�&��E�W�L-wٲ�(`�i}6�ۂV���	�?��HK۟���)�M�;Bs8$��ۃH��X��͑!v`L ��?�L>�'�?I�i����4�yb�32�9��Ȝ�@�<X�b����y������������O����3"P4Q�hĶ����B>�T�d�O\��O ʓa��b�b��'!M�^ަ���V"H��5/&��O�y�'^��'@�'f�f� [�� z�`��D!��O�q��E�{	6M/��	j����O4)x��\�V�TX�A�3R �"OTa�爑SBQ�PK3�zM@ ��O��	�0Ժ���Ob]o�\�Ӽ@�S�S��d#ׇ0	��q[���<9��?���#�� �4��$�2]��)��O�����iV�=��%C�Q<tJB�'d��y\�����?]�	���	��;�b\�h,M�0�ڏ`�&q�5�nyrBg�~a�&)�<�����I�Op��Y	�.g#�;�x�x���crʓ�?������|B��?�,ǵk��m[��#T�]��P%1�h9q�4���W�U����'*�'m�	
I�JQ�E���o��\@CҊ/�����Ɵ���џ��i>	�'r�6E�gAX��M�$	ri�T*�8[�^19G�T^��$U����?��]���IYy2� (} Y�r`�
RT*i�-,U�!��i��I��$)P�OS�<%?�]K������nb��i�:7"4�	^��  �g�63NQ�w�2y�V�;A�M����	Ɵ����'�����|BhW�M:���Óed�Ԋ��/6��'����4(ş}��v����h�w?��s2�&+�|��AY��x��O�O��?���?i��L�>�ʣ͔:bZ�av ҃G��1��?�)Ov)n��@A�	͟ �	b��5\	ئ�.+�>A�t�5��$x}r�'��|ʟX���Q�b�N��gT(Y����u�E����:wi߸}��i>�%�'�6�&����{� ��Sa�-\"��,W�t�I͟���b>m�'հ6��o�
10w�X2=HI��a�V�\c���O��$SǦ��?$Q���ɧ�M��CK�Z��,#���//� ���şpV&���'���҉��?���� �=)��A�72��#�O�����G8Oʓ�?���?��?�����	I?$=&����	/�MS���)��DoڣPF�a�'U����'C�6=��g
+/ 0Q"��2ު!薇�O0�D ��IލU��6�z�x g�+m5H��C�zV�9c��i������O����a�Qyb�'��]������~������>HFr�'���%���0�M�������?!��
{���%�?�|����?�/O���Y}r�'�O����� .�����3fϲ�1s<O6����V�F�ԌQ�Z���S<Y bFM���!宊�x%���E�ڵ��;��^Οp��ɟ����E���'��[��/�.5�aیr�AR�'uF7��+|�4�Y����4�h� +{�!BK�q�x�1OR���O��$?O�6�#?���Z;��)�� 
LH(V�M�A���b�J�,!�H�H>y-O���O8���O��D�O�����e`n]�q�]:�H���'�<��i�f��t�'d��'��Oerb�Y���҅K��O�<h�o�2<X��?�����ŞF�h�r���+�� �R�>!�Z������MS�O����^��~r�|_��re�N<�.py������N�����ӟ�	��Hy2�d�`�Ѵ��O,��gbQ�_zxh�γ1}H�aŢ�O6�n�M�@��	���'e��PR�ڗbȴ�bP�8� ���A0=�Ƙ�@ ,ϛo ��%�J���-��CJ�pb�����L<Se9[X�	ş(������Iğ���y��6�x6#ǯ�j$�@�˙�N��(O,����M�g>9����M{I>iR!�&y�
J�d��!޵�䓫?��|�Q�,�M#�O�T��玺�
��0gK� #�L�Q��D���#�'Z�'x�i>M�	�L�I���0PC�K� ��3d�y�a�	ǟ �'B����-�	ڟЕO� ���h�R]�����Б:�O� �'���'�ɧ���(w�2���F�.?����𯑷5�^�r����!$B7�Bgy�OU����P@Ԁ��/*c�i���'{��y��?����?��|���?�)O(�m�K��3/&u>��*f,Ђ
8���gf�ٟD����MH>��Y��	����)O?__�T���L3�ʌˤ�ٟ,���S�@o�<Q��>�	�?��'^~ V�Y;����q#I��9�'��͟��Iџ��I�	���Z{�a	�;I��(��']�7m;)1$���Ol�-�9O@�oz���n�f0�@�����x��k�ޟp��d�)�)%n��l��<�P��fcЅ��/1�[6��<q6FV�ZK���@8����d�O^�$���|�����^a"Q��,
�R�$��OX���O��^��)K<0���'b5S��� z_���E莕;b�O>��'c��'W�'	t2�%�^H�7�p8�]������ !7�|�rc>�	r�O�D�5-_$�3bo�,�:�z1�F�z!��ڠ<��X��ݰ@���+ɾDb����ş��7��O������?ͻ#�X����'?�xU�äz,�Γ�?���?1�cC-�M��OB�2)���d�<C���>V���AK֚B/�'��K�'R�ɋՂ� $\e��`�a��O �I�� ��OB�D$�ӝ�^h���Z�<��*ۭɶ���O~���Oj�O1��m��e��G��J��V�(�ޠ�0Јs��7�ky�ŕi�D�������$Ī���F���t��t-��@�`���O�d�Ond�3�r|�ʓ��i^�^%��>j���/��p��[��[1^b�m���D�<���Lg����0�'Ed8���Z�9ve�9J��(�7È$��f;O��$����X��<$����)���IF�s.�x%O�Q�r`��?I��?a��?a���O����F5["99s�ʇd	$�B�'���'��D߼��)��$��ѩO�c���8�d�W�Xɣ%��@�	�H�i>1�0��ѦY�' lt���B����O�c����d��g*���䓲�d�O��D�O��$J��������y!�G�=F ����OZ�Sڛ�Tl���'�rY>�Յݾ�©��֤b��)X*?��W�(�IΟ�'��  �|9�ӽ{�(�����dǂ� �ė�.�����A~�O,I�	��b���yR��M�=ZjI=vA.]��Z
96��'��'�ʟ��R0��<�"�i�M�EJ t,�Z(O΀���]��"�M;N>��'y�	Ο�Ò��p:pq��̊ �L���������Iw�vm��<a��|�Xt��?��'�j\���o�����Ə`���'��I����P�I��$��P����$1̵��� �����!2�7�� |Q�#���O��D�����O2��J��wΔz6O֖#���$ˊy��	��'sқ|�O��'h�P�5�i�����\�p�荒+x���PN��x��E
�� ���֓O���?��.��#�퍻O�=��D� A��?Y���?�,O0�oڈC����'Djȝ2 �����!�BT[�M �"��O�5�'@��'��'�Ʊ{���A�����K�O"���!�7�Ta�S�	F���O��FL�84��,��2��굉�O.�D�O�d�O��}���^dT�t�5���j֧�8!Y셊�W���\�Z��'��6�4�iޥ ���傑J +2h����q� �I����;M>nZt~2Ȋ<�i�g�? ��cr���.�� Jti�/$A� ��2�D�<����?����?���?�Ef֮:޾8y��%>V\I��\	��d즱���J۟��	ޟ0'?��I�w�`��EV+$@�`��
�,�O����O��O1��$;`�0/F�9�'�>��b�/F�Q�̈Q#h�<���>�H�� �䓒�䛣4�VD:�Ԭit��l�p{���?����?�'��D�릭R�J���c��E2���ʞ{`qP�e��0 ܴ��'듍?���?ٰh_1�hJ�C�	#-����eJ�um Q�ش��dK�>i((�	����:o"��*��ݳ�zX2w5O��D�O��D�O���O��?)"!� lt9��t+��; 'Kџ ��՟p �4^x`ͧ�?1��i�'ČuI��5j�y�V��
((|R�'��O�����iu�I1cs�9�͵J=��r�N�auJ8�a�ɠAc��6�$�<ͧ�?���?qQ�ڸ0�x�r�)M�9�6���?����$����agH�ԟ���\�O�h��$H���j����a�����ӭOn�D�O�O���yNp�@�_(bj�Q��^�DA��䄞mTU#� 3?ͧ5
��� &��e��ث��� $m���T�
�Ii�<����?����?)�Ş��ğ��q��$��"��ӑɌ��y�D�8 -�'�$6)�������OX�!��
2?Rx[f�S�l} ��ъ�OT��ƌ$f6:?Y��ďߞ�ryB�\q����܇#��۔u��d�<q���?���?Q���?�)�xM*�"���*�H� 5`���g�����$�埀�	۟�&?��ɞ�M�;P���a���QN�A�@��8~:���?9M>�|�5IE��M�'��m`F�8gL���
E�q�'ƈ�r����hQd�|�P��Ꟁ��"�j�f���B	I�:�Б��۟�����jC\Xy2,��`�aA���D�O�̐V䈅���o�`Z�W*�O���?	c\�����%�d��MȊ��x�g^����@Je���ɓ'%�jE ލ
�E�'M�������:��'v�!(���	�#�n	 ;�4A��'4�'�R�'c�>��I�p�NI`�C �x_T�14hRሐ��
�McQA�*��D�����?�;���?j}rd�7WI��̓�?q��?1f&��M��O�7]K��� =A�@<[S�	n���Xpkx�n�XN>Q(O��D�O��d�O��d�O]��lԵq������#��6�<1��id�\���'���'��O�үB+s�Ir%\RI�v��|�4��?I����Ş5<Dej��� rRPh�ca���x��f�8z�(�`-O
�2���?��<�d�<�(�3K�เ�E�͌ ��Ş��?���?���?�'���F���Qh�����D���r��C��|�Ta34N�̟`cش��'���?���?i��(2�!��i	���2M�>��)��4���������Ol�O��Fܷcr��礂�9���ӳ#A�y2�'|��'	��'A���U�y���ea̸��Ē���w�T���O��$O��h�Iv>9�	�M�K>)tEϵ:):�P�H��%~M��ia̓�?�*O��Z�yӮ�BW�\c�T�LX�B��.���l
�4D@�$լ�����O����O��d�)2� �E�I��<�f���*�����O�ʓF�v������'lBR>�h>z����b([4˪}D<?�wU�|�I��'������S�A<S��@�#IE�n��Y�q�+@�B��F�H/��4�*=3��&��Ox4uh��G�\Mi�̗�P��e9W.�OH�d�O�d�O1�F����ڪW�DqT�Z(0�(�s�ɭnl�s��'�Ҩ`ӄ�XR�OB�$�K�|@gK�pFN@Q��V�R���O�`��GkӦ�Ӻ�e��7��Ͽ<�$A��Mè��w�܄��u����<�,Ot�d�OH�d�O����O�˧>b�J���6x��:V�\� �iyj�ˀ�'V�')�OUr�q���<i�z��P�U�,�(�T��u�j���O\�O1�Dٺ�}��扨'9� ���ߐ),����ꖵ�l�I��Y���O>�O���?Y�0g��(��Q+\�J�V�����?	��?)OplZ}{|��ɟ���C��r�/PJ �b�)��.�ȴ�?i#U���	ʟ�&���F�4U�āѷ��q¨��B<?�/�`}���"G���'j��œ�?�3D�n��18�@	�J��S����?a��?q���?aI~�B[�|���$Z���'B����#�a>2M��Vg���T�>��'tb�'��I���7�ְ�AeX F���QI^0Di�	㟸�	��\����ϓ���L^5En�mM-+^! M4��U#���y*2�'�P�'�b�'=��'w2�'�b��\>zZ�j��QXT�KR��1�4=ތ����?����'�?!q��;Vn �R�;!?�)�v�ˏh������t�)�[Ov�p��� g%��*�[&kL�q�gP+7�"(�'C��0чޟ,�0�|�W��c�a!RO��B枥�������	������hyrhg�.��f�O~�dĜ9P.�Um�&f�*9�&7O�o�g��v�����T��ퟐ�r�XJ0����6d���{VnL3+�^%nZM~�ٲ1+�PF��w^\=�#μ3�Ԙ����JkBlj������(�	���	ğ���덺q�|�
���5�	ӱh)�?1���?��i�a(�O���h� �O���A�3;Iƌ������<(���*���O��4��Q�7&y�j�+��P� ��v���aWhUb��N�A�lp�͊��~ҟ|RU���	П���؟�*�&]	:C���3Ö�p�� �g��H��Ly�z�8��.�<�����^m�hjW��m���rW&Ǟq�ɸ��$�O���/��?��%搟b������iu/J�ZL��v �	��FA?	M>g/ �(�QDY�R�D|C��
��?���?q��?�|j,O�io�(c������4D�����BJ<�┥ΟH�I8�M���o�>���a$6��	��D����6�
H��?����M��Ond�Ǉ¼��O>�Y3���aT� �˟�V�
�'�������ܟ�IƟ�����ӽS|��oD6�Z�P��2J��4$j� ��?	����i�Ol�D�O�n�7�6C��5|�L�*rM�[A��d�O
�O�i�O��d�"R��7�}���# �2 ���C���(u�j�
b-g�,����$���6��<�'�?A"aG���%���ͣ|���A���?��?������������T��ٟ�"f M.h��W���J̾��j�o�\�I��	J��I�I+r�$�:�O
�n�j�V�I
U#S�M�d��4�Fg?�����<ː�\�����p\�	r���?����?��?�O5b�9E�'�K�2*v���q+��,�����z��$��yچ�<��iB�'(�w&&��dd@�D�0	�&ڳ�@j�'�R�'Y���]���3Ox�M�}	���'r�"44�H�ʩA�CX%v(ͣ�"���<ͧ�?y���?���?��̸E;� ��Dʆ١b��z����M;�eH�����O�"|�$�*M�0I �D�c��L�����D�O��i�ɧ�O1�9�BO'}��y�%i~���� �2}�\��O��(���?�t%2���<�Ջ"-�	�%H�i��\�(A��?q��?q���?ͧ��DW�+�V�@8`��"PN@��P@�}+2.�ğtz�4��'�@��?����?�"���;֦PQmB'?F�`,�:!��}8޴�����M��؟Ғ�����]�5{�-6�����!s���O4}����OH���O����O1�p����	 b� *p�T�S��MY�(�O����O.Uo92^I��П��Id�I/i���r�ߐTd��F�F�v��&���	������+C5o��<��^�8I9T�ڂY�r��C8��\xs,R�F��d:�����9O8�X&���[D4��c-��?u�M��ɿ�?��kП`�I��4�O$6 �U�� 4Flc6�ʞ8��O^��'wB�'7ɧ��UV�r�в�T�_�)p�Z# N^�`)Ίc46�Wly�O`T���k�܀��U�EF��UeF���EX��?����?Y�Ş��d���� E�r��jT�P$����%f8!�D���J�4��'�L��?y��4�����u���a.��?��X�F�!ڴ��dưPC<��Ot�	9�<Lb��ʬ+6�T�⡒=bz�,��L>턼Z�BJ %
iCg��/0��#�Ϧ?̴2c��3~BČ�SN�{��fC�x����4�z�@sA��v�$�ė<�P1Ѣ�A#:�#>i�O�5�P�a�h�"| 8�%ɏ:.M�X���8�~xbW��(J��xC�狊!� P!j�,`9p��ʈ0:e���G���G��iC����`�£Lh���T���8;��� Jr�jťːS)�)¢���\��ũX@�\a�b&dS�M�!zF0����T�j%�Ħ��ɟ���?՛�OD��Vc�	M�Zy`��F�:z�@�i<2�(`�'��'�3?��	�TH���@��]H��A�@պi�R�'��`\���d�O��	�\H���Ǣh%eHDJ�� ��}b��',I�')��'w�'Z�z�3�1-WK--��y�i��*[�-��ꓣ��Ox�Ok��lV� dED�l]t�)�@��	��3`t�l'���I����	qy"J�} &���	��$������m��M؇�>(O��d9���O��$�#ٖ��U/OZ؀��T<R� �[���O����O��ǂ�'>�^��h��M�Bu��c��$��(1C�i��柨%�h��柠��A�Y?�0��b �p'��yTtc�BG}�'JR�'�	
�f�#��"��-����-G|}��@&�	g8��n�ßh$����ß��$�R�	��a �T�a�,x��i���n�Ɵ���Ey��p��꧉?���bS�g�D�^�n9^IG [W���3�x�'��`E3{���|bן��hrI��W䩳gOƀ("�([�iL�`Wh
ٴ�?A��?1�')"�i��f��|&e�[�t�&��@eӮ�D�O�l
0�OȒO&�>�V�*X�AP�#T���(a�d�:�k6�����	���I�?Ѡ�O
�R������.�8�Qb	�+R ��i�x`z6�D(���Hh��>����ͅ�; ���'hٌ�M���?Y��c��)��]��'F��O���e�9���Ӆ=��ar�d���P�O����Ol�Ė�X�rh o��D���� ��{���mΟl��N����<�������p@߅T�nH�T
�pt�U���G}hʠCT�'�R�'uR]�	GZ��3K�7p�=��g%|6`��O�ʓ�?�O>q��?)"g� ��`�+�<Y,Ih��>�B�H>����?�����x��u�'"XK�=)�P���l�61-�~����?�H>����?�B� B}�A�C@�ِT��-�"q�p�ø����O���O��G�`���R?��I�CJ��;^�(�H0*�%�
�U�۴�?�J>���?1N�ĸ�� qe�T�d��K70�6@jǷi��'��ɹȈ�K|�����N��>����NЮQS��%�,�'\��'}��yZw$dYb��ĒC�ܸ 0���d��|۴���D�>4�(o���I�O��ITr~R%Ï|~$�CbL\$i���(�M�)O����Oa%>m%?7��Lz���Ŝ7v��0�*3��F�ü��6m�ON���O���NV�i>�`2MC|��8�"��U� ��P=�M����?�����S��'�b�7f��ш5��@�H����DE�6��O����O,���_�i>Y��k?q4D'2<�s�ؙT펙��iSڦ-�	F�ɭ�������a?Y��D=���Z;�]��$�ڦ}���{�T]�'��꧉�'�0�b�%b�@�㇛�p�p]�m'�$Ј$1Op�$�<��S�hm�SbN�e����c+״@:½���ɶ��$�O
��+�	�p���Z#팅y��l���T02�@lZ�'�Zb�l��Cy"�'*a��֟б��ǐ�	�(��"Ϛ��!�b�iir�'�O,�d�<a�����q�s�0w�dx���%�<�"�D�O���?y�����i�OZؙ!o�=�5�Ŋ��hJ������Ħi�?�����dP��'�Nx���(,`L`�v�1epvt�ش�?�����䚒u&lt&>���?��:'��1�ߦq���`���J�rO�˓�?1����<��*�������TRd�c҆!U���'�r+ܚ�R�'���'G�4Z��	��EKS$��y�|�Qb�5bY*6��O��oDR�DxJ|�s̖2gR�P�l�˨�z�,������,��ӟ����?՗��閲~���q��:yt��k�HE�3�x�'�(4X���I�On��7���<�>	�ã�Y�,����������8��t\�CO<�'�?���2θչ�"�=p�Z�Br�ƼT%d�k��i��'I�I ��)�|����~� �A�>�,Li�R%��۴�?IP,�����X�������ЊJwYD}3��ȁc$x�'�t�� ?)���?����䑎?��ݓ��^�/�j�c��:x���
}�	����H�IqyZw&^�BO7tC�-c��Ԇlm@�4�?�/O2���O���<��hD���i�#�`����> ����H�Q���韄�	����'�V>5�ɚK����U���dvb�#g���XUF�j�O~���O���?y�Q�����O�����V��8y�oڸi�Z�Qǫ
Ȧe�?����U�'���z���3!ײ��a�Ι�8��4�?�����kĈ��O�b�'��땧PX��UM��X�t@I��Ĩv���?	���?aa��<�N>��OVBB�޷ ����a՗�>�ڴ��ţ=���lZ� ������Ӂ����i* ��G�̸��D'�0ꢽi��'�ڔQ�'^�'�q���q@H ,�r$zJ�-�����i�X�
��q�d�d�O����0�'[�B��M��ۧa���Ǩ~!F��M��(��<�����:��ߟhE�����v�!x�$�A!��M+��?)��x�����X�ȕ'���O�8�1*�> n�(+O�m�`���i?�W�<peeo��'�?!����4`D�� T�r$�VpD�`�g�3�M���6�<�Y�Z��'�Y�S�w��a隭CW�J )�:e\	�'*@�'���'8B�'��X�dS���D�R��/;n4�R�G�l�  �Oh��?�(Oj���O���
�%��P�b��*,��N��)=��xw>O���?q���?�+O�S��E�|jUÄ�l�@Jք�`�d�'G����'��V����ԟ��ɰ����
e��������7,�� �ҍ�ߴ�?����?����ެc�X��O*"�Ǵ)1��ZFXҵ��^�d$�7�O�ʓ�?)���?-�����ܴ?��(���-O�(�l�;�oןL��By�&��b�v꧁?���C3m����GÆ�C�@�[�IƟ<�I��PZ�)s�x�Icy�Пle�V÷v�)��Iϝ��r�i���5#��Z�4�?���?y��"�i�U��"E�Dv�P��_C\H �d�R���O�2f<O����yb����J�@�C�/�5z��{���,s�F�K>z��7��O��$�O��	~}�T�����.d� Cݒ5�\�a���3�M{pJ��<a�����-����`�� )9�,H0e��;1���R��6�M#��?y����Z�H�'e�O$ͫ�@�#��℃ Q���i}�I͟D�%�~��'�?9���?��OȺ}�� v���6X�HӒ�B�^��F�'|^�9Vi�>�-O:�İ<����"�5��4��ˊ��T!���U[}"䗃�y�Z���ݟ���kyB����Ba��j�0��C������>Y(OX�D�<Q��?i�����f^ry�pk��z���Ҥ��</O����O<�$�<i!S�]N��ƀ)��-aP��8v�n$��	�yI��U�4�	Dy��'��'x8�R�'Y<A*
�7M!�qPr�P(W���r�{�B��O����OL˓|_�,yUX?��i��r���n��Hb�ju�
�Ѧ`tӸ��<����?���4͓��i�dQ�0��2)����ߗ7� ���4�?�����$K�_��]�Og��'��D���kj>��V�X\��yW��Hc�>!���?���
C����9O����o� ���ɃLa��QЬDn7�<��'�2~��'���';�ĩ�>��;�T�[�H�5`�h1�CϛV2�m�����u�l�	矤�'rq�� �A;�@��
��gG�CfD�
1�ifLͨG�pӄ���O@������'���/�f�e��0K]^�c8&�a�ܴo�&�ϓ�?/O�?��	�XF\� �^���K�-H�C* 8��4�?����?��bNz�	Ny��'%��̗�:(�L]�R��Т�*ߍPX��'���'~$�������Ot���O0�k�'�(s�n��U�J��KЦA���6��mɨO�ʓ�?A*O�������*�*�h��@���h��R�0��B}���	ܟ�	���Nyb���@X
.�C�><���BB�qg�>�,O����<���?)��k]{M(s��`%.�3n'��"��<)/O���Ov���<!����U����&<�(��cA�h���a�*��FQ����lyR�'��'a  ��'x$�R��E�����92$���`Ӯ���O��D�O�k zu �Z?��5$��	�+q�
Q�m3**��4�?�-O���O����_��$�|n�?r 8�F3h>*�Zw#Ly��6�O���<��L�M��͟��	�?�� ��7f��xE["�D�pB��)����O�$�Or=8�<OT��<!�O�`�Q�\�<!f9�gZtW��X�4���U�7�ޭoZ����	�\������t�w�����P�� �'�L`���i�B�'�R=c�'>�_���}�Ul�f��Փ�/Y�{$�A�R̦�X���M����?����zV_�ȗ'�01a	\<��%;E,�U��*a�!#W5O��ĥ<���t�'����+82L,��T<M��mr���p�D�O��DBa/F��'2��ܟ���j���H�+y��E�O�:P mnZ� �	���㒨l��'�?I��?)��k!ܽ��0k�.�ApDPk��v�'�I ��>�.OR���<����l�we�ݣ$,��P����a}BcW��y��'���'c"�'���(E��� M:��c� ����&� ��ē�?9�����?1�Kd@5�.)&�S$�V�3}< ("Y@��?����?�*O^}Y����|�d�uR)ISP�c�����n}��'�2�|��'�B�1u�D\>��͈�hܖ`F8a���-��	������'YX�Ғ�(�	��
��@3tPg%��~���irӘ�D$�d�O���F�i���5}�j�6��q	��S#kϔhP"���MK���?a,OT��[�ǟ��6L���,ĥ_9Vy�U�lw�II<����?ylN�<�L>��Ocbp8g��	V�9k�.�9��ش��d��^Ȍ�m������OV���\~A�,JD����L�>��p�[�M���?1獄�?AH>A���Ɯl���rLlR��C���M󵯚�OP���'���'�tf*�ɝlR���)o��}�&]�N#|���4F�Șϓ����O��@=�h��Q��'[��%`@D�=��6m�OH���O�q:�gY�I���\?)vM�/�H�(e�(Ʀha�.[Ҧ�$��X��x��?���?�1�I!Za��
���_��͸U�#u3��'�Ęp�4��O���*���Fp���06V�@aL�6���k�Q�X���g���'s��'�O�̥��C�*��ƈ��)"$@_5N�D�H<y��?�H>q���?�V剁ri�A��ܦ745�w� -}P �����O*���OT�����7���b̑ (�0 ��Ɉc(���W�T���X'�P���h��w�� �']��]!�����6�Z=��L�'P��'��U�|+���ħ�V�)�˜�t.u!J�_@�a�i��|��'��J0v!қ>��(շ��5H_�s]Z�ٴL��M����?)O)��(w�Sٟ�s�� eI�=0��D�AB�c0]0d�3��Fy��'��O뮜#6bAᘳ]< �0�	
��v�')"k�6��'B��'��DR���{���ӗ)�jl~ِ��|<:7��O0�K��DxJ|�%d[KFT���u�hbƞ�=9T@	8�M���?����BQU�(�O�z0Q���-!���ɓ�K��H�Gq���d7��䓺?�BK�#Y���zd̆�K�rtK4�P!��v�'��I:JѸ@�'��	� �<��ak��I�+�m���U:�I�ħ�?����?9�-� Ҡ��ě!I�N%�1- �{K�V�'��):X��[��6�2�$&Ύ��so��05���䇜,/b�'���f&0?���?������B�)[��b��-C��a ��)H-j�ӣ�Wn��T�I��?���k ,|��d@�d���1��I���<�<9��?	��?A�O
6pH�O3��ϸ�	��ҧ6i�[۴�?	��?yL>�����%f���L�o&E�T�CW�(�R�Y	��$�Od���OH�>jM|��oN�B��Α,|��<
3jZ?U��F�'Q�'�R�'ɾ-��}Rܔ$\��ZR��,axn�Y1Z��MC���?��O"��K)��O��iH#��e0oׄ8��HR�	�&��Iӟ����>���FU	Qߐ���b�lޙ7N��M#�O"1pG%|�е�O6��O���O��Ӆ��� ��c���] ޔm�������G�\#<���'IJ�Ur�B˳J�X���?р�߉�M����?������x�' (�3����xq1�
A.*����+hӚt;q�)�'�?	�A�#wMX�bq�A3��E*3����F�'-R�'E���1���OH����x���h*�DAb�X�M���o$�I�|�c�X�����I΀ ��T*�9R��'��&�hp��i�2�[�~�c���IG�i���=����Qm��:�u���>!�aWP̓�?����?��O��h�n<�<�Cv�Y�3�h�K]6�c�`�IA��ğd�I4}�l�ڧ�?
�}ӵ�W���%xf�8�I^���b�˚#F^�E�to���Xs1�^�()��"(ͱ�y�`�>S�&%H � �@�k�����'���S��ێ[汪����wW&( Ek�>������.͎$H�	��'�(�8�
@9l��mJ��ȹ����	!�a�DX%:�^�	2����i�S|Q�%BkGkH���wq(����'dc0�gV�m�A�Wй=��25i��=�m(S���P�e�3E�_��Z��7H��Ct�
 K6��rWʉ- ������?1d��C�@XrÌ	?&z�k���wYJ�S@���ۘLl"L�ԥKۈ�*�����	<|�d��V��'���شr>`�V��^���`��uĆ�l���P%1�>q���'��iIs�'h2��џ,Q�7r���!�
ʐNN袃 5D�����"�D��c��)m7 "3.O��FzB�n3DAb!jôOB<܃3��?���'E��'yb$8B-N��"�'~���y7�M�&�cuʚIhDc�T 3-�X��IN�bYn���/|y��3"�|�o�y�*}��2�y�q*�3y��l��ޜ���dR�#������L>ņ�x֢Kb�	O>L�'b��?�Or� ���4퉖=J���;8�AR�_>�\B�ɼ#�J� L��4"��4GJ�%đ��'����0��j��M�,
�d�Ʈ.Ey<Q+��+H�����OF���O��;�?!����DH��(��t����)F���pfʹ]����1F?>�\�k'�'lOF}I�/D�YgM��`�,jf4d��꒔,������܌?m:I��I>������jZ����*�$��O|�d9ړ��'�N !�,2{��`<S�<��	�'/��fͯ7���f��0��y��>�)O��
��]}��'[�А�πRZ��Q& R�	��!��'j"�!e��'a�	�h+N�S��^#/����F �h2�쉯GA2(�2�ý+����I&�̹��.F%�l,j�'@�9��F�C� ��kZ�n����Ǔ2Q���t�'��1n�� w�LP�D�$6UZ�ҋy��'
$�˳�d�fxa�0�*��'��7�K�u1 ���OSS堬�"�>V�$�<I�M��A5���'��\>�R��
ԟ�*���13G�p��o��z�ퟜ�I�  �9��4������#��WՂ�s"�͏��)�N!}� ��(y ��A�-]��s�-�D �e�J~��&mY��P��2�Y��B��Իecb�'�7m�O&�?$k�+�c���/1����kd��'��V����C�p8��M�'��9*�����p����޴�?���i��k[4<�óC_�?���у ��듌?q�IR ���?����?�׿k����5tV����E�直Q��S�A�>�5��

��1�|&�|�l�nຐ"t�^�:����,"���X���#���W�q��'�$���c�VY�E�R��p�U�'"�ɭq�N�4�,�=їm� �T���N;b� ���m�<�F�E�?�i@W`[�$��\hQ �h~rA?�S�$V��3U&X�K��AX�G�	/����i0���j`��ǟ��I��@�	:�u'�'0�;���2���6KK��k	_�GT:�jC+��U� �FB5�O�L�5��^���m�?#$-Â*ƠKq����&'�O���7Q!e��T�͕+��q�Vt�"�'���'��I����?B����\���F鼹P!nO�<�"�_!]ߘ5�e��
x�X@���P̓��uy'G�:ꓥ?a��\�a�b�1�}H$ʴ�?A�Z�9����?��O^�|�&��*W�I���>A�mZ#4�G')$ l�S�#O�1q7���l�\�h�u?QѭʳTS�����s�[�N�I8�P9���Ob�$�<�c��bъ��'(�����p~̓��=��HS�}�v��a盺u�����	v<�i��`���48�H�����3YT��*�'��	,ƞY�O����|"�I��?IgH^��8�-ڈ@(���-�?��y�dE!� �.�S���*���'y��Ce�_)І�_�ft�@�O���S�\�^�$����I�#}�ꎗN�xs�m]3W�(1CQc��f��'��>U�	�h�
	��	�~�R�ԧ���0�Ɠ�% ��E`�Q!�T������HO� 1�����Y%W�V5�)�ĦU���<�I�kgbAUm��I����	��u��*
Lر*O�7t]Y�S1O��8��'��,*G, ZF�T�S 4��{�-����<���XO$��e-�C[�����<ܘ'\����S�g�'����AI� ���\��C�)� P���C�ܠP�l��������Z����n}P�&�N����8���x-�$8��?v�h�Iݟ�IƟ�^wV��'"�H�gG�x(Wܢ���R	C�̂#OD��4�Q�J�t��TC�u�� V�	�0!�тJ�:��hۑC,�40g� ���y:��'&�';��'*�O�a�.	-��q���s�B�"O�@+W.H ��Ӂ�Ra�P`D�d�x}��i>y;�ϩ!�B J���7�VqZd/:D����Y��5ؑ�ӑH~l {�6D��x�@V�S<d�K��̄1�^�(1g:D��Y�	+
�]k�I�*@ST,9D�4c�oV$ @���C�h�ay��8D��0`�_(v~<5pA�6lܙ�s 6D�Hڔ	Z�4��0aߑ
��A��6D����,`<��I] `��!��(D������>g	 I�)��t��IU 'D�ț���4����Y�d�($D�\���G����9��\�����"D�\"��1$Iu2uDC"lD��b�l%D��!��M��Xi�'p�Y@V� D� 0Eb�>s 51#�*�$Y�d�9D�@a����#�|���T�l�H-���)D�p`��>�`�; m�U���[��2D�X�U�C�Dp�Q��M�f��͐��2D��ᄅƷ|�>��D�K� ]��Zrh6D�4 ��N�}�2	�H2��H�3D� *��h�Xd{���1Ί9u*2D�� ���;Z�Y����~U���0D��1��L�g�@] �IŤgXI�4�"D��ꅨI�M QTK�.Dm�Պ�"4D�l�sdōjnBa���o|,��k0D�,BQ�
r*��(���-����,D�|��
�/o4����`��� e*D�HK�)�T ]sF�R��إ�)D��t�Q�v�ֈA��D6.��e��&D� ����r��P�G����Ub�2D���IN[Ґ)�sJ�\�8`/D�(�0��E��#'�F���,x�(D��iӭ�=��3s��i~�4�4D����C1`($aE)"l�|Xx�#3D�(�do��B/����^.��3p�$D����N�;py�-��a��h��ms!�!D���u��!n����O� z��)SQ	 D�`
��V��a�p�!m"��;1E>D�D���Ä.jRģVc�'`v�ӧ=D����bB�4S��q�EL.1n��$?D����Yp�x��y���i�e
$�y' 7�yp��Q:p�����`C��y"�ӊ1�x�9����U��D��S?�y7 Q4�� �O�n�QR`��yB���N�n��S%�Tx<%����yR��#㮉*3�ղҽ32�U��yR��6Gnޭ���v6^���C��y2`̝W2�p�U�@"Œ� 啱�ybl<,!�,B�ۊk� �˵n�"�yB�E	1cx�� ��c���2&"ʅ�yBgQ�4�(�`�&ۑ\�]ؕ'K;�yҠ�.FJ|Z�M�O�\U	_��y(M�?l�t"���@�ɹ�(G��y�(Y&��9be��Ѝ$+��yr�R5 :��FA�C���x��G�y�b�&T�{�DĮ?dP�Wϣ�yb��o��aI��	�I�&e�!��;�yN$F�3�U#F� �R��y
� ���3�O�g�<k��G12@��"O~E:d$FZ���K�O� ��H�"O��Iah�����w�@41�HD��"O�(H�A�D!"��e��O��tQ`"O�X�W/�./$=����k�t��t"O��)�P5>�$T�O�7���q"O�1Ru�W(��!�md|e�"O����#�!��,�TcvPA�"O��(�J�U[XQ��D�z@��[�>A"l�D��Ho9��i�?��rv�<#�L�|�T���ϊuj�����-����s�OM�L����|h�b�\��4AԌۄ	�N�"~nZ*�D4@C'�p� 5��3��>1�HE�<$@1��4Ě�S��B�jU��:��)����+yrߓI�dX�K0P��� ��Y��`��[���Z�+��S��$�a�G�-�Y·���L��l(]"��yǬ=D�xK����p����@����zRF;}�@�L=2]qu��/�v5�FP����~�����
T�<���8�H�h��ҵ*ߑCXa�s�ص$�ک��-���U�ֈ�}/�|	f��_��,O��z�-(�s����V�\PU*¬V�r������	�f�(��Sb=:����A�E�A�=�X��Bم+r�X��ÊŗPJ.]�D�S8�xkR�
e�t5��-�;��{�A��&��aSrGGc?�OԱ�?��t��k��4jj��C�J&C R!����frh�������O J�$�#+˘ȣ%>�Zu��Ò	��5��Z����\�~����H3A�V���Sސ�g�$-�}�%�
?p�2�i[`�� kPcO���'h�!iTk_�J������S�4�S�O�8c%��j<�qe��Ǝ��F��!r�Ȍ��g'���:��QCn~+8�1�`-#��D��=��y#'k ��1�#�_$��g22�Ce� ��9��FB�0V�lt`d_ 	��H1]w �	:!��F1�2'�W5��h�'����a3m�RHrQ��V��8���U 2 "F�Ƅ)'T����1l$���)Ψ���)B�Ȱ+ L�H���VD�>Do6�8�H�h@ "�Ȏ<!ń�A�n#ړM��!!J%PH)�;<x|�f�J�+�F@;���?&���O�Af.D���C�p��c
A�g?�5�>|�z�#☗rH1jQ�i�$0Q�3�ɦ)u$1 U���}��x�%��V�.�C�� �Fϖ}@���H�(r�f�I��<,tlؕL̴�#�OX�ڴ#�t��hCb�,��C�'m v+��8,͉�Eɕv�ny���! 7���Ǌ��xޔ]kK<Q��Y�<)���=�~r`��F��k�'r��4��c��~rHM!xY����A�^��	9�J@���4�:�7&��2��C�Oֶ�	�E2>�NO,m�
ЛD<Н��@:�{�p�d-4�p��3��6�teH��VBA�
֝9k��<�ƽy��iAG漫n�';}� Y�$!�9Yp(T�
��y�I>Yr,\H�OK��I�������&��a#\!a�.,:�yb+L!.-8` �*�`@�`�И'�v	�f��&�L!�� -Εp�4!���ێ}2C�gl��ja�-h��i�t���';�MH��IC��(à��}Y�P�rظT,�52�g�Lz ۓmU��p7G�7J�	Ӗ@��?�t�JrF��pp�@��@B��;��G�sR��'��hI����<k4٩��%qaj0ZT#E��yb��'jgX�B�A�&����rE�%,6�|�r�E	$���!�+��'��#�k�\��w&�y�Vhγp�L����а5X�q��7���c�
�B5(�V"oX9��a�~��c�8��i�'>��*P�B hd"��%扶o�acA�� ��L3w��"'`,�>�B�
Rl�B� �3�,p΂�/��T���	,�v�V�(���ӧO(:����a�^p`�V�,LO�"׭��F3D�1Ea���;�']�9+�K?�v�*ufK�sM� ӭ���D�3A��_7Uj ���)��X���@���-d!��C�8�A�)#z��ʣe���na2@��:T�P�r"�ά8R1OP�p&�ތx�&yx�4�):��[+����X� �P��'�D��"��,�@���X�\�:�٤'�X�x��<٠/�5Ux��tT�j͎t�q��̓>ER-2��>A�|�wfA5U⼄D|үY�A�vԙ#�̵/{�-��B��P���Xd	��TҒ1�࣋{y�i;!jݕt�XI!%	#I��鳓/���?I�������x��) ��9�>hI$��s}���b� Vxx��'瓶2�@9��O��C�|̓�޹j�mY�/@@�ɖ��G��q���fX�T�?E���D5�H���@Q�2rHIVC�A�NUAE��)��)��i>咖���e�杞dG<{���.O1���C-Q|���[;<�B���� H����c��d���T�'�hi
�*6�'44�p��Dh�j-K�$"<�AS>�DU�8�h��Cl(�zT�a�?�T����D�Q�C��8LЎ���-҈��i� X����hD�0�GefI!��!L$����9`����̧^�� �L�0�L��V�{H�}��?��?�����Q��=`�g�n̪��DdD��@ 6ҼD��@y���1��� Ԕ}KR�{�� �7_i���<@b@L��)� �,I�dC&w�v�a�A��,�5@D�ɴe��m����0鑗��F�M�����6�U���csÂ�ÈB䉲F��ɰ��Y#L�0X`D��z�d��-vL`@��R�(�)#KI�)rd�}Zt�R�t�0t�g��Y�$I�v��}�<9���|Zd ����r�lX��ώ�1ʣM����H��		���fhSp�n��D��J���T�C.J�"��-�.Ȉ���v�h�H�D�O�f��6ᒬH��9c��Fi��t�e�5S�rlZ�/_4f2�ʀ� �\����6犉#�6�ۓ':s�Td��:X��]cTe���	�)d~��"O�aL;8�:ɘs�ўD6F8�`�i���b۠��s�/��Q�(�Af�(�k�\�����	lD�x�"��N!�5B�DEI�mҶTO��K��Li�
X!pGD��lI�,��4Ε�BT?��2�d;����G��҈Z���(�z��קt"0���Yl�Z�,N�tP��̊Z��#�.C�u��P��L^'%�έ�ߓF�q�ś0�^��
L�8���<��\�?��ݹe�
�}pP�7�P��O����J�/P�9sU��]@8XS�'6�d��%c�\p�uc��S�si�6�X0R���ȈL�����)�<���ǡ�)\T9��l�<3��4�s"O��6GU8[;@��t�3 � )�PG�9m{D��1ݙW�8T�L���2OE��㟼���S���qT�J�3���C�*LO�9�u-ù�⍣D�M�g]\�)#ɦmm�����[#n�+�����M�R.�<:7���ɺr�Hag��j[^�#%�b��+\��X%�ݠT��)���,.�p�� ȸ�u���=\tw��6!D�124%�+�y��G��X�%� [L������P�r�M_�5�I�͔�n�,�B�C䒟<�Z�w[�`6F��
�x�)a� �1��'?�dB�/�+�Bt��˛�/��"pI7�9�!%���͘%���<���Ѝ\A���ԓWo9�$�@��$!��ͫg�N1�'���	��W%+@Z ��������'f2 ����K>:���#ɂ9z���y�/Ѳx����a*@�OU�(�̈́_J˖C,���A�'t4�&��}��7M	/ Z�� PM^1���O4���3?i��]�J9.$Ar,؏d�� 0��v�<ၤ9f������ʀ̊�Ѧ~��� �`A�i>.���I�j��g���)�KX(eF�ի�n>&�P,� C���Z/�!���:"�����6B�5H�`�!�ս!�^=B�Ɣ3 Kb�<A�ʍD��Y���0v�E�	�.m��C�0B�B�	�,'1I#��.Ű�cr�EI�8����	�Tr�fR�PG��OPK`gԷG8�����E�,)�5�Q"O,䊒F��
o���+R�\+T�[Q�Z�H�t٩��U�p>ѳ������V����#C�j���k'�0.�~��vS����l�3jv�d�>W�!�S"O,ݳv�D���<0U!M!2�av�$U6A�bp�����&��a�B9Otҥ2���?R	��"O6Ti����v��'�
�s�:<(�g[�&�h%�<+��<�R�Άv�X\ '�O(P_�1�TFe�<�hQ�T�� ��K�!SU�5���i�<qp搼�yq�@�
%��w(Bi�<)B&[OP��O��$^<B�J�I�<)�N�S� "Ąu
(3e�z�<aeI�4��q�E߂=�0��*�o�<�5�ώ	�VM3�CQ�6)PX�g�\i�<��(P����B�:a��jš P�<�6*J�t@<��%�H�0�atv�<ٖ@!�29����1T���c	o�<�$�Y�9���c�,1%�q���`�<��#cI�1)�D�'=�r���)XY�<��Γ$�n��ώ�4���K&�S`�<ar�P��vd�� [�
�� 4�B�<	�M� kO��(��H�
�svc�@�<ѣ�P($�b��"aғD ���{�<9E�̑
�px�-Г6`�	!�,T^�<9��s~�/Y�:!��̈́��B䉝V����Ч)>�l��H�a��B�)� ��#`���Q��9�� @/%輪W"OF�S!@�FnJ�f�Ɔl��"O����e-�K�'�]��"Ob�2A�Y�]6z�
h��S���t"O����G^�C�,�tǍ wXR��`"O�@zj
j���¤8C�T��"O��Ұٟ2�Ƚ��C�;=�"O��!C�Wm6aR3C[<= ����"OdQ��-�'���qL��7/b�b�"O��Ђ�]�6,���E��bs
�J�"O�H����hQ2(Sԅ�䖪)�f"O�zҌԉ'����+-v�6��D"OB�S�$@�nH4��+�Z[��;#"O�����;n\%jĈQ�uf���"O`�D� ��ɣ�0K~|��`"O�R��09zBe8�G�S�*xj�"O���O&}�%�FeX()R���"O�����>T? ք�,
�v\�t"O��A��6��a"%�$����"OR�c�Se�,I��T�V�ll��"Oxp�kQ?^��Pp]}ڼ�y�"Or ;��U�e�%�߬|�\tP�"O"D0��eP��2��YƠ�S"Oݳe����<��o���z���"O�QC����
�x���D$f{�!�t"O|�5&��\W�!p#d��;��Ua"O��[�#n�~����:��lCe"O�P�J�d��P�R�_�\ �"O*�xX���*R<y&~ �"O�����W�쩃�hD�m>
��"O4�p�P2>]��3�}��I�"OR�!�lY�$۬�6��:�� �"O��񅫎�6~�i�!�D�6>q@B"OF��ń]�J���ɤ�J�&�܅��"O�hA���r_*��@ Px�� F"ORD�G/�<P>��� hZɛ�"OXHy� дHaO�4F�h�"O<�p %�$%ʹȑ�d\F�-��"O 偅���D�95��-�Up�'�!9�Q�W��!V�e�\x�'��\+��V�\І�VY	0���'7�5��FZ`�_.Tj|@
�'Q����e=3�H{PN�\�C
�'1L��5��r~�H`FB�[�����'N]P$た\�
0Ii�P��b�'��Ñ�F2|1gН1<�|�+O6���J�!�:�`��<dKUꛐR�!�A_��Ԉ�.�.������6,�!�$]�ty88��N;|����ʧ�!�d�4wYhIaD[7?>����3�!���L�d��4�C( �H�ek�]�!�dB�M� �
S<�Ы�* !���I��	�J��)+�(p�I�F=!��<R��u� H�l�=(3h�J!����q�6+#m�� ؠ䙏x!�$F"*�D�b����N�\i���Y2�!��bI8�IeL��N�l�Z�� �!��9��@0C)F�:� o�!�$��:�@�P"�_~5" ���O�!򤑂J�b��&+	�q�nP��Щ�!��R���!e�c�88JdGQ!M!���G@^M������(�H�*g�!�DD�E"��	�nzLtP�(�Y'!�D�P��5��ŉ�bg�Ⱥ��L!�� 0�ui�"z !��Ε�{>EI�"O�P�0���;3&H3V��.xul���"O�Ds��M�4�Z٨�N��ogT|��"OȘ��.H��|���,Ua:���"OLy����k01�`���DU�q��"O,-��"F<c��܈�d�>'�J�R"O����
)�1�c-R�9� H�@"O�]�k��i�~�ƍ��W�����"O�XQ���������R����"O8����J8t��
X�xz��D"O`��bO	S�t@U'"rfV�R"O��S�aL� 2�E�.xF�e�"O0`�Ǐ�.q]�rC
SH`=B�"O�\#0 ��:�*����E�>4���L���X�ue��jp&#��H����!�!�䗱8ɪ�c�.\p���1 	9!�$
�B&9���N�R�� �0e)!��;N=}���8@n2%R��O5U!�$O@y���(Z-_�arUa�8^��φ �|��ߩ~S�K��1�B��>ctY�흊4��M��"ȩ'Y�B䉒_>�[��P5%���@s(�q	�B�	%Q���F��	H�-��%-/�B䉣P��LEa��Kל%sՊ�q+dB�3;V�S4&��*LA$��PaC�ɳ$R��? �н�V�R�	��B�&P,K`�ťM(�!kŔ�x�B�	�c%`b%�=`z��rER�Qk�B�I�D�b0�@�T�2tȲ�L�{��B�	�
��xQ�l��"�
��J���HB�I5h�n����2r�AZ��_,r�C�ɻ�B��w��>,K�qQA�&�B�	�#���q�Ħo!���v�T6	�fB�4i��}0e�N7/�NI2��p1C�IMF� t/�W@:��4��,�B䉒(���C@ͨj��0z�_5w<>C�	�j���0~�Ĩ���mp�C�i�j"�C�B���a����"Ї�O�&�3Ɗ;}�@���"�'}�ȓ�LBT�ڽ\��c�(��(fLB�ɏ<��U"�o��{���b!Ϗ�!-lB�I9GN̬8td]�h�	é41��B䉨�f���Y�+�1q@�B$GT�=�
Ó&�m��nПK̸t
�ʌ�vR0�ȓE_p��4�d	�*%�C�	�g� �r+��n��T��nl��8�I ep���ԽbW����#7��B�d��b�K�"m���P-7`.B䉲����w�ɝ>��"�� �Pa���E{J?�C�m�w��*4�]���%3��&D�8���G�mʠ�'�6y�)Q�M%D�,h���(��E@pJ׌:1~MV�&D�@�U* ������2!�09�+�>.O"�=%>�bc%���)I�酴J�8��Ĥ �O��|�,e��[�m���H��L l4��9oT5�W�1c��Z�U"u4݅�2���tI�q-�8(ק��( 9�ȓF���{��+���i_�h��чȓ�x-AAH��YK���.U�s�z-��U}֘)"��?@��Af��%y����H� 	 �,�-9}L�k&*��	F8��s������a��\s �./
���	I��!0�
={��58 !��X�C�ɺ$Ӣ�r�D�|Ҭ<��n��!�� �l��K!uG�T(�+эZ�l-��"O�j扂�qZ���L�_�2�K'"Oh�a�ʨpP�)�K��_Z1yf"O �p���%b`�,0*R��ku"O�@��ŕW�laz�!�0(ЈC"O֌��ѓ^퀍K�Fղ"� �"O��Xq�# w���ħ�Ȕh"O�)!�.��0��`PC#�� �"O�`��h�J@��
#-��w�L���"OV,�v���|1�L��&!a6"O�1`"���Mf�H P,��9���۰"O�0K�N�9`�v����!p�X�x�"O
�)�`�Ahi@lB>5��S"Oz�p&9��tJ%�YS���X"OL1���/ I�%Y��Y�B���"O�A�g�m0<���dt�|��"O��* MЂ�>�!@� 9쥢�"O�hXS�D1rO���S��a�x�b"O�
P؛��c#��T����"O��٠�"̬Y����R�F��'_^���`;&Uh�L �xҪ��
�'�����ϗ5��� ��2~�p��
�'�0��e@ MP-����tj��	�'��ɹ�A#�`���h9����':�%*�!�g.�:�@�6�q�O����T����j�	q����C��h!�3�TE#'LH4	���a�;ng!��_�/|���.ې<��]�&��:0!�Dӡp}[a��NHtay��L4K!�T=LMYԏ��<H�	kE�O�!�^�0�8e#K,N<�M2d���!�$�:�����k�H�0�07�B�K�!�d�<됉p0I4���R��ĸ��yR�]� ��r�C�}��%��ğl�<�v �	��ɐ��?.��a)�H�`�<)�C]M6�Z0'�$Jy�Q���N_�<��!l��V샫c���0Q)_Z�<��ș#T��q�b�}`b��]U�<!W�t�ZAAg��&e��|ȅ��V�<�%�\�m�"M�@�K�g^���'�U�<qs��#k��#(G�W�&5b��]�<�RK��"�^A�QB�n�V$jD�[�<�5��q�X��5���?�X��M�<F�J�!4 �G�H St0a�GEH�<Q� 7��@�wc��T��Q o�@�<�7�$���ǙQ����a@�hF�C䉸K�����W�>�v(R�S��y��+&���M(l��(�y���K3�(���J�XI��c�.�y���������$�=R�4��	=�y� �0#�
�as�ة����T��y�K[�YL�"�<L�谦)Y�y��b��ܪ����U0F���y�gZ&�=�惚�D���c/�y&�-j��z��z�L8!��В�yR�аh�Z�������^2�y"��LR��ǎ��<���c�V��y.�9Q�7K�:.�^�[F�ҹ�y2�������a���"�Ҹ��G��y"�Ľ&�H��$lC��zE2aHS�y�f��/H�`���M�ژ ġ.�y�I�/FZ �w�N$\ږ%Rd"�y�	�l��S��_f�֌C�y�L\��"���WZ*�+�$N/�y
� rPaա�=X���z�
?�Ҁ"�"Oҭ�4,ƞ8����C�l�.�"O(-��Z�l��+6��G+�XiC"O�h#��~�:V�S�<x�`�"O�Y�qmQ�,=B@�IY�fe|U�"O��!@+�2.�)�I�ad�{u"OP�(g�]!P1`u*C@&<8=Ȕ"OT� !��S�p� s"ȵNr�("Ob��+ۋ&٨E��+�$]騬��"O| ��BCw��@�N2	����"O��Qi�)�h;���y;>���"OΩX�P�;�8R�M0�U��"O�u�BQ7a�u�K"U�*b"O��B�[��}�R �-Z Z�"Ovu)�K��E�j@a�m!(l�у"O&��f"��L�LH�ČNx��"�"OL���,� Z]<�1�lG�E�5"O|1�ۆv��R�$����"O��&c�>%��s�_�p�(F"O`H8�ʖ]j1��D^�J�� "Oz-h���u�ISf�IR����"O���f�+[6�x��n���9C�"O�B��E8^��<x��r"OLH	�DN/R�&��ӂ�G��@�"OT1h��"�0) �݅�^�x"O�TRp��j�3�I��2iCs"O��+gh^8���f� k���s�"Ob	(��Ce�\I��\/ v �"OU�CN�W�^� ��/v��}�@"O��dhS�4?��h��F<�|��"O\���Zt`,rWв;�F��"O,�a�g��D�����p�dc�"OT��ǚ1&7��p �Ńtq��"O.�#��+�6��"�9{s��"ObH#`��!��x�!�ƢD�6 ��"OPb�
"9��p�������"O����i%��!��hԣ ���R"O|Ջj�0�aG˓~ �Z�"O�,��j	!Hx� �E�!{��\٧"O~��� ��0=�P��	)p���s"O.9�W��?�H��Ղбi U�$"O�db���+S��Yu�ȋa��Q�"O�L��GZ�O���R���MG�`��"OJ�v�U�!����#"K�U�j�"O���V��;1�[B"�2TLݚc"O ��$��8��|k4�$0J�y{�"O���Ԭ̋4v|P����uF�5P"O�Q�FM�5
h�m$!9���"OTY�:3r�#�
�k�D�0f"Oج�f��;��Q�Z	G�lq0"O*Q�rdW�dT*��@w���"O
��!�[���䆗*,j���"O���j�l��I5#�6U^\��"O�d�W�[�k��H1p���X|� Cg"O����g��B�0`ӏQOez���"O�h�$bJ8`��y ���-^�4b"O$���l&`��l]�Ma��{D"O���ŀi��tx6ldS`���"O���� UC	~j5��;4��R'"OZ�K!J	y_�dQ�I�T��I[v"OpĚɋ=^�j��%���~����"O@�"�Z��lr͜�c��%[�"O� 3��ޒ\`�E� l^]��9p�"OE� ��5X !�Qʒ�6�z�R@"O� T]�a�k�^-��&\�8���V"O�X�h�$S朒5�?�\��"OL�[ǀ7in��ac�Oh�k�"OtT��˝�|o|��U�U� ��"O:���Pr�&B�X�&��v"OZ�XΒ�?f�*�+s����"Ol�{eρ�)˺�sF�ϔS�2!��"O���Z�p�d�؁oWX�>x��"Opi�F#�|�\x�dP�F�T�s�"O|(JdaV+Y��0��)g||��"O�Y�R��JUp']�4ZZ|K�"O`:We@�b�ec�-d3r�u"O|�j�W�QR(]�R�f0YP�"O.���c�;Ld�9�d�O�]���"O�`�̿^I��hD-�p��Ȋ�"O� �W�5a�"}c�*ۭ�*$�v"O$b@�ڨb[��q���U����t"OP$�c&O</X1�'W�${�d#�"O\��t!W� ߄)i5,�4&מ��G"O �#J�we�����
�#$=z�"Ob�����3t�|Bi��@��D �"O�x��\0"e���+���"O�|J���$zҔћҡF<i<D"Od$�7 ʴE�rx�^pR2l"Oz��΄F�]zv/�@���� "O�D{0�87[>8CT���p�0��"O� ���ߢzN��P�W1P��"O�P3�Ο>oB)�E�ʺ@�@<P"O�0fh�5�JC��P��>�b"OTeK�Z���)����jt`�"O]��ݒ�fr�-ɪM�Y��"O���a��?�6�X�L�J�>��s"Ovmh�OC�SV��U�Z�A��%�y�լ9�±��hģN�X�Q�߬�y�\�+΅�C(N�|�n2e��'��i�r��%�<��O�#Y"j��
�'���9���+x�@D#�*@��Ѩ�'���ݓeS���Z?+Hԉ�'i�U�c�ܢZ���
�h�;\,���'���VE	�S���E`��8O� @�'�*h��� 6�����5*^ѐ�'f�M"��������w/M�XR��i�'3,���-�2~
LhDŐ]I���'���BQ�����H.QY���I�'0�e��I!y L�S�\�O��'H��V
ގ���@Ǟ�u�0���'ݠXC�$O;:5Ps!ȋ�8��e��' �����UʆdS4fЫY�|(9�'|���b�Ows�,��Y�M���q
�'�R�BE	�)�TJ!L��m�1S
�'0�Cc�%Q�ع@)V��M �'������G��ቀ/O�NYX���'$~y����k8�s��A��ih�'�d����r�hx��3>�}��'�FTCd�/ZV�jG�M(-n���'�<`J���i�>xA+�*z
�!�'<LQ���?{:�Ѩ����$wL��'����%�/�0�
�H!�hm��'�:h��L6\���ɡ�Q�?��� �'����ٶ71�b��<�T�
�'�B*�@aX���7� ��
�'o
p�E(��|�5OT8'���	�'K� #4NL $�l|���-�F]��'n� A�Ӊd��ݛ�%?_�l����� 𙡂�0��Da��R�r@q�"O��;�䇁��� �#���vDk6"O�t���g�@ �ԃ�!��a�e"O�`#E�$̙3���;���"OLa��Ie��� � �3k�4�ٴ"O.���^�MJKQ:j�XbE�4�yλ��#�� ]���)��� �y����m�G�D�N���%�؊�y��,O�t�bg	�L���,�2�y���g1�0	�ȑ�7���1CM�;�y§�=|���SJ�3{O��ӣOſ�y���T�d�U���W�i�ᐲ�y"��p�TX���%q-�)kfZ/�yQ%Vv8�1��N�dZ|a;����y"�%_ ��R��k����vfF��y�,�$��VJj.� V�Y�y���2bz�VgH\�)UFץ�y�� �q���`��hBDoŷ�y��_�u,F�@��G�Y/���
1�y�lU�2����0U$Ԁ�	��y"�;wq�����S8E�`�9�G�-�y�_
2�ր��댁l�D��!���hO\��3Q��@���8����F:џ�F���0R\Z����R��� �����hOq�ܘs�b��S#�d��[F �j�"Ola�W*|�=HE��)g�6I��"O.P&K�-�$��Ą˙s�j���"O�Ġ�m!�^��EiOYpTi�"Ot�@C�7U�:U[(�ak�y�U�'��Ⱥ����[nx��Ve	�ܬ��p�)D�x"@���6@+㣈�)u�б�-D��0�b�NdNi�Ҫ�'��xk�)ړ�0<!J���d�������!z�R�<1P �;*:���E L���qd�P�<��LȊV�����l8�9��P�<d��i����UM�I�fe�t�I�<�-8tC.0Q0Bԁ+����G�<1 �K�j��9A���;sL�+�j�p�'�ax��.OoD��Ƀ$o�8!:�#����<���G�>R��� ��6��0�ΚZ!����V0xbK�8� -�v����!��$:AD�� �h:�k�"�!m!�䗴v ��jSoB�s��!��X�Z��'�ў�>��1pw�x�H\9`��@�Q#9��7�SܧhL ��ԧ�l56ZF���g�H#��͟d��5Q�ϛ%��=E{��OȂy� �;e32�ڞ��y0M>�,c��`�Ӎ-��-�gO�V~Іȓ`X��'6��}���"?~!�ȓF�r��%�"jO� S��ڟj�
D��S��xĸP,��6��D2�k����C��$��y��;j�B�j����x��C�I#n���Y����|v̈1����?����) ?��+b[�KED���I�<����;��Y�4�{r�mS��K�<Y`O��X `�YЦ$SPnũQ�F�<�2��{KNA����0I  �m�~�<OխC�*���[�K׀�#3��}�<��UvF��$�^ AmH;C��A��0=A`� �JlB�9# _�O/���U�V{�<��q��x�l�9jv��P��z�����O0�$��N���
�nU�����'���S�%�g�p���<�(��' RYl��;<��B�Ԟ.k�%���� <��b׎ }(�(�Ý�F��q�S������|�&��CO��P+|��"A�-6�C�IN)&��P��6"��5�t�O��x����x�'�d�D��l�Q�S+�x ���x�
��z�u �R9 5r"F
�y��Ăr��9�M��*����'���y��]�wRIaf!�r�0DF2�y�i-�`jDjq�e�R��y�ƅ;Y�|������ 3��8��'Gaz� 	y��%���4 ��KAn��y�A�� :�&Ʈ) y��!9�y$�"���5���'Bz�#P썋�y2m@�B*J�C�3{x��4��yr-C T�Xӱ�Ψ�����y�g��)����e�_>o�0pbC���y�J:�0�3��LQ����T����0>1nR38���ѣݥ?N��R-]d�Ik�'����<aD��Isuj�!A8���[a�<�V��v������on`AkA�x�<�T�1|�
8�T�:K�R\�C��?J\�YB$��Q����E՟B]�C����b3C�:Dp�eC��Q� �C��/pu���!��*�q�^1Tn૎"�)��lN֎�"���#WX^B&�Y��y򏀰<�j�S�lQ#Kn<U���D0�y⏇=}�
����Ќ>� �����%�y�E��ZĴ�#me� ��װ�y���eH��t �"U}��hQ*���hOr���@+[���kakŭ(��TK�
��x~!�U,v���%	/+��hC�nF�)�!��I#�J����@����#��2O{!�DǕp	�£K�El�}�`�MI!��kH����٘Kh��Ӕ�Z!a�!�ċ'@�<}R$J3�,������!��_z��Tb�
|8�:3*���!��W�b����I�p|-Q�
��!��\C,�|yvN�U���cB�7��O����xg*Uh��:E���O�${!�đa[J�;��@�%#TJ���S!��@6��tI.��[p|:��"C�!�64�jL[��I�h�1ɖ�!���)�`Pg�_�"9H�'O�!��5I��x���v�8�c��r�'Vў�>��>Y�a��6UʚT�§8�$*�S�'�Ƒ��L��^A �Θ�o �t��	b~R�.���.��җ\ @�J��
�'��#G�� p��f0��	�'k��ImQ�=�aS��D�2<��x	�'E���/Xǂ,s��#�����'�`�0����У H#ZBQ�I>������1?v�k� K�vXF@Ƃ��+2!�G+x��z���
{AȘ�C A�,!�D�!z$�5�ƤKV���<L�!�J!�����%��DK���A�
|q!��U`�d��@j�?\B�P���!�Đ7v^T�WJ՘!Br�h�/G�!�I�Qi�焦j�lhq歁$.!����4@���V��)YWBƍ<!��L��1��Ց:{䍑�Ւh�!�C�0���t/X�Wu ��Y�!�DĚN���nmb�SO	�!�$	�gy���g��`�`���z!��Ta $��OE�p�N�BUI@��!�$Q�e�p1�g�����a�`)ȣXo!�� "�ʎM`h��lDj��@�"O��Y�LN90#Z(Ɂ,�)���Is"OZ����IUR�È�;?�d �b"O��Z�fQ�3�j�����k����B"O�
6���1����0�W8�T�p�"O\��3C/w�dʄ-·v�>�1�"O����.��P��A��'��'��6B׆��􆛜_��@�ȪB�!�Ĉ�G]�rdB�
����흄*�!��)g��I��D�������&�.�!�� �)f`�i�m�>w��mC�LO�!�G3� L�g��J����i�N�!�K2F���-�0�Rq�o��T�'�a|�E�'�<���'X92 �j�P��?�(OL���P� ��`i�iA�X
��6d�o!򄘔V3��hs���y
F��6B��3|!��D_�\J��Fz^�����Mx!�d��Y��u�vJJ�
����!��SPnm�En�0��-�6P:�!��j�$D����6�r R�횎b�џ�F��M��2��p-�<O��v�B:�y"��>��ip�+��E$4k%@՘�y'ԹBo���g��<�P�)�
ŷ�yB-Ln�R�C��A-k��TnK��y2#����!c(  ��<�'
��y"f�2-|����$�Pˆo���y�e���҉�1�Ѽ"�As����y�	ՇjR��#�#=�ƍ��ɨ��<���D4�\@���#�V�X��ǚ*F!�DV*L��0��RF�0S��,[+�y��	� JmX�&�WHf��*]*"B�I4�e�����iX(H���+'B�C��6q��qm�c����va~C��1R@��A�����p��OE��h�=��'���eZ�u|�[��Zܰ�ȓYa�S��>�h�c�FIa�Zȅȓt�>9su�B�m���5� �r�4���鶨��F�A]]��,��F��ȓ_ЮL��	\t0ؖ��'𮹆ȓc�l��3,����[@�A�Ky�!�ȓ7=��IE	j���EdF�%�0}�ȓ��-�rd�(�X��s��=�DX�ȓ���h�G����cs�<i�x����T�f�F�T�����6<N��d&^���#�����*s����ȓaP���2��9���7����qզt���c �#6NM�Q`v���$����m��镎�3����ȓT%��`�8r2s��W��%$��G{���M�v"8�;�\�>-��b�X�y���V���<x��T���y"F�T��z�㌮~�t	�$�E��y�&S�#( ���B���tɇ)�y�j]���
��;����AG(j�)��#%|LR#�϶5n��&K��j�|��ȓ!������Ի)�: ��q,XY�<�ǌ�0���@P��y�ҋ�T�<1��S�F ^�䁛�FsМ3b��w�<���߄mP��1�.F������p�I}���Oܚ���ɗ?��´�:�pQ
�'<z���Ƃ�Ϯ�Aw�^���$�
�'��5R��8.+���(� �ک�	�'|` ҖGр�,֯.�d�I>y�z^�I�V žDz��RfEI:l�p���S�? ���
 9�FPk��l3����"O�������#]t=�w�]"D!}��"O��&֞�(���Μ6n�ű�"O��Ђ���v��(����c\D�""O�Qc
$T^|X)w ��E�x���"O& Z�/߹')SRA�"6T�p�"OU��+L�oB�(���Q��"O�ɓ�%��(���!�0|����G�'����ʱ�iY�}����Y7T\B�ɵG�J�(���4����[	2B��7
�`��E�$O�q�%n�����0?��Iו6�z�pUbY1|�:�*����<a@KZ!�&���
.O�Z��v��~�<�Uo��B�(t�"��	��[cN�}�<"'V3{Ĕ�J�/=M�Лg�a�<�5�& ��l:�l͹}�l����`�<��Ŗ��!��H=�2��І�R�<9G[0)���ql�UmyfKAP�<�Ч��@r���	�B@��NZK�<!�@���䀐��	Yj�@D%�]�<!G�	y'���BgQ:�F!�*�n�<QBF,�.�el����C &�l�<AA*�,�j�`�/c�l�K2�l�<�aF#����G�"{�.���͈k�<a���@��"6���+�0����j�<��ܤ[P�J@����D��e�<�#L��M�����DЬ7�� ���`�<�BE!l���#Q�Lޒ����Y�<a���3h��c�G�-Z郔'�Y�<y��3M�!�c� OA����U�<���*��p���oV���N�<��˝9_C�ة�X�nI�y9%�M�<i�@�s�^�I�*��9$�MG�<�o[�r�,�@d�d�T@Q�Hn�<9�.��E���i0 Ô~V}	$�Rm�<��F]�S��H�sĜ;E ��*&̚k��hO�':�!J���;l��g�eI�ȓ�M`Ʀ�)�(@T��!�r	��K��|��k�h�I��Ɇ�D ؠ�ȓDI�E�J�ʅJ
��!��|�<�V�ι\�p���7�ؔYâv�<�w#�;Jz1��.4ROd�I�]r�<�+ۊ`"�=化�Rg�:3I�F�<I0b�8.�1!���N�����E�<���Ő՘��D���:p��DC�	�F��-b��ڢ,v�UkEOW�(L�B䉘?������i<����V;,e*C��	h�P�7��D~UkQđ�N@ C�'��哳���/*�T8���2:w���d$?��-^�	E�l��}��	���t�<�K�
vŎ�cal@���Pƨq�<�&��?>w�t�삁W��`�)o�<���M�w�l��Ũ(?�J֮]A�<��K�z���xg" 9JV� R�<a���v�He�!
9ȼi⧛K�<1؛x���᪛!X��a���k�<�m���(	 ���!�Fi�<) �¿�\���--�xi��Ky�<��0pkH	�*D���bNL@�<iEK�� 6<8��R#p��J�I�d�<�R�P�V�~�4�� 8_��R-a�<)ck�X}h(�6�0��X
VT�<��a20�mb��:�
�.�S�<90�3eD���U5t�����Ux�`Fx
� �)�W�ϓ{?D��`�݅)ٸHW"Oj���L6_&� WC��*�vtI"Obe���y�� ����q��jC"O�Y����Аj�D~�t���.�S�)�b�6{�Ԯ8���G[�{=!��-v'��i�� ���1%��5O!�dߟH�
�A����[fEL2!�$� �$0�ƃ�:�t��d�!��Ob�=���ukƢڨQ�>Ts"��4_\V<�"O,=k-�T��d!	A�W�!k3"O��C�B��E�g�;@�~���"O�����H����MJ�"�SC"O�)%���W��|�7FE#��RD"O��D��[��� ���k��@�F�z>)��`R�r�
P�r�_�i'����Ĺ<�+O ��7�&�J�bOC L@a��p�8��"O`1ƃJ�E��x°�U�<n�b"OJ���DD$���&�/Hk�,��"O����
��\�-����f��KG"OBI
�7v �M�񯙿
c�mb�"OTP%��
�����JK�h1"O� qwjİ&r�Vj_��
�����Oأ=�'X�x�0ԉʌb��Ԛ%H�6d�L��Pa~U��J�?��zχ2M���ȓ%��e��'��Y��P�߮3f8؆�?�\��bʄhGN'G�D�ȓ\~��$$:�y�Q�D>\`�ȓu�@P�"h	�{���3�J���l�ȓ�T�a�׏S�TY�んu. �ȓ��M+3 �-/��MC�ꀕ;���ȓ/�2��������sEm�i�✄ȓM�e�T朅1D,AS �%v����ȓ4�4�����0q�+��!=X�لȓՂW\�!��=�� �<O�x�P"OLa@ ������`ƅS? D��"O$�@�HZ�0+��-(��"O�qb�/$�vD�&����D8�"OX��U	��E�.���
�����"O&�KtC��u��(q���z>��E"O`�{�����ʅk��g�P�"O1��M�c�N����7-hL<�'"O)@r%LY��p2 'ϖM]���q"Ov���C��O�D�[��P+LS�dI2"O�|�!� ]s��y"*�%�>��"OJ�Y�S~�X�`@#G]��0��'��	�6�����Q+bp�$L�4C�	:�v�bi[�W������FdC�I4_��@����)hX��.O�DB�	1#_�ѩ����J� �B?H�8B��*.��eR�b�r����f��(�"B�	+Xk q���ڷo!�B�ɚ}o`ȊW��(�İ�$�\RivB�	A<z����	 '��d,��O�C�	O�8����՛D[�FF�`��C���%���{%�8�|��"O��O��a@FXaB�P��p= �"O:�r�Г:8�z�M�;��ʲ"OL���k���Z���S�;�HH t"O`�cb,U{JQ1��h~@QQ�"O�� 4ĝ[�q�L�k��c"O�mj�̕
N�ՠ�JH�,�J�Jd"O6��s�]�|�:��ށ�tt`�"O�@�TH�02�IuGK�N�z�"OT@hb!�4'��M*�-�Qj�H�"O�  �r@�P=�|��5Ɯ�S{��a�"OH��古P�,�4@]�A�da"O>�HD�c�u��Wx����"O�iX&@��	�غ%,C�Bd�'"O��(�Œ.�@����1+���Z�"O`P闇 ��/�/�TY�"O��X���E��̈:�.Q�"Oȵ�0C�7�6AF��l.��(C"O��!g(�M�6��!h��H�1"O8QѓҒy�L ���Һe�Җ0�y�ŝ�b�B82gb�	@hZ������y2�I�o��EI�ď.Mdc���y�%Od�}Ycˈ%��DQ0���y"E��5�0=hu#�O	�tSd$���y�۴>w�M�F�E�vh�S.״�y��?w'�4:�i��:��8��)^�yB�,{�`	�$̎�1��$��f��yRG�#��L��$�te�ä�����!�OL�H�%��T�Z�:�`G2pq^���"O����K:�$�QW�Ę`"%p1"OB���u��X:�-E�NL�$��"O~\h@�4F�t��FT� V5�"O"�@��%%T�Eo
�U��'|�cF�D�[ ��k�	�R����'5d``��uQ� ǂЌF��)�'v��JU����&Ը���'�R��
�' <��SF���(֫P�1B�
�'.��7�(O~T�ȥ��*+�L8)	�'���*pȉ�.��Aش`� p�h�	�'? [��,I�f��qX�� @	�'�l�эNL����AĠt���'�He��C@q�3Kքp�R���'�H�3�/�-,�}�[�lY�-y
�'�X�h� ø�����Nxr	p��y�@��<ҕ�C�=*���[aDI��?��'���F����,���Ƙ
L�0��'�Z����K�_~�XYQ���|Q0b�'S��)Y�?��e��,=�NA�'�p8�I14������*�T���'qx�Q�Um��H@�E��� u0�':���eV�Xࠨ�b	�(1��'(f�2��FĂ5zu��*R|f44"O�����;tV�z�HL�I��"OH��!IK0��	S�N0.<:�I�"O�(Y	ͭO\�3��G�rz���"O�|���ÆcZV<2�D%\�H���"O�y��@M?u�]�t�+}.�˂"O�2��R�"�X��vbI�s��Z�"O���5�������DBk��R���D6�O �;�Eu;B\�g��G��a�1"O��y�HW�dU�e�4%�����'�p�e*W*��B�D�V�9�'^~d���<�=�1FN�B�y�L�edPi�A�;�ވ:��P
�y�	T�M�
����N�:c���Q&�y��?��!�i��+��I"�4��'Jaz�(P�}� ��eω#�xs����y���Z�B�D�i��lZ�(G+�yr.�.p�v #W$װY�R�3c�O��y� Ҥ1��q�P�Ь(ب�r�c6�yB�S�efACǉ�P�l(����y���B��4Q�HH�H�ƭK��ݫ�yjkh�� ^u�x�0J�y�U;��%�2g��ӇF���y
� �U)��-wy���T����"O\
E�6*���I�*�>[e�U��"O�X!6LЁJ�&������{"Ov	�Fg~F����A;;�����"O"�[��?S����&I�]'��"O�hI�R����bfF�l� Bd"OP�C�\�&q�h�#U�z�Q"O�5z�/�0{f���fc�<-�ꍂ"Op�
�G% nd�#T85[��4"Or(��ʓ@� ,٠a@I����r"O����#�;Q��x�31-����S"O(��Aa�q��mT����o"O���#סK�^`�&cD9%�� $"O\�(wI�2J�xl���O�b�C"O��B"-u#J�
u�L�L���1W"OL�[�O9�lڒA�C��0��"O���.L1SنB ��y�D�Ä"O�E+���.n�T �a^��b@#"O���M��z$�����8q�D���"O�!�DL�}���R�-
�>���˦"O�@1VeE�7(j�����/;��"O>���l�Τ�����$<h7"OM�ӊ��25��:�U5��D��"OH	�rlF+g�x���?Qڌ��""O"p�Eꑍo�P%��aײX]d���"O�V���/�Ea��@X�B�"O��R㩋� � 8�).,-��5"O� �d��0r 1�Ph�$^$L�"O��p�I�&�v$�I��`��E��"O��*1�\�
���*y�z�cU"O��fF�i9�ybP���2����"O�����e�4�+�^����c�"O� 1�Ō
<�P��DUx��+"O��bV�DrB�1��)�9y҂ �"O�̪uk���I���&#f�dp"OL(��nS<j@+d'�4����"O2�93��o���p�����5;�"OnT �L�d���W#���W��_�<�HS�"�9<�E �-�S�<��=>҈4���܃DЮ9Xc'Q�<9�n�$w�$@�T�CV`3�^d�<YS�bj��1��.:��T��G_�<)��X+[�ro�)-����!�B�<���+�e{�ʋ#}�KUHOi�<�`�?30Kd�
�xt��(i�<yf�Q<`�ѧ�P(~7td��K�<g#�?b�H������ � �-�]x�8�'���"c��5�
1�`׳[�|��
�'ۮ��D�'L��r@M�6F1
��	�'s�p���Y75��h�į@�8z�z
�'M��D`�+c,�aHܧ4h
�'6R亳e0$����\t����';>�$S�Y��A��.<u�BP��'|<)�e'J5g�n�2�Q�j[b 

�'�*������֠��D���&��
�'��*�c����K���c%Д3
�'����g�,-�QfGA7' *
�'2�!pV<H��9���	v;	�'\�9k�A�6�.y{5�W&����'���A�?&�$49�ۚ���'�(��������;���'���	eU�f������-��"O��3F�V$dn�ȦCΫ\n�#q"OZx��'�z"�?\�@�"O� �x��S�Mt�R(��j��D2"O����Ι.w;Z	���(~V4�W"OB)r�gM}�FQY��S� VR�X�"Ob�xŇ��b�����D�Dd@*�O`�T��G�6A1U��,^�:�xT��OPB���&��PփRA��m^�C��4x2%RP_�'�����2�JC�IQO*xQ��:����d�~4ZB�I�k�(��o"$i�AӦ!��R�<B��&E�|pb��T�m�&a2A�+ �&B�ɋw����^� 
%�U�$-0B�I�~�RA�P��%Rl.��ՊJ��<�&�D{���+�����g�Z�1��,�C���yo�����j�"�p�3�Q)�y��?nb�hEc�#h���B�W��y�삽R�� &B�;a�~�9�bݘ�y���ff��W���*�x��T�1�y"!͔S� )�G6kE��Th���y�	 G�T0R��j^�i�5.��y�'�:m쨱�h�N�KD���y�J�Z��U��@����)3ɘ�y"Ϛ+B*,�bT���%�r,
��y"�X�q;������� ť�y��V�c~����Q1l�(BPKC��yU@�*y�1G�Z�x�����y���H�����d�e����5�y�l�(bX`9�'V4��('#�-�y��8B�0�K�R���B��y��3�0-����*\��	��y���gk�E����k��g<�y���2K��x�'ò�f� �AǼ�y���D?hqG�U\�,H��G2�yB�@�+9 �cd��a�تvBօ�y�WM�ޜɴ��_�xI!q���y��ŎI��˷h�?DCN�Y�j��y���S�t vd�$�b��+�y�����$-��~�#��^��y��͚��c�>	&�C"KW)�y��H� ���FQ�hR	0"�̉�y�j]�6J�x°�X6���y����y���1]�o�$�t� ��	#�y2��;^��}�Fď3<�6D����y��;�.9�e?.6huP0	�y�!	BnF6�0aEH����Yi�!��\h�=��l�[)�]�"�	b�!��>g�v�d/3.�Xa��&�'|!���e���x2���n�`�"�p!�Ǳņ��J�W���	v��Wb!���f��iЕ�N]S�b�a:wU!�D x��8jV� J�1c�`[�H!���7�F�;V�G=jE��)s��:�!�d�t���z����  n��F�W5�!�$A�\5�=�pƻN���m�js!򤁲0K�� !��c�#j�	=�!�����`��DM�N�Rw��	!��.�p�EY�z��8w*B�	�:E�9���"Df�� ��:L�B�	$@ P�I�<}�l)��1�C�I�b�0b#�+�8��A��F�C�>'Bi�a�@)%t|S�$'z!��D�F�BMCDS�	3�A�����&�!� s�\���(��1���®+�!�D�g��bV�!l �.��O:!��'6�J�hքS2*B�a��.H�!�� �d��.0w�\�{�Ù[$Hã"O��[�Nߝ2��`З�W�A$�'"Oe��.��K�"e��Ce� )�"O�p��ߔf~@$���֨K��}��"O�"�k�qRΥb���O����"O�!�1�X-N�ȡ�4k�(�"O�R�`ڪY��m�q�F%�"Oz�z_)n�KBb�H�r�+��t�<aPa�3r~j��1�3d}V��[�<	v�ɓ��e�%"�1�`I����<i3�����2fB�!��d��Jq�<�&@N�~sfQ�#� ~�J���/�C�<@�R�l�Sw땢U��9�uz�<�S\����ǝ���Ш_�<�"惲8D���h�p2\����Ea�<1sL\&J@�B`/D �!�/�s�<Q�֖dz$13'�'3����.Ll�<�+�4�4Pb�c҉cAE�#Ym�<iw-�2��͠3+[�`b�#2�~�<�d�;'D�D"܀W���Ox�<�� ���q��LQ| �"�MHt�<��@M�d"}� _y81�VCBo�<��G�{�N(AC� �D0���i�<���[��d]	n"tBE�l�<a��Zx�1!���w��l�eÆs�<Y� :R�ְbE�/c�Ƞ� �q�<I�C	��1 �%�?;�����DMo�<�A톽nh{T��#|���
�g�<	Q.�<b'�)�	�&TD�y��	d�<�UfL�A��	���C#��@U�<���Ӏ,3p0�A�ӥ#��հ4N�R�<97��f�:T�֋ӇG����f(�Q�<���|�<Qѡē�t}f�%�S�<IEɃ/9V�02b�0u:�z��R�<A�iD�НX��Q(K� �@CTE�<I�o�O���;�&P ㎜H#�w�<	d��@G:l���E�l�Cchv�<�#V�4&&�22�R"�"�"!��q�<!�(��%��\A��/m �)�b��l�<�t["6��њ �@)Z �]�4�\M�<I���Ӿ���K�	/�+C%�J�<�BMM:>�tA���"������]�<�W�#��j0�&^|r9Z`O�X�<9��Q"
�VD`Q��$G�F��o�L�<a���@��h�U���QP� F�<QVe�-���#�Q F:�P�A�<afk��,��:�AB�U�v鐵`�y�<)��ȍG߾�;Mɶ<U�]���q�<�� -	��R�F\��J`�U$Jq�<9\N���c����`ĂF��!�$�2c_Lx�$�����у*�!��Ro��	���+�-х���p�!�DG�F�(�dS�8	�}1�=�!���N�Mj��90��i ���!�D�sN^$yB�Z4Z~e#D�:�!��W�jp�"�(O���+��Z�>~!�$�;<�Bȥ.��"g豢T�N/A�!��?d��j C[�d�颴"�V�!��ϋ���r'�`F*t�c���!�=
.�1b98�ؘ����lu!�DO'p�� ��mߝF�E��Q�pg!�d��h%�Ԙ=a ���AO!��R�
������xARX)�/!��ث_:$9��a�;0X��ĕ�j!�� L5;�cW/|�C���>0�P"O0R���-aӦ)��e:�:"O��@T,��e�J	Xp&��d�RQڠ"O�����VÒ�S�n÷�"r$"O��� �����l��,�*�"O��ԥônL�A{�m�	f��H�"O��7�p �ݸ��_�Ph�:�"O�SF��bąH� ��[I��8�"O6�b$�:]� Y�͂�$2����"O85 ���%��h�`L_4_,���"O��	D��fHW�IjJ�)�*O.�I�k]���eO��)�'.�hǆ�7����
���B�'~��t"-?0��B�H$
2�Q�'2B�@1'��B�:���d$��
�'frY�v�G�$d�X$';Vg��A�'�68H��KK.���]�H���
�'��BǂӌP���Ίt�؅R
�'6(X�#��-T�a�#Ѵo���
�'��ՑtmOr��ˀ,Ѓ\��H
�'��tZ�h�R�Cp��"(
.<b	�'>0��d߅$Y�t;!�~t���'ͤ�Ӳ(����Yj#��͛�'�\<rEL�? Yk���@xd�'��azЎ^�d��,X"_�� �'Kp�A`�E�8��ɸĒ�
�'�0Y�d
G!������ݳo��k�'_ Ax�B��t� �&�Ǥ7/�m3�';H�����;W���o�_�9z�'|=���A�F�
�8�=�	�'�R-Jt�5�
ȹ��p@�:�'�^����6O���)�Z���'1��{���-�`�SR��!R!��'ᄄ
��Dmnv���dS�'h�8�'������% K�6d	2�0��'�!PA�Π;���,��r-~dY�'��y��&M�2!D�[ŧ�=v9����'h�x#7��(<�|h�΋#n2z�*	�'���rSN�'�������e ���'z��"���k���(��ʊd����'���Z�)܂V��<���6c�jA��'eB`��)�Z�|�r��֊�x�'䔽j�NR�M�z�3��/���y�'���hQ.Y@�Ӳ�͑,�8�'��@p�������+Y1V���i
�'��5�⬜S��5֍P:b	��'�P1�\l��[�,W�Eb��',��V�S�wM�LJ�bǝD��I��'�6��cZ�s"��NΥ<�q*�'����%a��psL%���G�=ޚAQ�'* ڇޣgz(p���B&3����'�݀�B]�:V\��4�@�0P�0�'�@`���6Y�&�"[f����'��$��K�c�Z�Y3��)T^�$C�'C�b��� >ڍ�bV?,����'�x��#��Q+��+b�&0�j���'լ��b�IS��x�Vi�#� $��'B�(\u�:@I��٪"�hi��'N8�R2��]X(���$F�`�'ȡ���.��w˓ HT:�'��1�Ǌn��!k��N:z��q��'
��gIL2%������@�"a$%��'9N\�RBV.q���g��p�'O�`h�S�M�hp�v� e��b��� 	�g)�&���N/��q�"O�5J�b�%#���E�D/m�J���"O8�� #EM�~�kT��8O�N�۷"Oh4�GrrcŪ�1�|C�"O��3��pbԩ 1�L�]�X�H�"O
`�C�&J��6�5�8���"O�ݨ`�s�T˷�ݥQW�Mr"O�Țp��;���3,`�@�"O�y� '?�h�щ��R&ى�"O-��� �8���@Q(_5�^��"Oĸ��a߿x){��]-H}�"O�PQ����;�
���Y =����"O:	i�j��x��!���RR�v�P&"O`hHܪM@��r��h�"OL$8�æ}L��2�@�_�m�#"O֝���I."(��E�A8sY.��"O�,{@/��ձE��
V��z�"O0u�R�-BC�aI�� 9Q�e"Oց;`#W.����%W��;B"O�����s�ԕX�H�B<d �"O֩���� )����M<*�p�G"O�Yɰ膩 �@���G�$Dыp"O��eGۂDĐ������>\���"O�if��f�z4���w�`�"Ojx�B	%(I���h�
 g"O˶&>d��[����E)I�y� Ͽ
���[5��Y,F�h����y�T,<]l�sg�7F�(Ŕ/�y"�	�)�	�	T� �g햩�y�m�#x::��(�`��c�O\��yA�_F��@����T�ʭb�Ɂ�y2c�	�N���!��\�CfFP&�y*�=�� ����?~��pɅAƼ�y�IUr�0C�m�Ic���܏�y⃂ �Bd���u�`$�`��y���!��d���q�ؘ0�.���Py�� �|p�D�X�~~R�;�EK\�<�E�T�H�p�cVs7�ȈY�<�F̛�3�,�#�J��2C!�\�<AK��V�H\@�H��o�RA�@��[�<��I��2���.K'\G��c'�Zl�<��C��(�ʌ��CO$Bye�q�<�ь�6I�!ie$,���y��B�<p�Q��R�D�I^֝��E͹!�!��>��"k�,u.���'�^$<�!�䍖?��Q�ɜs!"��"�P1!�� �̉`�B&�8���!�4c�!�dD�Y��1���̫����*�#>O!�d\#X�$(��v�X/�	0!�P�-��L	TC#V�M�!��P@!�$ޙiY܉i�7 Fv�bw)s!�$.?D��2Ŕ!4
x`����!��2.<�w�S�@��1��A<�!�$��hb�����N�lά��C'�!�$��5U7ʃ�s,ۂk:�!��J�o+���6!Ƨt�q�#ߢ�!�d��K��Uj�Ybl��@�8x!��,1YG��p'��'�N!�$�0B�dDq��3�ts@j��^�!�G	����&3r[�(T,!򤜀Y��#PHV�Jyn�8�s!��ݜab�4����m�^` ��S!��0%D����"$Up!�R��H!��>�(���C�+���b��>]!�� �	�G��R/���3jX�;(N�9e"O�\3�(�TlC�� ���(��i+ў"~n�	:"]
�g�=�Ȝ� K��?_F�OP����(b�lJp�[�$k�d2�,¯���^�� )0#C0�X@�I9uD�8��5�.�S�'T;�L��h�!�P�u� gBԅ�e�L5H䩞�6ǜQS�+t��Q�On���ˇK����93�\��"O�2��ec(c��ƨX0��`"O�q/�R�J�W��	?(֍k��'��	6 �"D���
-|����YqB�I�&>Lб�^�*�(+�O�g�BC䉔� |�DL�b%���'杗V��B�	�eP3 ��	���!�+?
�dB�I�)-^���)��drs�KR��G{J?%�2c�/�@%�ͼ+yH��g�j�=E�ܴ��@��S/(p�qw��X���D{��'3�ؓdO��QAn
?/�a+�O�����X"��mݹ`H=����	W+�	�<�J�ЦOq�j��"
�2 Ҩ9@�.��J��7�'i�!��؇dl<��{@�V$�D�MH�	Ex��)T�r�R���� ���P�DY�=�a}>iC�C�Q�p�ްf'��(Ɇs�g��rD�C[���iƲ����f���'h֐G�tcv��yu�P4���L��!�p�A�4D� *H#	�Z̲���-}$�P���T;�4��SF{@�;fIؑxR ۟<f�|*�c ��y��{��ѹ��U
j 
��3���y"�'=0A �O$PcPd2�I8*4p%q�'mڌ�R�*��k���*�����'m�(�P��=\�&��f�O�"�li��'>%���N+�!�ך.6�)P�'���a�/�<ƙ��O�z���L<�r�"|OU)� d`�L ����DH���Q�O�U"�c;S_�	�e�]-u�  	�'B���g� x�B�L5����O���D�4D)�6����	!#<!+A�C��y�"$�z��G�$l��D��yB"�3�����gdv��Ə��x��'�IZ�N�2-�&��Lʂޜ���'�a��ȩm�)���.춨���N��y2iLO�2h8@���<MA����yb��/�� c��	"��wI���y�nΥ#����FT�O;&�/W���'�az�n��`J�9�, BV+�N���<��k�*#��<C�Ӱ�*l�$��@
�B�ɣ.Ԥ,Z�hf�=5st�@!LO�X�>`�Wr���Z��Y�q�� 3',��<���&"˪EksLP`�jYZ4��y�<�U���(���a���Ф�V��t�<���2f�(����4H�9	ap�<��c[�C�,��W��0������k̓�MKS��>IO|J˟�m�!�����D#��?���q2������'cʽѥO��D)fx0��2Z9P�6&2�S��?�&j��c�! �N]D��"'ȅX�<�(ΕkT�E9��؃�|yz�	�?���'���`cT�Y�uNU�͟�L��� � 9��ۋR!����F�"���ȓyl��2�J0Q��Tj��ٰ�B����O�'�Z`3�K\����j1�$Xz�N��3��'����E
�i��\`U%I�O�K�t�Ik�����>�6�ϡU^VP)�'Q�:�ّ��o�<�!�4�0!*���<��ᱠ�7؈OH����(D��ɲ��ԕ5@`'%M1!�� p}z�C:*��p� ٦sH���%"O&i��U�I*(-c�\kB�����Oe���i�Of���@Cn� � ի߰w%ȥx��x�We�����̅Q��Ӑ�|��Z��-� �=���'o�S��?K&"U���Ucb��@h?+.�C�	���r�G5^��)�-�% �P�,�S<��}�pd
�M՘@��D��Z�xQ����Q�<9%��I[�x�HȦIx�����c�<YU��*k���AɞyM"I���J̓J̑��'�H� ��R�B���l�"ap�q�+"�Dܖ�0<a���MVB=��� eߑ��J�͙�<�L>!*O?%���1����BK�_-�x᳥=D�����.Z4���bLK��J��0?��O�Ósl$rG�M$r��"�ߑR��p�ȓ*����G!4Q�4C��H�<�;�4s��oDC����q�:�M��y��X�]��!�#&�8:�R����e��D�>��!1���fV������az��=	\\��?)V��d̮F�!��1�g��z/�9��$ma��"O��Чm��*�R��R0̔�"O���
®�@�{��V�t�5He"O�u��HGWwd�qw&^(g ��6"O,��[M<���� w�(��"O`�t�r�:Q�r��vO���0"O��b2�-e�pm�*]>�H�"O0(��H��L�&	���	~=0P�"O��r�;�8���E
�:-4�"O�Y��1FL�<I+E0E���"O���B�Ƹ4�b� H�`����"OFU�A�V���dȚ(���P�"Op,��. �q�$��1	�L�c�"O0�2
G�z(`��0�����"Ox����m�`4���  �^E�!"OD Ys�ԗF��5:�A,Z�ne�7"O���� J�;��4����*�z��'Nў"~ZЏ�y�ɢ��

k�O-�y�Y�">�b��S!_lTS��@�ybDPn>�+���eϚ���"���0>iM>�dn��-J��q6��/i��H��^�<1���?)d@`Ri�)`���@֨K��hO�1E{��Y*T�kbg��k�Z1��+����m6Uis��5!���W���{� ���$;�O:�PCg]DRڅc�,̏e�t�(�O���&_^����f�3e;d�"D���,�R��R$�t�S`�!D���W���!Y� �wj��/�ȱ2	�''�܁��� C��!���$�C��hO?���5v��S#��5@\� ��<��ضT�<�t�O�,�	��NV{�<y�UC��<1�BJ$��u��5T�X��ث٢a��-&�|���:D�`���{�������Tlf��i&D�����\(2�`

Z�t���8D��S� �@߼�I��l�BV�:D����A�;pZ��dȉ�C������7D���%�N����wd޹rD�4D���q�G�b#~���N߹}��1��M(D�`� nO�`�d��-�{�l�� '&D�̐�!<e.hb"V
U�h��4�6D��1�"�:b3�AT�y��\*g�(D�l`�`ӧ��|eb�m�R,S�*O�]I��0y����Ǒ�Ȣ@�"Ob��RL��NVi�էK�1�\@YP"O� Z�2޴bz������o�^鈲�'��/���9�G҅@Y8�$ �27N��ȓn������ ��5�C!��l�$�ȓfy���rJ#"��F�$|MB%�ȓM��`W�;4��kš�
��1\L)zr�\+J~�y��!E�cȶQ�ȓN9.Qq�Ƶ�d�W �#|(X�ȓx�蕸���3�2����$4t�t�ȓu�x|�'Ý n?�h`w$7�i��yGj<3���.vH��v	ʞ?+�ԇȓF�F�SݺV®u�� +�1���T��u@�(r�͕�[�]�ȓL���@��s�I˓��
j��ŇȓC�Z�J@a[*�J��� Uin4��l��Au�$<�-�@F�{�rU�ȓ	���@U4O���%G3�ȓ0��pQ��2y��U��l۾�m��F���(Q"��(��=��l+�h��p��|��)Eh��:�l[$��@��v�d�##���X0�D*��Ԣ3}Ω��V.8 NJ�������Q�i�ȓ9�.D�s�FZ�4�F!��jk`������ʦ�Ė{8�A�D/[�4U���Y���g�n�Vcؠd:\9�ȓY�Ju��cٓ-���B�����b�(0����!A�H�p��1�K�<D��9�F���K�/�$��C��J�<�T�>Vf��ad�*�<�k�A�`�<�&,8'����.	��ࠀ��^�<A���%*2�#r�� �)X�V�jąȓ������KL*�!���L1�`�ȓ%�ֽp���$Nvyat%�,{�*�ȓ:�D���d� �Q�mơ�ȓN,�KE�H�<�0�"*�|�ȓ�α&ߟh�t�p�@ԟ!8Ҡ�鉷M�~��
�fNH�n#�Z]�i?Pn8C6ဗj�FC�	�xT
��􏛑<�D�X �ŗ,kC���`6�V�I(�C����B�Id�Z�`�#d ��^���C�I	�!B)�6&&أ��<<2B�	1$�T�����\��̂�e��C䉕/��iuH_� $�1��>	�C�I9Pv�:�U�I(x����0DzC�I�=�"Vܪbep�K֣�a�B�I��T��X[��2fiԅ:��C�	��F��M�>E��:�cH�'��C�	��lX$H� �)$�ʬj�zB�ɐ z�hp���=Ghd���F
nDB��-�&"`F��l0�3��+ �ZB�0�$��H��p�����i�n|C�ɹ.w������0p>��Q��V�8[NC�I�h�Ѣ�=Y<��!AmT�UZZC�3=�5��F?�F���s�6C�	�!���[�g�8���[Q�Ԥ	�C�	�&u��*�E�H���x����b#�B��1�A�0�V9X��d�%e]=x�B�	�]V=J��ѕ�p �M،L��B�	!Pu�yP���f�ba`t��U�pB�I{��� +�M�z9�U�̞$;<B�"���g�P	�2AK1o7�C�	+.�3�nD�>Q*�@��8��C�	#txص��=%'��Xr��
]'�C�� ��YH%N�8,r��C��C�I�v�^I:���bU�]p�	y74B�)�  {�!J/)B|�!�XTR�0w"O�XTG͋#7d�HR�+]^�G"OhAP�.�7 uz�H!� ���%"O.��
Q��e�1) Y�f�z�"O&��7��0a�9xC��ɪ��c"Oij�D @��[�!�'I�8P�"O6�(�K�!?�ě��]-���5"O�����6%&�����i�P+�"O��oͮ2��q���K�GX0�F"O���<w����Ɓ	*p^b�QW"O"\Pw(ͦJ�Q�� �Qd�S�"OؽFk�4�恊��W�'F A��"O\�"�f�2��I���$$��"O�!a5��$k{�$��Z�O�Qz"O$����*"h��qԎW����I�"O@ XG�Ø�0���+����"O�P����ݶe*d�Ӧp��h�"Oz�C�.M��;Q��('0HI��"O�h�� Z�:bb�Q���X� �u"OJ��/��h�`��E����E�"O&-�4���0��4����.i�>�sQ"OBTx�c_�>8PZ��ګxd�Q�"OHd�u�ܗc�4��Ao�B�� �6"Op��Q�۸1O
���N�1��}ʔ"O�*�N���r�{��ʬ�Z��'"O �����]�H�cю�}�<ms"ONX����h͚��*L$�!��I�8|���%��TT-9��]�oq҇�X�[U�|���<��U��JȕD%ƥ0�6'�B䉦#W ��-~8:�f�+z�On�x��`�(4A��d�#f&����K�i�x	�G��<F�|2�_4{)��H�!5���`�;9�v�H�b�on� B�[�J���	��䨲�qD@@xP��).V�<A�������rM�pGFL``�
���i��]����F�ή�˵N� !�d#o��!I��K���@�왿�9�&��"f�X�t�f̖��	��o�Q>�����II�邬Y��Eʆ�E�Lf!�1(ƮI�ж�YzT�#LВHp,X�aӦx@�#L�A��T�Ʌ������'����b�.`���#3h�@�r=*
�i�5(�5z���+]k����$u���h�-�-C�ܩ�V�]�O�xͅ�	�E�z95,C�um~y�0�Z.?h�<�C�@�n)i���venY�Nڟ,;n�R\ws�D� -�_@ĩ�Mnf�M��'WNcB��� �zWʌ����wń2 �ӑ耮t������|PB(S8���$�!U�P @t��6J50)�"O�%�3N»>��<C�+f�-RT���9�4�Ӄ�"r4��R&�� @>��vd��=9掐�H�<2�A���"mx���6bۭa�Yc��P�]�<�DLW���*ƮY�B�ջU.I�I,� -Wz�z���qh��tnκ-�,� Ř���O���+��vx��A�,Ϊ	[B���K���@�:f�\���aR}t���Iu~d�s����Js��h���wI|y �j<bb`<�'���c�˂�Sg�-cÃا=ML `��{�'e@��V�։I�8PR��C�2��'�J\��f����zB�B*F�l C�W!O��1�faH� :6�:���1�r	�d�߲m�,rb�ª���P'r��y�����FLU�Y��z�ʊ�9��D(j���?y�ثk��8�q.�3�5Iv��>��Iq���%B��[�`�>�c�MP�!�8����}�'{��� �0H�O� ��Wj�g��(���ɇC�dj�H�=W8�ӕ�Q��Q���#j_���"�9%V��#��ĸ-�v%��)}�sB�<��Z�r*�Tx��.扯_�T	X6/�<KK��A���Qʓ]� �G�1MlR0��/S���e��dr����zם�t�,��Ã��z4H5{��ѽi���ɟj�ہ��W�az�ě1@������I Zj�Z#pD�9;4�J6�,�� ��2+�h!D�C����-�V�!�9#ن	�c�3���B*�������t��@;�#����]�q�Bpo;2c�P����]�uA��(��s����z8j ��L�q
�r�O����CA/b�N=��]�T�#2E	5�d���ɤtJFu:��	�'�f��E��	P�(P����$09������1m̥��Bo�mJ#�I*}Ҁ1�V��P�,RCF��&�(�"�p�ɓ(�R|)��3A{`ʓUKDQ�� �������r�4Z��Vl�	1Dsl8�Yw�51��lB(V�d�a��<��I�'�z}h����<� |!r�V'&n���F.AV؄mא#lqA�F�J�d�����K�r"���$	ƮG�S�<qt��0t�T�[���n?�� ��%F�~b)Q c�L�LU�0y6��s&B �۠nϞ��0�BPy2��U�V*�D��|[�lZ;]��a�?kT����M�Y�џ4,36�����ͫ�ħ_�l8���I�|�����
�'���%/�$�����M��?�`�f�cG�s���ə'^�����)����Q�*�<i�/�<���1}��)�'S�j�Þ�(�I�gD_*d��Эu0��A~A���剷J,�:��W|x���N�pq�L���2Ǧ+���&?���G�sKZ&
��q&���y:�0H��,�Չ�[��|��V|Nm�ǃC(x���bG�X;e�U'x�'F�H��%	r,���)_�Zv�+��J0�AsaE1v-џ�	�	�\�>q�p����;?�|���*��C�M%�M{��׎!0�Lh�^~���isf�1 �)Z�ؠ93b��0h�)Olq[#f�;X�H��|�2"��$;P�%iG-Wk.%�0�r~2�X��LZp�'s�1�1惭8>U�`�\��@Bc'=}�aܸ)�5�����O`j'���:0��Y#V�}*��X8�p�
�/�6!`�g��l���͉4��a9�cC�Hr����� �OV�Xd��`D�<���&Y,�t��ɭFm�邤�R��O�b�i0�V?��4�&��{$�	�'��ZA"G�G\�[���>����O�$��lY+O~�O>�+A%ȵa��Uc�ԁ,.F�g(D����u��(W��9l�ᓤ�&�I6b��A�Q�'�*�p�&�GL\�9�͞>	΀�	�'@Zt)!eѶO$����bD�� �'{�Ǭ�v�L0���?��M�'bP��,F9
.4���V�e��d�'a�1�0o_2�s�KW�X����'����
.H�@�d�78Ɗ��	�'-���E�P"D�.�af+1欀�	�'���h"��\��@�s�$ �"O�8��R*���`�,P��"O�m���6R��˄�ƥqֺ��"O���A�8VXT ���!<S|�Y�"O*�:u�Z)%L��T�Āy3"O���7��+D�\� `�-P���"OF=�)D��H��V�9�>H��"O��kP��MC��� c�8چ��#"OX ���,Bp�"�".�R1G"O�D��H04f6a��)qs��@�"ON):2#�3@n<���݌SP�d�"O�u�6��*a��5{�-ٯp^p�"O����oA�1'F��@^*D�P!P"O>�H��^�S,H=����>Ա�4"O~$����/~"��fƂ�E�< �"O��SaI�K,°ڄX�I��(ܾ�6��i��Y�\c�H�6�� �P�H���	4�-D�k�OַV�k�F.��5��ͱ7�bqsH�g��|��]�tʷ�GI����V��<	�/O;�d-1e��!����>s�r7�i����'�~�!��D�X��QٕzI�]Ys�Y/C��)��(��F 2\���('�ߵ�H���H��Q�0�z�Z�E)oj�<�"O��!���u6�e�I,gL��1�Q���{'����j��A9�q��'J*��%�@�
��%�"#@�+�d	p�'K.���R<=3��fE�����a"K��"ٓ�C�mA\��1+�h��|*�*��R7��Qǆ7H��`E�>O���-�>?�i"'��*)�6[� Ǆ'��[e�=�x"3PwE!򤖏I0�R.\�T'P)3 \��	�q^X�xńM�qwf]�e����G�$O�)8�� "qO�f����W��y��
�}�&��è��A0S����gOC9:�B@���[�"mI~��y"��c"���@�Ӗ�>��FG��?�^'`>$L��Q�o�,�p
 �6�`6��FAɀ��A	ӓ/0��7�E�Cs��A��3Wj�G§ށ���"��a�t��Ċ|j5Ȥ*Q'L�Q��Al(�Z�"O8��Sb҂
�fx��$���<��^�p���ړx�\��ʸ������g�π ��a
�>DΖ=q�$�h��Tx�"O����J��߬l�5��N�ĳ�
މ�0��m�'Y#��`>.��O"1OB�I1AWb�ۄ![v����'{F�aQ�Y-�����ȍ+y�Ȱ��C!dy����J�=�Ș�)̻i<az2i�&��}�r�7|˒D���-�0<Ivo�� ߬�V�˽#`�����g�,���I��2LD�һw�I���`��#͆�+�u#ӏ2P+H��'V��f�`�N�0A Uz��D��l��7�~�K!���ty��D��y҃U9f�P��!�){fV���?
5L����$+ �D�RK�ᓈ�L>)���j�����ʹ)f���H�F(<�ō��p�i��J��=����Pg�|�	��[��=�D�P`GL��w��?r��K�OCX��j��}��5r�(�����+��b eJ�ju2Y�*ݾ�y� u�"EA�=>���D� ��'<:���$��
DD�dD��r�	."\R�-_��y��V'[s�P�Cl������Dt�%���\ܓ:Α>�^�`��2���q�:�ӱ�\�|z ��\w����͇F����c,�:_�L��ȓN\���2 ԋ��5�ɘ}����m�T٪��؞cAq�h��������!I��эlǮܰgj�}5
���ڜ��w���]�6T �J�<�j��ȓM������M�=pL�&��݆�XH8!s�#�$-h�(��A$) ��\8��0�&L�}�)emU� ����IN�{!GG=#��Y�HI�3HB����bգ�!�%�����: ����)�9�� Ͼ82��7C�h��V^he�U��1	P�Q"r�W��Xd�ȓ!��	��G��!$'L%iż9�ȓ� ��Y�;��6�T�OV2\��'V�=�`)�54�j���i3C�J�X�'a<� ʎ���
 �
���'���3�X��u�
����!�'I�\�Ձ]�MC``4\+��[�'�c��Ho����	j��
	�'f\e�X����̎xe����'�,{s�U
K5	a��вogQ�	�'��!2ֿ1�~�c�lۨc�.���'��tjP ��X�.�!3�ޫ^��8@�'�v���M�*ffNt�CN�Snd��'�B��e�>Ev�sl����I�'Q|p��4$k`9���X�F5����'�ruq�`[
�h�Q�.��7j�y��'\��i�ρz�^8s#V))U*�'���s��]<,� j'�·$g�Ԣ�'�� �d��>����6��WC���'��q���Iv��LiX�'S�@Ys�!y!�U#]"D� 4
�'.V��,�氱�4l��Nk����'��҉��L���H�6�Th�'#���dזj�R�J���7��U��'�v�ʇ�Km`|S�iH�g�`�'� @F�1�d
�(�Mk �a�'�t���ֶwn��@�ν,��p�'�8���H�'D�@g��v�#
�'YlE{0��>. 0d��3
!�`
�'@p��
�H�T��4a�� �8��'�4Q�0%T�k�Аrԋ[.�Z9��'���DN�-F.�+VfU�J�'Ԛ� 	�Am΁��k9�	`�'��nJ;���C0�J�<��ݘ�'���Ǭ;�Pp[C��2����'�r<s��j��`�"��2�
��� �A�
�qIZ��G
��'AL���"O�����MR\5�P;
Nh��"O<�����/MƬոdF�J)d�h"O�t[bgʀ I"��`�-+�x�"OX-xP) � _�X�@dU�7@�w"O��	�2�yh��W;�@��"Oޘ��e�>&��c��F+*��`�F"O��)g�3�ne��%�Hc^�8�"O���E�*����'��9q"O�5 _iW��q����P��jP~�<a��˦cX�$�2��mqo�t�<� �	/%U���g����#�_q�<)�
�5/�;Ą�f��)P�/G�<�G�I�\y�́a�4�cA�<Y�Ɖ#2��I &䝴0:Q:��|�<iA"̫}�A���7��l�΀x�<�'�čn���z`/�@S��	e�|�<���RK�,:(��� �D�<����T�\[�H?�\� �B�<Y�*@�sI����ǻjr� p��U�<!B�ObA�֨_�F���h��L�<y�!	Р�hх��l�v�<7��0�,�J,ax�3�n�<I0��*�|lsnD_���{#Dr�<9c�"����+/hRT��L@n�<��O��?v8 �4d-ǀ[��So�<���\1F�Ll�k��x�ıå�HA�<��X�u�gd�*u�D ӑF�C�<�&W�V�87&mv�c�&�S�<!̉�pT�H��n��2�l���J�<y$�Ϧzr&�����N0�ݠ�Z|�<I'��`����C9�t)�� ����ppH��9J:�$�"~F�6鬉a����X����=�yr�y*��Z$�*?Z4��L����T�"�^MЁ"A���<�1' 	d�����l+#�U2�o�t8���	>^�`�9bC)H��ɱ�MȘdta��H�1�2��ēAd�YC2��*O}�9���"�b�Fy��En�q��+M��vd9s٫5s2�8��#x��C�"O�DMԌ ��`�7DZ���Jġ�c�P�h�O�zD�-����2�W&t��M�r�I"LvxvmI�y�a��z(8*�Ń�r����P�~ba��+��PP#�.�ayѦA���0�$�%fC���#_'�p>a��H�z��u ��*�]bUdL�T��ԯ4l~��	�'H}��ϛ]�pp1�A)1o>a���M@U�AΙ^�tb?ɐ!�ھ���C
��`b��3D�tiS]�E�- �\ �C��<M�u� R�T�
*O?�d������Д=�T�H�l	�Z !���N��d@���z���+~9�O�-��4�j���` *W�h�ɠ�`Ϳ:�@ܳd�'�DԣDM��K�4�H���(�L	X���z�<Ћ�"Oh�������{4n��mK�Qk �'�H����37�V����$x�T.�
ynD�I�;B�XX���5��k���`��U����,*��F|�&qYC�&�(��O���ia�	_�BըeL�Q�r�ON��D
,a����$�r��Ac`�T�h���H���]5�{��F�,��!�h��s��O��	��D覽��#�8�x`� ��c�G,��ڳ��"w�J�҆��E�\K�"���<J�JĪo�~�j�@�A"�x�񮊡p�Z���4���f�9Z��D/2Z\���?%B6i��Ǵƣ?aQ��H���p�E.� @xKv�	3CL�"������ �
�{6GQ�3;��pbI��y�Dp��8�C�j��c�ЂŔ�mMr��PE�>�{��<ف�Bt��pk4�ݾ. �HQ����$TGk�@���� kݑC�T��b���8��������Ҡ��c�d�Y��'7X:��Y0�#���8D��A�"�E��]q�#��`Z�3d-,;@,���?�ݠl�,`鱂P�($Z�8��Z�0� �5�[i��
*#N�T�.X?h37
�'�S�g Dn���×�s�P�(BAO9fzZ)84�K�^;`WZ�4�4Js�7� f�@��4�I)�!��$|@�W�	��d���*H��A��(Z?�m�2�o����<Ǌ�1
�(G���F�ќTE���W\�L��6T��B�>�%-��2f' I�`�w�ބ<˓`(I�ߟxZ6��D�x�3�l���E�O�%
`����6)�҉O�:�2<���*���6O� �c� mS.�b��!<O4��DE,�<JR�ݐM7E��%���"1�A�%V�����J_(��l��.���u�Ij��넭G�nk�-�S�E,/4p#�lF>�p?��o����MYw�O0h�|m���@k�$@Y�tG���X�d� $A�bU�!����#�ħBʲ�#s5D�@#�F M�u���U�'�V!�X>�&>*wi�pW]q�gA'z\��"�N�!p�Rc��Q0q`��O�	\�AU��Qȟ�d�>��y�AƝN�~��L�6.��uH(}�Մ�2��S�O7� �C�_�,�J}h����pX2�'��-���U���� H',O���.�Ew٩���7faR��k��C5h
���`/��4m֝�;AF�1�柄d+X�q�z|�Y�b/2j�����}����+T�D^xQh�&'���1�S�,�N�[L>��/�Z�dE���O��a5�
<�H�Cf{e��e�'�WƎ��c��2a���<1�e�O��p��g�#q'B��ig������u�Ds�O?7R�<�ʽ9�+�>i���Gg�?��I/n+�f�KH�S�O��!׾�E(��1�Z����g~B �.g`�p�'.NPPn�8i��ı�K%_<�1��$}BmǖO�`����O�Ģ�� ��S��"CPv	��Q�]dZ(�
��+�1���D$\rDȱd��.$T��[d�Q�'2\d�e$�O�9Y �V��A�!eT�1jB2��� Z`�EXw)ƕP�O�d�,0�P��U�V��tMi�'u��1��+<���*��:7pX�O����v&l�O>հ J)`�҉�J��gr�d�;D��p)F9S�&a��)Ȱ7  ��+7�Mȅ�'��y���Pw:)��� ��p�'�Vt���5��L $qZ�l��'dv���KT%?H0Bѣ�_�hQ(�'�J�;P)
c�|l��GD�~�P�'���� ���1|���Dƭ�%%�W�<��
�(X�}iSL#0��iS$��y�<A�^�>4c4,����a�I�x�<��섚\\��YS�Ԗj���Jh�<6"�H|��a!��in�E8���N�<���:�,�����<�D��`A�<)Qըh����`���.��D�B�<1��ܫ/|�9�!�5oSfx�q�x�<�F��LZ��E�D/�6��AL�{�<�WξA����Ɨy�f���"�}�<)���C ��K���E��{@�y�<!�C9E�xr��[u���f�r�<��($�:Y�_�EZ�j{�<��;,� ��;"4%J���X�<1�O�>������A�:4H1"�	Y�<I�� 
r����l�z`=Z�gNW�<�&F�rd��h��:y�b�Q,�S�<1�i	�F�Se��4}�����@O�<�t'J�:]x�ǰd�DuɄ�P�<At���fN�+��׭Dp�l�ƫ�k�<Ib��B�(���+31p����x�<�&bH���"ή:��MB&�B�<y��_3v`n�t��.iL��z�H[x�<f�#y"&�B!L9��|�<���ޭX�%3����l4z�y�<Q�%]�Ɣ v)R���\����v�<Q�]>ob��GG�x�.�ǃ
q�<A��J�z�3����N����7kXi�<��ٶ�����$2��(A��i�<Q� �[����Z�j� _r�<��'��ҹi��!#P1����m�<�F�3ڹ�6�հvA4XK��d�<0/44��`3�
p�z��A��f�<���4�b ��&�vD����J�<� ��
G��!ip Y�s8�'e���N�KX�h�b씎!���0�L��;�d��F�$lO���%�ԭp�*��#k�dḊR{�=��@V�$�NB�����sI�
8���	�#T���� �A�_�h��V�o[<� �L3�4x5��1J�C�-��D��-�39Fx� 瓝𚨀R�M6j�6�'�-E�,O�P��1H��U�䃁�wt��0"OȌj���j:Ȝ�g�ѭC���C�L(tx�|�f��}�a|"!��c��M��+>k�0��T�G��p=�/�6
�*=؁�x�9t#F&x�N�B@�Yu�Z�� a%D�T{��Z�5<~��х�X�ٱG-��ܸc��F�?�#2�U5Q��8!�u��� 4g.D�@��+�ʂ�����2�x���6
��y�l(}b�B���`:z� 0DX�v`x�B�Q	S�!��z!Y�P鱴��9���A�_b��U��JZa|�̜�K�l��L��Uʳ���=)�)�4H|޵�'Q���5hKz1dL��g�"�¥�	�'��a���-�%��-O�^�q���\+7, �G�d���'\���bƖ4�|3!��!�y�H�������* �M�y�*߅H�!��A�v��Bc�L�<ٰ
�4=������O��qI���}�<����+9�R���,G�S��а�]z�<�D��!"�\��L�[��0Ɔr�<a��>l�	j��ޥ5[��P�)�s�<ycOZ�[	�e����)?��p���g�<�TmG�~���CρAɮ|HN�k�<)��&v,�AV�@�G�j�c&�	{�<a�JR>lTU2i(Φ)��oPq�<�R�
�V=�bGDROĔ���g�<���`�j0Q' �#"R��t`�E�<i��D����J& �D]��NAA�<I�	�l��-y`��&�����d�x�<	"�X9*1A� :Z8�Q+Ʃ�o�<Q嬘�/LdY�alL5~yڭ��N�h�<IW�`op4����7���D�R�<A�&	~�
�`G-�0 ���T,�u�<y�s���;��Ev�s�<�A`_�v�B�i0�P:(��Ӧ&
`�<qď�5G�j�q4��8N6np�`.�G�<���O5�B�PA��ED�פA�<9ue�9�@d�ҫ�4��ax��U�<�u�$�j���*���"�Q��4!0��G�L�f�-T">I���6i�	�k�W�  ׄ'D�T�!��x\�uc@ꐳ9)���Dg)D��i�!:��	[���/�-"sH#D�أ��˷%�
��c�x]F���g4D��A�F�(g.���d�(iZBIS!.5D�B��=�V��5�V�Q�EY�5D���D���;�p��%o�`���>q@��W��H�<EcC�T�M��hBg��X�,��imJ���R��@(O���T��DI�W��7m�(h
���'%U�]�M����z6����oӦ�"�����ԧ���	-vm"u�AF���q��e{r瑦R�"~*2��I۴����R�@:6휖"B\�Ey��	ƻ"���AI�1�@��_�zTQ�P�W�O���3!$��B<���gQ�7^-X�{��[���'C�b�'���b�!��U.1�O��ڋ��i>a>V4��g�)|l�u2'�����5�hOq�����r$|��E��t�A��1U�b�>�O'dc>a0 ����)���=}O8A*��4?�CO#{��t�D�/}�𩈣s.Y`g�ϟ'���hL:5��f�������$P: ��)�p���8t�\&c<�y0��S�L�G�^C&�a:6�s��8u�{>U��O��~4�۱�̥mE�3Q�X�&��W3O�X�F������	[�@���mI-1^z)�o��s߲a��hJh���kY�������� |�bR���Q���]�Ƶ�3�'Čĉ�.�_�S�O]�\�ə|���1���,!(N�����5>���|���.u�`m�<Z��hC����(����{���Ipa�DL?,�ر`�`O'h|�z�̉���i~�r��)�)k�.��R'�L9@�)`D�9�PB�I\M�x�!GB X`�l��FCBB�ɫ8^�:)��pW�m��^�lB�	=�P�B~�������b)B�I�aqrk�G�>[N|��T/�)P��C�	!�F���l��0�'��_G�C�I�e�$�¨�<����É5JjB�	�C�Ҕc�g�>��t`�R�B�	}���'ŏ)��5�ņ��c`B�	�{ǘ�ٵ.J%B��1���\~*B�I:m���W��O�h���_,PC�I�%֨ɐ��D�<@(s#'�3/"C�	kB`��H;,�$��	cUC�	~<���r�E
?�P�aQA�|N�B�I%N�<\@C�O=p�zm���=e0xB�	:p� 5SgNӥ/��<�q�Z'{�0C�_��}Ad
iF��w�Y�?8*C�ɣ*H����*�J�8�&>@5�C�I�_TQ`Gȓ�Z���Rӂg��B�	T���e���,���,]�OtC�I9~���h��C����T0DC��zJԉWΑ�H���b�;J�@C�I>#D���H[��"Se��e�RC��T!<�5K�^����vՆB�?{�9�� �4r0��*U��B�	��0�"c�|��A'J�&VrB䉒F�I3K�I�j�jpe@0sddB�	���躅	3~�L�q���}S�B䉫wY�Hr*߉k�6d�m�1ѴB�I"g��K���"u��{b�Z:6<hC�I����n"��]�1�vfC��t{���W�ʎ$`�QqE��,4C䉯F�P�Q���pi�p��?�LC��&-�` �Mϊ1�4٘���y�.C䉟^-6�@�įq;u #��dIC�ɍY(��0�9O� J�ˋ��B䉪]_T�p�� Wm���q�(B�	�H�S!��[��a�4o�(B�	� �x	���	i�0 ��6q��C�	�0�<�+�J��7��� 1j0fB�0�t� ��5R{�ݫ��P.}MC�-"�B�)[�ta��b&.��B䉺4Q��Z>1�R���[�|N�B�	�@=�@+���1XH%����?wj�B�	3�ޑ��N�J����/��B�I�\�B0�<P����g��B�	%�l���ɾ �n<����1O��B�RE��A��T�mJh�4�̬w�bB䉘E��e���_�6�"tÅ@L�C��2\��Aq��>Zjf�o�|C�I�L
"�jq#8���)c̪	KFC��''BF,IǠͼ'�z!��\g-C�<G��9�$Q�v.��� \��B䉸*�����X5� P��M[�_q�C�	�H�T1�H�@�� xT���d��B�ɪJ����%e;aoL�rW. �y`B�I�ӡIW  ��P��X|�C�	�d�0��c� �g�`���ͣM{B��sHI;�J1�T�*���qi B�	2a�^���/�!7H* �u�yC�)� �yR0�/d�ܥÂ�m �!�V"O��R"_j�&���'Șz�%؂"O�P����S�"���f��.e)A"O����g41t�I�rE�h�nTAp"O T$JӦ9�2���#��X��"O���H>u2� N�T�T�[�"O:��d�^�!X:�Yf�ɀ9�P� �"O ١����%2�����r-R�r�"O�yB����N��#hԴ^����G"O��Sm&`:�b����H�"OXMW�E",�sg̉�U��@��"O6%�%e�(^,��`
K�H���%"OV�IPB��@�4lkd��1����"Ox���K(2�`�ڕ��JV�`�g"O���󈄫#r��gk],n��5"O��#�in<X˂���*���H�"O�I��_=<��aJ��G>@���"O�LYrI[�#޸�qe��71��98�"O�<��%�[�D��eЖ? z�"On�#r�F�hH�Y��^34<��"O(к�lZ]�Xq���Ĉ�6��s"OԬ`W��0 tH�BE�J�F"O�8����%<�z���12jļ�q"O@À�ƤiU�.�1,2� �"O����ѯ%m�BV5I�y��"O�	��c�/f_����8A��z�"O�H����*"+�9P�"���t �"O.�����E
�9bF"I� Y�V"O���*@�LƖ��!��zW(�{�"O��x��c~�����0c�l5�"O ����v����C�X,�1"O���Q�)I8�X��-5�4Ń@"O���5G�o�ųe�u�j�"ONXv�״_K��;��D�:h��Y�"OB8�6 ȷ)s��"�(�iN�j"OV�Y�S�I")e�̉o\mC�"O��� �0\���T���:8�/�!��B� vЁ#��(����!��a�tp��O�0�ά����8�!�T��:,˂L��	R�I�!�$���<���@%h�HDФ(װz�!��*��)��̐Z��cQ�ё@'!��Ê|��L*Ā�7b֌�Q����/!���)~�ˀ�Q�0k�>!!�x�����C�I�RA"P/F!�zKnl"�}$ъ6����!�$�14#��X�!'8b	ru�P/C!�$=
T�x;j�6Q0|��ߩB�!�߱��90��.}��|A�4�Py�E���x1�N��=z�z@Ԝ�y҃
9\����ǎ�1Ҧ}�m��yr� 3J���fލ&�%����*�y�+,� \�%�$�:q؅�
�yRQ��	�L1~Ezu ��yb+ػ�2��T@�p��4�I�y2�P1m�P*�G�r�YBT���y�I ,?����8Yu�@�C+�y"�@ �U�"�$XZE����Py"��,lF�#�E�Y�������S�<�d�N#!BH�EK�5��e��@�M�<9���]��β��X��K�<Ɇ���W�Fux�l@+6����O�~�<�DNY.`��ő�f	�K�z��I�y�<gH�B��9�,:j��YrH�L�<� �����((°b���#Z7�I6"O>=h��
Y�!3WjY 1>�x�"O���E��:�4�G�!Z'$e5"O���φa�&E���!�m	�*OF|�n�T��%)���K�\X�'A�ʧJ�%)8Ȱ�Ƒ&4~��'�����W�`|������Q�'��x;�@�l����g'�	
��d�	�'�l��ЃZ�V��4'�6���S�'bh�!�ț`x�I6+Q�0�����'�q�+Ee�� z]V(;�'����J'5���lo	���'�`%��X�ڔ��Ya�����'����`j������
T��� �'< yk���:	#DD"�K�0��
�'0�u��$�K�H��B�M(�o@M�<�wb�	Z�dd!��6]�*��T��H�<�4��B)��g�	;Zk5�Ec�|�<��B�T��P�s�C8�Z���Q�<��$KA:�Ȓ֊~�X\	���N�<����p�=*�Q���|� *VL�<�7ˉ�9`�S���Q�O�<a%)�'r�
�aٛa�r�E�<a�搐)x�1J^�%V�II7̀Z�<)�I�k4>`3%�Tp��� d��R�<A"�M��x'��R]B@iqiBY�<�p��9W��a#���|&�}�s�U�<�c�AD�%�b
�+�� �MT�<A"��*��#���#9�l�k �.T��K(k��X�ժЛ_G�Aڶ�(D��p������ӑ˜p�]I��%D��Z�`E�~ia;��=R����Q�#D��ZcfY���;�!�	v���s�"D��S�* <K����JM2�hj�#D�hy�g�u8xͰ��	+u��e�?D�����."�&��B$ǔ�y2�=D��!g@G�Eon!�׻2�PH&����yrG�0��D(f�ը~������yB��c����'
�R�)��X��y��˟��� ���L�}aa���y�`T�b�*$sR�Ĥ"yִ
1���y��4:��h+���I��I��J��ybnH�¥
�;E��ݪGƑ��y�#Q0�S

�{@p���0�yc0%ṑL8_����i��y��uE4*ޔ�s����y� �*`��d��-HLQ$%�.�yRk_wk��S2b�̄�ق���yB�:�xd���򈫂�y"#�i�`$��O9|����&R��ybܺ6�Ќ����,��X��喷�yRi��R�p��8n5L��r���yR�I�q,�$��Q3p�@��J��y��8x��dyV�ȝ<(��Ф��y��Ʉb �BRiH�58������y"i�����k��0�q�/A��y�G>�͐��[(�5���E�y�ㄧs�:I�v��Od���ʟ�y2��-�D��@��I���(�*��y��"^b����؁luĠ�	��yg�D���C�ǘa��!:�	T:�y�f&|�@A�F�Mz�ލ�y��+eR�m�.� $y"dT�y�%�|��Õ8Q؄�q�!�y
� ���/�F�b�2�ʃ�O�a"Oj�Bb�!M��$��k.pֱc�"O���,�%F�`1�� �Rk��"O��N6al��S'�Rbj����"Or���B+K%H��BFU:�j#"O\`QA�3k@q���!oҔ�"O�m"���p/�]iZ5V�!"OX�j"C����E7H�
���"O�b�	   ��   �  i  �    �*  �6  }B  !I  �Q  1X  s^  �d  k  Fq  �w  �}  -�  ��  �  `�  ��  �  &�  f�  ��  �  i�  ��  ��  q�  �  a�  ��  ��  ��  5  w � ^  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.�T�DxB�'��PnS�8�2 �f6Q��$��'#j��G  �?�	{7�>� %k�'A�)0�˲e!>�i���%��ə��(Oz�J��_�c�q7(�4GW�ȱ"Oр�Hr�́a6-�E�	f��E{��i�dI�hSm�?�4��Ń�	O!�?�[5)ɂPɌIP��vY!�D+q#b��@^����A�芢
I!�� ���2iR�7�`���R�/PFxe"OP���]���A(�1�4AV"OPձW
�=~�����T�Z�[c"ON!)�fi�	5 �H�4 ��d,�S��:6T�����x�d@�PoxB䉆��i�7�Ʌ4�0�sl."J�"=IǓ�VUP�͎
#nDc���0���ȓu���Т�1�Рxԋ��B�J�<�指�$Ҏ�3�Kh|Y��B�<)��ݧ|@�����E�D��v�<��胹����g��>6X]tg^n�<a�B��m����w)�C�ɟ��b/��C��Y(�r4b�O�����7� ���I��&�PU8�.�x�!�F�3@(�Q�K?<�X�pG+1��	@��̫7�\�Mİ��nW�_UTyKa
-������~¶��k�%^��L �f K"1m�O(<���S��3F��e�h`WGK?i����n�NQ��N��a����$�@=c�C�	�EP
���cJ�z�̀�C��_;J���<��'����O�3�I9Hj)�.@P��5��8<�DC�	� �y�cbN*B�{����M�C�	o�������9��%Bm��Z%�>��)�#Q�����g�^,ц��[!�Q/�$�p1��6a���F���!��1&�̉�"��'�zDBcFM�	!��H��Q��Q�qc�;�$�%7c�'�a|�O$�4��&�Et�2�	/�y�F\�r8bf��st�4�p. �y�G�2:Ѯ�15�a�2,@�I��y!U�p�n��7��3Zcb@c2ب�y�K��*��U�N�`V<������'�ў��ȍ�E�Z(
��2�Pc"O���R(�/(�z���_�{��hB��0L��x��;Y�ȍH�*W��4����y�GO1�DՃ ��2�j�# 3�y"GL5~X�"�<��H��yR%�|����!5��H�숝�y�埕t�\�ƥ�GfU!���y�&֗���9 �O+D'��R�b�y��<s�|y�T
E�?���rʔ0�y���lV(-����%ېP���	�y�f<V��v�T#�����2�y�윖t}HI��/0_|l�e���y2'   ^"���*E#h�RqoI��y� �60 ijQ�>�>���H�yB%�s��h�V���=�V�Rd���y�G�7<0��!�mS(*B�PDB^��y���xQ�D����a��Q�y���9P�Z�����ty�F��y�M�'e�\���R"����w���y2�.+��LyV��~�@`�!B��y�b�2���zb�3.qj���)��y�C�=F�o�#S88Y6�Ƴ�yRE�t/�@��<U@����U�yr�٩,HY9�#I4W ֨�d�ݰ�yrB��Cl��uiO,{����ʑ�yܑ*vp3%'��K��P���	i�fO@LD��0��ƛA(��ȓl���ce�}�ZP pʘ1q�Q�ȓ4 xI���c�,��D���A�ȓ *�m�(�� ���
66m�ԇȓAW^�2e���5A=a!�� ���J��!���l��������S�? H�ق��"c�����s��!�"O
����M��HP�� +t���1"Ot��c��'O��	�B � ��kg"Oa�4G��T���dI�$2�2�"Ol��Q)sN�c����'#�-�t"O k���,b&��5<��t"O���T�#$?bl�g��1��� 6"O� �pa¼�0|Sp��03��Y"O"����|�����V�	���%"O.P�b�ۯ/v�����k��c!�ڂ/ov�AFl����I��+@�6�!��u��x��d.ƘUʏ� �!�dW!=~ �����]%0�(��:�!��C�j�C$)Pa�G	�1�!�D��w�6���p���(���C䉆��x���X�	�ε�b�EV��C�ɷ<}��;0EL�j�	I3(ޗW�C�	�|���v��g��-���APC�ɭ\���C�͊�4����˸ PXB�I�(u"���dDP_|��R�ɋJ&�C䉊5���*���T�DmKJD|� B�I�t�xMz&��8�.ٺ�IA��^C䉡/�n�.6d%*e�@> }���sSD3¥�O�q�/	=z����ȓp�\I�E�P\�сN7n�� �ȓ4�zPP� ,"�|����.]�(��V��VE�$��2�%
!}��`�ȓ�2�36g�"v,��*		W����t-jv�1�2����񎔇ȓk��
�eׂ5�����J��X��Yv���N�w�
���Z�;{X�ȓg�Zx�5�N3�f���#L�%����#�����J�J�b�{�K�3g8���Bq��t�	�=�N|k�H$fK�H�ȓ
�B�Ba�D5r�(e٠$�B��ȓ\}L��Q
K�G^��Xp��#��$���8-Q��جJ��U�¢n'�y��`��@�#�^!v$�7e��(&���K�ɚc� �N\;g,�<a�$����,��Ǡb\�ď��s.���S�u��O��^��=����?q]�݆�!.���U���җ<:U�Іȓ�6���	���R���;y��L���������h��e�tQ�ȓS�H�2�c��Y�!`Za��)�ȓ���)�I4�"7ɔ #��Ԇȓs�~�#�/a��┘U�|�ȓO����Ȓ��)c��>Y.�ȓO��|��]��`q��5�de��k��x��LāG1�LI n�Gp�X��\�V5kd�L�6�:©ݾ='����\�T�؁ŃO��P�$�Y�?�Lx�ȓ���ů�*~Pek�f�6;�D��ȓ1����`^�zt�	[u��(�>��,3,=i�ą�\�*���-�=��G(a�7�ݑ+���2M 0��!�ȓJv���I;�q �ϗ9kx]�ȓ�4hr�"=C��A�Iʑ=͆��N�|�H�j�hD>�����^��ȓ5��{���1(��v�˪d)�ȓ�Pm eƇ���T'$i����y(�13��3\uT�iĤI H��X�ȓp�<E�V�-�0A�MtK6��ȓ�6�A+�T���KW�ü=�~���S�? P�k%H1�輣�+C�B��"OV���U)%�"EhD�Ow�l�'"O����OB�UVE���!�|Q�w"OD%Z��l���&�:k�<tH�"O���0k�����aH ������'���ٟ����	韨�����I,tvɲ�NE�E����'�|�I�`��۟��	柠����	ɟT�ɨ =���V�Î[�`�Ƈ�*N-vd�I֟�	ҟ`��֟���ǟ����X�ɕ#ﴠ�w �4#p��螄p}��ݟ8�	��P���$�I����Iğ���_�
 �t�M!���b�G��]O���I����	���	ϟ�����P��ߟ|��9}B��a7�Q�l$X�����z��$��L���\���8�	����	��I�0P�ea
1� z&�T<}8���ڟ������	럸�����������I�PA�q�ӧa��]+jD,�������	� �����I�������I3�$AQ���-B�m;�W�8 �9���,�	ȟ�I��	П����I(c3�qS��^�B�@��W*�=_'(�����	����������I����I�)u�T)vB<";��fLħ.+RT��ڟ4�Iǟh��䟼���@�I�|�	�w��)�Ɏ6(��1�M�ff���	ן��ş����d�	�h��ϟ���	V���6f��(�,@+12>�	Ο���ן��I����ڟl"ٴ�?9�}D�K�n H� �ON�-�QWT��	y���O,�n�:�^L���ܮ*����EK�0�RP�"�%?y��i��O�9O��$j�HCv�X�3e$�a$
<���ON��$x���$��|�O���3��L�[CJ��r�J�"В=��yb�'��^�OV� ��	9º����J�+'�D�h�Ƽ�5��*�'�Mϻ;�P�6�T�!L�R���:]�	���?��'�)��<���oZ�<a�P�0}bA�g�ƦVy#��A�<i�''h�Đ��hO��O&lög uD�EfX�R�lВ`<O���,��������'+p�s#�P1F�����HO#Zv
9j���c}"�'��9O��k)�*H�G\�a%���B]~��'�`��5 �ݘO�b���]����$�d5��h�$rh�0u��Pq�Ibyb�����T�Ls��B��N)\�ېq/��T�Y��%?�@�i��O�I��k��J��*�0�`��|'�D�O
���O� +��a�H��D$��t���աBtܴ��dB�i���#��U����4�L���O��d�Od���h���!�?
���N�,<��ʓMԛ�E�u^b�'���t�'���z�.Hzn��è=r�t�q��>�f�iL�7��n�i>E�S�?u�c��(h���Ѕ�;z��`����G���o���~B�M�
�4y��Od�'�<�'F�����݇BHx0����~��'�R�'+����Z��)�4h�L���.�-i�_�+Od�r�A)F��̓=v�V��_}� cӘtl��M�d�̯C�hJ��\'Tz,zZ�̀c)�٦U͓Un,�Љ�9\��)���y�'�:�������nUJ��w�L"lH�����<���?���?���?Q���jU�}�t��ЋG=C:Ĥ�4i���B�'��i���3�*��@ͦ�%��eJ���&u����ٸ�gF���N?���z�$��_?;�6mv�X�I�\/���sC\�-������˘=��H�0.R<="��Y�	Tyr�'HR�'{2"5�����$W2�%�5*�
R4��'��I��M���Q�?����?-�U����5uX�k�OJ./4Ljҙ�\P�OtIn�
�M�u�x�O���e���4C7��� �+�+1H�`9�e9nI��m�<Q�� ����b�_�V��i��\������2�4��֟��ǟL�)�@y§r�NA��x0xր�y��S`Ps!����O,$n�u��V��ɨ�M3 g�>�f�2�� (rl"Iz�CM�r�gxӈ%p�wӺ�ɟ��T���I�@y�OX�$� EO>A��`S��	�y�]�������(�I���O�J�(#
˟ �d�W/,I�%8�q�l�C�O����O𓟀�D��睌];���W�U%�
��k!\Ǝ���4��v�%�4�f�����(A{��I�B�B|Swa �1���eD�E�<��6u���Ħ�1�|b^������(*�J� ?E���5TM�0�!䟐�IƟ���Lyb�jӢ�Q�A�Ob���O�����*7*y�q��-|�|�ː!-�I��ė�U��4.��'�8�{� ���B&��,HJ�'����dNV�R�TY��	�?EA�' da�I�I���{���;Z�6e�r���2��	������$��C��yר����I.�\a�nC�L���mӸ%���O�������?ͻGB���Gɺ-�G�2L"`Γ+|�fy�$�lZ�Pa܅n�<��c �u�Ӥ�?5��yh=�J���q���A�wyR�'��'���'"�[�D��ѳ�	Z7X��6//J��	2�M��#\��?����?�L~���_0:�AE�?s�h�RPA@�,� �S����Ŧ	�N>�S�?%�g��HZr��#N�8�"$	�H��hQ��%(4�'R"����ҟ���|�W����@F�|)F�(M�+� �֟(��ߟH�����JyDo�T�J� �O�x��V�T�� ⊃pta���O@m�x�\Y�	ßhlZ�M�Wm��!D�!*�O<�(��SCE�-��4ٴ�y��1Aj�"-Z�?YC�4O�t����=� �8f�b�t��N��S~�)�0O8���O�D�O^�d�O��?ݪ��,���ڒNY%s:H�������I�,c޴e��Y�O�6��O�˓0Қ93ק�!3?�(�W��?X:Ą�|r�i�p6���]	��`�
�iݥ	uF�g� S�>���jY�J�X�y�@�ԃ�x��<��?����?��
��B�|�W!]��,��d��3�?������æ�`��^ϟ,��ϟT�O�ܑ��!FJd��Q�ۉ+hЉa�O��'�¾i3��O�
w�||����{���%d
�P���p����	 �n���4�4I �'h�'�lq��,J�n��PIO�v�ek�'��'�"���O��	9�M�����{�m"�@�Y�*�j�%f�l����?��iC�Ov�'��7��ir���.
�D��Ip�ԌW�f�mڜ�M;�m���M�'~���uH:4�����#+��U.Xtrs#
%M��$�<����?����?����?�+��� $D̳�L�X'�V�Ьz��Ħia�@���	ٟ@'?���4�Mϻ;� &�+��ų���=0����'�i`�6�Jg�i>%��?���n���̓#,���GX�Q�fUK���!}�Aϓ"~��ɕ��O�*J>�-O���OD$����{l�q+Q9���1�&�O��D�O\���<���'���b���?i�,���R.��"��d�$?֤ъ2Ϧ>Q�iJJ7M S≃<� yJ0��1b.Yb�,��I�����Us -	Qy�O�\��I�$2�n�)v"H�G���fa�&R�'��'$�Sɟ�S��m�N�	 ��5�H�z�c[�����4Vrܙ���?�2�i��O�. �e���{˒9)X�Z�FϾ2��dӊ�o�/�M3�� ��Ms�'�҈U�4c�����2�$��0�-Đ#�$QJ>)*O����O��$�O*���O�5p��ǘl��X��#��&���<A��iI��Q�'�R�'Y���b&\�,�@��R�ՔYM�}�Wi�j}ne��EmZ8���|����
��	Ϭq�&���"rP)@�,:<��,���A hE���kS��O�ʓ׎P�*�$��d�!"��?���?���|/Oh�m	t���I�Fv�� �A�.�,��,Y�r}��ɢ�M;���<����M{��i��؀�ǝ=PgD����+X;���#w��6Ot��59�d����|�Zʓ����oҔ��D	֖`�X���fL 	��̓�?���?i��?!���O�~��J�TO@�u��,q�0�'�2�'���������'�R6�:�$Ҏp�VC"D4���B�X�����x�~��@l�?yY� W�����?��c��^({��'Sh��)��Rn�%��
�O$|jO>�(O����O��d�OXha��V�}O�m���)���#�*�O�D�<�Q�iP�Q'�'���'i���O",=2"gИ3��TpsaY>j����O@�'�7M��	L<ͧ���/N+\5�,����) (-�U!��U��z���M��Ry��O(�H��4�'6-ɲ�U�[}����U]_"D:"�'�r�'�����O�剒�Mw/�L�Z�9��T\���7j�q�Z����?�P�i��OJq�'��7-�d�j�V�*F�cj�J�X�l���M�g�MK�'12��rqV���S��I�[_<V� an\���I����@yb�'S��'��'J�W>��aÓN|�
Eg.!h0Mh�8�M;�O��?����?�M~��T���w��xȅ#A�|چbTj�	E�4{�Lo�0 l����|��'�*�%�M�'��*P+�)$}R�Y���>�ve �'���@rF�ٟ8�s�|2V����P˦kN�_��0��lϻ.��J"�������ڟ ��fyB�r�dxK�G�O4���Ot	2����v?�\+�'(2M>��j7�		��d�O�7m�h≹W�`��eE�{�x��΍�5T��I矀�ǈ���&,Y�kyB�OT ��	N���Kj<��b��[^��CX�(����?����?���h�����:I4��1��;^��@�E��ut�� ԟ�õ��O������=�?�;n\`�àf�-���Q���?��Lk�&�y� l��2�n��<��\iӀ�j����S	m{��7'��$0T�2#Ŕ�䓦��O����O��d�O��$�i�VL�Q)Y�5d� p*��x�ʓM뛦`S���''�����'��ca	��f�� ��G�V6���>ᕰiz~6�Fa�i>���? w����Vp�U��`�ł5���8���UyRVR[���I3r�'^��dP���;������] -jxe��ß��	����i>��'Rb7�����پm��A�[�ܔtۇ�!$����Wʦa��R����d���!+ܴg��F�O�C����'M=C���E-Uh��'�i��d�OޱȶJ՟��3æ<A��ڿC4�F˖���n	��"
8��'���'���'�b�'����(2��HQ�E�'�S�:41�Tſ<��do��M�2��T�'F07�9�䆈{��ؙ��U$9�{�bY� :h�$����49�&�O��5`�i��d�Od�(a�]�3������: ~�����a5��'��'���럤�I����	�@�dД��@��eH<������'��7�H�L���d�Ob�D�|�o��C�����_i��ĆMp~� �>��i��7�Pr�i>a�Sy}�M�DbPZH�W �t��G8t"�EFy"�O�� �	qS�'����Ѩ�0LV���5!�ҸZ��'�r�'�����O�剴�MSW�ݨP�1���#�T�¤�n�*��?�g�iU�O���'��7-�#0dލC�!��J���1��׎,�V=nZ=�M�c�ӻ�M;�'��N��D����� z�ر�ZD��l��.HD�q!�>O�˓�?Q��?���?����?�F��e%�4�g�%S�ЛF$��^��qc���Qt8X"��?���ڛ��d�w�|�$c�$���!U����P+	"U��m��M�`�x�OF�D�O�>\�ƽi���ml@�z��5{g0PR���ĩ*�"]���"���O&��?���]��5�6�?q 䨑�Z-sP]����?a���?A.OR�o5y`pL�'��H^�F� �+�e��7�yp�M��O8��'l6�[Ԧ�hK<I�'Ynp�Pa�g��azg���<���X{�$h`K<M�&�+On�,�?�
�O�X@�����h���M	����t�OP�$�O����O��}Z�zǮ�K�e�d�=�N�6kj|���Yp�F��.g���'O�7m7�i�i`Q�V o-$G�
_x��fBu�ڴU����b���hƈm���|��"ҍ�4�:QȊ�Dxд����.]��S���$�����O,�d�OB�D�O��D��6zF� E�&b���BB�#{����֡Ƒ�2�'��O��؟�i�͊��>�@��b0��C�6���������4[������O��T�H;Kr � �ߣZp@��w�̧}�f=�-G�i*�ɬ2�1���'���%�(�'bF����R`�A�^0T�ر�f�SП�	ӟ������{yKp�֐��	�O*���?3j����[�/Ϙ`rӉ�O��oZb��o�����n���M��U0� 	���FZ���Ε�U���	޴�y��ȉv��i��IS�fJ��T�s��$�>l0%���]�W����Ml����՟�������I�����b�(7VY�����.%z�P��şX���M�����|���09��|"I�16p|Y�'
L�us|�6�{��O��lڔ�M�'Ӵ��4��Ē�.l�Xaե�/h�a3�̋!S���9FaL��?��8��<!���?q��?)�I�)�<L���R���;��Z�?����ZĦ)�d��ǟT�I��O�t��7ke����u�B���O�9�'�@7����SI<�'���B(E��D���ü=St�T	E-�"��N��$�*O�	Ǌ�?��#�$H�ژ0Ks��D�<"A*GP"����O��$�O��ɭ<���iR�(ؕ&�	� 	)��G�d@ؠ%�]mr�'�7m9�I-��D���Pg'7.�JUb O*L9�6�F#�M3�i��=�d�iG�d�O�y�@�����<��G%QՌz�aΧp�ܸ����<-O����O���O����O�'un�#@��="G�H�ɞ�oNl��i@�$��'L�'���yb�l��a�,5[���~��e��@���qo���Mc��x�O����O�Бy��i,���j��+��T�ʪ���36O�càP��?��n(���<��?q2��c��$ҏՈ^t�2����?���?	����$Q��)�wOD�|��ߟ���$T�,Z�@Տ�R9���Q}��:���̟�m��l��9�%Ȋ�"���� GA�a�0�Γ�?1�L��VJ1�ڴ8����?���O���ѲR_n5`D�O@=��&�@z|���O"�$�O@��6ڧ�?�E"�`�H�ÃN	)f��T/Ǥ�?��i�� !�'��e�&��ݞ~� -��h�'�&tj�
:(�	���`ڴX/�& A�Dۛ�4O��$�v�h����A�DTѶ�Lh���.Ϳl߂U��*-�d�<A��?q���?���?���޶d�ua�CͲ�r������ēĦU��%�Ɵ8�	�,'?�	(����Jǉ�8�rt�	<I��lh�O�lځ�M��x�O��t�O�Ht�b�_E��'Z�i>(��-��1���(�[���0lJ�z�Ң�}��~y�N�H!���0M1���'�Ub�'���'I�OP�ɞ�MK&H�*�?�b/@4G�}�"E�HĶy�A�)�?��iV�O�'1�7-�ͦy�ߴM,���7$â��)�@Hm&�sJ�/�M#�'��Ȃ�>�P����EC�I�?e�-`��`�g�#���30�!1���IΟ�����	�l�	l�'9�jp�c�͡H��\`�lJ�\Z1����?��)���\�����'*V7�+��G-9p@`�[;��A ��>6z�$��m���MC�'uE��4�yb�'9rL��k]_踝8V	�%zU�T�Ç5\����	�c��'�������I����	���এ�[�ك��Q)r>Q��ǟ��'��7�:=c6���O��$�|�oЉS�Zæݣ~(�rCm	g~��>q`�i��7�v�i>��4l'f���'�>0��!T�;���J�q��$��Ziyr�OqΩ���k��'E6����#y@�-P�@���	ş��I�4�)��yr!fӖ�
�')ވ�(R*[�>0H�m���h���ON�nZE�N����M� *D�WŒ�x�	oXXU[���F��v��O��#�i���OVv�͊�U-�<��HI/=/&�dؗ�:e��T�<�+O8���O���O��D�OF�'U�ܔ�E�ٴ1d��#d�p0�7�iI$�w�'��'��O�2�x��.�$�&���D^�f)��m�|ߒMnڼ�M���x�O����OC�t�w�i�� [^�r�ڬ3��հP"G-��D+.q���'p�'��Iܟ���8|d<�Y�A_���q̂�v�M��ڟ ��Ɵ0�'8B7��Mi>���O��d�G�湘1��Ă���%O�E��C�O��lZ��M��x�醿�&���Ωflx|9K[:�y��'��`�_x5���@]����}G������-�~�X�#�#�F��]��˟�������I�D�4�'!���EE��ff ��΀(l<�H��'�7��$ ����O4Io�A�Ӽ�%m�`��	T.TVe�AP�&��<	��'�V�l�\(��&g���I�:�5^�d&� �@"E�Hc֡��A�|�dس�!(�$�<��?����?��? gX8BzX���1�Jl��M��D ܦ�HB����	ߟX�
��8x����4�d���(�M��	��hoZ���?]�S�?��c��+��Sc��[z4\�vÐX����"`�hy2eZ]��cE���y�8�Zv��5<zA�cCV�?X �[=z��aF� �X��E�?�ybLŕ7V��& ]�X�ׂ�,��'�X��l(g�*�̭�P)R�*Rܾ�`2g��y���A �m�R�����"�������4H�0V���3n��U�2����Y��q1r��<;�NH�5Ț9c�Đ��@,��pJe�5�)SǡI	4�����c�6�@Rd�AhpL��f̵4�2ؓ��َ@F��	�!X�!�-٫Q��2�HY�V��?������?���)����,���nIw�h !d�	P��aQ�\�IßP�	Ly"J܅Ȃ����L��4��4������̦m��e�ϟh�I;"�\��c��\gH��4��,�>�q1��k(��'��U�D��I��'�?��'Tg��cӨ.,j����E8C����x��'��4a��|�џ��(��і@�=ࣚLu|)��i�剱&����۴��d�O��	Y]}Zc���Г�ɻF����LZ*F���ߴ�?q��{ؼ���?�����5V�ȍ6���!C^lh������M��̕ ��&�'�r�'B���>Y/ODd ��5�M��	K�b�@�����K��d��ӟ\��F�П(�	 ]�1��%�Nʨ��&���B��ߦ��Iڟ���My���O���?y�'�ԑ���qWȕ���?m����4�?���?��-�"|a�S������\�'5�8�٧�\����Y!��J��0m�܂�ŕ��ē�?������� $�j�Z�HWN�cJN�1�Iw}�ԤbR������$?Ţ"����Y�$Iب[��rӆ�d�
-��}��'��'���'�b����3e�J�����<�2E2V��������Xy"��@�v��-7�~	�q�T� ��c���%+>R��?������?��z8����B����闫�2yy!��_~��X�L�	͟(��@yr���/�"�'�?��	T�xN0�h٫%��I����nz��'����p�'�Y4T>M��&'��Q�7�.x:B��֦�1k���
ܴ�?i���?!�Q~��_?��I���|�v��a�D��9:��F;Y�~dèO���<q�,����	�O��D�?��-Հk޶�x�&\��:�mӼ���OM����ߦ��'���O����p��_�\A��Fϒ�)	s�Eئ����,��Ş柌������^�S���ڱlU_n>5S�l]�jh���4@�d��Իi���'g��Ox|O�)Վ
��ЈΟ[����"Z���n�%M5Dm�	�@����h�S]�]>��EM��f04��u�7�����M#��?i�dϜ��*O�Sb�č�8�E
�"������� ���>T.�y�'���OjY�	NP�֬C��ʫB���iz�u	����)-�IH��U�Qc�|�s��N��h�4�?���O�'��Q���	3�r�"�U�
��`�1��A �.���O4�$)��Ɵ(�IXp�#a�J���뱇�(���	@+x��?�.O����D����:X�����t cB�	ae*7��OX��:�I�H�ɹ
���g��-;�,��[�<Hҏͱ+\1&�h��Wy��'��@�Q>����e�Am���KgJ�X�^��۴��'���'��s�|�B���>�R��0��-ST���6��Ol���<Y��A4�O42��5&�й6��5�& k��Ӌ��ē��]+N���*�)�?�%#�8N�(�Be��V� 0��)�>A�N�"����?A���?������&�I ��d�hh;7�S�u��)��i��'f,ል���Lrn9�CH^ L��<#5���-��l�g�7��OJ���OL�	a�i>��p���s2*4� ���Q������9�M��C�?���?!��b.��D�<
x�ㆅ,7L����@Ȥ�� ����U�<q�O�Z\��#P!Xj\�0Af�O��|PţA<�1coϡ	z�a�6F
_=ba&:�ެ�a��uWLQ��$X���lȯB����D K2؃0����v��J��z�
<H
�����,`���yaf͢MXY B'W�a��|b��
�r�\:�a��)�]���N��� '�H3_�����^�2.ұ�T��O��$�O��ɻ2�����O��:\JP��btBAi�$� ���9�,�C�d!$� �'|�,!pj�SDН!��T���4̀%l��!+T�^�I�c8�����Oz}m�Hb\tq��.dQ�0r@�^�6D<U�ܴ��'�"#}�H�,�M��f������f�ȓ1��Y��o�%Ҿ�*�-47t�����Gy"�.6��O�Ī|��
ǃ��$b@N�:���a@�=���?��t���T�D�C�f�=I-S)�.!붢��a��[�*ף֐����	)@H����$S�� s�?-���%NUR4,\� ���Ŝ�1��<��ğ,��_�П8�R�N&" �H�P"^�z,ʀ+�џ$�?E��'���ʠ��3C�\	� 
&+z�(�{��'��Z5E6k;pu��H0�V�0�'�2��#w�����O ˧i��ؠ���?���T��āLe(����	�^�;��Ȓ{T ��^*�"�S������ >��P���p��Be2l�)�:8�x��ㆾodFyY�O?�d#u�6Q�@��	&V��DЎBCv,r���O�b�"~�Iw�8\3U��!@B������}�C�I;W�FI: �#A�X1��	�l"<�V�)��M�x��qSkG�C��`Ю�G�<�c,ÎyLP�r!F�N��(��n�<a�k9}?=!�iX�fׂ%�YU�<��lN'Uj�p�g���R�Q�<�2��?JVx��턍@Ju���Ka�<��iH$�z4�0o��S%����+Nt�<��)��.E�u
�$0�E�`�Et�<ɔ��J��r5J�#nL���f�h�<Q�m��G��B!+\�X`��v�e�<�D��V�L`ҵH@J�`ɺ�ƞc�<���7;��"��\d6Y2�c]z�<�Ņ�;6����1m�����a�<�E͘49���4�0"���iEK^�<��H5	��g� ���"J�V�<yӁƗ)b�@aW�S(��Y�c�H�<!�NE5uhr��f��䨚f��C�<)�
	����kR����~�<q�)�$�f�y֮��D���7~�<��Μ?kLB��	Ěr̛O�~�<�Ej�:=1����Lޮ!�2��/�O�<�����f� ���^N\-�5.WW�<�ΞJ�2A�g@ $�t(�HX�<�F�e�0a�O7=����K�<�G)�pT�pf
�`y"�[�hc�<Q��RHZ�Q�#��+&9����]�<�6�ӝM>8ˀ,öe�r� S[�<�H�Fv8MP��߹I�$�:���a�<���U��
�P�o�0|j\�a.[�<�шP5?����M�=���q�,U�<�0C-̼����>@%�- �f�x�<�"��w�^�#�6/t��L�<y�	T�O:�/[rlX�dE�<�/�*Y �HQg�^ШP��g�<��I����P��+���E�e�<� 'H	B�Π)��X�P�x@v��I�<9c��e+v�Ѥ��&9�H��H�<�򎃰BwjXӦ� �L�Ju�B�<�"gN1��]�0IɞN�08�`��A�<�Ь؋9��9�S���QBA �A�<�D�
5R���$��}�9`C�{�<��Ȋ'�n��HZ�N}�G�k�<�"�A?y�&�)d��97�\�cc�f�<)dnȅ�3� 8\�h�aB�X�<ɇ���H9�v�M�39r��3U"O��Pӧ=-� @'\+����"O�!!⤄�pr�D��?p�0<IW"O��Y�A�
q��e����[�tQ��"O�p	Vd�.+o2�I�`��*]9�"OV�P�'��fx�p'}*���"O1$n�0a������hz� �"O �Tˑ�B�6�q�L]�h�B�"O�|�c"=o��p�DZS}�D@"O%!��Z��|qP�6 �8��"O6�G	%��D�OB��Ҧ��Z"C�hӱI�����8$�^�Ct���%�����"O�D@w&�(R0�ɀ��ίV ���"X$4�r� ��<A�+�@���d&�̌S�N�� *(9Z��0	�!�B�xh�$�d��oqTp�G��"#� ��.Y2�p�O5|Op*��6:]D�{ ��R�J�3&�'b�㪄�Rj�����,ֺ$�JG���{A��.N�4���S�? �4����(G�HdCN��p���^1D&�q���]^N,�}��&l�nZ'!�O4��J��C�<ɵ�E�{��� gM�,zQ:!�^��^�SC�.��䔠;!>�O�,T`Ѕ�Y������<Z|ࠆ�1 F��D+Z�	[�HK�C��h=4�ԙ�횔��=� �*j��pQ�Ə�P��p�A`�eX���"��0��M$H�-
Oߛ����yҢA�,8QS"�x��)��ȇ�HO>�kըH6�h��`�6��ND�����?z8��"O�i@Ƃ�1f�:T�`o��D=�U!�iHX1¤Fg�S��M�mƖv�l�jf�Xa�J��3�o�<y-ƈK�R!�Oi�NРw)����"1{�����m��D蓎�(}y8�ڄ썬!$4�k��,lO���1���?���/� ���t,��R\RҡL"{��
L���
���=�Ь�'nhژ�D�9i��>�cF��0$2	��S�>��矄 �'�>l)�O������=d���[�'&ĵӶjD��:����*b��`�`JL-+FE�$����9-4�!�D�	���K� VӢ���M(��OX]؟�·�Av�l1�iӿ������V�g~�ߴ��m�f|S�h�ܯrc���f�Æ?�f��1i)��a �&*V&o�c%�%lQ���!"bDc��.q�R�[��O و�55x�ru��{��$���H_:QP��7Wڀ��"6<O�X�U� �t��cмlr��G�O ��^�d�'ǈ:���( �O��2#�,tРe!N1!6I����z�A:�`��S����'a
�S��ͮX,�l�t%�T,���Uy����O�)�f	�PEd���jOv�6`8 ��"�a�;Y�DKZ4e�� %�Y*U��I�
U�:`�Z��~��Q'�8yĉ��镭ex,�H��8=5b���C��H^�X��J�T{~��U/�(x�ĒO��p ��?1�z�`�ؾ(�$@�T��.G@��W�G�Mƌ��G4	��S09X���$J8L���çB$�0����M�"���E�
�����σs�~V#=S����-[�Hz�ɐz��FN=,YZE����?�0ja��.��_�N��cZ�o�U $卖'��<+5OW4��xR-�p���d��v Y+e���QU��3��A�Hj�Ot����	6p6�~�72�`E[�O&$�����J""�&�˄"O���L��`��DY��Ι~��#�i��il�Ɵ�;�ȟY}D�� {�E[����?�
����[�$\#!`�0(a{b#��+�m���?���ԇ���8�����	R�HD_h<1v$Y;Ө������R!�D�1�*��d�X�6��PA����b�R��U����%쓾\!���r���B�x>��թ�V��A�T��=E�ܴ'Z��K��D��1�o�.56R8��NP���Ց1�l��u��#����'/���`��O����@��0��N'<�$�:d?�O`H�q��?��a��BP��FZ�\T�M�cĉz�<�4	�&����&%�F)*40c�l�'�d|��Qs�O/�đ��S����G�m���s�'P�H�r�U�/\���m���v�C�4I��H��;�)��]А�Gt Ei���т$�A6D�T
�W�"֊�i@���=`x��'��>�R�^#J�\��d��]���kg��:�����a}b�+(��,��8Î��S���IB��t E%6XC�ɐV��8�e2s  2U��y#=!4`X���}��	.oԀ}���?m�P
U�`�<��K֕'N��f%R�Fv��@�Ʀɸ���WPqO?7M�,�����J1&`�oî7Z!��e>�d�c���z� @�`ʂ/C�%��l��w��+N��t��E�*$B�ɒ,���#�Yt����A�"�B�I?̱c��J���{��߈3�B��3�/�:c���1���J��B�IB�4ѩqJ�5+n��(��L	#Z�B�I%8ͮ͛�K�~�T��#��k��B�|rRe��V�1\��vN�%ƀB��;/L���d�"zN^u���ԈwC�I�'�h��MW%s�Z��@��Y��B��$$�z�$=(�(EQ`BѧcdC�)� �P��/D��[A����ne�d"O��#w.lh�1��1.ڈ�F"Opݨ3��0����@��x�xe�"OT$���\kp(� C�<u@�(1"O&i��=fBlIWm?	S$	x�"O� E�Bv���"�+�$�@��"O��"1>�$�8 ����5"OX�B�뙴=<������? �����"OTܻ��H�|? 9Qj�>�|p(�"O��Z�)r|�$��q�8��E"O�Z���;	��bS��1X*K��y�ᓴ6���%�лYMxp�Q�*�y�J�~�����m�6I�,y!E�y�'0r���-�yTu������y�]����������BǄ;�y�l���N��c��Z���HՀN��y����d��mN"^-�p�dc��y�)A�eJ��ʱH�U������&�y�b�z�)B�ĵ�R�P�Զ�yb'� �����ޛ
̺�p�.V��y��Y�:�lYZ��<D��e�?�y�c<M)4�P��T���M��$�y��h�A���k��i�FA,�yR(V�H@����L(EŎ��y"MÍ4�8���U5X>�Ĳ����ybJ�2428�aU6!�~�r7���y���HIpT����.�Y�H�yr�̽%�4�v�$;�i+q�ۦ�yb��	Mq��������"!���y�-ĩ���#qG��{�T������y����vZ4U
�I߫g2��S �Ձ�yrm��gIb�[ (�)�2LP�<�y�	�<ך�@�lF�@!! �>�yR.D��P��C%&}�WJ܁�y�
�/��Xc@
��IJl�1W�ח�y���yx��*s��j��#��܉�y�Q�>x�� �2�jh��S�y�"|#�UbA��,.Q`KF�נ�y�BV�zE
dI'�G5�f �_�y��Жz!V��&1��yr���y�l��|z����O�9$�R=22Ɩ��yR��*o��Z�L�gix��hW�y�k�[���k�&��NH�2
�<2�'� Yd�e�("�J���dx��'���S$�'A/����CP�6v�D��'t��i!�8>"q(��3%��[�'�zu��3���{�E�90�'����%?�V�
���t�)K�'��1�%O�5*�uP�*�F��a�'$�yc�'�%1"���G�J�@���'������\�yC��ASА�'�D� �h�< _x�1�!%_0E��'�LA�*��h��4)QnϤ���!�'�^5� jÜ+/�q�7d��l'�]��'�I�6��;Q��`�#�ΐ����'�Y	��W�T�z�j���	�pM��'�\t+��Ai=s���J=��'��-k���8�ʠ�&ް�e�
�',f��$�-B@q�D�� |. ��'�fĹ!��c�pA9�&U�'�s�'����!C�ڰ��ME�l=$�')�`���=O�&���T�0���
�'.��2�H�3��ݐ��
q���
�'h4��t��n�l�CP8 �e�
��� ���/Z��PyP�D�-3OT�@"O,�C���U4=@�M[�hKJ}˓"O. �ҁ^E:	:���P���x�"O������0�	ũd��6"O��Sp拟E�6�K`!_�iZ��"Ob�do ;5�����M(V_hu�"O���ヌ�m�R�k��UDX!"O@Q�gʗ#���	!`�.j&ZA"Op8U ��"hԐ��n=r�e��"Oy!@�C@�md�	�(�"Oؘ��A�2L!�Ɉ�!l,�̡e"O�i�f��p;����L���"O<��V@�ynle(���[ �00"O����i�.|4��@�w�Dz�"O�qYQ��D��d�@ZSy�}�"O��`ϟ%-ø��5h٫�~+C"O��S��)�<+�E�>	S��I�"O"A���Chw�_B�:��]�a�!�H��"��d��0:84�ʠ�@��!���64Ԋ=*v` 0dpP`%hɓi�!�� E��#���3�ّ!�%z�!� ]��a&AƐؽ
��|�!�Dլ}�����X6�t���fZ�Fw!�D��l����.ڏv�v��w+�@�!�dª#�N�NQ�)�'--L�1�ȓ9`Ha��o9�ʰoR!LIv���D܈`A1D�?��	�5Ɣ(&�|��_�� r�ոr　��C�.�х�HPJL��)$J��M��D#����G:}��j��o#�!���I.ɤ��ȓ!�������r0��!��L���5*(�0��'\�6D�^���ȓH_�d��eH�*�qB�Ҍ\~*	��Q��P;%n�=K��Q���		���ȓ;�>,� ]X�`���b���ȓf<FX�`�L0[ݮ\��a�)3�P �ȓYt���J�jo�p�ŋL)P|���;�L��t���T�<bEdH�;���YX��12j7zd���T���������58J�(GZ�dQ:T�ȓHG>L� j��/g�x t�K�&y\]�ȓ,f8��&���qפL E��\�Ѕ�s���J���Swn!�3*�;]�̅ȓ<��h�D 1��0g�
�+�4E��#p ��ྀ����_-4��q�0ܚ�̙�z��'KK6&�����z�R%;�)�H�	�J�9�> �ȓ	 h���X�*����5&�\ݹ�"O45D�U�~��p��#	.!� "Od��U�Z�Op4u�D��T�0hQ"O~�`D�]�1�i;�e��PQ���w"O��[
��%z㉏7N�Z�"O�����)a60j�\?��v"O~��H�/9lx��}&*���"O���УO?�6}���0`���h�"O�p��AV� ~U�S� �Ӵ"O�QP�Ĺ
�z�&ʁ1Bk@�cC"O6Y!��X0a���)��
���#"O|l���kX�iFL7�0�A"O.k��3O��F�~�9dˀ��yr�\@¡Q��r��cC���y���R�.���C�oz��2�.�y덌\%zu̘t��K���y��  �6M�A�Mz�&���y
� �	�\iX�S�$:��X"O��m�/'l�#J0h�k#"O�[�	�*���$�9 j��"O���S�25�D���E��e�4"O�L�v���m� !��n�m�j�j�"Oq����&)���	�w�����"O��r�$�A$��aB>a��:u"O��2�*[��U�C Ů��`Y"O����KU�x|�y#�l��&��G"O�T#���l=�q�ށ��C�"O���#Ԋ+�\)4��X��,��"Ol��F�.�S��Ѕ��Q��"O�!J��f0��@D���	����""O�H�3hΰ�z�C�	�%s�U�"Oj�1h;!��h ��td��Y""O��S�d���pt�� ;4�)�"O 0@�K��h�
�^|8�"O�x"�L��M2�)1Hd)X"O@dԥ@-U��$R��Χd�j�*C"O��c��I�~�$�2��^�^���2#"O8臎��[4�1�(Y2GؙsG"Or����P���щǉX/���"O(8�*�.'�M��.�y�œ�"O���-A���@���0=����K�Z����e1e�4�����y2�Ύ-{�L�-�_���Y7!�/�y�O�3�Z�"��֓KV��F���y��5���i$kS���8�ķ�y�EʾG�(��c�T$7�������(�y��N5�����
5�$]r���2?���߀3�<��Dб'N���W+s!�;vOȀjRc1yJ�-�I_-`!���=m�|�"�ѧK����JϨ`U!�D�8�|��'��!Ւ �5�1�!�O�6��P��?r^p=F�6>�!򤎂.v��S%�ކ��M����g�!�dǨb0HL��wFB�bq��!Z�!�d�a����!��{D��&�+0�!�D�oR,�ġ�D��@l !�!��ĥ�B�ЌƄ'.z�z��6>j!��jNz8��?9�	�F�N,\�!��<M. s�C;,s�A,!�$�1bY��7��3�|�(�%N�!�DR?z񚜩D	!�&I�ED��铋�>9��7]���bKY�C<I��V�<�@�قlމz��J�Ql�� p�U�<��ޯ����"GV@(6k�h�<��'U	s�`Q�$Z����zg�P�<Y7#�e+4����M�6����ƀ�a�<���0O<�����]���Y�%�_�<1� @�;���5%
1w�V�I�@�<q��?x9 E�(���{R�Lu�<��B�S�T �v�57�<hA�\H�<q�ŸG)���DO�:��{��GY�<���	t�x1�PI�8:���	�A]y�<q�!G|� -�@D�e20��nBt�<	�e�p)J��&{���A�T�<���O5<w~�s��7t�Y�<���@W�0C�f�>�P��X�<ɐ�:=��s�Ɇ�}ܸ��!�U�<y,:D�h�($�J�|�4��"jZV�<��(ԁ"�8&[64VЛ�iIV�<�tn�6���H������H�b�j�<�S*ݒ)�|`�m�&R����O�O�<� �j
Me��sFO�?���P"O$�%n�=f��H�v-�p%�Xx�"O�T{B�u�
ɪ���0��H�"O�(�wρ�{� �s���.)�:ː"O8m��H��]AQM�,Z�c"OR �����s�F�����05�"O���mA-IQ�P)�H�	 w����"O�j��1����M�prh�ѵ"OBp���&�v%�v��%����"OxyҍW�F�}�f�,;�^!
F"O@ Z�"�<B�R���)0p��hB�"O�p���SŘ�GE�j��T��"O�1��2��L���F�Z�R((U"O�e����ob�0ui-r�����"O�S�LW�R�FU�E�6 V���a"O�c��/����T��pA�p�2"O^T�O�:IJ�$C,e4Ȁ
5"O`M#�O�g�&�A�-!�03Q"Ot�NՁg�؁����\���"O y��IJ@!�@�I}�m""O�Uy�b\��D����p�$0��"ON�IQB�$��5��F�p���в"O���$��*�x�7���@��Њ�"OԜ��$ͻG\�H���C/X<["O&��p��&*���c��&H��!7"O�lhB�2Ily[�0=i�0"Oj�'�\p��q/�8��1"On�+4"=s��Xc�O؞@�� ��"O(,b�5r8I���/L����e"O��9ख<��L�� w�� h�"Or�������p0�c��n(41p"ONkdm�> :v z#��&T�Y#"O@E)�o�_�B���5�]�F"O�h��l4d�I�CĠx�b�x�"O�iS`�Ĩ5$Ճ�/�=Wخ�""O�ܹ5dÓ\ N�H�oʮm���U"O�HR �Y#��� �<��x�S"O~���#x�a;�M�����Q�"O� ��N�7D�l[tb
<j�ڝ�e"OԠ 𯍈9/,Y [{H�1q7"O8{�+�[��hh�nR�42M��"O�l�D��Y��ȓM�%(���"O ܃nGy�ԄH��ȵ/ȌZ�"O�aht���N}���X�f+~��"O����1ຍ��( �mw�]�"O8�*�A�EgT�@�"&Ԩ�R�"OȄrB)9��c�L�d��5c"O@�Bt�;\1@�f���az"OʨP����bZL(�+,Hfy g"O�0�G�x(��@�%"�^�3�"O�u1��_���Ţ��)��p$"O�5K��c������P�"O��e(�#L2���N�N6���d"O^�3���9 $�`���W ,��t"OL�;�B�5idApb�Ûn $i��"O0	+Ԁ�39��8Ї/y����"Odms�&&w�@���+T��`�C"O.t EI).<Axw�ٝ8���B'"Oxf�[.|�����F�:��`"O8�'�]/�ę� �&<��e"O�t[#Gú8k�M�� �~-�%��"O��x�g�8:�K���?>M��r�"O� *�&�}Ƃ�PqA��>��%Y�"Oz:�O�vVH��`J���7�!D�� �=ȷ-7�꭛p�ՓjynQ�5"O������ %<p����RS�� �"OXm ���0)z��ː�b��w"OFdH��	F1V<zb�$t���:�"OT`9ti
�3Cb��Yyx�
�,TK�<a��K3C��iq�$F�b}:��Z^�<)D�յ	4����\_�H��\V�<9L�"]T���/��~E:�b�U�<�u`�Q�Hdh$��5\h
��J�f�<��Z�a�l5���ڱ>�@}�BnW]�<)�oP�SG�hCb��+/F�x	w�U�<���m�F�Y���(0 E�か]�<9-��|�~�1E�)C\���X�<)TE�C�$X��%atU�נV�<��4gT����·5(.��c��P�<i �޹Tk��à%XN �*��U�<Yĩ[,�p��Q��T'��Bvl\m�<yk%7��-k��{M�t2"��h�<i�jH�*GR|��g^N�\b��d�<�D(wW�I 'nD-GmA��`�<�թ_6Q�1S��:��R�PZ�<�r��&�Z���� ?����X�<�r�	�'F^i���ض^�tR��\�<)��V|�
@pDն�,�1�RV�<飥�6C�D�@� �7N���#O]U�<�ق4!�����ݎ.�2@�	K�<�##��"D�8��Ң �ޭ�"�b�<YDg[�l�� Ab
�d<J���HLt�<�Ӡ�J$�i��U�8�.����m�<Qb!ӫ>������:8S uD�i�<a�nO�)�x�Ƴ&���R��o�<���7���k8|�sqH�l�<AɓUʄY���X3S(���l�<!7�
�]��e\2�
�DcTs�<�4��@ px0ϛ�+>�y���T�<)�U&Q��#�V+j�8 �J�O�<��*2Rt�Fd��"��'��@�<Y��$ia~�C��V#]�B�x$�E�<��d�<� }c�S![ڸu�0��D�<��-ݿ'���"�*����g�I�<��D�~5ѥ,;��@ `��{�<QAH�k�젡Ѫ�Uа��F�x�<ᖅ�/���
R�R���A��\�<�R#W�~B������{�Q@�Ls�<���V��]�	����!��k�<�)ب~$^�ȕ�� � y��h�<!�L��K��"3��(<E�̠��Tl�<�qG�e"�`anD%Qs�i�`	h�<�A	�<ѨՓ���|]�����c�<����p�"����jA/_�<��KO/jԁ�EN�o�.LR�VB�<�.]"7�(�pwH�	k�|��#Wz�<yg��m $$���ɺ;_�����N�<��ī#�4!�/ K���`�e�<��`\���<�Q	�'�r����[�<U��v�ȳ���+�R���b�<�w$,X,B��eg$�����`�<a6�	(*8<��^w���Ob�<�A�uR��bc�={���b�c�^�<��7I�)���R�E��$ip�LO�<�F�0K�D0�Ve���M�s&E�<!	��\|��]ú0y���~�<d��.�u���	neDiK!��x�<��
f&� ���P>k�BT;�.�v�<� @ȳ?3��mɃ/G����w"O^Q@,
��¦�D�5��0�S"O��a�gĲSe����mQ�Μ�"O� 8���<�� ��L݁f�8���"O�Y��� J!"AQ@��$���!�"ODj�D]�*�<9!����� "OXL�2��G��`�%��.���yu"O�5d���I�SaA/u���҄"O�99����3Vh�!A�6P{L\�"O�5�B�<U:�Ej4����<@�v"O8�1�NH��Е�5Ϙ;�x��"Oн����"b��X��M��a�,�'"O�<�B≛n~����Ѽ2Ym�"O|k"�V [��	��ȧnG`�IR"Oj!X�G=ƅEo�Q����f�!�F�$�0s��p�����֭=�!��R�q�<�@�T#���Y`��J�!�Ưa�Z�B4jH.lGr���.�(�!���sy�d��br� ���=�Py��<�J���{#4L���
�yrOϖe/��udȔ\s>��� ��yR��/���D�?j^lZ�ݸ�y�a��y�>tqL�<��4�Һ�y�)��[&h9�#݀7f(�$�߬�yB L�B���C�m�85t��$��&�yf9jX�J���'�Ʊ[gm�/�y/�b25�d��' \���y��%_EB���L��Ip�W��ybe�2�B����f�ADĜ�y��H�`x�ЄZ1U��2����y2��*��������p�ai[!�y��G4ά��y�RE���y�Nϻ�\%1�D���gʟQ<�a��1�J&#�At٪�L"�2��x|��*0��@Nv��&��J�Ѕ�]�=�E	�#y+�򥤟�rzP4�ȓr�ҒOr�| k4��	�T��f0:A�5'·.����i��Y��`3�4��탮d�leRqQ�m��f=��v��	�tz�i���d��$�p�׏�/k��%��-?���ȓ�,T�n�?G8�г%
[&!Q|ԇ��>�a�K�-�j��U��%.��	�ȓ#�X�@�O��~P>dS�f	�B��{�<a:? �t[�s,� �c�v�<�0n��i��|�a(T{��P�&�v�<!P$N$F�f�[�'�w����.�s�<	7�Y
���Qe�CI�!�Sr�<���ى@�A�a �?Bg��Yd��p�<��F�-@!�	Z�(�?��;�"�i�<i�@�<��T�@�N�v	�ELd�<���F���E�,�X2D�\�<1Ў�&><$1�E�+3LP�iU(Z�<�ԃ%!<�R�*�)dqfѱ��U�<	'�Ҕ44������:r��P�<�}޼�b���� .8��3�O�<�AI���}ӡ,7CJt��⢁K�<q@ʂc�pgF�(FXdL��l�J�<���ѤsH���%�� dm�E�<QQj���� ,Y�cf|�U,�C�<��IJ�?����Ǟ&5��V	�A�<i#Ϗ+��Ģ��Z0�y��\@�<)uD�g��z�NB�xzd���[V�<A���@��Ё��D0&����	�R�<� ���N�T�#�aO=�vAw"O����b�&Y1h��@��EmL�"O����(��p�4��e��BĶu�"OD�����`(C�Q�A�,@�'"Ot(� +I,���s�\a8,QV"O��f�K�y��4z��G�l3�ɱt"OZ��M�5���ê��N�8��B"O��zE��/n�R"��;^\��A"O��a�M����(I pY����"O0��� �$7KZK߱�P��"O�M�:!��Q�]L]�"OB��1��IN�(Q�!�f�8��"O����ŚW1�rP��6W�2�"Op�g@y���K�*��"O�S.�,p��1ʘm�"O���@HHtŤI��i�S����c"O(���) >�X��Ņ�9��h�0"On�j�V
X�Ve�`�	w����"O^!!"*��sV ʔd���"OD�:T�Χ3wJd�r�_7?PL�ۀ"O�5�2&	�4k�Uk���(]N��;�"OX���-U(�TI����VU�H["O.�I��Qj��P�ޕBG���7"O�=�І��4�dh�b��#>X�#�"O����^=J�I�w��j0�HkD"O���5Ώ��b�Y%J^44�acT"O~�j�Lߒ8A�0AHә:m��J�"O
u�G'�F���@A_d�&"O��7��O����؅0^��ڂ"O�Iɥ�F� .DJ6��Od� �"O�ѕ��{��Т�ũE/��R�"O��ч�p�9�fL��E�����"OС�H
�I�B�r4J����"O,���7x�A2�j��"m��6"O�$!�&�� ��1 �HL�DNL�sQ"O.��*ËQT��b�ը4/&�"OFL��#K=Z� }X6�O�f.�$�"O�@4�\bȶ�Dn��{�u�P"O�ź2(�j��pM*n�T�j"OԙѠ "Z�P�W�����*ODa�U�
�2�n�r�ꕱj?r�[
�'N�D"ƌĲ(Ĝz6o×cD8�
�'�4�Ia�`�vu;'��$b�H=��'5��A�(�m�n���&U¢�{�'��r�/ަ'pDp��O*��	�'�v�%��=9|�10QA[QX��'}&�ꃏۊm\H;�ؿ�NI��'��I�cɍ5id�b�H]�nnT�����?��T]>�ۢC[�(�,�{��3���#�YJ�<9�iV�c5.���_&H�0�@��B�<��jO5b��`h\$ U*Y2���z�<ׅ	.h����J�k��TB��y�<�g��6���E� "?��[�a[r�<�Ӥ?5ΚA��o�F�@�sbbl�<9�ǥJ��Ă�%Ղr��4�i�<��
ҡ	~LS�)� ��4���c�<i�b̪JZ�st�N<��%a�cN_�<	�-�R�� �8G���bBRQ�<I�	�u`�i����/�|��g^N�<����$Udb��0�ЖG��+6�H�<��I�^ �� �3���A-�E�<Yj�5&��q��Fz
�#�f��xG{���%_A�р��ڝ
q%) m\=uAC�	?S��A�V��9�C��	ʾB�)� :%��.�-!g@?�` 0"Ope�!��!l�dy8�e�%6��P�"OJ@X�d9>;$E1���=BQQx!"OA
�(�8~�-�C��D�l�P�"O�����ho���,V�W?������O����OpL5��-A;�B�%�Εb{��	�'"��&�=Ebh�1�"�=`���
�'-6���`���H�^"mꨈC
�',��LD�#y���qJ�0����'
<h �<^)L$Q�32=�eI�'�&�u��vi���Q�� U*����'q��e�ME��Ia2��#z����'�]3g��O���1m�g�����'�p ��B�F(푶LԮ	���
�'V�d���Uc�-�)l�8p
�'�R���ͩ���Ӷ/����
�'Q�`�C�O�ж�ۊ�J�	�'��u����� �v�}x	�'�4��S,,�D��叕�+�y��'�� $b��W�`� ķn��D�
�'��I�녕~Q��!�Q�BLT{�'T& 8C���l���,	5t
���'�8�ue�8v}EQ�k4� ���'>�K Ր%ج3VfS(xP��'�e�A������ 'i�$R�'���H�!��ܥ �ƙ]%@��'t�0SQG&�zĈ� Q��M*�'��e��!��F
(4�oE\O��3
�'�z`��M[�a#@�#~v�� 	�''B�EE5F��ivM �}��k�'���c��� �T�Uf�v:�@Z�'�1*�
�I}��넅ݥn��MR�'����\FH��F�YD���'|������+m�1:oΛٸl��'n>5 ��U0j:���ÝFt`�'PH��$C�1i�Ƒ`0��������'�B���8�Du� �	�K�z%1	�'	����l�;��p ��!B���`�'vB}�ōØT0�Y�׋�=�2u��'��(A@V3,��"�
�Ah�0�'$e �
���r�K7mBu��'�,�A9]T�E�P���"6�K�',��S�D1^� ��G�^��@x��'T0h���٢l�z0�ģ��dq��'����F��
0�d����
���'���c2�� s�|�a��/L��$B�'c����,Όjs��XD#�P�<��'��P�[�����_E6~I+�'Y��Eޡ`e�	�?%,���'������U"<�ʡ��]7����'��Y��*I���E��*+�A�<�dnݠ0�.�x�F0 ���"�|�<�����񰃡��>v�ip��z�<��h�04��M��	X�}K*@�3%[t��?�çe1����KY6D5�`%�P =yb\��&�����=@�ݸC-;U5����g��(�������s�6wLdهȓ{�V�Y��ш~H�����9Z2 �ȓ1�����HG��D9H�mӹ\���ȓD�m�dHT�v��-#p�ȓ+�rv戗U�L�F��b�,����r�q�L�B����d�I�,�zL�ȓ�� ��Q:Sa�����h$�T�ȓK�ƹAD��X�z�cWm�3Ę��S�? ����a�E������K$��Q�"O���&MOa)�}C�� �:��C�"O�es6��<�J0x���;?�l��"O��`��\�po��@#�s��������O�����b� �a�J�ooR5ѫ^)7�ў���	*S\��S:β����,̒B�I/l�d[Si�~BlxI'^�ZhB�I�&�xH���a �\6wRB��;�j`��&]2p52�fމ	�B�"��TC'C�F�d��f�9����$|�����	�X�F����P$�&�D�7D����
�5N:qiO�7�<I&k6D���g�	�����ͅA���Yn!D�@۶,6]~� �g�ˠ$���iF�>D�l�3�K�x.=P���#�Լ�u�<D��he"�\���i�:���6�,D�]5�0�	 N�@�h+�a��xFn��sj�:yt�[q��.9�	l��� ȁ7*�֐�A��O�Y�2�(��0�ObI��sP13�dR��<��"OĽ��U�2��q��b��3"O���F�so�E�bCɠ{�j���"O�4���ƍ#�L�:5+6�q"O W/�+oj|�3�*^�q2h��"O,<��`ͻjF��	 @�c悥Ґ"Ob��g*�Ӕ�Y�>E��d��P� ��ɂ��3�/��f�}��&2FA�C�	 j�bȚ��H�F�"@�$��%9�"On�0� �%*U<! �N;s��t2"OҬ�������EC�:��2"O�I�t�âku��ҁO� |aXd `Ov��t����ْ�ɘ,��бUI/D�l��G��f Y���IuK�T� �+D������2ps=XtG�?i�LI�!�*D���qᒗ%���CF��� �)D�,��،V+pA�4��1��Iɓ�(D�d�C<��У.��Mb��x�,%D����×�r��WA�	s����"D���"�7���;��3��qГ�+D�p[Q��:�|qّ-�a6���%��9�O�8Ȇ����b(�� Ưi>�y�"O0�q#N̽L��2�T�܎i��"OF�ʵ�ݿqވ8*S'�,0�B(��"O���¤R%���i�Ƃ7O�J��"O�XU�ơ(�@��$	1%�z}��"OB≃�;Vj$y$Ⓚ�4zE�B�0��G2k�v�a���*��,�g�#D�X@�쑚
rN��CdVV,�D�g�#D�H���g*�� �RK�`���.D�4�B�>#��Q.��`4@ D�0��bT!rڑ��@~��D�:D�d�Va�"Kfa��Q�Y���3�J9D��ꅫ�QI���G��\��Q�we7�O��¸ �BAZ}�&e*g��<Z ��Qz�,#ˋ���3�R�j�܇ȓ�l%�t��=;�\
�@6t��ćȓN�1Ir����L��	�aW�ɇ�CpF8�"F�6�l�	�C&'rZ��ȓ�!3A�6�aa����7�TE��
������	2�𐠂�53�0�ȓ!l�]PU%�r�(�2D�SL�ȓi���-�I�����耆ȓu�N����3g��8�H�sᨴ�ȓA��5Q��H�@\8<��	[�ơ��S�? ��j�
@<dSZ���* �c�"OΘ�D
|^tY�H�,�,�j0"O4A#$ă6�� B'D�M����"OJ�󲤈85T��z��0�2���"O<��r�\� �؀ oD�Ȃ��"O���2�ֺQ蘤JE��>7T�y��"O:	c�+B�&'4A�  \� h�"OL���.((�����!Y(œ�"ON��+NV@.4�S([P�[�"O4오��m����eݢ[m9�$"O�����F�̔8�d�����X6"O��A��Ɔ):�-Ag��݈l9g"Of���l�X'r����8]�|"O��%IB+1D2=�!�6 ��K`"O`�y��T#��C�f�IƠp�"O-��,Z�d�.l.L(��X�	!�$I!Rh�tS���:"w�L{���I��O��s��~��$X8�H_''���+0�H��y����C���[�Mуn�6qQ Ѷ�y¦�d����ҏ� ����)҆�y�S� iޠѴ!D��US��^,�y�E�V��p&E-z:�uR�!�	�y��CL��E��@��$B ���Ȗ�yB� �pM8��T.�Ή�D����?q���S��l���0�֡����_���C�]��"C�/����|�����`_��I�ȃ7���X��V�1M���ȓ�����I�[�ݠ���n����*���`ͽK�n�0�MF|��_���R	*4b$%+�X;x�-�?.O�#~�vm��s�!H��1��+�B\y��|��<� ��D��r���v�A�o&D�XhT��]E�IHrcA.	>%�%#D��[D��N�L,�d�/>�Ę�t�!D��� �M&b���P�^rrа���!D�x����,�v�!J�0\^@X��?D�T��[E�4�!��%)�"�K�<��Hy�^�d�O��	*ߠ�22�Q�Q�T u/T5�!�[�������}�A_j�!��U�h��0���D� ��K�;]!�$�*G_v�˗�۷.x�bu�-me!�0}`���C��]���腤)e!�$�1<��B֌i�Y��$~V!��ӲG�xI��Aӕ:D���7$
�T��O�ʓ��|�O�©!-%ͬ� "k�I
���'���Q��ˠDp{�엘?�v�q
�'�|d++I�!��߀?���y	�'	n�X�� ��q� L4�2�:	�'�*�Q%�-vn�(�E99�b�;�'a�qUd q0��W��!a����'��Y�@�f��f	�6f6V�C�r_��F�D΂�"5Х%P�jjL���B��y� ۖ:;4!�S��cXM���޼�y���-+�(���M*f{���&�
.�y��SM>�d��G�R9�U
ܠ�y�m��1t��p��B�l�9�G��y2��>!��Y��Ù/������$D���A�ID�hQjC�w)��5D�T��K_�q��Aץ=�8���4�O��m`���v�QF�j��"
�E� ��`K�u��A#� D���E�\]*̅�6��0` @�+��B�S�d=�ȓTR�[��'/�X�B���p��ȓC>�c��N��H����N%r�ه�S�? h���!��}z�|��cE�K�����"OL��BV� S�a���
pjt��Q�x�W�Qf�fC^�4�a!D�dk�ƻL��x�@C�*��9y1,!D�D�&��*Z=�&��T���S��4D� [�d�S&Y��c6�B��t�3D���h��<�N��с@,)l0��4D�\ ��� V�31¥~�����F0D�X�E:{�d!���z F!��.D���íյq���×�۲�l���-D� �ӡ�m3̡�A�ݒ�4���G*D� r���5"��f�@($T:tk�b3D��8���Z��r)ܤkf 3�;D����ȿ)��$3�N�;[P(�'D�h�)��80��"sF�
&����g'T��ʰ�C9|tIR'Z_j|@W�'
!��P�m{�L����Z���to�5�˟t��I�"��V�גXP�P� u�JC�I��\�q�+U�����- '$C�I1>����o��dn$L���ԟ* C����p�Ws���j,K�&C�	R��H"�
��O��pZ���Jg.B�0`�0��+^j��9����T�=�'�a~�L�$f�[QJ��)�N��H��$,�O��S @��*
�����U�M+��j�"OF�A@�?t�S�eB�o�X�!"O���a �$��Z�gAp�P�"O6<@�"S2f�Uc�%c�4�'"O��D��U=�E2��V&q��@"�'����Pm� �;nV(,`�W��!��V�qx̃Q��~�B�r"ڧ�O�����F�~���1�j}BQ@	1!�.��2g�5r��ĩ'χ0KT!�0S�pI�W�'��P�2�ËKE!�ąW�>h��F�v�*��L�,^'!�� �M���j�8$���w��(Wk!��\>|	�8���;�0С@��O!򤞢<� ͫ⣈�p��CT�V+RB!��RLŬ�XC#�?E��5X5靭e�!��8y�cuł��!��I�!�˳X����hE�x�~�P��W�d�!�$�;���
��Ңa����S,@}!��Б
�ҕ�$�Ƀ8#aaŎ�Zo!�D.z�2(H���6
2�JBE��	n!��ɖn�:����H;L브+cE�KY!�$S��p�P[�':ȍrg$�c�!�$���![�CÇʈ����%)�!��{��	H�-J(ds�d�M:a�!��[3k��!@$瀇xj���P��;>�!��*`��d���Fw�p�o��?�!�d�=�(�-�4MD��'�Ҵ�!�$E�k��'+�'8D6�3�K��!��1`��"/��J0:��I�sE!���FD��fL5�QCÄ�7~=!��[�B��6�R�{'��!C��(!��(c\Z]��nC�g$�q$� !���j��҆h\�&���O�!�D�(�8YG!���4�2	�+OB!�D���q��#A]�@L 榐�&!�dO:΂�pd��U�L��`Ɩ�p�!�(
��@������-�F%�S�!�D\s���c�^*K��M��j�p}!�X���=���>l�"|I�ۮ�!�P^���atOU�5|��ٗbm!�� Z�%]�D�$�Ae��	��H
�"O ���ʐhf�Q�0�3X �z�"O�5���b�L\��L?OVVTkT"O�հ@+G�.����_�w�\I�"O��9F ��Ȯ�0��+�
�s�"O���2��t���bAL6[�^���"O��D�	mD�3��6d��X�"O(X�Ag�3)�"<�Э�+۾�P�"O��Jw���4� �L�vg�C7"O����`�ͺU+�
ۜ �^P�"O��r \�r $��.j�N�P"O ��#�L,|��B ��T�3"O�h�'���f��䛙���3"O�x۞�����;Β�)ɦw!�D�cXp\hBN8�� �(�=�!�d�(|���Dfƻy�`y�D�t�!�&%�)H � �&��IP0�$�!�$��(�^	�6� �*�$#H�p�!�d�	.��aԧ5r ��Ţ+p!��rY���	2b��Q�o���!�d���L��c��m����[�Vj!��4$b`�S�K]�t�B"h!�$V=t���hEe�u�b[1O	�V7!��m+�̙Pwo�BŊh8	�o!����e���:�ٴԷt!� ��@ A7e�����+U!�d��lh2�F�;�b{���56E!�d'~�x�W3?���0q�	�U!�-�h%q�LӶ:}p�R�f��3$!�$�%`�,���?ǔH2�V:!�ЫV<*SH�4'��Y.a2���	�'����AN>Ә�e��i����'(��� ψF;�ah5� �n����'H,H8t蝍z�<���G(:%(Q�'���yUρ�\+:4k�C[�8I��C	�'� Q��H�,b��@�2D7�6��'�V�xAÚ�["��d��Rrq
�'���@w�^�^pܤ�4+K�
v��	�'x���' �D� M`g�I���(��'<�1��8}���S�"�+C���'����ۖ(��@R���)[0f�y�'#n�Qb�CO���ѕ��5>� ��'>��5$Ӌ,x��Q�=QΡ8�'}.�%kո	�"X�3��-u^���'�61a�*�O��a�5�7q���'r��P�@�(�Rd�[�f~E��'���u���Xc�6,J,���'�����'	.X M��	�v���'&��i�QC��Q�@��j��'�PԓWa�1l�j,����2uHT�'r@)5D�A�<��>���
�'h�Ds�"׭
��EJ�g��5�l8�
�'SZ�`dJ?b�jsf�-"h�
�'g0}�%�k~�t�R��o�
h�	�'l)��eB��HeG٤��H�'�HǣW� ��1��;$pY��'��]C����eܶI�6&�=g���
�'8��P!�O&LI*Ȩ�`�dj���yR���T���B�4�D�p�Ш�yb�'j��L�! �9&����H
�y2��7ąR֨��5[V�Z#�y�)��?����a��"2Ț�����yb �QM\�{�l�`� ���߱�y��K�Gj捉p	�
Y����fվ�y
� ����e5m�m�RB��v\����"O�d����Mw ��`Oy%@Qh�"Obph�^2v&|`/\0n~Q��"O��b"-��t��#X,dk.er@"O���߬7�p��!Z=hb��2"O���&��?r�(�g}]$�	�"O���6�?jt�4�:A�"O�\S��@�u&$�j�;6���"O�d��oO$v��)棎~銀�5"O0�H���4fXl�Z!�#]*�u0g"O
��O	l>�$��j�tD��"O8��w��uL��9������l�"Ox�F �%c�Qe$��J����5"O,U;c*ĶE�0I�S��#5.��g"Oa��k��3�^E���4l(�8�"O��m���p�/�&7x���"O"��F��O~Lyf�0�H� �"O���f���|?�	I���*�a�"OL��w���_����,@�S؀�i�"O���a��H��M �ˮ�Hi��"O̥s�C��7q
���L���"O�8ss�O48���HR�&�x��"O� �IPr��Y�D�
*h��S"O���+Q�^���P�Qm^)+"O�AAwES�!���P˼wW��r�"O�*���`�<�ҩ�+hZbu"O>(2��%R
v�XfoӖ=f�i��"O���рȣw���@�.�9dڽP�"O�m�PB4p|Ԕk�\�"4:��"Of��G�0�� K@0M�Y��"O����-�0�ZL�96"O`Ĉ�g���\\R0�T�Q7�)x"O ����E*%:���$��� @��R"O|m!e��Q�� ��� F *��"O�}�#ٴgb7n��`.&��"�%D���G @�$;���'L,e�� �*#D�`#���!o~f�0�gHo�Ĉ$�+D� Sp���
�dŤ()H2�N'D�LqmI� @����k�ր�ë$D��	�0-��x���Q��Y�&� D��p��J�cz�`���ډg��쳰�>D����O{d��`�$�(5� �g7D�����T` y��ϳ1n�+�*O��qP�'��T!��$-�X�(�"O�r��Fht�#%N�s�v6�?D��	&�M�{h^��`�/s�XQ�>D�H@��h:`؋@���!UF�� D� ��AR�"���R�l�-�@���+D���ǦP)���}6DLâ�'D�D!���ce !�.�#K� �E$1D���T��!x*��s��Ă<C*���!D����J�	W�v�� ��7k7b�x��>D�4����[��C�BrO^� �7D���FE$G��e;�.�4$-�X�7D�,cR2Y�`���L�L�)"�3D�P"�ˉ2y�MX6�HFȔBSb3D���J��m�Pԫ��5F���K'D��3���" �"��\
ؑ����/!�$S�)�Y`�	�[��x$!_!��U����t��/_>u[@E(�!�
>���:U��Uv�˲oO0(!�ރ"i<��Z�KD
��RH\��!�D��Z�c�b"5/X���a� 2�!�dF2(��m����E~p�S�s!�� ؅IrOB�Q�j��3o@�; J��T"O�h���
q�����B=_��Y5"O8IB��^o�L��0�T���*�"Ojy��NI9X�H�̋4�
X3"O X�Wjܔ2�P�
*54��"O|l9��w�x1�^~b9;&"OY{�K�7A輁�jO�#{��a"OR��2I�
^��9)d鉙7����"O�0�V#X>�p=PaiWX5Ӥ"O���#�
,������4^�̃"O�TYP I$4+,A�r�N�l�:X��"O��t�X�x�l��PNO6\�"��$"Of�C�<Jy	3���T�q"OR�:BO݋#H�*��2a��	�"O2�CԂ$�J]Õ�Kp����"O84p"jR�D�ي& �(R]X"O�LCT�\�u��aEY�%b��"O�xP���3Bf�gM���]2u"Ob� ��[
G4%�:N��v"O&�S��:k�<ıc���LG�A)�"O���$����p'MC�v\b�"O���S�M&z�j�b%��R5^�
"O\���9��85'K�3 �p�"OJ���#Ĳa����f؍8�X��"O�y V���[q�� ����2�$��"O�(s���1|y��ʟ%k�~�`�"OH�S�Å9�0AR0��	��q��"O������9Z����dI��Iw�=��"O�!��̠<�E�F	�k��`"O��fg�BcNE{�H+8bv�I2"OB��%�1TC��s�]~��#�"O6L [��i�&@1i`�� �"O����# @��p�D�����!��7���P?7�Bl�̑{�!�d�G/���¨A+8hp%�{I!��gil�3����+b�Q�:9!�$@,'�cO�F�lE
��2�!������D��Y����Ɩ>�!�$D�4(�!���V�?��c�Kޢ �!�F/q�� � -
x��� �!��ȸ:��t���_�y ���L�y�!�DK_ǬX�-@'I��sKD%�!���'��4S���AH,��ͽ�!򄑔<� ��E��D��#R�� �!�d�9}.��u$�0P�b� 6|���&�b�уў��섊�y��d�d�s�T�:��ْ!i\"�y�ˑ,�J2��҆��-[A�@�yB.�6o��I`��.�tii@���y⥉��P�o�
[�$C�˓��y2,�5C��\�d�̤1 9���Ȫ�yb��ԾL��S�}&�9I�F��y�ₕD��0ڠ��l�ֽ�"*���y��0bD���0�� KrmI��y�aH�E��"C�[+Ǯ`1���y"��<- r�h�MC D��!�V&�y��р!���am�:0#�uaaJ��y���q�*}�ƢZ1x%vb ��6�y�	�=6HfcV��o2�A�'�y�E�~%�����~+�J�o٪�ye���*3AS&t�l��P���y�����B�<��T�pf��y���`(h����/��E)�yR%�A@4��_�U�ZYr�D>�y
� th8�Ի}���)G,^  F"O�{V,ڎ4��]JE���D��"OLi���8�B�P=?�P�"OV�`�Y�d��3��T$��Ust"O6Q`j�!�@�9�H��O�KЧ�y�CM�b�@����<Nd��Bg�-�y2E�h�6Lh�o_Iv��vjR��y"��98Gj�[�o��E�Eb���y"�� n���";�䝠k�yBWR��3w�]$P�
��yBfH� ��rA-Æ^	�����I��y�`��m��@ⓤ����n�w�<��:��9��_
+8�8�$)N�<aG��V�!fk�ݚ�Q1��M�<�"���{&Y�_�d	�����PT�<��M�0?_�!�������W�<YqN�#f�s�g3�,ui��}�<a�F76=Ƙ(�j�L�@�I'�Ho�<!�!ďgn� �L',ܽ�f�Am�<��߶�(�S��"@���Ph�<�р�D����.S�U��<�"��~�<�blI�u%R�s��G�#I��@	Dq�<�� �7DJ��Wl�%o�:-괃GH�<����$O�$)!�6?[��i��A{�<��dNh!*���۲�\���a�y�<�@]��L�)R��z���"x�<�a(�0=�0�{S�2 ,��r�<B��:�HUŁ�)�b�l�<�V�������D'y����uH��yEz; ���
��yF���y���Ib^]P���`{ �_�yRƼ^�D����	���A@bƂ�y�	�b�@��˪��*ݐ�y"��F�.�3���{�����I��y�)_�P}R���,��x��,
D���y27;gp��D�t���sI��y��\�P�r�J4e4AU��yBȉ�y��B�hp>!"�j>bƱy����y���.N i��!j�Rt`BE��y2�!2tx��B.qG�]��bއ�y"��x���c�*ʡdc8�CQI>�y�!W�w�ġS�F;d�z-����y�釿*���T�l��^ �y��Q;2�\ ��	�R485$U6�y⢇�k�<�y��9)�r�8�)F	�y̏�]�����i<J�J�Hr�B �y�n�8;� ���ՊC<@�e�y��	����#��-�h�C�O��y�]�y��e0�B�{ѧF��y��4��5��`u���"��y�͍";o���R�S����0�yeQ(�}��h��Y������$�y��ӊ+Y h��φQ�6����+�y�X����e�N�^�r��ݎ�yr�^� ���P���ءb2E�=�y/\�; B=����a�*�h��Hj�<!#"ٓ
��"��5�px��B�<�i�J�F����&\����(�@�<�eφ�p~D�����[�y �|�<�!�G;IΩ�e�+2kn�a7� }�<��/�����3�@�v��R�Xw�<ёAX�erN�1rQ�E�p�h���r�<�5@�t��s��A�~͈��l�<��oҧD� Q` �d�xy���g�<�  ��6��1'�əo�S(�P�"OaX��ޑ@��H6m��B 1�E"O��YņZ�)�l�p�(����"O�-��0t�mE�s��4)�"Oġr�Y rC��;4�ͿuCD%ې"O
�q����A�\9F�B9J y�"OD�[�[�f깲b!BU:ei�"O��%ߖ7�V	�� ��$7D	Ƞ"O%i��ߗ���S�n�P�"OH���,
3`"�0I��Y�V��#v"Oā����[g�5��l@�Q��LA"O�!�L�?f�0�R�F=��5"O��x��K����2 �'���a�"O��[5 �n�|	R�!�K���9�"Ox8*��ɼh7���ekɦO�&��"OZ���|�6̓6�|$�i"O����FE�<5����uoD�&"O@e�r�$|4�2#O �,ek"OT�IG% :������EbdӴ"O:���S�NRU(��ݟ}U�$9"O�%ȁ��"�h���]�z�a'"O��sF�;`��D`CV����"O�m�&�U�t�9�Q*!���"O6� ����a*ed���J�"O&q$��8tF1笂����ط"O]���	�V�>d�TK�9u�Ԣ"OԈ�.�n���V�/�R\� "OP��ĩӑ7�0-�`�)0s(EK"O�}sn
�w�K����F^Ԑ�"O,$�!V���E�y�FTr�"O����Z�B�Q�P�ٸ=��D��"Oh̫��X?i��C5���~2,�"O8h��� ��Y��D�"B�+�"Oh�S�ۓk{�mX�F&�P��"O^���/+Fz������HyV"O�B�B� 1�\$;x��� "O:�"T�fo�D�fcʙj>��*�"OС��ގ ��kB�L��-��"O~��Qo,l*�-
� �2Au���"OĬ���WG�X��#\X�`BA"O��'��vk�Cc�8�إѕ"O��4��>jX|H�r-C)m���S�"O�}����<�ʁ�˃.R~�3�"O�p��ޔEJDxZ�i��H�#s"O|����ǷLC�A�3��T ����"O�`�bޢ2k�܊���/ �p,�&"OnM�2G\�W6ntc@�A�_=��y�"OBI�儫�mq�G�.#.��AC"OV��l��c�f��FH/J�2�"O2u����K1��;G�آ58�l"O����{eb��"�+h/�u��"O1(�,��03��%r(4��"OP@���CE�8�/�;.�ـ"OD��M�I>(�'�)h����"O�\���#u�ш�戍}ml���"O�$�p쁻.�Ԙ�Tfћ>���Ӷ"O��r��4-- �+��#(v�1x�"O�|���D1*�+�KQ�lt~}�"OL��tdQ�T���#_�O���g"O*E0*�'Kz�]�a�g��"O��3��ļ.�B��vo�*�	'"O$Yc�
�e��j�J���"O�
i�/��<: �CK
,jG"O��8�K�p̈T��/T-]0P�'"O� ��R�d#�|�"���K��:�"O�P)��B�Uˈ��
��Z�r`�"OvЫ�j�S"�bV��6��-#�"O̛��� }Bl��fLL.n����"O���B�;p�<=2e�W�"2���"O���ơ\).�<�u�ʢX>RL;�"O�TpC)��(-B��
3( ����"O��	�NIq����e.a��"Of9��/�T E)�}�P��e"O�a��Z�^�>	��AҾk]J��'"O��KQ�%q�7��P���d"O�``E����3r�÷K(��"O�僧e��f�!�3��)g.i˒"O�����W�E[*�-^��%"O��C�Q���j�)Ǐj"5� "O��b��=iH,�E��h���"O���v��K������&K�U�$"O�db���$A̕c2�: H��["O��i�ǜ�P�*xs�,IB�*Ob��+�3�̴��S�(Q�p�'�Hyt�	Z�:	9�㕑j.��:	�'�p���&�<Mf	�qrBEQ�'Ǯ�s%ޒ&���b��Ҩf�Z���'����>4������+d`� �'���3Gꀺ^����˫{m$I�ȓht�9�w�]�V��m`�	�f�D���~��PYӠ�+��m25��
��\�ȓI�P �V*'e�pc���>N����Ɲ#$M5�(�q*;/�F���+nq1'�"�t��&�X:0`q��
�h9$�ӂ����g��d;����Lr�}A$��#+m�9�� �M�n	�ȓO(����To��!���_�8���?��Z-L"���x ��cЂ\�ȓ�\��h�3ON��G�(8�ڈ��a�JYC�k� ���SbW&q?d��ȓq=LI*�)�(��z�jڢHK�l��!-8Q��Q3ܩ�0f�39�m�� w^�k *�&hY�UA��+,�B͇ȓ �D���B =急�"��2=�(�ȓh�nr&돕>�\Y��L�pYj�ȓ|���*6Đ"=�)Y�B�k��e�ȓ)�U9`�C�q��,����D�h���XalY�$b��.��s�RwR6��ȓw@v�R�퉞�vӔ�J�7v��f�f�S@	�6�~9
CAX�WP��ȓfl���@#M0^���Q��W3��a��h��qlJNY��9'�C�x+t����T��7�BL�`���,��Q�ȓ*nH�eD@��R�#�
�U�Jt�ȓw�.��B����H �G�+\XV��0<��{sF��s��)I{��5��zilxX��N/P0y1힉b.JȄ�o��@Ā�-�
���k�-L̘ɅȓJᬍ��C�xPx�ad"P-e�ц�'�"����tU*i��+s���ȓr�I1��V�B~mQ�&R)czȓ$q4`��ϫ ،�ǯ�!�r ��b����NT�)"�}Yk�E �$��:��ٳQ*��I�ܸ���ז?�T���`�lC�P���$��$�.7`���W�M�M ��<1��5_Ҳ��ȓHo�0	�H��J �d`�ċ� J<��Qp��)0F�.B5rah�!%uR�Q��S�? ��xv��hz�R�bW��A"O�D�C'�3Xnt�"!b�d8�K�"ON�1�cY�O�J�ʃA��j�(525"O��"�	�	o�B������fǟ��y��C�4�R	"�ϪX�Fxa�S��y�+ܚ �N,0�0}�tظ ʟ�y⊗!@� ۔!M�p�V�PՊ��yb�Mr��x��f�n�9�g�>�y����Xh���%W��P�!B��y�#�B��d��cHe�: .���yB�]�z��	w`�v�x(����4"���S���G�9�,�k#��=r����h2�yR�ݧR\���
n�~��!���y2BؘI� �q@$	�c�F��dɭ�y�E 6�����LD1���Apd��yRI��>]����+
K�H�@�8�yr���7��iwe�Vh�U@'���y�����pd� �����d#�yҭ�M�~!�	���MJ����yB�,7f���U#��
a�N��yB�� (��Xp��͞�ƀ<�ybi	W������_i�����yR&�D9Ĝ
p��3�|=�4�p=�}�WP$q{�@Xm`]��gȑ�y�P�q�$�$@��O^�h�b˛�ڈO���A�7b���+2c�)\�blQ�� l�<90͢U!�-����#"Qt	�p*�|}��'�45�!�Q�6��ӫ��j- �'J�c��.�TX۲*��V$���')��p�c����!���(�<���d;O>$0Q�]j�� �[2&��s"O��p3�Z#���vL�j���&"Ox�8e�1rx���ul p����"O�(䁊�8�RH`�*�O\.er�"O&�8G$Qm�𠐩ũpД�b"O��PAB�6�X�6�ĵ#B�(S�>�;Șy����@r����քbT]���<�;�jђZj�A��P=m��|r�0��"� u� q���M�a1�=�>�דPN���\S!
�b1��(OG�h�ȓ^μ�؁ϝ�"ix\���#WbM�ȓ w�ȃ6�)eR��j��̖. �t��c��
a��6���R�K�@Z�5�'~�$$|Oj���:w��$*Ɯ@=���4"O�k��B�T0�1�Z/Թ9�"O�y��B�*,�p�ҕa�)�0�"O����$ݽC�:Y9�Q
�n"r�	M�O�m��&̡1�z�:w��"�Fip�'���Âl޻!7xq�v��-�]�<yU�ڞ�)k�2M�8yذ��_�<1b僸?5�qZ��I�8��07J�Y�<�2,���$kz8�k���U����W �y뇏��[��P����z�Fz��O$�}��P!2�����^�T���"��eX���O����X�$�����̌	�B�jd"O�	qDƲWZ�م�U1{�J���Q��Dz"�Ӌ8�`VE
l`��1jF����'�h��dޕw"0�{�T @������?�hO���Ч_�&�h��Y�9M�48DI���yB�G+KD%rsiB�}R!yT��ɨO�"mB�~۰E�`. �rZ] �Y[�<����H� |�E#A�@��J��<���ٷ���ÓT����P��}�<�ciHFB��`��)�l �˔U�<� 2�(�!��Ae)�*�@dQ�"O�!�ыS�'�LC�7��i�"O��@�O���2h�nХ"�"O�hs��B-R��`�M�f$��"OVq$E=M@���T�4aHa)�;O~�=E�ܣX{�e!b.�]DvX�*���y�!Q�=r��R���6;���$E��y�m�\���fRq� ���jÃ�y��U(*V�*& I2~�:eH�N�6�yrGDY��zF��EUH0���%�y��Ɗ|��1f�|����k���y�e�76��Ly���c	6�B����y�P/����͆k.~�(S����y�Z�f9�%���b�>)s`����!�$Y>2�,(B�E�@�
��FD�)3�!�d�,��a�
�}��	���%O!�&!��\��֎>�XYP�g�!�D(Td�*�B�"I�h�g��y�!�DJ�]=P�jE
Z�ػ֠OO�!��X�;�8I�f��0HYcT�]"C;!����&�����疥 �tr��f&!�$ӴS��\J$�l�l�nv�!�$@=^�ڝ��E�?�0� g�S5�!��p
B*J����#i>M�!��^�B�Z��A�H^�&|` �"O����/G�t�H|`�GK��X�ʇ"O��b4��6�x dG�4�Xu��"O�$���1)Ep�C� �5��hp�"O:��Q���h{@��eM����"O�9�EE91�ٚQ�ĜD�1#�"OZ���#=��������`�:�"Ov�rӇ�0r����F(�p���"O�)��"�=t$A�R����HF"Oli�& �*5���h��9���)T"Ol)��-�&Y���ڐ�B�E)�H�'"OB����C&M��0kF�� {
~TH$"Op|�c@#t5�B��͌4�N�a�"O�M����P���cIM/A�؄q�"O"q��G�(B�X�V�&m� %q"O��RL'=�Pr"-�Q��T�&"O����<$p%cqi�M��-`�"OX�ZS�3�(��E��N��Aq�"O��n�i" q4%Z#���"Oh����=q�f�#�d����+�*O@�KW�R�},��P�8�I9	�'�.�ɕ�'���  3qBP�b�'ܐ* �N�u
=P'�C�t��1��'�D!�%eW�Y�nP d��=�&xa�'s�\�7�����x�痺�i��'̀�)����D� 6�� tjԙ�';*M1��L�k�� Ye�~F�m�'*�U�Y�Q�m�t`
�z��X��'��)����8g�x ��k��1��'�j���Ϝ	M�E��Ȣ$d:ْ�'ND}�ph� ��P��΁��ƅ��'�p�	�M'140��!�	��a�
�'��):���O*D�R�E��|���	�':x���!�6b�N�p$}�����'a�@����b�����Ilz��{�'q�����zu2��'+�4_��r	�'t��9�ɀ�d[����@H)]߮03�'�e
����u���`�*G!2R���'��1R�!I��Ya kB6��q
�'�T���!m*=�G(���`
��� ��q	�6 0�T�r��+Jl��"O"1�C��:Z���B�dΆFj�*�*O�u��	@{Qi��}�z�
�'�H�+1�Q=Ѩ�xA�ͤ?�"̡
�'�"�͇�-}j�Ɲ�fΩ�	�'p�ȃ�N��H��ĝ��:�	�'Yf9K��c�B�a�*#��*�'A���&%�0���[��9�
�'��c2�+&��2(΅&�� 
�'��ʀLW�y�z,�qal�0���'�h�	gkA�@�&��0L	6322p��'�#'�	<`�����/o�8��'���	���Gd�-0��,��}��'@pغU��$�
!Y6���M	��!�'��xЂ��3<\@�H<|XjU��'�]�Bl�s�tq٧v*�ɫ�'����υ�֥��iNa����'K�	A�
�!��ŁS(�2[�0��'����GO�	*I������No�ի�'��`�_ z��єaH�H�D[�'X>D�2�$0�xKaCu��k�'�a�u��;5�{��k˜=��'����Rj��#&�	0�_��r�'�ZG�V�I߾��g "W�X�
�'�򄳡Ȓ�}�A�҅�Z/H��
�'���Z�IM7�\q���W�����'�T���ME��:a�_	V�8��	�'�z|R�Γ)+�B�cF)6�	�'	\�[����]4Й�s#�Z���'��Y�2J̠�	惛<��'Q`��`���5yޑz�cC�tO"�J�'�JLP��ζZTx ��͉@� ���'�^@��� ��aIr69��,	ħgu.%p
�N�ԑ�C�]�^l͸@l>����ȓU-���o�(i%������!r��ȓ|�jm�CH!*��k­I
9@��ȓ2\�=�F��}R��K&��[k��tR���K�mZ�9AD��L����ȓ��4�V͒�Uu\�P��a	~4�ȓ_�ƹIB�Q�_6���Sɋ;CŰ�ȓ#(�"�k?O��Ljd,�0P�8 �ȓ/���O� y�R�J�E�|�|��ȓ;.& ��T�8�X��+2bZ\���l���4o���B��ƍ�� <��n�:1ȑ'�4)d0�5L�D�(h�ȓ[|	� l ?�6�i��R�X ���ƕ�A���F�q9�I��p�d��ȓRY�tRtJ�e�>$!�c��,ܴ��ȓT�ʂ�
	�~�PR��htb���?],�+�ˠ)]��X�Β��0�ȓ^%� ǥ�1�^�p��	U�^���b#p�&�$/Ѡd�� ��l9�ȓX���h��D<� ���Xў}��x 4��iŽV�BhP���yц�� �����EaL�!)Y�9�ƌ��"��,#��[9Rm%�է-NP���;�h�8∗�{�Ή�dM��;�T!��56�4�pNТQ�Cc&^
�|a��j��o��>�耱-W�*�.���|�R]�tn�|�n���&�1�"��m�"]ر�8GN,��G"����X��m�Ð6�PSA��4��ȓi�hՙ��ܟy���ٯ{��ȓ!zM�F�^-|�#ǢW&4<=��S�? �ݺp-^�]xy�����8���v"O��XG�R���eW�V����"O�)��`ز�50e�F�Ƭ��C"O:��EAV	-��͟2g�T�ɠ"O��3�Z2�|-(�[�����"O>42��L�g����ū�44�n0�F"O6ZF��J\��1J��sEl�b"O۶ _�|j���( :��[�"O�ղ��77%N�b�胟Z3R��e"O���I!Gw��:���e-L�{�"O��աH�7C�4��v"O��T"F�1 N���
ɻ2�.�Z4"O� ��Z3Tt��K6�K�g(�S"O��+vk�8Z��"�.{Z�9u*O��W�W���CЀM�����'�z\�@���i^��bR9n�'�$�K�a�x�u���Y��-�
�'���a�VtAv@ Dy

�'�6�ҶCO�,)Ĕ �J�M�4��'��|��	����\�Tb��E�(���' 1E�(3ɶ`��F[�A��'ֲ��3��]����B 	��1��'^�7�S<h��`��j�s�'�4�e�<P������c��B�'Q ����{,
�LaÈA��'ҹ� C@dh�0rl�VY`YH�12�	T�6�)�1|Q�E/?2��D!)	I�Z��
�'�hy+iUl�D�S�eO=��Y1�'��h��^�.y~��I�x����#Ƙ����C�%��s�h�>�w�?9c��$�?]WF%y���	�R^F�a�	Al�.tɔGG��x2c��$���V��rb~��(���?1a��l�A0����d��!��mZ=��O'T̒E����jb0i���ߑz!�V�|��#�l�eɶ�ۇGET`%����?A˼�Y�4z��$R��?�+�Kg;��O���-�..?��b7(X�e�5ZD2�O�$�@,�����Ff�3.�yłٲKgʤq��D&p0N4aa�T+�����d�@h�'��0�YR�֌�bE�0fp��Љ�$�> ��g�ba"J֛^��#F,O�08��w�5�v��pOذ\čCh�: ���IOb��񨒬k�)��
�Ay��5m�.�&��A��,�|�;ħ� ^�v̊A�Ӯo�=��*�~��w{h 0�J9"Њ-�L2���'7�P�'G�(w5�dC�[�^��ӣa�=��h�$��3������8N�È�eJ�$3+O,�B��Q�����OV�R���'~��bt�@�6�u�%�Z>5EL��c��k��m�#�,"j�k3d�8�x���ݕK3��
��V|�'�4���g�&k�~8b�aɫd	P��}�JY�|��D��������(]�!��0� W�He��o��\sn�z���K�h�I'-��[��͇�I!�����N7s�$)�Dɗ�()��8�(ȓ.��L[.�O�vu�"�K�'��$����q�"-�'U��1*R�j�%܊�4V�qr��D}&�U��>�a�	�[�� &P��q�cE��U�%�	e1�a-܅9Q>�]�q^rpi� �GJhHgQ�0 �hJ�#T$L�CV�8Bu�k����к@GqO�1=EQBh�.)��#�
�px�E½��%���0r�����3W2�Q�_2���	@��\�rJJ�J@êČz*D�e8�H�ƕ��X���S�mUXa�H iP����8�(mQ�/�Ȱ�V��[S�,�V����d9��7QoJ�g���4��Q[�$T,j�TAx���&h��1a��71AT��ViZF}�F�ޑ0��qcӄT�k�V�'Y��n���9 C@ˣ;���� �� 3���BC���gQ>}2��
�u.fR�Ŗ�n�6� G��&Q�8J��#T|	��(Rv���݆*�ܡإ@]F�5�O�-:��D�IJ�V��$��,"�1ON0��@�0��)��]
��Ņu�ք��%��yY����54B�)"�T�iT��K�'�+��q��#�L��d�C���:b��5�X��$;�Eh��`�	�Jq:�H���8_K���ϐ��FIN�!
�3rIr�2����U"T�x�+��#�!�_Q�dhT�ص8~�Tk� 	-A���)eA��@�i�S�I7E��
�k��P�lxD��4�w�IQ �[9]�ha�O~�ҭpa4D����R���iT��y�t��a x�*x	EH�C"���{,��2
_@Zf�0�I�~EVy;
[�(����-�*x����Ҟ<ֶ���:A�����בh�H˳�%�:�"��W�+�|	ᡦ*�O��a�^�N�f�sD��Y�Z}	r�䕫-D�t�SF��A�$�AfH��g�? hʤ����	��t�ڱ��"ON(Dc��zS,p$$~��"���@1J���SC%�U�w��0,S�>�	�*������G�j|s��ϫ~B䉳1|����);zu�K6$K(<���_)(����)T�pc��s�'��VE�L�Q'`��(~�����`���P��Ka�%M��C��:��Ő�b�F�P��93��"�M� �lL���J�\���Gy�ɸ80��9bn��nH�|�2��c��ɋ���s��Y(-B�<1���\M�=f�k9z�G͙_0�D��'�+�e�(��)�y�c� @bi��O.;�ap�'���Q4�Q���!�'	��8�t�O��K�oR�paz򯃏g}7Dиq5B͸N� �y�kA��$刕(��M�.NFX:�'E����H�$��� ��&��X*�'
̼h ��p�R�f��1�ݫ�'4���T�%7������'�Pq����;��X��L��Z�'L�O��<	���sB�-	S$hH	�'�Q��LA
l�n̲ЪT�8��'WP	t�(0���
����8Q�	�'m��"2��:_��l�D/��r��0	�'�$�B��@��zdi�?\����'����G�>�Q��W�B�5�'�����L������8d��'c^�1�k"�H�5'�:�R�'.�j�OOR+��Ζs:0�ʓbw6���i��C�=��BӸz�D�ȓsd��;&MF�c6P]�r�ͳX��q�ȓt�
Ux��-�ȱa�.�4:�rx��OV@i��VD��H`o��9�*�ȓ[o���S/E�X�鈁"K�a�}�ȓBx2M��ϫ'
%���/�Ɇȓg��x����$�W�c�v�j�'�:��&�ŴR�:|ГKڔR�lI��'}X���./3�h��k-B
���'M��6!�7&��%I�> $�:�'0������Zqi�7��Wp����'�4�3��<��!����AǆX�'w��� 
�
�R��03��0��'�(d����HQ\P�)�-��'�pHqE�]P��)f�P=#ڼ��'�2ْC���	Vڍh��ێf�K�'�����35�FYɇ�U�(�T���'"��扳HJ���	�*N6m8�'��Ʌ�^�r=Ĭ�A��2P|�5�	�'1|�Z@��Nтъ `[�\a� ��'�$�3�(|*E��E�+[�r�'1��Y�&���駨�#a���'��0@��($�(A�3�X&!����'�
�uױ4լ�+4�ɒ
.
p��'�x�#�%$�j�U�0��0�'D�����CFX�G�^.� �''�<9�/U
`;th�wOQ��ѹ
�'�ah��w ��f�{���z
�'M8@S
Ծ)���|چ�i	�'�p5
��ڔZ�ϭ~\P0�'6F4��O��ji�I�$�1h�����'�xԋ��Xg��%r��ܑ>���'l����9-�N@�󠅴�H���'+�Jա8N���#�/��В
�'�ʁ`����z�
�k�;�ހ��'Azy���abԹ��ӯ>=��2�'��Q0!�I�X�Ѱd��4U��'e��^��}�&�ʕe������ ��;���7���J�In���"O���«�^�؃�@�&qa�"Ot���Sl���a�F��5��Q��"O═p	^�t�(p1��$O۠,Yc"O�	w��1	4z������:�0"Odq+rd](�	��%:�(P9"O&��Ǩ�+�N�0��8��Բ�y�B�{2 	W@L*��$�ц�ybn��\���B�>F������<�y�K*~x(r菢O�ɑ@썊�yRS�Y�%Z�+��R�ܻ�M
��y"���Ρz��:Q�l����y��"�.J&�X%R�����ä�yr��f��J�/��&��Л��yR�<I��y��I�e���@�H�y�̐\>Z��l�Q�H\``L0�y��K�-��ī �ГS�PH����y�cD�J�͹a
_g�iс�S�y�T�����hD�\8 �z��I��y���2�\�r#J�,|L\��O��y�ü\b�QS�C�v���Sp\��yb�Q�x:�����y�2i8gNƦ�yR��2X`T{�dz�	��ω�y�# b0-I�(io���$Y�y���?o��Lj���	>԰ȫ����yBfߚi��*���3�>%D�P:�y�	�6jx��#N�%CU��y�n��%ը` ��_���y#ج�y"l�q���a��+hB�ړ꛺�y�Ó$]��X��M�g�P����ȶ�yR��-(A�8�`H\S�=h��"�y2���:]��GAX'�i��Ņ�y�F"!A������&1��0HB�y2ȕ�c�4����W�,sg
X��yBF]`�L� $�H??Jm3��گ�y��ލ|���9L�� �C3�N�y"a�8A�nM�&j|T8�-P��y���B޴�r�E){��3�m���yR�ޙ]æ�:�eI� 7�Y�[��y2BG�r��0h���&Z��0�Aӝ�y��J��(#��2�R����y�(\ ��q B�T�'�-A��*�yRf2J���b�8"49�+�@�<��֩W���)6�<]�D��P���<�� U�������D�j(� B_�<q���BK�\+��9<�����F_�<�q`�VC����l����9s�]U�<�S�P�����1j㒑B�dL^�<A��� Ԍ��_�~`´��X�<'⟄eZ����h�Z�`�A�s�<�'���Xr$"C�9Q��A��^n�<I&�ճo8��)�J�/0��g�s�<����m�X�(�!7�`�P�i�h�<��"��T-��D,_�V����BF�h�<!@쀲oJ2)x�eԤ'�N�"vnCe�<iES�\P��Ê
�����u�<飬��S���б. ppȣ�%�^�<I2�+z�p��J�ԑ{��W�<1g���h�ȭ��ދL��i���K�<I���<�Xfʀz���A&�O�<�a�V#VG<�K�G��:@���@�<2��c ����@��I ��EG�<���V|����D��� G��2 �y�<�6͐"|^Ly�D�:���S�̒t�<� �Ź�@��
G���E ,͡�"O*� *����Z��ȕRT���"Ol-�T-_%y[��rP��C�$+�"O�}���]�M�@����s�<5��"O���Vm��aQ�3@��0�"O2I�U"ݫ{
NP�f���V�T���"OZ @�8,��9���O#KaP-�0"O�("���?o1�m��K��{ʹ1�6"O�MX���t��)ITI���.��"O����m
O�n�JS�[8~�~���"O��:���Fr����"��O�ε�"O.�8�%�<cI��Su���^�FИ"OF�Sd�S�1�����w=��K�"O�!A�F˸"�����6 �a�"O� �t�"V�������1����"Ol0*���2_����u%V�,4�s"OԌ��G��z�����2���bq"O�����V��� �D� ^_��"T"O��RC��9wd�Q�cӼ|�f�Z�"O�y���+z\p`"��~�h�r"OM�P�2���a��&�W"O�|0��-=i���ߍm0�A"O����͌-�>ٹ ��s[&�q7"O���$tq�tj�
Wx���"O�pHiV�s�Jd)�I�7o��Q�"Oz}vh��3�a��O�,z�9�1"O&�z��s�ġz&�;*f��Y�"O<��K��i�N8�pL�&]�� "O
��s��%%�U�0� 627i3�"O�P_$�`:@��Z	B�"O����d
�NxQCr�ޘaJM��"O"�&�S?r��u:�Y=u���X�"Ox�p�[+jUJ0M�9K�<}�"O�	R�	O8]��8 �*����"OR����g(����(� �Sc"O<��H�@[��V��e�Ƅ�"O�PY_x�� �C��46w �(U"O��(Ԏ')��F�Dxj��"O|�!�]�Q��F`��Vm&�S�"O@MBcI��p�.�W� 8o��"O1+���9d[� +ǩ�
9��K�"O��s��/,˜5�0h�;sZ�C5"O8̠��f�-� ��n[�݉�"Oޭh�M��g�Fh:E�	�����"O��T�_�;����	�^Ɗ�(�"O��7J��0�[7�F_��Z�"O.Z"k ��%�(O
>~���"O��H�nO	1/�3b&C�pTle��"O���e�F:�p�p�_O`���"O�vo��|]C�B[�L\$5��"O�a�%�O�4궀I�jHZ���"Oƽ{T�Y9?�Vuk�O�@t�"�"O<t� G�fA�u��{���#"O^Y���]ᮍS��C"�H�iU"OP�y�!P�ck��I'IZe�lJ�"O�y�M� �r�#T�@B�05�v"ON���H��u�7ALa�(Y��"Oj�#�E�]zf��"`YsҶ��"O���ͧc�2E2��Lͨ��"O\x�e��%]��(!a�N�6	i�"O�pgdD�A{�5�E�Gn�(M��"ON���f%M���n��V��DÑ"O���'��f� 
��X�hT!��]"D��_U�1�"�!'H!�� ��r%�YZ��� �TTc�"O�pU���r�|�tE� ����"O�\�%ÌI��)���ͣm�fA��"Oԩ)b�E�j�*�$�-d|49C"O"d;�ǄS�e�¬��`oh�"O\0ʠE�_�v�iQJ�EP�@�B"O8�kq��j�|P1�W9l�>4��"O�8FEޏ��34��3j��� �"O �TET�a�HXJ�dI�Y�Ԝ""O�j�]C��z�#���M��"Ohha`�������s�)`&"O�ar�e�I[f�C�!E6��h��"Oh��J��y��jX�w�&�St"Orp{u�!�X�bp� ��x9B"OB8*�#=&��҇�(���*6"O��:3��ub�1�,͓~ڬ���"Ofl�4�×"瀉kaLA�O)�i�"O��cc��:/:Js�BC�p��!"O����R�E���S2|�Pb"O����,ū"g*�JwŅu!��Җ"O��+��ӯ�\ʣE�("��
P"O@��s�C).(���F
.8F!�'"O�5���W�p��ǐ��1��"OT�Uk��Y7�E��C� uI3"Oh��qLV�}��T�2'D�v�J�(@"OX��ѿt�4��e�	c��� �"O��hM4y�&p�E�0�lmC�"ON�ƭ^-<&>�wG�L�ʀ�"O���vN��U#Fu�B%_!T-,�4"O\�J��'MERx�veR�/j	:�"O����� d�-�%Ś�k��XA"O@��4E��xt"�kڝ1�d��"O�9桂"L�a��:���x5"O0�)� ��h~u���	�b�X5u"O,Q!ÁK��Jb���u�,t�"O��@��v�A���ρH�0۴"OY�#��d >d[s#��z3j���"O �����"�p�Ď�P��`"O�!�ū_?8*D�bOs��Y"Ojxkgo����E3׊�F��}BP"O��0׉T�m��U��H�s,]Ӆ"O�a:��U�|����j4���"OFx[��� �52+�	SeF�J�"O\@!`�7�bhs�J��5^��*"Oֈ�#�¦/J���	T*1
%[W"O��5�� ђ�(��K�x^@s7"O�j�!	<D�E��m�~!��"O�����^�1��64��b"Oj��sU�~6%��Y7RY��"O�] 7�7.-��b��ئ�t���"O��2��Y�oм���)ꮀ3R"OF�	 ,L�N�0�#����@-{t"O��:�J7��F$48��z�"OXe�)6�tm�AC_;L���"O���G�u� jt�&r�n�*�"O����aػ\�"H4 b�P
�K�o�<��`0L�x@�QFU7A�R�i�`�<��o�Hp�S'�V���˓�i�<�Ch�mψE��g/U�n�$d�<	bJ	�-D@���o��ns8���'�f�<Yt�Ҟe]�p��@!? ek���d�<�' �I@�DZt��!tRZ�2ց�O�<A�I���MP1�a�M2�-�H�<�"��s(���㊚.&YJ�
�I�<� ���AP:���l��-�`D`�"O��A�۠Th��f%�$p(�{!"O��%��!~0,��꒲*xt%�A"O�SQ�C�J�C��Uv5�E"ON�I팂h �1�wA؁v��P""O�h����8|�9w*�;(ɖ��"O,��_� h[��1���s"O�Ԋ��;^&�)&j
[c
�"O��y�a�,z����a*�^�>#!"OܠT+J�z�h��qlN�~��(��"O�Њ�Ꜫvn�L�ТB z#Y�"O�|��i2X�A�aF|X��"O� �l�9�,�1�?Z�Rd�$"O��R�f/6��$kۖa� )Ѡ"O���&���Xѐ�U2!���:W"Oة�#GاG��h"�|���ق"O��)�ޥ ���B���c�Ba�"OdXاό�$�ā�	��*�ԩ�p"O��5-�9�|E(�ƚ
YJ� �c"OB��3T\
 ��$K,h5���%"O����&�9��9��#�9C"8dq�"O2I���Is��s̴P"OԨ鲃������"���x$"O��r��;, H��c�DU�ă"OK�a*Zq�#/n���� ]��y�i�n/�DZ�S7'ڑY��Y �y��:k����k�3ޠH f�P��y2F�f��;	G��H�O���yR�э!�D1�qnQH���P�*��yB�Q(7*`5����=RI��O��y�Ńh��,2�ٞ0��E�`×�yro�5D�&�Ht�ɂ3�n�;��Z��yr��8"��;���,����0A�,�y�e�8zn�P+��$�vQ����yBQ����+��+h4a��!�y���"�$��0-�2 ;����/�y2.�����U�L�Nd8���-�yb�U4pZ�h�e�,2�.06�X#�y��݀`�$% tK���@I�����y��Z'���a"��e1�4CUi,�y�
�p�,!����`��\A��M���p���0?�6H(�(9�
*oҎ�[FX�<٦N�7�B�ՈO,7@�:���[�<)��.D����ǝ[���ɷ��p�<I+�Rv��q�J�
q�3T�^�O���a�L�T�1Oq����b�7E����n+Y�hUS�x2׃[:U�b��|����c�F�
S��3pHrhx0$ʟ41N�-0T�b��~��*W!(r�kAl�'=q���c�{�p�W>�?�W����Y�wj��"���}�j2�'�UpG��)L��ǩV�CzyX�ޟ|"}�D
P�"�t�c���$a_�a
pd�2I��!�mG;�H�Z& FT)�ᓡ}�. Z�ǝY2\q��^�<2���"e~ލ؀��'����3C*��|)�a̞� ��/ߛٲ���n�r��Q.бJ���+����~rK|R" ni�1iŇ1��:���'�- ��Đ��#��s��nځ'�hQ��B���Sf�[�p�BC+�%[c�n}P��4&�����P� -��2�J|"d�+&�v�yp��0W:�P0��K�;a�v(�?�~�u�ؔb�^4���T�T���u�n�<9�.�b�x�(��O*�AvkE�<!�� C(�8��N��� R���<���s@b໗��5+��q�sn�w�<	�,�Y�m�d.X�%�0'��|�<�7׻!}���"���)06n�{�'�ayҥ�&L��qB�".�<�`�F�yR��#v`i��O�����&U��y
� "���o��/xc�O����p"O��2�[�t*��0���"ª�� "O�D2�	;Q
թd���dИ4"O$�/�
�̑��/ζ1�v� �"O|q�g#]0_[�:�]��)"O��!�(F"W���k�Z4��Aw"O0đfI+ؖE�L��-���	�';ܸyb��~m8!g $
�Z0�
�'�d�rp'�=	e4�Q%ƺ5�f=�	�'����ԃ� �pd]0x��	�'��ȪT/�<�D�G'�&E*dy�'M ��!=�.9j@
AVt` �'�P(���=z���,[�;��Y��':�"���2�&߃�f���'�j��A�RX"`��� i��h��'O\ &BY���cv��_ٖ�j�'Ӧ��Ă�F�
�{�+�6']8��'�0�c�gە:���1b/�Hl*�',�C���8�.e3�Q�n��\�
�'���`�  |*���I�gC����'��x+�+n´s�ūe�Ly��'����D4
�$9ҭ�d^����'%�(�)E�fg%h��*R(03�'��q�Q ����12���U��x	�'tl�)e��r\�IZ�焒<�X��'�R���I�=����Td��&XZ]��'��
֣H1���#.�q� �8�'!��
G		�p�2��V,�?p�BU#�'���E��'<�ZR�/˚k���
�'�is�
:$�آl�v�(u�'JDC*۞(��ic�G�=K��I�'R�%���Β)�K��F).F���'�ܝ�r΋�Mb��̅�TRL��'SD .�+_�u��ʘ"���s�'����΅od: \%��� �'mZY��τ�}Ku�ׁVJ��TZ	�'7"��c㓕gK�`�%��1����'#6esW��+�)�(9 j���'����e� �
9�#�A=eRܨ�'*�e�tˀ�
�|سm���s�'�`<Z��8���hАY�l�X�'l4��Fd[��X��cD��>	����'>&�(�eN+G�*܋$��2u��B�'?$��UF�$\�����"̖1��'�BYز������Oθ_����'\&�0��,<��+�(̇c�h���'v��D���I��R�Ckx +�'����bΑ�_���R��<��]��'pl�����K�h9�2�����'A��PEB]:>\�1l��,V��Q�'�ι�Bƾy1�諁E�(��l8�'Ed�2 ���hJ��+1A��!�L��'v.�B���>(>J��&¦���"Oxp���ʦA�IbKA]����"Ot��C�A�1�<�I���u���"O�xђ&�+k�%a&i�g�B��&"O�a3��7���I�!F���;t"OI�ĉ�*�jl9t��:��l "Oځ�B,٦�A���n$>%c�"O܁�%��qn��5I<7��"O�TY&Ꜻ4��d���˂F��y�e"O�xxv���6ێ�k2k�=*��E�#"O��Hv�K6�>\��N�c�,p�"O����P�z~�A5���M��dj�"O� 4�"��[�i�4�&�. l�"OP8hDd�?�9�O�5_��`�"O�Da��8Ը�C��Hw��#"O�I�N@�t����kȐo��y3�"O�E�����H|��*ڠ � �"OV���
��s�,ATI�g�`�S�"O���S�%��h�gѤ{Z>00�"O��y��o�����>@EXk�"O�E�s"]�([��ɡ� "qc*O��s_ W�����"؍����'�0%8���` �H�܋6�i��'a���Eg�4I4z��&�>�a��'y�h�a _DsB-*�_ 0)T�A�'�ν���f�p��*�"3��[�'^F���ɻg�Y�	�(JvH��
�'S�iJV�S�gs���wE;-��	�'^U���k�Ʃf��,���'�V�RD�7>tHh��N%2����'�J���Hh����e�[>��QY�'�yRu�J�U|0ar(�g~�*�'T��B ��7gw���NS���x�	�'��QK �˜��}P��)B���'v�PYgb%R�����P��ZQ+�'>z���-�'Q(�� ���)�$M�'B�3'W�:1�������$@u��'4�Tk`ᒾ;�VD��͑���'iHB�J&&\ִ�qŉ;Zp���'��\	1�J�7.�iP�۷@5|���'�d-k�c�J�|���Ꮑ$�j�	�'@ 1p@Y#Z�tE*2)07�H�'DD��"L3k��c\)�\�#�'2P���L�Y����P�k�H\�'�\\��Haq�pR����O��)1�'�Ra�FK5V�@��U*S&TX4�Z�'C:LB�a�6��8��Ҙth�{
�'�0,2�b[^h���#J9f��@��'V@0��^�w�UIr��>_��x�'8��u
��ʝQ�X;%~P-a�'`F�K�..-<� �JR����'K�!����i%�ɐ��
G \��']�E�M F�)agNs��H�'�&�!b	5��u�.	,.�=h	�'��f�P`R �+��׈��P�'t�غ'4x45��_�t�(��'�*\�qM\7Z.�$���_H@�X�'��bF��t��#��4p�  �'�(�!��yΈ�C3g:1��
�'P�hQ�ES#�$����a�S
�'|����΅�H��c��X��B
�'���x��#3�� K��-S�Xc	�'(4usD��i�hLJr�ʩP���1	�'����$ O�\/�R��K�~�0	�'%ح�uFYY��0��`��q�1	�'�,�C�7ѢX�Ѡ��y� ��'� ��)�#V�<,jBJ���P�'���"�^��N$�� ]� Dy�'�)��&�tuAL�T�"�P�'J�ȉdEؑ4�Zp���Y�PX�(r
�'�ie-���0�I"�D�' ~���a)y�AAR��<Y�t��'b��$��0!f��
�1��P��'��%X'îD�2�b 
<��C�'��m��?0�.Y�4�P1$���'�<�{�U���%E#�p���� ة�)+�hHh�hZR�,���"Ox [��;:���n��#����"Ȏi�	�4rz4�4 P6G�DA'"O��6��>iܙkV/̙{��=�c"O���Ǐ��9I�eYc�]1*����"Oj����_!:������O�8�b�B%"O]�V�04Y�fs�8�h�"O�%!Re��9=x|����B�L��"O��CD͝Mm,*EHn��C�"O��Q�'Y-F�r�#�v��aT"O&�Q�H�'?dJ�Ȑb 0R�A�T"O�l�d�4��S��&T�4hA�"OP=!��̱a�b���/ܒ|���H"O�4�����V�ǉ"w��A"O@���G^�X�ˬ-QT%�S"O�m�	�=��`����?D;r�Q�"O<Y�KQ��sd�a
&a>D�$����%ݚ ʠ@�[��U���<D�HS��
+�؁bÌ�#"\Q*PK0D�ЉC,�5aBP�#K�Q���"��1D��`1Ĝ�;XIJw.Ԣ\�:y���/D�("uAM�rD�JR3b{
qQ�1D�TX��Ю ^E3C��/:M�3��1D��b��/���e+��E��yC�0D�0:��eh���C�W$p��Z��!D�8Ƀ�ȇL�ΈD�V4|����W�,D�0H� q��J��
H���q�&D� A0�d�q�a���:r*&D�q��-?Vձ���?1JX|b2�)D�k�Ê�1^��r�W
F�R�	D�%D���2���p�q�wb�q�bm��1D���v��r)�yp�X�^��ƃ4D���EbP.����l�=FԬ	�=D�L+��/*�ۖ ��`��ɘ�):D��NǦV�Rԃ���7�p=� l8D����Q���P !����1D�4��͝18$�a��):�����-D��"���/b�y�q�KD�ΐz��+D�<��E�u��i�T�Ţ;�I�,D�py�K=Y�� ��ĕ|�l�Sn D�����|�0BO	,ۨ�� )D�|���	tOʌ˷� 1-�`�Xѩ<D��r.��t,����fB��b��s�<D��1������@:��@k��:D�����$:�$�0L�7nd�6�:D�P����,v|^�3u��r+,�K 9D�@��o�)q�����W��4�"�d!D���!mɂ	����'%
$0q� D�4��ݡ`�V	�`�Ӝ}�8%�!D� �2�	�d|Tإ�*��n?D��0�(�1keT,Ҳ`B�>a+=D�����$&���Z�Ϛ@"��H;D��KK9T�Yp�H��pr�!��i;D�����>k?ܘ�˃j��A'/D�$*FD����x5fBNd)�g-D��ZL-����u@U^LV����/D��3�+4u���@cK�j��� �a#D��� ԱS�Fe�GΉG��hp`#D� qc�j���p�J��Ĥ��!D�ԃ!"�R"|��I,윤!��;D�"�O�>5�\�C�H�n�j�9�D?D�TJ�k�T���Z��D�T$�l�J?D� iP
G�+KޭZ��Fk�䨈d=D�2g�ZQ����I27 ���`�<D�� 8�t↵=��4�]=D#��Ї"OpMZg�K3?�<� ߖU8�$�"O�����AQ"�$�Y�|��͘V"O���F(d�f`b"��eZth*�"O2��e@
�VJ��u��0*�Xu"O� �Ï��|�m�v��4ta�"O�L�%	   �*ot��R�Tږ���'�n��-��Y!a9>�T!�G��6U�@�Is�t�b%
 e}��xk�j45.�y7lW!_� �'
6T���}��neV���q�vPp����'�pDHFM�2���ֆU��*�	wLg>�YS���k��X	��7f�����C b�p�	��&n]#V�Ϩx4��D��K��� � R�-� ��K�'�-ꄎ�7 2=�B�o�ԠY��,��'��M�R�h#��-1`X���Ҹ�|�B�36I�à� � 0��*j��`�JP�lWj���7�����e�庆e�:Ҵ9�ъ/a��pJѮi]x��S`̙6��'c氐���վ��!-"ِM��$\O@�/�tE�����m1`�;8�6�S�e�*<�����5���3.B�_�Y��N�-�|3@+��{r��40閁�V���g��AlY���'r�� �����i�LTu��
����T	�+˪����V�r� �#���N�@��aLۍZT~� wM"\OhMK��8�XR0 ��$\ikb��5jz�c ���?�"���H([A$J#hDFł��i��4۷��-���A Zk�Շ�C�I[D�1�i�1�n��	�ɴDV��� �6�E�J[J�UcT�~���vC"�i���T:W�D=;�z}�'.��"�/��M�g�a�$�e����ޤxg(�7Wp�ч@\�\�pKM�v�bEW��c?O-�ߙ2~��ë���h�Of�:V�ы*�%�4��?|�*ѹU��ac���nY�HER��ۓ'q]�0�S	R���s�X�\����		Q���/��_���i�i�0���)�\�p��><����',*��W�ܶ����m��Y�$��y�-M�\�0��"¨{��>���k�d8�pNN�|j�`$D�<�EE� ��a��R�>���Qb��[W�@��1}���E���$A(	;�hA��4� Pq҆ſ6�!� ':��*��	U>�8 2��A��CʭL����;��HCևF�6�*d�%[<C�I�-?�(�CH�+��
C��Br�B��)5TT<B��̋V�Z�a�+֗v��B䉐{&xM���J(Z�>���;0�B�1O��AP.��4��Ԁ�;.�\B�I�ҁ��խ_ 9�p.�#N
hB䉟��Q�e�]�R�����FŞB�ɐ"���sP��+��}�Q'�$.%XB�I>y]�A��"�9uW����޴`�VB�1hՀ��d�� ��Q��<@!B��&����*��v$����!�j��C䉺^f�Q0�	��φ��6_�C䉅�H�3P'�t`R�M�l��C䉰']������#��(: ��4i��B�u�q��P�2���
�̰B�	:,���O����r5`��r�B�ɂ6������X�8�����e��B�I
m�2��p��)A���4e�5)�4C䉞%7�R@H7p��tˢ�ʛo�<C��=�f�H��т3t� �����C䉭H|���Z#D(I��֡*�C�ɴi`pYy��U�(r�Jվ`DC�;�(�Dϑ� [N0s�V>9C䉍,p��K��H�T0�Ei��<1�B�8����� �:lB/�C�I7
=Jq�Ƌ)98�es���7BC�	;k�0Tw�5s�9P�fB�g�^C�ə����qb؄q�j-c��=hRC�2l��`ҕO^������:�tC�	;��@{
�	�-�ţ\1\ZC�	�P ����*)ät��A�x� C�[rX)���4 [�0"H��/zB�	�`�n�����Wܸ!�"�,"��C�	:Xdi1u�G�h{���F���:��C�)� ����S.n�dH�G�,Vh�s�"Oa��E=� �q���=OX+$"O�ي#dG�AC�tѐ&�7���Ȅ"Or�x����W-�س&��I�$��F"O܉�P#
�8n��!�Z�!�洲"Ox�����.a#��9㌇^^�09�"Of�`�Sڌ�(��,'iz��f"O��VO�8d�����M�}U,��Q"O����������-JiK���"O�����Y>S����	��0Ry3"O�487)�[ �r4o�;��8`"O�aЮ�.#D53���x7�'�ڦE ;P
�]���a j.W1�A�� ���;减�Q�qO�>1���^���7����j1�E$���� +y�c?���*Ս��t�P
ro�8��'�<��i��UGα�Ì>,OPH�Wd��tܐ(�q�ڮF}ƥH�D4~G �`���3c��b�4��b?1��E�%-��ↄ)QA(U�U7,�����*2(mL����QVx���f@5lJ���+j�*Q�Cŗ:k hI��;i�n��F�%<Pv���� 6lF���'�,�ͧ���/�@���*��?%b��	 "��	Zq.myD�x6 �2���Q�)y(ؓ���b|�ىuJί3�r���
H؄8�'px�D���l�౉.Ӈ%���pʌ�{�ƴ�OP8�A��.�A�R>3;�A����s�O*�R��gFR�Ņ��/�Eb��'���S$�<^V���X%G*џHB6�Ew�b���-�0!
`�a�A�&`�T�9�KW�=�`,3����%�b>	�@�!�x��DU`z��g���8j��
��7�daE�|\�=)�$�Wav��S�X�p���2_Є��SJ�
=��A��<������?����s�X�Z�p�#)Z��*X�?�(�
ݥ(Ty4�E:��tDv�X��!F�XL���>���$�����#�7:���B�b�8^�NQ@A `���f�vղ%��B�A�	m����\�?�O���	��"�~4�,y�,l9�.]b� �(�'n�R��e##?�1��/K�Α8����4G�L2�fx��3��K>w�3�!�kN�	C�Y$s��o�7`�0d��m��g�2�d.A�l#JF?����q�s�6ʌ�i����#H3�.P�%Mr���̈́l����c	2�<x��]>�cr˛�u���%Z�"�(�
۽���y5�`�t(K�[�Ψ��a*�S�n*^�~�4x8\�����4i�z�zQ+�_o��E	2���C8v���o�,1�bT��Em����[��B�hǇ-�L��֠A<r����[D�@:�i�ym��E�ٙT�\	�e�H%P�`�wN2[���A�O(��D B�6{�����+@��r$H8E�b�u�۲{`��
@6��6-�a�]���[zD	�f⑑r��(��7d��8��G�h.9i�Q�FIz ��C��xr��)w�Fbƨa�O�̳�eL;�TZ��M�':�}�qO�<8_̜��iģ0a�&8`��ed��O8�X9%�NI�tr#8_B^����LP5�T�T��&$0v�����
N8�L��Op�H��F9]ADt�AD����"C9-�e�3AE;H��AQ,*4�Ò��:N`��!D���b"�/�Y��9��K�+�������M�W��$�]�7�詢0��+	ڜ���L'��+S+_�����y��-^66���ɛX�&�+.O"\���O�]��"�@��]k+�t�����|/��q��^��ft,@Z�3��,�|e�r�91.��s���Afj�jn�)��;ӂ;?��@ܭV(37������*��8����W�ŧ��e��f��J����Y~ITp*@h^me��� �:����'�ĥ��m�fFZ!J���kXcq ��#	D0�W n!@�+�>i2=�D��w\?5R��D{ ȱ�"E?aw4���#t��U3�4,~�qBD=L�B2'�۷6bju�R'�-N��tiĢu��m{3�'t�q���I�R��Am2Dj���*g�Q$O�
���'���"D���6(: Ǆ�� !K-O��nâ t�����P�>���c�]�u���t�2���S�]<��	�l@���I_�i�^�����C�s�浹ơ��U�A�	3p�(a��n�$� !&;�{��u���hu\��F�&�ʍϻz���K��H2`�]�"I�e��o�t� 0�L�HT,EС�'������P2 ��`�"�P�{q ؼ�~bh� �p��\������K�*��yP2(c$Ѕp�_�;��H�@Q��b��Ђ`�ɉ��'2D.�#�
 ��k֕jdh�"^gr���H��(~6�ҠE�!!�A!F���:����r'B/	RfAIR�U�	/P`MQbb��Dٱ��M��Ph�d1R�lOr���&H d�V�r�C�*?�^��@aVj�0`Ɗ�/%3@�
��ćPr�к��P�7���^�$�ZXXu�M�:�1OX\HU�,��'�TT������;!�(����D�6:����N?1,�R�(
K�ZH�q#����s�R)�����w0�u�fAϕ'Ժœ�/����'���jD�.&P�p�も7�lH��!ЫG?*����2*$pS�|�Z�#R�#
F�8p�5�d\ᇁ��,���M9s)\��
W�N���c1,OP,��k,<�� #	��GW���ϋ�_JH�����Xrm�VF˜|����ę�Z͓�@w���G��.q�$�"´Y��\�|Q`��O/����~W@�wON�O8�12l۵8R����A6{�� ʔA�4+���EEQ3(`8U� �gsdA��
*ܰ?�T��/��dy��ֿU�B$��c˩N� �ʂ늖}�_D�?�'aǭ�8x�.��v#�.z#:M9�'���Zv�V<2�kV� 0pːh1i��f�b��sc��g�L	���z&6?6yݕ����`D�Σ+�6���.H�K���뉯L�t�"�R0$f�����hx��%�7n��P6bBl��V�׈;RDq��9O$��1�z��K��g�? �@���:��y���φfD�̳���H�x����Z�w���Ba�ȂD�WmA�?a:��G��N��$mQ,	Yf��ϊ&2�t@ !J��L�˓�h���O�aXqÕ�Xv
i�7����X����0PU�gP��p�s�+�e�}ҝw���S�!��LRc��o�h�4@v�pBR$�JlQ���!<Oh r�ay�"�@�<�PW���Y �C^'M���$�P��0���T<�e�$N�?J���G�:�;��Z�����EH^�9�-Г�{���Î:i��)q�ըof Y�ۀ!E��7B�b��y��&ѷU��-X�d�!z'�E�Z
e�.Ԡi�8Q�h��%�֡�E�Pm���4�@ru��	�J�S4 ?��?S�-�)R�g��У�Զo*r�so��<�	�	�Ӟ�H�;��_�j�X���j_�~B���l�=5���̓|��m�����B�í���߼�"t��RC�I[��M���[��ʪG���r�d�7 a��� �ɹլ�
$K�/QD�]s�&�����k��K�h	���pNW:p���ף�b�Z�����`��G
�5�1&�	�c�^����i�t��E��
4�@m���N#I��A��.ZM&�(�L'��(-��V�d��UDC1�^]�!	�I��I�i�&4Aw�S�`c���4D��P̊�	�S�YS6M`��L�+��6��k�RAH���Bʩi�e]�x���h&KR�9A,-i�=w]ة��o�a�0�����w���[_w���#梘.Mj�$� �&y��Q1N��p|F�@��T�����Ś���a����T��a�Î�iI��B�ݝJ �+��T�p6�H�f�^/u�ݩPH�:mnB���~�f�Ч�ȃ� Æ&(0�����};�(����idT�J�!��}��q�t}�k_[���¨A<�D���ז.��m��	:'��YDc
��dY��4�0}I�а �fH�ЏQ�/Ws��\�$ |cH�hĺ��"��16��Yb@C%	0�����H~�@�Hj8y'�ؕRt �&�3�d��=7�P� g]-7����ÞM���c��ŏr���RS�_<4�?3�F�p�۟�ؐ�Oͥ>����\�K)B�U�z��� �T�"P"�+w�օ�t���Xڑ#Ʌ)%v�n97������}:-F�@����Ō�+LȈ��S"Z`�l �R��	���R��si��2W6-۩[��r$ͫ�E�
�V�Z���#D?D,ѣH�!3��X3��++B(jD�E�:��$Z�iJ6T�P�����A6Z���� 2�����gI�|mb����Q3[P��Øp��7�*h
��%�O2��@G�yfz��f�0?����=�ӥ�3�$� �F�J$�B�\�8_0�AHS	wc�X�T�C �)����&� �&	K>�� �0=V�����{w����8�LȂb9Oz��G�� K����I��hON�E���Q���__69�-��Du�u�QAy��	"W� �HP\/�vL�#��?����@�>�	W�F�9X�ݳ7Ȝ�m���Пs�0�#Ҩ�:�V,��o� ��O.x0$�ٔ�<�Y�_�~I�'��DؐQ�Pm��BW��i�K�ą\?pBIk��_0:H~�#��v�q,�����؜'���3i��u�k��jܓrD �!�\�r��l#��8;wh�S�����x�K7g�����vC��'r��tsv*;9vd�o��"��a�50*:�˕�[�y��T��(�RTL+�S>]���䑢<�yvD%y���)�0�\�a�Y�a@.�!��K�r%�KA�y
&�"pШtI2�x��D%dJ@�*�A=]�Nu��+̷D�(-��'���z��
�Ym���i�" �~��0�@
9�TQ��0I��x�f�y�������D�d��7o�=�����<�|!�ıH�)\{����ƭZ�!��J�N�F�*q��'�@��i��%��A,Y�9��J�K�R�Xq��
�t�ڻR_Z0&��.;�* ��nX?t���3�ŀ`�6�S˂��0=e�GN8�6%�]%����-U.�M� $D"kT����"�#gl�"%��EL<�;$ur� 2h��]�B�xG��E�PXK/҈T�ij¨�V�X�Rm�5%� ��Q��'��Ec��O�RP["��U�hD�ŻK�/o���c�h1V�u$]�j��)?2��9�pa�TC�ѓV��m���#sH_�F�C��i4>�)�$�?Z�ؐ�B�ZcF�:w�CJt��͹!/�c����k�8#*�E�e�T�u;"�Q���1D��xB	$E4vi��h֬4�l�	%"��h�� a�X(�6mʳB��prR?�I�jU�B�ED�L�ؙ���`2Lz#EO~�a4@b%ϾZP���j�:WDh�@6��5W��{���@Q��4�/FGb��D�F
YhUT�B� �R�ֈHAf�����5AU��;�Bo��B�X�
Iy�Ι�w]�(��Z���|S�@1r���s�eK|�� ��4c$	wY�sU��gNZ:���X���B��FIz���D�d�RŨ���%]�H��|�H `f*T�~7�x�ug�&EAj<�7��'�@|����	(<9���!p'�̠�섖+���`B�Rf� z�"���t�uRR
MC�F��a˙�*X
�&	L)�F��HG�~��sՉ�d��>�R�������3ғlㆡ�DH��IzJ���
A\BM8Ej%z�%�s�E="�� D�W�<Xr��0=|N��"K�G^�?����
�	�b�K�Gx�ȑB���{�j����<@����򮐜 z����._| �{��R�k����4��	�%F�=-w,]�Q/(u,t{ ��_l4��ҥb�����?�
s	��>�4�@sA��h�����M@�;X�!�2���~b�o������"Xf�� ��[Y�ՀV -�x	ⅆ�
kIS�I� �J�ꡨ@'k�YT�M7b��r̔��P��A��CO�@{�Ȯ&�T����%��k �G%�`�~!21'	P2��� }^��c�V q��Pe8n
��ge�:b�jJY+.(t�����v�#� װ>���Dg�.�qC�-_�W j9��9K~V%ɂ�\w�'	�}S�M_2U��d��X@��VEl��}(��i��s1˃Qٺ����4	̂%q���%A�~U��2`Jހ^�:�pQ;Ѣ"#�����V��㟰`�*�<3v���B�&ANPQg�O��p�c�G�<��Q� KZ/1D�:'#F8"�X���K�����d�(u:~�KB	��9��7�׶:Tv�P5FrC>��g� >k#K)%�l�����o��q0b�04�Ήj��^�ٶlN�(.8+��+�?�5n�i��4YP��	6�X��M#gb��"�O?���� b�{��Q0?3�YQv�^�]ϐX8���(Qf
%�cU�I�b!\	I$�VI��/(h V��gBV�m�fc����	�\�R�,�+:��(����+�a&P�y �
DY�����n�PXH����D� 4%؟'@��E���'�@����P5�`��ѕvL���N��tL�P6�N6S3Ui�D ��$K�@��`.�\{��rA�����J�X���P2Q	�% ����<�J�SSb؅�|U�<Ys��n}R�n3$=�3�U�7&�U��h�$$�|5y���(T��2(0���֐P!lС��D�L<�R��d`~)A��G�y�89S��D3*0���Q"��8�JK�@���zc�%}ȥJV��7���i��1[�h�����f5��(�ꋚD�����J'yƹz�̏2�� (��Q!�6Rָ�႗{'�x�B� As��M
~(p�Wb�.2�D6PԼ��"�D�b��ǡ�O� 2�������FxFi���Oܕ�'�`��g�T'I�4c��z����AZ�o�4�bb��#��-ه�-I���_^I��d�'�t��<�5�<$�`���iT72���)�LT��f&��]�tSP�#|��)�d�og����oV� m�qB�IR��vf[9_�l!#��џ&v�e[$.J'?�T�Ca-V�{�`}1f�;�	�z�jaq���4C�@���9�ry��M�c��usT.������bv��ra�z[nр[�?�y�0�Of��B�H�E۞��I��':/������J�ظQ攨-��I�c�H�i$�5��@K�l^��Rk��{�C[
d�>�R_d	��w�`pH��3����G�2U��ٴ�5�c�0�)�禭�����=~��TmӟZ>�H1�E~t��s��2H�6��� ӈ�^���'ǋ8u�<��-R�_*�AE�|vl˧��).m�0�w(P�$��1*�>LO�d(��q�!��oZ<A4rɂ��8,!(<����c�tXt��/���"�/l��y�nB�bղ�����>Af���\�4�"��wn�YCU{̓vd��h�bK�ըC9"瘅ig0�T�k�@ 1�PUH�j��U
n�1�� �N\�K��f�� ��Na{2�C�C̈�yQ��"!�iKm�h+(,`��V	Bb^�UѠ��^w %��SN���mT6, ��� �Р'��T*q�Q������+#XC��I��)S�`��o�L�26���}<l؁tKX3 �����D�d}�'��L��!  �j�\�v�Q�|>n�ӻ[��aA��ĖG|�� ��Q�]����.F�0oG�f)�w����n��b@�Ce��j��]�6�P�"0�G�(�%!dF�,5t�E8c�4��{b��4�ðo�>0DV)���G��'��Lѷ�O�p���ᐠ]F��r��)GK��8o�E��f�v����q�4��#��cUIg ?\O2}� V� ��S��+Ѥ�z�BӶsj���m������|��'÷
��|��M�,����\�Mf�@���
��hH��B�I*68���rI�$s�\|�b�X-v�6�H�.��A"�&+��:�Ҩ20���R�i�&�����
A!8-�f��*u2�j	�p>�ĉ��$1��	)rO�Sf%,��h�KY�k� �rWdM3a��A���'��%�f
1�3�dD$�L�	��@�X��eAC���d�&rƴ��G�
1�*�kg�33B�IB�L�;r$�(�/����=���>@�ոChƯ,�ܠ���Bx�Шs膮/�Ҽ)�da��&	̢"r���A��M��]8BM���y���)J=�2	��9hn*�OG��'ij 
��q^hU���ӨJV�l��bW�M��p�P��S��C�ɝZ��LY#K��N� �!I�M��ѱ�i�4���'���G�,O��)���V���p�FS�iB ³"O��Q2m�D�<�s�Nߢf����'�D Q4��{X����֦Tx(#�X�}��8ەA4D�h�t��Q ,\ˢmٱH�L�g�>D�pK���[��q*�J�]���1D��ہ�Y���,I�h�"� �.D�8K�T�5wZ}h"G]F7�j`O*D��a�쒌��Ȓ���  �����(D��1��"1`m*BM��V�~9b$k'D��𡔅�j`��Ǔ2�TUt�9D��{0͐�
�P3pjN�S�\��/4D���ԁǺ.�t��Qf/�
���@7D�D���G�݈��ˁwKX�i�i7D��YC��m*���ߴS�@$#A2D��16�#��	Y��X�@ �0
3D�੆BT�u��M�9Z+^T��0D�H�`G"N�}pЈ��F����.D�T�Ŕ'�D`	�C��Ql,D����Y���C��Z�Ĥ��f*D�H��oK�t��,�f�����B�4D��Cp��0f�*�v����M��4D���d�h���C��K(IF��*7N3D����#K����a���S�n0q��%D��JUh�
BZib��!��A��4D��	Q,T�f�.\!&��'[�D�y��4D���Ro��x�j��Qˀ9�@�c�0D�d�e�;s�P��f	Iv�=�(�ɎNy��@(T��K�T�6a�b� �戏b�4 �CG��,�bQ��.4}b�ΒX�����=���8b������tD���
p���H�W����0bM�)�'Vp��ծ�^w��ʅcçDH>��w%�.\�H$�e�)���/����u(V)Q�����$҅:w�5󢉞�^�`���?yN�Fǎx>�rp�@�!4���I�mK�����ڭ��b ����M�V�PX��3� ��BӏǆG�nQ���@I^�s��4�zhp�OnB⢈�0|c�2N3�u�c]�y֌���S�1w���ȉ��F�$�P����!�"L�=J�ٷ�C�75�$ɗav��A�>]8�%��?��v��*_���kFFD,	�ɤ������j1�$jI<E�$�՚`�܅k��W�C�ly��%\rZ���8Hz !���"��	(�m �Wo���MǧBʜ�*������d��0|���+@�Z�:��޿B��U��@��
D�E-s���3 D�^4�����ӶP��&Ծeo��j� ˚z}�u�!MKxn@�S��)�?��'?������yOP����%�\��5��	k\Bd��$���HX"��	^�a���RQ�&���M�X֭���n�,uKҘ[�� ��@��a�j��ç�ȹ"wd��b"~p"�ūr�� �1�|{F�� 6�G�~R֟�8�a�IU
��4�x���D�"c�VQ萐x�ɄE�a�䬑�`.T؈".:����ۂaω'u@���#J6�a�d�$)�1MЍ�
<X�E	LN��'6j�"�@�%92O�OO������*`m+!������4MҲ��a�O*\�oM/�~
ç��в���Ʈt�`�w�čϓ-��M�p̪��35n<���4�ܯ#,���-\��-YsnY�@���2�'��q�S>�Y����$)�F֧����`!e=�	��~�����<�Oe��c�f=I�d�#r�pU�s��� v!��ِb���RL�k� Q���	�6I!�$ڤ�P�F�4i�ڤ�ͮH�!��'t�^�8�K�,Nڈ�7�:z!�D(1���h�O5PAPm�3F�?o!�J.@�)O9H�|�f��'kc!�d�<���y!NX���p83�R�_�!�DC<���2��3
�,9[t�L�u3!�$�<q��A�/��=ߨ�����5K2!�D�*��bbET:��PΐG�!�d��1�F4�P�@�%�B<�s�K72�!��ZP�@C�e8x�!H�&��#�!�d�s�HD
�mK*e��[qf�'�!򄞻_f��L�?+YQ�״"!� e�2�(��6���c�N!�E�P<)�c�D�@�^��Ǟ:!�_�cbų�M��:�T�@�!���!���Y=��Q��&az\H�G)
�!�DѮ{�����z.��.��c\!�d�Bv�P ߀i����Ԃ N!�Ė72�"D�u��,~qA�H)�!�䚼O�,aɐ��
wb����	'j!�T�j���'%j���c0.�O!��E���mΜf�����hU�C�:B�ɫp��!s6-���W��hB�I9D�40���s�H ����TB�I�M�����Z$f�x���"�rB�I8p� �]j<e��*ɕ3�jB�	3�$�[�'�'���шF!	�(C�	�?X���Eҧ^�c��5V�B��)V�48�� ��L�a�*��B�I�Q�>u�H��HV�̳ma�B�	L~���F�x|�&Kw6�B�	�NĐ��%�1H�X �%ƛ-\:C䉋'�!ȖG�W���� -���tC�ɸ!��D��+f��r3 B�8k��E��ĘY�u�-Ha��C�	�F%	jdm@%��Q�  �;y��C䉋qi�02v����Z�V�xB�	X�v� �C�5Mp����WRB�I��I	�A�'<<�C���$��B�I,h3�4������=��J����B�	�Q��q+`˗�f������ 2 C�I�B?�������Y�����tC�I�}�l�0�ƃI*h�� Ɖ~��C�	�z$YS	[%I#�{@ L" @�C�)� ��!5t���>a�8�"O�][�iwv�x�΋�PU���"O�<��"�?l(��]�GF�(ad"O���Q��t��]��K�1F��H"O�0��&Ӄz�8���ʏ�I�@���"O~Q!�b�E�P1CD�`�$��"O8�rԈ�x�N�+bjD��S"O�0�=[ ��L�xƠ�"Ot!󀌪y�f����̹!ݢ��v"O8ݒt,�0`9�p�A�M[�.�9�"O�9�s"� (��5Q�НD��-I�"O2] #��#��������f��"O�s6�<���sf�ԭv��xp�"O���A�E�tZHD
\�4���"OV��ġɔ#�$��MP�c~�|��"O�EpЌ��mHtA� LĄ x��3"O�T���6�j�YB,�S�.�1G"Ot����K�U|�P�*<i<�Q��"O04ۤ�ƟA��(�oHGT� ""O�II��^�K2Bm�N?D��"O�p�G��`���IW�Ky-|8�"ON�s�BC�e4ҥ��Ù�"F| "O���G�ޏ6)��IA�=�8q�"On�[c��&IUH�Co�'2a90"OT� ��;V�X�q!��m�1a�"O��E�I$ބ`'N@76 &"O��3��=Hs���wLαy�L�2B"O�L3WL�2E����Iu޸��"O����!��c�M`cH��9w6��`"Ol5��$�7�-cr̎� N	ړ"O0�Y��߳J'lZ/R ]��"OT�5�<6�;S�/e�M�!"O�	Y��A�$k�j�)U�L�F"Oxu���5,��)93��;S< ""O�Y���M�i�FE�'��;EX؈"O�<�cF�o�`E��&A'E�XA"O�8H��J�!��t���65$ތ��"OD40�%
?x3�)��I��(� "O��s���:�C���г�"O�ȸ7��xzൊ D�)]�FH
F"O����E�h�n I�c_�0��B"O0���jROy�Y���� �%�r"O��@×p^b����E�@��e"OrUj��Ԓ,j�-a���"~�0�B3"O�x&�Q�aX9͹J�bT�G"O���C��~�
`��o)o�ٚ�"O�4IB�;LB��P�%.qZ�{P"O8�
D��tUtx ��V7"Cʌ�4"O���v��n\���&���_���!G"OT�@d
��X�"��Y�k:T"f"Ob@���œ2���:a��#���"OX���]5;��0+��X�]\��P�"O� �d�p-��Q/���3A"O�����եuLp����sԔ�s5"O�L���S�H����恅|�ܨ90"O�d�w��Ff�3� �<�!"Ov�`īN <\8�B�P���	�&"O��j��ۅ=���Ibb�1$g����"O܅����o^���0��fPD1�"O�%xB!�.,�(�2dR�.Bn�a"O��c0�v�L �J�wN@�"O�͛��Y
%�R⨈3l�bX��"O�E�s+�)a.��1h���S"O,9���>>��ɴK)s����"O� �]IA�գp�~��q�{��9��"O(x���n$���E	/?�BM0�"O�`��Í_���r�dF2|uj"O }� ��N~��Zv�B={�	"O��HG�H�uN�<Bs�g����"O��EV�y�d0"�N�/i��7"OH�Ӗ�*;��;�F"2X)"Oह�&VW@ 9
w������+D�D�4��-R��qzr�μ��� 4D����̄�ZQ~5�2�߻- ���)%D��0��֙{Ȥ@��A�1R�L�"a!D��9ul��`gV�j�'�P��9��"D��y�T�".��(ۤ#n�q��?D�@��ȃ� Wn}���/�����(D��b�CL<�2�ە�
�?�q�(D�t���ǯ-�~��Q
3K�Yk�1D��3����jyl�؅�F�v$�i*��-D�dCqK��q�hI��~��@ D�4S�I*_���d�}�p�2�?D�h�E�A-|����C�	ez$���0D��X�B>���Z�lB& z|�B�+D���F�ԥ�����Z�(@pP
t	7D��	7�8L�x�b���34��c6D�P)�k�"�p��W�D,j�� D���d�˥?zP�iR+h><�9p� D��Ӗ!�_= 8���3N$���<D�\9��.,�>t�MP<zb�{#�;D�,�� W�Z�Qֈ�J�>�b�%D�h�!<ޖ�G
�+A ܛ��"D��1UF�[�>Er� X�p:�i���;D��Xd۬(C�� 1�Ȋ���,D��Nʮ	v�P�e�C�Xm���8D��0���S��P 5�UE݊:� 1D�x3�a��f��*�ҹ!�6�7d4D�`P�L�TX ��N�3�� �"-D�h[q^k�N�$-�N�����7D��C���	w�j1Z�B�w��d96$;D���c# p��xS��9Q���ul#D�,I �	"�(1W+OF���C�<D�x6O�>?e�����H���
�7D��i�C�K��9�WB�7_X�!�E5D����D��H�4e�b�4���G1D�����)	%�=�0 T�r�8(Pl$D�|���ˉE�����O�(�W� D��9ry�d@1��=P���@+,D��z����ؤ��Q'���ұ�&D���5f�f�ĊS�ц.�,ee?D�h 4I=]�6��a�N�"��`)�#=D�؊5�кp�^X�T)�&?l�� �<D��
 0�`��	!D�P��2�=D�p;"�`m�5gO�E:D�T�&J�<�:=��T
-����+D�<[G�D�9Ÿ�82MH�O�ze8Qk-D��R%H\�(.f��F�p�zi���+D�Ȋ!�S7{�>�bũI�p<(���<D��ZC�!���k��1��C�*<D��zD���+ﺜ8�.����(�7D�Tc�g��)9�V�m�X�{�5D��Q:XsH�A�-j�8�{u�5D�<3֤�X��hyAAӃ�(���j1D�� R�Y0mGd���{��	��A.D�4a� �;Ԕ	j�؝E�v��E-D���R� �
�������f�Y��,D����c�+$n�Bf�߄|Bɢ2�)D�� �Q	ui��F�P<I5���b��ak"O�2��������n0|��"O��1��a� ��@
 nYH�"O�@2��5Ɏm�%'Y2�x��"O�	P�Qr�v���	��Lzy "O������nx��c)[����%�Py�NΕ]n��k��Wp|����X��yr"P2\�$��@n�la�аa�I!�y��N k.�O�	fBz�Y�̠�y���/0w��b���H�J�fJк�y2*J$y�V)5)�Fu�(�MJ��y"�B�w����'�n��(���ynڱa`�1*�.�<2���E����y����(�&�Y�9>�yDf݃�yR�X>	b������0��D�R��y�ƅ2e6�uA7��h*���c���y�(/:H>\K��ٰb3`q�q"��y��HƝIB.�^�~QRԆE�y"���U�D��(V�f�i�-�ybF���x��n�a�@�*7�L6�y)F�
�ʅA�f�3$��������y�Q�Z�\{��ėQ�҉�p����y�J�
h��L������yA����Ex5�[O�:��gG�y2�I2 @  ��     �  d  �  �+  �6  �B  �M  �W  /`  l  rv  �|  �  m�  ��  �  4�  t�  ��  ��  E�  ��  ��  (�  j�  ��  ��  ��  ��  ��  ��  � � &! �/ �9 X@ �F �L /N  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|`I!'G#\���%�T��'ItcbꀀK<�k��̥:O��'������Ǝ8�ݓ���"J�S�'y`=c �d���	%�BPiV��o�<)E�I�M��c�Q'��I���k�<Yb�`��s4��/~�����M�e�<Կ��رD�E�?�t�Жgd�<��j�aZ����Aّ'�F�r�b�<��"���e�ďfe��ѣ
�[�<Y �{�<Ԑ�[�0�Rѳ6aE|�<�ǆȕP�,x��H�o���ۀj|�<��\��!G	��lhP�qI}�<�cێ�,����ޣ��@�#��x��G�<��Fъ��u��Z�JQK�%v.1���� ׋� ^:�Bэ]lr"�&���I�-4��Bbʴ9[��g.A�$&��$@?�vĥn9zt�&D��v�����Z�<�5��@e�
I
p%j�a�L�'�Q?y[��Ph�d:�
�Z�bg/D�$2��q�HÄG��R����I�r�����䕘!��8r@�P�Fi�	� ��!��̲��u*4%#\l􁦪��,�du����	�j�����
���k�h�7EB���˃���.*����u$ML�BQ���C���C�I
|����d�2�y�e#Q�B�	�� R��g� �t��B��1�s�Ee� "<E��'�����?l�i�|����y2�6�Şw}��̞�� `�d�ǁ���a����dE�D��p�i^�;>��S��%+�|�L3}2jN,m��+�lRu��iT�y���>�����Q�g�عQ� ��Mˌ��%��|ph�9IV��1�!�;qu��UA؞X$�>�XR��V�ԎPԜa�g��:]&���d(8a�МA��řcYx�h�G��%ڧ\�ƠB�!3]��`��G�44��^�Ȅ�-J�S�d�Ӱ%�'
<�'Bў��$��Fa�,ʕ0�i�9j.!�$�!i�;��@�f�I�Iſ+� �牰D�-�Dk�;�Q���c�C�	;<�4Qd �
����'�4��'��Bm_�K;�HاA�H5���|�����Hȸ-&�tbr�Žp#��v�/�yb(Ͱ6��9�L��o�(��^��~�!�S�Oaƙ�gh�[8|`c��e��e�'% �;?ʡ��� J���
�'��s0i�3y�Bd˖��Vy~9�	�'�F��A�^_8@�D_�M}F��'����7�[�Y��:C��JF���'�*ex��N�d�B��9;� b�''��SѪԮ4	�#"K��7cL�8�'����d �el�0J�g#����'�HS��Q��*�р�	����'a�|@0l�9�0�p�A|�`<��'/x2���93�]���:%���`�'W��P��҈4�����)뎨2�'R2K����y(J�0�D�Z"m��'�~���j�$)ԡIg�0����G��O����^�E�� �9rdx05$?��{rɚ��I�m#��Q��Lm��$*Ǹu��ʉyr�'q�x��H��t��ѯ���r�H0ND$��=�3U����"��M�霂���.�69���ȓAR�L��/�B��ǭ��-����=���?Q��Ӟ6 ʝ)��^�%x"T�&��~�<Y���7?=f` ���4~D|9qM{�<����J�Fa@o�`Ѡ�sS�Q�<�[y|�d[� r:���`n�EB�`�'F�|�ڮe��)҅��F��b�O���	^���O(���b�>�bI����O��p�	�'eF�Js��#y��L�Ǆ�U�
yK�}�x�鉷4��9{�ɐkL����N4Z�rB�IlZ6�+l�	<�ؽ���Pdֵ����'] �cV�`����jG�%��9�'jX-���_�"�ba던�Da	�'�bY��R&��l�� ���$��˓�(O��5,��N�R$�7/T�j�~�J#"O�BS�]9af�K��G�Y;b�s���=lO�A��ydVEk��ה:0��"Oȑd<$�X���$Υ|����"O���t.R9ǎM�1���S
nj`"O�:AJ���,������eh�ha�"O\�!��שn=Ҍ��$�	'�<Y
�"O��#@E�U��C��W�9���"O�؀�J��}:5��k
:�P��"O�D�G@فE5ZA�Cj`D����7O���df��	Y0i؀}�~��)I�5,�,���'���ɉi����AE\���z�&I����5�I�|9������?& �S &�T|�B�	���0p#� ��� �<}��B�I�Jz��5B�% dY��T�A�6�F������ ��A��ƛRTV�BpH�>���6"OL�ke�I�Z t�A��V)(��2dU�p���h��Q#w��
T�� s!�F�H�ZC�I,A:� Iv�CQ��2�iħX+`B�8P��(��_�!�l�s�H�3
R>B�I�T=dX�!��N�ZAz���._B�	,$��rVk[	l��-q-�)
B�I�e|Lru���Z%��� $��>r�C�	0����ThW]jP��-B�6Z��#��c%O�>�ȉ0�F.`�����4�O��$�QԅƪuJ�AK����>���0ƈ3D���� 	F��AƂ�5�a �M2扃5���?�|b���b�c��$��iIGhd�<�0�� T�4+	I����a�`�'O�yB	Q�$�� ��>;L@�cc/_1�y��%&�&aYF.đ-�E �Ј�y�C���v�Pg:��P�7J<�y�n 'Ǻӑ%�0�؍qbC��y�ώ?~�Pt,(t������	�?����v\8���,�H�Pu��!i|���ȓ@��-Ӥ@+n�P�Sd݃B�v,	��O�����!3��q9�(��D���fcҖ^����)"?��,�;�2%��۷�����(�f�<���H��z�eZ�j�
1I�<��l����v����¡К3^lm��	�!n��M{�O��e�k�!�"��"bN؜�"O$Iǣ�W�$�����w���S��D�O��s�{����P=j��1���{�|x{V�D˟̄U24�K4�ҔT�X��CDP�(��:g(I�&�ݱ*�������>�rԇ�,�*I�K�J��f�3��!�ȓ%�M�adT/J�������n4�ȓ�Jt�0o�zB]��j�b���^=�P������[Ôpc���ȓSܐ�bɇ,�����ODN�ȓ&��MJ�� m=j�%)F@�م� �]Y�Fѫp'T�C��J�[@�ȓ?�,�B&@�����1FTl��b3�Y��N��z�	d�.n�B�ȓ9����[��䪧(Ų!xPl�ȓI�@��Q�(]�r�I�Z<��O6�dұk������@�]�(��׈��H $��<1ѧԗk����n�hU�ݢh"69YŨ�<�\�ȓ[�p�Q��L�r��a��_p&ȇȓq_Mb�o˗%�@$�+�# �����<_p�+3
�h�F@�3$����@ua���7���9�'A.S�\�ȓ:����<%�.��P)��(����|��6�Ѯ#���ޠg��=�ȓ-�E�� '��ߓ4�� �ȓ"cr�@�0!{�	�fΈ�
@�T�ȓu+�,J�$��P	�)+vN6Utz��0܅�P/ٮr�\��v!�h��x�ȓ^��`�$5)x,�N8�f�ȓz� 8��O�]1l�RT"�39���ȓ{/������-��$~(�ȓi<ش!ĭ�_<"c/ק!а�ȓi�Y�&T�w�^��n�%4P��ȓ*�f�K�JB�$
��R�ĩ�ȓx?�W� ❩3 �.��\��`�Y Th.���)˯vD�ȓM��R��+�:v�Փ"6E�ȓz #U�$ut�A��7-�4q��S�? ���*E��t��Ś���(&"O�"&H�8��U��e)���u"OnQ�A��r<x�D+^�@:8�W"O�h��&Y���k��N+/���"Ob�p����U ro[�[Ά�[��'��'��'��'&R�'�R�'Ӡ���J<OT���ʗ/p�4���'���'t��'�"�'A"�'�"�'�4�Q*J�$BLc񧆈aR��!��'�"�'HR�'��'42�' b�'���D��'�� �1�u�3�'��'���'���'���'���'h�v��k��<"#��>2\�E�$�'���'���'vB�'R�'E��'�Dm٣��"D*����Y�r<�f�'���'���'>r�'���'��'&����
���`}�&�ȐF.Jp��'/��'���'e�'1��'��'"�����5`�P� �R�F�RC�'Z��'{B�'>��'ub�'�r�'@����k5c@�A�*�-5������'���'�r�'e��'or�'���'��)�ը���e��Ȓ?'�=�F�'�B�'�2�'#B�'7��'���'_dQWhV gg�0S�M��˂�'���'%��'��'Q��'"�'���AЂ��t��!�,�W�'{��'�B�'���'���'+��'u�� coK==�vlz���f�R�*s�'���'��'���'R�a�����O�Ձ��	{����rrgjm(*O��D�<�|�'dv7��%{�l�ƀ�M�hX6�	W�~����d�ܴ�����'���FnM2]i���5�T���*G;��'�:���i5�	�|*��O��>et@2`�h6�IC��s@��<A���$)�'~K\�9���[Uz�	6iǃfc���&�iW6�J�y��	����]2T����l <Px�G[�s�$�I���ϓ���i��6�d�����	P^j�p��?6���S�lc��̓"I�~�����'����J*�h��q�
�#�Z���'~�q򉗤Mw��N�	�|��(_-��h�c>����>���?��'M�I�F'Uc�M�7h�X��E�ԢQe���?��۰Y�Ȝ�|���Oʜ`�z�:��/F	������G�&Ѫ/O˓�?E��'�bi��	Us�ZȊ�#�O�xi�'�b7m��r�I �M���O�P�Î�3x��Ǭ�Gঁۛ'�"�'��$
��v��T�'h���O?Z��B�{��	B1"��;e��'����$�'z"�'���'N4��� B�U�ȑa@)?�9IW����4e���)O�� �	�O��R��T�Ttʓ�̽6}60 ��M}�*s���oڇ���|��'��2o�S�]QsF�Z$"5i" �6 #�հ@OS��� H�Θ �B=֒O�� r5�E6��#'mF�:f���	��M�ЄV0�?�$Ѡw5 ��6��&�"���I�!�?y�i��O���'�7�_�i��4r��(H#��aU��*��Y�4ǔ���b���MS�'�"㘥8���S>p���?��_cpv����P�����%�z�����'M��'��'7��'��O��1;�'�0X��f5V��].3��=��'��Af�˖�3��I�T�	Uy�AѠ)�8�J�,�1��B�#7Xg}¦|ӎDl��?�x��Gɦ%��?���^h�P󐥂�Z��U�ԡ3P�wn	�Y�������O�n�?���ߟ4�� ):0 C��up�1��]�N+�heN��Ok��ɤ\�"4�CM )UC8���џl�	�M#��&<,��X;(G�s�`V�y0��ϓ4���_��yB�'"�f��	Q��]k���OP�i��W�Q��s�i L����f�G`,�xW�8��d쟒x*�D0�O��R�K�J���prCT��2uc�D�O���O��D�O1�
�l��J�l>��#�/Y��ԑ��A�/������'���o�,�R�O2XoZ%�t"���-���Kŉ��SX�)r�4P���MS�IN�f7O��$�!0T(%��'A6�I�<D�3=Ƥ��plԅGfJ}���D�OZ���O���O`�$�|�̏�Tl�x0��ڿD�⑑�É-^Л�dT�d��'>r����'�X7=��P��ǇK֩CEOۢ�f�Bh���شw鉧���O��Ԭ��s���>O�	��-���T��Ân�bpw7O�Щ�-	4�?,.��<����?a�兎l%*ёP��'��i3wl��?���?�����Ϧ�*��S��t��ƟL��(M�h΢�3gCQKG� �����'����O�ToZ�MKR�xr,�'Y��(v�$^����Υ�y��'�N��0�(\l�$:eX�h��r��!�i�bҦ��c�_6N�X[�J0D���'"I9 �Xa6/۞RTD�(�e���$��4�a����?9R�i��O�N�xC�!��ك���?4��\��۴U��v��s���2O�D^=&iX�3�'wC������.���.iW�`(r�&�d�<����?y��?a��?aD
\���	0��.{��d��?��$����FMЂ*���	�?���PyB�� RL��s)˨Y�h��[�d]��5�M��i`�7�K���?��S�n��0�'�%m�TC�'�/:���ք����N>dvčA�y��O�˓l��L�ER��tnV.j�ƈ��I.�M�ej�?1��@�a!Є���Z}L�����?C�i�O���'U�6��H�4x�r;���,x8b�N(V@����'�MÞ'�2�
�7�>��S Y����?��\� R�;��x1dn�	6��B�6OZ��$��(=���цܭDϠ�#�)
c��d�O��D���e�� J"�i��'��ęf�ŧ
d*�A�	�7H�D�G�*�̦��4��g�M�'��ʈhBF�2E�x� 4(�lA�=*���&�����|V���	�����ҟCcٗ^����r�=:�ؼ�㈚����	xy�,m����O���O�˧k��5��$��lА��k�z��'���[��v�p��&���?�g�X�L�h�c�	$1t��Sg�qΌyZ#�V�tE�'\���Mǟd��|b�= 4m�06�$ ZIO�?�b���O.�D�Oz�4������I_B�S��ր�lZ��e�ײFٶ���D�o�8!ȆU�(�IB����$�'-07�B!v�
�t��[S���Ѧ�	%�nڰ�M�&�E��M;�'�
�37�N�_���H��'"����ύ>):��DmM=��lb ��d������ϟ���^�4�t����6�ش�����3`�ܙ��i&d���'7��'P�O6��~��.��Jpn�W� e��J�ɏ�7q�yo�5�M���x��$��5qƛ�1O�D*�&�2.�j�ЯՈL��%(�0O-�S�-�?9t�2�Ģ<����?Y�a��wʄW�:3GD��c�?Y���?����d]��eR�/PyB�'Ъ���[�SgƌB�F�; �a�����Y}҆{��mZ���[��4��ԖP&�\��lG�^�`p��?�d"I5sYt�1�΅����q���n����j�Z�c�`Vb�@��Ѕ��H����O$�D�O���(ڧ�?aTk�"Gǖ�2*�0*_\�:��?�?y�i���f�'�d�\�;�4��@�b	6�`3�Ԇ��x�<OVpoZ�MS��iw�͡��iE���OXa���&���K�;��хe��k�c�0�O�˓��O��� �8|R�Ȼ���1��D�P��`Y�4X	:8����?����OZ��@c�_3k T�K&iHC-���w�>��i2�6ͅR�i>����?	Ǫ�����='j���/D;��b ��Myb���	K�=9�͎o�Q���b���ܖ��A��sdyk���5N��1��8j�X��L�4m�#e�Y��<�&��__��*G��&>	�f�&*}�)5�^�}N�<iu �a�Y��.Ò/�����Y
-��R�=P��B����ɒ+B"c��t�_/It�0���S��}s�a�3�`�7�L��h�Z4/�2-
Ψ�S���r��$��
���j�2ag�Ѱ	K��C�#��x�)u�aF&�dh��2��. ��i�5pH
9����"/򽢀�ty�ǃ$���R�F�*�����J��x��#��t�!��r�d��O&��<��O$�$�#]���J}8����pc��r_��T��>����?Q����,�y'>��@��X���i�(e����r%X�Ms��?-OX���O��� �,W�.48��Z��VӳϏ,!$��oZʟ���jy���>d����D�k��Y���B�	�^�1��G�6[�4�	Ο�P�h)�Ο4�s�N�3�"�PH�E%h��A�iy�ɰ_o*�I�4��S����!��D@�en. �C�1�Icq�J�@u���'s2���x-�i>��	�?O�<	��ܥEYl�H��M�Z<�E�i+\ŲTEk��d�Oj�d��ze%�擪%FznmC��M�MGz�R���M��JS3��D�O*���1O~��W�8}F(�v��zO&	�T��)5$ml�ß����*d�����|2��?q��y_�,j�
�;}k�� ��
;�	����ɰ@�Nb�D���0�ɼ/^�I� �,�����.����#�4�?�֫
R�����'�S�Ln��]���z�Ǎ�q��
�K��M���=����<����?����D�N��9q�E�"Ih�M{e�ۄi��J��ES�����	˟l�'�r�'qH�	���*U����0�P1dT,��'���'�BU�(i�mD*��4��1\@p�s��^a2 �������OB�D�O^��?��Y���O��-j��̤@�N�3O�D�n�Y�Or��Ot��<�@Ɠ	��O�ژV�2R�*�u�әZ�ޘ`6�gӊ�d>�D�<��s�'���K���5��&�ӖFČ�lZꟜ�Izy�&�G��0����k�G�+"���A8ig~�wD��G�&P�L�����I�2���4�s�� �q���J5 ��qF��Z� �i7�&A����޴%���h������<T�U ǯ�+GdB��e�Y���'�ҁP
5"�)b�g�	�kk.�
�fީO/b�d-	<R�6-��u ��o�ޟ\�Iԟ�����|ri܅��u"G
Ʀ�2�~h���??@��ٟ��I�?c�\�I�}$�ՋD
�^(����.r�P��۴�?)���?��Y�v�����'	"*��;�8�S�պ9-�X{b͛���?y��F���<���?��'�ڡK�&�j��h1�Zut�Pش�?���З���O��$�O��ܺ
;~&p����8�Q��>y�JF/?{�=�'���'j�I˟�*���{��f��-8H��і�i��t�'���'����O]R�s�j��1e�ac�k&��А�����ԗ'I�М_��IJ�`�X)Ec)W��lK�K�e����'���'9�O��DU2HSj�ie�i)^YQ�ǐk옼+Ђ��U.JT�O��d�Olʓ�?�hR���O��Y`jY�^���I� xѰ��%oݦ���O���?���]�.��$��@AÔ�u����t�^�^d���v���D�<)�;�B��)�|�d�O<����'��	H�oʃyS�x`,S�?����>��[r2��ώA�S�T%�-"����dV6ũ �����D�O2����O��$�O�$�J�Ӻ� T�c�� |��ː)Y*a�#P��I�b��5y��<�)��3
6Mr2(�)m1���Q�'��7���IO��$�O���O����<�'�?!��C6!]\|9��B����s���:��(کآ�s�y��)�O
tRGFO�����"Xy���%�æY�	؟4�����`�����'��O��F��s9�J��~��@Zwe�n̓M��u����t�'��O(��t`�(+C�ub��*��p�r�i�b��"P�՟x��� �=�eج�� �R��i6]+U$B[}"J)n�����O����OZ��?�n3n�Ti�B�Т]A�H�G+V�5k.Od���O���;��۟x��薍I��l���p�����Á�u��%c��7?��?y/O��č0 ���Rע1�����W8hp�"L�Q�7��O�$�O|�`�I�2�����Nk�pa�DJ����]���8a%^����ş��'�a�;V�S�@"��R�<����Dߕ����5�M#����'%�N��E����O<����2&��!Q��@�4�Ȥ�Ʀ-�Iry��'Ɋ ��]>9�'i��L��S���@)ȵ�(��&X�R���<i��x��u'�:@_���)���T�`����$�O4Ha��O��$�O��D���Ӻ����uQ�	¨}N�{%�Tx}�^�`Q �/�S��>Y�=�WnbqF��Ge��s�7��J�z���O�ʓ�b-O��O�3�㍶�f �����2lQ`�l�q}����O1��$�6$j�MS1��)\'l��6-E�R��n�����'A ��V���͟��	\?!�k�"3�"5#�M �8����MD1O�]�-�]�S˟��IS?Qr���Jp�FP��(;�J����I�(r�L�'3��',2���E�.mZ��&T���(2F�`�I��R]Y 9?!���?+O��dP1	"p�� �+�h�����m%p�0 �<���?����'X��Ͷ��4�5	H�RK���3�5V�� d������O��Į<Q��m#��Oc�� C�:D��cL��)�۴�?a���?��'����W�'�M��C-"$T0Q3�b�3�U]}R�'@RX�|��� j��O�¡V
|�pL)R+�/2�(��P�Q�6M�OJ㟌���n�dYW�=�d/h`5`�@���S�� ��F�'5�ݟ�з#�W���'��ONШ���V�K�(�᪂??@���=��ϟ,���G�%��b��}�Z� h��i��G\2�R �'j�g��>���'$��'���[���Ky��D6A��X0��\�B�tꓷ?�v�F�y���<�~�U7Р#'�Yb��袀��Ǧ��F՟<��ן��I�?�����'<�bt�X
	�F�y��=I��aӆ5:G��E�1O>���
b��`��(W��ܴ��6v)�|��4�?����?�ˊ��4���$�O<�ɴi���@!��)�`�h���*��`�y��*�~���O����mJ� 
���y%�G�m6��OR1x�C�<!��?A���'p�kӬǚN�P FK� eҝҨOL"1�G�%��I�H�I^yb�'���*����:#f�'u5ʁS)/B��Iޟ��	����?���<��h���U�no��kgC�p�F�y҅�=D��H�'���'��	����7j�S��IŖ�j�04'��<"�KA�	ۦ��	쟀�I@���?� "� X���m��"	Dͺ�m�_>xa���n��?	�����O���«|R�'��h��H�6t~6�ڠ�ZhcLd�ݴ�?Y���'�Ȍ��\�����hօ��"%�w���`�H1o���'l�$R�[��柼���?=k��̊��gB�-�=CR�α��'�B�2�̅��y���A�i\�p4��a�� 4��Gp}��'��$�'sP����@yZwF�P@@]+=�`��ٵB�HS�OX�$��W�P�a����I*&&� ;��V��3��&x���f�`���'{"�'�T[��S���1QH�K$�aQw�o)��6	�/�Mk��N�S�`�<E��'.5BD͇
QpT�Ά3gyL�a�jӈ��O��$۞\;���|r��?��'Hl ��H/r3�A3�ɽ�`�t+9扼6,� K|���?��'a��a�H9B�P�6�����4�?A�,Z����O\�$�O����;Q�����\�4�j�	gH�>�Q�+�Y�'���'��� [rD@3GF��[�]!uI�䳕���vGp�'���'���D�O<2��G�`���g�]�1-	:!٦M�������ԟ�'5�@�iH�iץ.����%q���c���&zțF�'�2�'��O��	
W�� ��iW����\�w�b{�CT�7E�� �O��d�O&ʓ�?i!�,���O�L6GߓV�㓊�\zƱyq(JΦm��N��?)g�Ů��&��P��[�(�S� K1]Tr��S!c���İ<���P�Ȭ )��$�O��)F�]E��c��H�Ƣ�'I>v��>!�7�f�����p�S��!��|;v���dɣu�p|��N����O�}Y���O��d�Op�D����Ӻ#�/�2�쑪���3}xrU�O}r�'��`�/L����O��uiӏ-&,vu�i�H�"��4����i�B�'�B�O�����L]n��0���<.����Ҝ}��$mZn2\#<q����'�H�K#hF��V�%.� �F!��Af�R���O��$������'��	���S�? ©G�x:$TX��0����i�_�T��@f��?���?G�٬ǆx;�G�"/Aޙ �� ���'OX�QdJ�>�(O\���<�����h��|a��E[�:�H�}����y��'���'o��'��Ɏd�䐀T�d�����0<D|I`j���D�<�����d�O��D�O�d%,ܡ
pR<���V]��E)�b۵�1O����O���<�H����J4'̺�H8>�9 $��0ěS�t��dy�'���'��D
�'6N41�o��T�v�� �>�@ [Emx����OX�d�O�˓Lj��7Y?u�I�A��̺tN�b����
Vz���4�?Y-OV���O���D��[?1�㘨	�&����
>����¦��I͟\�'�����"�~����?���k�6��$�y_��2��m�.O���O6�����IXyRݟVt���Y0��Pp*?�bR�i���{�V�R޴�?����?��'#��i��A�L��dXIU��P�XREzӚ���O���d<Ox��?1���U?t�xE�G
���@ɵ�V�Mc�cR�/����'X��'��t*�>�*O����'J�'��T�]0�
)R����U�Bl��'�H����;U>X�B�ۥa���k�ɧL��ݛ�iz��',�0{�$����O���2'��80$NI|7&�b��=��6�6�䄖2K�?9�������-0w�����wL�=C���WN�A��4�?��cϰ��v�'&2�'yrb�~��'\b\R���)rT���'vR�O6I��;O���O����O���<�	�2�0JOR���<��d�0z%���S�L�'��\�H�I֟PΓ]~�}�B����~]`�mB;w�aQ� u�h�'���'^�U��;�����EL�pm��'�2}d����M�.OR�Ĳ<����?A��-���n᚝#�4b$�x%	у���U�ia��'�2�'��	']�p���~��Ɛ�sg�L�S'�I�4�	�i�zu�w�i�B[�H����8�ɑ)Z�Iu��<`	�!�`��F^��+@���AG�&�'T�X�ȳ,
����O�D���%��(Ggr�I����'r&��Ћ�u}b�'�"�'�RQ��'��'7��2pڬQ9�Q"�lջQ�3>��^�����=�M����?1���zP_����ZM(p �!�Xs��	�:7�O�dœ`��>� �S5G���Qd!�F	D(XGMS�P�(7M+)��ioZȟp�	��H�S�����<��'^Nk��J�-��?��(҅�yB�'��N���?�ॏ&p���ш�	U�!�kC�L���'9��'�а��>�)O��D���#��O�r48����
�S�6�Oj�Kbr��S�T�'���'k��Y2ɑ�-{��A����囕T�&�'S@IW��>	)Od�Ĩ<��{`�D�q���Y��R�V!�@Y���T}�K��yB�'.��'�2�'E�I���e`(0��˶@�#X d��۷��$�<�����O�$�O��e�X+yH��!_�^ä��SHL��������Iӟ��Iiy��B�,�5
,Zp�N-lHaR���
�Z7��<i����O����O�t�2OkV�>5Xf`�?K�&8C@�&/��V�'���'��U�t��˟�����Ok,�	��]Z�N�It���b���)��6�'��	՟H��؟t��+g�@�O�%k4���s���p�kƕ!2���"�i�b�'o�ɉQ�����D�O��ӴL~�ċ��ڥC���@�lP4p�'���'ҁ��y"�|�џ6�+vn�@��)z׌Sl���
 �i��'�h޴�?a��?���|��i�UP�#�������?=�T`�t�r�$�Ol�Yb7O\���y��	B��X�8ք�Qz� a�
6E��Ĉ?d�6M�OV�d�O���SS}R�`xgAʟ?��X�$n(l����/�M['�<�K>��t�'6�TRU�B�X�0�J��R�w�r-���n���D�O�������'��	���������`׭	S����N���QnZ�'���ٟ��i�O����O�q��7�ы���4N�]�AȦ��	�Ʋ���O
ʓ�?i)O���8���N_N��˃-A�w�}E�iI���y��'���'��'(剗&�@p�ݩojfxaf�I8��-PP���Ī<Q�����O��d�O���*§xnD�gh��0!��NY��D�O"���OF���OV�@Ԅ��d4���&�E /�6L��:.^�+7�xb�'e�'_r�'�.���'�d��sĖ�Q�`�9W(߂ h$8��>)���?�����)���'>���n��(	�6rT� K"�8�Mk�����?a�B*A�>9�脍$�+ �.2D�j�a��ʟt�'vLA��&���O��醍V~Z�i�m��b��Ÿvn�\&����˟���˟�&���'op������\�Ҝq����ml�PyB)�C�6��F���'��K/?1�ŝ6P�*jǖW���;Aj ٦��Iʟh¤��$���}��&�`�@A�ã�io� 4Cͦ�fꒄ�M{���?1��R�x2�'��<����J{�i��3l���2�M;��<yM>i*�V˓�?�p��,�rdr�CE�R�u:�#yٛ��'��'��	k�@;����l�"���Ŋ�0x�h!�F����>	֫|��?Q���?�2�Ɍ�V�G�`N��r�b����'�����)��O��$%����0� K1b	�e!�c�Q��\�q]��xdŏq�IƟ��	����'�b}�c��%0$q��c;�(�pcZ=?N�b�@��W���D��ǀ Vl�p!ȑ��R)�t�fuSQ+P�<!(OX�$�O������M��|�S�T' `�'MΞ	�7�TB}"�'B�|2�'�H��yB�s�0s�L��E�}�b��;0	�OH���O��d�<ѥ�נ[\�O�\�b����3�-	$	R<Z*`�"�$#�$�O �$Q�Aټ�d!}�՛=۠�3�36�9�D��M����?q.Od����^�۟(�ӟ=����A[��Yk�(+z��J<����?���^���'k�	T�hz� �4+�:�}��Kh�]����̓��MK�V?Y���?���OD�)G�@�	��v<�~�K��?��`�������OӪ�#�[�$�ҷ)�#M\rEi�4g�pu�i���'S��O�:O���=���ƁV�cL�-�
֤jŴ�l�˴��I�Ė��*��_�$�4y�dl=3�"F<M���l����	��d�c�����h���'���U�pH���f�.e���s��U��Oxa��d�O���O����G���0%��d#� R��A}��A�(k�	zy��'{�'?j��4��`b�IՁ�>`�
9pű>	�/q���'�2�'��X�#�_�	��X�e�0P�2�;����.���C�O����Ot���Of��
�Ƿh��u��IH7H����ri	 +$@'����ԟ��	��p��6���I�h�J�""E�+v�"XD����h	aڴ����O�O\���Oe���,ڛ�˯S��|ru�W%lKls׬(����On���OB���O�P����O����Ov�zSf�ɀ�ֱF�pY�M���d�Iڟ���.B-�!G �$��I*�,�7eP�>�bu���ԛ�'��W��c�Ϟ����O$���f��'��~����!�%7۪Uz�����?qRl�"��'��\c���!�`Ͳx���S���F�ZQ�ie��'������'�'�b�O��i��2��
l��!"C����/yӄ���O��z7�C�<1O�����M+f�d(��A�ibr����'�R�'5"�Oo��4��n�\Q�!G-{Ŵ���Ɉ1l��6�F�8�S�������r%A\8�J�ʅ�'�0�r�V��M���?��"K��Je���Or�I,��$��	 J8p _(oc���+0��ݟ���ӟ��ȇ�u�$�˱f�'�¤�C�_1�M��Y��h1S�xr�'�R�|Zc��)�#�0a�mqP��l�F] �O
�R���O����O&�)M��r )�#+�D�p rr�	�I({��'?�'��'>�'��80����Q� r�k��0ܐK����'N��'�R�'��H*D��	�� c2U�E%Ǜq�2]z�h�(���'�"�'��'�2�'4��:�O�E�`鏭b٢����/>;�P��:��K)u�N� cn��<��e�g�+���4+v�W4ct��thR�7��C"O��b�[8jJ�p��d�
]
��O�@c���@X� ��hiw, �Ӭ�>2Rh�D�p�n��E '�X��;f�I2O;m��P�c�0Dn ���9i��@2��85O>�"'�%*@�s�I!Y�t032f�&h"���b�H�(l�5�G�-c	��ˍ �����RDĀ4��%� |B(���ų(�HC��'sR�'��H �c�2SȔ��;P�N}�ǝ@J����nQ=���S����'���gMT{NTW��I�@D3�A�O�d�ж��)GJ$�S��?)�L�6��6�s9�wfћr���G������ڴb����"|��WL��4��o����s�@��̇��5.v�iW/ƅr��pA��1#<���i>]�ɀ{;ލ`4�V4
�(�!�,Db:a��ٟl2P�XY7B$�	ʟ����!YwX��'u(�f��a�1��)[�% �	+�a�O�ܹ�G��]�~�1�Ө����$��*ot��S*0ehep����Н�?yq!��l��@�����3ړUN�ҍ��JC�Q�����D��|�m�d���˟�F{�[�t���M#�Z2,!��q���%D�4p�Ԍ8"��uf:~ԝB�	���HO��Ny�\7mD	��KabN�5���2���ef���O����Oh���@�O:��d>�K���6)-���?2T�A��G"}4�цL�@��t����Dx����k܁w�Z�2
54��Ё7�C%e�p|�!�AZHj�"PO�Dx�`�!��O���Y\6��@�.~��m B���-:(�=���3U24����0f����^�;!�$̧v��sw"H�t(��Lƚ;��@}�Y�lB�
���O
ʧ1�ม ۟d��k��άGc$@fN�?����?�4�9U��a@��^�.�����i��L4�X�̇�R��4�4�˙�(O ��#�t��+f�,4�' 9&:Ţ#��R�`=ză�3Xt�Ѣ�(O�,#�'����Ł+��hl^*'n�ԲC���I���Q���
3a�_d�C �Ⱥ\�6�3p
=�O(%� ���Q)Z��U�WK�zt���y�P@�J�����O�˧:�da)���?��^���դ��,kv|�"�>j$U�`�4k"ع�`õ��E���	+��O���k�b�NL�A"܇!��4��	�TZ�I
l�yQ��
@�:@�Pl%���q���I8�=���¦KK�۲��x����Iߟ���'��h�V�	�hJ�|h��@lH�2|x��S�? �4b�%\J�Hd!ߟ~���I�ቭ�HO�8�t���˛�u�l(�F�%T^v���2��¥d�>�	�� ���<�Zw���'��H�5�P�@�􁰍=g+.�R�'֜�k6fZj�R�o;O։�q��^d<�ӔcQ"���%�OXI�p���(x�Yv8��H���emܟ>gJ��E�����=g�r�'TўH�'B�h���M�'�F�;BA)�nu��'�d�2T�%;|ΰ��L�� gX"f�)�S�TV��{"	��MSu�Rи�"����p�P���?���?���b��Px��?��O�`�bu�i�B�A7?�Tk��L����F�L/�p>y�!W��dΰ@��)���פ_ݳ���%A�|b�
'�?9$�i�:H5!�yC�l�2��6������s�"��<	�������'u|���b+�IQZ��
�!���;n�a��)>~1*�0 �̕1Z���I}�Q� ɂB�M����?1*�X���;� �F�K(8X`�J4+8���Oz�DCPOZ�ڒ?�|���-r�n�����
?iRe���Yb�'�F�c�E��h��500�*H.��Kbb�6�������:��J��b�4�?�*�:L�ӎ�6(�!��a-�]H���O �"~Γt-�tåw0eXg*�D�,��	���X�s�����l�i7%�R�� ��+!�i���'	�%xNʀ�	��͓O�f )0&�>���`�L@�Dy�.)�6m?�|Fx�,B�L���sg)�� %���I'yϤԳG�2�)�矼�D�ta��eM�#����B-«_C�Y�	ǟ�*���'���6jͲ��4k��E�8a�౟'���'� � �h �x*b*va���Q�����:~PD���ڂx�(��ߕ>����O:Iɂ�
4B��$�O����O,�;�?!�!��P1��̨G���"a�I.G>P��� 	��e �T����sdU�P���z�(((� Y��FJ�#a�����?𾤁�R F��h�'�*�B�$˚xq����O��ԟ�	�<�'�:MGJ�g��A ���
�����';�y��<��A�I�4��B#�瀅	���dͤXf������Pu#��?��i8��4ܚ����?����?I�b�-�?A�����4I6ܻ��i�м@���cm<�p�UR�����vO�=�횫�M��B$oj�	1���MnVU���{8��QU��O`�lڷg.�F+��QḆ�a`���� �4�?1(OL�� �)��M�M�@es���x8X+��j�<I�	���Q��Ȕ"�Bآ��<A�Q��'`�A"Oc�R���O2�'j[�$j� �5���@���`z��!�V��?1���?����z����D���ݮu�І�<_�S�\����@ 6����>zv:�<��^͢#��$���gQ6f�(i�O��di5`�� �#wY�@����$��Qs�%m�T	n͟�OL�0JAdΜt�� �3M�,	��'i�O?��i��)��aI�Z*���E%'cP���O�I�sf�LX���(-�4���E�=�2�I:�D��RN���L��H��4!���t�I����1a���R�����f�&ų�B�"F��(�)�3Z1�hQ��&:��i+���0т��5�rxy㕙%��4<���s��uVz�����2=,L۰/�<-����EE�*�*���)!J,wި���:e1l)�猒A��qDx���'�j�s�G�qu�cI�)��%s�'05	�$6I�áN+��b����F�����'�l�6fF��`�v�BG^0��'BrO�cO a"��'�2�'��"l����� c��׎����]�=i�,:S㥟��O=�Zx���&�ȓפ� wV�t.�OA���/?X���n|؞X�6Wt�3�O�Ƅ ��V���$�=3�t�'�r^�x��I�LZ8�)�*�~\��%�+D����J�0X�4y�IX7Ű�H�Ȓ�HOT�'�򄝆+Yx}o�%N����9y�e0"��V��<�	���Ip�����I�|" aU<B���4le�)��CւW���
�Q*t`����*}���0
����5���v���Q� U*�:�OP���'
n7m�B��`�Qhӳ1�J\9UF=cƵmߟ<�':��?��Њ��>���dF��ER�JbO$D��94�i�H��!Ϛ,#����a��j�O�˓����R���	}���H�!�y������A�$�jb�'#��'��˳���7�b��?0���T>mhq�!��a(WQ�`�e�=�x� �iX��(�7+L�3atX��c���離&`v��3�W��2M���H��Q�8Ѐ,�O��m���O�`t���>e��T�K!vl���'��'��a����g+��AD�N�qz���-���� ځȓ%�7M��u�$���}118O�m��o���	��O#6eH��'���'�<tr��>FD�A�+@_��#�	�w���y�b�b�0�ņ֐�������Ͽr#Ͽ'5!�EEn�%��M?]����iDW��� �Q��������X0q��4�Ͽ+�S>���ںx�(Z��D�2���s���?Y�O�$��O��ð�F2h�`����Eh��9O|�$(�O�Ұ@�0.�W�H8&�	��HO˧}.My򧜓vJ�@��D\	dtR��?�GI�&�*���?y��?�Ĵ��d�O�|h�,	e!<Mz���?yl�3��O��O_�$�,�@�'|:1���K hKU�AjW�}X�x�'܈*!n�B�hR	��:���$$̥ ��@F�REZ��H:��I��~��Y�L�	by^#z��=c!�c;(�b& /�y�iR�+P�l`��-]4���6���3`�"=),���O�N̲���ã��2�ЊU�W�u!�$,�JaY�D�/��Y�ċ�'��Ј�ݭz����@�L>�	�'r�ՠ�d�'�$Cv�,HX����'9�[��ۻ7tҴ��A¦�r�'t�R�Gٿ'�����ɪ��L��'�HL�#��X�R�8c�_yZT%"�'��,豧L�p�4$S�b@z��#�'˪��u���!�s3.@�EM�9�'@ͻ�Cǃ{�j�s�W��HE��'�2�h�*z��r��	_��i"�'y�*Ǭq+��
��^z"I�'eL4ä�yy�L�ыТV�����'$�4(%�L2�)�F��i;�'@ް�g!H�~'
��9<6���'ʰP)�$���,�'��/�Ƹ��'ib�ˡO��v\ 7���/Ɗ���'f�=5jSpK
���V#��L��'���X�+$$ykF�0��d��':F�ir�S�$�H(%�ʏ�de�
�'���a N�:7�����"� R��
�'�<p��IŜp���;�
��B�ډ
�'}�P`Q�1����'� 8��	�'��pz�OYP��7��,ZN %��'��b�U>5�6�E�Pr}c�'T�!贩��@H��3V��Nш�'�b)��V��E� Jb��'��P�Ǎ�@���a�ȭy�p���'��:lˊ&�(	�1k@
�,R�'�YeZ�Q>�A�ں�H!��'�Be����LA$�À��qO��h�'sL��CC�+)v�0�>
yR�'R����L�;H��w�3/����'�֝!��۲U�4���oOK��*�'쌡��a$k9�D�1���K��	�'g�u�e�1o�=
6���mR\$v�C����*�� �"�E�@�6�~*4o�$W��ݛ-ʺ�b6�E3u�T=��Cɯ�B�ɻmJ:������h[�Aa��	�wi�ۯx��ic�X�r��E�G�p�
��b�"l���D>_T�6`�%g��b4g BKax"�ʔaˬ88b`�y�`YD.�a�|Q���A*
hʜ�EH1}<�A�5Y����܉>��{B˾;6MJIH45�ҝ˕i����(꺄x'�N xA��lߖ	��B�392,�������rR@<�"咱��;��  �"O�!�!�1+�yr+�:NiQ� �*f�BZ�n��c?�mࣰi�$XG(Sj��g=A/���wl�B"�/Sv\A	U� 5�TA
�'�l�@E��58L�����-���6H�(�?�A@�('ΘӴ��-ԭ����\���u�d�+d�y:s�S&%�p!`���Maxr�é[U��S�3?���k��*v�����oK5l6$�!DI�X�$�y"�ܭyu�u��nSZ��{���5�f$1�GPT����4��(��䟀@h*�eQ-5��pA��®`��)H"I�2��A.�"mԍR�%@����I�����*�"O �1JL�����Ɋp���x��|cD�i��A�{�(A���3&!�5B�|�&�P�޹λj.�b����*���c�5+�����x��R�^{�X{����+lCD���ڿ��GT
�݃GK]9x(��S�ӎ9��d�$��<<Ĥ��x�:�D]����K\
=p� "��T� -�n��F��:oTɻv)���O����N)4꬀�J��W���ԫ��^�KQĝF��Tp�&�
k��h�Q��P�@�k�@�O2������Z����~ʟ�y�f!'@���jM�L��r&���;�"�>kX�� �@NO�e�� ��%����FNd$�ӭi�bZF��M:N��GB�W�^ݘ�'ց%�X�ڠ딿8���s�D�R�עE��=K����<z��dI$JU�,Y2#ƃT�.� �Q��c�|ҖO?}����u�uI�
8V���`G �y2�KD���
OfpF}� ��Xb`��I>'�2F�\�B$���M��!��\TQ2b���R�J��>ͧ!�-���i�|`#4��(ZPi��6y�0Q#�V�'��i��M�6=�`��b�k�@pg��S7
�(���Z�\��"<i����lá�O�)̧ �esn�>@���3���<6`�	p��J����9��U�`۵"�����0�%��8��O6����G�4�����d�� q�'�I1�J��$	�[��b�D�����g>}r'����G�V�
	�U:#�¡i��+1���b�}Z�O���B(��y���) ����R��O4 �6c�+�ܼ FCO��O���j��?V !{�J��zY�i顉��
��Su���'V�:T[��i�N����@��>�[#-Κu���p��H�'��)�ÞuR�[�񧿫THW�t^��筙^����e�'p
�ϓF����s�Ox`�I�!��Бd��w��鷧�|�p���n� ��$y��r���"� 3��|}���=y��%�T��H�(�NY
$j�YIz�IH����'����2O�*ap E�2',I���vh_ g:����_�Xd� V:/�批N���&�p��/-�l��׼\o���RCYZfe�+�p̉q�H9k�0e��m&O�-@�h��(�ޜ�E��S!*���"$�ى��ݩT�	F�O� 5��fp��:sBϪgޱ�P�R����fb��s��~�;}R(�q	�ML��jǚh+P0L<!/ĮuQ�D[+>�g?Y���i�|�jφ�\<��#H7;�l Yp�YH�:�ꑄ]����cآ+LB��cK�
U�F|cq�	(8XQP������5?���I<Q����/�n9�JJ��'[�5�͂9#���%�����J����C�+t�@T��m�>�X2�h4�	>GSv�#�i��3hjhF��X�l�B�:���6 �,1�!�'�����#�����D�yشS���p���3!�}І��o�P,���<�$.�	YWʤ���G�
L�z�R>
b"B�I�D����ɝ�$,�d#�G^�m��I "H ��?��'��$�K��5U��;�*��I���\'ga}��ۙ��ᣢBO�pW�h{%H�/J�T��b�y�������:a�u��B�0yޔy���5}���P^��"�vqx�j�K��hO�%@c$�7E㰄��M< Z�Ђ�O8�(	/b�e�+i�t�8����p�1�)֐I�ƽ��A�hX��y��*9b@d�2�J4*��M/?ɰm��N�hUr���uO��C!Oh�T>�Y�f�K9l5j�Nɣl��Cc,D���eY"���#��,L��|�p�V�hٖ�#v��+x�x�䧘Oش���Nͼ��	]Ė,r��Yn�����[J�<&�(%V���+�"0��NN!�P�-O����@�y�1�1O&E� `L%|�F���A�r�
��mR�M��U�CdD+���"#�_?M���,h���sL�1<�^|"�)[b\Hˆ�~G$��	S"�j���"2�\����H5E*a�5-��V��, ��9�U�T�"�&����,Ox�	���	UW\�x'Q�#�kS�'	�\e�H�J<��W#Z�RZ��p`��=��a`�G����'��A 47O�t)��;J����&����W�'픰��G�e��z��,Ą������p��(c���PK<���$F�m���~��s�%$@�L��E��<%���G�A @h�4|�D8��J�?>���E{��2LHl	���L
��� A�i��!"G�մ��� �
x�e��'�Hm���+�����O������0�1h1�׫c;�h��+��&�,�/�OJ�C�A�xn��W�3>��s �T����:l�d��C8�ɭ|
��qp睫R�`�7O�
𼋵f��:���M�u�4 P�D�Dҩ[�Bڧ:��a{���:|
�y� +��a��H�Po�,϶0Y�G�/�d�7�Q̱;�(�"_AL�Y‏8?@�"<��2|'��#�@�A���0���<��*��&oT4�L�g�;V�|X�L�O�=Hs�'x�ћ�읪܀�a�dJ�HN��2(2�l�iA�H�D˦����)2 ����̎�I�4O��6 Hsl�kE�O'!�u!� X���)d;�aے'�;_�R@Zj���@��'�"#�<�P:��˺
K�����yr��g3���0����~bLI~�����`�0� D�Q%�|��s',?�O���2��9eqP:�d�	j6�Q6A1�^���T'�&����O������^���DQT&���ˆ8�����j܎Q�<eK�(Z>{s�D�cg�/u ��	��ĚY+xȒ`a���O�-B�-	y�Dri�:a��8��E�O�m��� :.YIʷ,�|�#�V�V��%�$��J�@��3�e�+�� ��JY+2�4	���<�R��X��%��ZQ?�4GV%� ��Ӏx�Ĉ�9elAq`hELBX�;4�'X�W�t�'dA��,T�:�F$�vɏ
�<��I��y2jU0)��x���ہ�~�_}�'��@p �M=�4�K�)B�Z����$G�y�! &\J��"�&À D<�C�#v�������Y�pE�y��Y�p����'�(q Dξ?a��G��N�T�áU*\��=b�Aѳ1���R8@��P H�P��;D���cr ڱ%E��!RZƊ����Ǿpx����A:�"���ٙ�h�i�/_L�����<�vL�xJPQ@�F��e�@D�4#�-GT삣%$�tHZ�T���ي�9�
���_�d�'�X�^����x�H�������: �
�?� ��3~BX�a�V�Z�v�a�B_��X8�/��X6l��!e��]�*�ϧ�?�O3|tcKP��a�׆�p|��X�N��*d��a��>��y�F��j��ҝw%�9��%6s�CBگNN�S���\�Ra1�'������d;-��q%4w�A��dƘ� ܪv-ш=bt%���O@��0���<A�Q�J�Q���H 
�|�B�.C(�(�v`�2��5X�� ���p ʛ.�6(�$N�EɈF��P���` �B5��Qc']/�H{A��y��(P��<u��T� ��W.�}��'ʔ��0�ԃ�#��8E(Z1�LY�M#H<z�I�8uz���NJџ c�&�o��XFN̙F�д�Vi�0��f[�%dĝk�I�(K��]z?�O+$s��T�dvn��΄;i����s��;gl�Ke�!jn�xB�ߩ��&e�咀EL�Q.��G��_����(^I�����O��P��� qbi���W�,p����/�i��X��k�Qq��P��;ѱO4U�%�^��
}`��B��Fă�J3��J�5����m��)�B�ծ�4m���Z'���OR6�ؖ&��*Hъ�<Q4䆣3����U�n�9�� �2�n98��	@ZD�2ȏ^��,E��O �Ka'S�%���j�	ְP�À
R�T�2dY��[�6`	�G�L( �?��d��`H���9���s���#/͖	����j̰0����G��<���~��$�p���MzI�T/K$	T��{��]%9i>��C�l4q��爠2�k �(VK@��b�4Iq����B���n�H�G�/p��'ڌ�"�?�� ��9'���Ks�!+^@��t*�AȱO<�@d�?o��xg'ܫ�yu�#�T޶%���5,�`���A��e�lY&��4���D��	�*Cr,��Ot�I'�$�B��-���f$�dgr%rIX�k�z� Ti�:.�r=Br&'�U?���йV�ՙp���ӣ�$����+^����1<<�FR;`k���dI�F��9rV"��oy��Iǀ�9��uh���#�rI�O�0����Ӻ�I	��H�� 1���A(T�D��2ʝ@�UX��U�b���$@�.���3Q�I)@�x���/,y�����6}���I����#��d��'̴��\"E��秘O0������e�k���4<�ڕ�jCV�6%|����%F�� ���Ȕ2R�EhK?ٛ�j�H-���d��3�p9�㗝)/��'��"v��|����V�t{J>au���:�0���WA	 1Xq�,w:��B9�l�S �U����|��O�T��&x!C���lb�x e�?%T��e�4؎�"��' �&�����sU���h5A�#Fxv��g��b�e��� �O�T� n��	��DpMJ�qt��D�
(��-�B�4��f
)��%�:Y�L�*!1�ё�S�6C�������I>��4H�
�?��>���&,�E����#�"�^`I�k��4:~c��X�!��@H@3lZ�0�Iy�-�N��{���1�� )f�EB�(�M���D<�s�@���	���'ڞ��կ� *�dApH�>f���噎}:��C@��eK����ԟd��D�%8����Ї9v��A�
��ɧ~��ʵk�l8������O�TI�p��|q��M�_��� D��H�����<����]}"��=� Y��ɄSw$�3�w��̇�ɉ{���������%kL�;oNV�Tx��
��~Bϑ8�r�'�.�S�s�((����U����S�ǎI�Tj�F9D��+���<Gi�Ea"ǐ�hC�@9'�$D��2����#s�! ����֭"D��J�a _Vn8
'���;�Z�3�H!D�D��́� [�hB�G�&�PTzfI)D����� �|��aÓO�$y���3�H3D�D���W=}��ء�*�m���{�!6D�8H�*�dT�I�B�� d���5D�$���f �i�1�6>"U��B3D��zb-���G$ֽk5D����=D�\1DB�7A��0���֨k��S��8D���p!M %f0%�U!p�$+�+6D�� eD�i���sl"^,
yP�.D��29HB8X�h��
���q��*D�\a�Ȟ�~�"�����L��f�>D��Ö,��h|��b��R������;D�0Ic�Ǖ�@JD�Ҹ\�<����'D�T�2>�Z��+�d�"�ԋ'D�0��@��>�X�!�3 T%P�%D�h�ĕ� �� �eM�[oм�G�=D�`��0h�4��A
2粄J�A;D�� FU&�QZ�\��eɋtW��"�"O�Y���X�y�*ɒ�FҰ�q�T"O|���![�=����6E>~� ""OlD9"E�|8�+�#�p��Փ�"OΡ� ڙH��%�爖3
���#"O���n�*U�ąsM��y���"O�L�uK��.��-�j�d��R�"O�$�n��	�H�l�4�"O��K5n�T����kP���<�"O<�iU*$&��!���F�y.d��c"Ob|S5�������ؠ/#Rl�t"O*!TE�)+}bl� �x��c"O�`��F]�f��c�O�Mt�t��"O�H8qaB�xG �a�?!tl��5"O�tg�	Cl��Q���2Uz�"OZa��!�L��@�ћW�r��d"O$�bs� �����vyZ$�"O4��B�I

��:�EC5�u0d"O���5͜�k.p{�B�[���"OFIٶ�]�V&J�2Q�ֻ�(@h "O�-�@�0��բ�8��#C"O�9�(Dp�
�ip��4YmʀY�"O��h7�u��Ta��ݐ;g�qV"O
��'˪P�$8���Ī&`�� "OX���c�\�~U�	ԥk�ȡ�"O�Xhh���P��ʵ
�t���"O2	��d@�,��BP�I�;� *�"O�Р��̆ � ��c�3/((�T"O�h ��;7~���K�8:�0V"O(,���)#n<����u�'"O�1��A#N����KJ���4"O8�e熞�܉��n�<E���s"O&,"���]N@C���ВE��"O�X$M�?H$���:�3%"O�@��.�Tj��_�J��q��"O�\��A�A�Z�'h��p�d"O0j�	�#+��f(v���K�"O~���mD�\���SA'p�h��V"O�8��-��4�����F�	� с"Op�p� �\ �h``U{n"`�U"OB��ɦs�.TC�ɂ�V����"O���I:rqV�Z`�T�87��ҕ"O.�ɑ��~Ѫq�I,$��%"O�H��H:�| �kP�v^p�"O���Zd�و��t!���E"Ol�s���9
9~h���+i�T�S"O����˖����q�D�U�b�q"O��[pG�7��}���[����"O�E��׶..0�$�D�X���"O����A@Z����4 X�ӊ T�@ ��G�����F��	:f��psB(D�Ȃb�_�U(����`,�*��2D��a�BÄ)�V�b/��ee^]��%D���� U?x����ԍm� �*O�����.]���QR(#�^l��"O�xy4N�B~��!0���x'"O}�ra�e4���`��xV�,�Q"ObIZ��s��t�X�j���@q"OJ�1��F�����ԥiyN��Q"O��Zc�lC���hH�DL�D"O�p꓈�50y�Vǔ�:��s�"O6��3�&TJv��� �"O�q�d��;M�0ՙ�$B+7&|�(�"O�Z�`�?P�B�b �?��� "O� v=������>���� ���{�"O6ȸ� L*�f�Jw-'��@�"O歐�iP;2�h'�:^R��"O4,�!N�mQv�ad�<�X�"O.x�� ,�6�D#��@"O������b����[�.�:�h�"O Pa�Щv<�h�A�;���"O��4�6�`a�����e2b"O��� #�%NuxXYe㐨��la�"O䩢b�]b-\��wO݂D$�Q��"O�p`��J���H��I6L�3�	y��$x�2�y6���W�Y�f9$���0���{�D ��T{�ڶJM�y�E�6����(�
Gֆ�MC-�y�";���I܏M��L�%��6�y�$�=|v%�1BʟKT�`%�G"��',ўb>mcB��j��8BUm(W���� D� � G*��0�K��4���F D�tˣk֭"�����o�gȔ<pwL?D�H��
j���z��|fpRР!D� Q�IB���0����y{8 ��=D��(�b���I@$�Qur�#&<�Ir���'zA"�ᗄ�
�\�3���f��\��y��0g��Q�`��F��i\ ��y	*h;qG�<d�e�Pț�@�ȓaƆ��Eϋ�^aV�*P�"l�|��s��M�gg6NeP�����Nu�i��~�whN%L7*A���DsE��������Q�)M�I�t'�<����H���R���`�A��A�������b}���,hjn����Q<h|%��o��y"�ģ������
�x�B�@���'���ډ�����s̍�#xr�(��O�oE�iv"Op})V &�cr* 6���z�b8�S��y"��_���C��Y��#I�&�yr	��0�\M�%�Ʋ���IB���yb�[h����JJ7#\ɒȏ��?1�'4�ږGC�Y�ސ� o5N�>x�'�Z�Js@�;�b��WkT 7�Z	��'��%2$�\. �廣iJ-EGN\�	�'M�Ab�Eڸ�P0��ʦG�T�q
�'2M2҉�&$Bp���6:C�4��'�(���OG
� QʤE�4��,��'p��&�(Mj~Bs�-,:�T1�'��5��WDm�x�'�S?+���"�'ԑrDJ/ ����V�Ȏxc�;�'٬���-!�v�*���0C���
�'��-�Vn)/��h�E/.}N���'��1Rh[%P�^\�`� =4P����yb�D�K�|�	D���w�8�S�b[���'��{rFڐ�d�,��i�ZQ�@
,�y�H*�D�AJIgY�]���� �y�F�"+�]�fc��Q��ŀ��g�<�͊��0:�X=D��̈b�N�<��&U�L���dƼ�U��h�p�<i�i�&"�����V�{^&�ZG�p�<)f�5m �*���}���[�%h�<�p��p����7Cn��@n@Z�<�a�M���,�} ���4MZn�<Q$�ĜNc@���� `��A�f�<a�V�{�+b�N�fX��A��a�<��/]�N@|Zү12N(�Dn�^�<���F�'L)��Ӱ|[�����@W�<�RX������Y0B��M�dh�i�<� ~�e
�(�:a��Y�}D����"O|�5k�� �\��H��U�}S�"O(h���.�4��F��6պu�"OT0ÔZ�	�@�+�l�l� �"O�x����;n]T�8W��8h���'"O�Qr�@�]&x�P�;� �`"O��:��[����[�I��k��`�"O���E�4��Ti���S��E�"O�x���#_ےu#5oQ�4���"Ox9Ʌ�Mb�����JM$��2�����ɫc�:�����iŤ��3�ED����-��ñ��Q#_��b8�W+B�<L!�$K�j� k�^�(?��PCː
w!�dI^JraQP!�"U& \[ظ~]B�ɻ>,$� �
;��� �'g��C䉛)��is��	 ��Ur$�M.@�C䉴;)�]�A�0)H֩��aF3+!�C�ɓ M��)>^X3�k��9��C�:>h��Ơ�9! 4�"�o�bo�C�	�:�m	X� ��r���`ש#D�Dq�i��ʌ�tO�[l�"�e7D��SS�Kf�ɻ��
+Zb��Ӄi!D�w�:B���S�1Vn��a=D�T��^;a1�e�r'Q2}q�҈&D�`��k�>X�40�a ЄRR:���%D�|�բĔ��i2P���E������/⓷蟊08�JP?EЅ�s�RqF"O����?F�̑Q�I��.�ɶ"O����o��dH����-Z�"O\���ו: Z���@�hձ�"O�h�F�O�c/&d(��t{[���'H�k@
45�D���!�-�H�[
�'V�=S!�>3)�aRuc#T�I��'�.�Y6�$|��X�sJ���i�'Q����*O�.I�����Gh8�'�\�pd/�:8�2��# :�{�';����x�,8YU��Hy0��O�eҲ� V �Yu�L�Q.��"�:\O���SkW�>��K�	վH!B(1"OJ�ZVD[ .�"e�c#ƥ"4|I6"OD�k�nA�.L��hEn�F*OF¢n�,*����M�|�pp0L>����߹a4�R���Dv�@�f�Tf!�D�	��H�ªN"yp�؃I@�"g!�D��-Dx"f�/+�ndـ�<\!��$���]�{�hp���vG!�DC4�A���	{�*��'>6�!��!j�=c�\�f�>]yCa"~�!���H=�ɘ6���"��i�%R�A�!�� RF(�r��<JP�8���h�!���>G�.�i�M^��S���^.!�D��p��Y�����V$�#J�6
!�L�_�0m����y�����&^�!�$�+�`)�A�6m�A��
	�!��L;$�d���I�W��j7� !�D/��m�G��E���<!�$�#4b��H� n�L�N�/.!�D�(v��1*�%$X�a١�R%+p!�D;r��� ��A�c��	��Q�fY!�dP� ^�8��L"R�� ��� pT!�):�m#�F%nǾD���ɑBT!�$%ր�%�Ѕ.6DI�o��V�!�D, �L A!ď8��A�7^�!򤉶_7^�J�ɣ$�Db��7!�� T��C��<I�L�Fo]S0hܐw"O>@;��Q��έ��˴,�-q1"O@hs���|�����%�=@洼q3"O�X ��� ��#����\�)�"O�[��[�"V���
��e��"ON�HU�Y)��THЅ���V��"O�@���6&��:�D����"O�� Đ ���kC�;5<��e"O�ěe��L��A�k�5>� "O�Ƀ��V6(Y�p2� �~0Z�"O�CH��ڹ[���5��A�"O��a��0yy��2��%�d\�"O�5@TlV�MJ	�4�
����"Ol0Y�`˥|{zL���4e��;2"O6�UA@$p���V.Y1O���"OF��2ɘ7,nPl�<3���"Oҙ��J߻цS��J�'}��"O�2�s��1'I�c9��"Op�A�QA+��%ܞ!L>��"Op������I������`�V�y�"O�� �!"M^��R'UɊ�P�"O�	+�U
*�I����![%���G"O
����"VD��Z1Nȿ|�T��"O���p�C& Ѣ!z�m_bl��"O z6-��> ��B�R
)8@��"O8hQU�޹f���;Ao!Q ��0'"O��gk�$w9�-+B�D�欥�G"O,IX��<�h����N�r0"O��#G"ԧ��Űb�T;޸��"O؍��cFj$�ъ��I�ꀓ�"O\A����3S�f����ơ)����"Ox,�UiX � ��֮-%l��"Or���O.���*U¶Em�"O�9H�F�h9F�c P�H�FxY�"O$M� ��	��ur�@���c�"O�0��'źP*�8���8E�,2"O�$�4�̒A�jD[�@������r"O�ر��}n��2E ԍA����"O�}�ޒWe���& V>0��S�"O����K�faT	�j~,���"O`�ĥY�X� ����-OO��"O�h��+R��ft���t�B��"O�u���{��@�7���~���A�"O�l0�ˎ5�Qa@�1jg���b"O� �� �!Զ�S0��)X^=Õ"OvyꉐG.����A.T`�E"O%�q!,K]>���C@�w�.�W"O<P��$�m���Ӣ�U�x�d"O������hb���z�X��"O
!3�'Bh� H�(��a�"O�`�ѕhv�Q ��Z�d��X�"O�X!���`���(�D�#[w��R�"O"�@�.��ݶ��ʺys0�:�"O2Y��#ح�bPyg�D���d��"O��	"��dy0���	~�C"O��Q�q����d�E??p���P"O��#��%gP�<�!"ڸV��!�"O<`#&M�Y*Z�X�+���ԑї"Oج�7�3���ь˖k\�!�"O�!��п[沈)��H8v��"O�d�T��JԸ-h-kaB�[ P;!���ge��Xu��9�8P#ÖE!�D��qpv���\=O�����"�P�!�]��:ġR,o�ĠT�#�!�� �@�`ڬ|'�$Ё��I�n���"O����ޘM!
��0L�>z�Fؙ!"O��g�� '�T�DB�
�
h��"O@���I�O;T��i!Kk��""O�����B�cȄ��Ađ���"O��� ���|���@�.4���"O:�zE̜#�*l�S�F|���"O��	tiO:%�p�cn:�d(�"Ob�����D��U�$AF�b"O��rӌ�b�h���,^mZ�\��"O�`r�63��U��63> ��2"OT��r}3jq�j\�i���c"O�ixtNG���J�Iɣ'��I�f"O�=�F�9_�(1Ί1rz�+�"O�Ѩw�ǩ2Ϣ��NA
0��@g"O�5�3�w�����G����"Oȝː`�|�hĊs��ܘt8"O&uA�%f��x�NJ/RqĬ��"O�\�sMÃ�dB%΋�m���"O��׬�0%A�l�jpF���"O�sr��lc~X�P� EdN�"O=;I�)/,�����,# �Y*"O�(j��O�l�+���	�'��P ֠B�a��!�gD�k�����'��m����B'�����	jX���'*�$X��V�h{ (�7�8\��	�'BZh�Ǆ�!|�"I����[����'�ʹ��` �!:�`v��M�����'Dh$iԎ�^�^�U� �[ ��`�'�f�
�l̑>��U�T!%d]�X��'�v9�(ͯe��0\��!AF��y2BP�"yY��PBV�L�S%�1�y�[�,�*�g�7P�p�9DD�1�y�E���&�t)�Ӟ��Cd��y�PE5��������� ���y
��Ԙ��i����pUL�y��T�x<�����wRz|ՁӅ�y��	e��肓�]�޶�H��_��yBbT�k�,PK����E"�t#�"*�yҩ�d��l�26~��A���y��K&e����k�>4�V�
�E��y�-�
���B�ɀ�)���a��y�Nڣ��E[�S�q����yr�K��	#�E^�����׋��yR֞$��Ó�"h� K.�ybkR;E$ʉ��	�9SZ4`#`ś��y�l�$,U��1�mȍG�3rO���y��Y�	�4*���;
*������y���$Tl�`�D�06��z�B�6�y�Z�r��c�)6qn��4�K��y���/6b�#���Y���sM�y2���jd|��ςIqf9��)?�yR�WW�	�veQ�*��3!�6�y�i�&c�)a$pEXgʕ;�yR�S�	ɫ2B��7I���,�y�E�"�@�JF�4�uk��y���kR!�*̾ 
,�KӉ݉�yr%%T{z-�r� t9�(do�(�y"���
S25���'؂u������*�3b���j&��thH4�8P��3xYbn[0kv:Ѣ�ojh�T��3�hř�L�t| �AAA�B�d��ȓ�tQ��$)�pk�T5:ҝ�ȓ,�XyS��B�8��5)1���S�? �H[�#��,�m�C�T�(��
$"O��)�N�n��X��âH�|��a"O|UY�#�)=5�̒a-ǡrK��� "O��ZwÆ#OJ9[�␇W�db"OР�׎ِ6�0��s��&U
�"O8��C)ۤ��E�a�턘��"O\���NK\�Nak���ky�,��"O*Bq�{�pȢ��5j�!��"Oꉲ֮�#-t`�XZU���P"O�l�0�N(P���K�D�A;̡�e"O�ahe֞�8��%J�p'����"Oaу�<>vL�Eb����"O`�kM�M�
�̍g$� �p"O�	i��ݙi#qҦDC�u0B�h�"Ofy
�N Hy��F.�ry����"O��@�˛\���a���#:P
�"O��3�^G��\@Q,C/+�r��"O&<��υ|�N8Y�k��T��`"O�d�gD��>z��4쀷A���aQ"O�s6�S�
��AZ�4*CNt��"OF�I�+�.S|D��wD$>�W"O����J�\0#Û�"S�)R�"O��b��Јy�lҪ7��L���2D������e���P1a��C��4X'�1D�A@0.�ɊP��b�r���:D��)�$ҞA��$���6f�+g7D�$���T�CĔP*P�K�_J,0	`4D���Ă��c��P�aD�P�$�8'�6D� ��1S6BT8�N�>D�2`n5D��� �B�W� ���$��hqh.D��{G*��1zc�Ҧ�$��T..D�� �)=T~�xC�N�O$�M0D�d8�$��{9~Bf�t�c�a-D�h��ʛ�w������G�Ҭ���5D�0�W�J�n�$���:��rW>D�D����#8L���# �`�C�D=D��L�-Y�� �Q@!G0*\�r�>D�Ћq�&o=>0��ˎ�)�^`pu	=D� �����LI�KN/h��0c��7D���G�q#~�����{��0W7D��q�Թ=ϼ��D�K%t[� 3�c5D�8�QZ�H�ᣡʛC
�t���'D�����7b����͚�	n��`�%D�Dj�'�VH �
ܝ,p�` �k(D��ڐ��B=�Ex���=Nr���h!T��S��,�v�*���}XN堡"O��r�`��N�Z6MHN�cc"O�hH�(��LQ�F�Q��"O��E	�?���
D�	
/6x$h�"Ot3�+�i2�qK�N�1 (���"O�xɒF����#m��F���G"O()��l"���W�\�U��"O\�W捰�s�*��講�"O$|��ab�<���1���%"O��;r+^~�D�bX1q�v83s"O Y�qo�H��p# ��"O���`*R+c,F$���K+=^a[�"O���f�"M����I,�i��"OP,���W�l)��� �]�xb�jF"O��ҥdʽKX��b�4o���b�"O�ꖅ˷"S�i�0��K���;f"OM*��*1D�#�!J�q*1B�"O�"E�=���c�*�/�iC"O�c� �9���P7bfuy"O� xm�R�ϽN�!��#��e>@u"O��sEьMܤԨR>I(��"O1����0"d'���"O�UqnW�x����6sF\3�"O�Ti'�%L��{C�7c��l1"O�a )D�_m.<pGÇfʹ�1�"OT5�
�	FA(2h�M!�AW"O�8�-Eb��uJ���g!�9�yR (O~(C�_z	�)?A ��Y�pp肎]�d�Ӈ�'�q�ȓHXL�3c �<T��k!��:M����ȓ(���J��t`��  /�Ф�ȓ,�=aƏ��J�q��=�bp�ȓhti0��L9�ڄh`�@NV0��j���8e��&i�������:)�I�ȓQs*$	�i��jn��,�
6nN���9��)��R�*L�q ���1��e��9����2'�H�L�y�`�k0��>��XH��{Vj+U��6�h�ȓ`�`$��_va#gL�<��ȓd��y@BC�XM��r�~���en4����[|�����id��g$<��#�'B�h0A٬ ���ȓZuD)ذCZ�غl�ƥ#Z��ȓ]�1[sDW�jC��)$C�si��ȓHW��n�0��5��-+xE���ȓb�2��Z�6I�󮑪0\⠆ȓ{��=�$ڞ`c���j�%^��0��^Z�jD �j�T�Ɯl���ȓ"�Aiɠpq:��R�%��q�ȓ�������`�T��� &��ȓP*i��/<&��w��$c+8D���FѺ
y��P��F٨���'D����g�%����ϓ�#v%�s)$D� �be �+R"��e�V0^E8�(D��BPC� 	��|�7��\Q� k9D�(;G@�f읻�'X�Gx@]C7�8D�P��7q����&.B>L�t��e*D�����@SHn�a_�N�~Isub#D�
�ǟ+g]l%P2�GL���D"D��e��;*�L|��+�}6K#H D�� ��T6-u�htQ��3�2B�	%3�a�a2[$�X&���j�hB�	���rV���Z���`tKA�2zDB�I�j��E��q܌+���s B�	��x�j�N�C��hU�U%C��C�/HV�P0j�6c�PÂ�7w�C�	-6��!f�WrR&�"�gM1i�C�	� ��i��MuZP��Ǌ�Rr!�䕯F��p�g�5)>`XÁ�K5F	!��*j`6��wΒ��´;6�Y>!��
�	Wʽ#��N;[�d���J�d�!�ی�#�M��D\�'�I�!��n~������q��p��!G�!�LRα�vG�/�ȍ�w�^�#x!�dT�j|23+±#�m��EE#a!�Ę�?��ت� ��Z�C2�� 4!�$'+����eJջy�n�`DR�!�#
$�=P�Cة ��@��+T�!�(TNp�نG��=�Iw �2v!�D�?e�-�E�^!$��%�ńʢn!�K2�4�0�פ/��$K�D�MW!�d�ZWLI����+\�c��&et!�L1�>��̮<��4���*a!�� ܠ[qi�M$x뉵6���"Or|��C�UU(9�R�Q(HPIU"Or�i�-H��ٵ�^�D�����"O���W��x�z�E!�(��p"O���b,�R������ݠ "O�u��O�%@��J��,b��}�"Oj��w��;l|ށA�mC&�x5"@"O��0}H�\��� pu��"O ۇ�1yz����Pm�H��%"O������mi�<;�!*�|�R�"O�``/ɇy���C&`��-v@9:�"O>x����,�%z�n��Hp蘀""O�ʖ��vh#��cP,�f"O��r��(T*�sg�M�b�qh�"O���gH�1n`az�C�2G�R| �"O.h`�@J�*�XAl� 4���'"OЈÒk �%�Z��e�P�xf��	%"O&�J�+B$Lk��	�hd>��!"O����F�#�j�P5*[=f�`C"Ol4�P+=<^��Qd�"}�^U��"O��z��,s�4��"\�z�8R�"Omk�7�TuA��4A��	Bq"O�ٙ��R�|������O[>1�"O��@�K �l )T@�6=2Ԕ+�"O��ƭ��S�<�Q'&D=Bb�"O(�0G6zE�X�� eJ!��"OB�tz�LDQk �Ax�� �"O��X"�J�%4�U��*�kaE �"O�|�p��s�Ω�I1Q�	�"O�1���Yh�H��j3��*w"O������U"@�X���h.�=z"O��Ȥ� 29��y�M���"O�{�@Z d�x��ƤA��"B"Ot� &��z��#�AB�#0~d�"O�P�ui[@��6��3��D��"O2 P!��Q�՘��?`�8�c"O��K6�Y_ր=+��+~��]�P"Ot����ҰC�W'�@T4�D"O<e*TD�X�t�%�#�eX�"O@���LM�j��ݠ!�4�"O��H�/���;� �>�B:�"O �����2-QP�O c@L�#�"O5�f䕑C��A1A�W$���p"Oh\��L�e�l�L�(��+$"OH1�6`����r,ċ-1^��C"O��#���(/����g,�r>�Be"O��	��K4*���ؔ+!e���#"OZp���%�nP�Q*�*j��B"O�9���p,�%�Z�p�2��"O�����gH���A��
@(�"O�9���H�V0g��
�`��"Ol���HA�Dd����U:#�́��"O��)��/+����[f��e� "O,m	H��6��x!�"^�{�����"O,DB�C�0B���RH�!'}�"OJ�a�J�u	:2$��?�%�"O�I���<��J�]�6��"O��'mM#BT� 2���8���p@"O4ɠ�6�*qq �҂G��T�4"O���$@ &7V��h�+%��"O�]���j�I2�'ӕ\$xy�"OtHx2��;l��s)&�,xG"O��R���↺t2�p5,��y��hB��Ȓq�LA�D ҄�y
� D(
��R�U��@���J>(���p"O||�	۬M��!
W>�)��"OZ������b%I���/ ���"O�\���	�8�&\:�Jǜ �ه"O� �V��(h64ԀE��FwP�"O��
#��\�⸻��#A2`zf"Oa�F��+�Y��J4X\
L�"O̽rІ��-~Ԉ��B�'U�]QC"O t����#	�TH`���T=�q�"Ol��#+X�vgnx�u�́5C���"O���"C-���Շ��|B�"Oeb�bԼc�#�ʓ%��Ke"OD$ v�R�Q��:�-ˍTTA0"Oz��&�r���cf�Z([V��@"Oe,��EJt�1��Z�lX�Hc"O����L�Q?聴f��t?|<�d"O��	�*+�=��F�{<l\B�"OT��	���P0z%��D��1"O�|�v�D�b��	���9;�Qۅ"OjeѲ��p���k�#V�L'	Ya"O
\��%T�%���P�L�'LL�"O�9A"Ì�1N�C�t�d��"O��Em½;������I��R�"O�p��L�3'�)7 ���"O���`�&��d�& Y;4B<Ҧ"O�ȓ�ψ-#�N�Ғ�Y�T �г"OT(�7��h�e)���c*>��b"O(�p"��1#�a�N�:#��@�"ONq�6���
D�4,�0Ph4Лu"O���R��:!8��pJ\-&R���"O�� +S��F $>� *1"O<�8�R
	� ��Ś�`F�Y�"O��Z�I޴Y@V��$.!�����"OZx�RFѠrt�N,7D�t"ON�uBшy@2��B�0IH���"OP52���1���� �~�hhy��I�<Yce�	_S�:B��t��� �G�<�ƈ�;Z8<p O@�Vj�a�m�<���K�M`�S�Jܟ#�6+��_b�<�+o*�Lم�B�YI�5h3��a�<�2gU+<=��`�c�l�S���D�<	'��RG��x�BP�).44�A�<YQ�U �BUPp�q6����Ji�<y��ܹ88�sIP2�cejLd�<A�I�9�"��g�X][���/�u�<��)�	_
]�4kH�	�l��`SI�<�&�&B<\!��LBvH*���J�<����3GD���f�-ЈA2���^�<�ǡ�<XZ�Y���O�B,r�ŔE�<���%�L,~��#��K; B�ɡ	ZR Y�+(��iEm�740C�I#u��0�e�,;�����j�RC�I�j��T'L=qP���CD�#T�C�ɿ9���+RG�� UH��F#"s�TB�ɚU��m`��G��0|"b�!�hC䉽S����w��?FJI��T�
B�I.�h� �n��+f�YuEߵ^x�C�I�D�50R��r	�`a��$�`C�ɟ`��)3�H*"s�-ha�\�ZpC䉇ac�ۄF�n�he�H�JC��zT6�Ȓ��EL� �W3�8C��?�0���7!�ʗ6	�B�	"NP��$f�� pR	5ttB�	�k��9����[* �� ܦ�4B�)� ����ʖ1���C ����hV"Oh�@�NۆF�ɐ�$��%�* 0!"OP��䇚�c"�2��ShЌm��"O⠐��-0�}#�(/���Q"Ol��eM1��2&��3F�*���"OЩ�QG:4�l% 1�?d�F�	U"Or�U�^�ҝ��LU�Y��D�g"OP�QT=P8� ���1�ֵ��"O��MŧD��4C�jM�K�x��"O��g�^TF2MzSCK�}�x|kU"O6�UL��d�0�	�k�X�B�"O8U�p�	8�:��NV\�["O�Y���fw�[-A:kh"��B"O�\qGP#9]]{��'gD��v"O�}��D0A�,6��;Y<F1�"O,�a����X�!�F �~Y��"O�}� �X�ب�Sd�0%���`"O��	��<?Kv�Ȯq~���E"O���F�	�W$Q�҂��0D� �"O�H�6.��cιz�B\e��HF"Oh}���Ex�S*
lbR�h6"Ox=cĀL�Q����V\p����"Oީ#���oꮜ���Zp�]�'"Om�R�/T���g�#=���8�"Oxh��Ps4��/�^q @"R"O�(476��$c5��,s��`�"Ot��)o@t��-��|xeZ7"O�MaRL�~���٩(\���r"OZ��0�ՠ*���Рb�>���8�"ORx���eJ)ো!@fB{D"O(q ��@�Cܼp@���#+�)S"O�:g�I�0�@�����,�8�"O0�{C�	���HFCϗ�<�PF"O���"@4{�t=Q�O0jϰ +�"O4͑@�ikTZ�$Q�=�t��"O~x�W��u6��:�\Q�ޑ+�"O�c1L�_o��qEB	:4�"O���4���8u��	g�j}	"Opٲ��W?K�r���ו@����F"O����b�6B�N4�iĄey4�Aw"OЕ��X5q����W��k��k�"Or��AG��_�����> ���"O�@2��ڪ;,���ϊN��ib""O������v�Zl#�M�Cά`c�O��@���C���!�Z:`5x��O��=E��h^�^��RW
�?6��Щ 嘠r!�D��^�D���B��;��l:Vĝ.&�!�$�I)�p0q#�d���%��`�!�	��<3�'I�q���	�3:CrC�IpL��!G�	"\gz4B�'ϦbrPC�	.|�af�vǞ`K��
�P[VB�I�O�� ��9vo�`�dȚc@B䉺L�9H�G�8X�α�*H�@��C�I�jRm��L2Ҿ-ZT���} �B�I�	l8�GiN+, ��) eO�ۤB䉄3�*�0Ō�vl�AsB�L��FB�	�o8�x��}q�-Z�˖EB�I;#%�h wgP�y�\3���:1�B�ɤN���el̥U����GI�`�jB䉻D>��ir�E�2��i� ��d�zB�	�D�r��Q�mB�(B� C��&���(@�M�F!�i�,y�B�	6p���M�	�Ţp�ǒA��C�ɷ,TІ�Y�R%Hh�QjC�>-~C�)� 8$��-A8��})$�<W��h1"O�a�� \O<ģ��IoQ yK�"O���פ�F���bK�%��˶"O��1�[2k�P����s^�(��"O�U�Z$^��J�&y�IQ"O�A��d�2��Q%1l4dI�"OHᩳ�_�\�� ��3n0�	��"O0%`�*��B���+$b�O��zS�D���L���n�z0�OC�ɦKцDLC2S�, ��3�C�	�$x$Bf�,�t����s0�C�Ix�̸�J+&�m�u`ݟevHB�
���ڧ��^+�0C�nΟQ��C����mc�O*h�����?R8�C�(P_x��IB�6��H;�bݳ3PC䉝47"9j���S�Z(����"fC�I�)'ڑ[�d�#h�:�c��[(q�"B�q��`�/Kb<dL:` �B�	>vXv�P�	AX<��d&�2,~B䉊u�|,bS� 6W/��i%Kg�C�;[a�92�piة;%�@0.�C��<e�$����-j?���Ff]�B䉜QQ���	c��M��I`ŮB�	]#D����ހ�8��D/�B�ɒ�T�nĢa�*d�p#�=s�C�əF��,��!�⬅���L���B�	�C	R�A5������F#��C�ɼ/�6�st�O/t*�e�G.�-O��C��,�@zeň�8qn��v)���C�	"M؊a�@a֌?�2%2#N�:g�C�I.���7ɖ�\�u�䑥V��C�-kyI�NȦz)�`��	�*iG�B�?�69H�
�[�@�Ѓ�F��B�	��H�a���
���v�H�0רB�	{���§g��w��)�AELg�C�I��8e���6�q��&P�Ou�C�ɇw��Wd*d���ǁ��:���"Onq[�(����k1&I`|��JE"OV�7�/s� tb%Ċl^�Q�"O�癎hh���Tg�*Uء(�"O����,��Gz�Ձ����2`��`"O�xA�/׉]r���LY���6"O�0�Aq �)q�a��{G�Y*"O�ݠ'/�>:�T���H�~6*��'w�	ß�F{J?�i����n� ��j�,��cg�!D�T�� f�:6��8Z;���3>D��e�4fL����uz�z�;D�l�0�Ӹ@���W���Cp�f ,D�4��EA����-e�J	JAl*D�p��"�7x�#�IL0%� j*D���B�-�<�ءa˝`�%ID�(D����,�(s����
�V
�Őv�'D�,��]#p#�48����7���i D����+*�A� E3i�@0Щ!D���d	+�`x�+j�Fp�£2D�8hB�:�Z�{ !G[/��K��6D��ju��q�(!�D c���Y�6D�x�`F� n��8��A�T�f��M2D������B8����A�4�H�E 5D��x����~�CF)C0L�f��e�5D�\ꓮ[�[u�0��+-�e�ҧ0D�����T�UF�A���&7H����k0D�hp���uOȵy��G�#��a1D�L�:D8��`9i$.�e!;D�� �@;��X~�ђa!x���"OΌ��/\ _��`�Gv1X�"O�����(k�L���/T=��"ODȻ��\�y J�Q�A��0AB�"O���
�M��D"
3,{�4rS"O�ĉ#�M����*Ƌ��
��X�<��%A~&�i�r�� T���)y�<�`�@�z#R\y#e�'.x�!��E\x�<V$(X j�:$��[ʀ�BN�������FJ🜖�(OFX:(�I�΁iA/Y���u��"O�9鱢�6:g�����Gq���"OJ-U�T4B���#Nu�!b"O�e�̗��`ș�'WҠ2"O��H�NY?�8Ě�CJ�b�� �u"O�� F�e��Z2���w@�8!�"O��XBV�&���S-�9Ƥ�u"O
E�6�z�B6Cƍa�R��T"Oj�v���~nZ�Aw���H�t"O�i��X��ۓ��#R�l��"OZĂwč�1_�E M�uO4m*�"O ��r8��%/>�d�U"O~�@tǖ�OKJsUY�@m�)��"O�M���( ކ��lB6$V.5z�"O6Y�6ֺxn���@�ڎ��!h�"OB5���" �hm:�*��#�bh2#"OZ}��	�Bt�cu�(M �[�"OL9��

7rD�8%j]�7H�8�"O��fF�1�HQX�J��I@Հ�"O4�E�(�N�0��T>f1$H��"O������ZNe+ �±6&�غ�"O|�Y���.g�شz�K��Xi�"O"��"eT������%0u'�2	�'G$P���6V����쟒;P)J�'e|p�e���pBd��tS�'�jYr�O<>�< �s'�'H� B�'X�"�J�(r��K�%ح=�j��'�����ڋH�ru��m��4�e�	�'�`}��6 �����:H��t�ȓY`^���O׿���q��M�[ ��ȓJ�ڈ�0E8L_P����Gh<�ȓH]�U��<I��-h"��*掅��O�Ԅ$�5��q���X
����xh(����!R�m�0>�ćȓOq�`�Έ�S$(局)S�^vPل�e��m��/+q6Ĺ��޶>�2!�ȓ!���q�l�6c�2�괣Up�L��m,8誄�:"n��R��0���ȓ� �;����0͂���(Q�a�ȓ"�*=�eHVx|���S�$$�@��ȓ���Ñi�'��P��X���`��-h0��ʗ�� ����ȓ�Ȫp�W��$�'a�F�z����걡��̀��E`G��#�y�� x�����D6'��@�_=�y2�CTpQ�Є>56�yG*��yr��F�x@)CÁ�zFD�2F�܍�y���im&9��A�:��4�"D*�y��0l4�T�(٤���x@ʱ�y��6�\4`p)����rl��y��S�%5~Q3"�آ�ؠ�fGG��y�OU�6jb
ط}�l��ڄ�y��=f
�i�H��}�v»�y"���852�*J,�- а	�-�yr'��*���ie��v�2!��ɉ�y
� ~�J�fF�rդ\*f�E� (m�p"O i#�j�9i:��s�Ԁ	l�k�"OH���fJ�B`�Q8�fյo�a
�"O��9��ÂD���i�T��!�U"O(e�g��;�.5��cһD���k�"OE�2I@A���α@����"OXQ*#��޺��B��<yq"O�F(�Ll��D���
"O�Tۦ���De�|�&�Ȓ��$"O�l��GJ69�L�3k!?�Z@�b"O` rs_-6`������6��CG"OQy���_�NpPs�՜Y����"O<My�ↅ6:tH�6�ķi@�d�V"O��3��W�5���tOl��"O����ۜV��yR$�\��`�"O4�Y4��Yhb"b &���"O�x+ n�W���Wf }t�)*�"O��ړ,[�:v��pdօ=frp��"O$EO_�'��R�J`�t�`"OV%�e��T8��K4HPb1h�"O���%�8u����+Z �<���"O���o�����@J�m���E"O<���<Q���w���,��|��"O�\3�O
?/�)0��G�@|�t"O��%T���3F�R�wA�4"O�	�P"秃�0	�����17!���<rH�Z���m��	q5ρB�!��[,e����?U�b�#��g�!��uO�z����y���W�N�`�!���^Q61��I�y
)@1�R�6�!򄏓S����a�M� �q�9 �!�ִ]a"iJ�X">ʍ��F�v�!��S��Ҝ��h����K��!��{�|���J&m�
�d�8J�!�Œ_����' � J�ޤb0#D�Ar!�D�hX�H���  ��0f��MC!�@�X`&k�,� �{s�U*s?!�7[ ���M�R�$��a�;!�d@���0	Y�WL�(����%V!��ٳrt���U��"q����47!�I����7l�?1����5w!�D�y-����
��)h&�Zlh!�DL�]˴(�b/�2�ƅ��B�&"Oƴ� kC�JH�@z\$<�u"O��(�Q�d��`�� �`�"O��C6�B�ݐ��=�$]�@"O��@2"K�/5*���K����J�"O�%�fm�4{����k�d���r�"O:a�	��@b�[���c��2�"Oz�3��z������C��${u"OB�Ѓ�]�8�Z *M���C&"O��)u�ݷFd�YIR���=�!"Oh����))��+&h�)�0���"O�\ȇm��W���hdɿ��YJ�"O���I�?^&^,����R��3�"O H�V��;K��|�t��"O��X��F1e�pe3�'ݜ;�Xir&"OҌS���/!>%�0F5_�� ��"O>�2�=�r���BZ�K��)!�"O$ ��ϕw����0 ��?�<�I�"O�륅_�t8�,H�n]2t���E"O�If�~��!W��y�:\1�"O�y��bK�@�����A1q��|
�"O(�+�i2C�\��"A��$�
�32"O� ��� ��G�Τ��"J�Q!*�x�"O��[��!M!h<����c4��P"O�a���g�t�$�'%�P)�"O�-��C^�`���Ġw۞�8�"O���1��j����N�	��Y�"Or a���N�X�ʢ͍�_OҜ�R"O��� ��|�@���.FV|4��"O,�����z2�@�>a27��A!��Ў����d�/e�0�øm !�$N
}����!�� ���箞?2�!�P*y��(��ȏ�o��!u��J�!�$��e����K;j����J^�j!�D�!{�����.ʹbb}��hEA�!�ޞL�T��1"�W�lbN�T�!���9Z�4��՞X�`�`&�7|!���7������sm�����,Fa!�Du�dGS1[\���KR�$a!�dN%h�0;V��)3s���֠�?;D!�$�)i�޼�SM�|y.9�4���j&!�$��t��DƀM���@G��!�d۟.N�y�ň�.`��)� C�3!�䊉��T��ڸU8X@ѯA�V-!��"��Eڲ�[)b����
	y�!�� yByy�i��);R��6�._�!�ĉ�ac�	BF����Z��T�!�43�
qA��B� ���!���!�DV�;	$��o�6��|Q R�!�1�h���&]���yJ�L
�%�!�@�sjt�y�a��+�6����!��W�&�±�K�Z4 ��M'3�!�$ _xpx�j��i���y��߭'�!�E�PPa��W�Z�`5���8'�!��ö_�<P	��):~V�R-ڸ`�!�
w���PsE �zt����Lխo�!��ٜg��E�e��;]u���ťP�!�$�3`�9F�C�8��Axe c�!��ք"�04걤���x(�!�$�)q�ac �h�(�c�����!���"��	��	�)S ����[n�!�^*NTtZ�@ �>�����N�!�U����7�M1��PJ�8T�!�$S2���se��A���(T(W=I�!�DŇ5|x�qwM�.��t �f̽q!򄅲\��ڤPol��&�'qY!����Z!����pT|�p�d��+��� "V,�d.� x��dNO��y�)d_֝P���`�\刡`ҳ�y�O\n��
�_�<i�5�y����!�t��&/A !v��IE$�&�y2 	[��e���Ɠ�������yb��12-�b�N�q0!�HA�y"�Ä?�jyݴ2%�u��*!�d�:���� *ܰ����"�!�$�n"��<wѤ���f!TO!�d�)5Ka:�b�<}�0a"�U�E!���� ���U9IȁH�$Q�Q�!��h�aqpbR�pD�92��e�!��N��ؤJ̰�H�fGp!� �+�$�XÆ��޸pt ąXU!�$����2�P�*�µ���¨>!�D�8�ys�g��9eL��HK�l�!�$A%ٮ���Y(X�Y��G"M!�䊌'`ÕS������Q�!�"��1q��1A�a�r�B�!�� �X�*��4Ӭ������n�\��"O>��`�N<f��t�-������"O�@k�*�q�2�8�,��6��A T"OX��ჴdS 1˞�Gd�Ӥ"O���D$�TYhRj�I5r� r"Oj���`׫X���؀)]K80�$"Op����-�����M2&��"O�u(�dS1djTD���ͭu!���W"O�u@OC���J�R�j8hb"O���ƀC�y�,IbBnN�vr��%"OJep$�0S�"!m�-VX� ӷ"O�,0s�ĶU�@#q�ȰL9�E[�"O~EU�@z���q�ɛ87*F0�"O���C�L� �f!
G�N14��E"O���2��l�
���W�-�LR�"O��{��͵/�
�(&#�$�ъE"ON��n\����Dc�E�<�w"O�ejN =��Q((t0���"Oj=qf�@@�(˵�-6"��X�"Oҥ�&�N)&+�À�������"O��p&',���� F]�c��u8�"O�`�����1� �=�L���"O��H�	����F-R�8�q7"Ol7!�U
�t@!KR8;�pS�"O^�0��("�5� ��5-6RC�"O���u&��/f�M[ǩ�9�H\14"O�:��R9S��&�ܓ/�x�u"O��p�쟑k�z)���
�7@Es�"O*�r�2�6,AbI�9|Q&Ep�"O�Ԑ��0MV�PA+�<1�`$��"OD	i�䌣	V����?�p�8�"O@!U��2A3B��A�λoq���F"Oʭ: ?��mR��˕hmD�"O�X�넪q>���q�A�U�#"O����N�0_�$̑��I�ҕ�c"O��5�W>���#gLP/V�� "O�x�@i��Z `R� �9ZG@uR!"O��6d w��8�7o� t�tY�1"O�AoL�.P���㈜�m˴���"O�I��"�bcgՑ�Ft�"O�ix���
Z��7�E�4� e0b"O�֎ �#�L�Y$F�Z��ñ"Of����+��8��E-���&"O��W�P��:q\���Z�"OLa��a$��1��b�%�"O��X5/[l��8C��-w��-��"O�/��a��L4/�:��S���!�I [d�r���X�:�-Z�V�!��,D�dE�J� oJ�Cv	i�!�Ćt����əgk.��_�!�DΗU�8iS"��'F�J͘Ӏ��K'!�d������I��_?-C S�'!�$?�F��Ǎ��aO
�'�V>U!��ɁX����g6�:����9�!��+�(�aU�ǾL�'�ͬ0�!�ĖW�!Q�i�>}��8q��,�!�����t��g��T��M�bÅ�{4!�d]
���.F%�����"6C!���
fcI��ڸv�u����M=!�D�t�x��3�Y�.����5!!�u�� @V:���,Ay;<��"On�p��K����]�@�J$�_��yr�ˊ%���``�L���8��b��y��FB4.<�`FRj�������y
� �<�r��{vbT�&�7�z�"ON2V�֐U�֨Bb`̏��SP"O�]��B_i�v�bp.Q�i�x""O�Y�a�>3n�����<&N�YP�"OB�۲�T�+�`dz&		��<P� "O:蹲L�}_�飀� X"l0�"O:�	�J��0#��y�f¥#����"O��dL!H&
�E�F�(]9�"OƱ���
��Hu��V(#��{�"O�Չ��P3Hp<��@�n��ؘ�"O�hDCز~v�<bjӓ^��d��"O��s�a̮KiP�RI�$k�b�H�"O�h�GR���]��	�b"OZ}���S��(s�J�"��i "O�Eᓈ[*�ʘX4(ޟ}�(��P"O������3�bm(�g�����"Ol��N�M���V�̍r��"O^���j 1�x afS+QT�}�v"O�uq ��b���#����x&�0p�"O\�9R.�3'D��j��$=i�"Oz�*��*M ��3j�4t@ܸ�D"O"���GI�">�ćX�v�2$��"O<]���g�.�6G[�r2a��"O��r m�>B�+�g�+Y�h�"O
<���ǨGJR<���'E�|Y�"O*�P��[\�`���^���A�"OP�k��L�p��y��Y���r�"O�apD���xiN��떦_�z�P5"O���a�¯xЬ�鏼�U�E"O��Hk�m��I�@Gԓf�ԥ:�"O��b�֟-������$��"O��"/�=x/v5�o�5o�����"O�S�"�(��qh���)Ȧ� "OV��&o�k6������}����d"O�I�H�<F����U!���"O��h��ա+w���dK׫�v���"O�Q�q%бr�H�%+�P��trQ"O�e�tj��.��@D�S6m��BQ"O�p"���+*^<�bh�Mΐ��F"O������vN�)&hޔ@�.%*�"O@�b +�8Sd���"�2�C "O��5I
$\�Ha��/[V��i�"Oݓ4��-�X�9�CZ�X�~���"O�d�@��z��U(�Dy��ye"O�}�^<6 ��B���gpp���"O�J��20���ir�4iY�����~��s��F�&&�9�E
Tp�!��Dkm�+P-L�n�Q7	�H�І�}�Y�V%�|�R�ǧ>U�A�ȓ)�ڕ��,c�ar�/�4لȓ0�D�D��+*�X�y�FЍ0X݄�>V����:��퐄*�%@W�<��3�\�z���O�J�!� �%��qҠ�MˉPlI��L�'�ȓ0��1UP*!��A!�?/:���%��	��*���8&+����h��B`.����G���1)�y�����&�j�% ��ՙ��5R2�p�ȓZԎ%�g�!�y�5*/ \U��v��z����B2��b��;_F��ȓl_���+�+f����")�Q�ȓF�JH����T�v��#�>�@L���<�cAbJ�i�z���m֮fK(8�ȓx|}���L=l�d)]`� ��S�? �t���Q�vtIѶd�I�I��"O��� L�꼃".���p�"O�8ȁhيD<�U�d�D�j�TP�"Oh�rhW�#R� �'�=qL�t��"O a��rcNU��H.���"OX(aA�� ��0���S�0~���"OhVJ��(P���!`F%����4"O�L����u����������Ԝ�@*T�)�'C��A��ǁ$6�����n�1i���ȓ"�^�چ�R9j+�8s�b��H��|�ȓ{��Y5�&db����kș����ȓ:����!��&X��B�)X����%;T@>��B�\�F�ȓm��ܨ��
��ȫ�݁"	"q�ȓ4K\d2%^|Ȥ+c�OA
���l����Q&2Ga���D�� �ȓ�5ꒂH"A�S��R�`�$��}C�����3{�ĩ�7@�(����r�'u�ֆ.B��|2uH^�wcv!�'��2f��	��f)1y��j��O6��'VAZ�� ��*} D"O:��V�ðO�y	���H�nM����?|O��Kf��
>���Ь,T�T2��IFx��8w.���da�Bi/+Ӳ|�`c-D��%��)^��C$�Q�!��ajSE.�O��5���`M��Df0���ϝ�D��u���J�';|u�e�H :|���$ߕc��
�'�����Je8	�)`@�E�	�'PYꕉQ+;ܜ�9���&\70��}B^��F��c��^��y�c��r���0���6X����'�@a֎�=*�t���=^�@|3�'�ў�>	�g8O\�Cr��|y($8�$E_�R��&"O��ˤb��بƣ�%WF��W������WL��`����>Y~�� �K���$?!��V����J�D�0�n�S,E�<��M�%x�4D�AF�1b��]
��K�Ą]���t���3���.n��Ƨ���t��C�<�I�����vQ4]�a	GG|q򥊓&a�4�"a!<O: �����xK�-K�US��3
O~��R��!Z�,�w�S�bn����.]��O�'�Q>�TC��٦5�qZ-N`��Va1O�eӌ�#Z�>��QJX.��4�t�%+K!�( fXa�d喵,���"�^4VF�'b>��=	��I�(E��L���"-# �q�,Y�E!�W�D�VIq�D�jJ<q��]	�!���c����&��ָ��T0"�!��3.�t1����J�B���KܶO"�&�Ӻ���s�dp���B�G����+
&a{B�<�I�R��B`B%�4�0r)��%#B�I<0�H��a��h>��T�<s�"?��	ٻWg6��(A+n&��\�@��4O�c�Є�xy^}'AMU��!�`��\4JC� F�q��W�Z`����U�pC�I�:�tB�=�J�L�3Q�B�I�Y=��"�X�������=��B�� �V]"a�]K�xX"��$�B����m�q�;]�̚�Ӣr+C�I��9AN4#^�y&����<C�	f��SN�-*V ��� �2C�ɨD���o��"�
�H�C�I�� p��³D<Ri��A'@��⟠E{J?��� 00(�AWMS&
��bgC6D��I4+g�$�0:ّ��xg�������Sg��{
r��r�I6i�*�n�8=��IVy�L7��� ���sɘ'~O��gnH� �0�"O���G5�4x�Ǜ%2�R��Q"O�A���ɽn�)��4��i�"O|���(��b�v+d�B�+"�Ɇ�hO��C�sd���4����oY;�!���3#Cr=�u�Qfet|YQO��vl!��S�;���R,1eZ辉Pq"O����� �`q�TQ�ե(Ŧ���"Ob蓧d/}�	�`��-Y�R�:eQ�|�	�qO��<9�hJ�
�d ሒ-|��8CX�<)oBzN�s��+�<�ÁS�'Nў��Z�i��L'1�~� w��=<��Ԅȓl��%�fd�W��8uo�:���ȓE�pP#�iQ `�:���nN9"��F|��ӛI����Qm�K�^�j���i{��IT��P���ػh�ԘP�b�6f@̨ 6D��˕#��wD� �U惣V����5D�$K� &ɒ=�D��}��s��h�4�'��' �	H�i���Y5$��X�!��$���c��"D��{�d�>'vT���M�I�$�֥�������E�fE���&s*^�У�#���?a��IL+[��j�	ɐ����R!�$iO.D�q�V+��7��8����c���l��kZ)� KV>�~�i&��!� C�I�W�Bh���F�&�fX�]��4"<ɍ��?Ej�`ǯ4PJ2tB��78�5�%4D��	Y�oF���F*S@N�� �)�<��哛!f80S
A%���#[��B�(G��h��ز$T�|���� v���Y�IVx�l+�I-3�m�$M�??�8����+�O�r��P�v
X���q`���N��ȓO2���"E�/$���G'�Q�^�mE�������yR-L�#�<��W��=w�eAa�yrON�{R,\X��JG�vd+4'Ђ��D"�S��ͪ�\9?�f�a�m\x� Y�"O�@j���p/���5̐?P��=��i�P���IG�� �S�̴���lH�r�F"=YN<���-��Y�h�@�o.xL�PbW/��Z�*B�$�ͳЪǗ	���z�c�=1����?�	�B��y"���"�� ��	i�B�(Z��B�J�9f~p03��^��B��15�,���
4'��H�>��B�I:J	�a�nCV��R�*G�02�Ol��$��'+�u����22�%	B(�t�!�Նh�^��l��Y�ظ�IFR�!�x����ؘL��80�hKA����'��O?7	>-m�R��^6���&�M�V�!�Ϯ�������{yPyJƦ�*�!�dʡD�y�t���<��S�ʎMa|R�|�h�2W~��Ȍ�;�
��cO������p>)%ۭaJ|AD)�THr�j���1�OV���gQ;<ul,���2{�c�"O^y���=y�9��E�V�Z�E�xbS�$'�b?��n�_�P��,A�]�0m�6$D�l¦��&Gd�`��+L8I���"D�I�AB�;��K7!ʩ_����%h2��p<�AJ�3-�m�G
��Z�.����x��P�)w��JLjE�C�
�y��
��Ļ2�@˪���熛�x��'�$	S�
�78{̸���H(G@��B����>A��$̘41�j�:� ��Z%����y�l?�|�����%�0�x�N�yr�9�h4���?�T���א��'�ўD�'S@�B��ߒV���Cl�5~0h
��� �<��f(/�9&'�
����G�Iox�d7@#��xC�@�Bf���c'D��Q��T�<̈́�h��_y�e�$�#D�X�a)�9>$r]ru�IoP�)���5D�L�@̣,4^�a�LF�+m�ca3D��3���	-h� [u�E
ʐ-��l1D���g/A).�����'z�����.D�0zQd�'=� ���@�8>�����1D��tk�o.HcĬ8thf���A.D���D�I�XVC�"��)��o+D�(jFJʗ!�D���͖�f�d�)D���!�Y,p+\�W͒�$��k)D����Ѣl+�@����J�{DM(D�,H�n�@����˺.�%���&D�"-�� ?Z@�Wh�c��pH��1D�l�M��h��6sɫ$@#D��[G
Y�b,�h�r���^޼�tk>D�,
�g�;yX)��OJQ����1D�@�+�Ġ#��҇��
�0D�t%�H�6��\���3C̩c#D�,@�hֵd�|��֎]�pp�eHE?D��cPoի2={d���@ Lm	�(*D��а%V�d�*5�a�p�I;�/+D��j&jOl�r�J�,��g�(D���g�W.0U�����3��@���1D�\СNðr�ޠ��Vek�|!�k/D�D���^��ʵ�E�̼�'�?D�8��F�*Q8�k��M{XS� <D��)��H�N/9�ʓP��)�U�:D�8!������IqP�Ǘ|Ct��W�8D���/�g�p���8m��@Q�8D�(���o�z`X��C%4|��9!7D�l����ma�1���
M���n5D�\���8
�QѦb��nйwL!D�蛃N��l2!���Q��8Sg�4D�D����`�N�B$�Ͻ?���z�L7D��H�
�`��E�E�Y�wҜR�!"D������q��<Z��Z|x��"D����$��]�p�m��`�Z��u(+D���) �
P�#��D�5�qL-�O��@V��#I$iyHQk�4<c�*/_z�sq"O�) �A8?q$��3�ݞVz�I"O�p�f8X:��FH�"v"O�X��l���JH�I=��	��"O A��KT�{qP�Q��;|a�z�"O��REbP7'�� �a\Ba�4�1"O�ݢ�C	\9��"�Nto(���"O@\ ��B)�h�c4���6U���"ON�ѥ�7-�|D2P(D�Jn�1�"O�[��ݪt���a�A��;8�y[�"OjS�M�MHaP� W�-�x��"O����p_?8$H)�G�
pν�ȓ�P	j�ĉ�fF)ۢe�%M�nȇȓ`����"޲(��XCt�Ŝ"�Y�ȓ,OI��&�/=|��r�M�3A~�ȓ�}�æ+S��� b�3i�=�ȓS�x�1�L�1������*<�L��e4��ө7b��i�I�N�4��Ku�A�S)3	���k>���wL�R�J�-R,�� �lW��`h��1BZ�6}�hD����~��Q��&��I3��3Q1�L`�Ȥ]�q��E�����&B���S�O�	C`��.J녁оFT4�p�'w��Xf�Ǵb Y5@�8��5�-OTp�1�(x�;�H6O� �1xP+	#����ǌ"C��6�'D�X1���
`�AW�I��rN�;��c��v��t��I-2�Q����n"�}ᓀ� -S �<�e@�/ <�i�Dl&�u�K|
���,��3��N,? H�x&�t�<��,e�H+i
%f��|���1/#��b�̀�V��p"�JφȎG��'��I ׆	�/�D����B��&��'	���*Q�I	�8R�+wSj�0� H;������!@D��"��׊a	��G}�`T�C���b�E�5���BP�+ڨODA)�H��(gX�CsJ�)���E UFS>���UH�:��A=y|ȕ�ZMX���I�Xb�`���2	�,@$��=�4�VWS��2�`H" @����C�zSx��%[�7�8`�?���B$1�|h��e%��unU}�<��☨P���a�n�~80�BA�4o,��Ju)���w��.��U�O��h��D��z�8�O�(+`�R)e�,�Y%�N����b��h�a��6��'_D�d�%�ـy�te�`LѮ�uz��)Y���������z ��&�~t��;_\��h��p��<�CX�f�(�$�.:�`��
J�1�'�f�)�
K�{9�)ZFIDHf��M��w���B�X�.���g�bU�5���,���R�?�I�^[�CgJ�'(�����E�Rf�&%+��;2�;����F޴+`�I�>'K��c�^�%c�u��&$ !��/@����y(�" V�)�#4Z-y�*Q�~����Nt�����W��D���D���y�h��/e&�;�d�\��y�Jʚ@�l1�r�ED���k>�a���1+o0�c$D_��YYt��AĜ�B"LYD|Q�i�M��8t��`�b"K�I3ȕ(r��`���-�,�`���>�A6���J%�G铟f�d�XT�,au��j,Ց{�&�9��F`�fg�+�T��)�<a$Ƒ�c|���r�� ����#��e���.Mj(x�L����Ϡ���q dUȈS���Q��ŭ+Ed<�!ۊ#�����3]e��� �)C��(�
�IT�-�FX:�?9��{љ�ń&-���C}�֝�����m��иU�\&�<��SÒHE-���Ϗ^]�� ��Қ>��4�D��o��ذ͟�N�'=����Z�H����)�%l԰yn�s_Phs��y,ݩ����TN�iD.IJ�O�?��]ϻpc4)�ȄHĦ���Lwl,uK���Ҟt��,�N���1���|:���Lξ���h�pl0IK��A#Pt�y��ek���!�|$��nZ.0�qЖ�P80eJs/��_N���^�����ͿId�r+�"[6yS�'�^��Qm�+�,��S6auFP���о��!jR�%W.MC�'E_
��1mK��"�IR�(��U���i���Gh�'� �hX7Nl%�'�R ���� d���Z�|��1cID�KE�4����0�1
ԯu_�����o$���HkڰZ5\�ŇI8 �X�P��w�ܟ H��&b����>-l
��L��WJ�r��>k�@�R��N��u"1%��"a4��fi�?/h$?�ݻszI�XY���ҒU���P��34��ԑ��]�R�$1�%��?C��]R�-yeK�]���
`ĔD�-7Ct��eI3 �m�P��B���R��X��(30��?:�GV�%�r��$G��dx�&�A� �0��А�:�0�Ů*��I�=	 -�7�J��b�E��l����%��3�ҕ�#��O����r�[�]�`�gX�<�Mⴊ�,s���e�6u����-��H�������U�P���Y�9������M��%�􈗁6W�,Р$Z�y��A´j:�d�4�������5E��"����L�!���k�[�@��
¿� ��t�[+K���ňU>6�6�ې�C-Jݢ��T���]�T�Cê?���weL��OE7zӆ4��i����(�Px��AL�DA	kdN���)ʥQ�N)����?P� !4��h�ir%���
�f�+��P�A��qʶ��L!��.G>T�	I�i[&m��\�'����OZ;{���pa����6w�x�"�i�u!QaB����'d�N��|���#n�Dbv�.*����$'�	bL�`�J��,K�H�Q�L!!D�=b����ʃemI(�A&7�,��P�ʈ"�̑���^. [3CH�8
8��x��I48qpB�$�Rұ��#Lf��4#��p?�R`�=�� �'��	c�LL�͆,����"��h�H���rаڴXqx�Y�o1���"cZ�y�͘�QbfX�p/ۭY�v�8]@0���[r��"쑃=��E#�HKN"]����/�1���شR����d![z�����8��ecU�
K4i��p>�����0��Ί�"1�Q��I�n�ǥC�:����H��#�C�w���,F_t����	�28(.T��g�E�t���͏L�%G{�K�`��!�4'�?�֠��.��'�д���̬"��YV�#Ktb���(L=����Qf��x���]�tS��� M Q	A�%|��ak�,�O����I�@�X�G	
��"@��:L�@j�Ġ~��tK��6V3����d$G�@ ��)�� H3�3�B�;r�y���P��U!`���1�"O���˔�n#��읜L����oI(Y�L��F��m���$������u�<k.�5��\N��1��Q�%��)^�`�UL��H�ԙ�Bn]5Y�~��%�K�YǠ-��l�9)��U�����FM�`��mq7���S:�kc��.4��� MN ?�����13N2�"��
��(�c��p�8�D�m�'#���a������ˋ_V��"�)�l��
،ؼ�ȥ!�>)�)�����A-�	[\��_�-�L�AÂ�;<�|� ��``J���lŚ1&�`��/�~�`()�2�L�A�I�8u!aݾE�e`ح_����A
U8��-[�Y����A܎K�lZ8ͪ]�&�A�Y�(��Q�Ɂ{>qȑn��*���H�iH⬴)I>A�	�J䢨���Б���6�؜�DnJy<yؑ,�$L5��*]�{)XTJ��޹��u�q��8����w�ĦB�𭛀l� F-����y-^Db�韻��7M�0J��\�d犟}���$Eخ0=)�J�7N~�ؙ�/�)NW��z#CP1I��T�$G����T��.1>�T��}q�!�e		A�j14�A
=�H4��g^\��0T�BK���hĂyy�<��'��kZ��ab�\��80RE�9ZS�D��U)JM��΀%X������aL���TZ����Z:[_�|{P�#d8�Ԡ0��x��9nJ�-:qᆂI��<�� �1
�
��b	;hA�Z�� ��#Sώ6�J���B">�ۇ�=5��L����Z�|Q34b��[��4�T5��+״@$.��
<6��(��I�Ҩ��ꐇ>�v݂Ēx�O��ub���)D�#_ �
� �0�F1� ��^�VtyR��,[��Xr"�E[ у�Q��\ɪݴJP�q�ˤ{sf9�5B\*]�J�;1����S�]!��	:j���C$T��x� 	̷xOn�ˆ���8KXu�q �$	��Xۇ9o�����6�P���̷zFz�N�L-��-�0\��ધ�5n4��t˕0(� ��+�/xI�P��f�Y�'�Zi�b��k~�J�3k1��+��)H�����"�j�|
�H�B��|���z���qÀ+di��iʤ�$:CP^R`Y2��'>�-x���"'���꤄�h_()a(��f�� 1$���{x�8р�W�^�*)��Gj�a�@��L5I%ĩa���D�6sl�P! �R�P$P0ؐ"r�E��ΎLL"�bA/0�����d�e�ߢ �)K�1�p��1��Y$�b�`��x�P5��%��!�j4[�ś�Qի���貭@�m4��(h��V
X+��v�9�	*j,f��ҨW���;���=ҁ�Fb)�be���8p�������i*n��R��'��sghX�>��N
C2����ٱ_f)BC��b����P$+< �1�`W 7�����r;ʝ��&� JO\吰ף��	���i�1�tD�
[jbA`r>�����"NEJ��شA-D#�G8a�H�[
��
��'-��h���IQPɻ�)�6b�9��B݉.�}��Qc�1 ��#���r)P�[��IQ�sx�̓(�y�u�O�3��ŉSDd�T���6^��ԅ�	�@4J��@nqON(
�)N!4\`�9P�E�-��E�$��"P��zc%G��ə�!ڂ/��L �ჷ9��3�l}�2H'�8�N�vu�y��`�,qO`�1� X#jN�}��%�&exvl�7#�"�)��d�|Z�hR�GG&}0b୻`��)I�!7�����I�̼�w��ZcrX���]�1���%P}�~��e�Ǵ\�		�(Y�S ���<��:�bX2Ҍ!���yV2���ՠv�������	��yӀ ��xT6�!`�*Y�:)�E�:TGfH0(����%���p=�$�C��f�tbB6����eb|�A�� -2@��Ȁ<_�7m.b7&����Dl>��c�1��&Â�]�B�8ز��a�������a�)��}�!O�(�&���͊?V�a��C?�α���.���`T2�"X�/��{�N�2��:N�1�=�̵��mD/��A�W����D�K�b��58��:yّ������*{eFP�t�3i� �����=m����,E&�V�9rc�=X�8�c���g�T�0rjD 1Nգ�o�9BtNA��E	��O��;F�@=A�P�{��=��Yy��O�bG�#4��?�Q�Iܖaf��v��=C�^�3��9��MQ�=gN���b�o��l�D'O0J���S$�%�����-�OJH��L��	� ;��O�7|hu�VŇK�=���35g��j�7mAZPؤLP� +���(1wz]��4�%,Ž!�h�j�f��cc���'�hf{�l����,d������F����a�&�rs,��[.6-��gH(�A�l��S`��kRo���a!V$C�1�fe5F�O��bো�&jX+P�K�A��)hV�ɺ��De�N�d;Z�����a�p�Pl�U	��"�A��d򕫂�)�
%��J�z(n�yM$Z�2����X���ׂF\�'�!:3mJ�]�6�Kl
Լ�2�`Z#0۲X��B<�� �mJ�%�c
6^�"�#���ܨ�J@� 5(ݨ2"�8=��mj�G����I�v!�/+��˓�'�����_�1�*��Կr����$)�x��Q3��4H�7(��N�����4Ko�Q�qfêz�	C9�8��,� 6�
]J�Nq�fuV�' ~�3���2TC�TV���F���`1hE�G�NST� ̈́
3��$a�Wvr
���E���\�`��c4nQ!W�H^�h�%4�L�JUmߓPFfd�FGո�O�2�)�Ncz� %꛼#���`�Ϩu�}�􆁯6�XLh��1��#2lU���3h��0uN1cѨγ'�Fuip� �0��PyU���ؙ�'�3r�v�d&O�V�d%p�	�,t�cnֳKl�t9%
�����R���t�b�	(U�8E��ѻW56`�5�
7̞Q�e�)D�kE�'SR�ѝE��ɒ�3X�aC�� �%�
�9��/ar�!Å5#Y @��ПB����FV�7P�y{�w�NRF����aH�� +'Lə	�L���E�7��}��b��~�PP Co����5ƴ[ �I���U*ĩf�XJtd땂\}��t �@k�����O"�Jb -jxU�4oL,2v�(x� �iܓ;m�` i��bEàK��}kr��sf@��\❏-�����<y��yȔ̆�B'�٨PY	Y���7j�O�j@"��$��n�{� Y! ��R��Z'5h>��Ӎ�6��2��wn�Q#���<�r�s �"��j�fZ%0c$��c��5��}:���jB\�:���)�҄�o\g�'.Ѐvd-apP�bZ�8�A�Z1�Z� ��W�y@⣌ ��%���Z��A%݄#<����۳�V���R�YB�m��I�/�s 
5���2!N�"�<!�$�8Ƙ 5L��%u"}����-(?�1�F'
�r�q��]�5lj4�"#�"r�`h�������cf,5�zǮǥ�h�)1��1dd�	�' ��)��:��8R�mH5l(ȀBb���~r���nD�A�6��"�ǟOJ����6gDan�l�Z$a�"�N=��	�$>g�I���b%
���T&U�#&_�hڱOKR?
֤�*�'Qc�M1a��hAh��O�Wv�p�]��T�Ѷd>t��ӏa�qq�JE�kHx�s!��R~%�+Ť_ܶa��)�&�Pzd�3b�^X��-[f�\,&ϥM�1I�#"�\bt(3c�X��4C��xb| k"b�`�� �
�J:"��G�N�rT�٢,,@����	6��qi�E�����/p<���)B�|���㆙�0�ʀp񅝀��D^�5�l�鄦�*� �$a�>s���Y�lW�JgB��	E�Iy0H�
�^mr�C�#�ܖ-{��h�$��x�*��N�Jj����E@@p�w�S�p�,�4�@-��l�[�|��'ꆕ]X̴�A(̿pKN�*W�{�hH��E����{gd�?�5
/)m�� Ħ�:&��rUK@�WH���Ϛ4dX�fÏ�6y��@E?j��e���ԣm<��03�QB��<!���[X��?V�)�+Avj�B�pG��Z珂�E�������GE>Hp���(u�<L	�
.Et�;	�	�ªܽ��qSMC1nIqẻ�jhX�Ia�_�@�$�H!�6�	4A�(� �×�R̎x�����a[$G:��xr�Ƅ/�6��MO�}z�����ud\�B��S����qA�����@&�,�&�!эxp��� 0�k0�ˇWR�U`E�f ��5P����
P�"S��Y-��!(`�B)
��b0� �R�� "Ā���� @�*0�E*H�@8�dr M:|f�0Hj��_��DhT#ʧ"���K A�"$�5ʈ�C=�h2�i��э@�r�4���!ɥy/�U9D`�� �	�8|�h���F�Ӧt�<<�T�D>/��&�e��,���ىt�r�{�m��1Sh�y�#Y���(�n;3� ,A����d��4�=��#M�^KVt �BՅ�n��6�Ug@�RRd�P(^M`p�o+L��$A) MZ`����l���b��eF�RB��U�ʍ��gۡ=c�M�"�@��x��]:+v�	�[�b���hsV�\�@b�;�J�*'n�=;Q�P g�FU����N�..I>�ۣ7wb�qtň��������9R��}K|uaB
»8��Ӧˢ�t�5�l$�2(�� �F�'j��P���C�Ҥ�ٕ}�zm��ُ`\ɘ)������\�z�X���V�`s����n���GJՈ9d�I�V�V��#}�w��9��96[�D",�:b���+�Kq�Pt��I���,��M�~*fi���y��I�P�����ߙN����K�H>�l�!��i����`�]� ��ψO�q �m�4c��4cV�[�����q���ٳ؄Ƞ�̟���s��a�Y�t��y���=h�)F�� N��q�`�*m~،�����=Y��3r���O;�@���P'>��P֏�+���{�/$��V�*���s�ı~)
q&?�م��b��낦Ѭ.�Q���(���+�G�6�`}�O?!Р�0��v��$9�~��C'D��0�>d��Ha�6�3�j�<�I�P�
���,}��	�4'��ؐJ�K0����@	Dr!�d�q�>h�5B0��tÖ�I�qO�e[�d�
�0<Y��T�C.���'
��S& Rp�<q�n��c��E�6���?��L#R*�r�<��/Gvs6����y�)�J�m�<���ՅdAV�����6$.8+D��d�<90
�q�LВb��:�E�f�c�<�-O�T��.��=/2���#t�<�B`�!��	EA�VF�+�#p�<��h��!���p��S�))(�vG]m�<yS��3J�|��eS�FE�T �@�S�<pL�eF*0�+2G~
��㧅I�<���	�EP8���T�]�LACE �J�<醇=2"~�0�)��P�a;���^�<)TK�-O�v��$Ϊe�����Y�<y�50��ȩ�铩\��&b�P�<�Wj�h��<����'1$�����g�<Q���NRbi��4ɂ�Q�a�T�<��ձ.�-[Tc�|ih)qPK�I�<���,#�̰`%ώn_�bd��@�<CO��Gz��W�ӉY��@�1�F�<�de@(?�`��!��_֕	�C�A�<ArkI�*YH��r�K0II� '�t�<1��Y�yvE�����T��~�<AB+�k�~p�!�>�RL)�L�s�<٠�A���Y0��2O�ݳw͝h�<�'�ZqX@�!/��L����gMk�<��Z@,�
f����2 �x�<�'�V<I
p�RR�V�j��T#�O�u�<�$�W��r���F@��Y��v�<y3��;M$�[�LF�}Vty��Bn�<y�%9g��	�$�*3vP�L�<Ar�E�(��U��J���X�I�<�â2��4!pf��V��t��k�@�<I0�C�/�̉᧨����)FB�U�<)�R%i�݈a�	���{&?D��"`�p���s)�6@�X�4�<D�����L={�>��3̈��lD�B�8D��a
Rr�h��7j$,�� �6D���	�xxD� t��?���2�2D�t��j�@\9V`��J���huM:D���A`X�;d5��+J�f��܋T";D���$Gj��1X�a��Q#�KRG$D�3!��-w4(jҫ��-}8q��+"D�<ÂB]�74�00�F*��e�7D����V�D��r� TT!,�9�&5D�J"�>���R�ԗ�{�A6D�� 4`Z�'��%H>w\���"OΈ�eI[�u���R'�	Jn�x��O��ˤ�: Nr�O�>����<����"՟m�V�b�)'D��Q#i
*�fp����G>|�2®<��!ʶOK�(�	K��0<��' y��P�@�i�b1�/cX��r 
�D:i�k�s��d(���5�r�"'Dӻ%���+�';�9BG�J
k���>G����ߟo?�2�9L s��;��ra�J�7;��c�L��Cg!�ěM����!e�yPf��7mȼAɔ�Z-Z69Їe׾Z��򧈟�� h"��q%a�):���tD�?�y�\��K�0/����HH'{���`$�~(��BO�)��\�G���|F|�B0GL]���,1��XB��*��O( c�����y��$7������C�B�64�Bb��`ࢱ�X�#3���OB�)!0���oXt9�� +ClL���G�D��ŗ����F��M[S#^	;�<���BP3\�İ4�3b��Z�M��p��͞����I�!�yBI�u����%����Bá�� V��b�ΊX^ɘQ� �5�5��N�����lp��p����ㆫ��}ȃ,W5
�$�"#�ɚD� ��)��G8L|0I��F�ΤrgÖ�4Ḵ�� ǧD�Qc�4T�j̊f�P�А��I�i���Ex"m�?3��X�Ƚ<5�<�%g�V�5�!��Dӎ�'�<�alY @۞��#�΢Zp�V�M���H�!l�x5�M��39"����W-O_(�P��VBڢm�?!b([5ObxPZe'�/��)/�N�Y�%Q�k����\�\����O�qQ͸ F؟o��ٕ��(+�Z�	'e�
l���џ�O�k�����6S���LZ��V�|����-L	m�h�
�'EЖ��7-� r��}1�CJ�c�$�Z$�~��0"��q0��b��|��!v��QQw�g�,�B$-I�#�����%�Bh�ЄɈ�<���b
�z?Qs�ON,řE%����'�8-��'�RK^ag�֡{c�I`�R/h���o��x�b	��Q�$�فbֻ8�����KV�{b�IR�y��{�p-����> �����V%
��	�pg^/E%��C"o	a��Ix��`�H?#t�A��B�qC2й���1����paD�I�lɒ�J�i���`��F��$l֭�d�ƇJ�����	M�z��@j �jz��i�Q�Ė0U�"���+�yC�]9bLC� KjkhS�~���ʷ��"ěd	�`�I
7��_��s��0�*�qҢ���I]�Y�,�GK���M� �Z5X$��k�b�j7=��A�BJ�v.h�S�l��y'EO�2��x��Q�!���"*X�)Pb���MbB!N�*�����O��l9@�P$'三�*,Z�k�P5&`EQ�F��'�2A w��M���,(�丂��$���#/٠i<J�w�2����?b���`5 �,�>Qb�	�U%�K@4R��rH>A5�E�Q��"���%�Dye�1V^\c��\�x� ��^�%�H�0�4�`�2@�t��9�(O~����A�=�M�wlÈ'�>���c��zΎ-	ŉ_�5˴����	��x��Wl�V��q��H��[�[���Do�d[��w��x6Hp�"XkLH�|z�o_ e��EQ�k÷R�~��4�������[����%�]>o�̤�f�0<��ŉE��
Y�����(��ksT=��/�����U�ܼj�֐򶧕28���ɣ ���05���n�8���ɶh���D�k�BU3G�N4+K�I��yb��(C�y�D��]F�IY"�N��Bq�eN&p� �`�D[� �����^�@@B�ÎeJ�iJ�����]�̚d�b�J�M$tY��ʌ	��10׮�h��������j��В�@���@���w�R��F��I�d ���v�������CH�a���
Q�x�Lΐ
�>E"�<8q�dl����Y_$0`�I&�j}�Dg&y�N%�E�� 熬0�,�N~|\�lԢ_T0 Ү�����w49Ku�A9Q�> �֮�e�����T%���o��ҧ��R]+F� ),l���7F����̜6d\ �q"Å:���r3d��\����� -&p�s͍.2K���%�O�����X�:�Q�뒯Xf���>��W%^� b��}{�*��͎�0�<
f�:Ov&�1N�W(dk��
#g�����'��@��!C�cT�$j��I�!6�p ���6R���"ޏ>���c!oU����A�N�ƈ�A�׿�n�a�E���F�:�NR!jb�^�r�h����7GF���	�  :w �?4�Ź�װ_�bM�P�w�A��#^{f9���W��MԎ�)uzȻ#AN/a�ɺ�wD�ɰ�)ʴ/�d�S�ٙe��+�'{�=�sjK� 6�8S��Nb	�vg =��\PK34K�E���2j{�-�j
�<�#$��Kv%���'��z�77�,��b�,rw��BӓQ@pqEO׻=�f���Ա=��IsJ�-ӛu�X;b���AҸ$gX��"�Z:K��&��s,�SR퉂t�T-#�i�?W3���%��3�Db���Aŋ�6�^ 	԰a�H�3�#,X�cE r�N}(��o�ִ@�I�E��L �f�����͋��>�u	��bX���$��Bg��`c�P_�،QV�YIx�i��
1N��	�dU�%DFo��hCD�߼���G���D���A ;�H��X�<!�
1�V�3f���& ا �%_���
�9cJ��h�|�P)%�	5�@0����,<�kA#R���*l+�@� ������#K��Җ 
	�b�B��������)��T:5�G��,N��k�Z,�����a�a1����#���
�)мWg.�P� �e�r�R�	�.��Gz)�$ٲ��%
��iV��X�I�6I:���^�fԂFŐ/|.����$L,�}+�+U_ݰ$�u/D1�0��st�M9g�OQ~ȋ�Ϟ;?Y�Z�g�y��4�I�(<��Ҽu{�d䎏�.%�q!��ٲa�0i�ǎ�7k�T$adB�ք�7~�T�n�@(�e9شc̎A���l�ȥP�D�/ X=!&D:Stf%:U ^�-�$��В|B`��/�(���b�aE(�5��Q ���B�B�	.\91d�ɲ�� �]���Co�
2��� L�?"��!��;7���@3A�ʺ��p"����#�؈6��m:� ��Y�G�9h�d���ȼT� T�A��at��N�����{�oC&W�i�'�i�n�@H�=V�,P�!dx6+$'ȄS���F�H"b�¨ �JðDy�lx�Icp�<F+��:k�')�Fx2,+�	�%H�`&�1xLIx��14�0�1�AEqn�-�!�f <4iҝ!T� ���OPqhv�3������p�"���M,z�>�;��@��
��c�Q��#V)�$dt�[7��2aTx��ͽy��;3+ ������T(���.��6��E �
.l1�>~��<KëY�!����f�P ��Ӈ�� '�T�G�ɴ	:8����$�ēh~lx���,O��{4�X ��ٖ!FE]*�ڔ�K�BFz�+��͏zz~��b]�S�ԈĎ�����/�F�sA
\���ъ�*����R1?���A�OᡄI�/+���b�lߨ�,P�M���*ab,'N�f�KL�����."��z"�iڨ���w��݉�J��~,`T��@�Ff~�S�
��K��bǧX]xt�8�£>�Djޭz��i���-�zS��%������ta����^�,�7�1Fa����/J;Ǜ�g	�j�36Kȑ^�f	�BcC`�i8�H!��<6%F� ɖ���PD_r%Ybk�&"��U;
�ldB䧈
��=���C_Τ�� ƦC|��0�\�'8����'�fxD'ɍ������H���z%�<5�,�Hs'R0H'�'k�Ib���e�Z�S��4�*�ϕ�6�>��S�K"��ɔ��H�2p�� �-ұ�V�7YAynڇ�PA��O��V+��J�LI�P�ɀ'Zb���R��O5ޅ���{�ܠ�!$Ũ,퐡��c\�%��Wk͈LL��2�x9�an��E �ۥƅ�".,0z�j��vȗ aElZ0������h�j!X��'R�y�($h4�L���� w�̵� ˋ('�Q�fK~��)27	܊����q�_�j1�P�׌�"r�¡l�W<J��d�D��9�G_=<�����e�4������$�۱C��'��OPF����B;~�$��п)E���$���G�� k�MRD���'P�h�����t��!�X��@�A��$.ކ$(r�҈��'B�`�D
K��rt�"y�D�
�B�� �-{�J8j��^��rQ�#�|����7�i�~O�-Z�^5��B�)ܸ'n�� � O�tBf-��UH�ˊ �MȄ�G�f��hSeA�1o��]�}4i��Y4;�\MX l�����Ɠm̢��2b�%C���:�h,�
�-'�U:���! _���dRɒ�rK	77���R�H�I�ZN��A%���]�dx�é�?�Ŵi�����	Jry8����ebF�1\vL4
'I��i�0��kf��L /Ś0Nn��*�;G����7e1�����,�!���K��_�yR�6Ɠ}��A�>v���Sq��!c0y��G�ywm��f֤�AL��4>�v����>	V�Q�=�@�Z��!LM�����R��:@!/!�&(�T�ɋ�,I��m� �<�"���IA���Aj�8Xa����y���#������!���z���HO�]X�G�A�B���Qvw|���u~�q��J.y��T� ��`��9h��\g����ˊ_f8毙�r��9@��Kl�'ef0�fL�L��\Z3�K �>�HTFր2k���d�
$6k�4
�O��Amh(�&LN��x
��
"�4�`$f6���r���nx<���h�"��z�/c� ����'af9P�E��,H�զA#`Xu���W T�mؑ���\mL(B��ij%h@%�&@��f �&iLY��w8D��ًctT\S��P�� Gx����6y�D 
3 ]pb�̪Gdb`�$��J��iMȩeH͏j�^d*���j0h�p�]W����V	')�b�+��P立 u`��V�"�O�}ki�8]> c����$X'�_5@�\`��� ��C�U�XͲ��.k�.ts!�C�:�J���J�_��$�F胶>�=9DL@�qp؝2�h�-u"�s��ĢB�XX�眪���
����B�Vb�L�ssҁr@��s/�34N�E�p��&��^h.`J��	)yv�zehA�?`�!��F¦��>qAf׉4��Âɟx�ڈb�L�&ih�8�ʀ�*��б�)fɠa2���ʦ��%��=�f�L���y���L�x�"���#������0>�u��\�n�"4 �<�θz&-J�Rg�./�fe�Ï�+f׬�ɀ�Q�r?XԊZ,͉���o\�L uhл%zY����ܟd��&�J4���#��a��,1,Y�=���8<2�D�'�MD�2��#N�иև�O��H�gǼYh.�ґc�fs&���J�0qf����-1F�Qv�Q�'��T�F	X�V��*�L�c*,:��Ll���;*\�w��z6b@�F��H�&�8U��1B�a������xg����ȝ$ϒd�G9ndܺ'�}�a~�O�90���$��3/�p��q��/���C�!�
L���B.����Q�"/��5ର��0)�dԐ��'�yw/�-g\��d�#�|�aaV8�p>��i�[�>��+�|yB|@c�5�V��HK�S�^�g��!:P�q΄����pE��<~L`xrc�7�B,��苊��D�O����h�uF�����0,6]�=I�%ؖ�$l�d�D�F�����6 T�Y� 郥Nܐl��c۬b�f�'�=���ɴ;0��z6�{��)I�ِ��O�D�C^�$�p�����i"�dω$��Y�
8\\X�V���J���ߒ#�`��u 5j%�J�Ď
"��9i�L�s����"��=T)���`#�l��D}�J�;/W��k�	�7��)x�0��A�7H�L��Ė�2��� nHۄ!H&+�FX��jS�}����6I�@�����$睨k����%Ƃf�r�Sr�ľ^#�˓	��1�	 �p�h�:�'PԚ��g�Ux~�*�����I��h�}��a�'�2}��1q��y�*���nߛSuh�rs'̜��a�W�����0�v��u7��c���7�2Ty����q%�ؚ��ͧxmp���J�P_��IQ� �S���	�5
��q�b��,f�Zl�WJ���@�����(�2����{��Y@	Lt�/GD:�-Q>L��ݳ�!�3F��J�F�	5 ͓�*ٿ~=Ctj �!R~8��3����a���B��R%��9�Ӵ*ɕ�� :$�)AuDݲ�d��@��H!"B��DptF�%jX9�ʗ�&��< �D�G�6�5O�GZ @8�#Lv��9kR^�FA*d��%l8ʴ�˞�&��O�CR0`xrR�N|��a�ӎZ�>Hc���oG2��q�E=����Opq�I� ��1ň��L��@A�6!������?u�`-�c��9�(��9�4TҔጓ$F<XP6�@�c�4�3/�N�4!��Cg��i&( :� x�DAM�!N2Lx޴
,�q��#�-�p�����}5D��`bڶ9t��_�2����Ux¡@�D�F�
t�L<��}8q�:� `L��Vt��T��#S�?�ܺWc�Y�f� 'k�'>5&a���.~?th�e�O�<~t��H��`�q��n,Lb7�8^My�-�%~�99��@$q�p�c���e� q�'��-�]0�Nd��5#���qV��2������-Z��|XR+b-�U1��ܞ`+�qas�M<;�xĊ�(�&��ɩ�%ӇIzU�Rf�q6ع�%/ZV*MX��+mv�Zc*Z�Y���Ffm����t>ԥ�E��S ]�VdP������!^�c�TXr��A}�ߖ�J9k��J�@3bh�E[�M���Գ`/*=�Ot�"��Xg��h6��#8��X�EѮw� �������UH��.۴]a��D�!f�1�#��Y�2���G���%тp���tn�=g��I%-*U5(�!��I�2좓�R�����?I����32���Y�#�!���k$� �A�Ɨ;��X�!]0@����2|X�H^P'�1�%aCT���`mE8h�-�o�/f��;de���[1��z ��� ��6�e�e���%��`>m��A3O^<Zd#�Λ1	D��p�^�Ș@OISp1�ई�T+2�i�}�c�NV׍��L�d�1	E��p�lM4#�Yd Jh���{SOR�1��d�`�јD�ЈF/
�5�*�X�,m݅ �fpɓa���	Ѳb�L�C�jG$)��ǟ)��	֊DJ��O?R%B��f�h���͉&&8���O�Y��1t���D_&�KT.�$L^�T)S��/M�iQ�!1E�>!�;�Ȣg"~�R�/I-�Flxp�i�ȭx#�N#P ��eSɦc?!��)DƼ�У�k�ʷ � V��/�>>Y����[�$B5���"�(��g�'�����!ZW@�P�A��J�aY��~""�;,
8�� �C�9O<`������W�P'��2k��ȒF�F�%�U?Ua{"+۹f�.��v �p���"�L0f.�@�e/h ��1��M�I�h��!���-`� ;H~�d�+]u|@ NN�BU��j�h�'�\劣@C�sw����~�7+�
"�I*ċ�i��r��	A�<1�$�3M�GQ
b�1C�ty"�_�D*��B�Ll��S�z�1��C=(	�9R�kÓV��B�	�L7�e�H�Ղ�`\�r1��DIn�9Xax��ٕ|P0G��U�
��7�G��y�e�8ohmP�ήJQ�ZրY6�yb� 3:��� �=s���9�$���y�-�5.5��7^��jb-Z��y���
��h�#�!X�М��`F�y2ㆄP��I1E�G����'��-�y��M��m �G\�;�x�X�ǒ��y,Z�g���!��Z��в�-��y��0?� �V&eޔu#�,���y�d��	WR��'��X!��(����y�f��o(��*rOW�P��T�$���y�O!M�\�A2f��8�l���	1�y2�<'��h��T2��u�A��y"8�s2�2'��	d�΂�yR��k��h��+̠�À��yr��7��B�W�t4� ���ȝ�y2A�-���3��=�,��pNM��y�NʅK�n��_�8H��� ��y2��8���qw��	�L�k�/A�y���[����doؓ�j}�C-�&�yRDȯb |��m �p[��#Æ��yr)�"MB�a�^#{�h�s��#�y��A Z�P���d܇&y�!{ C���yB�͖b~0��-'蕃�I�y�H_	f�s����X�2I��0?�T�C��t���&A��2����{��R�GܓR[-�Q��w��1R-�1Uq��ٰ�
�	�� .G�a��$J� ��ı�4A��  �D�����$N���т������h

�H�4%R�c"5��Pm!�d�A����:T��KȚ+S�8a�NV�8�Љ#}Ҫ=�%��蝔1���3�*T�@�p�������'��&�)�IƗ2�qe��M���t*ܞ]��'$�LGy��d�B�y�TA3D�T
n�H�t"'��$ڡ�(O�>͢!�ԀLO�D��o�h�����bӦ������J�%+��,	�e�>sR@���^)lP�*��>�v�O�$�k!��U�2�I%��..���@�k�9��USs������0|��DB5�n���)B�5Ub	y�!�{O&�X�8O �RC�����Op>0�֌]]�� E��Q���C#h����ŪQ�P�)�'R�H�P�耮qP�%���E��4(�����O8�a����d��.h��Tz�DΗ>���2�,�zw슖;O�6�R[G�KE�~֧�S�P����KD"��
SDC�A��`�>��@���0|�$���u����~I���bN�~H����'N����3� Z��Ȏ!#r}�3��+Q����O��'�FO��a�S2Lf�����+:��T�T�C�%�t�OZչL<E�4g�%l;Də7f4��Չ��y��v��S�|�a���$}�"5���H������Ҟe.�OpE�ߴKz�c�b>� �$�KJ���h�pe;b�3?�)qӢ�ʍy��)�<k@�ӱ!�K���@�ƾX��$�������56����d]`Þ�$'�>O,R�xL���y
�'��0���2p.���N��: (��
JS?yQ-w��	��?UH�LY���C��?��W$ N��a���y?�)��?,�!�y?J�X�܀ܑ�*D|!�DI+u.�:�	CJ'��*���!�d0s���c��~�x".ϊ�!��F��@ڴ��[�(�B�g!򄍯|�1����
��@��(��W�!� I�>$�V��|��e(Ua���!�D��9:`q���ɯkm�]2� ��^�!�®9����h 26.Ec��BC�!��R�v����,d�f8#��Y� �!�d��>"�Y� $1&V�C��Ճ5�!򤜯
*X۳��#K����Sn^��!���%B�t+��>�Й��l��g�!��S�7�z�ݝF�P=�U�ѩq�!�D>d���	(Ԅ�*&�499!�d�ti�eKɹu�&���YK+!��[,Q�d�g�2@������<m{!�d	,J����#�`�(�,Uo!��'��ňE�_�qe*�������!�d�:M*��T<	�T<0 � �l�!�$>}�	�C��*g�a`#ň�`�!�d�/&��Yba�5w�j(�)H8!!���-��QX�!Q;)��A1� ad!�$Ö`z���j�3���v�Ʊg_!�D�:l
��U�0Gl����^aN!��u�jʖ�R�cX��P O�Ge!���#"�f�����HF$Mz�����!�$ �AG ���S�:�\���3t�!�� �J�`b�ϯ1�.u�Kߓ�!�R�rW`��6 W�{2P@�ˈ�L�!�6K]�V�z<��K
�!��w:��R�DU�W�\(([Q!��	EG�E���	Cܔ�
�A��!��$:���Aճk����c�"!��8Bք\��T�`&/!Y!�D��2��D�c�ZN�� xU�I%�!�$GiC���&��u#��;�"K�8�!�D	�T+,�` ��d�����x!�&4��p�#�	G�`d��nžl�!� *� 
Q	�(<H�%�՛'�!�Dطt[\\(��(K-�������l�!��9���!�ʎLy���ܡ@!�D�'N�0$�?Ll�A
��_)!��y�� ��?*�y8�ǃ0a!�d�"&�ڦJ��\B���C'}�!�d�5ta�gM`*��(C"�hz!�d�6:�´�ׅى�(|��N>�!�$A�V~�,B�JϗO��	���w�!��3vf�8�A��yvp	P���0c�!�����S1M�)F���B�aW�l!��F:k��(1e�P�4�"4[!�M�pM!�$���IP�F	}�\)Ҁ�C�!��b���i�l�(L�~���g�>�!��#F���I0�	�4Y��2(�"V�!�D��z���eoݡ��Vd�'�!�dE��tJ�b)���!eb2*�!�� Xlu�>B��s��B �i"O�e��BQ�|�h5T�ͅZ�`�"O�:���=/��r�B?P_�-�a"O(��íW�d9d�#5���ib"O�8��Lj��*0������"O���f[	��I�7�TbZ򤺂"O,CT��g
@(�#[="	�"O����cP�o�(���%J$#�� �"Ofu�b�X3V"�`QS*Up���"O���/�8dr�5�U��+� *�"O�t�b�йtPB5�T�+	�mI"O�M��C�d<f�+�4�8X�q"O�L(`,�(f��KN�}�JՃq"O��zb^�o�pP[�*�$P����"OV�۲Nʏ��  �)�Q� ��"Of�rĝ0A�0�r�°�^l�w"O��H�E�xA�i=.R���"O� :�l�6��x�i�1�റu"O�HV+C��00��QE�� 3"O^ah�E�yU8u�'��`?z��0"O� 93��kh&�8�F��)�<ؔ"O�M�WBM�W$2(��/E��蠤"O���%(�e��k�n8��Yٴ"O6]3"֎�N�sH3㔡h�"O�%�sCõ+]��`�(�^� F"O Pbș^έ�`��[Į|Q�"OPzs��k�A(�M�AS�"ON`P.�;8)�f��Y�V��"Ov��S�X�"U,	;��8�t `�"O4���.Ο3|����"�(�"O�{F��ry��+��ȞK��XB�"Ob5g�	�L[��X�6�
�#g"OFpA5��eʤ�g4�����"O ��4'�(j���Xæ�K��a�d"Obu�c�� ����gڶ^�z��*O2YЖ�Ӛ<)�E���+]1ޅ��'������"m>���	K
@�6!�
�'��A��`]q���D��7�% �'߬s�M�֘�(݈;�r� �'H���ƍ��%�E	 b���'�؈b�\'W2	#��� .t=��'A8a�!g<Kb�Di�r�	�'2�@`��v��	`ǝ�#��!#	�'	���6��3[CD�;�L- +�I��bN�Ű�a�a ��άH9XI�"O�����5R����d��֝"O������J�R�Xc_�Y,a9�"O�C���P�J��!I2"�ʄ��"O�-H��
:	�.��f��h>h��r"O8-�u&Y�O�x,0r`�����c"O��zWG"��a �bx���4"OJ���>C��	Z�E7QA^؀�"O$$�3K[P�AF΁	�A01"O��0Q)�M�J��r�R?vSz�Ӡ"OX���P肝���	L5���"O ��&�{��H�F�X)5X��"O ����9.���z�c1PP�i "OF)3u/� J�(@�oR,J0["O��)`*G�����-02�٫"Op��(PL[F0�-:��4(�"O\D@�E�9x%�kl�T츍J�"OJ����6?�$�	(�FX�5"Of��B�W���æ��t�N�"OT�r�]1�|�c�dV�v]�	�"O� .�j2Ȃ"�z�`b�>�՚�"O��#Ӆ��l��U+��!Hx��"O��q���2(���@�>5/����"O��+�������%o[� .��g"O��S�O;lY�8b�=_����"OX���BRv�n$�k�+*(-�"O������8H��e�B낈�L��"OL��EĘ�H=�	�'��e	&�E"O��B��],N�\9h��$h�t@h7"OHՁ��r�܁`�T�A�>�Hc"OXA
�$�=����c(��A� �)�"O2ث#��7/(0ِ�2��z�"Otq�h� *�L�U�@h'�La�"O)X�+���qRN،���q"OpUP�.ҝ9���Ҳ,\�r�(���"O4剂nΏN�~�I6)R��:��"Od����ޭ%����(M:D��,�&"O,L�̝=�������\��K�"O�
#���V!�"���"O�x:Cj��a��낄V�B�� ��"O:�[G��Q@��0*@bX݉�"OLpR��d��8��H-_7̘�4"O�8S� �&�#���r$ftA�"Od�X!	C����A3�ۡ!$:�H"O:@�6@C"�}a6ƞ���"Oވk�/	�GkB ���7w��B�"O�����@�	�x`�T鏟?$q`t"O6���gV~;ɚEc!�LE�"O�,��˺�<m��\�*�L@�"Oބ���R���D1g��<�B�qv"O*if�B�pVx@��cF�4�sB"O����B(�c���|q��"Ol1*�(�m��m(��� ��h�G"O�ٻN!4��[�dG9�� r"O��6eӊ?����)�� ��Xф"O��WGV�(OD���a���aY�"O��jբ9 Z�ʀǋ;�$d�'"OH�(wc�"���FG�O�(�'"O���3�\1a5Rac���SC�Yb"O�e�u荗L΀@S�^%V:�Z"O��P�#��v���c�F2*�H)�"O�-A��ʈT�:��G�t� ��"OB�cb�k@�D��y��+"O���=V��Eȶ坦#;X��S"O��戲�
�	c*tѱm��P�!���1\�`� )���Ye�-~!�Ğ���:V*-+��
��ـD!�ā/������B�f�r����%�!��O�x���a�b�Z�S�^�%�!�$Q19G��(`!��@�~�ɕ�J7�!�d�*B!�\�!M�lP��G�ǃ'!�d :<��Y12N�F��*��}$!�D߭�����(�R@�p&�<`!��!t���gH=q��pѥ�28�!�̙-�	W���
a��K�8�!�6-(��]�T9�!��$˪,�!�D�8,i��)Ӡ�X/⁸R�@�*!�F$���󠪎���0��Ⓓ[!�d��@@G_�O��9�U�f�!��̚s���ذ���5�@��'��!���0~
���V�R#w�,���A=L�!�#a�Ћ�bP�S�X�nU��!���f������F����k�(!s!�ę�d�6�AE�K?-R� E,��5Y!�� �1!FFI-<`Lm��çPϖ��"O�lj��ϊy!�
X<,��0p�"Ol����M�ڐY�J�3�^��4"O���+X�_j� g�Z�Y�<���"O�1y�l!:f���CB@�1�"OhTrB����L��aT�j��@��"Or\rU�ˑGp����N��ز�"OT��pn�J�4�+dDű:@D�R2"O��r��.��ys��!V2@iʐ"O���Q��o��ܡ2"��*����"O4��.)|&&�E1�� "O�(��T�ҸMc�HB�Xa�A"O0���`� Ґ�qЍ�2V�2"O��2   ��   �  F  �  �  �*  �6  fB  M  0U  >\  �b  �h  o  Uu  �{  ہ  2�  ��  I�  ��  ̡  �  Q�  ��  ٺ  �  e�  ��  �  ��  ��  ��  �  �  V O	 � �   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R��I^>�Z�l�)N�HI��S�6�CJ.D�Lh!Nġ ٳ�fݒ!�҉��,��T�I̓L��@|� ]	r"O<��w�R9{&m�7 �)Aj��P䘟�F{��i.[�����N�&�6��Х�}�!��U��0C�/��10.�`��s����<��-�|����G�� 3�iC�ą�IH��?�������O�3: � � D�<�%L���.�����%*4�U����h���� ��#��]C��5'�.��"O�у1mF�1�dIU��'i艂��O>�=E��܆5�>=��ҡtN�pH���y�mX�~�vu�g��G491ŮK��yR"�0A��٧�K�E9(ʡCI��yb��!G��p�$��i�^����P�y�eɯ0�<Y�(LO0P�3��P�y2,ئ ȷ�ɼE.x9u�yB�G�6�vy�*˰Q����	٨�y���TN>aJ�������"�!�y2+�e��[����,�ű�hV&�Py��G3h  i"��yD�RAXv�<AU��{1��s�-�P(�A�t�<�4 �xA�!A���O�hH�V �n�<�6J_�\~������Q�W��t�<1@�]�)p�bI؈k�FE�F+r�<Y�[.i�T�9Q%@+||����.�U�<�1��i4�T-�dym����v�<�`b�� �����*�K�y�<0��7qz��ekM y�p�#�N�K�<��:g�����+J#^��)�a.[F�<���ׁR��!�jI�\H4!x�<Qb�ݟ]z��۠�ۙ	H�P��w�<���f[�%!j�?���cl�<����E��iH�
�(fU��Ti�<	�!]�hRU����, ;�N
J�<��ÿ[�F�:a�#u.�G�D�<Y�l�&w��J"ٝL�H���A�~�<��M��(P�\�*�1&����/ZT�<)�����L
!*5c��q��N�<�S�]9�Xt��+F�yFiSH�<��E��y�t�׆*	Y(L�É�M�<1RB�VrȲ�.]�L,�`��N�<�Iƽ2����C�#�^Q�H�M�<��jr�, ش��uX|<�)�]�<��#,�<��嬌�roܵ�u%�Z�<Y��V�-5�i��Z�Ҳl	BœV�<q��2 �d�k���T���[��O�<	�+��>e#f	ڽ��z�L�<\�"C�|�AE��5�F�n�<Q0�|���`��T�*�����@h�<9�.K$.0�hV �BW�1ؔ�m�<��L�*������Y(i��j�<�A�s�"ء�ɐodA0��d�<� ��*c� m����T��+�I�j�<��m6$�4���6�F(�vȔM�<Ʉ�ɃRԀ��DO�����j�p�<�U�ǣ0����Y\!T�����b�<�6E�)b��m��$��H�#_x�<!�Ə/Y��j��@2`f��2D�v�<�F���PD'�-?��dX�
w�<	���%&TKw�Z2G5�Y���s�<y�Ņ;ra�i���­-,�*Ԍ�E�<� ���vcV*w�Mkf�G�<:eY "OXU�B����4\�ǭ�M 
}��"O�T;UaN�I��q� �R�D�B��r"Ox,BKW��X��
M(����"O�쒅D������!�����"O�YAd%ϥ^ jY;IGJt: K"OlDx�Ҍ[�<�8e�M�@\# "O� ���@*`���I�?UM��8�"O�E+��	7z�y��K�>M�A2"O�ڠ��>t5>l�4FȲY1
dx�"OVT���H�p���#� �I���"O�!�"�~��)[U$����C�"O0���Р0��ϟ
��:E"OF-�c��p\�娥�=R��(��"OH85�N�n"���&�Lk>�A�"OlmP�j��i@�d��*d^�j6"O����(G��@����.R��2�"O�qKeđ,����n4��`�"O8dbElًf��0���N	0�Ā�"O�ubQA�7��}؇˔�_/X]�!"O�쳲��@�D�/)�4�*"-��yR�ùF-,x@@�!7�,������y������1Q*a{��4�y�MS��H����V�~Ё�1�y�i��+<!��\��|q�/P�y҆� V��(�r����ƙ��ѽ�yR��q;���B�܄��͉AѴ�y�珳Y�H�Ҁ-E
�B-xQ�7�yb���p��U��\�9&�{���!�y�O��r�:vj˕ 1"!��j��yr���P��F�F�yA�-�gV �y�#S=V��a[��9r@:��g%�$�y"���!�֔��ϫ6����	�>�y���k���״0����K-�y2	]���`Ɗ]�T�2�A�m��yB��4�4�;�ǊNhy��8�y���>^}��8�[B��ųt���y�l	S��ئ�McꚀ$���yBb���8��۪W�؊t���yBʇ]h<e��K�0@9��+E�W�y��
<��=���C'_�yB�֡3��ȗ6��T�CQ�yBB]�=İ��ܢK�^������y�I*OM�$����H��-P��J��y�4R4P;c��1��}�a�5�y��=������|E}I��V��y¨�X�U06D�iEr-�Q��y�)Й3��|x�K�6g���p�I�9�y�k͗)q���qgU.1�F� ����y���Ȁ�"�R>7*&y��%/�yrCƆ}'`��M�,v������y"�L�jd��C��;!�q��a�<�yrLͯL������BQ0��0'�3�yR��zPY��Ҕ@=z]٠JԀ�y�*�/j*p�+#5�jP�[�y2Ȝ'��Y�.P�(�TI�F��y�aQD"`<*��7LF�̢����y�Et 2�lU�D\�Z���y�'��d�,����]�@9]+ʍ�yrD��~��Ň�:$"�֍���y2"܈e^��Rߍ9j
��Vg�y�/����s��1"pP����yb��;Sr��CA�$Ѷ}�$�ś�yB���1F�.1Ȁ�x�*YI����S�? ��r�/�;.�8m���
��lZ"Oj����e@�9B����X��v"O��ȶ�J�DVb�x���ABx�zP"Oư�e%��2�T�O��J;�dC�"O�ð��%'
�:�A]=#���T�'���ş���ܟ��I��h�Iʟ��	,#6��B��gb�9��n@$�����8��ݟ��Iܟ��I����	؟��	>,D:����8�;�N8>Am���,�I����	ן��	П`����D�	� ���0j��F9
X8Q��	 ���	��Iß���П��	� ���8��,@��Pb�OG�Y�&U��`ƌyf��������۟���ޟ�����h��ߟ0��9��S�e�(���)2MO�+�44�����	ʟd������ퟔ��՟�I-j�J�C��)��p�b%%� ��ߟ<��韔�����	џ���ڟ(�I�d�ڐ�S�I���J@"=ؐ-��Ο��	�0�	ӟ���˟������I�egpa����knA� b�X�N����H��ʟ����I����I؟��I*]��)�T`�Q�U�s�[h�ځ�I����ß ���@������џ��ɦB;�QAέq���JE�@<�Nx�Iן(�I㟀�IƟ`�I�� ��۟P�ɔR�*x�E�8r���j��_80����I���������	����������3,X0�;s�, �0�G�M�{�2x���<���P�I֟�	ß�ߴ�?���"������Y�_(��7��'/�W�jy��'��)�3?aG�ii:�����x��Qi�+2���Q�Ǉ�������?��<���U��X��ڎ3x>�KTe�%�2�Y��?���W��M#�O$����L?� v��5P@���f6���ä*��ҟ�'�>Q�g@�8வ��-m�Xke���M�%�u̓��O�L7=��<#7�f<Ѐ�1J@iٵ
�O���b�ק�O�xC�iW��֯$=�hĔT��\Z 	�<|��$j�LI���=ͧ�?�q�x���*Ō�3����M��<�/O6�OnuoZ�7�c��� �C�p�|�q�7�<���Cl��l�I韜�I�<��O��Y!�N���9U�������	(O�34�5��(N"�U⟔Z%'HjpB��ҜJ�"�X��iy�[���)��<�u�:�pP�'��h�bb���<Qұi����O>�m�R��|:ѪR'B���#�;ym�4�+�<q���?9�N
���ٴ��d}>��'JI���Ti��p�	ӎ�$��Pӄ/���<ͧ�?a���?I���?�wi�\�u#��J����A���Ħ�jp��I���&?��I�GٶPJK����5� �r@!�O8Hn�2�Mk��iQ
#}bDL��E�nˠa�U�~���]I�p��4/�~bc
W@F����'7p`�O���-O�q�pd�?�(8[�-��3���O���O ���O�i�<1V�i� pA�'휤qU�IK4Z�:�O3�X���'�6�$�I���OT6mӦ!�b/T6X,̤��%� rø��PM�_w�9o�f~������3h�O����7��&#��w��ʃuez��T�	ݟ��	ߟ���]��U��Q8��&Rw���ȑK���x��?I��i���D_��T�'��6�:�ĒI���kEK*F=!4cL�i(E��}}2(iӆ\mz>m��
��Y�'�$8�N�
up��EW/
�)�PH�X�.����~�'��Iş��	���I0Pɴ�s����}��a�6P�P�I��'�7,U[*�d�O���|���
svT��h]�N6�P���z~⊰>�¼i��7�\ݟ�~��&:h�����=� I�8i�h��jC%`P�Y2*O�˪�?�gi!���"o�� h���k�
��A�v���O��$�O���i�<QҺi¾5;7��x=ĔУ���@�L�%�+s���'��6�4��-��DV�=�E@A�SN�Q�H�3U����;�M�@�i���h�iw��RWJXq��OK��'�X`���`Y���/C>��ə'����(�	����	П<��I����]�J�{�bH9G�h��h���6m�K�P�d�O��<�	�OH�nz�5H� ���D�v6"�	*E@��M��i����>�|���M�'���P��m5ԉ"���B<��'�z�����8(4�|�Q���󟘫�"X���A�ɛ6��=a�����Id��UyR�b��|���O��D�Ob�0FϼBT,ɘ4-G�Z��i�6��)�����ٺٴV�V�T�qh�#�Np�5� ���aVd/?���1	8ʼ:�lˡ��=����!�?�3�19�*�S4�͸Xb�㱩��?q��?���?i����O8��τ�B[@ԁx禁P ��Or�lZ�>� �����Đߴ���y'�\&0舰��� f�J�P��H��y�Bh�:n��0 � ���q�'�J�r'�H�,Ǌ��	R�L�U:'
�(v�<K'���#��T�ܕ����'��'���'ZHL10	U�
�ԀG��/ Dn��T�h�4>7~1���?��"�'�?)�4n&�Q�!�h���T�����SDV����4<���"t��E�d����j"�[<v8��hf钸A�0o�X3�I�KE<����'�b�%���'�)��!< ��T��I�
�n=���'��'�����S��+�4x�@C��#�d��F�1Z�]IC��+k*Y2�yj����[X}�Jh�,�m�П�#�L[�!�`�3����q��˸tN�5l�o~b�	�,�
e�E%BBܧp�k� ��#O[1����J�1YV�-�R3O����OV���O��d�O��?�6ޢ/�L��j wA���B� ���I�4qZ��̧�?qd�iB�'® �J��4

��Իh!R�� ��O��l���e���_:`>�6�+?Qv틹f�ˊ.�Z����әr���%���Z
���{�Iyy��'C�'���97/����D��F�� ������'h�	��M���қ�?Y���?�/�Jl�P�օ=tZ�q�Ö	 d�Ǖ� ثO yoZ)�M��'x���L��;B@�����
2o�@@e�4��DK�C&*��i>]������v�|��(�ԅ1�,�*T�!��	1(�"�'���'s��4]���4R���s��E+U�L�[1�ݏP�8@�FG�?�?��;śf�'��i>��Ox�mR�d:��k�ą3�Q= j���4K��&o@
Y{���t*u�m��ԦmyRm̀b��9�7`-nb���"��y�_����Ο��������ݟ8�Ob^�;���U�`PӇG;IX4�*@a�`���
�O���OԒ����N���:$�(9!��D�f��!s�CQ"Y�	�4gM��8O�S�']{n�Rݴ�y�(�9�=���WA�w�6�t�|���TAɶq��x�kQ�	vy�O�2��� (���m2ت��Q�B�'�b�'m剠�M��ʂ6�?a��?��J�-}����F�5Zwڼ8Q@���'
�]{�m�b�IC}rl�('@��V��^,���Q���Y�q�*��٫F�1�P� V!y��2��;ڔ�1�b�;ADBŲ�'��p=̉.�M+��?����?�J~����?���h��B!%�7b�x5s�ɓP5*��5u��+L/f,��'��6�-�4��n��R�|i��
,���ӸI�$L֦�h�4-��v ��&֛&��D��-w������1p�-��l����}�����'f��Oyz�4���T�I�\�I:7�Qc!�	Q( ��I�!Rq�=�'a:6�1�
���O��埀��=���I�fB� k�j�.���jl\'���'���i�6��p�OȾ�۳��8�Vl�A;F7<� 5��C�>�iDX���p��\&�q�wyKK�L���ʱ9d���C����'���'��O?剃�Mӗ@��?0�}+Vű��Z�y����+D=�?��i��O��'sd7D�	�ش�6��/HT�9%
�.�X�E˱�M�O���.���r��*�i��s���4�F��J�=P� UC�h��<A���?���?i���?	���'E���B o����GV�dl2�'-�%k�V��<����AʦM%��+�ܫ6���vDF1�~MX�W<�?a+O���e���
+Gw�6�9?�W��83��Q���CE	�2o�.�,c2+�Ol(SN>q*O����Or��Od�O��%s�lw�؜LB>�V���O��vћv�
(�"�'��Z>��Ъ˲^R����4��2Ģ+?q�Q���42��L�O>b?z&_�V�lx�2f�Y��#ܣw<����1O�����JПDі�|2+�*H�!F��4�0$�
�2�'+��'Q���[��3�4$ؤ��@^U�@m �NH@]ޙ�����?I�r�f�$�{}B�aӨ	Zp��j��9�cn	WT*��q���9#ڴ]nv�
�4���D��)��'XT��O�F�,U��ݫ�[���Y*�`�\�'8b�'�r�'���'�哎^��%ô��-m˂A�[J-���ܴT������?����OT>7=�Р���!�2Q�P)�)ւX���ۦ]�ڴMW�Q�b>��ŖڦQ̓`�ұ�BK��+��c��N��<�+� �3H�O�đM>�+Of��O�Ż���x��肤q6�=�ׇ�O���OL��<AҲig��[D�'�B�'y��`�&:�P!ӢL(�����TC}��a�&�m���M;�P����挲c:��d/�	Fҝ(��:?�C)��u��[P����'b���$��?)ţ9Y1���jB�`�ԝCO]�?����?)���?	��I�OTHq@�r��pi 1Mw�*���O�0m�1{|,��ן��4���y��`e����	ۢl2�j�Ʉ��~��'ݛCo�Z-�%k~�z�z⽹%����e�>F�V �KJ�p���H>	-O>��OF���O��d�On�)�œ�l�\a2FJ\Q�2�+dŲ<A��in:3��'�2�'��O��Ƈ�*(藁I�r�D	pw�Ł#@j�LH���t�j��	M�OT��0q���6Q��)����P97l��)�0��Q��C%	\:S�")T��zyB"��{D0@C�m�NdYcȐ	��'��'��Oi���M��C�?Q����6*rC*.ǈ�k�ჾ�?���iD�Ox��'<�7��Ǧ�jߴ?�Q��P�J�1R�9z�ī�ǐ�M��Ot�1���J��=����[q�_Ҏu`�H�oF8ȫ&�F�<Y��?����?y���?A��>|C��U ʄ0���í	%R�'Bjo�J8�&1����֦�&�HC@��1�. �U̕*?�P����?�ODEmZ��M�'L����4�yB�'��yg��f!dKu*]�&C�+v��/p�ĉ�I�T��'��������쟄���oL(��e ��{2*l��ʛ6U���០��P}��j��g/*	��ʟ���$�M�'H�
�+BI�$���b6M_�@]�|�'e˓�?�ݴ#������Oy�fKY�/J`���͒�(1�$D@�l��!��g��Uv��?ISf�'XV�$�RW��,C*�Ȗ�RpE�e����ퟐ��şD�Iߟb>Ŕ'��7��<iVƑ:��!EWn�2��	*']���u��O�����?�Z�t0�4��A�{���X"����yV�i��7m	#t"�6M`��@o��nT�|�'�O����?� ���ũR?xr�#��XY���g�i�2]�' �'`b�'�'e��%���9#@[�n�E��IIOHYb�4?v�l���?����'�?�Q��yg��='K��6���&�:A�a��95&&6m���E8���4�0�iꟜXs��v�,�3���%x9x�r��;Nh�	/1,��w�' ZT$���'�'1�)�`�P]�!a��[,F�Ne�@�'$��'��\����4P�V4"��?��	;
,zPJ�1
(u 2k�9�hͣ��E�>y�i�66M���'�:P�`'öٸ�o�2���c�O�mSS�"Fq@M��8�I�#�?io�O���.O 8�Z��F�*h�m�CG�O��$�O����O��}���d����*!,i) ��[�Z�!�f��A�-B�'��7�&�i�1��+�0FCPQ2�Ŭ�� �V�j�A�4
"��b��+� o�Z�\�eA�m�JEA�$��	��P�4KʡH$u��IX������O|�D�O|���O���R:�����Ȍ�(�z�j1:Vl����Ζ<�'�r��$�'_ܹ�7�
�TTb1dE$H�� ��>���i�\6��韐G�d��s��4�#�I�?�q�P�^�	n��gϴG��I�z�"A��'��&��'@F�C��6XҰA�s�5|�pU���'�r�'�����4\����49�lq#�~�t�#G���	�uX\���-y����\y��']��/`ӄiy��^� ��`vmB�?'�7M"?����u^��	�;��'`[k�e3~�{�`�`�8�����^���O��$�O����O"��<���쓔@NDUisfI�
�I���I�M�%H�|�����6�|��]�H��`�\4��t9u
����İ>�Q�iG� �'g5��4��$ԻD��p�'0D�X��U�b�$TD`N��?�$�(�$�<)���?����?��䘊F�ތ���i�L-Z���<�?������ަYBjE�P����0�O](8#���<nv�	(��*��D!�O���'Q�6�Ħe;���O	�[�+'mv�p�M�#X�s��$,��Be�	Y��i>��`�'9da'�P���#�(21�ԕM�D4 �mGٟ��	��	ʟb>��'�7��?j��8��3j���h�U;�����O��DKϦe�?�cS����4|:.)�����8���A')uPM��i�7�P�=�7-,?��,��iB'��d^y�T�� H��W`
Gc��r���<���?����?���?i,�F՛��ܶI�12%F�%3j��$�����X^���	Ο�&?��	��M�;N�f�͙�&��p� �p�t��e�i��7mAɟ ԧ�O�~��iC�^5)�!	���o%r����H9U�D�~ڤ���B�O�˓�?���L�8:���Ϯ4�� ^I�,!����?a���?�-O�,m5`4��I����kTu9&τyr��`5l-a�F��?ɔ\��ܴy�����O��a��9�1��G5�CEХSd���'�j� �(�P������4���|�$�'�a����qr�9���S�Y��'���'���'��>��	e�BT�Rƚ=8�ʽB��#r�D��%�Mf��?y����6�4�P8���Q�uL��m�>����A�O`��jӂ�l�\��Tl�]~�rFv��s�y�*BW|:d�1�\4i�X�Su��	����d�O ���O����O�dnQҵb�_^\�EO�}�V��PU�d@شu����?1����Ou�آ�n�004�)�U�-��ڀ%�>���i5�7���@E�D�G�W}6ԁ֊B�0�\��U�7��R0d���I?H��J��'uX�&��'�B�Qb@&2���@B N�{�l����',��'+�����P���ڴf&����vԄG�Tw ��dЂ8M@�s�`����A}"�h�"%m��MCa�̝�l}����.�Э��I4gD��Aٴ��Dъ	� �J�'T���Tܮ1)ASt��-  ��2N��u̓�?���?a��?�����O���[��Q͞�fc@b������'N�'|H6�]���O�m\�1�dT�A*j>bx(esv����������|j�X�Mk�O���H q�0�T��;ȑ �o���`��GeғO���?����?��?(^q ��E�u�P�s)M�&D�����?I.O�m�:T�����R�N'QZ��'�^�pM�X�ɲ����y��'v��E�O�c?���'D�� ��&+ǵn���`�N F�"��n��m��������*f�|d	�6:�eR�a�?M���qb��\Tb�'	b�'z���\�`۴N���2��b�����I�T�`�D�?!�-T�V���W}��w�4E�.	�n�(X���9R�X7I֦1��5�oZ~~S�O(.-Q�	�V����D�̑����aB2�/�:.��<����?����?���?�)�ح"�Js��p�FBYk>�y�pI㦉�F)ӟ,�������W��y�_�X��Hȕc��6J.)��T.�7�զ�����	��6�j� ��n͔AD�Cw�[-qIDePf�}�x$��2u�r�FF�ry�O#�{�����ǡ+���%� t���'���'5�&�MS�ϐ��?���?a%�4d: SQ�G_�~j#���'@R�``��,x�b�oZ��D�4F��9P`�Vh�<ZP.O6��	�#�D"a�T�r2l'?�B!�'l2l�	<o�p(A�K���4GF��GT�l��Ο8������u�O�R��*<=H��FL�BJR5B��I(8�g`Ӡ)	Q��O���ߦ��?ͻuO�A( �1�Q�1�G1p�n�̓A��6�b�z n�5hT�nZ^~RИc���S� �Pxr`	��ܬ�A�çA�X��#���<����?I��?Y��?a����7Ht1� �3`���EP��� ˦x���ퟠ��Ɵ�¢�M,M��q����A�:�����M㴼i�D�8ҧ8\>`��.($,dċ��n��h!D�I��q�-O������?���?���<9�M�9�ఔC�-F��QF�?����?���?ͧ��¦I������l@vE;${0�(V�^�֤����Ɵ0�4��'��H����v�0,oZ�
��P�O�G�DA�q��f<��`ئ�'6D��� �?����tD`�1��@.cU�=��,�0�n���p���I؟���矬��埠��aA�6\��Rv��c�a���}���?9�*D�V�U#����'�7�*��կL=�<�D��8t6<� �X#W�^���Cy��'���O�>�*��i��I�_�~#� ./�����dOY��]���` R��N�{y��'~�'��bV�Ҝ)���7���WVR�'�剁�M���O��?a���?Q*����*@��2#%\�A9И���O�m���M��'���v�P�H�56*-UE� ���ZsaV�ؤ��ۢ^����|2���OF��M>�&�Ԥ����S&/���2�듾�?q��?I���?�|Z+O.n�|��%JT�\j|����7_��K��x�ɯ�M��"I�>!��iĝ���?8( ЭQ��iJ��|�2Pl���rӖ���� ���ݘ*O<��Ш@�_����go��> ű�8O��?	���?���?������)f92�z�昽6P��� Q�q�nZTL��	��IA���r�����a��Z�q`B�Gx�T�জ=�L���I^}���N^��:O\-3F��*i�z�r�B�]����>O
�rD����?)���O^˓���Or��P�e��	�į�t�Z��v)P�`�Z�d�O��D�O\˓Z���R�n���'�g{Qr-���/s�ԉ� _�N|�'�bm�>���in*6���]��O�-I�#՝&}$c�l�":�d�×�d
�ʙ�&:(���n�S� .r�����+�+PU�A��j\BónO���� �	��8G�$�'���Ï�E�9�׎��F��<@��'p�6��6�����O�Eo^�ӼC�N&BSB����Lp�h�A���<!e�i�^6M\ꦙ�s�O����'�R�����?��܉#�\	WeQ�k;������]�'9�	ן��IߟT�I̟��ɨR���rD拻�;���o��=�'�X6��5lǘ��Of��<�i�O,i����3���06�Ҕ5���)�lWT}ed�jYmږ�?����<�|�/ȸ{����`;w��Qȱ��n ʓ=�d9���O� J>�.O~T��m_� Q�i	��O��XH�L�O��d�O��d�O�ɺ<�`�iK2(Z��'��tj�+�[��yBi��tOnxS��'��6�+�ɬ����립��4O}�F���1�.P��x� �C���0Rq�iZ�	��0���OaL�&?��[c�~q+��,;֑x�k��z�֨)�'hR�'���'�b�'��%�ENݏ@T���eR�X���<9��+�*�.����'�7'���GT�3a/H���!���T^p�I~}BbhӪ<nz>IYp��Ц��'%>H{`��(���o�C�p0��Ǆ�3��y�I�x��'��	쟰��ԟ��ɾh��Ae����hR��ðK]nL�	ҟ��'�`7mC�d���$�O.�$�|Ba���4����: ����t~m�>�Խi��6������~�F,ae.�1���6��ԠB�En�ɂ�h;.��+O�Iâ�?�sl&���� �s��; �<)ĉ0�����O@�d�O��I�<�1�i����f��~�P!��C����&#K"@mr�'��6�3�	4��D^צ��b�!�Lp blU�e��<�B��M��i�Ҝx��i���� �H� ��O���'���[�SXi��$+�!�'��	��h�	�0��Ο���@�Tဟ���E�̢8�H�Ra�GS@6���@�D�OV��#�i�O�mz�=Xen�j���*W�����2Ѓ�?��4Z�BR���д��"���	/*�ة�q��*�R@�*�扈+XU��'+ P�IoyB]�T�����Ćȡ7O�z��:-��u�S#�՟���� ��ly�i��5��A�Oj���OpU��(�&Z�@Y*.~���5��3��$G禽��4���l�>Q�.Nb}�0i WpBⶪf~Ra�Ӣ��h�42��O��@�I32�RB~a�0A�o�{�ఄ�\�(	��'�"�'���Sȟ���8P�+�㐖>^ժ��:�4\�����?AG�i��O�m��Q�fo�-l��J��I40*�Ħy�4*��������f��p�UI��jn�DLQ�]�:�z�Ȼ1�� ��	�Am�&���'�2�'�R�'�B�'=&�:X�F[�,�t�(��RAG����Šu'�ԟ\�I��0&?Q���F=p� �O��)	J� �����(l3�O|Ym��M���'��>B��B)"ka��#Q�CT���"��#R'Uyb�o�V\�ɚ8�'�剢+��\r�哪ZQ����V
�ڑ�	����� �i>�'A�6���U��$U�Z+h�r�.�Rq�x ��t�T��R�Q�?�%[���ش^���nӢ����:L�٣�E\W��$��hςe�6�<?1��Q�|����P���i�k���[srebPK� [4���鎋aQ��O��d�O����O.�d?�S3� s&҇�Ɯ�blSa�j$�	ɟH��(�M��,M�$Cb�B�Ob!�J2��VBA&]{��hAa�� �'�87mΦ�#:���nZv~���� ��( �Mu���*r�e���\;���`ܓ���'/��Pʘ�?�dH�#!B�k���B5�}A��h�<����79`�W�1F\��>),1Q#@��2vf�q�$T��t2�#ԒbIB1��!Ө�KPB�!P��G��)0��
X�.��SJ_H�7��YIT `�k��x�Fb�{�"�qU�l����AsέP��9smVLkUFL�~]�q�:p��$B�b��o,@Y�"�/%��T�dDܴD�6��OT���O|�IO������ߴ'��a�@ě@N�	'����ȟ�(�
ԟ�'����sQ! �JȻ/�ȅa�iP�4�U�ش���_�`�x�mZ��i�O��HZ~�.H����! G�68r����ġ�Mc��?�/?�?	L>q��Tf��<�rtS��=?�p2�
�#�MӠfHa��'���'z��F,�Ɇ<2F�ф-�@f^	��ݔeR<(�4l}0Ő)O��D�OΒ�����O�h�@ɟ��й����~Ǟ`0��䦁�������;C㚀����O�Ӈ
�JHɡg���N���MP�S�yR�ͲQ������O���^	u$&Ac����is��qO�_��`�'U>���'�U���	�$h����ѢǞS��@ZVo�up���O��q���	˟��	ܟ��	ٟt��dвc�Aʇ�»
$b����W�Ce�I䟬���P�Ir��T��YV]����a0l�cb9�\�����Q2��?����?	��?��ы�?Is �q��c�g>:�=؆k��s[���'R�'��'B�'�,z���!�M+��.T�>�PA�̹d�j��w}b�'sB�'|�ɍb-�0"O|2�+�O����36�������ݛ��'�' ��'X̙��}R��	ш��c�^�����!�M���?���?��
����O������c�v����n�%�6��3���&�����0���1<��c��F,j!��q0���'n�nZß����8�r���Ɵ �'����'Zc.���<Z-@`e��+J���ܴ�?���������M�S�*���C��2�`@�cP��6 n�(vD�	ǟ�'��4�'"X�$ねL�h�|��4�"]r�q��^��MsBڴDg�l�<E��'����#�	�B��ű#�Q%M�Jy���'<��'3��'(��c���	m?qtJ�:�3�(��B�y����p}��'<R��%#H��ǟ���Ο��{�nAh0H�Ũ<)������n�Yy"E�|�)�[�a��N�D�p�h�F�.�"Lj�Y�x�pM���$��?a��?�*O8�cKN�S��Tg��prx�6% �4y'���I�d&��'7n��S'�"`�`X*��b�E�ͱ��'��E������ݺ<?���#�8½�d@��y�)��U}Zh�e@�J��C�$��'9ީyƠL����⊬����2e��m!!�n]-n|�WaH�M$\���E'�Vl���R$q	�d�������ò��Bҵ��gE�%5Լb�J9&����_>*��Ȓ��e)��)7d<0�S��)�@P���Ԝ��r$ϭ�"@��.��EAN5p��
� �2��z;��;4 �k�d|���ĜS�������?1v.Jkc�LI���=FTA:��Z���i�Df�@q��R �$#��"��V%��Ɍx4ĝ�F�^�Zy 0�R.����S@҈F娅�Oހ��暧7�"��.1`LJ�X b�O"�lZ�H�6�)���X�iG1A(����Vl*�B�	�r��c�χ+�FxcE+UJd����g�'��xsR [���b�o�-��rej���O����?���I��O��D�O���WԺ�FfǜorT9� ���bfHY �	]6�E��>��3�h���L>��J�(���QjQ&�t�A3K��p�a�/�&�9�J�ȴ�}r##�Ty�f-��Ȑ�v�0�Pe�+�x%�	{~Z`L��S����	���cA��7-�jJ�(��i�ȸ��~h<�q��-T��h����,&n�Q҆�a~҈4ғ��	�<�ń �m�vѫhh�t-y��E��dT�	��?���?��h����O ��p>}�.S�c�mR��r�*}�"���<R����?U��l�>|R���w�I�m���,�zȆ(���^�iE��)P�X��&����æa�6�D,w��b��T#���K>q���(�Y1����]I�F�B���#�M�Q�iTBV�D��F��[�$���)�����cH ��U��U�B�ؗa<A����B��K���<�#M���$���N|*G�>u����\)/2�|3��O�<	f&05��d+�(N�GLār$��K�<�I�2�8$@	�X[�u�Bc�~�<9�-������.π`�Pف' R}�<��F�>���Z��˔<͒�)�kB�<a�%�NJ�I'MD�ka��C��|�<�5oثrĸ]����(�8(jU�|�<���U�3b��� Ȍ��pLB7l�u�<i�$��M��&Ԅ��T�%�y�d�	h}L�J�΀,2�r��W;�yB��)z�R|�1�2Ft|��0N��y�B�X%v�����J`^U����y
� ��Y_�gt����T,��}r'"O�L�òA'00ZA&ؔ0��}"Ov�����f!�Ef�(8�%�"O:89&@�`��=Hv���7� �V"Opr�a�j;8����ۏ$��"O@D�@+�P�t�0��~b� b"OT��dN9Y�	{u�1��"O�q���8�H3@ڍ3�^qq"O,��āB�aXX����ȞHN�"O,`h��*����#��)��"OJx��;%Ŭ����8N�x�"Op�#��ըB�Z�B���	k>��f"O���Nk��8rp�\��
u�"OB�2/�
�XSAҍXK5H"OL z0"A�&(A���:K�0"Om�`̈�D
2q��@ۨSH���"O�=0o��:���SVo=���t"O�� �+qެ�G��)B�S�"O��"��:�~��Q�Jlȣ"O�������g̈́�z��"Oh�P���<�X鳔V�e��"O��1��e��  KA��zI[�"O�񺰋�<���I� � gܞp��"OVh
���d�I�@n�	:ܤPq "O�8ڃ,Ĝh2�m�����k���"Oj�B7��3�n��6�1|^m��"O$ ��U�\M��R`�f�4��"O�SeD��	��D+t�X�t�1"O��@��^�(t��@^��"O��R�18' ���dK�WI,��Q"O<���Q+�d�Be�HdfAyf"O����&�D���cR'pVXHf"O\$
��XR���dF�h�p�r"OL��!Ȑ4�ĩE&�zaF��"O�,�U57@&�"2�R�)�LM��O��2�$�Oԍk�%M�4zɻ`��q��L�7�'�ƨ07����	$v��c��-N��P"�?D����Z#SĒ����+{�%"�+�^q���)+�ar n�t�	�a�U�Rg�C�	�~[*�b��	t���J��Ҵy��0鳭B	v�1Oģ}�4��	2Fl0Z6�q¢I;
zZ5��)��Y���d�fi�s�A:��)K<ў't��W.U5v�Xڄ��L�|�J��1e�'"������<�,U���b�����|I,��ԋL�XpG ��v�Y�7F
C��Pː��!7��I�d���=�����/j�đ�h�;C��×�4r��'����2G����		ָ1H����Wnp�i�� k}�%V%��DB䉔�ʴ1#���	��LK"/�I���\;Q��h�xN�%�'�Z��O|�`�Q�A���/0NHP�Cѭ{ vĻ�N?D�X 7��8rz�X3�@ X���kD�%�?�!�_����A����4
�����j�P�M�sɎGY�ѱ�+�o�
8��Iz�p�C�%M!'>��+��+2�!���8MdV��5��:`?-��.C9B�̌�Bj�^���h�#��t����tb刐 7�	��"%����t���a`�?�7-_�dy�5�_&A~�h��ʟ5<���钑�!��<���ę .�����F&�\��1O+L��*\n��Uc2��%�0Q���yW+kpP�[Ӫ�WD�( L��y��8;�����MN��81����l��ADR?^-^���#�3�<�+^w`��҃O�w�qO�8�Q���`D��(� B=JTh
��'�A�Ca�*vXsV�@0Z͔�z���
o,X�{5�eK`��D��G�ب���݈7��zR��l(�A������G�ֻ��'>�Ъ��O90�hJ�D������:/~��'۞z�=�t-Ŧo��yx�%<}�C剹|��bI7�JY�`�U3OI����g�v�r7���j�4����=��aM~�<���z',U#m\���
kPR��'��@K�c
�:?�1j�G_9 5��U�����@.��	p�a�r3l�S����
�1b�0�8"1�>�I��-q�P�VY��� Ԉ�<	F�X�M��,s�	;~V[������ �0��H<,\9TL,7������)���q�ʅ� E��q�.�8��O�G�<��`�Uu�=l�4����K�gp� ����G�I�3�I�䁀�@W�t��}�iɾ@�2�"O� H��݃t�"ق�͆��\$��/�$<�6�F��O�a�%# W���ͻb�(A�fmǓj��5b֧j�jl���0�f|���ֆ"H(@0�L�=`����'bN.}X��G[�	�<���ïv���"���>@b���q��W �l�%靲#Y^���7��+RW �`��޵u. ��`C�%ǲ�?��%cC�J��+�`�},B��co4D��B'���@V^ ���ʢ�&"��4��	`�"l	�-xtf� �����C%F�-^�b�zFE2UȨk@��r�<�V�H;z{"Ay�c�3-�~Њ���4(��	�W�68�����M�S:�"�<�,,h$�ϙ72��%( ��R��ô$Q!=��
�R�<q8����%���(��Cm�f��/�{�\��	�*eh@4h{�ʠ��"؆ȓ ���[_-����A,P`��ȓ�@+Qa��w	Z��t��?^Pq��w�&ؒdE^����[��6$��	�h���*=J� KN�"0��ȓS5N$'ϙ9|�8�6�@/`M$!�ȓ0UF���ŎH��@�/w\�@�ȓ�����Ûpil���U>U���ȓ.���{0��<���i��<	L ���h#s�ƺ6���©��{��ȓ\d:8 ��˥hc��!Ū�	ܩ��{���xӁ�+BvD`"���Ze��ȓC�\�K�e(PtǁE|���mUԙb�E�Q����Df�+rjՄȓx5�Y8!���/r���*�
8ھ݅�vA��Dg\�e}�M�P��xd����	`d���dڲ[�F�Zr�74x��{�|e�gg۴��yr��ع3�깅ȓk0*�K��]�>�:Ub�a��q�ȓ �-� ���c���6�Ӊ"�����T����<BGRi�&��+�l���k�|��	�%}��J������C|VL�G��	^���q��əE,<������7�Ƈy)�� k؞��-��-������N��܁Q (��)��s����S�DliQ�Q�gaɆȓ4�2�![d��@WL��j��@�ȓD< �S%6%�p���//����ȓ#|PWʆ�|U<���S.|�Q�ȓz\M��m�*-��P� �F,�J��ȓy� �'둑B�e�w)
)t7Щ�ȓ��Qփ2/�n#u�D�/���� �&����Y�'V>�B [� ���ȓO�����HE Hi����P�ڰ�ȓ7���qN��VN�I{�iH*p����U���&��D�(ň��G:�0�ȓV���2,�:�^����\$1K֭�ȓU�[ê�N�قI�$�� �ȓ��˵	EgB���ˡ6�9�ȓzL4Ng{2���$^!�t���P��rF�&vb\���kѪ��ȓFpZ1����*ܮ��򬜴!x~�ȓz��	�`̎X�q�0�D�A��S�|����ͥ"2%rW�̌t�걅ȓ�n��p��3H!e��	�����9�$���J��o�xء�H�>9C�͆�`r��'�M�R4�4��7\��͆�D��PPG��c� #E��)vU�ȓF���R4�Y�V,
�YF$)��
\�0aiI�H�(A���T�̅ȓZ����Q�h�RE�ʑL^�A��S�? ����MR6��j`�9B^�"O|͸mRyW�YHEIV��r%"O�@��NZ�DRh�!��'@,|Ԩ"Oƌɷd[{�j)���F�T��%"O���茬F��E!�L�HU{"O��˴c�s$���B����xh�"Oj�b�G�0��M�U��G�A['"O��ٲ��ej�I��!S�άd"O�������ʃgݎj�\�ɥ"O ��Ao[�hh}�f�/� P��"O���rD��S��s�#H�#�fc�"O��+6-�>X ��@M�8=F2��Q"O���[���JD̊M�J��$"O8���-З߰1�
&@���V"O�#�\~��R��/l���A�"OJQJ����f	D1'(�G}��!"O|E�2����JxSǦ�rn�ٕ"O�\��B9�d��M��hc"O�KQ��59��0ze�Ֆ!4i��"O��`f��=�踨f�M�a%"O�Tk�l��X8����[�]J�K"O�P���K�o�2%P��XR,�%"O�L��O�R��m�JǇ:W. �"O���Aʶ,ʬ�hjOtdhQH�"O4x�u&
�=���yԨ��n\u�"OpX���#�*�Ӷ���n��X 6"O\5)p��#G���p����qe"O�	�a	kQ8�)G�H-~�y��"O�#�
2S�"�r�(P�R�"O����A�/:+ʈ!�^$!�\Ah"O�ٹ�gǸ',��ñ�ѣw��AH"Oh�*h�q��P��(t�@"O �ơ�D��t��kB 	�~�('"Olhy��6:`J�HU�J�t�"k�"OP1a��c�t�Rj!��"O``�&g�{\Հu��C�b�"Oy@䂥u�쁨f�_U�t��"O�M�-���*�p�GV$CF��"O�:2�%��PP�_�i&
]�"O �0��\'R���
_">hh�U"O�qS��Q�(�Wi��L(�"O������s)t$xPHW�_��I��"O�|���(_��d���S삜��"O��sV$O�}ƒ��"�&|� ��"O�h��
��zd마v�r��""O����i^�f��L��A��X�"O�����D[6Nс=��={#"O��D���8K���������Ye"O��{Z�K�.��.B.	�c"O>����G��葶��$>H�"Od$C�IEq����!�6$����"O��k���h⬄�fKV�R��3"O���PK�8 ޥA�
떵�"O�`�I�Lh`5��R���+�"OP��7@�)�dEK��Ė�l��"O��B+�-2�l�a/R�6�8p"O0aկK�����B�<�T�G"ORl��Ҁd�
�͘$j��EXu"O�H@��,my�@��NRSF�8 �"O��ce� �,��D.�j��HU"OHE���\9���kY)y���U"O	��&��a��!X��FN�X�*�"O�t����7�`,�h�C�:g�!�$Ԗ3�̒`��;Q7�偒i'�!�� ��رE��\�3��7{Pu��"Op+W��uI�u��%��$U&$"T"O�p��k���z�E�$C88T:�"O<�c�) �p@���O<�M�T"O�:�
W;j��FD3j�@��"O���«�#X��"�c�#h�(a�"O�]s�Q.B:t�ѡb�Gߞ�JA"OP�jG'�;)]�H0 "]�K����!"O�`PeB_�C٘51��_�x(x@"O��jGAZO�>�S&\�H��"O�1i�
��� P%޹	)��b�"O�]a��X%(��|a��I�8Jp�"O܈j�É�4MK�>KL�e��y�\�"7�m��ΏI���uh���y��"ꈒ�"°�f1�䄗)�yi0����
Y�x"�mD	�y�%ˁ2Q�l
4F��Y޲��S�Q/�y�ہh�N�+t/YQFnqV���yr���9�,7JLKm�L�5eI��y��S�]�Xe0� �2�~-Y4mJ��y��̗G(����H��%�ӫε�y�mG-)� Q��t�
d�c�ŭ�yB�-l�\e!��pG�x2�ⓝ�y�"v%@`wǗ�9X��;⍈��y2dR�$������+���;T@�y��L�\��� ��q�{f�Y��yB*K�n�6�r�����!�ܘ�yrH��|������ԛ&��p2`��y�Fl�䬸�d�~\|�sF����y2CH�$�@ju�ɳ@!�8�թ��yb'�o�Le�+��2��UFP�y������Eлz�Z�G@K5�yb���7�=Ӷ��q�
 ��B��yb��i58 f� :>H�%)��y���J����]�,xN鉵���yR�#hv�x��� 3������M�yBG!�.�J�$(��=��ۉ�y��M����+�)V6��� ���y҄8v�4��`�T�X<s5��y���u��!i�}
D͛�cD>�ybZ�V�KBIzl�*C��y"��
T^��PCa��	�ԔY�f�	�y��WXfL�
�����k���y��&:]�d %�9y�x��4BȔ�yEϢZ�zĀ�u���˱�э�yR��7��������,� M#�yB�X kx�8�%�\?v�6���I��y�j�9<.�Kf�­?��űe�˘�y�EX>��ڒfʿ��䱳���y"��N 22���
�����W�yR��
���Aj�64 I�)���y2�R�QY^�[�̑G`�RT���yB��&�u����=f��4�c�K��yr
Ӷ�4qva��YH"�1@����y��ȃ|�uكf�z��[@�Ӹ�y���+;*�ၣ�?	�`Iٗh��y����Ab�������|�,� �C%�y�G���yq�EJ|���1w���y��[2>D��P��&l6�G(�y�`˭X���4	ıS�fl�v戛�~��)ڧnU��[�LߦUj0���կ�8P�ȓ�搃F�N�k�L�
�)Ozy��iІI ����h���%�TY��me��Ӣ�?�f�#��D�mu|���S�? ��yTA�+C��H�L�C���zיx�.�D���O?�Tq�(" ���puk�2Oj�͘�'|~�;4l�av��	ÑF|��a�'���zsϒ�-#�$�@m��E��TB�'���,�,��( 픥I>*X��'�콱wƋ�LX��-<X^���'pd�B�s��0)�@S�~$B��'��l� 3x3:�
�R�x�pZ�'���@AԀ
��]��@�
G�q�
�'f�pC�;j�V�e�͡C��uk�'Į��Vo��]d��Iը6��1r�'�!cg����L!̩2�p�9�'.i�nA�B���K(tyԩ�'#��s%�/jqԴ��aA�����'��9ҩS7P���P�R�xY�	�'5� h�A��#y��&�ׅ.����'a@����*�~�x��/}n�U��'d��Z�@���]�?���k�'�X,Y�E h`Z',Ėf+<�'g�l�c"ڧQ\���A�,�f�+�'؄,�rLՠ,�lz��
{C�d{�'�B̪w
O�I=:��#�ĩcqŸ�'���y,P$<"E�SmĪn���'0~A7%��ze|tɢ@�Q��'U�{��=tK���QbI�"A+�'���Ae��P�X�y�n
	H��'W��(��ϚB�� �%G�3]:I��'0���!�a2 i��^�(~P��'��x!EϯY��\@���.Nt�
�'��T�Aӳ=��4�Q��Q�ث
�'ZB<�U�$bྉ�	Br���'����-N�'�F�h@韾P~B�B
�'�Rm��E\�H�h�P�a��I$��r	�'�$�`���n�tK����d�	�'� z#AI�Ma��I��B6$��E��'F�$���^<Y\���̽+|���'ִa��+p�](��I�!��R�'�A�5�*3�=s�Wy� B�'?d1j�<��=I��K���'QD��+",��ű�+I)jچ���'	2H�o�m���!U9\�m��'@�s��:�}��e@�K�'�ԼBB�W�Z9��~��1)�'U�8Y��%�ɜ	x2���'-����ٳ*�Ő�c��Z!�'�\�R	ۙG�Nq(%���jx!�'��ڋ8'&�3�f  D�	�'L읭(U�ְ �K�&� ̫�6D�z�� j@X��(��!73D��a�ń:>N��C�/�6H��a�1E2D�,�Ec�V���.�>��|�%�3D��	!�ye�S�ܸf0Hz�a1D��y��ߘ:�Y0�BN�$p@��<D�4����
T�@��T�+Aʹ�R�'D�y��JT��)�O-q��-i� 1D��Q`,�4��1A"����0D�0��Ɛ���E�v̵1�k.D�pa�XÖc&�*����-D������Y6�lڔmϊZN��A?D�� �eX�Z�D��cLVjIC�=D�|��)�*B��P�Yx���?D�0ir1��=Q��"�p�C�#D��s�aH�tY�1d��4V,���<D� 5�
�CHv�CA+B�F�Ց��'D�� ���2@
j�dTR3���xqp�)�"O��P�'
lƢ�S���h�"�"O� ��"aiQrB 0#;���"O�!+A�Q���Q��S�c"D��&"OJY#�Ƈ1I���O»U��R�"O���+V6**��2�$ab"OdܫPh��h>t��d��E��h�"O�4r��S�����I��T���"OQi2ȉ�n2�	Ua�j�t<�"O��s�L͙j"�Ep��ˠ:���`@"O^���K�@�P�@�M���U"O�������y�j���M�y�� �"OLu��n�;�4���
�ra��T"O����R6k��PBgJ�wx��� "O��g.[�{���c@�ur�`�"O�xj�0�Z���3P�9�"O���dK����j�/O��"O}A��/5�p {� ���4�;u"O�3��1k��@�-K~�u�s"O<�yN�x�77��EZe��c8!��Zo߾Ĳ �M,( h4-�1
!��Y8}T��G��m�@��,
C�!�$Y�|�x�jT&Xy�����!�dZ�\��i1��O�-,��ˊR�!��˜n"M��ѼY>��fh��e^!��&8ZW�ɝG�H�Q��TS!�ă�?1Xc3�C�4�&�B��S�.J!��D"��M[��I�ld�fB/
=!�Đ�%ļY��jLq@G�!��z��M�B��h�>\{�ċ�Qd!�䑡^�@�@� ��P�a�!��r
�c"Y�;���x��M� �!�]�k�H,dI#�n83��?G�!�DD�t����+d�dM[P�V�ny!�UC���k�5fܢ��({^!򤒶"�~�$EWyxl�y��;%6!�D�7F�p�ۢ*3�<����_q/!��4zu�x�&�U�u�ܐ`�煶p�!�dUj�Nա�i�4Uܬ%�Sg��?�!�$�-F�� � Ή���RťS�-�!�$!��q���J;f���S��r�'V�����y�2���Gŀg��C�'�xAA�ňKI���©�<[#�T;�'�T��!��bHJ�Rg�\�XJ
�'
r�@��ԬX�b,b�!S4Ym�lr	�'��@	�T��CG
U�tl��'�6,I� �1buI$h�2_=�p�'�@I
���)Ed�QaT�B"�N�1�'�6�g��;?��[�oF	�jm��'�8�����8�\�1ő�φ��'ި��`f �K���+R�H,��'*�{נO��f��P����k�'�&��p��6ļt#�e�w� �j�'�l�37�FD��0w��F��%@	�'�l���"1VͰ�����6E��#	�'޶}�MkS�L��e�9r 2�'���C�T$NN�Bɑ�.V�z�'���H.AN���C�Z~)�'��T���W�t�T���G^R��e��'V���Cl�^�nh�#�s": ��' ����v��*����h����'P�푥l5!i�|���T�M�8D��'��-)�EY#$����A�xx"T�
�' :Y�'Ԟx����
kk
Ph
��� - abZL�%��c�=2���c"Ot`1�dư	'�͗)Y/��Ȇ"Oj��&��+Tɫ�k�WD\Q��"Ok ��"ř�ʁ
4b-�5"O&̘�FH� ����C�TX�b"O�9��n 8PX8I�"#'�p  "O�y9!NB���ć��5���H�"O���띊E���zw��<8^��s"ON�"ĆP�"��#��!B/X��"OBl3oܔ%�dⶁ�e����%"O�]��I�&��I���~4��"Op�����&P�6U�WA�x��,;�"Oཱི�A!F��qcM^��Ve��"O��b��Z{��˽&��k'"O� s����R��S �
1�$"O���5�A�Q`����Ò"F��Pj"O���].T�XM�BH������"OP���h5�ٓ2-�%w(�k7"O��q�aC�Vd@\@�!u}�
Յ�@�<D+7�<��!�� 4h�"�O�~�<a�ÄZ�� ң�&�B��!K�}�<q�553�q%�<E3,�s˒e�<!��ϊw��W��R A����G�<)šW4O��mؕ˔ u���2�OB�<у��E�ZM� o!��s͂d�<�ѩQ{؆��DX"$� �c�<ЕIt����0fб�%�^�<��匝+4�g��h��}c�&�q�<�v.���<5'�
?��9�Kx�<��"xP�3"$�L��F��z�<��/p_ԙB��zơQW��v�<��j�J���Q�lԞp�&�D�[h�<	b��c\>q�h�6��{%�|�<1a�W�,".y��Ά����t�y�<�פ�.x r�I�L��!�VP�<1��+Q��"�
4��У6EYJ�<�dG5_Lx\3�#�G�i#��Qb�<�'P�=d�SC`�g(����c�<�W� 8�i�;2��T ��a�<�t ��$`x 	<"��!�g�<�׌�"~@b]4��:)�x�i�!Ba�<���,nR�1���(��!2W�M^�<I��=!�9��Js�� jE�VP�<�1aK�Nc��q�X�E�ܨ�#.O�<���Օ)A���N��9�LK�<��hO�yr�dmێ#*�ق��q�<�0&�!_��X��0z��x�̕y�<I-��{aѣU�,<�5P���r�<	'@��x��ţۦ�:�C"\m�<�bј(��
�&Z�<'r@�1hm�<A6d+�=�a��<]�!P�ă@�<�fL��N���f�8H p�lh�<���"@<4�S��57��<yU)�]�<I�a��\L];EŖ-2�H\k��D�<aRm�3 ��R��+Gd��R�%A�<�t�1l�j"�F+Tm���F'�@�<	�lL
?��u�VJ_'Xp��𶣞{�<�W��1
��R�_V�$$������:\� ����&�H !�+�Xg�l�ȓ/8F=�Ae_4����BeݷF�4�ȓ\Š����Ӝ&T�ċA�ɵKR��ȓ�|%�U@�otX�Ԭ��
ْd��2����.;l)P� K%Z���U����$ˋ&TZ��!�8�~$��S�? ~|�B`�7�Y@4��:F�y�"O�	yk g��	�7��)�.tڇ"OL�r�g�oЦ�����%��DB�"Op��@���s�M���:�"O����AR>Q�(���摼R(�)�"Olث��K�&Ʉ�5��5{[4(a"O�X"Q�
=咠Rp��&h�����"OL� 0_v����<X�B��"O��h`��Č�� 
� ���9�"O����hN!2������'�΍�%"O���j֡|���
e������7"Oơ�RoAV�Vp�NWu���@"O�tIթ�tҥQ��Sj�Ъ"O�@�m+uX:eHsc�)gl9�R"O"EI���ډB���u�rq�e"O���ǓX  @�C�%�fbw"O�A���w���6�(��4v"O�h���Z*.TȦ�		eX"O�{RL�3�|If�6Nʼ��"O�E�F:("6<cӀD/r8h!"O캃iL$?�y�5������"O�e���)��刀eM� �|���"O"�A
U�)-��r��D'�d-��"O�Ӷ�m�"��!bN*K�p��"O~h�Qg�+��c�ʟ��~ ��"O ���E$Ay`�G��9�MA"O��i�Ϝ)bb��R�-VH"�J""O����D��o��(���.5�p��P"O�M��;��KV!G9��y��"O^�[%�Ԛ~�&���!My�Q��"O�a�g��ل��P�@9pV1�"Ov����K7+\t��,�''�(`�T"O���#fC�^�����%��/��1"O���� ;�KĪ����rE"O�l��i��i"�����z��)�"On!h��yMP���^a��U"Oj��) �/	�"#(�9?,� �"O��k4��)~:�𶦃�-vc�"O�� s�Y;-2 �4喃RD��"O�m1eKP�c4�B�51��P"O�<�6f��LW��&�%lV(A�"Od�Z�ї`�!C/��:�a"O�t��o�}f�1��ğ�j� Ёu"O�i�Þ #\�TÃ�F�H� �"OX���9��Z��PN�+�!�D�@k����d�� �rH�C&�!�dIv�M�����}��d,[;P�!�$Ե	�����p �E�y!���
����F�R�A��bI7J!��D
Qê���	C���!�ۤ�!�D�$`f����+>h���^t!���6��"N�GGl<r'��^!�˘f�`(q��_)X�)�VcZ?!��<6m��p��/�j���Ò4�!���P�Ag��t��	�!F�=�!�ʶ<�0�!J����� Ł�m�!�Űu!�	h�gZ�~c��CO!�䙵<h�Q
�f�i����܆�!�d�$?���!���cTl�(N�!��N 
�h$8P�Ɋz�UX�M\�;�!�䃆*��أ @ྐ4&��>K!�4@>u�d�hk��@r���!�U"j�U��$�L��
"	L�!���.N�`���X�L���\�{�!�� �`��Hk@�x���[�Z�"O����-�q׈�:gJ�-�Ԅ�S"O^�v�̂&5�R��ͩ-���"O�\RR�OXRQ��ܧh���Kg"O>%]�?���3A�Q�/��U`�"Ob-�4��XT�y�	ڢ6�0	 "Oz��G�0"Qh6O�39ߺ�$"O���B�͛T�����n�&͎uBu"Oz������y�:ّ��'	�T�kp"OV���ͥvb�C���f�����"O�]�tZPy� ��%W!�)����$ړ����_1����{R�Ц�o��'|a|�BA�(��كE�+2�@e���y���k촄Ig�l`���B��yr��.\�*�:D��)^Jp("���;�y��/a�:� 3��Y鰄�O��y"��̐��ȀR/����H��y�.����-J@�I�?56p���S�y�b�	o�J}b��S=B?l�t���?��'�Q�g	X�`9 �l	�4���c�'� <�f�:N�҄���
'��1�'v�3��'v)��XC|I1��_�<AAIȲ6!<${%/C�9�|,[t�v�<9��11j���[�� �hS�^�<d㍘?��<+�]5�: �G�u�<�ҥ��(��E�U�ӠXr.œ��A]��0=a�FO�;�t<� ���p�˒E^�<	F*�-O�. ��� ����X�<�0#�.�������H� <ӳ�H�<I�%2z���PcgU#1�����A�<� %�(���b�c�e�n�p4"�B�<��!��/���W�b���05M~�<�u�� _ ��)��V�{ ��3�eHQ�<���'�p��c
\N�#�K�<IA��0)����&�!�1��_�<I�o$���3�V�6[ʉ^�<��oW 5�*]��_|<���@P�<���^] ,tX �Ur�6�J�RQ�<ACLQ/l�.�gD	U�����L�<Qq떷���� JQhj���f�Q�<	u���3dIat	V�Z>ʨ�`�[K�<���B4o{\;�
 �F����FA�_�<	EV�$8�����xk��]`�<q �V?�̽##f�>I���˲�f�<�@K#3��	�W!��v|@Ѳ��G�<��Κ?|~�y��óP`��hpc@�<iWBȼfXa�U�줰�^���'&a|�H�	�Ԭ�3%�wp���)�y��N�$��a _�@��Y��
��y�S"&��E�ʹ~�X�.�%�y�솴1	B
(�l��P���y"��l
�t�MO�+���7  �y­ϖr�H+��XF�{O_��y2M�	'�\���W06�{a���y��� �b�0�]�G碹�!V�y�O��U��4*x�(�w�E�y�9���7�БKr���/��yrM��M��EU�-���JY#�y�nK%ZCD���I�9BV���Mڲ�yR/ߘa�Ԁ3�l\IŲ�9��y�$6��"6%8I��U�u���y����v��X�8�"�φ:�y��3f��I�f)B�����K�y�`��{�P,��D_�C)�I[�͐�y
� $����/]dՁ!��J�I�7"O�������s�F�$=����"O�ez��B_�1����$ui��'C!�ªEA����y�JhQs)�)c�!�D�.sZ�A�B'G6lc�T��W�g�!��T�Hɱ��X�-D�H�'0�!�d�B�e� F�)����f�Q�!򄆭��q�%@�ycT�
W��9:�!�䓿)�$�0Q�[<;��%.K!�D��k��C HO"&G�9;BƊ�-i�O����$�`σ]dГaC�2A����
�'�|l�"�.c""�˰NV4(�d��
�'�lpc�^�@��D���&/Z�	�'�6�����^���Kc5��M��'7�\@ ��6�E��2�:��'�P���,_�1 i����S~��'h�#��ײ(2b1K�mҗaj���'F�<`��El�R�y�O�*���#�'Yܰw�Y6/�ꌳ&kB�'�&�
�'(遥��T(<bVBG��&U�	�'����^.v�zI���ܝ=0��2	�'���a&� :z���6֐��'�젩�ʗ"��<B#�^+;���a
�'��\p1���h��Mӳ3o�=�	�'�4�p��ck��p�L&Y(&$i	�'�jɨ�''�xaV5X
�+	�'�.%�^A��)�J��E&�5�	�'�riq/F:.�
���X�R��e�	�'(���wb��Ii�02���G�8 ��'g��*��}@��ݫC� � �'�qpc޶-�
��R�J�0l*�3��x�ѹ[����I:� y�=�y�Y0^	T��pOG���&��y�P��9��P!T�P`E(���y���jٸe�qc��{\�	ɔ���y��W(5h��r�bR0{�"�����yҤD�n:�<��:w����W,���$.����'��p@����	W� =�6A��'�z}�g	~��\3�K�'9����
�'^m#���Ńb`�2 ��!
�'��-3���l�n�HY�)�(m��'	���ʌWn�|��8;��)�'������5�[�0���iR
�'��b!˚�򀴀0�WX�Ԩ	�'��tc�'@�c�jLn��H��	�'�T�"�A>(�t�XW#�{n�Y�'�@���,�?eS*�����|�r
�'���pM�uY�f�J �d�	�'s�13,44� � B[<��'�<4�2!(#E�sB�q32�'��ʦ�O>e=(y����iCZu؎��9OvM�%�������!P̼%jW�D�Od�D�O.�$�O��'<�N$�Z�^�9�&���e"O��H5+�$�Ne�f��9�� "O��IC�4>�d�+���U)v� �"O��1��<9v����;\���"OXhx�#�tD��j�
�pz�"O&�@��ǋatPUŉ 7^����"O�lӡ�» �Xy�g�G?$u��P����ڟ��	ğ��I�\�IG����=1������F07�d�����y�.�1*<n˓爉c�h�����yB�T�w��鰆�b> x���yr� mZT����lߜ�s��+�y�mqUD�O�.b	d�C���y
� L��bX��>�`�K��rU��qq"O�=�M�<l�AK�2%�u�7�|r�'b�'�"�'�?�7#�(B�yz�kU0]Y$4kG�%D�\�d� T�h� ���B�R�$D��󰁌4�����@:g<�QE�7D��F��_��M�R�\�"�4D�p�'�֬x�T`�N�	F�֭(Ҋ7D����ߚ=9��gˆ;T�U@D)"D�t����e|�1�B'�.�ЂL ���Ox���OR���Op��4�D��Q.�dk���9�h2,��<��Ð.|�xx�k�wդ��0��p�<Q�K�`���p�N�@Y����GXj�<��"
}8FjZ��n��v	AN�<i��#�A��^: �9x�b�F�<�'Zx,�(w�܊R`*ы �	yh<y��� [�,ar���7p�
7�_����?����?	��?�����)�5�F4�5HH�B��Q�ѡQ�!���}	@���J�@���ƪI5�!�ɥ�nݸQ��2$�q�K�,V�!�d�;>gz-��d%��(��&l��'q���bF{Z\(C�K��w�p���'��*��eR��ql^�i�p���'��T���U�s��2��$B����L>����?���?9���?1ΟxQ��S9HO�u�pǞ�_�ٙ&"O�����D�K�e��c����"O���4�X�� JE�><�J��"O
5cFN֙%��8��	�.�X�!6"O��E���zP���0!��	v"OH��gB����:!M=P(B|�P"O�eQ�/~�]3�䄋$�|�'Tr�'�b�'��?	���B�|��V*K;Y�졊0�#D� �0���*~��	���?���a��!D�|��-�~�@8���9*�\%9l!D�����U�/��e��n�s��ץ�y")B*J|z���pg�M���y���M�L4�T�� �N��#@Ҩ�y����v	�,ׁq�p��թ�y�V��f�/q�pt�u�X�<�`$�#�젲CZ+g��ڠ�[A�<)t���X<p( ����/q�$��j�\z5ϊ.kX�e�eS �:4�ȓN�v #q���V���$$C���T 0�Z��4���G'$�Ԅ�F��CJ֧Bdn��g)�%��0�ȓ<&�10!�9,hI�艕B��m��-�>��S��?���ʤ"���q�ȓN�M
צT<QD�K���6s�`��R���0S �f�R ��hʎr,Єȓb����u�ݒ<����h��<�n���o_B�6ȝ�!.�!�O�o���'�џ��<�W��$��p��M����wn�ٟ������w�[1����M�^b��ȓUa�j�G��yBG(�����*R��?` �����p"Odi�"�^�b�Nu�d��dB�X�"O �r��8%��p�eK�7(�`��"O.II�"�?	2U�L=?!XD��"O6)�V��;K>�k
^�{��-+C"Oj(�K�� yEC��0�> 
"OT�[�IC.,ɐ�Y��A5[b�}Q�"O��)�΋�0a��(��utJe3�"O�aC��ܲa�A����"Ch^3�"Oℛ���G������<���{�"O>��f�-�<�&�N�f	��:"O� �B$w�� '�=(�dH� "O�8�-:�N�a��S��T"O�@��'���~�kq�9U�D` v"OHM�Ly����2K�����"O��r$��<H�xٳPn�����"O$!�a,��ED
�0���c�L��"O41��']Y>������w�\�!�"Oֹ"6��s�씫��<��B�"O�Śh
>�x]a`��tL��"O�yq�% s��:�OF�!��dp0"O�|���D�r�D�CR�ޝC)0��"ON<�$�@�j���إ0����"O�I�Fl^s�f���./uT�F"ORT���ЀQ���Y�s ��"OJ|9V��-±�glQƺ �W"O�QRq&~��p
�ʐ�g���4"Oz��E��M ,�8�ʞ/
��I!"OP�ۄ�N(���� k����"O���Q�;$qI����$���X�"Of�`�͇$g��r�:��yI�"O�C����w�\I
P"K2v,���"O�Tr�I�ZqfUϕ�L\(R�"Oč(��^-T�P
E�\SM,t��"O�8�qk8[}l BnU6=��"O*dBu��4x_�P+�R�tdS�"OU��(��rZ��0���H8�"OxT*�ŕ�K>P��'�J�O����"O©A���2#R�x����(�"�"O��P7u��Ö[�Fovha�"OX�26�	�`#p�P�LF�,A�x[B"O�����	 �\A�W�Т:��h�"O�hy��V�S4�C4�Ƌ}<�[&"Oڝ���@�`b��8x)��"O�]��!bN�Y��9r��y�a"Ob)�2���Z��K��m�l-��"O�!ie��K7<$�5�j�5y�"O��r�[)Bw�٢���4�2"O�(h���4%�H���r��,��"OƝ��L���YqN� /�n8��"ODE�$�E�O��c.�(Y��UA�"O�Y��~\�-�4A0�P�"O�M��$(T.h@!�P�
��a�p"O���!�I���;3�� MD
���"O���!�
��Ttd�B�� c"O� W��J�X��W䎽T7���"O��X�@C�w�l��Ë�<�pUz�"O"�q���)5G�2&�("��t؃"Ot)��ӊ$�NP¦�\26��4K�"O�� ֮��]�\�@��B.̄��w"O�A�4�����(8Y�v�s"O�L�@�(@�����<�R�0�"O�	�,ȿZ���J�)f��}"O��$F�8a5hѨi�,Er��"OJ�3��֒dt�����?��(�"O\P���'^5�UIc1@����"O��i�`Y<�s╶q����"O4 X$H]�\�0�K��˒ko�d�"O^֠ �-˰�x�bЯ;Y���"OPu�;Eh���|F�A#"O�%[���ǎ�@6�!I�"OVɱ ��$��2'�?%�	z�"OB��%6dB@�:<��@�"O��Y��2G�Z(�1�6����"Oj�B������F��&<R�sc"O� \T`�HS.>X҄�Va77x�V"O� b��v�@J8.+Ra`t"O:}��/?��pcB��".��F"OD8sn�3E�p�)<�:ѯW�<ђΚB����*�-ext9�Mm�<yf X�s9S���B�,�2 Q_�<I�(E�A�x��ʩj^<�H4��W�<����<� jSiN�2~����o�<)V#�p^\0o�9E"�-����a�<I���#��}�*
5 /�i3��v�<q!��T�NQc���/'�Ӵ��yr�O`d�s��áYۂ;�"�y"���|�F-#�j�=O�pS��H��y��C�|����)P�E�}i��/�yZؕ���ɄB�lڳj
9d^��	�'��A,Q�Dʲ�ѶK��e�	�'�@��!ͨ��E��'vBܓ
�'Z�zӁö^s �3VEC�ͫ"OlI)����R&���r�ޅg@z�bR"O�#l��rYqr��5:�"O������9!$�9�d�2p!"O*�qEY.r�8a�b�J*�ن"O�Y0ԧ	���#SA�)v�eH�"O:]�2Mk -�5�J	��(w"O�t3�ο)Yt�;&&3zLN��"O@���"N�/�"��R8j�9`�"O�ժC�&o���B��H��"O ��S��+~>�ys��1��̳�"O�!��t���H�OZ�nm�p"Of��.#-2iz����9����R"O�UY� ��-p�qq��,�\��"O�Px�M��SV�jԨ��&�1Q"Ob��%��V<DY�m�
u���I�"O<QHY?]C����DXNx��"O���K&Lzm��A�S�"O��v��;Ո�ô��kX�"O����(��'Q�h��kas� ��"O��"�ϙ�.tIҪC�6_�QD"ON��b&��Lx������+%t�23"O<QH�fy�Q�A[�AW&���e���y��+R��)b+H+0��y��W�y�%�%5̦1�)@0"Ӥ�	���y���M��s��ڬ�g��y�Yz��h���� �I�'�џ�y2(��pM@����Ȟ�������yB!�!�T�Z�'B��#����y����HŻ�pL�" ����yb�*�@%��T6�(�Р�Έ�ybbʎv \��ֵ~r������y�L'P��eY�lW$��>���ї"O�5(rKS'd_,�
S�	�=�(!�"O��#��	-Fȳ��S�K�����"Ob�[�D�-�A����\zB���"Ox�����k�<;�VY���kB"O�(�s��:s��K���O㖅��"ORy(t��>\�PD�c��	�8�*�"O8�cn��(�XЫBN�2kԨ�p"On �gG�hK���#@�Q`��X�"O!�#�\�[]�廗C��=�L��"O��R�j�O����ռ�͙"O��uNKK��YS@��q�R-��"O�U4�&YUȑ &OԴp�H�0�"O�E�'	�wH<���Y��(Ja"O ċ��
�o��YXvL��ݘ"O� ��q��628��rRk5@�j#"O���aG�>�ΌB�*� ���� "O�1Q��~�����(�}�"Oe�V�Ɉ��1�M�O��w"O����72�ԩC���B�p���"O� dd�b�|1��x�xA��'.�੡f��9��Q�U�O����'�D�s�jIwC���ț�C(*���'^0�@A_�QJ�m�#ى>�q��'8���T�s��`���"Lh�C�'v��; �T>g���捻����'Tj�bR"ǽ���肢M=S"�(�'4x��"��13��9�'��D���'ܒ���N4�f��Ү�,�X��'��!�l)��}T��	�'�^��s@׿��P����1G�I�
�'��9��?u(0�DR1��'jp��1I_:���$c�x1L���'-� 0�	� ����&/U�pp��Y�'���Q���#�!���1#N���"O��b�gO%l��� F��/��3�"O��P��T��=��g �},�!"O���Q��&p�`x2r�R;Q�i��"O�Mc�	�Usn=0o߉6�P�`S"O�d�T�[Ot��d��4��ڳ"O��p!��2o8��
A悪!�4P�"Oܰ;q�B�l{6aq�E^�T�c�"Oh��HJ�}�J4�&�לM�Hِ"O4=kË?�$%�'��5�:�5"O�0�)[�4�<�&Lɐ{=Z��%"OT!@����u:lJr��w6&�YP"O�(R��<G�=��$/���F"Ovx*�#�/c��`p+M�2n�"ON�[��%�*(�Ϗ�;���ۖ"O �P�"^�D�酥B��D�t"Ov������(��2��aE��V"O@�ٱ
P:k�YY�*D;�l8Q"O��#�eI[t])3�Ȧo�vMzD"O�L�0(Ԡ�z��	IX��2"Opi�Qf�.W`�m�� Ut����"O>�+����	���#�a�"O�9$����h��D�eX�]3�"O����(�,p$у�¿QKFtcd"O�`G锗&�I˵M�ZIp!˒"O0�H�Ұ!Yr�� �
�=4n�F"O��I�BL'm*f9 bKW��T"O�9����Uy�q����&
�x�"Oz��� _�zg�<�BoЩc���k�"On �V�<���ӳgP��tq��"O�蹔h# i��'��X�$�(#"O���(VGjV`�oԐ �hD��"O9#�r���P�n�nU�ib�"O�=��d���DB��֙L�rs"O��P�T��)���+,*�)r"O��qP��*b��@@v�H�T��`��"O愰'EE�06f,QĮ'��`�"OB�Iw�)5��B@�H;@�^��"Of1I��P�'�P���v�|i8�"O�r�L��|��x����:crn��6"O�h��ʄ5�01���:I_�y�"O�L����<��P�BLA�XG���"O�m��Q�����%�653��y1"O�M��ݏS,�T��0A!��"On�����rGD krn�>u�� �"O� $qC�I��}���ږo r>|�2"O��aI�T{�hҒ��K�&�#"OtmY�U4�<��ؒ9���y�"O��$��y� d�7�
�^� ���"O^�٦`�1%:@���JߦȚ�"ONܠ�O�v6����S?K�Dq�"O������(����U�{���8 "O�QK��1�n]q����D��"On!�E��@m����B=�"O��q*�'"8f%8J�
J��
 "O�Pc㪙-*S���$��#)�F"O���`
Sd��XP�R�,�Lĳ"O�ħ؏c'�y�@��>}B*�+T"O��G��F��%,1iHX�眬�y2���J�8�&o�n<:��Q"�y�I�_��[g�!l��ջ���y��)Tq��E:�V��A��y��H�~9��"��",��`�JV��y"+�>�P��T�*g�X�@�^��y���5T���c�J""��(wiB��y�/�|G�y�B�K��-Z<�y2,�
#)	��?��1�VDǛ�y�À5��Q��ؠG�|u:S�д�y�R�N�*hkc�	�I�
i���yB�?h�@�!È�@T{�	D5�y��R�	�ց)��V�f�z�S&�D�y�kB`���\�/��2Ɲ,�y�h�2�!3�g� z"�)��W.�y"���n�x���.s�,��q%��y2�%l��v���m����P���ybF�Md�L E-׮[)�ف��y�*�CT�#Q��aĜ�
1jɸ�y�/M�Ru�Y�W���`��ya�(��1h�z�>3������^�z0�؆�%���I@W]8Zs̆�b��<��[��@#�,]d!���:N�\��ȓO�tX�$��J���b�d�4['���ȓS���D"E�F����Vc�+$P����~� MU�+A�5�,��-Ĵ���qd�I���H�
+��SC�ݪd�ʝ��)�������(�:ܓ���Y�^M��x]RP�R�_`d�3��[=�Ѕȓ���g�՟Y-$��`	?VO܀�ȓfx *$,��$(��� 8᪁��1�^R��V-��0[%m��rȆȓ���IBޯ~�P�%�R|���ȓt���)G�^��� 8S��,|�f�ȓc���eLŴ)���r��Q.L���#����e�W_ްqE^�@X��<T�-�%W�*,�Q�	�'0߶i�ȓyJ<IG'C"N�����8�ȓ.�0ׁ�5W'~豬�d�L�ȓpȈ���ݮO�0��$ ڔ.TlՇȓW�^8#��;�I*��	p�>��ȓp�E(Wcň"o�!�bG�t������
a��� y���9�K�w�R��ȓ*���I��W���A�{�f�9D���!O�	L�-ˆJ�y.��06D��kUk�%*�ٓ��"MR�r�3D�s�nYJ��0زI7h�Wo%D��s���UF�h�E��ґ�-D�[ʋ�`�fĊը��Ӝ�P��9D��Q�ƃ�n9L9���1`Ә� �8D��������y3�, �e�aD*D�� ��r���+Y�8�0�� -�p�js"Ox�����)t�̕�d�Us׶XD"OB�
͢u�6�1�^�d"b"O	����OH���Y�Ă�"O�*�n9N��P��U��|�R"O,�b���5��uj�A��S� �"O�4zbk
�&]�T�`����"Opj�.�O��X*U��4�~@��"O 2�'��]O��9�iƎy��X�""O}4&��DP�$"4c�!%b�9"O�����)h[� ���Ň$��"O1�%�\9�vݪ��;?�@�v"O9(6�MuR�������&"O��8��&|����CE �6�꤀�"O� ��NV�j�H�CR�Ytb�q�"O����\��t���A��aY "Ot��em�	^�)0���H	Z�"O�ͳ�B��v욇b�>:R9yp"O��J�&G?\\�{� @ 21��"O����؉$��F��Q4nš1"OV�a��1�R�Z3��#O~xs"O�����(���#F�/7~h0"Oꠘ�ǿ!��S��3y4H��"O"��!�ǜ`(}Z��?b�@y��"O�(8�
J�
�����T�Pĥ�"O��#s��s�"\)��	�d��"O�p�Т�bk|9"(�H��h "O4�ѱ�ι*w��#wg�>7�	R�"O�}��狫1r�hh�K�� ��"O0�LA��n���_�:�jV"O m�2��;�ܡ�&
�9\�=a�"O���l�"�4�dϽO�va �"OZ�0�٦6Hj�ru�]�7�V%YT"O
�b�:�"!�@�X<f���0"O��[v��J���9�0-��"O\Q���	�d\Ȃk�:_�F�(G"O����՞��|��G�t���"O����bϪ7�F��J�$&����A"Oz���*�Ti�`��0B0�)W"O\D�ᯜ�#L��)�1c����"ON��"�^���0#���0Xt�AG"Or�y&�j�PZԡ�_��"Op���AƏO@�q׉�%:��e�'"OD`5d�j)2���$K�p$"O�p(�t�E�$�=��p"O�)�b��	0��×"Ԫ	z�P�"O̩�D�
6-�sSaWb".���"O��`��ٿM��5y�O�Dr��r"O�h��I���\)֡o����"O��r������V�G%UR����"O�l��X�
đ"��$7����"OX5*��֦v����g�;%�}�"Oh���.B�`�\)���J�E|�� "Ob!��E.l1�K�Ay�!��"Od����WWv��Y�h0�(%"O�)��M�p%*A�7�ɩ��;""O��yE�I4{�h@a��]�jpg"O���A��H	da��<s�j��t"On� W�
�U4��Zu����t��"O��1�D���y�7��_���3"O��V���=��M�&�2P����"O�ȣ�
���T@`��q<�F"O�� @���I�&l#k2y�""O�4�2�� >�<LI�J�4)a�EC�"O� ������`LD:4��`�IP"O��vN��D0�w�O��X�
C"O���Vl],�&����T�bդ)�D"O4D����ܙ�ӧ��x@�"OP�d$�%¤qA�B=z.%(�"Opm���C,h�����dM6z�hrp"O\`9C��'O<�;fC"���qD"OP��!�F��8t�7`G	roe*p"Ob�K���p��a�s��ɼ=õ"O�p�F��v!3⇒O�z=�R"O6�Z׊�m舼5a2&yz4��"OZ���j�y
�X�Ѩ����"O4�����Xq�c��m��A`�"O��a���p���CU�"VA� "O~� ���Y[�P�¢Y)A���"6"O`k%�6�\�r�^�A|Ƹ�""O�dK�fغ��=ӡ�!M�Y�B"O�!hqĕ&��£`҅1� ��"OH�q��;���ӎL�e���kd"Oh����	�P�`�<L��@�"Oj@�CM߅D}�w�ȁ+��4"OPa� @=9"Na{�ΐ��ѹ5"O�e�S���V��(�P�.� a��"OR�Sa���vQ&�ۗ兩C+�1z1"OzEY�LX�E�����A�����"ON�:`�Y�5��ջV�F�"O���EޥM�x[�-G����b"O�xcq�ˏ8ِt[ cΒP�lы�"O����g�''7N$bBƠH� 4#g"O�Px4có$dh��f�|��`�"O�|�ag� ��\�1�\�S�"O 3�∳/�l=X�
ӵeF%�$"O���u$��5��si�5UHa�D"OX�i��!"z�U0�,6�$�� "O4�����3l{^	�s
��E�9Җ"OΤ۲l_�`��#	A�Ro����"O�I�.�'��j�蜆�� �"OrJ��"��
3H�.QZ�"O��%�xT8IE�,Z�e!�"O��C��	3b��D��jҢ$q
���"O���"�,'4@QƩ¿Z]@�"O8�Sa�BD�l��.�?Y��4K�"O�e����8s����+�(C����"OȐ�G�''�F�7��?��9�`"O"1�FP�nh��b�F�B�"Oz8a�L*�n�" b��L�jW"O����`F\�i[b��O{�Y:d"OLiaR������}pl��"Od�aÇ-Y,�x&�::ilQh�"OJ *� �;H"�)����#TBP��"O쵈%DC�_��a!�Q,@�NX*C"OҘ���4����(Z�^BD "O�4ь�<`�0�g��L.��"O��Iaę�{d~�05&K�%��ڇ"O�i�$�-s��A����/|Г"Oе��k��|B�Y �P�Y u�"ONP�R�T�)�BՁB5*��:�"O��BR��$�:\CS�	����"O�Pj�X�%=`��Aߥ�NY�"O>1�s�D�
F�x�e �#{|��w"Oΐ�#Ulġ`���'`�%��"Oz  V E<L����6O�0KU���"Ou`��P#H��:����X=@�W"O�u�NX�=X|��P�D�$nXs�"O� J����V��hY�4��1"O@�g�[�@�vh2�ē+��;1"O��0O�̑S��=͎�"O��9R+�-R����e��@�F���"O�a�҈<U�)Q����)�"O�I8����I[t8�0�䍲v"OB��g�3$_"�:Ƣ�9W�L�"O��zw�ΊPˮb˟���x��"O�q����/�V���X(5�pQ�$"OR�P�� �a�r�b�v��"O6����@�^(����[X�1Z1"OI �'G4�V��|F�h"O����IH"8�TL�Ag�wP��!�"O����NЫ6� ��&�3]f��"OR��A���`����_�z��4�"O�4���ߨA�R�pw$
+�¬ d"O.�hC@�VƲȨ2ɇ;��6"Oؙ31�L<Wt��I�MY�X���"Oꨱ��L4�*=a7zؔ��E"O(D�B�G��Uf�u��0�"O�h�w�[����� �I:䬸G"O�����tK��s��+\3tQr�"O*%��+�1(D�JP�D{���"O���o�"��l�aE��&"O����/�5$�D�#l�P$�L "O�|��P�j��q+%	�D
��'"O��H�+=�!�bK�`�*p"Ol��u�ѱzPDժ̛=i���"O���"��#Ħl2�jC�5��xI�"O�pP���q���hK�|JL��"O"�B���P�
��#��j�l���"O�� ��װHWv��"��H�&�y�"OZ��T�(g��ĳ�d�<�h��"O�XRd��>�0�s�;Ȅ�["O�q�r���0f�̚��H�QerȂ"O���E�X�W��8�柃[
$J "O9P�_J�@�Z���,@�-�"O�Y���'p�iZ�,��g�.;�!�d�Ms��;S���6J���e�C�Yu!��'@PIfCY�6����2FO�5i!�ֆ�qbV�1��� Ug�Y !��V#x��-����~���E�b�!��E�09���-vF����ɑ!��R�}ʝ3��Z[��0��H!���X��e����gp��)���P�!�$Zy�9@g�P� �,�"/K�{�!�';�8l���56�t����!�DS�a�F��ޞc؊9�����Lr!�)S���aI-s��,r"oӎF�!�䌃$+��CУ߱E�B)�T�U"�!���O�>��E,{T��9��X%�!�$�A��{'�'YH.��!
�B�!�$�({�r���.H0Һ��p%��!���;#��Kv�E���p��-!�$D{��$Q�ǀ4	Ÿ��a� !�!�D��]�Qp�G�[����bG0S!�U=&�Nkׂ��y� �!DD!�$�i���qR�+N�8	�@�a$!�DN�g9
��Vi��jq��'�!�dh*�����z�D,a%/��c�!��R��\�̉0 "��d�k�!�$�f�X�P���5c5�|�T��%�!�7!{�!ɯ'44�V��7�!�]	~�|ى1n�<x@~�)#B��!�� z\����s�S>D����"O����,�w�d�
wn�(����"O����C`F
�렇%��P9�"O��2����]h� ƹ�Ф�"O���@
=x���C�
�^g^��B"O�(Z�̟>K�v{bD-r�\�f"O��i�5\����͇b�\�xq"O' �,T�tT��6��5j$"O~9�� @�
z��S�"�xA"O���
�ii�r���-����&"OH*uGR���<%�9i��s"O<h S�SV�H,�¨	�� q�"O����"o��=��I�(��tqG"O���H��LQveR�JU�`wNU�"O���3n��#>�P��[�o:�	�"O�D��C *B��[VĜR:���d"O��K���&�	ғ"^�Y5@�13"O%��(ğw�E���)����"O���F�?���� Z0}���F"OȄ�Y�fU��S��AKg"O��Q5@\�A�ܜ8�$�r�\��"O�]
GI��8��`�*�;B�"O>|Z���/F��9ei�7~Ӥ��"Op}S��]ULH�r�^'[&��A"Oʕ��B� ˂	�"�$�&"OD��gk�v�ީ3sV��48{%"O���'�;R�Y�A��\�04K�"O6l�1DB!��1��E��'��I�6"O�P ���R�8�q$	�2x�"O����0�M��D@ {�Ҩ��"O4,Aw�ӿA>L
�ep��s�"O̐x0'��Z%��q$�<�@١"O����2MX��7B>$���"OĘ�C)��q]���¨�\B"Oj���nt�<���JHXh�"O(�Tٲu����AV�&:���"O���$`\]{��CO� �u)2"O�܀����Uъ|���pu���"O�k ��dx5���j�5b"O�3r��9o �]xB�W,��b"O�0K�l�1do�(Ksᑩu	Π��"OH܁cb[�
b�y�`��L��)��"O,��@�n�>h3g���(���"O�$����^��ȡ�m�8B�ܽ��"O��#��	#���C��
0"i�F"O�q��*,@8<ZQ�#�D��"O*̉w��)�H-�J���"O$J���1Q���5"�E�Fu�x"[���<�~:��=����  �L������f�<�RB�z m�1�ֱ/��M+$g�_�<�U*� "��僑�����)V�<I�a��.lL��ǉ+��d+��U�<����*�da׋�0�"��4��T�<i'@�3]Z���Mv>�Ä�=T��i6��[5qՉ�c�v�a_<!���6P�U����*|�.��R��\#!��ԧu���
t�E����vAW"U!��_5g��AwH�=zL;��?!��'z��h[��/v���Wk�!��F��	ےEX���;v���!�䂂;�<Q�AGت�~x�IPA�!�$�4k�����ȱn�NE��GV�s�!�$�4h����I�F��`8����!��Q��%/�,ovT�s�&0�l���� ��2D��T��=�e)D(H�J}(C�'���>z�1�� �)���@��W�X0		�'�d��_?�~0)��$VP
xˋ{��O
�}��hl� 3FY�pGLtZ�耠*� ��P}.�YыP�KZH �Q!�3��9�ȓYz&ؐpJX�x�%�`k�+Jޔ��Vmb1��nä!�p�҃J�T�ȓ���ڑ	�M�s�ܮ"�X���`�&� �	+d�I��͒�@�ȓ��d��a�z��uB�5Kb.]��	\�$� ^�2e���.�ahQ,ãJ1!�D��$��r�/����7��}-!�d��z^���3�[8L���B�N�}Ҝ��%�S)pTL���#�Ch!C�#%D�h*F�[�~tp�'m�`���%D�T���68��2&Ԁ�VQ���a��Cተ|	�Eb�^�*���KmҪwTB�I5I��L�6�/.nڵY@��8�C䉪CT�P��͡L�f��D��/N"C�	�r<� ��4wL	6��<D��B䉏!BB퉆��~��y`ELWMU�6M'�S��M�AKJ*W�B�b���S^L�2�
XQ�<9\�J�R+	�4)�$2���N�<���o�����ƍ6_�f��fMJ�<�u�v�� 1�P5�
�@�G�<Q��M\�[�"�u��Y�Oj�<��,�
�T���^�̤0/M��D�<	 o�q\ƕi& Q�Z
��T�ğ �!��Z����y�k��3ؼ͢S��~�|b��L��Θ�>m���YQ�TY�L>�yB��8ZT\J���;���hc�.�y�
4^XA�  �2�6 ����y�ă�	6�M�0 ���d�8�y�LE&rB�h5�W�(�Aw��y2툀x�:�
���J{ m�G
��y" <uh�aqf�F1�%�v@���y���`�<�F��'0t8���;�y�N �9�&���Φ3�� ���D�yǘcѶ9���Y:[}�5	pgݖ�y�N�L�\��C܇W�j�Sp�Y��yB
�,��a�‴M���Ԍ��yR�@��`�`E�(1WI��ʜ��y�E��8�T��2���<8
��#���y�D�5n5ڸ`�&԰�����	�y"���<�PĒ7S�>�˲�?�yҠ�1$FƄ���H�Qаn��yB�Y�L�}:��&)�[� ���y��"ytPU�ui��4���N��y�Ŝ?{c���ce����צ_��yrG:A���"�K��~����F�V�yCs�Z�2@,��I�M+�ʖ�y2
�(�X4`��2tT8�'��y��ϡ�����$1��*�@���yr�b�JuX�!1�6�*Ѡ�#�y��]92��b4����q�W�y������
0� �J4�u���y¨	�r٦9*��J�fW,"r��ybE��]K��;Y{hi�A��7�ybG�O�䀀�H}� �����yB��{�� S�����BN��yb�H�&x.Y�S��p
�)K����yR��O�4��bM�l��Iz��H�y���9"�p�6`��+�%���y�c��A^��i��F�nT��;U�8�y
� ���5,�9j�k�̧I��a��"O ��f�5�� �S�����y�*O��Thö��t#�悅/�����'=8�*q�R?UUD�rN_%�H�'�jy�g)���䂫!���a�'�Z�[uJ�)� #�-��=�x �'.��q�*�: �%�^)~�����'���@#�ܦk^��^4^y�UI�'�Z�Rf.�8U&�)�����	��m�,)S��F,'Mb��"%�]<h���&�P��=F�A���۴D�]�ȓ`�Ī���9���+�Ă:E�5�ȓ��l�7�Ĉ~J2 [���m�؁�ȓ.�L� F$*h��I**���l��xp���`��@[�K�#���ȓ��u�
3Ԃ�ʴ��#N:؇ȓ.�d��2��?3�lIu��*I70��ȓC�t��Q�K�8t�*��.t��)��L�d��$N��أ���(y�r��ȓQp�+v��,k(L�b@
��{jV��ȓA=:d���-	b�N��T�Q�ȓQB��Xw��O0B\ф�O"$a�ȓV9�Aɓ��

��m�Q>B���(�P�:�.�F��Ԓ6	�F�Ą�t��a`���0xAf�츄ȓO�����Z5y4��q|,��ȓ����0/�IkJ�pȞ�9�n���s|e���<$�M��@�/���ȓ &q��ۣo^zc��.P9�ȓrX<�R̟�~`���	�7��]�D0�Νx��]b�FF.^#����*@��"�)�hJ��֬8K���ȓ,f~Y[#�J�洁�Ș�8�PU��ZY P����9c��7��i�ȓ2,����[%(h��f�`����ȓ���H��oa")76�LH�ň�b�<y�E6]�\���6 J���5�Y�<)�N��!R��7��봁�y�<�7�� C�6�X  V�L3e�&�<�2J��U0�+E��0^�R2I�d�<q"�	�N��,Ђ.Uе��x�<���A*��	ֵ�k=l*�)P�<�d�L
~��S�3t�z�)4��g�<预>N�	��C��$)LYdI�o�<��'V�!���"�b�)#\����j�<A��ڭ-Q�`����N0�!�a���<ag��;zv�3�49�xG�J�<A�D�2{[�y��؎'Ȥ��Bi�w�<�v��w�`��a5�IS���N�<�DQl D%�B8D��P�`n�M�<93���!��4d�ƈ����m�<	f����Y�)S�y �K��f�<�u��� I�����+:?j��ˍx�<����
���0E��n��Wn��<A�X8h*� iOs�a�T��|�<� Q�uq2JU=f^zc�A�<)�`�Q��Uqv���V� �/�s�<9�X�-S�4���*9
�90oMr�<Aҹr�y�&�X�X0ţ�7B�!�ʌ*�q�b�U�d�^в��<�!�$��p�N��@���Nۈ@�W�-:�!�$	.]�x�φ���AA��S��!� *w�d�R�OM>Ӏ�y�AL��!�Ԡ��=��
�^z��GK�!�� n䈱n��HX��ޙ+m��S�"O��Y'J�)]*���
�3�.	��"O�0���Xl�����B84P���"O�)ɣ�ML��w�:Tm:�"O򬹣c�_�3�˛�~���"O((�"�FK�f��l��g� B3"O$L�3G\��y�-ͷj؎=ʗ"O�\��I?&���*V�T�U�� �"O���"���J��8&U�"O6��6ͣ�FL��it��"O*a2�R-(o|u�R�H 3��833"Of�N�/\�QG��
����"Ot�xv�H�ue��`@ǟ�%n*虧"Oj�����%jlX���W��,�f"O�-9r�=<���Aɐ�L�ݻT"O�ᯔ�s��Mh�ِ7A8]5�'�8�;s�	'�����]�xk�8��BӋ5Z
�P���O�8Ei�'���s�E�
����u\d
�'�vmHEoɈl�Xq8GFZ�ZP
�'~�)U�oCb���!�]�I��'I�%2��A� �~�R�3Qǒ(J�'L*b�P1���ɂL	J�����'i���E��Z�B�G:9��ݹ�'s\��� /=����-V�>��%��'���7�z��{��ܲ�����'�ʍ�pk�m������ $�z�H�'p,�Cr���]s�Y�q$�
�"O���P�bӆ0�懘
�m� "O$ݒ���V�z�h�f��5���´"O��KC���]�M!'\�*M���"OH )#$�
e ����E��(�>M��"OH��ʅ�_�*��v$�2t�R�"O�����ˈ{�ڰ�W��3]�H@:1"O6!�eF�1����@�ʽO��6. D�����R= <��"n	��HU+�$<D�d�4��wPb�	�P�K�=��;D��y҃�@���`
L�V�@�B7D����1^���d��(c�x��j#D������:'��11��7/�F�{�!D�8�Ba�z��Ĉd8s=Ne�r� D��A��8)tx����~���/=D�t��B���81��.T�}��@(�f>D�lY�ĄlʴuC/!TɈ��"J!D���t`�5a8UDK�MT��p�(D���E��,����j�a�h0� 3D���G��pڑ�B,�%C��g/D���F�Xr���([�EveI%A!D���!�D��H9bd� ׌�V�>D�4:j�px��@1�[$ y
�!� =D��vN��$�P����E,u�2 �� ;D���	F�"Y@�8���7&��c
8D���Gɿ�	h�e,V���SI*D�H�� ٬:� Y�8B ��jp�/D�ؚ�e��^2n�����&M]��3%,D���#b\0��Ĺ�"ڱlC��d� D���&BؖS�Y;�/č%yHA8�a3D��sH[0|��C�j��}�:�Qr�7D���iϽ|�J�����1)<��Ǫ3D�@��B[�a���&S*RT�$2D��t�@�:\�k����qz�Ƞ�1D�(k�C&�<4h1嗌f���'."���d����j�v�b�eBި�ڵ�J��,�<ѕ�ʈ��].q��K�?aI ͘�^8��J��� i8��V䌿�ƹ���Mm(<I��B�<W�IfᕸH0��$o\9v*�����Q���Ȧ{���kP��(��<��j���d����� 2��A>����!�Z#/T0lpO�)k���H9cG��m[n4�L�f��=rѬ�25|����F�m�Z�C��Ӟ�b&�Oڲ�X�O��%K�"ӪtC��� K$����'G�M�&J��@t�	�3�t� E���]��1h�*��By8 �Ҡ�W��`�u�i^y��N�EY�����",N� 9�yh'��k�h XrM�,8�OX�xd�_~����0�M��N�ם���!��B�R� 5$\�-��"Ц��l��
uӀ��*O���WcM�U�f�
���ѨZ�Vx�'�T�(l��a%*rK���)�OHѳ2A�*Yr�RG�Q(X�BH�爕=*d��aE��M�1La���B&Ɩ4�ȳ�k���P��&ʈ,`j|i �I<z�t��$�S؀��򩊐izd�#��S�?��	9u�I�)���W<w�:)�C���M�1�Ҕ"����7�'Ev,q[2
Z��꤉r�-	�4X��	���T��`X�ز@L_�P�R4�'��ɒl�H%6��*�{5���c�A1;˛6iE�WB���5}L90v�ػ�Np`Yw�|ɛ���P	���NC�W���P��JC��3���Sհ�%�Xs7��
<��us��'�m*3�4u2��S67�u��'�����OzW���3�R�~5nD���+���w%^(:�"����G���"!��'7���1%X�RLb�W:33"����~�"I�؍y����?݈2I�,B+,�4�ܚ����X(� �E���D�y�!ӭ�rt���Y��ad)�U4Ն�	=^����N�� m33�!5!F���<��	�{��y��_�b��yH�B��W������Q�&��V�R�;����d��wU�a�W��%',C�I�0���f�_�et��z/ѫQ���Z��^�or��CG�s��ju���5��&��jWҼ�Wc؊{�A�E�M�p��q ���w�<�u�ʹ[H���t!{�0���Z/[봼�E$�I����O�����e���XO���$aK������"
Q�F��c�+���	�So����E=�~d34�	e���U�E p�<���-g� �@O,ZkD(R�+S;���$�&1,�Y`o�n����
aj�e����d��vX|0#��S���G��5H�ص9�%�20�8�iA�S1�܈ ��Q��M;��|�ayZ�p��͋f�O8sAbʹOQ"�)k�8#�.�ŭԁt+�d����� ����3Y�V9��̷IU*�1��<�t��S܅pcmS�Q����?|L~�Pb�U�.ߺO���$�*S[�}��U����oIH.��۷
$��"˝7i.,xᓣF(�,M"U��3.��I��BB8;f6-^%K��0fֺl�Dh�b��	Q�'�<+��r4CÎ8ɼ�b�@�`X�S 5; ��L�(S�4�H�t> ��i�A+EJ�f�l�ƯO�K9:%*ED�cV���lb����4�R QBNA F�'���9��P�	�D�C�	M��H�#��%��)��4��hɔ�	&};��mڢd6�aF�-�j��O��>.�&�
(o�)c0L��j,��a]��<A��(I*�pʡC�O�D9#�39j���.�v ��ze��8�8pc�F��M���D�[�x��2���nnؠ�'�Nԛ5J��*t�Y�f ͈����8���Z��H<�@�_���HV�?)���-|"��'of�!��A�aH�U#3`͠>�h
E�߂X6|�s 	�52���!�?�E�G>��I M�?�l
�{R,�^�2)�F��&�nݸ���3�"d���'�!�׏=}ưkSl��]�*�� ��uWcΞ3�^c���	tC_?�V,dV�(d�mP��A4���S��@Cd��� 3�����߾|�)��ɭA�|1#�
I���;Q�Q�'Ӑ�:�� �6��l>!�js[�X���F2O�xfH�YFr��pÉ�QخE���'Gv�� c��P��䛀2��.�=Y{R�Y!��.	&� �Ё�(������B�0��T 1GX�|�f��.,Ѹ�bfh29Hg�f̓fj61XG�<�d��6���M�&s��!�2ĸ#*�*C�yz������[�P!�VI�4�ڒ�:z}L�E���%h^���~r�B��U%�@�0fȢ5mM�*a!���P|�ᒒ!��P�)��؎-S!�G=@U��HS,��;<e*���23!�$�I��h teňo�$m�G�|9!��_9�y����/*�(�AE�'!���k��%R��u��s3DT	o!��@�Z���� �0I"����!�Y�α+�������ɲTp!��3W�R�R2nL�#d�@X��	_h!�
k*H豴�Ք8L;r���!�DKH�D���{j�yr*[p!��""*� ����4X�{�jE *�!�D+F'��s�O�� �n�k2)V#!��
0���7�T�p�~"C���<�!�$�#^��
B��
���BӢ��!�D�FV��2�*D=M0�,�g�v6!��:Jv���-?ZXV�gr!���-!�
Hi����2���3"O�]pf��34���R���2�"Ov�rʋdѺ�x	y�l��"O6e�%~4B��_,+$I"O��1��U��i{��e�Ð"O� VȂU���U����*['`~�d��"O�D�u�7|�TY� _�FSFq�"O�P���\�� {%�3?E<e�a"O��X�IT-�����^2����"O,,�q��I&�LzdK��\��"OP���!Y�3�V�B#�$B��q;�"O�h��	**���G�9�"OT����V-s�hu�eO�  Ny��"O�
Mn�B4cđ��QSS/D;m!�6R;E�aGK�n��pS1��"r!�d�
���sӴ�,��m!��֏|Ӽ�X ��K�j4���3�!��Q�~Y8�v �d�"̺��6-j!�R0|-�$�R&�?�@�IvÀ�MI!��?�����I�E#�ɹ��H�B�!���Cl��C�g,
`Y��S�!򄛥fqH��]:)�5�h �!�Da�>�AECޛhͰ��!�!��P2)��h�oΥ�t�?y�!�
�I�a1�Ŋ�^<|ò��(�!�$H�{���`�܀1����ߑZ�!�+R���T��,5n��Bo�v�!��U<9�X��934��3��)�!�D�#��HH���W� uar��/�!��H�z���S�X5�����!�D��:nH�f��	r`���
{�!�ߕ�A�.�?�Z����M�!����.�����ȋ-}�!�G�/��@�`�ɨo�葹�i"�!�?^�B��̈)Ƙ�XRS�|�!��o�:H���L�=/���>+!�ڟa�1��EԪ,�QTo!�!��G3p�~�!��1X�5т�9@c!� �����6_������-x!�dL�+�)�O���w#C�$X!��8&Y��0$��-���V���!�"&(r����S
zM��^~'!�DY�qF��c�˅$����!� !��WsA��
�*��m t��P!B��!�D "H9j�Łub��s�� �!�]�RC�8�ₓ�n�f̓���Z�!�d�.�M�%Aڎ\�5�SC[ t�!�,8�ғÀ!�
�g�
�!�D� ���;P�:/��2A`��L�!�d��yE� ��j�[���+5Y*G�!��n�`i0���Rժ��KV�R�!�X=S�M��M1?�-�6KB={�!�$E�y&꨸��O���h�2�PyB�TL"=C� >BV�ƙ:�y"�|����ƥ��GPr�Bӭƻ�yrH̅c�AK[E�0�놋&#�B�I#iL a#��T@�V	x�A�n�B��e�v���i�8�>}��KzB�5+�paAɛ��ԔC3	��@� B�RƜ�B@Z;~��S�`L8,�DC䉴n�����.��AI4` @�M�-j^C�ɱ:1*s'H�l�v�'�K�
$C�Ɉ7zʼ��ɛ�|�8l@C�8��c�HȮuC��`�呲BZC�ɡX���9u�
1H:HL��o��C䉯0�v|���J:�9��׵)�*B�� &8�<�'ꖌ= �9G�Q�ErB�IFb��r3�N���WHȑ/�JB�ɝզ�A� #��9�A�?�
B�)� ����@Ur%���̴<����0"O@0�bM��$�
�s��� ���"OX$���S\��(!�>*��R"O�� O�H�))6m�Bjl3d"OP�X %�C���c��r&؄�`"O؝ŉ�%+���,
�^�^t�"ODp"S
��&�%�*�L��A"O^���Ĝ�)��`i^4K�)�*O�DYEl��9H�4��A�#�'�pp��j,u��s�e�B%�
�'͔��iƜTJ��K<XLj�
�'�:<B��]�\�H���#�^9�m�	�'�X3g	?�B- v Q���	�'�vM[�/Ir�|u��O�U�x)3�'a�勱�� ?²УጘO,�[�'�J	�炱@�D��2��>;���'�}3�aƱj�zX��>+*�z�'�܉��,TMJT���P�]��'���eZ'8"I�MŪP<\K
�'����� ��l��૛?O- �a
�'q}1&��{zH��Èx�@0�'����quN@���w� !�'�=���ݼyk�,�2 \�[���'@~���^�h�D� ��Ӑ���'�\�����m�n sb�i�T�R
�'Ԙ@ �V�&w��ZscO f4�@	�'s��h0�
*q|y겈@Q<lAA	�'�n=WdC�jFP���H�4J�Jq��'=��y����Z�,�.C�0�0	�'�m��'��(r`�Z4(>4���'D�-�Ӣ�a3\)@��ҀY���h�'�0�����m�Ri�!.��_A01��'J������P�:��1ꃢQ��x+�'8x}��J�'�<a@�D�Kh�@	�'/�i�9��]��ܘ~l�iZ�+&D�Pa�"��/TY�P�4Q�Y���$D�xp!(�s�|���Y�f�HL�e.D�pz�̔4"�	Y�│+� Kw�0D���A�RFz4�;V�1Z!�$D�h�R	����:tדC�hU��n/D���&��]�9�Vi�;e�^��� +D�h��Ǒ�#��L{��F�{	<��u�&D��a\&8�U�uH��ux���'D� ذ�޾_�D�8s���4��D���"D�|$FDH��
Q"Z��<0�i#D�`�Ƕ��;��qqn���'4D��3$E�jf%+r��7iC�2D�$�M��X�`\Hd�?�aðG-D�0r�@�yۮ e��nUu+��+D����$Q ?˦	�@	M�X!�,QÄ:D�\�4�F��<)��	F:�<���8D�8��S<\G҉���a�O6D�THF���*�Ĺk$ R.PB<X3��+D�dY�_+yy�LX/ 7Ԣ�6A4D������<� ��#��"~NH��.5D�����Cl~�x�9^�p�9�7D�h
'�/;���%N�8BryW�5D�xi�)�=]�t�)@(�4YJp12D�8x��E#F��!5(�*C��@1�<D���1H� ���j׸C3�ŊL8D�|H$Wz�@�A�&׈��d�*D�T8!
]��r��L�*K��W�>D�|i�ІPt�(��<a5!{e?D�8���_H�8钖��(���"6�+D�� ����=iSLD�3a��"��H$�|"!�#�����	96H|sV�0Z�Fʔ�"c�4J�J�
��	9F
T�؟.M�pgF|1b��U�i�MQ�ƫ��)��1���q*�2�n���� 4�� ��î���(d���ٟZ|�(� �j�B�Bv�O}����� �����!hF�-{ȃ�qP� !O�1�qI5dGT0����#w�9r�>#�H{6d2h$jyr2�� 0r���iӂ�p��OF���Ol�A3ճ^5��Ȃf�OM�!*��'�b��1EL4p��L�	�:n�}��A�r��T�ǭ"`2v|�%A�^d�
׼i��	��ǍJ�,�ቐ��kd&͙=�f��`)	4`*Oٸ�ASn�@ �c�Ys�Q�[(��2�,��,L��!$W.G"�U��W2$Ѫ���@v���1n�
	l�xxs� 6�",���П��fʆ�0�`{���1o�,iӎ��o�|h[s��6�<�ݻG�H	��f��`u~�.M���C≵P�}s���;�n����  <�9� [4Q�zd�#��#}�>s����!ڨI?��Q�'M�-` 	L3ݦ�p��#�J�؄�[%
��Tx�l�mX����	�Orщ��'慃��81�Q��X��l$��"C�H��f�4�t�bXG�ZpHvI��tj�Aa��I�L&@�8�-]:\m���۸.!O� ��6r[H,����s�KP���	Ģ>�F�*�ʋ	H���E�HC�q�����P����A�n\���	)L���J�it�Y3�烊�R��ᴟL�o�?T���O���c� �8�)�#AZ.�n��,���&�rTc��!򄓕8>�MBd*r�" @�]x8Q�ã_���Dсx��вsi���	"�n������Q%/����ݡ7�^�w}cw"O0!�d�Y/_~�Qv�\P�i�
��M����%�>��5�gyrE �*�����H�{8�Yz����yr�1'96�#�5i���rژI�[���jX��W~�|�1
��#�p�P	��Q扄�I�$� |R�m��{ �$�-e�0)-Q�Ul���m۞q�!���;u�(��2�ĝ&W ���
A��Cg����DI/\H0"�G];��	\�� ���Э��K�9%H���E��-=����%�'I��C�,<��Dռ\�F�+��N-�ѨA��3�IE�G��r�fh!3�� �L���?���L@<@�}z�Y)Z<�����$�$�3P�v\	!�	�?ᡧ�=L(�-e��R��e*ف�>�yG �q��q��"���X0O��r
�AWj�q�@�K�f`������*��h(W큦��Ot\��"	^I4��V �Y��,;�Ň� F7m	�u��2'���@u,�;��	1��98B�I�!Ȯ,a��ڈ��q��� }�j�K Q����rc��yr'�"pɛ$J7�2�i><J�kt�Y�#@��VMQ�N�>���ՀJh!���'��a�玘�6�����c߾�pM)"�DQC'T22|n���2���i�N�����p���QA^�<!"��X%�)� D*Βh��� r�V9���iB�fF2�9 p��c�Һ�0��98,�^1ܖ$k�lG�H��i0V�W���-ɲg�t��$ <����S�l� ��H���c��O���VI�-k���Ƞ+�����ؓ�ؙn��[!#16��;w�NTKE�ʳw�>T����J(�����~�{��B�:��G!��t`c闺D���)D�`�qPK��5�t�C�4>�dq�7
n�Q쩈P���Y�Gl�'pf���$�r�&���@���XW�1;���C�D���͆� �Jţ5%_�d(D��:�`�B�'Y����^��ѻ�cתc~�X��y�#W�b|�\�'l`<kg��O�2�2T�  �'W�w��iڵN���Ӊ��Px�"����ٸ�%Ҿ̴�S@���O3u�@�~��!���tܺ�5�ƕ17�SB�<y���/(u@�e@�5�$O�Q�<��+�5BXkG��(Cd�C��A�<�V�׶���O_�>���d�d�<��G?J���fJ�p�s7cFI�<��H�>?�|���
��I�؜ʐ@�E�< �ڞ=��C7��-��;�)^�<vNÞmuj`[���HR� ��K�_�<�V@E��R9`u	X#l�h�)��C}�<�F囗^.��Y`i���	�B�A�<���M&.iZUAӛ&#,5p*�V�<�F��07��r ��(�| ЦIV�<��"�	X�$%��J�>hj��B�V�<!���S#�<�`��-\���A�F�<�/�>�V���*o5��*g~�<ɡQB�I�f^+4���iԦ�u�<��a�4>PvܻэF"~Ǩ����v�<���RI�DA1.���(6�
r�<� �􀓥��^Pqˁ&��(g"O~�;p
(�x�k7j	j2�L�E"Oܼ��J�'���B+�S�@�"Od�I��މ��CT%�3���p"Of ������c�4C�"O��9w��'�е��̀Ƣ�á"Or�d)�!�I
��ڹVB��S1"OxAbe�+xlT�pо�Le�"O^P�t�� ]dN�n��ȸ�)P"Od�����@��	WB�$p��e��"O�X1R��:p�Bg����L8�"OxN�eO>|��H��,���"OFT��
ˢv���C��=W�Z��&"Ot�#�
^�i�zq��%�Vm� "O`�+��M3z%�y#�R��pyU"OV�2�)�83Jy������u�4"O����H�/i�����ԺE�e�7"O�u�-̙n���Y�V�
e*"Oġ�ÑF��d���ա*��lQ2"O�AB���$/^����]pCw"O�xC�,�_�@�y ��Q��"O�4+6HK;jf�tLp����B"Ov@2T�^4Ddqm�0�����"OĘ���0Pj�e�`-	��P�5"O��X����ry�=H
�[��,�"OdM:��ߓ.!�mȑ�ȝGr8��"OJ��D��4�l�� - v`��"OX����<A(ٱ�o�4|,z"O�XIm��	b�Ы�(�gT��"O�Q���	
6)�6�V1>@I�"Om�� �X[R%A�Ȅ*.tS�"O��!F�`m ���g�4�Ɲ�!"OJ���l�B{�X
�݌7N����"O��P����ъz�(Wa�`�K�"OlYÓM�)}b���d��ݒ�� "O���QZ�%�H衷��E���1"O��{��@�Q��\�X�b"O>�`�m�E�Rm#E)�,�i�"OЕ;��A-!�`$��5����P"O��s����"��`s ��"Ox���
�a��5��"�>x��ɻ�"O���2�MR�}�PC�-mĚ�S�"O��pwAE2*��jw�ǭ*�����"O����m��W�� �B����"O�AK�X+ ���K(b�0��V"OX�r֠F�uk�d��@��
�|��"O���6n��z��p�Uۍ^��R�"O�@"Ec�/\R\���Q��(�"Oj8�1�IIi�`�WK^�r4iy�"O�Y�/�-_}�eDX�M��� �'�4	�eҐ� ��((2M�'�T�[���1A�<�J�@Q#D�L�c�'�f��&�F(�U`ajзl���'� :棕q��ܰP�ׄYP�Y��'�D����˫;<t�a�K1HC�Ip�n-Ӏ(+�2�c�lC:�BC�����\#n	2Y'�$�B�ۤ�Z�-�/*|1�m��`.C�ɇO���� ��*��4@څQ��C�	@�@Iz���3���Z���n��C����|*dI7;��t(�cY{��C�8B�@P��7$w��[��5��C�	w�"� �.3[�th�F
R��C䉣V��2kI�w�m�F��}�C�)� F �dV�a��H��L�z^�!k�"O��"*C�O������?51ڤ"Oj���E^�
4�|����=��:�"O!��1xU�� ��rZ.%"*O� ��ᅛ&�tZ�)W�J:���'+*Dc��^%k
�h���/B.���'�@� PKU��$d��Y<���'jrc��Þ|�J0�F�)"y��'���3(�
���h!%�ZE.���'r�h+D���;1V� 5��r ��
�'���SՈ�f�"�"��
iFA�'���zP�Q2X�m���AP�Q�'�ܫS��B��i�D^�I_>���'��
�ˏ�|P�J���S>����',�գDJϠu�(���!LAx	��'�U�@-S�VĵP��$;�XiK�'���p���\�b8��l ܬ��'Yt<�"	ډ7���օ �w5��*�':�dr'�z��(VL�)y$*�p�'�B	"�(
�\}�h˝瞑�
�'W6ѹ����@y���ӡ���B	�'���	)��b�����/{Kv)k	�'-�p�B�l��Y"����iE���'GlaGM�C-(�U�i��U��T(�1�7L�4�C��ҥ~���K`�	K������4� @����<�$C�73:�y@A��c�d]�������ԹM�4eS��Ύx��y�>���g��ħ=H\�P5��LrU[#�	jN�'�ࢦf.���|rre�S��$y��6����j�P�ʩb4�dl��L��%�ܪFR^UH��O��-���ԤV Y��J�T`ʳ院�NI"q�@U�bt��蟈�įK�	�咦��j�����L��0� ��i�����0|ZV@�C��h�sc��_7���q��e�-9�+�f?�,�{nd��)V X������vH����%S�F�`nZ���]��.	���`B¨8�LȲ�g��9ᶂ-t��x���� ,*��yF�ߓn*��JW;Oa�t��YA^*�ňD�\ � G�8h�%��%?Ia�q�a��ח;��4�g���|u�gƎ��yDU�)g�@���U��<(��ڮ�y�O�r �Qزc(h���#��y�DB�-T�$��ι
�^�����y��<rT�!�܏x�~��!����y�C��F8��8E�6��+����9�S�O����@I@23d!@:[_|���'3���i��B�$�$�G��
q��'�4	�)�@[@@
�,+�BJ�'Fl�)T��p����eG����0�'=��𧩌�e����C�3�!��'k�q"$a�Q��a1'�!�5�'�f�����%�	� �
�2��Q�'�&e��n^2hĨ�:U�'��y�'����υM$ƈ�G���r�'��x�L͛-t�]�1O�%<i�'��	����11^:`)��Z� ]���'�v=���633fq�dK��'��� ��'����7o �PBR��	�'�,��*�t�zw�W�0��	�'�Ȁ#��7Tf@�SmL)1�΁�	�'��t�4�K�P!m��툩q�����'9����a6�2�11�ɐV�Z���'��A1�J`y^ ����T�V���'��i!4o$tzJ�0 	F؎���'��v��$;��U�'�ѧDo��P�'|d] ���6+� �C�+����'��I3��cIf\`u+�3�X)�
�'�vup��2.�R�2������  �!ਈ�/3艻�c�]DF%k"O�,Ҕ�J����QC� 53����"O< �HǂlX���Ѡը[)��`�"OX�ѣ�k*xx����yY�"O�d9'�ܚw�"�B�,A���"O��U͞[�<1뀱5����1"ONE�5� �xT	ny�I
F"O����a�v�PH$ȅ%=��ȃ�"OY�bN�-M;�511��&S�H,�"OH��˒�d+��`��\���D*"O���s*V$9ܼ��D�I�X�ʉ`"O�Xyӆ@�yJ���B?�N�J�"On ���#r������r�6�Y"O�Ɂ��sNN(@�H�ݰ��7"O��3-�3@��#��I�y��\��"Oj�r	F��q/� h��`�&"Of�H��ʑ33���.�=X{m�4"O�p�'/]�]^�m�R��J B"O�]"��� ��A��l�8yg2;�"O����?�V����6L93"ObD�c�� vµ���ֵ@�] "O6"��Y�{B�e��AI�qr|w"Oz�hlZRȢ!�e@-k��k�"O$=@�.#�8r��  "�Y"O�z`��{�贫�̀�g�J���"O��ѣ.��3gf@����"OhJe!Z$tr��c��!�hq�"Oؕ���#5�IL�!���"O��y���8XY(P�P��2����"ON�9'�K�V��,`R&�<N�=�"O� ����gr��j�'m��k��!��~�����nhQ���ѦtN��ȓ[��yA傆0���S!�&�����_�����"�����S��p��A0��%'_:P�ER���#���`�Zg቉V���Q�i��p�x��A2����J+V�v聳I�K.0���gl�ٰ��%g>�cg̔GI���h�:�Έ�G�VA�b���I��w���e�*fId1"§�:&U�5��N�n�3� �&a�2ɢ���[����Q��b�Q���I�o�<y�ȓ]=�� ȗBa�	q�$V�9����ȓJ��;�&��N����^�@��]�ep��a�Ȁ�]�j��a��FVH�%(�>`�X8�64�n,�ȓ|B)b�K�&�<�IU��X�D5��W�f�A.N�f�)�6?�4Y����L�x.Ե���0n��ȇ�b���Sn�?Ch�ԈW�cy�]�ȓP�;3��&�h9j�֧)A^L�ȓf��P��F�a��t��5�T�ȓXzx�h�J+���a(U������!X�Ur�d�u����~�L��8<`#uċh�*j۴
�j���\����6$ρg4M�$%�J�ꁆȓVSh r"U� �V���N�V�8��ȓnRj�KrEٺ�8���Z �ȓo�,Y�s��9ǒ�ˁ��>n�H���]���֢H�j�����lɽP�ڼ�ȓ?�e���g��)�ֳ\��T�ȓQT��!�J�n���S�^P��K�t(�pEͷW��1 �!H�$E�x�ȓRc��(�N�;$`���^�jх�S�? ���gdkw�2�P�tTD͙�"O>�I#��YpwG|8L0��"O�p��#�xtk0���{1ҁa�"O�hTNM���hD�SN`s"O��a��Ϡ#����C�=��e��"Ont�0 �D8� "ƒD����5"O��[4n��"�F�P�H�4u &"Ott�K�/F����ʛ�h,˦"O�����[:^n*�	M�@�=��"O�M�ᇛ�A��|3���
�^�� "O�!��C1V[�X�H�/g�ݸB"Ohy;Rc�h@L���FQ� af��"O�H4�I�_�F*�N�=`.A"Of�ڣ��Rb.k��@lG.i�%"OX;�N0��- ӄY��B"O�]�2(]��Тd֣A�4�
�"O��˱�N,���!����,��7"O�Y�Q��֤�b%�$�L��"O�����Q�9�ҡ�� �X��"O��1Pc̦.�lkAT%7iNA��"OZ ��ݸ0�����'RKf�xV"O���jU11����T/��A0�x�"O�h�p�02�&L�#ɖ$<8�&"O:uP��o�m�.	�x�(�"O�;f
 �/��]�c�Go�rt"�"Oޭ�`LM7}�lC�JE?��m 5"Oeڐ!_	dzi�`i��B�x�w"Oj�:R(W&k�f�H�(G�AhV�!d"OFYzE�-t�d�g�;DQ��G"O���r�F=zh�"lG#=ܫV"OX�� ��*\cP�5� C|I"O���GN�$���u(�|�8"O��J��H(j �c�οs��%��"O��i���+v�XE�N���AW"O��gä6K��ڠ,;�.�#"OHXs�h]=^:���#iۿ��xR"O4L�a��(���Ć\�F�s�"O^�)�/�#$�,U��/�2B��ؑ�"OJI�1�B6^INܑ�m=!��;C"OD�j�e��s�f|{�L�G|�$�"OL�R5n��0� ��3|��bW"O�԰�8l$ ��B!a�.��"O<�C�+Ux�a����<F�D�z$"O����T>� �ҥ˕�yo�,+�"Od *��R�6A��´PnA9�"O��a�����8�R��٩qV�E��"OV�
��q�^��3h��Z���q"O$� ���c��G�y��x3�"O��U�ĵb,^�U��(2�T�s�"O�cjɼ|8l���՗W�dhv"O�8��V,g��I5�Otq�s�"Oq'F�6Mh�1���C�r���"O�@ 5��:p`��ц&P��X�"O�,*�B�792��1��بF.��#'"O��{��Jzs(K�n��yplAq`"O�A�CJͯ �;�nZ3FF���"OZ�a�E��9n\���deZA
�"OX��gM�He�	 �=n��"O���w�Q,�Yғ)�\� �#Q"O�0
&�<=�X�UiH�X�t�p"Oju�C�n����HD;?#F��"O�)��H�+2���ȼk 
��"Ohj[�.|����3)���"O>���].5��2�.40튑"O� �ŉ���1yw�� #O(j�"O�@��@؜M"(��.H�'0i)U"O���6b�~,��r ��.v�kW"O.dR���R-;u/Ph�T"O2��7/B&U�1�t�\9r���jF"O쁣`�
�L9�E���
oz���"OP�W��0����4o��Td�ՠ�"O�t���͍0�A�dl&+QraZ""O⽉���mT �t̂�=B��D"O���EA}>��&��	{��܆�_w8��uj�=�q����<A���ȓM<�0à'�k}f��Ө@�>y�ȓ5��p��� g�*|�uI��N�ȓa�6u��n¶Ƕ�3���F�,�ȓU�8t�d�-,^�K��E��^���6qЭ�򄗷<�p��a�6�&�����L�#� #�mc����/�i�ʓH� G@�%`��� ���+dC�ɗk���FN�+J�����U^\C�I�@�& BJ��D��q���#r�XC�	�V(�ck�x��m����U��C�I�DeD	e�#YI�ips@ScY�C�Ih\�X��^�X�ဲLQ.�jB�9d��(�SFR% ��iT�.)��C�,vO�,�V�
�fS�)�7r&B��??l8uG�#q��U��AX��DC�	>�L��N� �U�!��u�TC�&;dB-������e����p�C�		Q��٪���V�<Es�k�� C�IAv��L��I�:Q�bc �B�	$<h��#T�
�Om`ѹ6eY�-�B�	�[c�U��׆]�$E��?�B� DD�c��D��-�
M�K�"O���C�w���S,�7��� "O���	ί3ΰU��ζd���"O8��D�B�#*�Es�KR$*���S"O`��$��T!�UpD
��<�&��"OR4cc��y�´sg'̤i�p���"O���wH��n�n5A%J�O���3$"O4%!��O�l9� ��A�3d��1i�"O�:�.�z��:��_/��h0 "O��KZ�x4�Өs7*��"O�|3�=�,��!���m;�"OP�"���:7>qpH]�����"O>�X�D3p��$*7	϶f�,���"O1ɡ熖y|R��P�b����"O(����̂9&��a�$���"O$���˙�FV���e��5>�M�2"Od��pĎ���$��K� ����"O�ͫ��+�hI��� e��"O$q+%g�$Ƽ�^-��mk5"Oz ��NYs�@�h��"J�;F"O$l��,/^��[*�S"O��S   ��     �  d  �  �+  �6  eB  ~M  �W  `  �k  Qv  �|  ��  N�  ��  ҕ  �  Y�  ��  ܮ  %�  s�  ��  �  J�  ��  ��  ��  m�  ��  ��  � � ! �/ �9 6@ xF �L N  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|`I!'G#\���%�T��'ItcbꀀK<�k��̥:O��'������Ǝ8�ݓ���"J�S�'y`=c �d���	%�BPiV��o�<)E�I�M��c�Q'��I���k�<Yb�`��s4��/~�����M�e�<Կ��رD�E�?�t�Жgd�<��j�aZ����Aّ'�F�r�b�<��"���e�ďfe��ѣ
�[�<Y �{�<Ԑ�[�0�Rѳ6aE|�<�ǆȕP�,x��H�o���ۀj|�<��\��!G	��lhP�qI}�<�cێ�,����ޣ��@�#��x��G�<��Fъ��u��Z�JQK�%v.1���� ׋� ^:�Bэ]lr"�&���I�-4��Bbʴ9[��g.A�$&��$@?�vĥn9zt�&D��v�����Z�<�5��@e�
I
p%j�a�L�'�Q?y[��Ph�d:�
�Z�bg/D�$2��q�HÄG��R����I�r�����䕘!��8r@�P�Fi�	� ��!��̲��u*4%#\l􁦪��,�du����	�j�����
���k�h�7EB���˃���.*����u$ML�BQ���C���C�I
|����d�2�y�e#Q�B�	�� R��g� �t��B��1�s�Ee� "<E��'�����?l�i�|����y2�6�Şw}��̞�� `�d�ǁ���a����dE�D��p�i^�;>��S��%+�|�L3}2jN,m��+�lRu��iT�y���>�����Q�g�عQ� ��Mˌ��%��|ph�9IV��1�!�;qu��UA؞X$�>�XR��V�ԎPԜa�g��:]&���d(8a�МA��řcYx�h�G��%ڧ\�ƠB�!3]��`��G�44��^�Ȅ�-J�S�d�Ӱ%�'
<�'Bў��$��Fa�,ʕ0�i�9j.!�$�!i�;��@�f�I�Iſ+� �牰D�-�Dk�;�Q���c�C�	;<�4Qd �
����'�4��'��Bm_�K;�HاA�H5���|�����Hȸ-&�tbr�Žp#��v�/�yb(Ͱ6��9�L��o�(��^��~�!�S�Oaƙ�gh�[8|`c��e��e�'% �;?ʡ��� J���
�'��s0i�3y�Bd˖��Vy~9�	�'�F��A�^_8@�D_�M}F��'����7�[�Y��:C��JF���'�*ex��N�d�B��9;� b�''��SѪԮ4	�#"K��7cL�8�'����d �el�0J�g#����'�HS��Q��*�р�	����'a�|@0l�9�0�p�A|�`<��'/x2���93�]���:%���`�'W��P��҈4�����)뎨2�'R2K����y(J�0�D�Z"m��'�~���j�$)ԡIg�0����G��O����^�E�� �9rdx05$?��{rɚ��I�m#��Q��Lm��$*Ǹu��ʉyr�'q�x��H��t��ѯ���r�H0ND$��=�3U����"��M�霂���.�69���ȓAR�L��/�B��ǭ��-����=���?Q��Ӟ6 ʝ)��^�%x"T�&��~�<Y���7?=f` ���4~D|9qM{�<����J�Fa@o�`Ѡ�sS�Q�<�[y|�d[� r:���`n�EB�`�'F�|�ڮe��)҅��F��b�O���	^���O(���b�>�bI����O��p�	�'eF�Js��#y��L�Ǆ�U�
yK�}�x�鉷4��9{�ɐkL����N4Z�rB�IlZ6�+l�	<�ؽ���Pdֵ����'] �cV�`����jG�%��9�'jX-���_�"�ba던�Da	�'�bY��R&��l�� ���$��˓�(O��5,��N�R$�7/T�j�~�J#"O�BS�]9af�K��G�Y;b�s���=lO�A��ydVEk��ה:0��"Oȑd<$�X���$Υ|����"O���t.R9ǎM�1���S
nj`"O�:AJ���,������eh�ha�"O\�!��שn=Ҍ��$�	'�<Y
�"O��#@E�U��C��W�9���"O�؀�J��}:5��k
:�P��"O�D�G@فE5ZA�Cj`D����7O���df��	Y0i؀}�~��)I�5,�,���'���ɉi����AE\���z�&I����5�I�|9������?& �S &�T|�B�	���0p#� ��� �<}��B�I�Jz��5B�% dY��T�A�6�F������ ��A��ƛRTV�BpH�>���6"OL�ke�I�Z t�A��V)(��2dU�p���h��Q#w��
T�� s!�F�H�ZC�I,A:� Iv�CQ��2�iħX+`B�8P��(��_�!�l�s�H�3
R>B�I�T=dX�!��N�ZAz���._B�	,$��rVk[	l��-q-�)
B�I�e|Lru���Z%��� $��>r�C�	0����ThW]jP��-B�6Z��#��c%O�>�ȉ0�F.`�����4�O��$�QԅƪuJ�AK����>���0ƈ3D���� 	F��AƂ�5�a �M2扃5���?�|b���b�c��$��iIGhd�<�0�� T�4+	I����a�`�'O�yB	Q�$�� ��>;L@�cc/_1�y��%&�&aYF.đ-�E �Ј�y�C���v�Pg:��P�7J<�y�n 'Ǻӑ%�0�؍qbC��y�ώ?~�Pt,(t������	�?����v\8���,�H�Pu��!i|���ȓ@��-Ӥ@+n�P�Sd݃B�v,	��O�����!3��q9�(��D���fcҖ^����)"?��,�;�2%��۷�����(�f�<���H��z�eZ�j�
1I�<��l����v����¡К3^lm��	�!n��M{�O��e�k�!�"��"bN؜�"O$Iǣ�W�$�����w���S��D�O��s�{����P=j��1���{�|x{V�D˟̄U24�K4�ҔT�X��CDP�(��:g(I�&�ݱ*�������>�rԇ�,�*I�K�J��f�3��!�ȓ%�M�adT/J�������n4�ȓ�Jt�0o�zB]��j�b���^=�P������[Ôpc���ȓSܐ�bɇ,�����ODN�ȓ&��MJ�� m=j�%)F@�م� �]Y�Fѫp'T�C��J�[@�ȓ?�,�B&@�����1FTl��b3�Y��N��z�	d�.n�B�ȓ9����[��䪧(Ų!xPl�ȓI�@��Q�(]�r�I�Z<��O6�dұk������@�]�(��׈��H $��<1ѧԗk����n�hU�ݢh"69YŨ�<�\�ȓ[�p�Q��L�r��a��_p&ȇȓq_Mb�o˗%�@$�+�# �����<_p�+3
�h�F@�3$����@ua���7���9�'A.S�\�ȓ:����<%�.��P)��(����|��6�Ѯ#���ޠg��=�ȓ-�E�� '��ߓ4�� �ȓ"cr�@�0!{�	�fΈ�
@�T�ȓu+�,J�$��P	�)+vN6Utz��0܅�P/ٮr�\��v!�h��x�ȓ^��`�$5)x,�N8�f�ȓz� 8��O�]1l�RT"�39���ȓ{/������-��$~(�ȓi<ش!ĭ�_<"c/ק!а�ȓi�Y�&T�w�^��n�%4P��ȓ*�f�K�JB�$
��R�ĩ�ȓx?�W� ❩3 �.��\��`�Y Th.���)˯vD�ȓM��R��+�:v�Փ"6E�ȓz #U�$ut�A��7-�4q��S�? ���*E��t��Ś���(&"O�"&H�8��U��e)���u"OnQ�A��r<x�D+^�@:8�W"O�h��&Y���k��N+/���"Ob�p����U ro[�[Ά�[��'��'��'��'&R�'�R�'Ӡ���J<OT���ʗ/p�4���'���'t��'�"�'A"�'�"�'�4�Q*J�$BLc񧆈aR��!��'�"�'HR�'��'42�' b�'���D��'�� �1�u�3�'��'���'���'���'���'h�v��k��<"#��>2\�E�$�'���'���'vB�'R�'E��'�Dm٣��"D*����Y�r<�f�'���'���'>r�'���'��'&����
���`}�&�ȐF.Jp��'/��'���'e�'1��'��'"�����5`�P� �R�F�RC�'Z��'{B�'>��'ub�'�r�'@����k5c@�A�*�-5������'���'�r�'e��'or�'���'��)�ը���e��Ȓ?'�=�F�'�B�'�2�'#B�'7��'���'_dQWhV gg�0S�M��˂�'���'%��'��'Q��'"�'���AЂ��t��!�,�W�'{��'�B�'���'���'+��'u�� coK==�vlz���f�R�*s�'���'��'���'R�a�����O�Ձ��	{����rrgjm(*O��D�<�|�'dv7��%{�l�ƀ�M�hX6�	W�~������ܴ�����'�B�3:*Ps��0vN�y`�*T��'����i;���|�6�O�'
,�=
p��m��#�ن.
��<)��� ڧL�`��.MZ�^�6�H�APP�iΞ�`�y"�I���[{�T�&Z�g���Y��ʢ���O*��~��ק�O2؜�%�ik�DB������0〉*!�
�q�K����=ͧ�?�S�*2C��F�6[~PR0�<)+On�O�hm��CX�c�`y�h=/7*��c�ޠ70>L{�aLV�A��	ퟀ���<��OP� ����.�y�&e#�����D�O��	b`�Kz1����KzR�d�7o��0Jϓ�܉ɥ���xN�˓���O?��.ht����'RUd���r�	8>��٦2կ,?Y�i��O�I[�f�Q�&R,RPX��K0 @��O����O����xӄ���$,����
"&�7Ȍ���Um��QPA�4����4��$�O����O����X��Q��I��b�)��\#��w���K8N[�	ҟ$?M�ɮZ��r�͌�\�$a֬$V�L�{�O��nZ2�M���x�O���OfЍ8\�i{ �	!�)~�(i8�g��{��M#�S�D�$�\s�Ҍ�^�IVyb��er�� `�J�x�6x�(���0>�&�i6��B"�'��xl)1��}0F���Jk$٦�'��6�8�I�����̦���4t���GZ6�Z���	�c��T�C�
�b���i`��O>U�w습��wa�<���>�k�0t���ȇ��8<]�R��ΖB$�D�O���O��d�O��$%���OrIb� �&~ž��ů!���`�O����O�nڹ_d��ߟ��	ß��'�^ #3N�0�nM��-Y�25�����e����'��7�ѦE�S�n�(o��<��U/l����L�T���0
)���2p	ƿ~���������4���$�O��䍳Y���Y���0!��dN�>�P�d�O(˓) ���,W��'���O(��JǸ�T@a䎡F����/�8�y2�'W�Iϟ�l��M�b��T�O݊��B�65*���S;Q=���u�ئ,Ɯ3���
�����n���H�OȄ��cO�
���j�'��`����Op�$�O,�d�O1���"���n�vC���f�T8m$�u��L�Jd��h�'���oӘ㟠 �O�9m��O�.iA�[#e�t��b�1q��ܴ3+�V��"u��6?O����
L�\=��'$�r�A\�ˀ� )��:�)3"V������O����Ot���O���|jdhǱfUu:℃�0/t1��[�V��։�2NEB�'����T�'ȴ7=��8D�P+
r�hQ��{���g'���-j
z�$��S�?�S��HmZ�<�&	(]%5��o�*��ٴ��<�U��3���D	��䓍�D�O���1+c�AbS�μ��x��.��|�I��4��џԕ'�7��"���d�O&�UK����e�1Z�Z��LK4ZV�d(�d�R}2�}�^	oZ*�ē0��y��P�A��1/[6
~���?a$L�/���J� �����$Z��_��D�$M۞�`����X��Gp�!�d ����@��Դ��.�����
��a+���۟ ��.�M��w����&l�"4�`��� �6.T�p�'"�7M�u�ش>QꔮX��D�Ol��ƀ��r�͏2%�CfL�
����,J�O��?���?����?���E)�pC���.��1���E�X��aH.O��oڦm-��I�`�I�?͕O�C� ��!��]�pw�=��削�M���i��7��^��?9��EV���"RB��q �D��e���؂?L��I����OB��K>�/OR��c�ܐ!ҋ�4(�0���'��7��$�Z�dKD~�Q�����U�%���M���d����?�!V�4�޴:6��cӐyA��.X��[0J� L�r� &��6rb�6�e���	��@��b�OB�T�'����k�� D�QR"�;&P���՛w��M��8O���dĚ\&A eÝ�AH*V�{@�$�O$�T¦�cF/RҾi��'(����#�4��t�MtZ���>��ۦyݴ��U
N��M+�'t��J�\m*`BV4p�
�j�I5B#���3���x�|"_�<�	쟀�	��t�S@�'/1&�;2�A�Q���7&�ǟ���jy��|��qB���OZ�$�O��'j5�pc�F0a���!J�bG)$?��Q��X�4Z1��-�4�.��ܯ-ՠ\����=�$x���G�|���s�Y$��)n�<��'w`�dO��?�)O�,A"���Z�Bu�B:h���$j�O��d�O���O��|2)O�HmZ�{Qh1t*5S& ����� 2���֟X�I���%�T�	vyHf��5�GLH�?���HhEZ��LҦ`�4 ���ٴ�y2��>bD��aj��?����:���27[^��E�Ǐ�TE�5�঱{�V���	矔��ӟ���Ɵ��O�R��kI�|B�h�(Q/z�f��Cv�ک��O���O:���dRʦ�]�,[���P�RH��i`�d�ڴO��b&��I\�<�7-`�dMA  ba��N\#o(Z�S�l�$ ����i�b��j��ny��'���P;���BU�Z�10��@�˻,*��'�B�'�剢�M�r������O�u����d����eN7v�H\�d=�I����Ҧ}
۴;މ'5�1�!�3+�����R�� ��'_���&�J�b�#t��?���'���	?�,�@d�J
2pa�/���Iğ���ٟ���J�O��5u�2t�5i��Yh�����:k\�`��[��'86m�O֒O��L;7�b��c�Q+E��!�'$�*��$����J�4LK��i��b꛶:O����l@���'�5�)��|�R��OԺH�f@�������>�3�5�7F��c�x$��+�n����'��7~����O���8�9*���!�\�d��,�vꂠ�JՂ�O�-o�*�Md�x�O2���O�j`��''�F��3焨9��1*���R�D�q^�B���L����q.�*� �2m�:S���a�I����e�6Ԉ������E��p�&�HpΉ�
� ����<_^Td!C`��X �C���y�P�S��G<�a(�5o!�|�0�ti
Y(V̞��B%�����]mڤǌ�;�T*`�n�I�^7#��D0M��}x��w��+%��� �؞J������i+���޲�	� 1k-��:�ŗ1�(P�Հve
@����]CDI�h��^F�acU'�p�<AH1�P$9���I%E1Xi*�'K"Ͱ�@��n$h�J6�D�*���L����P'P�P�E�1�W9pj=� ����?�H>����?�RHt}b��.�b 0f^>d�*��S�?��d�O��$�O��<`Xȋ���􋁉x�諶�B5yb���r�L.�7�OR�d�<����?�`C�ţq�Yy5��-ly��X�C�>LRr�{Ǹi���'��I-5���O|�����1H<z�F��wg��"b��moy�'��4��O���M�#��zJ����M8��@f"�¦=�'@����ddӎ)�OZ�O�@�e�,�f&L� (���N�*���oП����R.�����$�'��L<a&e��6<`<#���(�����C�㦥��;�M����?����2�x�O��gLD2]�.���n]�E�
��%o�f�Q�ϳ<���?!�g��?�'��?�ni�F�ְ/��h��
>r�6�'���'g��@).�4�L���O�`E��<��\��E4;���Lp}B�'."DIߘ'��'^�@�T<p#�M����a�0��(I��7�Oرs�Ax�i>���ßȗ'=h��OUZ@��"�"�`8xCBz���$&qB1O����O����<aĤ��{I����^1�L���3��=���x��'y��'��I���	�玙2F��kD��ʔLR��R�B�;�ߟ��	��ܕ'$�IBdu>5����KY�,$�4"%(�P��>����?9���d�O ��
/}+��$>��`�d�\'�&|�T�:� ��?���?i,O��V�D�S;6ȼ��"�"URН0ㆇ7�Ecݴ�?AL>�.O}�C�iB+�̓�_3��-I��̈G����'�rV�P��5�ħ�?!���P�գXs��c�6Z�KB�~v7��<����?!�Ŗ�?��U@�M�ֽ���s \3dzӞ˓S��s5�i���?Y�'#��	e�vH��k�g��(QU�.-"�7����'D	�E^���&���5�\#��؀R���:(��)u"w��v��צ��Iʟ��I�?1�J<�'��e��U�f��,�>2;@t���i���Z���I��3�	埔D�ڡIhW�;2�6��6$C.�M����?Y�k2`�ҝx�O�2�'�&)ʒL��:d]���>R�,,HTM�>���?��Gn̓�?����~2K���.�kHU0�>�sC�%�M��e��(O>���OV�"�;U��@��s�xG�4�0���g~"�'O�Z��I���@c*ߚ|��CE�A�w�t�	�Mpy��'�2�'��O�D;w�4�js��-B�b� X~l�a�I��I�����_yR�'�lt��ӟ��#���T�I��ȯ!�浂Z\(�	�����T���?V-�W��Doz%�+���8�mh���F2�eʮO ���O�˓�?��dD5��	�Oʕ�p�Q�3�HAJ2�P�>-Fԁ0�Ȧ��	m���?�bdN�="I'��;AI�H�� ��'{��R�EdӘ�İ<Q��r��,�����O*����U(>}`e��/xp�����<��y�>��P��nJz�S���Ɔm0D9�� /Ew�j���9���O��Z!h�O��D�O��d����Ӻ� bx��,�uN�pQW��8j��mPfZ���I�&(� A�<�)�S�~��;P.�;>�����(G6�7�\D���O���O��i�<�'�?	�,T�`�`��r���Q@�6⛦@J$3D���y����Oy��H�57��)�*�8��9�lJ�������h�I�I(�	�����'�"�Olq(�"^*A)�p���1?�J�$�x̓�����T�'U��OBH�b×<��H�a�[�r�~�{1�i��^�)/�ɟ �	ܟ��=aC-]�p�S�eV;(��W�>���9<SB0���(?9��?A+O�$����"l @P�KǊ��_�,�s��<	��?����'8R-�*��[�E���`lC�G�J��.@���Ol�ĸ<��g%j9��O�<@h4ϓ�+�X��B�����ٴ�?����?!�b�'�j����[��M���ռMP����@�On�]��
�E}��'��\���ɢG̖O��jމ�b<��o�
����C�6h��6M�O�����W(�ܫ�M-��I:`D�AꕽvV����ޙVZ�&�'�Iԟ,"#]I�D^�����t:��M�3�&�{w�F�t}:)C�}�^���t2�Ӻ�T�@Q�6��h´D�<�k`�V}����P������ßL�I�?	��u�S�	��m�P.J�
*�mrcZ���D�<!)�K��ħYD�����˅l��}ѕ���A>B`o�;{���	����'�tQ��ȟ�9!o�9*���xW�F�*� �)G�չ��$��b>!�	>*��0���͡S�H����$�,�+�4�?q,O���w)�<ͧ�?1���~R��*W�H hu�.DD�5	�D�./�`c�dR_��ħ�?����~Bg�<Op,��B�>7R�i��ǔ��M���O��LZ/O��D�O��d?�	'N��<a�o
U�H}HC��,\t�}��d��e~r�'��R�t�	(4e��)�mN <z1rAᎺ	�9���'�2�'�����O��Q�kR�R���,K���ksd�k��(:֖���I��`�'X��[#���
*a��TJ��ּg��I�=��'.��'��O^��5 
1@u�i? 
J�R�����d�/o�&S�O����O��?�T�����OR�C�h��1`�e�Fi��� J¦��Ir���?q
Wr;�X&���F���pAC���66CHQ�~Ӵ�ĳ<��-�l�+���d�O��	��$#��0@��N��4��BX%Nl�>�k�	�u-�~�S�Ĉ@9Q�e{�˝�)=F!{��ȸ���O�	�#��O����O����.�Ӻ��E�E+r���Z�T�{E�Gn}��'�z\�W������O_�))!�H,MV8��1+�*+���ݴ�a��?��?9����4�b��L�d�(<;�a�#8Oʠ��"�V�pn,CiZ���6�)�'�?���e����3���%b��z���m����՟����Vzy�O^"�'����	M�ƽr��5D80"��2D�e�<	��׳m��O��'���Q�"P�3-Dv#�R�@��&�'��!�_���	џ��I{�.[� ���}X��vk�U����'�Ե�����$�O��ī<!�k�d�@�J��� &-K�6t:@1b6���O��$�O$� �I4z؁02��04t00��s з\\��?������O�Qrl�?�![�x����]|s��Ђ'~Ӷ���O��d,�Iޟ��ī�!�7�C����)�joB��Dcχ�����vyb�'�x��G]>�����]0��)o\	������!m�� �?	�X*ĉ��@�-j�"�m@x�Y �d�n6-�O�ʓ�?ٗ@I��)�O�d�z�r�.�)e��+d'ϭrT��2��L쓸?�!�U'wXj�<�O iz����M,`L��V�R�:�Of��T�K���d�O&���+O�N��0Fܵ�w�ȠB�~4��Q�)��I���9�M[�8stc�b?�c0b8m�򎔞Z����t��`�P�OB�D�O&��럂��|�����/Y�EJ�
߰8�(���Mva�-7���<E���'��`�f��@R�hr�'D�¤k
h�L���O��DޗZ�b��|����?	�'x}:�����$i9���� qa�o(�I�"(l��I|����?��'�6���!��/�^	VgM�m����4�?Q�������Ox�d�O�➨)�<0}~�sNV�W["̒!�>فM�M|@�'R��'J���������� ������*��́
���Q�<��?)����'d�@� ' h@��<5*��a�_Hi�u
��>���O����<��'�*DB�OFn��4a�'@1R��R�iK���ݴ�?����?!�B�'�D	�ÍI.�M�^�ez��w��|���ʆ��j}��'�Y���	�,<�O����&v٢�$�[�s:�#��o�H7�O����	^q��a;��}AM��� ���f��4Sn�6�'����(��%�~���'���O��З#��br(+�Ҵ��dZŇ*������v��1/Ѹc��R�ti�:������U�'�".�M�R�'e��'���X��]
l��₨,HP^��nI+-��?1���
�ܥ�<�~�o�+��IC�L%4�j=�������s ���M����?!���&]�Ԗ'��`�ˁ(�� �p��<�`��WMi�rس��o�'�?���\�>@l�G��I<��� b$x��f�'�2�'E�􈄀�>�/OH�d��� �
�d��c��Uqv(���W�ib\�(
�r���?	��?��90�h��MS�`Ԓ h�-��V�'o1O�>�)O�d�<���{�hL!$�ܭ�ĂI=Fp��*c}����yB�'@��'���'%��noR�yT@F�a���� ª �d�S��%��$�<a����OT���Oh�C�搀eV��Q!$S�6�y��bKj1O����OB��<vQ�Y�)�.En<!b反�' �P�1`U�l�&X���IHy2�'���',���'����$I�@x�er#DB� ����jgӒ�$�O����O\�$���QQ?��	�$�V� $h]��F��r��)Q"��4�?�+OL�d�O��$��aG�IJ?	ǌ�VF����;`�Q����Ħ�I��P�'O��j�$�~����?��'ZR���'��n=� Kg%Y�	�r��_�t�	��H�Ɉ_ ���$�?��q/E -�H\���N���#A�{���S4t*�i���'�b�O���Ӻk��?A).2F%�.^�Ф��������P!g�ԗ'�"�I�I��C1�Wu*����ԛ�I�|�6��O����O����T}W���v�s�\��0�(e{D]��L�$�M���<!M>�����'�Q�v�F%&��"�N�?Ch!#�!eӄ���O��dB;Oeʩ�'&�ܟ��n�Zh�@+S�a�Ek��4HU�5l�K�I&v���)���?����10f�*�}�Aʐ�@<;��iB��*.$6�Ob���O��ćD���O��1��D	ij�8�FO��8�<��sY��"�g����ߟ���ßX��\yb��#�:)�)��8�(8i�MN��d;���>	.O���<���?��'���1��7B��)��fV�(��F��<y��?�����X�Y���ͧ$�Ɉ�mN8$�Ђ"Ɉ/!�0�m�`y�'U�����I̟`2��y��!�
Q� �s��T5a�@U�«߳�MK��?1���?q.O�]�w�Gp�T��5V��l��4�R����Z�O3�M�����O���O�XY7OV�'����N?2HV<kG���U����4�?����d�)y����O���'�����wn����c��aU�Sr�˼5�&득?���?��n��<�I>��O�<M���H�\U}�sa��$n���4���
� B�(m��h�	��������2�x���,T"�tF�p9�� C�i���'���<1K>��4�Pn�PT�d%O�s?&�{�'_��McR�Q
m����'�B�'�$"�>�/O�pKж(�ģ& T8~�Z��Q��ՠ�g����Ky2���OJmòE�3�Z����3*0<(�j����Iɟ��	+�X�ɭOZʓ�?��'.�3HYz�X���Q���y�4�?A+O�TI�<O�S���֟�3�BƮGb�9F�8$�"풢h�<�M����°T��'K�P���i�:�VZX���k� �����>q���<	���?1���?����D2|��,��̛u�&p��k�b}�Q���Igy��'ab�'2z	��L#[ux�Hu��hH�Z���6����O����O����<���Y����S��Uذ���)���0w�"Zܴ��D�O���?����?aӇ��<��8{�Y�HJ�a�`��C�}��`m������۟��I]y�F�v��맾?�1>R��U,]&|2t��$H�^/
Tmҟ�'@B�'I��Y9�yB�>�"+I�F�.���V� L<���Ҧ����Ж'y" �J�~����?I��,ix��e����I �Ӟ8[RT�QT��	��	�Ez�I@�	OJ��r��P)@Ϟ�LBhU�fNZϦ�'�n<��j���$�O�����*Uէu�4r{$���I̾(zM�0�
��M����?�4���<YtR?�	~�'f����AĘ6b�I� E�9v�elZ�ca*۴�?��?���=c�IJy��W�h�4<��)�Rtc�.{�6��?�:��͟h� �ؙl6��SF�����fW��Ms���?Y����*CV���'Sb�OZ09�3�E��_[̩z׻i�rV��k�y��'�?����?1Cӿ`�μyԇM�c����.ݗc���'�H� �c�>y.O|���<q��D��J'l[�L�0�S��V릁�I		�$�	ğ�������D�'�r���lŊ�D��NL�z�֠0�#.\5P�����OLʓ�?���?�eA�e�"D�e�I�p��Ä��S��͓�?���?����?�-O�`Q4�I�|⠂�;o����A%26��a��Dz�	�T'�D�I�0wm~��r�H=;�  k�26vQF�	����O���O��4����v��T�N���Dfة���"� p�~7m�O�O�D�O�m��D�Q�^�H�&�/�=4��-����'q�U��@D�֒�ħ�?���Y���d�D)b� l��*���q��x"�'T��\�b�|�ԟ��	E
ۖ����w�o2�hr�@�I�R�{��i�&�'�?���[��I��		�.V�seh��#*6m�O��D&&��#�D#�&|B��q��{#9\&ڨ�@�a����C�殮��ɟ��I�?u�M<�� !�ᢆBǟ?�*�4�ڂEP��q7�i��ۙ'��'���dy��'�Pdq���XU2�sD�-t6B�j�'q�H���O���G}l)�>���~r\+��Г��'6��a��-��' ����y��'kb�'�`�*� ¸|��`*1��	�Ӌ�ݦ)�ɀR�H�M<y��?QO>�1_]� 25�H��B㮚�>��|�'E���Ƙ|��'Z"�'���#;���*Q��D ��
�ێBm`TJ���'�b�|��'���8� 
yBq��XVp!�V�_�x � ���<�-Oh�d�O���BԻ�Q�|񂄵��й�
�.uM(L��.�I}��'�B�|��'���?�yR��IU0-�r��P�,
e���?����?!+On���p�Lq�ы���c5��3`�9�ڴ�?YH>y��?�����?aN��B�m�qiژJ`�K2�x�j����O�˓�J����D�'���l�>~z�)� c}JB�a,��m�tO����Or�:o/��r�@D	x�Ƭ���	�A���.�ߦ��')XI�5�h�l��Og��OK��/B��Ҁ�=h��T��o��|-l�����ɝ���n�S�'U{��8�5-�<�Jr�>l��lZ	@A�9��4�?����?i�'3ԉ��Ĭ�<t������R�4�	�\�g�6�������Ob�S�O�2%������'b�%��nL�i��m��i�B�'V�����'N�����Ugv����Ѳ3]6<��$C"c[���>Y�/�@��?���?�q��J�I�r�#f�hM�v� ,G�v�'�>�z�]�t9��Z��9���+EKХ ��!n�e��"�8y���'+*����������O����OP�D�ZX۠�/}����!S?�q��ʵiY��ʟ�������~�KPh�:��(;��ѹԮK@!9挊&�䓒?����?���?�6�^��?I�A5	�b�2��ʿm�T`[���&A��f�'d��'{�'e��'����<�M+6m��HH�6�4���v}B�'���'���'��Q��'@��'�@�fE�@����%5�����z���=��O��,vMHy8T�x���)e�I�.A������M��?A+O �!ET�$�'��O��;��[.�F�s(ױM�
�cE}�:⟴Ф��D�����R12s��)Vq� �υ�aឌo柰��)p��!��ݟt�������FyZc�@��c�V8�8�3�H�@I" ��4�?�@�Q�ǖ{�S�'x��CD��'9��e�W*{f	oZ�0���	���	ퟴ����$'?1�G������vc�1��_��MS��>'�q�<E�T�'��a0���Q;�4��m�+)���p�D�O��$%w2��>����~�$.N6^ݛ3�I�'x,Xp�����'�Ҝ��y�'�R�'�8��tNю��u�J�ye���on���dB0�U%����ܟp&��X>U�fԒ*��R��Pp�GR���3���<����?���$��T��}U��@8��X%I�Z�H���w�	ӟ��K�Iӟ�I��q���p
�%P,��QR� �2�I�H�Iӟ�	�;�UL�C���n�<�k ٤U�j}h��O��$�OR��4��OP�ąmV��7{C6��ą[���$�j����q���b�95�U�!�ݻQ� )�f���ZDD���5煵Pi>C�I+�F��1�]�i�t�E�mi���a��]�G�-(&�]#N�{1\�����2f�""C�>$���V��1ad�䌌)�~��F� �&��|�SǄ�F$9���R�Ã$%34dP�'�Zv����;6d*��q�E3�l���M32�T��¹s⤡�Ӡ���		�B)`��x��i�4*qP��5"@�XoЕZ���?	��1� }}ڽ���� !�{f,X�>g>���ᓣ�µ�)O�k��p��H)��}E�܏"E,�����ZtHDC�nѿq�A�)O?�DN9v�HY5��t{ ɟ�]X�s�k�O�l����O�>�:�r��V�(t��[P�R�BH�d�O�����{���5�J�9��!�D Ґ
����4����37���+�`V*l-��cu�\�����O��b�gɸ(�����OR�$�O�ԭ��?���{k$�듇�2�,�I���~����')6yh@�C� ���~F{2� ������J:�x3��={}��dE%)ѠUŇ�E�Y���hO(��p��+H�6L�)�Z��F�O�P!0�'����Gy�燛tل	�t
"Y�l2�d��ybIY*)oX��6MP\(sMX�gij"=�O"�	?5��MRڴv,L%#!��5L�����c�ʴ����?���?1#LR�?��������5��P��HLH3k�*z�(`��Mϑ:�DD�C����y������ 
�p�N���A�G�-�dƌB�*dnI�/�yeƌ�?�� ��I0aH��c�8���iWS�e���D.��9+N��B�v2��F��iڼ�ȓmf�c��Y�_{�}��a��ҊYϓI��IRy� ��t�.꓊?A(�����9���CE�n
���W��:2�L�d�O4�DYKюR��qLY�Ѓ�ȟ�'�D3�
eL�I%��h0�Fy&\�&K��/�8V�K0X^�#�.�(<h(����3v�9�J�7���Gy�k�=�?!���O^�H(D��Xm�` ����>���''�2�_�!>,!�f]�J�yB#�� �0>�E�xr,1Wt�ے�#�dK���y��@�-<���?�/�2qYW`�O����O�([7╌(2`�2��)pyRf�&BW�u�!�K7�:��Ɗȟʧ���?� -+����s(S)���ѐ���ANE�!P��d�${����0��7�Z1/��xG��?u|W� Næ���'�r�����O���nYWpI���#ܨM[�"O� ©Br	ԿH�Fl�̤f�AX��ɝ�HO�b�����̔l1��K����ڟ�B7��^�y�	����	�x]w�'�����v^$�� �|���'P e�䔮0�Ԃ�$O䴘d��[p0��(�x���O�a#o��UN,E�x8�<�v��_:�,*#ѦnG	�Q������OR��6���Z��zkC�D?g~��:�g���!�DDZDik�ʗ�&>��5��� ���FzʟN˓M�
�Z�i��U���ͺ�X8��Ƹ.av���'��'���^�r�'��)�#�r6M�OT��w�ԃW¢��0o�>:4����'�0T)pQ�����M4E��c?:�t�¦'-�O���a�'�27����XѪ0#�1t���[�F�R��m��4�'"���?�iGc�lw爺K�X�:�`2D��ꃁ�L��� R�!�4A�0�t�l;�O��l�hf�i9"�'���\�T�r���2�����,Ұ0>F=1�E韴����L!E��u7� �<�O�(T@���V?�H"�;�8tr���K�w�����퓅��aK��j��Z�NZ�Z�<�5��՟h@�4R�6�'P�S�D{��%&�R̆),�5Zz��IE�S��y⅀�{�`�yT�̬�}�'�:�0>��x²،@��ޛ�z��׳2���SH�h�i���'��VE�y�Iǟ0��(egȨV�F$D~�h�g��J�`��M��y*��<Ȑ%�Y��Ţv�<W��B¦�-5�t�����'+�u�i�<���@3G�Д���ڇ!��'T��:#|�	�n<���4�
�P�`%�J:vE0�	�����ɣ uvL��@�-~b��`H�F1X"<1'�)z6��#Y@UkJ"Wr�xwC��?Y��p�����΀��?����?���Ss��O���F�V.�#q��d22��g�V�]��$גt�>(���'T��� $���@/�Nj�3�'H�))��̹��=����C'\pC6�H�Zn�Xa�0�?	T�7�?y���?�gy��'��I1���:c �	k�Uy�n/L�VC䉵��xRG�%D���a�-v*�����ـ	�z�d�<�V�5o�[�w�����gcX(��Lԣ:z����O����O�����O���`>!a#j��Q;L�oڟ�q�� ��q�R��p��R4��$K�`-���v�jӬ�#	E<W�y�Dd��`�����'�X�_&� z,L���2����5:V6M�O���?A�ʟ��� ��: K���c �%B��Ec�"O��CaL
�fK�|�@!P�{�F83�6O>��'�	4J����ٴ�?	���T�US�����Ko����oP"dq��2E�OB�D�O&);ŁP�:.a�#�ɜK�	3 ��y�t�U*XTbE�,P30�F���J2�(O(�:w.��l �Ÿ��^� ��}ZD!�~"�c]��ȴ��'���{�mN_�'���	��*����o��$�|�P���)���cA�/��GG��?���9O\�r���?}4vY�r&�K��!�A�'66O��Q*�t\\��VO�z�4�AC?O\c!cV:y�����O��쟎\ZP/�O&���O���&͖9�n9Q� E�b����V+\��E��.[�0�pHoDl�8��O�1��)�ZU�����{s䱸a�>`�HD����F4�ga/Hp�Տ� j6H����I ���eɖ���w~ܴ�cB��7�To�IGx���'�.��D�,7��!�à]7.���B	�'
�!Q��B$oj������ e�	*��D�I�����'6�����z����(%"���'Q��ή ��Qa��'	�'�2�cݙ�	���x� $z0�2�))A��m�E��ؠ�۠]踝��I4I���Y�mء0��	cmH#�R��\����J�A؞ء2ЄQћ���0R*| �&�ܟ5�ޟ�0�43ޛ����O�ʓA�4�Z�ɺ8�he�I �M ���ȓU�j��wo֪*�H8�w-C�A�X`/�HOj�'��$K�%�F!n��=��o]�FO���덋S~���I����ߟ8�����P�	�|����2b�4nI�	 �K��h&͐e�&܄�	$zaVq�a�˦����7d� �pb�ۊ&�ޅ�#�O��{��'�6L�B�&u(pDur��dDE��ym��Д'2���?�P�+�`
�a!ra� �,D���(R�<-(!
!Ԙ���i��٪OP���娢U���	j�TK�23���Dm��ĔC�Qt�P*��'�"�'a��9d��@�j�	!�,�T>�8�"Ǚ[���(R�7]�la��L;ʓy�j=9V�ˑ�%)s�,g����*W�?����J�b�KR#B�(7�;FL/�`����	��M۠�	�=g=t�:f��}fV�@�/_B��D�O^��dR�4���f�ƋK��Q�ň��Z�a|�a%�� &�y��f��U�I?MON)�0ON�K����}�I���O>��t�'�2�'J<�"��g5��M��0-��I�r<������x�T實�l̈�ܟhb>��P�`Uv8��W�w��Lڳ�3R9IbE㊛��Rdo�$+�"���Y4��9i[�@�(��Ͽ�R�V�$��[�)��	�D�@� �,dj�a���?I�O���OD��9KV�ĭ݈�l��1O��$2�O,��)œlrz��r�)z��՚�I�HO��'��y�ϖ#u�Z��f&ڞB�����?�7FA��L�a���?y���?�v�� ��O��J�T�n^�4b��!Z=r��O��bу��]�`��'p�pJdL.*T�ы�k�ktE��'����J�-O��ϓM��D��h��/t|b���(\���M��(� �v e��Y�l��Ky2�C�5�z�@1�Ĕ &g��y��A+r=�4��q�X1dC�'D�#=	-���O�n�F�Z�;��U� �N�C1f�)8!��R�j)!�H&U��� %f�w@!�䃒p�X�I�$-w:�`:��άM&!��B��`��c��`1d��pd�->!�D�:(B���H�k�h����* ,!�T}7^p��
�T��	p��N�(�!��O�-��9��%
����C�=@!��
�1��L��d)f��� �Y�!�݈58�U��NB���\B	^�3�!�R�%�N��aH�	x~�Y�� �!��\RI�$�$�M�sg@���
,�!�䛁3r*]�f]f�j%h �9V!�=^0Ԡw�ڡҔX�%�D;�!��S>5�d<�􌏚;���+�m�!��D� X nذ?�!t�/O�!���;�&���-z>z�넊жb}!�$]D%��k@��&#6h �L3ou!�DjD|�$��1d��Ș���Z!���B��`���H�~��` �,׹on!��"}�&��w�$�d��"-�Py򡃘9RZC�ˈ]2� ����"�y2 ��J�H=����V�d���g˹�yBĎ�
l�Y4o2CD��Ag��y"@�. R`ɂ��
�){�0;��W�yBoنC��<�e��g����
Ǩ�y�ܳ�D`���1\�1ХM�y�e��sT
�(�M6"���@7EP4�y��F��=���Eņ:$��y��T�g~&�0��UTЂ9r��K��yR웦H��ts�愗J],��d(�$�y2
ԙn��x����&7�$�G���yb�U���Hr�/�@ 6E�6�͵�yR���:42�IС�N�t �ML��y����RT3 ��K�P��v�I��y�I� w7��w��
>�� ��5�y��Ksh��r��04р8�ֆ�8 ز0�I��@�'-����h��'`���b�#v�M`D��|k�P���
 Z�X�k7�LbX��g�)�hA���@���qa,B�P&�`l(��a�y��D
�;LҘ⟼�R`S�w�5"�G]2>���*!O*�i��	9_*z�����6�^y*�e�yͼ|�ƥ�>^�mf��"X� ����(�
�q�*|O*���0Ժ���oS� �����<<!n�*"�X���A�D^����'�K�*G�!���H�bd�2@_� ���?i�)�ȓP�B�	V�ʔ:$�q:�#L��N�J�%M�$�<M���	�w5�$mڹs!6��T>��.x�y�w��	�iL�F"б��ޥT�a�
�'?� '�P�[̫�,7"7pp� ����?�2aɮ>�"Q ��J��y顥A�j�����d �X�h�(t���hu���u/ax��T�'QP�0r ^�_L�x�mS2�Ψ��e��x�
��OY� �,HR��|�Ɖ�#�P>=p�{�*��j"I�/
�@�*�2��$b��L.2��sV�Xd!�a`tMP1L�P�S�'�&����.Җ|�W%�e�����"O,b��3��8�u.[~V�Q�� A��9����o�Š�e��;�,f��|ʒ���u��̻y� 5C�C�A� T,Z�I�E�\rh8��"Q��J��d��=�%�G>} �x k�2�P8��ӡj���uȽgrFD��w�*<�#�_ǀ�d�0 �px#�ң{b� �%r�$���`\xCc'_�ب��J��O��޵W�VQs�ɔ�Z->2%LS�e����
N�`̦D��×�$�r%P�\"�u
�d�O|DR�a���!��~ʟ�]!�d�	�$C��T�l@@���$@�.i�Mچ��Kd�C�*D
tɓbҴM���~�\��Ƨ��4����76۸��S��-���[d�Q3z	��s��zC�����x� \-6�d���S�W$�(�'��'���7�J�#SB�|���+}�K�(dti���ԍ0�BHr+���yBN��
�Z�J7%�71��G}�[�hF �``_$��(an�J�{�4 Q��*��w͔33��"$��O�	Xr�.�l��m���v��"ZU�y*�E�+"	۲�ɭ �^,�Q͊��d�!Ԍ���7NB2So$��K��б9F�ӈ�O�d��`��h��]\�è&c$%1��) }��w�_PMҔP��1���֟Z ��+��_���t2�_B�'GhE���-ʆ���E	q�,@�#iV��6�	�,T��P�'3j���6%C�E㦅����H�D"��8�VAS�U.s������Q2�nك�f�q%Xb��=K:X�/҄I�Tt��`Ն&���@y"L�@FT�}�Vlj��1�K�X�H���j�B�#����A���'��#=�O)0��q�:��*Ď����f�Q��)(F�C٨OB�jt��)�ְ��O��^�x����5(�V�0���5�qOrY��'�Z�0@��HY�~R��S���^O���E �;GZ��Nԩ{� �'���:%`��w8B��':��{���M�m��(��-�hCCHD�T4O�x˲��`?�D�'���ق�J�lk�)�A���}W��`�� p�P�b�#�`��s=O��	'��1O�����H�#����Ŗ�P�+� g� 9V�z�HME՛��xi8�x�al�IF�A�����Q���<QF�p�(O#|B`�K�N5H�0L�B'�:XW�E��iI� iDP���߭���	}ցSd�6^�E�.F^��s�ɉ�'��!x!o�?�	.0��Q���0%Y.�r[��Z�N�Rk
��$٪0YH��ƅ�}�b�XW�ڢ@"�
f�#1�h�9�&7��A:45O�R���^�I$A�q N�y��#�>�e�O�."v��
I�3�tZp�T�$�.�U��h?���M�.[��O���@@E�ajR�ٰ�7ul!3OTE�.E�M�hqQ��֡�p<ɶ$,n�U !�� $Y� ���Ł����J������ x��e�<�3扊�$��Y�hi�OP"z����
O`�"��=0������T��0��b�jܕ'�Rt�?��'�Lz�wT�6^�q�b�Bg�S-]3��i�:fyKׂZ C[�h��LM1�p1�ग���,��$���$�����n� �`��Y��m�д; m��a���/[�S�F{@�tmI�%b�'}F������%�~��O�XT`
s��*B E�%����AM�p'x�`]#�D���YFV@ a�)ck�@ʵ*X'����'F�a��cE��2 �%��*H`"�0I�ʧi)�ej�cA=dZ��A��\&/�.5�ȓ;�ā �F�S��aկ�?@T�7A(B�h�8�Ƙ?���O��5�r�ͱ� ��DM�H�찻1',D��S��e9�$���.$a�x!+�;:1�';��S����Ϙ'Eh� o\CD�'˚:g���3Q�֨@r�$3@�π12��q�[ӈ����D�wn�E�u	ۨIহ�GA�.HEz�J4����� �4����-Kڑ�GG#�b$B?9n��ڶ���]�x�s0�?�!1e�|�'d���ߊ]C@��tJU*Tt���*R��'�rt��F_�t���"�Y
��l�	V���L��'���J��h�$C�&`����t��z�\B V�����7��Ex�{i��[� L�x �J����$��j�Q7O	��lxʷO�r
��	�0s��;�Ŗ�<{�b#(��*�=�a�>'.U:�oܖYo��a�I�ZV�1fj@�Wu�L�q.Y9F4q�g�T8�g̶�'��%�' jO�S�b�6'R���p�I :�`q���'���*&R)j&�q��-q�\[ �I��y"fS�\����ٗ��Dͤb��	�o��d��a�I�}����&�a|B��O 0�0^V,���֦(�W�NyV���mр��O��Bd�4t
�%ǚ�X�,�Ϝ!�.�ZDIÅ�K#�ʬ6��\��΍G �}�1�����N`��1��̞�� ������a�� CKT���i��(�Oh�h�f_(I�N�W�+��5<}h[a.%-:����0Rs�\��O����q�T�Y~!1O|�hYe&~�֪	�n������D�O�}jX;r��,b���*�㞝��eڻ�9v�5|O�a�V᝭{��R���L=c��,����@���1R�����������]�Cϰmk��x�Z�%�|��qc��)���;f�S�5�<;���Gl���AnҸa�T3ˡ�8`F>��?��Ef[��U7�Qyu6��.�?,�n�KqD_|�#<�g�ߙz��Lj�EL,;���h���<�'�ަ�2�ca�T0vَ\���F��=Ț�\��!+C$���r��L��'JB���R ^H@�����Qlb�!�,D �8%�� 
=[�.9�y��B �@�
��ё�~�����R@NH!&�#�/�-�D��`NEd�ebj�"y"!��E���Oe ���8nԢIi�&I;*��d{�A&b*�$��r႔�RJ\�w�D�O�9j�NL*G��T����-g<��d.��h�����'���Y�.��`� VUJ���:'�fL��a����foD� w�d�.��Ɋ
	��gd�?��4�M�,vFu
t��=�R1c�(
�lA��B9Iu�T*#�^=.&C$b�
U:)چNYe����	7�.D��]�h9�� �/v���r��S�8X�4�T�����`����<׈�<��AFQ�l�TaҦ��1������=�d�G-���9��h�SL�V��=�t�#j�I�s+��~E�kA$ͱߊ��H��y7£?���We>��`�(|�K0	S1��xU �怈&ȇ�D0��˟� � 5�`�
5�D���m�s3:P��IF�X��P�@�;��<��AV����λmo~�j7�D�#`]P��y/�\����6J�
�@��<��ۥign�*��E��`\ L~$�
8ߦ�9B�$~}t	����K�'�r=y5@X50��L�w�	|��6]>��5���0�dt��� �`4A'��IK�BW%[5�	0evq��SCyR���Z nP�.t���C�+O��T`a�����=q�`����Û�h����/G𰁒�V%`�qP�����r0	;h�lt@��:C�<�t�O�'6d �$O�tPYD�"3 ��RiS��A�G�� -0H�/�u��O�7�t���z2�l��_�-�@�REEّB.���#��V8�� aC5%�
�:�w'�5p�@,U��3�-E]:�p�O#W� ���y�h(�։��
�(� ��jr���O~r��G%}���ޞ*��=�G�Hf�>��"��/^\�{pk�/:����K?E����W�ra!
�4C���@�N����81'4F)�M1�`��N��#|/O�$1�Dt�l8@W��8SX!z�`X2�N�BƖ#4�
�!4����>=��"�jG�<��=�4�K(3����(��6�x�Ç��3	c���6K����O|uQ�ׅU��]�Ta	��j�f�G�%|\Z1g͕���x�� ��n���?���郍I����ի_�,��8�$�K3+>ٚǓ>���ag�"jE�A���%P�l ��C�ru��l#�nx���y��K&��"r[�t�s�QN���VJШ�viF�>I��#�薅@z�>�a)�ZJH'*ʇ]���C�ă����;�*)�R�Z$_�(��$L��ɹע�B~"�H,�'kU�D�R�?A�'g�i"��
"P��R)�]��͑u.�b
��
?jR��a"���O�����'�01p2}���f�&���H�J��/�o ��k�cB�N�%�Óg��`y��Q��d����%m̓:o�=ad���͢L8�J�~Z�?Q��I�I�^h@Q�4Hs���v"�����)"�1ѠZc����`��\�R �7���/��o�	Q��r1h�ȥ����y��\�Rtؕ�ECT����@��T9saF8:���N�U9޹K�}iE�7fB�8��ݧ]i�i*�gU��'h@��U.�av��BE�]bdŁ2x�$��I:�Ɉ�O>ʤ�3�^H�'�lhB,�%V�L����<��1CDǖeL2x �	�6H
��G�3��O��4���T�5����Z��a�@[I�Z�Cq�Q#X^P	���6J�ay�ɉNY�U�'��9D��X�E�0�9��-N<ʺ����5P��:�S�� �?�&X���&韫4ZE�UE�(���:�/U�+�yRM�=h��8�'����17k�'.J�XvB\�[���@!�<)�j�)1�n��'��ҧ�s�f�ѧ�4���m�R��_�ƀ���oV�N�|	�p�W3/��HI?Q3�#� L���� C���Ɗ՟�H�8���?7͊V�`���-}�L\�~Q{��$%�l���%MĴ���w�IPf܆-q�Y��,O�)��s,�{sf�
��(�#%�ZV]9�X��
�MA<i��Մ㉞k���4��:Ջ�
�L=�軒�N+c8�A��@�8-��S�,O�e�'�>���ŊN �W�D�w'tX@���ԩQ*қS�,��ݿR��Lc��^DuB�S�ℴrvNP+�'v�!� m���)��iS�c�BX)^�� Z1͕�a��Y3q"O��m��#SIS�ѣP��+�"O~4��m�=-��,���y7"O±xE	/6�p �cH��>x|�r"O�M��'_��L�6A��K[�Dc�"Ot���kR�H��O� �,��""O1��.��.��Q�Ɣ*��Ɇ"Oty�O"DΝ��]��´{�"O~h�r�W z
�� �dL�|��"O�T(���E�������P;ıy"OU�'i��~��%*퍍;��9&"O��"W4)���w"��V��"O�@�&��)��!A$!	hܸ�"O��S��e%@��ّ���""O
ݪ4J�:0�fm�eo� >�~� "OzXA�́� w$$+��C�D�����"O� ��_�"��|(�Ɨ22˞T
�"O,ĳ��.D���єc١P�=h�"O�l1�Ȫ����P��F|e"O���		
�i���E�F�>-��"OAI���=P�I��(�?'{�E��"O� �dަI��-�)�au˳"O()����0m�@���AK �Ha"O�Y�����`n�
��F?�x��"O�i(%F��K���c��N+hU"O�Aa�!=~ �jҏU�#|���"O�9��Î3�q'P
��qb�"O���E�҃3H�s��>NՊ�"OB�jp������9��^�8"O�����̏��ZؙW���!򄟏�6L3s&U�q�\�)0�~!�D\d�"�A@S"$2�xA4^�|!�$��u�u�+,;J@���9q!�dV8r���x&��317�=��@ f!�@�dYNq
蛿2�.(�ՃT^!�D3UB@��g�u��z�'��Py @�9#��p���.x����b� �y��Z,!�
Cd�mZxp���.�y�+8%�- �M�0i�^8C���y�Bx�r�h�fסj�������y��F*��fǆzͬ	ڷ��5�y��E4c����>odȤ����yB�֔-�>��4��j�0 �&����y�)�~~n%�S'�e��8����3�y��78WP̳� �J�>�`����yR$ßSj��F�ҙIE�5�s@إ�y�JƷ/3^����P�pT����y�
��LO��� $�5��U�/Ҭ�yR��)VOt��F�Ж&`���V��=�y-���Z��M�-��	���y�ke:,�c R�(�xYR�"��yRǞ�T[�	�V-��(��Aѡ�,�y↖�8��S�/Ȍ����
&�y�FF)"����CiIv4�7MG��y.��Dm"��%��@�6E_ �yb��m%��A#H���t4��0B�B䉕+���c���Q�7/�5W`���A$j��#jC�#�=��K5t���ȓ�(��nP�W����@�/�@	��1 ��D�y��5#,f��&:
�q�gŰH�ׂ��<�|$�ȓ@~|��u`:@S&�%1�Fi�ȓ�v)�����_)����
��Wu�`��<`1J��.�ڰ�Շ!�n��ȓ!$�bs��HK4=��烠@ٰy��caX(����U>	Z�N�F��e��^���"�؍s��,��G&�$%�ȓ="�i��=~W*)����f���ȓ%#$�4#�1BRG2xp�ȓ_�e�t�Yp���gdɨHP@�ȓ6r�1����4r�2 x7-B>b<��g�%Q3���N�;P��%�ȓRK~�C�Jԙ.*`x��8 ���i����u��xbU�$i�����ȓ;2��Y}�2c0׬P�� �ȓ_D]Zs,�� �7#؎Csz�ȓ1��+%rt�d*��F$�j�ȓ}T�����"��0�ށ��N*U���^.�	��L@ ]�(���V���G"ԑ*�"�d�VT�ȓ;��Hz5O� N\�9ceG�2�6�ȓJ3p���JǾo�������4�ȓP�RMS2c߼9eȽaj��K����ȓD�t�K�l�~��@1�O�B�� �ȓ� ��-�1|��ǥC��Ʉ�S�? �4З��?8p�z*V�a@v��"Olˡ��!)�}�ی]+l(��"O4�r��Ag:�)��"l]9"O�=�0��PA�]ZTG�K�q!�"Ov�����7�h�%��!�j&"Oi�-�gmf�Sg\8(���r"O��B�֊5PV�@�f��4uH�"O8q�.1�2�A�^*Ȧ0� "O��@�,!-�`d�geO r�L���"OZ�C�*	/!���(W�F�2��p"On��VO�S��(#s�D'�y�s�	P��"���]⎝�Gi�r�9#$���@"��KXx���H�)*~��0��3�y�%A7(�I�Q͞
	�~Q"����y2抔R}����M��ܩ�+��y��W�a^�IP5I=3'�;掊��'_ўb>���L���VśO�;M�R��s":D�����q[�]��cԭ\y��0�l,D��0p�_�P�M��ő�
��lA@�)D���̙�uD5𖥐?&2�Aj��'D�|)��e�C���,�Ex�'D��6��/���)e/*>ql��1�0��E���'g������=w/�ivKԐ�����Z�����#C'���B��Y�RO~u�ȓrB���3'�c�J��$I(**%�ȓ�v��TH�8�`��n��'�"���q*��0/W�L5 �#��/R��xG4Q���3�VMr��ΓbP��ȓl�HhƇՇ΁P���b��}��Zi���E�՟+/��� �4���IP}�Aؕ&��b���m�@�f�Z�ybNȾe�|$�d,M9�L�k��D7��'��D�����D�q%c�6z��  C�0�`�"O� �J!(��:Yr�\ �ў"~�;#(<ےN	��uI3��p{Ь��PS���d��Ss���`T.4JR�ȓr��:.�1׃�,�T�"U��e؟ ��a��Uc����`��v`%)tXH�ȓ-��i������q��դt�(��y��e�%��j�f��d%&7��OD���n}���Sj��'�<I�ȓWNȘ������o�q(�ч�-�atȇ+Vt)dk!��A�<	�
����d�=D,ހ�&ɉt�<iEfA(��Ppcw�>�k�nm�<YD�V��PztN�5����
i�<�0�W$1��ύhL5���^�<��)B������Ev�x����Z�<�p&��i��a C��.��<�#��X��@̓	��,2e��D��!	�#���<!�u0��⯈�|�X��E�r�vT�ȓ��Ȓd��{�Ԙ�B�q�踄ȓn���Z��CZ1\49K�Uf�ȓ|�������*x`P�� L��%�ȓ���U���,p��ϳ����ȓp"�թ���!��;R�F�%���g�d�{Ư���Aʶ�ϱT�fu�ȓX�8�����p|�P��iʨt��m�ȓ=6����&�8��
�Y�h��ȓCBB��'�q�z���� ��)�ȓ��$`c ^")��I%�*/���������/����$�&��C�.�#�%W4<p����&���݆ȓa٘����pp g�	���h��S�? ��s�v�*M;�?
`��"O�× E�QSvXx��B�%ؐ�V"O�D!I���F�C�/�u �|�"Oj��A��n@9�S�M�{��xH�"Or�#��Rb��rU$aێ(�&"O||�`,ݙ]8N%�L!p����"O�Aqp�)/����1b�|��"O"]c�BZ�f�h�C�;���V"O�5 �.V��@a
�xx���"O8x' �1R���5�G0ktv@S���ą��7w0��zG� Q��m���X�e:�d1�,�@��,/���*�N�u1X�6M$D�|��ʉ �֬*qN�Sz�h� D��)��ȩ>�XBt�$o�.m�k>D� Y���4l���ۃĚ�lL
���N>D�0����;�P�*���7kd�h?D��!qg�=m�z'Rw���fl7D��: �,j��&�M7F��8ʷ�5D�d[u��=v\Y��^�[¦I���2D����,R�,���7�2E�0D�T:�E2q4��YC�!HC� FJ,D�\�6"EhP#K��؄�(D�0[�ٛN�\Ib�ݑyEl�se'D�����nY��9�e=,9��.$D��� �q�6�	�jY:�p`	&D��#��ېB�qR��k%� zqN?��蟤#@ �95�R��@��/Z,,��"O
\��ϋ(�3�,D 'CHс�"O�=�QY�6嚴�I�a"�"OF%J�����ܳÁ�>`aK1"O�Yp��2
��+/Y ��!r5"O*
���*,ԥs��'/�fu�6"O� uj��,���S�%�6��"OPH��ʛD�Z�[��&\�T��"O��P���P@]��݁�R�"OlL�3�		��AC�Ƚ8��8Q�"O<��v��X~R���!+��iB �34��
�o%j,C��N�,�hw�%��`����↳{��#�e�,���"D� ��,�f !�6����5�E3D�H��X�]~���Dk���xŚ2D�Lg�Rc��t�m %t=�'3��.�S�' �(h `��+J�,��𠙴	.��ȓ^VD�@��gf������]��1p�1��ۉ"@�v�
|B���V��sAT�}j�<���a�F���x�r����%O��`E/�
L�l��\bq�d�rض���X{���ȓm�6��6�ʞ�H�YB�.��Ň�V����a��}XF����@<~$L��ȓ����"R�Nm�x)����K���"��P��ȀM��U��D�8��܆�H8�����?�H�@��Y������)� ��n�u�3n��c�h�ȓ
^Pp� ���1ؒ��$B�F��ȓ7����AD:��%F\�a�ʓ�$i����h��x�� '>�
C䉱M, �r�S@��
�o�9�BB�	�b_�$���v`TH��#s� B�ɀa�
�A�C��c�Z$�a�C�~��C�I\�E�UgE�R�3%���X��C��8eQ�YҥJ��*!4�[���(v��C�ɓkV�x[rF �|QD�A�I˯��B�I�O N|����,~�l���7|�C�)� �I�DX�\3���Lm��%"O�٦��# ��21*�=O2b4�'"OV�ڑ�/hs$�{�U�'>��Q"O�9`�Ǎ�!B��GDG�&0�R�"O^��e�
����I���"OnIآf�I�.ʑ9�� S�"O��S@G�lFD�Ч툪(Ӥx��"O�Y�Ő�)��h1�`���&"OJ��P���l<��+V�T����"O�:�	MN:��S��5�xi�"ON���t�$����W��`Lk"O���(U�E�Dh��V����"O����.�VY�(�,�T-��"O�A9"
��G~њ�G�m��"O��j���6����F��4�H �"O\`ae���$=XǓW� �H�"O���؟SI"x�R:�L�	""O��#Ta�0��B$�P\�k"O �ze��(3`%��eN
�)K%"OhD��59V�@�0I�(�"OrȢf 5]>�JW,ݬp��1x�"O� &*0[\��C��p��"O�)T���R��tk�A�`M���e"O6�Y�� �����b��'1\��"O��c�.�P;P��A�d%�U"O&��'��Je��!���:�N�+"O���o����"[k �X��"O�9A��HET��e�_N� �"O$�*�'L�"��	�e��N.�
�"O
�R�E )lܠY��l!"O|! d��f���a�i�)0�P���"O8��M
.E,Dp�tƁ��pY"O<��g�M��"�d�/C�Hg"O��A�V2���#��o�`�"O,��"/_� ���2� �M���rt"Ot��w����(G���8n�)��"O"!��G!	���0e��4X=� �"O���"W�xΠ��IÄAV<u"O��逍��©b%����
:U��ͅȓ!%� ��ឮ.�<!�0�8F��ew�iHu���= ]�bÚ�ep�9��}���I#���6�l�*f��9j��x�����DD��;֐ S�cΜ!x���@�á������ࣛ./$�}�ȓUjF�h�E/A��`����F�T��Bo�(��اd���%��!K1�Մ��D�!���?�&�	v/2v���KG΀�p�@&E�d�9sGO0�6�����y�gĵLm���T��A��'>�m(EHٚp	ty	'm�7W񂄪�'�V�8&�́T<�i��疹LT�L��'/����-L�v�˵&D�?�z���'����@O�R�x㟁?����'ά�Rկ�����Qp�hAxyy�'��d+���rJ9B �M� 4�I�'��r��4�HaǮD�wb1��'V�����s���sgG��v���'�p��A�/(4��c�?�����'���#/ў �t�ranU� 6���'��@2A�?���k��M4(�	�	�'utY�,��f�x����]�M�'Y�ukW�%bn�=��A֙\vd]��'d����+�� T)S#O�̙��'�a���X���1zc�=|9*\���� ��J�䁹�R4�F�������"O:�@� �T~~I���J��a#�"OX؃��:��k�O>��]ze"O`��&�'��,(T�'�D]��"O��ː(�U��1���Y>�RE`�"O��#JN��#�G�8�p��$"Ov u,X������
"��w"O�`���"S�ic%�K";!�$3�"OT�noX;��m�P,��$����`"OX��S�B.n̎�A���
-�5Z�"O��2�ǀ�Lc��3�MB�'+�ȠF"O0�",�o'�D`Ѣ�3OL�"O�`�P��$Y�p\�Fa]�g$��"Oq0`'�pD�9�t������9�"O@�`f�̾U]���9e��B�"O�qs%���{�T��6�����"O\,��@�vC�X0e�>R��DA"O�<�ՆH�^2�dOA9�>��G"OکZ�m�+
�
� B��T��"O�A�S�L�'�(���]���r�"O>�	�J/�z��3Oݠ��\H�"O���ꋭ�L��t�
�@�a�"O�I;FϳԔ�A��ެ�9�"O� �ש[�ի6������"OB������+�F��D��d��mH�"O�����.@� ͪR�)sF�15"O����!D'>�Vɗ]4N\�"OBňe��I���<d)��`4"O@i��k�&q����vg��F=S""O8�(�.� ��С{��I�""ON5���J�,F	96�0=���+�"O�L�m%n)��ŉ�=��Њ�"O���R�ǜ{�6�іnV5?� ��u"OR����=dI�(��h�!�@���"O�|� fʡH���a��ff��X3"OH�'�9�F��n@��L�2"O��Z1��':v�u�U�,���	�"OJ1p�&*�l�[��%�l�p"O�<!�F��	�gII44��Y�2"O\� .])Z�  �ZsY�ɺ�"O�M�b�F�<;ꍀ��̠"<�-�"O z"��9L6����
VA��"OȘqb��y#դ*���q"O�$P�ZlY��W�Qk�R�BG"O���R!�@�Ҹ�� E���Y%"O��bd��7$�ȅ�Bo ���"OLp��	�iFL9�k_H} ���yB����ʡ�¨Q�����(�y�$ٽ?,���v�V	���!MY2�y2	ZGP]�v���D[d��y2�
�M�|d珐���#�+�y�h�1�
}"1mI7y�����
�y����tf�{��v��x�lI�y�O�Mx$)As��#�Z�"��X�y2ʆ���"B�P���i2�y�l 0cm(�*��X��XP�a���y2.�a衙2Ɍ�0d�"�ϊ�y�@҈L��`뉫s���cg��y�����ԝ�+hV�y�GR��yr-�K�<3�a��e�ہ��,�y��/{��8Ү�`�V��q�]��y��T+^zbh�akީ4��!	ݍ�y2�_2a������T�Æ�r+zM����#܃K6���F~��S�? �$˰A�%(Hm�Soޏ8��9�"OTt���߻=`�h`���2=L�3"O��{p	� pJ���l�j�z�Kt"O�@��8�^��%��c� ��4"O�`:�KU�t��e�e2F��J�"O��Y�E�3	b�)���13�k�"O�9h�/�D5Ƞ�N�!0���"O4�$*T�Fj4��F�u����"O��(�Đ"�� �h���ޜ��"O�|Sg��8��%*T�?fL��#�"ON���٫e�@	Q�!%/d���"O:���a�Na����G��6-����"O��s��$titFN��9� "O�i�q U���PC�Ԝ[i(髥"O�=��͐�$�0�Z���oLꐺc"O|�c6L�(5�R휮i�m�E"O�`.�}h � m�8H .�"Oj�+�Z�$��L��U1N8EY�"O�q���5oHqb��:0Z`�"On�8�ےf*�"���S��7"O����(�9p���F�z-��"Oe!d㗬i��pǤЖy����""Ot�����7E����dA�Hw�xA"O���.pն;E$��k��"d"Ov|��/gc��h�����$�""O��0&!�03%�Ȉg��!�Ұ#q"O��,ղyք� F�)]V�I"O ��匇@�ℝ�FM��"O8)(��߉g��	3T#�.q0"u��"O�9��m� s�=� �&�� ��"O*h�tK��Yk��څ�0qΑa�"O�����7h�YC�$��G���"O���6�̽j�욯G)�Đ1"O���w�PX�ì8=p"O�9V��#����ϖ)����"O��dAǅ)�H�㖡�)?'`�s"O|AsֽT�}���Ԛ\-���"O�������e}Zi�g�"�3�"O��p��O��ؠ��v�|��"O�@ժ�r��b&��4�c6"O0E�aZؤ�g. "#�X�"OBm���(?Zhq�W#Y*�^ĐR"OԴc3�<Ru���#D+	���D"O4`���c��h`B�X<y�v���"Oꑁ�kҎ�v%Yb/� 8�2�)�"O.�@埁���e�"&<�1R�B�<y�%��nO��jGmP$x+@EAbD�A�<����^d���ă*I�~�t�}�<�%��� �0q�&zYa��w�<�fcŜ0h&4��i�"j�uÕH�N�<	���8VkR�	sLˣ]�ze�TB�<q�NH���Ѳ�:̼k��|�<�D�hj�캲��9��u{��r�<�s�˺Eh��Z�)Y�@��٨a'�l�<	��wY~��Gَs�UX�&_j�<9T���� �Jցn�z�����\�<�7���D�1�D>`o��eA~�<I7L� 2@��5 
![6�=�ȓ8�Y���^S��	��m��O!��a���bC�.F�&�1�py� ��U���s��R�rf ����*�a��~>�0`aS�`6���X9%|v)�ȓ5Ƙ�"ĭRv.q�g�C`R��ȓl�<��J(���P ����S�? ���F�Z���8�iK�A���A�"OVy�vd	{�B(����d�<���"O�q�'�L(�c��"��s�"O�����i1B�F	SQ�d�P"Ob,3���p�$�`5)�+4 �Y�"O��1E)̳F���wǍ�E ��"OBE1㫞%%��*qf����c"Ofq�a'� Dx����`;�͠u"Oݱ ,Q�J鈉ٴ�&�a��"O~y2wDIw�6�T��&�N��7"O&Q�@���@�h �gJ�d��U��"OhX1 n!��2`��|��T*b"O��� k�����㟴v�>-qF"Ob�ZW��3�A�����3�F��P"Oƌ�2jڣR�b�q��_u�PzF"O.�f��/>c�%Ʌ�à*ɮIt"O�1�Q��1Y"�Ԍ�:�R�"Ox{��ѐ0۠C���T���"O��4iТ"��Q�5��8\�� �"O�m�(��I�zu
sJ�\W�]a"Oн��,O�]�x�J� ���`Q"O����L�R���I�1�إ:w"O�L`C�yb�	c�JX���"O��#�dJ� J(	�P���5�0�  "OܨqB@�G.��DE8��l�"O��!���Ph�p#���P�ƥb"OJ���O(�t�R���  t���"OzR�A�w�����h߻,�ͣ#"O�dj�MJ=C�ҬPdI�(T�<3$"O�Y�6�(_�y��'�3kL(5�"O8�҇�7�܈P�-��E�ܬ��"O±+!`τC;b4d�P�/�� "O<�PCe\,}�B!���B����:w"O�P��F��FE��-ى,���Yc"O`�D5`�s��΋*m�Q�D"O΍YשV����ǡ��w�u�"O�Y�l'a��峰���`�����"O��#���-Ҹ��S�	t�Q�"Oj������&T)�#�@�JVҬ��"O�Ԁ ��҄�0qy^0��"O��6ñ^�f�qbǆs��h��"O&M:���i�t"%GJE���"O��D��MP��AeG�6���"O��Pc*ۖ94�x�#�9Ik�ep"O���w�l��;3#F� k���"O� ��O�t1�1��!T��0"O��`�X��H�hR�Ίj�؃"O���&+åS�x���OB��A�"OfEД"��c�-P.�,�~���"O����D�7+A�Ap�#K��Q(�"O ���g��zc��P".] t� �q"O4A�B�F|٢�U48�ƙ�"O��c�B�&J�A�7��� ����"O���G�<0���� 	Ӣ1��"Oj�¢ �'t�fK��-b����"O` h�C��&���aC�mkF�"O���$�Q�$(H� ���g,���"O�������8XaW@P�j[nMC"O (�E�K�>_�5��΂v��Y{"O�"�'O)��}�����d�V)�v"Ovp���:Ǌ8k.û6$�""O$��ec�b��;O���zH��"O\��Q�$�d.ڄ#|v�y1"O�48�ɟ�4l��"�F.^Ԑ�""O� �՚W�H�0��5聏����t��"O����I:X)�1���`�<0��"O�Hx'���%���bR*�����"O@�4�0"��dkPO�b�=h3"O>la�C7M�8��s΀#(A�s"O�]��Ըua�!ya` 3W@x "O��� Kx8q����+	��
�"O�	ӕ%����ЈPh�� "��"O�X����=��� -"J�S�"O�����7(���U�N/a-�`��"O8�K�,�P���
���L�Xb"O�0��ȾG��XZ��V�*j���"OP ���t
D �����OΡ�w"O"))��Ј�n�bv������D"O��g�ԋ{׸��ek[�l놀�&"O���aC������5ѐ\
2"O��Ke	�+w�`t����4�7"O�z�&
Cs�(��lJ
S��zU"O\$����>�$hV��% �R6"O:s��R"G@�eEJ�atk�"O
hA��$g"x��ݷd"�Q�"O��ɷ��0^�xi4�?y��%x"OD��q��~:�0 ����I`"OR� �CA|�P9�`iG�y���X"O!Yd!_�����"ޒY�dڳ"O���G��'%-�R���*j[b�z�"O�T���9�H4C��pHpH��"O<����&t׾\H@���'-|a�"O@�� ��0r��@��
�ũ"O:���bt0��!�1!�2"O����Һ>B�u�׆��B��I�"O�,c��8!�i�cC�T��@b"O�e+E��)]��ȅ�W�!�|��"O�[�iދ ޡz�M�p�^���"O�p�	7nT�"�D4�4���"O�D�`)D%ٕT�E�g\!z��\g�<���P8d܆��7��5��YF�b�<!�b  
B�w�m�v�_f�<Q�+ʲ@001v��}.�����O`�<)t"�e��9+t/X xr�,I�'_�<a���/e \�(ULH��=�$d�c�<�b�^S��;�F@T�� ��c�<�bJƭ(\��D`(]���6OBD�<y��ɳi�,�b	l����%�G�<9�ŀ�Y�쁴�A�O��L!A j�<���O��rrb�D��8WgO�<�J9OmNU�«I�5|��`�l^T�<� ��#4α�V @�f3���A�O�<QcA&#S��aS��C>��0��D�<ٓ�7���g��"�X�㡄V�<�`HY��%%��E)z=A�nB�u�jB�� G�F)।[;��]j�-�C�	�4BF�t��5;5��b$9�B�ɜ0�p0tD�Y-}�R�R>�C��I�����s3 T�cQm��B�-"�v0���K/�R��Ҁ�0e��C�I�c���;���)d��D��RH�C�I(���:��f���c��A��C�	�*�h�sG�ŨqĹ`eFԽrnC�Ɉd?���I	9��"��Q�C�ɏv׸�z��":k��T��D�C�ɤC~\�۠M�=L�ʦ�E�"،C�I=|��se��H�؛`o�mCrC�IC���"��C� B6���e�>C�)�  ��e��B�j�C�,4�Y"O�łHM)UBS�̋F�lܪ"O2d9�H��5t�0r��/i�H�u"O�<ZQԷ+3hI��ԯg*d�V"O4����@!V�
Ha�N.z(�tB�"O���"��"4�@а��E�x��s"O�\��G�S��I���B�L�bT�C"O$�x��WSZ�Œ��K$E3΄Zd"OB$Dˎ�����g)҆��@[4"O�����F�n19s�T�xs�t;�"O�œ�G_ lb�!&�$N,Q"Oh%[%IB�qmH�B�D�4�J���"O<p(0��X$j|�c�3,u��q"OP�	�C 5:�thA��]W�`B�"O�d9,Cr�9�+]7SN2T!"O���p��V�JmzÊ�!֑�E"O4��R�ܶUV��a� h���G	W�<�$���  �,�dk�-P-���~�<Y��O�j2�ec���2� �'�U�<	S�M�C���U+֑�Eh�#
h�<����>m�4��o	v밍�3��`�<	�'�
b�� ���
h�`�$�S�<q��M�{����玺���C-D�<��)�70��!���H����aA�<9E�RN���P&t�ӣ�R�<�$��;r9b����(1]Xu� gN�<����FFڄBal	� ʨ�8�H�<1���ώB`F�&�8G�G�<y�a���P���cNd�6%H�<��H3
�(��~Bh3��A�<y3+��*��qX�*�7�"(�S��|�<Q�άA�p�(Ө���<ʴ��x�<�oK*�^9�D�1UyHtY�V|�<i�*�l`أ!�5L�T񱤈x�<qE�0?2Hl�q��V�T��E�p�<9Rm�Y�j�"��KL���kǍs�<Y'�P�K�n:0��\��"�K�t�<yF�n�`�3N�+ ݪ���o�G�<Ʉ@�nH&Ļ)H�֥"���j�<���
w�z)!G�4���C��i�<�pm�J����V�5�-�B��z�<�DMǖ���O�#�n�@/D�\R�!���|I{��ԋ>�Z�Q�!D�Ts����{��5�֬R/.P��� D�pi��_�\�f��x�A!# D�p9�KׂW���� ��{�"Ͳ�b8D��c'���T�@A�ݬ���E�:D�|�'�ǹM��H{�(��}��R��*D�t���P>%-��"��)
�咴-D��q�n�'.�H����߼3}$�;��%D��htH�&�
B�	3��1.D�ȃj[�)<�Y-��a�����. D�43�Em�ui������̓��(D�4�Sm��pԭA�o�
�t��l;D��6�E��� F�]!R(���h&T��H�
}N�� �Y,�$0"Ox�s� =���{F�=��r"O2��M�x�4� F�	�$�x3�"O�X��K�%V�椠��8x�`v"O���v�������$	+N8�z"Od�R�eF�8D�Q�>N��ԢA"O���V.��v���#\)�D��"Oh��@�Q	�
����/��Z�"O�p�"�فK�J��%
?݆"O� r��l����eOͅxePs'"O�[�#�`��s�$*p��*q"O�|qf��0pJ�j�� y.d�`"OY@Q�������K�%Ib!R"O:�a��Y6F�eFV�]4�	aE"O�]!�,�r�ڥ$�9��(�p"O��(`�G"]ax��5��6�@\Z�"OpE�kٽK�26�'b�+��yr�?|���W] i�~c'W=�y"h/8r��9��-v|�SF��y��N� �Z$"&�ԙ.���Bn���y�43z��e?.i�" ��y�/>���'�v^�HH���yRO�:�<�F���k-f�H�#T��y�/�/��Q��@�i�@P�a���y�%�-8��dB�\�v������y2Ɛoj����QL|%����yϋ�=c���� U�Huc�����y'A-��ѻꁸ8i���#��>�y�@	�|��ĺ�A� bf-�B���y� ԎD�B@��dʫc�20�q���y���%O�z$��îb�R��FI��y�o�v��yB,�>Pۤ��$J�yRgJ�F]���#i�F��)ub˃�yr M:J�@�%�؈!.5[DM �yR,*�ܠBQ�
��<����y�Ƥ2�bH׏��Y��5�yR�0����B�o���Ɗ��y�հ�@s6�G�o����狃�y�"Y+[ۦ�J�nF&hUH��f����y"��?�~��5!ĩ,r�F���yB�/��P�%EE=#;���X��y��-A��	G,�H�0�'Z��yi	+ ' .	��8b�Y��y�b��B�zy���>�bԸ�>�yM��$X�Q�ɔ4z"I��"��y"�Z*F��2	�s��p�5�H�yr-�(z	�K(���c���yr�Χ ɮ� ���j����!W��yRIڟ>��,X7���~��˥�y"b�BR��P��O�u��%���3�y����u�T0��Զ%�����y�i٪&���3�ς����f/	9�y"τ*9� 	����#U]�6�֝��xB�_:l�3��d`0Q��B��ds��)�'#��B�x��\��� Ԯ���'ߨ(�dM�xF"+ѠOy: ���'̈́!�a	R=��|Y0Ζ7mV4��'����7��Qg�]�͇|��)�'	��A@f�I��=b+��d)+�<�0CJ�Th"�`To��|��őz�<�BK�5x�Q3ul��Ir�	quK�x�<�CF�	X1���ڻz2`XPǗs�<�.I�E͎Q�&��M��ĉ�Bp�<I�YA��p�3%X*J��i�<��A�E�Hba ��S��(W�1D� �r/I#-����" �+j��!1D����M�^���1��QN���0D����ݏ0��Pa��Y�Ytn��1D���3;g��s`%41v,���-D�L��M#"N�T��F��dJ>����,D��;�ϛ-���K�'L�V���%�?D�l�r��q&A�ui	7<8&j��<D�L�"I�k�i��*I���A:D�� zL�ԆV|�@�ц<=��B�"O�"Da��3�%ѳ�O*9��p�U"OT��܇|�<�jd�X9*k^$�"O�*�.
"�� �um\�}L � T"O����g	�^NY�f��*���)�"O�����	4�p�y`�3op�8b"Ov�4�[%j�2�4�C�?6�""O��ыК]*��聎��[H��vO�e��ݷd ��C�P� �ؽ���O C�	�'��cQ�'*�5��c�B�	#&)Q���*t��׏C�7��C�I�'L8�BcJR>��5Z�m�=x�C�Ɋ	t]ᇧW�)��1(�,�	��C�ɏmnR��5$�k5��4��L�B�	?4�&M!��[58����O C��B�@�SnI&�RPc� �XC�	6f(M2��JͮT	��Er�B�I�B�Z!) 4�������@T�B�I ]X��s���	}�h�*
�kB C�I���P*�-@�`G-Fu��B�Ʌ:*ݠ`��0�"�
�䞷T��B䉄W�}�5닶)ζ���l"�B�ɤ^��h5��_e�q��,Q��lB�	�::�0�4�� a�ii��5PA�C�	�.w�X@�	@�x��so�BS�B�ik��C�!.�PTJs #R��B��(&|r(��Z<
�X{���?"�C䉹W�LB�`�$m�$�6b�
b%�C�I�B} ��F��Wꑸ�O�K��C�	�p�n�:3�P����	��C�ɝ+���)���$d�yR���3!$�B�I}N���D��,2��"b�˼x:B�Ir��Ӱ	T�3C.h�.�(ԺC�	�|�HeJJ�~}|3�C��u��C�	�6٭:D)|�#��L9^�̄ �'��twkB�am<�2&��]�4<#�'`�Y�GF�&�hMY1�G�pΈ!�@"O rF`��V����jǪ�ç"O��"�Qhf(8�)��y�]��"O��k%�K�� �h�.���2"OPH��IR�gߜEH��V�;(F��"Op݋2��7F uY���EDX�7"O2�aԙ�t�a�\���qg"O|�)E�bu0����BE���'�I��HD{J?�`6FH,B�h�����09���,D��r2�88�a"�F`���vF D�8�w%��o�v�b���˸�Y`�9D�$���Î�%!���Hx�,���8D������2��%�DH�df��Xt�6D��PPbV���tRD��"c��P��*'D��p	�Z5��K�x��q��#D�0�hT�����͝�qQ���,D�81#�C�J4HL��&(JLy��*D�4�#��o�$,[�nޣx$��Jh;D���!�1v�DKg��z���w�+D�<b���h�L�B,��l+��ia(D�(z���l�(�i!fm� �@C䉬G�ny8�eJ�n�d����T�PC��!n��ۦ�M-���EҧeblB�I�h��rjC�E� �+��R UBB�Ɇ$��HӋ�p��H�I5V��C�	�Kc�D���H�+�>�s4Ø.SM�C�	 &���PW��0��JD��"O.�;@���Zy)�b(0s�F�d�<� �e;3�]�n���Y�V90��![S"O������\5<b�B	�(d"O�Pb��)@Al<��- �G&�-Д"O,�0�H^ M�Ђ$��F|�p"O0\#�I�rS��gE��w$UH5"O�a����i��A�C�L�G i#v"O~� �'��k�h�aA�߅�����"OT�ҷ�[9�%IR`ѸC��"OX���â/�X��s �!A�J��F�' �	Ɵ��IM�3�I�C.5�éD���РdT�*pDB�I�E�v\�`fJ�/���!�P<#\B�I�{���2��ϜF�j��լP��TB䉲.�,�(�A��X�|"Ċ�7тB��+�ș�F�A4�X�.�7I4�C�ɠcf5b�y�P](�La��C�I�yhu�4�ßtU�k$�A�B�I�6!<h�%��;��"�N�rB�ɱ�@ZR���I��dP�HU��C��~$�@�(A8~��R'L�|�C��9
�����(�1��a`�� Im�C�I6S�>�p�BܕTn�a��Ȇ�=
pC�I78��x&�RI��� �Fq=RC�	 ��	�oJ3KΪ!��oU�C��r�L D!�x%8��e�"8v�C�:&����aa��Q�d�BL2�;D��	��31��8�	��U��2�n9D����T<p�5��IK><6θ��a6D�0j�뙭]�` ��S\^��7�8D�4�c�ǾyF���TH6rD	�&7D�T��`?*�蔢�ᐭ>�[�2D� �`K6��
�iκk�@�Z%D����D�:=/YX0g&���3��5D�`��	md��� f�q7�>D�T� Y7*h�;蝛\�f�C1O=D�L�w%��RN�$@gjְaQh��TG:D���de�""���X*�@03sm6D�
�� k1�$�a��(�4ӥ�6D�0!�	A(U��ٷ%Y�l�x�5D���g!
0�Y�"�V�*&�|Yn.D�@C.��JX��M/cg�tu/8D��%�Į}�h��u�'A��4���(D�0 A��Dպ�qP��7Z�;�d$D��
�B� ,y{#`R�<<��Ǆ!D�`q5]!jH�;�a��Q4�	Ƃ!D�vf^��.��Z�&��d���2D�|��a 
l�,�H�W�w|�P��2D���v*�J��T��I�Jר�)�`$D��c%۬V.�K�*�T���o'D�����P�<@$�7i�8/x�D��7D�|ѫ]!B�J��f�2"j��s"9D��	!/N���:��R�J��<ȧo:D��ђ$W<7�B����(1�D�7�$D��[���t�P�8��
#8����("D��-),j�p�FE�~��
!D����I֨~f���'�	38Ieg9D�p�2a �v7��3�D98�M[� 7D�t	 "ro��J �@��	�6D����O��/��"���7*��p��>D�8�gF߷K�$���-�\�b=D���)΃Mf�K1�
'���%F<D�t#8U7Z����N�0ȃ'D�أO�p,1󂉔B��[�J!D��(�I&f�~1��FE�.�٤�=D��h�"�.7ha�эD�$��2�- D�� `�9%��9���Q�*c���8�"O<���Xp�N�R��6tO 	��"Ot	�Ec˝5��<��BB2'����"O��	 ^$��TY&�V�<��7"O>��$��$�>�ψ�KnxKR"OvD
���*w,�)@'�97�j�"OX@�C�%t,��*&a�4TQ��"OD�ЍR��@+�bù'&]+"O����D� r*h(��!>S����"O|XE#Ȯ�ij�.C=NN��(�"O4�8���]��Җ��5B�<�e"O����ņc>Lx�rk�X�p-�W"OP��� }v�a�
ޞx�9�"O!ڲ��#O�`5B�hF�<c@���"O�l"� �$"n��ҧ�wa��%"O��:�I�n�t��@�L�]/�0��"O��V��'5���&��2%���A"O��.�,��5�O$i8��@"O����+U����N[(X��@"OP)��&XP_���L��M�噖"O���EFW|������T�&"O���#A��x\�C[&��`p�"O�9�d��((�S����N�x��"O24 ā�9ϼ���ߣ���f"Ol�*E�B7N`�1	&
�H�#"O` ���-�ҩC�֢0|D"�"Of�u�'-ض�g-Q� "AҒ"O0��BE�?KVv�ӕ̘�^|��P"OL`[֪�y��u��KĨ�
�B�"O����͉+d��i��Y�:���	s"O����엋�\!Bc�(�Ψ�0"Oā�Q��Ȭ:���$�(��"O~ݺ��N.F` �a/,2�y�D"O�eô��)Q\���m�S`X �"OL��ԩR�f	�p�&4P�"O4�C2�nq�!cS�ުdI�d�@"O�a҄b�,Ma�P�&Hu*���"Of�
�ǝ5w�V�r��
D���1"O@1 ˕�b�R�cE�QJ$d�B"O�TqBl�;Qߴ����ܢ'>�L��"O�i t�X+NP�`���P�$"OF쀇 k?4�(�Ē7!^��v"Oz`�a��X�pM�&Gx
�yq"OZ�b�ΘyM�Y����Bl��SW"O����+q�PÀ�6̘�Ӱ"O��� �&,�Bl�#/�$�M��"O��r�+5R��`BLM3<��=��"O��H�J�ܚ�d���Ĥ��'Ӱȸ ^���<�E��$��a��'������,�N�b��$hĊt;�'XaF�ϧ.<���0��W_�%r�'����e/�9P��{�i<T�
�'��Y@��K���"6Nȋh^�,��'��X��J��^Լ���%�].���'.��Z�U:�^= r%ܾU�9��'��	������sO8N�y�'�8�s�4_�x�.�:�b���'��ع�� v��PK�ME���
�'Ն����m�&!�I�o�؀Z	�'�^�	�:���;�F��ib@���'���@#��w���� 	�Zz��	�'sNɊp ���%0d�)˚�-D���fI��O���jէ��QQ�-'D����M<7a�X�#j�7w��0���"D�� � �6&O2-��C�E+3:�(F"O�#�O�P���µ�"p�TBU"O������(�L���aS6z�t�a"Of��W-Rj�L�g�y�["O��a�v`yу%[4ڡ#0"O^=h�.aS�,�dFF�S�4��""O"Ip%�,t��	Iw��`�"h@�"Of�@"��k�p�P�ߵ�*lh"OF�	1�^;F-�8�7 A�Ne��"Oе"�E݉8B`	A�lJ8J�4�3"O�Q��(G%f�) jZO@�x�"O��Q���P���b�N&�xq6"O�)S�=;gƔKA'R��4��e"O�aP�aC�t��� �6<F�\:�"O��(P�ؠ���R�S@d$��"O8�cpf�9}�8P�F��+(�Z�"O�tP�l�4=�y�u��".��"O��1K���� �z�IS"Oz�:�ȏ::�Z�����G�P��"OL�SM�5����fCR~���"O�
g��4s�E*�o�/���i"O%X±}��SS	�j�$M0�"O�8���.����G�n@��"OR�@wMMIr�J3�պt���"O��[��Y�3�x�E�t� -� "O4���*�FYX\��BϚ/>����"Ox�j�H̓u2�a ��s�"O8�r���*7Ǽ]y6�����z"O�Y�5+g�����Eҝ���е"O�Ys�T�c���1U)�=Q"OȰ�է� *h)���]�ljb��C"O�AxQ,�
1�vYZ'AZ ^^�$�"O6�XR�Փ#�QQF�İ|!�`��"O��K�O����$Ӎ	���۠"O
�W+W��]�.^�$���Y`"O�Ԡ��A�9�-��)Ag�\��"O<�QT��j ��`q-�6��j�"O�H��T<���w*��{lr"O�� �%�6u�J��qJ�<0���K�"O>tI�HҺs�V�"����|I��"Ol�j�)0w@Ӧg�Pz�"OAj#
�����3ㇽ�NL�"Oh���_r'�����=?x�h�u"O2$�ócf�C�"hf��J""O�9�',�:��8�&b�T	"OhL�A�N[@zA�aj�MUfI�"O:L�$�2C�Xi�D*�:7G@�"O�ٸ�#�~�l}rQ��u)�ض"OX!C��ϫX�2��#���$�x�x"O����s����S�|��mõ"O8h�0IāOJ�h�f&��S�`�1"O"�`%M�d��M5��	�ȅ9�"O� QF��Y�}�b�W�-�T5�"Oֵ�& ��>�1FW��� �"O0A�S�Ǌ���"t��R�i3"O���tm��Ut}����U50%�1"O����$d��a� ��=!��"O�%�gn�yo
 �@��Tu��"O6Y3Ɗ��y�å]�7��!"Oa*�Y�S���$���l-�"OJ��W�Q�aʼk��r����F"O�C4���n�:v����f"O�����>�
8s%Q�6���8�"O$�ڀj�;m�Д{f��K���"O� Є�%HD�Q�%�	e]��sB"OZ1k,�~}�0#�%�	E���"Oꈨ�«;Y��E�[�7D�(1�"O<���ź,���Pd
�lQ^5Y�"O��z�Jb%߸u�X�+�&I!�M���\� �Ύ����c%Z�O�!�D�>���H�HϒP�8\*##˾-�!��&�d�?�ܩ����!���1w�>ܑe�H�4՞��s�\�!�d�+t�Lp �/,�D!�!��o�}���a�����-�!�d�~"l�Q�ů>�����;U�!�dB|R����G��jBg��Q�!��=zB=3�- N̰�CgeH�P�!��	1>��*(��F'Ռ	�'�vaZ��J�,E|:��������'6�-�"νZI�|c�D\�n����'7Nl����e>\("g�	�j*"���'�89d�ӈn$�i)�OS0��
�'ئ�G�� "��9Te\^��:
�'Qt��5��$x@�X�c��RT1
�'�x� ���)��l�R��;���3	�'�hA�Ɨ�b�	��u�!��b/D�� �Eտz�8���"W?��M��+D�p	u�ȡ�ʍ�7#��6=�Q�@�*D�ē��ɂj�d�𧎒�+��1���<D��������h���JZ��je�'D���r�X`�xhbI��V|�J�A)D��B̝'��i��\�j�u��G,D�����A�;��H�F�ئ���	7D��2S�ٶ:N��R#����� �6D�T� 	�M����K 8���HEF4D�<�0��(��Z�"�9 �S  3D��a3
�B�⥺�g��8-Z�XWK;D��䕪k��Aa֏�A�F鉂�<D����#��
ơ9�ܙ��P
�l D������:�H�c6��,i��*CN>D��چ葨R]L��� �j��q�"<D��H�fK�ar�ү�8�Di1��:D�0Ig�͙=�8
P���{�-&D�0���\�G�i���Jv��Ua7D�,���ڜ�d��k(��:��9D�pؗ���z�� ��GW�R�`���-D��a��]+c�:�K�AH�������.D�( m,Pwl��C�:=���-D����E��EG�1��;F�հ!�-D������6(���Kg[4��1�)D�tE�_2̤�#�p�K�4D�̫�#�^���S�ɥaS�\��2D��3$#^��,����iF<�8�G+D�tQ�/$|�x!6`�)��p��)D��PѡO�3b��[��;l��Qr�'D���s)	�=��KF�G�@y���g)D�L(�G&Lx B�F� ��陖A2D�8�S��Ylx�Ad��wgҍP��"D���@�J6Ti }��Ķ{��
!D�P�J�IN:�a!)A8P ����+D��)$	�)`]������ ^��ix��5D��k��˵n��" C�;S���T�2D�܂��9s��T30`;-:%He�1D�`4n�e4��]���d�tA#D���W���=���Qj�c��P�- D���ب<NX�!�#�0_�P�=D�\KDA�;]���`DT9(�0�g<D�� ��x��^�-T`��I�8Z]й�6"O��{������H����PFt\8"O��E)̯t�N�*s Q&?���"OXC 	7/�j�0Aϒ	���!"OB���N~��C��e� ]z0"O��PD��W�~8���
�l�H��"O�$`��	�%¢��=J0H|��"O�"�N�	�F�[�Z q#��"O���2�
-�ԅ�g���"O�� c��E�x�;��Y�P�z�G"OR��T��<c|��F��ڀ�T"O���L5E����5jڽqF ��&"O�|���_"�K5�G=,�@�"O��k��e�^�32j^��+2"Op,��L��d�lA��k�7r""O��;q�>:�p��$��$����t"O�`H�(tLVY��#�I�P�c�"O9�d`Ђ��\��g�;�ܽ*C"O�(�U<�0�ufZ�a����"ONUP`�X�j��c��7���B"OHha�DzΤ��X4K�~!p"Oj�Ǝ^Lt�����͜Nu����"O�8s�,�@EF9�����d��`�"O���'
Mv����F6fj�,�"O>�H�c�;��Ĩ���$3eP R"O��(��:3�����+�p^�=��"O^�2��Iu�ث�J�?\�ц"O6� d��4J:%cI�/,VTR�"O����3#֬�A��(H4"O���R�W?]1��D���zl�I�3"OHt�@�ξE��IO.Xg2�"O$PJt�Ք�\�Kr(Ӓ(g���"O����A,z�vi�"e�"p-A�v"OV�����X��΀�L�C�"OH� ^�w\va���5_D8�2"OV���K��`�\�#�A�Z�	9�"O~�k���*&6,�)�/���r"O������|-Xsh�]�� �"O�d���PW��˴i�98�p�"O&��`Z�H�xj$_����"O2Y�K�L,X��h�0�zy��"O�U��e��&U%"�쉱�"O���K�t��EıT�L=@�"O�|)E =��X8%�<]ΰ��"O`�� �I�"���Q.�*8�DA�"O���wh@#FV�� �ƛ$EjH��"Ob�a�I�$��h��u\�9��"O�@ږ�=|��CN�;t�F|��"O6Mc�U3,`ȩӌ�?.<|M�v"OP����  �5LI6-�2�p�"O�Ĺ�R��/і~f�#�F}�<)ċŊ'"1����F�m��${�<IB�Ҿt����7J@1�t1��Oq�<1v.�{d�C,��s���YsM�Q�<�j!V�Pj��<�vI#��	V�<Q��<!h�rT`P�H������R�<��ښc����JV"Od��3��Q�<!bV#<��l�v��,�]0$�XJ�<AD��f�,<�%�d=�����C�<��d'.n�B�y[@�s�B�<���
5]�6C�k��F�R�P�_G�<1b�Y�w$j�b��(��D�sh�i�<��T1_��s���`���@�}�<Q�K��h��Rϒ�o�D�(!��w�<� .M��kϾoYذ�e*;B�b"O}�H`TD����4�,�'"ON	��
�{��كP	�p���"O\Q�i�"�t���(��El:tZ�"OS�B<r#�������٘�"O&�uN�M�&\@s%T�h�"OR�s��R
 �����\�x�B�"Oμ!��M$\:�yj���,:��cw������)�'b�.�z��D�5E,��U�T+-���ȓG|����@6��!ʉ�T4j݄�d��Ց��L�Z� �hC�� ��لȓ$P�h(�C�����*8�����m~�`�I	F���{Q�O�k��y�ȓ/�<�k- v��Ce��$���ȓ�$��`��C@�to�YO����v'�,�!;[,�cR�L>j��ȓ|�Zݺ��: O^�Qa8Y��=�ȓ�~L�p�X�f`@�k��EP	��X�'���ˇ�ދf>��r��[wߦ@�
�'E^��I��.�x��&��kl�i�
��O�]� ���;����t��N����"O�آd�T�#���IA�C�(���R�D.|O(9�e�(,�����F�M &��W�Ix�P�֪Kq��ՒػHʂ��  !D�01�dJ$t�i��Us:*��b;�Ox�ND!��ș(m�*�r�'J�'A�����i�'������C(��L�doת,��	�'U&К�Y�F|*�"�.�9�'~.�sDE�^@ �
��Jh��}2[��D�4�;�i�ω5.ot ��"F4K��l 
�'��	�0NޤBDu
a�R�={���'�ў�>��60O�l�vOύaB�PR\�Rh����"O"=���Ʈ&)~|A�/r�(��U�x��ɉv�*�!�'\,��h3�ӆ��4?�RK�:Zd�q%^"2�]
�K�b�<iH)"�U�F_�R�6�P��c��o���T��<s +؞]��@�MXvHqH�H��<�N���뉃_L��*؛g��Tr7��G��➴��!<<O.��2��gdİ���50�K�
OQ(�(�(���P3��Z��� �?�O��'@Q>y�w�?%.F�Qr�W�"��sj+O�P���^Y��.3����P��C!��K3C�Q�N߹��j���<J�'2\��=i��)_�#"���نiѠ��� \!�ӵ[��q�BH+�lpG��
X�!��W&Q.�� �ѱ��x�g�G�K!�D��*z�%�6�%RO������tFbc2�Ӻ��G"�2`y��֓pTI����<�a{��#�8�N�r�AO-x<q�֧E�?�C�	1��]"��1rY=����n��#?���	� �҃4qn@��C�Ŗ��D"��OX�X�G�6�Kǃ� �< 1�g6D� ��gìP�n,�!�%o��آ�2D�̋�g -�d�XF��>p8ё�N$D����*{隬B�#}�����"D��rt�w|�|X�o�8>�Zy8��?D��4��/WBp��	� D:6�ʷ�<T�ܑB֠a�y�V�V8�"��"O��"RE��4o�(Q�2޸��"O�-R*��c�@{��~�VI�g"O�tp��3���wN���{��'�S�)��Mנ0��������!�dD�Q��T`�ł;%B�r�cAz�!��� I&Lm#$gZ�z36`�'�έo���m�RY�y���� �mk��%�����y���9�"O4�J4�[6LQ@�T�$jc�]2�"O�p���PZ�z���,U�YM6��E"OLA����
�J�p+%5(&�A��hO�	�I&
�HêO0S��S�c�#t!�΋z���#�+vx����H-k!������&
`$�ba��W!��G�l ��zM� X`��?+3!�DA��p��<1(@ie�*���������;�IfVaa��'qTZ D�[r�=��+!�,�4
�$B2*��v��Gxr�)���)E؜!9�/���Z���e�<�'$�*zY�Sh�AJy��c�b�<a%�`O��b�&�\��D�`�'��?�	&�D�|�9I�L>b��� �x����@���0"�ci��H���h\^C��,-�y����`yl����L5B�I�7^~��(L�vV�B#�$����o}b�xRW�H%��]mi���ܭf��A	WHɒD�B�	Gn�a�t��T(UKBI�u���l؟���^2ϸe���P�
Ljѫ)��刟���B�P$<�R���`V��6"O���nN$_a����b�>Y|��0T� 
aX���O�>���4�ٙ!	,����s$;D����È dF� �ǢS8�h��9�hO���_!>�x���'@-2�YpdABxC�u�p%[Bȅ�t.�1�-@\<��hOQ>-�!@�*d��w�;R���eh$D�#�¹X~N��Ek�t8K��`��&�P��ɝ4��T@��P'g��@S$$�'���D�<	�� �B������P�<Yq�
�,�I���؅��0"�^�	�O��)O�Ϙ'�6r�l��Xm��2IA�L��'y���ʂ2�(i� J�Y���+O"�=E��BR(�(�d�E�{3�%jU	���yR��1���5K��`A:ըL9�M�1�:�OfQð�9I�h�#����3���2�	@≵;1��%�4Iˍ;��HǬS3D�~\"Ox82ej �'l�a
�K�hb���'�qO�P1�O�/��tX`�� ��lk$"O�@�f�X)un.�C���5j>mQ�"O��٥� H��#J�'s�2䱐"Od��1 ��z1�@w#��:�e�x��'������x�P|b2 ͳ=Gb|�
�'����,��)3�H"sɊ��Ԑ	�'��<���+���p�㖙EBn	��4�?q����iE�(� 
9"grtja.ֽ-Ԝ���'��L�%��(�x�db�>+'���'�x9�6"\�dƹ���(�e���D��u�S�Y|z����|LL��'�T��ɀd~�0��y�L}��ORVB�'�a}���n�B�#�"�����	�y�!�O�����A��Z��C�����$.��i�U��@"cK�&t�H�+�	!�dU�=��I��ɖ�:	Cd�Ԓ�PyB��}h��0fE4T�hi��*�=�HOL��$I0K��2�A�(0:g,�+9zB�| �H��-�4`>4t�D�h�vB�I)V�xx���٥{T�0#b���a&O��d[�w��@�B��@K !�Ыԩ#����'x��D͡լ�E2��j Ep�zQ�f"OŃ�Eѽr4Jh�vː�r�ƅjv"On���%��),"ݩ�J����A��'cў��'�`�4�N�I�. `�͏$kP�	
��� LiZ�`��8��& C4rV��ɂ��@x�$��ק[��M��]��b�yQ*O ��O[s�8��F�6ˬ�"O��Qp��0RX�B!�1��m��"O8Mc#ĸQb����L
36H�"O<�9w#	���;���=0@��`�"O�@R��%74���WEa�j�8`"O�Q8��̈\&d��$�R���)�"O�`p�=�$��E��ch��+�"OذSKN�{,l�PU��W9��"OHY��m�j�b�0����\�i�"O����L�Q��`{&aG/6)�@"O�L�!^���h� B4l�:�"O,���E>v`:wτUTب$"O���4.Zl�Np$m�P��(�"O���GGP�.�I�mгz��8J�"O���쎦6�d��lƌk�H<:�"O�4i��ݻO~��Zu���,�e*O8��@�G(\��d�߱nHT���'ˢ[ե-9+(�񣤃�e_l@��'U�h��V�L���r��3VU���'�d��'�I#==���Q%�Q�2�'[�Y�PF�mʨI;Xn&���'*BY���D1@&�\b6�B)S`�	�'���kd��@����-P4vj2�'IZΉ5n�=H%A��	Or	9�'?4uZRl�	R1�S�|��UP�'l�b�yP(�ss�Պb���r�'�Nٻ�'�?L}�b �� 0Z���'�N$MݿI!T*`�E�����
�'ȁ���ߨ�����T��6m��'T�`y�i����@�l�-`�,8��'X�!�ʏ)"U�����ӧ]1�0s�']����Yq�!բM�S�ܸ�'mqM�1X��ԂěF�T��'~���ƄR���s�j}��'�x`�@g,?�TIH�o��-l��S�']�Lc%-� p�� 4q�`���'"��:qK��s�i��A<:�B	�'!R�I�=B�0�а�.4�tІ�ə_5v�ra*N�Y�h,A���<l|!�V1N\FC�I�ph����n	3��s1��.1U�B䉤P3��jE(��:5X�s
�.YfB�&/\��6C�<�Z����[G�B�	�K�l��!��#L�p�fA]�6�$C�ɲ(Ȃ���R�4|Zq����.C䉯J<�����#����ЅM�>C�ɴ^��+6��by�E��Պ0�C��@�艛1�B�9@�$��J�9��B�I�U.)��-�-Mq�8��L3l?�B��4gb"l3qM�I�����$��R��B��!mh�mV&��F���)C8�B�I�/	HRW��"t�\Ȳ��# ,C�ɔW���񁋓z+̴8�	�g��B�I.a�&�K�Ǔ�^�웕.�J��C�ɺ> ���V��j������C�I�'\*U����� H�#��o�C�	+?mz�Pd�0U� �'˼[~�C��0A!�)�8?�p���I
`G�C�I�c̹�TO�6�"bUZ�'E|C�Iq��IH��'=�$ڐ�?TB�I�$7]2�`ݲN`�*!)ہc��ɑ�}�I�)�']�^�!���->��|��lh0��hN���7g�UвY�B��ڎ�'PI�V��1{�`+f��� NMѴk>�ı@`C�=E�Z����'�j�`�k�(+�|�X�B�%�����c��$��'�.p���"lgpX�!��%����b��S�ޣ<1U���na~D�Qc�'����J|b˰;����'\<�<��KUh�<�w�߼Qb%`�/�+lJ�:b(�.���a%W B�R���$-"���F��'s��zք_�m���'A�l�]��' �hY"]>kv�Չ�H�I�J�CD"��D#�����=������F �lE}�( p�͊��.+?d]�J��O�@�,X*쪲㖴C���(sH�u*8����w�9s�F�3RmL��R��>���ɰ3Ҹey�Ջ5�Q���ԋr�T��ۖ6V�@Ӂ�5{�D�g�ղ6٢Qs��0�E��?q�cD��B��ҧZ>izabU��~�<Q"NC�2@z�f��T@�q�&�$i�.g쑣��U4����O<j��/�(����O洉dSN��;�+	�bH�����?0&dz���o��P�Qs��OV�З�L5"��=2"�̥(,��� y��|s�ϛ�%��p��`�MS�H`�	ʙw�|4��.�1z�`�jv�L�`׬ǃz��'�P��Ɓ~� �Wφ�b�T��D��p�b�'�T-���3��ǉ��1z"�۲��#*Z�OԘh�K�db��'�3�t@G/�d J����u#�j�?{p�:@NG�a��' @1f�2�ӷ��-�p(6�@w��sL̈Q�t�dM޲$�8e�W��e?��ě�i��9���?�,��� m��E�a;s���E�݊*�^!��ݗ"�#g��2\�̽�8��I)�aC9v��0�կ�)�N���R	�t�T��G�B=2�΋>xF�2��O\0�t
��t}N��S*�|�I�EK��i�G*^�h��K�A�Bٹ.�<��+!O
4{Ǭ�AT�U�|����8��@�G�
�E�X���nq��!�J�θL`rEW<_�-�B34�(��F#^d��u��by�'�H���֪C��y�p�ހK'P\�1�I�[�8�V�V[�\lU�L~\�;�a
j�d!��.���^	���'� ���ב^�t� ��yZw�}��mW�0Ɓ#� �&k6���
P7�x�z��]�dFM��܌�M�a-�6̑;� 5�;aVx s FG�E�������v�iL�� �M�L��w�զ�S�	f��*0�^���7�F����
1�E�`��.Q���tfU�弐i3��$�z%�C`�ʛ3�mѰ(�V���q�f�撝�D-_�R�!k�^� E]��i����@�R�e���� I#-�ta	�~yҏ
�'������E'm:8h�m&\}�A%��@�b�� cÇ�f�1���S��+�*-	5&Xx0-�&XE�q��@�lՂ�#�<��Ȃ�0����٫8`t��j,:�"[�P��M)��4Ґ`�E�bXPv*O�橲@뎗b�Y��᜵_JD��S���t9��7y�i�e$E=;M�T�q���a�� +���&⟸�1K��QS�o���x�U TN�L���	]�����F3[ H���ԹH��I{��K���;ճPq'E�j*!�蕇�bA��Z,s[j]q��ғ�Vm�Q�W5�b�W`<�aH��r]ϻG��)Z����i4�Y�qn�M�L-[���#���'�6e�$�r���W��<�`��%L���W�P,|>:���Cٸa�@4	�(��R�G5��[`���d�jB/y.�'<x5���]�(H��	�> �40��2Cdi�c��h���"�I!h�9d�9�p�&)='��H�ן6KtE��/ n���땨�90;���RB�bDTLx���>Z�Ĉ#�#�o�I7|�
�9�]XN��s�H
��|�gp�c���-@�Ľ��P��ht�#nZ�7���J4*ݨ}5)(�G�?�!CڮE�ҕ����9�9D,?-�6qq��.0��
��'����r	�7�|��	.p�=T��l�hm!�O%Z�,��E��x+�d�F�&�m�%I�\ua�7��?i1��[�Y�>ē�'ч~ ��	?g��蹣���k�2�+�a�l���'��m�w�~�Ӻ�7�ÿ<���',�6$Č�� �<����@nHl��\!����(�(�c�\�� ����0(ܢ>�4b�0ha\����"�+�%�h�p��r��&��iS3*T=%v\$��\�/yP]ra�'&!��HAn�M������
[h\2�����~"���r=�o!j�p1`R�$ ܱ'-֑E�tQ��⇎8�롲i������.`#a�Ƌ���̻s�I�u)J!�1��G8�Ԅ�l�vɈ�I�)e���̃g�jȠ��V����R&�/
�� V�Gl�~ݰ`iK,o��� �M�b�|���Wo��x@H��i��Bp�R���9��4CV p���T���:�o�0IZn�RfO�5���b͙('�0�D�W�`��ya���)ڊ���ɲMPx�F{���gD�9ѡ@(~���J ���'��噕
�0/trA��T��'I]^�
 �"'��L�3	'W���ތW�R�)��94��eRU�?�O���B��X��͙�R�h4ɔ��3\'Zm�E���݌-y�HGK'�	���6_�H혒Q�j<��2��Q���Abf	��뙵����"O�99�����0i*�(])�j��#��4�m���s���-�n��	�1�q���%w��ٹB���=��5mZ%E&�a��ͺ1� ���f�v�,pAr$�G�ܨ�H Xh$y�����I�ER����{�0B�����zG�	7k騡���=g<�!��ۯqވl��ۨ6��������Fz��h|H| v�˧r�����D?V��U�Ƨ�a$�p2�n�>�X�#EoޗmxDd ��ʥu��Ի n>S��q�Fa�+L�@��1��ܘG�(B��Ja����#=�լ��hld�;��a�)ޑS&V�c�dAI�K�:lCÇ�;c/z!H����9�Ԉ��2rڅK޴$ژ����:a�y��FϺs��q˰���<ؚa��ē�R���Ԗ|��S�P��ؤ&�6����mY�*O0��i�Ln�uې�
���Q�ϗx�<e�&șIg�Dj���D��|�'
o���񔦊&��ado�{�4i�v(��Mm�ln��I����{Y\��̭VP�����	�|����HH��
�E/�E��IF8y\V��DL,VS�ܺql�	)xP��k����t�N�gDp,�P�f���E
�Z`�ç�1&0TA�3�6�	�cC�z�� R���+n�Ո��Y�;4���7�J"25��2�I����#ލ~��<2s#�O��T��<8���Ӊ�F-����|\Jga�?�b��A�1ʓG5���ͫ�dp*�!ڎ9�� T4x��:�Q�)pb��ŀ �:ݹ��R�U��w�0 �H�$!� %��+vr!�P�#��sBo�53��1aږxP���3�xB�Z5.��8Cǝ�eC�!�b�G:.�m�¯��7u�����9`Ƣ1i��E�( ��	,�ԙ޴'���`re�6?B�m� T;wʘm+Rȉ�$S�1@�	,b����Z�Kxl;���4V*�񊑀��N嶅aA$ƵvD�h3��/l��$��GnDsGD�4T#��FL'8�Yf!�il@�m�>�<��ҝ`�U0Ƈ%Cބ��a�S�'#.��r͙����s텤Z(����K(*ҒI��L#>�P�(��t#�A�{��tS1iv���j�n����a�¹M��a�S�C�s$p���'�ʵ�"��S�^�B��H�{6z�b]�[�8�8��͎Ff�t ��� �����Bg���x��Ά`ͤ��!B�\�*�$�En�Dh���(�%#�.ے?V
Ex������h)�	
)��y oP�an�MR��#�Ը�`bۙ�9a6FܴVm��PoJs_�q 'G9ua��i�E@.�5�?97N�'��(y���T�y%L&N����>�PyD�kX�D�t+��L8�a,�E��XȆ��'L��ȃ�d��pY$Ȯ��A��]��k���.�^��#�9k� �e ^�p��2M����<�E@ٻ7 *`h�&�4vx�5����e ��k�d`@hC��_�|'b�P&`�:5&$|Xf&�s�7�,�4K�F+O�Y�W�\�x��|P�`� ZazBn��r~4�[���
XpAr�ͯC� Ao-��	���<:��jQ������Ƃ %�D̮B
��g�QEjx�� �J8
�=zT��!��5�K�����=^�y�(Ѣ;�H����P=^X����k��3�ĺy#j��H� b�$��4te�'O�)�����
�.�Hܓ#@L�D�KXGDh
@	�2nx�B��H��x��ħ��,[��A"�Β�/j	!���$3�\�a�5�P�@b�,�����+K��h�3%�������伺��:2ax2ƣ5耬�*��8
�|����DM.R޸�I�dB"���+A�Qڟ�2ݴ;�`4���y!d0B��φ%�щ��
�@aQeΘ"9�`H��1\OV�#���?���@�-'�QI�c�i�*�*�㕼t4�ZR�[�M�PMR%[�n��N$ZJ�a��lG��,A��NF��T�V�?^�]�d���M4�z�@ax��j� ءN�`��q��L'�}j�c�L�0:�k��Ʃ��bZ�8���$���S�����ܛJ,�Y*��\�L�<���<!s� a�T��)L��~�aZ�'�Ԝ�&@2E$̩����P4���j�����V�t8i��M>""��8�f	����)h2����Fxj< 3���+�8�F|r��]XF(cE�Ӯv�pC򡋝��Y����U36�Rw �"����jX\ZB8K5���s�T����u�5*�vQ�5 �&9P�9](&�6Ű��^�}b/�4m��<2�'��K�tcु��He��)�"3x��dH��Z����U�n��Js�K�@;p�@	�y���`���u�]/�NܘV���0>�Ub�5A$�0���2%�Ȭ��dM�M��E�d����؅�I�2j�0m�E�2`BY���Q�DDn�T!f��@�(T*�ʘ9�J�I�q�����BA�������^h"<9ᫍ�J�,�ɳ���b��ѧ-���.S �𪣪�J���y�@z ��Md�9�U'x���g�#!�P�$�^�'�� a�בX
tp�$&�4�Zu�X��j1�u�F�JiQ��I��!81��[`\��е1�NE�D�ق�Y�5\��,
i�6Wp�����p�RE���''��g-�4/���a�$u���}�0}����<+N$y�gЇ /���ߴnR*�ᗅ
#G� ��4�"Fe��s�b��g�Tqڤ����'�̜���#�%�ҮǒC$���oԒY��l�щE��t 9t��/J�B)�E�˥�F(Bq�ƐF/���t/�Z��x�QɄ#����||�Ab9�wi�0��$�4 ���#B�	;\�awT�2�$`{ @ɪF2�uy�A��tT� T%&od��`o�z��QMF�ER}:RF׋�]a�ɚG� ��'K��w��I�1�Md��i��/y� A*W	ޖ���&(��C���w���r��}����� ���N� q�ʌM�m��BM�Gd��d��1a~ҁ�
�zؘd�̻t*�X��K�8���F�O(ʄ;��� ��pპ�j��t⌸r!�%@ ��y�ݦf�@X!�aՒA���s!)���p>�2��%*�(�y�Iم/��-�s��yA�%yDhY�EtXm��	�!9@��7D[B�����T-��1���	|K�94ș�����f����S��*����@�J�9��{R��/8�HQ@��^�<�$������S�U�b���4j+#tT�HS�H�����+эL���r�ǔ���E� Rf�ۍ��ƦT$��@�j�Hٌ�r��}T|U�wb�5��5���X�%|�4�_�8�c�Ɔ�SÌ]�6�U>k��2�?if��e�6�<�QQ�Tj!ӄ�L[£>a�����z�`������˱{��3p!��I�l;�i�1��0�WNK�
e҄ �7r�\Q s�
�}��s�$H�`�i�4��N9�N� 5�!ecb���|k剌�����4[��T��s9��D�-��=C7JB,@��f�M'"pْ�ߣ"4 I��Æ/i|5��b�+��z���5OH8d��O`*�i�/vQHBh1�~m����a����C���wk�����W:�<Yt- y���Q`R�J��u�bM�;��SB�M��e�0��5)��s���86) ��i�	��U��}�)�,dҶ,07DT�rR4:�d%+�� �M� vIPi��"JXp�����2��pBzq�E$"��Xa�CsA^��d�? �\ �g@��Rkh$)�,�:H���#P�EB�`q�	�Vb�?	�#���g�I�Cv�jÎ	T�5��4|TN�yԇQ�2� �8U��
-�u�g%��D�*C�P �!ː��6y_V�)DgO9N��� ԨM���`k��L���y�HMZgf߃]���X�ǜ'^�ve�Wʔ�rn��'=�0�r��9]-��oX�hgH�i�lQ��Y+���x�h��ff�d��鱪\�v�N�ѧ�W�mlR�6,P���7m�"Ӳ�B�� q%d �򎗮6t �@�[/u
�0�,�h��ןx�k�:?\g+�8	Q��!C!JΔm��L[_2L@u$�K0,����$ZƢu���QL �TB#I˘c���B!L��<�L�1zK�U8�Ιz��|Y��I�K��8��� ���w
M�D���4L�|G�E0 ����%н <�P���	�`)�G�m���A���#VZ��@�V��'W\����׀y���o ��x���+�:��MO��Q�oF�l���âo@!3>�����'�j��f�>(�(B##L�H��yZ��F�o������ � 8$DE�=^���BEV:.$ձ�S���5E�,�V�!��O���ɟ�Y[H�Ȣ�D���S�M �S�%
�[G\�	���i�`X�g�=AS����ub���fnM�K�E��ZDT�9�ތj�hT�Էiݚ�s�銛8F����d���SMI:5����!�..U��(�*�)?����XS����Py�!Q����e 2� ��L�I^@�!Ă2 ��sf�C6�ؘ�TE�fJ:[ �>d8��=�&3�B ��	��] ^���$m�v��-�2:�,�%�Ū-1Xq�f̆{�N4����]\��R#զo�x����1?5�RlZ��k¬�3n�e�ѡ)��n!�	3Fh��"$�5�f�7|1���y:p�c�-K�������qL�a�'�G8�Тd��mm� Gd�ug7�<�҆K[���ڢSb��V?A���ŉU����
 A�듫#�TTs� ;�8��A�:�'8�T+Eb\"g���e�'C8�ђA�Q#�9�!fI�Y�h��٭�H�j�_��a�쒢��A�C
;��t�ݴ?N�Ijt��:j�q�uӱ�֤��*i��x�A�&M�5a-+ ��ڠe�f6�{�d�T�H�"P�L,_l�3�4&ʭ�gM�W`!���F�5Zjqz#�\j?�=?ڌ��k3��'{z��&5$Ρj���(P�bO��qJ�4���D g�&��Ш"lOܐ�Y8d*���;������?A�֬b`�'@̬��K>i C'Aͮ��O�A��O�,�ڱB�E�$�I��ɱi&�B���V��<�vaLM��O���&��-@ʖy���<����'<zYQ ������\$'��Y�-O
�j#�²s����N��|G(Y#t$�8���%$�(K�lj�<��;h}H4��)�.��Jdlgܓ_�n-"&�3O-�"/�UJ��@D�#@H�9�"On�U@PMh�
󁑇&�9�3"O�x r,L�GtfRQ�x{���"O�X�RBF��aG��XܪuY"OF��B	Ϟ9��%�v-�"O�pq���)��l�eN؎{��)"O����<,��A�l(N�X��@"O<���
��Z؊��dϱQe��"O��fe�����c�-Yݘ�"O��w�G*���w"\�P��hl"O�W����ȗ���h,�W�D�<����"+&���0�����F�<iU$�)V�A�$ثiOte�G�v�<�#��8>#�l�c�l�� ��H�p�<q
/�)��ϪvB�����Uv�<Q�e*z�6\���YH�r��@�Wt�<�c�ǎO�J�Z���*~�r�HRv�<IfhԠ*#�!� M�h���"���p�<	�� �BD@H���0d(t6aV�<ѣo�D���M�2�h�f�V�<�En�\;M'/؆��qЅ&�Y�<q�I��u|:����8;l�7KR�<�u�S����O l��8���LH�<!p�j�v��Pχ�**2ܱe*�F�<�L�$=�(Xqk"[P�u��k�<���^�D�X0C�ŻCm�.��0��d,�a���P�PRŰ@獺M2��ȓ0��U�BR�S�2��C̕5~@r��2��耥���C�L0$�<�$E�ȓ.�HU@aNR�D.�3v,�4�ι�ȓ8�	��
X�}�}�����9�ȓAT�M��&M�.�ҧȎ-,�p����Pc�b�W�t��a���8>���ȓy�v@+e	ɦ`�B�P�N�ȓOF�%���H(i�
5�b��� �ȓ-��Tp�)L0VD�r�J4]yF��ȓr��Ȋ7O��7BR�S�_7O
��7�� `�_(�CU,_�j���C5t�����0�#Dn�.B�hQ�ȓn�V���NB.�kB*�k��ȓrB����X6�� #�	��t݆ȓRQ�ɐ�l_�<i���~��I��u���:��W?@a�eF�<LF��= ҵz�Ջ(�Dm��l�3IT���f@x�b����1��.��m��S�? ��O��z�
��6�JA���B"O���L�U�T�0S =�L��O��R�����O�>͚�C_�Z�4���A�-��pQ',D�K��XC��)�e(�c��	WF�<A��W!y<�͒$ܙ�0<y�J�&A��{�ՂI1�P��oX�D�v���\jV��$nķ<;�q�eL�2t�����Կ'�Npۣ�'zn�E�J�q P�j�G*�8���~d�)5�r
@�J.���7���p�Ȍ�Ao����!3!�X�B�2Fe��dLl���G 8�=Q�(g\v�F��k~�)��H؂fV�p1�EmǮ	vbkD�%D�	���� sƏO�nyi�)ݑ�(`�^ 6n�Рt�וR���3�	}��j��ٰ:�HQj��x}6G}�Ǌ�ޞ	ϓe�\��G'�3v��B��޷Q��Åi�=ckD͠��3Qb�e3% +�O�L�t�^�>���¢oO4H�4�'v�]�c�٪-���m��Hq�I�>Lp���?��ӝ~jn���K��W��%/�oq����D"L�rr!��[�d��@�3�DPb�.#�����A4N^H�!�OD��-H�A����}��,xH�t�LM���`
C`qOH4��H���OOByrLû;9R ���Uê��āX8����$�Z�}�ʘ�V�.$��G����@cfO&h����dF�VO�EcA_� I��3�̙�Re2�{�d=��Y�Pc<�;Ud\�3�I�dH: ��As�F�;Rm\�2T;a�T�HA��,+"��t�T)@@���?!%h�5t��p��T	��S�L=TDH��ɜW9*��$���ٔㅅ `��)�O��qQ
��H4@l2���S> ��4ޟ󎞉78�q�ӯj�MS�&T�i���e�tMcЌ�7��Ekç��Ys�Oۚ#�ljV�2��s�Ꞵd���9R��d���ySHJ�|z��[�'�x 
�J6��k��5b80!1g�T�F���9�� 'cZ�)�c�R?��LN�o(9�ҮY����'c�)�d�9`�hL�DnL��wCL�HQ�I���R�@P��Ď*}3�|�d%�w�R�:�j�nM���L��y�l�Q�Rt���5�Z̃��876����S"�u�a�=.�I+N��e"mF��p�x@N�M讱��h�E�v rW�<]�x� M�jk��G�O!ug����φ� ������J7�߾Y�H� L�in��iݙ�'�
$ >�τ�+����gk2��T����X�V��ۊ��V��I3Fp�k	FV�s�	H�&X5F(�M
UD��'�}�T  �M��腵O���`UdN�h�6=���v�Ԑ���Y��R �y�LʽQ��Ĉ��Ԉ�
\ ��CE�`�	M���ژO�*t�������1
�	´�[U�O�9���R-P�@|+�OA��M�C��YȤ	�Q���i����E�;w~˓{)�=��@	t����F�2k2�H��84*�v��Yj^!1K>	VnGZbL	af�0�$�s�­b�t���T�P(r��T�ͣR�@�r��2M�<I`UB��J��0:-O6U�D�\=2eS蕿R�^���J��ReH �8�K�\�x�@�.�:�6�Ӊ5�Pi� `��r�X�����ʄ���wR�����͑9��3 �*{W"�7��;}��8�S�2e乢g������-8#�t&J[/�h�a���+�̲���f��]��j�d�"�.Wf�t�ñRҾT1�M�sH1H�w�H�� �!D�R1�Q�Ňw?��!�'K1���f'.��O�y̓g$$�����:Y)�qS��� ��)ғ��H���&�62��J�� ;��q�dh�j
J|�n��P�1���V��_�%�Ý9P��qH�K� [��!��Ђ��'Y��� 9<ƭku�]�q4��Xp%��e���� U���Crd�D=+ ��_xJ޿�ē�*���=}MH�x��i�6r�I�W�<d���S��Ț� ys�'&~	��#v*�� ��	���5~�y���>g����缫׋C�Y0DM�cR5k��0�B���%#�!; ]���>E�H"S��Y��^�<}t�c�͝3k��j]^<i�F=����f�ط��&�
�z��^�j�u���бCV�d�𑱏&Q�O��#_��اu7�<(l�CR�q� �Ц�׌9^�u	��:*x Š@�Ék�`��c�^�5 Ɲ�BGQ�	�8�D}�AT�^��6J�.�6-�V"���'�XA��K
��*G�M7W�n@�f	����x��H)x���1@��z��r�i��b;"=� �� �����⍨bi��6�x��ϊWM������.���;#nȃ"�� %����e!�E0vd�%	�$՟��P�;T�"��w�L��n�)�� ��$D������su6TYdǂ��\H��/_�=�4qH�'��Eu(̃1OD7�셲�	w|"|	�ǃ>�H`�A����ʏ��
�CG�_��*����<LO����/�L�m���Q�Sv<� ���T�V�y � �E/�Eq�M{ JT�z�t�� O^�,�p$�<ړp,����]�qv�^=?%���<2N�<;/��sѧ�8K)�i!�A2%����#��;}6���	V�t�衢���4j��F�HR�~����'�V�qd�7̊�sW��e@T��+T�Aɪ, CL�<t-�t	�DT)[�X�!��
�1���#��M�gAP���whư;w 1H
�`P�
]�Wf��'����D	�5y `Z$\2M�΍>8K�Lc��'&D����;����3�63t:L
��N�_:a�Cnl����.��&{�f�a��|��i���4��IB�FhT���H7K���O�)b3*N2ZK�y��`��t��� �o�ee�����M����PU��6�Hp���^�������
S���H�$�RzX1��øAD��"�S�ԍ8���3�>�D �-��e-�
Wlp�	�9DT%�!"��V�ޥh%��}L๚5Y�#x޸1�P�����_�\���"��I<l�+ �ÎTmt�#�T��29J�͈� C�dI�)_���� �� Ոt
P�@���l��47�ZH	�$��S�	����Y'&�pQ҂�t}D��ȍ�>�.d%����H;=� xYr��&*VMz��D,�����o�'�x)�"�>پ$A��	g{�C��f$���˒dzR� &皲�!�B޻<ܲ8y�'�ex�{��c.�� ڈ�U-R���Y7 G3P@}�#���HH@�b���q`(�Qe�4;�ʔ�DdխS���qg�G�WLy��(MD����}hEI���o���q��	~�p��G�f$���
����w*ʓ|夜JU��%4���gΔ���&�*Rw�y3�c΂kp�x1�J�m���j��ܵ!=�4�&��O�<�毊�U{X�8E�������A��� nEPB	Q!�*ʓ���p[��,y�.�
V	p�S`b��r��1��J=
�<���HG=+�A�\�;��Ի�.r��+����v����ϊ<�,�� H�</Ё�wIߠ@B��^��Kqn�}��'��*�<;���kuOS<G���E�ܢw$���#�X�R�>��e��*�)��84�H�2hR�M���#cU�F��#_Q*����j9Z�rq>�*�Ű�D��ǀ,<��US����`�p�ULQ7,r���O\�Cǒ	Y&�N�X�u�R'�-?��}D�d�p�����A'H'[��mq`ŕ)C"�l	�G��r�P�u�_L��J�Q|��D}G	���1a	�D@�h�ǉ1es��˞����<	CG߯}qVlz�ЇR'�6ز8n���O�){���
>(bx!�T#��JRay�CU#X��P�G��� ;���c�|軧�g=�庠"E_
~�#�F�T�q8V�߯
%V����G<a�~��W%�O�� bD�Yd�sf�ڐ)�I���5��`�6]�BOmK�o�"i�ح CA�7.��� Q4�$�&+�7 �q jW���#�KA�Ź�oR����OY�aPR��9��QjQ��-8���a&�%��'!�%��g�sU�\H��I�=�:`���Z�Zv�Z�EH�0��,�,��)�=˕�-w_�l#�H�?�4|��;^'Б�W`��=��d��JC!2���@��zbT�s+�>�>*ϓz�IGG4#�Y�FJ]eh��လut`L3Т��\m�d��&�?,�a'��5+�q���j�����E�;���ӣ'�fyB����r��2�' ��؆L�J��]����>�����fкX��S(O���z�i/(y`�IV-K%_/6��4:O����'VZ?i��T&R�(J�tQA�D6;25ZHK)-d��ҷ'
oܓ2�P��SE�3*�Q�iыAXNe9S,U�<Sz)qC�[� �Je-� Kj��~�"I�4^��'���t����XM+�j�R�)�As����yݼ9e�>t� ���X5����K�2P��Ka�ʢ)���"��a�2��"�Xܡ�8�\J��Ŵp����R�E�&�ʢ�U�e	VX#��-f��Y.*,{axj�5X���`ƅL>1x�y�邜��$�3,c���3O�:H��3u���<��42~�e	���z�"U�%��f$ ��#JP3����6Κ�MQ,=xf""\O���F!�J��u��.@Q�V�ʹ-�xA@`�-UNR�BT��M�֥/	et�%ʈ�AV��`-�i[b� &A�+7ō�w�\�1̔{~\�Rh�ax�X�r\!sP�0rV�]�<}�A֝@��y��l��`D����R�gf�9To�=�~�1ƀ�[�(Y�!�@��u���W�<Q'�:&��q#���I d��1l�[�'ڤ�C�]Nr֘�f틧9�� �:9b�m8�!9�Lp���-9��h�bư�СLشĪÉP�b��t f!,�%�h���
v����mV�+<��Y��H6c(�-���[�~��cJ�!�d�B]"	~���uMW(9��a�	4���"��b$e9��	�)N�-�	O"7tY�	�r���Sz(4m{�◤j5��A��5O2����R�g/zE�F��v�X��$0i{BV&n?���;J֭I񥁅+P�ȧ�Hk�F���	>TAHDS�
�  ����'TK)4���B��Uj$�S#.��y@�ܴz>@HXT��rg؝�EA��&�F@�Gc�C��T`&��?����e��Z=����On�'������%~9����l<a�I�_�ޕa�"�C��AbaB)Ei��
'�~)8�H��'.p�2Tf�,v~ȍ�bE�ўPKg��$T��ѸCkU� 3��r��5usPm5]=�L�[��H�1�
}���U������9&8��"#��q}D}� "H<f��@��U�E&�YB�-��	)��3F�Nx����M
 �\�k��W �Y&G	�%�Dc��#�(��Ȭ���WVc�FL?f��)� ؖdz��]�*yb�	�e9�C�e�-RC����ت-�|�B��G@�"j���/%�t���h�|�2���!W���j���i�t]��,F�D#6)*���#�\�vV�j�l�jB�OT]ɲWz���TLA,m(�tr1�	O+
��2-�><�� ]�F<�d���)\���(Ћs@��\�p���he��L��P�AU>+hЕ3W�L�R�&���1�# �]*FJ�-�P��"���m�P1:"��$a�ֹ�ID�+��9��O��'(�A�ܘ)�F����S~V�����6�^Ay""\�G��A�'�O��0?YqA��$�Tu�$�	m�8��߅		�-T�I���v�M���e��Q�!�B}�a�h�Ɂiļ[�9|þEa�G؝f��\�C8�H"C�H!?���NJ�& h��W�FkLA��n�_����$u�x5xdF�>�L�rP�
�%
t:�ցCa^a���h}B�B�F��1dt�2 B	�|Q)C��D�]�����
ѽG`!%d��Z����}TA���c���9XF��G�O�B���H=7I����Ď~6��>!�ϷG����dkPf�,\��Q�^`pch?O�iy�iX��eGǵ@��ԳīЗd�"@�H�Xrz\3��Ȳh,$�A$��*t@�L�7�J8���	E�Bɉ�G�Xb�0�'�Tpj�o#|tԅ�G-�+�Ʌ*��s�\��'�޺�r���]�B@2GO!qЉ�wM[�(�8��w�v�@��8u�`AX�@ڝ��a�(O�!�E��jplx��!C<�H�����.��^����Ӳ^��h���3&���!,NH<1��a�r :S�!K��D��T��1X�87�ñ�~"�\�o=�� ��+J��� ��|
�m��c��PHb̄lW �ϧ�h�V	T#�T`�ƅ�>�"Q�Ј�F�ʤ�3��<yzȻG�"��aHT�͸8���0�F=9tn<�@�ZF��<����򍳷��$T5h�zf햧9Z�+�޺xIb%���b�pE�5����7`ЦP2b�2��W�?V� k�HˉL4���F�I�s�'i�����`D"Z,���@`��{&<h�lS�x;>M��E�Q��ƁB)��SQd��c�1�ȳl:���	��H�]0VN�rX�$�F�C-��51��a�,i'eI1h���c�-W���/�Y�R�;�O��r�Y�yl���4�0kp�)��*w���7F�?I�#h��*��5z����Z�>1�dT-�j!�r��'H��Ս� IN9���#.��*"�Y�*9Y2ĕ(�d5��4B�:q��eEz"$)��E �QH�B��Ҷm\R�w#*]|Z�%Eoꂢ���m�"�S
-#j9R�:� 4#g�B99{�-x�'�6-{��rq� 3ue"��#��!tH�g��cF�x̓�#��C�#,�3cc�6~��̂5�E� �I2�871e��N,_lDh��@B�&)�#��4|���]�0����x�����"`��nOJ�㷨�+�N�qA�N��^�!��j����$D�}���*Є��{���ڶΊ�F<M9�
<B��׉X(i��(t!S�`�j��D�~����Fn��C0Q9��W�G���gN�'1Gh=�@��7|>�0�l�P}R�Y5}���SA�+b���+w�'��uS g�=f��O���ٱfܬ3)�xpc��"= 
�p#Nb��Jc��0����"�-1����,2+�tP3K[�>'��@��ݦ2�51�B�f��"W�t����`k.L:S��u�U�9���a�?��K*
y(u#�0�*y�/�	t%.��k�#x@�K�'E�~� Ǣ2m�rʧ�;qt  a�Hܓ:� ҷ
�b�RIc&NL����3�aX�.�����g�!0HJ�%�ź��A`�^Uc6n������خ.�<X�A��>��Qb��ٖ�R�'���P�C��'tc��;v솈_(p{�
���)_��1 ��t����/�b晐�D��$s�� �>���"v!^	+WB�Lcݵj�|��M�GR> ��o��FJ�3����$/}���f1���iyRk-e�5��j�1��	�O��q�F*���@�
�t4tݣ��j��h�K+�lx��+��>U�;Y��%`�ׇaIp��%�5	;����i���@,H,t���F���c?U���Xм�e�/Vd��bX#6��R%%Q�ZU��zA%Ƌ(�!J�!ϬWW�g�'餩y��G�Q�m2P#�!��0K��Z��~2��f�-���S�9OΨK2iʱ&ꠡa�/B��4��@@$}�8�Ѯ��M�$@��c؞P↩� �����I�L����>���ǋ�lO$��Ę|��mM&��Ԉ�(i�ܒ��*&F��8s\��+K�p q�1�	10A�б�@R.]Zց��NE��G�2��1��ɝ,S �}x�"O�pI]�앹/ z�"�57��ɲV丌3���=��S�O�:�!�,�S���1�iW�l���'D�샱G�
N�ȇi��H=X�{"-�G����	�s2%���O�T�6�$k�0�B�	�]�6���kы=�Xu�k�#��B�I�	e���ǯ�6�:�ѲfR�C�	�^�
�� Y�x�U
֮Z��C�	@��h���Œ,�ՃA�j��C�;t���u�X��4�ʅO[�nC�,C����3�я̠�a�.AiC�5*L1��f��O�����ٻZ��C�*�ȱ
Յ���^``�)ՔO�rB�:����u&�b|"�C<r�:B�7���d�t���*׫Q�1�C�Ɍ,�0ԫV�ԥ��5����fu�C�	� .�Y"@����h4���_rC�	�xN����U69�j�����][C�iS6ȑ�ήG��]`�$��6��ȓA��g[�T�>���\��]�ȓXlt)pTJB�48��V�T�L��t�ȓ����=0�1�ǦW �:�ȓF2A�.A�H]�$� t��X�ȓv\�3��	g4!��MK�
��C�I�a���ɳL�"1����\�uG&C��BIܼY��_�b��r��SDB�	�yw��Q
��ht�q����C�	F��d��Q"���;t�Ò}|�C�	o%�Q+@M��st=ab��U����$�n�.DS�O:X#�`�&��W��0�VtqO���GC:���a'�0����}j@_�2u����!ɺlx�[%#<�� C�z�8 Q��M�r�f ��'4B��3#�Ӹ1T;�bc���K3�o�fy� �
b�\��sP4�0|"R���i��U�=���� �8"4��A����I��0|�ԋ��3T�K�E�3e5	ZݳL���#I�nH��ħN�F��ÍC�BX���W+�*H�&�Xy��)��.QZ,��UF�"���
�@���<E��Fb됹�%�ȔP?�����McSL=�S�OE�h��֑7���zGk��.1{G�ȶ �hqØ>i��O2Ԕ2c��?@��q3�!OlU�	7c�3W��$�|���Fe�0|���U�z7Δ�b�;Jo�L3�B�
+ZA�g3O����F��㸧�OJ"%	![��d�kv�� h�9I��Q"QnF:f�)��Edq����YݪQ��㇋H���AdV>�,��O�����TO�W��<!�ؠe98�Ur�:O7D6 ��)�~֧�� ��*A*��)��=cŬ���z�>�r�@/�0|��&I�C3ځ��	��a��ԡ1�OT��>a��Щ�'j� 2$�3� .�B5 X8%�DxӇnk	�4s4�O�-�'�O�H��X�.G�1��	*t
�^F��0��O0��M<E�Th�Manq)���2�(,p�+�$�y�VW�D4IHa���R���i3I=.�� xC�+;*O��Iش��b�b>k���n�nYxQ��79�j6�*?���p��䢍y��)��q@�9S&Z.c0Lʂ�� %;�$�ܟ`�"��S� ����D�b� �3��ԓNL��
�Nʓ�y
ç
�KS)�<���A8��䚄���q��I&�?�J��E�� r��ObPS`c�
G�F�i���e7�)X�"O�5��F�JI̒s$Ķr���S"O��9P� B`������< �"O�E��]~}�Ԁ'a[uli�@"O`�Q� :]D�R1�S�f J"Ozpp��t�*�rC�;)zL{�"O<T� ꛉLjH�^�	:��@"O$�� �C�B�rH)2�/*՞�B�"O�!b��lt"p�$��#'�Y��"O��JH�b�H��׍�Z�0��p"O�`[S+u�RD8�*���&�S�"O�p�C�1
�Zx�4�N�>�6�Zv"OlP�F H5B(�Ѧ�.r����"O��KG�;�J5��CE�U��A��"ONA��eD�"&�l�@c�J��!��"O��@�)B���IK^�Q�e��y���@�r�X���:x�	��7�y�&�[�Ɯ�"F?*n��U-M�yb��X�q3��ש<px�1g^��y��~z���E��ۤh� �)�y2�M
P]T\�����du(a@-�y�J��`��*��>W0���%�yb�Щ-p� J�m� �y��%�)��D">12U���y2�X���$�P��1j	���E*�yr+I�Pܔs0G�-3Dx*ׁ��yr���B#�Be��@�l(0���'d.��-ӈF1
�	����d.d[�'��� 1
ɨo���k�d���s�'�F)�� �ZT܍*v@�F<��9�'Ѧ��`�U�Nג��5D�DZ*��'	dx �i�N�>�u,R!-¶U��'.��CKF��v��$�� ��%��'��0�c�l6
�2G�UC)��*�'�n��j��5-FYI5ΗhS��Q
�'�N5R�G��;�v� �
Ǿc�pU�	�'��ȱ0��1:]*q�6(K�(����	�'����
�b��x&L�o��-b�'c�b'�� v�a�$I��4%��'��d�&���0��ذ3K(1�Y�'�¤� ������a�@�}��-��'�|Y�A�ĵ%~�����s������%�>X�Z�:�j�
h��)��,�]�<Y�eO�1�$�"7��c2K���Z�<�p��n���Z�Nǋ7Y.;�LOS�<�e� ��1#Z4A#� �M�<)C�ɍ-&jhA�#{�X�'�H�<Ig�T�6Z���C.�$�%OK�<u���驰 ϩl[��R��q�<!��ܿ2>Ցm֧s�L��@��f�<Q�*͹m���ʦJS-Ww����cw�<Q�Ƕ7�����Ũ<F���R�r�<٠�!h����M�n�1*P@�p�<�p	З}�D3N̠ܦ�2B�q�<��5`F��I�2�R����l�<��m���FD���1^t��.�f�<� ����΄�RU�r$m*��q�"O\�u�G9jB80em��%J(Ё"O>���̾J�zх�
� �"O���Ãثjf���d��6�Lq�"Od�r%�0[�fT 3ᅙ�`�x""Opաv�v�fD�t)�f�>y)"O��(4�x�hj�,g��9��"O����'x�0����\��ԣ"O��G]�5��rD��[��"O5E,�D6� kE�X�,�C�"O	``e��T�c㩙�]�x�J�"O�Ii'�ب%/^ݑA�B�(��E`6"Ol�h䬂�>Rn,y����`�UI"O\��II/0�a��֚#�ޙ!�"On+�AԤi�mWn�)��"O�ስ�ս�֨22��,A�q�T"O��(��P*hz��A�X.��"Od4��*Q�S>���X2*S����"O�aPF��)A8IaT,χ_�^�r"O��gC0���;e�6R����"O����hؽ֘�uJ�;`X��5"OX�� �vI`��iPu6�a6"OX�����z�豐�i��hn���U"Oj��V'�AИ�FnM9z�
M�p"O@�R�^�%���¬يQR��S"Op��T�D�W?�y֥ߧ]C� !�"O�Ԉ�ՋnD^�� ��bG� �"O=%�0P��ir䁑�oL�})�"O��R�A=�$��!U(��<�"O`�V��+Ts>���U/^���"OTY�R��Q���6Oå:r�Y�"O���ֹ��j���4|V����"Op�n�
y6�,[��NE�mhf"O���`0��iIp�J�p"O��Q���%lK����Y	xP�@"O���؎1*R[��P)dO4��"O�X��(T�.QP�+� ;����"O���`$ũu?�m���!K�IcV"O.�ZDoR9U.�: J�=}I08�"O,}i1̃�bY~h�%"	�!I>�"O"��tX�	�.��#씒i¸j�"O���g�&ԥ���KeT�B�"O���`�s	r1x�	\^T�"OHy�b`Z5x�ܸ����e\!�DBN;b8Ö?D�@���T'9g!�d��v�x�p�غ`�ѓ̛�WP!�d�F�M�b@��z�
�	/19!�D�D߼��w#Q�g!4��ߡ36!�$	�{��:4@�;j����J�!���U3���Ă,�(\��o�S !�Ă�0��l��K�"`Լ���Յ�!���W ��Kʩ܂1��X�!�$^�7:�	z2/����ӑ�N�!���!+�jE5�){�+%�%�*���9e 4�W��W����v�L�#�x���&<�20f��%���l�9���ȓ,�A�6a�L��F�cl���FIvm��C��,�-_��m�ȓRh6��3�C�( A�!)H���ȓ[>���B]8VY�F�RI��1�'�`��]�6O�b@�aTA��'閤�E�F'8��=�p�]H���J�'b,�a����{�LP:WN�AR�́�'��\¦a]�U� f 9� -K	��� �*��6t*��PKS�P���$"O�Qf�W��Hia���lc��p"O�8��5 	@�sQ#_X`�"O�8�2�K*V�����>LtEZu"O�)���9� ������E0���"O��z��5'-
�3�ef$�0в"OT!{�!|��!*ٿK����"O<l�P��29Qp\ٗNP4>����"OT��R� �De\�`1� L�x$��"O��Sl�> ��PR�,�R�Pi�!"OH��V�T�v����R	�~�2���"Of-0Λ"/<h(V&�5
g�=BG"OМ� /�8��`��Ǜqܡ"O�Tڇ�ϊ$���g�)U��0�E"Ot 3��������9+���F"OL8h��]<v�PE�ĭ��4pb�"O�3�	�	VL��`�	�$s�"O�H��X�F����` Y3$��X�"O@|(ǥ  r�A��������z�"OJ���2<\䐑��C�L�� �g"OҡK�@�hD����A�8�r"O:�{���M����c!�)nεJ�"OB���a�>y� Qp���8���s4"O����cT�7�(����?AJ���"OļyW��(�j�"A.j3 �H�"O̸���̬4�f���C�.�銶"O�� ����㣯ĶE��H�"O��2p'�m�<La��7X*2u"O���&�@�qPȚ�K��qNR��"O6�Ú� ފ8�3� A>d��"O0�Y(u�������t₇Ec!��D�H��)����|Ra�3C�!�D�[z���;�ҕ矦�!�$T%3>c%F���Ii�I�B�!��-U� 1z��Yw�ݹ�A8>!�䎍S�&�ӋM�qn��8!�ְK���,	m�`�QB�#(!��2%��jel��L��}bM

!���͢�dĆS�>��S�ȡN�!�D�P�j���?dbR�"UJ�:�!򄕯I�D]�� C�$�0�;4j���!�d�@^�;�U�<�e���E�!�D����@��٪�3�� n�!��jD�aAsB�:	�>��,�t�!�dC� ��a��N�*������{�!�[ K՜Iq`��4��� �g���!�$�_�IXwk*�:��$��=:�!�D��%��ɔb�(<=qTHT��!��C�8`E��D�/'�EJǇ�$!�ޅf���͈�"�N<��T��!�D�RhX�ƭ��9��ؤ���i�!�		��qR��ϔl��V��!��<�l8�r#č��Lz҆R�K�!��K>m�s�����ͩ�fH:2Y!�F!6E�%�/�8�j�v��/X!��C��*6�-N���(5�1nR!�/�D�%C
G}�]���D�H!�d
2����B�$�BQuR31!��L�)������M.~iz�V[($K!�DI�A��J�_/[f���\�^�!�D��W��d���E����C�@�
�'K�Z���a���Ç�D�k��'�>��ЪJ�qx��Ad�����'iJ�y# ��R2F�f3�l���x�<� ���B2�(tP7�	�>��(B"OBD�bL_lt�o3)9��9"O�t���^(�c��](>	3�"O�����a`���U���"Of�[����eE���)��%2�"O<�Q��v�z�uiK�b�%��"OT=x�A��6	�(R
���ړ"O�Q0�G�e����1%�%{����r"O�C����pqjH�g"��R����"O���g�<��<��� J��iR�"O�t����<N��9G�҄?6�ȋ�"O8������\��oö=�A�"O8��/�\�8�EN�+�v�"OTu�
   ��     �  B    �*  16  B  �M  SY  e  �n  ]x  �  ��  ^�  ��   �  c�  ��  �  U�  ��  �  s�  ��  �  Y�  ��  ��  .�  r�  � � i & �" + �1 U: IB 6J yP �V �Z  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p���hO�>U2��F1C4ӡ%B�>��eW�%D�����9]����"8�
mS�#D�th���*��6��4��$#D�\��2~F��u
�!.���sA D����ýe������[�<�����?D�@�w%��&�f�SS%D��8a!�(D�HY&N�1V�ȥ���V&D�A�`!�	�#��yr�C>s|D劥o^2;#y�Qk��Px�K�{�T�:���(8��+�#$����>iS�'lO�m���KTѐsF�W�ճ��'�铤�$ũN���rć:5�@3"��)rm!�P-s�h3eH�r�xb⪙�j�!�䈾�Bl�*ݎzp��a2c�1Y�!��8$�N9�%�D#f?��
�#��y�!�$R*l���2�Ɵ�1���8cǈV!���+ D�
�dV�e"⼐Fip!�$�8p�,�7�֐:$��`H�;�!��vM��­�@�0��/Et!�ĚYゼY@!҃&���K�f��l�!�� ,.�T�%rd$�4�]<~!�䛱���kah�f\삑�M<+`!���8�e��2G,%s�FS�gI!�� ~��d�)b4��ci��.�2�"O�a�L�I��=@Dg�0��TP"O�1���F�nؘA�5^�
���*O��(�NB4)�xt�θNy�:	��Ms�O�ݒ��hҊ�Q Ў!�ZM�"O�������@K�ux6Q���{�O˦�l�+E�x�Q�đ2 Na�	�'٬D9e��91��p�X$>��a��'�б�Q����i�&D ;? $��'͢\"�b�^�@!`�A70uش�~"�Pc8�@SD�?(31���T�j	���?\OB���$�`s8�Xt�����I�f�!�D_�)��#��R8�$=[���F��'Mў�>]@EÜ� ��9z#Ï1�̐ .?D�X�h�%;��hK�ɚk���F D�*$J�)" � I�3*�q'�9D�L��l�K�d<�7�1<�5xү3D��q3O��%pafӀ)R��p�/D���f��J������Ib"���-D�L� R.أ#�	�D�*u�7@+D��8R&R�2���B*^,�Tk�k5D���3
L0�,��f�1(��xC��t��=E�ܴe����Q�0�Z�(�N˖|���ȓ[��}(�h�0"��_�Y �0��j��s&�O @�B�I���@p�P���F~���`F��%�^�7��H�ӳ�y��9P�����:Dql9�F���y��N�'�4[�IE�%ߘ��E�̥�y" h�^�ڇ��5�-�'�yR	 ����P�S?`*y�����ySc8P�{��`���'��y"�U�S$�R�$b��z�K&�y��X�rm��"��\}&�I� +�y�)>1��E���O�H���؟Ǹ'�ў���a"QF�D�A$���;�"O����7��<�2��5c,dts�~����BAH�8�YPg�rhR����y�$�ޘcF�U�n���^��?qQ)=�ONa����ph6��F좱pe"O�e�/���Ukֶc�I��"O���茰+�j|����vp�d4�S��z��X�W {E4�(�&�DhC��2z��iH4�l%��7|�\C�	l��2�利@��MR���z'HC�I�)r�(z���$㠝c��+�FC�	�L��<�����Wl-s�D�$2C�I�]��%��� �X!�BE��ybgH�(�L�g�� �&�Prm����d*�S�O�<��� ({��Ar&�T
#��t`
�'�<M2�g��h5�����	�'�0`!�(��&��`ժ���� 	�'%���7�L�RE�Q$FB��"�'��h�Wl�B��	�qO�+K��ea�'O��Ȱ�H�j"�y��W�>��z���'*fՉ�Q*y������gӄq�'6Ȍa��5��Y2nϤTTh�8��Dp�ޣ}�qb��T�6(��Ob��u.P^�<a!��Vp��ᨕIF��S�GbK$P��O?��B��*h�w�ۿm U�6(Y!�\s����?s��!��$�����>��M�+�����*@�Rm�#�e�<�b�5q�������1�|0'"O4t�2�մer2�/�(i���"O������<4}B���M��!C����2<O� ʅ���^#7
��bQ��];bOx�����&PP�,[��=��( �� $���`8��2����7Z�����>+��;W�=�O��A�'^�}��(�d�X7��<wR�52��HO���&��&X+�c"�r��$I�"OJ��`S�l�1O�
���W<O��=E�t�܉k�Z(ˉX��0Bd	�:�y�: +d��)ɰ\�`�� )T���Cݟ̇���	7G�I�<}���������<IR.��h1����%"�&���n�p�<�u��0Am���4�D�e���yĊ�e�<�W�J�I%�a���
BRV�١AF_�<aTE�TԤ)���=0�U!7�x�F{��逯L`�!#$�˯[�&e��	�"|�B�	j��e��޳�-SET��ɧI��I��~��hO����Ǆ�$L�rs�<8oڅX�'�d��'�4��b�d0Q.Y�f��n�W������m� `�z�nZydN�V��0=A7�%��$o��<Rŕ�,��K�肍M��듚p?���	c����e�E�mhb`а��}X�ԦO�<q��ѷa�pz�X�L���"O<p��C�	R���y�-*g�|B�'��O�c���Tyƚ����Z4�����0D�x#� ��@�:��������d1D��!�[����g��r%p%��/D�� ����7x���ʕ3Y����&-�	��Q��O��좷��'>i�`��o"��	�'
�A4i_�f�\ѓiD�3L�ّ�A,ʓ�h�����t��|f)*>z���t+�m�!�:�1gI�>} e����)�Op��r옺i��h�&ԠXw
"O�p�A/EJ��E&��Wg�-i"O8���R A�	&e��d?N$	0"O��C	qȜ8p�!1`�V"OlUAR �;I����.	�(h��"O6�$�ܻZqd8S4�L(��e�F"Oڥ"`��?bH����t�(5�s"Oй�&ǝ5n$�`vkA�"O2�Q�!�Z�|�o>1���"O� �r�E�1ಸ��͔�/�1�"O`,b�m؜��H�&��8�`��|M��jȞU�ƍ���Ǿ^o�8�ȓRBL�j��@>A>qKv�N�pńȓP�0Z��E�
C�s��!9����ȓ�Tڰ�š<����s�T7R���ȓ-ъ�J0�O,B4^�#�a0|�ڴ�ȓ5� �+�!;ЌS0e��Smf���G�\���
U���dO��&�h%�ȓS�Pe�4DTJ�Ve����*p��m�ȓa@�����[��q��G)�,��ȓSIl��+m{B�ѳ���H
�ԇȓm*�U�#�>;�`p��S�y(�������Q@M��}��-S%ƻ'*Ra�ȓt8����������P�>� ����@�A�A�7#O�S7D��+	���JR᳢G@q`�[��\B��ȓR��;�n�iP��J�:{ņ�?x$I�6	E���L�ES�2.���ȓk�`��3Oĉ�7G�p�4Q�ȓlA���Mլ9�ɳB���$4l��l�*��T B�Rf�P�̇+D�$Ņȓ[z�akFk�7tv��C޲C4|�ȓZ��5��^;d��;A��+��|�ȓ���G��%Lժ���[vhɅ�S�? ,�T��5M�<���"8=�"O���Aٓ8.�ᡧ�7B ���"O�%�X�F�+��B�/�F"O�T� �/f��\u`�89��Q"O��(q��uJ~�	6k��&���0�'�B�'U��'�R�'�b�'���'arP�$@�[��9�,�95����'C��''�'�2�'NB�'���'��lX7F����ȣ��ͷn��H��'+��'���'�R�'���'���'�ik��4+*��'C�|/8DF�'���'���'�r�'���'%��'�t��I��[���LV�+-�?A���?q��?q��?!��?y���?q��ؽ�����K�MX�O'�?Q���?����?����?����?)��?���N���p$̂�s�:��D���?����?����?����?����?q���?�B��*�~�i��Z+Z�Ő�����?9��?A��?����?9���?!���?�S�F�)�d9�C�ab��A�����?����?q��?���?1���?���?�0E��g��A�Q]0,-p̙q�� �?9���?����?A���?��?���?��!3,KHI�4��/M.������4�?9���?	��?���?A��?���?I��=�X���R�;rr�$E���?y���?a���?q��?����?����?	P��)n��LS�ĕ5>F���6)E��?���?9��?A��?���aG�6�'n�x.�3��|��p��@�-8���?�*O1��I�MS��Od�=���ް
�Q��(bL��'"T6�*�i>�ܟ����#x��1������E	�ߟl�	3'G��ng~r9�@���j�I�}�n�	�,���T۶,8k1OV��<���i]+\�̜��$�+J�!�ь+��un��B��b������y�� �d�ȵS�옼iQ�ܳ�E8B���'��>�|�Q- �Ms�'rZi�C'M�Y��y&�M#-6,�X�'x�dٟ0�r�i>��	.l
�TFn-��aI��y���	ey��|R
~Ө�9��d.X��	�^�{7z8���yk�<;�O&��OP�Ia}�w�@`@��S�wX�CBG�����OD��d�`c1�D���`c~��/:zR�@1��88�������;��ʓ���O?�,L�����g�g�L[�N�l�J�I��M��FQ~R�uӘ���R�ہD�%n�0��K�j$�	�(��Ο�åݦ��'7����?�KU닿	�dY�pK�*N�4�2�	'A��'O�)�3�I/uXj,&o�$��(�e �&1w��Q,�&
@�(���'F��	\!-���3l���`��EF8_ ���'��7���� O<�|'ȓ#И���+�cV0	��O��}��3-�;��^>!�b�I�f�r�Oj�s�l8IAHX�Y�����)��9}b���	�M[�GJ�?i�CR�,���E��8$��?9�i��O�$�'��iMx6��5������(�Qj�dZ0?_�@[��kӔ�k�X}i��?�'?��ݿn[��pu�T8xaP͡���o9��L����#u\@�FӱJ�\�������I֟�+ݴ^�<8�Og7�>�d4$����!۾@����D�efP�O���O�iԙsQ6�9?�;��+'�PSᤠ��J?Vr��!�*���~��|BU�h�?I0H� v��b�xk8�q�K|�'N7-<4����O��D�|
GI	�f��T�A`E��!�`My~b`�>!���?qN>�O��+��/E�xxg��>�"�[�J\�x �j��i����|����\$�D�g �;����IO�1�.��E.B�,�����ҟb>]�'��7�ū/F6X����0e��BƬ�쵑p$�Or�D����?)�[��I۴rV$=�t��;'��Б���q:.�*#�i�*6�Ĝnh�7�)?�TA��6�������D�.�Q�3��2| � CQ�� H��<����?Q���?)���?y,��p�	\���̀�RhS�K�ܦy��Uy��'��O��~��Ǽ�LQ� J��Pb0�]�W�8�o���MKT�x���� 6�V?O��0`�	�v��f�ͯ1]b�r�:O�	&�d�'x�'"�I^y����#��N���r1�N�0<�w�i�����'��'�|��P�"9!H�*�ˏ�X@�3���e}R�'A�|2)L3I6I  Å
=Ɔ*e&���$�"z���Hvӈm'?!�O$�d�,��D@��	�{��8TF a���d�O��d�Ox��;�'�?ٶ�H�DiRq!�- >��������:���'�6m'�iލ�u�Ϡs-�uI1f��f���8��џ1ߴR(�v�yӌ� �+f�j�I�`c�EZsol��7.�&���H?k�ːA��< jY&���'�џL��m
�o;�QZ� ؊O�NAå�3?)��i>�3E�'R�'��R��$�#0�*Hp+�r��x+%�Cf}Rcr�2(mZ���Ş=!�q�&��V����_6��J����Ms�W��I�-���&��<1��ЬU�l�kҩB�R ��
����?A��?���?�'���Ħ�Z4kL��8��/������/�P-���Q�4��'C:��?Y�b��_���Q��J�4�蜛���4`hɆ�i��ɋ?`Ґ���Otq�b�� �DYŃA�KTҸ���F�~Pec�5O��D��-�b-��M�3Ơ�Pa�eP��D�O�$Ʀ���)*�u�iR�'/	P��%O��E*�M�}��$[ӂ1�$���-���|���[5�M{�OV4R��+P��p�DE;8�C�ڕZ[�=���uIƒO���?)���?9��{d	����1��i�I�/2�1����?a*O�l��.����'�RU>YW��[W�� jn
�P@E�-7D�ɜ����O�7-H{���I	�F�h�1�[9M���&��83���F��A�.��䛟��8Q���W}��7
��(ɶ�S4�tY���=b���ٟ���ڟ��)�SQy�dӄa��ΨOC����m��L��FӖz���OX�mR��MP�֦mP�˝�yV L�`��O���d����M3�i��B��i��d�O��3 �H��RR��8��+�T� u����1����f�t�'
2�'a�'�r�'Q哪�(!I���?/����ta�x�Dl��4 ʌq����?����'�?Ar��y�cG�6�<���\v5��N�w<p��sӼ'�����B�	a�H�I�fgl�Ѡ��)\��.J���mJ�XP�'���'���'�2�'J0҈N�y"a��˻>�� S��'�R�' �_�"ڴ it�̓�?��>d>����`�Ѱ�"�#2-A�2E�>����?�I>qEA�)+/�l00��3���0�I~R`�:g6�)��il1�Jh��'��*�>-���-3!�`����5���'�b�'����"�iTR��'%�-7�j�r�E�$�ٴ�*����?I4�i�O�3L��`��<��9y�ރ=m��O�7Ӧ�)�N�Φ�'�|�%���?uj`��I��A���[Gb��u̇?8��Q����T�'���'���'h �q���.@Teu�̅S�	��S���ݴg ��z���?!��䧟?�5�]'NS��8v��C�	��DʛFT��ɟ���&��S�'\1DI�D,�3f��15�O�vb���3,�;�(�'��P��&��D Ԝ|�V�\	Dɋ%	��3��
:]��Ѳ�C�ٟ����d�I���Shy�Nq�
���O��s�	Uq� f�-K��H��)�OMl�q�X$���$�I۟���� 3�ڰ��'9zd('�ҔK=p�l��<i�.�dQ��|��'^���wԸ�8�A�Z+�E���'$R�Ú'��'	r�'���'3��W%�N9�`4f��?=��*a��O��d�Odmڐ1h������ �4��Z��l�≁%8f�x�!#H!�A��x�-f�̱o�?�kr��ƦQ��?�%/�v�r\�5n�?pn�Y�BExy`���Ot�M>y.O@�$�O����Od��g��3S�}z�^�hH��xvj�O���<Y��i+R���'���'����O�]���� D�B9:%`�J����O Y�'�7-�mjJ<�'�b�OC�^N��3Bߎ`�$⤪J�K��0�`�#��	,O"�I��?�8��T�P���i�b�Xwjh11�]�?��$�O4���O���I�<��iD��X��
Q9��-�" @^u��UC�'�<7)�	�����¦��Ҳ�t�\�_|��e�R��DMmڇ�M�LU �Mc�'�¤=;����+C��	-.��h�Q��s'��iU��.&�4��Fy��'�R�'��'`�X>�Ydd\�u��D�#����srC��Mk��T��?	��?�K~�dy��w
(aJvI�)Q���K%C��9d>����rӮn>���|���b�*R	�M�'�4�i�"7�l�Z��F,1��M��'��qs���#�|2_������ c�	 5"|4 �EJ�Z���â�����Iʟl��uy��nӚ��1��O����O�qQ�!��y �酋|l �*9���O�ʓ ���c�L��'nBFR6���1K�
T�@��y��'�Y�4)�>|��V��<1��E`��Iٟԫ�S8:ߚY��-%����/����	��X��ǟTG��w�Z4�C�SQ6�x�����p%ДYU�'X7�[�D����O�ilZE�i>��i��L�`,L7A���XТm��9OfplZ?�M�Ժi�N�i�i�	�Vy�=à�O����cܫ#ܔہd|zt�y�z�	Ry��'���'i�'��.ߗ�e�ʖ8j�P�f^���	$�M#T��"���OD�)�|��7�z�XQ����vh�6Hɰ�*�{}"�wӆho�����|J�'�Z���1%�,-\pp���d��\XBi��M ]�03��J�$3�D�<��%�a�~ KEF�}ZP��1K���?1��?q���?�'���ڦ%;��䟐��A�[�����	M#*lq��Cٟ�4�?aL>�s[�0�I������Mnz�2(�=�\�VNO�h_8�"�Ŗ̦�Γ�?�-�<���Wy��OsW�W�m5T��0"ӄdD�� Ǐ�yB�'R�'�B�'"�)��w��jPk��[���c����$�O��d��Ef}>��	��M�N>����-)��m����	'�Q��M����?����?�@Iʚ�Mk�'#�I�-PZ,�(Ķ<�ژ�@&�A��Q�य़�$���'1R�'��'�>y�!�v7�)À��`J�����'�R��i޴4�8����?����Z�gL<l��oJ:,�����iZ��	��d�Oh��#�4���$F#)�� G���Y�P\#	�y[^4��o�s"7-Xy��O�������r_�Q���M�!��C��,��DQ��?a��?Q�S�'���ۦ!Yg�g�Du���U�♚R��OT�',87�4�Ɇ����O��C�A  X�T�a��2%���Fk�O"��DMJ�7�q���'7X�P��O��)� ,왕��""tϊ�L�$Ҳ;OBʓ�?9��?y���?�������)��J��� h�<�IG���9��]n��zP��	����z�S�,
����T�I,\�|�h���c�i��bH��?�����|����?	�B��M��'Tԅ;׭�D�:�c	}v�e��'�
�Aԉ�x?�I>�,O|�d�O�]��
�t]���ËK�:�r���On��O��į<1��ix�M��'y�'����톗���9���	X��]�C�~}��'�|r�B�t|�%�߯X��%�4��B�w�D�#�I^�ln1�`���in���[�9op�;���5��9���~l��$�O>���O���9�'�?��l��x��m*�
��ˀ�R��?!�i5��Ƞ�'B�Ӏ���'H7�P��'�����]�g#��	͟��I�0y�	���e�'��qǙ�?���� "7�R�Qe/D�I~���,P��'�i>��������ڟ���_P�*b-��l�𤚐^%�'�6m�Ԁ���O^��6���O����$�X�7'Q�-��yA�'NR}��')|�O��'�p`CEN�)�X�!�Y]��q��
�24-�l��Oj�cVmW��?��A;���<���Qr�4�B��G!7PT�`�	�<�?����?Y���?�'��DئU�Vl^쟠
C���<�$a`�M�X▍Z�Tp�4��'"���?����?y����DT�kg���w*]�cM�3n�^���4�y��'a��p��I�?1��O��)��\(Q5]�y依C�9zF�>O��$�O����Ox���O��?�@�W�3��$#��6ӌ ˑZ�����H��4txE�O�F7m*���u��d�UH�a��0Xd��o�O�$�O���(�b7M�l�I=j����&�5OϔebT�F�}���:ǥќLhRLf�I\y�O*��'J"l��g4�� *N�<��ib�j���'����M���3�?����?	)��DqAŎv� ��/D>@�"������O��$�O��%��'Wr���ݭp{��r�L�y7�he!�
�U��Ǚ}~�O2��2{��'B6|��7!�y:��׊r��Y�7�'�r�'�����O��ɜ�M�cƉ�+��IP�_�K�$�ɉ�%ܠ��?���i��OD,�'���[ѾXY7�Xj9N�Ũ�c)�k��8ˡ�h���ޟh�b`ݕcX�tH6?y�j��
�.���BH�8�V��gF�<�(O��D�O|���O��D�O��'` E��ʜ#i�fLKB��D�����i܅z�'�"�'��O��+w��6��a��Ώy��	�%�X�p�d�O��$��S�h��� ��<m��<�#c�W�f"2$��b:� ��B�<i�n�!)AH������4���D�*f~���˅�,����D?TV���O~���Oʓ+ƛ6+��aL��'�R-K��E��L�dhB8�+�%l��O��'f��'`FOv�"ҋ��9��T��Q
'�V��b?O��M%�BDY��-����?ݘ��'^x��	�dE�W��.S,���I�lʀ�b�'���'�B�'��>)�	9p͂��A��V�ɛU`�v��I#�M��n��?���iכ��4��]C�v�d�H$'òad�`+��Ol6M�ϦuI�4p.��۴�y"�'�M"cF�?5v%4P8A��7e<5P�́#V�'c�i>5�	՟�����(�I��� �$�2Ӹ jV	����'�(6#It���OT�$9�S�i�x�Cq���NV�Ud��(�ry#�Ot��O��O��O��d[�K�ؕ2&N& �8$�B�	P�"׏J)f��	8|���'�P�$��'ܴ��ҿ5o6��* c���W�'rB�'������U���40����iB�yu�
�I�D�d 9WwV�ϓI�V���Iyr�'v��am�6$��Ɲ ��\k"jV�ѱ��1@H6�2?)D������ ���u�C9��"��ƶ�-���w�����������	�(�JR$��X5���مX/ZX�P�T��?����?Q��i�L�ÝO�B�w� �Ofr�(1$mA��@P0m��iq2�`� �MC������ۯ9i�&����ϑ�.�qr�^"�R��m|����'9�!'���'��O4�S�!�"��ǚ,i
����ɘ�M�,=�?����?�*���#SN qU��	.z\�͕�����d}��'Y�|ʟD���^�\��r��J��s ��
��d�`ԗ��T��P?�M>Y��A�z�B=b���!� ����>�?����?9���?�|:+O�=o�E����J�0 �H��F�����Gj������,�M+H>ͧM7���D�&�}��<�&�V6"��	I!Wܟ@�!zpl�i~Zw�� �Пʓl栳bJ��
�<l��JN��<�*O��d�O���OJ���O��'p��x��N�VB0R�@_�ŉ&�ipР��'�r�'��O��cv����R�d���Z�`(,���G�hI|�D�O��O�	�O��D�+d07m`��"�G�/��=j2��"" �i��?o�
1��'!�'��	ȟt���o��Ls��")f���c�7`]��������ȟ��'Ƽ6-@fN���O|�d��K��pړ�Z/s8:1�pMB-x㟔��O0���O<�O����c�V�|�� 8
��Di0������O(0�pQoZ���'Tab�	џ|�Vm� /)6$�稛�'�$�hV��۟�I��xD���'���إ�J,p�������
���Z��'��6�J�*�\���OJ�o�r�Ӽ�U�+1~�uJd�L�k>�����<��?)��v0ű�4�y��'�|�����?yc� f��Ҥ۰S�g*F�{�@��D&���<ͧ�?y��?����?)���3��|� )Y�`5b�P֏Q�����2ǅ����۟|$?��	s��ЩA��.8D����C�kH���OV���O��O��O�����ap(2���@j������7�xuj��s���'̾�Q��K?yN>�-O=Hr	պ2߰�1GIϬ_z~e1��O:���O��d�O�	�<�2�i����B�'�,UsRϋC$� ��Á%;����'��6�%��?����O�����r�ͻM�b�y�ʞ~���1Ó7K�l�^~"��O`����rܧ����-����c��yٷ$��<����?Q��?��?���9A���X�G���[�R�k���'r�"l����d�<aR�i$�'���FI�}Ebה�A�\��5)�|�֟�������1d���9ϓ�������`��;���$�B+yL!Ґ�O��O��?���?I�5�����3��q���������?�*OnDnZ�jO���I՟�I@��o�	�nEJ�eI�xd�h�'�=��_}��'}2�|�O��E�U�|��Ѫ͛Klh�#X�P�[����-��m�<��'=���@�I3c��� `�Rw���V�Ao7.��	ԟ���ϟ��)��Fy�b�ViZM��(0�� ,$,_��y��&d���D�O@�d/�4��˓��V��O�.1�!�>[`x�%�G�,�7-��A���ݦ�ϓ�?�f�����:�'����=Į�)fo(j�T�X��V�'f��<Y���?Q��?����?9/�Hl�[
 鮽�rË+t���V��ڦa�&
}�p��ӟ�$?�	�M�;��P d�'$8.�8@[qdڙ���?J>�|�0A���Mc�'l�����I�	��m��mB�~?|��'j�L�pO_G?�I>�/O�I�O<�����kW�������Q����v��O ���OP���<�E�i�%��R�����l�`x�	$>IV���$�Ҹ%��������ۦ��۴S��'G��r��pm)�D5zD�Or�T(�v�L��!����?9���O�`ci�(.!�X����p���¡�O����O��D�O�}��
h,,#d�ۦA��0�r��YK����^��6�[�&W�'#�6�6�i�9�ФRv|b��#�괛��x�t�	Ο�(ڴ/��Jܴ�y�'�l��/
�?!�t��i���PE�\�?"%����'&�i>���ğ�I֟��I#2�D������P9Q%B�Z]�u�'�6��	��d�OL�d4�9Oza�feU.5F��aƀ-<�yN�[}Rm�L<lZ'���|��'��#��c}����l�2F��EGTGM~��45~�):p2Lb��On�O.˓t��邌O�S@ 鲅��3�f�h��?����?���|�+O��m8yPp��I�x���)}ѶiȂ ���@���M3��b�>ц�i�\6����J�I	�f�2���/N;n��d*4l �H2�xo��<9��B�"��?ݕ'����w<�pR'	G�^)��+�a�
XL��'���'	��'+b�'>�4M�A�2z@�q�Q�0頒��O��$�Or�m7�i�'�7�7�dDq��a�hñP>��駀­{�@�$��mZ��M+�'`���B�4�yB�'&Z�h��\�0Q��S�T��N�G]zh���䓬��O����O��$CMLJ�(ѾV�tS�/�5��$�O6�X����N�&��'�"X>u�j�D��b�	�5"Sq��o8?	�_�������qI>�O��@�v�
Bf������m��Y����0k��b��i[���|��H���$��8��Q�[�$p`	�9�51RŒß���ϟ���֟b>�'.7��$<� ����=��3`�:y��M�P��Oj�$K���?q�_�d��4We� ` �4U2E��N\�gGns@�i� 6�6YB7m;?Q@̴T:��ay�� -|c��:p�ږ}�P��挲�yrV�H��ӟ$��П���͟ �O?,a�N�e�0��WR��p��f����!�<���䧪?�#��y��S2O~�mDrEi���k*87�ϦaI<�| ��.�M�'�Vm	p%�.f���	ޱ;��C�'R��a&��n?�L>�,O.���O�Z�nо?pɈsH>�8ÓJ�ON���O���<���iF��V����.z)��"��E�@����C.I^�&���I���$�ɦAKܴ[��'w% �f�Q�d�㕘d����ON�'�T�^�r �G�'�i�)�?�G��O4k�OV<a��<б��f��1)���O&���Oh���OD�}λ;۶r��5?&L]au��l��a��<'�f�R<+�"�'_�7.�4��7Px�㕅Û
MҔ:�H�h������s۴5��v��\b�����!��C���J*4�D��o��lrp�+'a�,Z��'���'���'s��'o��'ຩ��+�mc1SY��Rd��g�剔�M�ɈP~r�'`�D���������C%Rt�1��f���?�����|:��?�5���&F��&`ݶ{���8����4B��ݴ���T�uB� 8�'��'J�	4�� �Ū��hX(�R�	;r�����O���O��4��ʓ:�v퓩Y�""]����>6)�fg�)M��O�)_s}��'6�'3,�Ӵ���I�*�+���cT����g�����\����K��i<�i�F�p K"��O��:�ζ|�� ���*�B�Q��ˡu刼kFφ� ����S��L�˼h�DH`A����`a��T0e��p'��+��|�&D
GdU�&f�4I��M�zjꈩ0&ҽ�����O��c�L6Q��� J4+�G@�A�"���BjX  `��xI|����D<yvD`rd�kWEE�UޒtR�)� �Y�#��a�ֱ���؊J��ؒ �4&8X����oo�}�iW�3=��� ��}ΦQX6�݀^�^�� zF���԰-����Q��<���i7��'�2��-�����D�O����K2�E�t$H8����6rb��(�oM�	��	ܟ��#L���?3�@�;"��M��?�D��QV�t�'�r�|Zcq�I@2Ѻ&�((��dYk��ᩨOFY��b�O���?����?�+OT���-�!d �ؔ�ؔ�+Sbߘ:��'��ޟ�&���ޟ���3p�Eb��ی��� '��$'���	���	dy¯� Zh��S�oZ<l J *���j�"�,$m�WyB�'��'�R�'c�]��O��ʡ�8��x� Z?`��T� ���t��Py��g�'�?����]�x��ԋ�/���nܺқ��'��'0��'�A������O0���1>�5�տw����'
2V����J�����O@���~��9��@��ąF84�hP�~�Iɟl�I�����?Y�Oj�x
��H B���w�K�%��)ߴ��dG%W_�֊��?���?��H�i�u�pL�@��k�-V;�Feӌ�$�O�:�,'��o�'m`��e	�{���K�<�Tm.!.��۴�?����?�'s�ITy(��r��=���ߊ!��q`�bH
s�z6-�⟬�R��y��8���9��b���"X�q��i2��'B�oF�5��듌��OJ�	1V8�}�ʽ>:� `���&�b�\bGJH���Iğ�Ȇ�t;���5��Vy��Ϫ�M+��c�4���P���'Fr�|Zc�&�@'�լzR���2)%����OJ�z���O(��?���?�(O<���(J"fLpBf�3�e�ŇT�˾��'��Iɟ�'� �	ɟ����
)�$�z�AA����%�!v��&�p�I����oyBmC=Lo��S�t$�BG�%k8[F�O,q��7��<Q�����?Y�Jc�ի�'&��BD�/��qY��Ьk".%y�O��d�OZ��<	��1Z�O��`@3jG |VD�B�]|�2#��f����*�ĭ<�@ҙ�?!L?Ykhʱs4�Ж�L3� �bӔ�D�O0�Q#x�I��t�'"�\cV=���D�`����4�ñ,+Ƶp�4����O���I'����;���k���J��ч-C~8r�.k��fQ�IrF 8�M�GY?��	�?!8�O�I��/f�� �f�|V�z׸i��	7
��X����ħ��禹��͉+
(.H¦�F�^Q�hۑ�m�6�!V!Ŧ��	ԟ����?ŹH<�'mN`A��]S���K ��8Hf$�1��i3�Ȑ�'$�'g��O��Sd��)�d�4��@�(^�$	�Bg]��7��O$���O�49�K�<�O%�|���H���TU$9�P���?��9����z8&>A�I⟸�I "�W�>bH��3$��@�4�?�3O��r�����')�\�����C��2�L�*!����,A�M+�J�������4�P��<������Bč+����#�$?#,����֛��D�O��d"��ڟH���o��3�I����M�0P���O��,_d��?���?�)O�p���|�H��9|�!�%C/��$ ���i}��'Y��'��	��`��>g
���#�h@H�|�*�AL0o��|��O���O�˓�?ip�����O&�',�4T��	H��h-v �W��¦��?����?QQ��%�^H'�8�'�i][R�@�~()3����O�ʓx�H�SE����'q�\c��X��E�;���x���.g�9ߴ��d�OB���2�<�D!���kl�9," :��^��@��"Ζ|̛6W����"���M��\?�	�?Ia�O��y#�&�V�ˁ��#p�-��in��'��M��'�b�v�)�|nZ�}VD�E��aK|�:� ��qXx6�R%h��pnß,��֟\������|��/Gp�2�+
�Fؘ�0�M::ɺ�l�Ο�������	WyU>���1�ǂ.q��2��y<���i�2�'S2��pH0O�I�O��X$�}Ȁ%�PD��ȟ�yL�oZ� �Iʟ�V!������������� (T�hqF��'�K�1��0
d����M���P�p	�x�O�2�'��	�hn`Ej��>M�����8���4�?ք�?)O>����?!/O��r��Mڬ�䝎$�qi��VB�P�&�p�������uy��'�⦘�s��M{tk�`F�*֩J����+W�'��矘�I�t�'\�\@0�j>�H� S檳� �U1�)��I����D�O���O�ʓ�?��!o�����lh�MI=�TY�k�$4;�ЇU����ş�'RF*J���x�V��.0���.�"Tl4uƪ
=�M;�R�'���]!t�L*K<�AN
*����^�D�ݚR�Ҧ9�IȟЗ'���ʠI%�i�O���Ʀ��`��A��ٗ��/������x�_��;���̟`$?M�'�
�À��W��y�b9J��'�Bb��2�'��'4�TZ��]#&���e�mz�0ᘔk��6M�O��$�t���h���)���� ���K*A���t8�6-�u:Nw���O��d�:y$�������Ø�N�<ݪCi&d+
A��4|_2p#���?�,Of�'��D�OJtZ��A;��P˂)�#n�
���u�Iҟ���1spR!�O���?��'���p&�
�s��q��7W`Ց�4�?����?Y���<�O���''�Ù<��Ԣ��P�N����R��r��6��O�$2�)u}Z����Zy��5� �ɹ#ԳT��ЋǁgQ���iu����yr�'��'@��'���	jP��aB=I�z��U��,^��$���ļ<Q������O�d�O����L�l
4D .1U��u����z���O��d�O��d�O2ʓ4�|��p;��HA��S�p2�5���Q�i������'�R�'�b�B��y�Q\v�)��6\2$s��N|�7��O���O����<y #IZ�Sݟ֘�e<����M����2����e]�\������p�	�����d���hm���1��D�ٺ ��n������Cy"�\n\0�'�?a��"��[	~�6,ćY��sD��/��I��x���@z�@*�(O���t��+�lJ��y�� �6͹<��.W�J7�&�'���'&�Ԇ�>��f|�
��ܒf�H�ҏ�bH�xl�⟘�ɤn���ן$�''q�R� ���(��)3��R��i�� HsӚ�$�O��$��d�'R�	� y7Nk� b�h���ߴD{�XΓ�?�+O��?�Ɂwe�=��%
+mݼ�e� S�P��޴�?!��?��J_�l��	ky2�'��$"Μ����T�(�P�m	 ����'��ɲ]v�)Z���?i��δ�Ȧ��9��i���Pu:�i����--���$�O|ʓ�?��B; �i�	�$s�hh��	O��=�'j��Z�O��$�O~�$�O��he6M�#L	scR�G Ї(2
�󌗔E���zy�'�����@�I��  �M��{l@E:�o�<H��fY:ZT�	�T�������ğT�'0 Q`d>҆D_(��ǉ'�,8���Ӡ˓�?�.O����O��$I)���n��ܸ##��k�L��cە�o�ݟ �	ɟD�Icy��5����?�s�>#s|=��O��ZG @2�"��v�'��ɟ��ɟ�bSn����Mc��UlQ�i�	^z`��u������Işė'�^�gD�~���?��'_!@ͨ񯈍x}x���G����[�[���I�x�	e���|�	r�%�E��$�M0Q�����m�a�'���|�L��O��$�R�קu��ƯQ�X}���K��LóAU��M���?!c��<K>Y��T�B�gn�	�$/�xjㅎ��MC�������'���'x�t�O���'���Y�Kn��q�,F4+�� �&��L��6���)���d�O��ĈZ������',ޙ��'x���&ŕ;�H�'k�:���O��$U�:Bi�''�	�\��?�Z�b!�J)�L�����>4mʟT�'.t| ���	�O�D�OX����ͦA	�c�H̓c��H9T�J˦��I�D�Ib�O���?	,O�����d���]�";���c�$�R�0��Gy����,�Iɟ,��py"B4���+ǁ��i��"
*V��ǃ�>�-O���<����?Q��?�~�F� [�|���" ���b!��<�-Or���O�������V�|RC�kf0�SA ��8�����i�'H�V�l�IƟ$�I�}B�	":�$��/Mǒ���O*2↸��4�?1��?������M%pH&��OgZcE&}1��a��iDn[�1�Āb�4�?9(O��$�O~�d�8e���OF�d�t��Q�¾t@d,��L	oZ�����By�ٳu��꧁?���:G�%]޾��',ݡ%��%��q�����(�	��WH|���'%ޟ��aBZ�rq>+�?/����i��ɢ_.rcٴ�?)��?��'/�i�UBD�FMrH�Y�$ՒF�����Mx�j�d�O��j?O�	��y��i�<�:؋�i�;etn�pQ�O��AҦ�ޢ�M���?����Y���'A���"�@���G�I�7#Pjw�b�Kŗ�d�'1�>�DL�)#f̲'ְ��!D�}��en�����I��Ђ"����<���~�쁏q��㮛.H4<ܙU�7�M�����a�?��퟼�ɏqg���':�Q g��1 ��}�4�?�RU"v���uy��'����֘�0,�%�3���p�_�:/��i�̓�?i���?���?�)O�]X���X�T���������VH|��'x�	ǟ��'yR�'/�7�,��+[: ��5duv��'���'���'��[�@/Y'��eۏ;w�����/r �!��ɛ�M�)O���<����?���@�wЍ@pfΘl@Dd�ǫ}ގ�+&�i	b�'�2�'��ɋ1 ������������ӽ(��!*��[�+ޜh	�i�"T�X�	����ɑM8�IU��482���AN�BE*�N�F,��lZ۟ �	hyҋǕ�p�'�?������#�E�8
w���L~�@bb� I�i6�O�����3?�O��d9�\<R����s�G�.���4��DYx�1n�؟@�	����S�����n1�P�u����[5��p�h�D�D�O<8B?O��Od�>MB7k!N�v�w�͋?h����d�٘�� Φ��Iڟ|���?�ۉ}rkԔuC���ܰK�xȥگ_�j6�Q?1+�D9�D(������M$@}&�c���U��̠eؒ�M����?���1!����D�OD�I/Ejn�p&m+/�X$2fk@�
6�-�Dۂ)}��d�<A���?A���Ì�1q�X-�!�	%��HD����!�	?O66d)I<i���?AJ>�1sZf�b5.�n�����矺%cr��'�
%���'��ퟔ�	���'�h@{�h�
�Ψ�G�P��9��!gpO��D�OO��d�O�؛��e�v)�P�A�6庀�ÕH�H�O<�d�O�D�<Y�HzT�I*AV9���B2_3�Q��1D�	��|��v�I��x��5Ĳe����� $hJUmoM�4�(��.�5��Y�`�	ןl�	oybhAf��PUp�C5��8�'���3��FB�����\��ԟ���9C+���~�dU�YIn$�4�<��I�'�Y2XΛ��'�S��C���ħ�?���QI��;��C$\�L�#�:Ѱ���x�'/R��y�|"ݟڅ�3�-�޴ vjO�)��P��iw剦p?���4%���ן��ӆ��������b��[�y�
��FE�d��f�'-����y�|"���l5���:N�r��&c��fh�,T2D7��O^���O|�IYh�o5�u -@���cJ�6qR5a`�i�@IH�'��'���݁�t%3�Dе.̾��֮�06�x�mZ������)����'R�O�5 �m�3R�1�3\5*VH���i�'c��Q�5��O���O
`k`FG�J$�u	aɜ�b�BU{������	'.y(�}��'ɧ5�jАCf(URf%����Va���$��et�<!���?�����d%ep���	!`*�k�Ҩ]7T�1� L�	�,�It�I�(��q	�����Z�u��a@߀L�ZH��gk���'��'��R�lSԌ������`C�CeK�\�������?1H>����?9�%ק�?�֣��3Y�5ɕ�CN��@C&]�W.�������˟��'�H���)��LxeBL���,8�-qs��:�x�mX�'arMM�>���'=�$;5��A� /W8�@��V|t�6�'d�Z��������'�?q��sT�J����,�wǬIK�c�\��?�!oU�?����T?��%@�0gq� ;wm,Xb�I����>��i��*��?I���?��������cT�"����F>NM��йi�"�':!5F�/����O���cF��[��hir�ɣ$��j�4�%m��M+��?	��zw�xB�'�؀���!qۚ��P�H�F��+eӠ�I��IR���?a���g6�7P�37�e�$\&k"���'�2�'�l���"$���OD����`J�@�[n�ԁg`�-�:�
>�	�CX�b�<��쟼�	q�\���+IZ� "ݿ)A����O�J�G�<�)OJ�D0���7s��(�G�!��5�p��6r���'��A�'A9����O����O*�y�RC��7�xcv��ڶ�"�!Q������	ɟ��[�d �P�'ԾG�T��N\h��xze����?����?q��?�B,ǧ�����`�LUA�,рh#Ĩ�%풲�M����?����?+Oj�"��ix�F�9���PGȗ�V�ဩO���O��$�<�1�Pj��S̟���O��&P�q�Ɔj�0i8��_�M�����d�O��D�On���6O&�D�O�5	 �D&h�: :��*Z(-�Rf�æ��֟��'��$�L�~j���?��'�������i\�
�έ���"f_�L�	������:��It��'��ɂ�m\����C`r��f�Rꛦ]����G6�M��?	���
�V���9eV�h�!O��@ �	�8!�
7��OZ��Ʒf�6�6�S�P1`�/�$�$��j�p��6Mũ-f�mZ֟��	�h�Ӳ��ĵ<هjƇs�%��ǵHZ���f Q�[��&ק�yR�|B�	�O�m���X�rt��E�a�$�c�Ȕ���̟���w�y��Otʓ�?i�'�zŚ��O ���Ab�)h����ܴ��f|��)Z��?�X�U�D$ѡ2��8s��Xw��!�i�Ri]�g������O�˓�?��L�DC���qR���B�p��'�蜳�'�Iҟ���j�(o1�Ġ�-� >��&�!���b�O���$�<I����O:��O�iZ��V�8�HP ,G�t�r���d(�İ<����?9���?	���l`�O
����!�w�,-��耸A�
�"�4��D�O�O
�d�O
Yb�ˮz��6��.�H���쎨;�c�@���$�O>���O��q���QBW?���.aFlʆ�gKQ�Y&l�T%O�m�I۟��?A�	��':%���PI(䊱[=[�^ɘ�4�?!��?���Y��pZ���?����?���,5L,5\�P��8�B��o���xb�'����K^�}��y��"���ˍ+��(b�Q�H��e�w�i�剩Z��8��4�?���?��'[��iݹhtM�+8��9@��3Diy �fӬ���OV�K�1O4���O8�D2�ӕ�d@�c�ƅ3}v-�@�M�"�ǽ8�n6M�O8�$�O��M}BQ������WNlQp�MUˠ��`��M����<�����d1�Sٟ�z�+ڸh�R��!�\`"ي�kX�M���?��>>	+�Q���'gb�Ox�ԁ��F4|y.G�0*dX��i��X��P�Aa��'�?	���?�����5�:�#�nK�&D�V�D����'T�1�স>	,Oj���<��# ��0-���A@�mH䬘w}2$Z��yb�'���'{��'��	E6�z�.�{z8(#bP�X#�E�����<����O��$�O:��m[�XL	��x��pU]�2��D%?�3MФi��Z�eX����	��4�t56�[.F*�Ć�Jn9�ЃU-��@jD".$��x�NC�)
$��Ƃ�uڔl8q�1�ɢmH0�����1s�� ��x��?P�1M:���*քc�^D{��1A,��(̫hQ@��kG��6�qPC��:LkU�
Wܮ��R�)���1.��bB�Xp�:9J)U�~�n5�V�� vj�s�E�$n�č�d�دP!�di�	 /"޵[Ǐ�9{`���L��bC�A����[�)��ٲ��?I�L#q�Q0���)-(\3�A �&�SJ�� �(�� D��8 s�L;}�v��$�>��`A�`QfK[�u��8��P�1rph�~���ίd6�2TC� d��Ub�DF)`�'��>Y��)F�����]>��(a�Y�>m�B䉾[�,��Sᑠzz��'��)"�'�#=��iϦL�t,��+\�c�v�ʔ��}������I�iY�@8`hS�t��韤�i޽h����t٨Q���#��9��O�U�F�[�\�ê �Y^\b>�O�l0�`�&Ϝ�҉	�r�x|�u�@CC��a�O�):U������vє��043���;�O\�<�����Ą:��Oў��C��?�ƅ;0��y�tq)s�$D��"���� ƴ ��
F5�~���=?�c�)"+O�R�O[,풽j7�Ӥa������C�r q�.�Ol���O��$[�C��?�O:�٫w�ǟ���"0d��GLbm*G��NȠ|1�Iݺ0"����'�~��e��;hV��j�O���0��h�<��f��.䋷�'�<�waӴU�KD`��8#(�g�<t�I�`E{��ǩa�ԐW��6cYd���X5K�!�Św�j� �f�kP
��'@��J�1O�\�'5�I�w�����4�?��Xǚ�y��[�59,ٰ"�!�ؐ����?�ˍ�?������$�֛��|"�/3�V �P���ݐ��ߏ�p<AC����'J�u����-O�-�PgG�Hd��Ǔ3�h�Iן��'TX�#$���3̜�j�$҆4��C�'$��'_�O>Y����^3��siC���Y��:��X۴F�:�PDI�'2Pze�E*C:�r�����<�L�'��W>Qr�lX�D�@ݸP�x$���bc�@�bY���I�o=�\P� �?}���fP;�?�O��S����mA�s �W�ĝwU�']8�+�h����E�8i�>e��	�(gZ�I�aO��H�.� ''%}£�*�?a���h���䒨Vؾ؃s�0/��L�p�Ѩ&$!���3� �������8ax�"ғb�~5�c�8!�R���b�|?\ƶisb�'�2��-�!i"�'P��'�w�zl��M]^ ����пC�`�$/�W�С�c\��AZW���|�1��'1�Y�&Bʂ,rH	���B�kl�P;Ӭ[Gr��q��*ߠڅ ˮ����d"������Hiя${�� �y�$�?�}&�������ZL�`�f9C�	 Q��蓐�NZ�٨p�Ӣ��SK��"|��^�b�X1B�"хpC�1Zb�۝?v�\Yaf��?1���?y��au�N�OX�do>� �C�k+��@�b��k�8`1�+Au�@��&�4]L�µ&#LO.a20�]�O�nL���ٺ2b�Ez4b��.����EI���tI*3��}Zax���/b���A�W Z 68�R���%����?��*Y1Q����׃�X��3��N�<��!�:t��邅�4iRd8G�_c̓K��O\�0&�Ŧ��I��|"�ĝ19*	��ĥu�h}��F��H���`+Ll�����ΧX�!#�4��O�䛆+@ y��l8�G$S�( ���:0� ��>����+��Hjp@O;%�e1���U8���#��O���O���
�/V�·�UF�`kP,ZC���?����K&<	wkي�Fa�ak�	)@!�d���P5#E�P�������
�.a[1�`���'��S�Lu�p���O�ʧ8h��J��U�	�3K`���

v<,I����?���K��?i�y*��I.�v��!΄a�dxk��C�F4V�'�yэ���C�-��4R�L�$:���
o��Hd�Ic�S�'KК���� � y�1����M@����za��lK(��=��F_�<�����	+�HOb!�����}�ȩ���Z;!���c��V¦9�	ퟘ���k@�d�DN�ß����H�i�!3E���u�\�*� y#�Xd�Fr̓ZL�p��I�H��E�Wm��z*r��`A3�Z�xIG&5<On�s��0�8M���tT�E{�2�IvT����|��HDI�톕
��t�O�6�y�*Y�3PP@ ��^���8@"�Z����^B�����|��$�xě+Ĭe�X �A+�8z�����b�'��'�z���0�	�|�e�#'�B��a��5�"m�J�a���sB�4��>I���$(�&��3Ԅl���J�B�ĀJ��%s�*Z*�N�ayℎ9<CB4p�EA'0$|8�f�,�������?È�0�:%�0�
�G0�5��x��&��0��YR��Y��>p%��d9�I��M�I>�`Ή���S؟��C�ֱ�8��� �\��H���\�]�By�	͟�'+��u��)%|FpA5����M�E��=w��4�n=
�K��p��xB�ݒ{6��p.�:qK$9�6�� ��EM�dFd�R��2BZ�(�'@����?)+O!����=6@��G#Y��Cv�d�O����Uz�:�9�| A�A�,�(G{�O�x7�V,�M0�8*��QzяY6��<)��G2eś��'�RR>QҳI���hp5��G��ae�Z~�!��N�şh�	�00��IB�S��O��FJU�]R�ԺA�K3L�e('�>�g�N���Od�%��gS:+%L��-C�(�6,�I����e�O����O���%���� �BB�LڼR�$�9�&c����Ix���bֹ)^�!(-�����d>O0HGz���ԛ��\-*�l�B�Al}�7��OR���OH�R�m��y*��O���O���W�m��� [KƉz���mهwybm�۴r`�,�2�o�g�&R�`�Z@B�`bZ`@�K5W��V,47Jl�0��i/$ш劕i�g�I8eU�<g)^)�N`�cH�[��<��cH���>�O��v#A�f�T}���)j?�Z$"Oz�xh�:S��H��.G�8Pd�HV��xj���S$`�(��W�J�]|�<0�F)'�r٫�72������������[w'B�'��I�|���k�W�j<��l͓�u)�OEq`�?yI���<�&)� ����)�O��c ���WCV�����r�� Y�B�'��q�����{ZV��� ��а�'q��A'P~aK�F�6HĨd̓90�O2�*D�N�	��ϟD3@�4LA�'�C�|����!��� �	.pe8X��럀ϧ;c�q���O�l)��J"0=(�AP��4L��	�f��H�浩�n8O�me�߁i�Iҕ 
�[ܰs�N���0�3ݾ �
F��p<�� �ٟ�'�p������ bFS���P�;D�8[�d��t[�l�1��<��9�<�Ġ�4z�F5���OXhF��a�J��i�<Q7�U�����']X>s�@����[��[�O�^<Ht��+WuM��T����gؐ,��T�S��OR�� ��oЎQ��@�}�Ƅr�>�bA����ON�԰C���E~���,��K�� a�Ob��?]�a&@4��`s�������H+D��cI(n,���:*X���-O��Dz��X�D����`m�/`J|�Â�>H��6-�O��Ov�c �5Q�����O �d�O�Ⱦ]2Z�yѢ�V���!�8's�b�ܘD�8<O��	�)�-�NP��$�7S�4���$S�~��y�*؁,��(�F��rي�9�%=�1O��9������o�ҝ�Td�)sj��F !�(��{��`� "lV!
��˂o���'�&#=E�Tn_7�x�P��^�Dk��P�0d��j���1e0��'�B�'a�Sȟ��I�X�2Q�ǘqb�}jN�L���PgF���?	���f�D�e�:�T8#�Tc�Lb��-M<D�����\�� 9��%3�|����si ܈�T#Ժ��ڦ�H۴�?i-Oj��%�� >U��e�F��q؜��6��hO�S/d����K<��1�c9���%��Y���M;(O� hQ�Һ���?�O7d;L�H�O�/H2�i E��?���X����?���d����߯��e�d���$e�j�R�c���\�㉾�Z�:���*���@cT�j�J8S����9��Q��"NI���q�'�����?9��i$�"��F(J�o؁^J.���H�#,����h�?E��OȨ�R���X֕�����0?q�wG�vj .���+ �`O����ცOp6m�<郎'���'G^>	ѥ�П��$��$�ڕ�է�i��#Kß�I=z�X��Q�S��O���c�P.��+T@ı.0��$�>�E��Q���OIĔ9�L�\�f�1Ǩ�8��كH�Ȣc��O&�$�O��d=��	 �(b.�#Hh�r�f�Dc���	Lx��
be�O%J�A���*s6.U��K&OȅEz��J�ք��נ��F7"(��.�6��OF�$�O(�(v��3A?��d�O����O���u��S�9L���4	�U�<$�@��O�Hb>�ON�[�
�%,��ᷯ�#����!Yf�ɼ�Vq� ��|���$r)B�:t��|9���D���'v�#�O���,O����3o��B�?tX�]�6h��;�B�I�y܂�B�m���ă�e�c���+����'��dہ$�li�1+�3>qⳅf�z���k� a���$�OP���Ofm���?���?��g��w��_�����E%o����&^O�l�X6NF�k���e�7��pa`�[p�FP��Q(�j](PY	F"}y4lP�%k�	��5!������N�'}\�� ��a�IŚ
6�)����2��m�O����ۦu�IGy��'��!�7"�z��'�6��W�3��"��No���'���' �fFp(`��)]5r���j��k���a�g��K}_>M�+Y��M{��?!�Č� 0Y%�?UT�MH����?Y��)0��3��?a�Bִ�Q�i��'�aJӁۚvo��faV	-�MQ�O-Hp&�I_~�٭O��b�O[�Y[�}����2=����'�dm���r˛�buӮ���:3w��r����
���"�hN��?�����'�l1	��ҍ|�n�Ʌ�MV���'I^7퍐Gf*5�+A�L�V�ڷ+�+ �mxyrI�uJ%��'��R>�+��|�w ��N�4 ��ʁ<Ub٣RhC����	��l��P�[$:��0j���^���Q���˧AӨ��\��xQi�'�<(�O�!��ޮK)8u#.�K�҉�e>�@H=���ra\Xje�ZA�F�'���h�����'B��t�'�đ�� ? � *�Ą��\R �'_��'_��'`T�R@O |�)Zq+��0�*��Ó]��ȩ���>]`�t c^��Jd����M����?���Ң�Q���?���?Y�9���3^,�s�� ����"F��x�Rb������Y�?�_;�ѹ!�
�0�Y{wF�<}�c�h���4\�q��'6��qgG��D,���ϸpz�mA��'���'������D�O�]�a)��S�9
,��k�MrH:4�H�$I�5���� ي{�r��5�"?���7[�d�<1�dD�Hw�𸦁�53S:]��-�{d�#�N��?!��?!�Jv��OR�D�Oj��r�A�G:C��,1���9&���oM�>(���d��/.���1�FY7Ҹ*�#��l��P1�`C��P�� �P<����'�}���H�d�&Tj ��CHB5Y��X��?�����f�'��	ϟ �?Q҆Կ#�h@�*M�r�`Ц��<��Qa�Tb�c�i��5�S��>���M>�L����R�4���^��u��'�"!��Zϸ��A!Ao�)qa�O$;n��'�.�4�'��0�aa3k�`@)1��C�`�6�� ����tmp=�h�\�xBo��oԒ����F2%���7�i�%���%^�xp:3!��;��x8�4��K�O��d�O:�dP'd%��˰�
�Ht��$�H˓�?!����\�A�� pJ<~3��r�.p!����m)��SW�Af�*}�� c
~��'�fQ ãlӰ���O�˧7������V�(8��@�uk80�EC�W9����?ч�Θb@$ ^�4���|b�k�*����jMaD�P�E{�D� @*�S茋f���p3�'b5���t	V�X7�y����cBU�Oj��'��'�R�	�I����(s����J�1�1O���+<O��h�&�1H�lM��.�v�R}E�'�p"=qGbϾN��e`�G۳@_�0�eF_o~b�'vZ�)�둾z�c��FR���'<$�b�ȕm�I(�,��T:hܨ�'-f���E�,�lC��ADP���'�����U�"��.�8n@�S�'�[1�Q�aeHh���L�2�V���')��'��N>,�SEZ)!��@��'v�ɇ�:1�����/B��`�y�' B����Ƨ\��ҡ	j��ɉc�<I��]�k%������5>�-(���_�<����7b`�P�H�
hp�t/
[�<Q���-�bX��`�1PF�C���n�<A�~H0�A�V�R��C���q�<yFAX�Zٰa)w��:r��'	o�<�`R�,x��	b�8H�ָy�D�<Iʡ~�B�Zѩ7g�Z�I�.�h�<1刳wA*a�R0x�|1s��c�<Y���a�H���v�ƕ���G�<��J#��P�����y�4�v@�A�<Qb���� `R=J��j�i�<��GQ#-
\���C��m���I��d�<����~�X���+G�%�biI	�h�<��К:�>B��H�)>>]�C�d�<�S�H�Iv�c��
}�Fa� )T��j��&�h]	�]'Đɪ��'D��8向5��	�0b�c�.U���;D�L��y����'�C�r(���0�;D�� N%�1�A�s�K��͋Z���u"OLp��M��`94���x�� ��"O~��0�U�O�@q``��<>r�QA��M�\�'����K�O�Ϙ'dHYP���PF�1�p�\�O�l,���%���(#a^���$ͻh���HEÑ�3��1 ��J�ҽ�
�r�T��#�"�pAY��q���F~���7XA@2�ʢ,��"֟,�E'��YW�H1��ƹi��pr"O��Ƣ��v��=����b�4̣q�O\�� �Y=���i���	E��`����ir�� �:�'���y�B�L����\F�f� ��'�DȂ�`�x��#0g�(r-̰sFB�H��1����*.b�s��=�^����N33�azrƍ��܃����&ODp�
ޜDy��`gC/ˊ���܀d-��K�O�<@�6e��'*',�z�Hy���	�a���2�y��e�дràS"tJr]�#��7{9�\	s���N�t�r�`Ɇ�>+�8X�g��y"�U*$��$[<8nK���(F*li5�C�}ǢāW�F�D���  ʇ���O#��"�w�Z��1+�:#���c��B�S���c�'�
�U�3)� 5�FL�6�az��M���C��ejd�'���լ1-�0c���E[�4�jF��5|��@���'LO`c��<Y{�� T#�?d�z�	���t"΄듌�pj�����P��B#�\�~I(@ד#�"��v/X2֐`%zv�m�<I�%Ô~~�Mx�.C()�$��i�@�"m�cOʦcb"�P�&ǨJ������/�<�F��<�t'_6������΃t��1g	�I�E󱨜�?F�=J�1w��1�p/O[��On�a�w4�z�ԝM%�-�7��(
4���'/@!�P�L�n��IM�6/��Rt
�IM���@_�pXl�&'P���M�j��$�=Q�A�,D~����f�9�`�CRfB������q8�i3��JJd�:��F�%�j��sL��c�� ǅیS�n�[���*{G�y;r�'�85`G͇>@�j�sg?&HmZ�y�g="XM6�Rr\l����g��a��Ć%+8֝�81��3�/�]���s�{�XC�	#1�Ѐg`
'5�TJR'$ABRS�O8��%�C�z10@J����N�x�s���R:�	�$���<08xc��]*�F)R
��{��m�2���O��P�	0~s�h����I
�(��a^a�� ��g��)�|oy?��:��I���ї	��)��iN�)`!��}�� ��MZ��8`��3�	$U��C�M�g
A0r�x(�g���
BYJ7�:/h�T;�.�w�����1���T�����wL+?G��r��:`UQ��lܚ��YY��D���.8�֍����
�$�Ƣ ��m>$c��*��v�y(�쬉	��Tc�K�d���;Tj�p��aR ~U������eu�h��J��V�`D�[[��X[�O��b��ź�d�n8��]C����#M�L��j�A
h��I/e������4G���*����u�<��E�S
��!V�'.֔�k��8aplԧ$�Je��"�+�A��_�f�w�% �O>\�ER;F�$��u>:��5��7�@ec1kU	\�nh�g�U�Er¨�VG��w�J�	��*J=}��P)U
��[�XGy"'���-��db�	f"ǟ2z�x!��вZ�"�� �r�k'/�5V�%��$���OQ ���&ݨ%P��L8.�L���%rϾ`hօJ"�p>YU+I?v�x)G�'9D�q�UkN�5u��!��� 4<Y�ôi3���X��}̚p�Uo�Ok,�'�̂�F�n4�t�U�O� �!�D���)1p�N�}��I�"q�	R�d�"���U8xb�(�yӌ]�WbO�g�R�O� �#����+䠭X��]�Y�^���2�-j��ל7�������T�)���?6�!CX�B���dD�r�aHN9rd��*#~�����&TXQ�H�����j��к4�1O��i��ȊT10�hF��5��Ӂ5��`۴s[��rm6*օ�pE�p;�m�lW�`!�jM���=�瀁ZwT����%�`����®[���sK�_a�	�7��܃w�P��~�N�	X4������ﰴ���[�vj�[�>@�\� �
O��ȡ�C��j)j�i�.gcl����1I�u����v�f�����H�ĥ�Pu���2C��q6�x�O��Ũ���7���"�N1 $�Ó5�<�S c� I�0u�-I>bb��Kb���"��`�� s��П�#rČ<`Ҿ��*p���C�~�?��-n��t���2�ب3@�e~��|�n��Wk�<+┹��O�nZ���O�dY��U;�`����"u0 �1 ^�:;$	R��� �Y*V@�8G����XCR.�=�DU��CI�C�D�YfE�de��qIM�)��I����x�.���U��7O��wÔ*^�\��ޅqM����-��q�ͷM���lֱ>
y�-ڋ!�|]���I==�<xf��_X��X��ƧmQ��d΁c��x�%ʫ����)*^�ڐeө2�JE%	�U�ax�.ͶHS޴
R&
�L���Y��.U�1xg�äz�>ȫ��,�م��3�,m���.��шRN�Yp��ϸ'�69��S�^c<$K� ���L��OFyKB2GѨ����@�>}��c|ݥQ�X&
�&�i3٫@&4��M��yf����J�J³+��%��Q^�T �h��dqT���Aib|�8EP5 IVxJKU� 5� �O�s�U�`��$����d?A��� ��cQ�=J=@e���_5 ���b�OX�`WN,z��,����w1pݫci�`M4��u�Ƃ_܈q�'��������N��X8����f��8�$P�Zl�)��"~"N���+8��O갢A�XKx�;�냞\`d,Xw�@�� ��:*>��f
Ѣr<�����S���!���޺�IP;�(O�`b�E_9 ���� [N�h��W� Rb,�<���q�I�.^���Ҧןd�j6Ȇ�n��[��i�F���a��S����5��U@�`>=�&�5m~8��Z��_#J�B򐨜 �zE�š�5�x4�`'�!O	J���_�~\
�X��o���R°�I���ń
(�:�q���"5�d�X����È�!e�Q��%tbx��Z�!#&�P��[R���N��6jb�P��)<?�b��J]�0�E(^�L��@�^��m2��݌��OxB4��`1��ٱ�����|`\#�,�bW�ha�׽V�X����~�L/=�H���y�-�~�T��"ȇ$�n��6D����I�O�h܃#�i~�������u	�O/�j8#%s�z�j`*	`}�E�F��r�ra3���y�h�iO����"��f<�-���MM>y(OFHy��M�U�4\2��O�=�\w��2'�ʻ<�j@��E���H��Y���S2�BW����-yi �9�C����#p-��ѐ���#�8����Oo�睲E􆵃`ꙫL������cЂ�4��7l3�)§
`�C�L�C��!y ���A$��t�O�#�#� %�w��*d�@y�'8��
P$e�]9+
+<���y#|���%�\;*�}�0��2�\,���ԭl6b�*��[�* +��բJL��
�Ӽ�/��d�D)�+�&<�s�z�O&=�w��?�J��P	"� E���ǾyԱ�R��\hc�X�[XqO�0y ��l��6M�ku,+�����o���#�� 9wV�s�A�b�.Q�RØ"�wo��t��-�y� p^BQW��.B1��тd�!^A  �-p5:� +K=-Ȗ���xhs�
�f�!Zt+�*R��b ���?iR�	�7��&�ɛa�b�ݥj ў�i�$qX�K �"{"�#uOp�2,��{rGP �?!����������ڦ)��)7�W�F���2Z٠lؔj	��hO���ы�l8x�4���'�@$9-zp���U
m7��`�'�e�ע7..^��O�8Ȥ�5��ƒ�<G�ː͛�{ьd�D�/!&��Jɘl�a���H���LY�(��X�d�P�m~r.<~�`�5��g<�Z���D�\���K�Dd��I���aXd��!��]�59O�\cՌ�
AeԀ���_�E���A�m�Mx�PN�J/�tX��K@V�O,}����ߝ`!�4f�䐔D5���Qh}�"��"˜�\�)�
ߓ\QP	��kȟif(Փ��BRe�䋕�b���?Q`�4�
: "��B`�S����8������ЁC�m$V^��u�jO�4��{��Bi�:m\Ȱq"�M��iJ�O���Y��qҨ�'?� b�-�x�����w���Kp-��G�Z	�<It%��.ZJ�*�ʈ{s&��@_���'3��H��4�}i�M�z'��a�O�R:��^��\+E�:���c6k������,@�W�ʌ�5�ԭ 6�ȳ� ��\@�yQ�ܨ�H�����'��Ӿ?���P�e�����䂮?g��O���쒎���G`,%�����$�(hp�0�B�X�I1�Eϧgr�����3�g?���6��]���]�?
�X3�+���>�b��Ʌ�����:�|�bfG�yעG%Ti�d��!B�k1Xrˈ��?A�.[���>A�⇭W�2�¦��2�b����V6��'Tb����FH�~�x�!Ӑh��I�g~��;1�e*�Er��!�b���<)�M:2.� �j�%��q��?v0���1��p
���Xݰ�a�� 3�Xwa�Pn�`��ҟwk�;�p�`c�#@@$� ��*7 �w�.v�n0 �T��EG�_�g̓(fb�Ge�� _�L�� \A{ꑉf.�:����s��%�R�Q�L��}��5�E�D���R��9/�CDI�\EH �k�a���T>)��
�򼳆Ă"v�N�bt,
!�|<"aQ1k�,)`c�FG��F��Rf��g?�~Rt%�m\c��Y�[�HS��U��'c�IQ��E?Yע�ԾvXmiR�&�)U}΄3�g͗Q��!wG����P��\S��}�2�4���|nڪh���d�k��&դY�6�G�6���l_�^1IjVE�(�zUh��'Qj���V�N��������p(Z�?aA�?�"~�R��z�`T"4�7�3�Dh8� �Ձ�^\�L�$� S!����-2B,@ kҦ;4Ō�e�Z��&+�"D26�%eJ�����i�9CK���2i��{dE�Xa��HdƖ<
]��'9ҍ���9��y["*�W�O_�UJ����Z��PYbL�Z�e���D���d���I�dJj諱��eF1O��"���w{��(�A����NR��=s��O"L-N���i_�Q�0!�4@���I]'3��a��	��f4�]��(��t0w��L��kB��<�xR�ͻB*���@
�rh��2f��qC�i *� ��1+C�F�k�F(3,@�F"�Ϙ'.�p�3툐^~���T��J>�pj�>ы{2噲����P��
��qh�'etᩒ��#N�`Zq9<�=XWN�j�><��l�U7`�E�hm��A�ޫ1I���Nɑ'���u��O��Z$*8`�=;v_ ���Ӌq���O~B�ޖ��*��-d��{J[bݮ�>����bn�@J�\��S�? ����
ͺ �L�+%KI�l�*��a	�_*��E�:�Eʂ�R�P��	ݚ`�\�k�KHD�S�X��-�@˜u#�����Z��,�ɂ1���[3Ꟍ\�S�ӷl�yH��iiRHr��̸ql�`���#�n̚�.�7�ʍ�.�+F���:V�֌٘Ϙ'ߢ�aH�C�&0�p#Q�RXr���OLbB�V�r%��%�Z�&5��=��%J�^��X�g�
qhLXy�CĦ����f�U���Δ�G�DmD}"��y7�}zt|�&�G"K���IUb#z��'GƵk�lb��/;_�J`;y)Jma@7����G��l&��cdH[�ɠ��	�^7�ɱ�Ŕ�;q�X����*L�x-ۦ8)y�ݓG�>Y�E(0��M�#��r�qZ��!9	�����5[¸��$M�h>�	(�P�A)���S�O�B�b��G̸]Ђ
F @lP=�'�Xs���e�S�O)2T�d�\\�D F��z���SI�ȋD�
 +u����	�w�	c&��>����b K�-�.�'�d�Ya�'s�}ʀL��Q��8�2A�%$W��y�'Њ��%�j)�PGĒv�����/�t�<IvoM�j\�@9��
t�<��KPk�<��^� ����J�[���P�Vc�<	�b�?p�4#/`�����t�<�G�U$0N���(E�T��]6.@X�<��E�*'m�ThE��_g,�j�˘H�<iD\?g.���`�>+��-�u�[n�<i�J^/ptd�S��h�_�<����<�Ҩ�w�Z;[���dM@�<��ӷh�a��e�e�|��s�FE�<�kA1J\x�ЭǚIHh���Ni�<i��¹Vchh1B�o~	��ECo�<ك��%crZ�Cl
�oծ��ASt�<15"ЧTO�|[��B�4@J�d�l�<��N]&օ҆��t%�D�%ʏg�<��@��r�LA�(�*/Цp���H�<ie��@v�U�q[�D�P�afo�i�<����5�:<�Q�]�-�F���g]i�<��L4"��c`ˁ=�J�#%�Tf�<W1??v�r镹p��`3���Y�<i�k��^<��cƷY�:e����T�<Y a܁���yUOD
C��I�%�R�<�eG5O+\ѡ�#ƈ8��a���U�<�u��/)��!�℆8V�x��HZR�<����Xf|ii�K�DR��K�K�<y�Ǟ'��`���t��1�L�<�����āPb�;_$���Ti�~�<Qp��3��Br��>J�� G�d�<�r���&>%�c��0��s��d�<Ye�Ʌz{~�a�&'��bt��_�<�Poʻc��3TN�B��5Y��Y�<��K��n�$��p	��SD\�˲nLR�<��CI�r��E(8�@����N�<A�.�70�&I����͂8���u�<Q�l��+2:�:c�A,�� �udAq�<� ��:���D̝>v9:�ZՍLm�<��� �B�8qZ�N��{�1���Cr�<��
��4v� s��P�`,���q�<��Aۻ)D,���D�xhP鲶�m�<1,ܛ{�(��F�P���
�G�e�<�J�
� �GQ.t4.�:4hYc�<Qc,��	^D�	��*?�b�1�c�<�E��w�`X�i�#b\T8 $Zd�<���-r� a�f�'6:��e�^�<I� B�#h
�-��I�pp��H]�<��X g��`�P��L%�CbO�@�<�rɁ<8K����Лr֭2���<�䇳b��t���H2c��v�<��F� )�,���]xv�)��v�<�rF��n��tA.xp�4)j�<)�Ҟ9WH]�b��%NR�x�vC�)� T)�R#%z�^DI��Y�m��=
�"Oi2a_H�fX����~H�x�"Ox���"۳L ���çvhtYʢ"O�����!�fI��˶X`�,3"O� ꠺ q*-ЃA�"4M#"Ox]ģI5Z���s��	q.t�Ç"O(���Η�L�Śs!�yê�J�"O�Y�uI��!�\`���Z���Q�'"Ov���
�<M��P�o�7
}zY�G"O,xfH�uv��D�$l4�
$"O�"Ё۴	�� _�X]�!12"O��(0"��Ĝ
 �#`@�P�0"O�7_	9�>)1�`U�{ͦ�Y�"O:��I�DJ ��`��Aa�DP�"O,��f�{V�|j� [z%��"Od���I7
�p�#@%��d��"O8I�N�C���@)S�~r�9�"OV�0t&�%_�f�Z@�Z��D�X�"O$R�� ;x,�:C�J�5D4Җ"OXPI���,c촄k��ߣ:.VI�e"O�h�EM	P
�E�F.E-�"O�)b�%H)Ԉ�r oԯ;����R"O|�a?On֠���)JN�X��"O��pWči�����m[$yN(T)�"O�t� d�+�8���;W@:!�s"O����U�+�t��_(�9��"O����!�&^#�E����s�!"O��Sj�9��� �p d���Oʢ=E�F �lU��^!��p�U��'�ў���ru	ːDN�PS���G)�S�24���"�-4M,� �O��R@�iM&D��(5O��;#�8%!�^�x6�6D���wl%c�vruC\'C�`��� 1D��8�i��y6,��C֙";�S��;D����+S����`IG�� "/D�ؐ`�]!D�1�_`�a�?D��ps�F)���[�˝�ڌ�Hm?D���� X��S�W��d��n;D��ӂ��x1�"R*X�'�����A.D� 2e�J~�Ń�IA��� Ug+D�z %�A�P�IA�F��Ó.'D�Pi��4�����Y�.� �$D�4q���Wq���3�ݮ�2$�J(D��d˔�J
�H�tƛ�k������r��D{��	���|��E(V�Z���֏6�!���yU^̲&-T<�r�P P��!��Cx���J�.�|D�Ců@=[�!�_�n�6%r�"q0�2���0�!����t��h!cT�x������OH���G"v)q���֚�*EO��VU!��\�+lPD�v��2�R(��R!�D����m[sոP��)W�D!�$ܪ'�b1���F!i��F�	0!�d��<0��8���E�E%fUў���	�q�-���F�D�P��Дw,BB�	�Ti�Ⰿ@tq!Wc	9j�T�O��=�}��Ȏ�:̢U�a�,�4I�D��E�<��+xh	� ����fe�~�<A�nJO�`��M96�� pT/�t�<���\�~8؜����	7��)Q�
Lp�<qRA%/&�Yb�Ղ���0�(Dn�Tya�"8��P1M_�^�݋�)BOn\��;�f`aծB�gb�4�g�@�u�n�'_rax�@��4bɧ(�[�uD�+;vQJ�E�4mRLxq"O� ���֮��	�
�K�呋J_�ءU���K���QJ����Q���]2e�PX��%D���'A?�������0v�>�1բ9D��jS��j�P՚��]�qF�xq�%D�x�C�I�@�ֹz��Z�^�윣�#D�q1ӌy�x5A�#q����d�#D�����ʸ2@�I4-�LZ��'"D��p��e�"M�`�J4&	�|#�2D�����1*�y7oI�t���!s-D����'��~��^B,��T��!�d�4`�p({��/y#XU��HE-Oy!��cΤ@g�� @��y��H��+a!� XH�����a�*�1�	��jo!�M��V�oD+XȀux6�$[��d��7�N\�$�9&�DA�0dT��y�m[	=Rt���
��4����.�y�F\�4�@�}�0��nѥ�?9�'�^t�uiSM�LZ��V4�����'H PL�O=`���S#3P*�'V�s�Ԥ�(�1�F� k�Th	�'��萌�% J��r��}����'2���Ì�^��D��Z�uo"e��'(>��FF��"	쀩c?r����'������?�B|��B�o��

�'?���h�}����B	��J֩S�'̸�*׆�|���2ge������'�B��/h;�$�\nx��O��=E��K�(#S.�3:m��k'Ƈ�p?�O$���E�R 6�� s�~D�"O"-+QǙ�htd��ő?|����"O�-��ۀc�E�⤐�e �Q�"Ot�T��)Vp̠�aҹ-c�C�"Oz)��#5ZkABG]D>���'1O�e���$�P���Ʉp.@�3"O��������Q��gL(`2'"O~u�%�P>����R�ؖBjbMA6"O,t���2`�Xt#�ݢ&O(
�>����I�.�B��j�(R���'\�!�K�,�Ul�QO�a�Uׁ�!��U'v�2�@+I;�4�M�#|�!��4P�4 0A�K"4����6�Q��F�i�:Q8f�R
�,���k��y���,�=��LΰzU.�`H��~�)�'qH��3o�+[F�c%��;͇ȓww��#m[1sO��3T�
{N�4���a�K�9���K��El|��'+ў"}�%q:\c%d�5>���oOm�<i�,�rƬ��k�1DU}f��e�<�5cҺ?~�a�珜�*�}����`�<Iң�!:��J2�O/!�ɑtO�D�<� �δI\� ��5&3�@Q��Kk�<i�g�}t8h��z�����Sb�<�g�@�H�tP!b
.,�py�F�]�<iJ��dB얦0�D��0AEU�<!��*L&�`�KA;j+J	�oDR�<�4bS ^�~�ē>A�0Js�FK�<��吔]�ȒU�Ddiv��$Um�<�KB�Zp�Qb����ITPy�b�m�<���e0��HF�Y�.�Q��k�<�5}abQQc��y���d�{�<��+�%��=9r���q��{A��A�<��eY�;j�UFΰ~*�[6��r�<�㚊T�>����)tNؘi&��Y�<�0hƑ0$��C��v'.��`.�X�<� r�d)ͻ�����>\�Q�u"O����^�I����S.�Z�N�r"O*�a�Fp��-�$�R!���#�"O �	�ء@F�,�S�Ҟ����e"ON�9��B2�v�Ʃ�e�i˷��l���	�*Q꼽�GX 	��0	�+�i�!�d�U�>BK��X� h�mV�0�!�X+C̺�K��_?I1k1�!�:X�b	�c`A�\��Y�`�'�!�DE�j
h���%��tb�iL��!�[�f�~�6o	�u�����.��Gg!�dU�B��*:,�^�u�
�%c!�dXx���Z���B���ڒ]!��V�6�ɐ���6'�z���`�I!�d�5:t���):w�!�OȈ0O!�䅉;q�=�d��l���ρ�!��§ ~��BA��k�bb�.A�!�䓓,����t�	UJ
A*A�r!�"O�I�E��B��wJ�5����f"OR�ؔ>@%�!�G0~��s�"OL$@GZ7l�D��BH�	���"O.��B��M|`V�C^��uhp"O��y��Xk���Q�m�1"ORD�C!S�Z�3�M	_l�iE"O�����(#hHXhr�]�(�"O���ϫ �z���;2p���"OJM�d�� @Ԃ؂Gdѽg:��4"O���^8w��#F�=M���1"O�iң���X�(e�u��)�rEc�"Op(2g�/MM����	+����"O��e�[����
�vo�A�"Om��_}�!Ӳ"O����"O��Re�������s�ڰJW"O��
�Iޙ`��L*q
]	#�d�y�"O�͘�)��o�l+ÂN�M�Tb�"O��*W�E�*���{��΂;��\�Q"O(=Тf�N�r9�v��D�4B&"O����X�h��F^�b�� ��"O�%��^	3��IPf�x,��p"O�,��B(b	BeY�g��I�"O q�&��s�Ruf�"O4��"OVE�Ɓ��\y�0�2�/�d!8
�'dJ���ڵ�쀫��HҚj	�' �ha���Y�=�Ռ�>8���@�'�,P2%��<$;�������� ��'z2A�'�H�P�R�ؤ�Y���)�'����D
6\0�;�������-�n�&�%>l�Y�C������eGx��i1xk�-qg.�8.���J�zzf�B��ya�zD�<�ȓV������_�����L�q���ȓ$?������u���i���ꊅ�ȓ\�,�Q Ü�9m*���޽F��y����m3�G��X�*�G�B�L�ȓI�QĨ�#'|��7�êX�:��ȓN��Y�(C-֨ݳ��ݤQ�P�ȓ{7^�I��	�A��۲�O�j&v�ȓ_Oeq@֩WĪL��H� 4x���f||�W�W�Ht�,;��cq�`�ȓD9z�i⁠8��x)��^�/�� �ȓ'�f�{ -�$`dI���#O�<������&؄ar�(Fؿ$c���A����rn�~�����gI�3/�ȓu5���.��n�Ea�G<m�d��S�? p�z"��-�����M�p��\�w"O�a:�%ߙ*�r��ۗ{
��"O@�07�U�HA:���r�#"O���cl�Ei���!��q���"O�˴�uC�t�ئ+ܤ�(�"O0ػvCJ��`�Q�.�a�b�ZR"O�H `��=�޴hĦU�8��i�C"O���σ�\�$,3gNMy �J�"OζU���g�\�
#kڙP`��8�"O�����߹7��Ea�	�KDZd�""O�0�Và	Dr�����@� ��"O���;b�m	W틤���"p"O�!(�eT�hq��B�Pf�$< "O�MZ��O�LݛP�<4�P(��"O�]��F�^�z���� �n�9"O�Xv��5	 �c�!��(�2"O��"�Gҋ���4��d�N�Sp"O2%��i�����[�B��5w!�D9M���X��
(�X	�ơT>]!��
�T���gH���	3�Ѵ�!�d�ϰt���Q=���aB�-v!���=(Y���;�����/�!�C!Of���bcʨe���0䞵Z�!�ă+� �a�	�R�. �P$���!��M�L�Qc��ā%nv(��%�"t!����"i��,�+{ ��#F� �!�D�A��+�+S�vp�1eN�!�D��*����l͗9]2����Ϡ�Pyr��( ���uD-#$M�W���y2�As�~\�%F�����6�:�y`	�zy�E1�,�.���Aw���y����mg�x�.��%����yb���p�D��&�({�",�t� 0�y�+ܴe|k�C�D6,�!�H� �y��;sD��(�1��\3���y�nK'�^��U�l9z2hQ��y�� /�|q��_'ZE2%�L9�yr��
�0���F�#
���
��y���K�L�b L	�s�T[����y���^��q��V)q��a�/�2�y2�F��4�A�:S����N��y��V-^PȀ�o�,R�I "O�y"-I�1~��s�BX|܌{�l��y�c�9t�!�T�&U�������y�k�"p��l�w��Q\����H��yRa;�H����EO5��:`h���yr�P�mN�6&^ά�ZG��y���=*M6A(��:z��"��Q(�y2G�~�4��śd�Y��Nˣ�yr�+;��H?r`��U-�#�y��Np˜�3���:L<0���y�K_;3��8вϋ�0Y�@� ���y2�39�lH���T9T���FF��y����Q~`%"�4c�8��v`��y�H�
d��S�6*�Ud��y�)ڼi���bӯ�� ��	 ���y�̃�C}f��.G!��i�R@T��y�@��ic��j��U��f胳$C��yB��4봡8!l�:�B	��IT��y.ۓBp�iGFKV��ő�y��(K��ŲQ��"���jF(�yr���paJH2'�nَ�SgQ�ybK�?kݨl�Û&_�pՊF)ڛ�y҈S��̹v ۑR#,��e,�y
� �#�c�a��x�j�*��I��"O|͋�`ڈ��H�=C�H�%"O��VE
6:x��$i#5�t"O�I A.] y��y��U))5�qb"O��	�+S�4�ud�0)Vq*�"O��g���<svBH�H
�E��"O�ЁD�d������Vf��pz "Ob|�V!8�k�m�?U4�I@"O"��c�?�D{s�E� ����"O��Cg��o.�]�F�.3)Ht '"O�L"�"�$[v�!c	/
��A"O6�dJ�B�\�Ц�&;��ps"O��DE+��Rq����l�6"O�t��j������ӗhm6��0"O�ՠ�N
��%��K��&��"O�<��C�&`��X@�D
R�`�t"O��bՅR�P�J3i�s�&H�"OV��D2�`��4j�!^�ph�"O0����[���'g%)�ݩE"O���R�T���Ħ�c�^���"O����)x d�5{�튢"O|�c�#4H��D��9%R|�"O���ѫB�!h�0R�]�< ���"OP*7(�	(����M�> ��2"O�1�0I%:��u�U���g���HS"OX���dۊ-���K$@>X��iu"O$�S3o f!�z�3Gm �{A"O��-�T��rOM�_Z����"O]�7bM�Z�Ҽ���){!b�"O�AهӎU,@����I�H*5If"O��jc� �i�p��&H��1��"O��R�f�29 ����'�lq�"O�y	��/[F����
�9T��"O�A�g�O�`�ܳ�H�2u1>E�"O�Y��
����pwN�/���"O��unI�$׎U��цK���c�"O����b�e�Pѕ��j/D�pG"O�EX5C�f�V�Z�Z'}�d��"O<|RU$
��T��t�3	j���矀�Ie�O?2�z���)`��[(u��;,O����O
�D6����Γ(���M� ��-���5:*��ȓh�.�D.D�##v�Id+̱b�x݅ȓ+�h�d[�dOT=� Yν�ȓ)(cUME�#*��+��v���ȓF�z	!�b@f,�a�*�%~��0��[���SG��G~����aI�8EB�)	���fc��j���gmZ�-����<�J>�ϸ'�����3A�х䖨��8��'�A��cC*Jt%����T��'��I����,̶2񥁧Q��A��'Ψ�R���&Z,!���O��h��'�Bm��g"b���{�햠E���`�'���$_�T�6m{g�ӷ=�LY�
�'�����)��F1ꁍ�6rY��!��/LO(X�Wɞ$E��KŪh^�}�s"O�ErGE��O� �[�juF���"O�y�'V+U��T:a�Q�Q � 3R"OV�I�"('�zI��G�1���y"O�BGD�?�Z��v�հVW�	6"OV��$a�dȱ���X8~��"O�r��Kl��%EM&й�G�|�'���� �^T��Q��	8Ҷ���'*r����v�%��E�9$��x��''� #��*/0�,3� eԨ��� �(`Ţ�9u0�bQk%)�r���"O����M�0O�q;��Z��U�"O:�(!+Z��A{T�=���&"O�	q��58x�xU	�;�t�xB"O^9ۦ�"V�٠&�Q~:�Z"O��qT���QZ,��b��?}�9�"O����вi����V͘�hz��q"O�� &��&Y`�J�|,x"OJ��J�RX~�+�K4`wr\�1"O�5�Bc8
6�P�w�Ԃr�)Z�|b�'22�ODjDs`A2A�ܱ����X�S�'D�z�ؓd�x�@��w����'���0�$4�<�U�P3hv�|k�'uX�f.�e��ԣ:M�6 ��'�<�s��{����W
�L7����'�*��F��gz&,�u��6n��4��'J�
�� 6�dѵ(S�t>MC�r�'7a��d�����ЍS�k�ȱ��O���yBF@�K�����2���Z�"���y"O�PK�@��.4���3c&�/�yrI]y|��e�[�lD��)U.�y2FњO���w�*^�0��# ���y�!ŲA�&Q�b�؟]$)r%Զ�y���9�]bdN]��!pNQ����hOq�:���czx�lʏM���&"O��+lΔX�� i�A�Xp��"Ol]Y��Y�]�
8�e��� �4�J�"OjI�@X̚ʂ��.O+f��Q"Opɳ��\�z��}�A��>\vu�p"O4�6��=;{P!�\��Bv"O�p��e��u����g.�i���KdP��F{��)�Cn�ٻ��[� ��):O�F�!�$Ł`��$Y�����Ȉ��Z�`�!��F�E��c��b��
oZ�U�ȓj4��2�5kn4:b��r'�Ԇ�9����j��<�r�m����y���I����ii��U�ui�%�ȓ}5,d�s���R�n�Y�.Ǒ#�$��	`����2q1�Xe��:��Ǔ�����n,D� *%�F@`���3@��f�fl+D�8�0���zhP����Z�3}Z���B<D���4��愁Tj TOz�s��>D�4���O��$k��I�>�P*<D�l�'��=gj�r���*h{(��5.9D���B�p�$̩"JW�*y��SsG7D� �֪H)�E#�5G�L�iGf(D�� v��F຅��L�7&9At�9D��s�F� qi�A���L�$J]���2D��y�$�#�^�xeǵb7Qzbj;D��r��G�9O8��ƋP���d��>D�|B⁉�=5�	9��O2Y�@/D�@������Q�H-����O��=E��&�� Q�U6QĎ����&I�!�d�
�P4IDN]�y��,�ue�z!�Գ<؀�a2!�VU��վp!��NK���qDfQ�u��A�Q��^�!�$�x��E���<ATD���ݩ�!�<C4�Kq��j�vP�@A�P!��4Dx��C�15T���K!�ފg�&	`�L�*.��R"�ֳ!�ă4zm� 4k]�;��Uz���!��?OI������*C��
%���/�!�D=�]H7�ɶ+�|�)pB�:<p!�$O5E�z	R�_6�������ez!�� Xy����h�蟶%j�d�w"O ,JߜG��!�'J�_T�tj��5D�$���[�:�8HQlGsy̼���2D�4��Жzrf�� �V@�EC��1D�X��팑�z�x�gB7�%(u)/D�|�`cBK4|�����S8�8i!�.D�(���S��5�Y�Ȑ"#�,D�kw'\�L���R�WT����׫'D�|"���y2��)��.\B���."D��D�N:ob����L�>'Wv���$T����!̈́Q�b8��
�w��A�"O�uD'^ /�r
��^�|�)"O"�Ƞ.�
w|Z�
f�R�"oT9�1"O �Y�Y�Z�@�Ɉ'Y���A"O��d�	t��B��Q*M^�31"OR�9��J�3>���@م.F����$�OL�$<�%D��᳏@�T��Y�XWc�h��|� Y���) �F���s��#�ɪT#Ҷ^���B� �\��#t���"I�p�ձ'�܃9�tQ������D.[�!�uo>JD^8�ȓWxDсn�X���Ë�����q���?7:��o�V$N�?q(O�#~
r�MZ\��Ѭ�H\��A�<i��$7�x6(�hcޑ�d�|�<I��48V�X�לK-��Gm�<���S�����gYG�Ek���h�<�Wʙ�\k*�j�'Fa-ۡ	�f�<�0؂b�@�{�I��m|�+'�C`�<�4��jn���`�6{�Ěvd�\���?���`}����1��1�LA )�D��"O�A�GE��o_&<���K-So0�q3"O�	�"��*�`@)z�HSs,M�y�͍��F@Y��Q�|K3����y�%G�c4�ab����0�R�]��y�+Š���
"e }�yp�f��y"-��uP"�E�w@���ل�y��.rM�)����mc.�ia�$�y�b��)@JT;��bΌ��pBU��y"��$^Ă���*BUxE8s@��yҥ���:�j�#�C���1 m�'�y"�X�+� ES�/H$l�ɫ�!��y2���v|z�� ��6 ��Ț'c��yR�K�o�M�&�u0Xg!S��yR�Ģw��$`բ�5�B�G����?��76D@�a
�N�\ՉA�A�%���30�j�m�95�j�A3Q��ܜ�ȓ/�
�8W�mw"=��I+ r(��ȓ ��fE��~F☩ �#s$؆ȓ1��(���O�t�J�C�Os$m��w":91e�ߤs!~�7&ϛy)���D!(Xj���/݀�X�	V:�p%�4��I�g��M��H�i�R@���LL	�B�ɚI*��Z�H�c�&����
;|�B䉠3!����@��!N	�0�B�I[����B�Z�t����ܒr�B�	_� ���`�ڱ�\��6B�ɷ9E��O��d�a�@V�C�	�jZd��5`+^^�ȅ<N��B�I(WG
q+c�G��P���	�,5C�I9k��*�
�> ZX)y�M�\E�B䉥eaި(4Ό�"N��� ��x��B�	�k�m�@�\�Ȧ����	�RDJC�	x0&�J� ��)��!�6�ǯ�B�)� ���Rg�nDHZ�
Ϝo�Q��"O\����d���+I̐��"O�]��F\ /4���3	��<��Az6"O$њg�җ+���3��*3�XHC0"O\�4"�W���A�fE������"O���cE:�:İEHMq�I��"O\	�ʜ�u��q��~�x��n�<�`@�'!&q��gj	qף���4��0?���[> ����m]���V�Xf�<���Z� Z��s�^� ��RBD�e�<y�ɷ,<�$���)���g�<��]4<�}�w���Q�~s�́\�<1� �*�����oPK����n�R�<�8J��H����Z���t/N���͓Dn���S���%�T�8�/�?�8��ȓH�y���M5�nM�6)�%0�Ԇ�YT��A�D"���j̒q&��ȓr�Լ��W��� �w��X��Z��%mO0Y傱jR�S��>��ȓ+�J�8��F)�Qz`ĵvB�ȓ#��C���R +�5)UB���HBH;3��9���棝�O��ɄʓtO�$B� �FQ��+���C���!×I��~xr�qqB@"=ҼC��M���`�4*JV)�+
2ʞC䉻ڤ��V-��P�(�B	�=�rC�	�q�%C��"�x�3S��TC�I B�(jă�.�.��b�^]���$"?9�ҿ��)+A��6<�Ț���_�<��$��U)�=7�����KYC�<)�hM������"��]F�E�<!$�m4�PPB����p���R��y�!���Q&b[����[@(B��yR鈈O�TA�'� :��"7�K;�y�F�c�X��P�x]�٢@K���=���?��'��h��#���(�@�X�%!P<��'~l�bO$/�ڼ�rK�2Q�43�'�Z� AGC�F�,��$Aw`^��'1^\�7�
�Q���Hrf�.��
�'.^eR��C� m�Q �B���Xh
�'�*��4�����f�M7C"���'�J�C�㗦&Q@e�V��bm������ğ+S@D��ގa�"%���¤v�!����u�v4A�ǈj�\����e�!�maF�N�<_���g�̑��l�3"O>k��Ma&���7'� ���"O
��&G��7��z3\�}�pW��y���<�j�VM
�&�(�Ҕ&�/�y��M���St�ц��PI�G
�y��e.��w�I.j�t�4�F��y�k�*�j��`OÞl�B���@��y2��;_�𚔢�%Y�����&�y�@��'���)��S�RL����ئ�y"�$hy���mԴFLH�IsK&�y"o�V�J�i�U�7��HY��D �yr��u�!�p@�"X䔁ʴ�I)�yr�Vf,)��k�!G;eO��y�@�'A�X Ae�^�V����*�y����RgtyGO_[hĺ���yb�ʖX�ĸ8-�k���U'͗��)�OB��Ηyw����G� "O�\Y��2i�lU��
�|����"O¨r�AH95ޠ�C ��`�j�"O9i2(6P�c&͗�f\vݹ�X����`�S�π J�C�K>N�jp��8ZJ��b�"O|Pd�_�!��\q1�|֬�5"O�q�a��W��X�L�h��{4"O:I��
��6����M�*�fY�"OF��w)�&i0��x$�K�+jhT"O����\ ��X��î/j��"Ox����c�&����N@H�u��"���D
�*��W�,x+L0qgζ{�!�D�X(���4�(�}�Q�[:�!���S�x] d� �,���"v���'�a~�c�s�6l�"��e? |�@-E��y�cCh�b�l��GFT1!�y�@Ռ>n�:a�yLJ ���y�ȓ��	z%)�)#v4�Ѡ���hO0��鈟]�k���:@İ��aP!�$W�F��U�S��W��Z֥K�R�!��=5(t�$��+�rՂ�I��)�!�Dב0	��w�K�(��� q�J/�!�J�jv��Sԇ�X��(X��/U�!��ǽQz�(I���>@ ���&~!�d3ld�e��e�J��f"G�'�O֢=��`X�SF��o�4І�.1L�"Oz��B	�3	ФB���O��ra"O��ge�6A���!�a�&�b쨥"ON�Ba�K�!]�̓Bᒔ	��k�"O0��#��yZ"��寄�F�8�f"O|A�ǈ�B�B���%?�,}��"Ou`æڒ�Lt*�B)n�|@S�"O���ÏG!,Ԁ���M�HCb�HV"O���\�#4��,�#��j�"O�pXGCO�f��KqE!����"O^�ا�6*V�KB�A��"O�U��/�+(�A�C?h&#�"Oi����8)���wGY���Ё"O���ň:岜*G�,aA(��"O�m�G�0���Zd�	A��v"O��2f�V�{v�������HYs"O�(yd�U*�̚#_��}�"OV@�G	�P4J����eI6��6"O�E[7�־=�rl��ءW�r�"T"O��ǁ@ꄌ�P��{�(Z|�!�$�2=R�[����o�<X"7'��a�!�T�'�8�0`ģʨ��5�!�M�3Ob�`"�u�������j!��مSG���bL�w�T��o��VJ!����Jr^��W��k��x2΀�a�!�ā�r�p	`GV���%�C�I�Z4!�DH�#�J%�1�~�s�ɇq!��ؔ��݂��{�V	cA+�5\!���8h��U�S�6��P�F	ݚEK!��lK���-4��rBʛ:G!�DC�O�:���[�[��H+�.�!�D�O�8�h��/A���/R*)�!��P�m�V��nJ-(xtk���/{�!���,WL@{IK�q�B�k����j!򤔬g8� �S�$L�ҵ��)r�!�j|�%2��A&mIz���c�!��M{QЕڶ,�2���3�Cv�!�W�uL��#v����r$_�a�!�DĎ*0�HY#�֚>��X��*[�!�DJ��#,x Y���_T �e)D�d��eC}�2L�"Nʛ1�İ�7�;D�L��Ht�3�$�1���o:D���uDȇ9D��.�;Zr��a�C9D�� �)pæ�N��İP��}:��b1"O\j�_u�ؔ� �<$�}J0"ObX����q�B|[�kH�z^�z#"O\��e�٫N+����Μh%��"Oz��B�A7,I���D^.+d�I;�"O�8��a���3�[&R.r�R�"O��ujZ�(��uel�h���"O ��'nҖ�v�Ұ�Ω9�l�"O�I���T�f�ųsԬX,�=�"O�5{�攟�TyN�G.��"O\�0P`@1R�"��q�^�V1�B�"OZ1iQhί
�,t�g�.a%Lhzs"O��r!�9\�&�Jum�$l-��"O.���^>*�qC�LSB���%"OR�i6nم%��+��̫9�<I "O>�H�=vdyfk�m���"Olu�g � Ƽ�c���-?�ii�"Oz�2"�;(3��)̝yOd@(�"O�8��/ǢQ��Js(�7B����"O>����b4A��_T�d���"O�qQ3j؏2K�-�!m2i����"O�!P�BE~�4�ۏ0�fR�"O�q�R�L;3ń�kU�M"���"O
�)�	�vvP�1�IOm�l�u"O2��4��r`��I��G��1r"O>�� d�,I��PwH /iR��7"Ot�ZR�Q?�ZI���Ҝe����"O�����А9e��5(��M��"O���[�BV�!%�/z�l��"O@�Rt@�U���8dt
u"O��j�Jߩ39\�s�ɠ+R�t�"Oΐ����x� ���N�� 7���"O�����\0_K�I����C�C"OT��Ey�ܩ���l�H��G"OJ}�4��l6��R�Tp��A�"O4m�ԩٌ_��<�5h�|���"O"I�0f�%^m�٫��Mp��B�"O���a��j�PT��Y�6Ic�"O��K%M��P���)uܸ��@"O��%/��t�Z1�BM�e"Ođ���ظjc0u�T&�#E�d=�"OBx�]�3����V�U@!"O4�;2�^�x�����Bs�xqr"O��ir���:`��o�B0��B"O
< ��Q>��@�a�>�C�"O(�'�
T2N� ���Q�H��"O����Z�>�i��ޛQ%!�d �����Á�@��(��+!�O+G��xÆL ����f&Y!�ˌ+\$!���ٗ>3����D�!�>A������D��t�Y!�đ+H��:P�#��e�� �=e!�d]�d/��W�
v,� �V+k�!��A�t�� �`��
z�r1��T�#�!��X2?p}[n��N�C4`�9�!��H�8��Y�U/]������8�B�|��'�������M1oVpI{�ǝ�C��̆ȓK־I(��H��dsE��4K��8Z�Q�"� '\^t���17��ȓOV���`J�a5%R�AP�[��A��qht]���<��@�  V5��9�ȓfM�`!��y�ƩR�a/=8.�ȓ�T�7��"�L3+�z��mL��ɣ���Y\n�4�F�B��c�<� �̓��/r����Gڿ:��@�B"O�!#��%8��3'H��F�:���"Or�,ƘZ�1�g@~ـ�9'"O:�@�G˦�*t"�H�!�;�"O����+^�ISN�*4����"O:��(E!H�U2�L�<c�8��"Od�q��V�Q�j�����+� x�"O2탖��l�0��a�$!A�"Ojy 0h��Y��L�A`	�.�X�"O���0i*��}���`q`��0"O|� яͫ)���Y��Z5n_�t3�"OPUh�Ɇ;����+�!{[j�"O̥�)�1?��wjs/J�#"O<�q`��)e��J	%@t���!"Oȑ#j� �.UA3��N�J(k�"O���(S�.�<�#,$>Ա�"O*�c��53�6����5���"O�a�̋&r�d��A�19�ɚ"O�ҵK0F��a��*N�9��i�"OH��2A�0T9 ����M
�"O�-�R���C����$�y=����"O������D��E'~�ژ��"O<����-�\����ȒJ����"O4������4h��A�"פ�Q�"O�9��B�C�L,��;Gv�A��"O��rsΔh���j��)Vg�A"�"O.CQ)V�:��h�bW,Im��� "O��D�>#��"�O�\VA�"O(�r�?7Ɖ��/��`h
�	7"O\��4oʭ~���a(KY�����"O�`a�%�gY4ͳ�fX�1뚹��"OB�;�� �$���̏9w��E"O�=/l�$�e�S�
��
�&�*!�� mj��e���H� ����=.�!����K���v��Q�ʍzF!�1-\���VmY�J��L�Qd5jC!�$R g��Ԏ�l� �!iX�(L!�-�4xH� H�1�2�H�(�L!�O�_ �Sԋܲ/]N��tG��u!��*�t�{5L�	T0eC��� '!�$S(:u��*�kT�4�K�dI�t]!��	�~����)#�8a�*�?�!��8\/�tp�Bȯ ,۰LF�D�!�D��-���&͕L�tb���g�!�D�I�ȱ��钡3a�t���>$�!� �.(���2BfL�+�O�5`!�ÿu�� �u�<����N�^[!�$G��(*���,~�jt���rA!�Ę�#��I �G�|� R#LW!��?:�`��S�Erh����+ws!��� ��f	(w� �TKʰy!����,���<&qXX����!�X�"cvh�uf,<���`SgV|�!��:a
���f�]�4!�eO�!���c��x�f�]!0e$QE%!�$��Xi�#%�$$�Щ�!�R�)B��҂�>=���IM�!�$�Kւ��U�,�D���͌4�!�D�?�b�{E(��@�:�@"GJ�|�!��	yc.i@�+N�>� @u&Z�T�!���n����C
e&n!�s@�(P!�$�BTE���5-��d�r��7H!���m�.�� �'�<�dJ̆D!�$�"rV(X�W�B3
�$ �2lDb�!�� �, �E�,:8�֦�I߈$�"O��z���g�B���gɷ%z5Z�"O2 +7Aw|3��{�� F�_�<y�#n�L)J҉n�2E�X�<)�hI�/���@��Kx�Z�s�āk�<yN�,XE6��h�o�:�J�
�L�<�rG��U49�ČZ1$��-XJ�<���ЌD؍p@�ؽN�ڴm	r�<�f�ڈ6�4��ɟ�#��c���e�<)Ц�J���tM�1m��Eg�`�<T�G�:5Kg��� 2���qʘc�<�e�ʐg&��a+�B��!��G�<i��*0tII�� 
s
Aq���w�<Ċt���1]8�0skBp�<)�g�YA�}P'����m0�%�Q�<	�bD�D���5nU)��1m�P�<�#�̓N9.4�)�QX ��D�H�<�KB��lR�
)YJ��T�A�<����4O�P���u*1�' �q�<� b-r��!�A�N�<��h��n�<��H�p�FA�M�o�Ā�h�<�#*U;B����� <L�Xt��d�<)G�P�`���h��7�����	j�<aP��9s\���rM[�G8�)dag�<��n�)��M0%�����A�Ff�<��^��6X�pmA(z��c�LN�<�%%��B�X &*��S�(�a�C�I�<�'�G�m�������;LT��Do�H�<9��NA�q��/�\�b�TD�<I�M�!i�2�ɒ���n�� � ��w�<i4	D�ʁ��M9?|���AΆO�<�4+��b��i;��ȱ~�<`��A�<����K�:����Z�I�'$E�<�֫\^�$U[���� I�<ѰI�
!.���'��T���1���r�<yRK :��q`�̝Wp�TaB�l�<9��L�R���٘��A���<Y��ޔp�T�ޗ*&1Ɇ��D�<���AB������I�	qG)�g�<1Qż���Q-q�J���d�<y��V��f��J��Z㺼 ��_�<��*Zo�r�Iv�zH�yX@A�^�<��T��
[�هG�x90�+^T�<��G�M�x�a �x�6����D�<�H9S����^n���U��H�<1��.[~��Ff��o�@�ڥ�@F�<䎘�ˀ���@�i�ݢ�FS@�<Y`͌�5ي[q�޽	i8ᲁA�	X�\��G41���S3�$x.���0D�\��I?hݠ6-̅$�L�cc�,D��b׊�S-���_�PaLy ��&D�lB�kL�O�6�@&�Ѳy���׬"D�D�c ph���"���Y-?D� x�@�_e
(n�ŮqCDE>D��*�	�&<�t��7CL��;��?�OH���/�lSTO�p��"O|=	���Dy�页��4/t���*OF�HD\^|tDO*i���8	�'�L(�Foe(��	D�4ڠӤ�(D��@b���(T���6ք<�ȓW�6ш3fP�B� }"��\5�XI��V>Nܸ7.ܤR�p ���~\P)�ȓHE���)Z�J�l�⣍k�<��ȓ3��U����W�N�D�Ƽ����S�? �ѻ�aZ<ƴ��L>�D�7"O��t�)z��cɃ4.�h�e"O����'�w ��9m�\��"O��	���s�ԡ�h,\�T�p!"O�Š���3|��H5ȍ*)� �!"O�CCL�����8Kr郳"O�!#��D�]� �Q�)�cN9�"O<պ�,V�^+�Q���_�\'�iI�*Op	"e��y��Y�4ɛ�<<�s�'cN؁0A�3�YJ$��A
�8
�'0���2��=>L\r���{;�	�'!ȱy�eM�p:���<x��2	�'� �j�J	�ȥ"��1$^N�	�'��I�cD=
S�!�����h��'�d���@D�}�h�� F��U�,�q�'�8б׈۶w���Y��>Mn]��'�*���W.(����.��W�92�'JҌ�1g&�@@{���$W*� ߓ�?��O�QP��U>S�6ً��$X�&���"O�4 �m1G�,��֩��o�p\�#"O`h�̍f)��dJ�-v,X�"O��Zb�Ǡ/�|9V,\�dA�"O�4���$"�9�㕇~<�t"OZ����0%��!��mҞC 4�`�"O���� �n��M��p��OB)���.�J��0Y� FdQ��N5D��ՠL�$�P@�Ɗ�0�<ق�A/D����̕�]�����>�
��VD-D�Бd��h>]�҂�-V�9{�+D�P`#-�.����-T�Oɞ9ǭ$D�T��Ń�i^Ļ�N�F2h���-D������~�(0f��n��P���,�O��I8p<$ad�<��"f�G��C��2}�(Ԙel�;) y�gGI��C��w��%����aFDHT��LͦC䉴m�D�B��7\�* k�L¥,<B�;��R���4Tp�A�@�M�B�I# �ؙ1�]�]h����_�6�C�	 � �RAX-*x��c[	 �pC�	*gLl�+�#��p,��E�9��B�ɬ3ct�Q0KB�r��]r� 8-��B�ɔ�U X�{y�����6m�B�$a@��@��*El$�m�69�`B��%'����IKHh�ܫ��f}�B�	'��XC2悧'�� �DFlB�K?��gG�2�;�
I4B�I(Z��c�Ϩ9B�9V��<~eB�;P a�'�k��s����NB�ɣErX!�81�z$j��:�B�	�_D� �BZ�+ڨ@����4�B�I �p�CP��y��HB���*yn�B�I�L)��G�*[�l�za�&<B�I�>���rc#�e�HP��j�B�I&t/��Cǀ�%F�Hv+��C�K��)�のK�����G�t	�C�SzM��cK�H���1A��B�	<}�Xʒq�����'Ō�BC�ɨ$���ߟe��·}��C��pr��	��%δZV�ҙ}��B�I�AG����4x�~�Q��[�vefB�I��>}�$�	d׺h��@X�bRB�I�fҀeb�f�Jt�F�8>�LB䉭/�|�D�-wP�e�d���Q3B�I=q��l !=�hd�ֆ
�"��S�? B\1EܢJ'hp;�k�#V�<x�"O�I���f�0xɖL��7�h�{w"O�P9�+4it�i����L(�"OV�+��
�z�Pҋ�$4LPsC"O>���!��(�cÀ�F�IP"Oֱ�Ӌ;!v�m��S)�P:"O6�y_z@@���b'xi�"O�,��R��, �� $\`|�V"O���Я^$17i��I�$P:��g"O� �ҫE�?�ҍC%�S�~��X
�"O��g
��Y�`�P:�̨S"O��#�OY�MC�0ivo�6Z�6�0"O*��á�,jeD��#Ӥ/���"O@��e��6��h�&�/y5n���"O�Q�C�I<5���Ab��DĶ�1�"Onl;�*R�>�&����}b�X�"Oh�3�%V
T���ZWFt&KR"Oh��t �8kȖ���#�_�!��"O���Z(N��P�R,$$Ɯ��"OR�@QJ�	�T8:7d[�| ��u"O�(@gd�`U��%�>:����3"O��	 �L���cN�n�� 3E"O&��ۆ9JƽA(گ����"O܈b3�Wg.�3�D-n`�r�"O���W=~�J"��<j��6"OZ���lU�a�&����H��	�"O��[PA�i�X�3�k�&��: "O*��G`O<|%D��é�9	��p"O�p��AL�Db��X�ϕ+�����"O��
�Cy�N�5F�h޶E �"O�(chҬ]�|�c랅~���!�"O��@����ع�݃s��P�A"OȩQ� �xvT�;��)D��1ku"O"�p��T1��Ţ� �%���CG"Op��s�	��¤��a�'rJ�Xd"O\�r3�R� }��#��؉b�e"O8�����x>RaF�g�pIc�"OZ���9�<|�VO֩*��{�"O<�ɲi�:UDu�7nS�K�|a��"O4X��R�>֍�v�P�K����"O ���ß�;�xl�6�\��>}(�"O$��'��6E�Ѓc�Ȉ�"O�d{�n(8N�h"��7B��,c�"O(�8vD��H�����%�ڰK�"O ����GXh�VC\9V���)v"O8�9%��|����D#ЌX|�y�"O>���
�-e�ڲ���"ЪB"O���L�H>d���D<c0�2"O셪R"���aM�y��Rb"OvL�)W�_OJ��b��g^l�'"O�Q@7A�/3��P��ΆD�^LӦ"O�|0`iS9V��8��]�E9�a�"O���1lȖ?�@pŢ��e�!��"O �PR.D�T14�ׯ�!O�n$""O*ZXX+�GU�@���C���v!��\/�ճQ��9dm�\ʢH�� E!�Q���I��B��lX $�UG,!�|cTP1aG�1��d���!��f�H1��P���s�!�а��T2�F ;q�d�g/�)JW!��2�����
B�0�S.X�M�!�C�X��@��y���Tk�5E7!��6Xa��
�[æ�5
Z.N�!�$,)F��)w/ܲt�d��tBU�'�!�� =��D٘,f��Qb�� 3�(�"O��0v˛D,�Bt/�}|�I9#"O��H0��c�,�R`Ѷ`R�J2"O^�h笑�RW!6�ՑO�`{"O�2F|�T� �χ)�65Z�"O�����/8j-1g.K�RQr`K%"O���@�rZ�RA�S>K^����"O��;��ľI���w+�4Q�4�C"OV0`�HM�>��}	��+n���""OdP� 5�`��I�;#����"O��qp
V9�M�@f�;���"Oh��X�^�&x��BQ�~���*�"O��KS�!=r݃�V�E�$�"O���ԭ�Pi���w���>�Q"Oh��˚}좭�$�B�Xa�"O@��h�}�(0�	�=w"1w"O��&K;:�m�Ԁ�1YZ��+V"O�PHQc�l�(�k��0�n�R "Oxe1/�&��=��6&`�S"OX�emU/����"�!D��5"O8,{&@�	Yr��f���$	�"O� ��ɒ�&� ��IV�b�t���"O�X�b�ͯJ%FEy��V�lEYt"Ob�$n0-�4�X7DH�ͬx�R"Opq���F�ó�)�r�{�"O��`6N�1H}��E�U��Qɀ"O>�3��G�d�\��f�R����� "O|����˗sѦAc��B�O���"O$}0��G�9��I�J�3�@4"O`]h��؜#0�xr&��U)�E��"O������L�
$��#��� "OA���ǊQ̬�󥎽w�t��"OT�E	+S
��҅ĥ��E"O>�@�˃*Aj�݁Cf/5zF��"O�(C�5u�(�� Iw>�9 "O<�*b�Մ� eɣ,N�
r���"O���Hǁ>���x���7
�� S"O:��!��r�6�C��%qþ	�"O�AS5/�aP<[a�����B�"OJ��)�<�j�4Z�g��(E"O�m1&�0�N�* Ah�*̫�"O���� S�#PܓP�W�S��A��"O��`�P8;��j�͎3$z����"O-z� -B��k�C_f:�aQ"O&(���[�iD��a�
�����Y�"O��+��ռXʠ��1�يE�08�"ON E�Qy��B(C~D��"OPEq���; ~��&V�Oς��"O�������(i��C�T����"O@�IJt>9b�љz�$� �"Ov���(4��ad�F�����"O��냽?p����f%��;@"O
Q���Ϥ%(���$E	T�M�d"O�P��ś!P���� ��j�J�"O�̫���H]��iACN;dd$a��"O�,��	+
�X�3��xt��9"On�YKC��֭��`s�`1"O�u�q+\�'>�|���Da�Ѳ�"O��
�FF�M�-���߾B*H�Z7"O�(r�g�4W���c0� �Rv�ٵ"O.4!�Cύ��l �B:��D��"O��20b_5<n(�BG+�t��"O�����0e7�E#��3�z�"�"O�����5�
��"�V	࢜��"O� и�ciS+��u�S"�bwt)�5"O���Qx��^�/(!��"Ol��j͸,��#So�2 ��$W"O�]�t�ݺfثg�/o����"O��{efI5O��L��Y��l#"O���V猚�F�7.�7ch,hC"O %�g���8Ur���Wy�1�!"O�)����%�𑑋�0��t"O:�y�`�(p��H4�!� XH$"O�1aӄI�3�F��4���n�g"OL��C��N�q�d��h��`+"Oj�dӝ k8&mވIאh"O�|�A,��T(p,� ��xX�"OZ�;���M��C !�'-(FH!�"O�A��Q��ؑ�ӒA�\��yB��P��A1l�,/�Vm)�Օ�y�P�i�j��GJM�.7�9q�Ȉ�y�_�r�� )��*(�|�A�Q��y���8T\ I�Fo,��� ���yrb�h�Ai�I�/c^܉X�˃$�y2��R��0񫚟c�`|��U��yr��PI�����a�n��+�y�,��(0�8à 	�oH�t�uk,�y2k%~�Z����4*xT+�̒>�y"+��.��i5$@00BN�(O�
�y��X(�02��=�����G7�yR�U�K
�J�*�""	���3	���yR���|'�I�m�g���D��y�Ɯ���H���J��p�����y"3V�!`+A!Vb�a�����y�"	&x�b�����C��9��B��y�⚴a�|}��c՟=�ĥ��S��y��=!�e�DHP�Mw�������0=�AI*���fK�I�P������K�ʐ� � ���v����<i���I�2��B&)�)D ,���O�b!�kaf�˵jO�r���[U���}!�]&?ۘ�D�	/�P`���!�D��`��a�RA\�UȖd�W �1O�=�|r�B�2-D�)�歀'(�@�k�<	�e�Nh���8����w��q�<�F��"@k ��_M�l���Tq�<9M(�r|���|��J"�c�<�eM��|G��y���?�T!C������+�)��<���\&=���S�B��`�0�:e�E�<QvkH.T�0�-Q�{�^\���C�<�����X�$��C\�ı�"Ѣ8]z���H&|px
�ѴR"�Dy�$Oʅ�%��ᆥ��޹6{���"O�Y0t��u$���G\���[�[�PxR`�@2�DɆ!�<!�� `�G�?������<��փA��R!�A�^��(�f�<�5���5��e�s�Yb	�X@.�c?���?m��a�5e	h�����6��a��;T���&�	)X�P��͟k��ņȓC!&�j0��8[P��"��ƸFy2�|:����'{<���,�_I�̓��M�<�B)��*U�	��,O�f-�u˜H8�&�4�1f=Jȅ�.�43V5Y��,D�p)D��!0[^�� G�w�n�$��OV����"�Ybb���� i�h}�����f<�B�	�}"Q��(�M��@W��.s}�C�	d�1��=NتT+u�T�C�=#o�uS�ރ2,�D��W�vPC�)� ��R�j��s�X �B��g���h�"Ot-X�KT:X��lc��E� �'"O
�8ac\�Z��S�K�$�.�[ �'/ܣ<�6hȣO��5@��@x��O_r�<)�A�?���(�$��-�rp[��VY~�"�S�O�X�ЁǢ-ZZ�#r�� j�jԻ2�)��<��E����'��%E�4�;f�N�<��g_� 8<rv��+�t��R+�<���	�VL1��6�-M�FܺD��`X���O(�kb��N�Xr@.O�6�ޘ��'U4��'�X]�3�#����F1~��1��D �S��� k~@U���p���j�bE���Ob�"��\�4�Ы5Ĩn�%#E�kX�P�O��@�/(�fh��E���"O�k�@-��հ�hӠ�p�a�OF�"T�\�~e��:���0������>��=n�`�Y膂7��};��c~"�'�⩕'�~PS6�6XD",JCY�m���a���$��!j8�W`��A�)���K"�Ia�����мW{��"8hf�l�Q�"D�xPv��<{D�4r��]1$s��Y3?D��1h���C�[�t��C�`=D����E�Kf`y�"��j�`���<�
� )| �0?`�Gk�l�tن��]���HY�)�����g��X^�ȓ�V�AFjS�|00\��6^&B�=��2�S��bx>��'�M,����hV�y�|#>Y�2T>-�� C�]���h�%Ư>�`��� ʓ|Ě��DԸr1�#�e/�������;�8�	v�O�2�c�E�rB��!a��P𖆉Ӧ��\� �@"`��Ilҫ^�T&��D{�����ov@��Lʘ.���ke�٩�Pyb/Fobb�n
sF�Z�C�Y���=��o�IA�Apņoz���X�<�kPt�&��E�
AF,̢0iS�<��ː*�X��e˹nစ��R�<�!ƭc(�m��d�1L�~���FM�<��(��Q��.	.��`2��~�<����kZ��b�=E8�p�ĕz�<y1 QHN����.;�Ƞb�)KoܓodD�<�M<y�&΢=�����hI/U�����Joh<�$��Eڜ�˓<I�&4�cB�	�y�G¼s�2���b�'F�*����@*��'�ў�0 *�s��E�V٥t�4��!"O�I�ㅿ#�8}۔F�5
�d*�"O�����r�È�h(&�P"O��(T@C�td�[�:hUi'"O8pX�皷9�ܼ���߇Z�4l��"O� ����3ސ�R�"^u���&�&|O�IrD�!D���-D�t��X7"Oh�aEƱHފ� ��ǀ-������'��;����Y��0��/�#���Ij���hs�ϥ
s���p㟙 ��H$�*ⓥ蟂�B@.ד`�q�C�M/�H0�"O�T�wi\$%^�7�w�� ����0�S�+8� ��Y�FHћe��jvNB�	=@.~qDN�^�E
V�Ě%odxK�}r�i>�#X�a3���;��)P �������If?�b�#j��%��������J�/�M#5Otӂ�KM�`EҎ� n���F\�W-`�9AA��p?	�~���`�5G�y7Kҕ�R��Ue2D���Sffi�L+eNdKv��g�ay�P���OtY�leJ�����QxyΠ��- B�Iz~J~�<��X�s�h�ӫ	V��JR�V�')�?� >9�r��?(e6d�E��-#�X�05O2���I�[����hį^Eh�����[����$?���
�^<�c%T3I]�P�[m<�~�P��#��fTp��DȱYx���&&}��'�^tR��N�������Pm0FTK�O&b��E����FnP(��Θ�B
S�/=����'��P`p-A�>����4�W���}B�)�^8`
��a+ʹ����.X(!�6RD	Y�/B��%�iv�܋���>O���c�Ԧ/�����P��(E"O ��O�"^����Q%�%Y���u�x���=��i�6�����(�)Ѡb�A��&�F�<�����~Z7�D�X��V�ބ�c�,�	]�C�ɘJ�ֵRA�G
9'(Ղ¢�a�D;��C�'����e$�-a�܀K��ܝ�@�'����uj�xK&�Ǻ)��XL��E{���.Y��D���a$���K��yG�+6�8��
H�`����1,C���'S�'Rўt�ڀ!�\�@��[
.���k'���ɪo9�5�Vg/�L1�%�Pb�A!D����J�2��
IRp��|a!�9�D>�&�ZI�,^+lL}����W��L��uH�y�#m�XI����J��	զ�Ex��tR���ÿEz�h��HVG�0��:D����cG.�6�5G�&%Nl8d�8}�%�O��J��#G-�{�KU�Q�"L*��'剤V���5��,qr%�eE�7Y6C�ɱ5"hl�$rQdBgP,ӸC�	v�Z\�6���k�x��1�lbC�I�.��2P���(�N��W�&>V�C�ɪF(i�&.�
S��ر�,e��C�	�]Oj�2p�^�b�n䒥"N�,x�C�I8dm�%ϗ,L<H���k�C�	�n��Q�FB�L1Z��J�6u�C��7a�@QKW&(N�pM
��c��B�6O� i��R�N�(A�&.D"�B�	)�xʣ�V}���d��2cQ~B�I�t�6GK[G@~@"B��,B�v����Z{Z�h��� ��B��7M��xff�U�8P`�a،#�nC�	�y��4fFA_�$�w*�	_j�C�	�&G��g(Ӵ.7`��,Y!� C�	'|�h��q��C�
̲�Bۇ"��B�K��1A�ƴ�&��$�C!9)�B�ɃtFd�����+U����@n�C�IReZ�xC�إD��bvM_,yO�B�	�"�� ֢��HT��j@�1K�B��D�0��
H�<�`�YdJ��x�JB�I�}�`��j��W�vp�'@k<|B��(,����U�̹.hL8v(I&�C䉠7\`���T9Sv�aY�k�_Y�B�X�00j�D��y��y���V�T
�B䉦G�p���F:x�u�a�:��C�;��k�Z�x��a'GT�\�C�	�b:����XT��`ғ|Z�C�.���5�P+��,9�A\"�B��&Fte(1K�;*r H��^hB�I�h������8UB|��l\!E�nB�  D4I'�E�"{��H`nY�7�B䉞�Be�e��%=n��DL X�C�I�UpR�I���9AA,Z��$(�C�	�5L�)�/��(��߁a��C�=X� ���/~��5Z]�s�(C��S(y��A�G��y
��2��B�)� 0���m鎤�.�(n�D�Ju"O��G���h $BL*���Ib/�*j~
U1��@�E-�����'�����:b����'BP��'ZH��So��UУׇ�77�	��'?���,ۜ�Ay���{�½��'����CݔK����&�U�vu؝��'o��&��<F�����R��؁�'�����` �V��ըGE�SG^���'A����
�0��I�b�>UL���'�pݩ˔n�2%�� �
%�� ��'�!��C휝�C���*ف�'����DL_�3��0��A�]+V���'��i�F�'�֨(e'Q4Nj,�k�'N� @#ʮ7�@;�bR3Ǭ�
�'�J��S�ǂ0�p�s�HuAx�K
�'�K��T�WvX���ޝP8���'8�������#&�9@4��	�'�r�.'K*�Z�j��r����
�'�B}����t�[�NѶd>M3
�'�:�Yǆ<K���Gk�e����'�*�H��=:�h7��(�����'*U��F0�l��m _��H�'Y�����"��!AF�1[�����C�`�"/��(4�s�eJ�Mێ̄ȓ"��'�C?+bh]["�F!G��ą�u� P�	�1Nm�ed_���|��
��T��M&l�I�N
5!�	�ȓz�L��f����Y��Ƭ��\���Vp��լ&���(�.��хȓR���cV�7P�@���-g�Դ��%�ѣ4	��/����aK�$Y@���ȓu��0�˅+z��b@%�T��ȓ6✹��+�P纅�uH Gt"͆ȓt\���ʼ:mDe��EŦgn�i�ȓK������&4��I%B����x�P�R���"�6�!�/ �KQ�d��O�BćV?*yD0���D30$��,E�͑Ԍޒlg�*!c\�=*��ȓ8G8�X#�Ù?��m���cwLD�ȓa�Ei�$F<8
�bF-ρ<}��]�� &N�.R@d9R�Z lj\�� ���P�M:<A�D��i@=��9�r� %#ͮV�V5��M^�:����ȓ{}��ѤU�F�8 �X(Slh�ȓ��%����4B�Q��BW||���dд��d�F9T�����_�
���R�����NF/a�n��pG�}�D����*�	w�^o�J�S G�����ȓz;V0X�IF�M+V��E��Q���U+�5�o�E��,kr [���ф�hFe�!�o��x��ͽ:� ���I����GW���_�����(�Ⱬ��#D�P��@�ZZ|�B�C�"1,� e?�	��N�����W�O��Q��S�d��;W�1;�H��'1�h�Q��s7�D����G����f#L'�̵�OZ��G�3?���߸6��A���}6.�1gG�p�<�`'�NF���ř�m
`�1EGЮr�a���ܣ_Z�����5}T:�8�✢�$���֧,vazR�	wB�u!K�V?y��ܖhqֽ�sN��cblI�c�R�<��V�hu����ȟ6 �l�
N�!�b9x���[�h�~�P�7 �28C1��M\�-���|�<�c��a���U�R,a��<�3 �;�"� @F:}2��	���ɇr��ԛWL�MV����f^�1�6B�	�.̄p�`X�Y=����'�>~��ˢL��ܐ��Χ� n����#���$�Z�B�(���'�U"2͍�| Q��(�sn�c��4�Եt�Х����TZcj��pmP��*\�R� ��=Y5.�}n� ��)�ZX՘aM��Vy��pvkIZZ!�$���ؠ`�ެ'�����C���(0���8�tM�������Y�4��MRX�a��6�Z+�#D�lӶn5%���Cm��0�:�$$A6l��)c�y8(�B�g�v T�2��4_#�l���ݾ-B,��	��
b�*}��lZ�e�����2��U*R��ׯM&E[�}b��)+"���l�x	����ܣ��Oڔ�ZZHxP�/=�l}�`^?�� ��!l9A�rd!`5&D�����0V4���V�Fz��g'�����LP�_�\y��>9�v�G���ͻd��q�"%~�ѥ�V7�?AƉ &S�!Z
�&�`,��ǜ��
iC�Ԫ
$�8Qb�ƣl}�)s�ʐ�V�B����Q�ܴC�RM#e
C�%D�����F�d|cG�C�
�ʬ8�(� �a~2�bS�zo_� �R�F�2�1(#����=Q��ϡ7ln�2`�dZ����$/T����,�q��B�����i3EV$�G{o� w�`�ؕd�5Df0M"���H���Ғ{^�C�M�l��ZA�E"7>�G%A?0�Ь�'�� D�,Om�S��dZ�%3G�ߵ��|*��'��Xa�E0v��m� �L�G�
u�s�S��l\�#L�.
�ui����]yF,�!jK7�t�b`��a{��Ҽ�h_�4-�6�Q�;�y�!͍�?������k��(���_w8=-)��h���i��,���*� ��ox����o{����*4y��㑴U�����[%I�D�4z6u;e�_!y_:\���J(2i�7#�<%?�A	�6?Sf5:1!�K�����hO����4:X~J�]ײGH]H���TPI��S����n�6� ��J�D@^MP5��=a�p��'WE�,O��q���\l��c��C�ډ���'授�F�;#�&4Z��*:��#Q��9O=䀂�-��<Sx�[B��-5��P��N){�<��CE��$ua{b�Z�x#�eƯnSZLB4�зWJ��� �3Yd��F��&A�Q�Oe��ؕ
�O�:)�v��O�e@)xP��,O>?)�D�c�'f�왡���(�LYz�L��_�n�sF
]�	j`3p�'�Z�ӵ�V�e��傰��6�\y:I>��P>��նjc��ǁY�9:`�3�Y���6���(�Q�C� 	�e��E[*AϾ�qb�B8
�6���_P�<�O�e��Ν�f���rl�*_&h�R��O�8�6Ǉ�`,Z�!C��<��*G�J1hsrb?��3�N+e=�Ј%H���Ptr�>D���A��z,���%`2~B���+Ǌu� G��2v@2vC�f���O#p�D�xQi`%���4��m35�՜İ?��h�")�d�%  j <�%��2��X���V!|\�V� �_>��)	eX�P��ۉG����'�{�� 6OL4J@N�<�p�C�����L��-)
a�����U6 u�f �`�h��ēYq��SP)ە&*��À�Ԡ"�'���ǡ�(C9@�#v��s >E��%��ƹ�/����&�h~�B�ɌwPVhR��C��ڧ͝(O�.]T`z�a1�˵�:R��=�}�O<���@��f&�錽c�w(<��T�.}��nU�r�N����հ3+��%��%I�Z}(�H�(_Z	�'�ҥ�p�䁒sd.4h#�Թ=&�!�Z=Mo�x� MW�n��p''j�0�i��\��B9��N�5ZhsR�L*a����'?`���Y���j�i�"��g���s�^��t�7}�o�8&�̍��I�o�O�8���K�	�~��d���N6X���U6x���'p��&�<̴U��g�Nu�������I/��ls�18ْ�`�{�w�j@Br̆B�phB��M��)
�'7(9�j�USv���	�;>�q1NZ+�2%�V=Mۚ➈���?§n����t���(e�c���'�>]�㉝o�f ��	ϼ'��	�8_����*�X%R��V�JȆ�"5<�r� +\O�@P�E�"wF�لH�����x�I�� �:��|*���#TFb��ŊFȥ1_�)�h�	q�8�"O*�x5Ꮧ:�j��0l� �33��Hܓ`ڑ���L�̚Ռ�*��as�.�%2z��3//D��b�N�>���Ph��[ht�y�*&D��K@��'8N��(��{�~QA�g'D��Z�h؅qx��#H�1+{BՀ#�'D�x9e`���p"/%i�(�G6D�ؐ���
��	��X�;��IH�%5D��!S�6{��T`��+�D�5D����g5j,J0qcK�4���j2D�� ��ѭ�'�l,�Vh�y�f���"O8����*���Y�Jb�y�2"O��1�#H2���J��&Z���S"O@!��ǱJ��s�ۤ&�u�p"O��	',0a�JQ�	CW�""O2����D�-EH7H[(_y�2"O��Cq@Q�AIp5�A��#j�z�;�"OLl� lB�&�����T�i���z�"OrE��!ӄG��zgB��|y�t�a�'6(�R���>4V�#B�
p�f$H̉[�-��n���@\�U��:S��	?.�'��"�I?y�č�皥�O>���}�P�Q�V"r%�Q�C�D�`�n��Đ�L�b�`��]>
�1e��4�8��F�<�?����PA�T�p�3}��T��<F8ܱ�×*�(���K5�I�a��V�'��xQU��\�'[�����C'wJi
s�[���<�'�8����͵R��yr�|��m�Ԟ|�OU\�O� ��|y��N�v5˩O��t�
��ēq�`��)�~��Kٌ,�ꡋp脡:ܬL�AA�~xx�*�*B"�J��
�8��>E�dH��4��f�7��2��cf��4Jc�����Yz���Kj@y�fۊ}�A��|���ٰ$�;=b�U
DG��I���y�)�8o�h�i˩P�� 
E�+p�:�� �.����'�Z����+4?(*�JI��S�QbpD:t�U�=Z1�"/P��*22eZ�s���1?r)F}�b�=/��6gr�d��j��4�F���H�AZ�c�(��j�P�Ꮚ�k����Γj����[����?Q�P�@�g����Š�u�t(���6��\�jͽY	��	�.�xaɐ큭��tc�i~��w	D���b�o�%�h!�� ����)�<�F��E�� �y#v!�!	�|���'�=�'(�FA̓q�����.�y���>��ኑ9X����;��d�ī�<q���S���S�%3,Ox]@���N�(=�U�<V��Kw6OH��i��[�2�k�EI9ve�&�q��bp�����م1(ذi����9��(x�H�~J�T�N�t@#�L�#X�=`�߰&S҄z�L�&#)��
¥��0�҆��fF0m�!X�)H�K�p�i>��JƆ� �eH(fx��E6�)�nt� �^S��.�ZD�ӍL��PF�`Ԏ���-�4�8�	 d�~XV��"K���ϓ�i.���g_9G��~�Y[�l���S�O2�\��!W�9�4*V�t��
�'�,��GZ%V����)e�pQM>�$�)d���䛳f�ʐj��8Rԅ4��1�!��%p��v��3@�Bq��
�*�!�d\��Â}z4�BvJ�e�!���T�ue��eY�yB)�j�!��7L��F���7B���@�Կ^!�ė�^�����/Tʩ3&X(�!�Ě�t̜I$G6}It�
��Gu�!�dA�8�$  &��J���x2M�	}�!�d�l���A��� ���a���8!��:�|�"JP�lVL[48�!�:Z�5A�����8��	 �!�'�:ժ2��/�4��Q�A�l!��G$$���a�J�R�\�@v��%>P!�!`��K��W�nd��-��>!�� zr�� 	
�� p���0�!�$~Ӯ�Hd�F�/\�Q�
%Q�!�Ğ3C	^�sB�{�ks��g�!��	)v��1S4�W�o��=�q.H
K�!�DC{Ƽ��=Bǎ�B-��(�!���<���+�Eݘ �^dQs^�s�!�DD�_�`�*�i�!$�rw��>�!���,�ʠ�5� ��A�����av!�$�Vk�8�ә7��)1�nϴ�!�Dϡ�*��+I/>HqSȌI�!��=-�6�a�+k12qD �#�!���p� 3��̚6!��h�z�!�d�;��ҡΨL���	���4�!�Ċ�#�"c�$�*a��@�k�!�DJvV%H�f�uw0�b�ʩa�!�V�`�jݫf�j=*� W"T�!�� ��u�QUJ�Q2�=b�id"O���kW�&l(�[�I������"O>�0�Ӹ]5�Aj�F�-�H�G"O�,iPJڄS��A1���3l� d�`"O�Y��/�,�J4�����i�#"Od�#h��#j�H�ʟ�A���V"O.�����H����%	T�>�9!"O�]3,ÔLW�-��ɴ|��1��"O�	cq��K �����ؼ-㘸�t"O� ����0㼽����f�N,�Q"OL�)AF�.�>���-�J��Q"O�UB��V�0���)�@)�2OP�k���2�)"�0���ȓ~��T�%�M���B2��fڦT�ȓ/�R�jD獩���Z4��hL����W�>[3��0H��;�i��"OD\��Nӏ,O^pQ��'�⨰�"OtU�v��>s5��D�Y�LN���"OFQ��c^)<2�H�jِg1 8r�"Oj�ㅆR+~�����ǣ^>zIsp"OiR���$8
*��Ʃ΄*�pC"O��a�@l���.I�g�T��@"O�L��ą:h@ER0��&4�ਁ�"O�U�s�54k�Y��f�5w���"O�,qFs��#7�_�Sl�,aU"O0̲F(��N���F�%Hv�#�"O����H�S���U!�TC�`�c"ON9YBԀ#{� ����&�4"O l��'׳R�"a��k6O!�LB�"O6�3�l@�)^�d[�I�@�"O�a:���UE�P̅-�R�[Q"Od�"E/G$E��e�J[8V؄İ�"O,�p��<wɀհ�?-�S�"OH99�ԯ]����5�Q�Q�"O~���޴_�8����,y6�q�"OBe��ʡ<A굋���.��D"O�Iq�����@'�4et����"O��uc��XĦt�@OJ�"\����"O� ��	}!�)�7(_�ސ�"O*�!�98o���Ί�@�:A�"Ov܈D����tض̀8>�Fi��"Om����(¥8&Q��,�y�"O� ��W/t�[�f��yOR!"OrYChb�ʉ�PE��o"X`G"O�,W��m2�a�Nޟr/���"O��Yr�S�a\�@T�Od�t�Yw"O�LۮK1@ad���z��@"Or�r���[�������D��d�"O``&ʌ�S�<��E.�L���"O(������JUjA�	�Z�0�"O&�"'_�D
�8,�/[���"O��Q@ 6�8}��	]�)����"O����ږp�"�a���DӖذ�"OV�q�8I�� ��-B4Rՠ���"O,��=�0��O=���'���Y�GYcyB'4�I��#L]m>�Xf�y"�
�P-R� qb��G=Z��@���'��X �< V�?}RP�d���фF�)52٢�@<D��`�����T����rj\���K��>aDTy���Y�E0Ĩ{ (8�̄��a^�F7!�$ǎ]��6o�-�V��S-3v��E!��m�J��
�NBp�	g�S0&,���79>�\�鉘�Ƽ(F�Z�j�d� (�SC�)
5�T�uLLk�!��X�����g��+.��e���^�1O*���*F�X��ɑ��� �ȱ���>�!�[:4#�)H�"O�B)	�h�B��ϒj�Vx� �Ѓ�4�� �>��c���$�	����4��Xkr��D�Zv!���j6δ��픃\Ma��^!S����͉�B)��h��]k�FX�x����-\����	<Y�z�A� V�W��d�4S��,�b#~*�4;O	%<$!���	��3B�(D��q�ߣ*qO���O��"�G�_�1(������YlD�<ё�<l<4��A�_]\�p# ���ȋ{�G �g}�dB�!~��K���o�صX󣈺�yb���B��xU'.w���b�Z�yb#�~�>�qf�M� ��w�Q��y�&_Dyxa��ՙ}��a����y��;
U2|���<��ܨ�M��y�
@�j����Š�F�Fu1$bt�<���:y�x����ۑ�B���t�<9'�`3ܰ���4;0x	���ʟ4��:X<D���<-8�3	�QV� ��i�8����S���'�OW�(�Sk�>��I8u�S��O�楳4�Wo
^C�I�ID�hqƅC�:N��qwN���7�/˲d�r�i�ޕ���)D�()�E�<%?�� ũm�t�A�X�a��t��=\O`
v�X�8�~Ip�',"D��]�M	�=����>#��e�Cb�\��E�Ԡ�<i�A/�gy"*�Nw\�[Bm��#~�x�������']����DU��}F�dAX�4�^5�����eƐɖ�3��s#jT l�2��&,lO�$��p�:9��(A2��1�вL�lD(��>q��9�ĈS�I�8s',R�Eś��@�,�ڠ[r��#L�tXq���y�ȗ_���hU#�N�c�n����h�uN�=9�X� ���>hKp�	�_� �S��]��]Z�I�Xy�!k`����DB�U�x����X-�y2�Z�G�����MZxؾ(�嗑u;��+dK��+ߠ˓^Bڣ|�',�����J�p�+ދL(�I��{"o�'�0�"a�Op�O�&(���2�����E�		��K�M)�-�ѻh�Z����^����=����! P�xs��u�K�z����O�ͳK|���O%�G'�Or�Ñ �l�:qR�c��p
.��"O`��U�><B�9��]����E�i��1�'G�4�����UP�L����:���V�d ��?��X��_?kz!��j���=���"[����5=%<=��߭oш�Z��Y&��"p�3$���Z"�r}�4����N(��#�x%�6�B�_6c?��ak�5w��iV"���k��5D�@�f��$�:(���]�ơ���O�X
-R�$����M�"~�B!L��Vl��j��p�EH&.I��y��ЅW[��qЫS�_� �pE*J���.Mwf)b`#U���<�����X���-[�=qdH*A�GUx����mۭ<pd@1�F�)�%HE$��|��-��MZ�V������VF!�� tC��0�J-�������'n-���.[,v�.I��^���jŞV��
R�8B4l��͇��y�%�-�i9��(�R8�%AY(	������@*3Z�(����xBHS(|@�ͫ�KT�UȀp�C!���Px���?C��<ҶI��-p��Ip����rdiL!i�<��"G����G���A7��KH���[~�(��I8iK:@�&˒n��P�ѡtz�)K�M�\˲H���	�Up�!�"OvȈwki8��j5��u,09���>q��52�@HJb)3�L�IE�.o��"�Vj�ȇ"O2�����,���+O�Y҆���f� �E��%aSA,�3�$�}0�;�Ύ�`�|�9$��*m����?�PF��Jg��a�"P�b5ޥɲQ`<���C8U�W�C�!;-tP:���	�^|�,Q��	hU���C#ìШ루P)m)tC�I�1J���EƗ1���8��û6gpOH�!�G�uo̒O��*�`GZ
C�1·@l�t�	"OR�r��;dJl-i��@"k;�B㞔��]�g����ar~��U�^d�^�aw�A�"[!�DݚM���5%ޥY�d����7N!��Z��UaB�k%q��L�D!�Ċ�*�r}PbΜ:H�V�8���(�!�� ~��ņӋp�I1��ܡQ�"M1�"O�A�T��X���/�&TH1"O��Q��M"v�h��h)@S"O��K��T]D�D�O���ٲ�"O���
֓T���'�8����"O������d=��T�\9Z�"O�*�u�������q`�"O����[��|�����'Y����E"O�����B�F
#�	Np��5"O�͊�+M?d��rG�ŊN2��{�"O\�v��P��ML�R?��k�"O�X�'T�>.$�b��-W����a"Or�jb�F��jŒ��]��R�'V�����7`o⽢w��*�`f�M�Gm|u�ƓqV<� �/PB&��!�@#UF}r������5�i�q�P�2�*3�*,��ġT�!�٠XE S�#�+�0�Y6O��/�$��':\��"���)�Ӈ.��E���z���7DUd۰�bę�X!�6yR��[�)�;kͬxAf$F1h�ɘuЊq�"�ɍ`0�t�f�
��>�%��SL�r��2�S-Y�hM
�Ǆ�4΢?�q�K8N�f�<f�iC�݌e�8�����' #�q���J(t�lTa���	Z�`:B�_�j��S�O&� P���?��YG��Sʒ؀�T����D��(� ���8ڄȁAί'B��>��4"Ϲ�ֵ㗸R�%��@���$]:}����%��<�gG�>r'��Qug��n�(�����<1'�NSz����+R�Z�th���dٱפq�z��@O ~���f�Ҽ@]��A� R�qN��"�a>�O�� !_�mV<YτPc6tq�J�T4v ��Œ�yƃ�:�5�a
T)�O�Sd8ҧ���ǷB�l��ѪW� :Ej"���O|hTH�?�tax�'�f�RƴG��h�%'�|�A��"ߒ'�`lҀ��Yw�9��
�&y(�ӧ��b�Bg��:����-W�~���ȷ��X�%P|�R�3O�p��%�
bxpj��$A��\����DaM�
��T*.պ��$�6y>��iX�հ<�1"X�3���W��Z����W��<���y^mٵ��;y��%��.���+�7w��s2��1�"����R�8�`����W�Q�}�/\�UX`��$N���*�*AW��5`2i��lI�\�T:�z�,��Mö$�
��"N>�'~4>�劍o�H��I4bD}R��[�����t}��?d�!�KEUv���O�O�ڍ;2�<Yt%W�{��㞢}���ob���G��}T�0s3)H}�� �>W���R�|��Iĭ0��AP:E��M;B��>v$!�d[. � �R��F!�2��� �3�'�6���D@OX����k1��r�kӉj<�{� D�\�s	C�<��F@P,#ȉs�� D�����H?-��H�P+.9�Q��-D����\t,l`�Ϗ?�nE��+D� h#�,��0�c�p���`)D��Z�"ɵ&�^��L	2IV!�%(D��bs�K� `�i��H�I4~��Bj(D��r H̩D_d
E
�d>"�&�#D����F	MZ"|ېe̠`�$�"�l?D�$��-U&hl�m@a��8.Q���:D����o�
�0��U��.@�HS��8D�سa(
%�H�A�ZP��O=D��y1g��\� 4�#W.#�� �8D��B���60���X)``uq�7D���R��9ml���nM���A�8D����N�h���CE�t�f0���=D� �����FiK"�=l�<�i��.D�D�F+� ,��-�� \4�(0�-D�`���߮,�I;��P�XR��D�&D�4��Dܘ�VgHE'�xz��%D��jT��2U6��"E*��w����� D�8{�n��A"�b0�R"[̤-"2�<D��5״-�b�*'o�~�إ��8D���hř}l���B��!8��S7�*D�0Q���`�%��1�����<D�*��%1BL��n]�6�����O;D�� "z�'ĉM?`�{��E�VOl9��"O����iN;h����k7l.�U"Ot	�uC�$�B")�s�z�˄"O��h�l�w�����\�Z0`a�"O��*�ݢ2��cf�VZ�pu�!"O��� �+��kW+�E�0"O,E�`b��	Hn���Ĳ*���D"O��bO��_�tr�+M0%�&%�P"O�P��77B��(���"ܤp�"Ot�j&_#"a�4kL��Il�Es׫�*a��	Z⦏0a����4&�w�h����`�|:�"�<5������B�#�l��/��'FX�"!Q���OF�O��Y��k�;u�B�3�nG���1�I��"w�(40�kT�O9�Ȃ�d�h ��1?�Ly��'�!S�`C8p���O�>�ڣB�![��k���/v��\ ��B-=+�*��[<��ӧ���@�OMT�j5&^�D��.�t��X�d�)VbU��ԟaQ'J
�0|"��&6�Ĺ(5��!�b䀿M�ij�k�O����F@��O�Q>�IQ��8�r�e#f*��%�d��!Z7P4h�B�P��'�(�P%r��"��Y�ƪ@
�
U�'�(*�<O��� �>����O`�AP�kR]�~q���
L���Y�u�$7m��n� p��0|�6!��J��e�a�ǡu�Fdcr��j�F�]=L7��	�&��;l�*�'"�W 8qk^M�`pg�U��%柫���'E2�;���ǿ?�&>��O-�U�V8�j ��`�-	�O���p(u�,D����~Zw,����=��b�.k@Z�R�/�:��S (?�T��<���h��4�QL�)	`�"퐔4�F9;$�xd��)h8�z޴.Lh[���΍t�M�Ī�>V���d�A�W���V$���v�Ps��	6�锼o��`Ӆ'jZص�F��'Rd�Nն6�Ze�S&�!&��e�R�N5��ZUG�I��0?�B睢�l���G�$+�4����a��hO�Oj�m�C�d��aTڹ)���K<��<�Uʁ��)��9 c�A����O%�O&��i>G���TOܮG]�p2f��X�c�;F>�ؓLH�dR����է0�D8�%��+O`�=�H>�Ƿ|�2O����O!?�Q��΀�Rb#�'I�CN�eJ�@`	��6��������*�!s��%AB	������ҙ2��qPԐO{�)Ȱ��u#Kg���Ců;��U=�d�/;���$�F'��j� Q�"H�ȂL�[�!��K�`��� f������Y�=�!�H��
�yr�]�G;P�@P	��R�!�Ď�tQ��Ôe'MJ�P��G@UB!�7�X��_,�1h$?b!��[�A���"��T�r耬b!�J�nrN�u�֮I��a�����!�WS`	�&�&���Xa��s5!�D@9�+@��6<SJ��Ƌ_O>!�\���}#D992T��LŠT!�d_�!����#�D87*l��Q<!�D�"{K �BQd����m�g`��G!�[�5}�P0�V!\Z�LR��	�/�!��%jo�9#�^��>�*�a\L�!�NK��	�F�D)�Q	����!�ċ���Х$"Q+�Q��!��+�$e�@(ݎ'��a���s�D�ȓqH0 �Q�ϫB�zL_�_\Np�ȓ\.zh7���.}���^UO~A�ȓ�|=K?1Z�+�R=�64��DZ�{#�]�w�Ћ���:�xM��	z���d߅ /:DcUb��z�@`��P�ƀ؊=׊�
�����ȓT2�x���30z`Z%Ζ
+:���,�l�adk8l�]�G/�]@�U�ȓTP�����%IpNɨS!��˔e��\"Լ��)�Tv����ր"���ȓa����U�;\���恀'\܌�ȓn*�H0���B\)�}R�"O� R����V힤I�'�dݢ�+�"O�H��L�7d���S��:ʒm� "O��ZA��Bn�Ѡ'FO�aɐ�:�"Ov�ʥǇ?\X�
�k�*2����"O���� ;MqL�9r�]�G�\��G"O���ўK7��0֯����F"O�������+�r���k���y�l@�Sy��x�
+f������P"�yR�	/y��4G=K�ԽpB��y2,[xd�P8�ŇI,Yp�C��y���j��!�K�;��ܡ�ҹ�ybT�(���F��#��M#�yB&�$8�D����H�(ג��bg,�y���
�^�@���Ihb�_:�y҆�yRN!rߪ�d�qA� �y�R7C��XS�1:�lS�ƒ��y���9KgTt!�&I�|5v��G���y�!X�[�Hr�Ȟ��Hؘ��&�y��~�l�s&�S�v4I�2�Z��y��Y�H���ے�� ,�"۴�y�&|� ��E�^� [�-{����y�mՒB�D|�wN(q��A��B�4�y���Z�$��EҦ^�`�H��܎�ybBV-eY��f�#!�H�A�ܲ�y�S�Sf]�Pi�#(ًB�+�yr�[/*،�K��$#TqyB��y"��u$2A�т�zx*��1�y"kڦ3ش᱀�xt�Q�l��ybOJ�L���̀����S�%���y��6�F]`���~p|��Ĥ�y��(IJ ��
D�}� �Ž�y�'�M(�2ro٪{0콒%c���y���"g�e�wN�6v*i24�
�y���?�иY# ȴm��T����y2%��3�PE�B�hF�X�	2�ybƔ -�`%��/s�*d�3�2�y2,�Tî�p��Nj�p](Z�y�oI�&����^x8-)�f;�yr�ʇR�I@��l�`��ujȫ�yr���$�D4���!`���eP�!��6�x��w��n�Dg/\�]L>Ʌȓc��Q� J�Y���n�/9�����h�.`po׌.�E��˚�r(����q��D��JA�AH	�W �L�ȓ<�h@�UD!/񬵋��^F�%��_e+qǉ
��ժ3�'I���ȓ�rT���L��R9�V�Z9�ȓM@��S��>���R���\�ȓs�x����QX��u ���7iE氄�ob\|�)Y�p��h�W.ƈq�D��ȓE��h'A�?Z�ĉ�BN��d�ȓK��91�>/��)B4�Dt��ȓn?�5��D':�^"�m\"]��͇ȓFw�9Ub���xtqa�50%���yN�U
WfϲNưI:сׯ�Ĝ��q��X"4ȵGj@J��+2ظ%�ȓk�PrE�ɀm�q{r@��YEJ(��b� ��ׇL�>$e�$�K��j�8���#n�{֧αf@Ɇ�9&�GN�\8:Q�4�b����r�䘃ThA�b��4�GY�c����f�)�.h�$��e�1Ӏ���Sj��2��4n�5(��+h�,u�ȓq}|�k%���2�c��)v�hx��S�? 
��ՠ�U��-b�:� �"Oi���M�h��U�5��"%�TQ"OZmo�d��&-I�J��MA"O�i��_�#.�!�혷3��q�"O��Q,�)q*�1Ë8U��9�"OF�;��S�xz��f*ڹk����7"O
k��څA.f��H� Z�@ �F"O���􊌴HV�&A�'|��1X�"O��QM�dsB��e�29�\t�V"Od���_�=����2�B�t���"O�0I3�>E�=��ͅ�͊|F"O�3S�$�"	�bK�%7ZP��"OehC�'Q��\��b=P�:"OT����<v��y���9I����"O��2��L�n��DX�:Xm6"O�)c���^�HI!�d	mh��"O������P�aY��`H_u�<S΍�;|`!AJvQ��#.u�<�߁l㠽ڔdJ�XR �P0�C�ɱe3j�8�ˊ�2�\2�rC�LOt��%��*�0dY�p�rB�4DXz�9UD��mۉ|nB��@x0,��E�9���6���Q,C�~A������I�n��h]1i5�B䉽8��,R�,2��l��\��B�ɞ&�h�&�a`�SrK^�|��B��0#����0ӄ�H@�\�|�~B�	�5xĀ°��Rϰ���8 �
B�Ig	l��'�R>׮Irf$W%|�FC䉺%���PC��/] Ƞ�eNG�a�C�!+�z�X�J�a�0��H s�B�I�"X�	�"�D�f�� s�G�V��B�ɇ�>9��	[�8kx�A��]ڜC�I k���f�<uA����"~��C䉱j�TR��&�
����,��C�I�"L
(H��ؘ^����&M!W�C�IO�*��U�Mqp��Cr�L�H��C�ɜFm��TI6��A��$�zC�	�h>X蠧�6��,�R��Hx>C�I�^}|�c4J�]9�S�Ń�Z�*C�I}�0SS	�|�t-)Fh C�I0m���dIa��H[���.!U�B�ɣ3��1�W�ЕH��@�4勔KD^B��4c�މ�0a�c*�<�腼c$�B䉟0d�U���]�@�n5���6��C�	�8�ġV K�C���F��B�Ɋjb���+ۓ�",ғi�"�B��50�T����I1%��2qΨB�I>j�L���8Q�ޱ�Ӌ��	$*C�ɶZ?����0O��u��?|dC�	3}���`̝���H&��5_�C�ITZށ��>�2�1�'�B�	�>�\�j>���Fn��3A�B�	�3�.�z@��rr)� �E+U`B�7:re�3AY�*�B��6�D;;�B�Ihb�k���_�ܕ�W�ߔie�C�ɿ$?��`e$]+O�U�2��!�C�9h,�@��Y�E+z1��D��D�C�ɼp�Ҭ���Y
w)P��&oS�m��C䉬Yk���E��:+Vpma�fҳ�vC�ɥY��:].DY��fΌ5	@C�I >�q� �#V�6=S���P��B��AU�r@m��Bl��PPdC�/��2�@�	�.)Ԣ�
�pC�)� |1Q��ڸ<"n�4���J1t���"O"`���W���zD��X3��[�"O4R �9EM�(�$I,2���"O�������1��$�;@�ȁw"OΗ��B�c��"z�,��Py+L�;-�%���DM�~�KE�
^�<��l�#.|��&K���(�d��V�<��fО�>�"�'W+[PPE��O�<!��Xp 1P-A���'�O�<��nȻ^]K@�ݚ#�]�vB��/kZ��#�KR ~���N��~L�B䉻��re�ZMn�G�M?ML:C��? ^�D���ϘgX�ڲ��j�vC䉫V.����|�`EBׄ	(WjC䉶\5�eM"�,}�K��<�C�I-�]�����A���dC�&#�Y:���3ht��V�'�C�ɪ�nx{��-Y�f�p��gC�ɏS�zف�mûlJ��1x��B��&$��9��'7�zp5�  �B䉧v��4�t�S]<l��Q�ʁ4RB�ɖ1��q�`	���h%`�,H/�C��,N|U#�%{8k�m�%b3�C�-G���7	W��8h*�	�H~C�I;��P
f��~��J�`�UC䉱&r���R�(��W��O��B�I����JU���Pa2���B�I�vY*�@9N��D�Q��6B�B�IvqY��-�0�iR�Yf�B�	�z���b���S�( �!ғ,�\B�Zp���7��I#�|�f�U0*��B�	=\�����֙5���b���DVdC�	�T 
�z��N�Ib$��
>�B�
=`��VoL�W�̙��pB��-�2�S��ܑZ��b��J]�*C��n�bxQ�Lі�������:i�B�ɽ$(���.ݜ�n\�Ā�8�B�6�X}��>/�T��(��qiB�I�B�ճ�N�����tK_���C�ɧ``,�   ��   M    �  �  �+  V7  9C  �N  �Z  9f  #p  *z  ��  �  ��  נ  2�  ��  ݳ  �  a�  ��  ��  0�  ��   �  m�  ��  )�  m�  ��  @  � m �$ , �2 r; 'C +J oP �V �X  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r��EQ�( �gVlɦ�M,H"�O��@Pg�9^��@9dr<8�q�"O�Q3c茟u4P�뒤���%��"O��$f�2����� �IY8�(��"�;�g�6��I؀)?D���嘈p�l����J)�4rŭ|���=E��4a^dX�(�7#!���O�iV��p���%����'HN�+���?�|��v��6��lp��~��˙}ּݙ7�I�<.��2���?�`;\O��'�LG$�4[����G '\�Lы�������I~���4��;���5M]��A��D�>���O��u�T�Ѓuk�a�V�ѸC�00�L<�N��E�����̲d��b9���3hY��~r�)ڧI��q�ȗR��z�	Usv�,�b$�j�����d�7JC:�H��B�{�L�I�&J8u!��L$���W�۠T������,!��/��H%,����P��/32d!�$[�)�$�`A_�-����2NŽ_!�d�$
�8����~�D(��B�^!���@.XH��ِ\��h�w'�4`�$�O��J�e� C�,�B3�%}u�	 �|R�)�S�PL�Շ�W�<��E�����B�ɛ����Q�X-7	����E
%�bc�䣎���W�	�5k*�	�E�¹a%�X��<C�)c�T �*�e�ƌ{R"X�'v£<Y��T>� �K$&e�QR��-7�<�Q�+8D�� �t����n|E�!�
�I�I��F�'��>��9�F�m��lP������f�bІȓXn`@��fI�Z����$*�9h��Q�ȓ���dK��:��p)wJ6%3���ȓg�0=��`��yM��[EeN	5��ȓu�ܜ�Q`��|R� ��e�G���ȓ?T��y"̔�{([U`�,s�B�I`�0�3�Ŷp,[�D_���C�I=\M������a���R��P� ">����D#sG����ϺY�$,�P	�(l�|�x�᜝sfQq��1Hm�uY�*�)�yR�V)~��1fb^:NNԺ�#ٌ�y���d�B̘��3ʾ�0#�A���'Lўb>��V�J%:�1o�RX��B'&*�Oh�� C6��g��D�j*���؎B�	��x�� V)3\\a�En�B��:^BD��l�*�\؛�Jp��`
�'�(<ZŦI�0!2=��zy�		ד���<A#�3����Ձ��D �]eB�F�<1G�^�=3-�a@=4�hۧƐi��T~��6{|�2��B��ܵ���(+6C�I�,Q���7g������	A�P��Ys��������&2�J���!�ˢ�z1L=D�T:��;7s� ���9@7���*6�#�OX�)�(R=o� $Яْ8�RlA�"O6 �Ӄ�y��ۘB��es�"O@Hx�%�>��0S�ߐl���P�i)�6�Oo�רO�er�Y�Z���c�@�,E��(�S�'e�O�6N�{<�H���L�|�9j�"O�ыF��07c��M)֙��"O%�Q×?<�dЁ�8r�iڂ"ON��S�j��\���+aT�"ODq�R��'Nr��O
�K���"ʓA��'�.ܹ�Ö� �b!$Æ�av�)����-��
�"��y�ED��IɈ�DA��H���]�]�X �ưo�jdp�e	2f��
O�h�C�S7f��#G`�9} D�"H>M���y�)��}�Bʩ6򌙗��D�=!����p>)L<�d�!=y�8{1(�4���2��<���@Ͼ��w���b��� �R���G�fzӮ#|J��וp:���W�'_�� `fTF�w8�`�S��/^����%��AX�!��O$D�D�'(ƼmxD99(�W}�D"D�t:��}�-rΜ�1����^'��	p���O7L�+7��.d"trU�,~�>=���'V���e^yqȀ�ċ�3{�,�@�'nx�]� ���+>��TȖ V�Ӹ'�ў�O:f��I*\�t�c�lE�|5`"!3D���	��rB yjW��$ZItە�=,ON@ʌ��c����ʗ,��t���yB���QϔL�#�V���2u�"�ē�hO�����7�4ry���a���pc"O�d��'B��V� �nQ�jg��!�'A�ɱOP�Q%)1$�!HS�
<<B�I r�H���
j��3k���C�I?2 � ������OS�|vC�Ii�r���Dݸ'���S�k[3'��C���$�������&(���C�/9̒��Ö*?�H�R�2[r�C�79߶a���˙[rHP�jA�W5�B䉑r�<�����VV4hB3�K?^s�B�ɽ18h���tXr�	tK�$�B�IS#^= �l�99h屴E�Z��B�I%|����%k�@P�,��B�\B�)� j�#0�'j
q��(VO}H�B"OB\�I�8P�����=}hI�%"OzI�lV�2/���G
Ts�p��"O�59�\*&4�����rX��`"O�����=C�`�G�h7z��!"O,eA�d;�D!��C�6�P��'��	�3ԚMX׍�9-(pX�#��!Qf�B�8t8����7	�!XAIB2" �">9��-�*�{�D�4V����G!L�^<B��1-d,r�,B$h�<��� �dD$���HO?����/D��t�c�g��a	B&!D����E-w#@�����7ڂ��V�??Y�Uw~ Ё��ML$�H�@Wby����	XyR�7,��R�o���Ĉᢨ��y�M��}�
$*]�l,3�d�8�yҩ�д��PO�2X`S�+�y�!�_�Lh���ƎNa$�i�(E�$�Gz���'hNQ�W�(�j��aE
ˆp��'8qA���_Q(��YG�QҨO��"�]j,As��ۗ$\���*۹u�f��	jy���%H�	/4���@dT�>sڄ�b�O{ �C�� o��Ȃf�Ɨm樐@��+W��=�I�|ZpnW7S��Q!	��c�%I��Y�<A�K��-h��P"�!�44�W̓��=��n&3�$xZ`E�C1)�FhPR<��s�0)�g�5-+�e蔩\��ȓW�b$�W�G��<���������	N�'�}��/X��AY�!:��%*�'	�y ��,�$Ԋ�H;9Ƃ�
�'@� ��ݹp�1)&6�0��
�'�$�j�j�J}X��N�!>�6��
�'CH��s�*U�r��5d��2�f�K
�'Z�L���92&r�5G��-d�Es
�'7"	�� _��c��Q�+:Bx@
�'�`�	"�"!��@#U���2�
�'S�a��Ȇ	c ��P�D��	�'�ܕ;��:y L�q4Nۣw�����'��d�@�!��ղm��h��p�'�v�@����)��0)d�X![����'ظ��C1v�aDG�����'Mf�H��f�;q��V��I�'�\KE)�2��� AN�P%f9�	�'B���ɝ P���;O�0�S	�'�LkR��\�x3 �G�%v�8	�'�(1�6�[�R�t�!�eB0���)	�'�"��ŗ�o>X8"�1[y����'��X��A�(����a9���'8�l��v���kD�#]E�ԣ�' FT��gd@ۓE�X�찺�'{t$S
D�B�P�ca�P�ٚ�'��HA��Ɨ%|йsȄ�N,��'�KO�2䩠��xF�uJg�~�<��Q�/�0�jf��4bF��z�<a��qD������Z�P�A�L'D������Kt���5�V�PU04�PM%D��p�S'C���@ʗ<A�봬!D��ز����Ƭ����y���ғm!D��9�aϚll��X��:	q�U��?D��Q�Y�k�Z$�񋔧s�x��>D�,�@o��R��h�s�=q�|��;D�d��#�V�:ipu�'$)V�x"B;D�0��n	��P bQ�J�
�p��-D�p0'd��s�!��"�"KX.-��./D���/ϑO�\r��'6��P�.D�� xxxe�&ԌLSCO H����"OV�J��Fn�h���*E��H�g"Op���dےO�jh��ǩ $��Hd"OfG�8I�� �@'ݾl@(�A"OtMi�(E���I���M�F\qu�'���'_��'�r�'��'���'a��k���3$�x���X�D�S�'�"�'D�'��'��'���'�8���*�:4��#�O's�"0h��'���'�R�'i�'���'gb�'||J��\8�v�@��B��c�'r�'���'|��'�'���'����ڕD��pr�������'���'7��'��'���'��'}��3&�L�#���X��H�,��s��'x��'12�'I��'G��'7��'oJ �ekʂ0�R�ѻu�-0�'��'o��'<r�'U�'�R�'
�M3CgLs��!����`�'G��'E��'�'g��'�2�'8	����Sʔ��,s������'�B�'@��'s��'���'���'O�������|����S��%+�E[S�'er�'���'}��'���'�b�'���Ԃ�34����U��&�T  U�'��'b��'���''��'�'��P���8p.D1k�,
_�����'	r�'���'���'j��'���'T��!Pj\>R��l�K̟E����@�'��'�'���'��ll�*���O�[��Ԇ4�Z�`u"���c��[qyB�'r�)�3?�׸iZ��;�l�8��A��-<$�:#"(���C���?��<�Nb*���B�W����'D�7�������?I�鈴�M��O瓳�I?i�vÛ�k�0�`�`)�d):�#>�Iߟ,�'?�>�z+�(����(*b�!��P��M�&c�Z���O�b6=�Y�Ӯ�%_*���F�: �6����O���i��ק�OS:��t�i/�d&�`h�F*��У%��&��g�d���Z��=�'�?�$����K>HZ���G�<�(O��OTPm q`b�(s5@�T��شi1�(*7��r�+���ğ��I�<��OZ���ʃ�=���&ѫa+�A"��8�II|�0�T�"�S�I}B�˟�N��v��DI	lS��r��py]���)��<�D�+s`!0D'<��	1���<�P�iz���OB�mF��|R0��	����*������I��<���?!���!�4��e>qZ��^�Ȩ�)C,F�*Hp X n���!��|�(Oⓟ��r�A1��L�!
 <�����t�ڴ
&l�<Q��TDQ�!`�)����.i�0)*���k�~��?����yқ�t�'�2��
4�*�b�h�9V�X��1I�-zHn@�R(����OJ|�Cb��O@�[L��Y� ��W5p�T�_�]��P���Q�P�'��	b��McEE��<!EE��(�&� aۤ��V�<�F�i��O�9O�D�Ob�DN�Z�ٰ�:2����`H�*C8����gӺ�I�q]������џ��i�*G:��1n ���.ۛ4t�l)��<�����?A+O��S�O��t��26��eࢥ�y%~i��y�fbӺtJ0��tI�4��48�D�V$W�=�Ղθ3�y'��I��X�	ߟ�����i�<Y���?���<J@��)������!�*���hO�<��-����f��/�4l���1;�1̓�� R�6ܬ��'w�S�Uz���m� t��a
�4{�<�o����$���<�N|���Eab��V�X�K��!b������A�L *@K�{~��'����0wB�'X�u{�K�J��K�g�e?�0���'�r�'l����O8��M��c���U��F�l��)ɶD�80ś)O\nw�h��ɚ�M�O�7M��%�W`�vl�� �!Y�J��s���'c��I��x¤�8��4l�byjZ�2����
7*��#P��y2Q�4��۟���џ �	֟��OG:�@3Qp�������g{� 8�RC�O����O�����Nئ�!:����4.��A�~�	���M���۴w��0�� ~#�ir�5OZi���7@�t��HO%h���5O�xc�J��?���8��<1��?�t.�s?���G �
}���2thM��?1��?����^ަ�CC��0�I��$ar��y	]І`5{5��*�R��3�����M���i��O��p��[*P�R���P�p[�0bT����E��8i4h�g��G��h���H@�BP&ੂ��J�٘-�'DП��I��$�	�E��'��-�T���COh8Q��/^ �� �'��7��H&�D�O`lo�`�Ӽ�'�c� S���
��A�Ȍj?	��M� �if�x+�O6��$�!C�4z�'k�m��ǂ�䮝��8�e�g�4�İ<9��DͰr�b��R��=JM�����r����M�΢���O��?��V`Ң2f�Hå`S���iю
��D�O&6MK�)�ɂ��ν�+�%X"H&��*@x�P"�`����ʓ����s��OxxZ����<��OٱH��u�`.ZB,��Aք���d�Of���O�ɴ<)��i8i�w�'RXb��4�:�rM3�h���'v�7-2�����$�On7MK⦥鵀^�KJ���,b��t��&�R�o��<�W�s�P�������J��
_w���� �Kd�I�n�FԩRDĀ*����<O��$�O*��Ov���O,�?u�'�G�.��u;1�Fs�ԫcf�ǟ��I��d��4
����O$6m�O*�t%�����?��{#��!o#<I g�|b�i�N6�������wӺ牷�$�+q�T'2c�����9�����ې:���'��E�IH}`�<���?���?y���?%�D4�T�ٹJ&&+����?����d^ӦaR��\y��'���W3�dل�I�Eɖ�B3��>/��Z��	�McúiQ0O�	��rb�"�T'�0�(p�3��!k �*r�S}���J(�O�Q����d�.5Z�<#��݉@�p���%ʢ�D�O����O0��I�<�¿i�(�ҍR):�D�����N1�0�U�-���'�M����!�	��M�`H�,}s���C�ӼP
�!���+$��6n�b�k�JgӘ��ݟԃ�� ���NIy�OE
Gń��H�H����Z=�y"\���؟8�I���������OL(J�Ԙ�}	�3�ȥB�� ۴pu����?����OKH6=�V�0��e���#�8^ 	d�̦���4)㉧��O�@�#�v6OF���Y��aj�'� �͓q2O�]QH��?	��OB˓���O>��6Y�nU��%%jƽ8H�#\`�d�O ���O�ʓ^����5�B�'�B�L|�jd���+C��s�� P�O�e�'l6��-iH<q'%a�JL8p��{�@�̕�<����h���.O�n!s)O`�)Q��?q���ODI9�� |E����΃�GF��O���OR��O.�}��b.�-	���'"6���5�� H��oțv^�^�2�'66�:�i�)���52f!JA+֢�`�Hb`��B۴-*�FKg�B�ۣ�r�T�	ҡ)��&z�t���ut8X�� �q:V����m�A�	UybX�H�I؟0�I�X�IٟX*oU!Ep�ñ�ըom�E��jy��o��4��O�O^���O���\�D];^��:c��48��!���kgl`�'o�7mۦ��H<�'����Z��X#m�TwHl`��4mK��)�]���@/O�-��nG��?��C�O���$��CX�Mh��'3�Z�g,�>?���?����?ͧ��d��EK�Ç�,��.��o��pugY�W�f}�Fe��Pߴ��'��B����~�DnڄF@����Je#��&t���Ӧ�̓�?�������)܅��D��(��e?����QG�4m�v��.^�$�Oh�D�O����O���6��m�X�Q�!�J�^)3HX���	؟,��>�M�'l����dS��'���`kH�
i���Ҫ*^��4KX��ēeQ���s�@��ɺe��6Mv������ K��Pcx�ȠgÚ4VH�r%�B�Vc�ܟ��'��ܟ`��某��B��Q�3&R�T��̓^�r�o�O\��<��i۬x��'���'	�$2��]3ĭ�4G�;�)\�;�Z��O6��'�R7����Q3L<ͧ�jůA�3���cT[=@xp@`��[�*���Z"�M.O`�iC��?�6M�Oʓ[�,iɒ�^�L���NPt��a���?����?��S�'��$ᦹ&싦Z�}��
5Q����Eˌ���d�'.74�	6��ĖĦa�5Z}�����3Jr��� ��/�M[t�i���ǶiE��O��*�S��Z3&�<9��3g �@!҇[~M�����<I.O�$�O����O ���O�˧5$�����- �2٣" �.<��"�i��x�5�'R�'`��yHf��N�S�ı�4ZPة��F�}K�=l���M��x�O��4�O��T�%�im�3v�
�3��)EnQ@���J�DP+=R�r��	���D�<Q,O����O�1�0�V�7F��ٱI
�O@N�ĉ�O���O����<���inz���'�'��uj�4#�I�U���]����x}rhӲn���)E�]Q`E@�6^1��у](����?�a�V�=����"�$��D���"�0����5&�x���	���L�eK�S0����O���O��d9�'�?��o��k��	��)ni
 1�
��?!�i<ā*�]�0b޴���y'�*		0}�� �X��%��D1�y�js���n���MK���'�M��'���]T\!�S,	~$@�3�G�|ܠ������l���'Q�	^y��'k��'@�'���QĘ�V+��8l(6� �A��ɠ�M��1�?���?�M~�z/��f�6Az���I@�Q��)޴'J���<�4�l�	�J�*qoXV𘸓)L����Y�cY$�$�5�<a�fi� ����?+O�˓zRZ��GLR��G�^4RLc.OB���O
�4�R�X6�V��i��H�)��)���M�G�p��dW���޴�?AO>!�^���ݴX'���h��i+����U� GD?p����WL�P7�p�(�I=�����O9@��'��d�w�U��X9H���aDj(dC�'���' "�'6�'8���B�S�{A��`i���ڷ��O2�d�O��m�.3���l�ݴ��E�ep&CU�����H/3�Z-�a�x��a�>Po��?}����U��?�Qd[!Zt S�S6w����jJ1-���yU"�Oec�����<q��?���?'��v?|La�+�+}9f�*�I��?�����d���������������O��ty�~��A���<�nU��O�(�'�R�i�V�O��O��|��c�k�����&@>��� I�!T�a�O�I����?5��'�&��	Oy�iU"BbL�i��(ѫsg�����'�b�'N���S��j�44������xʠyrf+�09@�Â��?������D�m}�ak��aᵥ@�y�Teb"hA�NS�����֦M0ڴ?W�\ݴ�y��'
���D��?�bP�� :}�oJ�Y���w�)h����A=O���?���?I���?����I��eb\��͂;���BC	�K^h$m���U�����@��б���k2�P1�0 �cJF2e���&lԐf���p��&���?���&W���mZ�<yҀ[A���j�@�Q��T8p��<)d,9���I��䓹���O���Ɨ}�5(D�>2PGJ�!|���O�$�On�CK��M�"�������Y�l�~h��"��h�J��DO�Y��z��I�Mӂ�iA�O(��g�Ch|X1�ˡ�����8O�`c���Lߦ0PE��+����
��7'pQ*_w��d�c�ݡ�?F�xY�Ԉ�ǌ���O6�D�O���5�'�?�E�ݘJ���7[�>T�F_*�?)��i���&[���۴���yw(��
��$�gwx�X��G �y"�`�$�nZ��M�7��!c�XU�'qz�[S��?��^�"�J!C�Ɠ�d�f����H��'��I��	ɟ����x���`	�\���q��])5oK7
]�@�'eH7�ԛ1Z��$�O6��*�9O�1��KF�Ķ�B`F�"ca.��s�BN}�mv��$nZ%��S�'>��B.��sFDa9�G-����dK�u� Z-O�T�����?I��<��<�Q�E:r����'��	��տU��L���?����?!��|�-O��l�;�$��	5T�� 9w�[�Uͦ%�ë	-k��	&�MۉB�>I�i4�7���A3�J�/�x�'T�K
|8�����=E��[��,?A")H�yB@�i��'�+��%x.��ħ�.�0����<����?����?a���?Q��E��C��sI� c��	�łTSR�'�B�i��ts�:��d�ͦ}&���� R�'e��D��%���Iv��ēH��dy���Z�~��6����d ��5}v=)�g[ @��4:��	e�yC�'u�1%���'M2�'mr�'a�Y��'�) �D���>8l�����'cr[�h�ش%� ��?�����i`�����&���M>C<P��OT��'�86mPڦ��H<�O�6�`#j� �r!���<&c�M��oÏ6��h�0
�1
��i>�k3�'�(�'����@�(H�rm2�-� I.~� V�������T�Iޟb>i�'�.7��d�\�j毝�������7Y|����<�ıi��O���'=�&��\��`z�#O�_b�E!���=s"6-�ަq�)�pQ��Sz ��Ї����/O^Mhsa�(3�:�2���<	HD1<ON��?	���?���?Y����*<����X8�$žQ�±o��&/@]�	֟��It�s��s���Kw
 %�*9�.V��,���H����~�J�'�b>͓�Ƞ4G6�	�X�D����5xu�R�'L@�	�_���c�'z.D'�З'�r�'T�x���;:<ӓ�ά8Ѡ({��'Rr�'Z�Y��ڴ%�����?���wr\�� �X�$�AD�Θc��1q����>	��i�67MQQ�<?�`�RC�I�����bᐟ���Ms��*B�n�Ӗr����p���䖄�!��1m�� �G�����	П�����E�T�'�.�%(�&|�}3�,E�+B���'��6-Ր'��d�O^�lm�Ӽ���29> M`G�_�����D�<���i�L7���d/�� ���]�����T)���}������1ĥz��-����d6��S��c�����Ó�X4��A�'+^7�)BH�ʓ�?��T`�OH��'U�k�n�#�G�i�,��?�ٴ>ɧ�zk~d!����&��y���2"m*����C���((O���v���?a��)���<YL�g��l1U$�¬|``�^�?���?���?�'����HE������JH!EG�ȫBl�CjA7'L��P�ݴ��'��C�F,}��Am�:*�@��5, �A:�4��U�PXJg�_�N�H����we��� O~J��0_$� Ԇ��}OH��&��`��̓�?���?q���?Q����O��i�bM��U����'�N��0=�@Z��I��M;w���|��
^�F�|�N%�!���Pt'��Pb��#��O�\m���Mϧ�x]h`(�s~�N�,aȅ!��5���&�Q$JM��2ƮRğlZ��|�^������8�	�c��>O�2D��'A�A�	@IF,	S�\Dyb*n�lXZ�-��&���O8������ L�}pk�B�/]l)0�9O��$�v}b�a�m��<�N|B�'!��#��36�HSr�ſ�4��b���,��}~�O�q�	zK�'=}���<}I��y'�P	�t����'���'�����O����M����sz�[��Z�P��d@��U��!/O�xnZX��V���զ��p.�| ��@�K�N-걁�̔8�M��i�l`�ŠS�����>V,���'�@�(�~��P��N����͋�=I�͓���Ob���O��d�O$���|����^���`g��M: ����$����@�6�'�����'��6=�Xؠm؄Q ��-%<HJ�b�Ŧ�شA����O��$m�&%r�'��pA1Û�"��I�7��uX���'4�I#�-�(P7�|�]�H�I�����?Lx�A�w ]�*����DKϟ��Iҟ���zy��{�J��N�O����OpVńǶ���S8s���(���'�r�eƛf/g�ʍ'�(�d�5^�LXg�O6F�=Qr�|�\�����'�	c��)��<i��&�����?��eL��r���bA�3GV��g�]��?����?����?9����O��'n��D�pz�e?*V��Q��OH�o�MԲĖ'��6�$�iޱ�C�].�t�s��!4P��#s��0ٴnw��Im���b�OzӖ�I�R�&��9��=� ��S��8 ��Qz�j�< ���h7�$�<���?���?I���?���ݠqL��h��	�L �a͝����M{�'P@y��'��nIrG!�D9���Ꮜ��5�B`�i}�|�~�lڹ���|�'��SƄ�"��Y{L��v��Q��EV����Ӈo���dKol.�;�o�O*�]l�����=�܉Ҧ�\�c�n�?q���?����?�'��dǦEǦ����Ϟ3B,I ��L7"��DsB+}���ڴ�?�N>�sV��)ڴ8O���xX���*Bd:��EP�B��y���r֐7Mh���	�2Ò����O��\�'S���w��pSIP�tb��F�|���'�"�'7��'�B�'4�!����=�N̡��2	5�P����O �D�OR1nZ
ZWT�ğ�3�4��+������. ��k�s�=���x"	w�x�mz>��E(��)����MƩ\��(�q�Y��0�Էv�v�D�������O~���O���m���Qp��!j�� �#�Њ%=����O(˓Xm�6L�MR"�'a�X>�H����I���ڒ\�q���#?qbR���ٴ˛� %�?�K�/��S j�1/ӕF:�pRjݺt4a�IT��~}���������e�|�(�V�ވBsIў�ͻQ�ڂ�x��}����"E�/��l(��!&xh�$#	,Vʓ0������a}��dӈ2w�B�`�^���$w��hc����]xܴz�XDr1�i~�Q�`����:A	�	�p�jm2bdˡlh.�c�ex�Ifyr�'9�'�2�'��R>I��*�	U�����5[d�BA��MS��ޕ�?���?�H~Γ/j��w���e*K�-B�5�"g��J�fE
�q�LlmZ����|Z���B���+�M;�'.������*-V�Prl�@��@��'�۲��͟�
T�|�T���Iߟ Q���z�`�ӧź^\Bh�����<����`�	Wy�kv�i��O����OV�h��Ȥ2_" )a=]�u��I5���O�i�'�"7-�ЦQ�O<��X�'ƞ�:3H:��e���P�<��,3��`�K�JR,O���@�?1th�OL�
�,�~Z��wM��:��t�Z�R�'�b�'&����W�D��o��\:%�K����oO�H�Z��K����SN�O��D]ͦA%���i�	:q��Zd�u� �׎>���`t�p�ݴg�V@c��L�����#���Ozh�g����҉�^c�8YѧY2BĊ�P�-G��
�O���?9��?���?��$����օ�|<�h�B䀫Y�X�x(O��m�E^]��P���?]����	�l(&�P��O:.����S6@��5�O�qn
�M��x�O��$�Or.%qVG\�}"�ɷ)�}H4d��[]�!�\���w-��R��a�IWy�8|����/Y�KN��P�g�d%��'���'+�O��	�M�4N��?1��L�X��n��]��[�?AB�iU�O(��'��7mJ���ش>�
����U�B��<�ЄS�2�T��s�Ʀ<[^=�'ab��3F�?�JӜ���w��Jt�	&X�ȅ��\3�+�'�r�'8"�'�r�'��<ـL^�%� QIV�� `�r 2��<a�bě�L�4��4�'\�6m8��
b	��[R�ʳj�}{a�Hc�^�$����4bH��Oe8�{p�Y���d
f~�۶���D���]�qo����S9�?�W�=���<q���?����?��`�!�^19t�8�fŪ���5�?����d����l	؟8�	ߟp�O��`4✸M�b��A"��{�|���OZ�'�x6-��� O<�Oސ�DB |,Z���I��d���>Aq2D����
�i>E��'!*x%��ɑ���$��%��H�����%�ȟ����$�����]:E�)O��m�T�"��
��dLy6��! !J�ʟ�� �M�J>�'/��	�M�Rl\�J�,�:!�x��Mځ�A�@ě��q��0Rc�Z�h���O&=�+G���6i�<W/ƽ�vU�t��,u��б��<i(O��D�Or�$�O����O��'4ޭ��� R�r0&[~�<@�!�i��d�'R�'��y�{���Y�Y<nٛ&E�@ӆ��T��M| oڝ�MSq�x���^�n|JlҚ'��8Ç	�N�F��%*��Pn���'����dK��,���|B[�h�I� "s_@l��p�ځUx��j���<�	ޟ�	Ty��x�pq`cm�<��A^��BF_�[L@c��ݱ IV�)�҉�>�V�i7�6�{��o�ri�GP�X,j&�,�$�O�����`���Ф�<q��r ��C�?�e�]�zP"�.��|!w]��?Q���?����?�����O̵�	 Y� ��cJ�mMιq�B�O�mZ�t�N%�������4�?�L>ͻBR�#���j(��xvN)�u�R؛� eӬ�o�"9��,m��<���e�dt����L�#��.i��|2t�^#}��V�������O���O��d�O0��ܒ`�����P�Npi���#F�W(���?!��?�������?ё��c!�x�]y�� �bۀ.�ɫ�M�C�i"VO���2�I�I��d��n8g\�堓i��-2\I��V�mϾʓ&�R��1�O�=�H>�)O����C�&��Jǉ�+B�c�O��$�O>�$�O�I�<Ie�i��ȃ1�'�L(���6P�B���i@�~��i���'`6M5�	/������� �4G%�fL�� �2\�����s#8�!v��Sh\Y���%��$=��y��'Lʓ���Z�qH����@�}��5SD)�
��d�O��D�On�$�O��d4�S�3�����?wxa��lQ��~��I���I�M�4/����D���$�d�Gk�726 ���ѳt�ڀ)���&�ē7��p��i�R��I���|��K"� \$�b�P7D��Qj]�
dDX""A#�?	C�(���<1��?Y��?��b�
t�6%��(c�r�ZW �+�?�����ЦI)�Ae�7��O���|�p��6X�ȃ�S�x6�s~R��>y�i~�6��V�)�v*�*s�q�@	1l[���Ҭ�m�r��C�D���,O�	C��?Q".;�D˫��#&�ѥn��X:�-(/��d�O^���O���I�<a��iW�����0u�����
dP ��G�x�B�'*j7m!��=����Ϧu���*Z���r��ޕ|4<�@�E��MSu�i&�i������-I[&) ��j�3\�Hk���T�hL��X����D�O��D�O4���Ol��|:��ؓ:�ؽ�u.���%@���hϛ�@�+7���'%"���'�v6=�du���:,�(e���ϼA\��hqA�矨o�%��S�6"snX"�"f��PcE<�z������wNt��sp�	I'rK�b�	Hy�X��{��
hZ��.QZQ q�0O�MmZ�%O2�'������^�B�ـ&]�Kx��+���Tu}b�uӦ�l���m~�9c���:R�,��Q�5byp��'�2y
u�F�B���d��tgƟ���'��Lba�ܱA�0 ���.j�Q{
�'MԬ���M�%�d䡅�ذ�Ux�'IP6�\���ʓH_���4�NPX���x;����3���4On�mZ(�Mkc�i��UKà¢��$�W��P�'Gz�!�c�=ta��Z��̾��$3�>�d�<���?���?���?!A�� @R͋�Nŉ�*{�����D��kP�۟��	ӟh$?��X��Xk��NSR�7�T!A<*,O<�|�&���d]����2$�SȐ!WE"�x�hX�v�x�S#�<�@�#rE���� ����M#`��.O�OD��a�'Ƭ�a|B�f�����OYa��żh!�(�G�'����c7O�oZX���	��Mcŷi��6M�#���p�%L6>���!� T�	�A
�gz��,�D���O���$?���J�ڬ�'֑ ����)B�q���z���xr`6hD�'�P1B���:ų������4S����O'�7m>���;�
�[���Rr0�rBNR19�8%����4yǛ�O2�Xb��Y)�����_�q�5Dޘ0�e &�
�˶L+;L���
�y.�k�J'Z���B�,tr�9���� ���4�?ʑ�����
g`�7D�n�`g(� Q+�/��Nz>��wn�@�l�C�c�;.�|1C��f���i�'�"�q����=���aO�3x,|	7oRU_$����� ׃�l���5�Q�3����p;j	P�)�mWA,�j�$#&�4J`)߮lJ�F��L>Jს�O�>�=�5'��[u�i+$"9�Ԕ��,Ը@G��X�D��X�-��ӆC�(E��B�1�L �IԠ@����gH܉V��R���h�F1�4�?1��?��'Z�p)5BJ�!Z����� ���I�x2�' BiA?���'�"�'J�i�3Dƾ0�Uǣ&:�@'�M�c����'���U=��'���?u�	��X4<a��Ӏ"X�\q��! J�7�O��T�vӆ!����	�%)�t� ���$d�Zr`A�x֛Ve����'N2�'e�T]�(�Oai�A��+��;��_�2����Bv��ić&x1O>��	56`�#$���cc��2/�#9��m�ܴ�?�-O|��/�<�-O��$���c�Џ@J�9��&X;fkt �٘'��Eل�0��OF���O��f#&}^%��C��Zjl��Bݦm��'NA|����P�����5�&V�"a�-F��F(2�ұ�'i�`1��(����O����O���O�5{��7%*4���f�uR�=����\m$�d�O>���O��D0���O����O2<��	Y�r[V<ȃf��6~�����Gb�	�X�I�$��ʟ���AOG��X�HJ�i��J<���MO�����韈��c��韌�	�"t��a{���c�ƙ$6l][��2Y>Fp!_���Iğ��Hy.דk����ٱ.�U�pQc!�-F:������Ij�Iٟ���
:Ӹc���a|�I ��6.����K}�x�$�O˓	Q˰P?��˟,�S4�Z�� ��V8����@@*q��Y@O<���?Q�+h���l�IE���	!֬�V����t�a¦}�'/��G�{��d�O����tק5F!��hVP  �Ο}����5���M;��?�#�t�'|q��XB�6Nc�M[fO#	}2t�g�i�D�Ȗl�����O��d����'�"zb����	89`�um��.r���i~�2��,�S����#����I�7�͙M�ܑ����M��?1�����G]�L�'���O� y�F����i̗s^��a�.sB֒O��D�O���<7�t��*�3;�%�ͥ �Eo�۟�B1���<�����W@̪C.,�:1#)9|��S`x}� �� ��'R"�'��T��kBN�F��lx%S"U�*pHG�Nl�fQq�O��?�+O���O"���6{p	����\Y����̵�!��O��$�O� <�r�6��1�Ȋ�.7���$T>E�X0m�TyB�'��'�R�'�����O�eCdD0��<��[/1掑��R���I�����MyB)�Gݘ�'�?C$�!	"�Q0���=>:��r-��[ �6�'e�'�"�'��h���DS�H�4���S�(]�,w8���'bZ����@��I�O����b�{��e۔����Dk����M���X�	���?��Oȶ��O�,� �q��F�H!�S�4��"t6�Hn����˟T�Ӫ����� ��@4/,(*I��eS0;��t`�i��'�`�d;�=J�tlx��?��DA�
w*|6- 7��um����ʟd���$�<��#��#s�m�#�@;����D� 	5��I^��O��?A�ɖ9�ؑK�_�hZR�Ё�.nG԰�4�?A��?�"�������'�䁟 �<Q�e�:)��i�x���'��	,W�xC���D�O��O �q(��Do	3�|<�BC����I�l�zN<�'�?	�����Cъ|ұoڤ"�1��C�,���oџ� �������'G��'��S��U*�"���B��'[֐q@,��7 a�H<���?����$�Ot�dI2r�f��!�Y�V���`B-�*�:�3��O���?����?/Oc���'e���a ��R(��NWvW�M�'���'��'��I�0����}�j�W��'!�QSTM��P�L<1����D�O�L0@��|���G��8���M��m92�orњE�i��Od�d�<��Gp�	d}v)���8���⩀"}�6��On˓�?i��O2��	�O���k�I�[�Jt�@ͯ2˲,P���9�'d��'<�b�d�6������y� �A "�a�8}���
/�ILص�S����I��(���?Q��u�dօ��`c5H�<V˔�S���4�M����?��I�	�H��<�~R�
Yk~���!��lNP Y7�ަa�������̟��	�?i���)Y<�Z��1�R%�D���CQ^�(oںBC"�Q�M"�)�'�?��O�6{Y�@��@��8C�!N�J��F�'�r�'�N����1�4����Ojeٕd�i�$����/̐A�Gd ˦���ğ<�	�v~�`����OL���O$�@�Qh�`����P�Dڞ=�6ʌʦ1�	�j�T��N<�'�?aK>��4�8!谁��E�ȵ��ჵl��'垁S��'4�I�\����Ԕ'<lZ��V3J����U�� ��5)>O$�$�OV�D�<���?!f��&<̩���٫$nQ��&F`������$�OR���O4ʓU�\d"36��X�GS5�H%[b%]0Y�@�� T�����&���'Y�AR�'���TDTVhUP5�=zr�i��>���?�����Ğ�C�VQ$>��'$3f���C�@p�	��M����?�+O����O��g`�Oz�'nHmH1ɗ NEP�qb��"_�4�Q�ig]���I:m�4��OT�'y�\c��;�*Ȣu�؈*1$B�M:�pK<��?��ȭ����<�O�.����fp所���S���ݴ��d�D!�Ql���i�O��	�E~BI	�a������'<�u����M�/O�qQ�,�O��&>}&?7M
�y�U��'ӻ�>�[Rm�'����*-�6��O����Oz���^�i>�˳Q�	قѱ�"�nD��P���M[�	O%�?������+�9O����N�p
���fV��B�L�62~�m���I��h"g�����|����~+j8�p`�A�Ze�h��	^��M����򄋝{���$�<Y���?����5>���A�-Hyh�SDNƦ	�I:j�0ȨM<ͧ�?�I>	����`'�Y�%�H�2��d�#.K{ �I�� -�IWy��'���'\�I�s<�P��ӳY�����"J�b�D��7�������<)����O����OZ�� T�.�`	��2O���
�Ń��O��զ5�I�Ж'��x�b/k>m��Ǧ)�1H��C*#�R��Nh����?Q/O���Ov����6��ޏ��1��3�L�@��ʮ	�9oZ۟���ݟ��Iwy�K &{�F��?�1V)X�8Tc�ܶQpt"Z)6�DoZӟ �'�2�'L2,۔�yB�>���(<�RC��h�x�9�����IΟ��'���`�~*���?���z����l�vH�CōG*?GPd��S���I���I�sĢ�IO��'7�IG�r���� F� ����u!*:�F^�$r����M���?�����wS�֝9����ʤf^��Ѝ�ER6�O��$� /�$�O˓��O8z�z�)^9� �z�-�� ��p�4��C�i���'$��O����$ӫhh
t�@#Ŷ37mq�Eάr�(in�*t�������I͟�j��#]x%�����(Xx���gl����i���'�U�q�:ꓨ���O*�	#bB
�	U0�`�å�}��7��O��?����S���'?�'C
� �`�[�l����*l�
E���b����a�@��' �Iݟ̖'Zc�Z'v�b��/�&(ݢ�O�m:V4O8���Oz���O����<����LkPH(f?-/x	p֍ˍs� �
�V�H�'�"W�L����ɰ D����GĮ'J���p��v�|pu�{���'���'8�[�h�����; f�	z�����^lBw�]��M#/O���<)���?���F��'���R���ta\1p�.�s��%��O����O���<Q�+r������b�NvZ�ty��4L\<���C��M������O��$�O�j�?	�NTtl�E%ԝ�%��?�J�m�ڟP��zyª�*Ұ��?���R��̪Y(x��/޳s�V����Pj��Iȟ���ϟ��C~���	yyrݟ2��D��I�ز ���nBN�T�i���'![D$ڴ�?A��?y��xB�i��R�l�1Wؚ�ې�4e�8�e�rӖ�$�O�Hrd;OY��y��)8bv�I�0
M4u���oP���I�@7M�Ox�d�O:�i�h}B[����	��(��Jٌi��}Cw�)�M[����<�����d.��� � ��1Xwv��Dء/J�Ej��X��M���?1��0�f+�\���' b�O� &�����oVb�KNBB��#�i9��'�"�ٱ�yʟ����Oz�$��eڪ@{��H�H�u��DZ��o՟�������D�<1����d�Ok�$Nh��c./j��$�֋Q�GC�	0b��	uy��'���'��	�~�6,���Ē&0���M�(a �J�M����?1��䓈?9�}W>U��$J�*: �Xw�?O&��3&�<�*O6���Ol��<q5+�>󉇸x�r<b#���r���G�9d��Iڟ�Iz�	ڟ��+�8%���j�&�S�@�x���X���Snhc�O���O�d�<�E��kȉO�ĸF��q\ 0�@ʛ
M�պ��v����)���O�����"�'O�<����A�	0����CR�nZ����	Wy©��I#v���������7
�L��L�cD�)~���Xk��ğ����I޴���X�Ip&��I�.p�B��)|��Ȳ�Qަ��'id��G�`Ӽ��O��O��	�]��,�h�Bs�J 9�H4l��`�	8@]�II�Imܧ]�24��� z)l)X�P5E���o�7=Wxܴ�?9���?��'��O<4�c�K�`2d����~j�(��F��9���Ɵ�$�t����-�H_X%i��[� E��c��{��V�'R�'ע�K� 3��Ol�ģ�#�Kެ=B�����_���"�p�r�O�q�6O�ן��	۟����"{ �`���*2fT��6+��M[�Q�@ؚr�d�O��Ok˘i/���&�J�EС�TL����P�r���eyR�'d��4Cp.v�U*{ZL�VeW�(������"����d&�P�����1��NN>�x��U3X�\A�h����Ny�'R�';�ɿ#�����O
���nX�F�V�� C�2j� 9K<i�����?a��U��mH���C��@	r@��m��/H2�d�>���?���ɳo��$>%a�I^T�P�ʅ_�V�	0/�.�M�����?��f������I\#���M� x]*�ۢ��0 �6��O����<��eĉOhb��5�� C�@CcX�?E"�@b�'��'.2��n��|��J={�BQ�xI��KG�  ��� �i��	%e�P�޴Z!���������	)?�� 0���!d|�R�@�\�I��\��������_y��4D���F�����7���$NI��M�q�ň(t��'r��'����>�+O�`g�ԫS�B��쉝&�����i٦��3?�+OJ�?�ΧW����� ��&J���ٴ�?���?1�o_�m5��~yr�'����	���(�J7�dMh`�нy3��|b^�yʟ����O��d�#N�Ԩ*�I	��Wg���($�ik��\7B"���d�O��?�1dօs��%$V����|�o�ӟ��`�X�I��H�	ڟ��ey�%����(fF�:��#"-츍:���>�)O�$�<����?a��[\��3Ğ�ge8m�@�B[z� ��,��<i��?a���?a���ĄAx(ϧ+�h �P�1_�>�� C D*tl�Oy��'�ϟ�����|9'�`�� 0@�=Bd����i�02������M����?A��?)+Oղ�LEB���'�)kF,'D@�آ"�� b[L�Z�/e�J�d�<���?!�pB�!̓�?��'�$��mC�}��y��@����4�?�����dͮ^�\�O��'��d��ֺ�S7�J�.�����$;����?����?��o�<Y���?�����b���N!�b�܊;�Z9��	��M����?�#NO+�?��?a���+Ok�K-m���Tn��i
Jӛ��'��O;T=İz�y����a1�mҥH�5*4]SU�$�M��M?(��V�'��'���I�>�.� #��8�F��r�)}摲֤�צ�SW �M���I>���)8�8�@��6j1���Di%�\��iR]�����R�L�Iuy�'���f`�BrDE�l�����e��$��<�iI&[�O�r�'�2�L<O8��stc�H������y�z7��O��+	\�IΟ��I؟ ��5�˱*���(�3���󁆃���	�1O���O��O^��,1�Pݚ4�_,���$L �=ΐѡ�L�<+OR�D5�d�OP�Dҍ��uy$m[�GSt�(O4C4�A ͆(8-�IџT�Iޟh�'��X"�o>5����5{Pɒ�1n�\��Dn�����O*���O���ĭTU?A�#Cz���A,E�V���BM}B�'XB�'�'���ȥP>E�	�G]�̙#�0�df��5hz<	Z�4�?�N>���?I6��_=�&���#��uKF�w�AM<@��odӜ��O,���OJ����|���?��'I��\��Jٛ
Db�$�H'i���t�x2�'�����g�Ԁ�y��@��h��:�*D� ����i��I�mނ���4�?���?��'6��i���nA�'-@4�W�Ǿҵ0T'<�!t7�X�SE����j��頥��R�I���ܚ"כ�h��b�'�r�'���^�T�O�L�`��.�Ȉ� g�Q���@�wӤ�Y��Ǧ.�1OQ>	;���//� ԒDn٧~�t�it� %O�{r�̰s�p���mZq����g������`��:�F-�$,�nQ��s�1�O&�b��=o$IH��ѯT�Έ$+Ҡ^��x6ǐ�n�DM*$j��[�Z�Z f��}GT��g�֡H��(Y�)תvȹ��Bw�@��v��*�!	>yn��е	1kDP��"_�X+� cve��H_ȠӇ��j3�%jE#4mZ�t�G�R&D�b�[4G�v��e�R� �"���'5��'�� j�R�'��阕Ƹ����3� ��+Ʀ�e�F[��7t myf�'Rl�EQvI���Oʓ�F(s��
���5Xaꇋ۪z��AZ�� bȄ�Xg&N�bۤ}�'�����?��S'7n)�&K�g �*���hO�?Y�熆y�R}�ժ�;"j!� i�<�E��a�0� ���uU
���<�QQ�ȗ'�p�0���>	����ɍ�m�(��pƘ8ZլЪJpj�3!��O����O�Ty��#$��������T>qIgMY%SyRY�Ĥ��B~�C�)�<�r�0�K�>`Y�ݫ���UGu�q˴�*�"q$	�,V4Q��zEc�O���(���%S���MZ�{�JM��JdO��Im��l9r��,zN��[� �J�t�'%�OR�'���w�Ѳ(��J'���~|�&�w�8�1˄�����O�''(A���?I��qp��⫝�A4�� ��P��a��
��yhWF��;`�qV���I0��O�{�W4$2�E��/J,�ֆ�%p���2!�ݸ�H�g	��"~�I�k	�,�5k��M�����C��?��e����ڟ��	F~J~JI>��J���L����`��H�K\r�<!Ō�Q�lKB	sI A�PHSE�'��"=�OϠ��g�cҜ�X~y��']2�^$A&�W�'���'c�+�~���Cl%��R"I ��1V��,+B�iUj�sw���~Ph�*�D����D�:O�t}À�҂G�V��Ƚ6�}�ɦ<��7��J^^Hjٟў�� �+���x�IΠ.���kv$�h�2hƟ�����M�gy2�O��Ƀ-i��.��$��-�2e�B�I@�~��'G�� ��Py6�A�l��ݴ9�V�|ʟ�ʓm�ԩ�ir��f�JF��zb��>댔 ��'y��'6�G�4`qB�'r���%{
����K�TM!'��v1CR/� fx@PEkُFL^��ܞTX��Ql��V�JE���]%3f�=Q�I�J;u�čY	HP���J��y�n]�CހnT#1�K/8�R���O��d�<����'�ԉ�����B���LaC�ڱj4���b�>��I��[�E녅b�� ����4VELX�*��	, �X�	W��)I�4�?�����I� =�i�����m^E;� ��}Y�@h�!�O����O �T� qz�9�v@G<&T�r��|R�%�)OE�@y�'�.:X/�J�'�\q��0_ �P4�%a���OzޑQ��7E��B�,L]��Q���~���_>Z)��B�2�T��GeQ*,TB��_�jtQC�	�[�k'O)���d�D�JA��V�Bx�����2���
A��#ش�?���򩀥GR��D�O��D�<[��Z ��uez�aӤ��^Ք!�pc �!��Qw��!2�|*���qB���1G�
=":Ē��[\��W`Ų)s8-Xp�O�}NN%ɆOܔ͈��ٺw����X5(����ӏ���{��'�1O?��]=s�������	u�(!b�U�T�!�$.,���)X��C�'ON�4���?�bhÍ8{&�h$J˘e�T�8`�����	 k���E͟���՟@���u��yWCs�:��pfJb�h�iص�~��A���>yc�_�b�˷��=~.�'`?��Rgx���U��j����Eo_�aR`�iD��H[�/�O.�����7�U�.u��,�֬�%'Q!���(tT�U._.=hd{B-ԭ~DҠFz��)�4D<Yo�"���1�n��e�`Ы�F�?Wl��Iϟ0�	���kʆ���	�|������I��� ���<�TX��O �2�P����$7��ɠ9�:R��O���'Z�$}���� �h���'9�}k�"�X�a�:	n�
�'7�[P��-�v��
�}:؄x
�'*��hR�F�`��ꔢ� u8���'��7-,��ND-m�ڟ���X�TU:m�)3ah�u�D�S�	&=vy�v�'��'�����'1O� t�@�
��œU���"�Mm��<��Y�O�ތiU"Նqm�M:�d��'����k���S<��k��:�\�:c�$�B䉉k.���#k	YS��C��R��$Ee�;6,����~4�Ȼ�-��Y�T�Iz�����4�?�����ӻaj���O���ڂZ�^��2f��$a����Ȃ�2�1іjɛ9"�&��'���?�b˗L�(<q�P�g֪ED���oh��W�N�Gv�9t+�t�P�G���1�Btk$B=0C�d��_��t�D��?��y���'J�HL��$d�Ԅq.�\�'�(�E ��[^�0D�m�tm��y��''�"=�'�?I�ᓒ����nS6��I�����?�y�u`4G�4�?���?�2`���O�n�M�΄c�"Y����NV�[z����!B����:����"ӟў� ��#'�
z��t�Gmʤ]�t8��+Dȟ���HA�O�x�۴J�+2��퉢WG���@C��+� ���K��^��I���D)|O(E�a�ȯrh�}�l�"���[O�����	Qv�b@��N��<qv��95eEz�O��'�r���d�N$!�/Z�&;�E�ҋX�9a<Xd��O�d�O���^�;Z��O�$���O��h��F5�DK��^�Y0��T�'j���/On��d�{��d�"�F�Nk�="F�'�2�Q���?��J�G�٠�ʌ)s���ӁRv�<Q�w�<J�U#��s�����'���P%�%\�����݋'���͓
��O�%�W��˦���۟P�O���T��?V}��A��c�U�[�O��'�-��hub��&`�1�Ǒߦ�'Vrd�	��F���C	�&9�Ey�F�	`$�R����t�0)P /5����.���@�l�<0�*�@`B�9�(Ov��T�'�����'��IJ%�z��2����.��d�'
�O?�ɧL@8�'�^�_�ʥ5BF�2������W��\��]+q��P�{Biגl��R��DHش�?�����H�S����O�� �og�=R�<��U��kʏ"(@Q���:,gh@S�5?�OG1��KW�n���'fDu���D�K��A�u'Ӕm�)�g��~�fx���'sl(��,H",Db͆B`~�0�ƒ8���q��l�؟�E���p�D�JEM��g���k�,5����?9��ly��D�4����ZB�Ex��7�PB��ɘ<�uIw��9�0�Q1ǃ" �V|��ğla��\�d�<�I�����ҟ�Y�����!��{��I���v�Y S�D�+6��L2��'l�y��\~1��*{6P���'��h���H���=1vh��{���۴�֚?;Q�wړ�?����=�?����?�gyr�'r�B�Nͫ���2c����I�4|�C�I�\�@zc"W>��� 5$V�Zkn1��|r,O��"�O�UF��1XU L����V�v#�O��D�O��d�$7���O���� e���@��R(������J�hTٰ�P"T���5�O���$.� Az��K�$;\�)�BRs��p[���?h�bqE)<O�x[u�'e2g��bHY�����3�v�R�
 �"O����O���'_�����!�t���Y�*��<�
�/�Y�(Z5BH<�)�h��ϓr��nh�jʓI�^a(��?)����)�
���a3��x�X�l�1,�J���O0���O�R̸t�xM$�L�O<��w
Z�*&a��^Xy���	[T|V,�&;�y%A��in��'hk������	C�N,xzTDy��G��?�3�i�87�O|ʧA1��
� �X�q(D�x۪����������D��;��ѵ�I�3��`�[��ibe�)�/�M���i����q^ T`��dh&a+�K�&�y��ջA?�6-�O.�D�|z
J��?����?��iU1����c� +^��M�͇�Vٔ���lѷ�����/�I�SάȄgN�Uj��WL%J:�	f�x8��<E����IZ���G�ڑ؆� L3*�#靤�?����?�����B��gm�!`.�A�^���!��yB�'��}���0h����Ub�	h�`�b����O��Gz�R>�z��%f���K%B)bp*����,���_�����-��T������	��u��'��K_�j��(bh:a���AsA�)@�8oZ�'5�FH�I\B�9���?�=irƕz%|���͗?>��`� (A�6�lA�4i�&�*�D���	!eڪ���,�n������26�d�	�e.���O��O(�$/�iP$~������< ��e�#��N�!�$QF�8#C���X��H:e'Z	���Gzʟ*˓kΪ}rD�is�8�� �z��-[@*O4�z&�'B�'���՝ayb�'��ɇ��'+lc ��{�B���@ܬR �2�R��ؔ'�Ɓ!�CԢf�$����*?^9��=�����,��aeTȤH_�PJ�,�4o&D�xj�mɘ_W��
�/'6�b�%D�l�F.ی�B��	�h)p6ln�0��}BKS�e��듚?�(�Y�@%HDyf([D.?�JU"��P�tT����OP����#(��*Dg�T0��**���M�O%��E!09���uKH�B k���˩J&L���4]>i�t�I��Q9��#�j�#�0��g5,HQ�Lۂd�O0��.�Ӟ�4���XkL�8��b�re&��ݟ���ɷ=q���0X�JT�,�<����]�I74q�a@� �Lr��E��$� nB�(ȨOT�ĳ|ңF���?a���?��e��RNPY��i%@�".��b���y���i��?y�|��/{~�t`Ѯ
<�!�7������2�!���0cPK���b鐵L�>�� �i���ҠZ�h{B�X�|,���[7lb���O~�S�Su�ɸ��� ŕ�gP.A��<\�C�I�.R�ҡ-^6��a86�e\L#<W�)���D/G��Ĳp"�*o �"G���?���6�З(g�$��ڟ��IߟLq[wEr�'���&�;:�����&�11����'j�2@��\K0�'��T� '�J��B�Ux�8$��)���y!��ǫB�"<�/ߞt����>��qQ�E�uD7/S�Y7Z1��+K����cq�6`f��Y�$��JyR)�]I��Q��0��1�ǒ���'�ўb>�w��m��i��c��-l���B���Mc��i��'��Gy����7��.�����K�+=@:��@�F@�$�O.���O4�Jf4�8��~>��f�1S4��D �|��Y�_�A���"Q7>��|�	� �&�;�\�hZ�� g���(�J��PL��Q���DO�9� *S�cvD��q��a��MH4�#�M�����OP�����i�N�V��D�CQ�6*���m�@�K':��h��H�tr<Γg�	Vy�d�b�4��?Q.����G
�8�t����D؀�\9|~����O���ό%��HD��-Yd��p�с�~�aLэ��S1��72y�� �R�'�����8�^�*B%�?Pm	�]?���t���P%�Q����e�)ʓXŜ��	�����%,F�J�@A f�(�e�u ��<����>�e�Im|j�i���2�z5K��UG�l�I<�d)9���¦��6	+r	FE�'�y��+�a�G�o����A�y�/ϩ�huR�� ����S��y�:"PX�[f��H|���y�P��*��JoF�Z�$��y�"�� cPMD�b� �	��yB���Cq�q1 D��Y��2Ǫ�7�yBO߂2q�����O,%�*|H�K��y"P)~\$�2Cm�2m|Bf�y��ܷ8��|�l�e0(@���Q��y��1��6k�9Z6t@ՀC��y��Vi2���� R�BQ��ׯ�yȋ9z�eiY�B�Vp�
�yr)E-SL���&���J��y�St�\8%D
�	��p��)�?�y�"M'u�fm�FfS?���Q�>�y��I�1a<r3ᒖ~Hk�M^��y2.�2j�	d#[�w�č��#�y���y�R�bTDL*k'�t����ybD�,U܉%�Ne�RY@�"���yB��<�  ��	�kR�؂���y"E�!@`z`h��R���C�j%�y�d����4i�� #��ybFT2^*��06T,jd���g_?�y��ì/ R����NnxH�(� �yrbT28Hr�TEX=x�${�o��y2�[?Z?��`�jd8�b#��4�yR�/̴�
�J��V RH�b-���yBȗ'Uʀ��� ��a<�X��Q���<��(����'�Xʰ�����x�Վ�)%nLPx���ٛi2#~:��I���X��P���E�O�Ɂ��������G�]2���d��	tq�̋Ղ�8���CV8?�u�=E��4xX�s <Qx��(�V�� �{@�hc?�O�Y��G�\��m*DAQ&�P��>(^�φ�dP�+1X���Op��C��N���C^�(9ȌZ��X�Y�4�X�{b��?�8������>�wTQ�-�s 81x�� ��8�@1H*�i���F�k��ɏ+�~2F%߄a�C���Pqj7�ÏF�@����y"^�_��'�h���1
�0��i�gG��P����^�ɮd���1��/}��?ug�B�YUBh�b��;]f��W@J�0�(��I>�SH�~�J�7;��84�����G�e� ���kƅ���aZ>l�|�[2}�Ӕ<X���)�$V��8z��չ1ii��`��y��v�ݚ0�OV�d�3�d�1�Q��&D�=�N���Ȃ��_�~l@�!}�9�{��;�O�#�NC&M{�����P�Zك�Dri4eЈ�DӾ7� ���v�0�;x�=��D�*H���+7	�#���=���;�Ӻ�v�G3!��)y� �Y��(�<u;��j�(�1b�|Q�xҤA#����� �Kv䛣f�0��'9���7B�4L Cǚz�E���dJ�����*4M"Gϊ2:���'w@�+�
�	^t�:SJМ#��tԘb)Мr�M��s%��D�)~v�噶E�.����������۴|S�)��-�<B�8y�ˆ�|Fy�Ǟ�Mf�a�мg�p��ؽ3��䉤s��"r'�,�yB��.	xP�UiBf����Ѫ<)�J㖈e�'jT��� 6t�hGzޥ;3*�o2`����F�hrE+�<�I�A9���W&-�<97"Do����.�y�|�`��H.P��O0�R�*� �|�%��3��R'�DZ3"���1�j��FV�,��k޶(d�4!6�z�T̳��Z��|̕'���2f�vi���͈� �:�k�)\�n㶽b�nQ+(_�9��	3:�}�#i��~-`�x����Ԗ7M��<�ԧ�P/�����&~���c�W�&O8倲M�Y~b�8q	C!|�l�*v�B,h[����}�2�>aujʑ(X���)D�r�P��'���M+O�e�#����D��'il8��M�6w��`��XM��,=�DП(ь{*�k, s�hz�E�0Ҕj�j O�ON-�aIB ��%Z��˃�D���!��_�n[J9�"��V6f]8�[<�?��$�~*�@���Zؚq���~� �� �Q���.?��=��J�0B�K2�=�d��J���lQ���x~��A������~-|a�s��?@�'�L����|�0b��~�'p�5dZ*�p9P�#�)pwJA�OP�˶�PT�cy�#�D��+�O�!�W�A���x+�M'=�
�I��"?�������� �}�@E*�����D�r� a�uˇ-�MK�|"��O��=��5��!�Bp�-,(��a*u@\���$K����{��?)qHL�?�]�b�#I��-���Xi�|8!�ݧ|��*�I^��L�:W�`�[�锬6�dѫ����ϩZ?>��@ |�1O>��Hp�0,x��½��ԟ�Ā/��cr�I{����Q
�"��h�O�u�s��/[%�"6Ɛ�(O�M�N�"�CeBa5F��b	�<Y��'B	q�&�'���Y��Rk�O�Q�'�le���ǥ-l���&I�~.�	�F�i||]Dy��F�l���.9��ҏC�4t�Q"��&`$��&K�ASW�I�_�Y�u�|��O��.A<���G@�G�` ��>cS��`������=F�ӧ��O����K\I�D�,J���TDT�}&jȳ��?��¦]즩�5�E}(��N|�O��j�d��Yi���DntsW�Z����=@	4���'�� j�Ɖ�F��������ɑ, d���/ƍY� -��eʴ��B�fK�npbݚ� ��K�џ@0�ٝ|�P�0Q�44�<��ƒ�A}~���'@��s��t����L�A��9 �0�d@��y'�G�R.%F�K }���wÐ�B���*R�Ӆ$C�q�牺]rn�W@�ﺋ�ٕ6%���K�P��ʻ8 �\kWB	^��pę��)B�njo�)2Іp��E� q�nn��dYAz`R@g0'ha�r��	rP�Ϙ'�6$�u�I*i�]��灚ex�aN>���?a2aS2�������u:ģ��l���N rq��i��vx��Uc�6I�L�� (�OֹiS�7�)��w�2�A9O
��{f�h*���#[���ʟw���B,���=�Oƾ��t �1,�X���!^��TI��� �j����P8$��0��"i��)T��.:q�/4c�(�r�8�|�W�\�.u��O�y�Hm/@5أGM�Y����íT�T#����'rĄ�U�ι=�ZU
͟��>*-*�X��jļ��e%��������x������ӥ�J�}N�q�3�*D���<ɳ�.L���
N�1�h�s�����` ��%���YC��t�	�e&��[G��}w�DC�(F���I�Z:�8� �̰�
�=�@���^�c�`c�4�!�_�g�p�� �o���7����B+_�]��P��&9���I?j4�؁��?��qt�Ƞwk��ʧ>������ h�@й i#]JX�ȟ'�-����6�%����0|*q ,�J�q�͙�7�IٕJG�R�P ¶�4�|�爋Y�p��#���yb�؟X���Qe�8�|�ZF�� ޚ�ɝ']�]����a,H-Rȟ��V$(�R�_��z����8EB�ؓ�g�T�ϓ�J�Q �)�6@c�FU�^z��<!DFT�Zj�9�oݗ`e���f�TC��F���]I��C�I�Wq�\K����8cGP$�n�	�8Lx�"��v��#E�(�qD<f�@�f�E>b�P0��C��5Bd�!�?a�u�9k�a�D*J0,P��b�O ����A?F�4�� �k�f`�q�T>��n��g�8�؄h͌	n�u�ń��<9ւ­	 ���d�Kĸy��S�;��(V,Ս�65���0<d���ީ"EqO�S�[�(lh�%�!�,-�M=���l:rd,�y���SŰ��n�ƀa���#5�����̱ZWθj�W5&.12TJ
�`qۂ�U�r�	%�qS�m\TY�)WB�.b�t)V7.>A�s%�I ���rO�u��Iu�
�z�"�Ӏ�=���:_"�ф�M>nwD�#Toȼ��Ѓ5:�@b��v*	���0_� <Z�+41�1O'+65�6x*'��+Y���v�R�Y��{N�ݢJ�	���$�E<�Y��l�Za�%����6,qO�S�R&��q�=#���ED��iV8�����s�Ϟ�TL���慂y>��U�C?l�تSmP�Sh1��˘�>��b�T>�Q�ʀ'�5"fh��<	cn��X�0e�Ƥ�<x�92�U�4�F�͓kDj��G��!g�L����Ā�4&҄3��\�}���jSLTs?�$���X��才vED�2��Z�;�켃�Z�=&�b��Ñ�[�9.�� ���e*��>щrk�<:s ��vK�Y���a�|rC�9.���e��h7ɡ7��~��Y�r�\�b		�L@� ��8Z��*��U��'�k�T�M �(7�8U��"'�,1�b�qCN����Ij�R�w&=wdT�+T(��xՀ�ʧ`�(�jg$߲~6z�a3��i�H�'b���2k�������|jc,ϒ��i�	G���<s�e	���8H��rt
(��a5�M�`kqO�S!1��)k��Z�8��}S��:��Uu2���$�-q(���'�g�,�IUr��	1����3�sђ���D?!k���!�MD��0ϓ<`J����Y��EB�F3Q��$����D�(�y�Ϗ��~YQu-�*17`drЧ[-��q�`ep�Wz�	��5W���~]j��4p�,x2�蚚m��!0��K�,H�Œ���O.Y� ��5��'W,睫6G�T �-��[c�i�F%ȈY�$�hslY%b^b��1���(Ԃ��aD����O���\�>���(1,#���$6O��g㋺k21��4_�-X�B9�N�C�A��~$���J�7Ұx�F��$�
��7<O�y�B���Ms��ޭ �D���7��������v1d��K[�+�q!�∘=��H*�kP��?���-�� �"C�� ��6D�������'��	����e��dI�] v���W��"���7�%�WC��B�:0ӕ�A�v�^�:�'���)@�����$w>��V�;$����d�ȕ�T��`}j���D�q�Le��=Rv��#4�����^��y7E�#U�A��;#����斮���0=��s�o����<a�������d�h�JCK�	FL<�sb�Na�`J��������P�QI�
J0~�����qw�ۨ4�a��[�S>�hz��'���xe#��S'��+t�N�	H`�0��1i�Tp��ˊ�bgh��V.3HP��A�},I$>�'�
��?��`�r̕-V�,�$A�JYQ�x�=��@�vąl,� I�5*����	0Y�);`(�*<t6l�!�<YC�c*��#ҩ�Go����D�>���m��B+��
������:v$��Gm��ȸ �ڻ�<�gOB�=\��V!��o�>�����~��,>Tm8�fҀ_w^�ӕ�P�RJd�'?�2�#I�:%�����p�p��B��W�i���k�����+I��2�d�$4
���ӟ^Ha��)F���R�Y>9�!U�W�Dm���b,j5�������=iF�W�kA*ʂ!��
�t�G -M T�
e�d��GW.;�`��r��0 �.�SpC��Jq�����'��PyS�̤/��uQ�I�;Y����B��6T����f�Yy��� ��H|#C�ڻ:A"��&_�W��$���%Ψ�,�Q}�-��O��O�°Y�c�LL�ߢV.Є�'�O���b�"!��p�.i��-�5���*��P�����'X�ѧ �5Y�y����y�A�X�R���E
�E0. �VX>���5n����	X���韴���Oݐ�cG@�\ƌĒ ��-"?�L�bA�f.䡑��InX����w��Wd�79ux��� 39l�AU�>}��E �r�Z�CV��̸��PWL��8󎊬A�ف�,�=a3�L2jƏ%r��\HB���ēe����SZ�ۢb�X�`C&I��/i�r��)"����3`����	L�>�$��/���s�b�+���P�V�����F`Mg���0���(u�`���#8�)�	1�O�v`�c�Ԧ\H�=�D�O�Y�6Z�&���$�p<Ig@��	ɸdL͚86!�BN�4�D�H#�:���J�@�#�ƽ�5�66���s ��4Kb�Q+Q�t�F��� �K��!3�'�J�p�U����c���0&)F� <0�#t�S	}k��9��+#b%��,��3�	�'aМr*O�PJo>͹����$SذY��ƌxy�ؚ'߼[J�s$J�i���c�+?Q횪Q���Y5c�����$��1Y��ZEΟ�Q;�̔'{�D����O��Ò�c��#6BT�6R�ɲcFQ!�,�:ҧ^"�D�j'm�{�ɧ�sޙ $�G�[`09q� ��|P	�C�Ojt���c�p0�&LO�Հ�,�2ḟ�P��M�mBURj�YJ>�eR4���}3��Z
|6 ��)�m=����0���*g*� 2#�iqN�}��5 ^�32�I�H��(��ID>W��9#���y�้�bݱ$���q�)^�sr�)�3��l$�=�L�<�'l�Z*�ƢIa�Y��ɩd�'�����,K���ER([h��P�F^��d^L��H�l�T�V����
d�����J��:Ȧ�u���i��s����W�ռt��kYl�P����=\~$�T�[7n<V���N��<�O��K$ϭ-���&%%� �Q )Z�DKN�b!��D8�����w�T�gf�,���A�KPH�	�l��ϧn��z�Bա:�6���z�`(H�@E$^�����=��\��K��p>�w%�=� (�N�:�t�����Љ��	΁|y�WE(*�`�h���8�z�~]d��'��fL�I��TZ��L�|�`��"O8�a�c{�X����#+ôl�wW���D�\�اH��x�Va���B�!`d
m�X�Ir"OtU� �V
�ܑ�#[x�F���"O.X!AL� ���hI0:qV��b"O*9�� M��Œ@a�vDB"O��ʆ&D $���A�4~�ܰ��"OT�L"|��1B��.�Z�)F"ODEi��y!��s�O�!EXC"O� ��Ռ�M��`�Dަj��e"O�)b��Q�R0�bĒ�	���"O�L	#���wl�TC���"g�S"O�倃��6,GLȃw�. ,a�"OV�#B۝h�p�3L����A2"O�P�K�	HT�d
1�\4X�\4Jf"O�\����`���(2��I�B"ODxje�z�FM��"�"m?��)6"Oآ+�"��z����
�D��"OV�W� � q9�A�0.E�1"O�鑭U1A�� CA��W� ��"O-Z@�Y���s��؆R�x�"OF��a�ѯZeX0� �1�L���"Oj����J.,���� i��q"O(�{%�N
�c��?P�;"O�rs�� �Խc�"K-> D�i4"OT��`�
�q�Z���?8hԸf"O4�����&,���o�/Az�l@"OJ%	�K2_p��:�-�X[0��"O���qn۲z�8勆���N��ڡ"O(!�4̃���*���(*�Mr�"O�Mi���3%��!eE�9&&����"O�qx`@ͤo������[!�骲"OLSթ�t��9�2D_!T�jd"O��q]:\����^9E� ��"O*:�K�tAjD��:���1�"O�� ��SKP5���� B�f�ɷ"O����e?2y��$	 (�Q �"Ox���_�Vr�y���ghx�r"O0TC�JW�\b��S�`�ɰ"O�*�l�o*�`���N�5�F\�v"O��5 �*'^�YQ�B�d�g�<��B\:2�i�#&U7Q�%@��~�<�`
D�>~ +�)��]n� ���x�<���<�t p��
CHMxs�s�<Go�H�&�!󇙃-���	�o�<QÉA�NP��"��?j�깛0l�l�<�R-�1 ln`��L:<�(�ij�<���$\����*�v� �HR
Pg�<�$f@J������<�������y�H� XVY���pn�ig�C4�y���:~ЄT�2ǀc��M�q���yr�Y����C�/C����S�y"��?����Z�3(���A;�y�&ǖ0���Z�C��vHF(�y���
[zXA�5�\+O��(��L��y�ؼ20���Gn�&Gg��'"ǒ�y��qل;��E�,�B
�yri	Va��MB6�����^x�<1�e�/8���˄��sԊ�0��t�<�J8fI�dc'B�8hB�0�@�s�<��Ao�  �N·yG�P����H�<�7�
9dF�dy��D�_F���DD�<�0i�1tF�P����H�Y�� F�<i��A���rE�Y�v�S �j�<�GJ	#FxR!.	\�����\�<Ap.Q�C���B,�!�i��<�E��+Ȑ�����o��#�@�x�<y�b�f̍c%l�0���RP�<���U�L����
VTHH�cP�<3����[#��R�^�s��N�<I�ܡ7GD�23ǞL80a����B�<�'�<�4�ŪB�7r�0TfLI}2�)�'S���c@�>�z �C��ࡄ�S�? ����L9Q���$�!���"Oޘ��ɰnG&M�r�K ���"O|͂T$�r��4�!�c�BG"O�l����@S��ω�[<���"O��u��HT�}x'(�-=X]�"O���^?
*^��'�F*�	��"OJ}BW/к5D���L��D�؜p@�	SX�$���T�����x�4�`.D���4�&V��R�F+vފ�i��+D����*� �vt9m�> ���zwm=\OP�IM~ƒ8+�RBi���ڝ(@��y� ��3D,����M�ִ�B	Q.�y��,)��I���B�$�Ӷ��yr@H<�F�z#BT@�@L9�Һ�y�V�3��r�딾87`�:#����y��9j
�SAZ4�0ĸB����<��$�PΚ�P-j��%��ăD�a|��|r��9g��!A(�:r:�8�Ĕ>�y�NN�L~r����%jьh�!iɎ�y���t����`��b&$h2$��y�mU�;��iZsFD=b`�I2�K˭�y��-,4�2�A��.�}C��ў�yb��V�8d�O�!D��)e�[��?��'Hz�C�@X:��A'
��ĉ��'7�	��ڕ_���B���>{F,��'�.����0_���*�:@T`��'c����T
ya��1*S:_� ��'�-�*�e@
���2_���z�'� �۠�H� H��Ag�<T�����'���
eA�<�pa�P���A0��*�'}���TnD(o��!#(C(q����'�~٨2�G2l���BfA"iB��'x��N����C��L�Lfv�c$`(D��jU�F�F��1&d�5����c%D���ĝ�JvU� ���mF����0D��C�Ə�8NQI��:Fdc'�/D�lK �ѶG�l%`�W�R�=y!���*4�-��'Gc��a"O�-��"'D���9�e��9a���q"ObhbBE��J��Z��GD0��"O )KB�Ş]����g�
�.>FXҤ"O�]�d�E����@¢E)���"O��KK!1�X���.#'���"O<� �h�{��� X/et�XB�d8�S�Ӯ¸�Ar�0PB�a�%Z��C�	�S��!Bvf��_!J�sS��?U^B�I�h��E�!B(m9<�`��ƌ�
B�I�s@���x�t0�.�q�C�ɕZ�`��6�ޯ ,�1�b�9��C�)�L�s2.
�i2�Ã
;g0�C�Ƀh�ʸR'�O o�t�&�� aXC�	?��:�bW�9��@H��t�HC�I��(Yk�EʗZ�M��4%i�C�	Du�t@�\�zH�l���7C?�C�	�,������	����@k�!ǈC�	&&���Ӿ.�������#l�B�	�>�^���:~��0����mrB�I��tC
��#��kF�vQ�E2�#D�܁jH+���ǂ�'�2(�aG?D�4�ui�3��T[6�Û�n��<D���c�K$ct����G9
�����9D�)r-��_:��pT���J�xA�V5D����-K6{�E"�"T�({zP�1�=D����Eɜn
�0�"�]V  ��9D�� ��0��:|�Hݩ!�B�5�9 �"O4��tbx�J)x�I�(�!"OTp���ǅ[����I�J�V0a"O����㌫`�P���Q>��R"OlX���YV|�gÃ$z���@�"O�H�@ �wD�H��/j�ʌ�3"OF��$
.
�ݠSbX�!	��y�"OzD"� _@nYA/�&L���"O��Q5_�-~�2t�Ҡ���"OΤ1��N-LN�u���/��uC5"OP4��,�04��c��"{��A�3"O
A�%)	b�lh�!��nx���"O�\�@��M�d�ą9�|�)t"OR��@'��5�D�m��2"O���Q@>#�@Q�`@̌,���O�(5癢V�&���߽,u�'�ON�<�7��x� ���ł�2�G�<apZ�j���R��'��j��A�<�F�X~�$��a��r �%�cv�<yQ�ƿV��5�t&R�vX��)P/�X�<�R�S��.�ᢃ��4H��YbEi�<��ƭD���;��?��"k�h�<i�n&Fɢ�Y�j:r4�����_�<9�-ׅ;X��0E&����aIC&s�<d�hC��� �nT��2G�q�<iVO��V�z�����i�Y㇌�R�<Y��Ȉw�l��dFN+F�TMK�c�Zx�dP�҄[��Va��!�(baTY��y2߰f��AɁȍ,]���3N�:�y� �u�Lmf�G�STu�­W��y2d�p�&QP�EΗKQ¹�`��<�M��'��4��n�Q�^e	$��*4¼=8�'>(��V��r� �$�P�\y����'ZR4��AoE��' ي Ne��'|�BV.�=KX�X���vmQ	�'���;�f�'!Q��p�	T'u��h�H>���	�Jx�S��1L����M�5 !�Dպ\]��T�}�PpRQ�2�!���c��5�$��TM3��&r�!� (8���3�
�YN� 
f�@9m�!�$G�Srԝ
���06A.��$<~!�QxƁ걄�[H�<R��6M!��T�i
��g�=s�(0!��n�$�sB昖�T��i�1=!�$E�`X�зe�^���#��b�!���?ɢU��d	#�@�pC�m�!�$H�W��)q,ޣ|sXs���8z�XB�I�?�0w� '-��̩�Л?�C�I:�.�Dn]=]�aqP���:E�B�I�6�13��� �I����U�tB�I�=l� ��l��M����gDtҞB�	Z�L�q�/��
���c��4ʲB�I�{�P�Qa�N�t ���':{����+}"m�U���/�-3 X "K�����(OQ>=�)�}U\��a�Y�f9D�X�g��]��ԫ�¶q�N��+#}�	�P�a{2�M/?"�M��,�dv* �@)��p?�t%q��f�$i�YaRj�F7��Q��0D��`#LғPxN(c�

���R`�-D���7ͫ�"�	�ɗP�<صj6D� A�Ɖ��ܛ����h��'?D�x��J�(h ߉.,��{D�=D�@t�	:_�0�9.!�R�.D�TpS,*gy����W#D���F1D�� l�x��Lx�s�� ~�H���"O�P��+r�F��R�E�X��"O�1{b�J5d����VҼ���"OcU,Yiq��p�a�Z�ڳ"O�1ʰ��#I�����:P���"O����:3��H�6���G"O��J� ނ7�F����&�|��"Op�R`��B��sG�D���3"O؄`0�
q�R����Θ_��Q��"O*u����je��j��9!�&!�"O�s_,x ��"P�N(�e��"O���"��)'���Tg8#r)R"O��DI�1'��8q�Tj���D"O��Z�܄W�eSRd]�G�x�"O�Pg⌆w)���P x�P�{B"O��k@`+2P�L��V�l'�8"Oj8�1��(��Aq��^;4�B�"O��C��C:T��լ�2�P�5"O,)��� ;o�}�aN��J�x�k�"OF�VN3_ n�g��Hs:er�"O�pH ��*t�hHT�)oDt� v"O���1 ؔ
9D��@dD�p4�� '"OZ�2�8{޸�y���N4�eQ"O��8 ʓZ��m U�;0��g"Of��6U;7<�xaA��؂0"OtI�HS�n��1�������ڕ"O�Ѣ�Z���j�HØr6�"�"O
Yp!���V�f� �C��eR"O^5	1n]*^��S�i�&�%@�"O��ҔL_�'l|%Ѥ��go��@�"Ol)z6Ś1|H��A�g��hu"O���p�,�-;�!�9G���I�"OX��E�#!xP�Ӣn�Z�3"O�0Q@̋���I�$�&e�"�r"ODJ1W�U�"�3zp���'"O���
���q�
�l���"O��E�-z}�f�
�@��B"Op}�tMS//�4(��F\�L���'"Ob�"�l�͋7O�O��KE�<��GiT�3���n��
�͟~�<ْ��v�N��a�X?��DAA�<9s��C�X�H�c����!+�ȚU�<Q䍜�q	@1y�F�G�%Jg��k�<!�C3C�rI�W��R�H�y���i�<�dd�s�@DH&?��		�i�<9R�|�$�*
�R�D��HYO�<Ӎ�B͚�[��H�uAd͛�*�Q�<�dY"s뒸�gd�n�tx#�� P�<�/#��
�9+!���QOM�<y��R2D�T��C���c��<�@(�H�<�� 
�B�@��r����FTC�<�AJմq�h��������5�A{�<Q1N��>&J0#A�ߑb��P�O[�<��O�cd6ɳ�'Щ@� 8��BW�<Qrg��t��(P`�Ѧg-����-W�<�K�Ya���k j&�ذ�yr뜄
��K�#��c�:�8עF�y�G"f�2�١��^�ĉ�����y�hi�< 
�-M<P*����,��y2�ۃE'� Q�B8>s�	�5-V�y���)qlʼP�iվi-��Ԙ�yBGE@qt�� �[��h9���ybo�j��(��Z]�p�6`
9�yRl�P��<�I��MI��z����y
� @t��FW0>��yI�h���ۅ"O��`@�àz�R=��:����A"O�����>����4�O��h]q'"O̔M�w<�����r��EA"O"3cȀ  ���&QdHT f"O�� li�Hm�r,FÊ � "O���ǷD 	�׫�mO�jt"O� r��RM~���ћ;I�"O��i��K�j��늲c�ٚ@"O t"6mT�)�b���A�?�@Q'"O�䒢ϟ=~��S���#�+6"O�ܡ� V�X{֥�BE�"~d
��ȓG����F��L�[&��(yrt���?L����ε���:�b��� �ȓ<�v�s e]?b�}������ܝ�ȓ_?&Թ��t3Xb��F9�q�ȓD6�`�Mf�.ApW���|8��ȓi3ꡒ�M��2ۂ��@�$�<i��=�F������6�x���f�<Y��@\wZ$�`�B5 �����B f�<����,"D�)�.�0Y| X��@c�<	K2e�ԫ�G�T~&��Dg�<yug
�w�©��-|��b�Qg�<)BG�!F�`�	�w5���f�J�<����4�ٵiߥ7��|"TGY`�<�a�@y]�lgA�$+Ly{ҭ.D��Cp�[�8\$<�A�CP*��U�?D���Z�s=()d��tl�a�tK?D�󗮈�y�iҶ�Ҍ8U�᠖o:D��b&@ęGF�|SϋI���C3D��iB�J��+%�>*h:�[�M3D�(�b�m6iQ�Ä<D�`{�e.D�[�-ڣ=�=��JM0 ��
3N*D�H0�����G��w����a�'D�Yp��!��e���J����$D�dH�@�kglI�g����Ă#D��[�H�$2,� ci��Hh���U�?D��c� 3M^4;r��
��M$�(D��I��B�զ��Sb�ݣ�3D� a;Jr���'F�$Uh ��5D��%�"p��1�be�8[�$0�)D���3��p�Рy�E��|/P(D���IG�yDM�	!��y���$D��kK�U�qa'U�3��r�� D�`�2.қ'I�g��5*����+D�����A�x���ш=8��*"�<D�����ܳ%�D�d�/�\Mj�H(D���G%V�0-f�`���N�@���2D�욡-��>�:��31I�{RK/D�$��Ɵ�iJ~����Z7,O����0D�h�E�2�� �ץ�(vи]�Cj)D���ًLބ5�bIE1פ�->!�$@�_j�')��t4�r�l٢q !�$=��-���'2$����ʟ2!�߃}����γ3�}��i\0#!�$�4r����
< �q�bǗ�1!��I2`�mA�2 |<H�eW�u�!���)fov�"P���pL @�n@~�!�d)n����D��w�5"ŀ�9T�!���@tA�ř	
H�'��<{!�d]�O��`�U
��Q����+T*�!�d�i ��u�]i�ݳP�I�!��43��u8ə��!� �S�8
!�F�jf&D�6�K�+V�����+�!�� �Qꤩ�G<$�c�$�L�z���"O4�@��ndg#��.u�
 "O����7i���ڴ��Gc8 ;�"O ��ȉ;�B<��k3W�|	�"OޘJ�Ca{�l�'!Ӑ_0`՛�"O )[5b�,]b|M�`��5,
��"O�5��bZ�}�0;d�����aڒ�yR�ȇ"L9ٴ��2�6��%���y��L59z$������\��_��y���Yh�e���,k�.�5+��y���og���6�]-W4�%���yr��<���Đ7�,�(t�Z��yB�û[��Ht(Q�;1ޠ�c._��y�O�� ]���A�"��a��ڤ�y�J�hД�'DӶKXT8�"-�'�y�F��XO�<��pG����yr�ѡ����R.��MpF���y")�;`���E�-�,,�����y���Ihm�� �*��t�dIJ
�y��4{9t���j�:g����ˌ�y�hю{ǸYj�e�'-�>�	C�ߋ�yB�N�C�^�p��Bbd���ύ��y�X&Nzز�F�"7Fx�!�y���j��F�o!�#�(�y���M�p�G�A�u�� �y�.X�<w�<*��ǆ)x��������yl|���(��XX\��s��*�y��."��څE 8�����Ȼ�y�N܃x��)�U�1�~��Y�e��v9��3�fC����&DH<تQ��GA���$��t7�,����Z'NY��u�@f*B2Z�Uȗb ���ȓlN��Ė>A��K���V���ȓ3��C��P-$��˧�E����ȓQ���:���=ng�Q�cV{����ȓʰMs#^�1j<�6��o���ȓW�t�a��_&J%FD��=5�,�ȓ!���7Ƹa���a���:zx��c�KGҺe_F�!��Źu�����d���i��Y�!��6G�8�z,��5I֔�HԄ���l� �Ȅ�H� �)EH��`s#�1��l�ȓP(��*S�W'D�6p��.F-KS�<�ȓOT*�h��I$�D��$3���R$��X�#2.5 ��&�$e E�ȓ����0�
�*L*f��0����ȓW���*�G^����~Pt��-:eۃ��bf�IՍ �h�@��7�
�+'B�']<�8G�� �v,��
8�ˡ��nX½E���T��!�ȓx��1�#�ІA�\��M��B����ȓe��]R�6r`��5�3A:�ȓrl��L��5sNέ!��`��+�n!	a�./��p�����ȓI��Sp��9qJ9��f��G�΅����MZ���iY����%-�:��ȓ J ��C 3xĊ�q��ɢH4����k4q
nV��	�G�(g�d�����8ѠIE{C$�3$�� �l���O� !�E�/MH�S HZ�8�A�ȓ�40taX<��!�6#
	2Ʉe�ȓv>��$I�j���*@Dތ��\�2᫂��R=p�Z'LE�(h�ȓV< L
�l&���b4��z����S�? 6�bc�W��| �jjݬ�Q"O�a!��[G������I;Z0Y�"O�s�V(g)������->a�"O�8z��C�4�ܩť��HR"OL�­��<HH8Ѥ���Q"O��[&NG�ei�� �L�(�Ӵ"O�T*֎�]�����[�rP�Ӡ"O���%�)\1H���ܶ
^�W"O��b%��6<�"˚�zA$�ʅ"O~q��&J�Oen��@	c4� #C"O�`�č-.�@@����΁��"O���㕉n������F�=�0�4"O���`�ۺ-�p;�#Õ��� #"O^�j1،$j�]Y�@""Ob�B�,�@12'T�˕Bev�<���N~���p@�[�V�Ȍ���MK�<!���;@̽�3�tmXt:�n@^�<��H7jO����'�;�M*v`�X�<!�ME������;t�� �dk�P�<� .�G ��C�Γ5G�HQ�@�J�<�s`V�0�d�Y�����`D�P�<�A��q��x#w"�1ܰћA�AV�<����.��'��ec�9cb��P�<9�>]�,��7[�.-���b�<iE�&{l��f'V�,�0�P\�<�%�G5dҀeB,«<���2�$�[�<q$*�#f�Z5�G� ����'NT�<�T*ۗ.jV�8��A5�P�W�<�0�E�����Ȯp}��;㧎U�<�SF��Nڜ�DA�.)�9&\P�<�G����AÃL�s��2�GYN�<a�k�\�&�Ĭ'(՜�۰G L�<����x��%����/���S�� E�<Aa$j�~���,![��3&�LA�<�'Q�=-}b%��� ��PF�<�Wn��X�����/e���`wI�{�<�Q&��(ݮu�kC0]%F�w�<���&N��`U	H�@/�x�<ifA�!p��� 2(�8lN(�ҥ�X�<)��*/l@��!g���L W�`�<�ҔL2�@�eLQ�k�`1@��Q�<9`f��̌Zg&�:>�����W�<!�!]��1ɥd�
/<��G�
Q�<��(M���"���A�s�ǇQ�<�En�SĴ��@� f�NQ+�Es�<��B͂E����\%o�6�P$(�y�<BI|���F��Gp�ź �UQ�<1�� N?�ѧƆ�VtA{ǬTO�<I��	�K�(���k�pH��'N�<�s���g�@�DU�bn �Aф^_�<q�#��
�!/�p�*IQ�<1g�oI�0Cpm]�E�XIy" JI�<���o�z5� h�4��"�Y�<�&a�2�� �åӹH�	�#%R[�<��dH9�(��|���ÂY�<���X�T�JYEjox(��)^U�	y�̋��حg3ziҠ!9xYx8�U�&D� i������e�)BA�0D�@��(��^v���Oךs�����/D��c0#z�����1�x���j7D� ɰ悼.{��FӞ.U>݁��5D��	 �ц���0��
>��q�8D�񠃉/3:ArsiѩG��S���<�	��ʭ�&��v�P��aĲ(����S�? 
���C�I��Ԩ�ꟽz'�iҢ"O�E�Pm��P{���u!B��"O�u�䧜b�|]k���4O�`p�"O��bG��$�(�Y��	�S6�ـ"OL� b�?��%sQ��|�HMr�"OP��d��Hb���B��W�$�"O�5�eh��IҨ0�#�1~w�!�"O|�*�1�y�`�e�0ܓ�"O�yxF�ѳO��#�T9I��8�"OFūOժ���� zx�<�"O���ѓuRҙ�ǪR8C����"O�i�HY
P��#J��5t2�"O,U�����`@ɒ!h�h��"O"�pH�,i`\��*�0;q�XQ "O��A7�5>�Y�郺d	f��p"OX���e��$U����Q�����"OШp�)J�D����U�v| �"Ol٣Ģ��rC�cT\���P"OAj���C�z�b$�hr,"�"O��r�җ�v�z�"�Łd"O�� kӃPd�pB�{�ua"O~t��O�-��m��O_$R�.��T"O�A�6O�R�`��Ч�Jp}b�"ODh e^z���CI��[B�	�"O<��+ǀa4��¢�^�q�R�R"O���I�GP��rP�?c��	xf"O��;�� *�L��P������"O>l����#rԀ,hl��(j��"OZ� ETڥB�=3�%��"O �Pa�
uzl���%<��"O$�K$v�R�^:/ fu%"OP�����p��UD����"O����.�&dRdY�j����"O�v˗DxtX@�%0%��a0"O���]�-��k�zИ��"O��֊;6|$�q���se0��"Op�DCE�U�BW��-	X$1"O �i���I���2a�B#:"�""O��;�"ٰ^y�e�ʆ�Fg*���"O`�ȳ�Q�*�³�ܩ.U(�T"O��Xb���y#�+�,�C"O`� �עO��E 2���)�,��w"OvרV�|����#��%�����"OZx	"%��u^JT•�s�8�"OH !�M'T��!}��"O2�s !�Hv,�K�!�>Ktj�"O������]4�	K����lDU��"O������4�H�ID3^f��3"Od `�Lה��0NK�e@2
�"OR���&��V yԍZ�J9x�0�"Od)�Z&Bưx
c	?��e"Oe�ǉ�,�XT�G�,�~�� "OҘaE%,�v���Q�~��"O��k�mN�`& �q���Z� �"O�0	��ɮo�9J0K��Xאыf"O�0�&��9a�)��lb��D"Oh��P*h���n�#Wc�t��'��Ј�E���hT*N��'oj|��k2S��@3 ��A�P@�'���1`쑋$��P+�(�
�'q�&�ʤ�;�G^��H��
�'�T��G֎{ي���\�d��8
�'TA�g�}m�M�TA�s���q	�'rv@��:E�ءĨ��#~4${��� ��[�'E=i��ͫ�H� bZB��"O��:�	�
,�'M��|�jf"O𬓕�ſk=���eM�=���y�"O�����b���q���R b�"O|-�tA�{x���b��$P9V"ORys�H��.�lP��N%}P��"O���$Aݓ�N��-	;'j�M��"O�ܪB�D9CkH\[vL��^��"O �b�o�*q[ָXR��fV�X�g"O�X�S�ِX�y��,´?A�Q�&"O�IC)s��H���5�퉆"O(�l��a�P	�+���ôl6D�(9�A�,+��Ղ�GdЈ�2D�T��(8ht�6*+��i+��*D��@�m��&��愄�$�ν��&D��T�Mx`Aa�*ƌOX�'$D����o�>��qՏ�7;B�u��F=D�T���L�}M�BÀ..`�a��!;D���A�à&�4���}C���!'D�`�'\�a<�c&	�.��U���#D�𸶫��h�JD�*�d!��`=D���*D�L�J�ls�xՑ�F=D����`[�H��e�ŀT'�xQ�a/=D� �d�Y�r�t�$A;n2�s4@:D�8	�Ȗ��`Q�Q T�3r���d/7D���D� �M �a�@���\&� ��9D�B (B�K�Y�@��z�9�<D��"g�D)����|%B[��9D���R	�-�n����0�%D�l��h��O�R�Z�%� i�WG6D��fP�~ƞ��$G��P|�aUG3D�<8ӣQ�F�N�"�Л ̸Hڔ1D�ĳ��^W씒c�O5\T9��;D��B���7��uB���<~��6G8D����΂G����s�\�/4 sD 8D������sO��%-�,fG\��i4D�8K���(V�+���
 � ��.5D��(D�
	h�-r��XO%�ȧJ&D��'�S�P�8�2ă.j�Q`�.D����0߮A+  �9{��@K-D��z���1�Na C e��(3�6D�$q'A ��pK	$�h@�U�)D�(�'%!}y�t��L�w��
��,D�a��_�&��ǈ�<w��tiE*D����bϱи('�����FL(D��"�7	w.8��ȏ!�80��m!D�@a`bK�L����g��({l,@q�(%D�D�t�÷B�=���&)-&[#�!D��kb��2"8�ig�R�2�2���N>D��1�%Q�gO��a���_���	�8D�(�c.
�I�6�+Faո~�3�6D�Z� F*��AIO2I�Oc�<�"�� і�#pf]1M��i�Y�<�u��75�l��+Z{�݃�/R�<��*��s�K�(��X�60�C�Ju�<�b˅(�n�;"o� %����o�<I����0^�	Į�H�ʕ�&��m�<i���[�P;��V��9{5��<i��?��S�Y�(nK1DNA�<�R%MmyF�cVNϿH����<���-v�-7B�2Z�d��G�~�<��߉--dP+5%��1����L�}�<��F��6�ޤxҢ	�'f��DS�<�#C	+N.LP*����UDP�Q���V�<� 6ؒ3�L02�Y�wȘ�6ELYȓ"O��j'`��K��m@@�N�=�~�R"O�3�ш�zP���Y!�2qA�"O��"w�Ρp��(דVh�B�"O�����c�B� ��M��9��"O�@�D�a���roS�g��<��"Op�(D+�'�.�i` �6S��qP�"O���4�ќ^ZLd�5�Ɯt����"O��J��OV��zr���`�<�HQ"O>����P�2Ϡ�.	vX��
M��yR/۾�$�X7I��O�|�D@X8�yB�� w.i�%s��@�	:�y�/^�gHrYi��0vÐ�ABEX��y2��K��8s��� ���k ����yҩ�����GF���v�QF@�<���&V^�K��G
R���y�@]a�<%K�]�M�v��s2f�s�$�E�<9��G>3Pk�ǎ�w�XH[����<	��A�ZD.�.c���"!��x�<��-C|%�	qE(�'*(@ j2�v�<av�Ķb�@ţ�b!sg"J��Ir�<钨�x�,!�%�c�($ڕ�WV�<��&M�$������K�2�T2�S�<�r��%��`n��]�4D1&�K�<�&�CZ������	q��VD�<�p��E���rᅮU�\�8cm�A�<���$IxVBSB�3�ԙآ�A�<I��((��mّ�]�Ծ�BYB�<�g�A�*�޴�a� ��=�3��}�<a֡�<� �zc��?r�E��_w�<�߃�q�4�H�	�l�\�<���$�Љ���)rR���]s�<�����0�4Y���S�����T.[qx�����IbN\4�ܓ�/Û�tP�ӡL� �I����	@���Hsm΄G�4+��N0x�xI�+5D�S�P�#�(��g�8v�^̻6�3D�x��k"v�۷a�"�b����<D�D*t�S�^c2u���0��A�7D��BW��?8~����lC/"F���WG!D�Lp��?/�T����TQ ā#�O~�D�O6������o�H���8-wdՈp��Oz���Od�$5LO��I��2�F��jQ05����"O`��J�;#Е�5iG/k��3v"O�4�vJ�44�3��X4 -�E"O����gT%�d��J�0G.(M�2"O,8¤+��_l�Qx��1�i��"OB��e
��r���a�'��7����d�'���'�q[`
+'+�@�Q	z �f�'���'p��']$��V�N$<���� �"��P�'�6�ꀫ�b�$jb.]�z�.x��'~x�����P��Ag��_��I��'?r�{G��=����@�=��
�'�ƽ
�&�XBP}$]q
�'-��bg�;�d1K�'
lٲ	�'i��B'��A&Qz��J�2Cz���'I�Y7�?Zy �r5�F.�D��'��p[��H;�����*vA����'m��K�P������F�H����'[j��&큚&��u���Z=��'��xB��� �D�� &��eC�'d`H�a(�k�������;t����'���Z%�G�5uxP�ӌ+\��'f�8�s#ڄU��0�5�-	�x�	�',�@I��I#R�SE��+j�PY���� ��a��2��9�dIH7Y$s`"O�5�eM_#�H�q�aD�-l��"O�P��L/H��ݠ��fzdSS"OJ��.�?g�����ܦ<�FE!��'��$C�(Z��j%Hi���h��8�!� B��1�ݑ!�q��e��O�=��r�I'cѨ�)��O�G_�Hp�"OD�-�	|i�iI���U���"O�C3k_� -���h!R ���"On���+�ze����t8�L��"Od-p��Q?nbl�'ƄXN��E"O���&�� ;a�@ɫ�"O�x��B.{�����X�,	0"OtEI��Q��!�0��*i�}Y*O��[<Pd�p K�,?ʕ�'��"«�\�b,b��� +����'� ě�Q7�܀t�ǌ"�A��'�,|c��Ϳ.pvВB�
�P%�uj�'p��15��*~�X��ӧHb�X
�'��7	g����0���G0�b���hO�#~��ǟ�6��)�#�S�M��p7m}�<��E\dk6�Ӏg��5�eE|�<� ���:��%aܹ|��a����@�<a�E�Rt^�U'+@lF9[� @�<���хl�@�
`Ɏ�m
��{L�U�<Q3�u@�!�	W�E+�J�z�<	'HƶY\p�!�ސ��ҡ�Dq�<a��
7g���Q�ӤD*�����u�<Ys �;Q��E ������l�r�<� ���Kvy���y����#�f�<i ��?]��EK�S4�64���m�<��J�y��d���^0���C�<�!lI�z�ĉ V��.s��2phZ{�<!@B�"h����:���V u�<���.�퓐(�Xޚ��$� n�<�D�ǝKR��Cg��ʔ�-�.B�	�2S����N�VmӀ	�7-KJC�	'L6<��,O�SIT�;���q*C�I�,���#���6�)F��iK�B�I�/���"�
�u�<`)U��_�B�I�^��@rB�/!�졐�B�&��B䉼vrU�*���
,p5jԛ[I`C�	";���$���E��]�RD��X�NC�I�7�� ɣ�I =�(���G��>C�ɪno���jV�ּ���&��R�C�	$Ol����|�ʐ�K�q�C�I�)�h4�2$�(7��@a��RC�ɬU���h7��q&�Xi+�3q�0C�Ɂ-k�`ǡY�:�V�8$�_�GfC��?"9T�!�G� n�B(z#�ȫeDB�	�jg��B�Ck�Y@�n�jhHC�%|����'^�.y
wGҲ\�O|�=�}��o�P������|@@�����_�<Y����W��\� ÉU]����KX�<1$�N�W�܉3�;{0�E��Pyr�'a�wy��q�F���O���#��V&�TB�oh}��M��P�Q��R+*B�� S*����+DFr�i�_=NQ�C�	!g��ea⌖�?�Q����6��C��=
(9آI5Q�Pɛ��Ԇ:<jB䉸9��YxW�+�bX@�
x� C�)Wq�c6+ ��$i؄ꋄ/��B�	37�.��4.�~��@j�DZސC�ɢ�B8�0).���".A�F>rC�)� ��P�퀊hC���3�7�,`ɇ"Of!�0.��4P���vTD�1�"Ol�*�],!���S;_��"O�i$癐1"\�*�*X
��:�"O���Isay�5H\<q�"O�ˢ�Jwf,��'�l�2p��"O@A�� ��ubL�Y��]�}���"OL��G�Θ3��`H�*[��C�"Oh�ф�Lr���q�����|R�"O�M1�)[�v$��ae��|�ܬ�q"O� �Cի~`�+�
����""O���&�9j��0�Mw��ҥ"OL�m�~v�B,K�_m��S"O�81⭜�[W^ap��,j�D*U"O�r��D��Ju���<]���"O�����X�B���ڗB�lZ8��@>�c�e�:.8��n��(/�D���3D��)�J%=!�MZ��lˤ�!1D�ЈEǺe@��U;A�<+b�/��M����"�vuؕCåƄ -,�!5�,D��3Dj��q�#6m�?An�q��O7D�̐oХ�
����?�X�W�6D���#�G�u��l��%��o�h�y6�4�D�<Yç�4c�K	&Y���%}d�Q��V�����D*R|�E&�8�$@�ȓ<2��BE��%H��Cd��jG�t��:��qS3��6a�%i%曹Z��ȓ��D�b'[<n�h0o�!v9�	�ȓ	t��� ��W$����B|��!�Rt��K�w��t�9 |!�����I{yR�'��󤋏qӪ�au.�����	5�B�I)/:�-3���o"uB �o��B�	�|� L��.կm��a�� 8OPB�$!R5raΌ&�� ��*C�ɻNł�
G��4%Y�E��!L�C�	&r�<%��ȏ�5k����eR�B�ɕ�`�!�۴Y���#��݌l	�t�IKy��Ip®��V9���H抝N�B�B�N��J��H��$  'I�g��C�I,a^�U�`i��Hj1�F�=h�C�?sl������IY�E��^C�Io����g�H�PO�PãA���B�I�
� %�#�^>Y2x�Cq�.�C��:t����G�D���AM�m���O.�=�}��H�#���z���{,@1A�Xm�<Q7GZ e�z��j?��X�dȋk�<�����1i�l�w�!��[1�g�<�f��SLBu�ޜ=s�٫KH�<ua3�H2�"C���p��z�<��$��Rx�ā�M!!U8px'd[y�<��`��3{z��Ӧ-���q�<�CܡS4�(�R!�~�r5��LJp�<��)��Kd�!�Bփ#�8�ؕ�Jm�<A�F�./w�y3 �
b��H#��i�<�u�0 �Ȁsd�@�h4��t�g�<)���%/(|�H]6	�A��W�<���?-��y��y J��S�<���ML0�qǉǮ*oH�I ��w�'ia���ԧ�0�emM�V2B���G��yRbW/4��)�Qo*�;�Lޕ�y2�,y�T��&�»GN��⑩_��y�J��!�l����ݞs ���m%�y���}ز��� 0fc�q 0���y��I"��p�hU�d0���G��y
� :�cU��t�(�嚿(P�ق�'����p(��8�����	(P:7�+D��Kֆ!(3���eE�7N̛է*D�`���*r>
:ϗ8[X�� *D��+Aő����� �_�$��$'D��AV�ޑxmh��%������L&D�h"wǒ�u�N���គRIJ�##D��s�(C�J���ZA�ٖS����Ta+D�����ޅ'��y�����ch4D�,I`�r����R�%[����� (D���a�"}Glqң�#B�щq:���䓤��G�V�fe�c�,v���/G>g_!�ɯrѸ��&/[(���+�!��,���z CՄbT�d�%i�@.!��Б7����a�%=���5��G!�d� &� ����/`(v��C@�_�!�$V�4��"�N��\��!�Ē�U�I!󭖩>o2pG��ўԆ�=�@��"�K=)���@�ɀp�NC�I�G��pv�EM��[�dC�I2�Na!�lǁx�6���h\jf:C�I5��9�ƃ2N�:I���E�g�C�Ir5�9h (�z&*q���C�ɀnΔ�9�I�.�쌷%.B��:\O.2��%2 ��	�d
���d�<��O�l���W�am�!q�.�/ApA"O�yГ���U-�V(��Z"O�|�7�X�x��k�X�PeqR"O�r�57�2���M��f�!"O<%hҨ�vNy�SJ��?����3"O8$�3 �@A�@*C�N�'���A�'1O��$�<!�R�¦�;"H����"O@�S�`U�<��WE(YWJ��"O,����6�L(�0��4w�|��"Ovp�3��.��icn^aeF	q"Of}a �K<76H�#��MQ �"O����șE�\�@cJ�<J^�9�"O�M��f�~{��A�Tbh&�@�'1O$As`�ќ��5��F��
YQõ"O�E�T�=�� rd�!#V�}�q"O*]�j)�I��^7�{a"O>�(d'�	r�b!J�2	>AQ""O@q����{s&�)Ta���8�""O��7,T�G�j�+��'\��-��"O��1,��/~R$!���7S�����'��W/�8�i���M�e��O�=���$Y�~�F���-D���9�B��:(B�	;_�0Y����:`�A����	��C�#3��@�rHY%~q��<�C�Ƀ|�9�eǟ�E�~!��G@CmZC��<�+�;�zݸ��^��B�	�#�&=�@n߉gH��Fj�� ? B�ɔT����B�>K��Ự�\!!�B�I�,�Б��c��^Y`	�m4��C�	(V213��G�tSNu�7��4r�C�I`@��A3i�8-������*C䉝?s��Y�h?_F��ؑ��F� C�ɿ~�Hsb?v�8� �a�B��v ĩڎ<f���*f^���8?���O�H\zA#��L(Mbp��oy��$$�'~�X�5�K#�����B�Xm��ȓU���B$��&��4��T��y��+�:b"eB�xZ5!��b�y���m�R�O'
Kl���C^�\��S�? ��aG@<fє��o�2�D	3�"Oj����5e�hQ��.İY���`�'2��@@�!z�
��5�m�ZըB䉁\��LHc��6Vzu��'�vVBB�ɧ!X8Jt`@�<�ra��M	V�^C�'Ԧ� 1����k�L^�N�RC�I	 �����G�r��QX�曮JC�ɔ��Q�1+G+)z���Y6B�=<�T(�sHQ"1ʡM`��2�I�e��Hr#�I�U+��\aBC�	
Sb,���+H;����E/�.C䉳!��Вs��>а���)�C�I�T���G3R�t=�#&U;>nB�	�T�������8$r���Tg
\B��)�\�p/Կ[+\U�E�ВX@B�8ݒ]2i�*��pEӼF����<�����fФ!�)�`ٟ\�ܹD"� �t�fD� ,���G�)�.B�I6|�a�Q���,(�FlKE$B��0M�,��.�$a��oǌi�:B�I�l���CD���r��D��0B��}���юL���YꕾW�C�ɊS�4�!�'u��4�#/��C�I�(� ���+S9����UO@	2��B�I>1sv8)P/R��@�u���h��B�		{�z������ْ ��P��B�	�`�,��/	(вXC�H�?aDJB�Ɏ@^|J#�����j�K���C�ɭA�*q�fF�D�b����!I��C�I�,q4`�L�4l�XH��5%NB�I72����AG[�=�GU�7�C�	9L�dt�(ƍ+�b��%�5��B䉐B�6h��a�K�r,i�JOq��B�ɤC�<�s�DY�Bta@*R�B�I�~��\���27�R��Ł_?_��C�I�u\vtb�QZ�h �tmJ�B�9)z�50QM�22���[58��C��3M�0l��	P��9��!=nXC�	�� �s�Qi������(�'z�ͩ���*(6�ABC�Zҁ��'�lD2�@I=��y�Ik�Z�'K.���)ӠC�����>@?PL�'�(�C@�j:昸p�<-�i�'�(��b�[zP�!hP�"E�	q�'�p` �r�<@��7(�θ;	�'����(����q���"'(���y��\�.} Xc�	�b�Da9fJ���yҎҬ3e��
�b��\�б�E���y�ۢ�`:6R F6V(uK���y¤C_����AI �;Vn̫���
�y���$N�`��[�/{=�ӇG2�y2�H�+(U��R�&4���b���y�Bqft���'��J�"�K�)��y�$�16tIH�aS�A+�ȓ�y��ľY�TK��>:����� ��y�i�ds��{4��')i�����I�y�cL`P�$�Ԡ�Zͱ��[/�y��}��C��߮�|Q�T�A��yb���-������-
�@� �i�-�y�L��Kt�T�����
��y :V�mr�� ��3�C�y�AR;lT"���Ԧ""��bS���y"�)�n	a�&��s4i	����yҨڞ-��&� �Ό�C�Đ�y
� ���G/ԇE�����V(��"O~��B"D�k]��8t��u�QF"O:D3��=D�`�㋡I����T"O`��G�,E��$�v!�}Z��"O"deC)m���(G���px�%t"O��0��,�J4�S]�s�di�"O
�����}���cNݪDh		�"OV����ȳ ��1"�^�%��)z "O��g�L%q�N1w,�% ��h��"O�e�`m¯~iYa��ݚV��x��"O����Q��S����v��Ȼ�"O��u�=*b|h�%�	&����$"O��Jŧ�6�af'�/R�����"O�9P�k�Z���#�M�*e��"O�0�[!�(У��%@�`�a�"O,ȱ�,�<��,´Nǒ��t(�"O2͓1�nnR=�AĄ�m"O���LYҡ�� ռ��X7"O���̇,פ�	vM�"�.\g"O���5�	�K�X�"�»G}�q�"O 4��A�=�J(i�&K�HW�Iѱ"O�!�Q&��gS��˄L<��Q"O�� �� \:�̂dn�D����"O|��bʌF�ک녍�-��;b"Oq�#���5���5#�"O��B3���3'���x���d"O`�#ӈ�Fu(K6�W"O�����39���%mC�I���1�"O2Yi�-A8 OpQk��+P ���"O�T��jT.A^��#៬x+�Ik6"O���`T�h�K&���q˄]�%"O¥�/Ƞ}��- �-׸��Q��"O�`j����̢(V�ܫd�~�k�"OT�Ca�G5<x�ab!HҶ	Ċ��"O:���땾d�2-��@��`�.ͳ!"O�8�(�D�f�C �~�F4q"O�$��"Ǚ.�tySUnI6��`�"O�H@���Pv^iz2�_�mw�ڑ"O� I6��g�����Hb���"OѰ�CXb�$B8t�RӰ"Oꌢ��<^�8&��� ���0�"O (&U�!�d�(>����"O�06���gY�]���R���"O�2�oQ�,�\Ċ�G�Q�P�""O����A��Rw%*������"O��ҡ���$О�u���f�*���"O�D�H	J��@!�Tqw��+�"O,��F�����fbְ;�v%Y7"O��A� I^���q���SҔX(3"OBabFb7@��B��X*�ui�"Od�A�(	���.����"Oۣ��y�:��A��\�ܙ��"O$)��_Hc@R�Șu�T� �"O��7n��dFҵP�F|�E"O")���0��h(#+{:�U"O�m[u�^��=+�П>t�8i�"O�%�EE G��񤔓V^�U �"O 2�8A��ʂ$�|I��""O��9CJԄz�1�Ff"fJt �"O"�ٞO�Zt����xsg"O�m���2��MH�"�09��Y`�"Oh��R�Ӧ-K:��C�؍~���""O�����D�<`s��1����w"OB5��n5;��PZen]�l�f}K6"O� �y$"�H�AN�u�@ed"OH��ޫ��d��M
�9WHu�"O$-�'��	C
|Iq,� AB�aP"O>��b��h)̸s� � ���S"O`!`����9��/�Q�Nm�4"OjeKd�D��A[��Ǻ5��$�"O��{'�:d���H�@֋e�q�"O4�2��	$T�����n̈�"O�|���H:u���Z�ze�I+F"O��C��	NА���*K1'�I��"OP�{v��7nM$\pҮE�8�(��g"O�p�ʆU�j�s -ʁ�N���"O�5r�i�}?@��rA��� �k�"O������: I�������F"O���n�Ŕ�3V���e�"��f"O��)��O�<��)
�RE��"O�]r��m�ޥ�2k��Va�"O��Е^|�(A ��Or�ݺ4"O���U�-^�$K\�uX����"Op��r��/
Řcj�	f�\@�"O�YĆ��XgB�����;��y��"O���I�*�Z8�d�v� ���"Oj��0�0(]�d3�M�C(~5p"O���E�I4WT���炤6:J�R"Ol��Y�3�6i+��L��Ig"O�2��_D�FQ��*��9��d0�"Ob,8�/]�{f|�$ �#=,�"O41S��s����B�T�%�w"Oh�I� �Y�VmHU�	�q���Q"O>�C-��k�$�TbW9 2�2�"ONdX�`�-�����KsR���"Ov��V �D3v` �AT(Q� ���"Ov��b�,Uh��p�J��&̠��"O �X�g��@ �	�]�b���"O�ݓ׌n��Q��I�W7(��Q"O��y4J�$�t�Z��ͺ0�)�"O��c3�L3J#�A�!���� "O�P�AƖ\��8�Q.�1#.�ٱ"O�`)D��'F/,�z�
��O���"O`�Q�Ո�R4�e��6�{"O��0l�U[����X�F�H��"O��Hƃ�A�bEɄd�|��"O�	`a��o���`��}� ��"O��2�D�8;��|� �/D��1�U"O��b��9w�<�����"O��'D8K�QcQ-πD�ua�"O��)�� 5(����\���"O��R�kD$5�X�"��$�t��$"O����.��U��⒙Rl���"O ����8$�,L>,�"O�P�P�x]�V�˲(n�K�"Oz<�&��7=
�yU�^tGp�*�"O�hʀ�u����5�^i��ӣ"OR�b��%~�@�C�Ǐ�<����"O4mڴ�\�c�h��S�T �p4��"O`i�G����%�4o� �+b"O\u��;/�Ȳ��"�TY�"O�i��JG>�p�&�C�%�!"OZ�z�o�0�I!e�מP(>�6"O�j��%A�nYHRn�����4"Ox\"��	�~|2C���@��"OҐ�� ��yO\����v�0Q"OB	�E$ 5�ʃ�#9���u"O�T��3|k��0��5z#>Y�e"O� ެӆ���VJ�IQh��j"���"O i�T�	Z6������<b���"O�!�'b�n�����'��a`�"O<h��R�Z��ɖ�U /��:�"Ot�I`+"G6�[��J"Ro��0"O<i��օz$Zؠ�JJ�8��"OqHEQ�dG�� �	M�|	����"O栃�'R� {t�H���� �"Oh��w�Y�aB�a$O�P��Qw"O��q�Ϗ2H����G��r�"O� �QJ�<(���!4��x�2@"&"O< �Q:}~�����F�7��u�"O�U	���q����we�!Q���H6"O��ɴʏ�p� �W�K�"Ը��4"O���i�C8����
�g�&�{�"Od`e�@V�)�4N�6$�4"O��qR�w��J�L\���xɠ"Or��1���\qj�E+���P�"O���jO$�|� �D��< �"O8��4@��F��!5br"O,��7�]�+pL��-q����"O��l&��1���,G=��"On���P�{����RO�2l��"Oh!�6x�M��Æ;w/�a��"O<��'�	i�i�f +t�0�"O:��v��Cy"a��S�'px�QU>O�ч��Z��Lɧ�ߝ*�0�H&I˛� ����O̒O�1�!-�kw�=h�@��EI�uQ"O�is��/U��q��B�E�����!�S�)ڳ,��4�pb 3��
 �zA!򄂉m��XX3X�X=N��!��%v_!��.FiЈ"��3d2��Pլ֊
9!�DW�X7+�N1w�|,c�kؾ`5!�$d�!���=s��Ȯw�Il��~��������@� ]�ܠ���u&!�R�|SnŘďƎ|c̅���V%!�Dߞ�����δ8JJ!�F��85!�DCk[
Q��~��Y�w�̼"`!�Dۋ[�<�� ������ɬdY!���rzh!�0U3��E(Ц:H!��L-N�5�A'b��`��̭@g!�ްe6��H�W&,��+��Z�X�!�,ABLQ��Ir >4dM��!��o��-Y҇��^8�EΟi�!�dE
LE��1 	B��u� �
�x���c��H��#Q��d�l	�׌M�\#���"O�<"�HJ����a�89u��PQ�Do�P�'�����%;z�&Q� �B�F�����>D�D���Z�,�9���u&��q�o9�D%�O6t�&V�7��+w� g� �2�2�O�y�R��-16�����ΐ-P.����	P�<�f��`e���;�ϛ�G�P�=��'T�F��2����	%k���@)+�C䉃��z���!(�e��`K*Y㟔���'�2̑O�(����0j̖'?xWxh<I��S�sр��8;�|;�oI)I�Hф���m
��9g�����$م��R�Z����vr��DjZ�=�ȓZ�K�C֠ܪ�`L��G~b�SH�tK�]�F���+ 4WBC�	-��\��,MJ�ht8#A[��C�I,}�9�ė�jLy1&W�B�'vQ?�; "�&B6��(����hŔ-��-D��b��$����֩��8C'@+D�� �"eiǽG�l@:���4Πۑ�	�<ɎyR�O3�}�,���%��N]<���'=���F�t.��dR
�jA�2f�X���gT���$9��h�:m 1�׍F� ��V�Cipe*��i��d�[���O"Q��}B�����%$��Y��'�	�s�tbw)I�PZ����. N��p?�6"��8�r��1 ����LCP��hO�O�8D��22π �� AT��	�'o�A�vjAS� ��rLţ���ЍyJ�q���']�`��a Ҏd� Y�TGO9rN�ȓ)�E�F�+3��f�ן�\�ȓi$s3,�R�h��˗ 2����,��HS�|�ꔳ�-����jƾ�I��ʣ3�|5�� 	rN��U�ܐ�C�+h>RɂDg�Z�.i�ȓl��x���%��*�D�4x�'��'jў�'Gk��1�n��P�d@0E�П�@(��	z��W�#a�"���x������M��|-D{���'t��Pfj�0�E{âפ<h�أ�'Q����GQ�b��D���� B�e��'׬�'��.#�d�B FE�mE����'v��h6�D.�-; �)_帘
��x�k-c�x��R���|�>��Ղ���(O(�=�Ojz��@H[!2��yJ7E�,k�(���'�܉R�i[��u�W�]�i��*4�2��:?E��i"�\�V�U'����b�7�~M�ȓ"��ufJ1K�=K���-��'H�	Mx�Dqpdt�D�ALY�"y`�2f`5�O��\�h�ʃ��c*:Ś�>I�f��ȓ\[����ܰ~[�H*�+ȆSؒ��ȓ<N��
b�U=$_�t/�=|nх�xPJ}2�F Q�����+�Bb�Ԇȓg���tkƳt��@�EG^$�D��	\�'넔����)��{�
�W!^�����'����lW�U�(	Ӧ.,x�M<�s+|O"	��Y%x���$.B.*0T�3"O��	�� �v��t��'bGZm��"O����%\��=(4�\���"O��s��0ژ4��1A���"O*����pT�p;��Ro]���"O�l����ܹj 鍤u("��"�����ɗP�R���G�-o���$W�e����Uf}����iZD�	�؞8S`0�ǃ��y��1Ԭ� �NN�8�"�kG��y�9���£�	2�z������=a�}N�$lxyC��aˈ �Q��Y�<����iAz���$5@���`U؞��=�!�(Ri"�!N�574��B�H�<ᗨ�0P��m@E��O(rP��F}BZ��%��g��|�|�bEKʃ��9�2!�./�B�榉�BfǙ�n���&
�z5/=�>q6�|*���'7���n�<c�}��@w��M�<�QN�7f �R#�$�H<JTSI�'��x��Y���A'�(���,���,�S�O�Z�����s(^�[�'�T���?�
ӓ�B|r�(��7y�Q�;w�b���I5o�則U�\���ɨze���[u��B�ɵO2�K��N���#wA�/U~��hO�>5�g
A�M�X���\�@:0�*��$D��#��|�B e�YC�6�j�#D����G
6YR��M�<.K(0��?D�Ȋ%�<w�$X���J.o��u�-?D�$c�ۿ#C������=0v�z�*�O�P�H�H�GЏ#.T��Dȕd�uّ�2D�� *ઢ���Z&=@��!O�
�p"O���@���g"��4N-�����'�>��?���@(:<� 7��)���9C`��<y�{b�'ڠX; �܅'��!auYZ��	9L�<B���l�S�'Z��\9%bM�<=�% -y�R���rᒔ9Ќ	���y:rmōNk&9����O"�S��|���!y~|C�,2 0t�@NP��yb
�sg�i�A^�,������d-��HOxL�D�.G"@��AW	w$`#��IU�O�pܐ�G�:g��%p�Gڵ�����'F��OH5'p��B9�R��'v0�@��-b.	B��
��T��'Tj�N� ,�����	MP��'#�0�7�G�H+�в+ �"�x
�'�R9IZ�꼰"/�qi��2	�'���+�=�����h�d���'j^�1j�5x���{U���*X:���'4�a1u�����b��� {	�'Ւ�z��U�/���l���`�'�~�cp��Q���&	��8�^8�'[v$I���`?J�6KB��lB�'(��@˧f�d��@KL�
�%X�'fp0{��O�9�<�pJ�/8�!:�'�Z�`�
u5�,B��)�|���'�<AƂ�Pr2=�sg���:`�']��1�jе���@cW���x�'� Ba�� /�e���rn�ܲ�'�Z$��o�Eؽ�����v_d��'7l���&X�,�L:`�ˈ\H�r	�'=`[�.r�X��ϟC�,�x	�'/��0�i*U�d��d�C��)	�'�z�K%��X���+S!xD҈�	�'�,�xF�R�B�(�jr"��w��9�	�'��(��d�6 ����W9k$E:�'�X����T,���G�N�\�'�H� ���
R�4����M�>�k�'p|���W�#�MX6h�-B��qc�'�h�A`S�@>*}��X�>f]��'��p��N�"�J���`�	2FHp�']���摟@� }��Z-b��'�GغC\�ͺ5j=�T@�'�~-��N�c�0��_G��|`�'��aKd�+]Dt����N�g���A�'��M��,� zы�nM�t#��'Y.�3H��Z@��3vN35-|���'RH��Uą /AQ�g�;2��D9�'0�Y�M��>�*B��K2{鐐z�'q�7A7ri�ex���o���r�'��kt���Uza�t�[2g`T��'�Ĥ��EօM���X��/����$U	Aw�L�3��D�(��b��O0!�DҎ^n�� #�C 9��Oq�!��M�TS�o�1.�2�0�]$4�!��^-4���W������i{!�܏E�L�!�GU�E��E룠��Iȡ�d (ؖH�D�X��؂f�J	�yR��3�8z��Q9�\*���y2��>01��b�V^T�jwi�=�y򮌁!�@y2�M5E踰�GI�y���2!X�G�Ĝ$ -�v��yFWW�
kC��w��0	��A�y2FW�D��hEg�h;�4�����ymJ+D����˚t!tn��y��m_,�R$�^�Xa�Iq�ɚ�y�	\�>�p�����&S��B�'S7�y
� 8A��m��K���ZBh.%���i$"O�};��H ?��¢ʞ��e"O��*�{��y��G�=6�J�"O<���D�Y���Zfg�7A%�"O��2�ꏆrЅC���v�p00"O�����S9��	:r�ٷ����"Op �׈��[s8���Ò68�m�$"O�����ґY�U)7�C;�Z��"O��KqD =�֜�@�	�hp&E��"O&�:JZ=of`��B%:`�1
3"Oh3�Pɦ�RԎĦer �w"O�w��
-zf���+O���Z%"O��p���_t�ׂ́Ҩ<���"OvP{��=mr��p�T��A@3"OL*fg���Q�'N#܀s6"O^)qA�L�I�ʵ��-�H8&uz�"O����ކ2Z�`�D7ώ4��"O��[�ӈ"MDd[rn
3~��j2"O5zvL�%(��9�dg�/��X�"O0�;R���zf<T�� �>����C"O����&.W������T*M�
P�"O�Z��	N�0҅�9Z(]�G"O
�[S���g���r�kȵ_�f��%"OА "�_��^���ʈ#�6	³"O���H
o38�jv�ϒM�x$rd"OڥR���<I�$r≷m�&�5"O��v�0X�I:s@^ZF��R2"O(���Z�&��@3�G�aM�q��"O��RS��M�	����L��S"O40XR�6l�a�P`���В"O����b����r&΍�;{z��"O���D��)}�q'◩gl��(�"O��0�*�� 9tCɆ!��ȱ""Ol�
0�/o渑� ,A\j��)F"O�ٶ��+B��31�F#yDN]ش"O>�Y���43h\���.�;Ox%Q�"O�q�Tb�1�2��:@("O�x�s��)Z��"�*��I��"O0T$�A;�4d�`�8rJ��6"O�ٰ�ܒ$���`Ï�>� "Oxu@��'�v4�UN��j�l�P�"O���N@�P��8�%�İ)���"O�d�A�ՏX�t�$�U̾�`e"O��!��&���ŊA��
�"OP�Dɓ,Tt�aRO�:u���"O ��č'����a�,b���Y�"OZ��L6J�ra@@jM*�4���"O�B���.�<��@ǖ)N�-��"O�Mز�	l����`S�|�2q@�"O�Hs#A��Zz���V��V�8�"OJU��͖Qܰ�z�e�}x��!�"O��o��G�V���D�d�Y{�"Ob�)0�M�Cqt!8���
�vi�"O����w
4�G�_�F���r��'���b�Lͦm+A�>p�j��B�IX��)�@#4D�t8�'ȶ,�@1�Ɂ��5�4d5�!�2��C���(�vicbE�duHЩ0�Q�h�,���'�$��+��y"p`^&^l\��ȇk����琧�}ڵ&�1�~ҧ��¡�9�2���F��W!ĕ�HO�������m��|��� >n�Dh%�āHrb�c�E?a��B)$/d�S�0LO��Z��#���1$�A0�9��.̯49� 	��OB��Şa�ܚ\n|8Ó��$�xD�B�Q"��l:D��T�V(D�#�� ���t"��(R'��{r��'�bmҖkU�w���S��)\�s�`8�Dn�Ny�d������p>Q��N� >~Q2��<� ��5[�yP,�s�( (\�`ZV��SԤU�ǅ�?d�������Ί�z2!��2"��ұn]��(O��BDNK�|<5���H� �z���.G�P�uA��6���u,�h���>`��!J�*��0�(��� +Z�����/�=���>�|R'���U�VEQ�) l�<��mY�l���9�!W_�,��'$���%��1�$ؒ ��I���K�'�$���aA� NdEB������r�[��~*BaZ80�)�/[�^b �Qn�U8��Ў�8FQ�L�F�[�3�A���,:X�P���B侱93��5e6���!�J��S w���a#b���T8 A"ٴ<ʰGz�%�:{��A�����O��TxN�1��qa�S�cYx�-O�G�I}�u1�*R���B�N[��1� Ѭj� 8�I)*�4ĉt���1�S�'Y��YH���Q����6ˋ$Y´p�f��b�<��p�+$���!�!��PHD�	�ipvN�<����!@\X��y���Q�͑Er �O�I��uy��Á��);&�6�I�4
�}-��1�I	�^ o������j#d"�*ΎF���	��*��&��ӡ�	%��0�F�
sIКv�p�=�5h�>cHR鱧a,��&8����E F=b%b�ΐ;��B�	),|Tk$�� X6�z��[%El����5Dt��2�œ/��)�'�6m�Ud�=F�b��T��cR�mA
�'�����a?#�v����P�]����OJ����Š�"���B>��90"ǣ��:FC���~R턡
�L�"w��x��T�ALε�4�_p��C�	�qz��W,yc*�(6��nb���]�ꙹ�y�/e�4���lD�:�r�ҕ�=�y�L_�,���X�˽*+R��G���	x_@� 2���G�!�f�P�b�}PЦ�?�!��A=LC`P�Zi�h*��!-�'h�xPB�")ax2 ��|<@��C$r���'%ƈ�p?�� �	+V�	`"C%ToF�����{��Q��ޟ!4B���p0@R5ek�`���+%��ā$TQ¸�F�<��b��\Y!�&�6���O���Ƭ^��"=�V���j����C"O��RmJSHI���C�A��*�i^�A3�Ci}b�O)"?��)�.E郁С
}��iB�{Ʈ�M����E�#-�ܪ	�a�J�PK�S������?d �U��F�&�B08���)��[-5b\Q�Ȅ� hF������#��P�D�C ��Թo�P=��<����&��x��,C�?�'"R;�Iy�*�� ��x����:��e�xv�0�o��;����D�4p
�8�BJ�#�Q�d�(o�$E+����h,�d+AB�ş��V�R�s���bK7%�A�6ԟ׏v��`\�#�58�h�	�Ѕȓ �1��ɇ���m���G��1  \�(�fp���B}XA` $����iG���]pD��E�>�&(�6'�i��Ik��\�h��'Vx��  �F��!R�5`o��눻X���@�#�T���8{�����n�d	r�=��me��H]�0�KR�'b�<����	ho�賷�i.:(HB!�Z�
a�ȈT�@Y�����B��M�(x`r�a�"�R�$���ɎǄ!� �����r��OJ�PQ옓u�%#���M��	#�%#"��2a(�)� ����
H�M��i�'jҽ �ڀ�ȓ[X
pɡ�]25x���,ž7�b|��%@���	�$�N�K#�7���n��>A�y�b�u�w]`u@2�''5�j`�kЌP�k҈X�Eև$J2I�v�L$QZ�@恋�"0�bĄ��hG�T:��Nd�<��¬@N6M�f�>q0"�[���,�XQ�UkS�S�j�j���F�a|BÔ�#NB�(Ȕu�P��G>- �<���F-'�0H��������� q�fS nP0�Ї�I[l��0ɈW�j�B���b��<1v�X|�ꐉ�S�f�bŠ%�I��is��3vp 4�,~���I�.4Sh0��I�xK ���c�L���Aj]0K~�Ń�dB�	8��AĚ����g:��"I67P�[i4�?�!I\'��D��̃$g�h]�Ax�<a�j*t��4�Y'$�ࡉ�J�$�d�d��L��mrI�.�`90��V+剤{o���%0�����̟iw0��GhU�_+�UC��'�Rг��]gz��c#Q�{Ut,(����_�(4K#$	/9>�ǅǃ��d�'���P�U�<I�@��k���(�)R/&�4��fjH�'!�$j�%!!�u���	u��-c\,,ZJ�+�� 
Ʃ�n�*�"�%B�#����2O��=�c��5R u� ��X���kPB?�"�C�1�����g'}��b`��5'��-�9�C�i�j���+*�Jq��������'ے ��E��,�@�
R�.f�����yb�[/e�望v���,Y��	j�v53�W?�Ó��$}zf)R 8H!�7��ѐe�=BTxY#�kL!r��Ԉ��+��s��7F���I�6 }�g�� V9���"=��5��g�i���4��s+ϳE��v�����6�ӒqY�T����7;�8���Whl^�0�eI �Ls��΂na{r�íiA<=�!Q�o4��Yr����$Σ�v03�B�z7前�M��� �d�'^���,T�,"b�h��	l�mK	��l,��c���+q� ��5&`��b��(N��BG�>m�N/x��r�U�*v剄_.��զ�?��!h�? <�hq(�.8IVa�#�@d�-�q�R�Fp�:<�	0�Y�j�.��r �MDrp7B� ��m�Fljy2@]1Pr��L��K�" ?��+�?����e�>���*=����f�<��C�y��b>B7���w\U��/��&�x)���u�eC� ��欇�	S��aC�"F&U2D`_p$0�'�j$��B���T�O�P�@�Ń4#f���)A��C3��/����m@�"���$Y�;7�ǥrw:�#�n���#���+IhtG���3gD�(U��$������#��o]*���F҄'#9�!�ɝ�na�"	�5��O���]��, �`�
���y��Y� �TmjZq�&T�уEz��ʓ'�x��`����S�O���AeΕ'�n�h%+�(���b
�'��}���%7Z�$�3GP>T�4i�	�'��Y ��h���:�b��T���A�'��H'j�
~��@�� �;Ĕ��'e� �tO�$6���c��+;�"�'�X3�����P�"������
�'����f�	t�)�oP��;"O�-I�.G�n�JA*_�a-����"OZ͡%D��uDpd8d,��;>b3"O9��ϋ$���p��I�~�`QST"O^1����oL�J lXPNŀ"O0�HPHF����"���0}�hI�P"OJ���왂DXg��Y�*�`�"O\�hrHʷ�V$a�
��Ƽ@U"Ob��2*J�20<����j�
]�@"O�<p���B�>���ǵ+F�C�'2��s���<�҂V�	��� �'����VM2&��\S��R�J[�?D�� �Q�X�������2���B0>D�pQ�oI#+'^,���	wm+Z�!���)|.�p��$�,���96l�T�!�dJ"�8��4 ��a�"e`˛�L�!��=f1�BTvw�M�IK��!�®=�L܀5�N2*j��;��6kO!�Mn�y���O`��KWo�Y!�$�"lP�YB��p��r��T�!�d͒X�|���Z�d��PK��	
!�$Z)y��`�1��'}�:��!J�!��U�C��c�NLu��5{��$r�!�D�<r�B@��-:b�99l�?3�!�^
H����'+d�Ej��ƭcq!�DK�0�8l�NY�>W�q�
	�.`!򤓵,,J��w�� 6�)�#��&�!��R؅R�O�µД�W�)��"O����oϖS��Z�膳i#b��"O81+�ʖ}���G�9y � �"Oh̨�"�9��!��B�<�r�"O`�`�uQx���ˇ>��lJ�"O�E�3B�����-T7F�� �"O�m r��)�X@�#�3	��)B�"OԬ����:!,\b�;{,�P�"O��{ Kݲ Ș|�sH�?jԕ�"O�찥'ӅD[^ ңI3e��	j�"O�P��JS(H �l ph���� ɦ"O>�c�/ +`?����D��\hz"O��ç�Z���P��Yb�q��"Ỏ�Gwf�o� !���Qq2C�I{2i"�K�0a�ޭ����Q�B�	�fnq��eP�?xִD�	�B�)� b�"�L�'%��Z�K�Ҭ�j%"O\PK���#Iy���U�(��"O��
Q�|N� ql� x�D�)�"Ol���_<�RPkMSΞ!�g"O8�H5���%aL�e٬Y�&"O��Sq�N���:���<�X�"O��A ƜD� �"�ͥ�z��u"O0`G/Ǐ�x��h�	�~}�0"O��X�o-4���M:��큵"O�}��j��Bپԉ�&Z�`�2�"O��i��$���Ya�ʼ�����"O�q����%LȌxx��V'�8�""OXY:$h�*d/��0�a���i%"O��)�l��m80 g�F9�xԁ�"O�=��ƺ�8�ŧ[��`z�"OQ���[*�D�у��
;�yD"O��׌O���9�!�6!�9�e"OĈ��͗0Pq)瀚�Gv�� v"OΨ��A�H�����CU~�P$"O��9��
����*&MD�;B*�"O
L�v/�6O���ΤVRhp�0"OZ�d�ʉ$�$�!�S1@dxy#"O���"�ʤx�2�,�.FV�lp"O�5����u����X�=EH�x"OP9B�ˀS���󧬖"2�M� "O�9�!�H�� h+&*Ħ77�Qi "O�[EN���Y�k��2 s&"Ol%	�R%Z�tej��"8���"O���#�I�y��T�Μ<u�� �"O�25��?>�%���=��)p"O��� X6َ�"D%�����"O�=�cI�7��	���U1�4���"O`�3#N4W��=d �8<����""OXEX�J��$M`m�n�9hvBip�"O>yaA�	�~=��4uS�T@'"O�ya7l�1K���K�_*���4"On-�Кz�����A?j���"O�=�aϑ�$�B��Z&ʄL)�"Oƴ���F�����o�S�H	�"OtE��lڰ]2�2%��P"c"O���4�.,����1���a�"Oj �`�v���1`(Q�f��!"O�}��A�&C�p=C2�̙&�m�'"O��V"@�QyD0{e�
�La�-�"O�apd!6w�Z2HK�{�M�%"Oz�3r+��L`$��&�S�9��C"O�ᓂ.��">-�.G8~h.�	`"O�89"	�K�����΍�)F�MR"O%r����u!(9�bG/F��yC"OHQ;��%���iQ,	�"鮉�3"O:!��߲W��9`嬙�|���"O���D�h�|�t*�dR|��"OFݫ�թAߴ��U�kYf��"O"�pF��G�FB�E	�s`��Q"O�����мh	>����Pr!��"O$Mp��P4�@:cDQ2Q~(ղ�"Oj�ee�5*Oԛ�-�)~�	+"O���s�%HA�UhEf��]]��A�'\��aHȦ��c�2@�~��8,p��%�;D���LZ�P�����-=�n8ғ[�JCv����(�D��&� z���T**N��
��'���
���h妚�U�t��韻5�t�eVl��`�!�6=��ӧ��D�/K�\���L�m�>qKPj�HO��!򮈖'L��|ʅ@,JmH$�Fއ HxeF�H[?y��"0�*$p�k3LO� �5��g� t�d���'��!
3y90�Z��S�'	K:  �Õ2e1�P��!�tިer��	b��#B$D�X* �ɤa[��sv�Ҁ$}.�{G����R���<�S�]�8%h$�1-G��S��Pƨq�fZ"=��A�Q�p>1p��AT��Cԑ[���`�h����$�L��ܳi>i�FM<����O�IwN��4Qau��J@��y���%��ys�M>	>��΁�O�  ����,+d��a��t�fɆY�r9A��OX��Rs.�-*���
���=�R̚��)4��²�(>�ҧ�O%Ʊ�Eg��Uf�T��>�f!Z��=(R,�c
(Cw!�DH���z���q�Ή���!���ղ[Ԑ�k�9��yu�T H|D�M)?�O<NT��E�'W"��c獪
���3�7� ��/�bp�a��'p�U��#(�d�������l:�	P���$�J�"~��
A� �2����� �HOѣ���%מ���ɑ6v(CV�]���}8ŭ��c��ɑt�V��WᕶHayB���>֨����V�� 	���)�?ɰ�8Mf�DY��*}���ٲPy�m���E8S-4(��Rb�Ha�u��FR\��ēc���9���Fʪ%�����jp��'45�V�[[M��m��c���x��b�i>����.,Pd�#1���zP��#�O~D���Xfpi��ܦZs*��f�=��]���'�?��Oc4➢}��$�1�T(� �^{u�PJ��s�'̦(���9,��~*'�ҝ|x�ZG��><4$¡Cn�<�AL��r��96 @CW�V������ rzp�s�>E�T(��a͚1xP �h�d11��"k�!��7�|ؤ�Ϊ<%����֒3��I�T}@d�s,�mx�d���^������V�m}4L�h?�O8 ʷmX�Z�xp�	�T�d����=���	�'�f!��!����-Àypj@X	�'SȌ�S�O�oM�����9K��h�'��9��6}d(=1ga�O",�3�'�ʜ�E�,��͢�ȑ�_��$��'*��1�k��o��i��lٺK!����'J�I�u+וG�~ "�E9� �`�'�^Ⱥa�,h"�����$���'�T�p���9i�H��ő'������	������S�O.P��efN=�d	 u/I�_�.�"O�=�d�'!Q��
pۨ[�I��R��bei�L͂V�'�D�P)q���aL�Y��1v��Ϻ!W�\�GDΛ4��JF� �LzK���x�n[^�.�ta�7߮�;�b£�(O",
w.�	[�:Ř4!-��9��Aa�.S�/-�h;"mN��lB�	0i����NŤT�0�1i��{�T �ƁZ�O�L|���J����O�1�G@@���iB��fE@R "O�,���V�NLR�A-:]9���O�aZ2�F��p���9,O�ѵ�B?BubȚ�E9x3��yS�'����rfL.n`1!�Q�c�6gż.����ț�P�!�$Լ]�~��")	#l��8 �O�{Q���!U�X�j��B��c�,d�)�S6Iđ��
"���M��k!I�D�� m� -�U�tL���|���+��)��`���1�نCR��j��R�?D�tY2��E�VX��4g@�稸>�����#� �ɤ%o8�_��Z2�ͿL
D��Gӿ{����3�O���S�$1� ��
�8�L�D��3DX	��c1�IW���pD�s�OD�`������4$��
�'�
��lM�
"P�{e� �V}I�Oй��\�H�����<q��_M$�v�^+!�nu`/AS�<�D#�7q�
���	 7�,9 �ԌH6
eS���<d/���I=[7M[cF�#u��Tr���j$D��ݱ=�� �dZ�R/
�]�>�(	�d�B���Ԇ�yB�-aނ9�3�R.�h K�(Ƹ'6���u!�
�1n��>��@���Lط�)W�P��j.D�$ -���ʂ@�7 ��Q��ް&<�2 ����D��(��	� F�Y�G�<�x���L�#��C�ɴ1��A�ƽ2$,il؂��L�@#B�p�K������=���V� �$U�1>���dXH���p��@�tI�̄��M� ��YF�.R������u�(���"O�	�PI?/dp�rdR"#��EX�yb$# ��u8������G��ܝ$�E�'ā�'�: �sa���y"�:Iݺ��Tʀ�ޖ���?U����5�B��/s�����L��1�fɮ�@T`�n��Z�-)?���&���?%��Y�	вa�+�
�myM��|-�e���Z3�n���'�Й*�Y�6�iY#C�"w䠩H>Is� �t괹(O>�X����i��T#�A,M�4Myv��+ֈ�!�O�%��n(
�����/J���z�I^18�0��	�������O���� @�O]`�G��cÀ��\'ۓb,��X���O 8���>ӊ{I~��21f��!gF-C`T����$0�S&�[yr�
�K9��f�h ���2B��9w52%�'�ִ�e(T�5����OQ>m��ǒ0���Q�ڹQ!n��GE,h�r01�A ����/�\�J'�G�%?䡙��.JzY�Ov��#T�Y�8��O���g&)b�2u��J̋6/�C���C���-`)��I�&$���̣ES������cH�ܚWo( 6�b��`��^0Qh�%���^DI$M�{�dsQ�FT���@�ɢk���WH��O��4#0��4���y D�"�`���'K��b���dp�R(*��5�+Ohh��!��Z�(�OQ>AԭR�j��eF�OC�$��1�,D�p1�q���Ã�&1^d�t�!D�|�G�Ϯ%�¤��E��kgF?D����F�V���:	��a~���F<D�X�QOZ�l�=�V,�Q��əbj(D���1�G���Hp����F��O0D��
��@�a2�a���2f��Bd�,D�D��K�}�*�؇'S&r���(D��8�e���nk�S(i�䍡m)D�4���.ΦI��c3��z��)D���1-X�a[  I�J�-u��S$D�t�檚
��h4
���C�
!D�ԡg���Y��FSf	�!=D�����̏n���{Q���|���C�=D�dK���<�6��c�7l-HX1s@:D���d�FΤ�!sMͪ*�V�[b�9D��BA�ʂ|b���ą�#}��r�(D����*Q4B}8&��O��L��)D����
�J���p�6/��Bb%D��9�9g���`�W�JC\Yb�.D�h9�-T��.HK���!��QS),D��@�bI�v�9!�[�w��#�
(D���m�q�����D�o�EXe�$D�\R�L/}��A�BF@ ���"� D���D�+����b�|n�qF+D���m��rrB��h�5��(D��!c�!VX"�^���!�-D��0�eH�8[z��qʗ�M�Й��<D��h�f� M�4�ޥwG���CM>D�`�A�1=	d􋁭F� ��	X� 6D��K�/Rj�B!	�놓(x� Y�8D����ݚm~�@�HI{�͓d9D�TX��&�
�I7S.��i�J8D��'���o���:���LC�,D��0� ]�Npq�L$��,�2�+D� c-��C�`�^TQ�:��*D����*�7.~4zu�ܲE �QB�,&D��2%���>�]0Vd]pz���mj�t��NQdKȹxW�"Ը�J�K�<)���#�~T�
�q�	�C�ɬtĉ�o��jdq8J�<�+��4���`�O�X�Bׁ�9�(��%��.=�@ʎ���\����X�?�5�������@Ƚi�1O�Ez��DC�"E�:�Z� 
�8�{T����AT���j	�E�Rv�8��ЫG�D�8OR@"u�̓Y��r�!}���ӢGiZ\���M���҂�n�[̓
�ްC�i1?E��-_�	�zP�7�	C[t��g��*�y"�G~R��ey��� �t	����)�q0����B�|=P��p>H�DzR�dA�oZ&��� 	�U���� T%�`�=q览��ҭw�<	K5��9f�٩��#I!��H0��́検IH�M����&!�dïC錍��++��{łQ�vB�I�f��xP'�/�J� Qk
V��O���6\O<!��H�~�ipp 
���A�"O�#�C	�/ݘ!��v���'�qO2���`�Pƾ�WC��
��]���=���?y��I kX����6��Bh1+v�޴x��	1)�T˱ҟ��~R�'�
�%�/?.t,i>��hH<Q���|�Oq��]��;x4H� �G���&�9�ʾ>�Q�D8>���=��p��6I]2j-�P)dI%3��Q/W<j��!�޴*d�(��D�0:���IǍOԎ����0$p2�#�b�v���4ҼY6�ĀN�t��B�=��iJ=<!���é�a눈�v���U/�)�r]{pN�:*�S�O�L���J� ׬ �"���:wo�$*��  `�J�P.`��M.�0|aGG# *ThFL�"����s�F���(� 
��	 � �t�g�I$W���2dkHsm	����qxC��~g��X$g		�0�5U0P<HC�	�u��b���W�ԓ�i��e�C�I6x�B�xUlъ׌��di̦_�B�I m�����@�:ZX��d�H�TB�ɉO�8�r�;]q6`���[6}��C��f�M��̆	M:9�3O7N�C�31�>��C� K.5��>L��B��"K��a�đ?�*��wƜ�eêB�ɐ'F����"S�?o�(�GM���B�	���Y��ֻ44l��� ԆC�I�C,��7�J�L��H�<x�a�ȓ��@֏F�v�H2�O /����2; �Ȧ��8t���6DڗQ��t�ȓ3�4��&M�vmP�/��f�!�ȓ���p�MH�\�������A ����K��uYP�X���1K��<�ܴ�ȓ�<�b�+5@Z��p�,���6f�d�Tk�S�Lu�D+�$�^���s�Ɓ��c���)J�5�zU��Y�]KteD� �d+�ϒ)nr���y���g�]�Q�SfL(�4����҄x��5Gڶu��bE`a�Ѕ�Q*F��h`��yz�p�RŅȓ;�	A�Eӆ*��Cw,��#Wށ��q��|I���V\`��tb�	W�8���n�h�D��'�30�C�$�م�eP��s�^RAg�<u΄\�ȓK��K@� Q�3�U�3.N@��`�ݒ�B)}Px���E�`U��Y��C�&M�T&4�#� 4G�"��ci��4N��N4F ���ˈA��-�ȓv��1��S��AbT�Y�M7����x�4���	"���0]�E�ȓJT��V$��y��D�T�� ��)u�y[AkO5{���c���(�ȓ+�ԕjRF�-VAJ�Fg��w���ȓ8�~�٠C�'R=��H�ʔ	E�لȓ_x��Wn�90���~�q�ȓ-GH���b�}
���`��X�l��%L��^�|ͩu)C�OC���ȓe,���𤍃#��b�J�	��Є�2@���e�"B��ЏT1��-�ȓ	$��RސX>Zu��g�9-C汇�[�l̳�C]kre�`��?���ȓ��U��fѾ'l�C�T`h�ȓ%��\��m�{�Fl��N�p*����S�? 
m� E]$!���) F
�?�Y�G"O������r�rD��E�����g"Oj��s��r��b��;?Gn\�q"OF�AD!u�,b���{-�a�"O*1�b\'u9$=��%w6*Q*�"O��Q'o�Y��(pWHƲy/��"O�x���כv��Q��� ��1"O�U��#@1J��q��ЇO(p�F"OR�Y����TL@"�揄+�H�V"OPԡ"��&��'�u`�Td"ON�ڕD5�Y@ 06:f|x�"On�K���b��*��a�Z��a"OZ�Zǣ�=U��t����#�* {�"OX����	�,��$[,-�D��"O��£ݣO�P�c*=.c�X�T"Oty�Vc�[��%���N�xG��T"O�1(@oȟF������I.<p=�R"O�+����t��%�.F"z�KE"OK�g��4Z�
��#� ���y��̥[)H���"�� ���y�#ڰN��f�Bļ�m��yҧڍp��ʧE���L�R֢	��yl��w�4�u����Qb5�_*�y�CD�nQX���N�y���M�y�aS�fg�\�4�"}�j��y'A�kTD��كW%l%���R��y"gK�Z�#s�W�K�E8ABD�y"�]�z��z��X�Ou���L6�y�i[���d ���Bi�bN��y���z@�9b�ؙ^�f���y����#�z��e&�}k�	�rfL5�y��"GvI�E�֐sfCc�-�y�b
;L�Ak$�ѥ�D���Ž�y���C� �ۖ흭B�I�W#�yR�!R�Z�Zd=#�Dx�д�y2H��^�H�AӋ�>!Y0����ߺ�y�F�f�
�kg��z
a�E���y�%U��uS�!WBE�R��y��ݼB�,)�v�|2����7�y2��*Q�x[0� qW茢��U��yi�Wr���%�m��0����y�"������Ӯla�=ȥ�B�yr��h��4��-�c.�D22Ό4�y�gދ\�T��`ڒS��R�Ά�yRGPs#�IQ���_��0kqE�8�yi�"�؉�ER�QB�G7�y����/G�ě! ȴC� X���P5�y��h�\#��αm�J�P��y�O_4,f!�C�da�MH `
�yB�S�U[P��&b� !!a��yrJ��{����AFF�T��	S�l���y�&��s#�-����N�~%�t��y�`�6���Ä	�G9
����ď�y��Q��Ec�%�$:��m�)
��y�@[��8�@ˑ�7����c��y���/pNᴪI�C&PQ"�.�y��oJ�P�O�;�D5��ң�y��>f��06�Ĵ<�J�X�ͼ�y�o��n|��;Fl �,�a�)�y"�J�h"jy31��M��Jх�)�y��G�qS*D�'*��Z=�(@G��y"���dP`�,]�Y*V-)�g��y	D�]���֬�#P�n��GO���y��;���P��M�������y
� ���KU3L��R���
5��{�"O��hg�N�|����P ���"O�0�P&�G[��H��$e�"O�PJ>��ݫc������
w"O2�q�)Mp�䈂��^�B�0و "O�]؅ �U��b1k��z&���"Ol���Z6G��jAd^0!th��5"OF����?fT �u��T�����"O�a��@ޘW>h
�bĹ`A�ܨ"OV�`7�\i���� V���"Oؠ�5��p\�p���O#���"OV`4S�I��S���G�� c"Of��'� +��I�c�#g�0�k$"OlU�Ìdʢ-q�'Yk��8�"O�,�� !@D�U���;S���#�"O:��A�㌉�sj��l9&�Zt"O�r�5�Xp;բϧB��h�"O�Q��ĀT0�dO]���`�"O"�S�@%KQ,qy�/وN����"OP�٥��(ot1��O�7@J�"O��X��HI^����N�!��@ "O�x�d��K�h,9rK��4�S�"O�lCD��R����.Uy�"OI��b֊�-!������"OV��K)��,�!�B�3N����"O|a���  �6 Hӣ^�;�@  "O�Pj�Ě����Ȯ=�r�ؐ"O����ظ	&-J���9z��x�R"O����qˬa�I�<�Xt b"O�*�E7G4X��P"̶:���K�"O�Eh��~#�!s���D���z"O^E	Q�u�!ʐi�������"Ou���F��<���i�V��e"O��� R|o�u�a��M�ҡZ�"OD)c�]iX9� ���$;�"O���qe��I�y1�(M	&ΠaH"Oİ��F��6�&𨠇�B���&"O~�bF��
8B�b�Fϔӆ`�V"OҰ`E��b��|@�@/^��I1"O��ɧdy��7DNC��J�"O�QQ��fm8�##hψ�z�"Oj�Җ�J�Z��%��b"X�E(v"O��9��4X�D�a���&;?�Iq"O�uy�&� 8��M��!>A��`;%"Oxxx��]>i����M�"r�J<�W"OlJ�ԣ
D�)��.p�"Ov���w��:�,~Kb)�"Ov����Շf�,��@k�G��"O�Eа��L��A���2+
�Z3"O�x��ąw�j���&�6�jR�"OX�HP�_o��\�P�A�p���"O��c�#��s�:��*�1P�!�'"O�caȌ�o}�9j!
�%��`�"O���܉XĠ��#Hܥ���*""O���rk&_)��8%���n����"OX�� �0~ˎ�����/k�t�"O�(c��J?S�|09�cR�P�� ;D"O�yЁ
_��,�HC��`����"OBͳ��:=���{�	�:}jm1R"O�a����g�0TJ �Z͸��"O�� ���ݻ7o3^и�+�"O�d��晆	E��K4�P�S�8D�F"O��ӥ�?O1��*e�+@���K"O2�1��.q�Nd��Q8��к�"O� 
�CE��|�h]�Cm��/�v��C"O���@M\�r����KM�
FE!�"Ot���
�,���!�H�lNx+�"O�HA��V�O޼�[@�ƖQ�x�{P"O^e{��M1��$�`M�J�@ ��"OVP���"l�qӀ�]���j#"Oh��C��5"d���݂�0P�"OVH�m�*��ztA���*�"O�L!"�� Y���pa<�YӢ"O��I���Zm@D���ۅc�b4�d"O��o��M��&f�%y�t@Rb"O�\7ݕ)!��P��\�k�xA�*O�혅(_�0�:_r�<�
�'ޘ��iD�Tb�=�H-8Ƞ�
�'ŀE��Α�D�B<�vGO�N��i	�'��L�a�͢a܍qE��0U��J�'�B��@+�hxJ�fP�38�e@�'�]��b�Rb4#�%=�9�'6�e�uC�-��x�cA98�h��'�N( ��3w,��H��T)ڰ�H�'�`y���'=,��A��?$�di�'B��F�҈�&-�1L�Ԥ(��'�<�  ���     �  B    �*  E6  'B  �M  sY  %e  �n  ux   �  Y�  D�  x�  �  J�  ��  ָ  A�  ��  �  c�  ��  �  E�  ��  ��  �  \�  � � X  �" ;+ �1 }: qB `J �P �V �Z  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p���hO�>U2��F1C4ӡ%B�>��eW�%D�����9]����"8�
mS�#D�th���*��6��4��$#D�\��2~F��u
�!.���sA D����ýe������[�<�����?D�@�w%��&�f�SS%D��8a!�(D�HY&N�1V�ȥ���V&D�A�`!�	�#��yr�C>s|D劥o^2;#y�Qk��Px�K�{�T�:���(8��+�#$����>iS�'lO�m���KTѐsF�W�ճ��'�铤�$ũN���rć:5�@3"��)rm!�P-s�h3eH�r�xb⪙�j�!�䈾�Bl�*ݎzp��a2c�1Y�!��8$�N9�%�D#f?��
�#��y�!�$R*l���2�Ɵ�1���8cǈV!���+ D�
�dV�e"⼐Fip!�$�8p�,�7�֐:$��`H�;�!��vM��­�@�0��/Et!�ĚYゼY@!҃&���K�f��l�!�� ,.�T�%rd$�4�]<~!�䛱���kah�f\삑�M<+`!���8�e��2G,%s�FS�gI!�� ~��d�)b4��ci��.�2�"O�a�L�I��=@Dg�0��TP"O�1���F�nؘA�5^�
���*O��(�NB4)�xt�θNy�:	��Ms�O�ݒ��hҊ�Q Ў!�ZM�"O�������@K�ux6Q���{�O˦�l�+E�x�Q�đ2 Na�	�'٬D9e��91��p�X$>��a��'�б�Q����i�&D ;? $��'͢\"�b�^�@!`�A70uش�~"�Pc8�@SD�?(31���T�j	���?\OB���$�`s8�Xt�����I�f�!�D_�)��#��R8�$=[���F��'Mў�>]@EÜ� ��9z#Ï1�̐ .?D�X�h�%;��hK�ɚk���F D�*$J�)" � I�3*�q'�9D�L��l�K�d<�7�1<�5xү3D��q3O��%pafӀ)R��p�/D���f��J������Ib"���-D�L� R.أ#�	�D�*u�7@+D��8R&R�2���B*^,�Tk�k5D���3
L0�,��f�1(��xC��t��=E�ܴe����Q�0�Z�(�N˖|���ȓ[��}(�h�0"��_�Y �0��j��s&�O @�B�I���@p�P���F~���`F��%�^�7��H�ӳ�y��9P�����:Dql9�F���y��N�'�4[�IE�%ߘ��E�̥�y" h�^�ڇ��5�-�'�yR	 ����P�S?`*y�����ySc8P�{��`���'��y"�U�S$�R�$b��z�K&�y��X�rm��"��\}&�I� +�y�)>1��E���O�H���؟Ǹ'�ў���a"QF�D�A$���;�"O����7��<�2��5c,dts�~����BAH�8�YPg�rhR����y�$�ޘcF�U�n���^��?qQ)=�ONa����ph6��F좱pe"O�e�/���Ukֶc�I��"O���茰+�j|����vp�d4�S��z��X�W {E4�(�&�DhC��2z��iH4�l%��7|�\C�	l��2�利@��MR���z'HC�I�)r�(z���$㠝c��+�FC�	�L��<�����Wl-s�D�$2C�I�]��%��� �X!�BE��ybgH�(�L�g�� �&�Prm����d*�S�O�<��� ({��Ar&�T
#��t`
�'�<M2�g��h5�����	�'�0`!�(��&��`ժ���� 	�'%���7�L�RE�Q$FB��"�'��h�Wl�B��	�qO�+K��ea�'O��Ȱ�H�j"�y��W�>��z���'*fՉ�Q*y������gӄq�'6Ȍa��5��Y2nϤTTh�8��Dp�ޣ}�qb��T�6(��Ob��u.P^�<a!��Vp��ᨕIF��S�GbK$P��O?��B��*h�w�ۿm U�6(Y!�\s����?s��!��$�����>��M�+�����*@�Rm�#�e�<�b�5q�������1�|0'"O4t�2�մer2�/�(i���"O������<4}B���M��!C����2<O� ʅ���^#7
��bQ��];bOx�����&PP�,[��=��( �� $���`8��2����7Z�����>+��;W�=�O��A�'^�}��(�d�X7��<wR�52��HO���&��&X+�c"�r��$I�"OJ��`S�l�1O�
���W<O��=E�t�܉k�Z(ˉX��0Bd	�:�y�: +d��)ɰ\�`�� )T���Cݟ̇���	7G�I�<}���������<IR.��h1����%"�&���n�p�<�u��0Am���4�D�e���yĊ�e�<�W�J�I%�a���
BRV�١AF_�<aTE�TԤ)���=0�U!7�x�F{��逯L`�!#$�˯[�&e��	�"|�B�	j��e��޳�-SET��ɧI��I��~��hO����Ǆ�$L�rs�<8oڅX�'�d��'�4��b�d0Q.Y�f��n�W������m� `�z�nZydN�V��0=A7�%��$o��<Rŕ�,��K�肍M��듚p?���	c����e�E�mhb`а��}X�ԦO�<q��ѷa�pz�X�L���"O<p��C�	R���y�-*g�|B�'��O�c���Tyƚ����Z4�����0D�x#� ��@�:��������d1D��!�[����g��r%p%��/D�� ����7x���ʕ3Y����&-�	��Q��O��좷��'>i�`��o"��	�'
�A4i_�f�\ѓiD�3L�ّ�A,ʓ�h�����t��|f)*>z���t+�m�!�:�1gI�>} e����)�Op��r옺i��h�&ԠXw
"O�p�A/EJ��E&��Wg�-i"O8���R A�	&e��d?N$	0"O��C	qȜ8p�!1`�V"OlUAR �;I����.	�(h��"O6�$�ܻZqd8S4�L(��e�F"Oڥ"`��?bH����t�(5�s"Oй�&ǝ5n$�`vkA�"O2�Q�!�Z�|�o>1���"O� �r�E�1ಸ��͔�/�1�"O`,b�m؜��H�&��8�`��|M��jȞU�ƍ���Ǿ^o�8�ȓRBL�j��@>A>qKv�N�pńȓP�0Z��E�
C�s��!9����ȓ�Tڰ�š<����s�T7R���ȓ-ъ�J0�O,B4^�#�a0|�ڴ�ȓ5� �+�!;ЌS0e��Smf���G�\���
U���dO��&�h%�ȓS�Pe�4DTJ�Ve����*p��m�ȓa@�����[��q��G)�,��ȓSIl��+m{B�ѳ���H
�ԇȓm*�U�#�>;�`p��S�y(�������Q@M��}��-S%ƻ'*Ra�ȓt8����������P�>� ����@�A�A�7#O�S7D��+	���JR᳢G@q`�[��\B��ȓR��;�n�iP��J�:{ņ�?x$I�6	E���L�ES�2.���ȓk�`��3Oĉ�7G�p�4Q�ȓlA���Mլ9�ɳB���$4l��l�*��T B�Rf�P�̇+D�$Ņȓ[z�akFk�7tv��C޲C4|�ȓZ��5��^;d��;A��+��|�ȓ���G��%Lժ���[vhɅ�S�? ,�T��5M�<���"8=�"O���Aٓ8.�ᡧ�7B ���"O�%�X�F�+��B�/�F"O�T� �/f��\u`�89��Q"O��(q��uJ~�	6k��&���0�'�B�'U��'�R�'�b�'���'arP�$@�[��9�,�95����'C��''�'�2�'NB�'���'��lX7F����ȣ��ͷn��H��'+��'���'�R�'���'���'�ik��4+*��'C�|/8DF�'���'���'�r�'���'%��'�t��I��[���LV�+-�?A���?q��?q��?!��?y���?q��ؽ�����K�MX�O'�?Q���?����?����?����?)��?���N���p$̂�s�:��D���?����?����?����?����?q���?�B��*�~�i��Z+Z�Ő�����?9��?A��?����?9���?!���?�S�F�)�d9�C�ab��A�����?����?q��?���?1���?���?�0E��g��A�Q]0,-p̙q�� �?9���?����?A���?��?���?��!3,KHI�4��/M.������4�?9���?	��?���?A��?���?I��=�X���R�;rr�$E���?y���?a���?q��?����?����?	P��)n��LS�ĕ5>F���6)E��?���?9��?A��?���aG�6�'n�x.�3��|��p��@�-8���?�*O1����M[���L��0� �1Q�\���ɇ�9���'�f7�?�i>��̟<Br�K?a]����):Yb�1W&����KD��lZe~B>����V���b�Xe��)K�u^�K$J�"m�1O\�d�<i��	D	������U?
����AY q4�m��"��b����׻�y���"m�@y�ȟ�>����J`���'���>�|���	�M#�'�F 2d��,$�UCF�������'*�d���Q�i>q���]�\d��"r�V��ѡ�>���uy�|®x������ɹ)GL����n����@�'(ڞ���O����O��	h}�h(g�8���ƳIyƀcf������OX�"�V�J�1�X�*�J��䅷'XD�GL�Z�����ƩN�\ʓ����O?��[���kA��} X�Dm�5e�	��M÷�ED~�Dqӂ��+|z �G(��P�H�T	A��	������8pr��Ϧe�'��) �?����U,��D8���3���@��c��'��)�3��g5`�1M�:�PH�C$ݸj��{3����t�b�'���)E�q1�$� _�w�i�,֥A�8��'��7mަͲL<�|BQ�D�Gr��YC�J�!�L��a�w�-�4'����^�)X�1�~TԒOP�=�����&W5�0���Ŋn�L��I��M��&��?��g�Eٰd�į�0h��(s GW��?�U�i��Oe�'�2�i6�6�Gh�9Y2�4"�^�{���0'4<p��ޓ%w�I(�ND1�؟ʒ����ħa-d�;��#�d�p�"�d6�O⁉�"�?���)٬S�Ҥn��O0���O��oZ,���'5��6�|��8coZ��DK��?�x�	�� �'N������Vi���O뎑�-Zν�g^�S�x !���������'�P�'��OX�⁊�0MB����"|��� �I��M����?���?	*��tۦ#-\�����=L���W��<��Ox��O��O��(��HÖ`H���5q�4�����F��4�Ty�OJ����,k����L'zL����oJ|���?���?q�Ş��dL˦I@GE��\b�ͫ2�,�V��g��"V�����$ ۴��'<�����i�T�!Gܟhm<L�J�-;�6J��q�����S��+�0��0n�Q/O�!���E"Z�P8��6[Qe��5OTʓ�?i��?q��?i���򩒫a���-L&������o4������E��h��X�I۟H&?}���M�;yKX�izf�����Xh�*��Mk%�i�jO1���z6��-P�dY��a���[��m3�i�&s]贘�'��'q��{y�!ɺ.�3F��3*�P *��0<��i��y3��'�r�'�\0z� 	S]� ��
�Jm���Pf}�'=2�|ҫ�Y�R�{��5%�$ZQJ�(��D�=Kk^���@�4QvꓟH���'��K����Q�R�+R���B�R�'���'`���P��ͱN�j�p�c�l���bt P����4#Ｈ���?�f�i�rT���i�@a�'g
�`�̌/lu��a�xy޴d-�v){�5�p Y 
��$�Ope;�%_0�����H���c��:/���b⃑3�'��E�',�!�ǅ_5c�h8�L:i<];�O�m>Y�n��I˟T��n����ͺ �N�L|���p�@`��q[���۴��6�!��)˃7�xQ;���}�M�酮qV�;��U�c^��b��o���'�Ȕ'̘I��V�8��Z/;���6�'\R�'�"���P�8��4�t���lP,�8��x{JxٲJW;Ba"u���<|���	P}��'d2Mj�� ����j��)6��K�����c�`��&��ԡ'+\e������� X��E��*R]v!q�̰&b&�A�3Oz��D�h5�2��P1ͼ$asd�9y+����O�D�æ�RJ%���id�'�:Uj\;w�@���$�B�qUm1�$g����O/�4�A��.�i���b��K�m3$��g)H��Tˤ@�<x���ҭ�����O���O���ϫ\��yf�!c��A�b�צ��O�ʓD�6��z��	���OZZ�O��]u:I�S�A��=�O���'�ºi�ВO�4�O�*�{��ӑ	m����a�6� ���ҭ����&���d��0t9��?�6�O�����Jk�������P)\�?I��?���?�|�*O��oڇ�H�qq%^�s�h�2���($<{��Dٟ<��!�M�"ˬ<q�4?�A�G* 0<���pg7�*�;S�i�L7͇�cp2�م?O��䞩, ����'_���"}4t��b�:l�+3�ԲX��Gy��'�B�'S�'�B^>źF7.6�� ��X� ���ߢ�M��!��?����?�M~��zΛ�w��(K$��#Q�*8a��9Z�����O86��E�)�IQ�2���;O21$䛅c4H��v��a��;O�Y�U:�?��`(��<���?��G["��a�єQW���[0�?���?����D ٦�2`@j���ʟ�أҡNF���a���L��I%C�O�)���џ��Ip�������x*�]��X�R��k�,�w-�1u$���|�f���	��|�jd�˙��h��U
p������|�IܟD��{�O�"�Y�C�f���ȋV
�-xFݮv��n�Vt��*�O��������?�;(������+i�1���5V�����?9�4;��bÛqyą��O>��A׬�"�/�t��l)�Fюp>����<9��$�<�,O��O����Of��O�$�IVO.�.�.�R��F�k$6ʓV��v��9$4��'Cҙ���'�f�1g���B��yc@G��q ����>I��?�#�x���IM�tF��R�G��EJ��7�D�o�4p�&�-��T�z9��A��Y���O��'jr	ZƢ�Y� א�q����'�R�'D��T[��Y�4L]���"��)�����3��@
2	��`��*�f4�F�$B}�'��'ܙ�EO*|Ű�:���z�-�Ыݑr���=O��d
�M$���Q��I�?��4����X�3R�eڶ�?7���ܟ��I��t�	ڟ@�Iu��?�0i;6�"����ߨ]$%���?��]�6C5���'Y�7!�����X��ήs���ˀ�Ԙ=SR�$�|�ߴ5`�F�O���6�i����OV���o� ю���˙Xƚp��MD�`��M�>�O���?y���?��Bh\�U"]&D�����Z�HM����?�,OV-lZ�O,I�	�l���?q��ԕ!f�U21�dK�O�3jˆ�X���M��ia�O��� %B�DXa���8���"M�i#�dAb�*x��*���O��yN>��ʞ1`����`�
A���Ù��?���?q���?�|�)O��oZ�BRps�+B8C-�tPcn�'�TT V!��		�M��A�>�^��Xw�U6D�f� ��A4�v�%�6t���t�����x����ʟ("ELǁE�$bgy�E̒_t����ɘ<�\�᲍Y��yRW��	���ڟ@��柨�Ot)�2e��Ib"�c�mC�!L� @����%��O��$�O����$ͦ��i\|���((��ɔ�Y��k�Cz�flm�����|"���"���MK�'z�6�D�G��Y'�P%#�Y�'WL�{T@Jޟ@���|P���	՟���H�	֐�\�8m��J�%��OL�D�O��|���Ә��'��ާ?@�+��
��L�q�@��>=�'�"ű>��iO�6m�I�ɏf��4J1�ސ�U���3<�Y��'��� ��,� ���iw�I�?�K��O|��_�:E@�_<k8��4!�_�����O���O���;��׆�~�|Ur��\K�Z`��,Ԓ�?)v�i�Ȣ!�'�b,jӎ�Oj�4��qe !5��-@ LvhD��9O�nZ��M��ig�=��+���hx����U�0{�́Q��H��a�'s�804%��<I���?!��?��?)�D�
���a�!����J���$�צ�7�̟`�	ɟ���P���'r�h+Gj�23����\�Z�0��r��>���i��7MSf�i>��?U�3��aP<ۀ)�0G�0A�W�thm���$	�����'��'h�I�I����Y�J��J�` ��П��I����i>Q�'�^6��2pr�d�V�L��d�I*� ���O�t��D��=�I`��+��$�Oz�4�tl� dE�!'fa�5 DF�� �I7m`���I�U����џ������gLԅ�4(�?��9���_9�4i��?���?���?����O��0i�A���h�|!R�ؗ?���'�/tӒ��7������'�,�c.�"3fez�KR+9�V�Q�R�I˟���۟�9i�ͦ�Γ���(�.B�i`u#[�L��(�����'��
�O0�Oj˓�?!��?���h��
�ЎyP�a_FLHRFE���	Ey��q��0Ibh�O ���O*�'Q{��3�@�g��:,;On�a�'�f��?�����|*��2�luHc�#.��2�Mض�|$�#[d�4�H�4N�	�?	+��O��O�H��� u+���r�ڋy�JqR��O��d�O����O1��˓-D�6&�I~�q��8||=�!�t?r雤�'�Dp�2���O~��YZ���9�R1n~ k�hܝ
�6�D�O�% &�q�\��SJ�H���Z�� �]�"�!g�-�%�FwF�2 >O"��?i���?����?�����	Ǐjr0��%ϣ2�B)��0��m1����'���$�'Ү6=��Y�2����0��3���O��d>�4�"��ODd:�i�4�<=`:�@ӆ��&&���T�F,{BV�		4��bB�O�Oz˓�?�� �D) ���G��C'�XH����?y���?�.O�im����	��4�I�Ii"LS�D]�q�D�GE�'�j�?YER�L�I�T%�t�ľBȾ�Ssi�p<p�&F=?I��ؾV�� �c�ş_���D�3�?Q5�]��Eh�A7'w��(߯�?���?���?ٍ�	�O~-���J�!�d �%,=[�� re�O�l��;ǆ-��(��4���y�������3�]���O@�y�'��'҄8�½i�I�*%x� �Ob�Q��Y�6"��4��f	��]�	Zy�O;��'NR�'Q¡��(���kh߃d|��bh
�ɮ�M�D���?a���?!L~j�x�JMʔ�<T��$P�'F��F�*�\� ����$��ȟ���*qb����Y�mN&d���Bzll�eŇK���T�H�k�O6�#I>y.Ozl���3)%�a��Ͷ'����O ���O����O�ɠ<�ӹi�����'��hs% D�/@q!j5,Z�3q�';86M ����D�O��d�OẍC��b��h5�ט6#\P��,e	�7�~�P�	,:��A�OϠ�����V�d��1c��p�{1ASP�Q̓�?���?���?����Of�L���=l dy��I���B@�'�'�l6�]c	�S�M�O>��σ8�{�'�(%��@�=���?����?)a/��M3�'���%�T���H8����,�5�-!�iUџ܀�|�Y�����8��韈����BH�-Zt玒LW��H����d��uy��yӄM�L�O��$�ODʧh���!؁[ޤ�aK�xrE�'����?��}����ŝMC�PP�bT%V������%%�^�Y6��3r	QJ��擾f��*\�II*��V�	m�H��Wk�+R��	ߟ$��П��)�Ty�z��5��L�3lM���5D�*0ģ�����O�l��w?�	�\X��S�L�욵�;�8p$i��ܴL��I�4�yr�'�6�s�*��?i �O��A�J�5=B�	"!l$^tQ�;O���?����?Q��?����I�+�L�K�vJY�C�G�T���o���������I\��(����[���A*�@"j�h��Q�Ebɤ�?�� ������'f�t�Q
�v;O�u�3BL)��@��g�,�z�3Or3����?�!�7�Ĭ<�'�?yg��?R��zǇ��$~t���?���?�����ĕ����j�ޟH�I���� O�+g��F�A?$�sĢ @�b��I��H�I=�ē��$�e)�?J����ib��qϓ�?Y�(�>H�l�C�~~��O��M�I<|R䄎#��H�+�uq0K�$��wkR�'��'eB��џh��\�;F\�UO�6d���P��[ğX�ٴcwp�����?y!�iW�O�n�;iB��� �{���C�Q���$v��lz�o��'��aoZ�<���}z@�����䤩P��/<��L�w̒�B��mx��8����4�����O<���O��+d����&���Z��0P���ʓ9��(Ir���'l��	]]����@2 Q��@pLƺu���'���'6ɧ�D�'+���G�H�V �bM��a�L�jQ�u(B�6�����(Վ���i��O��?쀱B�O�h����UL/'`�8��?����?i��|J*O.nZ+r}n���-�T�Ǜ�=�b�D)՛0O6�ɚ�M���e�<���M��i(��r����d�	�aLq���,I��xHi�O� *��G�������wF�pѣkǮ*�.��A�߷/�0���'���'�"�'wb�'��,	�B+@ d#�Y��\:X�U��O�d�O��lZ�I�������ڴ��d�ĨPa��&���Q��G��*�c6�x��o�nz>]� HYB��g�*�(T)��IҼ;���;n�|�$V�Q����1�����8�	 #��җo��\C�u-M�`��#<s�iX��'�'�B�'[��>��MY���u�v}3�G	Z�����	����	T�)".ņY���xDgU�(d6���iC� �l`d�SuVu�(O��H��~�|�lͤ�$��o�"PK���֦�=a���'���'M���V��kٴG�&��T&S?PD@�b��4Ќ@��cR��?��>����|��'Zl듛?ɐf�>}��xz�Z���|j�/X��?ɟ'^����n~Zw<��TݟJ˓l�l9Z�e�8���)��M�i��`����O��$�O�$�O�d�|ZG	�P1n�аh�V�e�I��hқ�"ލ��'������'�F7=����6L�@[�`� D�����O��,�4�����O��!'b��	���Ih�k��tȂݙB�"�F�I�F��C��O��O�˓�?�� L��Ku)���`)e�S
�����?A���?9)OnEo�-���	ɟ��	�c�p)�Ʉ	2�4�Btc@<m����?!f^�p��ٟ�&�����\2[g�ܨ�R!~�X�9�;?�Qe$|<0�4~��O)�p���?��E׌P���K�+`@���ո�?����?���?���	�O0#�*/�q�A�2=����O���	�"8.��OZ�o�T�Ӽ�R�U7�ڽ��
Ë~I��㐣L�<q���?y���t �ݴ�y��'��H
� �?��� V����](f
���G N4�i��J%�d�<ͧ�?����?����?	#����#4$�{��{��ۨ���W��YHr��ʟ@��ß&?E��� ��F�? Z`�R��8�����O|��OV�O�i�O��܊B|hY�Ս >|ui���8
r��!�j��q�'���#�Q?�L>�*O�ij֨�h�4���p�a	�O`���Or�$�O�<�i��Թ��'�*<a�,��dh�J��_�i hR�'��7,�������O�D�Ŧ�A��h�IZ�ϜX�A����4h�d���5?�r��T""�i=��ߑ��T�`�~�3�`�A�gl�����h�I��X�I��d��bK��H��E��O�a��c�����O�n�{����䟀+ش��'���է��L/ic��] <��-�I>a���?��:��#�4�y�ߟ|��0h�
K
5)��ܲh��a0�!�
���	s�IDy��'�R�'5ҎN�A�x��ь\�|�E��r�'��	�MsG+���?����?�*�b}�ec#����)�J�2P��l�O��$�Op�O���O��I04!���q+7TD���.��l�q�e�&e�'��$Oc?�L>�ҌҼ`7>Lz�J ����r�I6�?)��?����?�|�(O�,n�"��v@�;v�$H�C�=H��)"FZ͟0����MH>1� ���&�M�PKai���-��� e�����4"��F���43J��'����8�@�'��D[������&)(�Ń�)��Į<��?A��?q���?1,�&�#$���,)�Jχ��چ'�覡Ѥ){���I�P&?�I��M�;@Ĵ�:5H�8�^��Bզ@������?�K>�|���S��� H���E�+U�x��d�NB��͓_�T�Ců�p&�Е����'�Rqy�"Э(= 8b�䔰k(lzb�'
��'l�P��8޴{��5A��?���~*Ѡ4!]�k��c�J,ۜ��O>9�?��	�Mۦ�i��O�D�)q�Y@��Ks޴����� �M ���a�F�S��B�Dԟ�:$OȓX=��3��ʁ	������쟌��������F���'b�Q*QoV!qPx��Y`���͛	i��~�����C�O������=�?ͻ�(٤�L�\*x���18��$̓�?I���&���'-�Q(�'���cdT��S� *����D��o���3��%O������|rQ���ڟh��̟���ßXi��̪��	��L�;kXr�ۢ�Qy��f�\]ہK�O��D�O����� thyEޗp�@E0#�G>(�0��'м6Ħ��O<ͧ���'&bD��pcU+c��@ACG�zgx��u�ܸ�MK�X��;�)#���8��<��Z.,��q���P��'�ճ�?Y���?!��?�'�������YퟐBf�9}��٣�ۦcd`:����h3޴��'���-���x�J�lZp�ܰ#É��R�P��*�w4nU�HȦ!��?����-<�J��|yR�Oe磇�!�~�G�Q�2��F,��y��'AB�'���'�2�鈕(���CE��,��p+��'<���&���'H47����O@�lZP�I�b���v�ٞ�p5�Ab����)!N>�ٴ?���OE)W�i��D�O����S/#��pVOI���m�,�R���'�'�������ٟ��ɛ5uvh����L^��3oә��������']�6��:t���O���|�剂�:�T:Cjʭ����z~"�<a���M�s�|*���$Đ%RZ	hTh�4�"�0'B6X��Al�B����d��e?QM>�FԣU��4P4 �'3�4t
�M�%�?����?����?�|2*O�Il��q��22GY.xR�@��9���׈�� �I�M3���>� �i�����nX�S�
G(�+��Dئ�S�4v�r)ܴ����*G.�ܱ�O\�	92Z�����jv�M҃��B���	Xy"�'z��'E�'��W>�B��ߩZ��$�U�\�?v��BQ�� �M�T�T��?����?�M~��H��w�L����+�B� ǬS�F���-a�pun�;��S�'m�8�В��<�7��)N)�ᖶqΒ�!�B��<�b���<f�Ik�	^y��'���߾EI̅(�`/ggXI�_#��'-2�'a���M+6lݳ�?���?yd�wq�%�2K�7�R4�R����?a�V���۴�f�"��W�:�ꀀX�y����ED�-��	�@;��SFŬT^�&?�K��'[�1���MQ�T�SD 6���DdB3j�@�	͟��IƟ���e��y����|��`��Ŕ�m�R ���M�xdR�d�bY(���O��	�'�4�iޙ�B�5MB^����h�"=��ey����4Q2�Fz�$`u�r3�	8h8"E�D�O�.\Td�1O��hf��(��c+�W�Iy��'�r�'�2�'EBG��WkH�CC�Q�8S�P��W]剻�M۵΋O~"�'��$��4i\�Ju�`�AÑ�*�|aKA.C{����?������|z���?��J�23��P�ˊ�����q�^:�4��$��`��J�']�'�則Y	��b�)^+:T�yc_.T���	�<��П��i>I�'yR6��8jn4���9�PQe��|�Ԃ׎��R�����Φ$���ɺ����O��$�O��F�΄`  
â`U6q{��%'&� ��CO~¢J�q�'��'i�F�x�m�02X3�Z=�ʜRA�ݸi®y��D'��e��.�$(�};go�:.`|�ز�]3��<��زE��Z>����L�ʹ� A�'m��Q�"Hgx͹5
�0�BTA�$]��di�'4?I�&��&~�mj�(U��jb��I��b#fڡ\�z��@jբ<rxz��/,V�ͪ4+R�~}*���]�����cѷ�� ��!��SH�iħ �>��;��6A��E&ĖPHb�I��}:���"��Opj<�E��*��Qe�G�uPp��t��Z��U�?<���i��'�r��'\������O��	E2�1i&�Z�.�}k���h��c�T⥀�d�ǟ4������'*��m)��&ng���JÏD(@�o�ҟDFHG�����<�����%�[�J��%���� XBD�x}�JB5Q�W���I����_yB�\�u���(��N��\h�ƛ1?@��:*���|y�'w�'j�'�vL8E)ίF�V�V!��1�r%@:\��''��'��]������/���d��i���7(��0�±�F��M(OF��)���OD���q&��������?f�����E����?����?	.O���F�l�T�'����Q���Epqɞ�?�t�6�x�h�$<�D�Oj�D�D� 㞔�լ�+Q�$��2A��8x� ��yӲ��O$ʓ��*�V?Y�Iޟ��S�6�ډX(�+L�i�)+y��YH<)���?�� ͤ��'x��E-,{0A��ɋ"^��pv�B� T��U�taB��M����?I����vS�֘-Crm�P�ׄ_R��W%;Ph6��O���P��p�}�����qB��r'�t�~��tk�����ThH��M����?�����[���'��`%cH�[�*�3Ul��8���b&`�f�3��3�IL�'�?I3�ėI�98cIN�eG`8j�������'c��'%��i�l�>1+OH���,9�-߷dv����ĜGZ�� ��O���v�(���O����O��H�.w��p�Y�=s���I�ht p�O*��?I>�10J�!K0aםa<X�!�hR�1,A�'-Px�@�'�	��H�IƟH�'Ĵ��w ���`�I�M�T��/�{�f���$�OؓO���Ov�9d*��2]��Y�,�{����hÍ���O��$�O�D�<����y4���Z0�ܑH�T�kq��T�[�`��C��ԟd�IM����F�y�$n��l`���-�h���'�r�'�"^�L)7����'}�j��ХQ	&n�hQ�V?CL��3��iPr�|r^�$)P	��������x�)�*{e���h�(>X���i���'���k�r�L|������T���� wu6E�ф�a�L4o�jy��'�r�K>����D��5&kX��h���E�,E3�&��M�/Od�:t�Nɦ�魟�D��<��'�\q��&� ez�O׌>��ߴ��$Ԝ�:��P�f�s�d�#5h��}����`��.-�!�5�ifh�ڣ�~�����Ov����D�'��өA/"��(�;3�^!��˚�f|��4o��� ���?y���?9�'���|�3'D,!��-�.$@@H�{10�ѣ�ih��'� 1{�)rJ��(�	�3H|�m�gJ܏D�n�b�2�'&�1��%��O��d�O8a�7l��1`�h8���u�J  �K˦�ɾ�� �N<�'�?���D��0��}�&����f��>5uvlZ��Xp6��D�����'��Ο|��*O�O��Ȓ�.p@��t��Ж'8��'�Or���O"�j�!{.%����Jn���q���^���E����I�����ey�*�d���JS&-J�%��1m>LI��'F��?a���?9*O����O� �A�O�LzF��uǴ�{��� � �i�� d}��'W�R�x��8i�V��O"̢ Ƹ��eǄ��e��kN�K�7�0�I��ɚG<��`n0�$Ń/p آAE0xД1�@[O}�6�'_�|Q2��-��'�?���Ö�C�ajZ!3�BU�\�(L	��ئy�'�R�'�buy3�'��O�\c8�|�poB�hR$�FŜ7RH��4���9�uv�if�'�?A�'~���:�������Gk$�J%J�("
�7-�O��D�*N��$�q�S�?���M�%�V�Z��
9^~�@(�CY��a9Q�ʞ�M����?I����x��5�jF�>�&�a.�d�s��M;���?���?�+O��g~�OHa�q���W��`ub�Ś�>�7�O<�d�O��c�G�p�i>m�	���'�ޑlW���ql֞���&�U,�Mc��?���(��\?��?��#٪I���]�Ը `�$ .�.��'�i��h��d�O�	�O����<��mݹ<���S��)u,ʹâ�-|6���'D~��f�'s�'^��'r�I.v4>�C�lϚ ,S��'$I0(a�œ����?Y��?Q+O:�D�O�M	 T
Xi�U��ǒ�{���`����<9���?������ C���ͧ$/���bذ�yЧ.V�t���'���'�]�����a#@�����Ҿe���hC6�Rep,������O���<��F��L�.�x���2y��s�&f�liB�hǨL���lN���?���vNEJR�]�	/+ʭA�a,�����排J"7��O���<YdJƗa�On���5V�A�<��!B-�����c�	����t�F@ʟD%?��'=��A¥��t�>!�. =��'r6t�b�'�r�'��t_���9���!J�LRZ���c�^^�6M�OF�$W�*��1�5��	��9c|�Y�E[���`Z�0eZ��
�?Z�6m�O���Ob�I�W�i>�c��� ǜ��L� �|���D��MS0��?����$�|�)O~��Z�{�@�J(i��9�T�ݠ[�F)m����������Ж��D�<���~r*wP٫T�\%vm��LK��M+���?��r�x�S���'���'M�0:�%*�4xh�� U$�"tqӴ�d�$����'/�ڟ�'.Z� ����J��Zm�5�V�]�Eh���i]��Ʋ�y2�'^b�'���'���k3�P `Jėb �䛖K�'|�Vd[U&���$�<������O>�$�OR5���6�QڒC���@���&J5���Op���O��$�O��>Gj�z�9�Z��u j?|�K������s�i��	ʟX�'�R�')2EB)�yB�i0ư筜�*
��ʃ)����m�؟p�I՟���wyR�̀�v�'�?��o� �J��U `x�E�-�mZ����'�2�'��I���y��'��$)J�p�UB��f(��Г�pc���'��\��
������O��D�����A�0�`X�☉p�и�aɆK}��'���'��:ȟ�˓��
3rC����4Ʃ�䐧�Mk.O2��"�����I��I�?��O��؎uk@!���M]� �� ){����'�Ҡ�yr�'��Inܧm�<H8�D�.t��B@�G�!l(����4�?����?!��#���LyRBK=��1"Kǵ]:2�C-
�a��7�߱(@���O����O�"g��G*��Ia�!R���H3D��7M�O��d�O4�Д�r}b]����R?y�C�V�0�ǥV?g/��	Dj���i�ICyr���yʟ�d�O0��cӘ��G�8k�� F��j�4�?�G陼k��	iy��'��I��+&D�H�>Q�i0s���Dj�{��'��'W��'創=�J����D�#Ȩ���-��6h���T���d�<����D�O��D�O�x��ǘw�`Pf�N.t��0�@��*G�$�O����O>���O��|�=�?��<{��>��p8��	������i�����'���'B��2�y(*x|���*<S(%�����Ff6��Ob���OH��<���_�]���ӟ�1� /F:��(	�D,��d���M����O.��O�{�1OF��Q`T�٠*����&ď)�`��4n��$�O�ʓ 2�4j�\?!���d�S�gp���.C�(����F�c�E�OZ���O����e6��%�D�?���$]�li1�ԋ������g�t�����i�"�'���O¦�Ӻ#��P�@��N'M����a�Φ����``5�x�H'���}:A�Ď�@��'v�ȱ�4-�ߦ-������M���?	�������?���?���3d��0�U�?�BL��
<���J�_r�'�o�~�H~
��5S�B�U�j��%*4S=���W�i�"�'�b�H rl�����O6�ɾ`�4L�0
ʵ'��h;D�0{j>6��OB˓R���S�4�'�r�'�4���Wp�PX�F�~',���n�v��4J,��'1�Iڟ�'0Zc��126�S:A(�8�C 9���O�S�9OP���Oj���O��$�<���kwdu�Հ��1~2��F(�g�\5{AW���'��S���I����	 ���p�e��1��EySa��5�ԅ�Dh��'+�'�O�&Z�hr>�2Rj_'d쨔�vD�	r�p�W	t�Z��?	+OX���ON��0j����>C22Q� ��k�-�>HP���a�	� ��ʟ�'Ud ��~���4��k��x4��gټXe��٦��	Ty��'���'�0P"�'WR�'hxT�E"�8*֭�1<�Ɲ�wGj�����O��_*��b�R?Q�	�����䖼�u�\,s�����+cu��{�O����O\�$��=?�<Y����C�f���k��ЕR㺨h�m˶�Mc)O<u��%�릹�	ɟ����?�i�O���"����oH�O�L��Z'�F�'S��0�y�d�~�θO��Lc�D7�.���؉=Ȑ��4Ԯ�8��i���'���O�4ꓓ�d+�ne0�≶����KV)��o~����6��̟�/1ڤ�fԕ�`-���/��oZ֟��I�p(2�Ϩ��d�<���~���o�剦�K�`_4ur&$B��M������AU�?a�Iן����$)�1�q�J$!�� 3&�攰ش�?��)�X��IKy�'��	˟�ؽa/����i��[�yb@	�<��	:ެ��?���?����?�,O��p���s����@脽���A�%�J��'f�۟ؔ'gZ>���'j�C7m��.��E��I�8�楹� ���y�'��'!��'��I�E?��ۛO�`Ő��N�=�r�����n[�M�۴���O���?����?�I��<�!�~�F���]���D�MGEd���'�B�'�X�0��ȅ��i�OkL�8!��Q��Y�X��A�\�5L�6�'Y��̟���ȟpɳ�k����Mc��p){�`Ԫ��9*� 4���''�P�$b���*����OL�$㟦t�+��ݵ��� ��\�Q��'��I����Ο j�4�'M�I$>~��B6��nM�� ������W�P��@E��M����?I����]��]3Z�FAU,M� �:U��s��7��O���˛r��d?�$>�S(���\Yxj����þd�޼j�4l|Z@J@�i��'���O�nb��Kw��g�l|��CӲC��![����M�����<yN>ɏ���'͞]@��Z�>��V����0�xӬ���OH��Q�P��>a��~R�>ݴT@g��Q>����T��M�K>Q��8�?�+O�i/b��5�Q$)�V���ѻJ �h�1! �M���)�8�`�x�'2b�|Zc�\���
z���!�hfR-�'?���'z�����ݟ�'������2\}��J���F��d��L�nDfO���O��O��$�O�4c��V�%8��"��>E^P�"�g�l�OT���O*���<��F�dX�i��A�sG�k�4�K���2K������	f����I%~f�]�Ɋ�� *��C��ה0���\�ܱ S�4�	�����Ey��ևf������@0��Ѐ���1�<qB�A�ʦ���T�������1zĖy�If�K&n ,�B'�\1~�����F��&�'��_���� ��ħ�?��'f �₦ӷmx��	D�ސ1�0=���x�'bB��;�yҝ|2ݟ�Ѓ��8�v�[d�$4�:��5�i{�Ib�"a�ܴt��Sݟ������7��Y��DW�C�(���(�EK���'1Z�}�0&��}�/5��u@��&1��D*7��ϦI���T�M����?���
��d/QA��'U�"Y�"-�At�lZ�I�e�	P�'�?�@#�"'���2.Z/9�f��u �>�V�'X2�'ʐ
��'�	۟��Zu�����5P��X�O�n��l�Q�	�m�H|z���?�� l����$6���@� 0ؚ0��i>�Z~�b�D�I|�i�UPv��7���]�#'��c7��>Y����<)O����O.�d�<y����f*��f$����y�b�Iܨ��x��'SB�|��'RrJZ�������6�)h�(�=Eb���'G����	���'�XZ�Nf>m��`�E���֍��Z"���%#��Of�O����O���)�Ol{�兀bE.5�G�TZ���̟i}"�'���'��ɏf��I|r!`2�PLZ��N����2�.V����ҟD���Pɟ�Ik?	�կyQ�p���gW �'$��]�I͟D�'���b�7�I�O.��Ƣ�Y%M#x;*$P���d�j[u��O&ݢwE�OL�d�<�O�����2.v��"e��V D@Q�O���O����$�Od��O����<�;P��e�'h�^9V�ɩ7�z�m�ҟ��	Z����'�)�S	�p��k�,I7i�<`1|7���0/�n�H�I͟P�Ӣ���?�A(4�v�2$mǗ8L��gF�gY��b���On�?���hid#�F�DW:0R��#J�x��4�?)��?�v+�3�'Mb�'u��i�q2��';�8b����2�O���$�O,��Oh��r$�M�ZXr��� k�F$(�˘�Q�I9u�<T�'�'�?)N>�ґ4�$����#=~J4�ӯK�<��	&8�R
�M&?����?Q���$�;k�R!��3����&�uW^�¤Fj}B�'e��'R����lI���M/�Ul�BX��4�D�O����O��$�O֌�s`�?�Z��@�ykH�Ö"Č,*���hӼ��O��D'�$�O����Pl�x�iw�ć,��q�]e	d��?q���?A(ON|I�E@��'x�°g΅-rV�p�^�(��eX��f�4�$�<1���?���lm�,��?I�Ds����)��)ZF,]�A��ŨC�i`��'���3�~�ҭ���D�O^�iJ�K��K3NCK'��
��D�x����'r�'%���y�Q>�IU�7��6[�0XF.�+b���A�˦��'�IE�nӶ���O
����էuw���8MX��ҡ�N������M{��?����<�H>���$���T��c���P1����)�M�mɼ��'�b�'��T��>	/O\�Z��AF +TB�&eF�}+")P��q�f��$�L���X��t�FdT1	 ����'P�6����i���':���uɘ����O��I� �R�a��=<�8{ jY�>��6M2�D��~ʟr���O���R�f��A�V��
i�'�#���lٟ�zCgX����<I�����Ok,�& 0�M
��1^���DP�u���xҼ�IVy��'�B��	�<�:���� #fn-�VC�T�p-~��[y��'*��۟��	⟼���+s~U�c��H��	�@b��S���	Ty��'��'Q��'����ܟ\A�c�"
EB�0!�W�Hr�PG�i�'G�|�'Fbρ&�Dy۴:�rtZW˚@�~9a�0�5E�p}2�'���';�	��]i��b�G'jA(��a��8p!ā�	%bΩnşx��a�����q�{��U�3rr$����.K6�o� �M���?���?Ů���?A����d�Z�2
��5hF��M�Ji@��Dh������	:3 ��	�,+�~��ՠj��I���w������\ڦ��'UH����`���O���韆�קu�ⅷK��I�""��u�p�A4�M���?QrgM�<����?q����O�^<�͚/R�6���������h�4�]cs�i'��'=b�O�H듑�� E�lB"+`��3Cw`��n]���	͟��'B���d�&��MA��8n���[`��Ub]n����	՟`3�B���<���~�B��3"q�i��%xT�K��Ǫ�M������,A/�?��	���ɍ��I��*��p�!"H�M�|a޴�?�a�U2?��Uy��'w�՟�X	����%Ϟ>���AQ']A��v,>)̓�?���?���?�(O�	�1�@�r	۶��WЩQ� ��%2��'�I����'��'�b�ȑG�h����$+px,�疭cx���'l�I�e��3�h��j�>hg�So t���͵,�lu�q!U�B�0�f�5Sq4\�V��.s!�$6{�0��@&�&҂b��;p�qOεS�O]9m֠��6�^5fq&mR>o���3��غeQ�i� �ђ at�!� �iN8�ǜ� ]���x�P�R`
�I	4ɑ��܈4	�@��'��yT��3�)9M[�q�~��M�O �ز��lۖq�'m��������12lv�peiV	D⮴�r�_�x��� ��'<�ĉ�̕{1t��g�:�H��'�B7&�y;�gφpIvt�d,�AH�u����� �@Bq$�+ А�/H�d�RD�>!�eK�h��u����xD\<@�!�,]��E�~�k��Y��ZԊ��N-Kq,Ai�Dկ��'0�>���,�Fe4 )JmTș�ϗ�m(~C�$�.|�tʔ�|��aU��8$�P���Y�':H��B�3r��rO�������>1��?���Ai��q!���?���?�;��x&��%�����ϜPW�ܡB*W���w ����N�g�	7n��D2f \̶|�l%K����	�R���{��|��2X�n��ă)�yЃ��B����Y=?�O�ў�(��qy��S,ȖXu�D	�5D��9b�Ѻ��!9�`�5CF����.?���)z+O��RPD �RZ�h� 	- !��Ѧ͖s?�5�¡�O��d�O��$ ̺c��?٘O-�׋��Xh��g�&d���C@�K҄آ���9N�3��'�Z��KUJ��3��-lQ�H�t�@
8��q)��O�Q�B}�e�'��q��(L!x��-��"��A�|N���?����6�	�@�:|{Т�#�����E��.�\C�,����Q�ot8@2��0�Jc�Ļ�O\ʓW:60�g�i)��'��`3�cjūF�O�^u(1�'3�&F�j���'��"
�6-?��ԣD�h���75�0�-ܽ7�x�3k��O����V�d���+�a����%I��'�������?�.O�V�c�&�{b�܅�4��B��<��?����I͋m����%K.��֊�G�!���	�$N���H�A	_��Em���'H[�B�>������Qh$�$�}'f�F�� M֘�0�CWR�d�O�H�_��e�ө̒\r�+�O�SF��	�r���RU��}ݲjC�8��I1>�h�z�d>` �8�F�O$�C�$߇J\���J&`>�(K� ���OH�d$�'�?GR�$���B���r8�h@M�<ѕ�D��訥�i!V|�`�o�,���$��m�z�80�o�Ac��>!�.�m�͟��I���DcV�|,����؟h�Iٟ�&�XT����"P�Pܡ�S$-�:�R��nU���Vj˝YN��ӢnOf�g�ɳ|�r ��J�0��Y�DU��x�J[�ڎQp1�?,J˷�c�g���`ӡ�oQ>�קJ"*X6X�<�J��>�O���r��@��})6`M I�����"O"K%�O%=n\�� �,t�ـT�� C��ᓓC��w�����F�
�Ko����j�7P�e�����ퟠ�[w��'�	��[���k��E�0 d�����$1�l �᫜6FB�ĘPJ�\az"��Il��S�G9Xbes��	!1&e���B�	������ܼ3c�N�����x���D!$y�C_*`����<�O��ؐ�Ѝ���5�.��R�"OPEB篜����pLѰ.ln1B��O�^��I�ӻi�r�'R� ���<����0�/���[��'�"D֤
���'}�F�0�7�9���~���
1c71Wh�8��b��xRH�l��Oĥ�T�α��:��D#6m�����'�p�����?����?�q�Y�+�H���bZ%T�B��Љϼ���O
�"|���9x.�Ȣ��7	-��K���v<c�i7�ٻW�ƍ{�hѡA��r�|��'��	�F.����4�?!����IB�a�z���/Ujt�
8-:T� �*�����Op��$�O�b��g~"F��T��ԣ�i7��(ДM���	�J#<�RA&770�I�4�HWi&0z�k`�����������OgƱS,Q�[��qҩ�Ib��'7<q��*>	��L1A%>�9�_(��d��Qq\J9��w�|Hv�ԧ�M���?��n�v��f"�?!��?a�ӼK&��*��qz6�M"0>��1_0�'yP] 
ϓ	�$�"'�ޢH��|"�Ӛ@`B��=9"�@yx���ˈ=Afh�"�G0�b-�D̓C �)�3��%d�z�yW,�
m\���� �P�!�$�(10�h( ǉ2]��Ļ� U:r�I��HO�	)���e�4]�r,�d�<��"�K�h	t y��N!S����O�D�O8Y���?������ нRD9������J҄�
	����"E�M�}R��U�7[�.�v-_�x�F �f���?9 @�T�V�Y�4�$�'xz H7��a��|��1P X��׭�?�������.�uÖ%2��>����	K���>(��r`�A�:.^����Z���'Ѡ7�=���s+�E�OyB�W^R�H��g	CM�̉�BR,q�"4O�2�'#�<� �9U�7S/L	�d��E��7�G�,���ɖI���!��(A��x�C׺r�|��@�0*��i���� |�r&������W�qR�t�D�']����?!,O`�#٦Ob`iSAM>^V���@���O�����[��Juk��:��@c���	���F{�O166�Y�d��q/��'�����]��R�D�<����?w����'|�V>����Rɟ�WLӮ~(�����/F�r���fs�6m�O�]�GL�O�b��g~r�
`[|��l�7Y��[�I/��lx"<��3o	:,9B}B�k��O� ��7�[}�ė6a�b�'���'`�zK���Lh�p���6���e�$�O���$�?[��Is�Ŷr�ı��ņV
axb`2ғhB���� l�$�[�5q>�,86�ih��'"�#)����'Q��'��woY��[ F���Fm�������u�r�����zb�S+��b>�OV����
L�Z)A��H�T�I!����
�b4�����M3f�:)��>�O Ղw �'Z�x ƪ���r�4��
�����|rmT=w��@/�<F`,肓d݃�yb�?F7��@�B�4�c��F���_H���&���&�X�p�q���WQ,� �^�wl��;".�O����O���������?��O� �W�O4 ,\P	5/���]D
�`D�2�����4T[�\Ӡ�Z�HI����'bD�B�I5V[�,�`�od��c��(`�~݉�c�O&��-rh�cHC�]|tU��.]�0�!�W�3/&�sUk��EƔH� m�%z1Oj��>f��Yl���'��T������YU��D������'�	RE�'��8�z!�ņ�;E�"Ā��2���0j͛+��{4��I������I��p<Qiܹb{d���!��)k`�J�2���sL�da���#~Y����0	�|�B�`l,ʳ��79l�ƎA��y�/c�����_��te��H��x2�~��"�O��&Y �ԯ�4\Y栀�! u�nZܟ��IO��i�1Pp�bO�b"��Q�:����Ϝ;M ��'��r��'�1O�3?��-��
t�D�u9ЍJP�Ƒu	"�'��:���Ƀ�G��A�+�d�F�҄F3Gu�I͌��II�S�'���kX����K�=:��Ѫ+D��q�&��u�|�a�(^� ���!�*O�QDzr�\�(Gtܰq��A$7QZ6��O����O�};��ׯA,��D�Ox���O��o*�G��Kh\���� @�c�Ȩ0.4<OD]�T�ָ;j�w�P�<�n*&�D��i��yr�O?`�|���[�w���u)�H�1O��5�����E>��@�P�#�E.}rj=��`��)��*N$F��ew��i�'�#=E���!�>�"t���r�6��g�I���xөOBK��'�'e�S����	(����`#r�f\�7a�1_��%�s�B2��?�%FA�vu�P�"W��h sH j�CT�`C��q#Lׇ�0=ID��,p��s`��u<d��)"}�,�	��M�&�iZX���	r����8�*)I,d�AP�V���Dx��)jB�ɉ]�8�V�Ք]% Ub]��w`8%��i;�ɡ&F�[wy��'U^��քݶ'pi"�82:�����']O!�r�'o��.�~x�|�H�1~nuP�X�_ֱ�qEډ�p<���@; F#E|ܪ"*|�� {q)��w�`�!ߢT�l��d�1O�M���'�rcrӒ���U�r�ȶm�O̠id�)L&$ʓ�?����� ��ܥ��Q$�Z)�Ą��a~�'��6� �]üE WaD'*Μ!@�c�E��-nky��)Ab6�O�d�|������?���H��9Aj��F+8��ă!�?Q���$�B��̘���`����s ��F���k$���/0}��·�O񟴍�!��!c� �k��=�����>I�-ʟH��ğ��IQ��R��ͣad�`��@;�.�Ӑ��<�����<q����n����'�*PBpz4H�[��h��L�jK��A���0��(F��
I�0m������Ο�`�K j"���	Пp�	ɟ����c��Z`݉L2PL��ʏ�%xQ�M>W,�_���|&�`�@@ ��揝��xi��	Q�_�n�O���׎_�����/Ad�ŃO��a�bn�%-�������?���.�Yb�S�gy��'��=�WH�=,6��r��q��vh<AG!Y=Έ<(d�>&҂�)���l~�'9�S��R��c1�N5/氬Q�j�;�⩒�/��Rf 2Kٟh���x�	��u��'��'����L�K��$���"�X�p�˻d�)��lE�
O`��Q*�q�b F~R�D�s�ژ�C��:�&y ��0Dn�S��*+��� oV�3G�
 A1E�(����T� ���(��I�2����M�m�<���O��ĕʦ��ITyb�'��J	|�`�'��u����y�l���>I��|�'��.���!ӯ�*���C�� �%�di����Z}V>�)�����M+��?A0��I�12P��$���#�&�?�w�� ��?��I�B��$�iE�'��aQ�j�kxz1E�ـ0jǓt�lq�&�H����O<�9M�38]�²�A��:�p<b�k޴.����'�+5O�5s]���A+:� ��W\�@�I@�S�'�?!0n��q�"���ͳ	����r<٧�i+􈪐��R���RO^ ����0�o��ʓdql�IFL��?�����L\��M!>"%�5�ӏ(���"W@G���$�O�)��6bj���r&��[*���c�R��S>�;%��zc&z�o�>Y���>}¡��NV�<��U'J�
�yA-�w;����ض闯+��8�����P���>aD�ןh۴�?�����?�E!R9;G\hkP�Q��\�Ѩ ��?���?�����<)�L��Nu�ݘ`���V��1%RF��Q��������
��K�RU�&=4�o����IȟHC�38��i��ߟ����pJ_w�1���&t�:�
Ļg�j��D��P�*�7��9[qV��S8)�*Z%k�2 �A�<9׭Q+���>c�T��.�U��ɱ���
j��˧��Of�D�O桨��Oq���̟\!姆=h�B#F	'8�6r5K]h<9��S�s����R�3�d$�&j~�!>�}��yb�S?"YEYaF��{�^eg5�^������h��':B�'\�ٟT��֟�7H��b�L�ҵ�\
bU/#�B��Q�D�EI����9>�Ak�`�/2��E2�χ%Kp� �ᑭv|&i#b��?q����G�'�n�k�C�w4p��Ң��Q�Z�P�%Z��?��9$�&�'���ƟD�?	1�D�xC
�R�͘c؞��FC �<���c��H�(
�=�H���Y�b���PI>��'Z�B��VZ�D��g��ug�'`���>R&9
Uj		��[�� �"�'��M�P�'-b?���sv��<.�������)�06ӐX\����K�l7��A��"��x�k��&_��:{$��o4V$<�����p7B��p<�������������$��r�¤yH r�W�(��]�'�b�� )A���D�;�X��T�F(�B�ɟ�MkDG8>˖�@�&V���`
 A��<�/OX�cH@Ħ9�	ϟԕOQ���'���f�U-|d��c�DY<X���'�!�3���Xv#��8���|�*���*�e۪.��L^�+nL��2�>�t��\wX$!�e��e�v�z��)\�n6q�����IE&�u��`��I����p�Rb��B�~�2�˙v`5q��`̓�?�
�x<h�+ЁM�
6�QA�\M�a��>�HO$�`sL�7/�� ��#�P���@���̇�	�ux��
`�Q$	T<����/��B�I6{���� M��Xa�_<L�B�9=�%Z���/z�8a���rbJB�I�K�H$ʠ�:+t�]�l��K�zC��t��h"�DP, u�J��=+ C�	 N :�DI u���-�1%?�C�	��@4���)"���b�P�\C��*/Y�E�C�h}BcՁ�5\��B�	 �.	eN��v>2͠��Z�NtxB�ɍ��9�F%+���C�V`"<B�	}zL�r���JB�8�"b ((��C�	�u�ʔs����+�nuH��()M�C��W8��P�:7:����ў}PB�I���\jS�#;�91�Ϛ�_�B�I)q��y��B�����\�dh@C�I#�PUKI�0MR�j�dY�C�I�Z�H�"��_�T�S�JC�
Zj��WbǙH� h�O�$�&C�ɐ҆m8�H߄ n. (%��)�B�I�;��5���[��PY�6H�N��B�	3=ê�Ӡ�C�-;�lȍ 5�C�	�Xz�a��
i�-D2-�zB�I�,�¬���-h2Ԝ�T̃�c��C䉄wj*)�։�G��L	�! �k`hC�	+Z�����ZL����	GTC�	!�^ ��aߡA���l�J:C�)� @�����(�X1���ԑ9�Nɋ"O"�hBH+c4JM��H,1�z-ہ"O�%����/�&�P��֍.3�s�b[*Hi�'6nu�`�O�Ϙ'�P`���)!�u���O+P�Z	����(��ٜN�}YSF �a� ����#:���p���u��
�"���0r��1��Ҥ�U�T�G~�L�� Պ5��-/��؟��p肑_��a�Y)�q��P@�<�Gd�+\f����T��<H�'|?�v�Ҙ���'i\����F�O=H0p�G[�8+vD�6f����'���"�� {߀��$lr��!�bx!�sI�0C�.��a���b$�"�ON���`�`hN�{�`�'l�|�{%�'�ܝ0��^6�R�\�F�(���g��+�X��A�\Όx�'��/���ƀ�~��{f4}�~���"�0r���3 M��'���s� L|i6`���+m�!s�Y��ł�O�C!� _��.`���q�!�y��!k<y+�"��E�o�=_g8�&���f���e�@4~q�����+��O�����w�2��&�)DPz�� ��81���'���̘W�:9�#Bܿ�tIPc��
bܭ;᠂�:����uC�$u�,�$�͚S�*c�)���?@��i%�O�
b�ӱo9LO�R`�M���ɘ7�YM ��r�
TR�U�®(r�j͂��Zw*@t#q�A%kl�� ד`\.q%�Z'�U�
�'\���<��
�%X�
�KF����Ru�O�{! x�a��� �.pIvT�44l�ɁH�N��J䬚j�<�ǋtWe�FBF8(.P�PeT'Eq���%A�.�d�����K�VT�ϛ<4��O����w]������m�a�A::�b	�'F�=Z���b�Њ!k��;)"�#�ˁ�*1x�.�\:ع�*RbN�u��j���=�� �_��L�2��'#pd�� a�h��h�@Ē<��m��H��C�)�$B<vxS1A�=����	b ��wh�U��3�'� U�❙=x��&��R��+�y���V��0k\�:�Cu��>|�lKO	�����0��S���PV,ω� �L	��"Ou��F���)z@��::.���P�~�F�!^������Q(�A�������O���;0H\��ܴ*Rb�Ё#�.�MC�0p�`��6`@�π�#n����@T�jX
��B���x��׉M�� U�gӐ���g�~�� �Q)zY��R�\s7�G:|�<�&�.W���/Map��?�!)�P5����i�^�0�� �r$!��� �.M�/ Л`����#�l���d��?$B��s�@�i�x�IW��+HtQ��R�`�nP� ��*P�@�m3��V,!f��	i)DxL�S�x�P�h�.Ќ!��}���8ɰ��ф$9��a6�@�d� ؈��8[�X@��	5X�r��Q�	"�T�e�;ONP�!#Ɗ[}����[��p<Y��XN
�j�ˁK}X9���նfU:��ߓ-�NM+֥��8F
�hT��8X�p�ŀ�o���(S���O` �ƍ#r��� �B���V���Cbl�^	��ყz�H���O�Wj����*J�F�dm�'u��8!Α:�*xd��5f��QD�ٰPbĉ�S���6L�'CB�/^�J� Xqw�)�_�ҙS�cޚH�V "D�=�6��.�;Q5�����a�4�Ӈ`CeҘQ�kκMV �<�ҍ
�/��4@L�q�(iAEAI�i]�q���Z#At��K�nP�������4�O�Ff�e��T�`��O����|��'y����?�1.���R4�� Fq�%�u�Am����e/�yU)���R C���HP���?��s?yQ!��YcR!A��r>�Q��λ:�\�����A	�qIrj�7,�Z���ɀDp�%;1�69������_+)�̲SD�#$͢�PA�E!}���.O�5�K�W\�[wb�ͰWL�C��Km�Ȣq��+��y����'+�p��<����kgp���.�Zg���g�^A� P�$T81����g5�9�"e��A@a���=1�l�!���Vo�	��x�#!I��F�)u&�$�o�S�����eY5m��F�����j�c&,��@�3���2�X#L���gLјt,QR��*�X[)Ot�1�`\�K(�\w~<i �Y,�	���Ʋ_�m�UᏣI��DH�6���``�J��J�6FB�����jhȡ��H����"�>A%�p�XgM�x�V��GY���ܥB��T�J�����I
p��'�a��H�huj��萔h�BP���O��3D�P��!���B�"j}�u!Ȁy��<a�H�a|�Β2�IIQ��n����f��q��-+Wg��T̰��,^��R��6�i	���j�����<)󧉗3�Q�%�_<^�d��x򯙷B��sw�^�\3tH4����!�)�3W�D��+Q� [�͂�J�r���uJ0��.L#��'m��A��baM)�ʁ��	:x��rT�L7K�J ZQ�����,�2�P�c��ԉC{0ձՈ�,nŲb�O^�x4R_�(�Ҕ?�H1���-L�y�ga�0��{0�,?��ҰC�<��h�9iݻA�Y֦YX���?y�����Kw� �qr��䦕4#�P�蚓0/�Z���0>���S�\�;4i^�
W�X���41�<3�՝�t���ּ� �J�hlN�3VO�-��ّWO�H���o��˅��3dpбya`���l��']�Ɂ��$�а{e��b�!�K�T���QQ'\#Q�XC����GrOU�0hE�g�&O iqt$�º;f�Ղ5M܋�S�U�K�L̵#v��N0��X��H�&���E�FyB�\�p���V&�''�&TP������DƗrQ<8�2��2��]#b&]����}���j@P����.ilƄ�d�r��ШU��>��ɧ.�x�XR��6�pȪ��^29r�|����e��aG����'��O���7<R��m����8d��P5�R��w�\�  R�"A��1���|0����|���<�����'�"�*l<����k� I�ҫ�/d64��\}��l��H�!��O��@bKC��6H�͓��)�$]��P��F�%��Ba
Q�Dj�I�a5�~B�*$P���y��ϧHe�a�f?= ڴ�񯂊���>� �����g�D�H	ݦK��h�QE�=(�瑡�l�@����p=ͻ'>���3��q"��R�K��K!0�oq�pyB��9�����"�~"��W��0���JcH�c�
1ˑgMV��� mF:�qO�p2�� %��p�A]պ�`q�C9�	P6`'[4P��Q��o?�bu5���`^�Q��k�OǘLs����PeǸGqO>)��������k�<Y��
0E���~∝<C`����D�iZ�.�?�ڢ<�K��hz���F��gL m̓}�cD0��m�Dc%&bZn���Ǭ_\�Ys�d�U�0/7A�ih���y�D-(U��x�K׽7�`�Q�̃|ϴ�$�`�U�ܣ��Vm�w=t�It��O�C����(�#!Y���� ƍq����P����	n�?b9��i�#-JH�P��3�` ��#Co�V!:֪�H%|�:� �2�)�'/:�n�gp ��"�]�4,���=��s��jr.]ۑFӲ),.�1U�3?�����P��6��FNTB�N�982ŉ/�ލcd�Ti���;:�=A-�$x���ߕE*��a4J�Ҧa ��D�A�C�I�'�y�*\%?���G#1�́��J�-�DS�kX>=�ў�J\3��Pdt��F�?9�NL9���9n)ΰhUI�O���ĴsZ���J����i��EĢ�8D��5~�T`E��+B�J-i�����' J,k��h��R��X%T��`��Ű���#gN9��)�!鬽�#��=��I�|$���N��<y��I�be��HB8����b�DyV#���U�#�O9�IaRiT�'�����dOz����ˌ"�V⟸�F�Ӻ��+ �>tT���HïQ\nQ��i�ɦ!Ӄ���#h�1�'������!mʡ�U�͉!2�a�ԋK���'��V�}�Ӽ�w@�2�EkJ�*�"��#뙇eY6�9�@	�
#�������D�uO�OK�m�;W�~lS%O�#-�4�dQ8TD@��4u�d9��HKq�Q��$?Ar!�ה���Zt	�Sj��˱�ڑO��#�I�]V�}�Y<.�Yc�4�N��&/�,oO��/Q!��!W͙)J�i�[�J�4h�CE�h^`��(O*8ФI/Um�x��nӁ"ByS6�F�?�6�Y���K/Re��%Cl�'gӿ%�0��*E�jQ���>I��C�<�(�����!�$M0l�9��"eD2؉�_���1��
��d/ޞc���@A#�I@�(�r�ȧ�^��@@d3�<�I �2�`B��K��A�V>�λ[A�#�뎰!jy�B
�U��Ob>�	���'/����'D�8��w�
�Rf ۹�-���Fi�b}hv� 8�0�X��Ѣ-o��͓�Rb˙���<Q�Ƃ^� �����HfL��$#E��'�L�� +U"B�,�b��^�g~���!�Y�#��a�eK׿�M#�'����a@X!�����O@�ː�������]:6�p��W٠�ѓ@��r�Pr��]!z| s�Z>}���(s	��� ���u�"K�b�:���� |Z9�rO]�l2��#�(�h@į�lw�b>c��9C&K)ȪK�g� �r�AAL�s�c�D�O��T9���0�t�2����R9k�u��F
7  ���A�˚�*�A�nH�q��.޸�򉐷u��杳Rp�R��!bQ����qf9��(�h�}6(5Y�ch��?�)�S
NrQ�3�
_ ��@E��&�n��<AA��Cn�"�,%~S���(l̓���DV%>�,��ݬT�Xdb���dT�'���H�)@o��4_��q$?��F�Mn���B�39����D�֊)��U��e����8���>O��!c�R?$<� ��K�d���3�d�����("H���=E��&qb�i2G��L�)��p<Ʌ��>1�xE1q�@�K��4�����T��2�fX�'n�D�ظ�g]�{?��"'a�8bqO�Ӛw6�ϻ{≮�DX�(�fK�@�-6�اO�j� �h�l��s��9�h�܈��Ђk���%�E�u��c0M+�I�5�a4E�)!
,�IX��Zc���	$a$��g`�"Q�8��G�{0AbH��4���Іx��w��$��S�P�l�9�-I����N	�:�h�
a�F�[��9u' Ka���$�/_�؈8$$P*3)"cGe�P!$������4K �"�vuS 5���1O�)�I�-v=�5���hDb�&.}��D�C��5��OdhE`�>O�,Av&I}8��g�[a��أ��2$�Տ��>&�����d�����&�5���h%�0(�F���!Bd��Ycd��r���`��?�5v�ح'?}���E�p�2���zi�H�MmQ�T
S"�1kX��O2��)� 293����_o�(���'*���� �#krF��&�0x�J�>L��Ўg�h&�c�VgX!�teI������(�h4��	�
ז՘��Z�,�S�SZ�xP�@�i���4�QHҥ̰[�0a:#��*��@ᵈ�$���1��Ϙ'\�����Ơ;��d��j�^����OL��i�0>=��
�s����=�����Y��K=K �p��A+�E����{�ձ �7?��1F}�JI��yǦ?	�0YP�H�/;ܜ�3$2x�����b�H�`ePbվ�rwbްH��uw�5j`��*s�����'	#>a��ޚ�l�pEm>��Z�Tڳ�;QT�x ����zw��'"���jC]u�ͣ�J�
��|3hP4�2��"o �r�zY��!��<A� C�lr�+c�'}����/{���G�-�Zaб�ï6��dJX�����{��Ɉ�t.x�A�݈R������u��Q%�aOW7��<��S�:l���c�5/\�����	�UW�q��Im�:0�A��8����SI C��9�\�*�k!0�X�K�I_7 !B�	>PPx��K�<[(Q̞ؗ&]��C�	�l�
̊���(��(1GȊ�o�C�	������x�\z`�\;y^B�(�D���#���w͖��B䉍i`���b�ݹ2�@����>*e�B��	d6J�{EA�
��4R�H��B�ɥg�����(�;���S	U��PC�	M���*�Õ�s҈�Bg�0C�|B䉧��Ѱ��/gZ����� !�C�ɭy�:�aud�M�
�:sCN�LC�I��P�9��F�)��c等7&�C�		F�%�B���c�m\�N��B�I&jf�� �옅BDp�b^9dz�B�
u|X ���}ʘi�&��)D]bB�� �]���Q�l�
�ꂪ|B䉃/�|�p�$ϋp�Zy�̃�X̪B��Eix�(-J��'թyلB��.'.�m�� F>@��t�ԝ\%�C�	><��I�C�Z��(�d@��	�^C�	����#�]=�ȸӫ�)�bB�	�J�D�{0HT��t����e��C�	�)��d�E�0�\�R#�8�pC� &TZq��'azD �b���_VC�	�a�ԙ�1�]�y$�(��N�H�C�/���g2Q�4Buၶ=;�B�I�R��i��;cf��ڶB^�(�B䉘t�͙%��#O �1�Ip�*C��!�)P�-2��a���Y�\�$C�	�pG��k�<*��Ȅ�&��(D��K��ʎ������=m>�+G!4D��B$���E�&P��`�*	��x�2D��B��L�t��}�$�?W�³b0D���7N�v�x�U�I/9��$�3�.D�lq�kٔ_%֡c!�ȼ���+D���/�V�zqP'̞wi����*,D� ���M�9�v�5ʇa�L�Q��=D�({��,+��T��d�J]�(�a�;D��+#]4}:~�h�&B
SNH�E;D��B@% x^2���:Q��qp�&D��w�)tޡ�ìl�a��$D��JeI��2�@P(s,��6�#�E D����"��U�.݁%k^;2��]R�J>D�У�(J4%�y3Wb��u�X2�6D��@�
�0d0i�F�ۥ-c�p��.D�t��L�P)��W�@
�)D�@�0���'��P����4ð�,D�|qb�	w�yB4n�+��=���&D�� _�6� U�]�_��5�Վ}*!�Z�z���˕Ś�H�T3�(��] !�$�X$ъAՈF��sҍ��dl!�� �����k+"��-ۿ`�X"OL�j��&A�As�B�+�8C""O0,�#n�|����<�h�af"O���cڤO��=
�F�?y.�[�"OE�eA�'m��!�z֤H�S"OR�H�GXl68��u��#�ju�"O�t���f�dx�WBG-.��@2"O�X�wʎ2i�8��&bɑ#���`"O~�!۳"D�5�Ъ�)(�D���"O^ܒ#��]`��E��+Jͩ�"OΜ��K)R^E�g��~r6(��"O��ࡠ˛*f�ˀ�݈vd����"OP��b*G�:���a�ϖ6p��d��"O^L��J�b� �:��5U��}�"OL��˓k��U�r-5�R�"O��(����Ғ��d&H�P�@�
d"O*��
*����H�=��a[�"O$�1vb^b�z�h�LD\�V���"O�ؒU�̟�4Qa�r�Xm��"O,S3@_���Brǰ�t�""O.\�BO2zN�	aц�Q�A"O �A�Ɩk�$��3����� �"Of$X�@\�T�}[�����C"O^ܘ�L<jbp�C�������P"O @s�֙!�P"��Ҹ���Id"ONA��e=E9�m���ڬ[��a�"OD4P�#�'PD��p%��+ho�Д"OP��f�G��ГSb�lx�h?i���S����H"�F�]�x�{�g�/M6�LF{J~�ש�8!h�<Cd� ��h�Q�f ��xr�Y�T8�ൄДT�K�)�0e��R��lCsn�4y)`��bf��uE���w6��p�X0:Q�%pD�,+�@)��<�(e���3N��k�b&j̽��-"]ǉ�m�Dn�/6\@��MF�|ɀ��9�*�9%䛣a�хȓ)���2��E�"~�a���1��A�2XhV#ʳ��I���QMF���h�A$Z0�P�!ib��ȓ;�ʄr� �!:dd�C�Fi�9��Z���a�hTY�v�s��;fqn�<�sS$(�
�A',@�>��Y��P�<Y����y٤�#E�p��I6��q�<��B&{�\c��M]����&���<����1
5�qs�J��l��(�G��Z��B䉡f��k#�M����bg��F`�B�I�r+�͢�f�2X��RA�/r`�B�ɚkT�c�!,
�,u�^C�i,tu�H�:��-p��Z�J
ʣ=I�'��)+�����̓,�0DC���ȓ�<|6ˊ��*с�c٨X�8ԇȓL8X�'H-mm���w�(7�Dȇ�]M2�����CA0Y�N;(��ȓj	�I���:H�����e���F{��'^��%�]>kv ��LU9.�%��'���1�՞yh���ΚZ����N>������P�ph���բ#��E�R�֯_�!�� �Id�I���k��֬Ąl�!�;�&i��#�	^ ��!�"O�cb�[�a1*u��o/S��)��"O���`+
)0dY��h�$E��lɰ�'*HU0��ĝ�\<�#򢁮_e�@�UV���@9/�P���(�.#��E��E���䅾mό<�"�哎I#&�zaa��c\��a�K�W�BC�)� ~��$�.2�AEb�BV�5Z0���I���'%�9}3w��$HHb��/D����/	,i�©FB��I�i.D�@�t!:�l�QCŷG�f��!D��S�$T|�b�� ��ZcM<D���7�M�i�ã)�8}�4£e.D� �6��u�6�+�AkHD�ek,D�4����*�t�yO���wF>D��q�*9!*[���(�Ƒ�`�(D��3 ͙}4>�R���,L%�(D�`�B�J��C4Ɣ:�x�U&$D��I��E̸pᰃQ�z��y� D�0�활6	F���nO�스�A� D����d�1���(�O?&\@d�1D����(lIH�0�j!lÛjJ4C��.�5�M�g�~ Q��'� C�I�&Lq9�(�}�"��99{ �d9�t���߄7�<���[�%?�R$	(D�l!�W.�~��	_�	(*,a�$D�|+��@��.�ps��C�>Y��$D��BP")� �GJ"# M��=D��
Vm���}J�"�+#s�9��;D�șk� l5�T�u-.g�q�t�8D��2�GLqG��`�q���DG5D��"Z5(�v$!��)�e7�'D�J�f�x|,aХ��&&�HZ�1D�\�ҪA +�ց��C��(n��ZÃ�>a��铓
]��j���4T�$�����6&r.��D�>�tf�=9�n���#D�^ƽU�|�<Yu�S�4�F̉TI�9�>�áo�<ك��N �E�Q�!?F,�0+�R�<9�'�>\x�9�����@f �N�<A!J�q�BkV/ZKb����DM��|�<Qt,T:<� �X�"\-3��Td�d�<q�C�<�r�)�2^ 8����_�<�T��h"�ЋƩr�,��dΆX�<	���?�.�8��M#R/LE��z�$(�S�'_$���H�*��|x�n��!���ȓ,�vJ��	�euv ���ڂwajY�ȓ,o���%�1{�~�� ,5K5ꘆȓ@PR�g�^��r���� 8F}���nV�1��$�1ag@��3��8�B�	��V��dkU�jt�#l��`�I}��h����%��m�>�s�J+w�6�H�"O�V5p�V�C�BQ��*9�`"O Av�N2Y�����%��| #R��F{��i�M��qs����'+Լ��D!�DY]&��eF�o>X���.)"!��܇4�4���ɹ-8Z�,['{!�$��l5x��A�Y�:�2�-2!�D
N0���B� �ޞ{�!��)a���z�JАMq�� G� �!�N���%c�%kQ���4IE�O!���1����w�	[K�P����=!򤅡P d�J�g+@�+�Kޞ$)!�DUeW���H�vz ����;6!�䍸tZ���˟O�2%�3j[0c�!���|� ��9%���+��RR!�D��5ݬ���Z1N�֕ q��HY!���4�ĸ#Q/����f�ړzL!�<}�K�I�e����G:!�$Q�NrQJ�)|�)�Ӏ0rE!�d\�S�G�&2�+��	)�!��Eتɓ��ơ�."/�5R!�� ���Y)^y`�{�W�<G8q(B"O^��a+�������MDn��"Op�D� R ("O �qN�(�"O&)�c���h�PףH;��	�"O��c�$L2z�|�R^-O5��Is�C����\�e�qa&�4s�A���!��<	�)�Aa{`h@�Dnv!��J�,�U�*s]��$�Bh!�d�/\f�"cB�<4%{vĒbI!�Զ��m:��5{8 �2���(
!��71Qx�Y���:6/R�����v�!�Q)Wp�|���!"�8���C�~�!�l�*I�2��#d�QP���!�A(SV�)A��͵7������Cm�!򤍊Y&4)�j��Y�$��p��>�!����X��#Q%j�u�D��;a !���1=��S��K��9�D�;�!�[�S`<�U�ՂF��q@�ʫot!�D�h�0���G�[4�a��6G�!��I����C�)F�Y��	�!�D�<�:@OJ<sd�R�Ď8{!�D
uöH�+ ��|�oIa!�V����3f+ڔQ�0�AX���$"Oq� Ϸ}�nų���>|��4"O�P3�0`Ńg!�e_*<i�"O�H6��46%����ˆC�@��"O��0f�Zg8=S��B�(��H�"O��+ �!$��<�Q�����qYS"O�E�@�2�v욗��-�^��V"O�}b�H��y�d�jedI:F�ޔ[C"O�:���K��Ç�V�,՚�"Oʠ�e�{"���ł��L<��"O�C��'6䤺5$�Dy{�"O���'���"�H ��jK,�3�"O��0U��>� tksD��F�� )�"OJmQd�,u�0Y�#��F��A"O���O�Q�{���`��%c�"O�J�o��VG�]#'�!j�@p"ON����X�Z�Ife��W���"O��)�e N�;�$�;���:R"O|X1lR̀K�cO�9�^<!2"O��B`�R����p��4u�-��"OV���'��~~\H�		
J\���A"O�=ys��-;���'��cZƹӵ"O�XPu�I�s� �j�
' kl�	�"Od��A�ء���C����_b���G"OIdI	�'�~�+�e�<aX���T"O2�-I �$����t!�����y"�U�klͻ�&2i�,�1��y�g�Y�<� �j,^
}�����yR
8��cFD�U���zQ���y�@۞?�X�y�^�G�N9 F�9�yBO-�D�!���<2��p��7�y��;�4�E�\;g�.�mB��y�*�F���6Ŝ�Q���Ȱ��#�yD۴P�22���-G	��c؏�y�@�4Z����݆�DL	�+��y����C�M���@�(�x%�֞�y��8Bĸ%� O5���D�·�y�_�y�0x*�N��.�jE�3�T$�y'V�Q�ܡ��h,)��YbV/ۚ�y�"�0��xI��ȶ6t�X���S%�yRi>��abeE73HD���֫�y҆�.&�����92°��kI�y
� �l9���,����e	���"O2���54y��e�W�MP���"O�<FH�vD.TX�D_o���"O��gR�f�
@�ac)OA��S�"O8@�mɰj~΁"d��C��x�"O�8MbS$�jG^��%"O�p;fo�:�vT����NE "O��BG���)���ʖ#�Ұ��"OF����ʉ)��7ݽ�~}�T"OH�S"�1- �W�<�~P��"O<i�6j��	@d����ǌBd"O�����)��91v�R�8���"O�Tz�1��S'���� ��"O,yug+X`H�3�K�y{�Y��"O����,p�Ҹ�0%�/L"ġ�"O:1�")F�]t�0��6<�,Ӷ"O,���@�_ -br�X6TW�)f"O��ĩL�uTA�'��M�e��"O��{�͍sȸ8��3r�NF"O��p&=$:��4'(��l��"O��+uN�\ۮ)z���E�nQ�D"O8���*�^�Z�qj:T�ڀæ"O���5g�4*_��"#'^�&����$"Ohp1E�I��*X� g��
D"O�~�Z�i4��4y���f�Q�$!�$�U�,	����"��$�S!��XO؀۲j���j�f�%l�!�D��>�ZxsW��F[��(we�4ZW!��=��3��KZpQ�tD�^G!��
�OaTi6�B{E.���B�Z;!�ŏe)�c4���~��$AH!�d��M�`z�MD	qi�Y���Ι|!��І+W�F���aI.�!�d�!E��ŀd���sgGƘ@�!�䅏""\I�,�F��b��^2H�!��M*r��d�M@�(��@K'@�x�!��˞NJ�U��ּJ�b`câJ�!��4{��e9͊��ܕ�Ck�>a�!�d�>9$�}��N��u�ǊU�?�!�$-Y��I#7G[����f��!i�!��L"t)R�o�+���eo�5Q!�Ğ���(����iv�H���D!�^��Ҭ�r��$2v�`%�@�'!�$�E�l�����*]��y���ެ,�!�$�t���ȗ�L�{�ψ. �!�dX3N)jQ�N�vA���W�HW!�$P��|�*@aU�	��	�:T!�D���P�P� :H�
�տW!�D˺v�t�i	42/ �y���(#!�$;#��A"dË�f�Y��Ԉq!���Xp�/��5ȇ�˖p�!�$̖L��=J�*���z!�ă�!�D##Z2����'�-�_�[�!�d� -6z8���
(G>%�UG�	R�!�X�>�8���+��Z%M��cZ!��A~�����g�ց��)^�[J!�$=���V%V��ڍ#�愄N2!򤌥E���W��a�V����g!�$R��h���Mާ"�NP�Ҧ]��!�$@�F�C� �^��6���E�!�D
�'���A
�8j��]16�ΖZ�!�D܁�l)z���\�Hui�n�7j�!�$NF~�B�Ƃ�`j!�G��!�B,;�8ᥓ+ה�z &�<!�� �M��̵y=T�iek�ML�-X�"O�aѤg��$�h4qAk� X9��D"O�0�l�:&���/dy��"On��`.�-c���2�ǒq4l��"Ob����}��q`#%�@y��"O$�X��S<7�`��w�b�5	�"O�9�ҕ?����3�K�oڐ�w"O��3��h;b��r���9e,��"O܄b󌗸3���U/�RS@5��"OB�Г�qW L{�m[kp@�ؠ"O�{�j��tz�)f��o2�:%"O0�g�� uX9���65��=K�"OʰaR�+<���j>
��!��"OD�	�m����!��[|�
PH"O�Pbc_kt�p�`_7T�;�"O��*F,F���+�͆wW.q�"O�� �AF�=�R�1"ýID>���"O��˔,�=�riFl� C?���'"O��U��<w�V��U��91.>���"Oj ����-}�t����h��"OX�4��O��]P�/MZI�"ODx��`��PI�ꇙKl)��"On��Ō��2z��C	�89�ZX�a"OV �$�/~X�RZbM G"Opjq�Lq�l@��۸^QR�C�"O��jE�A���%C^�@��}Hb"Or]"AiI�0E��BĶj��1%"OfpR�!��������y�DQ��"O���5�ƈe�0q@�AO� �X�"O&c�i�#����W�7�詩�"O�}j#�A$PՔ4���ܓ*�h�@"O�,#��D�t�A��H��e���*�"O�F!S�6|37)�2)����"OZ���&��cI ��ώ�B�6�:F"O���9~�nI#��Ӫk� )%"O�M�g$z���R��Tߺř "O����_�d��IC+W[��T�2"O�i�F��O��"��\&%�>��`"OژzWz�"M{$Ț!��!S�� �	~�OJ� Cc��b�Jв�I�,�!*O��D�O��$.�����mY���@ͽ|��h ���7��}�ȓQ�Fݹ��M�36�(d���v6�Ɇ�~�) ���Y�LeyU��Jb^���P9"��Rǒ�Q��̈�(�%���ȓ1`��aj5Q��	�"���4P<�ȓ|{m*A+A-Z�F�SwAM�RV5D��S�0�:�)4�D)]f�1�A9�����<�H>�ϸ'ktd ��t}qa"��Q�ֱ��'���u�V�8 �l�L,.I+�'�8��ѡGq.�]�����Ku�Ī�'2�|��\��mH�=��d��'撸�aƛ�9}8��I	 /^���'lr��KV)>R��
 �$\"Y��'bș�̈.6	�-G�O�@ʠq���'	�P(d��a�艫�8L��#�'��y��K]5L�m0�ʐA/f1�
�'M��*ض}�e���Af��
�'c^� r�[�/��5
5cV6�����'|�e��C�N��]��w#���' �,HUc 
Y"LE�T�D�9ذY��'���XwfyK�< �J**���N>�=d�I��i��L��$¥JFz,���I��t��KlC~�A��V�RfE��.(8X�FN;%�,�c��T�U��S�? ���J�
���M�-��"O�=�P ���f�yB��$S�#�"Ot����І.,:'c �@�F�2�"Ob���� "za�U���-�h9�"O�(�#��1V��CϘ30�D&"O�{�
�>y�	�M�Tm�d�@"O����\#��cw�N�Yl���#"O��k��H%|�]`N]*���"Opm�u�A"D��8�@%	}�d{�"O��w�I�/����R`�@b!P�|B�'"��OT�m`į:(��Fe�}�2 ��'�����"U�H~�F�A�m� �b�'���[ ��v��Q�>v��Y��'�;Ƭ�?'�M�7."q#:q�'�(AiV��A�~�V�;{(�#�'c(\�Qh�45�޴;`���x�BtQ
�'�dQ"�P��FMe�R ��Љ��'a��N�j�My���A0�����y�HV9#@RE���<c��y' &�y�CI4��)��9�rDj#�y��R�,���g��B9����yeWmc
��Q�6�q�U��yRC�&z��� �Z6)1�i �ʫ�y��B3&X��(�oEb�D`���䓖hOq��%�B�ЀR�ļ����*�j�;q"OD�q��
:�R��g��'U-����"O�8��ֶa{��'a+IK���6"O�J�/;�0 aѠA�홦"O��!�4�p!�A.6J���"Oj�a��3��y���5wXq�d"O(�B0h�63�jM�6��kR�S!W�lF{��)�,a䪕�0�ѢKN�iqA�!��N=�$��@�	N蝋�!�;\!��^� �e�6y8UP��Z<�!�DS�S���B -^
��R�ũ�!�ć�7w���3�ѯ_*��[o!���1q��1s��"%�2׆ŀky!�$L�m64��	����)j���P���)�i|��������uI�>.�~�;�'�ԁ:t@]C���-$Ԁ�Qdٓ�y��H�����Z(Hy�%��c�yC�'�nԛ �J�,0�@�X����'Ȍ��g#�ry�i��I�|�9�'R����D�%��Zb%Q7R���Y�'� (�T��
m��P	Ϣ2ofH��S�蔀T�۟�8tC�hGE�V`�ȓ	WU ���-y6Q��R���O�(��!	)t�ֈx���_Jl4��'��-�倓	^��1��AK��m�ȓt�0��)�B�S��W�aT0�ȓ5�y�E�f&N`��+�#��ȓ��3�B+
o0%qIԌ}E����o����¹���M�cK�l���F�+��E��b9D��2/A?H�d��C>'o�]b�)D�(r�af�^�t�ܿ1�Q9�!&D�s�!�~T3@�[�L8�q�T�#D�� �ڲ,պEjF��8G:h	�N/D��jr͆���12�)'N�H�dD.D�8�(�=!���;Ё֬<��=�6#+D��;a�H�1���$_�y �1b'�4D��	��KN����Fީ0	�%JШ?D�4�į��uЈ��*�C�����;D�x����M��@p�Τu��]1#4D�,P্�n��k���Bmp��3�2D�� ą�V.�(�>�-Y�H�!A�"O|	C�  �ĐtǷ`2N��R"O@��0,�c%��`�� 5�$	1"O&�����80��u�O��e
Y�t"O�	���� 8n��[�L�� ˱"O��R�M���\u[���g�P	��"O��ٰ�U �"U�i�a��0�"O�M12曣<p���H�	�0�(�"O��y�
��������J�8�"OŚ�mX �Z�`�D]��bm��"O���jUC�� �"��"���"O|)����%ĚT�������"OE��]�U"���QHD{�%��"O�����R-���S��rD"O����C,�k�� � /�@�"O�P�fƍ;^4 :CaD�H*"��@���O8�$=�'hˀ�#d��e����1`�9�ȓj��+��S��Yb��A�ȓ	WȘ�� ϛg/LTP�BF���ȓPB<�0�K�q���1!���j�j4��^��Y�������Y�a+��".@��F��YK�f�9�֋#[d�u��v��`��PͶ\�b������?)/O�#~�U��9^~��F���:�z��!˞l�<�u	
f��%p��͍s��T��@�^�<	�ʱe�j3�K�
'[%�$�R�<�@ɍ(d$Y�,J�wĞl�S�Ec�<)��7�����V�=�J��1�f�<!�˃ToR+g��hؖѣs��[�<	1���!"��Ó&�����NRb���?!������e�f`Ml�lI�$	�{:�PqB"OrlJ(�soƅ@�! I6�P"O$��N�n#4�8e��#x��"Oz�ei�qT"����'WT(�d"O�Qb �	=bDp��C��k��[P"O����ȡRÄ���[=/9�A�1"O����nC�q}��`DC|.�09�"O��#!�� )2���[	��uyQ"O�dXT�?Rec���5�hB"OR	���*:E��F^�w�$4�e"O 5XƋ��3e4PQ��;i�:�x�"O��򥅊��2�q �QW��{T"O�T#��nWj�s�.���2�"O`Q��L�y{�@sу�P����"OذZ�n�&mE���	�^�܁Ɵ|r�'�azB�A��T���ժ�u�d��yr��/?f�­��w���9tI���yB́�E	�l����o�,���EO��ylI)�Vt�R��Dyʇ�1�y��ř&��J�	X��kPh�,�y2�H�� �x��B���w���yRT�)���?�q������0>��Ɖ<�nl�b��KT�D��Mz�<��l�(B8�(po��c��l�C�ɨIwb<)4%��~��/�C䉵B��Ad�3U:��c���
&q�C��'=�h #'I�bj+p��r� B�I�b��8��ȟ	~�2�J1 �(x�C�	�IlƱ�F��N�mӈWZ�C�I�xR��Կ[,���[
#�nB�ɝi�&@��Bv�(8������"B䉲!�0�r��#el�%���Wx���S�Y�*�
&��c��%x�P�T-!�d����jt&E8��ԈA �D�!�� 	��̇#����4�v"OT������j�h�N!=Y��T"Ofs���2����L��&7�āe"Ob�3�  SM*%;�Ē�4���G"O�p!f�T�jRR�j��s�	3r"Od�(1��� ��`!|�x"O�e�'(��n�s��D%,?���"O6�S`b2:D�8��A�>$։��Z����	6�R� "bV�j��b��A�`B�ɂBv$��@��j���ȃ�C��XB�	x�$$�C�ٍqM��9�)��6NB�	��r]��\��Ĉc#N]�4UBB�ɊL�h#����X��5�"B��:A\����>8�p�b��v�>���i�L@B'S�[���oՆ��8�#7D��ѠF��)�8ӡQ.-�;��3D��!�!M�V0����� J�4ק6D�����K�fhp�FO�<J��8�7D�DC�	�I�Ȫ�̀~�,��d6D�|�פ.��8$L��lZn��,3D�t!ri"x (�X5.	�"�Z��5D�4�N&|���@�7=�T��d(3D��"�B�F7h`D�?^3�:!�/D�@A�� ��{��]e�T��(D��S��
#	�e�N��lDZw,(D������V�9�T�L�:s/$D�c!�	(���[�*�1Wz� D�\�� U"�r䀛�B���t���D=?��B<���t/aBxj�hQS�<A6j�&?p'��*hC@�����M�<�t���=�4�p��p ���	M�<���N*PY��3��N�-���j�F�<�؃7��2��B<����Ak�<IЌ˙@΄���ؽ+~���a��g�<I�+{��y�KL���!�������=����?!�'$�h���Y88$�"GL�4%���'p.Y��BF��`0��f5>$��'�]��"͙R�-�ֶ_�`X�'%fZ�gG�����A^kN��'E<��!�� -�੩ ��?	���
�'���b�(ȶ��4
�{���`�'�D=3�A�
[ȱ�뗉w2�����P
z�RUĈ	�t�V<jGl�#M!�$֐f�D�qVN��h+ASNӟ,�!�$�2�(a����$g̠�k˕$�!�ݯgz<�anL�e��I��	�y�!�@*<��a0�W�9�B�d+[#1!���7�@�J؋y��I�Eʔ2j�!�D;��t��`��S�8y���4S�!�d��k�TA�wN�ĵ!`jZ��!��G
x}�ӣ��
�*y2`�C�!��Q�S0a�BbŨ8v�ا'2s�!�ğ�L:���U��/4h9�փ�?�!��E�La��8un�_y ��(.!�ĆLq�LQE&̴g`@�c�`��_!��Û˂I�Վ�N�Ȣ�80 !�$�/U���3�.ʇ�D��EP�q!������[�
��,����</w!��P� dpp0�/��g�:�B��_�!�� 51 0UJ�}Q�|1��D�b �J�����C:j��͠?�̓6` D��cbQ�v�0�x�L���Ģ� D��jU�"{�9�փ ���̻&�>D�DXu�2 C����A�5c~]"��<Y����(�� �xS�쏪.��A4�zHjU�s"O�X8g(��J#��2%�0@H���"OD��tM�R�����/L��"O�14'X��8Ip5�ǟn���7"O|�aa�/"�u�$�@�/���h�"O8�P�����Ti2��q"O�xʕ��G���	ͤE̲9r��$3����N#?�][��ҾW��	iB�X;NA!�N�[Ѐv��<X�ބkdk�~-!��6,S�<y4c��X�'1�2�'�a~���<�n<BH�7I|��p�앢�yҤ�4!��3��I���"��y"EL�	&��R�@+���b ���y�&�f��W��%=�	�'L��hO���i��x��5ٴY�Lf�KGGC�!8!�� |�D"uLʀ�\Q�gƟ.C!�C�t�x�+SIL�@�R%�F(@!�V�?}��+aE���8q�D_�B!�D�_Ѫ0����#oL-��(ݻh�!��]P��(�i̫P_�y�c�;{�!�Ď�6<�d���	I� ad��3Gd�OV�=��nmipꂿzNб!A�FI@%r "O��3�[��hظQ�@�5-H,:Q"On���#��&X�"WI8f�YS"O8#pk�8^��XG�0h'bi�"O�e�*[/Xu�hwf��{1��[&"O�x����1aKV;�d�0����"O��jE�_�����֢�5�
ԩe"OH�@�I�):��J���2>_*( �"O�L�L�32�S#�ϡe rm��"O��¢E�u��XH1ʗa��@u"OPa	@ �H x�ьߢI����"O��"��W(X�~��Nb�B��"O�\� �-_��|�`��l�&�z!"O��L�|c�曁fq��"O��b
P���,�E�Qg tH�"O��JV/��h�\5X��	SEl�U"OƩ�F�>B#���(�/C<f	�s"Op(�mʶi������7A%X3E"O��;�e�)\1������/5޴��"O�d�7��\l���$AT��e"O��("޷y���9�֤`�H	�"O�U��M�! %���fɜ|�晳�"OxT��jL�d.�}��Z
;F^!"O���P@:�t�NޯT3�8x�"O��R	�"�੥l�#�$R�"O���O5�H��кUlڍJ"Ov�ʑF��j�� PKNd��@1"O�i�`��&B�&e\9|��"OPmr�;cpR9"�\:/9Q�"O
��� ֦���X+C2 �ҥ"O�L8&�112������l�R"OFDic�PX��@�A��
�E��"Oʨ[ �Sw�0�K@�HI��"O:���$W<Z�)@ψ1*J��ғ"Od�Hg�11l���P<��'�.D��`W�R�v���h�I)M��|�� .D��r�=��Xk0b�3*�2D�*D�d��2��<Aqd���0��,)D�X���Z���2���3�$D�0�	�_�ε�c��-|�����"D�� �@��w|:T�Fa�6u�18GK=T���	��W�l� g&���I"O��s$��1����@�M;����"O� ����Y�6~��sa�Z,�����"OJ\a�o�A=��pu�Ћ}إ�"O��j[ 4�RĢ�$k�NAY2"O�]�Fh~��-��o�=*���"OV��v�QY|�rN� i�8"�!��٦-  �E��S�N�ЮF�!��qB遥i3bt�lj���=�!�ʌDf��Sc��$(�l`�e�	=^�!�, f����Ȅ��2��UN3Ca!���,
�͘��Z&p�񫓊V�#C!��$��D���m���5��4S(!�dO4�`u`T�A�=Y�@Fi·!�P"c�Yr��U$ę��Dn�!�Ŧ
�`M"bm��^�U�e 1�!�DL�e�0J�N�2
0�r!�A�!��W,J�HI�7kͫlr��)π,y!��8*���a�͏m�x�T)�\!�D��'GP�����9@�<�4��.y.!�d�T�tI5ʪ^q�X��i͗e,!��V7hD�pEA�59z�v�W�@�!�$�;9.�y��(P�>*>�آaѼ{]!�H�BԈ�gJ&���!��w�!��15ry21���z}�LS_�!��G?U$��e�SW�J���(B=)�!�d�u͠h+b#�ҵp���t@!�ӻf�P����Srpt��LH�-9!�d�0���S'N�iZR�)�`GG!���6b���Ù d���v��G!��ښz�6�pu-��������!�$�<Nds\�������g�!򄐸Q�,�T��71��YK�ĵ�!�T�4����@�יX�H��V�:T�!�d�6{�
A��C�d��@�M��!򄇗´��#-p�8�Z���,Q�!�dP�>��`��h� ���+Cȃ�Y�!�$Y�R<\����=�R�@B�h�!�D��0�H��׬�&X�*q!���T��HS�2fB�ԉ��B�!�D�3���iYO,�hv�ґ8�!��1f8J0e=_G�4��O�Zr!�$�dn� ��U7{�\('��=[!�%:�r|�qW��i`'�v!��T�� �Q���.�蕆�0,!��Պn��=�ҊC��v��0H�/t�!�$�-COvHF��X�$�k�aӒ~�!�$��_�v}��D��5JF@� �!򄗻3��B��O��1�Pm�9:�!�$I�\���
QGM�H���;b�-Z�!��S*���#�X�;o\��L��oB!�>&(�O�=X�0�B�\�!�d�R$��E
H�_J����a�!��-q��H69*��aM
Q!���x�>�#0� jt",���!� �w����휜t�n�ˤ"A�!�P�Sj>����|��ʶ��@�!�dF!+t-�t�Ǽp�H�:�@�U�2�|��'�����S���*[�ZR@�[j���ȓG�m�'` } �	�Ɨ�����dc^�&"�̪[�DLDل�Ĉ1�H]k��X �OB�U��Մ�1��I[�(�r��PN�!",e��
.�=cdF�*o�i��N�q]����[�(h�	�Ppx�1�O״?N��ȓ'^���`�A�ò���(@���\d�<� V��#������E:`��l�"O8��#ő8aҴ�P�����"OV�)��_N��
#���-s�"Oܵ!1�7_p����6��-"�"O�Q�8b Ӧ+qR���"O�8c��\$"̨�IQ��<ZX|�"ON�*��%O8��hW0 �I�b"OPi�D)�<����g�= ����"OpTTA�C�:��+.�qf"O��ش㍡Q�b ���{֘�Zq"O�@RE͠yM"d���3AbB�k"O�(�6NX����}�~�a%�&D��I"�"��P��� e�#�&D�< �g»i�-!%�L%` ���$%D�`J�-���a��b��*H
�c�i!D���I�-��@��G)
=�B#D��S	̙;�`L�K�����a��!D�si� a�t]i��>ր���2D��R3�4mdB̉��
T����-.D�<Hσ%0î�a�k
�[��%��1D�0p4��o��P��qv��.D���G��w���u���A�>ջ�,-T� 8b�˻vXx-K�刷j��M$"O�eCêJ�{�
�� eL�Ol��0�*Oƽ�TE�>u�L���i�����	�'�Cb`M,i����Q��	�	 �'JpX�
z��فA�yZ�=Y�'�L�FƐ
oj�8�Oɿ?��K�'\�sp�K=�F$�BK�%���'!�p"q
�n8�S7�0EHp	�'FҨ��˖&�� W� � M��'	���5ō�'26H+A�M��|9��'�n�;�ҙ&�Ā���/~Sڨ`�'�J1x�-@+zzY��!��|�6L�'�T(k�.��R�hu�t^�?i61��'�Jd@]7o	p�(�ΐ�" Փ�'�~�A���*M���G�1�j���'z#u۳[&���
�6�YQ�'"��/-�*�c��T���Y	�'����Nrx�e�ü_L(	�'MR��瘲#&6X����P���8�'�0)��l� fot��0�S>E;�m�'�֍x'mC:��|�#��@ͮ��'�����"srj��'�T� ;�`�'�p#��#Bx4	W�K�{���'d�l9�&[�-
�� c�ʥg���'D)Q�E�j� x��6U���'�xa	�b>TC �"agQ=_jR�'l|4�4FG1Ts���*=g�q;�'�``	�)��.�vt���&]�$a�'�*	�@�ާ�W�_�
X�'�N��ċ@E��YǬ;]�JX9�'Ӝxq2��e�@dX�٘Rq"mR�'���7�څ.*A���B�����'��D�Go��xϖ�`2�ك	Us�'N<Y�G@�9��,㐪0i�z�K�'G��c"�4C�hЮ��p/�-�'~$����}��y7A	�.�
�'��8s'��u�\`�&�WC���@�'��}�/�/52�{�ɥOB�S
�'6&hK��^\�!A(Ox�	�'���Ɗ,&�R��u
 >l*���'����#� �(�`@DDe���'�%��ҡM���H@C��r������ �ٓcK@���$�$o��Rv��*�"O��Y򮟈>]hP �Nן1rT�2�"O&�S�7V��� �{�$�h�"O���;T�i���}����1"Ojy�� �-�FM�TNȐ/"���"O���0 Y�4�'�a���1�"O�˔�Ε*�n��$�j����P"O0���*����e�)�r�"O�J�ꘖoO0a�g�] 08 �!�"O��P���e4(��a�F*�ٹ�"O�vOϗ��4#
m#��1T"O4����Y�xoґ�䁈5	��I�"O����X5)�@A��@٢� }q�"OȬ��Qh�Xࣲ��B�✚u"O@�(/��x"���T��|	�"O^@cp%�{N��EP"��Q{�"O�%�3��A���ƃH�C�r���"O�3�̒u�l ��A��YV"O���gJ$Ru�&��'��m�"Oʵ���4=�4� �S� �b�"O\�(���.	���^r
4J"O�i�!.�D��XE)��o���"O���&A-K(�}ң�]�Y^$LX`"O$�W��}(eGmٗZ2"82�"O �BT	А`*e�.}����D"O2��G�~�z��dȁD�0��f"OM*��N3RH��G�[�)��p�g"O�"fn���Ny��E"t���S"O6����j��ݳg%��0�e2�"O�hc��k8���S*XY`$��"O�$�O�9����f.�^*�p�"O�)d�]bh���3Hj��!�"O�L+�̗�"�I���!M���`"O��;$$s�0d��lK*��U"O�=(�J�:vS��̙<>��"OtdrB]���J��	Rx�j�"Onj3�������#;��� "O�P���R*}�ĽS�I�\~̹�"O�Mɇ���!"��Y&�6���"O�����a�9��j�+f�:�pa"Ot麇�W���p���e)aXE"OF�saC N�Δ�$W-l|^L�"Op��� �R�a"�_9yԆŲ�"O`!)uQ�HUB|օ�o��숧"O��ס� SF)�� M�^d;s"O�]XƋ]*����wn��"O�ՉW#W�9B���A)I���"O�0�C�Λb�ГD��"f� �Yp�|2�',�+��/+�䜋ЭE�����
�'i��� eF��n��7��Nٰ
�'y^Xt'�������5[�`�j�'_���������D-L�$���'|R��fm��nt��àFz+��
�'7�ݘfl1_|�� �c�\��q�'f��DӶI�fi�　|<��3H>A�26�����T�O�E�f��U�X�ȓ4]Č"�M��	e��a�з~X��M��!QG.b����6J�B����7�(Y�ōpK�����շ>�pQ��hd1K1 E'O]�]i���3Հ���Ċ�ZB�۷d������.�� �ȓ�b�D�PV-��V%qx ��M. �����3�:CF�;tU��dk65��E��
SCW�Yy�ɇ�S�? ��5�	�~��*�v9�Qd"O�	����H�0��V�cY�	9q"O4��@c
mzh��,�6K. �bg"Ox�2�E�B���߳[�h!�"O����e^2��(;s(�f	V�Z""Oh�ʢ_�`%ȭ��,���<�2"OL����&g�l%Bp��3H�y�Q"O���1� ΂m[J^H�qp�"OlB�?}�A0�՗>��
�"OЙ(�O �
�+m֡_˞� Ak�<Is��/� �ROQ�d܁�P�I@�<)q�8V�昉�@A"0��%���N�<1w��0������/y�[�e�`�<�P�0O�ȋ��6��	�ţu�<�%C�S���Y@$[��c�^h�<yp`^�)��X2��ٍ~�R��B��<���ı^���pA'�qd��	T�<I�oQ>�n9��؇mP]���R���	c~B/�%m?�1�1�B�2��P3�A�y�ϕ!7�^ţ�-M�(��Ջ�*��yR�5��Y��hΧ��G�Y��B�	4D0� 8��Z�2� ���}>�B��)`��G5� ��r��y(�B�	'C��Pm�|�0�6�BܖB��.�����'Z*Qr�ubB�	�id�,9F��$�^��E�A6��Ն�1Ϩ�s������bƩ<FT>�ȓ9�	p߳o��lb������ȓ��ES ��
Cj��L�hC5��[�"1��#T�?�XZB%ۭV�T��ȓ>����	ڬ.��BP�R�4�ne�ȓؖ0
T*�b�����Y(cdx����<�#hU�?t�):T�ü8�D���Mq�<)WE�/<�pP�7(j�V�s�<�bD^�?Ed�!�`שk��ͪ���u�<񄅘�{wf��6nţ{ b�JDJj�<��m�EF� zs���s�b�`!ol�<���4�^��AcR�#�qpt�k�<Gj��&z4�b��Q�	pA�o�<Ym�N�&4������=��$Wl�<9�C��"��A��P	�́��_�<1F%��M����/��$-;v�TR�<	@�WUL��@�
K�Va��EZ�<������q�פBn��8�5RX�<������W�L�/|�Q ĎR�<�n�[��d��AJ�oM\l���MO�<q�b'i����U�^D8I#�g�<iф�q��&bP�e�Nm�� Uc�<Qr`(Jo�kgg(l��a9�I�<a�- ]ق�@�B$"]p<���@�<����!=T�4����S0����M�R�<�� �c�"!re&Ǹ8�8��ƍW�<�ѕt�FdZT�K5��9�OVx�<����FZ�(u��^:eZ6Rt�<���o)\��e\40|�2�U�<iwĀ/V�V�Y�M�	�t��BP�<&E���J�r��,n"*��&@L�<9c �*~�*�O��]��(֩�R�<�C���vh��Jৌ�U]tm�5�P�<Ѷ���ss� [2░-��ԇKJ�<��Ptj����=�-�é[\�<yS}�aӺQ�iPF��V����ȓ	��Q���
ߺD�&d�2|Zp��.^�Yó$0>p�1q�ݱO?nl��S�? @b0L�s���Hڍ�B�q�"Ot�Rt��*
9�]b��e9�E)r"Or�21% )VP ��O�M^��"O��E+J�>R�bdm9W=�0p"O�i��a�,\����KH�!"��2"O>�5�P�g�lmA�AI�\�eC"O��Q0�ٖA;$�q�O�W:� f"O�eiDN,3����ƊL7
Ԋ%"OF�Z@�ۨld%�VJ04� "OM�N�,wm�]�pF��"��`��"O�H�e�˞ap�L�k� 皡B"O�%�ㄫ4�̋�$�E���"O���W@�
j��ӣQ5��!2#"O�d0Q@��&�X��Y�VI!"O���ĎN/.x�ţ!��D�d��"O@<���Qo�Y�*d:hĪ"O�0�Bש2�<0���09�}8"O8(�.�`f�a�獛�#��Z1"ON��sc�u�,�ۑ�*9AC"O(,�b���fO^��FD�FH�	�k�<��98k$W$^|���֡�!�Sz�;!�UvKtȓ��Y�!�\o��8���ڟ!,�G�!�dū{\�ʥ�^	_!��3VY�=�!�$��t,�����=cJhR�#eo!��(��J&f�v�V�;�,RB�!�D:)�nH���b�.՚�쑥M�!���`�Mh��A)V0%�v�{!�U<h��k6�$)� Z �ي [!�	�!a�=b��.
������� :`!�DN�F�fM8#�E�m~X�q+A;Gn!�$��z�:d�"��8��e������!��=0T��+S�>���x��?�!��(z�]�g]T��!�P; �!�$4$W��C �K;Hj	`6O� �!��C��4+w�RD2%d�?v!��x�~����� 1R���؊#�!�ɀ�I�ŃW7�bb
�6"_!�F9wUR�X!]�#RD��$�!�dմ1Ƹ���L�-g�<xG��Z�!�,�b��C�'Pf�U��mU��!��Dx������0�k��!��`����p,�?_Xt�`���U�!�
BHՒ0�D�WF�Eig��q�!�$�<�X�r7'^.�t�fM�)�!��/K,������-�@z���0�!�_��8͑�i7��zW)V	�!�DM@��J�v��cѪ )W"O�	5�9@n�"ci��`�""OF�H�m��-��jÍo�H`�"Ob�j��Q� s��;T���+�"OTQ��e:r���Y@�̕e;<Y"O�mqdLߠnm�i���D�pAbT"OVY��Z�M���H�@���i�"O�ʖ75�]�EgW�Gu�f"Ol���'ǣ�L��acX�E[B�+U"O��y�A+)؄�R��tz��	v"O�X� �
^�T��!���di:���"O�} GlT:TL@` �
>_nAG"OJ���ɐv�<�B�_5eL�ڄ"Ot����["��m:�c��xg��f"O"<��oݼM��]
��4T�D�"O�*��kָ�@ � ��ʵ"O>-����V���Ⰿگ,�da!"O� n!	�C�0TjH��N��Ik�"O�Pr�c�(`�R�����J"OԄ�JTO�H����YP�,%J3"Ox��.M� e��!���"�VT�U"O
Ժ� *U�I�Nģu`h��B"O֥�!���*5|�"�%}� Q"O�M!�J�.!��R%(9Z�n�"0"O4q4�V�[�iClY�2�@IP�"O�-�C'@�æ��2#����"Oȑ2��5��!�D���Q��c�"O Iz"���9�I�;	��� "O��F��n���3�
�(��z%"O�M�t*�d���zs��*`��B�"O�|�$��)o��ɂ�&�^��܂�"O���t��Y�č�p��M�T=�"O l`�#SÐ��C$��^����"Op���!��_!�ܡ$��)#� t��"O�5J��,,�(![q�ت=�N� 7"O,����?y�:�:�m+,N��"O�p�P h.�%{�_�a ����"Ox�`���RU�ˋ�Q*h�3�"O���o�R�Eʗ	vI`"O��Dʎ�7��82d�p`�$9�"O6�Ƞ�C�*����Jߙ7�<3�"O|�	r�4�=��㝇��1"O�]��'�(G$�S #A�m���"OB���K./�� 	�b׵?Bz��"O�ݵFցj��G-� C"OF��EN�8��hj����Dö��"O���2�\���2B-Чy�n�y�"Op�Q�F�Im�8C������@�"Ox�{��ɸ�t�q� �2[�V"Op4
��T2I�T�cOP:U���"ON`
��E2Fo��K��$_��K�"O<ubF�B�oA�iyćʜ"��G"O�ڣC��1��$�F�;I�$"t"O�ms�J�!�A1uⴼ!Њ6D��+�$ƁQ�ꨋt�߷X�6EJ�!D��#�������r�@6{�$�b�A D��X��C�P�:�?�(1��'A !�䄿5K|ℍW3Bu���Km�!��8pch��se��(�j�Ha��N!�D�(������C�`���ҁيn�!�D�;���H�$p��*s!���+C��1B��C�|¥eͮso!�DO�$/�᪂���e�$u`�kI?6S!��>���VȐ�O��l{Aj{I!��/<$Q�c<ں��I��H!���C�H|�u���3�L�硄�"!�J�\@P�C@3_�@d8�!߸Jt!�D��Pﾨ�r��:!����C �+�!�S�1��FV�|�	�"���T!�d�:_���4B�� w"TC��68n!��nN��Eo�Nn�L{���&Td!��U�T�r�rΙ%�@t�`��#I!�E�*O���F�<nܪơ��v�!�G?B#���c��T(0HSa�4Y�!��+*p�q���(|4#�b�4��g;�$�3��Sy� ��M+͸��ȓaH��y�F�#I6�B�{0j��ȓ\�NTYŀAǄ����p��݅ȓdM,����G�tcd��o��$�ȓT���D#�T�@�ZD�����v������͖,��ɉ�䒞��`��S�? ��qE�0]5<i�w(�+9���"Ot���*����6� >/P��"O����. �.�PqD�&�!�u"O��ݰ}��h �M�b��j"O6D*�8�"����ԟ#��qJ�"O$9d�ĥ/��	"���}�"O��kT�w�B��`a�6㖼�""O�l�h:4p��+t�s/�Y�"O���`�T��(p����t�T"O�q0#�)���b�'>��"�"O^9��I�F�:��]�8mv`�"O���׀�Q�� �!k te@���"O����B
=2�aL@	q>x��"O
m����gȒe$L��&��Q�"O=��T��@�S!սa�"9)�"Oz4� ǔ
[���B*��ax� ��"Ol=Ab��3�Ԍ�F��3Ur���"O�!�$��9r��5�� 6F��av"OhĘ������2�,L�2JI�7"O��n�5��X��@#$�	�"O&\���9��P�M ~@���"O�q�G�t�&��fg�;��L��"O���� #�Ւ�Ǖ�*Ev���"OҰ;�L�tX�'J=+�C�"O�W-SOt�(@��1���I$"Oz��6�9wn}iSH�#���!"O�U(���ڐA�g�(�tx"O4�8q�A7}��#��7����"O8�mXE����f�<S9(%J�"O�(ҁ��.]L��%��q"`�k�"O���w�V�,�`��9Zn�J�"O����)
�NT�AE�#"O�$m��N�9��'� H[��'��O��Q7�#��@� c�;H��J"O�LQcA�3]���"�b�1g(ˣ��?�S�'@~h��h�P�d+������S���d���pssb�pFȄ�*6�(A���.H�Pwō�5��"O�YA��T��W��PgjU"��"�Ş>�����p<�!���:g�t`��Ro����(�
��1���=J��Ն�c1D)�wl�\������ԓ1� �ȓ���B�^+ �B�
�+ۑSf���t��+�E#"I���s��N)�x�Ojc�"~ΓAN��a!˜
�p��ϕ�}@���)�(�1�ͽa�~�Y�b�.A��͓��?cQ_��}2��3d�l,�%F�K�<)����@-�}�ЀƆYXڴ���H�'�����5p�B\xRJ�'o���󯇛.!�$կa �Ī@��J`�u+�+WWR���'Yp�璢&�4��QCX�%�Ƶ���hO>�̓3�6�;�G�+\��p4iK�Hk m�ȓ,a�_�-�0P�I��p-���?",٘g�|���4**��%�d�<��1"�4��Яڸ�� �G(U_�<!��"\�شD
S7A�P�``��Y�'4ўʧ�b٠���x�U��$A���نȓLM��k�m��lI���� J�$��w�	�~2Y��`�?��|I��&��B�I��8�B��j��T ��XBIB�$T(�(O8#>yW D-�����7_|�%�Io�<���Q:L	�i����+ؽ G�j�<9�ǿkC�a��|�tɈb�d�<�-�b���)TO�,2��c�<� ���n��^�.,��H0\b�s�"O:MB�2-�d���ԟ���"Od!��B<W8P��C��nT���'��<yB��W�̴Ct���ix��@s��[�<Q�T��
"�I�_Z,\��B�T~�a;�S�O�9�����t��L}��}y��)��<�u�p	 Ԣ�f���D��k�I�<	e��Ljq���ƃ�̑�ᧁ�<��lz��fT�w�z�;3f��6��IF�D�S
�)ԩ�2��u��4�a}r��}y�.7��@Rt�׿g�ظ���HOL�=�O�.�Ye�B�?j�ܳ���#v0P��1��%.e��!� sN>UP�BۣMȒ���	{�DG '�мS1*@�3��"���#�!��6?rF$ҥ�ş` �d
g"J���gਉ��KD=�� �� !��'wa}RcA�Q�9���]����C�N����8O�\I)Oh�*��B�ˠ��!��\�x"��'/�I*5I���:�B%2"�	'&�듅p?AA��Ȥ9ڠ�MC�*���+U�<��Cͽ�B�C��.*P�U+�P�<�(-|İ�WX�He��GWI�<!!%�>�d��%�JBp|��"Ky"�'Vܨg�C�a�nAKV �8J���ۓ˸'��a��(Yhk�����_7"`��X	�'T��ӧ�h4��O�L�,�؏{�Jt���'_��F.(U�$1�bQ����G|����|"bǛ�nƜ��5�L�� 兛i�'*#}�'kx�I�"�R���M��bd���'��O"���`�?&5h0X�@d21q��Ʀa�W���ZԎ0'�.���@�iZ P$��G{����_̈���6 ��:�ɝ�y���S#Ft��B�Z ��d��'4�{��W |,��πtxj�1 L��yB�[Z��y8#O/j7�xC����y�A]�^xI�L�<��0�FŊ$�y*i������#��`�$G�y�ѾHW|��G�%�T�Tχ��y2d�>>���pdªz�H�!$	�ycR+}_$막�� �8�3�٘��'q�1Gyx"E�(Gdt�@�x����⏰��x��7e�Rq�(�O��(ƈܫRB!�Dּ[R\m��'sN
h��n�n0�O2�=%>U 2�&U�,I���� d�u��%$D������<�F �2��=���!!.<D�l�E(��v7J 
�c@0Qf���c=D��"#/J�C�!E埠Az���$�;D�0X�Iٳw �P7��l.E�b�4D��17�E4>���30Ϝgê	�pn>�IN��8`���*@�B�ka�����?D�@�Ӫ��lnM���˳d���sM+�O����%*�A�����i�
0���̓��?A�*1�Fd�'lĂLծR��s�'W�?)k�K.��a�d�8bȔyW&2D��!Ci������S�����0��\���'@�2Dj�,@� ^�a���]H�ȓZR|��mыH��yЎϺ|�2�����xӬ"|�'������?&z9��$}�P<1
��~�h��V�8�	����VS�m͛F Sæ�!�>i��d�6Z얥"�����6Ii��ņ&�~����<�4�@�Pzԥ� �ƥ f�A�<��L
*��ۣ#O��E�I�|X�ܔ'��Lh8d)f�g��C"Ѓ{)�ԓxB����1O�E�t���t��-βa"~ę4�	y�π �P!� B�S$)ѩ�<���R�6O�̆���>n"�FʞY��1�dTJ���$$���&τ�%�� Vx)� 	�!Q��~�\�pc��O�@�	*��	7/F��/}b�'�kF��-$�P ÏR�+��ODc�0G��ˀ�  �f!�:��XRD�9@�!�$\�*eT�(���x��u� �T��O��=%>5�"��GCJ�I5Eߛi` d�h!D�ȡVA^8W��i	�*�=?��m	�F>��p<A�BG"��s�*��pa��y�<I��L�'��h㇇�4S>P���(�u��o��HO��-Q7%+�iB��,�<�xB�O)����8Ot�	:H0(�c�TBl�q�C��'�pC�I~tm����n��1G�d7X�?B�$.�	d�'e�p2�dRY^��0��R�C�B�8�'^��rƙ�:̢XpE䗯B�H �O��E{���e�|,��T�fE��LO�y�蚌n0&��%[O@FUHr�[�'��'TўH�3[�Kk�3u�>P��Г��5�����,��	b��fS�	�b/F�-]�B��,Rж=�@̴~t�ȓ
�q.O�O�#�� E
5sD�� ��-}�h���ZD�<Y��	f��hR�D�'Z �[����hl�\���Oq�( ��풥Hj*U�&g��Z��B��f<$����2�٠j���O��	�(�>����1k����!вy@�����<�Gl� jty ��|��i�l^�<�� z�XsT�CM� �CkW[�<��ꉄ�1���א�|l�v�_�<���@��Ҩ)��I	80A��Y�<!AW�~�T@v- 9�Zg��^�<Q�5{�L�9$�Y�&���g\Y�<�#���Do�l7�i����M�U�<��I[�].BDp'�U����ҍ�O�<AA�˴<��%yKD>�E�C%T��ʄ��0����1V �ys�5D��KdM�,[���P�%j��A@�4D��I@��2UbA�%���flP��&,D�`8�NRV�{d��N3z Z��5D�|��hϔ�ȁ�戞f;v�P�#!D�ؑEH 7
�	�@.��b�@(yB'>D�8@����Y�pz�[�L��p�;D���F��G"�!����X�ք7D�D����}���§�O�a�n7D�\�ubP-e@�a� �A�Az~�Qv�4D���W��|(<��wF�-�
Y14�3D���R�\>p���+!ʺIv�5D�l	�B�eRF�4Z�c�N=���4D�h�v,[�s�b�*A���`Q�\(��0D��x����"q�I� cX�#��,D��3M.)Y��* ��,H�b--D��X�F��Z�Y#a��To ����.D��"�然7Rp�pbi�Q��-u�(D�<PcaNۘhs�$F�W|��A�,D��
�郏x����Q�X�5P�	�F�7D�Ȃ@K�r������݉�� D�tY�ق�`0�㠀�G[�i"�"D�x�#C�]2[d�J�k��r&D�P��m�X���B�n	;6b"%Z�:D�(�]:`o0�ᆊ~�^I��9D���e%d�f@��ƃ`�rX@�*D�x�� I)���&�E�	]V�u�*D�Tc�@�	$!J�e^�5����)D�,3�&�3	j��o�,���)D�� ̩���(2����Cߧ�J	 "O�[ҀH�1H.� BY�9z��4�P9"��as�/��`�'{�c���VJ$M�W��:g���Q	�'�%���
r�II0��4Y�Q��'�V��b�*^�\��� HO(�'�`b�'`�J��ڀQ�|���c.T�|�/��fW����B�d�ȓ#+)D�H2���H$a�Q�T6^<B�%D��ʵ���b@�B��(d�qw"O�1�����C��6���|��{�"Olh�e*���%G�)5 <Ļ��N�y�[�J}���tH<S���@t��y҈��X�~� �ߐQ�q��y�@ݏ@Wl`[c �9KaV̻�䔦�yR�H7Vщ@�)F1�U�Ҥ��y�L�-+�c�H�:�H��A��y	��&�X�Heɔ7R�������yҥ!#��eX ��|�䰨& Y=�yb��-d�V�c��֮:F ��Q�δ�y���#hoFhA�'*ڒ��Sϙ��yb��E��C�"\�pyc���3�y���
ZV�A�&�]iH�%7a��y�=.@	�@��1�neqTh�8�y�	ޣ;|y{E�G�M�  �f��y�]�!���7`I:Q`�5�y�c���ܽ�e�a��(8��	�y���d��!i��
�fBlT��_��yRO17�<���˖�\�#�JE��y�B�]�@-����!�B�ۗDX��yN�7]ڎI���O)U�&L#Be^�y��P�A�LC��	�A{��P5G��y2�HmM��E�Uj�\)T�	�y�lP/,�#��V1���.��yB��C�@�(�e?N�T��Rd��y����(C�y��G�dYa�(���y�\��0�r�K�<��$���y��I$,����G<-�0d������yBm��~x|ud�� �t���ȴ�y��]}x���S�[(��*&�O�y�Iƨ�h�������ڜ�GƊ�y�!d����)̵��t -�6�yB�"RV�9S�cN���0��Q��y�Z�&<Ij���S�����	Q5�y�Ă.��`�K��B��8���+�y�?|�0�"�D0jիP�Ȍ�y�,*mx!�3��4?Ƅ�9��ի�y�� �<��%��K[1�-�4ջ�y�aZ/0�H2%�^;9b�Ō��yr��)z��l(���&/���Cb��yb@������wN��8cMع�y�b�Ip�SA-�At�B���=��cÒ!���] ٲ4�@�Xen�[�`B1������?n3x��a��#Zׄm�V�k�����0�ȟh�)�@-C��jg��ro�$��"O�-�scU.=����A^G��SA381\��K����B.�g~�B�Q��H��a��ԎN$�y��y��APc1I~ލ2�� �7�H��KY 3n��I�r2`�����$~}\�2�ΨFX���$R>=�L�`�"�~BLӓO�Ap�� ]t����_�y���6�t��w+���v��q����'�|���!�s�0�F��"ұ5v�)��V�z�&���lG)�yaг���Y����tE��ʗ@@�a��ʎ\�d�c�>�~yj��4F��Kc���Tl�_�p!�ȓ	&Ԑ3���oڢ�B�[�_4� �;f�\��m*�O� :q�#�P�[rd	�g�1�ZTH��'8��ëCp(.�����qC`Dv�TX�fMD;i�9�ȓ-蠘���=~���CN��~�z<�=)L>B8dI���� <$��r�i�+d�~���8t�!򤟾M�*F��21WN���lC�r���T�2�	�H��ɕT�f�O�GG^�5d�>�
B�	�Bz�ђ����%�
(aÇ|f�C�*2IB�w� �Q������+?�C�I�ю�ŌZ�b����u�ͽ�B��8dÈ᱀�G
��<S��M�s�fB�g����+Y�Z�(@��m�'(�XB�$1t�Y�n%Z����$i!�S�eت��؈HiNq���Y	@BF�K������'2Vl�c�&	]L���L�+��)�#E�3��T'>I��2)��9�6�'G� B�O(U�0T���R%�\x�'��8@�E��9̙P����\��ݴʺ�X���M�ǇE(hmB��������T48*����f������p=I�F$) p�a�w��fE.o\`�E`�(w��䛲�W�m\ X�r���$��(��	Y�����jÄ��ͱeM@V�P��&�"
���z���]�&��C��<���q�o	"e6��u���8h���é���=ar�8Xhp�����#��pH�.[ #K�����Z�D7����n9�<���9k��m�U8��{qB��n߻Z&C�	Dh�,��B#T|ґ�ܿ9,� P�N� �*�'�����Cg��(O�OW�����X�S�V�!0H�)b0b 8דTb$��
���?*a3��P
^,�Bf�/o�؃��4VRU�(O`����Y��S�FN�-�D�U�	ҖhdN?�Ik�b/#5p?e�#����VH��efD�[沍�A�{B�|t�@m؞�b#Jғn�A�A��J� ۇ�L�5�*%��@�$���>b�O�M���@�>���I�S��8H��h�Уs@��-M�܅ȓ��b1͒�O�Ҷi��Hm��A(�M:��]B�<}�b�()�AL>�R>�p@�=u����ɍ�����&|O��-cL�tH!CX� G\Y��U��Fa��$! �A��EH<��)
4k4�j���^�n�I�'%�e�"EL	�R	�~Z�־a�����B�&� �@4��l�<a�E]&CM��I��Z]� p���l��X�"&�9���>E��I�?h<�I+N\:*�$)AP(V��!�D�)�����̀���YzsH����	�)R|�����ayb�נD�6-HM��b�h�A$����<A0�c�j�Qt&��E�b%rd*N���Y{Ղ���"���	u��B�I�AI܄�=	�V�B�)]j�Op�բ�*��-�T(�ut`ق�I�;=x�3[�Mp�h�
'ݢ�
W"O�0*d�r[xxf,^ L��@S�oL�C�$��e@�d���M͵v�q� Of�)�*��	��y:��Z�7��YZ�
O�R�l�/lJ��yg�T<_���� ,]	lòђ&d�t�L��E�ʘ��I�7���>�4(R�6g|�v쁥L����̃x8���!�۲�&yp���,��U�-(�TTnQ&�֑���v�I" K��'$�Xv������5;ָ�K�$�UF��(fb�Y��	��u��@�B���98.�T6b�)�>�z`�!E�؜ �ń�y�e�=�:H!��<Q,T�&	O+P���#	Õp��A�#�B4o��4���:�4X�O��i��f��A��Ը�i�iH���T�)�|��:��,� ��T Qsɹ'ʨ�3��-�]�1Œ�u���s�'K�l0��M�R�sW�_"k�<d�u�0l���	�������	Ǡ�S�U 3�\SP�a�T��c$��)��X�f5$��,=Al|�ד3*����Y/dj\��#� `��%��2����4�{�"�>��%���M+�����1�G�~���a!�ɐp�pi��G�!�J&H=$hɓ)�Yl���n�tp�x�DC9��е�� k�`PYW�	]Ly2M8xl�"��%/�Xa�6!ψ�y�'z��KW��.�
��{��`��S>e���q�x���ϖ��OTY4���e^�̙3 ��Rظ���'z��1`�۫iP�} a�K�-X��HE&��b�#J��2�%��\��h �U�>�[���>U�2��Tb1��'�4��$b��|�)��ҽ!��K����<�Z�ɅeB�L;����yҌJs�xg��Y"��Ch��yʸh���w����U�ܚ0������<�[�$�@d�ǌ.+��pW�{�<� �� 1	�E5:��kV&kKMB�bXv���Â��pM�6��%F*��?�0&�;O�4Q�M���Q����J�� �iN�u�:q��5��-Ӂ�Ư �ba.]4����$c����a�7�OtMX��?W�9��*�e�c�DU	E���q3+C�*Nd䉂n��Oj1X�*4(�`i[�H�E��'+�-�W/R�<Ȕ ��Ŀu���z�b^�~�2%�����F�S׏[*�(��I�kF� F�o���t��( WpC�I0`��3��.dB �u�\UH7-�v{l�����	�$�K�� O��5ʏ�8*�!���9�����'���@@���R���[���r���~D�5�1��)�%��
O���AZ1O��DA�[&^(ꗜ|b�[�%\ �lO+ �ۄkt?!ɟh9�F�ǻr�F,��@�D$�"�'���J�-�#%���i�k
9�N���d��1Z���'�j���*Ԝ0�)�'d��9B��˞S�Z9y&(M��<�s�@�|��"?٥�1Dn��?���eW�iB���ʞK������<"Κ=,q:�;g�Hzg�p�E�� �ɧ��d/*�p�J2A�6'��/
���'��`h-I@�IO�`-�0\?� g�\�[���[��"Uh�JLٜ+�$���`Y=7�N)z�`V*WǞűJ�"~2E��!_��I��O�	]k8Y3CѤ��d�5_@�*S�[��?10-[��y���D�0���i>e�rꁁo}�� ��C� 廐�<�C�8}ri3ԯ"�EJ�Q���l�-CGE�� #@��P�J�䟳w^�Ը�ω� sR���$ʱ�^�g�.,���4�Ôp^��FőD��EJ4#Q�)� X���U+2iP�'Q�Y��C)\��0C%B�|o1E�W8�h����O�<٧AU�f���Ƹ
]�H�e�;h�SrRZ1�<q&E\v$2ը�@t�''�	����bU�͓+l��۳d�4�Pҟ���(֜%Ӡ�s6���4ͩO�S��S�O���*��$W�h���*b�U	��O ��@�8,X� �'Fl���	� ��}�#%s�ـ�%ۺb�*$�LCyB���h����L�pX����H
�^N����ޗL�Baq!q�;�%���A�4���d�O�ūRI+(�$02�ѕ:9Q�jB�G��mh!(H�@��M�ާŢB���`��W�iZ�ŃB�cmxH�6 �+�t��(�	C����E���
k^�$�擽R�l �GG>#��������>!�h�}s~��M�>����)G4F���-��dJ��؆$�� Mt�<Y��ԱQ�qO�>1�F�c�Up-�=W�6���ɻ>)p/�j��BO>E���U5C���0	E"B���S���y�ቀ+N�#�(8Њ�b9��8Ҏ�7B?,O�ȩ��[�F1�G@�D΀E�"O|�ZY��Yq���J���yQL�RH�`�(y���1#��y��J�P@,�V���BI���C�'���b/
L�XX!�<=.�A��'4L��ѤqR<�$i	�,�N���'.�9h��A�'���s%��%���{�'>�8��X�C��mr���y���'�,2����Y��`��{x���'��5���ɾ<��8��X,�as�'-tJ&�=+֘�r'�*�8}
�'���s�N�O&��9��*1�1s�'���%jF.f�<[%%ӬS3Wx�<�2��'>��`"�ˏ8k�$�9���k�<1�C�9sT�<����jS�} ��o�<�Ң]�n^H(!�V�E�r � �g�<�0,��D����)N���أ�'�a�<�U��y�Qj��G�G�4���I�V�<1�Y�FYFeK�X|M�)"`�v�<5��$h/�B✬��D)m�<�2��3�ޝ�t� t�Y���L�<�R䝦C���� ��@`�M�<Y4n�4}>f$�:$ڰ���VJ�<9#Q$F@��"Pm;}�6D�P
HF�<�F�\=�RiQ�A��Cs�d�т�@�<�ď�{��;F���/l��rI�}�<9�#�.t׌h�s��H��T���z�<9b΀�NTP�&���YÖ�xc,Ki�<!s��#�|IPB�S�9��� �b�g�<I���a��Q�tU����kVb�<� ƥ�������g���(9�&"O�� 䒂B$���G�z�(��v"O<�27��V�Th���T9���"Od�B��P4J�4���	�N��15"O��xr�|tHQ��gI�#X0Ԉ�"O`IQ��3N�� "�ػJ���	�"O��pF�W,�N� ��ȮI�0 "O�)9����&]�0㓺B�L�*�"O���¯֝9v�h��"��X�"O��R��B4C�\�3$�)K�����"O68�������kǤ�����"O��ĀX�{Lm�씧z��i�7"Ox9J��/�|��ō�9Zf���"OȘH�g\�l�� 
��T�xF�l�"O���M�IH^����?�ؙ��"O�T�%��5�]b(��F����"Op�!���$!��!��6�|��"O2�*Ě>%ˆ�Hŭ��O�\i1�"O�db�eD�uk�X���.,k<4�R"O�pz0�����ȫSFT`�&"O45�ю��o����d֮Og^���"O�LpG�"L�9�"ZtS�`�B"O���WY?��Hd�ѯM�� �w"O(eKÇ�	<!CR�پB����@"O�H(��
�W*f)�e�8a��A�"OB�!�߁7m�=��EY�}\�=�A"O ��p�\š"���05bP��"OE曔p%��i��N9^�#�"O�4�$�E>K�,"d`U�P�|hv"O�+�@��n�(��ˌZT��"O\8�6���R́�N��#2ji��"Ol@�q,%%.���m�?<�U�"O����f9<��`��ܒ��ZC"On��� �H��GN	5�J�t"O������R;�=8�L�^qT�q�"O��6����	�)9v2��"O���eU�STthA����nd�(�@"OY�e�6_�Z*6̆'*W���"O��2F����L�2(C�^�H@0�"O��*�#� ���(��W�����"O��x��
:Հ�"s	�y�r)�P"O���ϋ=g|�<�&�Ռ��I �"O�0i'g�5K�FP#�
�?f�4y�a"O�T�A"Q���Qg��bV:�W"O��C�9�p�1�fG�Dj��5"O����aؤw�^Y#��ƱA�q�4"OF���(�7��\���$q`c�"O����g�M?P���AESiZ�""O<����N����B-�9C��c"O� ��ڑ鼬b��=Jt��"O$��է	<��`N؅i9���F"O y���J�p:Sʟ�a,D�"OrDp@���$�K�l�j�^� �"O��* *_�����+X�l�Y3"OL�����T���`ɕ7�޼`�'X$��F�[y"/�d��@ЃD��n�&����6�yr��jP�w��-4�:��_��'
tb���
��?�r�/��i5(ĸ|0�p��"D�Ly��� �U#VɄ�R@:���t0���>��C���d��6o�|�1+S+eNZ�z&W��!�23!�\���k |e+�	�&l9�"K'52ࡪ�h/\�V�D�F}�S�!�`�(����#<����P˞1A���ٻ����`��^�Z�*5�L��!�Ēch���t��,*�:�z�M[_�1O>�Be͚Y�"m ��� |hZ� �1�p�H2�����	�"O�pY2��:I�(xZ1A�2�\uҰ��#����L����!8�g~�F�
re��ɒ��F�`���Q��yrgK11�Z��b��q��}�,5u�S���&n����=m������()��ϲ;2���Ĉ����[��Y��~�l�mz����+Ѯ?����%N��y�BN4��1��,ه|I�R�#��'�T9�#*�s�?���f@�wN�h8�oC>�� Pf'D�D��6�4�G�/62��R��4Ab�%�=���>ae�@-!�"�1���@0\��)^]�<	����o�X!�-�(DtT��B.�s�<	�!%��u��h��R���x���w�<� �ݜ���B'�\���� 1��s�<i!��"2v�Q�_[����f�m�<U��-T�	s�̆�_ՆВL_n�<	�®x������mj���'^M�<I��,IP�����K�$E��[-WܟĂ$�	�X�����I"%t���!͠)��)3�m�8,T�,B� G���'G�O��9�͋�.P� �	�-WH᳗�L�e��Q�2*Ⱥ(���^��d��ɚ!��͡��B���.�H!I#�ir,0q�%Bvi"�U���>S�;V�8��@�S(1�dx�!�'>>D�d��0|L�H��3cM<
:���$	;���$AM=6�ك�S�����<� �+h��� j�@��t��t�ik6���D[z��"~�Geё�h��^`B�o��xV�`H��P��|�5�'Ί��p��?I>Y��Ù,!J
�BF,�m��K����~�4�a��Y$ٲ�M���'���e��0��wd�D�<�2�E	C�,e��+�'1�|�b�)�R�`4.S���q�6)
r��nD�D��)��IYL�+|]��0nT4�뉃n��a�����V�nl��rI�?4ڡ�d�E�~ݸf���,�<�'|�G�,O`=�a㔱��EB�i�����D��PP���+����)��P���`�c�$�Kҍ߲.�I	AI
59BM��ɻv(�@l�L��(�ߡz��������4l��8�Ӝ����	Z����t��.K�+4"-�DT=VE�y@f�6D���ׂ��"Ebi󵌇dhT�@�Ki�X�2-o���ӌM
�r!a��o�	
��Z�r|��2-F5p���ءHE:��{R�͍�P�#�i��qy�@���<`'�2a�yy5��%HTH<���$ю)� �P� ���GDJ�'+&]��jȶgL,@�~����	`<��Pb')\d�I1��|�<�ƀ�.X�P���%'�0I�i���%�6-�@Z��>E���ܝ42L� �P�-��a��D�!�d9��('�߷v��E8u#ܔC��	 |�Ή�סrQayrhG;�l�q�AH�I� ��cH��<y�ȿH� ����L�n��BO'~I:a����P�j%��KP3U,�B�	[��ze�0]�n�B�;d�
O���ՊQ#tʢ"�S�\�9���^;yt`i�o�DT1#[}~!��W�}����V�h�ؘb��
Up��׌_�o2v��F��(sf<� ��&�$Ǹ��E��5QrE�)myz]p�
OYFb,4o�ؙ��6��恈�,��s��h<��9��S.m�yr!��EU��K�:�꨹E����p<A��,"�P�����U�@�|ю�ۖ$R�S��A�R�=��B�I&A�\�"�5p�x�����8\-f�'��Pգ¨t�PĄ�ӓ&����Ԧ*�p�SA�P�|�:B��s�e[���{�v|y��L4� 4	G�>}Ҍ��m�1�}&�\�1��.FT��̈́<���En9��8��Gk�����^�����?�l���[�\sa~B�V�BF*$7d^]��K3nF��p<���\znzI�2-?ǃ^��"�X��C	���7��r�<�t�߁2B��BC��x�k3�YP��?�x/1��O����(1L��
�,m�L��N��'"O�r#)R.X� �
#U�pZ�h�*d<%��L�	�&Y-p�r�3j߉b�0Vn2D�D�`4r���Z��˦-;�0D��(�	�����BǱ_ٴ��1D�����?�ht�B2�l	hs�-D�� ��В#�rs�0���\6�I�"O�U2w��`��I��/R��;q"O4��P�2f�8�)�$It�f"OBI�MP�F%���F�+b2�zg"O2��S!�uF����Y*u�2��Q"OVYUe�7��XcWHzp��"O.M�S$��{zI��"-x@��"O�H�dlS�h �� ҒpN�zd"O�!�\t Zt�ۘm5�ܹ�"O�iA�* lT �{B�A�]�~��d"O��t��RP	�1*�94 Y�"Oj䱢���(��I9q��%HM��"O�A���)�x���Q|:�2��''�y����!HlР�N�.��(S���+;����J���5�
u����"� h@�F}2��=]&��@���H�cK"4j���D��
��v�!�dM:�qꓢ$g���&)��X��d�'</$]JF�>��)�ӐY�Ҭ���D�[,ݺ�(�-C�q�I^�2A!�$G�|Ǽ������Q�r`B�܏"I��W�x͐$$��G���O�Q�2�$��S�4�P-�Gg��n�0�h�e	�>�?I� ����U*T��j9%BsG\w��7h�-&͑�C"5r�yI�ʚ q��S�O��-(� wZ=BrFe%J�PV����JQA4n,��g�i��@\U���>�S�jX�X�`����·M�@�����<�U�>"3A�*,O�y�b!m��r� 	z����1O25)r�-p^��g@;z�]�1���u�$0S��%�\��hV9$v<�Tʖ��I
���"ɀ���dk�(�qpYB��2ɸH+Q�h�9@��s��<����5��Xa�����?��L��@FB��A�3��!3�,��*�i��Ւ|.�2ڸ��S
'B�A"E�����EM��O!�h�Pb�'�Hd�I���)�P]�3Fkh Ĳ��Dku����'�:\����� �Pϓ/��9�M�f�>�xD!D�w�(*ƍ��Vhѐp�<�Dh5`Ny�",O���FQ�JR.�[��9�(�:C4O݃D��Df9�C��.1F�|��b��_d���S͢3�DB2�	������Fɣ!�f$	� �jR�CB���墘
��)�4�Our0�Ƞ�T���%3;D|nZ@��ѥ��M�i>�a I
� �µP1�[�*_q�cg"���81��܊Q��;�8�E�>-�&@����~/�}�Bf��p���I�.������o �	c�Ѽ5"da�Y29
����9q�����S�OO�� ��ǆ=���)bM� :�\!
�'u ����>C8��k����HJ>��+������"pv�ڶ	F�C��h�G3!�w��� ��Q��"!�d��_M0gi��u�s���b!��A=�.�2Q�D[78d�!�''2$0TA�&l�r����f�NL�'<�٠��~��S�C��[lj���'�
t�ENB>=��a�����hP��'�t|�2l�6)ԡ������'@�))V러�
�C5T5qB��'e���Dk�=J�� q���m�Ft��'���2���s*�@�k�v�\�)�'�T�(��ع>��Q;��Ҽnx�ē
�'�8
������3�>b :�Z�'��y�+��_18����`�( �
�'
��)�uy�x*��?d��
�' �q��L�9Sx��2�M�/u��5�'
2�s@�;ݜ	!��0f}�Hp�'Y.��挡',|���ӄ^����'��A	�D\1� �o�Z2H<X
�';�)��b�-p\�;�`ȇP�ܭx
�'t��qq(݀w,��4hE�J� �
�'+�d3 P��=�c�^�A2<i
�'':�{��F�G؄���lߎ;`�
�'sR���b� Z0��c�:'ܭ"
�'[~��4i�=�r b��O�B���	�'8�tʴ��]V�
�H�*��]���� $y��ʜ�==����ߌ:���"O���GC;I6-�2��c��h�a"O.��Qaʬ'����B�NV��Y�"O�XB�к�Җ$4��3�n���y�G~�(�kY�p�
@�����y�@�7q�x�sP��d`lI)�K��y�LՅ	xL�x��!N����� ��y2�8qu�Ӕ�N,(���HQ�G�yҫ��/`Jɠ�'A�r20Q"c�ن�y���VL����$'����AW0n����'?��<2�b�/vQH�V�J�O�8$�Z�)�@2X�=�e���,� �K�>qF��'X�E�|rN~�qd:u�vQ���CTL:�$�Z��]�J*���d�	��0|z7eX>�����)P�����Jn?�����?J�*Ul=}��Iʭ>.�S�F�c�%���Ť�R���enVD1��>E�d ��R��Z',-�<x��(`ڴ`��uجq��B����� g>����!REh���nK�t�s��
<�u� &o�D
';�*��#�~z���A}�TH8��/:>m�Ѡ���@��s�%��Ó��Q^?�G��&�O�Ι���4v������?�4�܉�,IqG_�(��)�=�2��#M�`g8a0���j�,�c�m0��f�S���D9����b�ROS>�BG��� rB�_,W,a�$�n?	&Г��L�����M)���
WbY�oW��T�q�n�"[ة�_�t��phE�G��I%�i�|BGl�F|O�Xt��v}� x�V'��yp�e�}�ӺK��jŻ��c�*�$���b�Y��ڝ��d�f���}��o�?%��ԛ�������BZi�ɳ0+��[��e�����o)ڧ&�@l�q,N�8�K�$]���b�Oh���H0�M�5�Yi�'�ħD��УI�$H��\�#����O:��ٴp�qO��x�Ȍ$�-��D 	�*�k�_���Dg��(� ꅎQ��������+��T�t&+�Ix���'j4ر�ƊH�t���_>n�(!%����"v�E��T(Shn0v:]�h})r���'^a��A���"Y����dT(7�-�O�I3�g+�\ p��@)wb��!��t����x��3��$��h�]>�ʚ'�^,��G��gr��g�[(o;$�x��?�`��}�����cR�\(F�t�Z*l�:�Ռܪw�h)	�W���T�&q*��9U�B�Z�O.0Ha��ΔEo Ӡm���f�#�@K<���d�+ӓG\�͉�[^6�[Èܚu@L������b�>Ut�P��w�f���*�<�[�S&��Y��� 9zԅ�(����Ű-!�=	7#�"Xh,��\��84� �$��� G�0����/i��i�i�D����xȇȓZ��<2��$H��AEH�%��-��c��=Bp��R4UMבA�Vy�ȓi
b��3���$�@���4!�z�ȓ98HрB>%�\%`�!�%b����ȓls�;�+Ҷ|2�e�pÃ�C^���j�b�	f�@�{W�y âO9A��ȓPJ� �� N9 9N4|�ȓW�`��%�(�\�˰g��+p,��VtL@�.A�S@��%��| ���(�1Ҩ ~K\'jBEH 6D��
႕.OP���NO�R�4D�Th�Y0A$�Dڥ��.A#���2D�4�1En9�$�v�}~jY��k.D�lJ�k�uAn�#&�R��:D���뉃b�`�y��ލo���#O;D�$�����>�V�2�%?ܢ1@E(6D��iհ���:��8;��0`8D�`Kw��Z�p�v��3A���"5D�l��D�� �L�D)4�A�4D� *�再JF�ф�?W,�(5�0D��CoҝIq)��[�
�C"O"D�B�E�<6��فA� d��d`#D�� R-&z��A��Da%���M?D�� ��U�U�Y6Q�ր�*�p��t"Op�(�
��K�T� �7Y�~8�"O�}���J(a� �!��2PX,KC"O�y�«ٷH�d�w��]񢘋p"O،�í�J ��m�5Sݜ���"O�|R��>a�D;�, �%ؒ�V"O�=0�C�K `A�7��m�z��U"O���CIE�!b��Q�[�}�L@�"O* c�˵%�	X��п
yz�R"O�E0�J�/#�"4�G�Di\�:R"O�hi��B�8�ΌbQD�hh�dc�"O�����'FNl�����M�n���"O���C�=?�����o� ���"O�d��\k^��Q)N�l1�"O,����(��A���J�H|P�3G"O�4�� �c��#�ًp��Z�"O,����P5�2���(FlҜ*E"O���H^y���C�U�J�"O|e���++���sv
�+$�C�*O�1P�\�R��X�DzJ��'Ӕ�k��si�`����O��В�'�e� ǤK�V�iQf�CV~q��'�t��'Kؤ(�����\�)W����'��g�C6C�(����ڽ(��Ł	�'��`z����n���%��R��[	�'sb �sg��g,�,�EE�Bx�d��'t�l(�@��$e�$i[�C�.��
�'I���D/BzO`p`TC�>�P4��'�v{1fZ"2����h�8.���']N�xb�DE�a)�ގ=0����'& I��FƖ��B�T7!&,��'��-i҃9�:=B2��ZX��'�	P���y�D�j��U�'����'���D�	5�^ ��w���'܈���e�#r�F��#��_��K�'r�0'���ch�*�F�O��LC�'��-w.�d=���!I���P�)�'#j10�]lIt�"v���¬��'� �˳m�wi��@(�A�$��C�ɐ^켘;W�n|�d���1��C�I>�41��V�t�z�B�=g��C�ɿ%
6��&ˀ�O�S"J��si�B䉾%�)�w��1ࡐ2hƽX�~B�ɐn���r�$}���A>P�8B��3=�JTpU#N[V������"�B�I�O.���Ĳi�䃃��H^�C�I(�,��R���W��-Y�C�	�a
� x5	L#
w^���3s�C�&p!J��Vİ�BC7_�B�;*�*�Z��d���{2��!G/�B�I4�L1���Ǘ^̜2�IN�hB�ɥ[���H'��瀅�"��0n�C�ɚ	d��#�P\�)A��F�.C��8�0�h�A�#-by{r���%AC�&�"	�u��|��<3����+w B�	�X�X�h�Lxޠ��):q�4C�	�:�V�Qt���m��ve�� (C�I�n��|B�� NO���5�X�G��C�t����vj-J�~�����4ƐC�	�Ֆ�6o_Dc`42��(r�C�I�C�N�x��ѵ�4�
�P8��C�	-P܀)(�H�6>����e"��
�C�:H��	�G�_*��`��C�`sB�ɀ*gF ��@�d L���:_R8B�)� �1�"�(4;�3�bG�p4·"O =� $�'��p:7�Y�Z�u"Or(r1kH�fClĳR�Чs����"O��c�S��r�p���|�(�j�"OF��SjEq,�� � �|�3"Oޘ�WET$w��m :W��a�"O�(Ӷ#�''��3K�(��v"Of�{�ث'���$�̕����"O���i�;S^��{�l�:����C"O�q��V!.��x�옽w���"6"O*�@w�x2,+%��q$���"ON���c²c\���D
��`"O,�S5�ǧBcz���*�2N��t��"Oz���. �$�g���Jq�"O�u�h�H��@	O<6�����"O�J�!�1��Yj�A^=��d1�"O����υWB�ɖM[ur�K�"O��+���kn�X�tB�2pXu)�"O�E�oV
I��C��!t�.��@"Ol4҃H9l���aN�=d�8�h"O<����B&���₆�	��"O�P�.Āx �a7�V$�+5"O>PꀅO�8[�h"�	�5�n��5"Oа��㈞u���P)M"�d��"O�������jK�m�D۷"O��[�ȇ-� J�XWФ�"O�QJA֟vZ��%h[�_7ʝ�b"O��@�i'%��Ap���7�
%"O��v����=H�� 71��ia"O
�QӀݎIbҔz1��9|��{�"Od<�"���=�F����ϲ|��Y[�"O��8�H�	���Tm�&m~b�#`"O�Q	�됺�2� 
�9bټ<1�"O���$�ȼ&z\$*b�Y Vӂt�"O���e��%~��r�8#�i:�"O�Q�Ќ�x`�и�G�`w��	6"O����`\�(Z��) �:g�j9Ӧ"OXY�J�@2��(��W�k�-�C"O"�T���F��*��	9|j���"O�* �Ux���RrG�Jk4��"Ol�z!d�*!�$�QFK�T�p`:�"O��:���C��*3�5��"O^��&���,����0�H@"O�m�1"]�Os�= �`]�_�pq"OP�V�2V�aЅ���0ur�"O�UP��MR%��RK�� G"O�Y"Xd\��D�%�>�8�"O��J�A��+�Z�Q@�ƒ/�@�"O����� 'L���%#�x���"O�`"��<[�F���M�yx�;�"O�� ��K#V!�0�A9je,�3�"O���h����pS�hL��R�"O*�Sp鏷�xs��I%/\�z`"O�$Bq(7:x�P{����2z�!��r����E��?hĒ��B��r=!��a!A{��.<��GelG!�$�3��`�žިa�`�ث.!�$>8�hc $d� }���!�d;^��S�N6.���Z��Δ!�$!S�Ȩ���+Jo��@��!��d�.�2���*@��Ű� �'�!�
(F��;��@�+�d�6υ�Q�!��K\���i	9��#�-]I!��6T�8�u@��d1ΕpS�V�W!�� ~Uj����[��-{F���,hE"O^����B�p% )y� [�T �=(�"O<|��B�)
:m��`��^, ""Oh��u��N;J���ԇ6oĚ�"OX�c��(�"%��o/q�^@�'"O�d�r�N�Wʸ#��1�};�"Ov�Xq��gi4ŚG���3$"OL��e�!�����AG/`���04"Ov��U�yhd���΀]!����"OL��񧁃ytT �$g��*!>�"OL�8�G�#AN���`�U�in���"O��J�+B�����˦r�V�a�"O|�ȕ&^%�����ʅ�XΌ�H�"O�T���pSn(k����q�F�S�"Oj<��<YP����Ӯ"��x`"Op����K�/��Ss�\/7��"O0����6>(:�K#��?z,���q"O�P0�Dtf`��bPrl�`"O�$��`A2"�H���P;C����"O��C�`V!5|�(�G�9� 5k�"O �r���C��tO��`�:�"Oz�����@ hUo�s�9��"O������1�0Nߚ�٣�"O���0�LhA2��˨(���`"O��RBO�"赹�H� �Ҡ "O��h�� �c��x�`�2����"O�hʳ�N;H�j�Hg��$>(�g"O���׿d���3K_)�~���"O���1MAR@�jE�U�vA�"O�Ð��'Kz����14p)J�"O.9�l���A�k^4�Jѳ�"O�%��χGs�X��L�:ռ�+�"O�"��X�)�(9%+(,����"O�D���AB�=�1�Ʒ`��"O
�s�FD'B�������I�� ؃"O�T:��=S).���0 vrUA�"O�he��N�n�����2���"ON#�V����a �(�p�T"O�@hwJ�n�^x��H.ndʀx0"O��`   ��   N  �  �  D  �*  �6  NB  �M  (X  �a  �k  st  �  ;�  �  Q�  Ġ  �  H�  ��  Ϲ  �  l�  ��  �  S�  ��  ��  5�  x�  ��  ��  t  � 2 �% s. h6 ;> ~D �J O  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h%���븧�O@��1�AE�8�QP��Z�	$��
�'q��&װ-��J�gI�H�'|�仳n޽�j�R���*[�����Z6����C�k\���T�[H~�B��D]HV��
	����2�W;���'�^���d,�'HW�ePU�K�D��!&I�� <��6���$�8x
�Q{�/gY���=��^�б3�)�+("�F/W�4}����ys���Lס8����R�%:������?��.ߥR������'/�F����j�l�L<�@��=l�{�nM%VZ�����i?���S�^
p�Ė='�:���l� C�I�HX���4������ݽ}z�C�I5n(]r�'oϋ%P:ӣ���?��Ob�"~���/Xr(+��ˀ*tv�	s�E��y��]Te(���aE1#ǒH��f)A���F��4�$�͌]a2u�0��@���q��"|OHc������Ţ�\�?� ��>�	�v��yh�5��dY�eݽf&:P*�Aޚ�Px���3:� \I
�<I�y6C.9�֑���>�4�*lO�0�±�
������ڨ����c~�>q-OT�	�F��pa��G�z�qf"O|	�t@1����v�K%H�J���"O�كh��<������47u�HY��',h�O�i���B$;��hu�Qzj�(�p"OheБ������ �_rW�	��HO��/od���
b~t�`��~�B������*� 5�d�h�!�(ǶB�3L���a5���Q��?�RC�IM�R��&l�����G�g�I���?	r䐃]Lx q"̖�G�flpc�C�<���+��XuF�/�}����}�<��){ji��eH�T�H��R��zX������ ���J��ZVvE�$���m���Q"Oظ�AQ�W�4!Z��۶7^*8��x��)��!WI�8�Ȏ< �����)J;JW�C�I9~@ h�)N�̖��臰T$����q��G�y��N H)�ݨ��ב5�b���+\܍8�X�`�J��0l`2�D|2�S/����gN^+z1jE��>�C�	'Gp)��@������;W7nB��+O��Qp�L�*�m�)�~�BB�Iz7�l�E��BMx�{����<6m�����'��\�Aބx�8����ؕ2��H����$�<!aA`}j@�'"m� 2�U�<�4�C>y� �R��ČF�ȅ�ULT�u���O�����@�V�:a���?�X�
�'�` �,�.��ujw��0s�Ԛ�'�V���*�^��s��Ŧ,N-+	�'g.%�$S6*i���Ԥ��]<h�'-�$��WC���R*7Όq�'��T{��%SZ�sE���ky�m�
�'������Ǝ1&�e	ˋW@]Z
�'T�,*bA��XS��ۅJO�X-Jt�ʓ���'ćMf<�g�L�{W�hm�q��������_��Z&9��	��yR.�'-dR�tN���86n���y��֎
��i	��VX�5����>��O%34IO%jC<tY���7�����"O��b��R���F�E��X+�"O����B0N}����VJ�rLA�"O��蔪��.���Dr�x�!�"OIK��"��})@�\�8� ���"O�a�NP3�z,jtL�3�����"O ��E�� �%쀗)e��`�"Ox0 NĈf��PT��C[t�W"O�R�®7ĵ�Q0W�!����$�S�J�r�����g��8pvH�^�bC��]�TI�dcT�Y��T9RaZ�l������O.q 3��(b]�$b�F�+0�l��"Oz��a�?Ml�f�<�4�'�'v6���e}�p;�CP�R9P����!X��C䉕EǾ��ʱ�B�aH�@��C䉃E�.����,"`���Dfx*&��F{J~�g/g�֕����x�hZ5�!��W/0�SLݡ'u�Y!�ꃟ�!���6��3J�A|f b�*��;�!�d�R��e�R�e���ў7�<�ȓ`P��g�sl�!�$�����,�ȓn{@�KE���RF�$[c��7��L��V�v�Qr K=�Tsv̆�VTBm�'Yў�|*�ʣ4
�#2�o���Y���b�<��C�-jM�#uƃ>Je}y�_�<9���/��L��� 9U��mA��Z�<�`)J@8��"	����I�c�{�<�1��*c��$ɧI>.)��a�Fc�<�s��mSA�һ}��QKS��(�<0J=ږ�a��D�v��)�'�C�<i&Mܫ���8��F�nI`��C�'4���S�yH��q�#W�=0�t�aȅ�<C��'�p��\�My:`�v/	�F� }:�2P��ۤ�x���'l��qo5Ttcp�!LP���'P��(���)GXe�g���F��(H����I$A+>��M�"�&�14�M�;m�C�	�b�b��	64Qy0c�.z*pB�t؆Jׅl<
����5L�6B䉮K?���#����<�ĊE�c!"<��S�? 65i��C�(�@v�J�c~��SO�၅��U�ݺ�Ɉ"8���@������H8�� �,�.|
����&%6}��	9�O&pj�''�XK���)061��B�E�@����HO�ԑĤ�P�Uґ�נ\\���7"O��KTh@�3�>�h���tDB�(�0O΢=E�Ԩ	��@z��X�i�̱q��ʐ�y�i��j<��P0*X�]����d������џ܆Qcj�: B�?5Ć9���/������<��k�=�q
�C�%�_�<q��g��uc߿hŌ�SЄW�<��Ƹ��9�O�J@��*�S�<�/S#�6-;� V�pZZYP�lʟ�G{��)O����񀄕T��A	߃r9<B�ɣwZ��v�UI��|[Ь	�(���;��	��~��hO@���@ph��B�FX��_���	�p�*e3��ԎatX�KG��\H�|�Ĺibў"~n$>q�lP.��R�j,�0DF82�F���[)Ӹ'ư`�'ǩ"gD�"�o�>_&a	�O���d�-M]v�a���HS@�4�a}�>1Q�E$��0B��O�!H�fX_�<�����k(�!�K�N�r�����u�	���?i�yrf^�C�T�[���.t�&�Y.��y�'�{ir��G'�*k��	�P��y"���x �'�ec��� �y"F�)-��T�v*�ZRݣS����'��EyJ?-���В}��)�j� 	z� *D��stk��}��ŏ�Vd�X�$���(O|�}�U^�*'��
q���2Ç�" E��r|�p`&�z���D�^*{W����?ƞE���) �ȕm�
��"F?D�Tx�Y�OϨ���B�}���4�(D��Je�A,��2�E@�:ۨ]X��&D� 	�*��w��2��%��9Y1�1D� BC,�2��͋p#X�*&P<A�O2D���ڹf��b�v�$���E1D�(�Р_�W��Й��&c���6e4D���r(5s����0�9b1rE��M.D���V+�,m>��9a�ʱ.�&=���*D�����؅6����&��"�N���'D�p�0��62,	QӦ+�ty�F'D�hГ�ة8-�*��
t�4�Ѷ�:D���4E�xN�y#�T,n�����8D��AkM�C4a!'��P+��P�$D�$)���<=Rtr5�*P�=D�\H���BXp�`._���4�9D���EeͱtV]��Y"`���9D��0�<��H��ω�t*�@�k6D�34�ճ3V�pp`�v�S��2D�H�l��X/���FA}T���#6D��P�+Oe�1��GH�w���GI4D���ܢ}���@qc�����H�a&D�hs��� "n��DB�5��L� '%D���F�%k|����J�O4�d[�$D���&�'��`�玏9z2����`!D�t����Jx���`��S�����$D�P����%(; �{�ɀ(<X�4+��$D����Mk䄠�I�H��0	� D��R�.�O�P�x�g�ZT���?D�\Spʋ�"���ьh��z7�?D��ض��'~�jX�a�:'[�I��N"D����J��~]�i�bܶ����"c!D�dr�CP#Y���y2�Y�Yi���� D����& �TCvA�,����2�?D�� �Q!����Iʄ<E0�!�"O��B����<�x�Ci_j/(��5"O2p�DY
q��QB�fD�.���V"O�0���ᰈ8bl�<* �q�$"O�Ļa%F��d�������B��'q��'+R�'�r�'�'���'���m�4�J�0^��=���'���'�'o�'�r�'���' ���t�#zm�)1tL	�H�P�U�'���'4r�'5�'���'O��'�KYm�%5���;*p������?���?���?���?a���?���?�S�,vZ!ɄS�tK�1�`�я�?)��?A���?I��?����?���?ᅀE�^��������C��H˔j�:�?1��?q���?9���?1���?���?��BQ�/�����+[D(�W����?���?I���?���?	��?���?��@�uC���g�&m��%��-�-�?����?���?���]*�?i���?�C:|@�
M��0��C� G>������?Y���?1���?���?q���?���<�P�;*�������8N
���?Y���?a��?Q��?9��?�����}r&�A�6����H�������	ԟ4�����	��l�	�D���#��+�y��G��2,x��6k�ϟ|����t��۟���֟ �	����	͟Dy�Z>�(q�,��F�֩XRHП��͟t��˟��џ��I�MS���?D*ZB�dѰ	�<#�h��o�6��柈������R����n�+`��$��$YCf,�� 3b�$�D����4���O�8�p�	�,��p:���}F���/�O��DZ�a�6�;?��O���I?����) ���wk�b
��P����'�^��F���̓8�b�:šګU�*�Sb��6�+j�1OX�?1���+W-�:�|uУ�](�vE�"ʯ�?����yZ�b>1��]����HF���ìG4%1�ѣ"&֞,��t��y#�O`����4�"��R�Q����!�"|ђh�¥Gk�D�<AJ>���i�,m��y2"%9*�Q HB�5����@C�?"�O\<�'B"�'��>Iਛi�e����O���Ƞe�M~��'�xd��C�(��E�OF�C����+Aǯ}�D�kF�ȥ-\NЈ)O���?E��'
!�v	�/1`>�c'a��E�ࡘ'��6��G����M3��Op01��K����y�Ӌ�� �'/��'��K��CW����@Χz���S�^Lze��)�!�d@R�)4�6�&�D���Ϙ'�<�ȵ���$V���S�a*Z@�O*lnZ,������X�	K�'~l|�ǂ�1چx��7H�<)2R����49R�&�7��IZ="�����_�y�v��eB4w�� ��
9	Hj˓�L�S���O. �O>q+O\����D�}��@��YVܪ�)�'�j6�.2aT���_v��/@j�aA��F)f���ަ	�?�qS�d�	ئ�K�4e�	!!�)���/+4L��z���+�����$i�� 2���)����R��EC,������_oQ�,#E4O�����!��F��5I� ���d�OR�$[ߦQ)A�:�%�i��'��(�G�Ϳ-��5�e�"n�r�U�|b�'�O��᪀�if�iݑ�G*ˌ%��M�E�R��d�&,פ���������5�	�9�d-�A\�_��=b!i�6P�8"<Q�i؜D���'�b�'�哂j�~X�$�	Hwލ����+@`�1���̟(�IU�)J�o�t�44)S�M�$d���U"E���q­���M#']�擐n�d3�Dۤ&n����K��fe��
],���O&���O���<Y7�i���S4�ø7�ܘ�I%	2�	���E��ɡ�Mۉ�I�>���i/v�pa�۲Ag��*1��(~D�dq��gӄ|oڃ6r�mK~B�/AD����.~����	�#x�LڀF�<\����qy"�'�b�'��'�2\>��P�k�Ұ%���Q�8�����M������O��?Q����cGA
]�	Q�H<! T&�-�?�����S�'t�J�ݴ�y��V-'~�����Dl�x�e>�y�gZ �p������ĭ<93eܕ#�(�Y �^Z�� En���ܴa������?q��4�2ՁQ,�]��,Uv���>1��?�O>��O�$^��Q����>`!e�MC~�N����s�iݺ��F)P�'���MCz�Q�JK a�8�a�)F�4���'�b�'����矀iQ�N�꺴hA'��js���s�	۟ܛٴ:Q�a�+O�m|�Ӽ� ,��t�Ud���ۥ��<��?!�UO <�4�y��'$b�j��?���@�-+�8@�%M�;�����/��'��)�3��/WkF�9��˞������L3,I�%��!ۢ3���'g���,��C�(���2�иXq�|���>鷷i�7M�\�)�S*��̗��l�,�.w��{7�����1)O|��C蝻�~�|�^�(�R!N�]���wL�jC����b���	�d�	���ky��|�@��#-�O�\�lφd־H3���"�F=0���O�XmZW�8�I��ɕ�M32�ӼF�扡��s����5K?Qj�4��$D�֤���'��OG� �B�(�ы�#D�\rp�8a6O�����E��	)S�� �q@6�T$U����O&��˦hq�*"0�i��'�\�
�IE�$f0�Y��݇pE
��%�$���]���|��*���M��Oع���$���-ɒ@FR� �nF>!4E��r� �O0˓�?���?	��X����OW���8�#�6%5-���?	,O�l�?"�$����0��P��gۮNs���N?[���H6�P���dNyb�'ڛ��9��Ob����3N�:�@ ��7=l�� �b�(��}���1w:hS�O���F��?���-�䑑4��H:�FPK�����b^.t3*���O0���O���i�<�e�i2 �S���/�xғ&�	*�#(N�E��'x�6M �����nӞ ��� =gd(��@��@�ljT�J¦�46��Q�4�y��'� �8c�?b�O�T#�C?Z��ٱ� 6$���V=O�˓�?q���?����?a���i�R��hroĻ*�z`��!p�t�����B�$�O���1�9O�emz�m	��M����+�Бm��3�J��?Aشxɧ�'@Ҕ�Q�4�y*]�\����*["<eV���*	��yB�����I�~��'��I��|�I�i����|X��Ӵ��?1���<��󟠖':�6m6\��O��D��l���C�˿z�=p���J�j�q�O����O�O2��Wo�a�f��`$�-���%����a�H8n�o�l�'`� ��Ɵ䫀�ߌ#��%[Մ���y����I�����ٟ�F���'� ��Ba40�;a�S`�L}J�'t6���R&��$�O�5mF�Ӽ�w��+2ؾI�sL�e:��qD�n?���M��i���i�i~�	0
�(r�O�\5�5��s�đ�,�>���ؖ��ӟ�'��i>��ɟl��ٟ��	�X����MV O�4�3V,I>K�d��'�\7��MH��D�O��D1�i�OB���#V�?�4cO��v3VY �l�h}��'�2�"��ɑ�y4D┧N)sa�!C�	6	�r��@�V�L��	lB���e�'�R�%���'T+��-=~8WeQ�Y��(�HQٟ���ß ��ٟ��\y�o�O�EXd�'�Y����[{�1A�_v�VD�'L�7�/����D�O ���O2`�#B��!̍72.ހmS�G�=&B7{���I�m��4Ȑ�OI�����,��Ճ/$�����ͺ1���?Y���?���?����ODdP�3ƀ�(sN-p!^�:<��'e��'`�7�� W���OҨo�X�	�2:��3 j����䊈a�&���	џt���H��m�<q�OT�@���ͪ�px����A���#%*��J���"��<���?y���?q3�ȇv��*�J�(�d��-��?�������i1����X�	֟�O���Zr����I�E�^��L��O`��'S��'dɧ�4�'�Q��F�k0pPP�K�Mk��{�-��8�d����i��ʓ��4����$���T	��� �2.M&�������	���	�b>Q�'�V7m��\�e;1�Ɣc����B,COe8���Oh�Dæ��?�T�`lZ����>g��ʥ���L� R�x��oZ� (�ls~���£��?ɥ���!���7Ir�t	) �׳�yR]��������������ėO����ЎΛYdhړG��|�*���o�b a��O��d�OV�����֦睨8f�8j�	S�Լ�$��(2���4'̛f�4�4����쟢�naӒ�ɖK��Yj�'E1��$s�χ�I@l牤6�R0	��'�|<&�,�'��'��R���*��C�k����'�2�'�"T��jߴMex��'�rΕp�R���� Y"�����~�"�|r��>���?�J>���$j�]y�čy1�aŔ�<	��ZO�A���M��Ol����~��'�jX2��9(T	�2�ܟ}G�Y��'
��0$퀐\�X�8��	|l ;1�'�n6mD�Fz���O 4n�x�Ӽ;+�!I���E
�6�d��3�[�<���?q�A�N���4����#�?�* ��-`h���_%��c�z��_y��'���'Z��'�B��2m2j���"�M��ӮA�T�I��M�7ŀ��?����?II~���+��ǂ�:I�]��H׏W$0��aV���Iퟰ&��ٟ �ɽE���$�?U-z�k��E]&llj�&�䦥�-O��Bb���~�|BY�\�V��<��#��S�(IJ��۟���\����Sfyb�rӤ�r��O��#�*�|;��O=r~��b��Oh5l�n�W@�I矐�	��M4H�7�TM[ �ф ��t1(�$Zb�;ܴ��$Ġ�*���׸O���L�؝�7
ة�|�!���y2�'���'���'��ɔ�a��#��%;�@T(D���[��O~�DBɦ�ɵG+?a��i�'���4	3es؅Q���)l��xb�|��'S�O{~k��i��f�(i��$ǂ<V��U'?��	1�ݯ(M�� �$�<ͧ�?���?�Q�J��(ٶ�X!}��X��_��?I����D���rpb�byb�'��T74T�'/M0"Ģ<�@iA����m	�I�0�It�i>��I�,��Ƨ�h�b�iTmۢ3�^�ʂh�	Wl���)<?��'A��$R���K�r���@צg�v�S��=+B�hz��?���?��S�'����禭*�,N6��w,�DبEBݬ��H����̹�4��'i4ꓩ?y��֟�N�K��6H����ڹ�?9��i{��"��i$���O����ۛ��G��� n��Pb�I:IC%�[?�6 8OL��?����?!���?�����閭yr(�ׅ�"������/�nJ�`��ڟ��	l�Sڟ�����[�OA�/Uv�cq�H=o� 3�g��?������|b���?�gH/�M��'�����؁o��wn�9U&�X�'���9a�z?yK>+O��$�O��꤆?Z$�.~���Z���OF�d�O����<���':R�����?���M_q�Nf�|��	I0��t�����>��?�H>��I�L�t�]�8�}���Xh~R��0��
����O�����82"G�!��Q3$��-!h� ��Bk�';��')���ܟ�[Ƭ��urv����9#2�9�����<�޴	d�8���?Qg�i�O���m�����6RR|A(�`[�`�D�OP�ĖĦ�Z�k@Ѧ��'�$TH���?}õ)�~h^�CCm������~��'n�i>��I�����ßX��-�h��E� <� �+ClY7\N��']�6�J�T��k����OВ��$P�&� �Kr _�Av����M6A�'y7m��m�I<�|2�L�)1Y6كԎ��J-�Xs�Ūb��(��E�	���,��q{`��q^�m���ܗ{]�a��bb��'I�%��$��n�1L��R�-�:�ȴ;#�N2�n���X.�:�2B�	���Ph�$TU�c*�$"�z���Uf�x�@��N R01�Gət��Rd	 ��̒2�c��I��1&	/�|��o�7X��p*�V��
�N��������D$��%�Ү.�\�[A�D5)���b��=KAH�#�d3B��pe�AST�@�b�ʱb��WCr ��C?Sx��Ū7�(؅�J;c$4�VI�q��H��d��b��0��+b�� !��ӒU�������D�R-yGG���m�'��|�'r%�;$h�DA� �R��3,�::�J�SE�=`��Iҟ������'���Zǩ�~*� �ʭi�ʆT�ܕ�R�C�9'�a�il��|�'mL�W>a� E;eV���lϧ���5)R���	ٟ�'qf�[̽~���?	����\81MK�b�>0��c��,�*�ɕ�x��'X�%O%!�Ot�S<�VA�#F
0x^��"ɘ�Lp�6m�<�aA)śf�'�2�'���ɸ>��F�J��TLQW
&�C���WP��oɟ,�	("<����G��LH�����y�r @�'�MK��	t�6�'��'9�s��'�b�X�V�L�h1ic�y'�T�g�F�P,g��O��?��	�Z�|Y�^yI��J��-8��\�4�g�x���O����;����'H�ɟ ��ޙٓ$�{An��t/�l޶,�>Y5�(���?���?qg�Lr\�$ ±n4�}��I7,כV�'�x�2V�>�*O���&���<�S'hJ�eL�D�p"�Cj�l*�R��1�D�������':x�k�o&BUFYRs��̈�a%(Df6����d�O*�O��D�O(�)r_�V�y�e�F}���%��]���O����O���<ae��N�	�n�X��g��\Xr��'�p=��]����U�	ݟ���`����?����1��'Ff�i��� pX��'L2�'|"P��
��� ����O���q��=�z|��E�QD8A�f�֦���G�I����" ON��	G�$��M�.�R�!�	9��B_2K�F�'"Q��J������O�����v��ae=B�����Y�}ΆLhr�X�I��I.[����?i�O���.�:+H&ݳ�(�1Z����4����*�o�������S7�����I���F"vohAb6�)]�� 9`�i3��'�|�����9�(t���U 3�lu�(ٔ	�Z6M:>�f�n�4�I����Ӗ���|�G�)I��1�2EH�|����[�4��M��vB�'���'���U>��ڟlKE��-fT.pJ��{��s0�T��MK���?���󄕪Ñx�Ovr�'��0g��_`�z�݋Q��|���k�V���O��d߹G� }��y��'��O�ł�N�;y�4a�q�鑆���Mc�gr<��x�OX2�|�N�#]Hq���>=FX$Q�	��O�\��z�A�����O��4�n�NYZ�i�)�fZ)�"b� T��M����R��'��'��\���	���ᖕ�n�2E��� U���c:y����	`y��'��T��ɎQh���'w�h�+��N*l�B�eeS70ö�o�˟��	X���?	��*[���D����	! AB1_��sX��i�O$�D�O<��<A�#B���O#D@`����+?0%	@��5w����ѫ{Ӗ���O���?Q�$VF�Q���	I�#2�)�MY9aN�mb�Ƴ>x�Eoޟȗ'7�G�E�����	�?��NR~���o�J��x���4�O��d�O"m)���	
1O��3�:��J�4��L���$�p7M�<ɢH�[�v
�~�����Ґ��K��\�&r�)Uϋ?�$:4,s�P�d�O�I'#�O�e&>���C�ܴ$A*�0dm��+~�� JM�o���oZ�$Ѯ��	ٟ��IПT�SNyʟ(���L�k��B:�VT�����5��O� ��b�"|�����0kϨ,�>t�'K�GXH+üi_��'`�OW�i��O�	�O���,@��:��z�X�ّΐ�4H�l���4�I�TEK������Iӟ�s��=x>�j�#�!�"	��B��M��.0��x�x�O��'C�=xo|�����I�DhЁG	0*����4�?��
Y�?K>���?+OV�۵A�
;�(�r$ċX�Q��m4�%�X�	�`��]yr�'�����z���j��ˊlt�x�B�&����'��'{�'��h�����OF�U0Uˏ:,B��̐`�O����O����<A���?i��?�a� ��&k̖x�*@,��}A@�x��'E�P��)B��ħo�h��(!��e�w��8��ib��'z�韌�	�]�	q�	Zl�g+L�8vi+�2a��F�'��Q�l!'����'�?��k3(�W��q�AF����RQD릁�'1��'��I��'��Ox�\c�|9(g J�N %�Ă�^�8�ݴ��d�N�l����)�O���L~r@Y���}A�Ҙa��QP�`��M��?I�/B��?�Ú��O�s���B���
�FY���R�uJ�	��i8F�ڄ�'�R�'&��OI�)J��9�Ҩ[Ƈ�J.eh e&]��v&��~4M��y��i�O��H�~���Q�T6!?�H�1&�æ�������I�WW�$bH<ͧ�?Q�'y�(���0/[� �e�K�~YQٴ�?.OZ=�K�J��O����<����=<�A�G�U�R\��[�ͥ>a�� ���d�<i���"^>�IC�O����-т&]��m*�ك���q~��'�b�'��1q��*��qGZ][D��?l>8x��*�ē�?�������O�˓A�)Y+����O%R2� ��E<;[�d�<���?����$�uߎ�ϧp��������D� ��{�6ʓ�?�.O4���OX��)��d�+1{�TC#	3=�HjD�Ѳ$���l�џ��Iޟp�IVy��?�"맨?�1>\hI1��\�d��`�${���n�ӟ��'��'NZz\��?��fZtx顭�8�h(0G�ɀxq�����i$�'��I(|o�Tˮ����O����6j�J�"�藻.&ڝ�R`_H'6��'���'���N�y��'��	F�΄3Sad0�A�U�ĳ��𦝔'�(��K~����Of��꟒�קu�`�/j�\����12�ͻƨ�:�M���?����<A^?�	qܧ^�^]�T��<hɸ��.?8H�o�;�� �4�?����?���|C�	Vyr�67��}0B�уWFT�/X�n�@6�m�$�O����O�"n](r�0�D-2;�< آ��,�L6��O����O�Ɇ�II}B]���	W?1��'vܪ�A;R�)�6�Ϧ��INy��D�yʟj���O �S�F�E�I$3P�H�GP6(��6M�O� v�B}bY�D��nyr��5�b[7?�t|���&v��PP��1��d�}��D�O����O���|Γ*'N4�b�\���*U*|�����#TU�	zyr�'��I�������	veDn��0���L�е;�m[ "eJ��ϟT�	��4�Iӟ��'E)Җ�h>�P@�֫bJD��d�Ky�X��h�8ʓ�?Q+O:�D�OX�M�ae�DC-2��x�/{f��V�4&��l��(����l�	uy���=[F��?y�B��<r�	��(�F���&0����'A�ϟ��IƟ@��H;?��EӦG�|�z0�<z�䜈bc{�^�D�O�˓S�m��U?��I埼��-]<���,� aX�枘��5a�O,�$�O���[�n��d�|���TK�6�&�r���&c2 ��1����M�*O�:�̦���ԟ����?ႩO�.�����	�����a]�&�F�'V�*E��y��'&�	Oܧ
uz���)O������K&Il�MM@9ݴ�?q��?!��\���IyRH�\Үh:���z����r�6�̰J���O�˓��O�銉k2J���߂vv�p#݆֮vZ6��O����O
Т�N�B}�U���Il?y�G�]�ʔ3č[�K�0�w˚ʦ�%��{���?	���?Y���e�P�f"�,��,K�C�7���'��em�>�(O����<���[�hR+� Y�E�r��yp�0yD̓��D�OB�İ|�����0"���,�^ij�,�Nf�\+'�T_a���'�B�'��*�~")O
��<j�&�p��C�w��EJ���D��:O,�d�O@�d�O��<���I�XR�i]�S̤����߉#���%V�BY��Z����ay��'�r�'�"�ڟ'��)�u�I�?.j��,Y����!|�*���O��$�O8�S_�1�T?]�	�&��!v-R�k��an[� �ޝs۴�?�+O����O���M��$�O��	�1�TՂ5!V�W�<�*E#�l^6��O��$�<��$����S���I�?�S%�@��x����Q�L���D�O����O����?����E� �PR��^�K��� G��M,Oh�3�l�������	�?�!�O�nԼ!!�3G��y���a�^q�&�'�2�,�y�+�~Γ��O~��睹[=F��E�;��|{�4+�\��B�ir�'���O�n듟��_�b��L-M���
�N��)�ҋ�f�IR8O��$�Or��-����R����>9�8(#��ɓ^1�u��4�?����?9čL����~yb�'6�D��y#� �@%d��".I;@�vS��	�a�2�)����?��p�s�*#�	bg��(r�\�u�iwbCH�A������O��?��U�p{A	�&��ls�@@$#V��'ߠ�ڞ'r�'6��'gP������$����W.rZ��M2u���P�Ob˓�?I)O`���OP�D�+&��d� L&BZ��U�H/{��������	ߟ@�	ҟ�'��嚴fv>��o�/UnbOג�B��bg��˓�?�.O����O �D��W���<9G΀k�䅁k*%��'�!OB�elZٟX�����{yr� }��?!�� @`N@���ͭJc�(���-i��'���d�	����vju���F?���N�8Tjp�άz��I٦��֟ܕ'+
(b�~���?�'?̾�Ksh��A&I1��J>��S�T�����P����x�I���')�� � �2D��xkʯY=��:B�iR�ɬh|��ٴ�?���?���D=�i����%p���̕;~�r\�ox� �$�O,�;q?O���y���/|�zL9f#5J�3@h���&)��6��O��$�OB��X}rW� C�d�*x�أ�H�/lxˤH/�Ms��<�����5�S��W��F���ҽ��8\RR�m�ן������3�JX��$�<���~2K�w�ҭ;��={$Ҙh'L���MN>Y���<�O�"�'9�I�)BD*��V��'܆B�B�q^�V�'��`�>Y/O����<Q�����ޚ/�~P�r�ܶu�R���]}2���y�R���	�H��Ky��m�D�$�ʟ'����P"J!aJ����+��ʟ<$����ʟ�¬݁$Mj,P��5[y����̌�&����Cy��'&�'�ɥ_U��s�O+>�� iS�7dj`8�팀��8CI<������O ��O��8���ORY @��1��Q"�P#O�f����<Y���?����Ğ!�8&>��d���hd��������MK���䓦?A���-���	�4�0�	7+��I0��פ�(gr�6�OH��<y��OIr�O�0l�@�[�}RVL��9ߺ��;��O��䟉\Ej"<�'H�� 1� �8�� �ˑ0}� �oUy2o�\Q�7m}���'���J8?�� ˯���%�V�BA�Bަa�	ן������H$���}5�B�"��<���PNe"�צ��+�M���?�������B)��I�Q�9|pp�����e�b�m-�L]��O�Iz���?9&IТ\ Z�CCI
SE`ؠ0��y���'i"�'���P� 2���O��d��4�U퓉/Q6(��lG�e�2 ���pӦ�O��*7O����	��P��iC"2��2���H�I���Mk�t6R�7�x��'��|Zc��<V�ʚW�!P�HO� dn�ȮO`u�`<O�˓�?���?�.O��JR�N��0�����6��	T���>����䓅?������E��'��!	�N�9$��$	�<A*O@���O:�$�<�&��5��)�67���d�G	30t����[0b|�'�|r�'�O�t��柗uTTa�o��D���� գ����?���?a-O���@��`����ϓk(Π{W�X/a�إCݴ�?�J>A��?Y0���<�M���`��
Tv𤒒�1W�^���t�`�d�O�ʓ% �Up��$�'[�d�G)������ܩf�9�`��C�O����OTV�<AM>A�Oqՠ$��:�i���	)�Rm*�4��݄SNxEmZ���i�O����T~�i�Xvժ˙0J�!���-�M���?�%���?�M>��T���M�0�С�� @�^�R���M���&9�V�'���'��dA'�4��m
'�U�m���+����@��a�f�Ϧ��f(�џD�IRy���O,Ї�Sl�ɋ��%���3�Φ�������+���I<ͧ��5>8W.H4�xڴ,mڟė'Tv	hac)���O��䢟p#�@D����5OQV�Sij�n�D������O<M�O�ҝ|#_(	���� ёr�ؔ�e���(z��e|��0IKP~��'�B�'�	 '�:�)3E�*��t�cJ�,<0<��'���?q����?y��J���D6!�,����H�j�@�̍_��?i���?*O�hH�|jqG,#l0�� �"3py0�*Hz}��'���|��'�B� ����֡/�Y���<{�V,c�j�d���Ο����� ��ɟL�	����I�x*��x�&�#�h� 2o\ݳt��M[����?Q�?_4��	RT�I6<���Mÿu���%�лM~�7m�O����<�CKj��؟x���?q 0��
������Ӳ�/d~�mZW�D� (Q����5�F�(�����J4��M��dѿ�M#���?�5���?����?������?��r���rp ː9M��P'�N	Y{F(nZ��d�'��5!���T�&~ V(1E�Δ&��e�����MKЩ�
C���'Q��'���Ǵ>�*O@����+g:�k�/��*>0\�D�ߦ5���g�D��Ɵ���]���?�B鐓G��B�=$>,9x1+�"_���'I��'��YY���>*OL�䵟���/@�*� � C��)�=�`�c���d�<�G�<�OB�'p�/�X��h�J�A��1��h�,5�6-�O¬�3h�y}�S� �	Vy��5�K۟z��t� �S!��X�'���Hg��<1��?Q��������H9V���~�� �;7抹���RT}r[���Iayb�'�R�'	�a���ͮ��\Ja��@b��@W���y�Y�l����,��fy�ԝt-��Sf�(�Q�+�"�&�/�H�6��<	����Oz��Oՙ�'�(�ۖGC�j��k���6n0bBG�>����?)����$�*Rl-�O~�GC�4�$( ֆ��"�0�9IO �6m�O���?I��?1�mF@��O�P�Sȝ8N�~-��b�q��!��iU��'�I%*a2��2�$�Oz�	L�>:��֞H�ȱ8BA���'�R�'����yB�|r֟�ٻB������$	9gTq��iV��'��"��'�2�'9��O)���5F`ҖsJ�}[��\,F@�����H���?��c��0��HRn�S�fެ	��/):U	�˓"a0 mZ?X�"���4�?����?i�'y���g��N�=+ �A��΋;h~XYa��f�,7�M(Є㟠��r�	�T�� F�f�E�	Bz����+ �@�i�b�'��9:�D�d�'*��&��͊A��i���,I�4��<�a`A�`B�O�"�'�����z�p�� �9W��S`R6M�Or��_]}�V�`�I{y���5v%��/=Ήp�\�c�������M���M3B]ϓ�?���?	��?�-O\�H�P��eH�pL����@�����'r������'s"�'�bc4o�P����/�)aN��Hg����'��'���'�RP� �rң��D�^5R �-���l�RQC�)���M�.O>��<���?��o2(�̓o����r+�-k����T��]0��iX��'&��'�*������$˭b��AzE�/ p�p��
f�l����'�"�'����y_>7MǈA�1�s�#r,��3�.��{v���',R^�yQGĚ����O�����&	H��=zk IrF� &ݺ����q}�'C��'E\Es�'��'�i"F�䍠�-5���ذ�5<�l��WmДM�0aH�j Ik�lD�j�P��l�8��}�����nS;7iz!���(і1�E��?!�K }L�U��⌅|S2�R⌂@�4�'D\� ?�Xiw�$9�x�AeH�mn�Ũ� ��h{bA�����x��z�G��T��2�G/F��Ǥ��OY��rʋ4��d >uq�[�$Օ:�ڬ�`�L%R:N	�F���Sa|)�)�Nj���ő2��`�j�4�q#a�6R#r}+ٸ�����O��$�O�`�;�?���'��i(d�@��0Z�.N1��=�i�vi"<HGH +��4:�O�Y2���%[�(ӧ�ыN�l���.a�䋦�έc�,��g�Ҳ��t��?�*�ψ<��'\A�DFIVX\�K�-�s�'7�H����?�����<iG��!D�P�:d�M?I�<����@�<YPhą:�:E�q&ף}������ zz���'��$^�.�l2�t�j3k�>.��h䆄��@�����Iȟ�C��LП,�	�|��bȤc%��P�N�~���:@�!'\��Zπ0![� ���'�>�Yբƙ���Z�
�"bT$��cG�"��c2J�U�b��d�<uk��'6�A�BC�u$J���Хe��tR!�	A�'V*d!eFRf������ax�0�'Ζ		r.�	��\���A�I46Y�'�ꓪ�d��W;6x�'uRW>A�uĄ2(�u'_+;]��Y�D��Ll��Ɵ4�I�}!eA��@4����Ҩ�?�O�N�"��=l(���L�*<	���Y�J��A#W.5Hx�)P$* ���i�|��`��;��a��m���Q��a��O��?�S����1�*R1p���92+D�X��0��I��X�ʈ1Z�n��d�>�Or,%����GYV^hj 	�^*eEr������'�M����?A)�T�C#�O*�$�O��)��!�B S�r�.iI�D�L�oH�S���d_?T��R��#`�|�l�:������t�S��?�fa�N��K��;h8a��k��k"�C���?1�O����O"T(�ND*v�\t� #T�zz��<ON��'�O8���O��w7�, T��0m�$#���"�HO�����:���[�By�J�� \�E�I埰�3Ǉ7^h�	ޟT�	ߟq_w"�'�x9җ!�mB]3��A�sL}��'>xI�9u
��V��;5��|hWH \��Is9��I6������1\6:�T��fʌ�����$,|O��;gJP��̐��FرL��"O���#��D�(-�s�)8T8KuH�P�������mKϦ�!a�����ȒjD�X�*�S�[؟D��ܟ��3%�����֟L�'{��R�,�8�P���ܑR���iĈF:�����/Y���%O�U�d%/��(�� ˴�� �*4���H7z��q�*��p<qwl��X�	�|b�D�Kܕo�ãI�]lB�W=�t��E@�E�]9�MX�q��C�	;����ϙ*�8%bd�õ~��	���'�\l d�g�B���O��'u��t&�ٝ4�X��/�|��Sf�P��?��?A�E'WfHq�u�Y���S���I�$t��)�sMĵU��L(�eHQ�L(E��$G����k�(i�p�a�(�|"�v�uP�B��x�@P7�K�'�� ��h��:7�؏$�h��m\'S.���"O�����bS��7�5	�[��'1VO��v�L:a��T��4l���3Or��1��%�I����O�x�W�'���'B`H��LK*Ky*<��\��,%� e�,�~6/�|Fx2��)�L�����a��uH��Tsf��h8�)��l��h�l��ա��MɎy4)�&�fp���������LF���ڥ��"܇n �u��+MA(X��?��-w
�9�M�Y�ȩ��Z�nӔXGx"�%����L+c�n�s'��>TL�����Ψ �����O��GOW���d�O��$�O���;�?���*X��Ƃ6����c �*�-�y� ��I�'ȅ�Ag$d�z����Xx��I�g���� �U����I�����b[m��)��O�]���'��{R�ʡu=҉a��#D�$�W8�y�k٬&^VD�$��6]��h$$ݙx@h"=ͧ��@��Aʥ�i�b]�		�%nԨB�/ 5:Î�(�'���'�2"���'^���.���'���yJ�oڭ��'�	!�R�
	�7H\�'H���mƣ'iZT�$�ڞu*���iz���ڟ�bPGN}=������H(e��<D����J l*ƕS7%N�F7�A��.D�<����}��u��7{ԺY�`�k��"�4��R���U�i�2�'���W�����E�'䅻�*)a�0x�ʟP�I���*��A.E�M>�O�J8#fi�'<��	c�(�f>d����-�J��u�;,� �z$�B��3x �A��ZT��� �#@Q��$�O�}��/�-]L��p"�,��@��S�<�w-T.H�rEZt�P%j��ѡ�g~�i>��I<���W��p���Z�B�Q��<�fɀ��F�'��W>��oV��͟P!u'^"�F��p�җ�<1$�{���jP�8������M��?�O�1��L]�vZ`�8��T#y8br�A�rY�T���#W��aL�I6���O2	�$�?BJ�0rd
�l�-Aa)S�M@0���O6�S�џ��'��H��̡w[p��r�׮4a�٠�'HY��'[�9咼���.j\�"�yb�'��"=Qs�iIb�.x���'ߙ&�v�Q���42x��'����s�I'ut��'N��'�t�ޟ��I9y��Ӓ�Z�k�i�#)*3�v��D�p���O	9H�qG��,of��N]	��d��K��}RJ�H53�)Y�,��;� -t2�3���'�����OJ�3^����Ս����Ő�
K�ɇ�S�����]/8����ǖv�q˒�m�4_�0e"��M��o:�y	��0�L���C1�?9���?��������?��OJ<����P�<g�!fh�'g�l�RH��i[����NP�:�;��9,O8�b m��
��,3*U�k� �8aH���=�؈��[X�l␪�O�d�(|�1�a6q�����'�!��ӧ[�� �D�?&
 ��"�B�C�!�	iz%[!�H�t�| !��1E��D�M�	E�!r�iOR�'>�Sb���� �­`!��>1j�U!�.���ҟ�+Q`T̟��<�OV��൫��w&� �\�w��aȍ��՝j2�?5j�EX�v�H�Q)�0{��zí"�4�*$��]�O��!���+<G���&�\h�r�p�'���NۛvNx ��p�(Q�;ى'�x�(�O�(�����c���R�'�b�)��r�D�d�OhʧV��\��?)��Yv !� �Ht0��#DP�%��-��
	
�l�'ש	'�5!op��Sd��L��(~@NԠd 
-���F��4�����y&P1Y2�$]j�~�I/zPHTь
�N����/�;R6��_Ƣ��>�)�� ���	��4���:$�´8(<D�*P��+����v��ZɦlYtM=�Rt���4�@|�# � ��	BOs	��:��?�W�3�z09���?����?9R����4��#��#�t��+P���a�OJ����'����'��N�c��� A���'��Xd��!H8 r��W*�}h���E��Iz��(��e��!'Nҟz�P�� h&D� A3K�QLܙb#�δ�rh��`٭�HO>5�o���MK��@(I�e�t$zӶ���Fι\h��'���'I�A�5�'��:�8(���'b¤L�XͲ�k��[8d#��ek���p>!��tyR�԰C��YIBi�M���Y�'���p>A�gޟ,�I.^��DhT�ۍ��h	t�M w��B�	����
(`�D����(7rB�	�A�����U�Ą��Gʆ-rj�	���'!x]2�'��'[�?.]�����Z%3�ڔ��f
�2�:��G�J��`�Iџ�8�� �M�O>�)���!e�F�W=�����X
]����V�_�\ �J0a\^<�%4��Q,<L~�R�����L(�/�Q�4SQ��ON�nڰ�MK����?r՜<���I�m�����M��"��*�)��<����#��0�#��?�hL���FL��hO
	o��M��~F�(��ڮ2��QY�+Y�zZ���jF�,�S��?����\�T����O8�䊻[�`��f�Z����Kh}��b�cE?woēO��g�'t��#g�H
̌�SES�O� C���x�U��<���G'�����,�{��<�`���Y
xc�._����G�'�"(`���d9��� �8"F�!Y3��p��Ë#���;�6O>��=�O�8@CZJ�����Rj��з��OLDl��M�����<y.|�Qe�+90�����~jP���ORy0�G���e�'���'��	l�)�I��ȹ!D,*����d N/H��\т窟d���3�OV�rb Q;�څ���'@j<�)��Op\Є�'p5� :k�%��'r�'���F�')b��,Ob�Ġ<�(�,Z�8�s�J,+Z�aJT�<qg`ƬUy&�%F�)8������������O4�I�j�Ҵ;شτ����K2}R�Y���
W0 ���?A���?�,��?������y��)���i�©��!��E�]�c�;BŢ������Z-�M#Qm��9�<4X�Α�j�^(�h�b8��r`�O��ĆK_�h���-��#@�ê����O��?a�ʟ��Wf v-䔚ƈ+��!�ć�nc��Z�Ȟ���H(��L����S}�_�`{����M���?	)�l��\/�h�	�g�q2�,M���O ���3G�����/RJ�z�I.��OG�ab@�J2���t��,���)��D�H*\�ca�÷Z]Hur�C�~8(wV<1���(�K�-pu�mZ�N��p�n��f�IҠ�$�O�QoZ�� �O�F�LY8������0m�p"��'���0Do��(�����9O*��}̊-�6,H�'�e���'D��v|�j�NI	����m��-�`x��c��.ꛖh�='�7M�O
���O"�I�%Ƭ�$�Oz�M��j� 4��`af�+;�����M����'����Ob�ar�؆>�ܙDi[�V � �/6D��R��|�P�����B��YXɦ�'B�� ���L�F�~h��'"�7MԦ1�	w��?	D�F���3���3A.h*��Z�<�����-�S�t���0�)�0���9NĨ��k���O�l�3�MSO>)���?ucT�A�W����A�]\���.������!-&��ˢ�ܟ��Iɟ\�I"�u��'���;(��&x��Eӕ#JP�i���"�z����*3{��0���E����u^���խȜ{�� �D̅UxPJC�d�FT���ǈs!��ӟ�"=��J�h�t4�3�ڢ
��@ժ̋�?�vlG#�?���i��'���')��ywO�!;kb��M�rZ���,���yr%γ
�P�@�oH�R�.� ��Q��#=��V���'��[n��t���J�p�4xtC�3�򜡣��O���Od�$��F
��$�O��)�Ly{V��OJh���M�0U �p���BX�G�'&��1bc�&�?��m�,1"������o|
h�`��u8��!���O��ă�L�x��'\�=�K�(h����O���?9�ʟ����Kkli j51�b���"O�X�X:Om����/.�P�;O<�~BQ����	D��u��'�rU>1.|̌;��K.C�>� �8[�Pq������I���AC��d&��Os�=�RN0E=�H���d�򄈍S$��)UP^�i�X�4��<#�"9���&w�t,XS �y��<��G�������MS���)��Te��h��H�y#��J�l	`���,�i>=E{B�R��"��V!=��#�V��0>��i�d7��OJ�)6N�Y7>��F�X%9�\h0�:OX	���8gt��d�Or�'{n�I���?)�������R6"K\|��)QN*�1-���`mR��Ņoq<c���(��OF]s0���A�JA�RŒ�'7�鸓`!3�>8�H�)/����Sן"~�	�b#�P� ,��`�"g� 2�`9&�^ן��	���	W��?��Ղ'��4�%l�h[���<!���>u�՜c ^�`��Z;+ƺmP�F�_�'&#=�OΞx��^�~IK�(Ҟq�@�'�b ش;2��B��'I��'�h�A�	џd��V,a���k����>\a ����D:vcS�dv�(ಎ/<O$�yeb'�t��֨Ј���7��Ɵ<0�
	���Q���D��I�M����h�>O~��ţM����Ɍ~��Y�����?˓�?�,O�a�A��d��R��M����"O��ҁ�S�cz������?(�2Wl�S�����<�� @�p��fO�O4}{̖/$>��Q�@n�b�'���'e�%��'k�=�8ErB�s�����S�<H�a�ތ`Lf!c�>(��|��A�w��	1B���WH����|���H�}l��$#d��'�NXIV�h�PM끤G0h���|��'���?�$#ɲ ���A)�G�e���5D�Љ��	()p*�
��LӴ��0Kn�|i�O��R�tI�ºi���'��6"PXA��K�0醌e��9���#v��Ɵ���🸠Q-�'b������"�n�ZეK��+�;V�K�sd���L�2�B�EyB�m1B�	��Gt�!�c�Hk��%˺iaT�`@ɒ� 3�0yŋ	�(Ov�P��'E�>U�@��*�� Eÿz��+&�'D�� ������.��)ŮF�yx�!��'��O$Т,U�t��	`�Y�xl�eS5O��"%�ܦ����O���3G�'�"�'74̒��P�@�:��� ԼbB��
r�7O���T>#<����� 4�I��E�kl��Ě�.��+����OhH�f�i"������|Q�����F�m���?�)�矬h�'SC����e2���#D�D�둕\�z���iM�� �@"�c,����^4rC�'/p�(�F�9K�L���?)R�L������?���? S?�,0��Ő�hɺ|��
>08ʷ뻟0G"S#j4L�`��'U�bPk�7!��P�C@Z#��H�'8l�H����9��х�ɼW `)�E�]�|��1l,)i<��	�?[�	Ɵ ��?��?�.Oب�C&��.ق� �li���"O���aA�x-VU��Z�"Z:����S�'R�Svy֭}Cb7�$��)!���
� ���ӣj�f���O���OP�i!��O��v>Ţ��O|��B6Y�$��&�Bul�q�	G�g�|�l���d,x��ۣ�IV(�K�.V�|��S��?��xFz!�&�]#.<�Ԇ_' ņ��M>9���?�ʟ4�����s�4��B�\-&�T2u"Oz�R��V�|a>����(Q�&�i�7O�8�'��	�M��0y�4�?����鞐�؅�Ԭ�k���k��Z�Lc�	3���O���O����`�O�c�ʧ�*���G-t��S)S�otEy�"L���ȅ��#��*�ԜP��4)�,3B�	3!T��-ڧbJ5��K�!_�D�+�C�r�>�ȓ
d� d��#7��3��ӆBvt��I&�����0�b��&P*�#�3V}�2��Xp�i�2�'��O�(��Iϟ(�� >l���"��S��*`�˱UwH�1�C�G2 :2Gձ4��<rf��>	��=���p �GL�9����q�QR?�����#I�\��E
�u@�FH���Ҍ��w�`�q�Z�
�|Q��*B�$2��'�b���O���GM�`��#'�tr��%"O��3�eW11Gzz2�C�K�t�2�I��HO��:5�S�ǶU�NxZt�8b��I���#d+RN���Iß�����`R\w��w�H,ʡoI�.��@��Bw�OȑQ�* l@�(T�����$��a0h��G�� � ���$:h��(N�xc�	�k]��X�֟ўl��X�8)#VOqe~��������ĉ�OH�o���M#�bl�~�ĩ
M�l�qrm�ժ��*ԅ�u0,���/,Br��-֢����:���<�F��v1�V$K�ZR$�?�X��`疾<H"�':��'6|	�C�'?�5��\I�E���M2f
�,`0xJ�M�-$i���Ơ�_gnԸA!>Ȱ<�aˏҎ`�r�K�_;�:��6�ZU���S(�\��V��PHay2�'�?I�S�t��Y aWέ�aB%�<-Z����'^�>��(BĄK�(��n� ��V�C�I�9�F�F��/]��X;����������1�S�'C�()zGg
�&4~�F��&mBf4���&�;3��J���s�ޢ�F�ȓD�(hR�M��h\C�.Ej��%�ȓBR����v:�q�U�?fp恄ȓ�jAb3��/zH�Y���_tL��|��Ђ�@(|��Qi��X�qp8L�ȓ��ݳ@��<dͰe��*��jلȓH�D��M�)�:��"�A$�̄�f�|K5�V
\��b���I�℄ȓ'g Xp�b3H� L�̢9�`	��h������"��pp��B�3�n��ȓ9L���=�X�OյnX���ȓ7>LD�@*�5&�
�cT�ɲ;���ȓ"[r�Ad�W,{�t�#E�0����W(�q!,��a����c�/Fk~��ȓVK ���H��I'�;?�d�ȓ'u&i����a����\����'� �*q��0Z`@A5L��E�24��'��\����*8��,Rd�)8�@��'� I�W�� ��E�iڸ��'xƑ�A�"�lu@T� &vo�@��'l܉��$_�M�h�B��P(aj*R��� d��'��[or�����H�n@#"O��%T�eL~��U�@�j��B"OD�y���
n��0�p*����3"Oxp!��T!�2y(C*�|j�h�"Oh��Qo�*N܁2jE.�v��"O�,D���@�(d+5�٥>��x@�"O�)+P
=8���AD�B�B��B% с�/@������) 5�DlL$��.�s|����Æ�-���i&��&=a�OPg���i��)*�@�̓$CV<�A��<�.OV=�E�Q �Y��j� d}�=J6�>!��J�g�>9��C�L�}r��v���5�B���@O"|pra��a�X�O|i��R��jң'y�"��e�1�.1�%�ʌf=�p�S"�/�p<a� �8R�p�O�}�6�O�&���!1�'{q���e]qQ��ϓ
sT(h���;D����*DrM�4O5���aFTF���&�U�+e�pv���M�ʉ36�����M"��)�u�\ YN���1L���1��W$a|h*���`岐�a�'��9�L6R��8Cgf�;!�p��F�]ǐ��S�N���O��z�D�'�Ph�N��P�8t{�D��'@H�ku
�<��C�Y������a:�BЌVn�?5���/!$f���R$_D�dn�"<bܰ���? ��dE�%7al��2��$�~���	֤]p�V+m#HQIַ�џ�pf��*�\̀�JԹ\����,�&�����,x*D���H^;�M�e"�&S]�؁G��71�i>��F�Ean<���	à�RD�C�.d  ����0��PS�T���-�p�H)i
��7q�Zd˅�ϰH��©O�O������졉�
�"9�L�p����	��B��0�O^��q ]h�B'*�����W잹zLH����k}r���&��!Ƣ�AL��LO"��i��]?"�����D�h aj�k����u�%��F|�@-�L,Yf%��8�ՠ�h�E��� Ĥ��%��x�a,E% n��w���
�D��^FRU�ƚ<w~�D��q�'�TEZ�+՜Y	eJIJ?���'?�0�Tŉ�&�E����oDdu+݌yK�B�>�"-���F���%[��OƦN�pL�Ӫ˝.�<���K�B�ۄ�d�7`��"4�%�3�[�X��,� �^��Xkƃ]p}bf����$�f�<�.|Z� D�&�P�
�6]it��d��t� �pI��_�,�i��~���� O$��'��K��N�tYРIΏ.�m��E@�j��K�	�e?٣�[�i0$�Mĺ
�=���g�'ڸ���S2PD��#��5`Y�#�Z�eN�%hsg����1@��. /�,bLZ�r�����I8C��� ��ڢaF��VB8wa�u�&O�z��P䤉-����t�Ւg� c�l�	�+��4ЪQH'Jͦ�R����#� ��Bĉ/�X��!n_��f���?��LԂG�\���$5
,�����=MD,: ��7Xq��?@���B�p�y�I� &��n���8kw�����Ο�x	Xi	�͕��0?�b�X�?����\�9%x�[�SA"��:s�i�r��	y�Q�H�So~a�K� ��O�*j'����C���Rǎ�P.�$��//�F~r`��~��0�.�<�x��!��#G��za��~��Y֣I�93���D�=��2pH����P?C|�4H��W�p�f�'P��E��PC�uצr���Od�X��
�r����� 5L(���&FF�aC��iW
�*���-4��Da{M�����g�ށ��I���ѳ�LI �~�{
Ǔm�Hz#N�&���h�77�L��r���G���C�bB�O�FX3��E���O����Z!'1��S� �6��]ZR�ϋ��>Y��ީ�V!JW�
d2ĝ�p���P*i�c�p��������U��)� a�P�p�ϘV��Mq�P�z�z���+?�{�J4�AշI�\�1���.]��H�kQ1�AO�p<6P��ҳ�ē�y���'�w%��c0����&��	E?�iCSn�����2��$���0L}�ew� �4dJ��Ѐ�̎C�\\ہm&���U�~)a�
�f�l$8�MW�M����e,\`��D��D����s�R(�bC�*����Z6M�^�ϓM�4���
.M�d�P�u�(�fK>Pi*�=f��R���Hi��7B�1<h	�҈� on���'���A�I�l� D���J�e����%�4��H{.�+O|�i.O.�W.I��y'�C(^1V ��hJd����Z��0?I!�5a����%�
�����/��<�FA�D׈��$�r>��Ei��?!�mE�g��I<;��$ف��^����,��#>�aK�D����Ƨ
�?����8���;e�S�.6ur�CH����cs쟘SV8���iC��Uy��vG��;��$F>r��(a��7�U���֌ �b� 1��"&Q��*w/Ch)h�
�%V2�)c��R��T�L��s�f�0����Y��y;C p��!���a>ttXN�2j���i *E��KW�U��+�"�H���P�$��=@(��ww��#�%J�Y����4/�#�`x���<2q	ک[d���E�{xJ�r� (Q\X�ǋ߸{���<�ÃϘ;��ɲ���o��͕e~��Q�wY�u�0k�cD2\0�% ��O2�U���\'2E�Bm�A�e�d [ ��4��;] ����?]x65��ő�?�� X�J��ГoB!*BL=��I >��\�$�һT���p���~�R�UG�'*���H�g�!k�(�� U ~5��0'�p�SP��zh��$%y%(EAw%K�y�9"�U�}ǒp��S�? j����Ƅ4l��E.�|�IԬ�,/l�LIA��<l��-�Ǝ� z�F�ϖ,����'`��J�0�r�q
��d"J0�
�hL`���'  E �7���;�F.� �X��5zv`�Ӆ��'!#�0� ��Qy�}��G8�}P�J!N: �Z��:�`���O�HcgH@! #��M��6�i��ɶ[m$�X���lX 2�܅��`ӽL�I-����1o�U�Jx"��6c�LQu���_sV�X��2X�`1�H�4ax��n9��xD�]�n�PTJ�� O��㐯�'�X���]�d��L� �(.���z@�M�./PU�O��e��F���y2JႻ�Փ]M(<�CX<z��\�!L�p�"�{t �z�Ģ5.��8�4� E+�gGqO~��Ɠc(�.�s�v�(GK��b�Z1�����DN0��PCUoO�{&6�G 8P�>�;V╜Z��@j$�S�X4�Ii?��@��1hb˧6GJ��W�	}��#��ذqd��|�x�*�$o(qOv�X�x@焝�.���;�MC�1���'/��2�a��-{��p����Q�ι[�C�?$<��۶�/��Q⌛5�t�AǓJU����3@Q��j�*ЩxF��R��\�N1 	�6/��c$��?��� Ѡ��c	\U��oD> �8��e
ZK� �"AS�m���@O�}��'r�$q䁊"z���ܴza�B�N�DN�QR@�i�$���',�H�K��O�(�OT��UJ�P��ꆏ٤3���	���ܼ �TO�0�p�ϩYA��cI���8�B͏ܲ�W` �+鮱���Z������5OḖ�*�)[0��4�|0��EUJ���ʁ��vC@�AW��T�O@�ק�����<+X^�y�ǀA/P����_�;K̱�텸Wzp�
��},���Ǔ`+x��cnʴ^�~T�tQT�̓yf�M���7���I�Ta��@Q�+���{2��!���PW�]�N�:̀ dH�g��zҤ�N� ��&��U'÷X�*�c�L���'����S��(XS�d�'OؠGL�笠O�9�% �(	���PQ�Bj��lr����N�,p�����x��+��Ɓ�0�K�ρ
B蘊�Ȉ�B�lΓd���$�������!�0��.� e��lQ�Q+ÈI���k�"}""=��8HW��/��!�aH� sb�8�F��4Ej}�&�P���
4/&�\����\e����,ۭ[-��5s��!�ٴ?U�d�q�5���Q��`=������ƛ&+J?�p���9i�؍����{2ўȊ��\���cF�6��l�ߟ�[�(��LU*�"�f	�4^�@�`o҈ٜc3Cȅ1y�,��O��� ��_��	��I���1*�=O���ǐ�@
��*�'�Y����?�֝0X4R�3s�K�<L*%/H>&��A+Es7����r��AdJ8�ɉ���W6LC�е/v$������L �HBtm�T |��G[��k��I`#���c �l^2�ű�u��J�ՆԊEo���jC�Z)t��UeXM�'��@ӛwY�8�EV�w�e�U�FSK���K>�Q�V6Sþ���M1}���(.�9O����J��3�Xԉ��ʳpo諱�3XVV�qN�z�]{�"=����eT�%l��P �>~׾� ��e�FdXv�ֽ��	;$Ô���'����s困H2� �'p�<)� �"���QF�Ȁ~�iC�'�r�#F��=%�����=kr(�=��'E0Q�4��"~���4)ߺ#Nz��UMk8�'ǜ�XE�N�qZ�炘@&�YK<���F�`��yxt��+b0IE����lE���C�j��?���S�'�$��jI(B�����&�ԌӀfQ,�� ��!�i�5@�X��ҜwK��!5I�|�-�D�N��LYO<Y��i�8t�?�LE�$��/f"4��0�Z	?��Icb4-���`"J#��~23iD�R�~���<(ZTѳADSbX�-����e�,�����8l�}�G�4�"�-ҰrKJr�/��a7ظ�x�� w{��r��<80��$����,��?�Z(�6��Ղ1"%��nў�K�䟕VʸL;�&V�`ÌIe췟�xDgB�?*��$L�DȺ���&���*ޫl|x��E��):C$��#&9 ܊�0,H�?1@��-q��ƥ��AC�3�!Z�S�dHŨiZT�����1y�l����Q� (�'8l����'$	DM�hx$u"G;H�⭡Dj�� TQ�=�O���J4�T�6��Y�O��7 F�82��`O���໔i�0�`�G)	Lv��y��O�*I�s!��HI�۽%�(P;�	�iy���T;O��YV��c�����K?5�I���'	B��%�#����Q��y�C���K�mM����ɗO�.��t��7�s��z�àrFD�Kq��=+�5�b�H��:�əT㞔1&ҟ�A�ӄ���y��Q�'��� �̝~�0�QƖ{�zR
�@b����:51`m[�Ϙ����-�H��OؖE��;�0@��<�� �O��I��Gȶd�%?�"5 )d��x����Q=�� 1( "i�qO哑DH���v%�).#z]ϓr�
�3�d�3��P㔤��<0�)'��W�87�������2:
�1�S�L��
�b�
��I{T��
��<�����bt匔��	�t�ٳ_z���j"�M`��It��4G6pE��$�&B�$�Ә'/�h1�G4~�rh �Dr��1s��7m�|��2F׆P{��qv�3)b#�":�tl
��<�p<��ѩL����w�~�[��c�p*a��	"�r�r�G���3��Rvژ"F w>c�ʧ_�u��P���3�&\t#����d	�e��q��<��1���j�"D~�� 'N d�+�T-)@�Ji�S�4H^�@�4�( HG_(��
wb$��_
	�x�qQ@�-r��2)WOZ�����9W������d�Q�3� 4�-��5����A�4gT��b�O4�S��̸O���8��6#���>�M��#�ED�ˇ�9��Pa�؂�L��8H�����A��! �MTɋO|ΓA���&j��H>�sFh58����	�8���*���'f2Y����m���S�>�n	H�G0
���6�S@���冠$Pz��H�	(,�;�I����IV�e��G�.���㼐[îDxy��=~e���j�RaX���>�?��.��"ֱ��H��Z��T��Px3��I	a�x��@���OJ�>i$�sy��򃧟�JVmܤ\�"�[ g8! �Z��R��'T�!D�*c&�)�"xK�+�AՀ��Nȭ7�KUA�+N�D�R� _?`�1OD�P�(O ��H���G�2c�|�2,E[)�� �hޛ]'Lth��صjCR���
�*r	��q�D�6k�\����'d����m�l��5a�r|���ANY�\vp�O����?e�ֆ��=����p�A#��}��!܏x!��зB�O��3�$�'H����JJ�|F|��l�9�W$�	O����� R�m.A�"&�9ł�F~"ŕ�Gjm�;���E��.lA�0�ޮ�ƥA��Qأ>�l���x�d��̣�%wp�x�0�TBx�rbc%LO�D��
��ɲu�<�(@b!{�(�Q��4����Ri:=떬E��*�` �@d��|���sK����'�䀻����T���{ �����G,�H �
�yB���J�J	�X�i| \����y��"Z��=Q�d1��H���7�yrcG7:�Ji���.W-���EhI��y��׭D�)��TF�	0I��y���6܀Lw�P<t��@B�f��y"�@#�HQ��_~բfn�8�y�NO�������U,����@�yC�J�z�CC>{��P&�Ź�y")P�.b�4����>`}"E.պ�y�n�&[���
sFO�9�����ԭ�yBS�-��e��HO1d-A�!Ӗ�yҦ�`9��@I�2�D�1J��y-� �A���[7b@ȑ#��y��1jv���PSN�:!*�,�y���E�~4�-��F|(����-�y�N�%
�C
6�`Q��y2�X6-�b����.@�:�9w-%�y���$L�4���,W�?�,�'E1�y�ܟ3�|���`�8�P}��	<�y�aM�@�f� �ݟ"�-Kl��y�X%��A�掟�,t��	0%0�yrǕ?{ي�0j�;��%�-�"�y�JL�T��D8�@H.��Hz��y��:x� h�
	�=3���¢�yBE��uO���c�;k���ѐ�N*�y2ƩI�aK"Ǘi��H���b!�'��Ux�I�:@w���&��S~�ɂ	�'���9S&2�2d#%�ME�h�8�'h� �eB�0^���BX�8�� ��'�2ȣq/�$�6M9Tj ����'����@��{�n�K������kL�<��=�$-*E.؉�l�T�I�<���ۗ\��Z��'��h`mO�<q�-9w%Rxk�Iʇ�nl��Jb�<����f�.ѪNH�*l����G�_�<�0�c#,�ha8M��)��@��yB�4vƅ�&��@@fiQǙ�y(N9AP���Q�H53�
��!g���ybD��1�T%�΁%)Y��*���'�y�C�'�@0[�n��7Tm��L�)�yRFZ�y�XA��_F�\a%���y����$�,�jb��7DP���F��yBf��.�tQfg�C�R�ˈ��y�j³e̼��ڢ�$��M��y2�]*��Y1A�0�~�r����y�C�0Oh�ؓ��)(.��3����y"��px z[��ͣ���
�y
� ��'C�ss��c�.=e�  �"O��B�XC�m"��D,��1�1"Oq���'`N`�B]��� ��"OH�Ke�9���/�(o���W"O��ʥ@ِ�U`��u�H���"O9Y�%وf���;�EL���7"O��C�.J�g�,9p�jڃ��Tȥ"O� �wF4q��9��<{��|[�"Oh�y*JA�&���i�R��ik�"O������)'��$��4�XzFn�g�<�cV�2��BE�G�u^�,gDx�<�N��}��mQB O#::	�@Py�<�q�ǝ3��yjŤ�A7���'d�z�<��ʂ'�XI+���`��i��Ŏu�<��`�/o�P
� �t3iAu)Cy�<q����D!Bq��jD�s��u�<A��ۤ�ıʧ�W/iz��hi�<��F�Be2�Ѽcm0	R��D|�<��H��JA����Q�4)��ȇ]x�����<�s���XHB�z�fF.u�j�	��_�<A�@L��6���&VlHeYBQp�<iCꛊ8:d�! �y)9׭��hC�ɛW��1�!,�(9��B���=��B��
w��闂�v��af��nB�I�w� p���<��@�!�6�Bb�Ї�ɉ�)*�#[�RK��Ŧ�\VB�I3h��ӕN���Nx�#�(B�	F:�=r6-�-F�R|���+K04C�	���c��Px�@q��B�ɶcDN��"kN�<D$
S�@6�C�ɨ7
�m��C�p����2l�DB�I�~���Ie@��
3�z�[��'��O��:Uc��-O0HP.I=yn���"O�d0��'1'��o�v}�Lx�5O6�=E�t�� -4X��O[���K# ��yRАiB�qP�#w��)C���y�
�cL���Np����,� �����(O>)C�`�M�(�*�H�!C�>�{C6D���R�C�4��y���S�Y��'0�4�O*U���	Qk��:b(�
��=rcO�Uy����%*�D�90����FD(_!���%}@X�ʸ)*05`�QO�x�$*ʓfv\�cFs��RV�"�:`�ȓV�}YV�3��eZf��>���ȓ-*���1W̝y3�G�e�BM�ȓz�bժr�N-!X.�  ��5gfz��ȓKʆ���l]�(�p����Q�*І�Il���.�.o8f%xS�կ8bL���	n�/6$(:�$ ?|�P�"�Ҩyld��ȓ'��Qc���=n������(n�I�ȓ0��I���R<S���Gi �U�l�ȓR���#��^M)�R$,��u1����)ǖD�4cɜ[���)�@w�G���G2����
X�*T��PU�U�{��C�2i)��J��9fp`�R�I,kB�	,�L���^=G{����o�r[B��N�)"ƈ42�
��7*ڨ�<C�IT��"Ç�d��8�卣H�Ƣ?���	�7.+N  �DY�yj����苨\[!�D�� ���J����H���Ņ�	C~�F�g4������9x�@�� ��yR�	n��P"VeU�-Ŋ��s�R��yb�C�4��Qĭ[�$�ڵ�R���yro^������d ��(��-���y
� �P�q��g���méE���"O&�X�i��C�X�uğE5:(��3O�i���'ڂ=���E& �4鉑`�5D�Hߓ!�\� DK�y���X��$S�h � �����	�yR%[�NXjd<�A��-W�HO����S$,34X"�h�s}TQ��� �5��C��%@�Ț�C�J�Jȴf�1E@C�ɾ]�t&��~`
h�D���Q��B�ɤN�Z���K�F,�z˜���C䉕>��(4GDl�	���N�|��C䉡W~0��S�Gĩ�S�B27�C�ɰ��@�W�	'�4	AV�Q�zC��6cB�8�.����)c���nC�	�O�@y��f��qC'kA�~[�B�ɥd�ޭ����_������{��B�ɩ`S�DAw�@1�PM��_��2B�Ɋ{�X9�`<xR�"Afтp
B��$a�J��-z��	cM�6]�C�	;ȩq��
N�ԝ(���$Z'�C�ɿa������ �p�����ڇ-�C䉶I��X����m��yz�� Te���hOQ>չ��JD�&��th3����-D�4g	�'�L�KWE�_����g	'D�X�B-Vm%�P�N�f*�QA��#D������	G���1��B�8�[CB#D�8[��WJH.��Qʒ=sx�?D�0�V#/^��3$#MȐ��"D��	T�Q���t�ƧH$$��0n!D���GCS�P�� ��3/�k�	>D�hu"�#e��9���m�yA�L:D��ó��W�[ea۝Di6-��6lO��Ђvi��Nv�Sz�a��0D�$����%� ��E�����y�&/ʓ��<�׍R�~�¨�#h�$1t�arbc�<Ir�['����#}��`�₅\�<	���.�m�" =n��S�_�<2fR�}�h	ʴmT�2�Z��`��B�<���M9�\ʶ�/�8|(#c�~�ܩd�Sy�0��*����[�L2D�)5)�s�\-p�]zB�AT$5D�d�'�i���e��e�N��!�2�OBO��X�̽[����o�*; �5p�"O2��s�0%F0Ta/@�z��x�q"Ob�* ���0��Dy��0B"OJ���kM�Q�x��AL!ep��6"O��3�� K_Hi���,�̹s!�gH<�����m)�b��M���+g�F���>iSF� i�}�%�3/L��r�{�<�cԙ8��t�a\�>���UJ�B�<Q%���:䪴4�7x4DU�	@؞p�=�6.C�#4�DS+_/��M�"��G�<Q�H�*�>��Vd�{��訃@�z�<aa�yR2�{��,+�v��PEHv�<ǈ�_��cAo��:��8�e�i�<����=o`���@�^��l�%� A�<�eI#C�p�Ju얚n�Ap�v�<鶍�#{��y���K���A�+k�<af�Մl� y[���`����F�h�<Y0��!�򕠤�T}��H�D&Rf�<��Ρ9�A���#�P�r�c�<ّ��/� K��4��%
gȏg�<�B� ��-j��pߜD��/�l�<!�o?l8r!p�T�W�|E���A�<�bm��1����Fn��	,m���e�<� z�J�P�HO��c�F߲x,����"O�Y�a��#K������*���+s"OB��U���#$=yC�Ƚ{�� �"O*�YB�[UfP@�`�3&zΝq"OxK�Ø�y��݀�/�Xh�`�@"OP(�ݤ� �����RID4"O���I�j�������o-)�3"Ohm�ש|���`#"@�+*6=c"O`�[C�>)MN���KE�y��Z�
O7�R6	�g�Be�Թ! ���%x!��]�6qiԢ��/�a���V��Py¯Ա\ ��A�<2o��	��y2��8[�\"5[0#���;�D��y��$\rJ	n�$Q�&�x3� 7�!�òu/�X��j��is�1s���!�������1T�\"��c��C�I�%²�
s��79� [�bZ�g�RB���
S)�
R�i��@�cOtC�	�~y�1� >e��qǕ�k%<C�)X�(���VE�LA� ��JPC䉪<����a�J�KC�8�B�ɷKm���Cإ��ptA��J��B�+@H���yܵ;�eͯNӚB�I�pZ19 (v���(4��B��4YY�}��b�9G��$����G�xB�Q|�iؒC2"5�M9����C䉅x,�x����(~�H�4H�0h<6C�ɗv�h����
^4၇����C��cw��b��̱�(��C"D�*C�	�4y��5Gqp�B�nHB䉏fsLD"�ğ��>��kލ:q~C��#+�Ĉc5��7@ `���f�@C�.�HA���
�+a�<�(�UNC�I~svIҖ�����	8u�B�	ẗ́� tgφF�*Ec��)7/0C��:�
,���8��3�H���C�I�6g�Y�B@�j�����ŌY��C�	�2g!��-U�L�#@C<F�hC�	�9\tQ�7/ɈT)KF(\�`bC�	��x ��ς/9կN'�B�I)ГA�T�4���P!�+�C�I�7 ����♘` ��1f
@պB�	��Ԛ5 
i$�C#ċ�oY�C�IV�\���;o�Ȉi�	��B�I�M)�5�Q%���!�ʟ	>��B��	z�(8Ð���7`�,C_�utC䉕_RDUt��'9��(jƥA�u��C�	(o�UA�N�? H `� 9I$�B�I
I/��ʡ+)J�n%p�MC�a�lB�ɔ=�`��&���OTlaP�[�C�>X�廃�9z��ɑ� T�X�PC�	?{�2�fz%��Z2�3qKrC�I�{�K�+]�@z���
��N��B�	�M��hp�1j72��g$Q�TV~B�	�aqF�`P!F�H�2weԣ+VC�	".��M��E�1!��y�E��\$C�Ɇ}�Q�΃�h�6��0��2�,B�;=�X�RK� GX���t@�'?B�	?W����Cη+�APA�@��B�	�V�µj�g��.���aSFHB�L�L��@��c!��Ʌ�P�GY
B��r������L��A��|�C�I�`��5�EȆ� ��e�d�O�O2B��;��*�͌�ʙ�fg�		i�C�)� �@YTM	�N��I#A��@Ȭ�"O�Ӑ��x�p{GhP�i* ��"OH}���J��$H���~8[�"OZ�[����HqHȗݲ(�"O
�B�&�/*��ʐ&ʼ���hR"Op�(�I�:jc%H/�8q�u"O���F���i vɓ/�c���"ODp3�
X<9��C"��W�d"&"Oԕ��:_�ԃ��E� #�"Od�E^>;�fѺ�ȞN�ڌ �"O�dr%�> �$l3��
�.̩t"O85���≉E�',���:6"O����Ͽ����}��E��"O�#��ߴ\�Ss��X�$!�"O�Ɉ�P�\�j��"$!ݒ%��"O�uI�ӧ
5�d�/HWϜ�@"O�y�I�6/.���DO���Tؒ�"O��C%M66�̻\:�=I�"Od]����	1�a�wFF�|���"O�}!BŢ5�ԕكC·j���%"O^x1A��~T�,	�����"�yrGͣ����H+]N�H��֑�y��A�eR>�{BC��MB�����y���2������@P�`@��3�yblT0wz�UO��'u����	��yB��Ao�剠癹!��QR��
$�y"/2=�j�M�RD���U��y���)�T�jpO�	�Ψ�����yR��?X��[5+ߤu�l-�dө�yҡI�E|���f�I�������y���E4Lړ�~���+�y����y���N�t�~$1򬉟�y�'�ZlY`@d](W�<@:L���yb�:zܼ$!�
�'J���P)�.�y��T�y^f�HV&R(C[FA!�@Ō�y��ݽ?Zz6&ҮB�4�K1b_�Pyܷ:Pv��v��I���`����y�������S��/�����
Z+�y���s���t�ޫ8GAґ���yR�Q� k��`t��$C	��A�п�yR�&"�L}���I�QX�0 N>�y���Tƈ�ׅ�P�F�`s�γ�y�[��u!�/��qԄ��`Օ�yr#W9}x00`a˷;�(ى���y�6k~�:�'�0�zI
����y���:�~ܠ�-5�l��D)ȝ�y҂L`� �`ʉ�%���܃�y��E��BukQ�W x�J���g@��y���<rfE��ݚG	�#���y�/L�1����(ArT������yrAҫ!wܼ�a��;2����!;�y�'�e&^��"̓1��A�ʝ�yr+'5�fe�S�\>�X܃��ݷ�y2���Tδ�ቜf��hT���y�V,o����� �3]���aT�Ģ�y2�R�F�\�E�ly���j���y�$^�j�L1�Ђk�}�S'O�y�gH���Q�EB�-����e��yB�М_��	iց�
^}@��%�yBG O�۔h;D�4� f��yrnx-��;���5@ �y�����yb�W������X� �d\�"OZh�4oC���鑦 /b��aQ�"O<���/�nA�p��Op���"O� ���C�gjD��e#�2/A����"OB็��a�9S,Wr$��	T"O �s��4���Y7˃%T2݂�"OJ(KGK��.��gH6� � "OdM7pWJ�����q[�p��"O�\°��#N�:���m�e>�:�"O6�;�iH�?W�lbd�Z)�v1�"O�a2eF����A�&�%/�\��"O���ȒUԺ���ݨ?e�a��"O~�X��C1 ;B��7��([T�I"OH�b�M��ȉ��-�d��"O�5��H�3-L�m�p	D;���0�"O����h��.�� q%h�
x~���"O-�BD�9[����f�#pm*u��"Ol��� �I�~\��d�md�Q�"O�����3�K%��hP���%"O|������&��TM7i�L��C"Ot��.�2�e��!��52��a"O5�!L�Sq �ٓO
�%�"O>)�� ��P �9��һNO�"ODU� �O�,l[����"�j0H�"O&�jDڂt�Bt"".ZF��p"O� 7@�v�����&��θ���"O|���ֿJ(�I8_�e�F�[�"Oh�ハՂ72�i�WF� o����"O����o% � ��E �љ"O���⊁?MV�ըb��"O���(��w.��¡犏Q�<�0�"O��AfG�j�|�Cf����,�5"O�(�<jB�0g��)���D"O�ٚCK� �%
�e��0����"O��pDE&p�R���T"O(A�a\=!�h���Y�A �	!""OvᲡI	��d���R�FpVٙ�"O���h�Q<d�KY'_$�P�"O:�EI �+�7ޫ1􌐢fo1D�|ӡT� ���ڌ!^,ᖎ-D���2�Y<^���rĉ��I�T<�--D����L�,P/�Hrj��l�@���-D�,��a�n)vQ��&4H�EK�C6D�ؚũX�e��2��{���k�O2D�ظ0����p��T�!�&��.D�� S^�d�@x���Q6F*�H1#)D�H0�,�# ��"dNσ<�n<�BN:D��V�R��(���$�F���=D� �Oa��DbAG)N}n�9e#;D��(�2\�.a��$ؖPMn�A�g#D��XUG܉~ H���ǂ��.��
#D��r� -����d��'�����3D� ʐ�ש8U �O��
F�̩)>D��;�#������D���0D���˔2"i�DP K���H�(,D����՗&�и�g�k��`��(D�\C%gX�7�zXh7JV�11؉��%D�H��E/vY���*j�d���C#D�lÀ`�J7���bJ/Df�sb.?D�P��:OH �4c��^���=D�P�AMI�:��eH�x A�:D�4�'�q6\��Ы��P�j��6D�| �P�'L�ҵJBr}�h4D�X��
m��f%������3D�,��:>Z|��S/L��q���2D�\�O���"8�.�
,\va��b5D�Ĉ�B+@H���1'�bk�\s�)D�� xXp3.��$s��{���,)��+�"Od�栘	�.��qEA>��*�"Oxd)���`�LܩV�>>�$��"O��sF�AN`�q���B���"O������	���i��!`��,A�"OM�B	CI��QbfO����"ONL�T��n�	�����n���"O�X��(T4�0d��들t�T�`"OzxKp��6BAv��UꞰ`�D��"O���"e�>HZi�Z8X�"Oh(�G+[�}���y��LS��%"O������FS8@�t�V9uM֍��"O�lIkP�[�*e���ܣi�x`�"O:�
q�G�d����WH� U��"O�ApV�D�ZŁ��֖x��P0"Od��fa�'2x�$�D �h�$�E"Oj��-�%;(ݪ%G�����"OLi��FҒ!-Z��D�Ep���1"O-�7#D$dZ�E�H�qY��`a"O|����خ8=Xa���)DX$��"ODe ��S2V@>T�G�^	_0��"�"Oj���|H����${��t��"O�:�B	=���7)�8[�x!R�"O��`�8z�&Q1�gS65����"O�T��řX��F���T����"O��ATᅰ!$z�@`> ��C�"O�9���>���APA�?6x� ��"O1!3A�.�H娓�ާ6u�w"O����4b��iX�)Z)M]đ�"ON�ٖA��3�����%L�%v"O�@"×A��`�c�Ă�Ԉ��"OF�hpGs�xx#q
ω)�h��"Oƈ�f� �m�b��&߬'����"Op�����o�X�h�%_�9��4�"O ��#�v\�h­@.���"Oh��.2ʠeJa���7�1sp"O6����Yt���A��+�P�+�"O4�!��� &du���@<Q�z�3�"O��a���8\�+֡f��у�"O� �pGY�Q���k���$k~l��"OP١Pi�aF� W��+7�`UI "O̴х�Y��QX &G9�h��V"Of4AS�ѷ7|����n8"İ5S6"O��ڔ�S�<�
(�nÎW���K�"O��u� t��4h����$+f"Oz��0:��u`�!	�w���C"OR�qH�;�ܕ��ݤK|Y1"Ol��蟩`��4��M�<^��E"O2�z�F�+'RȲ�Z&�@�Q�"O��' �
�� O�r7"O��҆M*a:pT��v��8�@"O^�!"�$tp�,{��ïa1J��c"O�����L�=RR��Q��@�	��"O>	$�ع0i��e�O#�| `�"O��R���Y�&ˬo߾�sW"O���-���V�M�f�3�"O��(���	�Џët.�=�b"Otm1��9�L�IҔ-)�@��"O���dL� � ��d���9#��pv"O�q�G� �8�Փ�L�7{����C"O|x�R(�0v�n��5I��N���B"O*a"Pfם��@P���PsF�5"O��RUi\�f��a`@�.f�� �"O`̠U-N(#�y��\�L](��a"O� *\!�B����7�,1�D��"O �稌�+�lIc���-+B�D��"O@���@�om��bK/:,IA"O<�j-ȊF*ə��	V.���$"ODݻ���[ŲE"îC�QB�� "OȀ���e-�|;��)e<����"O �N�$W~�Q�P�X"�5�0"O5�c!�T��Vn��s���I&"O�l�񤖇_V�
�+Ѽ;�,�ڀ"O8�SeC��6����b��(8�"O�@��F�A`:���ʀ�(�r��"O.��S�O*7g��bҮY7n�,���"OD��"�2؞�Z�Q0=��0K�"O-jR�دh��=��^��٠�"On�B��м2�p���矜i��`�4"OD�t	�@�Q�;w��0E"O�!*��-#���ѮK�
��1�U"O|8
�<JG��1b��$��Y�S"O|Y#�4O�و��ڂ�bT�f"O�`H�oX�H� �W�A�eWp �"O�٘t�u�V�� �M�80�If"Ot�`6t���$�$Dv�]�"Om��Ɩ�{'�蚦fH�F��yU"O�T�%\��o�X�LT�d"ODL�@&T�b+���Q�
Axz�7"Ord�B�U�f�̛�Ekt�R�"O��P�/#P1��*.�]kV"OP)�S��#�FA9�`C7�`��C"O�]�%��O�0�`A�R�f�Ae"O�D��ˁ�Yg�̑!�Φl�>��"O�, �-O�� �@E�	&1���z"O�� ��&��1�ttR�"O����H�t�F�(��Ū{q܀q"O�zB/�[�P�*��H^ ɱ"O�I��M+��y��ƌsp��""O*U���:o���ƮnY����"Ovt�FN: \s���=R����"Ou�1��PX�,s��_�+3 X�u"O����N��~pB
�CF�l(C"O�a��`�?B�ӏ�#],r��E"O<�k��P��J ��Љ����"O=��H]���
E�i�*pLB0�y�6X
���2�L'j]�dक़��y�����mт�ȴiܜ��7e�yb�[:$<F։i����6�В�y9f�X4��oY�c���h���y�l2g��5���;p/p��gA$�yR靗otF$آǥo�D���\��y�3`�I�p��o�>�	���y¡�c�u:ʡhŞu;� �y� ��H���Q���_�Hz3m��yҏ
�\�yG���F	�����þ�y	��Ao�IBnt�h�DM��y�&��L�^�bW�ëZ��`H�IB�yʜ3Èt���+L�p]�R���ybe�(T��ł�|Z���E1�yҧ��Z�4 ���ep�$Μ��y��=��;w/�����e�6х��������Rh+�F�7�
8��D<�H���K/Z�:C���ro�І�^���8�Ixr̕
�I�+4��l��S�\E�B+ N��@�3�~�ȓ�܀��[�eC�D�]:!vJ$��	�v!�Q2a�R I*�7&e����S�? q�7! �6 �"��A�Ν��"O`��F�J<8bjd�D"�)_ö� "OT�y$�Y�.�D��o��0���$"Oޜ��Oǘ!N�H
��դc�l��"OxX1�(n��� r�^�\B�"O�<	�bd� ���P<^����"O|(p&l*�>x���.�Ps�"OIY�j�"�,��f��4���#'"OC��8t$���!�=|Ϻ��"On��p��+n[�m��[�F�8�"O,5x�̸Tu������̾��t"O���Ƭ�Z�!b��Z�V��kr�|��)�S>m�x	�TJ[:F\��p�\'J��B�	�Z~����	7�N�PA��l��B�I/I,֕��&����bA�"1�C�I��U�f�o�=��\+16>%��'Լ�Ȣ&��v���P=U�tb�'>��s�eP�'R��U��a�,���'J��� ��T4�X��-i�������0O� �����K��A�/H�"Z�� �"Oj���J�5�FTe	I<7R��(�"Ory{��*)j���)�t"�E��"O���BlW�s@�[rg�"Ud����"O�DSc ��c��X ���Rbrm��"OL��@oR��"��� Y�a^:  3"OJ%:WM�E昀4�#��%k!"ON}�"��L��p�%��	`�Ucc"O��	��P�e����e��;��<!�"O�}9qE�n�H�c����,��9E"O�L�*�h�I�7D�*r���[�"O�}BWC�B�(1��F�p�
��"O�ą� s�t��=D��q!�"O��1a�#nzf��E%]�-*v�����+LO�ꖃ�C,���eR�T�t<�e"O��
˛,Κ�2��A7݈Đb"O��G�� ��c¡�C��JA"OT�R%��C��	��oG])2��W"O�4Є`�fh��V��:�P[U"O�d�

�W�D{@�0��ܣ�"O�%���I�^d(�HV�	��zÚ|��'���'��t�$�*ݶ��MGU�N)H�'�$��!�� �Pv��<�r!�
�'P �EP]9҅�Y�9&^�
�'o��{�.	"��%�U��0�M�
�'���oC-��u�s��?@��P[�'�Da�U"��D�Sn]�1�>���'1�<�6jL+/4I�%���4X�r�'*�9�$ 
 ��tS��� &U��'�D� m�+hU���g�&b:���'��52���=M��u�6��\�	b�'���t�b��P�3��1Ht��'�K�9��@ᡅS��=��n�<AqE�8A�-�P�pP�a�q �P�<	V���a�"��F�O��݊�f�K�<	�+�2ΊL�s�E�b��
��G�<��m�_̚] 6�Դp\	�e�EF�<� �H���a�/U�W*��"Y{�<Q��ΊBd����(Z���$��t�<q6��\��y��Ň8�zN��y�'����_��С�IS�%��
�'�.��
C�1{�6�O+� �
�'�Z�K��,���f��T����	�'M�-�a��K������a�T8�	�'�6ٚ��W�����4��O>i���� X�3#�J '��t¡*P,�.l�'"O �j��Y�ik��Ӛ8��y��"O�|@�� ^p2���L?a�fP�"Or§`O�H�~Y�cK�s �D�!�'���P�G@2��X�F R,B~��1G,D������
O�ɰ�d6mĂ�x
)D��{Ą�) �*Q�M>�)e#D�����({�M9�.��<|�c�@ D�L*�	=Q0��@.�9"�n�B��<D�`�%ϩk��9(�YPn��P:D����ҏ}��)��I?d�<�aGm:ړ�hO8�	�  �	��k�>����ҵ�C�	&�dd9�HE )���Q�%�xC�I�0f�	c��X��9�M-%�h��?����	ى�qb��́	*IZr&�,�Py2!	�k�T���k�
'�ZQG��y2����&aU��XUp��]��y".��b� h�p!A�En(|�'d˘��x��Tej�L���]8
���P�NE�c�!��Ad��y(�A��lZpĜ!{�!��Ҥ!�.�F�#iid��g�&�!�;UB髐
U3Y R$�2�!�Q�V�b,��I�5e錥�
 d�!��LBnHbE&Hv�Z#�̈�!�G��I�6nRX6L,(5�k8�R7O�H����Yړ'P%n	:�"O��
���
�� ֈ�80�n%4"O��01�޽����眤Bvh�"O��h����p��]����5@rx�"O���"��SP@��ċ�ZoVu:�"O��3��PЋ�Զ3[�0q"OL���m�J��U!梓�m9<�j2"OR�c�f�qM6���aޗ,z\�w"O��%Ү	�0�cӊ6o "O��#�HӚ����'�U�(
8%a "O�\@�B��|��ti��[6~ �jt"O�X��µ8�ޘ(Ro�� ���"O\H��ߕ�n@
Q %���J@"O��r'd�?Y�����P��!V"OE�E#C��4��VA_�;EVm�6"O�l褋���h|J!ױWO�|h�"O� ��)/��Ӂn�#~<�8��"O�X�kҋ1r�P�_�;vI��"Ov0�3��I�x̠!� '�>��p"O�(Cŧ[�	��i'N $znt�"O �Ʀ�3^|Q*�nV"#qp	�3"O��!�F�uC^��E�	{����"OP�P��4:� �3�GK�-|L<�"O��X�ƈ+Q���b�U}W6�'"O<Œ�^�_�����־z<�[�"OZ��R�k���A2�<��(0"O�ppd�Y����ƯQaf���"O�X��ТV�ahU�G0d
��C"OI8��m�*�Kg��&}$0�rQ"O��{����4�2���p�9"Ob��Iǰ., I D��J�2U�"Of�U䊈(8�;2f��h؊ؠg"O@��ENP)*Z�����͂�6e��"Op����m�%�n�
p��DH�"O�c�'o���v&�;�Ӥ"OdhS��D�KX��eEV( �Dsv"O�����E�U��0 $�$\2�E"OP$�FŅ�'،K5���Z��#�"O��k��A�Ԥ��W��#y��� E"O� ��Zpgސ,a:�``�
�|�"Ort���ް;���@�
� A��$�"Or�6�W��(�%�A{���`"O>1��E�q���z�c��`���"O�AP��Xyl�Y�hմF�.��&"O$!aA͹��t�t΄�k�ֵ��"OFD�"��?�T�h45_���"O�iO
! D*&��#:�(
G"On1BC!)f$��qf�މN�X�j6"O2e���׽1*dY[���Rv�	Br"O��1�#�@s�Qp ��þA6"OXt�WE3�x��5D
�(���1�"O��Q�V�\�J�r����	b,)r"O�J'�
�1� b��'_�
��&"O$�P����i:�I�e����"O�������r�g�Z�}	4"OX,�%MިHQ�U	&��4ۼ��c"O�)��iJ�r8sgj���|LR@"O*�R���<^L�玝�4X��f"ODzX(w贠�@*#��Z�"O��c�b�4o ��"m/ ��zU"O�(�`,:�ũp.^9�T�F"Or���ث8yZ�j�
�`,�$"OF!4�2˖����$B�����"O����)ňG���[���V���"O���B��&C�L�QfӐF�|l"OZI%+�]���D�6;����C"OH�"��l�*�$H�J�P�"O(��IPW2�r����t��s�"O4���K��C��(ƉO�bZpmW"O�eX���`��ȉGK_+ T�"O�xS�ŗ$"XjqX���+u�FY��"OZ� 4��G}4icd��^���k"O���GK�~�RUJ�>z�>ӂ"O�X2��Avw�qO��@���!%"O�}����r}��i� H���K�"O�E��� #r��oR�z�Q�"O.	�6��
U��D��*_�L�"OH���C&��|`nph%"Oa)�n��W�b��S�$F`lA�"Ob����8Ar���I�QzM��"O�Y����e�`',^4��1"OZP��ْg�^q�JT�a��	�'4�Pc��b`8���s��Y�'�܈@AҵT^�D�B�՗;�`��'�eȐ�#X>� q/M��^mZ
�'7�9vl��m���CAC\�|9��'�ʱ�V�(5�|%х(�)_�@#	�'�B�:I�7Q��40r�� W����'[T�� CIڵ!� I�h�S�'�ۑ�ݍ+�����@ِQ�"���'�,Yke��Z�\�h��F�p�}��'C�L�T�e<��Ȇ8_g.)�'�1[�
lIVo+m�z!��'�40���V!Kd��ehI�6�@|"�'����e�Yb�T��*�.9�ظ��'��u �ϕ�B'�Q����.H�S�'�n����L�O�&lH����x�2E�
�'lD�Z�B�/��0FɅ�j=��y�'�愺bn��%�|͒�o�^tٙ����O �d"§ۖD���Y:)��A�WbJ/^���ȓ/���J`o�Rj�����Pb⌆ȓM$��a�D-�6���S��0p�ȓR��r��Ż$��4c�~����S�? `yB���o��@k��OW�ī"O����+X,<6�� �,)L(��"O�@� ZB8���&��:�U)�"O�=����}�� ��̜j,ȵ"O�8��fJ/|�zd���\��P�1"Ol r�jW�&��p	#�H����"O��@�ƚ/:�'e	;�M�p"O��Ä�Y����q�W"9D�D"O����[;)�)fhP�'�=��"O��1��Z<,� �{$ȝ�h8[�"O(��׹2~��q�Ȟ:����U"O�8+Q��SΩX��[*5��"OBAg�Jc�,���4�Ҝq�"O�DCFoB(&���K��˂w�j4@g"O�)�F7e5<��CW�/4���"O��#�Z�b�$��C�)�̨�"O�x�7Qn��y�a��/����"Oē$%�y �[V��8Z���b"O��9R� 2@��7���:ej@�"O����&��M�"a��:��%"Oxl��G�=k��u	�闣5� I��"O8�kB�10�ܓt5(�d��`"O2�"�GtxV�gG�z� ��"OH�.H'��x���0�����"O����a��|��hgŋ�m�~��c"O@�j3/�gTX-V]� �4� �"O~��C��H�C�5� }��"Or�
熃��(ұ�(=%Xd	�"OT`5EL�Z�H�ɦ͊�K�|#�"O�]��ME��� 0��/�U9""OtP���CM��p)������X��"O,Q7�Z��f$��/@�K�!��"O�0���H/PH|����8zx@��v"O���ݝy	������,Ȭ]I�"O,�ń;/��]��LǤ,c�9CG"O��U�N\d��K�i�"���a"OB�Ô铉0b�#f�V�@DZe"O���-b �-:E�_�F$�!"O��SI؞Z��{Ձ1!-�Q{�"O<�	�cĵy�r]�7�I//��"O�%pr�V ��j�Ҧ:��t��"O�xZ� �@?^�Y��[`��]j�"O<	���Y�F!��q/+U�Xw"O6�5�Fc4&�أBS�tQ���s"O�p�5&��&P�Q?lN.�"O5
��,^U�@,�diXȲ�"O�P&��&�� 8�Dϙ8�H�K@"O&Y�3�\�c�-zb$�9�:�� "O�(��qP0�.�vp��e"O4e���Ƥ"�uPDQ�^}���"O�9B�իu�<��7G�4w���j�"Oݸ��fd���L��un "O�ː�D��&����AXȬ�"O:1�7�������8&T��a�"O>�rf̏T�&�ٳ�+�P���"ON)P�DQ�S����ËИ>�૤"O�\���(m�B����N���ا"O,�٠ۋ1.�����\vz ��"OL�ۄh^�O������Xr2�*c"O�@��ߥr�>xj�@18���6"O�U�sme6<k��
� �J"O�i�Ci�4 팀	&�#f���1"O|81�	��w�4D32B�G����b"O���Dn�Xa���Bc�.��e��"O� N�ׁŢTv�T��̂s >��"O8͑�X.i�y0c�=\>�1q"O�а�o!�"h4�D. �d�"Or��-�e�ri�����"ܲ�"O��%P=F�t�y@(�K�J"�"OR=H0hP:�8�� �;$Jhr"O��Z�D9�f���L$ 4��"O�H��	�6J��ԭ�,�Xw"O4E�A���w0�lc���B�X��"O^����I���A�$��`p�"ON@�3mW�J��]���ȟ|���YC"O���@K�n���%��̐��v"Of��0ƁVՒ����'u���zr"O��
A�zW!(GE�%z�0�4"O" -٤va�q��D�$�ڨQe"On�`��G!��Y%��>	�6E0�"O��z�$�T��)@ �Ɨ)nvq�E"O��& 9;)���1���C����"O�X��ֈh�lL(�K��� �"O��+4BͺT���wg�5O�rP��"O�����T������G�&���D"OF�!2j�^׸A;���<��G"O^L��l8,�@���l�1��"Ovx��)U�a	�8X�Am��[�"O&%��`Dy�&���HD�w"O^��+5#6 �g��1o��}�B"O�,ydʑ�y����d�"���P6"O������/TL��F�k�<�9b"O|16�&��՘�,s�qC�"O
9k6�>�����LѪdK��YQ"O�pԈY�S��}���0e?��"O�`��.i�.�c׸��=3�"O�8/�-k�b�4!�hav�S�"OFy	�`�;Z"xH�E�� 9��"O��REY�G�0=3u���Ԃ��"O���1��(1�([ED�np��"O֝��KFdo���׃Y/���w"O<�@���K�B1�Űv߈�"ObUxv/ͽ)���dƻ2fmX"O��A&�H8j��@��O��"O����<]��R��B��ٻ"OH}��&ި@�~�j�C��P��j�"O:u�F��8,�ԍ٥)�V��u��"OP�h��΂-��X�DM%zخ�h�"Oj��A��S�\����}��"O P�s^�%�x�Җ��8�� ��"O�l�s��DY�� ��u��"O�RV�A����u�ؽrڪ��F"O��Y�)CN�
M(c�6#�8G"O�D� v��hz�k���"O�}:S��h�R�bB �)b�蜙G"O��[��Ձ_����u��23�R�4��#�S��ی|�4Jć	o�Z(G��F7!�P�|��K�>�6c5�W5v!!��<40E�� ؎{�� �P8!�*���i�m��Y���Z�!򤝓�B��b��s��1�\�{�!�ҍ�Jݨ�	�0O�t�����,�!�dB���t��:	���BA֤k��O�=���ä��g�fe0��ŃV�h-Z�"O��	�O�E��d����L��D"O %Re�ݱ4,�Z���<Vf��"Oh�9��	�T�b�q ���"O��J`�6�%9��$��P3"O� �k�;iuR�@����H�q�"O���ōHvh!@�A&	��"OX�+��Q�n==c��,i���"O�Xb�-�����I:M6J�ʷ"O*�p���LaӓJɪI����"O��c�˅�T�I��P�U�*Q9�"O��0W'�_,8�u��f4�T��"Or�C!B�c��[A�&��"O`�ā+n`2�%��F�vQ�"O��p%��u���4�Ě@�*ձ�"Oƨ���H8]��̰�.�0�D��"O��`�Ƌ�@A~x��n��&�h�`@"Op�KU!+�J�gc�B�E�G"O6��޸oQ�x�� {�4�3"O �R�5"�@p`1c�p�"O0���]$,$�|A�-L&�h2"O�dc�1N�]�7��2��"OyX3�ƿiJ���(D9"Ol�Q�3w���h � "!K�"Oj�z���j�
l��ρ��؈�"O�$�Q ��l٘6NP�����Q"O�Lb,��6����ɦx����1"O���'S�_���X���KM>��|"�'�az�l��KN�9�hG78�x(�&A	�yr�_m��Zb�ۇd�Q�B�2�yBf�)s��L��%:X̙�s�Ϫ�yB�P ^�0��"�;T�X=��☾�yb�+,����O�R�h�z�&� �yB�X7�FջdhB�F�BtɧmJ��yª�r%���X�>�\�����?����9ZFz��*��a��	��-A`.l��E��H��L%U�45��隧@��J@��1� ޥ/���������ȓ]�j�kC0^gt�ِA�4X��ȓY�b؀QBԹFg
9Q�dL�6Ǧ���,�~h@ Y|�x�Q��<2v�ч�Aq�1�(�=�0���5G{�'�b�c��Ιs E�F)��k�f��	�'�AH&��-&�j��&�P)��r	�'�&%��F]�6�an�
PHɢ�'Y2�7��B�d�MF}ʸݰ�'��e��$�0<�|(	W���p��x�'{~(�7ʧM��Q`� ƐW��K�'y@#@	˂D�%{�Ȟ��8��h��a0q�R�,5 AR`e�Gs a��WfD���Ń,BPj�la$��V�<���[��>\�#�['kB����e$V�%V!�4-�c�	�gBȆȓX��p��e���r��	�I��%�
M����P��]
��Ƞ3T��ȓ�P�r����7��D���ȓ�5p5+�?�v���v��j���ar����uHUL{�\��m�V�JaM9�ex�D	�C��X��(�P4cH�/7��G�P6Ao��ȓh&�a�n�3
YdJK�Bqh��>ljX�%���`�0�d��S�<���
%*�S%�$uĔ,h��͸0s.�ȓn�4X�@���x�V<�$��84���ȓBi�]�F��
KJuJ���K/h�������G䞗��({ry
�O$D�\�IM9W���x��� ��8���"D�0;���..���$��j���5�>D���t	��j����ŏkd �;D�� ����_8=�)���S"3)v�"O�5�!�C���KtE�>5N���"O0�P�F��"�<����R� MbP"O��Af�7��Hg�"z�+�"OD	`�J�dY.�P2c��	Ta��"O�#�+ƊZ�ᕳ<��l W"Odа�n��\6�D)�f^"M~�c"O�!#"��J6�3��ɈKWR��g"O\�#��f�&%A��'d;2��"O@ղ�`D���	��I6p1���3"O Y$�A%u�.ȀV*��.&≚�"Or9z�@�t�E��H�.t ����"O�	���8a���U�r2!�`"OJ)1��P-̀�BB�����"O�$y������DBo'A��cu"O�0���H���@cmͺ`��"O���GZ�`A�SN�;���"O��smX?i@�{�Ν�$ƌ�Q�"ONE[7G�%o$y+���B�Z��Q"OV�15�]�,B���A�XI��"O�Ħ�c}$0I#�V>n�n���"O�m�A��*@J��F��?��E��"OR�)P�X`�ԡ�.h!��"OvTJsi�dl|�W��>m󔩂�"O`A��`�9o��H$��vI�b"OZ\{��ٱP��A����`^�Ju"O�(J��7fZ C��D���Ч"O4�׮�r�:�S�N����"O��SQ�\:��l���x��}��"O����-ߜ|K5 Eb�{�e��"O�)��"؉w�F�3'bF�z`�Q�7"O:t�Ѧ��0!��2L���"O�X���_�|�|Z1�ɗgޜ� "OB�QԉB�-���u���!�M�"O��A��s��Y�B��R�|E�a"OZH����&$1��"��C5�.٢"O|�رHJ5e3�q���on�c�"OLi٧뜘F0������FRh5
�"O��� �O�F?�H١nH1DF�!Ks"O"X�Q<GO%9��G�|XRx)d"O��* MJ�n֚q�n�dMQh�"O9Q�o�<
x����l&d��"O�����;n���[�r�(ա�"O Dy���
#F�t̃�D��M�1"O�x:���_�ri�C�,h龔��"Oҡ#���"��ucVm��<�k�"O���˙qʌ�S���wӮ��7"Oր㍍�k�ZY���Î\^���"O���HP�j�FP��)R��S�"O�1U(!)25zr+�}�H��"Orթ�
�Cp��CAK�P۰�jU"O���&�
>�)���'-��92"O�Pq�	L�E�6h����*��e"O���]�` @T���4"Oz0{��up�Ű4ʒ����H$"O��%��y��P�c�$\���s�"O��C��%A�^y��m�@���"OZx��K�j=KA��&�"�
�"O�u�C���$�6ċ�8�D�h�"OJ���X���٢e�0|�� "O����̆5p�,���\-rv�ArQ"O|�0�N�a�j�a����_s1��"O���q�\�#G���t��X ��'"Ov����6kd����U�S2��"O� B� �d����љ�-��1�]��"Ö�C�R�[z���J%��y�"Oh ش�FC#�i��aQ+����"O�<c�@X�K��2�ꕪ�"O�4	1�B.#vR����<_w�];�"O�4�4o4m@}[�A� fNaE"Oځ0em�`��@�"K[�٫1"Ol�w"�:6؂RD'1��&"Oę�r'
�[����c�-Vκ5��'.0���k��bC���B�d�����'0��������Q��X��	*�'Z4�8�DD��.�`�4O� x�'��e6a�r�F@S� H�?3r���'�6lG.�		�Bj�:8N����'��l��!L#Y����VCž:'R#�'���M�ݸ���LA�|��'[�A���V!zX�FT�<fP%��'��]�P.9d�%ׯ�?:�LP��'B&i��0zfX�����.|0�+�'����P��a�L�`$ �=�&�;	�'P� ��	!0h-�c�L91�R�'��0�̒
5l\���ҭ3$���'��H���\?�(���E$_����'�l���K�v�5���
M�m�'���`���2��pp�υ	
�]�'fY���"cI�!���
��$%��'͞�������;4Mԓ�h��'�6d���Nrz���!ёz@
�'��X��Hc�5�3NOr�6���'�t�t*Ś_��Y�@cȚo`����'��)j�M�`�2]s �N�9¹8
�'��x�To�3p xKد!��q	�'�D���B" <&P�6����9��'��@R�	�6�z��� �\���!�'�� �Ҥ_<%�� rQ���M�ny��'RH�8$S�1��p��,?r<��'����e�P�@��������'�HD�3.�5��F�w>���'���)�l��`
ȟ� }��'��3�T���E��ϕ$d�My�'B9Ц�z&USϞ���
�'v@�ş)j��Y�-O�V�Y�'gr��i�B��T�sG�rHʁx�'���C��԰[���ɑ%Ƴhm$`k�'��pr�#G@{̜3&cѨQ?���
�'Nй��_�^3ȑ`U��C|Hix�'G�P6-@.b4$YuƊU���	�'P
�2d�U�dl�GǊ%!�4#�'�� a.ܽo���z�EUb0�z�'̢�C%*N�H(����>��
�'�Ĵ��`�a��,�a�����'ULc6������ğo�2�3�'�\tk�D@�@3� �Ҋ4�H��'O�u�VH�oM�i�'��)��=��'�ұ;�-�5fԨ�zBc��M��u �'T�Qç�+Y�����'�G�TU2�'&8��T�yR,�`(V�BK�|Q
�'o��PRʑ�Vj���ګKN���'���$R��^Q��h�;I��1�''����H�2V����.ZG��5��'p���� H��C�";/`p!�'")� �Ά;�D�j3��.3�*	�'��aFܨM��,��*��{8^M;�'�"����>Ra|1C %�I� -:	��� F��V�}����Ǝp�b��"O�!rb��(��m{a��ct��"O��3U'ǋ;n ء��7<_�D�#"O�1a7n͍'.~5���ܬ��=�4"O`& ��Y�A��ĕ��h�s"O��K�b�^Hj]��d�L����"O,�ӆ�Z$*��X��վp����C"OTYc�i�7aZ��"�PT�H#�"O�P�T$�4j0��`�H%d46x�d"OHls�+�-��yt��3a��]3d"O<\�ʘk���T�M�gF( '"OLMce��N���B��̍/ �iɒ"ON�[r�W�J>��[NL�`�"OTl�S�ƮaJ!�B�8�nQ�U"O����D��TK@�ӹm>|�i�"O�y�Q,�//��i���9왐�"O�<��M��%�ԕXՋ&�r�b"O�Lck6J<�����r��<�a"O�9(�h8��tfɦv�|B"O��c��U1\�����f�p9�"O:��d���wq6�p HQ����"O��ӗ��	m�
@��$y�4d�u"Oĩ�'�
�#lщ�!�+ A`Q"Oj)��́�|�<�W.��$L���"O��i�g��K)(,��E�"O6� l^�Q�ؕ�P�ԀL�u"O"|Z���	GR�q��LF0� ��"O ��5�Ӻm�\�x�.�[���q&"OB,��Lގ
I�U������"OXDA�M�zf��(��-}���"O�X���F+|���"*�fs���"O�%��o�X`�rIL�!�� ��"O� sB+�#@]�	�3��1�E"O,�����Vx��)P�7����"O�9�2�Ła����'el-Q"Ol�(�Ν�,�qc���)(Z����"O���Ƒ8��Q�J><P��"Ox4�K�p���U��eD
�PК�l����wM�"�p��09g�S!�X��$�<�ũۻl�pQI�iHHrP�I[�<�����.!z@!�fT4Z�
�n�<��f�U��8t�Z$x�B�$�i�<Y�$@7xEv�a��S�<W���TN��<�'��K���J��/B���3
�'{��R�o �}W>�`FٱM� !�'$��e��l��(b��о���0�'&�x�W��"#Y�"��\��y�'aa��`�2H)��)�%'�QIÓ���!�I)(��
��ȩ�l9�c*�H�B�	�#'�1��í9�s��S�-l���hO>�1A��~�^��G� �H��I:D�Ċ��������M'[����C 8�9Q?��0��^�n	�.O:,���k�/+T�0�e+W:�p��&�WQN�!�O��Gz��	�3j #�b����0��X(�y��I>Sth��Ѥ�*��(��؂(ړ�0<i�����iZ')�%���"�b�o�d4�S�'|�Ęqd�Z����
��(>����hɠ�a`�'y���yAaO'I[��ȓ$�P��LR5�^��U�ӡW�u���M�Tn�f�H��ŽX1��� �ZA�<� @i���!��73pb��ND�<yc��?�FX�ƮL/i�p�`gƀtܓ�=)�V� � }i'�/]X���pL]t�D2���� Lm��CԘi��H�H�`M�b"O���!\�L���2'̙�Ly2"Op8sԡ��b0��[���z�"O��fB"*eb��Y��hY�"O��!�*�Q�T�2�xA٠"O�
�%z؍�c�ػ�,��"Or!�Tn�'Yނ� B�2vg4��"O�Ͳ7�/F,��Cf��e"P�s�O�]��	��@�;P��UL���~Q��$b�	�(���)��[�6� �(�/�7J`����<ړ*�~iч/��F��M��σ7Y����4��Ն��*j��&N�2B�B��'~ў"|��X?$�"[�
E-Y�^ې�C�<���ZQ0aҡI� ��a�!�t��p=��)9т�CDV�S��Ś�L�G�a���������r�<Z�h��KU?h�ȓ6�{�'��{���D�E�fJ���'��Pu b�����}�`���}��'�FU�B��\��@/��CB�њ�'�����Y+}|	�r��3|�8����Ij����mae�-����E�bp�<Y���K�N�t�����(�
8Å!^�I�O.����.���>D8f
���y rp'���¸'3qOl����'z, P��!�>F(^�cd"OxxR+�A��-�g�ߵZԹ!�"Ot9��	�11�,a�
%[$��3"O��p��N7o`~4r�D��}�E�q�|B�)��DI���Σ-Љ�A[�S�^C��L~xlI���\X�/X%lцO���dY
)	�]�`��$�>Ѐ,ܠD��~�,�<�����GG���V���|'B$Ҁ��c�<Y�MxY���@� 4�R��X��'�dP��(O�J 0�� �끻2�Xl(T�K(�0=)��ÝnH"�S��_H�T1s�6{F��4�S�Os� �dƆ3iH�4 �
V��R���D��@/� ���#�"e�#=o�!�$�@��P� �$qv�
���8 ��E{ʟ �K�ၢNFD
��Z:eTEK�"O��:��T�S�|ك	ý<�䝘�"O|i��C#]�T��ơ�l���&"O��sP��4��UB��2f���Y7"O��&mo��XTk^Y�7"O^QhÇ?f���{D
����Z6"O\��nU,~*�����E�>ek��j�'����U¤:r-YS:1������8B�	W<� �r��*, -�)� ����'�S�OK��ۑ�_�.� �T
�.�kW�'��$ӝ3��l�孋2l �i�f�>O�!��G
@KVy���X�%뤱b��$v!�\/M?��6F�t~�h'�	l!��B�?RM/�WǶ�#�Iϱ�!�$]�^�y���,%R���jܾ<r!��ƺt�p�+e@R=\��B�ŵ
n�E{ʟ�,ʠ��3EL�2s��etl+�"O�HQSiӔ��z��ںWW��R"O,5�D��87��֌[�2b P���T�'�ɧ����q�N�p�n0���fꆙ�m-D��*E��A�ؐ�B�<�xKPEKwh<9S��S&XC�a�t�M`EQ؟��ZĊ�@�M�N�$�`��V�^��@�c].z�ઈ	'�z�G|b�i�$E���%rEX�C��C+��qq0aG�yR��+>�c�޶mX�$
�lS?��Э�Mc��O(��T�g}�� _�0�x���1U�FTH��\��y
� ��(\!5�������2��I��axҠޞ��td����@��"�y�b�<Qh�"M�ys챀�@���$�<!A-?	O<�O�t�b"(�=ܔy$�0[~B�I��0�Lk9��Sa��p�tp�'$ #=E�DhVS�^M[$��4-ʺ,z��y�┼�4�����|\T�������'P�{R"�D ���)��M�vn���'�R�$>�$�>)� �JB�y�v�CъM,Ya{B��$!w��:���3��DY�H�7M�p�� �iQ5��������'9��$���g?�nQ������S�fc21z�$EQ�<!C!�A>�`2��&�>�r� t�'�Q?����#{�f�T�7^��V-8D�p�*T J��FL�$�e,7��q���'J�z�*�f�f��\	q�F1q�����O��Q�ybA
�Q=r�/+���$����>�D$O�h��i��908�h eI�m����xҦa���=�~b�CL�0~�e)��9^=>1���e?�
�H�R0X�F+������AJli��IG�I�D2<c�@�,�$�x@kڤ;�B�ɋ~鬽��B�6���a�;C�2�<)��T>i�3A˽//aPc���ri8QR��r�L����'Nh�p#��*,��CvI�9� �E{��9O��A �2^x�2H���L@��'l�	�!�g I�9���9gB��
��z�O�cI^�>RX�[t�ɦ{}�A���'p�����8ἐ��½Dl�F'+)����I[ي�I�@A�z�
A$D�%� ➠����d�$UrK�Ɇ*G�٘���|�<)��TP��eZ��h�fhˠ�p�'�y$�W�@E]'xA*�(�y��A���û�.)KbK2�y�ꑈ<��,i��ҧ-�Z��a���y�����mZP	O�xl����b���y���b���;�NP�t��!c��	*�y�B�-?nYyDÎ[RBaAô�y�����X uH��}Gr8��F��y�,��>h�daj�{"ب�vH��y"#��J��!�?q�#�I(�y����\�0�d<�����R�y*�66x�D�K3H!zE[�y��)8?"���A@:4{��[�W��y��NX��%��$؀��Њ#�y򁙋d��]+�`^�h�$zdE��yR��0��$jE���vY&� Y��yJ�?{��ԃ�/�q-X]1�ʖ��y2)�-~T�� �.~#|�;QC��y�\Yițx��}��ڽ�y�cC�oЄT��iǰZ @�K��yB�_�{R��#�LR\�K�.�yb�َ{����Ԧ�9O|��W���yb,|
P}�T� &�T-2ǀ���y�瀛G�F��СQ#<�Xl�Ꞙ�y��
=l�b00����0u���FD��y҆��y���V�M4┴zc��y�f���m�"�T'm�[��F��y�(FEY4 �"��u�r�����y�+п@�� a-@2o�TM�����y���/p� QO�{..���.���y�*M;_� �J���vK@!�2���2�"Dy���ܰ��$"նa�ȓJ,Z�L�V�D���BA�5�ȓ2�X�@��¦c���8s��"Z�Ȝ��S�? (ё���99qG��p��u"O D�G�Q�45�ufD0�L��"O�MBG���D+��Z@�
�h7"O��赇a.n�s%`��K��}s"O"<�d�
�Q�媥)@�>�j0��"O��q"N�0C\,�`���+�J�ȥ�I�0A�`V�Ibr�*����
�	�#���m	4�Dd���:�,B�ɇ\-(1j6���U���@ײ"B�I�O�hl��.R'f52��&�I5�C�I�a���BG�+L�*���	�B�ɯ��4C��I5� qq��Y%TC�Ibn�2sJ�@5qv�N)�C��<p�&����wuҜHU@L \��B剱��P A�LkZ���F�!��ޥ�1)��|Z:������!�˨=��	�%�W�D&�2��A�!�ԗ=F�]
��1S��ɵ�
5�!�$�;i,ڜavE�1Q<�+L�!�!�Q�m�nEٱ�DA�!�p�H?X�!�R��R���L��Kd)s�!�$ȹR,xR�ڣ[K �U�Ó2�!�DO��TT��	" $gM
�b�!�d�$���8&d�/v4}��j��D!��:'���arh	WΝ��@/!����F`��^8�xEy�j�^�!��úm(��*Ņ�!p
|�9wbZ'o�!�X�+ �`3J���۱�2D!�Z�d�j��V�-��a�	�)8M!�֑p��s'ϵ;c]���S7+!�D͒{�亖HF�$�t(�L�k!�dј_(�a2v�S�A��}X�M��Z�!�Dٲ����0g�n![��^�1�!�	�1��9W�Vc�p�З��@�!򤒬.ژ,ҳMӥpX5*D�P�[�!��Y���ۃ3��-B��ɂz!�DB;w��|Ɂ+��DezRA���!�L�/sx��s��c�ҷX}!���b�>(�<B�����
�dE�ȓdB�L�3��2��ɀ��Q�j�ȓg��E�u�Sh���A�f�M�1��EG�TY"	:3�|�ƃ�=~�ń�a/i��9<�(1���&]���#�0���K
X�4	Rr%R�?��ȓ�8Psu�d�,R�n/�h�ȓkl�R#(��<�����`���+��LR���	5 )_�J��)��0s)
���	��VhQ�ȓS�����]t���;R�G�) Є�~��9ȓ� &�P�1�Е0�H���)t$��v�Յ2���H�B�7!�5�ȓ#���CgǠ#����	w����+!��4��$N+*��L��r�����vh!sڀP���p��?]N$݇ȓ^Z$2��F�N0$��
T�� ��(�<�x2G�	��9�`��w��y��4�`h�|pR�	U�Q�^Xց'��R3�T�w��y2LE�x��i�d"������#O-�p?�s��x�aᤍ�2�(���]�ɢ�h�љ��xBF�� �5ڒHT�:xx�+�!Q���O��9s@�4E]��d��37��KRa57K�0"e�B!�y���cx�,�^�t<p(��\��y��M{���R�� j
��F,D
l"D}à���h��B�I=LԞh�6��m/�l�B�>a���4�P���K��d��Dڈ;?X Fˆ/?D���,
�#]a~2%�+�X�	� ���cG�Q�vT�w�ڷT�T�C���Px�,�F���&(ƅ��pj7H���O�1�v(�;�
Ѩ��d1~y�vT�ü}�'��yr�Q�ta���-<����-�yҧ�r�h�����m���f	�D��Lۀj]�c'(R�1bnB䉖��5�a�Z�
kʀ���ф{z�f܌9wE_"����Tܨl�)]:s�v�)�G@<3��~��\�XasA�J�j��5(R�����B1�!��U����X��
/Qì���ƒ�B���pP�OF�%V�d
�K/�r�'Z�(yQ��$B:��0ɏ�M�r��Ls�:䧝�=��}�S*D�8��\Fx�WJ��x3T�{�O$d�h�艋�U8��O/��B�'Fz�($��2)�HA#��F-�$	D�׎@�`8�B�10�	`����������V�|�;4�3C䉰	���J�$`̡�$�I����	�~���R��hI��F�>Y�@B��B��h7�\G9����	�}���'�"6�$Aג��m�JG+�]�6+ϥ6r)�P8fP!W��6��S�Ok���2b�i�8TxFBθP��1�yR�R��q6F�8*$J����Eܧ{Q�!!��"9��
6�*18�O�zU��Vgz$H|�>���0���Ԛj���
�c �bk.�Q��
(*}B��FiY�q8�G�4.G�?ab��|F衧�P|\�X"DòA����WA$�O���HC��ȁ
Pi�	|��[��O��8ȘA��*����7�0w����H���ȅ`��
���O[ ���

BB.ɰ�&I�[ӦYS
ϓBA&݀4�5^߾iE�9�:��+ա4z� TE�Tæ�&i�H�V	�#�DY��xe,�<E��K�7u8���E޸Tht!��L���Tk|59���g������R��j̧�~I#�πH&��{p�4򠘒�]��H����k^����~�?�'�>Wi⭰a�Lw�հ�hA)Dp��e�߉^( ���z����Q�q�)�S�^�Lߦ�+�� +Z�d{���'2��T����p?�R�A�O��� �87!Pu��,�T&�äj�w~���T��,dZeB:�uǃ܁Z�ȸ0-O�4��j��I*��@��a�W�E���<!� ��I�D-A9T�F���\���xC�H.E���5A�f��5�5"0��%k]��S�OPP�qsϑ"_j9��.�<`:Kd�u����愦-�Đ�g�Q.��UX�-^p��fP+Q�h��`K�Z.�xUl�Vn�H�Hr�
��1����'i�E7H�]mn5�7�;Rt��F[�t�Q�U֢}G����ELh��ȰiͷI�B�a��Z9�h�[@Pz��!e!�$� :ԌIE�ߛ�L��ֳ��"��WL�y�m@+;f)���!>ޔEz�o~͹�R�:CD��b%�Zp�����a��\�d֝h����+�X�f}#K7Z�,���GF�[����+׵2� ��D߲q��i��O#�R�A��I8qO�(Y��ܾ���ӧϓz�HUꍐJ��'�P�CI^�zl�"O�NL�ȓ�h�;g���U�z�FL0&��*1�V�qbHA��W1Hg�4B�(�>5(�w�6e+P��4F�l�6�����'�R�6 ��o����H��+��Ū��b�p���	\����+����$@*ғhR�{`�M$p�E��[�p+n���ɷi�\�pQ� 
t�j���O#R��UK&��Y�lV�kp�R�`%�OzQ�)�VN���B�U J��6�ɫovM!��S�WO���2c�ł��k���V�(
a��D24�z�K΃�y�� �� �Gfȱ.��3�.[�}P��;�
��xl�������?!�%R���i���:�d�9m��p�Pu�4|�ȓ]�b}�0�̀%�"�(	H"Y��,��m��������6��0���LR�'o,Y$����&pTʸ�%�D;e�l�82/ 7	N����=�<xX�\�3�N��@HQ�[�5ˑiӃE�U���M�#�>DD��O`AҤ
B8(�����@%B��ɢv�tq�dJ��:>����ԍ5g^yŞ_����"��
z�T�`3�'W�MSŌ���d�GE�'FnȲwE�5V�|�!��L'���|WfR=/U8�''(�� c݅k�� �q�-C:t́�'�r�C+Qm�� H��R8k�Y[�'��|c��m� �a��:�	�I��!�.I���oԨ�{1X ��:�O`8�P���#�,I��A$O���ᩘ7e� 
vh�%�O
���Y���#��62�����@.��T�կ2�J~�@!��,�'t�`@KA��8"Dt	�b�-r�L�ȓ2�}A��
<�]��G�-C��ϓ�hO?�%�ªA�0Yj�����:D���`�C�W����gE�,━�g�'?9	�S�? �R��� �N�����:��`�'�剃3c  ����N-�Pk��@ B��X���*�x�� ��k��
[�#>���	�8���Q7�B�@8��H';�!�W�@mX���*>zLi@+0x��$4�S�O_D�(P�"uhP�	�D?[��D��'$y`���r(l����S&�J�OR���.%6���W��L8HزŪ�e!�$Y�r9�\ "咥��բԩ�$�!�N�=7D]��V
z�)r����!��˲'���I�n�"�`�����~�!�� �5�0�z����
�-6U�	�'�^(�fE���h��JV7M5�4c�'VzRa�� � ���M��I�!��&qO�D��O�� ਏ�u8��9���yv�r�dBJ��iִ*|Lk�$W"1�J��t�R:;fI�b�54Nv!��	���K&ݸP`�nT?+h�E��7�T��=���?Upծ��(d�u�O�]k�6p�2j�/3�JumQ�h0qO����Y���&�'�x�����
5K6 P�mӂ��Pd�.�?I�����Q�m(}���)m�����_(kk�`[�/�3�����Ѫ<�Q�����4��	!cE�p�� >F$��(2�k!3�"eI�d:��������-Z��dǓ L�!�퇐RZ(��'���BَbϞ� 6D�& ��`�}��4y"��Of;r�Sn�R�1 t�š�L�N~r1�G�Jn+0�X�m����g�}l�\aaF����)�ӻK \�{��/P t�h4�	�#L
��t`�z~�(�@�H'I��|�U�,���!�	����A�+T\�����(	~6=�U����b�>i�K�#����!� �h�[�DIx؈���
b�II"��w����6�L�P3��m�\�k��~ra&}��)F�L��
�j*xb�! 4 �?#�z����Ϊ��>q�% ��)���~y0�˩7��	�� Cd���%m��R��#-&hh�� _�ȼS�(����C(�XqZ|q!�%N�8����	�][@�aςm'�d�:T��1%î3��KL#ɐs �?[>�Z#߁t����L��iڀT`���0��4}=��jQ��(qOf��M����'L��ۑΖ�Q�Ȍ�'q�P�7�ՆwgH,)��J�/�؈(G�A���R]��)��L�0r�Cբp,0�s BG�.�q�`!b2@:�B����5�O!=�b��d޽sE&�/Q�z��f��\)P��O�;V`��:�_x�Z��".��Icp���)�!<�4�bOQ6tr�M�)�Q�q����Ã8q �	6rB�����( L�ڑF@d���$ �V>��@���@i�U�ve�(k�o�2rP�H)�+D���׬�bFl��RB�.:*�8��/5�	&�����Ӹb���,�#��wNM�m(�B�ɳn�@�bV�H��\R4c��=��B�	�w�4�+cM(��h�sf�8��B䉜Rה}��'��a�n��MI!J�B剳w��l`g��j'JQz�F_:�!��Q�n0�`� eH�,e�,j!�͈!򄗠4"@�7��:V�#�7�!��W�HIQ�DԖv~V�0�� w:!��3�����G:Ol�W�6�!�G0��i���8cLA0�Z�|�!�䘦6 ���g�L�xh&+�)@�!�ԵCF�E�ϓG�2t�u�I�!��]�|�|��w��Y� �p$ξA�!�dӳ`ݐ��s/���D��c{!�$ܒ�q�ڿX���#s_��Py�/O�i�P(*AH��L`�O0�y2Ǖ�H���Sj�?:�r��Ŗ>�y"ĕ�SDaPCD�6�T�rBE��y��$+�qQ�i�.�
��po�1�y��Ⱥ|�,qɣ,]���D�炀��yB��>?���S�F�ΰ������y����.��]=z$s$!��y Ne�5��K_K��:���y2���fl�Bf�!O).{�	��yb�.�4�B�ߥ9����ɱ�yR��32��)��:�����y
� ډP��"��AE��|bc"O��Kr�`�����ċ��L�"Op$`Uĉ37���X]r�Ap"O�M����#Q�d S+Ь1�6�x�"O"����1+��\��kΥ(��|��"OP� 4J΄Pn~#�ꚓ�@] �"OT�d*��(2xxx�ۯ? *E P"O�A�".T�:X
u[с.�4$;�"O��q��@�z���fɹ�I�f"O�X��r�.�!�D�J.���"O���`��G5$���DMP`&"O�,��iC
f�`�AÞ�Opba"Ob`����SS������.@�T"O6��#ߟq�Rd�ul0�<�q"O�����9_$$��@ku��ekw"O�a%��f���(�KT\^�<3$"OLe#�ث&&��j��
"rB�A��"O�J��ƭv1��h@�h�F�V"Ot ���ρz>!�eL;/ۊ�I�"O�x��IS��*�R�k� y��c�"O���!	S"�yYA�B�_p�� "O� H5a.<��\"2H[�[58�"O���̮Lux��4FӁu��"O��A�)��D�4L��ޤc����*O0��RJPA�l�S�I�ø�{	�'����H�#cr��bѷ�t�s�'���2C���Ua����� z��+�'��@S����m̶L�1㑡g����
�'b���g(�[\LLc`M

^]�
�'��22(ݨa�$l�AM���p
�'���
���t�@'��q�����'JJ�C��K�R�Z���� l� ���'B�d�a�Q�]������c-԰"�'Rp��dUkU�$Q�L��Z6,��'i�)0��0��B�@H�?:�Z�'�l\f%��1dΩH��^,|J <1�'��]xs#[�Z�f,P�H�w��)�'���T�J; C�s����D1�'?����	�d����f޿D ��'�2�`��Y"r1�]�4
߭QM�́�'$��FH�(����Q&S/� ��'��]�'����'d͋X�4т�'<�%`�AF7Q�|��R��4T����'���C�ܣT�*0Y��B���'^i J�2�N@A ��Bz��
�'Gle�BDE2K��p9�
G4=]V��
�'׬���Y�Zy>(hT���-mv�	�'�Z�۱<y�<!�nǵ!�l��	�'�:�+�.�7pʩx�aS����'���"@�/w���Ã�n8h���'�Lu��T"h���J�H��K�'~�)�J��9v�A�MG���	�'��Hq`+�-gw��J&.ƾȅ��y�ō��X���C"�t ᴉD �y�q6�X�c�7�n�xan��y2�ȉeB�#��'�H,!�*�y�lI�`�JP9')W xL���0%J��yb'�/5����̪u�Դ����p�<���)��}���zt�/W�<�'͗�>�h�c�FҝN~�5A�K�ɤ:��(�'�D�����I�f�¢a]j�����-"6d:�c� �zuP��DH7��x���5� �	�'�J��N�%ide`���p���	�����,��O�=sR$I����L�xR3��� ��x�hԆ7F�pK�`��B���9OB}H���A�:L�"~���hƎ��C�>�>��C ^�<	kܒFVꘓ��ZĦ��+�c~�,��}sp��~8��2ӆ^Ol"q��B�9xh��z%.8�OJ�*��V�0�$x@��z���jw�m5\�1Ƭ¶�Px�"�e
X4��'��r}����KV���OV��� �`T��a��T�. VX��Al�$��ؑFF�#�y�gA!Y��|����fX� ��y��M�6��1Q�U��S-m�`��1J�1�R�`E��>Y8B�IF'\�!���;9&��#�
{�.�w<xT:���?���׵��s��O����MĻF��~��!\�|��4
{��ɘfF&9��# �L�!�ܑ;K��*D��
z�D{�l\�t%���IBe�!#���*�j0��1�,�/o��T�3"O��Rg�D8�tir1�B��^�3�"O�P��Z)MFA�� 
<�!��"O$Q�&�!������Cw.DS"OB����O�>�J��7ȋ�@�U��"O����(M.5@xFa�1=7�ps"O6]�፜�� �`�*�7�Z0:"ObL�&i����	P��@C_��[��'A;*�'��|S �#\%���KW���E���Az�'�t����n�3Kf�� ,�<9�4�!@��
J$3K��yp���}�X N|�>�B퉀S�t��IԼ8��S��HK}�뗎J���`�|J~�e��iH
�h1'�1I��M{��˵gif�*7�DuH���<���R �:g�F)����)��|�O�z�+[�IU�����G�8S�G^�$����?b$* �\�B<"s$�>b�<�9"�;�O�Æ��,(���`�W�
 �Ag�U�(�EB�mBEB�.�xnYc�a�<E�d䚩U�Q�$#����yE��ШO��b� �H8�e�����fm���t�H�T�����y:ʓ"0\q@�Ӱ*����'9�HDC^�z����$ȒvP2@��'�ɃE�V%D�&��O1�6T�2Ð�B���;�jD匁c�U+mWn���*+�O�Q1'�N�dM�hޡ	)�ͲC�>�d�Q�EJ��5�3+����`��M��K,O��&JCx��: W��0��c�9�p?�2B�-k�rA*�#DwP�;U��(��U��.��=JT�U;PrP	!B9���>@�ni�D�g��[ ���N5�>	�HVeJ�P��۾�z�'xD0�5L� R�q+ ��.80��O�,���_ujh	N|�>I�b�{d�a����7X�����o�H}�M�6=(�ђ��|�B E�$bI���ճ�n�j��$T�TBf��y��=j�!�dR,M�<�G&ШA^�=���&G(���SP?�r�I\->!"H~�=����~}�I�g���4�BȓQh�Ah<�3OP�8q@���4a�dH`Эͯq��۳GU;C���A�+?r(����bLiᠬ��b��y�Ó	nTY��n}R���iDn��!ކ7�b�`f㗣�y���y� ݉ě�2�*i��.���3�$A�U� �o�,"J�!�YJ��@A�1�\bvj�s�<ɖ�ăq�d�R�D�^� @�$%U�j%Z 0'N�*TmD�����NUF��(O*���	NIr��3,��A
��$�'�0�T�!t0dSA�DDEIH�
��a�*_�2 ���T���>c�:n͉��3:��[ǫ�y�'�^�+a�V;kə���9��K�[?yC����Q>�}�%i:D��b��h�4+c@�Rz��&.�T�!M�5�: W9ie��F��
����k��L���1�$&��5�����'�Ŷ@���a�LF�So�` ��
}�Rp[�JS�n,:��\AF{R.B�<�~t��ʀ,��$�s���p>��N7h����gO�Wzy�@Y1G:�����(D��x�h�*[�	Y7�G��S�A&�j�u�C�)^�#|:Vܱ�S�m��S��{a^u�<�F������ɏ�7\`C��N�o��t  I͸$�� �O?�$�/�����&�����|!�KL *vmȘI���r�̓dZ�$�1iE�PbT���0=Q6LS/2�q���=C � �l�WX��H��-΂m���W|.WhB�^�t��a�Q��y��U
I ����b�ܩa�Ӳ�hO��q����H�� 2��8)Q��봢�H�P�"OZ�P�"��W_�k�l� ~l�}9�"O��CeO��cW�� �-�,1Y`�"O�`HhB�
A���ZR&�5H���y�E�"|�E� ��0pG���yB��
�Z���yƚL��e�9�y� �= ��1SV��NB IIbo���y��?2a�8"$�<A9HU-N�y�"�$��qU�I�G;�����y��[H��2��?;.�d�����y�JР�[�Ç�ѥ�y�e
�X4��yk�ld!�e�*�y��L*8;��!f��i�  �U���y�JM&1��%i�a�3f���+���y�L�Ü*硏�[����-�yB"
:dF�u ӳILU@$E���y"���m�D���j
�Tc��S��G�y2���XXy�jYF~�H TJ�%	1��jQ��D����I���������y}B K��Wn!�I"Ad2eb��wZ���H�g�� �#�\����$i�d�SjQ1k+��Z��Z����5HJ���A���~�۳)R<rW�Y!u��F�΢[R�5��{R'Qm���dr��%S��C55D��iן�1O��2�)V��Z�1��)�@'^(ꃉ��7m�2fL�L��y+$Bţ<�j��dҰ2�a�Q.K0Q��y�kB!.�>=K�n�� �' m��'s�4�0��)Z�2`�5!�>��jA'4 ��`�U�)�#!�a؞�z���c`$��Xj���QK�3�2����H2%�2���FȸJ���hS{˜�*[m�S�'P���ʷJ�!IM��j�n\�n��i�=Q�ֶa�:�
dNv�@B"�V�s�vi�ޟh�[�A��&��!��\�	������P�ѧO4��1�%�3}b��y�R#wJ��\�B�A�f\����'�U1�yҊ�A`�%��x�p�b�.^:a��ԳfK�3`�j�*΄VO��+.�>m��D�*��,�� k�NI�P�^�:1��R���=id0�VL�<�CØ�*��0����l�Pq����196�	>0�(S`I��M-�-Yc�
0ޤ��$�wA�����6�yH/,���n��<(��\-j��)�b��$�"���íWb���v�8}���G�*���	��e}X����-�'.B��6K��:�^��`��5ӳb��o�n�F�t)���X�
vU��lA=�X�����-��O�}iT'
� �J�� ���-�	�p	X�C�h*��O�eI�� �Jʼ�?�9�^�ڃe�p��l���ߧ}I����?]�)!G)*�OT����	Gdd���WNT�L�G��N��H4�F
;\��?+*�|ڀ4OP��k����d��Tx�h�� ��D�,M���Ͽo�a{�Ȕ$�����O<��`
�w��ݪ%CH�|���"O��1%&C��8�e֝)�`!��� -��)��	ӮK��U!�ͰL/vIP��!�Џp�Ds�J��AD����sh!�	��`��Ez�JA۳���*t!�Q�:�P8#��0�)�7Ã�S!�ѵ'�8��L�joT�B!�9M�!��M6_R������RD�ܨ-�!�+�����G^��=�L\�*�!�d�d�r���-�H�ؓբK��!�O�`����o7U�(�r���d�!�8e�$P���R�����$z�!�Y/w�0qӱ˨���w�\�!��
W�x	����K����И~�!�dX�@a�<����4��h��Ĥ'ǡ�D޾�d�&@(�8�$Q��yoB�l������V�0 {��׷�yR�?�<R�NV!	����R`��yF˕~���y!���4�DT�#A�y�&Q�[
�9��S�3�6������y�M�%{�0��cM�4R𰐠E�y�	>x�x���+��0,�3�I]��yRJ!gf=�eX�>���O�y��6/��aV��(D�Z���g
��y
� ^�
)�@XȊ�h��a�D<�E"O��4j^���K$�C�E�4Љ"O�c���!���S��m��Y"O�@z�P*�d)��ER�	�P�S"O���d�K�	����	+~�N��"OȱS��[�H
�Ap��[w�p2�"O�P8'��7 	'��Y~�i"O�i���WmE��Y,��rVf���"Or��
бs�h�
a.�.9���"O�5���͑Zoj�є�� ".����"On�zDH�/s���r��N0��"O�����	�@�3o�Co8�;�"O��!kź)�hP1̙N�e�"OJ����r�!�BL(L������3؞�cW��-<*@�yeɚW?��2���C��t���:Z��2f�U�z|F�V����fױ#����#Z��|�v�s2p5�r�d*W	��07cP�W�l)'@
fy��	�|��e�r$XLSV'�%f(���G
��?!W�%?�|���.��N\P|���M�:�^Qp�e]-Eb�$����.�h-�ᓵ��2�&Ǥ���.�=&�\S��J�.2�''��'��&)�V!���`���� S�H۷MҒj�' ���O;��@+Ņ��{��h�a�O�P����x��*0�<
��+�Zyx姖�r&P@;U��)�����yr"E4S�b)���ZQ?�Z�E�Y�)���kg�;�����Q՚ѐbj�>vpD��S�O���aS�;�J�H1Ώ�4 ��8r���@4���T����Q>�3$i�.1r��ˀć3$�xc�m��C���O`� � �F3�:��O��T
%��,�YD�>�
�9��
%P��䎢Z>��1F��|���j%0P�ehG�9ϲ1b� .	��	�C:ȕ'&�~�۴?!tY��_�f`<�[d��{$�nڮ+מ������H�S�S�iu� :���W8��T
�%�VQ�F�O`?�1��'Ri,m:�)'�S�+ܘ�ӄD;���7nq �<	�&l���=%?)�婀[qZ��C��:W��3s%=�U���O �i`seċH�l���������~���fX8��Cn@
E]���I+��'�ў��(B�3|-:p �!�H��a��'�<5�ǂ#�)�'.
8<��/ֹh��A02f��)dM겠���'�a�OG�>����C��p}��'�'M�Ox���i3��G�Ɏ�_SԠ�u(�{�F�ka��P�'�rO;G��R�ӝw���26�J-BO��`�ۜ1�2��3i��c��DѮ���	�>�$���/�4x0�S�CѮ�c�f�(�O b:���7�~D��J?�`����]dBdJ܆u��&�*D�D��/�?��L�:�$p�%))D��Ť��\��P�Ś�d��pm'D�h��)נt,�E[ǈ\�buÑ�)D����x+���n���c!T�!�ߠؚ�(���z��[rB@/�!򤏸Z(��*�(y� ��"D�n!�D�.,>�d.H�*��iPB	4b!�DZ.Pm`�lS8��uk�,�!���/� �XT����U����$�!�$�	�����5v�TU�/�v�!�F:4o�؇(��O�+g�׻/�!������`�,�U�Pj�H�!�$@���}i�-G��d�0�ɧ!�Ĉe�|�"�J�8o�0 b�N�n�!�DWR���9��R1�,d#$�C,!�!�$�p�{C�T�]��T�ϼ�!�$L�f.�5� h��� ��EϱP<!���;D�V<�@G�#�L�M +�!�̠L�:� _�Du��b�n�R�!���'p�xM1'�e��P�,!�ӏR(�)�1���J�1�Rg��W!�DĺU�Qs��ՏB�y�g��*	Q!�D��^A�є��t���Ө�I0!�ė�V�$�Y�)��o<�pE�0#"!�� �T��S�@�����52lH#�"O�b�Gr*`����.an�Q�"O��!ER2PR�}�%�n/Q��"O`���"�YV�%FB>"b�KF"O؜BQ�.6�����D�su!�"O4H j@��<��.ų �@�"O�`8[�V��i�ʜ�@���"OP$�H ݰ�[犔�q�y�"O�l�t��p(=�'ɚ�hX:�3@"O��eB��@^Q�`&Q4o�V�z�"O���լ�]�r�"C��m����"O ��f���9��m�CG p´`R"O���o߸\����Ƿ=���"O��0��6R�[����z�d� �"O�	��S�\w0\�îP	�(��A"O�	��B�7���T.�2m-~8K�"O>�Y�o�+y�������`��X�"O|9�ׯKH!P<�#a@G:B�u�ȓo�re�Ћ��Z]���uj-FTA�ȓE��ea�N#|��ʅ@�,�Z���j!x��6$I����zq��6����ȓ@��Q����.PZ�JB�ו�n��ȓj������թP���q�iUڵ���4�rtc�/��2H?j��L��CQ�X�re� 榙r���Ny�ɆȓQ��}�b����"'�L)5����Q��)c!�5I���4�G"<��I�ȓ`z�tH�ŝ�m��X�"A��>eN�ȓD�8�aA
y(�+^;A�4���u@l<[�o�;�fkd��UT|��U�����S�.�i�Iޱnd��mc�,I�.P�HV�H0�-\���ȓ.�xc7�D�,(jΞ�^���	| �
(+����D�J�i����m�Yh�����[&T��}��#�@���@V�0͌�J4��48��3j��B�3�X�0æ��(�j���ŀyR�'�0�T�÷1��1���@��o߮����o�H6ꩅ�u��9�� S9P4Q��=!����?�����)�H�p��,�̆ȓ!�kǭ�2"� \05&Ƶ%4 9�ȓ_��p�vߏ9��[uiծ��q��,O�}�/�7�8�B$ڦy�Lԅȓ(���Ȁ@����"d<$�ȓE"ȋ!Iԅs?�y��#"PH�ȓc���p��Kg$�c���!>6�ȓep�c��m���{1�m�Ԝ������@���s�\i�ƚeo�p�ȓv�:5Zt������(WNX�Ar4��*��(�Ue%�<(Z��UK��|�ȓN~����xY8��dS�4��ńȓ 㾡�3+�֍��4l�$��L��9!N?.�l 
f)0�V��ȓ|/<��̆�P���	ƀ@$JĆ��ȓ�(��S@Ϯ��2
GpR ��cL����
I|��1��|Z|��[B�a'O���Ǉ�!�ȓE��hb1B�_�M��K ����9|L2B!��tG�(���)�I��S�F��ᡈ�7��DyR":fP1�ȓ},�C�O��1[������(��ȓm�ā�4�8�.9a�ϊ ��d�ȓl��ETMYW��Wvp0��S�? �ii�ǜ�&j�8��$Ft���"O�����J�{d Q���8d@���"O�t��eZ=.�@�3 �>Y�D9b"OPP�6�� Y��0�A^>�5rF"O��U&�m�� 
�g�r>5ؐ"O`�I��O�_�RHStg�7P�LaY�"Ozp��� <D�ĩ�T�O8N��5+ "Oz��
5�>��"ʘ���m
�"O��"�0~;>��q	�|6yjB"Oz�m֗a�|�2'��c0N�Rw"O�Aӌ�2�]S��@�4�l)� "O�mcՄq.��@GҚ@k���"O�)�T=
����piN�r"O�(�'�@���1�e�4�J�"O��8!BёS�"����/<Ur���"O�He�(�����|F��ȳ"OȱQ'�<% � �-~>�H�"O���d.D�_����CE"¹Jc"O�!Q�R�}H�h�Q��P�~��!"Oxp�D��|�C�I's�,��"O4�p�^N����V�ݿ*��G"Oz�V��r@�YW���0(��b�"Op$"��Q�_� �#XJ�
!�v"O��z@aU��
w"V�S�E�3"O��j�O��}R({���6��P#"O�qEe�;��m�0�%��D�F"OF��#�ʷg�<�4#D$k�.��P"Op�Ò�K60��ʲL�'�����"O����Q�	Jd{p��Z{Dp�%"O�Q[撚P�t��#�Y�T�"�"O���w��:3��U��n\�"O��r@�M`��F�,�Y�"O�����_;��cCeu�<��"OBȒ4��&rD�ă>*H�8�q"O�Y��쒔EGl<���A$W�섣�"O�4I��(M�)P�H�"&,��"O�!sAA�`�&=c�$�-^�P�"O2/�*�H�e��)�`u�`"O��'�$"��p#�OvI�y�@"O���J��TP��B�)5G�ȣ�"O�1�"�˅@b=E��21n��C"OX����9���c�m��S���c�"O��
�J�o
V��Q�Y�* �"O�d9�a�`ڂ��
 ��Y�"O�P�mS�E5�|h%^0� S"O��*re�IB��{0�.x���"O�m�e�_>&M^�t
�*7c�uz�"O �A�����B9ȕSE"Op|+tL��a_�`8A͉d��q�4"On��v�M�%�p�	yMtAY�"O�ɲ��#�`�-��
��� "O��ߞ�qA5�Ӱ8�\�	�"O5rG�	�(����+%��� �"OV�g�O5) ����i���P"O�H��)�.��I�R'�:+Wv9a@"O�P���
B��kc�@ )e��T"O�L(�bE��0�s� �pZu��"O���n��Q�WG�ma��(r"O�@U��u��9��&��JJxP{�"O"����:�e[��0H�c˟
Y!�D�H"�mRcB�=k�y��C��Y!�ٟN�h Ӡ���qZ*r�B^*�!��T�'ĺ	
'o��cK����Y.�!�D\<`l�4���H�;�ؤ�$�!�� �ܫ-�+�n���̇��@AR"O&���
��q
aN�g��H"O�1K�^�C��Z��	m�E!�"O$�����bk�E���M.h���Y�"O.�ȕo.D�<�p�煰&����"O2h�FK��}NP(Q�I�*h�2�"O}�`@$pUt�sB�q}.�C"Ox���/ ��e��G�%}���"O�93/\�&�a�0NRSk �q"O�4�o�R(���n]�	�"O
:s���>�&T�VE5T��Ag"O����b>Y��W�4�V|"�"O� "��F�͢"�A�y�"Oʵ+'MX�J���j��_>n��K�"O$S�-8>mz䌍�o�u��"O����A�z� �5%��O"k�"O(TyC��Ԭ��1,(�`)�"O�EHҏ��0xM9V�؄P ��"O"�kAS3j�.��R���W�
�p�"O�l�&K�uneر�KO�<(b�"O�uqE��f��SV� .|����"O��YW�;-n���::j:L��"O�aa*Z.r�\�t�Ժe�5�"On�� �B���F��/�5q�"Oެ��g�t$��ES3Hf��"O�D��̴�V"�(g�� �"O�|	'�GO�I��
�-����"O�l�d)�,UҐ	�*Չ����"O��+qo��|�� �ɕ ̈m��"Ot0� ��F�|�v�G�Q��0�t"OHj�,XX�p�f(ҚC����"O�4B��ԣAl��W
P#N� �r$"O�����;wB��v�([���°"O`��$DE�z���M�f�"O��j'��rQ
5[�Ғz�����v<i��R�/oNqV ����(�ȓB'��@uE?��LigI_�z�B���E`��QW�Q�D�$�"�P9ըЇ�2|,њ�.Q"p���@ң��H�ȓ�@��J��S�hB���6N����ȓ{V
${࣓`6�1E,�c@p1��\�4���-�4�x�vR����ȓn$�!����n�ɋ'bĈu���H�V�� @�?�   I  %  �  �  �+  27  C  �N   Z  �c  Jn  �v  8�  U�  ��  ��  l�  ��  �  3�  {�  ��  �  �  ��  �  j�  ��  ��  :�  ��  �   N � � �& 4/ �6 }= �C J �K  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r��EQ�( �gVlɦ�M,H"�O��@Pg�9^��@9dr<8�q�"O�Q3c茟u4P�뒤���%��"O��$f�2����� �IY8�(��"�;�g�6��I؀)?D���嘈p�l����J)�4rŭ|���=E��4a^dX�(�7#!���O�iV��p���%����'HN�+���?�|��v��6��lp��~��˙}ּݙ7�I�<.��2���?�`;\O��'�LG$�4[����G '\�Lы�������I~���4��;���5M]��A��D�>���O��u�T�Ѓuk�a�V�ѸC�00�L<�N��E�����̲d��b9���3hY��~r�)ڧI��q�ȗR��z�	Usv�,�b$�j�����d�7JC:�H��B�{�L�I�&J8u!��L$���W�۠T������,!��/��H%,����P��/32d!�$[�)�$�`A_�-����2NŽ_!�d�$
�8����~�D(��B�^!���@.XH��ِ\��h�w'�4`�$�O��J�e� C�,�B3�%}u�	 �|R�)�S�PL�Շ�W�<��E�����B�ɛ����Q�X-7	����E
%�bc�䣎���W�	�5k*�	�E�¹a%�X��<C�)c�T �*�e�ƌ{R"X�'v£<Y��T>� �K$&e�QR��-7�<�Q�+8D�� �t����n|E�!�
�I�I��F�'��>��9�F�m��lP������f�bІȓXn`@��fI�Z����$*�9h��Q�ȓ���dK��:��p)wJ6%3���ȓg�0=��`��yM��[EeN	5��ȓu�ܜ�Q`��|R� ��e�G���ȓ?T��y"̔�{([U`�,s�B�I`�0�3�Ŷp,[�D_���C�I=\M������a���R��P� ">����D#sG����ϺY�$,�P	�(l�|�x�᜝sfQq��1Hm�uY�*�)�yR�V)~��1fb^:NNԺ�#ٌ�y���d�B̘��3ʾ�0#�A���'Lўb>��V�J%:�1o�RX��B'&*�Oh�� C6��g��D�j*���؎B�	��x�� V)3\\a�En�B��:^BD��l�*�\؛�Jp��`
�'�(<ZŦI�0!2=��zy�		ד���<A#�3����Ձ��D �]eB�F�<1G�^�=3-�a@=4�hۧƐi��T~��6{|�2��B��ܵ���(+6C�I�,Q���7g������	A�P��Ys��������&2�J���!�ˢ�z1L=D�T:��;7s� ���9@7���*6�#�OX�)�(R=o� $Яْ8�RlA�"O6 �Ӄ�y��ۘB��es�"O@Hx�%�>��0S�ߐl���P�i)�6�Oo�רO�er�Y�Z���c�@�,E��(�S�'e�O�6N�{<�H���L�|�9j�"O�ыF��07c��M)֙��"O%�Q×?<�dЁ�8r�iڂ"ON��S�j��\���+aT�"ODq�R��'Nr��O
�K���"ʓA��'�.ܹ�Ö� �b!$Æ�av�)����-��
�"��y�ED��IɈ�DA��H���]�]�X �ưo�jdp�e	2f��
O�h�C�S7f��#G`�9} D�"H>M���y�)��}�Bʩ6򌙗��D�=!����p>)L<�d�!=y�8{1(�4���2��<���@Ͼ��w���b��� �R���G�fzӮ#|J��וp:���W�'_�� `fTF���w�'!�O<��a�O�H��p �R���"O�L��͈|h�q�QO޴A$����Ex��#�φD
H��" M$͙���	~���O4�5M�3@ɪ����r`Zbۓ�'ՠ}��c�D/bd8�)ôS��ً��'�����%	"���˙&�M�=����~�%�&��$/J	Y��;&g�!��ߣ+mHU�cn�t�$6��Way2�k��G,�,Y�q��� #kV"��KC�<�!G�(0V�aWI��1��k���~�	a���O��R���!��i�SA>�dCߴ�Px"aƄ��`:�(��:�n	�Hɻ��>��O���ѧ;��]#FIO�0��XsP"O|\Qa�썩����?��(���Il���i
�������2pF�4�@�!�Cc~��%�U�=o�H�G%U�x�6�)�禕j��ظr�����>An��8A�-D�ܑ��^�e����P����-D����iȉ o���� �E�bD�Ӭ*D�PPq
ʿ'q�)w�I+\e�� �F%D��㕏��R�|�-��F#\���!D�L;�L6gfv�z�� Y��zl#��}���'p����(۽U�"D{3e��;]���S�? tQ9�#_�W�:(J�+R�������	B����d�{_�ء��鎅�u`"D�,����:n�T!��Z8(Uf��C�}�>7-'�O���B�z��)F̔q���P&�'!L�;H�����y�� �f�U� Vv3 4D���@��x��8�ggU�^�8-���2�O(�5�����N˕LRȂ�͟�P虅ȓ0�T<�4#�C�1�BOQ�a���F|B�$�k�L�CS&*��0yef�(����ȓ4�`�JQ��1���P����B�Γv񑞒�&�f"�T��f��@97�'F��ȓa�44�J����rWl�l�LH�'��	�A�n�?�O��X�NЌj�h���ηL�������G=j�+1~�X�b�:)�!��X�-{�M��#�����Hт9�!���hd�0@v��%Tp�D�~9!���;� !���R��	�r�A��������Oxp���Z�?������)��0�T"O��G�x�%0����n�$ �\�t���'��t�3�I>u�Fd)�F�$w$		Ó��䕊(��˓�q���_�N�4��Θ�@�d��K<Խ���3z�q��$�:i^AE{R�&�����B�Pc�Q�
�
:|�u����yb�F=/u�I�T��G��Ӱ�
���'P�{�}��d�&#�:�*q1�����xb�'e���m] 9i���2��+^-C
�'cΰ�%��!h�b=;"�Z���)
˓�(O�l:'�-r��'&K�g��-�"O�Y%dƻ(� &TA�8x�"OA�#��]t�R��:(�{""O0i�T�=,���!0e_�w5p-pr"O@E�/X���8�nēG8�S2"O��xwDV�#\� ($H�� ,lps"O���+�2�p ��!*�"O�|�r@�h��@�w��E"O"���$5sL�⯁�6ΐ�"O
Ъ�丕�'i�"���""O`�*���иp��G�R�HD�"Oh�2���?��,y��)p�
�"O��f�կIB�ď �\�l��!"O&ɪ�D��^�Ё0厀�H��܁�"O� �O�~�� p�Ș^.^% "Oʳ�B=G $Q�c�%�zq;�"Of0�� ߗ`�4�A���.q�+/�y���t��JJ3��(��F��y$�5��x�aϩ�.�'I���y"��8E^ Zq�4p�}c�#�9�y�,�����A:�dY҆�@6�y"�FWP��0
�$z3����y2aտw}��S͌-m�j��B��0�y"M��..��wG�^H��jO��yM�s�8�!)�[:T��K���y�fU\
<+�d��Z��pD��y2�E�`�b<3�Ċ$T���*@��1�yr�٣7J>e)�`�/M��)# ��y�k� ��L��I?�h �#J9�y����mi�m�7�"H��ה�y�K"eh2,)�h�(6U����.��y��.x�MR"ɹ*�$�gG[�yb$�/;A0�ӂ�\3�HI�FW�y2��1����d^�j'J��ƍL��y���s���"�$6�l�Z� U�y�H_'+��m�1)���k��_u�<��T�1X8��	�i�~D��'�t�<� l�����D�b���G�|[Re	 "O�uBG/
8]�T!���7\����"O��ZD�̏g"1���:��\�g"O�q�Vʇ�p��
O���1"O�J���\�!�͙I*��zW�'�"�'g��'b��'+��'��'.n,��&O	I����ղePcf�'q��'F�'QB�'���'o��'`� W9=�=�"כ"r�_��?����?Y���?���?I��?9���?���Oqj��ƫFI�JPH��Ӑ�?���?1���?��?I���?���?��J�g��xK�_�SJ���(���?Y��?I���?���?!���?��?1'��>�|L��� '.�R\��OL��?q���?���?y���?���?����?��kǿ�Da �,K�V��@h1H��?����?���?A��?Y���?����?9���76,�
v�A�k�����D��?���?���?����?a���?Q���?�ɔ)��=��^{��a6��6�?)���?i���?����?����?Q��?!��TI�ށ@E��.)a�H�����?����?q���?����?I��?���?��D�~_H����MD�jJ��5�?���?y��?9��?1���?���?�f���kH���N	>|԰<h�`��?����?y���?Q���?����?���?Qi��a�H�@RK[��	�ǌT�?����?Q���?I���?��g����'o���X�Ʉ�M?�:�h�O�DUH��?�(O1����MkC�U�B� ��&�+�>�5�ّ*����'6F74�i>�Iş�t`��#�Li袌�+0��������	��o�l~�0��,��v�	õu5���#�kKX��և̒�y��'��	W�Op����nUB1za��&<'4�Pcx��y��$.�ӆ�Mϻ��h 2"ҵG���҇?��e���?ќ'�)�S>>TlZ�<ISN�316��l?�dM�j[�<��'���dք�hO�	�O6l+�-�u'�MQ�����3O�˓��kn���I���'$�!�D�L�f�.���l�5CZ���U�ČK}B�'��=OX�q.4���ӿ1��X��P;���'o��FVN=����Ο8%�'vj2 . Ik� 
����:� ��sW���'���9O�+���+��+o�:h|T8OV�l�p���[����4�F�rpoۢGN�(`���(Q�hӅ7O6���O����7�7�8?�O�v����"`�hX�L�u��И�Z��h�!��4�����':�qA�Ǡļ�ȧT�b��'�6-��1Od�?i��	U<cFD킁w�\t�a������O��q��&>m�I�pX7i�
-�AyQ��������2��>��@��d��) �I��ҧ�'�283GI�Z�B��hݧs���[��'���cy�|��u��퉤0O��FҝC���ҭPn�Lk59O\1l�T��|Γ�?1��?ٴ�J~�( [�O58��������4�yR"�x��	M�?U���2���Mik���JI7P }ʋ]]Ԟ�#�'	X�T����0�3�f�b-v` �!R���P������I �/?90�i��'�ܼ� �]�|��qKc�[�F�6��<O���?��?!#��M˚'�R�'�в��!I*b��Ad��<ِ�@M����i>�'kܖ�ZUJF���tS�#R&�y��|��z�����|�@�9jB�-iRdi�9ѨWR~ǧ>9��?	�'<�O���$iȘ`;������@S�`	+��I�v(�d�D~��'�F����	��'
���44J Bc���&��5���'�"�'����OG�	��M�"E����L�e�8�T�b�lў?a̩)O�o�K��<����M��Ċ./�� 6GDX���ZS�C�*M�V�x�lI;�l� �Iǟh1V��69$�TTHy���D�P}Hw��]Ν�t����yBY�p������I����IƟ�O���P�(x�D�"B�-y�6��haӢI���OF��Od���ئ�]�e���@�a��E�T�� ��YTI޴Xj��.1�4�������(� m�t�	�����k�5q�j�"�K�P�jѤ)��'G�$� �'��'����s\�q�P�e�Әe�����'��'�]�3�4V��.O����Xh�٨�K�*�^��m��"|�d:��CZ}2�f�Do�� �2t��i�0�hQ@;���?	��1/j�h�c �������i� ���,#Rh!���6�`�Bmʌa�n�D�O����O�$&ڧ�?a3�������sn$����ժ�?�1�iz�����'6c�b��]�:O��pBI M�8dӇn��u����M��i��7mV�W;"�y2��|�b?t���d c<:5���C;RP���7�%%�\�'Hџؚg����\1j��.^@��/)?ѵ�i 4@�_�,��a��ecg�"ɪp��]��0J0V�,����zN>%?�H��G�+3o	6u�A�tm�7!*x�k�byB�҇1�v��	���]� �'i^�C#���Ĕ�f��*`���U����՟\�i>�'`�6��mW���!��1�wf��+���eDЄ0��d�����?��X���	Ħ�{�4m�2��,GA��
Q��O���EbȞ�MÛ'jh��DJW8ĢU�$���O��nN��� �`���e�xXu��+��pJ�7O��d�O���Ov���O��?���
"7�p�p4��eDU�fm�͟$��˟la�4J���O�7��O*˓c�l��ͽ_��Y s�\�$2|,�|2�ibl6��qKV�x�L�I5��DS�'�ZX"*D�f���r� ��hZα[�'�B��	l}Bn�<����?���?�@c�M�\)�.1���������?���ĈϦ�Kp+Nhy��'q���֕k�Rmpq[��U���<��I��M���i�\O�i��� z�µ����qǏ!W��m�@E�6�PMŻG|ʓ���Op����$֧$vBa�aL�"XpP�'�2����O��$�O���ɢ<9��i��ua"oJ8
(���'+ʔ9~���X�&�� �MK����_Q�Ɏ�M�1F��A�\�k��X�Q�5`�6"�����u���I՟���	p��TŊ\y�/W� Mr<��1Hܺk�n��y�T�x�I��0�Iܟ��I��d�O�� 5��7�
UysF��|)��0�v�&%�&�O����O��?UP���S�l�	e, y��J)�.H��oC15ɛ6�l��$���?u�S�0$:oZ�<Q�Ŕ�M�m�%O�ה����<�4a�Q���dZ+�?A.OJ��?��C��HqTj\�!\�ha3��'b�\Њ��?���?�/O�o�1ѶL������I�].v*�j+d�@"#ӃAB|��?��_��0�4����,�$Fg'b��#�\�{kF��+R�(%�D�O�5y�����%AR!�<���n$r�$J��?9���<G>�4g\�_�4a���?Y���?A���?�����On��VN���z��2��0����d�O��mZ5)��u�	��,��4���y���	T��8-!n/b9��KA��y�im�hn�M��
N�MÜ'PB��I����T�XL�pM��kv$Fm�*��$���'���ty��'�2�'��'�BV�]>��?���GF�R�C(O��n-~���Iß��^�ß��$oE�S���R6��0Ua���iے��DL�	H�4Rۉ���O����	+�ĨHc$��+�AsLD�aod��EǏ,�	0q�ٱ��'*��	AyW�pJ�.ד4�ja�U��a������iy�'�����4W��+�4>�|���R�D�Vc�Ng���DH�n>���tN�v��ZM}�z���lZ��MK$oڸWi�����AѸ��hY<pN�܃޴�y�',M�w���?�94Y������%I�Ȝ�T�X����P$#�
|�0�	⟠�	����I��$��e
&M���a)ƽmi|�(���?I���?1��i�~l�[�hߴ��+�>�R#�&�8�s�F�'Z�A�xRax�xm��?�qbB��ϓ�?���ЁCD�2�g:L��Dc3�$����O�������$�<����?1���?�#��kv���vbʭ6���DE��?a����¦e�������I؟ ��?	+�9Y2�'Թ|zv�Hw�=?��S��i�4!���.#�4�V�I��u"� Pa�;"� �#؛j���7R�Yh4��
�<y��DA~��(�?.OX$��C�4eQU��*R"+Xĉ���O����O$���O1�^��F��7�p����G}��jsE��B=z�Q�4i�4��'q��v��6���2�{d��H R���	!ux6m�ƦM9W��M͓�?	���#A@�)���D�[������Atx�ire[=��<q���?���?���?	/��M+�J 4�\�c�A�C� g�Z�I�AoY� �	���'?�	��M�;���s$��x����L�%P<�A`�i@�6-_x�i>����?� '�Ȧu͓toL!㳂L#>�&�[���/�)͓=+�0*���O�	����D�<��?�b��94������ì���K#�?q��?����OҦ�� h�ȟ`�	ڟ��G)C� �@%x��G�Ra�P�)�~�T!�I	�MKúiELO0�f��h��0@�!7���6O���M v�0�D]Z��Ӳ_w"T���(-��-��Vl�U�ν}!����5"��'���'�B�S������׶'���y�%�-�	襢����K�4o�A�(O��oZ{�Ӽ�3�D����j� �4���F���<ľi��7m	����ā��eϓ�?1Ï�oP���G:E;~aRD.ܵV��sS�-h�֘@���$�<Q��?����?I��?!�f�o���	�HL�:�0SG߯�����u"�؟�����'?��+%�qKV�
�=��#�C�sLM��O��mZ��Mۑ�x�O����O�:ʇ�.B/*Y�7�Qi��B�.9�����V��9�EK�)���V˟��'��	�A��)� B ��,DAt���6y���'��'?�Ow��M�4���?��]Q�`TK�b�&f-K�'A�?��i"�|⪰>�S�ii�6MY���#eR�k�Xq�Cv�`���[:y/<�o��<���6rusU����(O|����\)��4y8Y��N��~��<X&3O����O&���Of���ON�?�!"��(Ȁбdg^�K�r�C  Jޟ<�	ޟ؈�46<A�'�?AҾi3�'��!��7Wܝ�#ۣ!}����8�$����ߴ��+�M�'r�^��=��Y�\
�pC�:,�l�P���Pȅ�'5�ty��'��'��H�%.��D��F�v���ʕS���'���:�M�`A�?����?�.���q�o�HB,�e�D*X�(p�星��,O0�$lӫ�|�'��e������(V�P��10w��S�ʼ�sb�%�P�	/OB�I͈�?��g�O�˓���ZFĉVE���ə���?A���?�S�'��$C�3��&E Hx�ħ ���QL��.o�a����*�4��'���=^��o�5l�%H��O&����ף��D� 6M��e��*�æ!��?C.
I{*������ �D$�3r�]24"��,�̳�6O˓�?����?���?�����*�����`��y���9@S�$mگJ
 �IП��	\�Пd��������魯Ӈ���
�^x�Fj}��-%���?��SVZ��o�<a��͌����F"�xhZ�P%��<�qO�*b �������D�O��R�8��yt�Ù-+NA�',�oX�$�OF���O(˓#:�v�� �����Y�mU�b��4;�b��x�~m@��]��3�I�MkZ�l(%�x��tH}"�FS�;\��xuf���y�%"^4�sE� T��i��'^�d���(�	���k��'��"	4�S�S	0���!�EQ�r�'P��'������eJ�'������r�q�ퟐ�۴nNPy+O
moZj�Ӽ�DB��Vl�t��x�VX`��Q�<��i^,6m����&Ԭ �{��Y����>�B&(M�
�� ��ٝE�ExS.U������O��D�O��d�O��ēZzrAC�W�����]��G+�f@�O���'�B���'CB��6���ZW����-K�Bf�8�G�<A���M"�|J~�֎/QLI@wd_�c�vx�B5�� e���$Y |�(�S"ғOx�3"4t�&Z !�Eɰ�Q<XF�دʦ�	ğ|�����Suy��o�4�)q��O��c���cr�x�DL�9~DV�y"mӚ����Ođn���Mc��i�T3�"H68v2�!3�6�Hl�&�й ��4O`����,d��'npx��Z�;Nm�x)�iש�i)bCF�:��)��?��?I���?����O�N�z�NQ�z7p���I�+���E�'���'(6-[?'��i�O�m�K��R{������@J�M#�a�;<(�)M<�g�i4�6=�����#
 %���R����a��DbP�����J��֫OrUc�	ky��'2�'��A�O"��*\�:�4�`BU�:X��'��	�M� ����?����?i)�~�PO��i1)���  P����芯O@Xl��Mr�xʟ,�!��/n�����87�|��A�F\��8g	Y>^�>��|J��OrŲJ>�gL�Og���gk]�^LԨc���w<�i�,
a�Ի�z�3�K	?|��X	,V��	��MÏK�>4�iH�{Bf�=U6�zf˙�+��9Q��d���nZ�|�T�z��,?��ߪ
�Z�����_ʪQ��Uid)bDc�q���<����?!���?I���?Q,��`!�9|�|��%W!)�@�c ���P[Ո�O~�$�O̒�����`V�3N�m+��=:��남c�N,nZ��S�'Ew�L���\�<����
p[5�[I��ل�@�<�)M7[���Ğ����$�O>�$N�X��g.�&�!�"�O�6s8���O��D�Olʓ\集�ĕ�2�'��'� i���%�ԁV(�h��♟0v�O ��'��6M^馩�J<���,zF�3v� �f H_~"��3H�����a�)&Z�O�����(&BJ��Zw������5F����f
Ѳ�y��X�Cw�m���4r�sV#�\4B�vӐ�+��<!��iA�O���-{"��Va��bSÅu{�	�'��7mD��hٴ�
M�e˞D~���uX�-�S>��p�l�*+e����ċ	u�nX��|�T��F�_=n3JaK��8S\�X�	
��D]���-�gy��'�񟴡:r�W \ᜥ���݆/�h����ty��'��d3������p\l�{5�;c��)�
я*������OK�+D�R��g�'�>	$�Д'�h@"�”��@� J�Q!Q�'��'����dS��MS�$C	�?��BO�\��,�a	`�P�{Ҏ�.�?A��i��Oh��'@7����B�4Sʅ� �ϥ^1dI� �5(�J��6+H�!���'T������?�T��T�w8�q��� ��l�!m��V.�@��'��'��'lB�'��Z�z5,Û0H6�FÙ��H��E.�<����=���W>�0��DԦ�'�(�À�>3�)��v/� "�"��,��h��i˅������b��%{�j�t�4�K�� ov��&L�2�?a�o:�$�<�����/��j�c��~���x0,��O��mڇ�|�'��\>�Bb	�2od2}�Sa�:P�����&?�P����4AJ���;�?�� 	�KB�i����	a���y4�N�� #���8�:����D��h�t�|��C/P&��P�+</J��� 8�x�Ak�r�Q�ج���#������3"�L��������r}�i�ࠂ�M�Q���uK�`���
��Q޴l�<u�Xu~bD�3l����S�r��I�G1�i�D�Z�'4$�X��+S���IFy��'��@S�Ԁe�z����ȥ7,"�h�/h�j`p�̺<	���O�6=�����b�8}\t1�d�7o}41�������4\���O\��Jb����y��)^8��BML�"z ����"�y��	)������;��'���P�	5L�,k@���G�0K��l�t5����8�I�p�'��6M]�/N���O�DH8L��(1bi�$hcܨ S������٫O<-m��Mk��x�Ew��*���%�T0s��א�y2�'X�Q�f�hW|)�\�l��yJ2�@��lRa+܂M&�zU*éQ���C7�@��L��������G���'�����}ݰ�����1�� �G�'>�6��v��˓h����4�h�$އ~e�O��N�b��'0O�tlڟ�MB�i{����i|���O�P���2�� ���T*Q!8�̔�`+ c��#u,%�d�<A��?���?y���?u����ҭ�R@�պ3L������u���V]yb�'J�2�2�#ǙMYH4@A��:�X�g��t}B�a��Un���|������	l�.�j�e V7FU�0�$C41�M����d�,m	����(7괰��[i%�t�U��0%B��cOξ'v��e$�:>i��)-�\�EY�[R�m@s`A�<�2-�1FŨ.lY�"�s�����T�_"dra�v"0�1T���X�1���ƽ\�O�٨�K4�TD:�(M>�4M�$晈p�4q�Gc����5Y��k'�>io>�PGj�85� s�N��|�Y�5`MO�n}��/m�\誤� U�4�l;R�~�D�X�!��`pB��3R� C�l,KP��o�=K�aB,}�g"���41���$� 6-�7@��݃Ӭ�,<��	�p+�P6�$�P��v�	��T��&�\�	�{J�M*p�� .oTʑL"5Q ��޴�?����?���?���j�"���?��'��4�${��h;�%G6v�8�޴�?L>9��?A����N'� �l���}8��'dp��#x�����O0���O�)��M�|����?a�'h��=r6�8a�0A C � z��0�x�'5Ro�H1���y��T�27	�%�f���/��?��C�i���'����'7"^���SRyZc���ɋ�Iʔ�p2��"��Q��4�?Y��L�`y	��NF�S�'�%��6?��:@�H���r� `Ӯ]��O �D�O���|�$�O,�'#�!RFɑl�:��&��N�T��׾i�Ji�p���T�d% ��dpE N����;��Sl�-m�������x8ů����	\���'��ė8	=���ߦI���hqI���t�<90��kU�O���'�2�7�^�Z6��8�ٺ�Ő�e��6��OF�2g�<�V?	��x����"#�>b�@���AH\T	��O`���杲9��I�(�	��`�'4�9���d��t�W+P��Bm�	C��b����e�	���	�f">�G�B�d�`Q����4J��Y�->�П����`�'N}��y>�K�f�&x�ig��	u|�X`��x��ʓ�?�J>���?���9�?�7�
�X���sM
k�xDhf�ұ[���ӟ6�i�b[�8��+���I�O`U��M��\����L�*�؀4�Ħ��Ic�	ǟ��I([*�b��b���x 9�$�H-k�2p[f�aӂ�$�O��+��5!�Q?�	埘�+��4�$ }�& �����|�~�[O<	���?������'���ΞMR6}�2(J+Y�,Ii�/_�el��Y��c0lJ7�M��?�����_�֘�M)��Hp��9h�Q*F�G�d�6�O���\	��⟬�}��D�@ǌ�p�m���6Ր��ަ� T�/�M���?����3S�h�'S��!t�b ��ɓ��! @����kӾ�Ze� �	Q���?Ypo��L�"�I�<Ɗ�P�fC,E�f�'M��'�L9aɨ>A*O��d����$��E�& �qkW�O�~�JMiӔ�O଱�b:���O��D�Ok��n�y�R4wU������'=��'�J�fª>Q*O��� �����9��!Bi�c�d��VĈ�h�_�$�f�z��ݟ���쟰�'7NQ���
�PƦ	:�Ւ�N�UCxꓴ��O��O����O$݈���Ipy ���@Ҙ���N�7�(�O����OL�$�<��;AE�)\#�丘b�O*�ar�&/��S�<��[�ԟ8�I6}tr,�Zڤ(�^e��!�E�y��U��R�����,�IEy"OɢDP마?��,�0�*5�@% 1j8a� ���D��'5�'��'w�B�$�ZG�i�&/ʡGL�D@�����'��X��)F�J��I�OR���*����4�Ȗh���b�-{���4�I�6�`#<��Ot��-��teh}�eR8�JT��4��Ӗ���mڢ��	�O:��\~_ i��M�G#~|z�#@�M(O$��O�p&>=&?7�̬#K~)�''�pթօ��:oZ!8����4�?���?)��b��DdI)����̖<y�ȉ;��K��(7�����$�O����O��)�|��?�T&�8:��y�M@8^Ҵm ��W�>����'=��' �#WI0�4�����O�4 "Ϩ=4�+ � �1�JI�qFHܦQ������ �b�������O����O��"e
�a��T(p�S�W��{!�Ԧ��	>R��qL<�'�?�K>	�a�1#��ഏ�JT<`/X*lG��a2���IK�I˟\�'�bFXc��-ޕY��ܯJ
�"��1��$�O4��8�����;�␉�hq�A�a��;C�R�n��M��b�l�	hyb�'�>I��ҟ ���	1O>��Zf�� ����T�ib�'��O�d�O
����x?���	9W�=)Pʕ�+��EqB
+���?	+Or��M�x���'�?�!��{�HH[��փWQ��I��:T՛v�$�Ol��P�&}��e�x�	�9�4�r(�6 ��y�q旬�M�������O$5󔤥|
��?���%��#ukp���Lm�L����h��柜��m�@��S�2�~
G�H>�T��j�
l�d� c���'	"<�Ոd�Q�O���OeN�4��@��׈cF!0�LO�nen�۟��I��h������i�OB�i�|n�>�����27�8�`�h@#i��7mZ;^��-l���,�	�L�����|��]�����ɳQ��j�:"�r�n:GԺ�����8��Ο��S��'82dL���@���N��Cd3W�F7��O����O����� h�i>����{"�Sz�J��@.��dqĎY&�M���?��Z����Y?��՟D�I��@`	� "��d�D�$�L!:�.ϛ#ZD�i���T�D��O�)�O��O(����$?*��''�7aJ�$�eoe}2I���RU�|����	Uy�"[�����@�.��9X'�]:o�}�u�!���Op���O6ʓ�?��F͌��A�Tl�U���G�D<��&\�?!,O2���Ol��?�AC����4fY4(�X��I�QЬ�Rҡ���M[��?a�r�'����iDq�ٴ�*t@�[�i�h��P,�
T�<�'���'�T�tpD��'
 �Xe(�9P�f�7�_Vx��8׺i�2�|b^�8kT�����%�ч۩s7¹X�ۦHz�Ы��io��'J��I�@�K|������d��9P�h�TK^mб!����ory��' ���bR>	�	�?��-���@8l72H��B@b6��<�'��0d�V!�~
��a��X)�N�4�vD�n���F�1�o���R�:�)��}�O��D?Y�%qC~}ZQ�͉!t�DD�ݦ�{UK� �M����?���R��x�O*(]�f�7J �n��QyKc"lӎ��%��O���<K~Γ�?�1��0�8䓴*H�t��A�v�Tp+�f�'���'Y ��>�,Op�d���Z�f��'�X�ެ+�,���c���$�<yr@�<�Oh��'J�fOblqn4q��i�"ٖ ��7m�O�й7Gz}bY���Jyr��5����p���\t�X��΄�M���}U����?����?Q���?Y(O8��DČ�"�J�I7 ��R8�Q.�\E<%�'Q�	�4�'P��'�bț' 	hݻ��0!M��#|[훚'����$��˟T�'ތm�7Kp>��/E���p8���hG|�0n��˓�?�*O����O4����i��^���d��)`�)Dm�*]x|�lZן$�I��l��oy)֏0g���?�1aw�V��q�pI�G����)qִi,_�������#tD|��͟4�)'�uKf�ՔS��pi�cK?�El�t�	_y�l�0-�맻?����֍����Y�E5>���cf��o���ڟ��I����e���Ol�ݟN�:���J�F��U�E�+8$I���(T��lƟ��	埐������I�� 2'�u脊��d�^<"�i�R�'���z�'A�\�x�}Z���<	S��J�.TJ��������ݍ�Mk���?i���z&\�\�'H�\c4KK6����v��)�y��w� �Ђ1O��$�<�����'�4lC�.��u�Ѩ�b�(��Fv�����O�D� i�X��'���ȟ��dv�	�#lQbd�3�|�R'o�z�O��a�4O��ߟ@��̟�Hc��."�`��;�lqs���M��,�R� TW�h�'92Y�l�i���'�-�x�wl˘&<z qW�>��D�{̓�?Q��?�)OĠ+C��(���A#�H�\�,{�C'!�|m�'M������'L"�'���#s�@Y�gd�	��=-�p�P�Ÿ�yr�'j�'rX>�I�WA�j�O�n�Ӈ�A�@�|��eMc�ؼ�ش���OT��?a��?�����<ѧoݝ_�����N~����^m��V�''�'-�]��S��i�OH|�6'� )�!:G �H¨(%�D���wyR�'&�'����ܴL�t�He���g����&,l:�n�����tyB��vRJ��?9��R]wW�A`@K�"y���TĹU"�y�'[b�'!�l>�y��'���|¢Â����*1��;���]�'k<̓��|����O�d���קuCT[UT-"tg�iT*�-A�M���?���<!��?A����O]�A��	Y
��I�Ek�!�֨#ߴd	v%�u�iB�'���OD(�����?/@a���5f�<���̓un�nm �IF��h�'�?Ʉ�=��呕+R-�` x"b�R���'�"�'_�$��4���O|������f��H���S�_�PMԥ{3�r��O��2g0O�S��������kf��Lv�`�� !���daɍ�M���x��xr�'K��|Zc|�r�hՊZ@�!۴��W��\�O(�B#(�O���?y��?�+O�E���
�-�,��1��&4mbI��9�\�$���I��&���	�T�$��N|~����7��DG�ї~="�|yB�'r�'��I�O���O'D(��V+���H݃b�40�O��$�O<�O���Op�1��O�u�Bk�[�n��� i�����ST}"�';��'���A0DZH|����1d�����n�/�2h�*[??5���'G�'��'����'�O�8XS����!�"!"aȔ-��lZϟ��	dy���d���N����X�TI�d>�u1$���<���5$�N�	��	�Xzh!�	q�	\B �ٯ9֨`�Qv��z��[�1�'�8@�&w�$5�OP��O�t�"��Z�Ң 5� 	����)p)nҟT�I�~��&��}bW�T�h�q�r'�::�5ʂ&צM#��@��M����?����j��DT8	xT�)�͊(~M������]���lZ�]��S��j���?��fUjx�,��
�6VU��a�=p�f�'�"�'�Ի�"��؟$��a�E�B��Z yf�^`�nc�I+�(�M|R��?	�G��|�G:o��i< J홑�i��	�:{8c����Z�i��1#i���S �S�>L�1�>Ys뎖�?�.O*�d�O���<Q©����)�2�s���b2�Q2^��-:����O,�O����O�84Mk�:kt����p�Q���'
�	۟ ��П,�'�n���{>� 2a����31�Ƽk%J�%$w����\���	{�'�B�4w2��	2��e ;�u��e�0�p듙?���?i,O\M�@C�a�S�������K�(�r	JB��� ��-��4�hO����:�����O��I���2��_�@�`�:cJ��4/b7��O����<�gʓ�4����?EB��6$�����c(�{�֒����O����O X��ĕ'H�)�D��a���:��y�	��n�VR��k�oϛ�M����?i����Y��]�)�0@H�oH.<�~�Y�"Ǘz�7�O��P�C��:�d?�S!N�}��K2fh\rfD�P7�<28n�ӟ��	ß\�9��$�<�S6M��m�����7*PWNȉ��6d���yr�'���'��d��[�b���`1E�:y��FF�K�n�H��۟��k���D�<����~�&�� �li�G
�n����k���Mc�����Q�X��?I���p�ɓ ����Ԩڳ �HM�� HJ����4�?�5�C�u���y��'������	�
�9e�y�R�����6��O�`6;O2���O0�$�O���<�uA��2A8	рg�83�@���Ɗ2B���$T���'�X�������I-k�4��F��L3&��	@ �f����Ο��ҟ��	y↍�l���H��5Áɮ���(�Ea�7�<!�����O���Ohtä;O.K��1h���jv�*Z u�BEH�I�IןH��������qɚ\�d�'���� d��-���4,U��׏�禅�IC�Iݟ��I��"�b�<�$�S�ɪ ��#9p���
�*F��F�'VrT�@㳮�����O���5,�\��GP�Q��Đ�OK".m��n�K�jl��ىb��5&Ç�4�ĥ�g��3B�|Tc��D��M���?��֏�?y����������Ok�	w��<�Qa�"H#h��5&${L���'7��oJ8�y�y��DL�Ol̹��דi���
���M�eN΍\���'��',��6���O�8p ���j�����K�ֽ����̦�A��^����<a��	�֠AHB�tQ�N�e��r�iX��h�EGyRX�h�	C?	MƉm� I��)Z9|�zI��l�#O/1O
I� �[\�S��(����81@ߎ=>��j�$g����^!�M��n"ک��\�L������O
�'�j�vA�}�4���w_�d��O<@`�>�d�O��d�O^��O�-b$�5�F@�UEJ+0ujp3#@G���?���?YN>����?��jK�2{������)��� ���	�l �DHS~��'_��'�"�'��i�џ���CV6W,�5�"RҨ��ip��'��|��'�� �'J�\�x�4i>8��W�3����"E ����'��'{�^�x�V�P���)�O<8R�H��]h��A��= �֘����	ҟ��?��l�A�*�.�`G4��]s��[��N mZ�������|���a:U�O���'N�t(�4~ R�$E6Q�~�uFU��jO����O,���5>o1O��)*�����W���ׅ�i�Ui��\�
E��#�+rE�Pb��S��� a�L������/ۃ_�$��F܂�U��q�<� {A�����]ľ��s(D�%�9��RP�v|q�mH�0�jt����jeF%����I����+C�9�`ٚ�ۥ!����_�� �i�ʢ7X�K���G|�5ha�C���|2#а%zf��$�
�TH)`ͬ+%(m���ů$�q2ĉ1 3$AP��k1O���t�����?���?�����O�����=e���E�
Sfh`ѥ�^cVt�AVn.�AF����6֟��Fy�Hϕ0Ƣ�Ұ�rL�3��I���p -6cbLSS-?	��%���?`�E��ظ'E�!�(� D*~-;��Fh*���'~ j��?1���<1"d�4������7c"9�rKEF�<1獋�X������mh�ԒQ Ͽ!�����Ğ9��ym�4Y1h�0!�ڿ�
���' ��	����L��ݟ���g���L���|2��y���!+9.�X	�E�\.��%N�U~5���'Mn`CL�'Qz�`x�ś�Ql�#2�B�"H����/W4~��䉓a��'�| �o�	���mQ�T�.i�V��|�'	Խb��a��[�I�����'�������jDۦ�]�W{z�ӛ'��ꓹ�Ds**E�'SBU>����J�Z���M��%��D���@����럘�	�d;�sGi�)��k2�?�O��)�#g�!P36� q�22�|(0���MI�`��ҡ�)tV�ti�I-�	E�<	˦63<xc�D�c�Q� F�OX�D$���@���ĮI�.([cI|f��I@��X�F��#
<��C	�F�Zc�#�O>�'��YЇN�'�@� �L,S�$���w���Wd���M����?)*���Jp��O����Oz���l�>p�}����q�L�*b��.:��iq ��)�Hp��񦵔O���y�AFG�>Hj�(F�p�$xR����[�@IgN�&�Ԩ��/t� ���O��!�ɭV٠@��,� ��cjɚ����}�nZ��<�O ��?A�
�r1> z���1T�P�0� �<A����>iA��]O��bMѲZ�d��+�_�'�7-LҦ�F�tLN>DJS*ӋhC�	hBf��3�r�'DH��.B�&k��'mB�'K���ٟ��ɬO�Bh���
.vX�b1="tt�ߴ�X1#uvl
����|F|
� p�au�o���Q�V�<��x�wĊd:��˴"u��� �ĽFG�퉴���b%�$��zr�L;�X���-W����M��S�'N�Q��;ԮOd��0C�p�<��<�	�\κ����Q���g�'Z��a$GT*L�*�\� 1�UJ�>���v~�T>Q�O���i%�h��ːˍ�r���P�&i0�Y�O�On���O^�$�E�����OH�S�^\zY)�	�$>� zE�!	��l�0�N�$!^,c��;c*����'�L4Y�l��j�FA�E	DM��/VMHj������,i�c|8�<���O(��[+A�`������&#�x���yq!�D�.���@V$��D�
"!�d���(˔���Hi��(g�SM�|k٣D�i��'G�:;O&(Zn�;̲��7s! ��kB�����p�+{���s.Ӊ
�j��S���<�x�eÉ2{WD�
���x�'ht<*	
#+I8��&䆲K;�!�/� ��vƫb����G���~�DJw剥v��d"ڧ�A+����2h"$ ̑N��u��5"l��Ǌɛ[it��P�H6�]���/�ē��@r(I�"T�ȣB߇c�F��4��kR�irb�'��Sjy~��I�|�	KS�}x�I�&��h�F�A%H^$0����ޟH�<��O�|�2d���$�wN�T�|7%&/~"<E���C�jLX�IA�-�hQ{U+!AnV�94.Ƅ�?�y���'!ba�`kU���5�5��m�uc�'�6U0�a�	C�$4�w��`7|���Y|���	6+R��(�CG*Vw�lApmd8V��O$4[s������D�Od�D�O�h���?ͻY��#�*�R���`�	-��u�w>� ���)[S@�Z2m�>t$Z��"
�nD�	^_<��d�,�J�J�kØ9!����V�^��'�V�JED]*hE�<���D�[��%x�'4]%��H��Q
��E�Y%~�xt�,��|I>y��0��f�
>�p���{����X�jn�'B��'��V�'k"2��L`��'d2(�%�����g���B�=�p>	�ty�DW�)�R��j�\��T�t�*�p>�������I�����K�
L%<���Ў"RTC�I�%sh(��
�Ɯ�F쐅<�6����,
f�JM�؅�V�[�*��)�F�|R�Μ^6P7��O��Ľ|ڡO�'�v�h���TN�� D�z�q#���?I��K�����[��ɧ�N$C�>A��(�)QP0Ţ@�΃�Q� Q�B�s����*�1k3�QK?	{N�#I��I�@h�<�`j�8�5����e�Ob�	�6�x��r"��w ���'�̤S��qtٻ򊃡�ԤOZ�=�'(�'�Z��cK
U�(т�l��G2Z��'��01g�bӎ��O��'G�@1��?�Ly�0R2�܉.�Z)�7�M�sB��B�# 8s�1��J�<JT��+��O��t�}��u��#|�j��r�8��$��+nbY�n�ş"~�	7B�(��L�4G��J`�Y�*XqĎ��4�<E���%��qw��[��A��K<r��ȓ�,m����zj�:@�,G�8%�<���8z���Οd ���O6Ą(@C+0oP% ��ҟ�I�-��0�P!��ğ��Iǟ�
_w�ww�!L�4�qs�c:�����'�~$�
�R�"�(T��I�y8�c\0.0r<�ah���I�i⪭#�OJ�m�Hb�o˯Tʬ�� }R��4|OP�����e(&�[�nJ{fZ��"O`�`l�_��b��7MZ�p��	n���V|B�
��7��4A��Ӈȵ�Z$�`
�ڟ��Iҟ�I�_����͟��'5���*�g��DV��s��X$��(�蒱vV�I�eMG$wPfqpA�'�vL��^�|�j|S%��Pm��[�O�,4TR�GMgRR�H�� ,O����'�L���1x4ς�Wi�%@Q�4_��'mr�'��O�2@����4�*�ޜx ��0jHC�I�;��aB5�"^�hCg@��r牟��D�<ifo�'0V�v�'�R>�"��"�|��)�$0�Q�SgӅ.��0�I����	 ��2ܢX��i�-]�0��� ct��u��Q������4d��  1��9 ��N?�b��C5�e;3�	�EX�qJ&�<ʓe��!�ɀ�M;d�iv�Y>�3���|�#�/TuI��ҟ�?E��'���EK�S��a��RQ�$�+�2k�'�V���ǌ�:9AT�� ���'�l�*�SD��'���a��Ο �	0h:�Ѡ��2�H��QDA�Œ�X����<�O��O>���ꝡ�^좤�J�%��i���C�O�:�K�
+�)��� ����$׌F؅з'��9��4�����>N����O�D�O�#~�	
@ �e��C�A1��H�3�0���|��	��.�c�b�Pj�Q[E���N�0#<� ��~�t�D�1����FV��BfdC�A72�'H���ň�dN��'���'��$�' 2Ð�j0ㅆ��g����&��y�L�n�h⤮��[��ybD�=X���*	��3�%�+#*����t^���F�'Sr��hO�K��\% ��L'��&��R��O(	I%�'�"�7�$�O<�D�<ɔH�O��q�qj�0K rC%n~��)�'G��iQ��%�Z� g�3�vT8��i>�7-)����i�<y�^��?#nyG��A���&�i!FDE��?9��?��2����?��&E�(��.���Ǐk]NeE�V�wh�L���p>���
�?m����ŗ�;���^Pu�u�4dR�Gڪ�ҹ��o����O|�A��'C46MR+a�p�f� _Ɏyȴi�+U��n� �'-B��?ՙ�C�<i���R�n/HD��4�hO��\�{B�\�0YҜ�	D�Z�"牌�M+F�i$�ɾ� @�4�?Q���E-�ꍈ2�U�o��� �h��+�OB�D�O���3�6e�,c�ʧ�6���jT�J�Љ2��X`(Fy2$�9*��8���CG �p�^(}l�Up�,CoQ��9�&�O����O��$�|���*�-0'g�0Z�Y��U��?ш��9O�ak�g��%��I��ꖺM��9��'H*Op�*�̬ �4M�q@?kEf�s�=O┉��Ԧ���ן��O�;p�'M��'"TqyJ<w�>��B&ԉ
:}b&#]��M��T�G K�d�>�M�O�1�2�S;%��$��8P�`)�F�:s�1��4�:L���Fq0����OZ� &)�*L*<ir��W�����a��D�O���?iG���X��H�Ta��Ĵ'�����?9�j Jl��@0 &1���2f��Gx2�+�S�4F@4(��8����;���Ń��k��'kHl����Z0��'���'�맩?����>w�Q�D�D)"*p�p�G�k3�����[=uY�\�:��,ϧ>4d�<dk�]ǰ�j��ܨz�����)u��e�˵ahjQ�ԯ��/�,�'G*Q���rD�cr�cæ�%��i2�'�۟`3� G�P��4s������O�˓LČ��"թ!���Z��ֽ��,O����ރ�6�zUH^�@rrT�Ϟ<�qlڼ�M�����V�'���a��aI��6̨�)��WuJ�T��I����O����O�h��$�O���v>�w*�\i��O�$,'0�,I^�F���� (/�,ܳ1%��<��mf2��dAßCM^Q�TB�Gd4�ڒ�I0�m7b[�|\ay�E�?��M���	U,�
CJ ,�pN�?s�A[���'��>�	�s��s'2bȔ'@�[9�C�ɵUb|k�Ǆ$'z%��HU�f�	���<i@�ES������O���GɈ�G����*��G.�4�z���'�2��y���f��a�� :s
t�c�`�x2똵Rؠ�$P1@��<���NU� \I1i�/$|�`�'�<
�_3�����ދg-@�q7n	C�'�0 ��?)��t+޾0��H�F���|�X�3�Ȥ�y��'��}��<afɈV"V�ur�p���+�0>i4�x2�ر����P�]���'b�k?9'�λ&��F�'nBT>��siWǟ���ğ��[�a0+��甠�c�5�Z]8��]�)�P`�'��Sf�la`E��	\-y3D��Vfj�&2?,]���
C(�iT#X�aQ?���6&��Gh�@A�}9u�Y�8��m�`��O�mڝ�Mk�������x��t�H�j�p��]��y��'�ўP�?��ᜑ	��P�*�� `Y� �z�'��7-�ǦE$��O>���H�t�%�b�F�	� =���'mB�	=�>���'���'�Ŧ~��+r�{b�]�}>�\�U� i�����:���b��v��T{��L�acdMQi÷�ʵ��h�� z0M]}it���Ō1�,�x�ı]�L��0�^�D�W���$�Ħi
�t�'��[�|��*1���+f���j�a�$2D�`#&"�2-]���1hJ�#� ��B�Љ�HO�˧��$4��o�/B�y`A�omv� ����/2�L�Iȟ���ȟ���,�ן����|���B"��İ�-J��tB#0�2z�OL�$�d'gyU�c���G'�� �c���KF�i���o3LZ@��*��-�
�&�X%�-��Qh���	����Jθ@9��޳^�lH�Q�H��,�?���9O���AN�+�Tʡh�a+�0`2"O���b%D7F���Q���X���D0O���'Q剸vdxh��4�?�����/�BE��JI�`6R2��U�
��CE��O��$�Oxa�s)�&c�	`��F*SSZ�"a%Zx�� �2S:26*�#̲ (��ڈ�(O
	��J6z�5�� �`�����f� ���&�jE��#t�|���(O��F�'�h7-�㦵��p�� ���sA��`C<8���{P���3��O��"|b.O��S�j�S��ۣaC�C/��g�$#ړ̛FE~Ӵ�D�<K,x-�EߘF�`��4���;s]ȉm���������qz,�����	�Hi��� �_%����#�̬&p�f@T֟P�<��O<m��Pn��T��M[�}#T��	��#<E���)�tл��>4[Ɖ�u"�a��4�����?i�y���'N �"�Ǎ76|��3�P�l:ze�'>^����)%!9��b=f��L����f���I�vfD��e���T������d�O��@ŋ@������O���O�P���?ͻi>������5k��l�q�F!�δӅEcӴ]#�K��]VU`f�Q�����d�>{����T�.,�t0���n��pz�4X�n]�f���=F$�� k�?�=�b�e7��z`Ά�:5��{4-�y?�A�ßD����D�?Y/�\���k+W��Š��R���b"O��K�N���*�;�j�h�-	�)�A����9�	�Rw�Ȏ{�Y�ɀ"IP0�:5"OB��Ы��^�-Y�>�"t��"OPIJwLT�0R�Y�,'b"035"O�(P��n�]a��["�Q�"On��CΙs��$�r¦���"O��PEUx(���K �U���"OФ3ЏI�HȌ�zc	��p�H "O�T�2�ū`!����i�j��q)�"OԄ���Z�� ���Ƌ�Tx���P"O0�(Ȝ�_=
�!�R#AmHm�"Oj���A�lY���hC.H`�M��"Ot�Y��#sh$"P��<hP��Zw"O4pS�/�x�D9؅�Α&yx""O(�{���#�V!#Ɗ[4 +~��&"OJ@�&i_�B��1���]4x�x�"O��!@�ۃ>�2�RFG�ڐI"O0���E><sX��=,�\5�C"O���A�[H�i�ةB���G"ON�Sg�@N���цd��MBDq�G"O�Ik�cS�<��Iy�@���\�B�"O�A��eR-x7R�Qu`-F����"O�	���Pa���S �EȾ�{"O�I��	�:�X�uo�*YTq�#"O0�D�ڱQ�1�4̊8#Qbd� "O�d��C��*x.rkS"OP(	R"O���)� )�6��l2j��"O
�P�ƃ�EW�s`�N�I�b$�!"O�F�c@��c`���"Ov��3� 3�� �# 6;P�t�����.sr��$��Hz�J' �����г}剠h�A��I}��((3Iڅ{���"	�U��������r�z�d��4�.}��	��$���68�*�J	Q(.����7-�T I>!�;h^�[&!H<&��
\�����M��%����'`��r>Aś~b�-H$���33�˜.�A[��̕�ēy�\A��1�)��]'��&��h �Rt)Z�sl�7�� 5P�'gؕ�O�|���
���禕�R%چ������өb�|u�'HIiբO����G�r>�C�띶T�`��W\:�{���;d;��B,T#�!��['8/rq{��(Ov�I�.ϐ|��D���|3��ʲ4m�˳�N��I���O�d��b��>�e �xѸ�#���	J�l�!�I���p��+�ng��a�B��V�` @�P
�����#�kG�`lZ0L���EI��Sb�7L���Ox%��5cO6J�hp�U� E8�@����d
q��.�9~i`��殟�F���i��:0��xUl�*n��ip�|Rdw�4�\�%�Ѐ����?�I�4v^A�`+H��h:g+�5>z�Ig�o��������=	D���v$�b�͙�FX!�C��@T(��cO�	f?؝�e�5�d�
�g�'��Y`Fn�aW�p1S@���BaG�!\O���y��(SҪ���Ő^(�CPOE�4�~�0!��x�'b��x5��Ay�Q�(}�1����[|������V` u���;�	p �#<�����ŅI54��*�k��$B��6r� $y��x���-d�@J�,��ޠ`g%F���'���aq�T>�P��1)ة( �q	�:VH�L�@�N��@�/ׄ '���O���Wm]'=��1�D��  �� !�>1U�t����	�����  d:ǢC6P�|%)��S�A<�]�u @Fy���7A�r�!�����st|���a c���kG�x]��	D�n�X ��4p�@\qX`x��OS�$B���T#G��G~�,?:%Cb��\%����A�#	ñ{Ɛ�Ǟ)1(��1!5�� �yr�,��(1H\.�>�ѓdɔG�b4��r�W�"���O�-���F�f1��Sf�2@��y����"P��d Q�")p�$�gܓ���^�>n�A�w(�!���	�
��W�ݸ�X�s��==��I!�Y�ē;��0�J��@z�˓��I�|�p1&n�r�dSQ�G�(���@+�QU�~��U�B�<pQ��H��6}Ѩ��r�!4�l��cJ_�$��A���[(kG�	���
�>1F@�zmN�uF�9*�� �ʝ#�����4O�q�d���\2fxpF�= \zɹ���R��Fn2�$�矜�{*�k��W���P'�ݴl�~�i�Ŕx���ҀO/�ē�y3!	�
 ^L/��!��f�z�i�0|~$8�I:�'���~�.}����}C����qzAm�z��]�e��>�\)�=���}�\(е��WT���|�':t+�i��8�(yyE �7z�`���2������x�C� j�:uEy�w;zQ���ݸ}q��@�C&+p.Q;��N܌���XyB�(��ɟ���O�hi�9e,V�r��
�[H��c����N�Q���O�V�p�{2*��V��eI�1FLأ!m��Ms�"!}b��ԟ�H�{*�k��.�xM��l�}Z�q��Ԟ~���,[�����T?�Jeb_�-�bn��(30�{�/�lh%8�*J6%f23�r�D��ް���ċhY�D�,QF���kř*�b(�H@D���$��R�G���y�+ڈ?<x�:W-�O�s���X"h�gJ�@"��:t����i��DY7��@ P�ޒ_���#��4�d��co�EYN@rbӂx��zE�K?�v
�3s�C�O��٠IA�������'?�A�;d��P4B��j�틻zԆ�Q��d�2 Qt	�ңQ���	�A���!2LM�5!,���U�B�Q��!ꪬ前P&�4�ɀ!���s�,���E�����/�4�T�)
)����z�^�PDp�rҧ��Ozm��H[�3\�B�+�<|kg �5bztz�D�|����צEZ#FM�J�MH|�O�)��R�T0(i	����;y�"1F�"��34� �)��w�n����ĳN�T�5GH0�*����.(GX=鐦X���4�¹x~~��>�OЎ���f�'	80ct��I�x4x�l;�	�F��l���q�?�U`�/,���Fm����n�yVh�7o�,��=�OsЩ��nL�܈��'���CN����f�j�Y��c �y��Z.V�O���3Vh�λ=�F���k�<��Y��-8@Γ\?��ʷÎ�nܘ݀g	Ā}CF���?c�l[7@����"�N$L��+�I �Dk��DЖ5��+e��2o��N��~�'H"6��|���9�����ڟa��%`�Dߧ��'�� GDޥ.�С�3.�?��"<6|��@�
��2]�`���b�I���U åH��}BT������$�.lh�\�(��+3
۟E��ɄB��ɢ/Ϲ6���DN0�j��h�p(�p� �dG�����F<1�\�{*�"Q��h>"I�Am��`�͒7�P�SZDʄ;uhN��Z���9O�	���M�W���Z��?˓�R,.<Xm��*Ձ@(�)kSBv�q#�R��y�¹06�#`/�1wb.Y�"šӘ'j>4"ģW�\�U��nQ|���I]4j�[���'Z���N>Y���m���n�D���@Q?r퀩�D(�]D������aW����Yd�e_��t�X�&y�iOm��!M� �e��� �����`���?	��K�*��Jd@�>M6ڙ��)]^�S�`R��0/������B;�扢Y�Ert!��*�:�S@I!��R@'�7 ?���䉁O�z��DG\E�B}�{*�~)���j;�#��yBF��졡U[�$�����ul���'@��5KӺ��1ϟ�ɟe�!�F�� ��ڔ&@#qH�(�*�X���̓�52�ԭ"(2ы�C̭@����<�!CͯD��j .��L�^\)G$(*��mS&f�Bh��P��W�	���T�Է2�R�����%����j�N�3FW�e��'�گbtƙ��Dp�tb����E4kdbG�:5
��'q1��a"Iޑ ��$� �0�D��	<f��CZ�A�QC�1����'89� �����p�ՓѪڻp���'VH7@Y]%��I��?�0|z-/9�,m	��D ?��8�VΆ�Qr�W�"�|��ߩ@��\s&��-�yΗqBHm��L�8��Ћ�K%n�l�Q�'�d��c��L�q�Ο�I8P�C�,{8�򱣆*k�l��@�>;!���_�j��2�V�L�����,l�8��<񗪚.h�(�@�EäC$���ꇊ'�t�"�!pW$lzT@[�0�$mxPH�*(~�z�fX�k2�����X=���ղF�$�����4Ű�)U��#[^b��iՄ�!_N+$L�I$��'x��Ê1O���C�@�s������@���`�~�U;S�*8���'{GƐ���xU��$��pdӝ'��Q��`$	�%E�d��P�xuRh#"�L=M^�ܛ`�Gc�
��S/�⸧�I�:�ɻ3�Z�fF���!Fʁcf��m��Zu�X7oMJ<"t�}� �T+ޫQ/�U�V�%�'M�X)�� �Ge��{��O�3<@�E˨#���Z�0O��;���!4ߴ�8�������y�����'�ԌM�1 \��Z�"�|��Ir�H�*A'�	�l�ƙ���O�-�ť�O�Q��c����X�#џΡ�'�p���1fnGRL�!W�`^�SM<��G���O���;kY>9���ǘ���Nу����3K�|��5	]l<Z�,+�>��'�� L��S��*�]�Њ��p����i?��Y@�7�ɟJ��Q�R!�*Xl.=3uL��>HZ�˂�Կu��������ا�� E�������?k,�ݻ%��� 7⛑e���J&�֯TK�q-� *,�ɘOe.� ?R,c�f��p�hң�E�Z!�l����mb�y�dуQ�l`� V�b�zpZ���yE�&Ip�j��Τg���oQ:�h�b�m�)���$�;z��Ǒ>��'�禩r��<0����G$�P�u΃
gY��A�ލ=�¡!h�>����!��?q�s��x �*����M� �����
��Ps�O�-Z���%_FX�`b�HF�L+�	�4
Z�y<�E��'�<q��i�R��4K��``�@V���	ðK�<�O��X��f�!]��[R`S� <Q�eX�pQ��� j&�`:&̔T0�3����hcW,T�LO:���if�`s��3-l��H�PE?����R�|>0�;�Z8
�O���H �e�d\��Dx����]�x�2���(%�p�&��"tI���e�O9#��d�@�Y$�8!�O�,\ a@��?�A
�3y4��#�2]��=�s��9�!�;n,6M�KM�*Y��I�jݾg����Bj�2�5��Y�4*��;�-�	
�l�GU�J��9�.H���L�wgHT����h������'�ȕys�T�k[@���_+�p<�'��>\�|@��N˳��1��i�<����6\�$Z�m#*�ƍ�'lla�CFʱ���O� 1ӄ���� ��4��Xcfr����,�k�ֹ���L�LՁ���'5�ջ�uJ8a���D=/n�xVOG�1��Q��;��Ob!٧Bl|�h�D?�t�6F�g|5��A�~�',��S�<:���e�>$���h��*�ⱍL�!��y��%JѲ �q`	�<�H��ꗇ+�Bq�%�pɷ�T�A(~x&?���y၈[�4A\�aCB Exe���5Z �T
�̄?v��R��A�X&nx⇄K�T���bE^>����u����rM�Y��4˒�Sv��Ə�>Ү�+3#LCfX0v�'���A6��;���.g�8w��?$�|���)
�{�j�1q�����R�i�4i �)��و�K� C@��N��X1����6,"�e�o���cGN#��y�U\�69�R�Y&�d�3�����Mܴ��IF_?�&@���4��G�LB4��M�:���a��ҨOZ�1���#��%f��� u�hqb�R�k��9Ӑ�G9`�2���ǋ4c�<d��`��~���z���D��y`X�r��).p�4ytGF�~���C�O�\Q�K<����lH��/?�i�c��q'��(���2�������=3�X���'	�hk8�D�'��)��K;8V��ZOȢ-�Ҵ��O���ve�8<�L3K��Ӭ1x�-��&\	8���*�g���K�wљ��Y4&���	ד���b���l&l%���:B���Z 
 7��"��H1h�!�ȍE���vk
V3�����8F����	����E,���5��b�"kU|Yd���lq��Q��I�|�Z�i��V�9���ȡKY��T(2T'����.�
pa�=@���*R�4
�)��Ӭf����2U	���'Q�ܓ���Kd���<��!��j��O���@§iZ9��9��x�Nѳ�8�J6.�dut%�@�'�kщ�`�"���'�n\(�/Q�jftj'�ОuBn�Ð�֥��5�n���O��bNW�2����GH�~|h��X�2�����U0@��q2B��-�0>�ц�1znP�S�@�%�"2�x�h�K9%v^ipC̄�eb�E!��ש?��Qf�$sL\���]v'h��'��1�O9�M�E�>S�V]ڂ+�GV�:���ڽ�r���a� =&B���G�C��a{
i1�jLIL�����O�l�8|R2��7����DĨ<�pI�~��~�G�;L@*#����L��ݿ�pջ�T�r�phi�ބM���iL>���nV�1�	k�c�����O^�����b0��a95`az���w�X���ń����f�]�.[�0xK>�b�M����i�5h[XMz� Y*V���6��s����Q�`0��H��P�e�"�j�`ui�B˯0�@�$K//0$����#?V��F�2���Kj��:��i��h�PA�\��?a#�IۮS�dQ�&��`o�E�Vj%H^J��B䃖'&ȠEģW@�}�'��m"��q!�т�9w�TP��%�֦�Z�.��F*qO�>�@�ChB���i�t��8ч%�T��3�.T�z6!K���3=�bݦO�Ͽ��o;
�F4�dƃ)׈��DF���[�1�������/ԏJz���f��AI����I5"DA��k�&��@�'o]F��d���y2�H "�a��vR����!���y��J �����g�nq�S#Q��y�� d�Ā_&G��y�u�^:�y�n� ):�Y�R�)N�qY���y!p�J��6�@��d�����y2�;K����iC38
�@�B��y�`�^q \8�-ٗCǮ�J7b�y���8-��#A�C%j٢)����yb/!Fq���цaITt����:�y∐!����2�X���,�5�y�H�`Kr�O�WJ9I�(�yBָV��Ds�
5cප"�y2g��R�T,p��/�P�����y
� x�0���|,e3��3o��H1"OF���_�kd��J�Tb4�G"O���o�nά���ƒQh [�"ODuܱ{m�%�#�ԏ��iڄ"O��ȲHE���e�r�4Bk,lA"OD��A�/7vsH]Cf̈�`"O�y�"O��!p�Bq�Q�W8a;�"O^�Q�8,�`q�E%w:m�&"O(-r�΍�)S�{��ܗh� Z�"O�<#�NѠ� �〈���"O�q�ק��*&��򤁁�v���""O$$��dW+:�& kN�l�n�#"O�]�B�}S�J0k�xk>�0�"O(��S��8{n��"�	�eO,i�`"Ox����ZgL��F�]�@�@��"O���b����t�B56��yE"O�8��
�RvT��2�A/1�Tix!"O��AŇ�|���B�&+��\��"Obx��g�*v�JhȆ �36�40#�"O�8��԰z�N�b�/	F.�æ"O�<�H�F�F�Q�O�"F���X"O��	B"Z�~�N}HV��.~m���c"O��B�)eF����F�%={�HK'"O� �w(+^�}Y��]&nk�� �"Ov(��ɓ`�0��P�(q��#"O���]����V^4`��)H7*O�	0��S)~_ƕq O�:J�0:�'��рd�Nn&Ⱥ�Á,;S�'(P
3��'���q�=?�< ��'��ݳ򈛟!~����(�*����'<��b�
�N̬�R ��<o~Zyr�''�ҭP������.6�����'.�T#��R�i��#�a=|�[�'�l�jࢁ+����e*}!���
�'}J�CqkW,Q��m cI�r�J�z�'D�a��X�>��Y�h��n� ݸ	�'<J�xt��%kɚ��&�B4hfQ��'���"h�@�6�pf��)y(E��'�@���ĩ2��qH�#�"=��'%�T�WQ�ohZ��� #T���'��(���E�]g�WT=j�0�=D�DQ��K�W��A�/A�`���$>D�� �N,v>��/+pWZ�	<D�A&kP�>~1qD�Z4g:�U�.D�T����`��a��HZ>f&x��+D��	�l���te�?��9(D���p�	���!b�џ��<�#$'D�� Ԯ�KY��Z$�L�� `(��&D�8c�N�ј���Cj��&�)D����g6�l�B���U��%'D�9֫\	�t��a�āI	��WK#D�H�R��<F�[��Õ2�4�6�"D� �w�H�t������"��%���"D�l3�U�'��Á �p�\��a�"D�|�1����j�j*�V+��)��,D�h %-	k����88jax��'�Ov�	�&2��@�*^ *A>�st��LB�I����bH9z�>���oӑ@�:B�Ƀ*��kt`�( ��c`�?6��B�3H��%y�bB$N��YK��O!4�dB�I�'�]��� (&<DP�Q�M[�C�+s��_$�v��ԃʮ5��B�I(	��nۮfF�+��J$J��B�	7;,�{��L6Bb��eω1V����=�)� ���ei-5��P�֥`5��"O����6N*�(��Ë,CZe��"O��a��Z�~�����̜ 2�в"Oĩ��鍆v@���ƭQ�s0,��0�'�ў"~��H5ae�T(��Od3H�h�h��y�n�;���K��Wu����\��y��ӕ�L2vd��M�T����[�yB��z���p�H�.?I���vjˎ�yBd7oD�R�NNh��K��yB��C�r3!C]�M�z$P#P��'�z2慑R�Ÿ�G��O�v]����ў"~� b~�T��v�������t?� �ȓ=�Y#�(~l�YQ�I M"ڜ�ȓn��9�"�ǁU�������<�	��
���`�Ɗ`bb�@���.P1���ȓ` ���B�<J�kBH�wH=�ȓ��1rR�ɍ!��kt%{=��'Pў�|rF��8��s� �4�:ՌU�<�D�4k^M����z�����h�f�<Y�D,|�|�;�o�=`)z�u�W�<a�́3��=���7V=��oJ|�<it+)&�Ȕ� P��D��d�{�<ir�Of��� "W�Q�VdO:D�(ؠC7�rpo�)'��,I7D����]�?����+S�J8ƅ�y�ć��v1ٴIǲ?f�̺��C��y���,I��R�So`"A2B�ӭ�y2��'��`��>d��H!���yrN�}p.hrv��\������+�y�)H���ںY�,p1�O��y��-�T��e݌W�^m�c���y�탾Ub�u���$�D�h�O_�y��B�\�ug@UJZ ç��yr�Ɔ<9��K�i]�f6�Q�e�y�J�c8�hwn�}��a���
�y�#FTx�DU�q`&p;੓��y�莃5ub�bp��g%h��Wm���y�aD#_�`9�PnO TL��Jܤ{�B�I�(t
5t�D�J��h��.5u8�B�ɴh�J��uJ@�����▎j8B�I��|�`��H�F��br-Y9OLB� p�X5%-?���`3��B%4B�	�����׆̰B$L�cϸB䉮@~��q"X5wݜ���HH�K��B�	���kɕ!<�0แ`�X
zC�I= �ٙE
�U�,$�!��f	B��q�^� Y�P��C��/l��C�	�s����Ɔ�OزhM*X��C�	4c�Y٠m3@��=��.��`C䉋:�uZ5�EP����ʓ�`�bB�ɓa��R�@�f�)�Pɖ���hO>U��Ҝ1�܁c�Õ4�p� 7D�{�f�7/ĒQ�5�� �4��� *D�|��� �,d��P";L� ;D���B�S#����c{�� )7D����e�Ys,x���M�9���!D�T��*Ǡ( =�ӏ<{e��� D��Aj��}Ʈ �w葅 n@���?T������j��#��[P���Z�"OԀ�",��3��+��4��"O$t)�g[�vc��`䄅�d����"ON��$F�N�xH� ��6 Q*��'��,t�l*b�)S��%X׫W)LPC�	��@E�Ģ�#H���X�ꂅ.>C�)� .��W@��ȥ0r���vXZuq"O��1cE۶m�5�#�FJ�(�"O��:o]�
 jX�ah��k_��G"OZ��r���8	2�Z
���K�<�QNdc����%"��{7Āv�<�$�0eRЉ�eY�b��3d�H���x"�O4:��T��8#˾��bǖ�y�JL�"�11fZ�V<!#���y��M�t1�D��/L�}HzaId�-�y¬J6<�2�:l���X�@@;�y�/��.N���0�OX��E���'>az�˅fb<5j� 0h���C���y�'�'T�ڱj�,�(�*cL+�ybQ���A8�(�(r09c��yR�I�R�䂣���5b%H��yҀ�"6u&�i���"��T��9�y�F�)+	J$㶤� |�%K���y�;Xp~@"@M9x;�Q�v�X!�y�G+c��b"
��(�5iD�y�ݓG`��$)�6z�A��_��x"�'��Yb�I^����w��&{JT����	'<O����
̇-�p|2��ߐ�<)S"O��[��X	����EeP��}؇"Oe"S&�jHR�h�����Jp��(�S��0����˨?����BddC�I`�(��@愭px�t���R5+�bC䉝 b�hƂ8T���C>RC��5	YF��w�Ɣ ��eم�B+yp�B�	�@�&�R".M�1�^�:R�[�&��B�ɿ�����.��o���2�%�!��A�ȓ)z(��`o1P4�d�*]�䨆ȓ�|�����<(�աw
1Y�E�?iӓw����r�L="Oh�� "[!B�T ��B�2$��)�~4A(V�&���ȓ# (Œ���=yzUҵb��b}�ȓh&�����7`t���&;�⸆�[� �
�-Rv�A�,y����&����D��i��4�W�K=����ȓQ�=�"ɘ1O���b�LM&	Gb��f��8r� �=�,�Rɂ�yR���<����I�O"�8�'�B�v�,����!�KP�)�v�C7��Apg�S'!��'&04l`w(��.�Cg��R !��� �����F�
���
R�I1!��8b��U�A�B�y��P�h�?s�!򄘝ZB�����j��4΍q!��ܕ�d1�D�i��� �>��)ʧ0�B6m��E��X�J?qk"�S� _�d�!�d�m�uӹ��R����Q��)	k�O>����t�V��Q�D�<��}{�'�8yK���B^�Xa�ۈ-=`��'���Gy���L�O�8��4�H����7�1UP!��K�&���˦B&��Ja��cA!��O�Q.7��}��Dd��_?!�݊[�4�!`.dΎ)r��_-76!�� L�����N�܍�r��+p(!�$O�0�`�{tNQ�q����u�9e!!�E�r��{"��d���k��Ǿs!򤍦"!�\�"F+n�T�@@�i!�dG]����Q�b����O҄Y!�D� Sۦ�I�O��$!��F�!��/-�r���S�=y鷮���!��jj=��!��QH�q!�޵�����4$�����߉$U!�� "�#�@ۍj���cO�z^�2"O��I!c֤7vXas�nE+ƪ��"O��) ��"J25�
�^V)�"OdQ�c�>H_j�HAC��43
հt"O<���
u�ج����!<�ܫ�"O�<�3A��V��	�@�� 	t��"O�<�� ��鄍sB������p�"O½[a/N�3Z<*֔;�f��F"O~4��LV�)R�a���̙i��i��"O��%M��v��m�%D5"	�R"O��� K;X�$H�b,C���"O�xf�P�J�H�5+��8�ֹa"O(��M�#.�.4�����tE��q�"OX kv�1TJ94���"O���$��8rl�p&�9.؈A"O�dRs��P�N��'e�=TP�ʑ"O�Qh���P@ؒCo���f"OX���O�D�$���]�yb00#"O�Yrk@s�����dJ���"O*P�צ�:dͳ��@&6�h�"O����J�*ddL�Q�&S<��%"O�-BR�˃.�P��"��:$A
$"O�y{ E�a}F\����C�1�!�$�E.�LJ�b�,K"�S�!�D#mO��@��+/��P (��c�!�D��+�>(+P�,P(�}wy!�ک/�@��k�:H
��Г
?
!���M���f�Γ}�V�P7|�!�ը)��$����C���sdP �!�<r���rmB�(�[3��a�!�ÚTH��+R�x(
lZ�+�!�I�^�à�ļm���BB��7B�!�$J e}8�$#ְL<�q� j��!�d��0VL���0�^���v|!�.}�$�G��S�R!#��H�_Y!���7��q�#h 7%�����fB�^\!�$�![�aAd��(M��L�ո2|!��?J$x�A�"�)DC�|�U�ICw!�$ִj���� Ɵ&t����5�ծxv!��#"�h��	�t�H��FI2X�!�d@�L�)S�E@(o#�us���c�!���*(�6uh, �� <0�d�ȓ+fdY&(C�}�8�Z+���ȓ���%;%ΰH�S#E/R�х�Mx(�3�R!x�d�C�� 6ن�]E��Oիz�%�6y3�!�ȓ2�&xK�Xi/d�"��
r҈��ȓC�1;���'#i��k��?�8x�ȓ[�����ڐE�|��@Y�����ȓR�@A�0��L�P��J� -��͇�H@󍎍D�B �U:C2T�ȓ>����u�ڭ�.Ƿ='x��@��#���gv�0R��S�Ș�ȓg�5��V�,��xx���"�BQ��6�A�A ;@�D�L����ȓBO(B+�8	�$��f���Q��,�L�6$��\��c�@�h0q���|	��+t�8�S�M[����ȓj�0xb�������ax�3"O��f1�BU2so��}	���"O�!rk��:�h��� ���"O��P��U/A��3��9 �1�a"OJ���g�89N��Q��*�|�1s"O��1�C�#�j�Ap���`���"O� jLZ���{*`�i��M-�<q��"O�Ș�ި)?.|��˂4�F�3d"O�d���(D�t��q�u2�C�"OvP�+��sUTX���|1$R�"Ovu�7kW��Ă�i�%Į�"O��0�&���fn�2
�h!�"O�Qx��@Q
"[�,�x��"O��##�PL�1�A >�$Ta"Ot�hR�Ýd�Z��
�ujD �"Oj|�Rcӽ]�f!�t)^rg��C�"O(����$-F�SI�5L��U"O�%p�	R�S�H!��_�`B�i�"O��Q-��$�uʅȜ YF|0p"O�4y��S�&�Pqc7�Pk���"OY!�������!��&}��Xe"O<����:V�U9��E�@x�"O���'@24 �$~ey�7"OP���a��6�ܨ ��I0,_LQhA"O`Di�,B��R<��NHx���"O���P��m�Q�/rg�t��"O��3mP� 
:�!�MR�I6�"O `��ڣ�"���J�KCx�*0"O�,��N�@D����B>���R"O��g/��.&� �Alů0.�X�"OX�+�@��kϺ��'B'tp�I"O�����"���B�t�Ӄ"O�UiǇ�t���Ht�̞oz,`��"O���k��-i@���Yv$a��"O��D�c|���f՞jB���"O�@��6а r�n�.��L��"O�̢�k��u��P�'���A~иZ�"O�Z��=(>h!s�m�j8��"O}2����*$و�-�H��|�"O�ɒ����do��#�<~L��z&"O&�[t�+��q��2E��� "O��R�PgY�A��EE�:DZx�C"O�;��Պd��KWjɓ3!J�"O�L�a�G�>�a� i��@�e�"O�H�Unπ$
DmZ�!,�&�+"O�e�怞�-R�]�@�̅!�"O���A� )\���%F/&�x(p�"O��AA���� ��n�s�H��"O��J�	f	0ř���6^�QS�"O� )����V��E۴kQ�r��-�""O.騠I�����E�C%b��@�"O�M��c�e��Ѱgǃzq���'"O��H�FZ2@�����q:]�B"OnI!�c� -�a�e�N书"O��0u�P�l\v����^�Z��"OL�(r[�Qpt�K�[��l�"O��[1��)a娜�$F	*sHJ "O�:��EaO��3Q��62�"�J�"O��s�X�x����V�8$����%"O��j׀Q�k�N��b�S�.�����"O���@�#�����L�$�3D"OV(�_ҚM��g��H�~D�"Om*��A.OU�����{�0��"O,�X��H"y�U���	d�l4��"OSuLA2�$ܲw�Ǎ$��	9�"O dx�e^�K��0
�1Qo0��T"Oұ����V?"-;'Ŋ�j�I�"O�m35j^�8%by�u�S����:"O�E /YK�� "ċ-$����q"O��R�kW�$Zl4�Fb��^Ԅ	�S"O� �Tq��è�q���;�h��"O����E0�'[�u;"O(m��B�b*~h��^�DY0��"O֕I���a��u"��1zQx�"O	�3c� k�@ �W�;$���#"Of��󏚙_HX�s��T�6]D"O��Ѵ��*h��у
�d�*��f"O��1hZ��T]��g�'��{E"O� �-T,J,�3(�����"O"�E
L�t0Ty�G
-)�="�"O�pIu��G��yӧ�2�-*"Or 6�=ji
	j�$O
����"O�L8`���^9�W
r���"O��bG��T�(�xg#�U��T"O�� �I�	Ҝ�v�ҍ�. ��"O�}��J��Rd(��s�˪W�$hS'"O�����+)~�K�
F��!{"O�ɢ ���b%٣�'A����F"O\��l�2/�IS�m��n�X	�"OD|�&�	2T�);�mIX���"Oƕ	�� �Z�P�_OȀ�"O0|�
��
Fa�e�V�_"`�["O���F��R��W��{2���"O�t�Qʙ<1�)��o@e�a"O�;��'�j�У��T�]@P"O@(K�I��~��d�7;U ��R"OXy�-ҭ,��xǣ�%7��t"O�� �ͺDz��b��5/�K6"Oqc�eKo�u����6&5P"O���M��˲4C��:O4A�"O�AW�T>!�\��a	�Ȋ@I"O��d#�R�l['!ǔR�<�2�"On�����<nۦ�a�BF�{��A�"O YH� ��E�q�Gn��i�"O�S�-a�(�����~����u"O|xy��ݥ6-N��#W�!�ӳ"O�9���>9E��K����%�"	�S"O�����`\�թ�G�	;�tj�"O�cv��K~�T�ʡ��"O����A6L�&)ف@�1"�F���"O� 37�U�20U�U��i�6�
�"O����&Eƚ��+����ts�"O�P��N�h���hf$T�c�4J�"OBȀd��>8�������8N|�Y��"O*`���θZ��,	W�6��:�*O�"�o��h��<��0��'�����-��Rp�َ.����'����6��.<P�)Z�#�Z���
�'��p�mRF���M�/TG��	�'|�ZGn��l���{���V�z}��'F��t�R!_��`8�@�R�����'����(��Y!�ڐ���}�d���'��$�E��\x��E�s<Nd��'8x@Տ�7fq\�x�
���yR��"
G���!H�Oh�T�%�=�y�Q$2�>;$�N�?:lX��N���y��)ili��'`�T�i%���y�)7e5ؠ�-f�
�����y��\���oˬaR�u���y���`�u#e3\���R��qq�ȓ0��l�?=��Ұc%b�,�ȓx���qLk��Z�g��$u�t�ȓ+���JQ�Y5�J= ���75�%�ȓX(¹(2���D�ۖ���h����S�? nE+�%Q�6<��gɡ��a�"O�P�7��t��qƋ	v�j���"OvL� p��0�f�ݿ��g"O,H!�eN�A�>�s�!�^��m2c"O��@Y}|��E�1��de"O4�3�W'Ql�_��k7�
|!�ݔ0�XE�q�?l�p{��[+%m!��E�P�$�'d�����ڞW�!�ݍL/d�b@X���+6���!��߱k(r�hQ��0���v��.!��\"V)�؂�J�D�jE�4k�!�d^*]̀�����;2��L9v��-]�!�U����b��0%Ǩ�Ap�ۜm�!� ��)��� ���(ĥ �Kt!��;P�4���ď�H��W+=X!�T�	X*��G-W~!U@�3dg!�dE	�*���K�'�2���.H�>!�dڀS���؅֯n-\�Hs�?}!�$לj�� �^�u�ly�CQ�!���7UrĀ0�/{��ݹ�a
L�!�D�EU�1�������(�̴��'�n�&o]�	l��C��y	l���'}h8��)
�S��`�`�6!b:���'�4A������E�)	 w����'@~���Ų(�έz���z�`(�'�ʥ[�ҩ^@H
��L8>M�(S�'����������E�hL� x	�'�e�,�-Qґ�]\���'C�y�
N-!�lP��8$Qrq:�'�H��S�[|��%� /;��3�'b�\2��M48���X�)J5Y�ꭡ�'#$$[��X(�^$��j�5=:���'��31�§� H{�,�j28��'K�@�'�a���ѷh�tB���' `A�i�(���/�4@��x��'64L�ԫN 0?Eأ&�:8��y��'��
n
fa�g]�{'�A��'Ș��f�M��H���/!'�$��'�E7��)`�Nm�c��tp�r	�'S.|('`^6H���2c�M=z�.�P	�'�Q+�E��b��k�"ݓ HJ+
�'*���w���;��c���!&H|P�'��YQgM�*t��!�-F+ <��'��*��F��:#�:' �:�'
Xy�3���d�(��Դ
��(�'8�q�c�lj�-�_BR	:�'uҀZs�V-yW�PJe�@��v��'�D|0��ۤ�|��m���
�'�������2tf�����KR(	���2�'� @��뗺 �Z�H3a��
`�ȓD�"�&�<o��xh$�	*��a�`Y�A��={,�@�	;U0R��ȓA�,8���Տj#�0`*�<����ȓ����0K#����	�y�ȓ\1���_��Ře$��%}T���5Ѱ�(b�Z�H&��#�1F{��O�`) �5h�2�:���0ႉP�'����f
�[B౻"*�>JN�#�'�* e`z#������>Uڐ��"O(((V��,j�\�"���{�]k�"Ot�K`� 0�"�K$�Uj� }�"O��RC�=7�B�1D�<�ص��"O������=K�B@AV![,�j�"OR0!l�e���AO��	R� bV"O� ����LX)g���f40IjQ+3"O��ʢ(�9�\m��셾%����"Od�"�͸J�P���ˎ�{RzQ�6"O	�6�Rax��r*0HJ��"O,�±n��>͘�S�H�-3,���"O�(r$��,6C�H���'.�z�"Oj-c���u��q�#g)!��Hv"Of�t����y�C��)��[�"O��X �":���I�8-��\8G"O�E!eLUX�ŉ�N+���9�"O�T1u�w�.�U��>���"OJ`�H�j��iR�G� EB��*0"O���aPF� i�TG�H�A""O<�!�݋B�>�A�d$S8XX�"OdH�QA�p-�P'���5T��"O���PO��(�ra⟮]�਀"Ox��\$��pGK/��8��"O�x#�OU=:�l��ӥ8�^��#"O�%3�j��i��=y�
�(]�⩀�"O��`��_�Z���#�jˈU�f�1$"OB0��2:��̳8�0���"O���@E׋x���˃��:K�.��"OD�{'	�J���dh�-���3"O�����ه)�ف'�gs�)�"ON�s�-85���ЄH11��)�"O�����d�i�U���O�h��"O�r����h:3�k�_m �j�"O��бgB]ô�I^O�!X@"OJ�SP�X��r�cD��03ި�"O`��l��BÖA
f���(��"O~\�Q�܅b�Pr4�^>i Љ��"O�E��N�w���CH?��3�"O�p`�/(.�p ڏ	�,�x�"O.�Ӡt)�5x�;�h��"Oz�i'd-yt���׃W<.� �9�"O���R��#�$�#Vzs�0z�"O�t˧�ĎjA��'K�cn�0��"O��FU�b��p�L3�%i�"O��2�a��hʍ�k2V�z�#"OB�)ǋG%F��J �H�<��"OXU#a�Y���,_�;�Ny+e"O�p�UK�}y��%,�r�t3"OJ�5�
?x}�X�$�׃o���"O�\Q!�`�`���0$K�)�"O&`���i��Dz�)H��"O�ɷh�=Tֺ]:6�_"c����b"O��qs�ə]	$�p��?J��u�"O�
C��|P��G*A�t�9Ca"O��Sp�yؼ2S�V<ur�x"O5r��L7N�ҩ����V^	2"O�J�A�1ذ��R�T@<4��"Ob�#�$Q?*|���l]�A7���#"O&�R ܮ>{�ar�-	�v/���"OljǇS�h��Ƭʚa ��v"O���T��?7�t�2c��N�`�"O8��c�)�x}���=�ș��"O��ڞ/V@8�s	�5��%��"O��U�߿�R� 6��&H��@�q"O�)2��?~�g-�1��e1"O��x3��\n<��P���	�9�"O�h�O�6���B�ď�0 �<)�"O>�˗Cޢj������2À\0�"O�1u�8�^R�c�t�4M�"O��2�Co;@���^����S"O� �0�%�h\i�у^���X�"O"����4� �9e��$�H2 "O(y��lƼIe�p����f���"O����̉�zx�d���4wN�"O�:���77� Q&��1qX�a�"O+kR�MLBh
s L0W�Zy1�o�o�<�V�6  �E-���p�┉Ko�<Y1V({�#Dn�^���p�k�<1h�0e�~��P
�B��YӰ�]f�<ABЈqʦ�B�@U�"Ү���Sc�<Y�D��N��9��� "j�x��hv�<q4��7��l0d�\X[����nMx�<Q�쓢IR$Cu�ڕ�eps'K�<a  N�l�B<r�L�*��P�GTG�<Aƥ�"*���2�,��%/`���y�<��mJ��R͢�j�<Ĥ�t�<�7EC[�8�bW&��@��^l�<�����]�F�=@ʾȘ���i�<yF�6N�&9"�L��=ݴ̉�P�<q��Z���1����,�I��G�<q �ʕ���B�,1Ri��@��y�<q��>uΞC���#��-q�	]�<	VJJE܈x&�|V,h�a�R�<	��!b�`j�׋q�y�ì�K�<�������;%.E���(s��a�<Q�-� 7�%�p�� `�	nR]�<��oľ1�H1!	�1�<h���Q�<Q%�_�%~:�L
5N��Ń%JW�<���";�U���3�Fd��%�[�<��عa(��2 ̵A�8����LY�<1Q)@YvEkvH,[�VECpS�<TB�T6Hd��şu�)TK�<12Kى9�A t�~'Ve�1�C�<�Հ��Y�D�¯;��i�C�<	�a#6kL�X0� 	n����W!Z�<Q-��n���Fßd�2H��g�<Aӊӧ%�~Ty�	��.jdM�3�~�<�q-�<�\3��H�p3��UD�<A'�I�:�"o�=��I� ƊV�<i�#Qp��<��bW�Z��"��z�<���ɴ`��5��\yʠ*�m�<�q똢 �IŎ	DV,b"�@o�<i�ب,�r�� ��{�֨*���j�<��/Š|�P�AŞ ����*Sc�<��	��E����I',j���b��F�<ᇮ�H;TQS��\ (�&��P��H�<!W�~ �D��O�����0�^G�<���:J.�X�%K ?p4�FD�[�<�a��hR|A&�F=�x�[J�M�<i��Y�����e��GMp��!n�<y县8��qeͷ�����k�<q��$p12�qD
�'p�R�q���h�<�cK�S�.�j�I�G 6DQ�d�<1#!�7`H�#'F1eҲ��#�w�<���>-]`)0c�O)H�l��bZ�<IB"ͫ(����F�;{�X�H��C�I�v\9�I]�9� V�tB�dj��Q�B�pm��(�BV�N`C�I2:�Dbٯ7슈s�`.��B�4o�	P �<L�f��e�1vB�n��	fb���2([��Kt6�C�Ɂ= �z5��1	Z���)S�~C��7 ���2m�E��x��}�B�	�I���S���B�'e DB�)� J�i��%�u�%W	�Th�"O� ď�"tC�-���,HYp�"OL��ІΚYZ"���F�BA(�+�"OR���hJ�m�0��ɽ],���"O�A��6C&� ���� F�z�"O�l� ���-6ؼ��Ȟ-?���k#"Od�	�J��7Bai�'�<�|-BR"O:���S�|T`��ߏ�y�a"O�H���q8���\�zN�"O����.О��\�	X��B"O.U6.V�g���`�����F�ye"O:�A�K���Za�n�"g��C"Ob��V��l������FM�"O�k�gN#2Z���N�����"O��$#Ԝ�"�ޠ�ȱb"OX�W[�;����͈'3�r�"O>�����yp�[wLĈZo�Cf"O0"RJ�;^S�KP˘(,��	�"O
=@#�#1� ��RH����5�"Oz�"s�� 7���G�'gO�x��"O�	c����k�&d�r��/X���"O$�0�L^8~�(��Ŕ�F��Bp"O���6/�F���ȗC�I7�T�"O�t�����t��-	��"O�a��#\$"*���-C&�k�"O��êح&X��A��ϸ<�j
$*O����8�x0�H��������?���?���?a����O���G��0���.�;<0IR"O�X;��?yT�y�#�y�4l��"O��K�S=myc��(
�
d�E"O6D��O^��9��+N�3�p���"OQ(Eo� ��YKu*%Z��i+�"O��q����Tj ��M���"O�1�T��H�j��t�u�$Ш��'��'P��'���'��
4C��9#-|PD�+�F�pֈ5D�$P�bJ"��;iřOsv�Sa2D�T:�SL���f�C솘9�$0D�xA��9r��&kU�^�C2�:D�d��C/?F��ȃ,Јh�}�7M9D��Q��@ P0h�����=�W�9D�lK@S<j�s�h�{�|��Ӌ�O��O:�$�O��d�O��?i�!هX`v�jEȒn�*D���T�<)�I̾6������7�X���P�<i�	N��EK���}��q��M�<�E��d��H��%���,Ֆv�B䉶h|h�҆�n?���Q(tPB��/cP؄B1m�i��APid@B��&��(2F��U$�`h�@=vjB�Sv��fgx���'/Æt
$C�0C��)-R%>X�`d�@5O��B�I.�6�(m�w!�W+�`c�B�I�.�ʍ�A�s*�TyU"�x�C�	:���(��9[4���`J��vN&C����8�FfI=l���� L>C�	)m�R��f��V��QTAK�_rJB�	$bZ,����õ/t��#�;N�"B�Ie��0����{P:����p\6B�b�=#f�@DV�X$g�E\�B�ɨLk�x%�	oT�T��E�)YXB�	�2�v�����R6����(_�6B�I�@��H �#ڊ:m(��\�qA�K$D�0���7��t�C08�Lՠ�$�<i����HZҽ!��%q�f`Q�[TC�	(xl���R.��(�h�i���C�)�  \CQ� H�I�D�oо�$"O����FL�[�6����Ā �"O�3gM�i�� �7�	(�b�ۧ"O���@ �(u�j0�	'CҨ`�w"O24SOݫ8�n � �
.�
\c "Odʢ�N�r+zP����=��E��"OHMSmD�>�J|*��I�j���7"O�ɀ&ꑮ��k��N�]�xT"O��с^d�[�d>M�.L �"O,�W������a��&8�,��"O�<��$�bF<E!$DR<<��Sc"O(��#�tl�Bm���,p"O�%�k�'#-D�M�� '��"O��hThM�.B48	�No�@��"O0,2q*M�����W��r�����"O��o޽3���w&-p���+4"O �B '����	e�Ρ�*�{�"O���R� O�as&�?4��;�"Oh�4��^��aƃ�/a�"�� "O`<��T�t/�YqRbRf�h�a"O�����g��Ģ�3#��$�"OB@:�C�s>R�hv�2CYdq�!"O 0Cs,ټLj���$\<��3�"O��rʕ�k�E�	��7�Tj�"O8a��(xznx	g���D�b���"Oh�ԟHWh���Ǡ;��� t"O�v�<a*'�44���	�-g�!����B�ByC�H��!���$�f,��I�q�ƩV�گ_!�d��mn��B�eZb˴�PnI�e�!���Hz�{ק4�(���ÒP�!��)���S� �u���h3,%nn!�$B:(��/]�[�PQ�R@[�!򤗇@��h�V�(ĺ@p%��!�̆>����+C����	.!��K�W{�Tӄ��;6��M�5`	��!�Ă�D@����.<����ϑ�O�!��V�=r��d
�?/�%R��Ca!���1,�:� Z'e��8B Y�1�!�d��'���*9h������N�!�Dj���C��ic� À	�X�!��ܾ_&�C�/�S��HՍ�K!�۶��cg�C�>�@��_~	!�$_�y�(H :�nP9B��Q!�� +��۲矻T���U��`�!��.?����0$�	��I�!��1���WFF�c�v0�f��& �!򄖪}���3B�ɴm20���b .�!�$D�~�p��%).& ��׉�!�$�;u�T��υ84��v%�	;�!��8&8b"��#�9 o�� �8i����M�"�-�Hӓ�y�cS76��d��ǀK�dȋӮź�y�i i��HG�$�5��G2�y�ˁx��Q��YD�!'@�y���!J���sm�b�A� ���yBD� -�8a�f)R�^0��Ђ׍�y�)�4Z�ږ-�+*d��b�'���y2
�?�Z	+TC��T� �w@V�y"���~���LԸQ���A�/D8�yRcL*k�ꉳ�,�.U�b��oӆ�y��H'��]	�J�
�A"��%�yB�%r2&����1P2���2�P5�y�DӾb.�d�R���B��ҁ��-�y
� 4�*6��$���A&�>z��µ"O��g]u}�|��� yD�-H�"O$���	�pn���e%{6�a�a"Oz�Ί!>xR��%�;; ��W"OƵ:� @��҃I
18�!�"O��rb�C��(�Ȧc1�l8"O
 �PAQ<<�H�rD�}@ !q"O����?M�Hq�I�_^ b�"OR�x���k����C) ��""O�X84�J>,�������8`'"Ox���=�\�D$�X(v"O����������3A2M��	�"Oh�������׀�O��TX�"O�9yw��+,"���E���t�.��"Oz q�WQ�9 E+)�����"OJ�
�)W�T��aP���lyV *�"O��aE]=~�>݉R�H�	df�bF"O�Ȱ�����p	Y0@h�2"O�a��Bl#�h�"�Yr�"O����ʐ��DSԇ��|A��"O��R���f�vHKw�S��6�"O|yk��S�9��`儁

�^�X%"OfЫrf:N;�ABS��,��@�"O���B��Db�Dǫ0�X�pF"O�b�aB�l��!(�$�?o�dh"O��r�%?��a�`�we>�Sr"O~���+O!h�M��Ⱥ^~�p�0"OR���B[y�TC���9�~8Ip"ODP9�*E$!�@�F����i*P"O����Ě|
9� ��Y�"O��4�G1����iç��4�s"O�Z�!�X�$lJ���,K�(4"O���C!%V��C��E�lA�"O��ҋ_<��s��(�l��F"Or��u��\s���p%J?!s �As"Ol�����"���L�QY�i�e"Ol	�O�.H� �x�_ 4��
�"OBT"�� �>4�3��&�@��"OD�d�$�rX򎔢dD��"O�Q!��ӷ�&�h�_�i!҆"O�y��Z93�B��sC�(�u�"O�}:�a�-h�9����NЄ{#"Oީ�aLŌRktMbf�-\\��#"Oj��tȇ�@���J@� #Gtc�"O��󖬑�x�:�aӤ׎hpiR"O�)�d6;�b���O��$,�E"O��rK�}yb0�ßG�J��c"O����(��?g��փ�T���X�"Oڼᦅ�`�^ yG�A2����"O�H�,�����
�OI����["O��(�F��	�
���5v�,5�D"Ot0(ӇI܈D��_�P *B^����	�� P��bMdi�tc����B�ɒq��Љ�*<y	��AC�I������d�Z�y��I�$e�C�I*�Z��r�Lt"�!��W��B�	�&�9!P�-�4u�!�՞\��B�I�T�S�[,]��`���~B�	�l�8�P���>O�\�GJ�5N⟔��	!D8�]@UDT�T��(�Yu}�B�~���6�A�Tk���Ë�c-zB�	�uAPd�t`H�w�@, �%Y��C�I���2���Ke4hɐE
HPC�ɱ;��� h <aF�	�O��C�)� N((���+!h�;#�X�} �"OVy��2�����@̪�ʤ"O �s��X��@#VAٶ`�|p�'�+�/�d/­���0�i��'� �w[JR��ǀ.0���'F��:BkݤYd���$9OܤP
�'P��xr+�!CO��S�`�2Z\�	�'�,II�b̠�����ߕ0�~���'c��膱<[X-0��/=��k�'�|Hb�+$.��0$S�+����'�b	)�)A(H�� �@��>�[�'l0A�5h��} � Ђ�<��'i2ZAD�{��@��={Gb���'���R��F�~D��b�y����'��c1AU��򬪆�$y��M��'��| ��77$|9��jj:A��'T`��g��2Q����5���Zδ��'{��k� ��^P�R"�%V�y
�'�R<A��K8p�$���J_�*%���	�'\*����8���#��ڵ'w��)
�'��	+!�Ϭj�l����mF:���'X9��g�>]{Pm�7f�/1����'@�hQ��kP�%	W��*��#�'Lp�3f��S�̚3v� ��'� iТڰ(xm��^$�2l����6O����ZͰp��[ ��k"O*�#���~8�쓦��#> �qq�"O\�;wJ�=?�&�j�H!�~=y�"ORЁr,�*5QBlPv��-M�Z��"O���4�+;�j�y$I��8�D�@�*O*U{���Z�Rq��͆*b�(�S�'M�1�׊Ҽw��|��T�Z��=���:O�x:�N�'}Y��R��j��ТD"O�\b�A�����AK��@��"O��I #��X_��"A6�}��"O(�BM�Bvf�	ԀJ:r�hqv"O�I8�f�
G�`aX��g�@i�"O�	y��j��@,���9"�	�b�!���$�t賴��1:�M�c�І��Ot�=9�O$�	�M�&f�"i���ܚ�xX�|b�'nL�x&�_�v��ؔƒ&Hlb ��'{@�:���(>�P|PMU�9L(+	�'d������_^�5h$�J#hf�=`�'N�l�@�N.���r�޺�ؐ��'��H3c��wy��PS�]ӆ���'q�x�� ؛rAh�"c�ɀ[�� ;	�'�x֧�K =:E�`-�1��'�nX��[8���E�Ǯ_�J���'G2ݘ fE�PQ��e�F����'�* R0C݃U��y�3.˶'�����'?����4��w�D:�*ȯ]�B�S�4=jRl5��`�ǹl9�C�I%c��A�܆ s�
ˌIXj�$&�S�O����86�S���&%���C$/�'(a|b�R,2� 9���4 ��Q���yr ۥJ�쵃�F�2���Jf^��y�+ߜ3���d�YV0�0&�Ŝ�y]��(�X��/N)v���٘�y�a�65?��".ݩ}��A��yb�_"N�ʅ�	&u2���ǭK#�?I����8,��� 锂"hQ3�e�~���ȓl��(J【P>��ڦ�M8&�ń�,溉��I����dЩ=J����7��MzS�WS JL����z�����S�? ٖ�0ϐ��H�D�$X��"O��jRb�?,� h��BL}*A�C"OTI@�D�dŬݛA��?J�l�6��a��1�h�9��ɡq��!]V����	)D����Ť;�x�%��`P΀���1D�d����	���Ô�Hq����0D��q�Gǝ�f�3�͇:��A��,D���Ve�M
�]◫�f��I��/D��'��k�Bj%�N'�Y22D���rn.nb�}�GA�5���%�,�	t��D�Q�L�vI�X 1��uX2�6�$ �O�Q �ʷu��ԻC�A�Yi���"O�aCT/��)ZAA$�ŭCQ���"O`�C�6�8 Ӂ����QJ�"O�}�W��6Lp"@�F��9*���$"O~�f�q[j�#�@��XB�+�"O\la�✿u�؉�掻,
��!"O�u7��0�6}� f�/K����"O��GD�H�PIG���w�<]�"Of�p�/C+ujdd�4�^,�0��"OP��7�*+��c����"ײ�P"O�$!�B0ۦ�HP��Y�@"Ot��7��s�$��ܫ9K��y�"O�� ]�z{�y�C�",��
&"O4�5h�6����|���"O.x�l\�6Gj�dۖ_M���1"O>T��O�D����"j�LA�c"O�t��J�;i�"Y�� =TkvqH#"O�SEFY�5��Œ���6[	L�Ȅ"O�4a���WvU���]1L릐AD"O���4����T��w�[A�F���"Ox�b`Q�p<X���ʛ�r�r�(t"O� ��	2'_��┊g��M�"O�-�piȼ-�|0�"i�~��5 "O����~���A���6�F<s"O6P���)h�ppA�9
v�b�"O`A�-l�=�����|��"O�p+��;Z�l@su��<�a"O&� 3ͳ�}`' ��3 ��q"OTE���Z_���@`�@�0�"O�Q�1F� ��9q/�N�̩Q"O�[sA�Os�a ���0#��4A�"O����і=����P!G���	�"O�}c�-n�J:����U�"O"��T���FѼu�Z�"OTQA�ӿ@����s��;�) "Oʔٶ�	�u�Y���ŐU�֥�"O������`�@[-�-djN	��"O�7��L1���#�Y� "O>��E� M��1�To���@"OlF�*|��� ,{t:aS�"O �a6o��{�^�KW�I�j��9�"O2���`ʞQM|���b�n�(T"O�,J4�&4
�hPGᗹO�BE�&"O�	��mF>�6/Hd�0�Hf"Op�I2�I;{b�KdR�p�-["O
`�����OuH��ǜcj�a�"O��+�$L>I<<�	���kQ�P3�"O�w��r���Y�6�3͗u�=�������H6�l(���"h'I���,�0��؄��P�EDu�채ȓ5!�9�ϗ�v�X�O�e�|���T)��ᔏYkt�K�'Gm,�ȓ_�$�s�� �H\;'+�X~���S�? ���s�V�)�B��U��-��A"O1�4���D�d�pu��;c<� �"O�A
���%Fs�ݰ�]8e
�u#�"OСZS�
7�쩺R�O�0�Ȣ�"OF���n�o�8P����|�l�إ"O��yu���i��E��d5�f7D�<��AJo�`D��=F�8EJ5�3D�AvH���07+Ğc�����3D�05��"@���P`Er�9�.0D���S�y($ͼ�,X�S�/D��Y�N�
9�dpF.^�$���1D�X	�bI(j驕�!`$�"�;D��B��P�;z�J�(�yl�5��a:D�T8���?�����j�jP�-�"=D�\���)��v�d��眍{��B�	"zE� ��R�Et��f_0T�B�ZD�(��a��dg@��WMݳ77�B�7wt���n���2�i�PB�	?]f�+�M@�4���)7oo=B�Izx)�G-ݤ[��T�U-�.��C��L~�X�� ľ%��L�$	,c�tC�	:���"��%>�F���	N/N�C��v��0�"��<�8�GI:�B�1�P�hÇ؛T�b��A(H	M�B�ɚ��UrQG��|��W�#�l��	�'�H P��@s������L���'��C�E=5�0��`��([Pl,��'�����XW��y!�ܗY
�	
�'����(0������%�:%J	�'��DЩ1SUh�!|h�)	�'�z�y� ϕp�h�9�S�_H��'������r�)&bֱ�V��'���P��Hx�=��̆�1�� 1�'��eѡ(:U�Z�ʳ�	 1�T���'v6�x1h�B�@q:��!��	��'�\D�3��-LN��O�7vE�'�i1��H0y�\=1�`�#5��'��U���'B���:u��-Z�<��'_d��Í^6D^轙#	�5X�1�'qE��=�p�2�b5�1�
�'9�S�Ӝ�*��r�Տ`�X�P�'N�iB��r�$L	�jp���.D��G�
�0�*�9��ٻ�'/D� B�n��QI�����aw',D��ڲ.I�!v0G���UG��B��5D��r�/�Zs ��EE@�C�\堢 &D�����7�ޠ�7�9"]I�1�"D����-ׁ<���2�b$.�*���,D����Jښ���1��|�d�B��-D��K���Q�)p5��a>岗�7D�Ȓ�eĭ#�l|���v�8�˵	6D� �e�j>�Q*�%���V4D�,�EM�)7� �)�S��BE3D�@⣪�-)�F�;uL#t�(i�1D�Paq'�F�\����3C\���/D���7a&J�S&(��E�<d� *)D��0�d5�$�U�|�2�P`���)#!�D*�������&a�蹂���G�!�ą <�!UHW6i��˳��4�!�D�*n|(p�'�0�Ƶ�B,�}!�D�1'����s�Z�Υ���_*Ms!�V%c)�=1$����%�wL߽)n!��6O�܁ۢ�ݩ��`!bC�B�!�$�"A���ӁK1J��)!@� Q�!�� �H�&e�p��XB#����1�"O�F� vF|��P4"On��U:f^ܒ"k�� �tIa�"O�:p�bcļ(e�G�"0b��w"O��u��0G:���(�$;,= �"O�04�hD a�Q��Q��"O�u�@�R�^��t� "�r��x[�"OՓ3��=�:�%�W�Y~)��'t@I�W��'�4�ԢԿ"%<�*�'XrTPtO��Ȇ�!��'�\C�'�����a�M�!�PE�=��s�'�N��.L{�}�҂K������'e(K���!�0�*�ܲo���(�'c`�[��˪f�J�[�Î�jAZ$��'��p���Y�diPW$ɨv���y��&mdJ)3/[�]v��&�7�yR�Y5,����,�.i����d�y�lT�yȐ�A��D?g���ie.��y�	�!dd��P9J�r|K�����y�E��R��k�'6��4{t����y� Rl��$��� A~De�C�[:�y���y0�$;��P��� 3d&�y"GJ�Bi�1D��R �����y���C�`ıbbQ�S���g��y�� &7��XѠ��#"���P����y��|�X�֣��h��X9����y"I�~@ԉ �e�8�8��3�y�a@4]n��pc^u��I�Mȳ�y�h�=�ms�A�����۶�yn&+��s��}eJI��$D��y���
!��o�}M��8S,W
�yA�'	Kx���kŠrT��"�y�JǑ,%����К=LN�A�B��ybE+�M�pL�7���J� ��y��U���p��;Xy��yB]�����Æ��x̂��y�0)�Y��� �4DX3"6�yB���T"�F^<VY0ӎ���y"@�T���P����w 6bq͌��yr��dU�`����
h_���J/�y򆕱�j`�O8w{��HΞ��y"���.W�㱈��g��m�1�y�Ϝ*cl��u��,쮱a����y�I�&)���4%�X����
�0�y2�����`ga�O�ʨ15���y�o�(#O(=�T�MK��5�K��y�3��,B��
�D�e��l1�y�G��$������
�Q�F��a�yb��@�p�q�N��L���"l��ya��I��);���LoP� ��y�� K=�d��J��>�ع薚�y��͚@�d�iPlȹ"՜	�m��yĝ(բC0-�"�x!��@#�y�dI�H~p��$��"j$�7M_��yB�@=|�6��0$����3����y�N�+��@�
Ԕnb��P��'�y��_8�0��%K6h9Z,2��Ŵ�yB F~p �h�H�;aH���'�y2 �.��K��/ˬ�2�Ŏ�y�	(��I��$�Vn�JEU��yr`�4K|�|iĮ�`�XQ)B�־�y�'�h��\)J[Eh0@���ڪ�yb`��L����5�
�{1Z��y"���>�x����"@��� ���y
� �i���.�����
�qx
�(t"OL�C��[��K5B9wT�á"O���CV�
#�-�fA�E��y�C�j/
���-^�Cpx��E�#�y�)��k3��*��@_
X@e��y"jK� ����=(L�4�:�ynˢ	q"Pç:j.�A1���yrF��-�t��S�4(D��#�>�yB	cq ����|�5*SN��y��ϓlI�pc�mQ���x+b&H$�y"������
��m֐(��?�y�`��� �Ы/�,��6�܇�y"#p���B&-/�F�[�y�&_.��c%܃&�F�0�I�=�ybC<�p��AC_L�݈aF��yrK�qZ���F�L�G"�PB�;�y#��i�Xj�cC�=� ��)�y‛�?z���O�8�U�R쏀�y2ǀ�,�\�C抦.���2%�ɇ�O� Dzʟf��p*H^΅�!�I#3F��W"O��	�m�{�d�-66��2�7��֟"|�'bL��,)q{2��R��!t�)�'���شNZ-�8���������x�Q��MKA��P&u�5��,�yүG40!H���S4�>%����y�H�"aM��m*2$pU��b��y��	~�������#�`�Jt̍��>!�Of{�a�tۆ�s��82��O��	M��HO�y��d+a� @y�L8��Y`"O��A�εN�L1���[�>�;�"O\��C��j�,�T�@:�u(b"O� ���*|����Y�\# ���"O�	+G���2�X �\.y�q��"O�LS��,�l����8.�d"O1�,���j%ܸR"O����<b��V��l�-�&"O`��BP�9��(���\@���"O��b'�]!_Î����V���b�'���ͣ|�"��1희e��Q�	��!�T#V�.�1�G65��� Hε:���lGx=�(��S�H�AQ\ @����U�j!"O������.P���2l�>��ZQ�'`Q?�(Pb��@��բ"O��C �1k(�Il���O���OܬD���PY����'��#=E��,�|Pƭ�Wᑀk攔��OT��J֘�� �{�H<�v&�M=����M���x�a��]�|��̛�N��`��C��O���w��}�!y%�P��"OT��mR*p��5R�F6HG�p��|��Ƹ�Oq�jTA@��RR��*���*�ja��"O�-�C���	
ڣ^��$p��	[x�\@�!a�<ʱ�P�f��� D�̐���)-Q@�0�"[-y��Drv�:�D(�O&wO�6��d��̂�~��;�"OPM��/V�+,���M��$	���'��I6ɦ���]�B�~y��Q5��O���dJ=O�l���M"1���ٱ��O�!�$8n�H(4c�0��]�3� �M�!�d�9V㘔J��D��yJ��B0��ɪ(��D!�II~U�t�� M�-�40r�eS���B�5�D8����+xr�9��V�,e\DZ)ðb
���<�.O��<IL?&�F�Vo��9󠊀i��4�$D��j$	K,:�x���J�j_<���C����<I��O�p]�2�Y2C����E�!|0���� �Բ�$H~~��d@�9�Jиi����ȏ�`� �\<B*ꭩa"W
?�axb�I�fn�)&
CU�����d�[F�6�%�<8#"\�*d@���3���W3D�|iң�3��
��4Z���"�*&D�����<m�H��鎕���@U�"D�h�o�(�v�Uf9Wb�ɡ$*4D�����.?T,�w)�mLm�U�4D�\�D�;�dD[RM��i@R9��e0ғ�hO�� sW,�rǉ�uԅhv�:L��	Y؟4xT�M�b�11JY��rlsӴ�=%?�%�8� �#|C�\� �=6B�-X`0D�|�;Lcr-� $8hypŹD�.D���D��s��,z#e�)�d���-+D�X��	�*&��Af�/<6y�O;��t����g�*Ũ5��)]��@P�,�C�I�np�R�%�'M���ի�C�0��`؟�K����n� �M�&�1R�"�O�O�X�Q(�5f�����.
o"�ᣉ<4�	�-�0���S@�UH���g-����"��3����ŦƼe�rhy"K�7d��B�	!'���sTǘT$��	��F3 �,��%�S�O^셊���7k =��b�o'�`��"Oެ�r�Q1\��� �z�"S"O��s[�zf���2+z%�A"O^]�*�,2U�9pvV
I��{�"O�h�P$	d0�(q�  T�$�;��d=�IU�'��e8r��P�n��fnQfҬ[���E�h���P�ʖ6騍��ᘝQ�F(�#"ODH�p��0+��]���ЉF�|���"O�cP�>L�N�HVaKwI�3"O@XC��ߝo",(0W�����R"O2�:��_��m�`� 1-^R��"O�\1Ba��L~�ytDX����A�O]�|Hv�b���c��I
6qR�[�'0�}8��ҝC�=	U��B���'ފ#=E��TZK��vj�1+�p4'�8�yB6C6\�#%�+�� a �S��y���B��1(L�{	���B��HO`��d�:/V�����'�RI@�R<^w!��E�L
����J�3��\��L�vn�����ɍ@}��*O$w\ƕ�sÂu����8�Ĵ�(��J������D� L!��:D���Vb�Z���F'ʲZJ�-	%8}�l�0[�P�+_*vK�ՙ"���\�����Z�0��	&˔{��_�a�^�܃Q�X��d?�ɉ>a(8B�m�(K�X4T�G&	V���D������(p�n���F>S���p@6<O�"<�n�朋5�[� t4�Q0��g�<1�/?$�)�MϪVBP-�kX�)r��)��%*ޠ'��0���I�ps�5�O��	�`6��8)ȌaR�J��DN�,C�7EF�J�&�L`.����+^n�B�I�%�ʐ&��[�(��2�Ѩ%o�C�ɂK�(�X�C?D��ȋ%�K��dC䉿q��y���`�phK�C�	�*!��۱J��.Mz�oʧC�`���)��<�cɇ�G�\}xPH�f3�]����@�<a�G1"��{W��^��<��F@�<�,9[W ��nޱt��a�!��}�^��➸������8����tu�`�O����9���d�>(��
*����c'$�4h��f��X*����X�jhZe�6Of��>�(OJA���}�D�r��v Htqt"O� ��!�G�c� ���V��aW�	O�O^�xT)�R�8�	F7M�BE�{��'���x��$�E���>G�N��L�@����0{"�9�!�4�p<$ѰO�C�I�F~x
`H&��}bu&�0ךC�I�"|ܬ��	߿
KdͩR̍4tC�	7|��
&Վn��a�)ޏJ_jC�I	�¤(E�ŝhE�I"#�ڬ$"C�IfdȄPSd�=�:��Vn���C�I�B�F���O�T�2���kK�"U�B�	�P��ؒG.$MI�DO>AU^B䉀ZШ#	2ip*Y��
O]vB���´�r+�"~����o�7�jB�I9f�$���ɂ.\[Q(����M�B�	�3�f��Bn1�tIV"�!�4C䉖)ꜭ��GЧDMa��ߗphB�)�6H�FW�u�0\���6 �!�DE�/��Y�c��R��Ac���H�!�DG�Pޜ,$�ӟ~N�K�h]�j�!�䓘����q�YH���T.=y!�Ă��
��f��3�p��c��[�!򤃈@�q[�ę�$���4���"O舲�OݩR$���
]l����"O�uZ!��l2*̚��%
�6�ʰ"O��9��ۅ~��MA�")�¬�"OD�FJ�=#��a��8H�|%��"On@�0�;-l�Ի�m�#.����"O��P�K58U���F�4���"O��B��Ub�q�k �
`"O,��Ä�(5�J�дq|N���"O�	��U�` ��P71����1"O&1ϗ d�ԕ��#�)�:eq�"OnE��V��1�Mr�� "OڙFIX(a��؂3�q����"O`)��͍�2�R�R@���J�N8��"O�Aq�]�b�]�2g��k��1+�"O��w�ѬFI� x"��
S
�
�"O) �
\.2 A����`��"O���	�^7� `�D_%m���Xe"O���c/ؙtSd��ʓs��Ը�"OڕP����'4����(���ȃ"O90���*>t1�p�خH��|!%�'o����(@
{-|Y!�GL�6�茠��]D",�I�'��AE��z�2��"�)���
�'�0x�恚�N81�,ݐI\��
�'���G��Nn�l���T8	AT��	�'�,�P͢b���c�ؔ�`��'o�̺`��ت �ț{����'\v�P�Ń�W�	� AH�wh�ͺ�'�L��g�i#��7�âj�~�(�'�ɱ�׏`X4�W�b����'�l��u�/ub��p#	����'0I���YLW�ɧ�B��0�
�'���1b�¦_ݚ�t�ՃiV��`�']���mk6���/V�qD�uZ�'_�]�G烥{V�����rJ�C�'�
�HvNݧ"�8�TM�� ^|��'Zj�� ��n�-�t�қA�l�'3����;L
��"e�Vw�)�'�p�g)ߘz���k��N|�ŉ�'����O�|X��e@�	h���'�0y�ƭ�9z֭�t��]8&�#�'Hn@x��$�f]rT햎P����'�:5A6�ؼ�2�F	G,fE	���  ���*٤Z�	�P̑*�"O��aj��F��5�e=3�>�˂"O����+ܤ�0&_���I�P"Oz�����0z�I��N��^�I�"Of�bSC2W�FI��È����"OJ��e/��T�:=������d"Ol���D	`}H#`�-M�"Z�"OHP5%I�N�U���$u��p�"O���h��/��дő!T qٗ"OJ(� f�)	EuH�Fn�"ODH�T]�h�f�!��ư!��@�&"Ozܰ⃤4؜�E���= �"O�AGA��E�|=³Θ�U���a4"O \wE�mc���f����	��"Oh�q�O(�}{	�Y��Գ�"O��c"�WV�����֝v���"OZ<r�)�:l��x[G朚Bb�ͳq"O��a�� gD�	@�Ȼ(��ň"O�U0�+-e��H��	/��+�"O��S���:9̭x�A#s�u"O��Ц؈V���rc̙F�xt�%"O� S��W4@L��y �Όgxּ�p"O8Uf�D�X�0��Cm�`�"O P
pl�5!�9��L�U�!S�'�~PS��e0%�� Ϧ�(�)�'Z��A�Q|�<���+Oⲑ�
�'����wE� �;4R�Bml���'��X�Ũ�a�Y��KM�D�F�y�':��$d���´;�a11��X��'���w��M�^,�ta5��hC
�'��L���640�]�FP�-�n�X
�'BJ�����"��5A�mX��	�'�0����v���i�`H7zYd���'�wS?��HbKǥ~�B��
�'K�قqL�3�L2a�߇w���
�'v5��	�?"Jh�5Jn�Rq�
�'58�;����(-`E�c�LK
�'�����(��Z�E�-f��#�'/���$�]��8���U�X���'��p��(�~mR�A�
H||��'�^@S�j%F����e�	����(�'�@�s�
�1��� p����'j
���"Q�+̂I� ��4�R	�'���Ke/P�U����5��rt��'��	��JH�Խ"/E�nw�,;	�'�D
�c�^�,�A�X	�4pC
�'+& HU�1�0����MPb&��
�'A(1��o�f��E���=��P��<�B��@&,�)�<$l���Y;)z�]�'�*���'�ԣ%A\�gI(�ƀ��+��1R�O�5k!�1�����
�܈/�!!�����";b��P��=%>��ܔ!<��`O D�.ْ����3�hd�Q#\!!���f����pI��Y7�0���Z�l�ɇJV�ْ�Qܦ��v�Kc����p�>�Ot��j6����X $��ZZ���@�`q�7h��,����a)�eR�9�4A�g�NՉ��ٙ��Y8�e�J�ҧ���T�^�s���[�8
��\
�(Oεp�OQ�R�c��	G TQ4 PB��Z��j�[Z��A0�貗o���y�*X�}��(N�h�@cl���"e۴O��P�N�b>=��h4�6@�E��7e �@�8L� T3MN�e�@]��jV11��8#�V�p�)A
(�����1F��MFPP�l 0���� .���T>1�� ^�K�@}*d�0����L��|!
o6*�2�)�<Y�d�)���&!�6�����SΆ%���a�Xr�)�Ki�)��p
�jܷ5��MЅ��$Jg�$���/ʓ^��PZF*ݵ6��I��7nD4"�,�����Z4�X�WC�U}r)�N?.��!$���<� t����Ѡ��4���կJ2ޡ�ACx�"0m�_X����O0ԽЁ�F|�����6#��X�.��=&fY��[@H<��M]�^-�m�g	\5E:|���K}�.�=H��a+��Q�XX�&n׭�>͓L���8@��P���,+b	jb ��/4a~�d��1z���#$���i�
5�J�j7�o��;R�r��`�j������%�U�^�PJ���<�E{���D.j�:��C�MT�}"S��-$� �'��P(>E�'I6ti���y���NFI;���\=��@�!�?����$�0�Џ5}��4��l�Y�SEƭ7䘐z�(I|�d���VT�<��]�����̘3��=a'��oyr�2g�pҗtX��9��	G �0�͂�Wp�VF!�Or�6�@�z����	�h�����0I>�S��ؐx��N<h�jM�� ��F���J�͛��O4ԩW��k1�?*�!�V�$��ҥ���ix�g<D��9�k�Yͼi�$o�9*V �E����z��%x��]�H<E��bȧf9&�b�נ�
Hx.K0�yR(_R��Ez�?u��A�����'�ԼC �Z����運r�y�&��@ߒ�P �(���T�֑d��t�E�P�x�*�K���/$"~5qFO�9xQ�Ag4���4ț~3fpk��	�9���g��a̧2 B�QSΔNb���R���x�8���F�?Q��CH��GHt��5��%�B.G�:ҧh�"��td�W+Bx�ÏI$0��(: �'�� * h�LFp]b4�͊%�U8D�\�w��0j�!�e?!���k�ҩC�g���I4-�͉�,(��� L^"=iҢA�����䡟��5� ��5\�Ȕ F=2��(ɫ�n�%m�/3$�~b�L
��9�O��C�<����'��� L�@�:a4�c�i"l �yӖA�:�Ͽ�1&���B%�6A�k��!�gcPM�<ida�KS�f�0;Jތh��E�F"ܛDe*a��	�s$��Z���(�^)�VN gJ���矴1mN"m�`Ƞ�W?I T8�Bb7�O hA(�[�Zd��`�H9q�ĂT��#�@�x
Б�c��B0E*�:g8��� ��ў8�Ѣ3fDV����ɝ�T��=ʓZ���!"�0`NX���4;/�:+_8B:L�sv�Ƞ���+ʍb�r}��%0b��lʻ��>���E�yPɣ�N��9��B�&\kT�iP��?,� %�s�i|V���+��9��$cu L	�7���ܰi��0Y �
#F�J@R�yB��02͜�`�HIl�C�EL�DE���ȍ �����>c_�TQT4���P������<gX��}ޙ��/�$��AT�V��8(-�OXiB�!7a��
�L���(@@(SN�3Sg��ɜ�Rpa���BHiU!E?4yP��ly�YD{ªҤ{�� i���C�D+���HOX@ɒ<d`�<�l!�9ա�P�:�c��ߓ��b�6�D�⎓@�!A!ʯ�ē ��;b�"�s�̑���`,RsF��FUj��I9��P�b��<ad%�<p�޹�0m��e&@<C$�����;�vyI��;lz�Pv��FI�7-Y.-���� �O�Xr�AU'����	�i���
��fX�1���~���F�,Q���'~�49[F�'���ݴ?�|]�&�W�0��7�<C䉓N���&-��!��)�b���b�
-��<o�jL+��0-�8mH"#�O�0;`���y'�
B#���;]A��6�0�p>a��ڡ\��(9!�х���a
��Fi��� ��T���-���'B���C�2_?H%���I�{3�8�v`ŢDd�RMZ�H�Z"=��"�<p`��ѣ0�\��N?ə��!C��<�����@�煜�1Rd�K���Yp�!�V����̝d_҅�ׁ.:%h(l�
5���L;r�0 �u�D��Sv��E@B����oZ�ft��5��%P����'�-؆�ԛ-����
�J�R챟h��%ϤU>zX��f�p�VZ���I_ Bh�Ζ���jE�×P��U�	�Kc�~b�R�;X|�2u�4�ܽ�ä����a��N�W��u�@�:?N�ILsܔ*�-:�3?!�#[�Ț wg�8"�I�T�'�nY�2KBX�2W`�bc	�KZ�IaM_e��d9#Ŗ-3����d�[��a{2aR<C���ʒ����^%��M1��J5L��=��F���J�5�L3V"7�C�p����-.C�tZ�ɖ9M�!�䃺r�hE�F�ʹ]
ܜS$��/�t���$���^"���@��JҢ������ZЩG���'޿I�5y�u�ǧY$U�$��L�)A�%�'?�c����.�JԎCb��A%ѻL0����n��A�2�(�O�q����q1��sC��C
f��M)B
F�(Iʍ�'�Z,�.�W7�M�'z�M:q�y̧=����&ɋ';�ek�.��R9%/J�d��c��0>��A2N�d��ף	T�����)��$�B(`���S	:��.;�PPe��K#���S�? 0��q��č۱�ҲZ��u�P�'M��C5X�`���Z�Q�xJ�ŕujy�E�VI}b�iY����#l��ٖ'8���*�;����J=p!�P֭�36��ITB
;��O�S��E3k҈���O��#���6���a���" �RN-9F�I3LM_����*_x��~�'|Z �N�:�A���I%���s�O:�y�M�JE>]�M�"}2E�9>¢	*���H��cb�S��l�#Na}�Ɨ�e�x0D�K�a��p����l�9�.��îh����'������ 4��J�z��4���|�����$P�D�k���.^7e�)Z9�L�'�uڔ
^�z���XU��.&�)�'�`�񁆀XnR�����+"���'t5���G0&솿;��A
�'�0���H���y�4�6rR]�	�'�t
C@I|!�9KW茶"�(��':P!���^v�f'S�.�ԕ!�'�xr!ȏ0NW��z��:kjf�
�'��y� �;V�V�HU�D	d����
�'��5:�ϐ��4�؅F�7Pt���'}^���^5.�ք�u�K�DD�	�'��J#�4<fF@��o�4�S	�'�>PɂG�$#�Le���ިb�z@`	�'� ��TD�
t�#�=]MŒ�'�&��CIɁ	� !ܖ:BZ,��'�ԉ�&,Y+�EJ��QҦ?D��R+ӟ<i����f<$�d'(D�Ĳ� �	p�9`6������2D� ��I�p��L��G��U��m1D� �g�J�z..xI�E4�r�1D�,��ë,�|`���ZֽCS 1D�̊5���^�,9��$������S�,D���LZ��D-k��>5W
�kǩ,D�@��&	B4#�[5"E�O+D�ĠuΈ%(T^ٲ%��u0N=���+D��q�!�����!��:qH�B�(D� y�AȱsL�4�֏D3���o\I�<�RjC�@7P@��{̸�e�[o�<!�b��*���M��8�"��lD]�<1�N�o�����O>p�v1�"eSU�<�%^Vz"lP�*Sb9��Ȗ�]P�<��,A��ӂЄw ���+�M�<q'C�n�&PBd�;�h8PQf�<Y�cO��DиW��T��g�WZ�<�%Gd�ft!��J0�RQ#�H�W�<I7a��6�B�ɬG��rt��S�<��"(W(�ta�k�pM���D�B�<1�k�#�I ��1�6(�7D�<)��ت=�1�2Āf�����jNB�<і�+a��yH��klbU��<�Ӌ\�^�~4[�j
F��D��oB{�<qT�Y�&������z^رBg-�z�<���0) X��q�E�j4�WQ{�<i����S�ڸ#։��D`|����\�<!��ѳz�xE�p���4�� JD�X�<9��ԜR��L+gĔ��T)����R�<�SO�ibSj�$GÐ��N�<�����i�R�D�oE>�#T��
SM�KP�Ez&
)f� �;��"D� Jc�;*p�An-
kX$A�� D�$��)�-Lf���/7����F?D��i�EU�n|Р��g��U��)D����*ų�0-i4�W�A�F�#Ӫ$D�L���~�2q��ُ8q(`�"D��sG[7`K�M��B&*����"D�lQ�#��o����T:l���҇�/D�� �t10�����+�oבA�T��"O����͋
X�Qa"n�	:%��a"O�py��ȟ7i��B�]���x�"O�A�`���ab����,�Ӓ=S"Oyc�Z{h���ɐ?�DAA�"OQ�E�W�O^2�A�)��D�.�q"O&YPWBN	\�@@bp�ק�z�V"O����q֚�P�:k����"O�u�E�SVzl�k���ax�"O.qZVmG�=�pT�vB���`[�"O�x��N,.��'��x j"OPA1��@i����Z7-��A�5"O�u�r�M�_�X���D��%�"O�̫�f�E��%�sB'z��9 "O^����ت�� ��#.͠"OJe�boő`m��^�x�z���"O�bî�:}�TX㠅O�U�����"O,��S�Ӻ}nF�{q*�P����"Of!A .�R�R ��
X: }� "O������9[Z^4U��4@�L��s"O&�!���19J58 ��nIڈ�#"O����Jm��Aɲ.�9B:��&"O��͙ؒzC�L���u;��v"OԴh`�
N$�|�vAL�d6�	�3"O�\R�Ê6K%ȔB�KA3'�!)�"O)邎G3P�	4I�782��"O��b����e!'H�0	Z��0"O�PBb�7����T"�91�@��f"O�Dp ��@E��p"��j��Sa"O� ���fpYQ��:.�[�"O�H��`h�t-�C����"O,yA�Y�2��j��8�PY�a"O��q6�۳B�̹ *p���"O�E���$x��)Da�@�"O�����$a!���C�3g!�a3�"O��"�J�^KdU�!d��$�*�	�"O�� P	:�J��B�ٻz�*ܲ@"Oҭ�U�K[�~e���Lc�ظx�"Od A�`w��	)�J��"O�0 Ǚ�:��1�5AZ��S�"O���� �?&�����
��0�"O�=k2�[p�.�Ȅ�O��E"O����èn)�=J�9B�a�r"O0Qx@�QX�`�veIre�4�3"O�8�DÍ���)��bY�� "O� ��g��GۄT�&��Z V%z5"Oʜrf�])��1�Ec�H�
E"OXm��� E�`��BD�r�ۢ"O���C h0� ;���#6� 5"Ol� �M�%���+3O&l�́"O��P$�Z[��듦U,�6��"OrXKW��=���(�[��6��!�'�Ա˳�[I�S�O���J#Z�{',�����|g�hBA"O@M���YTBpB�㎼ ���@DY�ȲR"S;s��퉑��)�1��*_Nx��a��Y{�������=%>��1.�Z|�9�@�$��5�4*6�DP3�Ɠ|!��Йn�B�#ʢ:�I��8ck�IU���(�����Q�d�j��>�O�5ұ��/���@�&nÖH�
�5��cR�
�i�v���!���H�c�ND|V��z���9\p(����@ҧ��2Īitm�Ӆ�wl��@J>�(O���KE� ax}���i��6x�W�˃Cn���ۘ!����=!W �˟'G��y�H�g�>������`���� �L���Ci�Z�]N�b>�AeG=������&;��Á�M8��a��犮B�̍��C{��hR��S?����.�����kε�Y~�1A����qr�S�H7 �RŔ��� ����6g|��M��^wt�:@�'�p���j2b'����ʜ�a����~j��A��3������xR4���Q�"~�	7WkR`*ƠF��
��#�>n���<�)5RaF@��D��uW���� 	NU�q��]NԵ�'�p�*�ez�b
������%�k�d
��� ����WL�l[�]���V�q;�)������+a�$x�EQ�'��Z�7��ݓ�b�XH<!ah	9w3AÃk��C�s}b�,
t���{��� 4����آH���S96��D(0�ݻU��Q����F#Ru��X5��f78��-֘3č�ROβJJ�xv���K�l��P�\���)�'y	�1b�����G=f�p�y���	�G�9b�l�<��Otz�y&�S�fԖH�CL�.%Q*���O�%��'إ_H���ğ):bS�b�3@QbY�3���w����00 �Sd�e��i]�B�H9�o��Lu��I�!���1��ڈ�y2W=c�α���ț~�P:�B���\9S��NaX���	!�j{ꗬE�~I` ���{�����%y��ʀƿ�� ��Șѡ��ETM����'���&��m���KM�i���bs�/&��:Q�Mk�'2�D
�۵n���"��Ij;�M�ȓ~�*�h��$W��
��18o"���'"X(�4�)�'F��yh��"Y|��.D(���ȓN�8�9����^Z�Ԏ�&k] �ȓ�&�@���JtZ�zv��#d*�0�ȓ���±$<��LB҈� &$9�ȓz02��A�]�2@��#|�%�ȓ7nD}�N/2�q3d�õk�|Ԅȓf�Ԕ� ��*0��v,�-l�
X�ȓMx���Sfi���*��pż���ɡqǸ�ʤǚ�%��ҍ��o��!�F@"r��ȓu�̰�s�PjT���.��)PqGz��ۻqc���áLh�'Y���*`�"; �qTN�*�($��h!Z�kW� �y ,��/�'0]J��E�u� ���ǀ3.��)���z��`��ܳ�T�0p�o!D����*�'cc��i捬M^�H$���;�̙5epER��bX��p��.���h�\[Q6�0�1�OhQ�0BY�@>���ҽ9��{�"g��]hG�5�(C�	�.�a����� Ӧ>���<�󬏞!�$"GT���O: ��7�\�|jPKD�G�" T]A
�'N`��RGI;hvD��G�	�œ�DV9.�$�C�Ɔ9~@�S��?�.Q�,��@ŏ�!ba��d�H�<�7!���5�I�]�px�%�E?���̬DD�Ī/��<�&zX�qR�i��IKR8���]e8�(Y�,�+t���@pƍ�R7����,�$g��#P��`���ē�\bd�
�t*:M`� �7u2MDz�)Bj$%'Ez���*�v��V�tI"��ɀ�0���B`�qOv�}�|�|Г1.�1 �4�vI>0!�U�I=���Sy�)�'zu���e	��y��!n���u��4�$�xa��p>q$�˲%[��B5�']x\�P"Εs��閉ן>��c�<O�����=���Λ�6�#�"O����QLĮ����)u�!�����; ��|�X����ШDe҄d�t��╈(��-��"O4���յB�[�+0��� "«VDA�D ?�Q�:�gy���6���EI:K�I���:�y2$�'^zĠծ�+zT�Ѩ`C�i���9W�X ��0lOD,y��ĒN	`d�Ta�E�^A��'[.IHF�P��U��DҦ!���i�(���>[QL�K�9D�XB��Pg&0��!�b�0�9�	j6B(�Yl��`4�'n[r�@�LT��柵:U�=�ȓy�Z��	밽���,!uʧIĎ6G4�x�^��C�4�g~�� �>,���M�h�� �p�G-��x@� g��A�C�b>��)� �6�BV�r3��q�C�^؞	竝�~�<�X���b �#K�,��ÿ	���@\!N� �4
��](�FǭL���;�!�Q������Q ���{d��
j�5W4zIx'�� ���j�f��0��Jб�Q�,ҧ<@-&�](
2BmQL�k�ƠG��Xu�&� ��� RHiVNN�V�DIp�F�)S��·ʄa��B5h�>�"����ɦArT�0�Ǔ&'�"�꓃�����<�:Ѵ	�Y�ӧ(�P@#�S?Y�2U+`oЖ{�2�3�HZ�3h&��Ŭ�7����	[�b��Ҥ-8:m`w�T!0��'s�\�0�*Hnʧ'�d��IC:;� 0��'ل\I��7�, �kP�4���	�@7�5�2@RA�	���K�d���"�P5P2�I��>yde����B�i̢v��>y
�&�=a�9'�B&&��#�1�4>�5�h	�L�����[��>IKס�]�V1�A!M���I��r��#�g~��x����B
%{� �c�����Y<�K���$��)ҧ9����W�E�Vm0}aTE#2"H�CiI�{�^\z��'��J�)�,Y���ئgu�Ⱉ>��M]0N���3����}�͔o�t��E�I*@�U�X���?	�MTn��%8�dOPМ�Db�>g�0������x��F,K:��!fݤ@�^�*�"�y2jҋ��<�VC��h��=�`
��y��ؘ�`��Gn�ԡ� dZ!�y�,��.W[�c\��" Z���y���u�$�s�K�,r�θ��H���y��w�,Tb�ϣ0�\����y�H!]���K�4��	[�X��y�F�c.(�h�,�"=������y��8�������5�1���ҵ�yL�<NҼ8�F��Z[�$1un��yR�Mڠ��@_�:�:@ O�y�ҍB ����Tvl�p�A� �y��^b��i8��װA�����9�yүL�Y�Y�6����%*�$��y��ҎK:du(���(�L������y��D�Y,��h�OB')�����ͩ�y� /r�>��@�%Z�`����y�C�3]L���n؊%p�Ԋ�*ð�y"dS�6:�)��$A�8JZ�����=�Z�zd�"/H��t-��(�(��@RQ�M�!R��@U,�\��T�H��pK��@W�-f�I�ȓz˚h#���f�F0�����n��Y�ȓ2F�8���r��0��˪x�(�ȓ5?�A�F��'��$��dX��ȓLB�� ĄM1��A�e����ȓH��Tp�j]�Ud�2��\W:ͅȓ�����%H��c�{fB���P=lۤ�Z5aɤ�k��C?i�ɇ�>G�Ѱ�	)�HC�@�Gw�Շȓd]R��s��(x��Rj'0q����?X<H�1o[�tWM�/`�2e�ȓY+��(7
T�.p4d�`��<%lՆ�yB�p��\�=F���ێDJ���ȓ;?
-`��	�c�~�*��=����� fX 넃
�j4����6h����:d�����H�pOj���C�6U=V1��I)���Qe��8����2N޴Ie� ;��U�L��������-��I�D+��ܺC���	E/.9��F�y���B�D�D��X���C���	�(��ɱ$�I��i�
:"��+3%ܴemL���HO?���h��4$!��8 ���P�T;�HOa�4�R�H����
d(<���
�?�O^EEzZw�>I��	�.)�9�#��E%b�1���z���B�c~r2O
���S�W�:�k�뎋{r�K&$�G�� �'6�d�����~n:��4Jf�	�v��2@* �c�j��<�,O���k}��I=���H�����K��T�5��	
�Z7�!�)ҧ��M`2ٞP�v��Ј81��qn�(<�uk��v�#Љ�$=|(9���d�<A7-H0o�d⣯����2S��U�<���X/�B�Ä�e��$�O]�'�@��	P���!�Ak	'%�ni�R.��lX!�� �Ih㩈�Jf��;n�*k�X0"O�x(F��3��!�׍"�t	��	W����3	
T�0�_\
�@��ȟx^���1��z�HQ��X�Ov�)k��*�<���G�q�*�[ٴe�b�Y5Ї2��ҧȟ�D⇅;�����ʟC�$��B�~YhԹN>}�C%�������@h#�+�L�B���OF��'���(?�'`Ֆ�KeO�
�,����f�vq[$�x�d�9��7MѰȨ�P7-�*��}����/��(�P�ʕ,R��5�2�dYJU�`�FU�M�"}�0�	�EX�a䠋32\BA،2�S��'�<k0�U�T�Ʉ��=J�%ɷaD1r`��4$D�X6ث�|D+�!V�HB@�u� �0�I�L�+{-J���)[3nu8"Oht�D�̰}���!SF	��"O�ݨ7�ډ�� �)ϕf�v��"O�1S4'�k<�d(�>b�Z�a�"O�(K��ĕ.��a�A65*�"O �*�@&eᜩ�잧FnXxc"O�1�6*�K$�@B��N�'@�d�1"Ot��CiZ�`�2c���a��"O�mZ�"�}�>�R�mkۊk6"Oܤ����5`t���W%�t�"O�k.UA��%7'��3%@�ѕ"On�XC/F:?�Lm�G��
6����"O|����q6�X��Pjș�!"OB%[v&��{��@�3��0�qx�"O$eZ�)��T�����]a0��"O䘻p�R�	�Q�
O������"O�bQ�,&8���J�vY�Q"Olh�Ο�: "��'^�u���pq"O2����M���#'�
}��Z�'K&( W/Ӆt�(+&�+��a�'�N)E�#Z���+��'�Hl��'�,`�C�*%hD�ݳ �^�'��[�!U9E7�1#��4�d�0�'�IhW���T�J����>Z$��'���فCJ�U?~`��Vy��Z�'�F��/�7r��jE�v���2�'{��QV�B�H�*'��C� 	�'|lh��
H�����F������'�(�A*q�|���K�&���'-���R�j
�6f�6@@ �s�'G�����
�Dy	íئ`��<a	�'ה�r"���i;3�ݑh[���	�'GE���;� 4�W(Ɖ_3���'�~�R��2|�p�Z�C��'	��
�'1 @�I�-ĕ��!X:�Z��
�'�ȩ�͌VR�q�%�]��Iz
�'~����ҮA�N�p�kO�m�ʓw�v1`B_+��������D2�a����~��\Ru�<�8,��"����=b|�͂vJ�#K��y��L��#��D�|�j��B}�����(|i���t�\%ڂIҞ0�D���v@L���	U1X�9q�Ɩ��a�ȓqt2���FH�R���I���!���ȓ=~���g)1>�0�b�K�i��9�ȓ:�t���W���pX���w�L���\I�)�c��"�5P!� �U�0U��H��e1Q%V"�d]���H�b��ȓL���Suk��r;S�Ɇ#�D�ȓj��8F����T���F��Y��Nj��`g �H�����pॄȓ(h��*$!�F���'.�0�ȓ���3k	�k�a��g ��ȓ@c|�Y4	�H�V�1kC��P ��S�? h*.աx�-K���Z�򭡔"O�9Aӥʆr)
�b���<^�XH��*O�@{U!�<a,\t���� x�� �'�hl"m��3Uj�b#�Nh���'������O*@\1cF�@�n��'��d�t�Y%e��d '��2�l��
�'p���`��{�d���[�(P�Y�'V�p���Ʊ��*pV�4y�'F�yH�Y�@��!�N
p(��
�'F|8�l)%)\� �N8W�|)�
�'P�����:s��b�ΟP�:�Z
�'�,�@��Ր�+c\O�t�	�'��|� \�t����"�YP�l@	�'ʌ����%�`�M<2��'��}{��-x���ǌ^<}�~�
�'�&�ƃEDP3�XLRz\h
�';�eӗ���z����ׂ�u/�	�'�b���&r���9��0t�b��'(JYy$N�0=�:�[f!�l��P�	�'���2`UF`�5�A�d���@�'B2��� �f	�d��fh�'nr(1����p��8�-�����'f,|��U)��a��S�zy����'���P��ߝ?�	�$R�HQn���'WV%�u��}�2A��ݬ@_�(��'����Շ���J`@�	l\��'�%�VhN�>��'�8x����	�'���j�H�)�H�lփi��b�' L���	�C�ѻW�N�\X �Z�'>����F�=�~�Q�E�O!b���'�"�+���5b\R��q@ L�R\p�'�8��g�P!+�l=��럀@J0��
�'�N�!֮Il���.,a�Jm
�'��yӲ��xT����m��+gaJ	�'�Lj�ڥb�ȼ2�� %�!��'����ّn� �v�'�&��'<�t��-	/D~�F�ˣz��s
�'Q|`���M�;� �Y���#�l�:�'yr��e��2�����L��*�'����j˃}S��+�+޼��a�
�' ���G�Ȳ K	hK�
�'Bz��1❑ o¡��Б_�����'%�e!����;��l�� Q�W$<-��'�Xx�"`��1��\�׌#��mY�'�R�ڷg�6?X��F'�W����'%�X�IO�l*�iH&����Z�A�'�\����Mjp��GG|.-K�'>����銓]A��hҖ	u�P�'��I�4E�� <Hb@ ?4����'Y�0����g3D�#5 @()k�Q��'�j��)GG̈�A�=%E|:�'�mQ,�F3�Kc&��q,��
�'Op��D <lȹ��4�,K�'��x��L�:w�z��^�;}t��'rD;T�^Bl��s�B6o>��
�'oF<�Q�z4����$hJ3	�'��d�Tl�	V8��ڢ �	}��C�'	,9JqiŅ6����ҫ5����'��T��DY.�,�B��a��'�<���@/"h@x��	���S	�'#<L	���t_~41�!�,0�3�'��-��7�hT�573�����'����̸�nH#%.��+��,��'u�3A��1#��tY���+6欠��� :���e+w�n�T,�(hc�e2d"O�:�*�Xn��VJ�yYL��"Ox�(��?xT���H���"O�}BN5n�
!��B�V��u��"O$�b��M7rn0`[�FL
�fQ��"O�L{�p�Uj�s����`"Od`���Z� �5GD�>?y��"O�0�7�\�aг�ޝ4��<YG"OX����Y;<�ش����/r\���"O��r�
�^L�A�!ˉ�|n<U�%"O|R���!�l�*��dt��"OxY�S��##iɘA�2Jd"tR�"OhuK#��7�LL�5N�4��\��"O� QqT�
�-�D'��^�q�"O�q
�f�[2��0qOY�@;����"O��c"ʿ*�6�RF�޺Vx��"O�aPD�+R���3@F�]�ŁF"O�hp�G�#,H�R�/��9m���t"O�qҁ�K�8]XOr!&!�d�
=0�H�%K�~����gK&!�dB�gZ$��̜5T�L������A!�d
WW���'P$e��)�#�;�!�$\ (�=�qD@�.���)aG��x�!�DC�z#�f�i�r�Ն�%�!�ŸO�@��-]2o����#�P*�!�Zy��;��<�^���H7Ae!򄀭�\TSg�/B�҄9F'ݐNO!򄔎r�f��G
B<
u5:-�:�!������a �8���#kץ�!�D˚~U ̲����PⷊB*�!�$ұ[i ;a���G�����㆗e�!��
6`�����b~�A�A(B�!�V��%��I�<�YB�留^�!�D��z�� ��\�K@jK�l�;_�!�DF�6I�WE�b-�t�gˈ&*�!�Z�2�B�ۃ'��"�(2���PyB S�T�v�c�	O���l[�Ř�y�h��5�h}ض�/w�:%!���y�M��<Ĩ���J.!*e���R�y��]�犼�V+��}1��s   �y�����r���o��YAP��0�y�P�\����1fu�X�D슏�y�O��X1p��q�����ͣ�yrI�.* �9`���
j9�ຂ'���y�f�k�ڡ;#,5b�X�bAC��y���4��m�T��ZB�pq�^��y"EO�Tq&	�� �>T:� �L^��y�DR,T�cr���=O��V�G�yR�n�2���D�GL*�1����y�!� q�n�8@�ΓF�l3Q*T��y2A�[~v��*�t�0p*�����yB��HNf|�c��i��Q���6�yB(�r^��v��]�=ÔMP'�y�D��~�~���FO�(i̠�cL�y�̶Tv��o��T@M�C�J��y�l��+�P��Q/
��J������y�NA�G���B��Q�����r���y⤊h 
���D�t��V�L^d��FWF���B$mV��Śo�N-�ȓfi���(Υ%� =0v@�
��q�ȓ;\ �yÉ8U��ٳfY�����I��"�@ۮm9vD��w!�c�<ɗ+�>T1�&@B�z� ��b�<g5N����)Z~v�ҡ�Te�<� Z9i¨�>z��i]7�P��`"O�t�p�D�2Wa�5� ^�RL2"O�t��u��1������,��"O���B>ft��Qiƃ�D�� "O���BOo� Z�͎1�ɒW"O�Y##��fV��`�B7؆�B"O��RdN
(���É_��A��"OJ�+�A�X�y�3�؞v�|��"O:8)�䇽h�H�3�I۰��%"O��Y2LM}2qB�.B�� ���"O�m��&�	LJZ� �3w�m0�"O��dW`0��ʬBd*�F"O<�0�蓋l�p��'�Q"-_
t�e"O(��Q���8�LO[s��p�"O�,K)M�a��*���"��h�"Ov�0    ��   N    �  f  +  �6  DB  �M  W  #a  �j  �s  i  ��  �  u�  Ν  �  Q�  ��  Զ  �  j�  ��  ��  3�  ��  ��  �  T�  �  �  j  f D �# A, X4 ; GA �G �H  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h%���븧�O@��1�AE�8�QP��Z�	$��
�'q��&װ-��J�gI�H�'|�仳n޽�j�R���*[�����Z6����C�k\���T�[H~�B��D]HV��
	����2�W;���'�^���d,�'HW�ePU�K�D��!&I�� <��6���$�8x
�Q{�/gY���=��^�б3�)�+("�F/W�4}����ys���Lס8����R�%:������?��.ߥR������'/�F����j�l�L<�@��=l�{�nM%VZ�����i?���S�^
p�Ė='�:���l� C�I�HX���4������ݽ}z�C�I5n(]r�'oϋ%P:ӣ���?��Ob�"~���/Xr(+��ˀ*tv�	s�E��y��]Te(���aE1#ǒH��f)A���F��4�$�͌]a2u�0��@���q��"|OHc������Ţ�\�?� ��>�	�v��yh�5��dY�eݽf&:P*�Aޚ�Px���3:� \I
�<I�y6C.9�֑���>�4�*lO�0�±�
������ڨ����c~�>q-OT�	�F��pa��G�z�qf"O|	�t@1����v�K%H�J���"O�كh��<������47u�HY��',h�O�i���B$;��hu�Qzj�(�p"OheБ������ �_rW�	��HO��/od���
b~t�`��~�B������*� 5�d�h�!�(ǶB�3L���a5���Q��?�RC�IM�R��&l�����G�g�I���?	r䐃]Lx q"̖�G�flpc�C�<���+��XuF�/�}����}�<��){ji��eH�T�H��R��zX������ ���J��ZVvE�$���m���Q"Oظ�AQ�W�4!Z��۶7^*8��x��)��!WI�8�Ȏ< �����)J;JW�C�I9~@ h�)N�̖��臰T$����q��G�y��N H)�ݨ��ב5�b���+\܍8�X�`�J��0l`2�D|2�S/����gN^+z1jE��>�C�	'Gp)��@������;W7nB��+O��Qp�L�*�m�)�~�BB�Iz7�l�E��BMx�{����<6m�����'��\�Aބx�8����ؕ2��H����$�<!aA`}j@�'"m� 2�U�<�4�C>y� �R��ČF�ȅ�ULT�u���O�����@�V�:a���?�X�
�'�` �,�.��ujw��0s�Ԛ�'�V���*�^��s��Ŧ,N-+	�'g.%�$S6*i���Ԥ��]<h�'-�$��WC���R*7Όq��O©B�ɖ�U3�C)G"t!��"O���Tc��t�:���Pέ�s�"Ox�r��f���&���\��8k���u���'C�ؔA��V���RBoشo=�Dn�R������OS9� A ��C.����1�8�<	���O޵C�
n沉ar-8�Ȅ)@"O�iS��#df���Fꂑ$��{��'��	-26pQ5%Jl&��%��ZD�<lO��<��h'��J��[8<�����9D�<���J>{y�R��5�μ�p6D��c∝e�tLڇFK�F��@�.D��S��xj���`"	�{�̹7G9D�d��G�6]��uL�. Xr����5D��s�c�d
D r��z�(P��.D��ؗi�7$��m�� ��0��|3S'2D�TyϘ47���8��B�&����*��j���'U��(!l0&]X4�2c����5�}�%��$W�ژ#��7K����)����`h�3�6M3��<aj����8D�C' ��f�t���C�sQj��/�ON�[
�1�5��
Հ��to-QML=��>De��)4@��"%ȫ|Zͅ�b�:��r�HvD0k��1� �=����D�8&$���i�e꬐���>�y�
�=����`��I����W�R�y��І���Z#FB+X������6�y�n�	h����P�:T�r�/y�����A8�x$Kk �1��P#Ԇ4�����$@-Jy!�#�G&�z����<$�0�T�sYx��C�Y���'�ў�|����#v�ᙑ'j�C�k؞��y��Ω�,�BT2t�my���y��Pb! ���#�<U�!P���'�ў�O�x`��Ku�˦�ϟ�ex�'Q�i�@�M�E6��Q�A�	�4�'V��QDJ;���94L�#9Oʰ��ј']j�3BNߨj�x�G�#��`�'���jP+�-gN��jP�X����cӮ�}bn̊#2�m�ǅT ����Zr�<�a/O(1�ޡR�'�Xy��	V
ָ��D{TO?��ݙ3y��$MN�!�d�C[?S�!�$G�y��qFb��0P��0�F�*����>��M�6
�P�ꒁ�.j���W�Nr�<1����03��ǡVQ.  ��q�<��B�Heb}2����2����To�<Y��+Q����`6XF��F@�n�'��y
� ��!ыe�he�1GC+9m�t�`O��j��0Q���F C�
Q���ج��T8����I�'9�p��e� ����+4�Ot�"�'��l�`�[����s��s�|j��HO$��-�3N\��2���P%"OޘR�CKe�lm��FW����c5O|�=E�t���\#6����/�n�`�N���y�M�fs���7j�:zl�������џȅF�:�(��4gE6��3ED�	���$�<ѧ��1$FH�xd$VNΠ5��a�p�<��A�O�H�2	 �(=��2�kQ�<�1ˁ�r��y�vʽYR6!p5a�M�<����C�\��J�9 L�8sd@��D{��ɗR%�I�e�=V\��O]� r�C䉲#J�Q��G�x�Ԋ��.B����	�7;����~��hOj���L�?}�4���`��K*���'�2 ߳
4b�얏�lՋ!�Y26HoP������� )|!@E�Z��v���
 �0=u�?�(N�Q�Q.�o��ݪ��E�V�,��p?q�F!���{G۸��ؖ�]cX�,�O���E�M�a@j�a�	#\���R"O� ӿ�Z�00��H0ֵԐ|��'��O^b�(#�l܁2P�*s�R�\��ǩ4D�4Y��y���h�Ι&a��0D�|Sf�94�,%��`��w,.D���K�o;�0����> ��b �'�I\kQ��Os`����4$��M_'>&N�P	�'Wf�# S	���8����*�NE�v�:��h��_�#�����n_�AF��0SE;*!����7� =� D�"	�H1R���A�'�a�iZ�UBج��S�Q�� 8���y"��zh��Fo�J�d��@�y���Ql�X�P�4��͂��Y��y�ܩ"Pɩ"�J�5Cd�#��+�y�
�����2��=Wk����:�y�@o��:pH�H���$ �<�yl�aEX�9�o�2H�\\rtB��yrGOWG$�(CfR�sܐ�6�ϋ�y�gJ7.����F�q�Q ��ߘ�yƔ�P��<�1�A=�`MYe)F��yBV0D��t��(�:/�e�"P>�yr�C�[
|�p���#$�4Qd\��y"bϵ>,�]�aW����#0���y��K%Y_l���,O� GNL�B�M��y�8c5:5��	�#�!(g�R��y�^�6�Y &�ӱw*1&		6�y�j��o=�����i���y�F
H7^D���*E�PѱaO�yr��*8�(S`���^8*qL��y�CE�UI����Р�p$�y��D��Cr��4n/�`�Q��y�I�1A~�"��s�p-3`�6�yB**t�yIB8o�q�'nâ�y�9�fȢr@�oa @ʖ�yB��8^Jd�1L�,�rk��ybF�l�8�)+ ��Aqf���yr�?p���1��p1�J��yRĈ%�!�i��"�.
DM)�y⣋��e2 ��	&R��b�A5�y��I5hb@l��ٗ#*�[��R��y�FD"?���-�<���H��y©�Li���-����/��y����e�E�S�U�)Kp�QBY��ybG��N<�PN�n�t���(X��y
� L�����S��z�ŠdrR���"OJ��4���C��5�i�j�5�$"OD��P%�pD�P�b-�蘥 /D�pQA�OY���JN�77�����@?D����Cͯev���R~ְ���O���O��D�O����O��$�O(�$�O�m��c�7G�M�!��x �5��O��d�O��D�O*���O���O���OF%��F�1�j�8ԫ�5jjP�f*�O�d�O��D�OH���Of���O����O�p�!L!8(ĉOH����O����O�d�O�4�?����?y���?AF��^���'FQ"Yf܍��D���?���?����?����?���?���?i�� �FI�tJA� H�!�'Ď�?i���?1��?��?i���?Q���?�"��`�I�1g@0��hdC��?���?����?����?Y��?����?�S��P��|��gZ�?#����_�?���?9��?��?���?��?i�ȗ2�l3���p��[X}�	ڟH��ן���ԟ�����x�I˟|���=O`C���`��Y��K*�~�	��	Ο���۟���؟��Iܟ���; P�,��J"dr����J�'g���	ݟ�����������ßh�������`���r@#U}�N����5< ���	��D������ڟ�����I�2� ���_�K5�82�͓<#y��ݟ��I����I�����۟�8�4�?���Z��Ճ��2/ ��c�	�(��^�8��Oy���O��n�%@aL]�F�C)9�0�0���k8`��$�4?yu�i��O�9O����*?�����s���wMP;���$�O���c�����������O�|"3ꛑEd�!u�Y�k�j�q�yb�'��h�O�:�/���!5Z�E�G�ںB��6��%!�1O�?u����C�E��~}ԋҌ�.\�����?���yBP�b>�,7mx��!ua^�(���`�S�������k�d�2�k���$�'z��(�8^~D�`k�)!�L��'���m�ɬ�M3#B�G̓9�b0�� ��FQ��X�)�7����2��>����?�'���9Nq�(2	�~a��F�^����?� ��X"V��|� �OT�;�g5�x�s
��(�Vi�tJ��'�{.O���?E��'���@�$p���IXtd1c�'7x7��E|����M���Or4;���I��4�rc_�i�N�
�'_"�'"�l�&#�������'R�����F΂�ʢ-��	�LX'.X�*l�$�H���Ϙ'��$�q��8�� �1��n=�(��O|�l�H2���	�h��`�'j2��S��6!�`��ED�k2U�Xشn
��(!��)ϘA���R��EҀh`�A2c��t%��)j
˓��{�M�O��aN>Y+O�-Ȥ��I5��`ٻɸ��'�R7� Q���D��M��ɹu�)9����N�p��d�ĦQ�?Q'W���	Ӧ!X�4DAt�SgZ�\����@#��,�d0ӖbM��M��O���,�������w�l���xo��J����Q�'���b�iJ�R��4s j���D-��'$�cn�`	���?���4��7":!�p��v!��4�0*ikK>��?�'4��`�D~Zw�\�&�ˇvC�ȶć��Mpf�E�k���.��<���+�[>2�������p���O��oڷell���ß��	\��GW:�ԘjS��ek���Ŝ'���U@}��'?�|ʟ�xA!o�s���� ņFSL�j�n�#����'/�	���|��b���$�X�`�?@7�m�#�D��i%ß\�I�p�I֟b>Ք',H6�X�Y�%`ʈ& 撼��%��%j����$����y�	�����OV�SFO�x�j�I6O�P=�y����O����J6Mr�����f��Y��~Γ˦�����vxx�g�2G�̓����O����OV�$�ON��|����?"�����kT��'_�[�v
4{"�'\r��4�'�06=�<� R��f�L��k�R &�����O���H�i>��	�?%�s��ئ�͓��<r��V�k5 )�AI�DEϓ&]̅0v��O�HL>.O�S'�D��6x�Lx���\$���dԦ���柰�	埰J����n��Ć`�9S4�Kk��+��	�	F�I�b0�y"@���(�un��e �0+� �ҳ�M{љ��@�d?��A��!�4
I�pG\+�-��N8���?����?���h� ��݁=�]c$�VI�>TK�!� 	��V�=�2�7?�c�i��O�Ε�7�V����H,7�� R"�>tS�d�O����OB0GCת7v�I�"Jh��ޟ޸;1�4p�h��ϭs#.�jB�-�$�<�|�<�"�^XS�eHq�̀5 d8�G�I~2!lӊŋ�a�O��$�OP�?)��c�_�R��_(
�XQɆ	ִ��d���ش+؉��O�d�wM�J�3�p�;�,MJ)���<᠀Ʃhh��IF��ty��:8��7�M4��0�&'?���'z��'6�O1�Ʉ�M�3F��?)����;����9FD�s�X�?)��i��O���'�2�'�26�[>�x��>?Pk�,�Z������G��I/X^ ��3�O�q���� d!�@���qʜ'�ּ q7O����$'���Kߧf�Ru�fmg�4�d�O����Ʀ�6H7�i��'�����
�PR��)`� t�\��!�$�⦡x��|�A��!r��'����A��1� ��oؐr�~���r-�I�Y��'�I���	�`�	�t+��h'�\��vxP 	_^|v���ɟ��'�7��:�J���O*��|���Z�!��R��K^�� hc~2��<��M[R�|����!O
�Q0����]�TrLyTO���0z7�Ou~���'��/ޟ����|R��9h�"$a6�� F�^�RG��l�R�'��'Y��\��[�4*>@���&�tt��0�{�.l!��ߟ�?I��C"�6���Py�i�x8"���_�v�`Eb,L�w�\�lZ�8�YoZ�<1��D.l�Z��矊��'C�a�g��4#��+�)�&I���'���f����U[�
�>u�:E��6��M�uE���?i���?ُ��	v��.��b�1�JG�h�ԣ'	�.2�$�Or�O1��EqP�K���䁮I���1�	�^�ܴ���'\*�T� <��'��'�	���ɶ�d�����<P�!�7�K�* ��֟�����ܔ'a&6�����D�O�$�<il��B��&{w� r
Rs l�$��O����O��O��Uc۷+��̉2(6;'��`%����scP�Y~NT���?�Yx���O&\i���������$�l�`u�0��O����O��O��}���<����s�ע3y� ��۪�,M��!�vn�� ~b�'�67)�i����*E�"L����<Rb��,�IƦ!!ش�}�"b~�� =O��L�S��p<x�	�	K��EY���0U�Y#��'���fy�O�R�'�b�'���ԯ�:`R�ʂs�h ���.I��/�M`Ă��?q��?qL~z�tL����(:��v�U�P(���R���	Ο��H<�|"�*�d)�㙹^1R9q�!J�k��d`2��}~҄C�p�!�I{d�'�剋Ea�ݠp�đ`�$t�cg?��������	���i>��'�l6�ȃxZ�D�%Y$*h��$��`W`�Q�I�0�����?�]�����M�I� � @'.Փ��U���7'����ݴ���[�"�hh��'��O&7&��<-2���  2Q1�T<�y��''R�'���'1"��>9Z CQI�2�t "����$�O�����E�&1���i �'�4�z�K�C\��jT�S) ��91�|R�'��'$:��ֻi"���O*i � �j<
Q$�[�5u ��q4p����EB��O���|���?���l���NĎ�0l�Ă]�`��?	+O �n�nh���	ٟh��o���ƁH ,�Ì�)*!rP�c"�3���J}}b�'���!�?=�SoQ�)��H��,��c� h�Wh�;�9@�+ˢJ�|��| (�O��XL>I��L'H���E4i=�q��� �?����?��?�|j.O&�l�lKԩ ��	5}$�q@vmӬ ��YRUa]ʟX����M��r�<Y�4t��58с��8��ơ�j:�M{�i�,�e�i(�	�tx}Ѐ�O3�'}M��X���!q"ȉ0e���T�4�� ~�H���yDК��I�P ��!��+e
�)��f�޶�赀�O�8�4�M��Q��XY�Z �3ↈDg�� R^�%�D+ �,48�dJ'hE��^�@�8�ɍy�l�3�	* �2�P��n��p�|�s$6Dr�M4��H�fK��%{Z��! E�7K�C@m��d�,�i�oTw��kQe�Z�4���L�P�α�5fY�In�
u��_�ܑ�tj@_�5+�g�F�DaXO�D����0K��N>����Q�P��5���@�s�F���OH�d���|�'�� Yjz\�ț�^�����ZD����4E����B���O��J'"�0y�記ǏM6^�PC��X�U�	ܟ��	�O��<�O�ʓ�?a�'� �Si�2�Q�vΒH���ܴ���`Pq���D�'("�'I�蚣�\%QxM�.�V��\�"Kq��$K9\R�'��	��($���#�
��VIװSxV�!�E+p]"�:Jr��K>����?A���� $i!5)U?<j\��T�y���SbHV}S���	X�I���ɴ\��nG	�=���#�>;�����#8���T����'s^�{��g>- ��W�E8�@ТV 5l��(�Ed�t��?yJ>����?��$���~B�D/Z�\@�`��Q���ó۞����O���O�ʓO�HsZ?��	/?�8�B�Y*�|)c���a�U�ش�?QL>���?� ��'�������,�
P�(�~b�۴�?A�����c�.�O��'��E�'�^�p�Fc�P#�A���`O����Ox)i��1��}�GGQ(�fPzb��n�|Y���Ȧ-�'�VH*��kӜ���Od�d��|է5�BP	F|���H5H��1�'���M#��?���V)��'Rq��,�D�O���GG�d'.��i%�`�b�����O�����L�'��	+j�쭪͎/m���,��y�F�!�4W��Ԉ���I�O U �[�z�!Xc�\@�Y1D�E�������I�ɪ���O���?9�'�%2֢S�]�25�3��;U>�A�ݴ��<�F��V����'FR�'����:0�}a�A:��Ov�p�d +�01�'�����&�֘�*c�� �)2���b؁$���J�$�I>���?	����dݷK~����nF�P�Iy�+�.�v���'�n}�\����d�	ԟ��I�S�m�uo�d��KV�Z�V)1�iF���������Ĕ'��R%�d>� �=hCD�[@m�C�+F���uP���	����	ny"�'R��c��Ⱥkw���LЙ�^{���gr���?a��?�+O���K�Ӝp`��9'^�pqZ����l�*�Aܴ�?�������O|���R�d��/��9|xa ��*��s���M[��?9+O��b�AH�S���s�a��Ĕ�{��ճ!�^��4� �qӘʓ�?���m�>�������O����$�p@�D���2�'i%VX:��i�	)I>�1ٴ��ß��Ӣ���/?�ƴjw)�
$d���U�����'��ș�2���j��}!E���u��c�&�b��eq�9B �O���O��D⟲�S�4ED�B�������-X�H˓k�l+�6�ɣ[�
�A���Sʟ {�@O7Hꚩ�sMP����áMJ�M{���?	�<M)��x�O9r�'� ��� MgU�B�-QN�;�������Ol��D:F���Of�Ɵh��3>U@�@[�T�ʝ{R�P+S�vl�(��/yy ~Z�⩂�9D���d�Xt� �,Qb
�uP4Y[dh�f~b�'�r�'.�	�3�v�ʧDJ4oP���R�N��3�KG�ē�?9���?�.O(���O�=����;0��a*�l8$���4C�-,�d���<���?a,OT���a2�S��\�2�ۣ>w��I�`ɐi
H7��O���&�������8~l~��"iz�T|0��	*ʰ�2�"J'kGR��R�T����\�I}yB)�#]N\�Jk�f :g(��,�(q�E��ɦ��Iß�'���'���k��'��'^u����O!D�BY(�LN��l����	hy��::>������klH� �@���4k
6�Xt+��=�P�\��⟈#�GB˟d$?�s�e�%��(4���Ҝ]�=Ç�o�&ʓ>�H�"w�i���'�?��'��	�W��=����X-"���&��6�O4�D�O��$_�s����M�'�\�8��u*��=��yQ'-�٦Š���M��?����R��x��5�%U=+��$P�D-e�4H�ڝ�MӇ���?���?����B(���.+�(Ⱥ&��-:��Z0�J�1�J��ڴ�?����?I�	HP�����'��"�h,J6$�;4歡���O�`6��O����O.yŎL��O�$�O��h�ᛁx3���Ɉ<yx�h�����q�	�"��O<ͧ�?a����ěeWN���Ƅ#
2�6�>Y���o���[�A͟��'���'eBZ��1�"\�F���M�83�|٠��	�`~��qL<����?�����d�O��$�,5&�@� .S�2��fb� Ry	�E�Oj��?�����O4��2�?����U�f� �#�8+����Hvӈʓ��'���'xxB�I��M�壀�i�F�1V+ϛV\8�čQ}"�'E��'o��8.�hEbK|" �=	>���o\�IO�dQ�lU�����'X�',剭R���Ip��t������h�+C��<g�f�'��	ٟ� 0,Fz�T�'s���5��)&m��J$m®M�z��R凶���?����(��2Kh�S�td�w��y�,�o�B1 G��M;*O�K��ʦ�������z��'{�E"G�ÂC����A���4��I�57��Eu��a�T�O�i(E���� ���w!D����iO~Qi��p�$���Ov���� �'��'*5��+��80��CLM��ȭ:ݴb�X�͓�?A��?1��$�'�� ա�L3�x��E�5I�mp��tӞ�d�O��$('�"��'3�	���R]v���*j�p�`��<"Xn�̟l����Z��d��?9��?�Q�[Utp	��
`��"∐  �v�'�  �Ԯ�>I(O��Ŀ<A���tC�~+�\+c�S+u��'��B}b"1�y�'��'=��'�剂~�����B�ywL� D9uLl0P���D�<i����d�O����O��p oІ8`�p䜾n<��m?0��$�O����O��$�O�Z�p�?���Q�Z6D����J,5)|�	�i)�	��'(��'��Ŕ��y�­u�Ԍ���^r�N��p@��s��6��O"�d�O@�$�<��A������pS�*��3vh��@��E®�K��9�M������O��D�O�u�V�?��j*P+�B=G	�����U<!�)l�П4��Yy�dM���'�?a����@�D�.����S�ÃcvH��dζ��Iߟ�	�� *6=".Ox�ӈ�(x�lT�; �F�%ư7�<���F�M3���'���'a�4�>��UN�,�P�C�|<�s���z���iB��'�6	�'v���<���˕=�����'C�<�����M3����#�F�'$��'���>a)O��K/:�B���DEJDz�l	�����~����Iy��)�Oz�z�;K��Th@�O��<��঑�IٟT�	72F�
�O�ʓ�?��'2 H�JS�I��m:
�-	�O:�SO������'��'R�c7Jŏ,�zq��X+[K�}�GBm�D� ��d�',�I؟��'-Zc�����N���%�e�S04�O��`�=O*���O��d�O����<qrC�*?oi��� ���.G���s���'~��ڟT�'��'j2���QBX����7D�ktaA�v�ɝ'���'.��'�^��R�@�8��� B�Cz]Q�'� �r�#�-��M+,OZ��<!��?a�� �-ϓC��51d#�=:���#E�Nb}�G�i���':B�'��	)�|L�������z�E�X'�R�	�h�179�0˧�i��R���	�� ���z�0�	[��� ��	(,��Q��/'���'��Q�83�+A=��i�O|������ &�P��T>TPS�&#&L�UQ����ڟ���7���g~۟ȡ����}�.�R���&.���i���'�id�dӈ���O��d��\���OP �S�L��a�ٞ��8%�_}r�'�}ؔ�'�"�'$�S^��Ng&@i��I[�Nt�C���=����H�?:7-�O����O.��g}�^��3�E�<TL��ܾ?gD��'iJ��M���<�����D2���슐I!(=�-#��"<f� 0�MK��?i�{�Ƥ��_�,�'���Ot��
�?v�4�HB��
}�~ؙ4�i��^��B�o��'�?	���?��
��:�Mqs �>?J�)�"�:�F�'�̔�g(�>�(O����<�����OQ6c��{2��7�d� s}҈P��y2[���	���&?��5i�OaƸ���M31���IƄ�O�ʓ�?�*O����O8�Q�@f�1U�-3���P7J�3O��D�O����O��D�<�w��6��ɀ���AZ�WeVy���R��n�\y��'?��ܟL�����r��97E�,H�*���$�
)+�m���M����?!��?�)O(h���R���'� qZ���o	����MF�̑��wӔ�D�<q��?Y�^������ٵ::�jv��F���tk�Pt��n�����By"f��uT�'�?���j�*Q�lЄ�q�%��E����ʀ��O���O����75�|Γ���n�	 �B�c�l�ʀeC��M�)O��ɡO�Ʀ�I̟����?	˨O�NK/����!l�(~�8�h�cy���';�������<����*�2v�$Q	�E߸V^�p��;�Mq�Ӥw"�v�'.��'��t!�>))O�+ʁ��{C#�%|`q@�K�}*��w����ly��)�O�(��"g���V�	�/|>�AT�\ܦ���ܟ0�ɕ݈p��O���?y�'��D!횲4&�,��Zs���r۴�?A.Oݻ�?O������I��@!����u�ЄH&?&��P���$�I�:���O��?�+O�5.д��A�9�6p�$IA�yR�Jq��̓�?���?���?�,Ob%4Ҭ%2^�� ��7� i�f� jB���'-�ԟ�',�'S8����Aݺ�aU#�1�����'���'��'�2Y�tB5)���4�12+j@av���,�����Mc.Oj��<i���?���n��8�gd���ŗ�S~
�C�V��ͻs�iu��'�R�'v�Ƀ6��p������,}Y���1z���%bO�h��iq�ijr^�@�	˟��I�VV��g}"L��)#��zf'ё��	j��ґ�M��?1*O���4@T���'���O��X�,�2`��@A��R`!�>����?I�_��=Γ����t����e���ڲ��BEF:�M-Oa����}󨟰����(��'�
*&k�Mʈ�k��٩~����4�?q��zpϓ����O���seN"�L`a�̼u-�mQش+4ȩt�iT"�'ZR�Om�b��� ��nv4��!�+�\�Q���M�SΗ�?IM>�(�Z˓�?���B���9�u��,�~��vFʝ$�v�'���'�t|���$�$�O.�D���Q援$��Q`i	!���d�ΒO�՘�DH����Iӟ��CN�:��S�+݂ vd<3a����Ms�t�ꡛ'�x��'�"�|Zc�Xd���p�d �KӸb:ĠZ.O> ��|��'���'��I Q*�sCM�$�����D˷T0T5XŁҀ���?a����?i���H�ٰ�A�d�EH2bF���@9��M�?	)O.���O���<	��B�'����~�$�(�ǩ[�ZS���L<������?���pn�A��}� �Z��HoD�і�����ؗY�\�	�����~y&>324�޸@@��a�{3�D�5��X���	Q�� ���6�b�W��1,�ꌓu p��C��;����i��	�q<��zL|b��B��HX"�$:�.�	O4$�P(V�P��'�b�'{�<��'��'��ɗ&7�p�#ɮ8
�ɠ��F՛�V��Sk�%�M�T]?=���?�i�O��cņN�$0�����H�*��q�`�i���'+��"�'�'zq��+4GH��J�����2��(�"�is
`�ҩz�8���O��d���X�>4��
��Iz ���1����Pҙ)�6b]B�|B���Ov�҅ji�4fje�[ƈ��gJ"Ekش�?��?�� ��O������hD�I����ٝ����/|��OP!�;O��˟x�	��(��W���p# ֢1B���,ȼ�M��4����Òx�'	"�|Zc(��ɡF�d!al��	7�!�O
|q&0O�˓�?����?�.OAIAbY�����5�ƃ���KBP�2%f��>��䓯?��q�9Z�oN5�>9۰��� ����
B=�?)O����O��d�<I5'т?�Z-��О*�ʝK�&�6�>8��Z�P�	B�'	��Oҡ?(d��)��G�̹3�ŸC�R7��O^���O>���<�S,�#�O<(ث�L�6͊C��0}�0,��'u��=I��,ei���?��'\�� �H�,]r�9g��)�"�i�4�?�,ON�d�&��˧��d���7�T�a�z�:���&]�p<�B�����?q��?s��s�Âp�S�ԭP-�v4zC�Y/��"���M�*OF��#�צU[���d�:}�'D�1c+Ɇe����u̺*�4�?��|��Gx��,�:N*��K�
�0T�W���M�S(O?*�v�'���'���-%�d�O�q� x]z�E�<G�ȵ0�1'��P��i��a����ȟ���C_�������?{_
<`��߮�M����?�'ٜ�K-OB�'�?��'���U�A��t�VG�J(�J�� �6d|�I|
���?���MC�U?�HA�㛍wj�i�x����g)�q�'Z�꧒?����Ʌ5&)R$�>팙��⚥;�3�6$�O>���?����?���*����̋D�r���kt�����·�����O��D�O�O��d�����^'�@�#u"C�,���xӀ=�����ϟ��}y2�\�o�瓃&be�1 ץ\5���яϭoF�7ͥ<������O���O��bb8ON�*�N�5r������2`͉3���A��۟��I󟴕'�	ku��~2�� ��ã�#�����Ē�/�ҩ��i�S�x�	Пx�I�>���	W��4D�HC��,�޵� g�,�8m��P��{y��E�ik�'�?Q����T ݠ<L�!�uG��."ZU�R�F�4���p��֟���/|��&����)DY;�B2s�}@��I�?i�l�hyr�bV�޴�?Y���?���<��iݍx��á&���8��A ,ʀ�{0�b�����O�j�2O��O�>�sq2��X��M -���g|Ӭ�QF�Ԧm�������?)��Ol˓?���Bh��\����D�ǎ�\�V�i+P���䓡�O�r���X�bb!`\��T����HU\7��O���Ot���Uk}"P�l��o?q�m�^1���Q� ��5r�#�ݦI$�p��.o��?������L����]~J����oȈ�M���9�h��_���'"Y���i�a���'P�LZ�o\�+gxd�u��>9�+�<+OB�D�OX�d�O��*(3���+�`鎘&��"��T15��<���?�����?���b��*�����(-��Ěv��!4��Z�7?Q��?����$+v_ެͧh^ 8 �֩=����$Q�=\1mɟ��	ߟ���k��wЦ�9�'��m+�ē,c�DYKQ�,".�I�Ov�d�O~���O��Dڔ���D�O��[$JJm�&�wjT qJN7*kJo�8&���I��%g�2u߰OiH0E�;7������N'���1�i>�'�	5D�6����$���O��)ÔT�4I�aꆺx9��iچ|�,��'6"�'��
��y��'���'��I�8j(-  �Җj�|��#ڮ0���Q���T��M����?)��J�S��]l̤ �q�P9$��9!6��3�27��O���68��[f��'�q�ʤ���ʢ(�}�nN8���p�i��P{ӂ��O"�d��l�'p剐t�T9�hΆe` ��'��w�
�4&����?�*O��?��	�SM���Ao�j�HW��_�,M�ڴ�?����?Y��ХUP�I_y��'��D���	6�B,{tycsHKk]���'��ɰi�T�)R���?y����h_5jQ6dz�`l*�DqնicBF�
Lw����O���?��b�����M�e:d���o�Vq�'<��"�'@��.>�Rƣ#*�f�y��T�B���E�^D���[�j�e&�T�xH"�@"�+b�(K��Mي���%$�S�Fo
����.QQ��Y�aA8�`d�V���i�r��1�͎/�L@2���(�@B׬�N-��	>G����-�70\�j�j�{��,����1����Dڶ<؞�Д��1&��q
��z�Z@W��2A9��ĕ�h��6HG{j:h�1��	���p� �E'� P� �S��yNv���ȴK�b����<��(�"�ުpp�����'��'N��aҒ[������R([�Sq2d�јK�T��  Jz%�v�y�'gPAz�@�|w�t��N-z�@���fЍ��+��X:��Ʈ�%��a�SG^�'rb����?a����I�Ng�mz�τ�o!$���o9�yB�'O6HtB��/�&!�+B���{�'�'�,���.�t��f´j�P�؞'�����>Q����R0p���$�Or�DI4m <�w�U�G���#Y��E�� Gׂ�z%k
��T>��|�	�d����DH�`/&����}�a���ѓx��q1������)������.��2��5zf<��˼S��\�	ퟔ����)���;�L4�ȑ��/W;>j��s�^�P !Lِ���ML,<FxBf6�S�TkM�(�`��E���ZH⍡S�'iBmE�'�q���'���'�rHi�%�	�r4eF�e��XP�ڕ@�~�F�û�?�̖2���8'�NP(��3ړ6�@����
�,�3��@�d�p�'�y�s
��$<И)��KWF{��ջd^)ke�ۙs��`:ʹ�~�*Y+�?����hO��~�ɢ�I	�;<�5"�ݗ:R@�ȓ(�%q�Ã�~B�bq"øsꢔqw�)*/O�=�A�Bʦ���u�������~�rh2������П��ɍ_���I����'_��X��4�?�a�̡���{!��.�z�� �Q8�\����R}rC�(z��y�iU!V������Ȅ�	�X���O6y9".�,g��RǩE9�b]{�l6�d�Oh�$4�)J�ɕ�H�^$��b �ּm�f�^v�<iuMC��.�cʝ[��q�N��<A�P�<�'�&|��la�x���O�ʧ`���g_�X�(<K���	O�hm��?����?q�k۝�?��y*�>\�t*G>uR��q�Z��K��)
{�?� A��W�.�0 x��<2��!2c��#1f�d3�'2����C��b,i��JI��Ĵ��i�4��D̎��X4�b�ZK����	��ēm��ThC��ELH%K�g�TGތϓK��hԼibR�'���*fS�������	/^��V���7��iْd�E���ڇg�h
d����� 
���k�t��'�� ��C�z��eK�-�Ra3$OTI<Hѓ+i�f��L[����R'�
��If��F�pr�Bu���@�'�1O?��4Jܳum�"��(ƭ�%8!�ĝ����� o
Y+|9%�=I��h[���?!ȷ#V�DI<]iW���[v��R�Yџ��ɯZ/tб�^��Iϟ��	�u���yg<wg����I��)��W�T'&�@l��+��kd<���!<������@�p�aU�ڰ7�~���eY�Y�E"d#�K�R���G��}Z �ۺ��ɚJ�(K$�	z���D5|O��AΔ�g6P�����"��"OF��C�Ϝ:,I0Ɩ=�T� Q��C������Tܦ�*p�Q3{��x�D��r����(�<��ӟ8���
w�����'[��!�۴�?y��ł���$������qɇ`8��AA�|}2gR;��P�NV�J��y	I���p>��%���d���a����U�,zb)��G<��I����'����?AA���6�&��,�6!7��%L4D��+�
�u�2�37N$j����~�h��O�˓6��ujT�i��'�ӊO���yԯ^:x�ܑ�5GA���-�@ANܟ��	��� [���.�|⴮�qnhCr��}%*Aڄ/�R�'�̜���)���6�4+J"�BT駉^�[�Q�X���O�}�F�Ǒ1iZ��"a�'N�m(��Ia�<aR���L �a�:8l���2J�g�<�L<��g�}��8��L�`�-q�4�	�k�^E
ڴ�?�������H}��d�O:���	Z�����㞒5�0�
�i���6��O�c��g�'�Z�!R#�D�� ?NR\Qg@C�C}�"~��0E���c%����XrbnЮG�~kD�����<E��u��gZ�)��Ma愙Kf��ȓ;=�`PR�H����㑁lLDx"�<��|���_P��5�X����Q�̿mk0l����?�b���"�����?��?�A���4�,UY�(щK�,������"�O�
�M��c3lO�+�.�6 ,a��:�~|��T��M{%��!�0�{օ�_l$�3�+B����� 
/�e��%غ~i��s�A�	@��dpb2<�B%£@s�yjsi=�����Θ�rCo�-$�R(ݨ(4�4"��4�T�O������ψ!�RZ�	T'�<DV��I���ߟ܈�kEޟ ���|�fa��\���8h?Z�EF	>|�y�A �'o-�ńț��<)sf	<8V��Ɔ��!�D�7$J�tj�� ��R+����̯��<9��럸��(Un�)�jI�bX���㐁]
���I_��h��.mN���WlG�[4f�����'�ax���e+R�9�, +A�,0�B�x�I��Mk���Ğ��o���Q�d��10L!�V�|��I�vh��C�p���'X��'��!7�'=1O�S3�ı20B�#|8���	��JȢ<�6� X�O�:��]9;�2��^�bB���<6$�����ڟ���R��%^ӆ�(��C� ����iNI2��s��r B�&�RÞ
o�����1�O��$�|9!�H;V f�(B�<q�,� er�4pΆ�M����?y+��)�O����O����6����f�¨}DFԸ�>k��� @
��}���C��M�Oo1�Ҍ�M�HIdd��jC$,��S�a���ԋT)�H�t�N"���a���'�P��N��(墽�6���x5�=Xq�Pʣ�'�1O?��̔;=��J6�ƄHȄ��aֽ%�!�`��AP*�dQbG�����+W�	��HO��7,���$
�?682�{��Σ�Q���`��*6��8�I���	��s\w��w,ڠ�G�?I�P�CAM�8X �'M yi	�H�d�@�@Vܺ�R��_�ތ��o� ����c0B�"�OL~���`��	�f�t��|b��D#|O��Z&	��s3��j�X}�T"O
`�N7HFi��o�7U�~�R H�����E��oP�]cT)I�s�p�5�(o�]+RM���0�I�P�ɽb"4u���ϧ NM*�D�,u� ��F��:G}���O��k��e� ���ҧC:��<���Uwl���mΌ�2���i�Vi��)�,U��]�©ݢ~�ayRCS��?�S�? ��C�2�: C��L���i�"O�i��e��Mz�Q��[�Z4��"O������&�������yd=O@4�>���,L���'�2]>�*�J<~qQQ��E^Ě"o��]����ןp�I(
�����~�S��k�9}�h��j��XU�-��� �(O�|���S�2E#Z�5�qQ�U08~�<��W۟�F��X	q	a ��é'�pУ��yR�e�4$0-@"��YJDG�0>�S�x�oܵK�<G���T6 ���-�yB�I`�87��OX�$�|�թN�?����?��
͐&q�<#���5{�9�ɐ�a��H�������%A�Î40��.�>~��i��y�����kZ,萠T��Q8x��5�)����'�1O?�$�==ꦩ	#�Ԃ`���91�I�1�!��J@��A5�^�3�P̂��
4��\����?��4hS�)��x6�V1A�Q!U
�ٟd�ɇ8�,aZ�/֟��IΟ<�	@��wXTUA�]L���r��֌s3�pp�'�TUȷ%�O�ز��F�QA�W#���� l� �gUD���Y(��,a�?q�G�$BY��b�_'
�<0�X��?a��Z,�?a��i��7ݟ��ǟ�'�d:4*�>.��D�JX/��2
��hO�š߅.hr��!P=|��=�S����4��1�x��sy�랿"x�2aUXq��]+W�R����1. �	��	ݟ�Qv`>��埔�H��W� $�	�aC����ɿ LD;�/�8a����d&�N+6��E��ukg�g�)�G̳1(��iG��+G/,����gc6��O��ŎR.q lhB�2&_��#V-^�U��Ly"�'��O�4b���� ��N,��I!NlC�	66A� "�gZ�+z.|Y %n4Nq�ɝ�M�C�i-�;n5<��ݴ�?I��򹀃a�ި$��� �eZp��#C��$�O>�D55T��<�|���ֿj0��0�II�,S�X���G�'=N�����G$:����A���� �IQ���Ԡ�O����O���|" �B�\P��I�O�\* �C��6�?Ɍ��9Oz��@�$�}�@�(\F����'%�Ot��a��S���GJ�(A$-A'5O�0A@����	ϟ�OK�, ��'��'�����d�e;�I�e�� e,Ą;=΁�ņ>�T>�|���hs��x�!�Ux�t��<���!F�=9&q�N>E���G}<��K����C��j�x��û�?a��?��ň���N�`��R�_�*���b.�<�yB�'��}iȔ$e�m8Ŋ�9֨��ge��ORqGzʟ����X+%���/��*��'�O��1'�x�+�o�O���O����ݺ���?�G��?Ol|��Z2}:y��!W
Z��Ͱ ',�-ڢ��Pp�%̧?��<�(F;)�R���� 'u:A`�� h�" �q-��*��8A�A�-l���\Ō���C���-a5 ֠r���#O�T9��W`��i�n�?�M�gyr�'����8����CN�����wiE���ʤ�����3|O�]
v�I�@K�����m8-�f�`}2O˹xz6��O�`�D`��,7��V�<mJ4�r��8��� YY��D�O����O<%[�5�����O�0��F�Y���kV�pɐc55U�Dk6.5
 D����#@�� hF�� B�B�	\ b	F�G)oNI�.|O~��f�')�6�u�d@A6��m�$��g�(f�xmZ̟��'v���?]!�7��/��w���R�}�T��	$W	�Ii'��:B���v��Jg\�	-z�h��4��U��U��C��?�(�h4Ɂ �4wE
�)vݟC�ܡ�����gx��O���>"�t {wf��V-�a%�ݗb�$q�O?jaApǕl���B�l�`���d��oY��9�QX��X+�D�[���{i����k���2�Ⅶ���Fy�/�?ч�i�"�'9��x~�P�֨A�
�{��P��l)�	���	���i>�F{�B�z��i;�jR Q��PR�N9�0>qőxbH���u�Q�Ǉ6U�@b�&D��yb��cL6��OP�ĵ|���\�?���?����B@��qɕ�/��5��"Q��&옧��5��"u݆�Kb�L�Zl\���	��(2%��44��<E���n=K ��1�np0����n�!��ֳ�?���?!�����Kԇk��Y��ϋ�9Lz��4�y��'��}� E��t��>��xv�G.�O�Gz���i?�H�W�bM��I(&O2@��?��!����w��?��?���$N���O����M��DIāM�$$�)C
�=�$Lsr�Z@�<|OEY�b��Dt�'n=�!Bn���J�oB�˃C�)e��I�6�]�%## �����lŏ%%���I4\3B��I�D�t�'�"S�� ���da�-\��&�҃$n@�v��3|O q�vCՙCU4��F�up�	u�MҦ�۴��D\���ey��"o���]�b��!ԯ�VK�A��O "z�]�	ӟ���՟��6��֟�	�|�h²T�nՐE/�J�Lx�dN��(v�U9AHH'0�I���	<��<�î�;
0:���3}�=�����E��͑���*�l=8�V���<���
����	���� T�_ 4̵ئ�<rX��Iɟ�'����?Y�c��K.�4�(�b¨1D�䋖#6�6]ʠM�d J0Z�c�ܚ�O��t�p��%�i���'�哉H�Sc�Y��]x�o�,`�x"�Y�@��ݟ��Ԩ;x���`oM~*�p��g�ɔP����KU�5:DT�V剱Zj�]�F`�P;v]���Xh�J�t�ʢg�9�D���O���<Ia�՟�	؟��	A���%���ic�ѥ��퀐_�;|���s��0��2�tX� ó%�L��E.�O`�&� ���;_���A<_�`&�a�Lk��N�M���?�(��!���OR��O0]�R`O�؉j �I�-J��jtLmZ{�S����qc��#���Lx}۰�X�y(n�p� b�S��?a���!g4�mJ')�a�4ĄF����?1�O����O��g@��\'�x��+�X���=O��d-�O%�F��8�l�(VA?�䀲��I��HO�Ӭ3��1��ª3rK�i�Yj���ݟ��'��9Dl��I����ڟCXwm��'����\^Δ�sӌ��`�J(���	�@	��J�''���h�K�����ē%&?$Z䯛hK0���,Me����E�3r�r��枡(� �U۟ў�A�fNp��L��	O9l�@K�ʲ��4��O����©0F�P��$٨m�ƅrDB�$y!򄓦Q���B�5K�q(&��>|ƔEz��ϼf3<mn�6���L�3ڼ�[<p,���ȟ�����@�͑���|b0�����Z�>���#�{���Cg�hZ����U:l�I���Ċ��$=X �[q�:�@�=W���I��L��-m����]32T�x9R�(D��+pj�0;�&��$�Y�� �5�4D��PA�)�АZ��Юi�J�$Ex��b�}Bc�0�Z7��O:�$+:�)�Fj$�V��w�:�cuA�
wbB��	��@���Ja�$D� <4�ҧ�74c�X�p�A=T�r�Jp�޺O�Q���*$0$�@3�S���Q��IW�E��=��B ?y$��<�W�Z��I�4��~��C�o$2L�B�@-;G��_-���s��)�
N�td\4
�`�7z���f�*�O@,$��	 �[�}ₕ��xB�t#�ic���E��M����?�+��AAW��OD���O����@~�a�	7vK����Aބ�
��?�|Fxr�Ӄ6���r�f�4X4��K��-ǚ�y��)�� ��K�<2e�c�@?X� P���)c�@��ԟ������'i��`��ե̀0iv"�n9Z�X�'fR�'�6akV/yqF�+&���7�X�I���T���IM�+i�+��)����Z�����Oz�L�?zA�$�O���O���;�?��@�\Qr�A�1l��W��8��=��,�T����n����ѫ	90 �͛F N�	i������<��%	��eٸ=0�ڍx��dE)I\R�'�*db7��(\�NA�UD��Y����'L���wE�&�pul�9U�<�b6k&�S�OɈ����yӜh�b��<ن@P札��c��O��D�O����@����O��S<:���xgCŘh�Y���C�k�8�1Kдv��X��>Ly�`�������O(	Ҕ;]�8������� sL�#Nz��R�!Y8��q��h�G~����?A�ra��ggܣ���%)�E����|XM�1�V�U?��I�	�b��h�ȓ�8 ��F]����Pnܙ8�1�d��O*�����d}"�'S�S�<&���3/�;2�����
�\��D���������P�G̈́�;�l����&"�r�j�S���T*W��ǁ�-!���`�%�)�(O&!B�wZ��T���t��8��!_t�LJ�"�QR.���I/K�b�$�ަ�����A�dZh�����=��	�E�y"�'B�}�/�4s�N���F�}�ΐ� �2�0>���x��6LU�]����x��u�`M��y��'���?�(�%���Ol��O~A��oݭxD�ᐐ�[-;Ը&�հX�m�Dƒ rA�pg ��M�O�1�B%�!y^Y:ţ]QbL1ӢOA�jT� �aa��CS�Xg`�(��@����'��Mi�bX08��ıS	�$WM���o�6*��'��)�	�O�ʓ:_(��B���R���9��Ir�H@��S�? �-Z�ֵ8ư�p���RW�x`��	��HO�S
�6�ȱŎ6&-�  ���Q����d�`�\����IߟX�I򟐀����$,[By�a���K(��*������r�����FL���������/>X��d�wRJ��*Vh�8�T*��%�/_����Wc���$�Oz�ԟ�I�@�'oXh9�쐘�&��.C�&�j�!�'���f��}�%s�C
,��8�1���	�<�4���|r��!$���c)�.�~Q 1���'�2�'#�Bq�'��;���ar�'�A[	&alI���O� ���+G��	�p>�@)Xyr
NKd���C��5bONp���W��p>�A�����r�.�2�j�CJ�a�"l��C�I";��бb@��L͸ ��� *�C�	���s  �s҆=��O"_���I���?y�ś�E20�����8�,�h���k�<1���9�'OP!#J<`��l�<yS�Q�:B �@��U�X��1�e�@g�<�W�R�%�p��g����@.�k�<i��L+"��c� �o�`|��Ps�<��j�a��jB�B��0�IV�<1�K�#®�P'J˫_TVi��#P�<!R	� ��y{�� �l��$е�I�<�$�è[��`>�>M���_�<a��*	��xC��^y"�ЂC�@�<	�G3ֆ�a���7(����dBa�<1��N�DX{eR�5��@��OE[�<����Zh^aJ'�N�Y�6(�K�<�'b˪m�zmy�"��"2�p�Ȁ~�<i�Ҩ���.!`�X',�z�<ѧ�U�SJ��7�DU��9��[�<�����7�pV�
)Ez��OW�<�UcH�
2Xk��0F��9��P�<DH�24_�|�m�- Z*�Q��H�<'a�$(޾P�#6��E��KC�<��╍-��m��w��)!��|�<ɥ`۫dzB!#W�ȳ����R�D�<!���L���`��i��`��B�<��EM=5`8j�*�-x��CRAA�<9�N�S��B��>+|����y�<��ŇX�tM(0�7YZ �1v��m�<�S@I)J�L`G��,����bGNk�<Y2	�/ ���
��5[��	s�\�<ɢ��4��ɛ�(@0 �a�L�,�H�a��y�'���O�D	ªQ����;+����C�ŐX�$uA�M�@����	� �HTic����Yra$Wp��0n���ĵ<	4f�R�J<���W�r���Z�ď|_rr��D
O �Svf.0�O�-a��?ex��
��M�p����>iB���o(���H\aG�ݸ��Єf�X�����
�$rL˭;���D�=DPᣰ��27�V�ʲ�H�
��>b(�PZ�G�;
�bd[D�?��y"�Eunġ0b�,l��L㦥�RXE�cG:	�����Ѵ]1��Ε0�%9r�i�Q07 ��/�.����>�OF>ػ6
֛�5�A��(nZ��w�+^���׹>X����9b�6�8ӏw�ܵ�%@�1�l�4�ֱ},=[��_
�iA��ٌ:��BT��AR�銥o�?�̪���@yZ��b�4�H���_� i�>)�
 �b�^�-8ҭY$!��� �@��EH�H��߆A��H#��r"X�i3�U�@��L.o���	Q,е��"7�Bpb��������`^��# /F,<��c5H�ZިM�i�����0$���˺>�'rF`�Jԑ+r>ȹ��N�#��%o���?A���.�����J�S"�09���$�x��h�'��y�
�g�)�	�#��|���.M��16GD��4���Є-�v����65��uk��7>�F���&�9��H�U���O&�X��O��	L����\p���9#Bdb�㙾A���E��%�~�*�61��e�%EH������	��OXD�g��&;�� �22��Xy��T<.z )���Z�K� ^�h��J+j�����Z�#}�0�-�ڬ��RHk�'d��ӁT�y�V�I��m~�t"�o��8��dDE�2ǐ�8u*�����(B���'�d��7�ƱJמ����aW8|	�.�	<cl�p�Ia��8���R�?2���B L�z�C�G��8.�t+ҳ=�<%�0��9��$֧_�S�7��)ϻb9D42��)Pvf!��5x�Ć�	O�b�%�!� ��8�6��z(Yf�<��d��O}b��1Az9bA�O]lxB�NFnA��c��H�*�X��)-]*��4��"�*hF}R'��J��С���l|b6��$.�x4�X �T�z�ΕD�AJF���%�@ōgN�]K`���pH��I�0��):�
�1z`�1��x�@������K��x4�1*R�-�=��98�6 �ğd
7�DE���u)�Sb� ��EIdO�b�����?��h#��F�
X��$�4+xp�%���r:�=",O�������pv���^�ɶ�i0�$�
bYz�0L��^���U�[7p̒���"AD1�j8_=�qs'�Y�}�H����Ȧ-Bg�'��7�mY��Yai4}�giZ����hLQJ�!&KV�+��
�D��@�I�K� xX4�M+pߐt"f�� &($���kCZ����ҫi��:�MZ��'ǲHId��+~V��8#IՅS��!I�,��?�%C5H	�uK�t;�	>-B�`@��:x�ٵ J�
|�J�@B�@��2�I����B#��# Z�(%hO�NLty��t�l:����E���'��D�Č'}���ejNG����T�[�Q��y�c���Y��40d	˘I-џ$��ʼ�墁�Y
U
Q�A{?�}�	P ?���RDү.�jA��²�E�O)1I4݆�	&G�d#ԃҿ�il�6ie�A#�:sԀ�@�̆���O��[��tc�pB�[�i��E
�6��`��,Ƀã��.(JO8�I;k�P��QȖ9A��y8��C 9�x�')��	g�w鎑���ʒb���b�O�=c�m��!�hQoZ*l������M�#$�,���~���U��ak�I�f��I��AD�������,mB4Kפ�)�4���"�d�۲bM5p�7 	aid�	�m�֕�U(1����>Od��R �vH���ߝPm\�
�m �`���i<)t�]9�a�� �DE�Lˇ�����v��^�*˓bҦ�Af	v���nC=6��,�Z����a�=6�Q��a��V6��'�̕'nP����P9����20�.O
�A)O0 �R�5:����J�<�$[�T$��)� �D��}�N�Pe Y�:�������IR�IJ{H�İ?�i"Õw�R��3˛����Q���f�0]{c$��}3��[�>%�n�G��?c �X,/Fȩ1(ƒn�z���/ʓ��O���NXX��O;;�z`N�!b�B�
Ǔ~m�-���m�n 2�]P4"·2<�����/NG�|��.<8�ȗ�q	ޠBr
�3_``�5����>���T�0�$z��	@O|���c�<X^��3OZ���J� شBΙ+�����I�c6��&۵H��k��s���q��%��m�dss������I���pIԎ_wW�ݴsj�I��6�X*�鉷N���녃T�{e&� �'�Y�� ��Xd��n�p<��H�AH���ȡl�tym���M�����'� �+H$#��q R�L�iN֌kR�F�[s����JX������Z
!�~����'�~���**�����׾�Z�v�D�tO��o�H��'���)���!��ba���-��C�Oћ&�×���R3m �I!�0�� ��6Eq��� ކ�8��H�#/C�M5�ɯE8�-��!z�)2dei��{BY�9Ķ˦˓�:H)!c ɽ3)����lZ�h�,����2r��w��ԙGdK�,:<���� ?1V�ĝl��lX�"Z�!�Fi#Q��#5H���ݦE���c���<�p�ҵu��W�̺$r�œ�.�<M�(\�T���=�έI&�J	h"��	H���)��*n�ȸG��^� ��']�0��4T��z��]-�����͝`���� J�i��̖�p��t��KuF���Ǹ��Po:M�J�1OI�Q4M�HF"��@B�` Ot��aR� ��s�D�֙����q%�T�Fi�{�h�2��$j�OƘ��L�+HcJI�p��_v��֝>QF��:�riQ.�[*�s%�Ly~�L�G6.U��B�2J�qGJ�O�8�Q��-����'P�[��2M�[��ܰ�e��+�+�����p<IFFJ
0� 	(0�>6ǒq�E��$䤥���B.��ɟsК8��I���H�!��0���;k���6)����F�w����a���X:�ެYS�7�4���
�K^��"��Oj���R�BgԊ�k�sRQ�H3#�͟��V�R$?�Ո�c��|PwMYD!�R���nW�,kъ��'�Z���䊒\B�;�n��k\��[J�)�C
q��Ĩp�T�sX�lcs��R�����'ND9���v�J˓|�*c�8�BH�Ph�:��&Z�aЧ�^���
q�֌C>~h�A�A��x�jR;8d9�"��.&��{T�-&Ĳ/OH��
ۓdhm[��
Q��H�OZ���ukE�&\O�đR!��?��%A�^�"Ha��W(9��*�Q�8�=�F�ў>7�T#�(P����B���)	����V��1Ǯm����ȕM�r��D�I�JC��	�7��3p�Ͽ.�n�XC��M"���>�uN��?��mq �С�1��jy�	�M�n�B�)vRyY��!|����Ɓnd(��e�����<A`�-�	�w[E`'5�l<�үW���y�iё��pP��ֳn}z�F|��	޼ ���E�Zer�J�)7�t�z��Rڦ)OL��ۓ�v���,�4G�Z�[�-�3.�H��$Ň*�<I3�A�V�VaI1ʜ��n�^z�ZÅ�M�h���R��J���U�xZ�0��Q��zy�� ��0�HU|D5�O�3s�" 2O$1R�OD�1y�81�'�!0���2��OpQՃ] 
��5�QN�8݀Q���3�	�.@(mb򁛊^lQ�2���2�l�O����/n�@�Ac�6�^�H�	�<��������Oh� ��-�d��OR�a,I(4�!6�G�l���!�PF"Г�J�8"�L�r��6��l�;u��X���lQ`��	�Q�>�%�pb���>�SC�>�@D
����O�@��T�s�|UB��g�����!hb^�hv&��
0�@��b�0¦N@�!��a@�Q�$��,[�2����f�DI�>�z�T$��Pʢ˓ T y�M�i���
�G�G�4@͓xP4���@ۍ �dA{ D�`� XʇE�Y�O�I�	�X���F��[mT��e���=��K7ک(���?1�$H8�i+8ډ'�t���	�(�ͫ��So��(ƇI^�1���j}���eW�B��x�"������Ⱥ+�0��T�n�p�V�Aji���6A�H�".+uQ���qލs�o�,A�z��Ģ��Lj4Yw$/�]��Ti��@�Q�|�V��D'�?!ȕl�@�y��^X�2sӇ�I&|#�}��� �BU�^0�d8�=@1�l0@��
p�za��)��0!WN�-#D
�5�F}��R��c?�`D���;�S�۴�ܸ���t,A1t��'�y�;H��0BS�4��|0��T�=�X���1���\��}
�?XNԌ���<<�'JԷ \剂C���t�_q���3u���#$�^ !�D"P>����"#=@v�0b��P#�#�� b�TQ  ᛻9X� 0֟�q����6�\��O�2MXTu8��'xibe��[y$(рME�c�p��{*�8=�A�zGҌig��E(�m�ய>9�'@�-Ab�W=p�ʟ �Z�*,�B#Yj����dS�2�v13���8^	 5��.+�|�ن|�t�`b(Ys��=��d�n�:D��DZ��@^�1�'�_�)`v�APC[D?�~��D�] ��A3�<􋕉U+���!@��!�y��S�X�P���:B4np��~�>�e.�#�X-����<16u�q!�N��d�<��;��۬K�8u�O��#,���6q��hQ����s��<2�`cg�O�sT������#�9o���λZ�mbm�3�p���"�x4�$����&fP�9Ǽ]�!�CkX�|�<�O�1y�i��/��3��q� _��0{�a2K���'*��/W�8%���]�nf4HJ�W���pчC������ϛ]�j� �<F/��<�lu�#±�t	S��3 pȁ�G%~B yBǰpe*9&�<|lt��|�OX��"Pd�|"��-c�hD#0O�B���r�>�0"�Vp�X���0`Lm�������y�ԅ�9J��	͓��ى$c������i@�ؒK{��?���SҔ��4��H�!�`�T�Q� I8!EYM8�8
����0�,����D���I%�[+^���%��
)�L%Ku�ϰR���0�1O哀eEX�2�Xa�ۥĴP�|Gy�ڕ!�Y�6�H8!B�|��БV��Rs��U��x0��l�
;dm*�|
��	+(���h��y�[�F�&���JQ�n�)��t(@IQ-��8%��~��$H��bp��`��/��(�J�l������J�V���T�bxeQp��g�ʵ(�H�7 ���2CP�ɜ�l��hX��ɡ!�t�	�܈���u���F�'r�P�[�ɝ����<Y��/I`l�s��0!vL{BmŮ5�h�M�$��*}2IϷZ˔�	���U;��$8��u��g/v�(�"��S�~A���M'���`Ӏ�`b�93���r%�˒Ub&��ߟUH�4�w�UJy�N�zwF�S ޑ�\��l���?��o2~����]e� �"[!䴣t�ך��5�Q�Z P���>Q�I^
�~��妯�t�V�>U_*���۵o�z���^%�'����������V��_]�|YQ��N�J*�:�� Y��J*_�1OX��B
�p���I!(�8�d~�;�@�0����1L��A��]�sp.P��#,	�����'��R  Iٲ������Fe �`���O䠁�?Q@�e���^��sT�_85��\KD�&m��Q�A>���Qw#ߕ�T�k���|F|2�ӽ�V!3"��6�Ԙ��D?�8ܙ�a0r���F~��D����;pj�檅"=��٠‫4�Z� ���!.Z�>�'��-Z��Hg��� 2�΍��&�h�&J�;�.y��?LOh5i��=��	$u���`-8$�:��?��Pu���MX �E��b�
4��H��G>L��xẾ��'�R�c����TB��<� �ƍ�
BD�,�2�կ�yRσ��`-p6���PJre:��M.�yr�ęB��xw"ˌF;�0!A�y��� �H��I�+I>n�� %���y�u��l��g>�Ƽca���y���z�$����g����,�y�޶rp����)_cR4�Q����y���f���`3��/?�^���e��y'M��̤����=hH�Xb�!���y�N�#y�9$��~�i�`���y���*kMD8`�O؊���*@R2�y��N�(�^8bG n�⌻����y�D�,�UB��H�d��ͩ`�P��y
� `(�Æ2-��S��X�&����"OL�9�-�0�vL�J�/r�z"O
����߾M�r��NQ�u��A+�"O�tB�*�04U��p�hZ�  ��"O��Q��J��X�T�r���"O��"ơ�&=^�UhC!.�(�"O���EG`�=#nƻA�(|�"O �)�dA��C�+��wXm�"O[UE�|�p
�!S&@JJ�x�"O����'��a���ׯ��=�٨�"OX�5g�6�ư"/�6d!Q"Oʽ�g�۟�0��J����g"O�u��bԕ]?��!D�z��cu"O]k���\�¨����AzL��"O��z7��U�Z��6m�t����S"O�]ФƁU�F���+����� "O��đ;S�,��q��w�"O4qC��Wj� i5a�;ab��sA"OP�Ӱ�F`)��1T�G�8�PP"Ob�1+FI�H{q��%��]3v"O�p��ǼM�� �T�U�2�Jp"O <�ㆾ����%G�7�ɠ�"O���ԛnÄY�`(a1�|�"O h����5|4��p!��"O84���УR�FQ��$+���"O"	�(H?��ͫ��~��8�"OT�4��tIDQ+�Lϟ@���k�"OY�fW�bK@�顂��1����"O�ܸ�o�;tڌAX1��<�xI@w"O:�1�dǴ=�pr� � t�IC�"O�8��([6>��v"�yctk�"Oj ����w,�q2Ł7pE�i��"O0H ��d�^ԊB/ɗ�X�G"Oؙ����j�=	�%���@"O�s�IZ�^�27/I�"PR�"OL�m�V�Hp�ɼ��|ct"O:�b�F�,��a��'\�S��=�q"Op ����y��Ƞ7�S�*���!E"O&���R:�ޅ�q����p"O�a�m^�0C��'�d�;D"Oʀ��C.L�1*T�R$��1��"OTy���S2n�r�p�M�7�B�R�"OhT1"B����0l�b ���!�$�s��\��J�Ȩ�2�.֩~!�D�22�tD�@ȴA�ni�F�ä`I!�DMVH��*�f5:��I�&�'WH!�DI�PPD��ÙS�jU�G�
�!�d�c����2얽#� e�d�"�!��7S��wEC�o�<05ǼE�!�Ń#L�Z�E5� �bP�L�%�!�DW�D��Sq��e�� #�/J?�!��V����w�ݬh�b�D	��U�!� ;�i�֯\�p|�11��F
�!��:�4,��Ƹ&_R	���U�}��'4�$�@@��ȆڃIy^���劼TD!��V��A�IF5�R��ԤDm4!���=wQ���R�HN6̓U�QXL!��WK@�2��<C=!t��	},!�D �/�tp� l�'�1:�
�.~!�DjL��
�A��h3V�L1OX��dи���8�Cj�NH�l�%Y!�$��L�� "��Ps�M$' �!�$�l�#�eD<+8p�6��;�!�$���)��苘zO��CÆ>-�!�� �T�A�� g)&����-Zv��"O�!y������j�.l@Qˢ"O~�҅ʕ3܂�Aqi��1W��˳�'�O�i��>w^ʬ�7�զ]1z0�$"O\AA��{���%G4+"\�B8O��=E�D�L�������FP��x`̟�y��W�4�,呣Kҟ=3�A�b�y�$N�U"t٨1�ӣ4�L������[��(O>��ʑ�D���$)~vtPR3�>D��bSc�P�,��DF�0�2M���0��*�O�D[J�(=�"Q�PdۺVe�I�O8D�
V1Y����h̔h#��,q"B]�	�'5�:�e	�*8����1mV�Ǔ	�Q��4���d4��F�d�0�L+D�0ɳς�l�����c=u��;�&+D�,�_M�N`T
שVB	b��Ҁ�y⍗�r�#�LÚG�$<�DkJ�y� Z 8#4�x���;C��賎���yR ϭ|^���f,���Ж�0=9��Ý�\`uC���U7}�KP�y�ƒ��u3PF�� )��C�Q��y�k��}
�a��|b���a˕+�y�
hBr%��)n
��1d��y��TN����H�
��$���xO�'���a����XEr��Y!��ѯ$�!Ҡ�wr������Z!����u,S"=�x+Ů��vb!��"h��ȱe��cM�^�!�ę�cI��;�͋�eB�Y<t�џ�D��l�4D�7�٣%=��"�?�y��%H$����|�y������>A�Ob�Bg���=Ӝ��t+1��a9"O\�;1+	����2�	,U����"O P'.ڿ _���C`
������"O�az".�, �%(f �j�Rr"O�Eဢ�3B�J�N�)|xq@"O���#߿��|a0M��V����;O����'�O$lȷt�� ����4ɸ�'�P�𒨝L��D�!|��,�$:v`����M�!��OH�K����
?�%���L�pv�
s�I�0|�'��@a� $�t�)���_�<	�`��MS��2���#^t	�AT�<!��!ap���dm381@��P�<I��@(2�Q�)�C���(u��P�<!�넊f���ʔB�
V�u���ZH�<��͘1}^<X�ǃ�3	v,�*T��`�ň�t�fCǟ	O�Y���#D�$"��N���`�)o?���'D�8q'燏b�f(Z�-�$x*���
$D�\���V��j��r�˩���"D�\��!U�[�%��nH�6���A*?D��a�����)�bŇ\{n-hQ%;D��h�#T ��b�G
}�da1A&D����K
� {�t�v�ҁ�n@�k$D�0���X8Ry	��Z�H�b��O.D��N��G��2Հ�2t����<���S�O4�B�'k�P,Â!K�R��C�I�^
���%k�:�� H�h��B�	!fͲ���0@(�te�N��B�Ɏ\�2�I��=3-�ap�o�bB�ɵ��h�ɳn��Z��&�vC�ɢ)� ��+��ux�;P6B�I�:Q@�)A�[>ja8�D��2B�	�v��XU��5�0Mj4M��*B�)� �� AG�,��1�G�5'>j�P"O���F,���*�C��;�� G�'FqOz �O� 'O��$D]&1���q�"O�#d&4Ԕ:Ab�{��'��oX�ࠤ%�&]���C� �'a`�c�*=D��VD��R�4k�9_�ȁ["1D�|ʅ/G�d@�m�W,N�dql8��O.D�\�֎}-��� )ى8n1��j*D�Б7 �-��B �ٵ!�&�A��'��5�O4�i�I��l�K���4�m��"O�)�c׀��|�Uj�]Ff@��"O ��@�N�A�V����3�5�OnO��J��� zi�\ৃ�k3�E`�"O���ʞ���з&
�l qѳ"O�0�R���n��rF#=1Zl�G"O�]{7o��z�����]~nTJa"O�����I�5�B�:���2��wH<i��P�6~HQ��W�
L�"$n����>��W�Q���k�M��.]��_k�<A&�Π \����KQ�w�<�Ba�h�<9�

�3?
���Ť���YG�b؞��=g�b�	�f�T\ۡLe�<���s��IC�N6�l+���K�<Q�� s� �VE�.f|�S7mLD�<%�\ ;@�*�
�Rd;�bB�<��T�A�\MC�'E�//�"AJGb�<a"*�v�hX��W�=O� fJa�<�b�̀
X� �w������ЈD^�<que@"`�܁r�TB��꣦Ys�<A�&j��QGnԚ'�L��y�<ɖ�U'.z��"����ݔ��cSr�<�@�J�&���EB4��]��c�l�<YE�¸x�D��p)���Pࣁ)�D�<GK�*q�pc��E�v����A�E�<!7���{���O� ,#���<9�C��V��S��%y��z!��r�<i����d���J	#.��}�U�Tp�<�SIv��=S����U4y��Ql�<�֢C�i�r�)��љ2��d�P��j�<Ӌ!? �e@�E]n�ժG@EQ�<��MF5����k�s�
D�<IW�@�#+�5r��
z�⤮D~�<iE��7`�^mHOSd��`wf�}�<�c���h4s��Ȁ9�&(�gD^y(<yٴ68T0�Q�5�:P��u_(�ȓ�F��K� 8�VL$$�� �����e7x��C�J�HP�����.'Tҙ�ȓBor9*a��yJZ�{1���B�
͆����
��VS@|x��^���܇�QQ.�:p��q�By��^/D��l�ȓxW*��3HXn�����)=��ȓCP��֨7a�DjSD;M�ry�ȓz�x:N�#�]�C ��)B&Նȓy��[�c�#F�!�bô{��ȓ.��X����D��D*�ҥy��Ȇ�:�B���.�q(�}��ȟ5'!��9�`���9N�d����Z�!��Nڔ�PD��,`�(Pg�>T!�$ŴC�v�2��֊�$�)�h2$�!�D��3�����f���0���9!��Ȳ4�fɓ��e��!�"�!򤟠��]AU���v�0�v*T�Ab!�*tB�-�,gZ�ƣN�5O!�$�}����ǟ-S&�`s,Y7!�� @��n�7I'��ᡤB3����"O�h�&m�5�P�2�A) ���I�"O��w�ȳ^ �# ��<lVu�"OR�疖U�J��%���-�z�a�"OJaZD ӯ|Fe���4��h�"O�U���F�c�Dx곉�%s�J���"O� YAnD {�!�gH��5����"O����N��Q>�4�'o).Q`'"O�K�Fü&��|B$^���Ist"Ohq�#DGq9r]���B{~��"O��
���,� 08�hƊ%�&m��"O�����э;���[�ng�<S�"OU0���r��(�*Cf \iB"OVi��B�|�,pT��1:��"OƑZ�*�2��4�#L��$�ꀱ�"OH�� lQ�U=t��3��?��1�W"O�9�K@�*���"\%5`�z�"O,t��dE63�TK��J�1�����"O�I:դ�(n)'`WV�r��"ODݒa��@
�[ĤM�o�(u��"O愸r�S�oJ��'%ً0br�s�"O��s�-��[F�M�1�̔L�!aw"O��I�*��+� (�ŁMzI�+�"On,:�.��r��i�8my� x0�(D�zD��tt8eB�l�wоE���&D�,{l�-Jp������O����#D��#�eW \��2�$�-L�b���!D��B��/J"5{F�]�e��V�:D�T)��"j�:�@_�7йA�7D��'˅�
��%���2��YiBa5D����S� ���6�ά|����dk?D������޾���J�_�|�i�m)D��XP*�p�ADʪ�r�A(-D�pS���F�:�k�CH u�n�8�J*D��ѯB�_qL�9)�;+@��ƌ#D�P�V��(�P9#�B�	n*�{(7D�dX��5@�LQB�a�B��*��2D�l3�"�$aZG#
���ՠa�&D��0��
=f1Z��l�n�f�83�&D�l��E�3 -�����+^W`���%D��5l�5@\�չC��
mF�Q�m0D�`:�e	+@8���A`�'L�J�`�(D�,  �^Ƅ�1dN��;x�y3#n(D�4Q�Ċ�D͐�\�_�q�:D�  ���tHy蜖c{����"D�XJ��
'gt��d��	�n����?D�Lѳ䐒+�x��o>��=D�� f��x!��M�?��)�B�9D����Í�{r��/�0��v�8D��ɑㇰ\�<�R4l�(G�1��8D��[��E�6Ջ�a}|n@C��(D��	�x��ǊA#]"�{��,D����I?_�M�r ��i�8D�|��1=�.�!d�>?��YEb2D���g#����RUD�P��8b#�"T��ڦ@/)�%h��I3�"O(hq4.��0EX�#�̖8́p"O� vl[�Sva�S.�:
���"O������VA�0"�/y.�"Ofi��J�d��
�$�R��"O�3��&-.��1m���T˂"O���O��s�]ψ�2����v"O�a���O�8�K�$�S1�\�"O��H��T"C$�e�R��'@���"O� D���IRr0����_,Sy
t��"O2DH�	:E�V�q5d t��k!D��W"#<.�������);�c=D��aD�B������_ h�I�/D��)�ʀ>I�9b1�A��veha-8D�8w�t�µ W�ь���7D��A��#@����1\��j$D;D��v���+�ѹil�ث��6D��b3@	0!��HC����	@PDi��3D�tX�T�~��r�/�8 �2`?D��BB	�G�Xm����
z9�T���;D����BA.t���`U�̺8ܬ��i:D����D�P�|�[U���aOx��Q�<D�hFZ6=� ��ȴ��ċ;D���o6D &���Ʀ>�$�"�k8D�@	(B
�&�#�" `��:�b2D�sv���[H��f�_�jɸ��`0D��ѠnOBZ�y���	)P���wG.D�tr��0� �pV�r����/D���`�la>�˴�Z�r��uW�8D�8�Weȕt�Mwo�>aD��B#)D�$�!�Ūte�4�Io��`��*O �0BIU30"����УCS��y�"O��)� fc�����qRP��"O���N�A���2l���f"O�:'�
<
�T�bPJ_;GH$"O����T}�����Cd�
�"O�ݰ�C1kR4��ӆ88�bɰ�"O���ODTi���2fԦ�H��"O���*ϊ ��pAe��!~@�Z�"O�PCL�!c%��æŅ89�d(x�"O���"�,?���`C�&0��q�"O��
MԢ��}�@cߓ�B��"O�Ū��E|:�eQ���B�6y["O�q�@��)�Ҍ����>�vA�0"OnE�B�6\C`Z�G��Lb�"O��)k�{�^ ���ָ,�ycմ@�j����(Sx��k>�y�oЁ+X�裌��hE~M����yb���=���Tbޚ]L�ȷ�Q��y2kџX� �U�#O�	�w�ӵ�yR�١v��(�J��n�`y[w^�y�5&��Q#)��0kDA��Ͱ�y�'Ӵa��BH(�PHӋT��y��jY�99����"�`"fF �y��ò5��M��e/�p�z�[��yB��$�l�PG	 g$Hr�I���y���Vt@�{@�<(j�4!B�y�jI	T@zy�@��1%NE2`@]��yBȝ���!�j�)3|��I�y��K*,�* �vf�����2�$��y��F��3��j�X��!�yRL�~�^��Ge[�\�v컗��yr"E+?��t@��=Y3�|2p�B�yb�����C���F�b����ҷ�yb�m�2�Z"���;��`Q�˂�y�`D�TZ��0�M�0%����y2�k$�dk�O"����!��y"*ւc:�=��
���N��y�*� x�e��fN�8��Mc5�ô�yr���p}����M�-hԢ%@�3�y" 	0!���g¢tb!�ߟ�y�!��[�-z���pw�K*s�!�d2>:b��c酬����Ca��!�� D33��Kvd���+�����"O�jw茼-Ť��a@͹_�\�g"O�]�.�W�ܰр�FE��"ORH�:2�F�E&	b����"OX%��@�?Z�H��S ߼&R��@"O�PXDG�c�N,!�쪑��-�y��^=~è��s�;�M	�A�!���~Y���5a�$��1K@�!��&낝 �ݎp_6�Z�	Z3�!��	C�`�`�]��1	 �!�$.�z!`�b�3r]�P9'	ڽ�!��9\9\Ց ͍�J[���WG��s�!�dA�M��he�FxK����ǫW�!򤞬�-�pM�I\Tj#&�b�!�D��B�z�
%/�%z����
Ĵ
�!��߉Y~�uq����.˨a A��#�!�-?+��C֚Y��� W� �!�Y�|�I���N����g)��!�dP�/��
���� �!!.�`>!�U�a�8����f���Je�Z�e	!��ɎM���P�G��N��y��"�P�!�[�)gH��iF�j��yK��ǥ%�!��2w1�]JB;IUJpp$ꟓo!��E� |4yJW�[�#B�y�!�C!�d��[�03�#R6����0�!�dL:<����B�F�h��6m�!�@r�D�ECjFvpyw�x}��k�$�Y�Çe����R�S�J��ȓ&�Z�p6N��Gv�,�FDY�I�X���00|�a�� BB�C�CKþ��ȓ#NB��*ǴH���3�
Y;rP���ȓb �����t���bC�!�9���B����ߣ ��kT@S�*I��r�f���v8x�"V�T�D�~���Da�m��䩚�+ָ4�X��l4D�pb#��R�𑡶�ҋB�Pf�0D��R���&PT4�XdƐ��ꉙ��+D���C�����xȒ �vZ��F�*D���'� 7�lY�်>����L(D�� 3�C�V5���@�v�"�3�O9D�|�ħ��p�*A�3�/L����4a2D�x�eD�]�8�u�OQ��D !�5D�Lz�)��i(�mJ��	����ab/D��)Ab��rg�պ4P�T!D�X���Ō�f�"�cްY[ Ub?D�X�jE1%$>i"�d܇.�� �=D��Rk�<=� �s�ZU��:T�0�fB	v-�!􁆒0�D ��"O��J2J.��3�V� �X�q"O�)��B6�>���(ɭ/��3�"O���#FH=	��[&X{d��"O�e[HN	@��m���ܑx,ar$"O�Q
��0�yP�R8���w"O��c�!��qr�L32Q�BJ0�"O�y����C��l��%���0"O
���kV�\�pc��>���[�"ON��FA<_�0�-��dY>��0"Oz�I`F��LYBlGI0x�"O�I�Q�,|Ydl�)���"O�=�w�˫Q�}bvć�A�ْ�"O�����;Z^pd$�K���"Os��[0"��$z�C�=d�f]`�"O��CԮ_��N�jT�ua��2^&!�9.�e�&�_�&�Y��^�U!!�� �);���1>�Ii�iY�6~~Q�r"Oֱ���64.�c�(Fn��Mk�"O� %�#W�*��� �b�yf"O�� �JS�y#&��K��A;@"OL�ce�^'e�8�k�J��PD��%"Oh@x�.9��106�V"0�n���"O�t)���T2AB��<ɀ�!�"O�LI&яO�b�Nq�.�q�"O6��3U���U��+�)��(Jf"Oz��6�L�q.�R2jS�<��lB�"O<� �ˉf�����_<Olʙqu"OHͰ��^�!]��A�O�WU��8b"O���KA7^�D!{���yL�{�"O�������I��� t u� "Ob�q o5$f԰p���3Q���!"Or1ɐH
Hkt��H��(8)�"O^�X��(� \���߂H�P�p"O���Ӥԃ
���b��;�])�"O>���Q�d@jb7�ι�"O�X�u�]��R����6ZR��%"Ol1�I��mF|:$@�?)5((�D"O�1���Ko��i �� L��r"Oʌ���C��qtB&U3��C@"O� 	4�ΐ��HC*�<+� "O�Ո�Gȝy�j���"�(�"O�b�@_��\s6É�X��"O@Ԃ��؞^��I��@Ծ.{H�j�"OL�h ��n?�EAq�ؑt�<�"O9�cC;o���kGiI�SϏ7�y�lƀN�F�R�.�w�&Q c�	3�y�J�O�����p%����y",��P;d�C6��+>��81�\��yr�ڂJM(%��hW*.���#�yr��c i�tL:&��[M��y��E��i�0I����V�5�y"R��a��1�,[VK��y��	5�,�A�����S�*�"�y�j\�r��� �֑jt݁P	��y�W w��!DB8�4��t��y��xD챊pY���B¿�y���;n#��uD�B����ə��yc���N8�sɊ�4����H���yR&��XS��ɥx��X"�
�.�ybG��U�	A�Ȝ�q�������y£�3F��6g޺j^6��G�\��y���!�B���Yz��Kt����y���
'4��9��ă#�X
'Ǜ:�y����Oؠ$p�@V���.C䉔&�`)�+�5�l��'�2*LC䉢��	���na*��v�.'o&C��%U�R����L�>� y
a�/B`�C��o��4�7�0f9��MT�-�C�2u�Z��fJA��>�2��
ԈC�I	@9�a��� _T�eqwoU�hjC�ɨh$����CY@u�	C@%�JC�	*ڬh��̄V�)��f�-1AzB�I0]f�pcNζ��Aqa޹8t�B䉕g��h�u�� ��'�F��B䉆d��m@-�0&;��*R���FhB�	$0�j��_=<�����Z�.��B�I�\�b5ś%3uP�R ��QrB����T�DԹ�
d�Ն˵g2B�	�^��s���Aw�]�S��,NfC�I�#�|E�`�QI���r��LKdC�)� 48���I���<`GH�x#���F"O��[�S�p,p�sf�"O,���A��s=��1#O���<#b"O�U9'��LJ6��m	(p�]HE"O��'�%2Z�B���4h�h�"O���G�7.`���+�ue���"O6!�ChL���p�2�ӛdH��3�"OPe˲$�8�xk3O��Vf�|��"O�	�-�<6�$K��˄d2J��Q"OH ��l�9���qI�(��r"O�x��
<X��a�S/7"
q"O�8"4	A�
�E�r@�p<�"O�u��KQ�z� �0oK%>h �"OpBw��}��0v'V�>�d�I�"OP�!�٭��zs	W$NШ�ӗ"O^`���T�^�LI�Gg'���z�"O�xÀH�W���{F��*3�qiw"O����#�)m`|#��ǣw.����"OBqI�j@5��q�n-%�Q8t"OB��Pb�X��Ǌ�;�h�p"O�Ah`�G�,�~P�ղIW�Z��+D�$����z޼��a��h����r(4D����#y�4��*��M�G�1D�LH�$L�永��KU�kx����2D�t��GRk`ʡU�.����1D����9TܲQ���Q�'ZL�$�5D���a%��H��蓲��?x��%��3D���UJT(RN����>,3�iYN?D� z0��9g@-	u���)϶��.8D��;Cҷl"��Z�BO�{U<085�6D��I�K�o��뒠I�J^Բ'�*D�����9p�f�8w���k�4@���:D�Dkv�ża��L��&N"W�*@��l:D�PWkƐ5iB��I Lʶ|�d�7D�ȳ���������b���f�4D�dp&T�ݬ�#�
H<3G`�W�3D����fD�A����F�3�0�R '0D�İ��)o3��:PoI}h��&�/D���R�ƈw���ဩܸ8g�1�"D�X5,�<H �Q'����"�=D��	6'�4*m9E@��9BE(:D��:P ղ#Z0�&O�C���R��+D�@s".�ޭ���:D��qu+D��I�A�n�v�ҎJ~1dtQ�x�<)Eh�1�r��v��3�A�AT�<Y��1]H�0$gФ]�,`���P�<��
K�����F�9����U	M�IG���O��ĢD#X���؂��'�٫�'��٪�I�"pD
�+#�'�0��'���B��!2���a�"�`p*�'��4���[ [���x�l	��j0��'/��˧iW&��8��J��pqk�'G^Ur��׺�y�$�d	[�-V�<����+[ 6�*��P;ađ� �MD{�'��e�!Ʌ#$�U�n�!��;�'����@�? 9z|��U�	��\��'Ǆ\�r�ġc�LUH��
�/L��
�'�>m����Hd��5���
�'aH�+��H�6p��jskI���%�
�'�9C�D/��sC.��<��u��'�9�'�B�C}2�{�n۶��	�'M�����h�BHH��Ӆ	�R=:�'L�@�A+�0�2M�_��
�'���s	F���UR4H�"(L�I���� Z��͗�:nj����82b1�"O�9�-��u�Tri
(6.���e"O@]���^dj吀H�^!Z��
�'��4�'!�\��H� �8�&EB�b�'ZZ�1WlF~UX�P���x���'d�T9�Igtx����n�N�
�'�B�heGWp}��-݋?�LR	�'��R-D57d]#�M�������'Ț%����6Hp�Ѳ¤��� ��'��0�W�����D���I�
�'}�	V�ֽ��x����!]�z�H>)���?aÓ0���4�� �*�A�,O0g�Ȝ�ȓ!�8��:#x#��w�p��g�����:�t�
�'�wotY��)��'�]M��Y���jkpY��j�0����Ȱ�qଇ�J�d��ȓYMrm��;�|�'mG�=����6��t!g�4	�%M*�he�?��h=ڹs��3 L<��RG�9${����%^���Q����@E�33��ȓ�4��R ��0pJɢf��PMX��T5�8󆤇�]&��2d�-<!�Z�Fa(đ&G�!F��rj��p"OQ��D�G� �*m�X)��"O���b7�J�J��I�D�D��"O>�a��ƈm=�E����hdB��"O���"�<R8�C5X�]��$-�y�H��8��ȋI�4a%��c���yd\�ӂ}Å��{�☚�̛2�yҏJ=T����$���z�N�y�a+{b�h)�fP�N�8�k�����yB��?l��	��G�y��M�E�գ�yr�ƌ&�4��d��_�"� �� �yB��.�6L���0T5���*E��yB�D;B�6m�1f�*G�8
��1�ybCG&z��� ;7,�lbGɏ��y��[3-��ɐ'�U�.�fUWJ�yr���Lo|`�!(DS��)�y�k�&u�@@"/�x(�"���2�y�C#�P���36	��ι�y�`f�%V">����3π�y�fH�<������ߌ��اͅ�y����R ���,��s�g�P��y��lLu����sSf�����y���:|� l�4�,c%̨(�k�<�yBeQ�?f�
�πg���3��yR�\:=��5G��)�ÍР�yr*�!����M�3C���Q���y%lq�q����8f]�P��y��,18�j��ڃE���K ��(�yRd�0����BO,E��A #��yr��)�vlAԎ�6�Z��2�J�yb�E�K�Hj��X�YR�R�M��y҇;'��� Y-�(q����y��@�N:���a�B �\%�����y��m�ډ��9 δqiu(Q,�y�a�D�i�扐p�P�񴥈.�y�o[��A�C)�Y�ۜA�!��^(�Ա�SC$U<���!D�"�!�D�t2����cO�t:��kԠ�<H�!��@*и���Б`P���t�!�Y_|IHdd�T�n�)C ��M�!��F�����&�]�P|@��f�]�l�!�D� :f̀PKġoz�K�ė=(�!�� x@S��ʃh����s���?�up "O�P����@��U�D��O�X��p"O"i�֋D������d�8b�:X"O��b�+�!0N�=%-_�8X���e"O.�HbG����qZFA	�K�	&"O�D�!�*Q��B�ODM��CC"O�L�b��79������7˂m��"OVأ�Ǖ
�$�{����.�@���"O�����?yt�X�ϰ��L��"OBXY�MF��6 k%�ߥ1�6�i�"O~ɰ�!sX��1˜.l��py�"O��آ/�,����wD%7�r���"O΅���F?�J͋򄊴Q|(��E"O t����lB9#�2��ыG"O�3�-X�})���u���x�����"O��BR���p�
#�Ka��Xx"OvX���4V��h�灎�}�Ha"O6�&�Ιec� C�@	�wd�AiV"O����e�U��u����LM�["O���oܫ]��A���IJ�8�"O�%�q��� V�`�WnW�y�ؑ�"Oj����%�u��-�]��p
T"O����2d㾕@�
ð8�3"O��*0Nn��*u/[,I��S "Oȼ��n�q����.ךT���"OZ�z��P, @�3̈́�4��q�p"O��S���)kT1�V��F��0��"O�P����&
o����K0���"O*�W/J�zBx�t�L�r1�)� "Obv��,ԊaT�H5,���r"O��)ѯ��,�H\F皕9�"O��;���Ao�XV�Y0?N	�"O�|���'?�"Y�"�-l��(��"O��*G��Y��g�g�d��e"Oby�$]3)���Tui��H�"OZ��S�
Z��
"a��5��"O6tqŢ�Qh�A�.��^ur&"O�za�5�8�P���^��+�"O�l��I�)1є K�?`;�"O�@�3�,,n��v��=!V~p�$"Ox���$��co��O�I��T��"O� �0)��0�
p!��%h�"O��b��#A�x;�MJ.R��0�g"OF�p�CV�S��PW�+{���s2"O��Q�h�'\Hɢ ��~�ƉҠ"O�%��N�f��r��J7Um���t"Oj��w���s��Ȳp�Ѱ����q"O2��,��8��X��"O�yk�B�t�l�zU"� ���+3"OX9����h�d��QW��ڇ"O���P+��f�pyQ�승&�j�kV"O�m�FMʅF��q�Qj��!�`�2�"O Dl�'F�T�i�HKw&ƹ��"Ohq1D�$�j�۷�%H@�"O�P0ŁT/P���{�<�JL�c"O��� R;"@!K!�F�54	2�"OP�a(ܛT��r(�/t�1�"O��` I^�)�|�B��M��"O�m���82t�;WE�n��Av"O�%RB��f���"�D�9���T"O��Ď��(��܂acؚl ��Q"O�����ψH���a\u11"O �p��*��@r�߈8�8@Z`"ObyJ2��'Q2��@�I �N���"O� ��2@�00�8h�o�}�x�""O���KG}JJi���7LČ�`"O���q@Z6� ����-l�s�"Ot�J���6O��"Q,1I���v"O�!р ��N�<9���+%��	�"O��TK.��I�G-(� "Olؑ��V�CeX��u�w0y�#"O�����T+�1����(�i�"Od(��ڠ/&4�!��G��S"O�,��C��� :P쐘)^�xq"O�-� �:Kbč"Eʃ�2����%"ORy���>;� ���:�	:�"Ob�SiV�5fxDfJ��U[�"O����P �`�0f��3�:�hR"O�8@1c;��H���,'��aB"O��UH\L��أ�Gni�"O���wjN&y\J��A,<�b��u"OR�٥��e���"��÷F�m�q"O�qAlO���0W�V�赳D"O�`��W�{_�*�g(^Zx!�"O������|�F�Q�'V���"O�A�hӭMհ؁���-�l�x%"O�<hV�L�*vZ�RS���y�>i�"O��H�C�7(���QbOV�R7Z}s�"O̹Ad%Z)$=D��&�	�g�)�6"O���2c:W>H��� �|�.\y�"O|�u��
x�)���D�6�t"O����!|y����X#!Ʈ��"Od��%�@�|�LyC�� s��܂r"O��%�A}�Q:�kۄwq�H��"O����(D�,l��`���3(fJ���"O�E��I%
>Դ���W�]O%-�!򤞓D��10V��"�:,#d�
%$v!�d��=>Ь���� -��p2��+!��`C��p���ު�z�	�&�!��X�2���юyRS�f�!�ɓbK�}iw�;+��� ���s�!� ���k���D�Є�+h�!�dt����^.�x��C�|d!�N%z������VDx��!R�X�!�I�J B�`��qIj4[ ��;�!�$��? K	�CʰH�
�y12l��'^$�s� U�!�6��w�)��'RUY�/�D��af��	|�0U8�'U�-� `C4y��p[��l�
I��'.�qdۥ6^�y�DjU��2��' ����H=j���!��Y�&Hq�'4P�s���X/����~�L���'5�����k�4l���H�H�Ź
�'0J��U?��}�`2�qs�'�8HCSMؗc-z�[d&6��m��'�&)�CcT�8��d:'�O�0/$i �'k@h��!�@��8�Z�-�t,�
�'g��Vj�<i�����M_�-<�10
�'R�%p��I�k6�h��>'�bu#
�'�L�����?�0 ���2���	�'HRS�>9�|1 ��2&'�(9�'p��������q)Q?�����'���-/;�~�񇅴[��
�'w�A���5j���g�eW.d�	�'�ހ[qJ�[�|�{�1жp(�'�TX��#w챴�_�
ǆ���}�D��s���\�X|iW�p��p��_��h����1_Π	9P�q8@��S�? &�hZ>AB8�3B�D��*b"OT��#Џ�d��G��.�9;A"O*�� ��@���A���.c)����"O^ar��C��	z��	�=�"OZ�*��O���E�Д܀́t"O��9d=8��(��R����"Oި���F	|&�ץZ�gg���W"O�<ġ�/!��<���`Q�I��"Oܨ�b/K� f�$.]�b? ��"O�@��ATP���-Ns.Te�v"O��8�'
����`��?h�"O�� �$�h�U����*u"O@���%A8}�yS��C�T���R"OT(����B^(D`щ�J�"��"OҘ#q�	4;���b�%*�f�"Oj�H�[+�F"�*�#~�Z� W"O�m��ܢ�>��f :6a���V"O6�"��Z�la��O��U~ΑX�"O��3��7)�viq�o_ll����"OLh�%�S�c��"_�O��"O!ɥ��o��L��ؤ4��`f"O�(+g� -6ݨ�kF��e�v5��"O�a��"��f<E�n��pD)�"O��� �.̲�K�o\���Asw"O���C/����D��!S�l���"O��a� 4X���Y�.K6K�����"O�x��Ε���r���q�����"OE�V�&����퐧��l�W"O00����v�~��LG�g~@c�"O\�ze�W$)���b �L%0�bh��"O6-��E��⌒Pg/
�z�"O@TyBI�/�`A����=:>.���"Oj���)\:�wK՚:C
H�"O��3�Cz�Hb��hDԱQ"O���o�.#�R��`F��+)D-�'"O��`6l�)/#�=I0%X�H�1"�"Ob,{&F�?>�Us�nʵtPQ8�"OZr�Dl���X�d�"T$ @"O��3��2t\b�P֣_�""��C"O�l����#n|H���59r"O�U�u�Q�1��
���� 4Y�"OȍX6�%"ئ�҂���\�5"O|�.�,u��sjB4{^���"OJ�X��Ũ ���UK�y�Q�"Opm���s�KJ�L5(4᷂D��y�%W�2z`�U�ƈ-eB������yb�_�k���:�ML� ��52�AZ�y"B��$� iQ:f��fi�/�y�g
�"�M�!�D45O�Xhf-V#�y��0,������Ҡ=>v��"�<�yR��x��!w��E8R�B]��y�N������`�/fb��%����y�f����<�2�-j�Pq�m3�yRo�,Z��i��i�:4���lR��y⯕0N?,ht� �(�k!h-�y҆N��"�3����+�M�y�*�:S��P�ˌ���!���̚�ya͸
L^(���Á��JP�Z��y���`
 ����٩%�8�ZvE�yB��d����R/J%g�,ua���*�yb�F)6	2a��b�`Ecu���y��S+
��aY��S5`UK��<�ybO� ��󨔒.�=�%�y�͵ZuzEp�+�	�8z�I��y
�  ]�%iMF4l�j �4��4�4"O$U���8 vЩ�dQ�=u"�9%"O���3@�ZT�2)��A[0P"O��yvϵ�tH�1pP���c"OP1O5�����E8nj.��"O�TS���hH�L�AEDgziYU"O�E!#�FP|�|���I�N����"Op���ؿ{g�P�@jC��q�"Oh�X�e;z�M����r;�<t"O�}��n,Q Ï� T̲a"OH%���4�(4��:�r=qr"O���T͌3}nD�@��>f�"�y�*O&�KH(B������������',V�2o�0yf�����>���'�H-[��щl�r���䐦)���'�,�E��*��3�b*'��P#�'^�$�T�8w�:5LD7T,�qI
�'��ҥT�E��b�K$I����	�'%�ЗL�<�|��Rc\3Mj��'c  � -ƃ1�bY��W⎜��'Z�A��w9�L�P�8Cn�$K
�' ����
��H��	:)�`Y+�'��+%O߉!���q"�$q�.�H�R�)����0b����'�phh8�I���y�ᘱ,>�ː��lV<�D�ɮ�y�F޻D����*�Q��.�yr��iS��	Ca]� R��J��yr$I�Q
Ulҧz��0#����yD�87� �(i^qՂ9K,��y���7)�����G+a|<�I��6��'1ў�O5�)�	��m޴�̓�R�4H��'�� ��^/H�TDԸ�n��'��թ���2�&x��˕<�6e@�'�F��gh�l5{c�ٰ!Zf���'x\Zr����b4s|���'��Ȅ Y$^?T}C2�~b,[�'Z48"#�;�<���\"?��
�'S�B�S�����]��b B�'�I���Ѷi�Px��Q!�d!R�'a�"�Ù<;ζ-��9i����'�ʄ`�=1��p��Fȫdf!��'v�9@�I�:x�sQG�<؊���'+"��F�#C�ܨ��Ê�T�diX�'��0��V�]�F��զ��x8$�{�'XL�� 5T^D�w& r�L��'�&��EA��0<j\�f!Zg�l|(�'���y�g_%
��S���oF�iQ�'�pq�V�\g���c�	r�Te��'��T�	/_�hP�O]e�ⱈ�'h.�2u,�Z��eZ#�:4$�̡�'>%�Q�6k����G�b�'��M)��LBb����H�����' 4z�ǃ�=��i�b�F�,Ap�c�'OL=3��	�ԅx��Z�#��$��'µ��!�CȰXq�@=�L��
�'��d��o٘� X�t�7{vq 	�'�� ��ְ:�2�#�LX)/�<	�'&6�T�<}��98��ӛm>J}ZM>���0=��lIp�.��j�*y�X�p��f�<a�
 4�p*���'Tt����Xl�<9�c�@V4��tnS`X2ype�S�<鲂V�S �$��2ux��O�<	�!N8k���"N�5�I���L�<y5�S�|N����*C+!θ[�@S�<� ��@�P�-����s��u΂Q
�'�ў"~z *˰J�����n�] �����&�y��ɽV�D��D�"�&�S�Ȉ�yR!�0 h���@��~E�gN��y�H!w��5���l�� )PG@�y�h�OH�ȩІ�1�8���y��-)Dd�v���x���[���9�y��f�8��MoB�����C$�hO*��]^=
����ȥ ^�)�!���)�V���犎��=���s\!�D [� �b)�R���W-	s!����tZ�
9�,\3��(|O!��I>D���b��Ȁ9�J�ѡ��dL!�D�4�Rt��{��*
�!���8K Z�Ar,�A�L*'�	��!�d�&BUб�a4w��)CA_,f!�dƋ^s�#�����e����\)!��'vFxRTi�K�V������!���7�:`�.�+��a7�U�6.!�䆪>ptoԐP�*m�PAG�g!�Dҽ&����D�:��`C7�I!�$�	���Ked�~�H��!�dQ ubh�3�(�>�h1���o�!�d*��
�.�'C���� ܩ[�!���F��UCЉ7��A9Q�DxW!����	J���
�>�$�L�lR!�ď�A0a�G!@#^�P$괮P.B!�d4����b��)�x()��ʿ7=!�d.ZZ�uXS�̠$y�<��H\�$]!�$F�=�$}��
4��U��	� .e!��;�� P� :}U~-�e�H�IU!�$��Tb�)�)zK�-�+�U!��ϱl\��HҎ?>lrh:a4!�p�Qї3?��9WD�:����"O�@�B�<]�s����D�,�v"O\X��
y��(0*�:I��	d"Ot=�w���8y�+փ�>�RD�G"O<�@���zD �H\�k��P0"O@p1�	ˏG��	�IZ��`PP"O� �a�C�'�LC���Eƺ�#�"OZHsdcM.Қx���$�Z �"O����ԭy52F#x��4�G"O.  ��^:?�
Q1�E2+� ta�"O,9@r��%_o����cثI�L}�"O4�x�A݄,.�A@J�eȮ�A�"O�ر!�p�4K!�N	Z
%B"OX�q�WH;�y��ĕ�R�xA�"O�ۑCR�8�Xy�c��ܽF"O���T(#��K�X=[+��%"ODٰ�K�r��@��;M	�ؠc"O�x:��ޗ��;�d�gL3G"O�$�
ɋT��� ��`=�hB�"O�R�Å{�t�4��{.���"OZ�[��A
y�P`3�۫(½�U"O�Q!�MN�jt��Ú�'Qk�*O���'�K���,ocX)q(�,h�'��e"���)&�S�[�B1��')XWL�t�8�gT��iQ�'(T�H�/9<�:E��kQ>@FXhy�'kN���G'w�p�2dHE�3Q^TI�'~� ֋�T|q�t�!��͒�'����o��v.�Y��'t�9��'ZrC� �Y� � �l��#�t���'�b��5��;{%(l�-��e4����� AR��45��M�A"��=X"O�[q���V`k�˃!9�����"Op����?;K� x2�G�H��qIF"O�}��f�NLP�{�J¨4Lnt"O�a�ۣ$/�3�'�v��H�"O�h���rҨ�'G!~�z�"O�1��EW�4(\�ĦV-R�8{�"O<	���2���2"G��aߪy�5"O��
1�_)T�B��V/+�`�xa"O�l�D�7�up�凷?�ҍ�7"O��a&�ŸOj�<����!"Od��afء>U���Q%��()�"O[T`#T<�eh���(����"O��ѓ���TUZ&mKv~T�A�"OƍŨ�5F���"-N	&B��&"O�ah�Ā�T��z�,�1a9Xpc"O���>y�|���Y#['�iʁ"OX�y3��� DZ�8D.�j%xdp�"O����3UVT��5�V�}����"Oܙ�GH�(�X��kY��ʴ"OH��'�C���*�<0��[�"O䑐��8i�ͳFG�)�Uˆ"O2m�5�ъ~��9( h�U��U��"O�:�	�i>Ĩ�g�HQE"O\��W@B~�Zm�%2^Ya�"O4��`�׊ባn�4�Ȕ��"O�$CRO�ະ9r�S���	1"O�E��#��1  )GG 2���+�"O"CT��-��+� "�x�4"O�)8���D'Й: �6u?���"OH 7�ߎ9N|��@.`8�"O�8Rʄ,m��("�׿x��iA"Oҁk'Ճ6�Lh�')��Pk�"O�0����.t�F�{�lG�k�h�d"O��t�B1�(`ڦ̕�e��3"O�R��Ï6b-��ǻrG&��"O<����C�-?�DsRKޮ"V.9�"O������[Hz�y�i�z�Z�Z "O�-C��~��d�bi�U�|	�"O. `���.#J��[��*u� �W"On�ʂbЬJ�h%GTU<���"O��r�V�F����,Ķ�"�"O���!J\7W�Yjv�&{�,Ab�"O�<wWh8����4�*�G"OXX�'I,���PSc�h�B]r�"O��g�RG������֒��}�"OD��aM>D��Ub'B�+�bd��"O�u�fe�61��+�@�s�ٻ�"O�T	Hs@��n��6m ęW"O�(S㭝<[|����$s�="5"O���K��P8�`B6\�rd��"OQ��� �_��y�,�|��@�"O8�B`UI�\��!�Jl �g"O��)р�
�dq�"���!A��!�"O*����H>Ud�%iD	�54���"O.�͝ ex����3$��V"Oe0�l�U�	���lHd� "O��C��H���KPaH�n�t"OE)�!�pE��Y� Z�1Ӓ`	�"O�U�Ӯ��a��@eo;Z���c�"O8P���X(��ǭ�(u���S"O�5kR��4x�r��ᚦU��|I�"O�4� ��n���`$O��LM�T"O��KD��mS60S.ߔ �T���"O� vP�W��*a���.A<�r�k�"O��I���&��P�uΔ�	��r�"O�ƀ�<Jt�)��^2̺�"O�1TCI;o����еa��Q""O�⌡:��'�V�}W"Ov\bd���1�Q�I�/	�U(�"OP��b(�^ج��)�^�a�"Od!9����x�t|J3f�ZОy��"O�aAJ�*VM�m��	t�<�F"OziY�i.Y����2�, ��g"O�S&�J(vV�0�&��hޚ�"OZ�±��w�P�;��q�dT*�"Oʥ�`Ӵa�2�3#�4��Yɐ"O2�J F�$�z�a�<k;�	��"O��s� sa0����t!~�F"O~���'QV�C ���8�%"OH��b3^�ڔ�����mZ$"O~��)ɧ6�Z�b���:9�&�8"Ob<)���9�Tj�����"OHX�N+b�H�9�N�6d��9�"O�봀�	C�(�3��5H�(�p"O�1��/�H�萆G�4]��z"O�di��!D�4�P�,�"#�f�Qc"O���g�< �N� ��+��8�r"ObՂ�ıp�����d���"Od- �-�*gw<D�aƸxT�k�"O+�� L��v`��MG�Aä�~�<�Մ�w)bM�-�p���A��{�<y�"E?V��&�^:�M��@\x�<���ouj����U ����f]t�<iåX�4%<����E}��GNz�<q�#I�Q�L��!��5����Q�<�A�$2�P<8�fC9H>]�eo�R�<�*Q�MZ�͉�J�)S����R�<�ǫ&M$neC�e��p���Ѹe�<������#�c�@����g�H�<ـ(�3Sj��*��F3_v*��U�AB�<APB c�rp�p��?M�t�R�3D���@�Z�td<{���ۂ,3D���f�1(^���1��q尿BG4D��P��g�f,�c�Qvs���J1D�@Kg!K�<x��͐'���
<D��2�هz��$��E�2:�T��AO9D��7���@ny��C5An�y�6D�`TV�V���M�T$"%�3D�,@��*���Ap��$�D��� 2D���3�H�Q�R���ԧj���d0D���A�˼�zĉgCζG�0)!".D�4�g�P [|�$N-��48�!D�<�.�l�n�+7�Ps�<�"/!D�0Y�C˥�0�O�4*���o!D�`�T��'�.��G��^�"�r��=D�� u�H�.S��@#M  N�M���6D���C�	�*�;�o
�+��}끮4D�l��)ݏ/���ԍ� �u�Ѡ2D��K�+Z:Y�~l��հ|DvZ��:D�p��j�&��!�d��f�KWI.D�����3cVqSD	^��r�h�,,D�(�惍�Xf5!&bPR���`	,D���'��Y���'d6E��?D�ēF�F�x[1˚�$S�e*D�X�5$. >� 
��[$!�p�C�D3D�,Cc���\�cb.��|�lD�v�&D���Y$i�L�*����f�nPC&D�� (e;2CT5?9")�0���m�&�0w"O�0����Z�T5 Х�	N�r���"O|�R��8m�@P+�� �&���Q"O�9��ĵ9�T�;ve2u� !��"O0���Do��B�N6�0`�c"O
�@�'F8�A���(��p"O�	q�܊y���Vn� ��a�"Op9��U}pT���#W�a�j� "O�ӷ���ҩab.A�nّ󛟴��I ƕqAmĞ]2�ÇV�n����$�<�&�%��h{W�׿-�,��S�<�B'ǧvȦ� �':�<0�Ǉ�i�<�#�ֳZ�Z�BC<@�A�B�Iz�<i@������/;b9"��W/�w���'�9�R�~�$K�2:0B ��'��!�k5G��;���+�BQ��'8��#Q!�%p�n���a*TlrQ��'	-���(�$<�v�\N"|��'�<�vK�
X
��ɵ��+(rZpX���0��O�r< r/C�Q8=K4�	�DXC�I)gl�:��Ə(.*%сg9?����xCJi �͔C���{�zC�I�@M�5c5�Źvn�ʐ�Ϣ�P�>�����d��k��ο����n�z��B�I�{d��Z�%ΈYO�e��װ{���	�HO�>����D� }���"� ,`�<<O�"<����g�q균]��|E�iOo�'�ax"g϶c����R�qn.%�$*-��	i���Ogr��@��">�t���#��3a���'QRx�V��{��L#$J^�'X!@	�'��D��+]V3��
q��>m�<��'z�6n��_@0�0�R��D�
�eF��y���9�(6�D}snp��e^��y�%L�M���@OR�|��4���Z��'~a{�EK=]D�ˣ��h�%���@����m�'D>�R&��.eG$u�4'צ1�2��5D�����Q��X��lJcB�Xz%�3D��Y�'�p8�=�W�̡ES����0D�ģ���81mz$���'%$�� �,D����)�����r�«�H��p.D��@��۱;�|}9�O 'B0B��w�.D�X��¬~�~@!c�~�"�� �,D����+�f6�i"^.�KH�\��R[��؊!� ����gK�hI�̈�%.�OX!&��㱣I'Fz���c�q"���j)O0�=�pፐ�x0c�ځG���Cy�<����$��L�F̨��q�q~��)�'g|�2��������ȝ(�@��{b�"���
�I�f��-p�8��>)�0Z�A�R*;(��d)���>���>y��>OAk�MP?40"eP�_�Z�z�p��GT�<�"I_E�<��c���������x�%�4J�:������y�����'C�z",ؙx�ZL:�c��sD�30ƈ$�y2^�����C�j��t�'�ܑ�?K��O?E�%`)m��sD�5!#�+tn�i̓�hO1��$k���62H\�ˉL��a+������<�vÔ'G?x�x� ��	V�a��Y[�	@?ٌ{�$�D��d�lK�.�|��r�J&i!�D�,l��)�3K��	���BCL�q�!�-1�y`d߼F�̙�b��`�!��	^P�`c��"������'�ў�>��!%�1O��Q�܉*����.D���R��{�䀊��^�t���G.�d%�O� ��t��5�9Z7b*Y
P�*��'�J�̓~�Da���:\��h����87��l�ȓ:7��F����͈'���_�0@���3O�����OL%3UC�9cZ� 8&��a�E�	ӓ��'HZ��a
�$ͤ�Y��P�Q�<ܚ%�On�=E�T���^׮�V�[	���t����>��O��0��Rx
�� 9 ��"O����H!"�:�H�J(n�ș���N���	*A���PMػ`���Ӌ�(:i!���?���ߒ
�hd��i:,P!�	�G�� 1,�v�D̂�ə�NE!��D���!�6R����N� 9!�D�+{r�t�m�(	re&	�/!�ĝ51��4�7j�${pMH��,d!�$�9:N��p%��!4e��S��^Zў,Fy�T?�`w� Q�|0X��f��Ep�&)D���O!u�`xg E�>0�aZ"��O(�=E�$��X0H��A
���+��h!a��OD��V1h!�� �@d���"O\ �� �P(�5�բeOB��6"O��Pq��yΈQ���m����"O�Ê�?	���!c#�J�&H�@"OL�tC�<q`!9�7��`"O���O\'N�~�£!�B	���G��O���I� e�tѬ��i.AWMɬW�!�đ;]�-��X?� 	�B��C"!�F�D1a J����+M�N�	_y��|ʟ�Ɂd�r	�1c$w_�1�"LӚX�B䉉Et�0R�Q�P��]Kஏ,BQd��R�xY��T�xF��%X@���	O?�vh�?<"i�u*5)�F���*�@�<� ��M=B��2bX�(��R�'(��%E�O���s �*L>8���^<8�	�'D�a$ �}s4��͏#9�-:)O�Q��4].��D���}�'���'DB"$����b�1����'}�@k`���R��qA��%6����d�;�0<��-1_�]���v�(��2b�|�<Y�eõ!�lu��i�>G@] ��SQ}�X� �0���&����	b����,�vdO78Ąȓ,��� �i�0	��V暸Y}�H`+Oh|Ez��M�~��\�D	���������3!�D�T��SF��3 ��AӠ�4c�1Ob��$Φ��ؑ��l�Vo[�+qOP�d0��f�4Zrl+�͐9R;�(	���y~���+�I�Ө\�ʋOS��P�g� ��4��'�& R�C-��i�q�k��a����~����[��8�雁�6e
=�y�,E�y��M�@��S��Գ��œ��O8�~����=�R�,�K�u���s�<)�/�/^��x���;�j��0��>�����g��:��E���4C�����~���6M41OB�J1Iғ*���`���^���9�X�X&�H�� /m����L�5�@z�d^)6�O�<̓����O��S'� ��3�(G�k�n���'�a�^���s� ��>zErv��(�p>�L<��&��3���Y���	 �ؽ��O�<�$"�=s��i�R�Њ�iR$�R�'fўʧ#P�\Te��V�"i���^�"�̓��?��F�O�4,PԦ�<��+s	��hO?�	�X�2aB���"~M3��]�&���d9}��� �ڸ8r�O�L�4��d�EzB�ɲwZ8���%ڼK��h��M+O���d~�2�4+ӄq��U����
+��˓F7��<�&��>\+�,s&%�	nR5;Vnj�'������ �]�g�&��-���+f��se"OD�GC-=>,�K�&�G
9ї�Idx�|���*=+��L��T��>D�X2lS8��[c�-O�Pa�.=D����Z�:?h��Z�\;J	i��9D�� CM� ܳ@@]B��U�Ҏ8D�DI�i�/tyx2P��{<���H5D�L��	íhb:�[��ܪRk�Q;�#9D�|ca&0"�K�4�v�A3�#D��2tj�f� t�ǁ�r��4qp,$D����Ǖ&��m����ztB��@�%D�X���H�P��I�qJ9s6i7D��1� ���Q���=�E٥�(D���	ЉLzeB����(�D��� 'D���$��:�(dU+��K5�:�#D�|*F�ϛ+.���g�t/�u���%D�,2�	�� 6,��"��0v/%D�!�g�8=^(kA��jYn���0D�H�+S9Z$p�{����р/D� ���L� �����m�j��6�'D�� 	1M��-� �Mn4��3D���`��j�=�Q�M�8��7�4D��i��I�}X	#�(Ψ��mx��>D�PBޛ$��� $��#��8�a)D���U9@9�]q@�!k*��0�#D�4�1�pU<����]+R�����f#D��BqB���"���eߦThr��h>D�:b�N�z�\�Ӫ�zD��G;D�XX���h���4���k8D�H���D���2���y�B�P$8D�����T:�bx��%R9#[RQ�M7D������.a���ӧϮ�l�u:D���*�d���3�N_�jq058D�Թ�Y�l>�]����/b�R�C#D�0�#� =�
�G�?��7B�ɔ]7z`��2|�i��D���B�ɓm�� #5��8S����si@7<�NB��&NV�iq���YRy�ς'JD~C�	9A���RRA\K�(��#�%�^C�Ɍy�T4R4�kB\a&f�g>jB��=�� �E_)V�F����]�$�H">�W��'Ѫ�S5
�r�.�S`���<%n��I@��C���z0��p��E�<���̉#S���O��� ��AF}�<����c(H�J��Q�Z[�@�oSz�<	��5k�,���ǋkj�ċ��S�<��'�7i�=����-��
 J�I�<A��1C������Ǹ�T4��L�<�.Υ����O�
�4�HL�<�w���dd��$C��U��Aa�<q�OV3
R��v*Z�+s�`3�CYc�<I��۩RT
�;�K��u�n(�w��_�<Qt��.3�����2Y����bL�<�3I���c�@�-:�:!ig&Dc�<�4d�H�L���g���=1��g�<!�Aɋi���ӄ��96Rj����X�<	�\2�;3a���R�O�]�<YtbS�,�,��BY�:����N�T�<���N+���焋7��i�,R}�<��J	��(S�I�T d9�"�B�<1���5Hn��(��N�� �O�<ѴB:����Ǜn;ڍѵ��{�<1�ݙy������f%�2��I�<�%˥D�2���(I�P�0T͂I�<9�#�C�LLj1�`��/�s�<� ډ�s��jsF)( 
��o�0|�""O�	�F�G�^�D��V)[V�J�8""Oʤť�+!�T1�J&\�j�@w"O8��ǍK�1��pAAf�^���p"OT��,$�|L¢웣t�~���"O��5h�N}�yZ��i�@� r"O��R�$��!]t�7`��ȁ�g"O��Q;�LDa� �fq&0�E"OI���U5���E�؍j��B@"O���E$I�>8�Ba	�D40�"O:9�O�W��ȋ�Ǐ3D���"O�s�f˞P��!�&,(� �Kp"OP�q4�y1���)C�D��"O��r� �rl��Pfg֥'|Z�٣"Ov��@D�#at�^f}p�"O������*����l�J��Q�"O��
� J�=ߠ "Ҍ�'r
�q��"O�X#Ѧ��cƔ�@u��Tɲ��"O�hR�
��>�6�چʚK�(�B"O�p�CǶ$�|9�iCw	�Y[�"Oni�E'����"1�AT��"O.��w���aږ���&ҫ�X��"O������LhԼ�w�C�Y�(�S"ON驅�H)Dy@1B$\:¹�"Ox�Ä���
?���E�4T8�br"O��BL+.,zT��&(ʑ�iU�<!"f�,h�����i�6] E�Q�ɫ$Иe�P�'�`�C�J�o�5�d�#��s
��$ꔘ.�X��``A:�l��,V������xW�f���)��ىz��D�X���O���̟�:��83���"��N~�@ Ε�Dh����yb���d<��q�^�&�p��FU�y⃊ =�-+ˁG��S�]?x�z�ΉR���WfR p3`B�IL[�fG��H�F?`o
퀷"&?	��ďx��<�Q/%ON��f�ފD;֍���Uf6�yw�'� �b5f�ts�f �P��$��m�1H�w(<�p�֛SX��R�@�|+���4,L�'�*���6^���}Be�U�8;���
������.�H�<����\v4�y �/[3Z-ɥ��<�%�C���Ђu�5}���T4��agF�M�bWC%!��A?	��Y�ŊJj���N�[9�I���⣭��k��xBiB�+R�=�uƆ�H	�-�#���p?�CmD$X�<S�&1S�X��R��yYѬB���x�K7`{d�CGY�A�4�
%�2��O�	�k����O�\�R�!F4�����J�bub[�'Ylq���l�h�F̻eS�q��'�
mBD�PM#Z����RA@���'���Y!z�D����yR��-q�-�D���R,�䘁�yrN�o��L(����E��JQ�yb�ďd}@�Cc(��e^p)�&���y"�)s�(�&���f���0�$ ��4OH���B�8��0}ӢB+u�Zy��V��ʣ?)�
��c?�8��N� 6�
a��)i3>��0m�H���Q�lh���Zz�3�I�T�M��f:Z�P2ȍ+*��=�x ��j��S��
K&�j�H�!
p�l��k<4��E\8�Z�Pg�F؟l۠�3!@���͟�_ D9�B�;}���>\�N�B���m��!��
P����[��)�9��Y0E��4�H����[��~�`�$�����81���@&��*4J,J֍�5<�HՀ3�ںhj	ʂ�#f��)ڧ�-��Ñ�Y
�͑S� ��TE}��m0��� Y\�''�\����דo��Z��Q,`�9Yr_���F(�-@e��i��~�?!*�x���իL�!�OP?��, �X���Xr'-}�����w��}a�!T�kx�[��M"\�$@1&f0Vy���'"D�2i̹W� ���ٴ9��M�H�iG�oN��A�jX6�iWj��"v,	��� x\��E�B]J�����Y>����'78��-�SlB1��;ʴ�� �T.at�p���#��d�Ӭ[��D�FQ��}2eH^�F4�C+R�=���I6e�F�'��[$��:�&�˓�Z^��MӃ�a�䘘%v��#dɍ�Q��1I� �h�A����'(<J���'���Q��Q19�H\٬O^5/�.��݁bJ&�H�4���hf����OV�@q����@L8lB�Q@�:��R����d���	�@�� s ��V�����'O��gD�jG�ϸ'|d11�Kh���K��@�'D<|Y��P_~�R
�o��c�NC�!{�a@�eWmX�D���:D���C�051�-"U�,<O@��P��33;�92�O$ ��=Lx���V7p�
��R"O��!�6c�iP�.M(2�LAD�|���)7�|4	�k�O��m�4��Z%��ְ}	��'�L ����
,0����i���c�H��o��"��@2z�舦��<���X@\A�4d s���C?�~����:|	\�#+�D��ţ`+<2�1��@�J�-k���>,����'�vY��I./*�MrQ��eD ��dT� �xE�rfɮ/(�UJ!A� gF�L8�`o��1�(�a<F�̄ȓ�M��»��ʠ�8D�9yѠ^�?�>��Q
�!H������)ԟ@��矈f�D�X�0��Z>O
B�sci)D���f=$�n�ӧCn��L��&�Hb��S�V={6�1�6(ȅ\oD��<q������	�D(dXpi�0�� z�[ J�p����m�0a��e�jQH��x:u"#kK(���fAь��٩'�ӧ2��ɴ�p���ɲ{��p!2�6�С�M�<��<��Q�}��XbKƷ�ĉ�-պ=����2*�ЌK�lթ^
�F�!KA�1��o��p?���Kz�����0_9ڄ)� �yz8��'��Xyv��C�����'�?��Cc-n����d(�[6o���&ւr�F���"OH�Rʎ�{\���f��1�H� 2�@,�����%؋Lg�sh�	%K�i^��yRoP@,D ��'J�B���B$8$ �����-04ˡ ��W̝�!P�.Q��@U� )�U�q�]�{��B%�
�~�Ȓ
쑟�[���	&���ˁc�*Tj���"�
����bI-/�d� *�Y����O ���%߈>�����+�.�h4��'Y ��Z���I�!���r��Ȳ�'��������J��.O_*	���z�t�J�k9+ .HX$o["fR0C�I y^ ���I}���#� >�b4�0��{���g��X;�9��'��G֜J���i�g̈́DP���� ��0?Q�NF?��xz>P��\e��*�,�5N_�Q/�cuo�7Ss���
ߓ@!�`:p2J^�=���Q�-D|HD�N I�i�8a����
8���Ù65��"�Wx�0B5f[��yR��'�zh���L����4π-�ybɇ'[�0��.K��b7 æ��>�
@fǃ}^Pa�r�zm*��b�=D���5D��N~����b�GH��0����XK�q��Gi(,�I�_�V"���'h�QA�PJ���
�,�(sF8t��ެ��'F��
$D	W#Ȋ��P�'�l��� �t2����A<�O��R��?Cvl��r��L�l���	/!v��Ǘ�,�����M�8Q��IY ALy`·:fEج�&K	a�!��(I�]���T�����*U����,;�T�"�4d�Z�ʅnT�O=2��g��6��a⍛Y�t��'�ԍ�E��uI^�!jߘ^)�i[U�݉X�lM�I������7��g�~���W.9P|� �D¯>LD8�?��I�h�����X���%!WjX�v<��b�l_�%�PO�p���I�4��|c��1�(h8!GH�;�@{�ˋ6��'Y��Sg6�\��D�"�$���'� T���[JX��*��Μ�H�%�'f�MG�,O A�a�+��ᲁ/�(+�`�i;�������[p�ʈ=��D!'?�}!�]��\��c@�#�� P��P��3�MUϨOxc���
��DޜU$��°`�96U�(���8S��9���/	���'V�]����ti@�d���G���ٳ��q2�)K�(K6���)ްv\�O�pڇ�ܖ��	�$����T/{�ӀY�6�dvtd�x���z��iV��`Gƴ#< �g�>�}:�΋�I�$)p*�3uVh��%eR5`견��O�� !���k��qy�OD�*fN���L��wf�Q��C/K�|�i7�<�J��>�'8�)$��>�	MWH`��!�� }��g")~���)�䦟�k@.��yPͣ��O+&3��O$��;ج��!m�?}�:��L�\d:�K�b����'�2�'�� k�i#s��\D@ѐ��w�1�F�7�y����6�!�)�d�US�a�=[J�^�:1pᨎ�*ڢ<���<�0p��	6*,�Ə���� >|�����b/\4"g	L���h�æ �zvE"s����.K�"�2d�Oq�`x�f�3f&�����;3pXQ"���ݘ;�0!��#�6�y"���G�҅���Rq*�	 J!C�
��5����.]Av�p�>�#��;����I5ue"�p�d�b�����7:�t�fDH���-b�%�!��z�'>��]%&\��S��0k�ν듀�n��Q2!bվ:���	=T�f��0!I� �u�3�8;�R�[Տ9��#2@�>�^w���(�'E@�'�K~R��!;�DH�5�!ya��+��=��fՠ&*��s�'�Q��`�H�x)	��E${粝�
�'�
Ajv�X�g�px�(˥uh2��N�bAF�4G�YB>����S*D>�H3�М�yR�W�kc���a6Q�²���y�h�]�8=�al�/��\:�%J�yB�˼P`(Y��ə���p���ė�y�@�a	�=�5Eωy�hy!$<�yk�4;f��%`÷w��C�O��y�
�h�ԽXA�Vnd|�襂E��yȬ{��m� �!aRd(j`�K�y�iڒY��Pe�:���V��y�J�ZL����D�HW���֩#�y�l�sԨ<:�":\X�f��y�ۻp��ȂV�U|����甾�y���Y�I�6f�;C��a�5E�4�y�\�&@B�&� t�buǪ�yBI��;��A�"{$����V��y�������"E�F��x���V��y"DK�j\�a��U#G�<98@o΢�y�
��#W�6L�+w��y��� ��xFѰ/�Ay�kT��yR@���ir���l?����H���d�+	���C�m�% ���G��yr#U.u/������� Δ4�y2eP�hRz���$Ƌ}C�d���y�鏄?:���-��%�0aٖ�y�΅w$�|12���l[83���y�&M*����e��Pb8�&*��yr,oR�rR���i�������y��	�Z.	"�`��=�E&�*�y�% }�p���(`S \0��E+�yRBT�J
��Ȁ�j�2��tiM��y�a���<c�䙞s�4)"h�:�y�NW;��1�+D/c� T[���yb/K�T�^��aոf�u+�H���y��g�5X�L�]t��cƝ�y"�.�FM[�bXU��u�%�ĳ�y��.���0VgA���1�e���y2@
d�Fe�W" <*��5*��y�� it���v���ԬI�kͼ�y�	�LC�0����|V�q`���y��:�~a�k�$r�F8q�T6�ybM��D�����k&|5����y҉���dy��� n�L@q��Y��yRȆ�}Z�r�g��]2׃���y��-�d�+�+e�	�vGՇ�y��
R��Qɢ�Y��$���6�y�꒣lc2q���m���tk��y"f�>%%.�pw�؆[~6�S�!�yBnY7aS*q�3�ګV���c�ˁ�y�
�4 ������U��T�ć	�y��W�_ ��f�x������yr�d�\�w퇦xȑa�A<�y�΋��(�P�1��f舂�ybF��lA�h*�C9vl�j�l?�y���= �(�ɑ�e��lxqm��y2��h��4�eДZ�������y
� �	H�
�&a���
����"O�鉃l@�8ZD<T��.-�*hy�"O|#�D�?	�8ppQĈ!�Z���"O|����
y*l����-�%��"O4��`ÙB�B���eS�nhj(�"O�H���
]L���C4[hv�"O����FSO�h����b'ș�V"O�5"���
*]���V�M1%~���"OX���@#T�`5g���
1��"O\8Q1@ߜc�j3���
�����"O��Rh�:x�܍���F�3=��{"O��TΉ�U?�|"r��<.�Ȳ"O�p��.k��Y[�E.z��J6"Oh��t*�0^pJd��k"��G"OJ��Ǯ��zm�����'����"O��!��"?���iD�T:6�Nut"O�y��Cմ+d��ط/\����"O�	:��Y�
�>��'��m�Dk�"O
� �,=�V�P���LEPR"Ox������	��Y+���"O���`�����C�}��p2"O��y���- F����AO#����"O.��o_-*axHBF�?�"A)u"O��Y�h(t6&Q��ƼQ��LcT"O($ZbN�p-XCV�3����"O�0r��!x��eږ�A�Y'`TW"Oƴ�@gF�&˴��A��"]��"Op��ˊR$�Aa0m��z"O�E�a�6C� �3̃�A�V�ps"OT� %��oo�1AT�{HP&"O���E���ۦ��W��:���`�x�2v���=V:.P��� <̠s����b������n�R��0,��j���#�����ŻS!.C�Izuz;�
lȒ�P�H4${�#>ac�`���i�-9��X[<+�[��;B��2�:C�����2�'�D P����m���=.�P�+2O�J�S�Or�a o�$g��	1O�=~~��h�'.Zx��	=hlmh���d3d���O���p���/�h�P�^���!�ݣh���A�3��	��	l�����'~Bi����u�)"�OT-2LЍP�
O���4��EP�j{�-����yD�@�U=
�q�LhbEk��Oc��Ӯ�xǨLI7"Oj�qT�n�ZL�&�-΂iC62ODe���D6n�`P�J�"~r�/�+|�Y�#6g�ZԊ@K�<�����6�|<"��y�(}�b�M~�2�"M�R��Z8�ě�F�z=�]Ѡ�E�j���r6�%�O�EAA��c p�)���B]ӀC���m� "7$����'�Z�0���YV؍a!�<��z�a0���\9�� �3.6���A�U��B�	���4l��j�֜��gؿWTB�:���
�G��h#�U�a�B��m����փ&M�x�!�g�C�I�P��)3�Y%R�p9��R-�C�	X�L�Î?>_`�1��F	i�C���P�U.%�>�"�~ �C�g� h�R�?�6����Šp�z��r�V�Q<�$��|�fەJ��	cA��18R=��D�'V.���Ei�]�*MaG%��5ĺ�ᄬ=L����M�pۃ��x�bM�K|�>�f��<HH4H�!h�S�r$�H]}�ʌC6��z��|J~�uN� ��Qɐ$Fm�f���Z�J!$�aS<<��a;�O��0dG�nk�%P�'W�$�9��>A�n�/}NZ(�0����t-5����/O�tEY�i��j��F�*)��B�	���p?�` �`c�y�w��z�`ɻ}�J1�)�5��`�L�Q ���wO����Ӗ �[���R�� 2;��|
��I�֘�@�A81�� ���A7���b�ZD�+bI�Ay�ː� vvYh��Id��ę.�r �VM�P(F��A]�#�D�7i�.�"��)��)��=$��2o��~\Xqb�N,��v��*-&���NGE؟D���i�@Bo̱d�9}2&A� � �i��h�9p�� iL�!P����)��l;�� A!�����R��~b&��\2b��q�V��\�2�Ӳ;�$9�F�8gּ��*��V2%�+O�>�Sl]�Kr�(�ߤK��ie�&�:�܍��W	@s�E�(;�Ф�=jTAY�#	9*l�D����	s>^�ha(���g�,���SQL��*���9"v0��'a����ԉ]j���	EV�O+��J�4�$]���߸�� �4kBi$IC!O̡�敢y���fZ{���C�`	iZ-�0��г�l����gܓ>�r��
�]Y�B˨Cܭ�Ɠ@��Ȩ1�A%z��	�_>*� �	���$� �'�ORɒ�ְ/ָ���E-��+��'Բ�� �(	��'�� ٥O�G(�hRQ�s��l��'��5K ��+|0`
QlC�$�N�J>�ß"�V�)�o<��R�C��b��XjS�|DZ�,&D���9~���D.��-:e�G�<j���A�M������#Pld�g�'NU+&�M�s$�I�+��>	$U	�?\�RBI!j�pP�j['_t�@0��%j�㒂�,��]���HX�(;&V�Kܞ��V�R�ܤe&"ʓPd(0V��Iޜ��6��Q�֬
��9z�G�$H:�m��6^ ��"O��R���C8fL��\O���A�*G�����b�6�<v�"~�	�1���E�w=d����~�C�	��yKU�Vk�fAc���1#>�������U bM�Fꗶ��;��?�=��œ/"j��مW1hDeC�l\P8�X8�M�0vM�i��K�,
� 0���F�g��-� ��p6!��N*���{$��r�n�3w�ă'1Q�4Pb�O)y�ԑSᓑ#�l-ʢ��1l�0I#H���C�	F��,2آx�:��A*�J<�p�� v���g�3}���'�r6���h>L8�skY.Mẍ)�'k��"��{��]�w���j�'���k��v2h���	46F�!l�.5�ά��J��6���2|<by�����P�CG�-��Ÿt.-Ø��2#>�;,�!x&��!��hp,eF{��L���G��&�,wDL�í�2x��D�=�yBm�7ߠ	� `�(dF���˜�y��	+9j}��az*��i�l��y�G��t9����bm;�/ʉ�y�V�Xhfl	��:�p�[V\=�y��We���ʆ�
�4А�奄�yb�԰AJ 0�mێ,udq@U��5�y2,��$q�,�PGC�4~���4���yIH�B<""�X�*�&��e2�yr"�*q��4��	/�VPD�8�y�b��]/I�íY2##ҁS�D&�y��d��a�4H
$����"��y��E;qu���M9S�*�Q�H�>�yc\&W�:l��3L;>1�9�y�c�1zv:x�NT;�Xb�K2�y��Y?��+�!��nP؀��1�y�fN�z]� �W�g� ]�Vf��y��۹;^R�J� ҢS��˧�7������Q[���d��Oe�
Š�>�ŪT�fC!�d�!����gT���x���=g�y ��Ѻ:�%���(r�Vy�Ӫ<��S���P�Z��DՊa�ݑ3�˨�~��܍eg6��Q�͌#�:ġ�n�YH��P�{"AFl���P;�uiR��29h	%� 1Ol!�A��������;z���&�Q�C"]Rr��)XQJ��רi ��� �
�ٳ�JR�3��i$Z;0����\<� �'�Н�����@%)P��,#-�>a�nԸ<����*�T���Tt؞��%�Hw���GU��ȑ+F%��ݢc��q2acŘ��z�h��]-80�Jw!�7DR�Sܧ�.�qPD��fYxv�E#/�Z��=���_��]U�o�<���M!e��ڟ�x`�΂p�\i 
b����f�3V�$�O(U�i,�3}
� �<�0�
	"���Ir�V�\���'�O!麈 ;Oh���
��~N�(����+�߅#Մ��:�t�$�N*BH�1E��PJ\h�C���OCa}��ȷ% uZ�i�5sr	�4M��6�X3�@Фs�(A�'���@�Ɉ6&
E*7i2j!�D��>	�&���{��Őc�F\�ѡ�V���IA�5�ph��5O2 'C0x�Y���I��|
1��! z�Yb�Cכ$:�)�D�J�E�Oq�^��3�'ud�p�T���D�m8#��D�.��T�ԟ�y��K�	��9B�(�Y"�@V�U=�T���T���B��QhHœ>��%Ȋ����ɹ)���P��<��0a��^K�t��/�	�n�I��D���T�'J�x�]�N��Lpb��>M��z��0.���댅%"z��I>w�U"$Vo�N8���Ѹe6T��qǛ�A�n���ͤ>��*_�:�&牶o$��H�����HR�)��B�K���o2lOBYh��	!���	$���t��-P7*Pa�O,�*C�ɩ�܍�goV���3��=��⟔�� �R*�?e˶ʰ;?~��4�;,��G� D��s�낚%��y95爜H���#D�̰������!F�&��Щ�)=D�(�C���F�>�+5bĕv ��(6�<D�H[��T�I���xB�r��q3S"8D�й�"TI�oD�S�R�y n8D�pZc"�G�d�b'F�� ��P��=D����M0��2f:��GP�7B�C䉜:|�1�qDEz�� dK�C䉥R����ߠp`�@�pȅ�DC����dㄼ>X�4��&տךC�	{��-��e��X�2��s�׾�.B䉏�x�86p^���i�[�B�	�^�|�6Ϟ�y�((���"��C�I�DYĕA�F�7;�r0��+*N�!�!V=e�RM�`�8[��+q"OZ�����<] t�IQ&5m�x��"O��;QE�g5��8��;/���"O2)#3���j�y�p�P,t�#�"O,�X��[��$��[����"Oȅ��.�],(�K ����'"Op���`�>���K�!��s�"O��S2�v>X�2��
�5
S"O 
�W�!fdc$�B�a�P�&"O�M�S�
4j���&.nLx�"O6�S
Y6�,A�kԌk�d�Ң"O(|X�"��pZ!�?ä��#"O� 2��	z��֫�t��"O�p�`��O��Px��ԷS��d�"O8%Û�~�j���l�`j��y��{��T��g�3�v�QJ���y��L�"dxQI` QZ��hA&[5�y�)T� U��'��Q)��H�៫�yb#R�L�dL:sc�!I՚(p'MH>�y�Ȑl�A�4��A�=+�
O(�y�)I�6e��"��*��u��iɨڈO*�%fM>'YXiC�e�)0&i��ґ]cXW)J�	�(U�B�*�ųZ�H�ge�(z�P������ӌ|$���_�v���gjE63���DX�_Z��`�mψ}�T�S�O�jXxV�#��)(�VC�P�p��g��]�IR��)�3��'[Z1X�̺0]��9��6]�*�e�'�¨Å����F7���҂����C��Q�9��i�I��-I�D�I>a�Y>UD�Ԧ�&�w � lf����X9Ml�(H<�G�I0r�a��gԝ���5L E��@5�ēj����j�a����3n���tL��M�Px��ýM��=ϓM�m�t+�W?�}&����.��v3\��S�.��H����O��a'�l�S�O�P��ݰ����e�շ,�� W/���'�a��aD�ȈW%R`���02����'#�H�P�'��?�L��{�0��4Vby'.�L�I�oh��*�n�#�?�1c�E�7R��Qu�Z�t����wJ�>��/�*��"}�Q��3<(����N�F�╬��Uz6��%YqO�?}B���k���A��Ҧ> R��ɲ�0|� u7� 8u��7��.{��S7�D׽�(O�O^�34Jވ�ʙ�Q
"hڊ��N<9��)�S"c&�Q�K, $>�{����}���������@�&����(�%����)5��i���'*9X�;fj�|�d%(1�*����I9c��Iȏ}���]��n����1O*ЊQ	�?��c�&�	o>�� ��TS�����95���¦�_�?鸴���T�~�a��EH0����-t�:�q��ly��'����p�	�P�?��`��)d��hH�d�3����׃�h�J(�Od�9S��/Z|9@ �6��|��h�qj�8��B�2�H��c�'�,���c?	T�͝����,��	P���c���rm��}�B䉪 C�P�&�'#m�m��.5��B�	�[�YybB[����獌�`֒B�	�^�zIk�횸V�ʰb�I�)mSpB䉵Rw��3 �ċH��������q�PB�	�t����&aǻN�P �	\�ndNB��(pT�0���Dy����DB�		=c2�%�ڐlq���&�u�B�I7W�P�`G@�H�J3jX]6\B�I'��@:#�ҝ~5V�Tl�""B�*����C�I	'����!� �.B䉩ΚU@��� .��Q�
�V  B��z7�}�'
��6� R��--��C�	�+�b䡡)�6wf�K4%�TRB�I)l��*�OA�R�Be`�0B�ɂL�2�
�3{�>A��DT��B�k��V�=�ba��F�,K'`�r�'��eӢ/?��ʓfO#���'�d ����3�i�;z�d��']Y��fn"� ���+<R�'�=[ӧ�#���R��̓����'�|����"Q� tMX
k
6hx�'YK§@h��� LёIa�U�Kz�<9!U�&��Tb�|J� ����y�<�+А�[��{_�]��D�M�<IV��#���.�Y�zQI��M�<�aG�* ��`M9/HR�����H�<	��A�Js\�
�<4�pmzc�BJ�<��*�o�:IB�荶Eg��aC���<Y�%�.[:H�rG1x�|��B�c�<�"��W����I��k���Q���W�<�!��@��m��`L�-�!9��X�<���7bP�Ds��^�j�$9rխ��<1C�Tw�&a� �Ī|��R׍|�<#�fCN%A�f��t���`�u�<ip��^����I���9@��r�<����g����b�C�|�$Uw�<a Bs�Xa����85�5!#�s�<��<������Z6H�D��J�<i���"G%ZS.J�QT�Q4�E�<�G�� �@%Ϯ?�@��a�A�<��H!3����k��XPQ�r��v�<yaw!��ҭDEe�pz�	�s�<��e�����I�;�������!���aUNH;B���p9f @��K�t�!��L\xp���M�	\O ���9m�!��X-n����6��.3�a�%8.�!�d��}N�m�U'�z�p����'o!�@�X��Mc�ʢ����DŻ/c!��Z/|8��e�J4���Bd��w�!�D٭Mմ����w&����ac�!�$ћ|:ܺ�/'�����
 P6!���/�:�����g�U����u5!�I)AP�ģ��E�J����!�� R0/q�$�;�Z�s��d$"O�8v熌3�q:NRE�P;"Ov���0)�A��B�<Z��y��"O�D�6�E�?�f�Q���#ZH��T"O��ӡ%��q��Xv�3"O\	!�H+H�ܬ�U�X8(���D"O�D�F&*rъRd%��M�<p��"O`UY�I���)
�J�e���jv"OX(p�ڤj$��1���B��4"O�Y": ���t�NX=�}�"O(�p�fҒ.R���#l���.y�"O��
S���2h����J28sl���"O,l�����
ٶ�KA끍K�.1S"O���Alɨq����r	� tY��f"O8��婓%�����4,.��a"O�x�0��en�ȋ��Ȓ@�p5A�"OH�Y�)��Bļ��6���,��I�"O8,ʓ��1R��KGI*�����"O81�D(\I��f�.��"OHTy�o����3�4b����"O��Z"�:G_X�3���<v"tI�"O&q�.Ѵ�^1B�a��}mx]	d"O��#�^;=	�p�F0y�x�"O�J��V ���g�'>�0$�@"O�<���O&n�� G��7�`t�T"ON�����h�)�C؟h/����"ON�Z� ��у�B9����"O�x�
��@��ׁE�{��*�"O�I�q���$��@����+���"OZ�`�I2>уƅ�Hj�L��"O��
��1ڼ��bփ8tH�X�"O&(q�@��Q��A� �^Z*E�"O@�s嗑<Mj]sc�D�Q&8��"O��BM��tsf���O�9<Ƒ�3"OX�:�-Ɓ!���$�Y�6"O���HՍ67�-K EZ�R�ZmC"O��+W���4(r��$�[� ���"O0qk�/
K�:U)�ES	9��`@�"O�eP ,7gW�a[w�J6"�){v"OB0�1A]�Htt��nD�&"O*A��$-">�h	��$O���"O^�۠��o����#A����"Ot��o�(u�����X6Rx�"O><�w]�	�$�M�"	K<�a"O�0�ĭ�:\�ys�Ѝd_��{""O^8�	"Eh�Z�W�$I�1��"O�EC�X/IO�� &�A�Z>&��"On:D���&1v�aR�-��`�G"O�����M"]�>���@G�qwd (�"O(U@	�=Z��J�W^��sr"O���'��3�*�ō߃vPEK�"O8	�"	� �ecS.I�w=N�;�"O(!qNJ2g�^I����.'4ܩ�"O
�Ѓ�S( ��`����"O�A7���I��=��y��7"O��*E�&.Ѣh�$H�]u�Y��"O��*�+�)�:�X���1F:�U��"O� ��
^Jz`���ۭy��#"O��G�B�bp�Zs���zS���"OU[A��!�d,�e*�,\<��Yd"O6D�0�ӹ`B*�x�	��*�~���"O�c�JA�K9�q�VoG+*F�)C"Oj̸��a��hb��V�t�@�'"O�͊���- ]�󡬇���ٚ�"O� 8�1��4X�\�$�μw����W"O�����eɺ���r�*�e"O�I�3 ����)S�ȊB�ڹ�S"O����GTf���x",L1^k��a�"O���r�I,��4\�4��"O�m�څj�<M��,�:>�4�U"Oi��e �U�v�آ+�9�N�z�"O�@iAɅ�V�v�J�)F�^�����"O"��ϑ�C��\���<w���E"Ö�v���Y�R�C#G�v��"O�;p��UV<9sV'�r�@�91"O|h3���9IX��G'�&4��(�"O�9xG��N�ثQ�v�j#A"Op��O�!����
=KXpI�"O~�V΀7%�j$#"��� ��P��"O��ɐ P�`lif�C�Z���@�"OJ��&��Hs��@�Ŋ��"O�(å@k̐��ӏ����"O@�S�ܳ[���qE��4$����E"OJ(!��ȑP
|�S��Y�0l@9��"O�x*wM �K�!a'� l��"O���Ȕ2Ax�t)��'����d"O�Sd�ʇ8g"d�Ĉ <���%"O��䏗{v����U -��!�"O�5����"� i��b�!"�\Pj�"O�xdB	;mr��4��L�	R*O"P��ľ*��0J��
:&&��'�`��Tr�(��oT�5+Dѹ�'j�]j����>�=�0K�:�a�'�^Ly��tN�G�66�0��'i`�0�ʓ'B 8�I�!=�4x
�'n	�&(�9`���%͉ۮ		�'H�mHGf�6 �(�dB�c�T�8�'K`�P��I���h4��bR��
�'Lp�-Q�N\Z�C1g�2%�v��	�'�ִ �`�;�z�Hc���q
�'��DJ�
��J�Ya*�;\"y)
�'Z�I#��֢Q�.	@Q�ҫ�^�(�'W<8��"H�o,@Cc��s*x%�	�'�������$+�����D\#4碠"
�'��9�d��e��
��T�WG�1 	�'�2��V&R�^��5B���Km^=i�'q>�	A�:�~a��I@�~:�'���S��4�B ����AI�h�
�'�x��r �QjU
`d��?�r�@�'	-�)Ѵ=ZN�����frL5�
�'�VH�q(�#k��-���T\���
�'�Ń���$y��SvjT?,��'�@��BJ$�`+L�HP�
�'�`x��̈́#���h�.�;�T��ȓ֘�jP�	B�:��2�ŧP`� �ȓB�\H2��ʦ8N��9g��*4B|��H)`i9S̑�W֔��,�&2wx��ȓG[4���H�O(�aif/�
h�|��$�bԈ�����t��T�v1��7&t�'^U�MC��U�䡅�Dc,|Aç��bet#�\A���ȓ`%�T����%���:b+ƹkVI��?X��h�IY<$����)'vh�ȓ�~|P5��W��l��JB�܅ȓs�iM29��D����q~���-���&� �2Oz͙ W�8j��Cd����&X/�8A����� ��bW\X�U)�<���#�Q'b���S�? 0:$�S�OxJMJҭ¨Fo��"O���Se�&j�f � K�9�"O6UK����W��8�`�$�`�7"OlM��$J�,�|PbԂ+ֲ�{4"O��hT��%V��q Ş?��Y�U"O��ZqU�k�8�Q5�~�P�1�"OX-؄+_
.�z��A��f5T�)�"O<���S ;�)q���bD�"O���SM3 FA�#O�N&$�Ʉ"O�8��E<n.��� @əA�TYW"O��³��]�t�(,�Y���B"OLi��"�,p��W$J�%"O�`��R5K�"Аu��P"OJ�1f`۶W�����BA�ę��"O��u 
  ��   �  C  �  �  �*  J6  �A  �M  UY  �c  oo  �z  +�  ��  ~�  �  i�  �  ^�  ��  ��  3�  |�  ��  O�  ��  �  _�  ��  L�  � 	 _ � � U# 5* �4 {= �C LL U �[ b Eh �l  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+a��6 \��	�<4�d5h��'�B�'���'	�'/�'�B�'��I2w��5Kk����e��U�D܃��'�b�'A��'���'}��'��'�>��5�\ h4tIR �>���'l��'��'���'2�'���'b�Iz�k�fVЂG�[�x.(���'���'/2�'��'"�'"�'�^�qs�S%V��c߁Lb>ıf�'��'@r�'���' ��'h��'J����b���@�3MTV<q�'�B�'�'���'���'^��'��`�$�͡9Ql�#[�=�"���?i��?����?!��?9���?A���?P�Σ9<�x�
�&�+K[�Jъ���O<���O��D�O����O���O��DLw�eȴ���ŢW�2(�'��O0��O���O"���O�d�O&���O,���ƏX���K�8�n͊���OP�$�O��D�O����O����Oz���OL,���0�"&�:3�f�j���O����OD���O����O����Or���Oؕ����JT�
�G�Oݨ��Ԣ�OT��OF�$�O���O����O����OH�0t�ʰ[O�XbQd|�^4�G��OP�d�O@�D�O����O���Lئ��iީ�ć/TF�U�ՁN�:�Z�34�ڂ����O��S�g~�i��ۀ]�j߈��'�M�Z֢��-�&��I"�M����y��' �U��)�5K� ���Ș]Nz���'��a��$��֚��'$��$�~j�'N)W=�9��3&S:�j�q̓�?.O^�}�6̡#ӂ�'��#������D��j��'��h�mz�ݱ���3�U'Г>���5G�͟��	�<��O1��t��w���	h[(}����x��h�p�@;mbh���<���'�
�G{�O	��T$n��zօժ7�.L�R��y�P�4&�XڴZ���<���ӞK���;Ҡ�?�:��Q���'݈��?9���yb\�PK����Z�ЁhW�%!��$B!?a�B^�t�uiG�'B_��D��?	e@!nFp�S�N�B���)]��<��S��y�酅0�l4��XN@�YI�(��y��`�"��Й��q�4����T��B�4X��9D�������yR�'L��'UؔKt�i��I�|�V�O�
-�P$=�����i�*d[Jؓ�˚b�jy�O���'�"�'��ݑp/nt���e���C���]��	��M�������O��?�Ƞ/_Q�X��Q����3� 
3�������4~������O��M�$Oώ�zh�t��� dF�6f\��dI�,�RjJB`�C���6L�.K`�I��ܛy��,��	�*�JEҥk� Ox����O����OD�4���b����[�<�r��	���	�HB<k~�yU�I�y�{�
����O��nZ��M��i�>et+@�;6�"T�Mp���P3�f9OL�PA�N�Y�Nqj4�V���d�����*��2��U�&!�h�.N�U�\|b0Oh�d�OR���O����Ov�?a�u$�)v�y���!垥� ���������܀۴,Ò��.Ot�nM�	�,�тFH� 
cFM�I�ډ�J>i�40����O�p��i��O�eY�Z�lJ������IU%��%؆����T_�O�\������	��x;>��A��H-v�*�$T�d�IAy��b�2hؐ`�O�$�OD˧XY�Pr���WrB�Y�T�8���'K��x�kӐ�&��'t�BDJ�2�)���"V��Q@��O�ȁ7a�T~Ҡn�%b�'I����y�F�{IԝI�W�6R� isoG�
U�'�2�'����V��@�4h[b���M�	�"}�B�V3�L�VH���V����?�B^�@"ܴL$
09#�#�T���.J�T<b@T�i�f6��j�6�i�d�ɡ��H���O[��t�h�z��ބV�z�'&B,m���c��i��	����I���	��0��`��CҠ �lj�Ô�5��ȫW�O�f@7�.h�r���O���'�9O�mz�-Xϕ�3�a�P�X
TC����	����6��S�'�4{�4�yZ��tׅUӈ��uN��7r��'�rYU�X�Px3W��ݴ��4��dE�X\��!G�P%���D�;��D�O��d�O��C��I�W��ߟp/		9�O��@0THV��gѶ�d*�O��D�O4X$���gi[ �b�Q5�D��(9�&n����UNT�F	ðSf��*��n ��?as��O����;Yt��1� ��2 4f�Op���O����O*�'��Q�ON��_c�p��Y�b��&���a���h
�֍����ɏ�M���w�(Y�7��{��<Z��E��t�'����m��lZ%A-��m��<��t.���㟸��V���!�W�4P@\p����$������'�r�'T��'	fY�զ��V�����2���U��{�4-��l�)O���4�S�>�U��G�b��+Ɔ��x�F��OJo��Mc#�x�O��d�O_NEJ�j��r��b�: ��d�f�
&���Of-I�폰�?�@�<���i}�6M�	��/�>� Ȱ�ڎF�"��������͟��i>��'oV�dJ)�r�qt^�:�m�/FP�e[�y��eӤ��y)OD�D{���mz���+�qN430<m�F1�`�64�V?O���(N�����''���$�u���� h���%: J��$\ ,/�t�&<O>�D�O����O\��O~�?����\m�P���nDP��B��}yB�'��7m@�0��	�O�mf�I�
��u#�lR��=b$����X�'��RܴY?�v�'4����i��$W�I��UX�L��<� �����pM�0F��r�~A������%���-O����O��D�Oް9m/��څ�_HP��{���O�$�<9��iLd1�f��7�O��'X �|#�H�DA0T�)	�G��$�'m�꓇?����S��)t�P�C���R�B##8���Cwkθ+�J�Y�O�)��?��b*���\�H�xD�D�b�����,i����O��D�O.��<yV�i.�a:*� � �0,���ga�4���M�"��>��?��5���'\+���?������?Q!��%�MC�'b�&L�����Ĉ7Ai�m�t�7���X�
y��<a���?����?����?�+����K��O�I�	�&�P�1`�E⦩r� ��������%?��	��M�;��%�v$O���� *Q�`a��'%�|�����'�����4�y��X T��lXBX�B���p�ִ�yr.̤u=���	>�'9��ϟ��	4��$�Ձ	����*~��y������#"n�П��IPyB$q��p����	��d�4��0O"�Dyb�SoK8��?	�]�$�شTFҔx�aEQ՚�KP�4�<��m�1�y"�'��H��Q>IV$� U�L�ӱE"b�BƟ Z��5�Kˊ_^Ɯ�0�\�,�	�`����F�t�'�8$C�5d3�8a�(Ҏ0��'`06��Y&d�d�O�m�Z�Ӽ[PJ I�����)q�@i0���<���ic|�x�\|9D%s�,�s�Ph���៪ X"e�V��#��L5���*`�'�������i�6M�O6���O؜�e�G
*���3J�?��X���<�6�i��=!`\���I`�')?�@#V71�Z9bfl�oNԳ�S���	ӟp'����H�I9y��v��~���DL6r�ey�	���-p)O���eh���~r�|bU����$;o-^�(��g���Y#"�l��ş4�I՟�SkyR�Ӫ�9�-�O�!Ӣ�67��t��hC4@9��
���OVeo_��'���֟�������[1e�=�$��S�׻�Po��<q�Ix6�*%��?і'����wE�X!e�F0<k�9��]�;�Lu1�'7��'eb�'�'%� y�IA�.#:���E��D[p$���<��;�����6��)Ϧ�%�\���ݨF
��� �;nc�T:���t�	˟�����A�릥̓�?�vc��g�dh�֎�|M�� �i����^D��I��vy�O���'�+g84���O6U,08�G��y���'a�I
�M�A`³�?��?��'�:2G�?0����H��Pk��KPG�T~�ɱ>I���?!K>�'�?�I�1�rQ�o��x ܹCs�b�������+�bq�'��$,[؟�� �|����0g�A��@|�vk�o�"�'>2�'���^�$��4`X�8`�?Z%؄NC/>6�� �Î�?�:�f�z}�Gb� h �"H)޶}p�o��kp]���ƦQ8�4:�j�#�4�y�'ENA�&LC�?a� _����K*��I��A�_�,5q�#{���':B�'t�'2�'
�S>~[�����X��]��r޴	�<����?�����<����yG$�,E���7�-q�z��P��7I�p6-����'���?���6Bl�o�<��G�I��@�"A�<&�ܡ�n�<��+$#��$�������O���?��i[��oy�Iⵏ�<ViT�d�O�D�O"ʓQ�&O�<�2�'�R�7���%�/6Ir+T�W)u��O��'w�7�����&�d˒�_��U�w�FK�V�S1$"?����n*$�Ɂ��'c/�d��?�Gl: L��Sh�I����#�Y��?A��?����?���i�O�P	�� =^�p6�˽JL9C��O����B���CU���4����C��Cr��X�IV�*�	��6O��$�O����;)�6e���	�
cT���O�|�J�'3<���(C%Ŋ^p㈊i�	Jy�O�"�'"�'�2Gؐ(�LAiU�ۧ����.Ԑu:�I�M�>�?����?H~���WGd��6��;?:2�;��.6,[bT���ٴC���#�4���	��sci˥�L���N�i�6�YÉ�N��]�`��x��S ����I�IayB9�(���LV4ڼ�����:���'���'%�O��I-�M+[�� ��
��e{��	1UG�� .Ҩ���M���i/���Mà�'�V�/�8��p��X��=�4	�$u��iA�i
��Oaؠ�������<Q���K�&V1�f��A�'�Pg/��<I���?���?���?����8G�j!����xd��,�?s5��'S�`�"�xs>�����e%��� -ۢ � ,�$�@+F��"�۫�䓪M�õi��4��+��1O��d�-������y.�B#��*^*��gM��?�G�;�Ľ<����?����?�`��JL����3&p�xa̱�?�����զ��a(�����ğ��O��Ѡ�,�-(,�5`��k�O�]�' r�'�ɧ*�'b��9�'�y�đ�b�=�:��J�3)�diS����$��@���q2��O艱�@R�t\N�q�bQt��6��O����O��$�O1�N�VP�&��3� r��J�%e~x@�&�\��H �'���g��⟸��O8l�r����H�*�)��߽BF�!ߴ����Y�F��>O`��&�&\���{��)� h�$&�'ql����2<U�Hjf9O�˓�?��?)���?����i��5h��Ӈ\�2�N%��"X�)�lڡ+���	�(��k�韔����+�i��62�* �X��l�g�K�b����f��%����?u��1C�Hm��<�'�W��u٥��M)E�1���<Y��NP	b��P����4�<���,L �y�T�[����o���N���Ot�D�O�˓^q�&�K`��'+"(�άE@u���PtLՙ B�]��O���'r�'p�'������17=]���F'&F�2�'�ѱL��s�#��d�����B��0`��H#A����?��p�Dm�OJ�$�OP���O�}"��-���g���|t���M�0��h��W���
z���	؟��ܴ���y���I��0q�dP�K&u{ӊ�y��'�1O��c��i��i��z#��P�$L�d���Oəd�Dѕ�T�������OF���O����OZ��M�h���.�jOX,���_�?@ʓ,T�-��&��I֟ $?��I4aQ����
gl�ѮG�d����O��$�O\�O�i�Oh����<�i[�N#�7�!��g���'z����-U?QO>�.O 	c��)}�����7D�uK���O
�$�O(�d�O�<a�i����G�'v\�[Ǐ57����S�B�M�aw�':7m?�I=����O����OBr�kȂA�2���S4e����"(8��7�}����X7�:�ҟ�˓���i^(pI���3O3�ӓ��'7��$��?1��?����?����O�$H��	8r:P:�ɡ?���z�',�'��6��#����O�qlZl�ɧOj�8�3L
�`:��J����]�L<1��i�66���Л3�s���	��h��K�+.T ��ƵXNIp���<7Rj,a��'�lX'� ���T�'���'�zD��ր;�*d;aI	q�T�7�'�X�0AڴW�^@��?����i�A @��I^�^ȁ��G�<����Ʀ���4TE����Ք�\��Fl��� ��S�ƸPM�
�;I�Zz���2v�R�U@�<�\Qs�'^zL��qN��.��	ٟ,��џ�)�S\y�g`Ӝ,�e"��N��z$˖�fj��KW�N5x'�/ϛ��D�s}b�'��-�#'N+�\��E25n���'A��Is���7O|��N�~*��?	S�O�9GF�� �8 ("(h�̀�0O ��?���?���?�����M8ZՀ��MIMxr��S#}�lLo�R�!���	Y�s�{�����/X�_�tC��A��|����?�����|j��?!4�V�M�'6�[gb	{��ĸw�Ԏ�����'$fѱ��
͟�X�|�Z��Sȟ0vB�>-���g@� HX��!�M�̟��IܟT�ISyBm�½h2��O����Of��bRVٴ���K�@J��X$E6�I���d�Ot�D+�d�^%�e�Nb�F$��&�2)��O�1�4���w�)�X�C���ȟ�˥��50��ʛ[2�G�Y��$��ԟd�IƟ�F���'8e#�ޤ,�B ���ϗn�����'h�7� [��d�O�un�Z�Ӽs�� 	�l��)�yh�Xk�/��<��i�47͖ڦ-a&�٦	͓�?����5J�l���
��ЇF�5zf�,�O���N-����4���$�Ox��OP��6T��j�,Q�:����drI˓h��&B&��'	"����'ִ� �.Ճ[B�`��Lǅ��*'c�>C�i�p6��q�i>i�S�?�K��HX1���ډY,�8-�E�1L&?9�BK�|Y��$������d1D��l��O��B��2�����O^��Oh�4���x�ƢΦd����j�*q�D��Y��1���^,҂rӀ�$�,O���v�Htn�6��`:D��3"�N��+����4
ͦ!��?� �!a	J�ɓG~"�O�g��v!�u:7�� 0��6'�y�'���'8��'k��I�&:xn��.	
m'x�9�KD�Q���O��\Ҧ��0C~>��I��M#O>Y$�F����Ճ]H<5��iσ%B�'[�6N���CY��7-#?y$��V�ā�!o�).�(�
E��v�V�u��O���H>�-O(��OV���Ot��k���tCIW�;E`�(P��O��$�<A��i���'��'5��.YÊ��猎�lR�hpd�?���C�	��M��'������(]l4K%�ݟ>�ࡶ�J79�T��eO=XԀ���A�<�'3�~��O���.��a�5�^)JB�gmWy�2���?Y���?��S�'�� ��A�f痷�ɀ�gӏMr�` f5K�|i�'�47M$�	����妝����~���:D��A�M��M[��i��h�Q�i����Ol���7�Z�l�<�D���srN��B�N�(��sM@�<)/O:���OZ�$�O��$�O�ʧ}晋�!')���D�4+����i��)��'���'���y"�r�� 33=�!C"[�;���bL�~@��O��O�I�O���
�T7m��K����M�\⢮�\)�֌c� �$e��.����R��`y�O��� �ҝJ�(HZՊAoER�'���'��I��M�3�K��?���?���X�&p0��́�&x��KC3��'sx듿?1��� &h���m̭e���[a㒄t�X�Γ�?�ָXuh`��4Z	���?�c�O���GT�U����������O&���O`�d"���ҭ��@���g���C���pD���?���i&H �0�'�{Ӳ��?��Ͳ���`aL�pP|�75Of���O\����K<7�|����GNx��π ��* �
2������8|#E"@M"�$�<���?���?!��?�7$�� p2�N�_Ԅ%��!:���BȦ��v
��\�	͟<���D�/�VM���MhD,*���zN�Iԟ���y�i>��	��8{�o�,[�^L����9��8;a0�>lZ����	X��'�'/��7S�T�� n�#�X���\%]\��I�������i>Q�'�B6m�Q������<�BFD�|625�&���Oo�D�æ��?q�P��`ڴ"��VHd�RL��Guyh�iw,Çu��a�ŤN�q|7�-?!�)��	<���Y�C�;e̅b�Ε!1<t�$g��	��	韼�	ϟ ��wAأ^��BQgΧ@���w(���?����?%�i�N�P�O:n�N�O�}�� Z ��*��׋J$z�[W≧�M�7�i��T/	�囖8Od���"�I�dDY�0�* �g�޳5� �T�Z$�?Y3�"��<ͧ�?Q��?�J2�١���E:���5�?a����@ڦ�) �ʟ��	��P�Oq� h���-Q��V�/A�y�Oj�'��6-؟�&��S�?�ۗ.�:�(�A�L�i��k��}a�Y�CB5$Ę��'�����ʟ,cv�|���t!�@Y����C }�r�'K2�'���[��bٴL(��㑇���$���1&����&^>�?y����f�$�f}-l�<�9�g��(��:���2�ܦ�bٴr^R�
�4�y��'�X8:S̈́�?�!�Q�Ȧi��f�x`���<#@e�E�c���'���'��'	R�'��B��3a�����n߬-:As��:�M��(@��?����?�M~����w���#+�1��=�#N$MƖP����$��	q�i>��S�?yPP�ߦ�ϓFf	�Nڲ;2^��	��3��E͓"�,[s�O�qI>q+O^���O��@�'ZQ��	c��A:��;���Ov���O����<Ǻi�����'���'k���* 8�����T��!���C}�'|�AR�o�Ё�U��/c�`E����yR�'z@3� �<��'-��	Ɵx�b�Å�޼���X�L`��eI���,��ҟ���ӟF���'�LMrpo��&��#���v�H�XA�'��6̓ A:˓4����4�`��`��-��ge9J���SR4O���O8��ӷ#s7|���'}���C�O�H8�&ٸ#��z��f|�T@b�|�\����ޟ��I�������k�T�!��4Sq�B7|B͊d��˓J�� DP��	�0�r!�G9r�\$'���k��ز��:e��	؟\�I]�i>��ԟ0�$�Ҧ\���p̓�{�)��1�Z�l5��$I/?�E�'?�'��ɟ	C�`�g�>l$�F��N��,��ϟ�I�`�i>��'��7ΐCs��$[��|�񤊒 ^�*�bS���Q�?A�Y�<����t�ɱ�@�6@%�h��n݉P�Z=���"87mf����<M��O�J��*��(&��iF	^9j�3ԫ�(o�l��?I���?Y��?�����O���Q��A��x"w�Z�\�@=��'Nb�'��7�B���D���|%لY��)�W�R�!y��5ʘMT�'�b�'vb��(wx�V5O��DJ�!�0=����Y�X���D-����ő��?�%�-���<ͧ�?1���?q׭�b,��g �-+0%r%����?������̦�'������՟��OhRm9�΍�-�X��f#A�z5C�OF��'W��'�ɧ����.�rh*��V�e��4�!Bۑ,��Ik�o	2��	����S�a�,ST�}��D�!�G�fd�wO�r6��Iџ���۟ �)��^y�$y�`%YpƔ�R^JA8���'`�B�% fH�nO����S}��'s��Z�G��)��ِ����8 0�'��2������� m�>*x���~B%B̡5q�h!�k�r��!��W�<I+O����Ox�d�O ���O`�',t����Q&| b�J�-�@9�i3&m3 �'kr�'9��y�Kt��+v�q'�Ʀqj����G3-��$�O`�O���O����':R�7�c�|���ܧ�v��q�.~�p�p�}�t�`nǜBRIg�	\y�O*�P�`7�ų@C�/x�%z�Co�"�'b��'l��M3����?i���?1�, �	��բ'Z8.DЄ(��7�?�H>	�Y�Ȫ�4:s�F�(��>4O�ф�Ŗ%��aY�g
-�$�Ol���٪4��𱓟��5TnBcGԟ����
%a�ji�у��%	lPsl�ҟ��˟<��˟�D���'2 e�7��m�Hۂ��zUl���'�6�:[���O�En�F�ӼW�L�,#r�
v�Ӫ0G�Pc� ^�<�$�iL7-MѦ�0�/�Ȧ��'l��V+��?�i�*I�,d�B�LۦC2��խK�S��'�i>��I�� �	���	�O�<U�P05��0���,K<՗'��6���a�b�d�O�d���˧�?�ׁ��'���Ӭ^�J��m��N��
��<nZ<���?q�S�?�B��ܳ;��u�C���b�$��$Q�9�1���;?q�)�y|�$�7����$��,��A��b�h�?U����O���O��4�>�x����"�$U:A��)M�l����-P��s�2�x�Ol�m�"�M�"�i� ո��[���s��>v:�����3?�:O��DN<4>
��'(����?}�]�x������J��j��:2B���$�	���I柬�	q�'SN�ڂ ^2U��P��Z�Km(���?	��b�v�Y=����'NL7�!�d��t�B�ዩߠ��UDH�
̶%��h�4Q���O>�E��i����#��� .��,F�Xf,�i0,�< 0Å��:�?�e�2�ı<�'�?����?i�"�t����GU�D�r�˵�?���?���q�@�H����?�(�r�nz>�����@ܠ;���I4�4��f ?a`X����4a���n0�4����-4N����	 �bk�hQ�w��њ�d�Z��{֗�����o�R��]�I�z>��:��0o~$��D:62|��I����	ş��)�SWy��x�2�ڡ霑X�	�'"�{!�J�!ؽU���d�O��mb�Er�I8�Mc�OӔ,D���2� �q& �^����e��%P�Ct�(�	��$p�(°5���A \yr@*|"���H�{�S'U�y�W�h��ٟ<��ڟ��I��O?��@']7P�2��4-�� ߒ�
u�z�Ȁj*�O����Oj���d��]7;�]���41*���c�Ī�.��۴{Y�x�OC���O�n�0�i��0\"p堗F�!$k�9z�!ڊu��W>i�:�0�O�ʓ�?y��-���#�d�-�����N������?���?�.O�mE�ة�'��Ŝ(g~쪄��*j���bă=.��O���'Gx6՟�%�|��[�m��S��5�d@���j�X�I8ud��K N*��\�'��$�A��d��'O$0�pNGL�iz@4ҮA���'���'�2�'Q�>�ݮ|3pX�G�K����ި'PV��ɖ�MF	���?��/����4�����7 "��� ��\:|�p�;O��D�Oh�ė1O�@6�y����k:b�`�O�F5!�"�t�8�b�Ν��0mC�|�^����ǟ��I��H��� �`M�?���5�<JD�h�QFy�q�N]�3��O4��O���d�}��zt.�W�Y�"�w���'���'�ɧ��'�rD�*�P�r�գq�p4�#�إW��"4�iW�ʓ ��}�B���$�`�'Q<���Ś%gȰ�r�'���ȃ�'2�'>����4Q����4{�����Qjq�«��/�BŒ�a�:IVA��_��F�doy��'K��jbӨ�J� �lR.���iе�@�J�fL03!6�h�@��Q2�4{��OҤ����Z����ԃ�#�Ry���
-�Y͓�?���?����?����O�,Ç�%"�e!����S0 I�'z��'\7�\._I�i�O��o�A�ɷel�	W#͊[~. ��Z8~\KN<$�i�j7=��$�|��m��Y��=d,ʩ�I �a;���$B��n��*����4����O�����S`�zU��+e<�A��bM��d�O˓7i���K0��'"S>�J�\�z#�xP"���,1��O(?��P�0�ٴH��>�4�"�i�s�e��� �>�s�h�/3��b4ǋJ9��ZП�������G��s N���͍&��]x�`��+������4�	Ο<�)�Jy2�zӼ8�G��%g������}ЗI�;����O��mZr��Ys��,�M3SAE"4:ѲT�j�ZfGZ�J���h�\��f�l�j���8���'1���k4?�r�(	��)@��M-E!�-:6��<�(O�d�O�d�O����O6�'J������DJ~JU�Ŋ����a��i;P ��'���'���S>�����Mϻ3;RU�w�V�W�tm #Obq��9��?aM>ͧ�?��g��4�y�-[���!�a�0;�YY�C��y���0������D�O���"�*��A·B:la�qf9J���O��d�O��<��V�����'b2�0}��X჋;QP��E����O@��'���'R�'l�pR�]5DRȭ�eM*jx�I�'1R�\_���h��iH��"Ǉ����	}7R��·Mj))o����I۟�	ğ���C�OV�gJ�7L*T��PJs&1[��nv��d�9U�<�$�i�O�.�=�����_�(x��w��0P8�$ͦ1�۴m�����!��61O����57�{��:̕RF�X:��G�PH5q"�5�ķ<q��?���?���?��J{D����@��	�������D\Ϧ�ʕ�՟��I���&?��	����!�F��xpp�*{�| `�O0n���?�O<ͧ�����J�y�Œ�RS@�d��OQb���*� NZ2Ai/O6EɁ"�+�?��4���<��� h,!e� �n	�DI���?A���?���?�'��$��!�&`�ϟ8#��J�e�&�sbL	I��@��Oi�(P�4��'����O�OL6�G�&�@���*�XJ��W�<0��`w�2�]E�e�����%�I����루�?c�Ly�A.>6�?OH���Ol���Ol�$�O*�?98ׁ�#U3����&.��R�,�Iß(s�4-�ʙϧ�?G�i��'v�P4%Ě$�~ql9!��0JU�|r�'��'��c"�i7��?�$'
cF���*އ4�i�O�$Hy ����䓾�D�O��D�O~�$����e�gJ�k��c����Or�44�F��/l9��'��S>��f������K*B-:Я<?9S��I�� $��i�X�q�ˀ %��;�D#�����]3����0Ö:DX�ʓ�r��OaYI>��������Hd�j4��?���?���?�|�-O�9m����pH�45vܱ��6C�2Z@�_`y��nӼ����O�����c~�0JgJ��,���;��G2a�B���O���$�g�^�I]:d�ܛ��tW���I]�o�>m��*�-o� ���a���'���'�B�'���'���N����W�h��(JP��)?Z�Qxݴ:|�����?a��".��d�ߦ��/ջ#KY��dG��A����ߴZu��6�4�H�i�V��xӲ�)� �h������~����"qNέy�3O�����T�?A��<�Ĵ<ͧ�?�HU�b�\H`攃VD�� ��׈�?a���?!���Z��������������*��N�O��Gm߳DC@8��k��q��I��M��i�OV�����-�(�a��
.��7Ol�$��W��I�*f�	�?-���':̨�	)	+3�HFg��*a�L(R�������L�I��X�Oy�G��1�$����ծ(�<ӑ�M�sqd��8(�a�O������Y�i�U����0�f k��*C�h��w@z���43/��p�R���y�p�	ȟ�"ā�} �T��05&�;Ca��2���(�`����$�̔��4�'��'�B�'o�M�sl�yc��BM�"��FS��h�4zOnh�(O���,��wJ4�#-�f����܁q�O ���OԓO�I�OF��E�y��P"E(:P�D#bN[����a�	3�	
��[��'f�$��'�e��I�h'��{�(Þx�$[B�'��'�����dX�<[ٴvX)y�)�D���H�Ђ)YB�Z�5J�՘������d�n}��'��'��QD�vZ��k�a��7.�R�Z5^���?O`��ťc��H�O��?I��. �8�TOLh�%Q�(6R������ߟP�	㟼��J�'
��A�J^�V!s��6�������?9�����	����'�7-�O"�l� ��,E�6+T��ý/�.��N>�ܦ��I�D���즵ϓ����;wR��U�"|���^�<�LP�S�O8�O"ʓ�?���?���sԚ��T�]#[>uS�A�t� �����?1,Ob!n5h(\��I����	{�d ��⹢���,1���z����dk}��'vB�|�O��h�?��	�m��!�YFmʎ}�&@B���4�V�<a�� ΄��C�	�R�Ї��4Q.�(���	d�v4�	ܟ,�I䟐�)��uy�`d�����q6����[_Kd]��"��vA�D�OfPll��k�I
�M㕥�k�hA�@�@*�2���2>[�&"mӖu�0�k�~�i�i�����Oy:�"��N�8x2��C�	�8ӊ��'^�I՟���͟���͟��	g�tLs��r�dK1�v�*�d��D��6������O���8���OPioz�iC��V�z�LE*E 4~S����ő>�Mkr�'����Of�{@�i���ߤG���R���Q@���Z��.Aނ����YJ�O���?���`|xiaD�Q�~�0�@�V�>�t}z��?���?�)O�o�b\��I̟�	���U�@���І%
�@H�?AUS����ğ`'�p97�F�}:Ҽ��ۥY`+�c�����"ަ9JxP@Q�,�Sz�AAן�k��I;_|�iX�N-1s(���]����Iϟ��Iҟ�F���'{��C�	vBĚ*Y���5��'b 7-Z�RH˓Od���4�`�� T7z+:�k$>�<�+�7O�}oZ4�M��i���ⰾi��O��7��>����Hjjze%�z��%!q���ir�!�d�<q���?����?���?ɠ$����C�]�ﺴen�����M�a��t��Ɵ<%?�I�q%��
M0u�"�n�'�Z��O����O4�O���O��Ξ��q"�
R.8�uy aқcN2M�&C'W��I�7��<�0�'�xE&�4�'`��SU��
���c5PD��R4�'��'/��$Y�܉�����ɋ|y�r�a�?'~�3 �yD�扐�Mӏbʩ>���?Y�;dK���J���B]3Y.�P�]�4��n��<)�;��SF���'t�4�w5d(J f��pq�n-��1��'��'�B�'{R�'���P� �bQ�|�*�k�O���O�xm��@�v���T�4��ª��R�G�sn��n*&�(EaH>���?���/���4�y�ܟv���a˃+�y2Q��'
�м�c�P����[�IEy��'4��'5��"Y��3�b_�{Ԙ� ��+3��'j�I��M[��H��?Y��?(��M�3oٍ|�Bt��ٰ$�p k枟�Op�D�O��O���Ov!�E�G!r��t�L�I���,�wD�}��nSK����?��0�'���%�`K󤉀8��x���S�';�M
S������Iޟ����b>�'��6M��%�>���g�M�&eI�Ǚ%�|�rQo�O���֦-�?єU�x�I%^2 ��e'm��Z���	>����ȟ���Ѧ!͓��4cԤm���<¦�����U�
v�ei����<�)O(�D�O��$�O��d�O�˧'�|4*�!��*�4DD��o��ԺP�i�6p��'�r�'G�O��C~���ϥh��j ϕ�E�E)�cU�u�~���OZ�O���O�䃂W=�6-v�$BԦ�R��8��KR �vZ� q�l+E�O�]���9�$�<y���?Ĭ��
�Ze�ec�Gr��͏�?)��?������9��ܟ������E�u7$1��"�ڱ������T%� �)O����O�O�Y�[�f@@�W�<3�y�e4O�\ :�ʠ3���YP
������OxAa��R���Ss%�q8�Gą�0͘���?���?���h�j�d�9H����&ś<$�i�T �j-���Ҧ�҅M����!�MӍ�w!�c���|&~� ���׮��'@6����ܴO֎}Z�4�yb�'�>�h�L��?�cQl�:e����#��	1%�3_��''�I㟌��ß��Iǟ,�	.�0С�Dk�֩��L�x� ԗ')�7�2td����O�.���O�m�uw�teq�[<H�P`�an�v}�ok�:���f�)��%~�� ��[��2	�,�Xl��Z��Q�Q�:b8�ʓrzH��O��H>�/O�|81�ǪL� h��6#����D��OX�d�O��d�O��<	��i�����'�N�[��.���썣:g�A���H2ڴ��'v���?9��?IpHM��m���|��ԙ��1!�(�Pߴ����B�O��O��_�J�tĂ���3���Z7�y"�'~�'M��'���ɘ�S,�sU��a.� JR둾V�����Ol����mˇ�q>U�ɶ�M�I>YE	�u�Dy"@	Kk,��Y���?��|�2�P��M��O��\��J@�
>MQ�8���B���EL��L'�ؖ'�B�'�"�'a
qsC��> �� �яe���%�'`bR���4a�r�!��?I����I�x�r��Q�,���id�;��Ʉ��d�O\�D'��?1���>�r��W݄($�-����Q!�9"�J����*O�IP��~"�|�J ��}IC�G�+�4��@�1���'X�'O���\��MCtC����U�� t��AB'�� ��M���?90�i��OƉ�'�(7��1$%�s�M29� ��H�3JQ(�m���M�D*[�M��O>-qwŎ���N?�JC� a��mCz����g��'��'�b�'��'O�;S�vY�l"��m:���AH~آܴ�l�z)On�=�I�O�nz�ђ���8`WX�򲫝 >�j� U���M�i��O1�!�կx���-N�By��*l����] �8 A3O6�F��?���3�$�<ͧ�?9歗�1}��vm�+m����K1�?���?�����Ӧy���U��d�I����4F�?��p�C��L
�	���H�3��	�M�4�i�6O< ``�1!�Ь�F��P��p1OL�d�
"��	
���:���?�d�'|�IG>�b1�D/g��`�R�U�����<�I�|�IP�Ob"�-
TR��0	�9�M�C.�8^��`sӶT�3G�<��i�O�N��\��Q�m��<�};&���qU�$�O����OHd*� l�0��П �vIN�q��4���X�*��
*yC>8�L�+��%�0���$�'���'k��'lp8(6��KZ�I���W�ؼ{�T��ߴ8b� ���?y�����<�"�(�v��� 4X�L�c�!*�Iǟ@�	z�i>��	��1o-F�~DJ�%Y=Z]tYc�,�/j�a�*%?��BS�W��T
����d֌q���1�A&FfX� ��>%a|��|Ө��@��O��i6G��5��[`��#{���j6?O�,m�[��IJ�I۟x����4�'�[Kn2L��9d�f} #Y^eصn�C~#d�A����'���Α���VN?_.X�&NJ�<�	�1���F�2��3%F�#�f��(O��dԦee.d�i��'L�Ii�N%c@���A�L$720��|B�'�O8�{T�i*�i��h��O�}�<A��B�"�9Ң����L�����$1��19F9cC��?M��-��K|�|"<a��iTp�\��IT�t�9e�У���%#��5Q4 \����e}2�'�b�|ʟ�U��K�l�T�2�T2N��i��]�<ꆘ�'q�J������LN?!M>����8X��1X��"I<)��i�z��\Ѝs��S����IL�I~�\��޴��'��듔?q, 76~�B����Y��u�d�?y�m�!ڴ����:�ʧ?M�'��uq���3;N��J2
�
<�I�'N�L��0{2)G$,6&����l>D�'��M�e����O��?����;p���KBA� f�0��;@$R��?����S�''���ߴ�y�"�X�PI/� R��`Q��yBՋ4�P�������ĭ<a�m�:�m:2��[�PH(�fM�TA��җn�lyR�'D�� r��ItD�B�#N��Z��P}r�'4r�|r)S�G`N�7�����@T��,��XQ?���U�q�l}'?���O,���k� ����×!<��b��c�!�d^,i�6�e�(��TȠnZ����ŦU�ZXyrvӆ�杈-��#�ҋ
���J����[�d��<����
����ug�U[��I����Y�$+�.��MC�c�)}&�O����O���U�00v � ��є� %����۴&2�@s.ON��'�S;X��	��Q W�t�+f�C�K�R%��O�D�OD�O1��DR6hD?;��0�����ɸ�
F&E�7�QyOFU:0����䓟��'�q���G/Q�6h�`�Pc*a|2}Ӫ��"�O\H �-��M	�9��G_��%;�2O��n�[�X����I˟��Q��~LX�(��-l>�A��B}Qp�n�n~2��j��'��'ݿ;&MQ+[ d�.�U�l��%^�<���ca�P3 �՝4�p��>�t.O��d�ꦱ2�#jD�iF�'�t���ꈬr�6P�OT�}�:%���|��'��O��(7�i�i�Y�ƭί L��kD��
{961������������1�ɟ>zb�Y����Lv �N*�."<Ac�i��|��W��IM�D��hs���`���>>Uہ�����D O}��'T�|ʟ� 2����+HQV�5&U�7X� 4OC8^ZT3�j�ꄗ��D�i?AM>9C@@���Qa��>("0e&PQ<�a�i��QS�BG�G�!����n�pq���Z�E/�	��M����>y��G�� ���d� U"gkݛ\G �x���?i�/B��M��O�N��c�$�S|yr@º_�N��MO6A���)ݧ�yrZ�������������П��Odx�2Pd޾�1��#���.��g�i���w�'���'���y,y����87o����㗹A�H0y�0-̅oZ��?!O<�|���N"ôl̓>x<	��gT�-1����$ޜ"c΍ΓK}V�0B��O��aH>*O�$�O��9�gJ f�2BPϚ�$4v�`�O.�D�O$���<y2�i�a�g�'�2�'26؊e�$E5��t/�6�L����I}b�x����H≞��q��.'�,P8�,�=���_N�XЁ�^{�I~2��O����u��2dA�(�ܙ��"�'/�"T���?����?���h����V0l ��[�J��u�&���x���)R��8�I�MÎ�win��0��,S���0P�ʝ'���'¯Аskl�)�O�L�/n��e��t���ɠ1�������-��\$�ĕ'b�'���'���'1��ET�_���;jV:�{aP�drߴR�����?���䧀?�7�Ғr��0S�)Ɋ/#�AP�$�	���ҟ|�Ib�)��50�H��AkP	%B\�D��1~g�EX��(�*��'��%��A�@?�K>�(O�Y�qƟ-\[^\�t�ڷXުP���'��7�����D�+ۈ����A�B���a��>��$E�%�?iZ�|������[U0���Z!72H�kX�';`���*A��O��*s�?5'?���$l�����D�\������+,��Ia����.=4088����dy0����Kkyr�'��7��,N^����MSO>A&���bK���E��t�h�fD�����?��|:&ߌ-QA�u7�̣?�R��v-��(QI	)�4�s�O^�O ���'%��`�
6K��LsBI�?
����D
ߦ�K"��\y��'�Ss���:g��L��P�.C;��A��	Ο��n�)���f�$�C���2%���.�(�����5g9n�`)O�iN�~R�|�畫Dߨ� 4�ڹ;��P2b��xR�sӀ�D�U�pG����V}R�=�E�z�P˓-<�&��WO}�'�f�L�:?�-{g�LY<�}8��'���'E��d!�O뮐wْ�]y��M<�`�j�=g{H�!0����y�^����ٟ��	����ϟЕOq�"'�#!�Mh��Z
}9��h��g�tydd�O<���O꒟�Ц�=1P.���_>"~҈�WJ�w �Y��֟�'�b>��#dӎw ���&��Z��g�
�YǀP��牯E*(xF�'Q$������'��l�-����T�C���?���?i����$�¦����۟�	����PF<�����+� :�`�h�}�~_�	ܟ���a�L�:Tq���
(4�qL�2:ir�a?�P0�,/auƼ�|����OҼ��@Q��IFĺ8tQ�1a��M�VtH��?9���?���h���FJ�t��ҸS�؄�4
ˤB�2�D�˦���n�[y'l���^����Ě+7Dēƪ�1���ǟ,�I��������r�{��Ւ����,�w��~� �Ƀ�DZU��"�2����4�����O����OT�����m�K	,�J&V�N� ʓ��d��0��'����'�(����xH䑃�o7)�̔Ab��>A��?�O>�|��7{��H3R�+�.�a�&݌b�n��.q~�M��6���bG�'��	�L*xՉF��)�F9��"A�cF����ڟ���ҟ�i>Ŕ'�7m���L��X2/`�96��5B����Տ�s��KަI�?�W�t�	ß��3P��`s7_���fŘ2L���"���w��d������2�>5��@���Q ���NA��	(�[����ݟl�Iʟ�	؟��IB��?�(m�8}�y��#@i��0���'f�'ff6�����|֛v�|��Թ`�ш'�:UiNHq���u�'����TK��o����O���U�X:6a�։�%*��ط+ �!�r����j���Ov��|J��?���l��5��Ԩ\^��!由R	ƌ#��?�+O��l�$����	ܟ���i�Ģˋ�L5��T6aȘ@d�F���DYh}b�'�|ʟ����_�(z�Ex�-ޞq�L��%#T�La#��2��i>���'o��'���,�5M$�@��ca��Bݟ��Iڟx�I��b>�'j\7-ث��x��	��֙�ׅ�1���ђ��<p�i�OΙ�'1r�$l�)�eњZ���Xr�ŕ@���'��R�J���������(r�'��S*�x�7�Ġj��5��@TUa>Ӣ�L�v7b|J��_&Rl0�d�<7��$�����~̒�BCSIYN��#�	�$�XX#�)'�nǋ�%	��*A�?V���i��*d�(;S������gY':�ŸSDM�<8�ZشZ�$���O�Jq���_�P�l�"�+�*F:ДHta��i�I&H�j]�e�J�^#N�Pq�X�L�b)ՠ%�h��ˇ�7�"=)��O,�	;
[�R�T(��іh}F�����	�إ�ɂ�#�r���S�{�^?���p�d���6H����nÚ])sm�9J`ul�˟��	����'Cj웗��ed֙ e�ҦJ;D��#�n�����)�'�?���  lP�
 -���H�
ԞL��c�i0��'
R�S�;��O���O$��8ypr����om%�D+3_�`b�p:UF9�	ҟ��I���A��F���;��F4Q�T��@�Ms�"U���x��'���|Zc*�< �$[�9 9�LZ>Cؼ��O�����O����O0ʓ22�Sɗ!uX8d�+��mj~�էZ�U��'�2�'��'��I-!Tx* �4{��C�e��tQ2(�	ɟ����D�'40`�R+i>��,f68ڴ�Ė[}Z��b�>���?�J>+OFyp]���Qd؃b�±�M�4+���>A���?����I�9�U$>����Y��4~GL��Ԉ�!�M������6(1�O�Y( �)_�@�q��ʖ����i2b�'�	�$m.��M|���*!�N(�n�!�C=wmX�(@��)7�U���'���R˟�i>7��]�p�z∋&S�TQf�X!��[��(��?�MR?1�I�?�(�OXq@�74Pe���D����@�i �	�`�X"<�~j��c`�y�ӼG
<���-�ʦy��Ń��MK���?i��2A�x��'��(:��F����3�F��OxӐ]�S�)�'�?�AN��1�C��e��Y����8���')��'Æ�z�7��Пd��f��iT*�QS"i@���~�&L�>��Mi̓�?i���?���^$�"�h��KB��A5j�4.���'�DM��$#�$�OJ��-���&��6��Ltj�Q��);�^u!��������ϟܕ'��Q�"���Gka��n��r4ld�ց\�/�~Ol���O��On�'s�a�TDA9h����#�9�d��}r�'���'���2�fx�Oz�lZq�B#�0`jqΎ�S�<U��4��$�Oz�Op��O�jK����&˯@��<�AM�~���)�>Y���?����d�t��O�2/���� ʆ�0��兡k�7�O^�O��$�O�[�D=�X#2�ٳAzB�х@�`��6-�O��d�<a� @�x/��ߟ$�	�?�`�����T�P/���ݺ�_��ē�?���J�X���ڟt؀qn��\��9	�!zR�8�T�i1�I:/rȈ�4�?���?��'}R�i���`�4�ܡ�˂�P��a�d�o��$�OJ�3�n�OƒOx�>�X�'��n};�F�A����cn�l%�� ���������?���O�˓'	U�5
��IUnͧjR��2�i�4�b��'��'=���D����$4'��!4ltEA=��mZן���Ɵ���V����<���~bF��#U�T�r��i��(��'���'��PB�y��'�b�'׎,�v�9r��ac7xN�K��n����a�'{�ǟh'�֘�3�����i
��hU ���<y�$��\����O6��O��< X���镘P��L'�ܡ:gʩ�@	�m���yy"�'��'t2�'zZ��"�	��i�Q�P�8�K�
�
�2\� ��矀��py�)t6��S�����ˁ-s~Ҥ��$� O�>6-�<������?���B�Z���pӀ�ˇ95�LL#�`h���P�h��ß��IVy"�i��ꧮ?��-���*@�X�?A���d�:���'&�'t��'�NY��D��U�5�Z�d��p�F�o;�f�'��\�\�C��;����O����ND�vF�/'Fp�	-$��u�KL�Iҟ0�	/�P��?��Ow��+S'\p�P��Ʌ�P�v@B�4���R*d/6�n/����O,�iNh~b+� &��3�W�D}$�#� ��M,O$���O��'>I&?7M�$��e�֡L9q,��攷훖�%,r<6��O���O�ISG�i>%��M�#V�Ʉ�ײc�� �k���M$�	��?����1�9O����FN�h!�(J.�bW���
f�5o�$���i#�����|*��~�O��(�����K�4Q��ӱ�M3����d�!�"���y��'���'S��p�o{�9�R�[�Wk8���g����F�LQ�q'���ݟ�'��]5C� ��*Ǧvna�W �D�X�4AȽ����?�(O<�������6�I���4M�9A(N�)�	�<���?1�R�'��	�����e�@X��_�P��|�dF�Ә'��W�d��G�@i�'Cb)��
rb�5k�8Fs��m�d��i��?1�Α��)O�)��;8���c*D�O
�mP'8��Oh��?Ad�ܜ��	�OV���ȓ|�!lGP�̵#�(��}�?A��?�	�3b�t%����&�޹�Ջ�w�8DAoӠ��<��R	I/�N�d�O���ƞ(�͞;ö�"�@^� �����xR�'@�K�*6F$H�y��R�r E�D��$��/���vW� �ɑA=|����d������JyZw�1�R��;f�P���ǤV�:E2ڴ�?q��91��`#ńX�S�t(>��eB�`�h5�p�l~>�l���N(�۴�?���?��'1s������l�h��T�}1݋��8�26�ՒL��D�O�˓��g~2��|��L���C舚��^;&�
6��O����O��$�<�O+�3RZ��r�J"8	J��&
8B����dȅ8�$>��	՟P�	+P�Eٲkŧ�	/T�	��@�ߴ�?���1Lb�����'��'P��J��/=���Vd�+��p�!
�>Q�hS��?�M>�����d�O�<� ��R�ۚt�:����P̜i�G�Ĭ����OF��6�����	���Ĺ6�E!r����
c��` �#�c�`�	wyB�'�j�#�џR����)$\m���x���V�i��'��O`���O<	Rd�+���I�4	�!0f�V\&��K��$�O����Oj�d������$�E�	lT8#�Ą'8��-�~�H�#l�X�$&�ħ<�f�[�?yH?M0ABJ$f��0�CV,��j���d�Od�Mm��`��t�'�\c�b��m��&��C���f��UXJ<�/O�t��O�O2��,���&3�X��\��@��b���g�dʓ3�,AB�i0��'�?9�'0��I�Cܐ�2g�9�
U�P�T6M�<�AM�?����d��ܴ1K�$+���3���'CD?�9lZ5](�)���������ryʟ�$���S#Q`K I�Jx��f����Z�N_��b�"|��Q"�@jU� 2�h��դH��jƿi���'���#B5�든��OL�	(E����v$A���a� �İ�6-9����,�?i��ϟ�I�y��0�ͽ.\(l��Ave֭)�4�?��CA�q���Xy��'��؟���ʹ���5���Hg��~���"_hH�'�B�'~"�'W�I1A�zuXAɀi��h�a�P�I�W9��d�<A���D�O�$�O^��B���f�z칰H0u��#�-�$�<����?�����0r��''���ao�xF´B)M+�z�l^y�'z�Iޟ��I��\��	v���@>1ZebӅƇg�@�B
�M;���?1���?�(O��cV�G�d�'��@6��bl���0n����k����<y���?���̓�?��'��x�ᔑD=@`��۵Y ����4�?y����d�el��O	b�'���D�'�%g� ��ի����/�
��FT��	͟x�I�)���Пؔ'����}�;QJ�?h�&IS���;ϛ�Q��;TL1�M����?1����Q^��ݳj��D����'4`���"F9Xf�7��Oz�dT*KC��myr�	��C!�@��)�<sV��BP���f�H�H�07m�O���O����f}U��
E:a��0��9I�L����McъD�<O>Q����'��9�$Z�]㞑Z5�O�B�6٩wOw��d�O��?���'����p����q���Ʈ2ĸ�Y6��3pM^�n��Д'�=*�����O^���O�qH�C�qąy�.t�sJ�ͦ���~~�!��O"ʓ�?�*O ���:4�0K�1Q�%TEF�>��R���Ш|�<�	����	�X��cy��/��+S�+V҉!rHK+=O`��ľ>�*O\�d�<���?y��d��|k���	?վ���A�5k*E�Cc��<���?Q��?�����=�,��'y<nd��a���sE�sM��lOy2�'g�Iϟ(��؟�V`i���f��<FK�k�9�b�jeXHlZ�����˟�IKy ��꧒?���!=5 	��rh|-1n[5I���'��ȟL��ƟЩ�Gn���O�ݑ��37���i��{�R�y"�ib��'��I�B�������O*�IH J�@�2.��ڸ|��E5�ju�'���',�j�����<��O<Q���D�S�(@�3[a�m)ݴ��$܅r�xoZӟt�	՟$�����~�rE	O<\J�z%Û��Q%�i���'�\�'���'����P*���"A��8�j�)�V�O�a�z6��O��$�O�i�O}2\�����B.eiJ��C��(s"f=�u@���Mk�(A�<)M>э�D�'��ٺ�ŕ
p<�C��ؿyv��&�eӊ�d�OT����~Ӕ��'p�I�d��(h��9��Nވ���']�oZ����ğ�`{��?Q��?!6�؇�T|�A���=xe" G(Z���'ǒQ�̧>�-OL�D�<������/Wa�TX�K��P}���~}Ҧ�/�y��'F��'^�T>�ɧl~�Iڂ!�,"��P��q���?��d�<����D�O����O�D��!�!�I	�Ꮀf�	z"N��M�$�<����?����d\�����'v�:�@�������jP.^.`�ylZey�'��	���I�$�5"n�H���:;���tF�Vs���c�S�Ms��?���?�+OF��1�k���'O��k���a'D+SP�q�lA��E��Sy��'
�'�Q�'*�L����MR��ÃZTd�o�ΟD�	{y�	s�t��?���J�cӶN�,�p F�{D9
'F��/��	ǟ��	����%`:���TK�>Q� ��D�
�.�B�J0�M�/O��Qe��צ��������?]�O��_
j �$� s,�[n���v�'��*���Ģ<��4b5<j���B�/d.Mj�"���M+���g{���'���'��t�>�,O�᱔Η!d�t� g��{���Ұ���	5lx�D'���J��|��9��ղD(Lm� �ż73�@�i��'r��74�������O��	 =�&P�l�+&�Z�لNW�J�7M�O��a���S��'8"�'�&d��'��^ e��cC6�I�y���dϽG��a�'��ƟX�'�Zc���#*ړw�8����"&J� ޴�?qr-�<,O����O�d�<�7.���H���`���҃�L�v[� �'{�\�$��П����L6�J�!M��"��GV���r�8�'+��'��X�hHrEE ���*>{d�1�D�N��P���M�/O ��<���?��k�Y�'��j�iգ&���֨5<r�4�?����?�����*�	�O�Z� �9@eI�Xx��w�ZRN�\B�if"Z���	П��I �6�	k�t��<4崔K��\�c �!*��4HZ�6�O��$�<��f_�Y�O���O��$ˣ���s�~���M=(�8<+v�*�D�OD��0��3�Ĵ?�'�CU��w̕�&l���j���%����i��'�?��f�	�*��qIe�W��\a���_-ev6m�O��FXz��#��=��2�2�I�^� b�V�.��K��i�Avf~�����OZ�$��>�'���	�L_��2ԏ�c��Ms!Kl*�EsߴJƢ������O���z�ܘ�p�9��lb�)�!P�6�O���O��r�B��?y�'ufA�kJ-xD�y���%|��Qش��F��\�����d�Oh���Ok,O�:����� ��Ђwj1{R���'j�5X�/3�D�O��<�������y?tI[�lէL��+��S}H&J��T���IꟄ�IRyb��P-R4�2�7[fحB�'?{l�UM%��Ɵ'����Ɵ��� 1C�8�wi/sX�a��Ӯ�$�	Jy��'���')�	4CF8M��O"8Hx�+[��3'	�G,�U�O2�d�O�O0�D�O$]��:O ��Gl��*��P�R83��ԙ0K[y}�'�b�'��I'2��O|���I� O6 
%&ι��l�Q�&�'��'M�'��Qy�'7�hd-� �(��)Q�fד\�̡n����I{y�o��4Z�~��D-��*!b`�y� N�\y��L}�	⟼�ɫ "��IM�	YJ�f^ E0��ӱ"�6��P;���ɗ'����7�z��i�O�r�O��QPp}z

C���(B�õ#��mZ�d�����|�	c�I~ܧc��"ĺl�b�81F�8\�mZ�
1�I"�4�?����?	�'5�O����Ğ3f����)
,RLɪ�oOަق�	z�P%������i�2}�6���	����
�9�ҩ��i�"�'����5��O$�D�O8�I�%�r$�e�Z%�8�p6N��L��70�$O�J��'>I��՟t�I�  �xd�Q�Ҽ�B��_A2���4�?�֬�+^�On��(���މ�,�(.� eH�)�����[��딨��X�'���'rU�P�R'4��s%�K���2�$�:J/�p[K<���hOV�	.���R,M���D&7��O���?����?�.O����(�|��K�7������/���$@�a}��'ў��'�2�E'\�a�J�_�4|��@�[$���?	���?)��?15l¯��	�OFH�h�%x��"لx�X%`�H�囹�	K��؟��'6�9@H<	��	�8��J�-߀@@\0'����!�I����'��YP�!�I�O���~�<T�ł'���D݀�x o�G��D|��F����M{U,�V[��p��33"0!���IЦ������I����I}~�'��ƨ� �`�!�b�8��թr��!P�i2T�h�b�>�S⓪q��=iҏ�v�`PfJu���u�.������I۟d���?�#�O��C����W����cI�9=uR�궺i�lXB�'w�'����Ě>�$(��
c}�1��L�AP�l�џ�I��@�$!�.���<���~�+B�j��iP�K����-����MK���?Y��!-"e�S�t�'T2�' ��J�$�".X��^	�v	C�`Ә��Ȳ
 ��'��ɟL�'Zc��	��ɖq1�4 �AJ+z��p�Ot(�7OD�$�O��d�O��d�<9c��9��93L�Ɂ9e�@��S�@�'��\�D�Iܟ��I�)���77!]�8�R�
5v�,��@(?a���?���?�.O�-:u��x��[:r,vݠ��/���(uc|�2˓�?A,O0���O��������=��8(��NH*�PB��'Y�7-�O����O���<I��Z$aM��ԟ�X���<��'8,nxҗH݂	�7�Oz��?Q���?����<i,��Ơ�o�H)v��>5&=��IƊ�M���?�/O4��FQw�$�'�"�Or���s,�s^\+���NӪB���>����?���aFR@̓��9O���#z$�:d�X�.	�l�����{4�6m�<�NY7)N���'pr�'S����>�;"� as��6+40��jZ�@�b�mZ䟔�	5(%4�	�L��ȟd�}bQ���sH���K
�_��	I&�Ԧq�����M����?����^��'U$} ��Z4�)aSU�tx8t#k�H\+�4O`�D�<ш���'��uBC����ϗ+Gctq�A�h�����O��d҉7X�'�������|} ��W��$�~�. %�nZ�\�	�<�0�m��?A���?���Q[�IĬ�;(�@��ܖB%�v�'s�0r��>q,O$�d�<y��;#�Ʒ"b�ݛ��L%	�X ��Ħ����i�����x��ݟ��	͟�OV��P\3$j<;�	џ
�(Z��ͣ
��'���'�r�|��'���N�?��XӨ�	&s�(�bAd���������O�d�O��;U q8�,�0!ȆU�����c���JDW���	�T�	b���x��O|XmzP]27���	Mh� @�O���O��$�O4�$ծ`���'�~���l�,�������]��j��M������?�/O�=#�xR�U]e ]��훍�r�R��ϸe�� ���6�g?�D�U!8��(wkX���B�<Q��5�`�y�k�*�XL�!倷I�*��,X��G >&(�P����Ź�I�;��� ���1F�� �d5J�wx5��B�.9D��BAk�\�P� X>��t�QEL�'9<�P�L�	/�U# �I�a��S@D�f�V��3s��A�d�7I�<ᐦ�Pg�����H1n�zn%\�Żr��Op��O����Һ�A�L�D��g���d��J��-����w�ɃLa,���MI+y��̢��t�$}rk2����OO�Z�F�W2Hت���M�:�X���dt����ԧթ�N��#�F��0EJhRIfFQ�%cl��I`~⬌��?�'�hOB���N3Kaj���ϒt�8tC�"O@)���2B�uR�A� k��d�Œ�����?��'MXI����z,X!� K�@3����F@���\���'*��'y���5��Ο��')���x�eI8tvx8e��DS�6d� 7�8rd%΋1a{ˇu�B����P�bZ��J#����0��6)Nq!E#2lO81��a�
$�b�S��?G�F-.9�'�ў\�?Y�&�Q����#]�aP��-Uh�<�Qh\�^�s���s���c�\̓b��Iy��]8!�듊?Y,F[�D��38��cH��?���>Y��c���?��O�ܡ`�51U����~2 V�ZYr��A��)�"��r��(�p<I��I�0=��c�i��$U�]��䂁�L�ngج2��K�?��x�k6�?�����F9op��q�H���c��1�1O���D�/P=Z������c3����ˢq!�HЦ��gOG�.Z�	��$3����Үr�Е'�l�$B�>�����	�3���$ݪ3�4�ZFY�$��% �,������h�a"-3N��"�b��|R-�RA�GI�z��iSn�
kIH�>�! ��{�����2�Q?I�gW��Q�)�4	� ١�4}�fS��?���h�(�$S�4�jp�0l�=S��B�Q�L�!��",����j�4���6�ax��9�a.�qhv<P��ąo�� �Z�(���(�6���J<���	�����Ɵ�]+,*(%�[���3�O�R�,󡣛b.�d��[��S��k�g�ɛ=��A�#6>[0 �n�Kuz �Т��tT���9���·�#�3�D�H
V4�_1��́$�B�$3?�3I��j�'s8��X��@9g=j��@�'��,IV&I	��f�[(l�p���O�Fzʟ~�]G�T �-�YA��a��3o=~0�RG�p������?����?��d���O��ӍRMT��0h��J$R��2�8��`h�)<�樀����
E
S�'.(Jao�84(��&׻2�0�@�%!��B�'�"�)B8�D{C��)a���^p��d��^<dB"�O��n��M3�Z��O?ʰ�d���Z\����k_���(�'��0`L0�(;���GnB q�y"�>i-O yq��������l��"K��@�E/a�ƀ��aQ؟0��&7^��I���I�b����r��S�" � �\ݟP��ğ5\��p���1$�ؠ��:O��G���zع�D,j���P4i�<<���0l����X�y�ax��ǐ�?������'�~eJ�FZ*P&�;}����X�@�	^�S�O"�H��)F,mn����2K:4�:�)�nC��� Ir,����Ӛ([G��0rb��R�'�0\r���5�`�����oD�x�	�'�h���AH8#���)4G�vW��9	�'���H�M�{���/�q�@�J	�'�B�@�*�us4dn[$I�'p�����0�R�	␎_2Di��'tN�*e��8!lAy���'�����'0�t�7MD���J܅i��A�'��"��Ȟt��UZS��0I/�E��'׺4G�U 2��}���'.%z]��'�lb�딠php�B⃳[wl=��'���H�Rh��B�֝&�ڵ�
�'7��H�Oa��y�˸o�Ѹ
�'��tCB�ՖI&,�U���7Aj-�
�'X�x�Q=S�թ��Q�)h&$�
�'�(�Q�$S�{��e�
�t�L)�
�'����.[&N����5Cx��
�' ��M�#d`Pd)զ�"����	�' �JD����1���"V��j
�'M��F�X�PlH���[	n%�	�'l�������.I�U�ؕ%;F��	�'�%�lV7L�T�K��'0"8�B	�'��� '�A�8a�h2	�-������� ��U��ᶝ9F韢^UV�ٔ"O.��%�2I���(�+5:� K�"OT�s��H�a���7�
�e�LY`4"O�9(@�S5\�xm��&S�Da�Dq&"OPK��Ĳ8i�����zEjl��"O��Y��4]�z�)���/d�1v"OR��ak������#H(`���"O�*�F	�=��8��Q	��Q"O���Kyv�Lz1j�w�*�*&"O��Z�O�L� �q	āb�(y��"O�9Un�-g�F�B��ڢ2�8�H�"Oj@�2�-&�Z��B�9��\�c"O�Y�� W�D?lA��[��pl1""Oj��qX�7-�E�敕��&"O�|r�i%j�<D�T���pxH)`E"O&i�F� wL}#R��jv���"O��Ju�E�a傀�cO�)3H���"O<��W��;8ȓ ����h�#"O�����ۄN"���.V�n�M�"OJ��&� 3C��;�,!Ｙ�p"O�H�a�����؀�Fmچ�3&"Oz0��i	.b|��R!�9a����"OD Itł�qe�� �_�N	�"O�H$���7K��j�"T�C.p��"O��p'	W(��	a�\=�Q3p"O�Y[Ю�j�qjP���O��S	�'���I#
ր�h���1�Y��'�p�Q���i�J��@�&��1c�'0�d(�'���`(@�,!�Pc�'�2%��
*s�DQ� �������'}������=�G�?
��8�
�'�䅠��Ʈe�T�bE��(�	�'Z�e��L�1V
բ!�+dѺ�	�'�6��ql	������ǒlN�@��'�\LcedJ�+:�9��ٻfzjȈ�'w(�����JZ^�sꋐ]�:�;�'o�
QGӢ��Q��ڞBJ�k�'Hx2���|-j�A2��7�P���'FP��D�@�3�Rę�&)^:<�	�'������ 4��0��U=��(	�'��hVŝ,��	@�"�P��-S	�'� c�M�)����,�=x��q	�'���0߰1�:��bE�u��8��'|X�ni��]9�+тu��(i�'A��+f��0v�є"�&W(Y�'���Y7.L�]�(�E�7p��'f����Mئ0=�P�ʓ�2�H[�'Q8��f�V��ա%�K5-����'֒�aǂ�_�H�T�ƹ�[�'��ݰG��C����eZ%F_\q��'.�]���:N�~!c5�L�-�Ȍ�b�ԱO��}�u[���x�FA��]�4���ȓX-�!Ѓ��R�x����D��t�	 5�h��'x���5�B:��MH�%G�"Xp�ߓ@Rbti�>yP�ƁIc\�z���/Z��qj��<��W�v�JĘSʕ6����T����r�6�����Z8��ٔL�pB�f�>���1<�M�6DͰ<^f��il�#<E���A$�j����["xPB�`b�
�y"&�s80�b��;u�|���<���V�D���=!�F��Fd���1O�'m���D 5��6-B�F>���C,Q#=�}�P���X?!��D�<A�P+�C��@6 E9#�+f-^���$	�60�	7R�J��S��F�J��`P����mF~SF��rb �5�RB�)� �M1gb�Oi�8{��@�B�q3B�w.f������
1��7턥0w��S�T�ć��e�ꍩ&�L9y�M�"�0=)u�Uz����&e�<�#.X�b ـ��A
�+BNI<b��$�M�`X�T��'��'Y�X�Pd_�zI~�c�DԶo�y2Dմk������yZw@"�Q�(�a��pz�I�1�Na�'R�Z $�Z�a��<G� )�F�7]���s1bܨ{C��3��0kn�U����|�n݊17���d 4$��bq蚓B���P̞���\��e�2c��;���:!��V�(�� Q+7^0H�3H�<i#�
-̒�q�	;}ʟ�Aj .�U�\�`�˨Y���w�'��}�Ee�.Y��{�'D�]HaBO�!�����M����[D�Ƶp�d�X$�Ο���������r�H�k�&[6p�u��O\��<����KT�cw�E~�OH�A#�?�dD�\[�,=9`��,����C^81ZT���*\O�� ы��	c5�FQ��3i�- ��Ǟ����
�?��CF���U3�E3Pf�စ�l]2����Zƌ�� 
[u!��ȃ@����/�e�A��Fff�H�I?z�⠻���m/��b��г v���44��b>������q�4M�sL��c)�Y���*LO6�y���B`��i��<A���kbv! 0P�tU�'+t�hi�jނp�b7퍎j��ea��L>y�,��b,��ۮQ����X̓Ӿq�w�ݚ#'H�E��<9wHݣ�!Hb΄�1ꌊܒ�w���E#�@P!#����Q)�����E��IvL��`ޕ7�ay2o�$��'jٌK�n8(a��O3x�h�c'8a�,�Vo��o�PC�	�2w��#(�uXxؔd=bO���!�z�� W��w��|��B
�j�E�>L:�)AdWT�<ɗ���&,��vY�u�ĸ�F�ø<y(9Ke�B8)���)D<���O�� E燸>M4��.ֱ
��]��O�!��m��1��un �T��*ԨZ:$r��n��+5�a��qr�CW�Y��&X�4�L�( �=�O�M0񫐀7��7��9��v�V)>��	���M�!�<v#V `�V ;����f
4i�!�dD+hd��*�@�U��u�%���!�U��.� �K��/������+{!򄗘-y��j�׵I�px���=!����bx2�F&h"���<A�!�B�K�@�Uf�-KtƐp� *J!��y`x�"O̣UO�wi!�ۨu��V�*
\��⣮�@[!�7� }x�L�&mʥ3d��ZR!���b�BS�"giP���E�@@!�>hB��b`�6o�f�!6e\3�!�	.�~�e��(תuq���C�!�䅟��c!*C1Ŝ ��O�%�!��-�(h���X��z�!��C�!�)��}E	 }Ha�`R�5�!�D˟]R�H�&� Vp7 �\u!�$�({�l�� k��a�@�C ݂7�!�sA^8�t�;{l�p�8%�Ę�G�����"6ި�X'ڕR��|{��]l*�����B�f��]�unE9|ڍ�3��(m�݇ȓ7��"�������'���Gy�ν?��~�G`�-ö�)!ˈ?%^�T��}�<qWF/G0)��!�/^`�]�k8w�pİ�2�)��t�el�?m5�ɘR┝A@��٣�7D�hS� ^jL�Z��H�T!��>���pX�xǌ��X�Ȩ�peE 1���K1D���  F�r�+�z|<�b�*D��3a�p+�-Q��
X8�&D�� @۝-�j��ÀE�L�@��)�<���A��(�vI�BY�x*�C�"�G	�5B�"O֡@p �=4|I��	�}���|r�az�g֪(|H
2
�b��ٙG����?�Tgר�a���xip:���h�(dy�'��	���=�j$a4F,�����$�N�"|J�ºi;��bC�[(� *o�<Q�m����T蕉�P,P�.^myҡV$Vl�OQ>� �-��IW�22�p%��\X�1�"O�m1��S����νT����3�|b�ϿP�az"��u̪���e�$KlpxZ�h��p>�aiĠxv�)f���ճ�O�+�Eyq�P)�hC�I;OC��)c,E+]��M��NS�x��<��o@9KK�#~:s卆n��E��l;#�Bp!��Z�<�@
�U�<���GE6�I$E����h�S��?��҃W|�qt�4��\��)�U�<���0B�6�MF�]S�M��N?�6�i:����@�<�"��D���f���9�e�c��|"���a{�!�J򐁘�n�@1^�����Ia�)��O����F2DWN�K���?��Fy�k@*K��9E��
e-�y�@�x{�@{҇[�y�Ô3Q},�2(P2?��R#ƿD8\SU��������yЎM�@��<�ޥ2V΅�y
D�m�$(F�%%� �IHS�~2%@3v@>	��	@ �҆H�]��Xi�-��at���Z	��Γ0�"�KW���zȬ8�'�>�ȓ ���#��M���sn��tٰ�����@wo��t��F�Ɲ�F݅ȓ1)�����C˖�ڹ�ȓ����@I�� ���v �6�jT�ȓi3(�PuEY͢U��@:
H^܄ȓ�8T�[�\������Ya�*�ȓ(�����C�i<�p7F	c��X��T�4���cۛO�rQKƎc|l��$Ӽ�;�ۀq�L���oۉ9�NɄ�;i�XG���+'~yY�@�C�~��	
����(~�����/lF�M�ȓe����'��3xwb�ڴ�)8s�ąȓ{�6�E�j�L ���ŦH!��ȓe�� �CK�6��������=�u�ȓ6^>xbp�S�<�~Iі딌Fӎ}�ȓj\��CdR�D�<�����k��M��C�`��U�;��HVČ�����k�5�p/�U��P#���rt��4�� �E_�7آ���~kȆȓ@�R��g��(8!X�۱f�Ԇ�&e�5���J��|�Go_9��(��v�ث�)��k/�a��$��g���/�����@_�lQ��_�} 4���-����r�0Q;|��v'�?aDzхȓkKМ0�/�3���&tK.��'��0���S�}Zȕ��Jĵdm��
�']���/� ���� I �ia�'�"D�` #���'L#=O�!J�'/n(�T�X�O'��i�1����
�'b��Q!�����s��t����'`dj�D�� �.ա�� A�P���''Α��✤g��Qyi]�4�~�	�'D�0�d�)6$b,K�����
�'ˮ8b�C�>�$!��샪9�5�
�'�:1s)�:��5:�H��z3ܝ*
�'_�;go�w��]`�Ȉ.v�4ܸ	�'tXt�r-C0m�x́�ǒ�W!�"	�'���� ,��������R����'褂G��^�θ����-7P4��'�:y��P8z)��Z0腧1�
�[�'5��[�*�#[�8=�P�]�'O�D�
�'��$�Ŋ)A� �1U� 
�'�45KA�(0�ƌ�BREy�'p ]�S'H0#=r�2GU�!|���'BP��ŀ3�!�4"W�I��Pp
�'=PjF�U���0y5�
>W��	��� ���e�0D��|Y� �2EOjeʗ"O�}��^c�<D�c���;F=�"O�� �ě��H��?>*T��"O<Lw�E	U��3j�O7��a "O�����6�L=r�"d"T�JT"O��
&A�9��mau�T��5"O��YǎR�T �ye�	�N����"O��Se�D�c��Y�a�\�Υp'"O����jՃlI
4�ѭZ���٩�"O�����lS4�5�ٳ<K���U"O^�CЄI��\��+[7iE,D��"O��	�G"�����za�cd"O^h�� Q�(HV&�- �~�[`��'\O�e0�G��qޚa��{j2̈�"O�, f�ѵE�d	B���4=1R!��"O�8�_=^wHa�0͈'8A&�a"O�e&" 5׾�1���.q0L�{2"O<�a�eޏIPd�@@�f�2��"O:m��́N�it��`R�`��"O蝉r۱h��a�!�k@`���"O&e��Z�y���bF���vPA�"O�����.e��ٙ&,H�}��]!"O���b.A�I.�����zԩ��"O�E����4�@]�beR1<S�A!�"O��`D솱K�2��EØ}>�X��"O\}�dn�(<�6��ׄ��a9"O����V6rV�sAᗴQ'���a"Oz�ڕj��L���J�3��=b0"Ot��0ivt�H�>s�L0��"O�A1(݈�V `�'K�^�8��S"O`!��Ϙ�,R�W&�����"O��R1�@�$(�h7��}�¤A`"O$]�RC	?MD	��j+&�<���"O��(抝j���2NʐHo�S�|��'N�,�rH�� Ռe��Q4Gz��R	�'Kby�V�.x�2��F�u��': 5�Ƅ5-�h�;��F-��h
�'LZřW &;�@|�Ag�69�&%[
�'��,�Qn��&�{2a/xj�s�'��dqR�#`�hE�W�v5����'!F��G AB����'��|�v:�'�1�6��#���b��JVUx�'ɸ9PA㛪0�RI�ƾS���' �L�pn�R !y�·BZ`���'� �+� ��5, �J�NT0=���
�'LIbg$�r�H�R,Æ6K��1	�'V���A"k�2@���I�)v��'S�M������4:�+l�XY	�'k����o�&�����e�F�:�'�PqhUi²{ҔM
GkЏdv|t��'���t�T�wL��BC��Q
�`
�'u��!�*wl�B��4�as�'E�4��j�	�C��К��	�'������Y	��`�Z��'�:Ydͭ���f����x�'Hp��t���V'/�T��'%zD�`�	Z����E	,�4q�	�'��ݑ�	�<>s�� ����RXB��'����KW�q�������= DYI	�'��x���
x7
�(Z!(�����'F}�F�O�\{���a�!w���'��d����#����!A
�~Z�;�OX�=E���.��d�=���@I���y�I�Y����u�[Ø͢`�ͽ�y
� ���hJ�7<X��H�=�(z"O$�:EAI�tuq���(a2��"OF�i!!"l꼊���;��Y�"O&���ŔC���/T5u& ��6"O�`0u�J�X���#��O�f�p"O� ���%\�<��Ű�����"Oz��g1�(�*��X=��"O4� m�2p�~�!5�4�����"O>�y�F�$(wp��Q��-Iex���"Od��� �~�ZE� )(��u"O�T�5c�!��I
�7,k��"O�\�R�j���jA�SO����"O�|�4�O� qP�����9H8�X�"O�iW
�����$	F-�4�V"O�
�%ՉW�Yi$I��ʈ��"OR��f.8�(c&K�ռ: "O�Xqs�[�x���p�'��n��"O<1C�=�LES�e�:�r��0�'��d�s����H@����e	ر,�!��js��9���v�b���
H�!�DB�7X����ߴ�ڴ�`�D6n�!�W <��a�4� "-���b�fV�]!���"�e3�l�**��]c�oQ�d�!�d�"5�2����-E�5��^�!�$�!�:�A�1L��1��̝�[�!��	Y��X���(<��HR��,�!� \��X��äG�MK�l�-�!�$J��Z��Zy�8(�Gl p!�DB8��)aRF��@F�i�5"O@=򒏎4	��2�cƓW��)S"O�80�]�S澙k��"H���@"ODE!�xV�ԉ A��E�"O�а�F��O�<�F�&a��jS"OL���J4s�I�X�O�N���"OʴY7��'Y�܁�D�\|�s"O�8���?v��H�A����l�T"O(�:�7'^X]� ��|(t��"O�ܰ���F�p!a�OZ4yJ)�3"O�Ԛ��X�i
]�!��X�@%S"O��s�$у'dvŀ'������"ON�w��9u	�1���j<"l�"O�0䯘40z�J�A;- ���"O���&c���t�7-*�17"Oؔx2�ޣP�6���w�|�'"OLI ��1]�Ehg�݉`I��&"O��A�����Ŀp6Q�2"Of��J�0S��P�p�\�k��q"O̝�Vd"��E$��}�2}�$"O�9�fO��B �h{Ě����d"O\#��PS��Ԋ�_�w��h�"Op<A5"@ j3�4b㖔I��A1"O�8���V� �G�^qn0�V"O����H6)���`��f`���"O>�3�A>M�>y����N$
��"O�� A�a
�Q���.KXY�Q"OND�4 ��	?��Q3�T�@,;�"O��V�z� A1��Եc��`P�"O��+�\eXU����z�Ir"O��Ɵ(O�ҍ�L#4]Zd"O��ώ�Uh�vꄖP����"O0l��U.�NaZ#�@*P���q�"O�p󦄱È��!�]!yz�Җ"O2h�CԊIyl9؅�_>peu�w"OH��A�۞�,�ѤCH�K���S�"O� L�q��ڷ|/9���_�	�F��"O�%ꃤY��)�J4q���h"O�E���3���K�A�8n�����"O�!� �-����"��)���(�"On|X�%�U�BH3W�K�nq��"O�i������ZvⅤO�$�"O&�5C�1t	�@AUvd���	w>�d�@��%5
�Us6�8D���!�X�d�ցذ7QjA��(D�80�d*PV^-y���0##D·�'D����ř8i@��B�L�V�0�B�m$D�[U�Z�0�v]P���2 ��G/-D�0�� P=h�b��
�a���sr$�<��2�8���#Qt�Q�W�\O��Y��^�Jl{eKa���nY����ȓ8 �a3�L?F�\�b�Ӗ[��Ey�'m)0�F�$ �̐fd�5;��-��'�8��d��5'���	q_�,�`y��'���F��E2���������'���C�&����I�0h(��ȓH�t���/en��@d� n5����F[P0��%^1��K1(:X�%�ȓ �BH:.�i<.�*�o� �̆ȓ���Sțy(PL
0���]��܇�IY���F�>�l���Ȣv��5��|5p�)� 6�Z,����Q�Pe�ȓr��+Ƃ�*?̎a;u�ҕ<�ȓMGP��*YoZl����B]��ȓ>t!���h �����HX��L��^�{�A���D�R��	 �P��"�$�j�$�~;>M*um�B�ć�p�I)����o�
����,H�1�ȓ~c�i�DT�9p�5��-�(YM�Q��q�Qx����'�����$��ȓ��e�S�J<tn�:�D
 �x��!�H�B�.��M�6�ѧH>����{����A�`��� b��Q6n���c�Tuf���y���㗩_�L�0 ��F4�qJ�O�Ų�����T�����p����t�R�ӫA��ȓ.�"Lr�@�B�`� G���"O��Xw��-XD呡0��"Ovqs��� 2'|x��ㅊ/ R`�"O�Tr�Iʬ�yK�(3W��a�s"O�Y��N1)���ÈO�vp�lh�"O�YAV�˜9�����B�}�=k1"O����7�vD)��Y
cy�|��"OFMу�	���83tG׮`���"Oh	HP�:5j�Lz3�W�1�"Of]+t��W	F9���119�DI@"O( !fO�f��\��fـQ#�l;�"O�ur�bI�|I�_iz"���@�~�<��έQ@�CS��c��U�y�<�p$�^����M@�\�`���<i���t���FB�.Ȅ�;"FAw�<��ʔ
/}䘊1��1����aw�<Y�-�3�|���F��  t�CC�x�<�U �p�a�e�Q��dQf-�_�<�b&����v�&i��h��^X�<��O��'��y b����D� m�N�<)`�E�lҢLҼDΉ�&hKL�<�F���3j|�,B�JE���t�XK�<��CR@nY�q&�/^�}q�&UD�<!p�P�*7���D5Gɂ��T�<� n;U&���dKN�\Z"Or�+��F�A�׈�e�ܘ�"O8�rF�ܤ��y(�铖hET�!p"O��tM�:a�ə0H��6�,��"O�Q�p%.y�V=ѵG��W<�`��"OƁÇK(.����i2a+"O ��`΍����1�E��LѪ "O�Z��i��M�&%H1S�����"OB��"��=jn���c��Sx
dxq"O�ܒ5�ˍ:4
,;�=hgH�Q�"O��U��.$�4��sOR�C"O���ǘ.b���W�Ѧ,9��
D"OBⅫ���q�@�X�0�r"O��ā+� pD�N;X:�I"O�zu�X�;d&��ԃI<`_�L��"O�L
e������)S$�w�L��G"O>8BU))�
$zc
��$��"O\Hsb�K�5H(Fc�r��8A"O�ݩ���ua<�) F;.��$�a"On�!��߸?�>EѠ$�A�0h�"O�E�' �9���Kb҇Vrlc1"O��z��	[j���K�5ߤ���"O:t��cId�3�̕b�\[�"O��h�
Z^l8�"(^8:�D��"O|`��N��KEʐ���X�8v`��S"O~�1g���Ie�ћfM�hl�ɷ"O,�����qtиsG�Nfh�X�""O&�(e��*N��J�뇤-C��ф"O
����5N>�aC�+A
���"O扂�Ï/׀��`�[�5'.$�V"ONx� ���裂5.
� )7"O�l��^33�8��G��<�
�"Oxu����%�|��f/I�8��A!�"O̰�a�'n\��E@��i���"O�-
����2d��".�$P�x(��"O�@+�:j���-�:~@0�a"O����׬K)Xi����yL�z�"O,Y�ѩ�k�<���ъxtl-[�"O&РE��7B��}zal՛&��j�"O>�`3�/	�&E*W�Ë>�b9q�"O&�)�R�#���BP�ۂ&��ag"O�`����6��AX�i7oh�@�f"O�;��
#d. �#K��=q uR"O"�c7�Ҟp~�cf�LP�u��"O蕛��B�~�<xrOG�j7@��"O�:��p�D�s�L˿�9��"O����,P k%�߸u�@�"OX��"L /L�ꤤK�&� 6"O�08V��T��
b����@�"OL���o���=ɶhD�~:(�w"O8I�g]:M�%�3JD�G��P1"O�@Q�D�B�����U ��Mz�"O.D��Kݮ'����A�ĭy0J)��"OTix�ַSgV��H/,��q"O�q�F�(w�]���5E�l
�"O\�zW&R�V��yP(�*u�|��w"OJ�;SN�J%�rM�Uì]��"O m��֧XL��c�L�G�p�%"O|� T�D�����B���by���"O�L�G�o ,�0%1QJ�ذ�"O��d�)B�12S����0"OR�@��Н�������5k|m�"O������*	Ԩ*���7�	�"Oz��Co�#8�|�q Ǜ�Z�"O� h{��O49 *��ю��+U�5"O��3����5��aP� B���"O�pS���$f�6ᇢr�z���"O��%�����B@G�?�fii�"O�Q��cJ�C��ŲF��\�3"OQB�9�d�pDP�	x�"O�L�b�5(Z�0@��
�@޼d{S"O�y�7o�2�l�K���	�2��"O��z��K��ug.�E�P\:P"O�E��� F�Cs��8��= a"OB��$�^<pӠ�F�G�z�f�p�"OnP�1��(ut���Hօ%��a��"O\��$��2������S�4��t��"O$��lӏ&�P��g"p�L��a"O��Q3��7f(`+���H�t%��"O�Ȋ�+�*N����	4Y$�ˤ"O��#�bD9;���-�)TR�i�"O�y3yf�&��BV`��'"O��0G�E�I Pp.W.W��f"OL�Q(��l�D��L=C��!I�"O�M�u��ÌP*�
�% �1r�"Oxh
�<�J4����|�-3A"O~%)����%�dZ7$�Hm��"O69K�&
M21!�g�C�,�Ze"O>|�	^U�<�`W�[�l�&"O�=��" ���C�O�;�B�Q�"O� BeÏ�b��(�tO��f����0"O`�i6�T�\�􎌱z���Y�"O�M�
�u�X����#:zh8�T"O�}*�M�K#�5����5lR�[�"Ov!C G͟g=�}�Dm��8\["O��RW+JL&���Eհ0����#"O�-����Aw�R�yL�3"O �PD#ʝ|~���������"O��"��Y�]3P1f�#_�n�i"O,�)��($����I�5� �F"O� �%�	w����7�U�&�p��"OnpeA��Y����O��z2A�5"O��5���j���Gom*,cp"O� �˙5x�L�b���g�4hP"O���"�V.L1�#�� �"��"O�Ԋ��Z)}A�0w�Zy�����"O����M����HTo�#3��a�"OR H��z��.��h���v"Oޑ�4�
�V�-��Ȕp|���"O(,���ߧ@�B��g�2cHd0Q"O��a�b�6[M R�P�[@}��"O����ǵw�6U��@0Y:tt;"O2)@gTؠ"b�ˢw5B	��"Ohh�$� �a����mT���"O�����L�L1rԘ5'W?AVM��"O���"l˼n���!q���c/�U@"O����H����I��޽lЀY�"Ob+�@��!����
ЮA��YI�"O@��'F����T�ߌ4T�bR"O� �kȥL�r$�����p��"O��c�X/2����CU��m�"O>)��B���*���"�4fr���"O��oD�:ص1w	�rXj�>i�IS��|ad�M*6����ŝ)�� E"D�@�(J�4�6u�d�L�1�1�>D�Pa�.�wr��s�V?_T='%)D��	���#?d}14"Ԉ҄ :�;D�$��b��u.�4�g��N�Z�{���<		�S�? 0iy�O4=6���qޱf�9�"OV�KG��+�@� �<-����P�8�IS�T�����(�/P�Ca����F�<I��0>YG��� �̅A�H'z����VT�<) ';Xn�`��k��c�� zG�L�<�g��3p#^!ѥ��	F�1`7��G�<���I@n ��c�(o�	����yR�'5���� 4=\[���J����' 4��'y8��R�E4�=�N>1���!�ɏx>�ۑ�6}�M�תP�c՞��0?�Cm�$w�*u�="���Aa�{�<�DB,L�`��h3�X���
�y�<�%��/z��@�
�	g�|��Ks�<Q6o��*�μR�[�Z����`ipy��'}:�z�/Y�I�狹\z��ϓ�?�yBJC.X]��C�U�H�Ȩ�5�B��yrd�������<�B�����y��O?�ޥ��
�
D��
�_��ybM�G�R@ئ��/5��eH�@��y�)�.%�9�DJ�>�bD��JP��y�Iݑ� �3�ʜ ���@sǞ�y��*V 4d (	 n���j����=1�yB!�?k��ܒs)�"q� ÎE9�y�,��~�g��. =������yBA�;^��*A(��9S���y↖[���a�r�l@h�,O��y2�G�\�$��AE�u� �!M��y2cϮv��r�(`� ����%�y�A����s��ˊp3 �rtg��y�o�dA�F�=l]<����y�%"R�PH �OT=4w���eF��yDD��<���)0S���և;�y��]�(a`�+ǋٙ"��{&!ɥ�yb�w,$B�`(x�����&�y�̅�>.F�y�%�%��I�,�y"L��?��!��텨'{�d�U�#�y"���b]�:�/L:"��Se��y��ܣax����G"��H0��G��y2�G0-H����m�A�8�yrNM�_��B�+�*=uP������yb��k�ܤ+�eU�:` ��T�yR�݂mb�y�HN�.�\�"��4�yB�)�%��}�rE@u��gn0��V) �F� RPcy��'D.ړ��OFu�f%՝dD�H���A����se(D�,:��L�p������a7�&D�P�R�H<�`2m�6�tRGi?D�[�Ḧ́W^0Sv�5ZN��4?D��9ֆ��I�$h��`U�,&R��<D�,�/-B��쑱{.$���O>D�x�s���d����sN�Q�R�h�"4��SVNKRT�v�E�|Ʈ� a�� ��Z�T<�F߯ �(hфW!`5��1[>`r0�Y�(�@e��;+YD	��gϾ0�S �;�ʵAą�X�2U��>�����I�~��eIfk�~� a��_b1�2�T�|����sLyZz	�'|ў�|Ҥ���L�p�RN�e��aC�X�<��H�$���B�3(*Y`vB�Y�<��cC�5��ЦWyƵq��W�<�se�X\4�8v(�$)yx�DJ�Q�<٤�Q9W�
��$'��{�UM�<ٶ���bN�yѢ
��L�V�3"&�G�<�C�̠#�6l��N�\{S��y
� ���i�v�L�����qº�Xc"O�2�� 2#^���EV������"O���d@�$+��;�Du��H�"ON4���==m,������#�Ҵ�"O�Y8�LT� �^�X���}x��{G"O���S�Vt�ƽ8��<� �z�"O(��!nL�D�S�@V2�(e���X>18�	���Q��8!J�m{Tl9D��X앹 �T�3�ܝh����!D�Й
�t�^1���Vv�UrTh;D��X��T >5($��K� Op�ࡌ9D�4p m�T�,R�Y�>Ł�7D����C� 4����b�΃#v���� D��hT�ة@"�"��%qH���:�Iz���S�T���(�DÜb�m��D0�DC�I [�~}ɇ�0	=�m���Ϛj\�O�$*LONT��N��o����a"h��@g"O�CT�H/��*f�S:|��d�7"O~=�jɖ.
U
�o�IºE8�"O����T�Ej�i���$W%"�"O���eo�
h�plBrjO
�bPA�"O�L�q�X�1́�q*�'G� -a��'O��U��iyT�Q%/�b���ޣPS�'�a|2�w�C2�ζ`���dN��yrI۴QB� �!%�VB�����y��*z̒�K�,�"�����%#�y�R�gV(褉��fĒ�"!F��y��?�y�@,�sk֨c��y2�^�:���)�&�8_�	0P�[���x��my%��^���p���i=�B����Cl���DE�bO0
o���B!0D� �qJ&E��$�d��:�V�j�@*D�@:����'�\ ���<;�b7i3D��!��D� L%�"�3D�\^�L��0�`�<:�*TS0�1D�����3L� �j��\@*@0�1D��ba��!A<�ePDl�WchXdl!D��X e�(�"�R��[�$���SB5D�h��N�,I�D(G���Q�sv�2D�����#�aK(��q����E/D�h邍˪61 ɰ�.Z�BϖaѴ�7D���g�4B��Kc��N�$� �3|O���/?A �V� &P���0o�e��]L�<aq�Q�5[TD��#�D�Q&^C�<Y!�[e�r�AmΡ7��!��B�<i�˘�=�I:u�_����D�u�<�4��a<]�וfЂ��wĈJ�<1U(�Z�P|��*^�R�kժC�<��o۬	�|03'i��l�:���ȃ{�� �<	d�?(�up�$sv�@�b�v�<�&#��l9�B��
cB���X�<P�T�Bܼ��1��äYW�<1$�I�~C�Xsco�?C�49�e�O�<i�EÆ�X�����[
HIځ��M�<�#�S@��h��m���xp�d�Lh<�����=S���p	�? 
���j��y�dɏ|2��!嫖0/.Z�����yr�~ �`�"+�͢���yrOAW�>�(A*T���Q�W�y��>6tX1�m֐�aE*�y��:8��`q��Ѷ`RZ���y��'2��#�m�m0�)���ybU�i�jЀL>}���@ч�y/̿j��PP%��e��$Ku�� �y
� �4H!c�0i���4J��^1��"O��Q#�>D �qh�i�10a�%"O�`+���ӂH�f�=tLa�"OZ���0t]�H�S�5��ɘ"O��U��D��x)���w�vYӄ"O��T��%�m���	p޲ �"O��a�
x�����*�&��b"OY Ĩ	r>J%�'[�Y��"O��@q��cX1��U�(�lP�"Oʄ��$@	��J��u�Pc"O���� q��\1U�ຕ�V�<���H�"l��:�k͕j1��B�%U�<Y��M������C&ݬx�DO�4�y'<�!7�7��Ih��y�n�.$kШ��"�rK����yB%ȗkU�T��G� ��rO���y�D&Ѳܷ>(�
���yRc$J\v͒ yƝ�f�%�yR��v��q�b�ÌC.V�S���1�yBO	0��UZ�� S��yDK��y��3F:��xrh^�^̼�A����/�O:��n�?@xub�G��]rH���"Otk3��U���V����h"O�B���p��%�R�2�R�:B"O��hwAO"S�T�&
�W���"O�jD#Q v���f��x�)�"OꙺE���]HΡ�tJ3�����Ot��n_.�P��D*3��i�"�<��d2�ɦ|��� ��Ӭ)�ū�O�
�
B�	S����1�+7� b�3�4C�I%jqԴh"�\�*��Q�&H\'vdC�I�,&�t�1�]'شc�0�2D����
Q�`H G�C�{S�iՂ.D�@��[p��C�E9�P��&n:4��Vi��la�"!YBLh8������f̓n&̑��W�\~��F�YI�|��ȓ�!��OI�qO��i���&C>}��
�!)q!�i������ vw0��ȓ$��`�U�iC�=1P��4/��=��6┑kN�i,�jV�H�!ΆQ��an
p����tH����u@���:��mK�� �Ѳ*mӧ���ȓ.C����T�{Z�u%&(j�Շȓ%���"��+�H9x���tT���m�9�����1րp�kU1d�M��p������'|7J�)t�^Q���ȓ+� ��ڰ�zI�q�-YEb���צ���?V�j�h�![ࢴ����\aR瑫k0����SplT��X���h��D˒z|�-y�e�"M�=�㖉(��w��)��NQ����Z�F��2��0D�p:�LB	(�R�"e���-B5�1�+D��sv��.��@�W=Y�,����<D������:i��V;xa�4��<D�4��I#r���9���\���1��/D�L(��]�:���T�	�I��X�r/4��0<qd��(k|�3F��]@�PѦ�V�<IUL� °)���ȶ?(�*u+i�<Y���s�r@�D�1:��*��c�<q�H Lb`�hc'�u�\��2cX�<a�BF#@޲�C@ ;o�왢@�GP�<at�M%o$f���b��*��x��FJ�<�S��|՘���n�ub��M�<��Q�%�h� 1�^�I/މ*�B�s�<� ��STʋ��\ �T�U1� x5"O���1��\����tjX�cx� B"O��UI�Zk��'HX�z�"O|ti�>^k���kQ�4yW"O���ǅj��$s`N*EVl�$"OrxA�`�R���S�k4�dKp"O�`%`	��|��M���{���$LO�dQ����H&`�����"O���+x�"H��G�=p�^�3��2D���"�7�ux7/_/9n�bc�.D��r���%��q�Ă�2[��� D���5�,����g:�����3D�P�5���gz�}0�"U�����-�O�扟��M飢O�I"`��L�$��B�DLb!B�i:���ym�B䉅?6�I3	��2��}��$�<C��S���Q�ײ���H��E*�<C�I�Y����.A�@)���!∶v��C��x\>p�Xe����p��.��C�IcqZi ��M�?�x��h��f���'?qď�FP����3��A� H�N�<&��K!>��Ӫ��=Y�E��hBL�<���y*޵{�� (R��DCG�<镤W�~(���2���lw���CDx�X�'$�����wv�״Fc��a"Ob%���s�^���k��-HJ�;�"O�|h�"۹1���ҕkK�},�,R�"O��{V@ɴc�̑R2(��2�"O2:$� ��9b��ٛ<zn��2"OD=���ٰ}�tdԼI�|4�`"O!Ƞ�g�:1�1A>V"M�E�'���2Zz=���\ThRD�2�!��_O�t܀w�_	r�&�A5)�{����"՜�;��ؔ
%�D�R�e�!�$�:��%�b�ý=�.��.�!�H$c&Y���'݆@���F�!�
t�� �EHJ5Ҫm ŏ3T�!��GU�l2��G5O�z3-��*�!�F�k̀iCT�_4n��ɩ -�'k!�$R!��x���&��T�c,^ CN!�Č 5��[�g�VX�b�ģ�!�d@��;����y��i�� �@�!��S]�X�b�F�Kh���t�ǵ0�!򄓟#Sd�Qqoҗ|3���I�)!!�$�!.�DCSeX�3��� !��{J��jW�[t*ho)�"⟬E{J?�J�I�e�P�Ǡ�<۶�!D���V!������%JA�q�^=��� D��SvGY~�9��̞/��`�#)D�ĈQAQ<�� ���8c���t�*D��{g�  _r��˙�V��a�5a'D�	��B�C�z	�v/̞5ܐ�"�b:D�<r��7��Xs�`˳9ٌM2�A:���<��'`��Q�����q`�u��k�(#e�����Q��L͕p%*Śf��>�d�ȓs��QB����tI��웽�����KҖ�!@H�;j<�����L�P��ȓ5��5:��X�z�2���E'
|���Ӫ	P�B���IsH׷>���6"O��q�j�$1jʩ�CHD�
I����"O�a��R�M���_-�]S�"O����6���a��ɱI7�b�"O���f��S¥��-5*	*u"O�u�����
LR� R\��H�"O� `HS�e��{RO?�d��"O4�k)1:f<��.��eG�Yq"OѺ��%�!a,וX5�ö"OFqb����"��l�jȄ�A�"Oܴ�#��r���� A�1 ��p���B�Oڬ�ˠN�ZȨ-��d[���	�'в�a��%y�.�B����x|�!s	�'X�q���%�¸c�+�Z��)	�'Ⱦ :��ύ X�i�e�)ߓɘ'?��C��ȸm��1 �]�.5�	�'wl��c�B�|Tɳ!�Z��'
�Z�@Q�~
�q!2m"�A�
�'�z��>���Zre�.~�x��'��lIw���~T2*�E�H��'HN��E�P$o���ⶪ7qd��'��%���,o-.pk6a��( �-I�'�N(�Cc�;�(M�EjID�5�'Hb�B- �_&Fౄ�ԏ`}Y�'�>ͣ6"	�o��y#ծ��xi�'1P��@�/��ZT��3x(0�'g"���@ cB��h3
W�P`��C�'a~y:�&�xpb�@�	 E��p
�'#V`�eB	#n�"A[:6�(��	�'8 ��
^�|�*}Ȳ��&�Z�	�'-�Ej��Z�Gw�B�Z&l�Ρ+���-�re��G�
�^�yfAH��(���"Oڄ����P�T� *�qIE b"OȔ��+F+G���(�� I���g"O\$r��0_Z��f�СC�ڄ��"O��
�:U�
�$	H��U"O�m!��κ<�``25�(���"Or`��M�Xѡ0����@8S"O,a�e�&��� �΃\Grp+�"O�1�W�3� 4��t4�<�"O"��U��8����ƶj��d"Opxx4*��嘥���k�$��"OT�"B�g$���7� E�>���'����6^,�v"D0~(|�	���Y+B�	'bYhm�#�4�h����n�JC�I<<���ТD�l��S�,X�wz�C䉱`ox�i6	
�l�Ta�§�B��C�ɍs�v�"��Vk������D\�C䉒�>�j���>
��#�W-�PC�	�`%8<�&	�k$��OՋr���$7?�b 0:��튔
�#G#�(_�<�`�Kΐa����4��Ljr@�W�<1�n� H@��e��$l�F8ʖEYP�<	"O��N���f,%Q=}��)�I�<9���M�4�_"qmn�е�[Z�<��̈́�3���(�D��kZezCb	r�<���ǡ=	\�xk')T�2�I�X�<)FJ^'W��iID��8�M!��l�<Y2隺���z�אh� �-i�<�D��W�͚�!��:��pI��j�<�
�&"�x�H���e&b�<�`חS�EB@'Ze�.4`��y�<�#��_�H����]�2� .K�<y���z��s��;$ �|�v��H�<Ѡ뛟/���-�U$Q[v
�H�<�W��!����	��w�z�r�g�~�<qa�6�=���N���B�Z@�<��+U@�!Aȵ@`�}@���{�<��d�3*Jp�U�3_�j���dSO�<� +�!�T�����#q�����J�<� ����;������P�v�Ԉ"O��:���E�N�b����pDҵP�@�'�ў�O$Z *�d�;Hz�P��+�+y9&( �'޲�a7�ۢ9�4kqa��s���p�'�hQ�r�% <U3Q����� 0�'�����ݺ<B����������xb��}�ʰ҃-�*9m
U���ӛ�y�^0���K"�\��Z.�y2�J#��"$d]�&e"�B��)�yr�ίQuHx�Ҍ��$q�eJے�yrK�~ڜm/�-#���Uρ�y�C�q6���eJ�%�J��5�\���'�ў�O�،��k�QX���-�e���r�'�0�X�k(Ebq@!�D�_���'��PypA� 5Ӓe�J)7���D-�3��8�I�8C+�ʑ��|�"O�=	�5ba2�GЪ���"O��Ё�<\���Y�h��C �(�"OƐ:��4z�����5�f"O@�ڂNQ�|�b��R
n���"Or%��'���(wF�,_X���"O���Fl���� �Z��؁��'�Ā1	���@��a8�R��`%D�@�g�R(q� �#��F᫕�"D�@q�)z"���Ь(U��Ѓ!D�� g �	J4� ��͍�k�����"4D���%��# �����
=5.�iq&D�p��a�s2���t�JV�`�!H$D�hن�"v|j�P�,��8����#�"D��K��_�pe�0 �(��m��I�O���hOq��AC��Z<|Dʦ��f�� i�"O,�����S��d[& ��f�ޜ"O�P�5��(�g.�?����a"OR�q���'&fq�S\)��"O���Ľc�|��I�L�^�aD"Ovmb�&8�IkH)�Є7��ty��ӼI�]�`�\3L�Z�aN�t#��$�O����ǚ�H����F���������8�!�đ�w�����\k?��ĪT+�!�Dܢ\ܙ�R��9A9�e�D�F7z�!�K?3�u�a�o ��`��u!�9�@���Ô%
+�DWy!�מ�`Ɋ��˿N��1D�;��y�	Z�v�3�U����	ćoz�=	Ó@�°Ӈ�4"wr�u*J�cy� ��O'��(7�@}�U��)ٷ��u��,,��أM�"}�|���ȏ0רm��/Y���2�ԩ.�b�7�22�D�ȓw�V�������B�k��`P,��ȓɠ�vI��q4\��*��=�h���W̓^��m:���$?b�y�A��+}&���t_���#N�0���!�ǳ`��5�ȓwi�����.ۤm#��֭!u��"�� ��c�'<�yՆǯD���ȓw^���SɵCl��ɖ�ݿ8�¥�ȓ2{>xw���С�C�>rr|�ȓ=�qZ�˄�6��0�+P�>&u�ȓ,��9�(\	2��s!L�~��ȓJ�V(�s��'H�����8m�.!�ȓ�R1�cJ�6w~���ďX�J"��g��
��)#*y��^�r��ȓ8�,q�&�؃X�e !ʚ?,���ȓ@7�!�c�D������ "��x�ȓql`��P0?`�bՅM $KJ��S�? ��$�]��$}p0j\��d���|��)�ӏg�d�A@���d+���0��B�6�ڔ��I	%e���3�KݒB�#��쳑�Τ�� ���T��B��7n��	ɀcI�%=�!��Ən<�B�I%{��	�M�)W)�����/1�B�ɤ?��`R� ��މx�O3tFB��8L-����F�1l�� 1 �f�6B�	�k���I
V��#I�t6B�	� K>-��K�LQ�r�� ?P�^��D*?��P�8
f�A �J�)�A�u�L�<I@�G�Dm��[p�"n�!eC]H�<A�ɳu�6�*��ԡ%��Fb�K�<����nJ����}�!��%D� ���#	�V���ԈA��7��O��;�)�z5zv��Ƣ�;�i�@s��Q�'(����� 5ر(.HC�x�Y���hO?Q��d� L���r�Ė�x�p�q�+�b�<a7@��.��s�a��x�-_�<Y�$�:!6���I�=~7n���Y\�<A�o[�y�V�s�˅9mN��Z4�R[�<�/���ĀU�̀i%���r�m�'��'d�	���<6�ͰsɁ���E�Zdh<�`^
�F#ƈH�y�)0�ћ�?��R�D�O�I�jn(�$��m��!��Y��C�	6V3^�QKN�JhYc��1vH�C��<����<d�9U�E�1vB��(b�)`+��ai��tmŊq{�B�	sB���Kؿ	��鰢��JsvB�ɐRz�1z�B�2��(�1䗁9�m��J�v��&��cxh����W�h���'�  ���<�@X�.օ?E��A�'�P�ZU�����=���!9(�!��'��Y��N:j��9:j04�>��'v,��TDպx��Aq*�$z�:�'�h�	֦��m�2�rW�8"(B��yB$Y�ג1��R���)�Q.�y2�� 0)�$'�\�Bm�4ΐ���'�az�É:"zH:r��PƎ���A1�y�V�l0�4z�>}iF8��F5�y�,�ԉiQ{^t�� J��y҉F�F1�� q�Z+r�� x�ℯ�y��
8�(p�
��Z%(4��?�yrF� \��R�W�4+}�D��y	  ���QhƂ� �6-U��yR���U�0�2��Cv����u'G��y�E��_�L؂�_�_�,)��6�yR�N�up� �燄�y���H��y"%Y�+=<�!��Ͷ��`@	?�y��ͅ7x�H����N��K�e�ybMӮU�]�El�J	��TeT���=Y�y��a�(� m�>U'|�0T�ҁ�y�h��0�m�c��´j���y���;+��P@�DR������ �y2�K9������3;j��DS�yr�G�����r��8J�,���F��y�B�$���b��O�B��ag�R��yR5v��U�$\>�̴�&
	��>�O���礏(x��SfgҒ$��b�"O��b
��g�@}�R�7�"O�����
��qH!�S�K���!�DG ]M�%!R�B�z��!�>p!�d��3����7��	[��	�w�n���Ms�0��k�/N��w!J hAN���S�? ��x�T��E0����nI+�"O���E��#8��$��H߮�A�"O`ٓ��4$��y�c@2N�Bir�"O.=���p�>a��v��lѷ"O�x�Tk�1H&��6��P�˃�yR��:b�q�4hA�F�� ��$�y"��/ɴD*�"��-��UJ�&��y2��u��u�HQ
.���������=��y���Y�����-"�Hz����y��9J��zg�Z�&r6Q9Vf���y��6WRjT@g�I�4��z B���y��+`˒�
cFԢ��ə�yr㒤6 ���皚���V���y�IZ�Pά�U�Ơ&<b��/�y"���l�%�B��[pv�x�c�"��>a�O6M�vdT)�+��,Y�8iχa�<� V:��]���Of���u�<!�I9yd�I�3.\<)B=��iGk�<�*��* 5P�R�_9�XAU��e�<��"�)\� }��^�u<(�����[�<���ʏU��X��@�X2ćW�<AL�1q�^U��
�I�; �Px�(�I�<Q!FĔGQ�H�`��25��Ny��'<�	-g݄Ya&�0c�l�S0,_�jVjB�i
x�p�ыG�H�X��
ӂC��6x��R�� (M9���J;~C�I���5ǒ8|LX��O�vC�	�M;�a�b�߻A\.�K@�Kq�hC䉏J�� 
���"a���e��j����dx�0�!J��U� �j�jغ+�*�k�e�O��$!�O�Hr�� 'zUa���m�p��Y�d��I�s��@H��*ͥiM� ��4��"O*��QNɅK�F�#�^�m��-�"O� ���zh�e��m�	�"���"Op´�@.0����K&1�.@�"O�ړ��E
����@J�����P��l�O���� 7Rj�wI��+�X�X��' B�'\�r���)&����d��c��9���?	�b��ل�ȥ)&�d�5̨-�^ن�"�$�C��˞!Q��\�Rs��ȓ���v�Ǳ�@9����ȓm�h���!��`��
j��̈́��hG�C�2e�j����{7ƘA����Ob"|�e�B�5�0�S�(BE�+ٟ����W~Ҁ�wr��
B�T�F��5�����?�'��a��U�qf=�3lՂf�����'�6��S�EC(=��,��
<.��'���[�Jl������qZL��'V�������W� 
aI	�'�&�b"[,q�Xd(�#��x�L-p����O~���61:�`�_��D��E׭D��C䉻9��D��X8"��1��&b�C�ɸ9?\cW�ɬ/w�d�5�'nr�B��4��Y2�O�
6�x�ģܲDDC䉡`]d�����T'8ɓ��Z'��D t� �:�;�i�&R\��}⟟�RF%�,��ֹss�(�$J |O�c�pCb�#A"H���甫Eb4"��=D�Pڗ+�Z]I��$u��@���.D�P�d��5MJ���-�cA��UH?D��2 ��d�*�����.�m�2�*D�0���@0~�g�G�:������;D�H��K�[���b���yv�]a��%|OXb�Ĳ�a�7IЈHC'̲f�����&D�� ��F���$�\��o�)]��<{�'�R@_3m�RŋQ�T�:G�0qg蛛a)!��S�8|�"7S�:��!Nۆ!�$B�}N�$R'�Ld���'cQ-�!�d^�������[y��b��.V!�d�6?�B8QAH��`<���#ĖtM!�M�!HI�`�2�r�+�!���O0��ΐ>u�h��G�= �!��@�~�BM�"��z�h�i�d�Rv!�DN,o)6\$i�$s��(S�H��C�I80K�̎$����&�HX�B�I�`(����"wqh�����'}_C�I�=��2�+�b���sr/�15^C�	�^�쀷I�����"a�#@�B�I�Rƺ-)u��5`�e���ǮG�C��-8Y�ٓ��D�Yuf��B�/^^i@P��w����7+ǮyM�B�3Q�u����I��3b��2��C䉟#� x��@	oFm�Bj;P�C��%\Upi�u�!6'
m	�!4�
C䉜:��8�r�7��1��Y^�B�I�皴�e�7�¬x�3�B��3R�bV��I杈qI6e��B�IƸ��F�ӎDh�	�k
tB�	`.l�pc��#F�h���fY\B�	�P@�z��@=tl�vH�9op�B�	63jA�!��hM4����?g^B�	(_ �8�L� 9���U�Y�r��C�	�	av�R;��*4JR�|C�IJ� ���Q�n���y��0�BC䉵7��hC�C�"z���å�0/ \B�	'!Dv��"�ג��Q���B�I3/�,�єI�OT�]���G�C�ɛh}^�ۅ�Ǥix��:���E�FC䉯nXb��e�;H��͈��I�)QDC�!;8`����ǈ&��	R�G�HC�ɿ�r����x�:铥�P�^�
C�ɟ_�P�@��M�+�4��ďϤ7�B�ɻx8��QB�2k�"�RN�?vM\B�*Y�C���~mΜ`�HJ'�RB�I�3�Xh�@���PI�Bj�4"O��y0�ȡ���bs#�	5�*�6"O48�S��)y�ZCI�9//^��S"O�L rAe���(����x�"O�9�u�%@)�HC�gR�3��� "O>���ϝfy�h*#�#u�v!��#k�*�qv%��G���@FV2�!�D]�>Xi8�m����@�Ϛ�Q'!�� �6$ʇ]�.��9�oS�O!��=��C$����DP�R!��G@aC��J���y%�!���q�PyӔ��'Z�F�Уa7\H!�$I��$I`�ɼj����&ՈA!��Њe�Y�ŎQ�j,i%A�9vW!�$��.A3ajҸ]�|`8R�!LS!��F�	h&���m�K����rd 7;@!��L�L@
B�P�Nϸ=��c�<N;!�D�4'�H�`���\��tQa�ï]!�ƥh�J��ΈV�z0����`	!�ҷm�`�k҆�/�d0!
�|!�$�!.��0G�p]��s �(!���4��eb��T�ݰQ�\�Ko!�]-��iX�Da ��@�q`!򤕊6O�,��T�N�����[E!�� ,+�V�}�h�p��z��u;"O�1z��89Zh@#F֚Pz�"O��#'�A$�0%Ӕř�?_i�b"Oȱ��	ѧ'L��9f�V�}F�h{'"O�ti���Ps0A#��"�ȽA�"O�%re��6P���(�-��F�Xp`�"O�-+Ve��`ZhpÓ�C���X�g"O���R��V���P�����"O��g"7.`���$�bM�T"OB�%iP�f��x��@�x�B ��"O.0�!
m��E�!���X��L�"O`��!G�<7g��pH@�)<��(�"OV�# b�&[��XG4G0<�p"O
�{u�P=O��p�E�v5��1�"O�<�+H���� �%J�lx��"O�!�t刹ȴ�����<$��5�T"O���`�q��0�H� �Y2"O�h/�.<��sq�����u"O,Ա����;~0�'�U<���&"Oh����]+XWL���뙣2&�	І"OFqxf  &T���
f,[�"Ot���E�*��X2S��28��"O@�􅉣7�F���B���!6"Ox�kт�3��U1x���"O�t�D1��\��C^�@�m�#"O���A'?�B5c�Cs�Pqp"O(����vbN����P�JH�s"O4M3��!"�]Q��T� ]�"Of��2dV�w�,�bhD?&�*���"O�����9F�I�&κk��W"Ox�F&�,?�y�A�a�m��"O�pa�*�v���h���p��(96"Oh)�3�H�Ĩ\�e�N��q"O
��V�D&*|rg�hϺ� �"OdÀ�̇a0��A�ѕX��1�#"O��@�f��U~��:3IY�)��*�"O:�� l�V�3�*ڈN~�ZR"Oz��UG��dP��s$�)5��[G"ODIB4&���Pr��7'�@�҄"O�1{U(��s`\�B�H_~�*"O�	��ڏg�FL����8C�z%q�"OD5���	�&X*P��}��d��"O�8
�kO6�� �%/PG�\�b@"O�`�eC�X�nX��F�Y��q25"Op�X�@�����Uh>Z�q��"O8����h"�AI���)7�� �"O����� j�r��o��s���2s"OD��a��Z�Q�-�Tx�9�R"Ol��$�G�}B�&ꂑw�Q�6"OP�3��И ^��#�(,I��R�"O���􉝘I*�ia�ɽrߠ�ф"OQK&'�)|����$�� �x9�"OpyK ��?��ӱ�N�����"O�=I�/� ]�6�sF%��ER41"O�����X��d�Q6
	P�"O(T�à)A%ސ0�l.��U�G"O��!�$<Aw@�p��HB��"O�ݹ"$A�
�2|1
��bX�"O�4Ӓ��4-�,�j�ɘ�C[�A�"OD���T&U�TY	�N�ȀC"OT<AT舁"��'�,c�|A"O�Ht� :v"J5rC� �g�"0#�"O��p�� h3X- UD�4mʱ"O���ǂ4R�����Z�rĄ�$"O� �1��6X
B�� �E�1�&)��"O�\���w����%�m��x�"O�H��I��e���"Ov�Se��Et���䒌W�F)�P"O2��;bD�����\ )�"O�( �-D�; ����,Ap���#"OJpK!�a�J�h����`���9�"O̍k ��-A�p�G�2C�ܡQ�"Oӣ�������t�R?g��\ Q"On}!�mN�XM\��aQ�RU��b"O��3oT� ���U��PF��"O��D��T!b#�Hr8p!��,D��#�*E8<�`Q�BA�<��i��"+D���`Mv����q��f�Д�y�Η+	��qKC�ʏ<��8hS��y������g�u�JB��5<��USd��E	�0=�XU�S�1N�@�ȓ?IP���ȣ#0d���D5Ko���ȓM���� g�?=�N�C`Іo�C��#)̈́�3c�)�4�D�[?��C�#v��d��Mϩm�l�6G[?�C䉻q����,�i��3� [8K�B䉃��i�f�I�"�&D Є�8�B䉈7Cn�xt�!��
=|B�I�N,�x)��S3 -�qꐾTK�B�	(rN���L�'#��[p���\B�	�1��h"3�I�v���R@�ȬBQ�C�=��i1虫C?�Hz�FǿSb�B�	;��9��c�}����V��/��C�ɈL���͓a��A���ĂkY�B�9-n�Y�H@�M@��)���<rh�B䉦ؔ�	 �¾7fXKM�m��B��u�����'m�*`����V�C�	>b.�+���v7�Q�!�=SHRC�	�ko�	� ������[U/�(��C�I;4����ɔ�}�A�T�Vt��!�b��|�S�ODh�x��,�佱 �L�|�`qs�'��M��ٛ{h��l;�p�'t�O���d�>U<`X�'ʘq��ỀC�'~�!�DM�m93g�/UB��rE�$QF�քG<a�)	zYΔha��W:��0��h8�P�ش��'�$�"���QJ]�$F���'�n��J'�=������:K�p���锜.� �J�Mc��X�E�IFF!�"��#��l*I���x)qO8��S.ߦ���B�>Fq�2"��}2��9!
:v�j�ڵIl�I�c�f�!�Q'E�U�S�2S\����ɁJ�ў؆��funm��H�H|�J��e��C��#_��(�Ѷ��I�`u����,LO��lI�K�&��AQ�K���:r�8D�(���^�NԲ�������]���$�IR}��(Xu�ξ)Rpy�ǩ�[���1fI&D���V��C�V5�׭�����-C,!�d�7ZwRy�PI_5dy�h{Ǣ^ =�!��ط6:��vD�(]�,��AؤC[!�߄���+�.$Q᜕j�h6C䉴,<��0�X ?�DE��+4�C�I7 yt��iZ�YT�|Q��Dh�C䉜����1�L�#��UOa�C�I)h^h���M'.J�x0c��Y�VC䉾``8��5v���PB�^�:C��*6�8BT�)L�������6��C�*z�.��Z�z$�(��m�2C�)� �0��U�}�r�T���R�"O�}(���+���� �N. �Dm�G�<!7㙘O^��p�^�Sy^�:g �S�<DS	2���m�-.D̫4�u�<Q눵!���R%G�!�PXK�Q\�<٧�M�J@"�k�m� o) -�`��o�<��J���x;E�3|,�:0�[G�<� �L,-m�i+�A�&-��DBV�Y@�<�vl	�
kȈ�$ �E�h�06z�<1!�I3P��0z��q�l8Ra�<�a���O�0`q�Q	],@�d�ׄ̪�<E��'��M1��l�؈�������'Y&��3
�]p�g:2(�'��`W�X�F�^E��M��z��[�'�Z����E͸��7�%Z�8�'�����I�]>!���(�6t��D.�S��$�;; �+��jk��q�Dө�y"�ؑA�,���H8T׾�a�й�yBFN,Zkh���^M����C��yB�&o�mx�n�v�hy 1���y��S�f�ԥ�㏘�f%������0?�*O�1�CI͎CC� "�fMR=�bT"O��@���|q��Ǣ�6F�h�(R"O4��Ih>����1��S"O�;�]@"��g�Kh/�pa"O��adJ� W�E�6i�2@���a�'� ��'PjݛB`
hJ�O��t��P�'�a���1��������Z�lY��.�S���?���R�F�m�X�S���y�ĩ &DzTkюXm�ڧ���WϤ�<q���Oܨ���J�wZbY�LZ=j�h@�G��F�OgZ���>^�(���ʅE� ���O%���>8� Df�'{��nɁD��hO�)�b�I�Yj��)G�48U$�k�bB�I2_rx5(tX�h��qc�Z��*�O>�	�<��}*�J��q�J�]H�H3+ȶF�6��W"OP�G�S��q`�Ů]ά,)�'�O��}�H����.H;md9��K�|� 	���I�5����O/Riz!��
�� �`�-����s���eR7yJ���&T�d_D�k�G6D��P�l�M��QA�`Wv��D����O����剣2�		Ҩ�ǀXx%�h��O�#=�r,�U�	�Ў%;����h�ぉ`��C�ɀLٮ<��	�W�BT��C7��O��	t���O�� Pc	(�.�3 ���4��#
�'qT����]�M�n����}�I�	�'&��ʤ��,�8x��=z��@	ۓ�~�-P�>qBň�
<H�$�;���6C��ē�p>q�W=�@\�jP�
!�p��Β|�'p��>��ODH#�X5t��QC��v-�	�'�D���䗽w�ЪG�E9d��\�ߴ��'���?&?7͑,�v��eDל_��"B���D�!��֒4�P�{ă�������K�(;��O8�"~b7���]�.�ipb�����0��r�<���	 &��@��E�;O<ԃ���f̓��=�ֈ��c�d%�m���8��M�<���]k�
J�(�br��	R���ɫX�1O�-�%Cf'�Ա�&�8�l���'�qOd�1��֏e]��p`Ɖ,mk� "��<}r�S�B6p%�ҍM
}�����E b~B�I0(H �)� S%ZD��"�^��hO>���ؒR\<�sB^�\�M*g("D���$oFPWp����=��0�*T�$�%�V'5�)qO�9JN��"�"O� z<�pO	;����c�
<�8JV"O~�ڄ�J��L�Go��a�T�'O&�DU�XT$�J�l\\�2@X���MnT��'�1O�3J�TАÃ�&:`���!^�V���Z��~���F�5ע��IB�0 b!)ʼ#x�I��p?I�d�R��5���FF��\?Q�m7��'���ȉ�,�a�Ƥ)����*�B!��p>	D.?�d�R�"6YAb
��,��fW�hO?��%0;�u9cDF�!P@00���pUp�<	V"�ȟ�5C$���"6�)f@��e�ِ�"O�q:�E��|"����N��>z�,32"O��ȔK�L����r��4TgH���"O������3̹9�iɕ^|Y���2�S��e�"�#��G�G \�F�SVB�	�A~v�V� K���g�z�#=q��l�I��BϪdC ���ч�"����AjJ �❢p�{�'fe���LT?�}`ŎO͸���9�S��B�\
vU�+�0WN��ץ�ot�'�a|&�(yG��2�D�WN����Dj`(�=E��<O�� �\�s	�T��3�
ݰ�"OV�8 �<<z�$* /`���@��<I��D 7T(R �_h�%͝4"�,C�	��� I�:�Pp�M�e3듭�4��>�HD]�¬A�MtP(7�б=�]�ȓ#sz٘�뜩De6���%�8LvͥOx��Ė�N�n@�ǇG#�Pt(���(
!��f��ʱ����k2+ˉOM!�6/p�UY��8kp��qgā(Q�!��@W���GhI P�|̋�ݻ�!�$%g��XW���Zr<� ၸR�!��T��L�ǯk��C�W�>s!���O��+"��(�\ !�ZȌ�C�h+4�,���E�
�8⠄�(O�]b
/LO��!f�k���A0�	�n����Q�,D���Sc˦M�y3�\�7jʅ���+D�!"�D�X�"��O�=���Zv*D�\(TcE�XRbaOJ�O�h`W4D�xb�hC��*����G�cE� �P 6D�VG�!n���3&�����7�!�F�[�B�J@�L�*��!��Ԉu!�D��}8U[Ձ��F&8h�A�4f!�d�s���Ye��$L��H�	fY!�D��)N�����Z�J��a6�Oq!��6>�nYH�f��d��L��+�5E�!���%��U
�蔠,�x҃�� �!��ywx#2+0����WdM�T�!� V0V=I�
��jrQ��1AG!�$A��|��&Z�oЀ���M��*!�=Sv�9��D#�25��OF.eI!�D��;���-�(��aQ,O	p�!�d�ܞX��E
	���kԬD�!�\�|󴐃�\?$�H � þ8/!�DҼP�M��I�s�(�&�3M!����U�� k�	�7T!��X�6a��)�8�B��"(^!�DWL�R�"�_8�ԭ!M�''R!���"z}���D �_�E{s�4~Q!�d���j �5�(}H��Z�O9!�P䌀�6э &����C䉢Cp>ecP����C��/�LC�	B#�̢�ITz��p8�jIDC�	�!�D|17��*8�0;�J�>q�jC�9jb�<PS�ėA��|�d��*�C�)� T�Bt��4�8@�p)(c7xT�"O��kh���gR=O>	�A"O����F_�Sf:�S���<R���k"OD���+[7|I�M�� ��b�2MZ�"O�UXsǓ�L܄,X�.�N��@"O���r�EfXq�.��	�&=�G�� ?�8���,*HD	�G� �1O>Q0EO�@9f�ЀLȃC���A"O���ѝij����%�"OdH�jR�Q�P���#L	��r"O��@�A�HZ9�)�#7ƾ��"O�aH�T�&�JEP1i��R"OTh[��T� Q�� M �t��"OH,r�`GL�d-���;�Z�6"OnA���
�����s�P�x���"O�Ir�J�e�Rq�ꅻgJD�a"O�A:�%ۑY�̱�V*�"�,Xs"O����e]�?�F��w��A���"Or���bԾd�jQԆMri��"O����P��mhD@T�3�:��"O�l���� ��5QS�ئ|�`}��"O�q������[4@:2�t��"O�QU�W'xxQ�/X�:�P�"O<  ��:�F�#4b<\��C"O�u���Ƴe4��2��)r�p�P"O*u��>=H�U��N�X�9 B"OD��S�B2f\�T�q��!e"O`�ćЖ�q���tŤ%�0"O��P�L�*� �H1�%�l"O�*D�Yh)򈰤/�:a�\���"O
�᤭T\)��h��A,F��|�R"O�t��	عg��a &*Y�1nv�cT"O�X���L�2��`F<�"OHX��0����šA�=�Q��"Oꈘ'�QC[Nab�I�h��"O��I@�MБ�C7n��ؗ���7�t⟒��Q���I/}�T���(F�]�	b"O����\���8"�V�N�hG��ʸ'�Z����Ԛ!� �<) �Os���3C&D��b�l�8|L$ոv�@�P�t|�j��%�Ф���'4�aqi��"N��ǟ�b���`	ӓ�f���O*}�#�H0�����
Z^�Ӱ�Z��y⧟�6lXY�ae��_��20��ɘ'���j�iNP�S�'8�����%���`�j{7�ȓbͪm�Ԋ(-j�0ǁ-e��\��:�	�Dj "|�'?�Xڂ��?d�F��� 9NH����'���D�O�,�&p2��Z�:8r�gj�H�����4ݲE�#��f�Yw猙o��|R�2d���J��)�P��� "���2uxC�	�q������9!��s�̹`f�#<)G,��m�8�~� 咻��X�2fR�$�1P���}�<9�gG�V t�3�]1A<ָbb �:ryb�;ua �)��<����,,��(+�xlJKB{�<A���RҶ�js-ݫ7@��s��<	U�(3�������5�040'@
%T�q���F�a|�h[p�<��;'(�����gXV�b&���}%(	��_���#$k�=7 0a���?��Fx� �Q�ZuG�į*y.>Y7n[9b��zG�4�y��6`�<�0vF�3��2�"�w��a#��3�)��Lef��+��T�2-��O{���Q!&D���S3_��u\-&i�	;�0D�X�3��^� �+���h$����/D��y� �5�4�*ħD�l����+-D���TH�)44P(ư<���B�+D���@(��{��bRE�0.>
-�"�(D�� ��"�jyLTh0b��e�&1��"On����J&>�ǢA$w�Hu��"O�Aw�I>.N��s��<�H���"O.�����p�`x�IO��"��s"O����V;�ޠy%/�	G�z�CE"O��R1m��bVk��(���U�LJyah/�'4KJ�	�D_�"kz�Z�!*�	�ȓ3�x����ڀX��js�N�Tp�t�*G()Ȫ�'�������A�;q���$�LߞTy'l/4�<�A�'8���E�_�~U�T7��!k��C�ȼ\��q��	�2�d�9&�o��h2�J�]�����l��@b��K�^���I�:2���o �+��)@FD+�C�	6N�h�@N�;[T~��`-���Oz�4�+�I�4�6�4	��([�-ϧu����N �R���q�E�ȓ¢�(�)",���$
;7C����[�L�蔖'�����A0iC"��ܭ!"-oީ����)|05 Ѯ��5D�ГJ,4��I�kњ?>�XKd�ǺZK��#�G�
��c�M6@Sp���y��1���h���#=�1sSZY�5$�#8h�!�(	�/����d� 0|�qph�,���	.v|�ȳ�\3�F +���<pC��r�G>~��3�3C��ȇ�I�Z����D� 1F51�-�6*�D�OD=��P�)�J����i� R��yb��X�d��$^~cȀ��БREФ� ,Vh<��
C�[�ʍ3$d���x�hR��++�:����|�:�W%�0��"
��X�#4T?1�au�U��CCs�qY���F��� G2D����'c ��a�o�����	� �8�F\�F/	-���0H��&a$����ɮQEX�)Ģ�F�����68�B�	W��q)tB�_�L��e��k�"-��A/Fy���E[��9��j�b8�(@� _���+F�T�(�bɒa�=,OhY	LP+[����ѹ�N�`I^�~�j�{#��=W([c��
��C��^�|@��H�,��Q�3و�x7�Uj|���?(qH K�\�>�D��v'W�2Z�>����"P����_(S�)	4�>\O�5�'犕���`��÷�m݊	ke)S�a��
=z�\�-X�V���j���5}"��%x���NT�3(bjcO��'���G�y�O�0��JËLAq3�
�>��ځd?�$� �`��1���.N*I�xr �=]Ơ�P �phA��	�&�B�B�[v�4&p`B��?kt>����x	�9C�"�:T�� J�YQYV,Z��Pxbgͯoj�����V�^�rUMj	��W�0��ul�]�J�mK�+}���&?�h��}b�j��0P8�	BD�/�pe���R������^����M�D�U��s��[/��*����X��lw���D�&�A�m2�3}rD�D�d�#�-P@����&���'�|�#0O���ό6��h�J�E��O�Δ{�i��r� )v��-\^����M�C�� j��<a�σ0@G�DK�AƤkb��!"�v}2eZ�7,Mc�>	T�
5Vl\�F&ڞ!�|pK�OC�IՐ�)R��*w�x�ѳm=\�4���'{j��-�
P0���g4Zz`�� 
�� ��mz�@+�凁%�d����P6��֧ε]vp�>� �y�����.�	S�_/M1���f�'<M�C��_�hHQ�2�DT��/oo��r�l��"�b��7�O)A�Ҷ�/Ȁh"l�t�R��|
�yAKo 0�Q2(J�i�n�����?�6�C$���f
��yiBE�c�˄m) �!��
�����.���bNk����	�"���dC�o+�`�&�[:J�d�#��$ҭpC��,O����̘0�D� �/�$�V��
�ؤI�������O�3j��4m�5�Z��P+�-�6<��>�$-C�	�z�ƸC�W_ �pF�� ����)Y�M��u"#��m6�z��&]�`hF�v� ȡ��E���䈔8�˓k:�B`�� W����-�`����  � �h�\��#��'P���!x,�#B��Լ��r��.r�P�`TG��W�X������U�V��Dw���^�����85���2+��g�p����g$�1�ih�fFl�_60ܰ�c�'8�.=	�(W cØ���CL�$�ՠZ�4Dj��Y�(Q�f��$U����#�rl��I�)��<hY���"�>�N4iU����*�o�2>%*H�+DT�hx�L�7�R�S�?�D �?�0Ė�-�	�3!*]����m�]�xC�᫋�I�}��
D���)�lq��
�) 3J����J�3A�<d9�͐)���>f��e�.�`��\��&��[u��|3��d�����ߝN�����&�6)�>U��p�(t1P���� A�*۲	�­A�
�W��U���l]X�g�G{<��R;����Æ�
$`�O����&�'g�aX��3�'F~2�� �
����#V?:�[� V<9E`)9��0�O$@��]�&�dI���PV�)2A�R�6-�mbJ>9aԟ6!��C	Ϧ���O� ���H�T��Y��1l��A��"O:��E쌂���h������|���'�� �q��\�k!��I;铞�π  �ӥ*�;q��� �B9�"O�	W�G� ��j%X ~�(�D�sG��- �`(�3��.phi ���Nt"���%��	�qO��᲎O��r�k�gߋr�D����B�j�;��#y����
�0?�c��+[���J�H�!�P�pH��?C���M>P��s�tmV�G�Q��>���^+6��`�K���H3��Sh<a�EH464RJ�5WFIA����`Z�\[3� #��QS%%J��>M��B��h����(:����%<Ol��E-2���O ѐ��V�`�p�jg�I&"\TXb"O�t�FK�>8�J�窉�uB(���|�
I�pN0�g)�W�O�v�Xf��J��[@����'c�����R�a^���J*	���J��[�H.�'�U��>A���Q�$-8�/ѫ"�~L��A�Uh<��"�l��`D䙼O��{jQ2S+���X�DC��o�t-F%Zv:O���(H3��'��J���%�t&��1���*����f��2��7�^���jȫSb�� �zJlA����k��6m7bN�"ao)LO�-�膘m�9���E:"��Q�|��A�F=,����~�j��&!Z=+DP����5ç�P0NZĢ��&�>Y����/%C�",�0��K�;x����@MZ<�"N�! Ρp����h	FP8�1t����)Ǡ$(�Ξ6��dQ�C��X���si�.!��ڃt���*�$�%c�+WU�u�1HG/�EF�u
��w�HG���u���:��O��O�8�߄ !�8�Ss�A��MI���XУ�*az� �+��k���DB�|'L8���F����F��6D*��ϓ_�<���5���A���+πE���9C̸r�U
A�c�d�>"�n��o#rI��*/3�4Yt�&4��pcj٢�h����*���a�<���ج&����2��,5#Ȩ"v�����P���Vi��$h�� �>��q"O�zL�+*�L����:V*�M��n��v���BJE=�SՂ��!8$�� ǂ�5gL"1@�<O�.�I҈/�O*�i�(O�r(��[�)���]�`+_�C�>P�%�?�5�q�Z���mztk�ux��S%�3H�KB���??@���&�E0��*q&٥P�-1B�i>T��H8V'ĸx��#F��eoR�:�����Kh<Q�C�N٪�兣9ʄ� �'T���bIڗE��@t���B�㇖Lݮ �~��UL�e�g�ʹ5;�Թ���?pb���o3 �J����R�	�C��	r��tY��`elݚ0�4`�P�������=�%��_��Q�+�T.,s� �vX�`Fn�k�|]�*�%:�J9ᠣ،p�.L�t�P,c��B��#F�*�@��%P�Ġ�N���"=��"I�jl�%�]R�CvP� C  I��A13��D��ȇȓ&ݬ��6NѪz~&!I��Қw�p�	)j���Gg��v]�S�O�D�%⁛*��tå�<�r��@"OT(���	!�����ڧ|�Ṉ�\�ԓ�7h��+!�'�\A�фءn�~���_#z8y�=�4�Z��B�8W(	r����ۼ���@��P��'UH8�a�_���1����ҡ���3d�MÉ�	Ջ/�j5
�-��a�*Ы�ӧ�ybϑ�$N>U�R�Z&]��#��yr�_3?G�MR��U�9�w⏲�y2Oc�|�rQCL���Q��䔍�y�A�1p:�B��~n	#%���y�EH�O��lU Q�2�!"�[�J�!�䚐	�p���	�G�*�g��$M!�!���Cah��z���˅D9BP!�9>��bEM٥ܦ<{a�T6!�d��F��Ȓ'��2];"�G+]%!�@h`�����}n�Is��~!�ď�1ܸ�[�%Q+sg��
�	}�!��
�YVj�;�E�������F��!�dѴl	hĸ����
�X`M���!�D�,h�쵋��I#c���r�"@�,�!�$Y����GD��[������K�!��I$�1��Z�"�p)bᏚY�!�fN�hۆdE�|.���'|�!��	�`�E�4b���PÍ�!�� F�&�0T�"��Ch�5yJ���"OvB�*�z.X'͟d
HA"O��%,
�M� �I�t4
�"O���h�	�����f �c$"O~�05��c<* ��eL	AF>���"O�� ��
b3�m�SE�:< A�"O�]�Z�?�*���#	(�x�"O�)��w������QuE��"O��	e���P����>d��K�"O6d�F���6�'X~�x6"O�u�t�٥����S
�>/�$�7"O(\�
G ���a3HX�d&*O�$�WSјiʀǁ�b��I�'����"���P�b��ŸQ/�,�ʓs���O�L�l���JZ<(���ȓ7:��F'ײaWaӠ�?K[X�ȓ��qE��&G�nk�+�3+��؇ȓ^��\��)RD�L��/�h(��Yߨ���P�ǐ:,4��ŝs�<��'�r̘��vn��j��'��F�<�5�!9�Ă��-k�
�:c!AB�<	Q�/-���bO��@�v�Fg�<тM=G��Q��Xxt5:Ջ�c�<")�2��`EVd�l� �X�<�B��
t������pP'�[Y�<A���3)�����,���Ń��XZ�<�sN�c2Ԓ�Lˇ�"��$�Z[�<!A�Oi
 PhL
8X�	�Bh_{�<)��(=�U`�.G�N�,+�mZ|�<��a�	&��*��]4�L��	�x�<���Z9_˜�S'��`������1D�ʐ��K:�=r�#׏5b��b�/D��XC��vq��L��+)px��i,D������e�b�Ԭ_�^������*D��.�5j2�l��E9r-PA�di+D�0&��lO��X���4m#� 'D������%b'r��Q��'�$D�@���_^9f̠B ��5���1i?D�(P�Ñ/�B�s�'Ť7v�80��;D�H��c����J2� �ڊ���':D�(ӕoU�>�ȁ�7�A�b]:����9D���҇��c{��H����<j���5D��!M?[`����	9D-�x�4D�8Y���6��j���1F<rD��"7D��r#7l�dQ�δU�.TY��2D�<hu�؍ͅF L��@�aC> ��C�	>U�ySanD�jЕ��-��C�ɐLT�!�N�~3�89��A �fC����(
Fa�)+���㰯H]�B�I��h���0O�D�e�ӷVچB�I�C�� � �ϡ0�^���j[�k�lB䉡GjXԹ�IF� ��A��Z'C�IH:� Ag��&�������r�$B�I�?���(Q�d<~U(b�W�f3�C�	�3�Эb�(�"�<I���R61�8C�&�hp�v͉�.ض�&+��@��B�I�
���J�T�jI��$��B�I'���C3AƈO������"�jB�	�cO�ݫ�
��ƨ�7��.S$LB�ɢb^bg��e��"��(CRB�Ip���ߴL���a���}#$B�	-?:�A���,���S�Z3�C�I�n�z��A#PA�8�����b��B�ɾ7k64��K\3T��0�����B�)� X�ug�/�؉3��9`�5`@"O <Z��#l1J��ơ�5L�̣�"O0��ц�/(�j!;#��8��"Ob���ɮy�Á)�#�T��"O�|��+�7i8�(A�ʰ0͔	��"O~�{�LV$`��0@�
���2"O�A��X�d,}{W�� �,��"O��x���s�:$բy�*��"Ol��6/�>
�� @+�2*��A�"Ox�6��6��A�ɗ�v�ѓ��ڻ{����+7�'1�ָ!�ϥ-�,��F�=Z��Q�ȓf����,�`�T���o�\�B�\�Z�P�'�֩��@12�P��H!�I� �m���/4�����8vBܵ;f���L��S�.Ģ�[W$�� dB���I�L�T#!H�� ���˄*�����#���Q���(��ɇօC�f����"F��H*��d�+D���t)]�}T�C��`w"}���'��>c}:M�r�H��#~��j�h0q�u���:XƱ��c�<Y�M5H|Υ���yA��O
V�!r�L6M{ĭ�'�45E��>)p�Ɋچ���ȟB���I[h<Ia���l���{��O�2��Q�A%sT��
��1��@;���+CK��v0=[�B�c�����	�p '��g���̓J?�0Xe�ók�n��3��9�m�ȓ93��vH�WZ��B��a�z$$�슧�L;b�t8�ccNo�O2}�
V~E�J�)�%k�`��'�|-Z2BΎ'X�-�i��%��x�99G'}�,����	tOr����5^�@<8G� LD�C�(ž��U���(Lx0�Q(����r��^��T		�Eג!��c
�"���#��8q��ȓq�VhX��
�[U�����W�1D��sdB2;����t'�3tJ���,D��YTK�`u��~��9X��,D� c���80�T��A������,D���F�	2��%�m�Y��;�'?D��c��ɽ@CD%H��&X�|=Z�G&D��I���4(yx��#��,ׂT�$D�샃�_�?R$id���]q�Q�wf'D�h���S�'Xq K�S����e(D��1'"}�0��ڀL���� J5D����V��^�:B��z��yR��2D�`Ct虚H��IVG���A�g/D�<`�e� CH��z/hc<M��.�s�<!q�46"�cb-ֻ/��R���h�'�lИ$��u�	s�J�f
�*�>IG�(9��䲣��Ph!�DXO~~X3Q�F��T��T�}��ɉ$�T��\��50@d	.�	��Q\$X��^�n��OO3{����� ��1�Y�0���:�@���O �ќ�IpoK�/�q-�<y��A<.
�`@�.�>��ȉd[�5#Æ��q`��NGeX�=0i��8'&�i�|L���I�u��֋�&T���c��tv:G�iyBdH��	dh�q�'�])r� $\�����1�a�H��xgA��9n��F��(B����E
t�Sƺ$12dR7?���(�U ��-���%O2i���'(���jJ�f��K��]%!� ] AR�y��R�N��Q2�HQ��ڇ�ʠ`���s��]$��$�r�ݓã�h\X$�%k��C�9C�d�`�Ύ|c��ӧJ�dw�� �`��4���>v�y��R	��9K���Ҥ؞��		VX#��O�AC���(/������<w1�b�Ҡ6�8В�B�t|�+$ V5U��X�gVg6�ȃG���$�Z�9�����O���ɫ?ݪy4��`�~��>1���>u�X�j���=|(,A�G{a�H�|��/	㶍 A��6����D'��UJ��0B�[�f���� -8�R*[#&��ʤ�F	-^�y��)Q��!JM -N�z�q2�:�rU�;���2w�P���
IbD���0@C�	�:~�f,�	\*:}�d��?m�
�o����e�R�O�@���(�0`���f�����!���_zԼ0a���[P�E�_�ayr���N�c�Q�����ɹJT|���8�#ؐ�pm����$(�� ���g:�3�D?̼91�k�GZ҉Eg�"(��'[ց��+�h��哿�� D�3p�B�A9|���΂˚��7>�8�1��'�B���HNФx�0`�dZ����3�� %�`J�OE�l��-�0UЊ	�'��ȪUϒ%eG��U������
�'y�if���`աY+>@x��aH(1�HL�R���@�Ć��	X�'	9�D��%7	`M"&d�56L%��@�#�l�z5s=rM�p��`�$�
�n�ʌ�L>Q I�*A��a�&L���F�qO$�C�A�����&�H`
C�	z��Ag�I�GVN0�W��?9�>������0?��@@P�u�� O�9P���cE�y�I>1p#�E��/1B�hR�>!A���K}� �LV*Š��kh<Yflχa�������{��L��kO�I��d &�țzSX��7�L�����>��B��4˔T�R���"W��y�'/<O�D����'_��i�O�EAe��6/xL��pH�8�P�ȡ"O�XX5�¡L�<�*��<M�����|2=H��<���	E�OQ��j�*�9c��p�K2�xJ
�'��K��� �j�#��G2�E��� ?W���'f�%� ��>��`˗@(�!�Pf]&+�@u�B�MIh<邀C�]w�0��G�T�`�q��P�O�EX�g�2l�����;���I�$I��!�I$z;T�yg� ::��/Ƥ��$�9.�J'�ƥ�M�d��8��z����P7�S�#�fP�s�(�Mc A���}b�0t&8��[a��(�+�+�`'��8���#,�tSg�3j���(��ьs�`(�Bȷ3r,0�Ķl52vB�)�L��Z�alLU��V�9��MP�e��0�D0�*$H�I��M���#�Ƞ�S���,"��l��Sj�![( �T���$�Dx�L5j�C�	�4c��a�N�4i
��e)8��P3��R�p�F��l[���S�4a��q�n��$����>/o�����	tl��Q��;�O�	�`*�; �r5�t�A�b��ٰ���L�X�c"�M�x{FȟN�R����p���6.�����Ѥ�,f�f�?iw�[��6d���F��1����u( �E�����aټ���Q1Oh���gߣ"`De� A��/<�:%[��1�)`Ȯ,��ԭYi|ݹWHH��Oj���bC���+�|����'�R<8AC�u8���҄ob���$EA 48G^	r`&U�V�ى���>�ĒOD���M*B�(�w �]-x����'=��ys��?д��m��3e�ϡ�����M�P.���fʍ3V��J��'���yf%Æf;��!π	��1���& m�E��Y�x$t6��t܄�4�M�A�𱢪I��L��'�*��'n`h�"���ʰ�+ܰ ���'-��K�����	/6: aQ͜@��&P@�&m��oa
���LU�}�t��'s4����Y������̾n |U1�'Qn��e�K9����V��>�S,Z^��p��b��;͎@{�@�}hY8�E!�OlM Z}S��`��ǫx�p� χ~1JQ���Πy�~B≄'��H��C8ye���у/, �=�wɪA-J��@>�ӥPS��1�X�M�ʘt��!<v�C䉽y��e���N}��B�������Y7[��|�P��-��)�'f^$k�I�z�T�*b(ފ��9{�'H�����~`|�;A�^�	����*O����y{,X{˓]����m� �Z "/��1mh-����7���J�%G@I�y@��
���2QH��Q�@�ƓrŨ,��@�3�����B�c-dXG}B�J�
МE��М~It+C�϶D���� �y�L��)������22��-����yR���g���Tm_+�P�9�㑛�y��W�o��ai�^�+��\��
H�yҎ�]�R-[���R�6��T���y����0U�L/u��4�0�;L� ��ȓu��4��jE"0�&�d�C4Y�`��	P��!҃�3}x-���46����%dxM��H�C��aAI�K��ԅ�-�x�j ,�DZ }(�(�j��`���	��M�!A&���C�=�Ȇȓ<������;u�2Ȼ�eS�K|�|��z�X � ��{�!�tGF0OFB��ȓOU
�S�ϛ' &Pr�)��d2I�ȓ�4!ab��)`�}b�b�g����S�? B�"�$"�Ƶ�	��]O���"Of��!Z I��4�'��) ��;�"O�uS��`�@�� �4��e"Oi�u=w�ƴ�6��"s�~���"O�T�@�#A�z}�a�8
}@%q "O����AȂ��i�F�͈���#C"O��C�j � S"}c��O�H�F"OJ<���Q��:�׉�lQY�"O�	��ѡ�ԉ0aB��^�\]�@"O��aVD%�"��oQ�R�LX��"O�}ؑ�P�e����&p�L�:"O.���@U8#q��0˂A��i�"O�p��e�&Pg0��VKMo���D"O��� �ԃ\���Sk��Q7��$�Z>V8��h�BZMV���ٲ:�1O���� Uy<�ꆥM�H�@�"Oz #PݗbD�Se��}���e"O:}�g���J!���IJf:|��"O� �ӸaȮiДƟ0�|`�"O�@�T�]�\���҃"ϒ(B"O��d�����Y�a�!�t���"O��UC	3T�p&@Q�B��t�W"O>�b�(s�	����i)�"O>�sb��z_�YP6�X��� ��"O�@q�+�+#%4��S�K=$>�!�1[��،����,��#-։\�ޅ �'"���C���>�`㞢Zb��En�P�׺P���P%z��O.�#e!�!�0|R�[A�\��@B:)  �eCX_���tSB"���0�0|b��	G��`!N�w�b�U��]}2HF�q�^�K�0��56��dk�L� 	�j/�����6&ʖx�� ��S�`XA��ǺZ� e�\�o,~�lZ�(A��P�9�!(��
K�h��動�u�8��x���b�۫'PB  ����B���ȓYn���EA�	s?C�E��r�<�Tɂ�{�h����xz�e	�I�<�^r�=��I�y�x̃�EJ�<q!.b ���G�<D�r�<�g��A�b�SOC?�Hd��Kd�'�ў�W_���O^��YTL��_M΅�ȓr
� ��E����+���.vΠ�ȓ;�Hh�q�Ԓ7�������2O|݇�4�0i��_<	ڔ�T�A�<߰Ňȓ{V1HT��'Ҥa��.p<�M��w�S"��^���XħE(�⁇ȓl�jmX a�+Nf���
L�䠆�bk5��#S�B_
Q��eU����#>���uAC3FA@TI
 
��ȓGf��H�� ��˄�Ȁ2�(��v�xJpaMHD��_�>���"�@a)w�923������Ʉȓa�:���$D�ū�t�q��'u�#bʆ,"~�L��iv���ȓ��qɤ@2.ɤ̱�x��0D�\�Q��+�D��Q���a$#,D����m�98����5	��yDxiA*D�����T�(5��I�Hƌ2o'D���$Uh��3�ǒ@���D#D��*芩2�$@V�E�]�\,��� D�<K�i�6�ā�LB IT68���=D��� )M%1X$�p(2��y::D��H��ˁ=L���6�OA��Z֏9D��cga%�f-��M��E���k�7D�v�ɁhY�KÆW����T�7D��*��*f��U(��
�]4� �5D��`�ѲV�.�˦FM�+�xp�A�4D�� ����$Qaڄ D] �8(�"O<��cJOC�bЪ ���"O��r3�,B~����L]/���c�"O�͇�+������$>��`"O��ڂ��74@�@@�a�/3���ɐ"O:9�2(]�Y�X�Ra�+�V�Q1"O<ؓ�isuจ@�=i�� "O^ݱ�J8~5��
�/2UxBb"O�DP�J�A��؛G%MVY�B�"OJؑ"KE\�4�bbH(�qV"O&���D1*7b�vF2JU`qrE"O�];p��98���`���"Kf �"O�s��.D�<X*�dӨ#�d}*7"O`��U  \T=q��b;2�;�"O����I~8�!��A �q"OF����-��0���*e��*"O�"��H�D�f왦b�p��"�"O8$��,V�y�&�{ �F�6z؈��"OxY�Be�����T�l�p�"O�`�'*��J�P(.�
aK�s""O ��a*޿ �D��A�%7&�`R"O���ǖ%�� Ѳ�߾e�M�g"O,�����	ypz��ʙ�����q"Oܸ���0>�\��q��,Zހ���"O�Xp�J��e�E�ӹF�2�q�"OT�0��ȔB����a&�MJb"OZD����f����Se��I�"O�%!��>������ѽDk��"Ox��c�L
:������7X�2 "OL�;H��#i�=d˼_����F"Ov��&��I&
����ٽC�d�pE"O�uS��J�p�^h�u��	v5fhrc"O�(����źs&;�(M�"O�qaq%[>9�ĝ�JݒM0^�{�"OT��:CuR@㵈A-@&�œ "O�����>�H0AY~tq "O���d��U �?k�`��f�Z�<!P�߀8}&��!S�ZSX��m�<	�l��x�z���-%xɩ�+Nf�<�׍�9)���Շ) �����f�<I�L	�E8콂E�)��i�\�<A�M�;'$�����e�$�A�C�< �!s)v�`�Q�E�I��Gy�<ׂ� \.Ԙ�c�&[l�k3��m�<A���|�x�Zb�E�  ݀�$q�<qa�ִn���@UÍ|OT�D��l�<�!��A`p4P$��$n,��m�g�<5(Č*r�%�1�Ȟ���s�/Im�<I�
�%t������0s� �l�<y���Oyp�	VkF<4܊��Qf�<��_��8	q�m���p`H`�<���E�*� �'[Qr�B���X�<�:H��H`u&�q�Јԭ�U�<�Ҩ��s]ĩ����j�qB��f�<�IӦqW�e��nĝE֜B� �Z�<�o�]"��d�$8T�qT�AW�<�Ư��;���2�I8<y�M1��h�<N�� a �0\t�]�Q�Lf�<��I��)+:���B�*��XBňU[�<�t��|���6kS)~]�iҵ"RN�<Q'��H��@��CA�b�dOe�<姓�W�^���Ř!`�`-�g��f�<�`�H2H�a��s��;�o�Z�<I�#�5UTA�n̛&��`�]m�<� ��;�	N�D���&h�8��A�f"Ox���*_U�����*��P "O��Ya�ͣM!
a�#M��8���c!"O�$W ��w����E��+Bf��Hd"O���	ч�:D{w�>e�\L
�"O֠:$� �)@ą�1 :s$��"O|�`���Y��A�!k�X�@"O�)����_������)3bD�R"O���éRCH̻��ǐMU�5��"O6�c�e�0���MۿN a�"O��6!�3UH��$�U[\�)!"O�HVg�1i�nAYP+n'V���'�e(c�,*e.]���ҡ��ai�'�.ս(�(+G��4r|X(��'lr��e�j��Z%��rOup	�'hܠa��Eف��-c(���'�u�V�η,x�U�`��`��X�	�'r�����&�`ģa!_�>(��'j����	�lmRa%��U��i�'� `RLQ��Ƀ� �$�i�'�pH  �
*@m�B�(CCFa��'M���PX�5�M����/Fg���'N8 RM��@5�Q��F�l��'C��D	�9��Za&\h1~Y��'��!�A vI��b�ML<k�t�c�'�����Cr$h��#�`�
)�'N�E�7�s%�ط�� [���	�'��9��D�>\����rMښMn䌓�'}4�	tL�V��T8� X�L���'�걣܊6_���q�\7 4�z	�'��y��,�j@ �c 'R�K����'�<S�T'$�h�Eˬ��D��'B����2}���k��<W<D�<�Vk�"���ݔ2O��3�>D���T���t���G��a�/D�P�1e̕tmxT�R��b���.�$C�	4wR���k��r�ΥC\q�B��' �Q��FM�@�"�8��juXh
�'.���M:Ag��FJY.3��
�'��9��\�7?�h��G$]�fa��'��hPVB] ���R���!�u�':�1�UIN���k�bޱe"���'�Z��TH!�b�3A@�h�&���'^��!B��>y������R�JX�'�4y�T.Z8XP�I��*�!L�Bx��'7D��B	ߦr��I$l[�X��`�'�J)��P�q�r`�� *�̭�'gH���:e�~9��`þ<���
�'����%��J
!PqG�^:ً	�'� 	�d}��ؑ��V#Y��� 	�'"���R)9��hA ���R�:%@�'�&�Q�9z��(�j�x���'T H7�^!B��|�@��w��\��'\��B@eA�;�:��FHV���'��dQr���,��3i�3k�N`��'���ɣB�h, ��r���d��L��'�z�S����E	R���aİ��'c�)&�%R�h����,,R�'�h�
��q�p���H��"^@��')^ �TMD6�l��t-W�f� ��'���p	C.
��ݐ��L�`��'�)V#
��,b��%�xi{�'x,��W�&��Qh�#� ��'o��j�"FS
�HH�C�6������ >��E��0XL�\�f���El��F"O���Bf���˄��2�Q�"O<���ۃ%�� W�C�����"O�a���˘Y��T���Upz���"O�	�fč�2B�8���\=ojJ0+�"O�D�wCD�1�UH���~�� "OL�A@*��]��"EdÀKfı�C"O��a�̖�0A؍bw��&a���"O�A����nC��wʗ�V���:�'�hI �T$|Ա���&J�-R�'�ڹ� �v\<;�cL8R\�L3�'�q����z|B�]-E'*��'���"��U޺�X0J�jt��'������R[� =�/� 0B渺
�'Ӷ��p�߂��ТD|�����'��@* �#�Ս{�tp��'ۖC�7�"d�r��q:ܙ�'N���7gX�Y���`�#B��<X
�'S�͘U&[O��c��f{�)�	�'�8ͲG���gR�e{Р�.M���I�'H.u��gB�sֲuba �*���
�'���'EB��bh�3��(�	x�'/*%����hE��Y0��z0�D��'���B��/����锳=�����'�X�jVfI
��#���	T��	�'��]�Ղ��w��B㪆%q ��H	�'"�i!���0"Mk"� > \�ر�'
J���\�{��B�J� *A�#�'\�HN��_w�y�1�_�V(��
�'%4Mh��j׬my����4��	�'�(}q㯅��1r��>b�I��'��d�a��9j��*Qo��.��I��'�X:5ƅ���xEˈxijTS�'�xy۰BC$4\|Y0b՝t�t�Q�'��S�(�Q�E�r% ��'pk�ID�d#�Q� ��&enݛ�'�@�����	I��ই+����'��1��c��2�M�P({ƘQ	�'�rr�P�Х��+W��Q�*Î�y�-����*�e��ld�hڠ���y �*m]� I�7m��R�떘�yRNC^�r� #g�d ��Ƙ�yBf����ÅǢDے@�Hܹ�y2fK(3 @  �