MPQ    Am    h�  h                                                                                 ȥC=�3T��)7K�|����<��괟��A������κ��X.C���TD����))��0!��W�b�����X�����f��[˙!-@�MNh'� {�ڵ����=4�EnyK��2�f��Ժ��,���U��x���S13-�@=�����Y���C ���.��&U��L�B=#GQ8w m_�����,$�q{TMU��͒�	�*E�}.t��Q4�9ꞯ.&kz{���Έ�S����4g4�Z�9�aX�I���Y�5�Rb��ˁ�W2p��ZbS36�#�6�S
���)B��ZԺ��c}w������K��/��	��3_Z��].��W4����+����e!�V�V�!����EO�@���<Fj�D��(����K�7j���*���[�P��+/5-	��]�H#N$����ҲU� ����2D7}��@��eX(�9\�y�ucba�vȏ�B��-p�	m��N�����#a���?����'��%�ᚍ�ٛ�_�Й����4��ǹ��W��)����"s�h�� �o�,6MT[�łkg��H�)75�}?ӥ8 ����]�iyp{�{l6�ۚ�������+�j�[�=��/�b�J�B��/.��x��o7�\P.��x��Z��%M���M�?$����9Q�"�o}C|F�L��ӄ�5�/LH�3�D�ӄ�\Z��Q���}�� �~�G�:8`lip�m����%�4@�F�c���G^�M�u�*�,�j�A�ϐrU���s��i�"<�2l [��܉�&�i�>racj�b�V��<�s�A��߳߇��/�y!��8���V-9w��C�V�IM�N��Y�\B��~��T-�u�K�����咶��֑����,c��A��79r[,-.�&��A��I��o��$Q��0�7�!`QdXOD�I�g�%R�� >��VA
�3[�#-m�[vlZ���!�Z�+�ѝ�;�`�&C�V�3�٦�W�b�1�U�Y��G0�c)��V�?�8T/�'�"���"��5�Ɵ����..�ݒ���F3,�C�l�1��A��+j�����Q��r�x�?޲9̚+�J�e�g��Kjjhc��Oى_&���%]�o�qU�wf�N����k%�����y?�im���zu|�1�w�����2O��D�T���r���QwV?���
����lg�<�q���ug5��ӭ���O%����Dާ�ڍj��U&��J�EfL�X�}T�G1ÏP?�!���+O�W���@NJՀyE���؀��CֱinD�D����Z�������'�@AzXg>��ue�.6�ȶ��}�v���0�k[,���ҥyV��q�^��8�f\�"� yQA ~��˧G����"��阯�i�7�3{�]U;��Q�R�[�i��=b�H[C��S����fTUD�s���Q���I��1k��>:������)E�Hǃ����oa������rpښ�_���t��5��Vב��*�ZfV����3���k1�p�(�4��r�XK�1Y)�	!�deC���p��ҏ
cQe��
�_Wv�9(�9�0KHV�7} ����%��p�
nr?>K�$�yU�Q��C���Bg�բ$�� �#�>�%�J�i��cV��+����R�d^�w��%/m���V�m H��m��q�W��/XYH�{������p7�}bã��8��n��T��y���Y��Mؽ���M��l��5O0�_�!��y	H|�A����簲uEg������_F���V=�LYߝ����~�*����UB�he��d/]�����3��Q��@�ȞA��Z��^���'�U�Xi��.@�T�N���O�VS��i��p�S7=6M����Y�uYw�!?��+[-�V:@99Z<~������;)ׁQ���;�Ev���2��a����u�?��qw��X�,F��(����<�0�em��X<�b��!�nYM	ak�z��-���ԝ�yO�>�#a�%YY{>�N���
��69	��$գ�d�Xq����j_���Co�;�͡^�E����B��:�ٵv�-h%��RC�9{U��U�������3�([x�(9��1i�SI��&[ʃ��8�@]`�۰�g�%�I}�$���X���Gx�ڥκ�N�Q��q,:N��v���7:شS"9��&	K��6�Ě6�3�k�W	�"t+\r���o��XӇ��?�!R��}��0QE�>��}��7��xg�h:��b��&ݿ5�H������+@r���e֠�.x�	-u���c�� Kw�(�>��6#P�ϒ9_a��2���.p���~Ā���U$���S�%o�#Y�\�R�l���/�ǅ�f�e�P�x�u�t�S��U�D��h�ȱ�ۙ�r��r�jo�ߙ#��70Ԡ�۳���%duF��>8v��H"-������G�L{�^��Nz��̢���ۓC�=�aePأ�L�A����ߙ@�Z��m���-�B��B�etq$�`4Ǎ��� ��<��������N��}�+��M�rh�����]���{uC,����0J(�Pe$�����qݗ�i0�ɋ�>�^�&~�#:I�c���b�G�����f���L{������M�Uoew���Jz�j���5��SX���p�U� �;�הk{�I��6Ap�Hc2a�6f��I��!O�B���&w	:Y�'��$/�h�6�W�z��9G-3�h�R8�"�K7^5���+CѤcMSyųh���ԫ��C�kb!/�9���;u���"ʢ�s��/ӗ���OӤW1�����RX@z�Y/��x�H#��5��Ql����6�g4�b�6b�;�Ý���7B�J�Qg>l��}��n�9��zb���>\�o���'��-	�c�l��ڰ�&�e�_��\������G���OC�0�6�.Ou͸��c�Z��j����?Ѡ���_hu� ��W+�zl�����G����~c���tk����1ߌ3U=�P����iW?��Ui�c���oӳ3��NpgM�%�`��\����r�2�e8�����m"�y<RݽN���wy�`��5��Lԏ:�z����e���4���/�Mw�K
6��v�m�Z��>]wô^�%��8�
�4W�l���2ȿy'(����n���*V�Y���ӯ�J��Z�$��+�5����T�[�be~���`Z��P�U�_EϨCcQnB�"���/���;�{�5Y_Q��ys;�&F�K���1~���?C�<��i���[$x�p�gΘ��4^K=r~��s��2��n�-���;l�zs���`���b�G���9S@�W1�}�)�\K��h_ V�_/	"$���S&_6-+A�
�+�/Pè?��Н�sn�$��I0
)�Fg���γ�<�K(٭��w���G��,5+�ʿ	��B���#)$F�4�߲���͢U#��78C�x���(���"�Nu�/��q��ics�ٴ�,G�F��)�#��Յڹ������	�\+ᵛ �ln������=��>���aWR�B��=lӄ�� q���WSIM�i��}�g����䃯��#��~�`��:��)��]#�wpvPIla�j�Uן��m$��|��6����l�b*/Ǒ=�/�p_�SۇɊ��\�+p�S�lǕ��%��ϝ��	?N��N'4�=4�}�ě�'�ӿf�5t�?H�ADH�Q��j���N�>pe��#�~�:Ӆ�iI���m8�ߠ�4��۰>�K�۰���w�u�΍P�j�[�����U�sj)l�]�+�g Vj]7����!i���a��4�dfJV�;l���A�3+�Y����y<U�b̈1�Ow)k0��{�M�S��y�B:�~�H-V�-K�6g�g��-���a��-�c���A��9�`�[D.�Ɯ�<�,�u��]Ղo��Q�݌䲚�`,�O����%����[c���MV\���F�#��[�"ɽ�$g�U� �,�/;�����6��3�����������|�}��!�G�z)�J��s8/��'���v�0���
���EO�.![���C�buF3g{O�������3��o�����^���ueF���m�Ƽ�`^�g��%�n��Ɣ�;x:�v�B�6]<���l}�w��t�׷���r�u����֏%	�m��߀u�|B���X��l+��G��鵶Hr��A�L5f?z���f3���K�l�Ԡ�L��װ&�5e����O����q�������[۫0����cE�X6TY�J���<$
�u���_#�!edJp,�y@���ִϰ���oEDi��g�̯&BG�2����'Gj�z����a�e]����o��#��F�0� �,xZ��D��yq��qE΢��BvfG�"Q�~Q<�A�_S��$�� *����[��ҷ���;]P����zR�������=��p[#������.aj��ٻsFQ��(I:tk�)u>ub��9��)@d�ޗ�\�5a�Dm�Y��p�P>_*p�!%5������*o��fqUe�3�D�kl2ͳ+���%��0�KPS�)�h1!���C[�.�@��*y�L��e<W�"�9C&�̑�H��7���X����˧�)�->f���g,�CR���T���zj���#b�@����Z�>c������#tL�_�w��I/(Q��!#��g\ #��N2�m�'&�{v%���M��0�cq�Ō���#p@��}�H��qŌC�j�{��ٔsI��?��(�s�.�ł$]s�{
�O�����ϥ|�4�eQ���TEo��i�_�Sr��Б�g
Ý,`	�Y��5��U��h`'�d�6Zӝ����ѩ�'F�̈́�|y�Z-�Y��Zx'*Z����I��Ti�а	H��H.c��k,�7�eۊ�!�tu�u�,���r��3,d-g^c@44�<��!�ǡB�V� �̪k��Zvһ�2>Y4aˉ���n������U,��ިF��?}�ˢ�m�U���[b`����J�M���k��ã9Oz(�=0�0U���a�.&Y�`&{'lN0�
W�9�/X����q��K!���^��o�r��<}zE{~��:B6�v�!�%<_�CZ�~{G����+��^�4,[3ϗ98a1���S$�w&�F�w- ;��68�g��2I�Z�܈��X���G�H��-�>s���T,*�N˒�����@�S]�}��Ӫ��T���3u�����	���+71��aߺ����~A���?K!mj����0,:yq_}6L���,���m��/�&�5�������a+{�5��qn�ӭ�d�>� ��9���1R���y���љ���s_�!y���I�G�pN�?��F<"U�p��N�o�ב�ݡ�,�ԭ�Nˢ��=e{��x�Ut�2���I��$�C�t�!��",j
���O�7��4�	�.��d��w��m�-P3ܥ���G	����:�ir��k�ޣu�A��	�=d�P��YLZ���j�&�[o��s�����'�}��BK^Kqz0�b��H�c��S<xR���ĺ��`��+�}��8�r#����;G]K�{P����U��(��q$�q��̶zq�;[i����U^�]3I���@���B�.I�C�'=����݉�MUj�F�n��J5�����53�S3j�B���Me2 �T�o9�k6pzI�"RA���cyd6�����:�!J�@�'U�w�S�Yx�쟂�h���W�97�2�-._�ϭ�+"O^PX#�@+?�c�|"�N����7��,C���!J��3~v;P�?��=����^!���O�~�1��?��@U�3/�劍�Iq��ԧ���p�6�c&����];�LR�W��2���5".������y�S*���I���z�9�o'`Z�	RȜ瞧����e�
��ͷ�C]rҚ���Q�_,�wuh��^K�LP��b�ѻb������:꾒�z�ѩ���G�;�9��3�t�a�n�Ǵ*=]�
��~�W������B�~���"����q���M�9�`�rQ\��v�-�8����:+/�H>��H+Rx<��I��	���p�P��LOg*�Utn��"&�썍̼/�	ЂR���gm2}C��<��%�5�8��4�o���n��M�'y��`����n�`*�WnY�^�!�s�+�u0$H��m���s���_ey9�`SZH���p��EJ��c,�y�]`���vq�{Yv�Y"��Q��s�$F�$�r�1y6�8ӂ���i����֛�x�9�g	}'��ɠ=m]��ζ�2��n��j֒;GOwsӑ���w��]�K�7��S���1�)+)���K�������p�	�7�Wh�_��{A�oԦ�&P�r�?/ϐ��`4i���E��
�tF�:���Oj��KQ8|�4�|������+���	�@�
�2#D�o�@���Q��xj~=C7�F���~��(q��]�Hu���l*��#$�=�}p)��{<딟U#��C�u;�jr��ζW�u��ɵّ]����N�M5��$Y�|O^W����)�X�ք^9| L��0M����x�gK������'å�&�Ǳ;�dD�]�|�pq�l����ϐ��\4�!O��߽�3�Nb�3�8��/���^fɥ˫\FI��.�:��Cr%�iD���?��	5[�X��}9-������ٶ5�H�oYD��~��k5�l��#9��F�~!$�:n�0i�A/#-��(+��;�46�|�n�:��(�u��/q��j{
�};U�&�sE���D-h�O Q��F���!�i� �aYs��?�iV�oabAȍ��i�J��yWn.Bw��VwdՌm�M�x��>�B�k~�J�-ѪK��Ѓ>!��O���Q]��cn��A�At9�6[�A�.���׌��0Ƿ��6ot@OQ����-[�`�GO�m)����%�=5Ƕ�Vw� Vw�)R#�BI[����1¤�P̇^K;H8�����3�������w�����G��5))yf�5�
8
�V'������+z�ek7� ��.<$-݈���=�3�r/��r����Z���*���q�h4�@m?�(�a=�[��gn������m�E���A�}�[]�Pd�g�(w�ʒ��	`h��iYӠS`!Um�r�p%�|�������*�*�(`���g�>9r2�ܡGR?�'�!|��Fl]8��'g��T�5 ������O�Xt�,}���E[�`
��T�%�E��[X��T�{����WZ�����H�\�.J��y;?D���k�����D}���B��a��1i�����'��=z�0ɶ�m�e�-��~�H��}�%�0��p,�Ά���Ey���q��s��lbf��"��Q7@���R����,�����e�Շ�Bl�iJ~]K��p�9Rx�G��o2=Xle[�����[k���P\�5���s��Q�B`I���k[T{>����!);e��9�n�a������np�&C_e���ٶ5�h��G)�**[f���]�3|�Fk��Y�NO�B��(�K�e)�!x}C6ء�����G	���ݖWy�9^����*H��}7�d��煯&t�� >�a�o����C�nr���9��rL�_��#��[�_ط�,�#����C��ZīwO��/㾧G�L0 �\��emDb��v��?�ڥ)�~�i��~㙦�{�}��b��ʕ��?F�6<�ٯn��O�����i�т�m��v.oO��U�鯵+|�tw�@*]�&{�E��`��X�_�!��oj���T��4�#�p��UI�\h[��d�/��X5��^�Ggj���0���%Z�͉��U'�~��ΨE�dntT�C�Ћ㶿�]x���f| 7󴉊A\�Ə8uO���g�nL�-�D@/O�<4X뫂g;�q2�Gˬ��߿v�2��a�o'�+��P�!	�,<6
�� H�zE1�f��m���Lb�����M�Z�k�f�t���J~��P���j�a�lOYObw{�W�Nk_]
�o 9�v����ږ�q����+�9z�o0�s�׻vEv����J:��rv�5�%���C5y�{��}݋ն��f��/[��
9S`�1_�S��G&ф�B�6�����gl+�I�D���X���G��P��
�S�~C�G�N�g��vmz��QS�ŵ\���ڒ�P�30D �u�	w�+d�>狀;���yJ!�PE�?I�!���s�0�B�
�}���� ��������&�&�>W���+����5�>��L眿	�zJ��TE�Id-(gִ6!�l0?��F
_������d(;��=uz���|UZr��I�o=����<��G���L��}y��5e
Ox�Ut62��ˁr��fL����O� �2��j�|'��7�	�Qd�Indk���׵�W�U-�u����DGd�O���ք�����Pm�	�H=���P�E�L�"�%��vȓ���z$�����B�v:qu\n�����p�6t<�G�w��5]���m}��]�ږr�5G��%]ƶ�{+;ͳ?����(ڴ�$<s(���q "i&\�����^F+�/��I٥ �����ځ+ݳ�����$�`Ue����MjJ���1�5�\�S��}����! �:)�ʻGk�=$I��5Af�$c�=6������!E����w��Y(���Qh�܇W	xh��$-)`���"
�J^kw��m�+�̫c��_��)��	p��a�qCc)�!e8��r;+)=zW���i������q�OIxG1--�ĺۊ@0v�/�Dq�~�#��ϧO�H�+w:6��啁u�_�;�՝�D�-죬 ��=������v���EE�9��4�koh�h'��	:D՜b�RӃ��e7����2��7Q�U4M-�꽕0,���;g%�u~�YG��U��^���*3�U����u���7�z�T
���9Gg����v�N��tx��}�;�V�=�����Z�W�Zઇ���6Е������ĨMm`�V\Vn��A��*������#z閃��R۝�DF>n����a�kH�L�^��0[I��Y����	�/T�(����im��p��`�*٘%=�-8���4w��zab�h<8y#z��28nA�*�7|Y�1��|x������e�$� ���T��&�+�5et��q�Z�(��6E���ct!��N��e�M���d{
�Y=��Q�Yns�6�F��1tL�ϓ�b����i���QU�x�"�gD��jU.=h\3�)�2MC n�����;"�Cs��Ֆn��XJ�䒸S��g1��)�Kd���ڕ��	.S���B_���A��[�!��Py\�?j�d�K-�d0m���
��F����y�EFK�hS��%:���S�a!�+`V�	��e��Y#߃����&A���n[��R7���/Iڬ�w�(L����u4+�g��U����2��<Bs�o5e#=F�����M�8�*d��s�o�a��Έ�l�����w��W!���s�!�ٕ. 't����M%���s%�g��Z}P��KW�t�%âHi����]Y6�pl
Yl{q��慹�ḵ�A��� ��nG/b`X�3m�/?�V�� i���\��0�	�8��-%�p��v�?5��b��sމ}�������5m(5���Hؽ|D����$d��ar�4�����~\:	1�i�ZR~e'��nN���4��)��[]�Q����3u�v���j6٩� #�U��Es ;������� L����W{�i⑭a�'���XVR�G�2A�X�ī�~ryr�;�A���Mw����'+Mǽ��j"B�x�~ձ�-L��KkJJ�y���c���a���c)��A�9|k[��.Pg(�rt,���*+o/��Q�7��;`��7O�X�8#�%��J�!2�V�"
�}3#��,['�����K������;ԩ n,Zh3hK�V�k�3��r�!�jx�Gaߔ)Dw���h�8塒'S�˅Q}��&�\��Qf�.W���u���3݉�=qΨסq�����"� n��㋴���c@���o��Vxg�.V�aV�@���`����"�]r%��b-bww�!�M='$
�kW��{���Ym�8��kXZ|����ΰ�Ev����{��Xh�y|Hr�.O�B?0�������5,�lػ-�Z��&�L5��j����O6A��pb������؂��g�`��E7n�X>qT"���ly�r�0�k�������J��Ey6a��3]�&>���wD�G�t �� ̿��'��z���ՙteS��Y3�.����k0��,.cj��ћy���q;�Гc�^f��
"�&SQ2 ���ƧxN׉G�: �h�@���T��x]F|��˰8R3�#��\�=��%[�Bo����P�JW�oU�es�wQ��Iѽk6��>���o�C)6��ǔ�t�dNaܪ��O�pk�_����E�`5�T�ע�U*�1�f��z[ϱ3Wfuk�\��g�
�.܃=K���)){Z!�9�C$�!�^�`�+B����W4ܐ9y&̇�H��P7.7Q���4u��`��y>������[�5cC�K��p�Ɗʴ�#��Xvm���u'�܏�^�`�Y3h�U�Sw�=R/�L��פ�� �TX��Gm߼��q�"�h���`B���ł�7�tI����}3����Cb��ס�����ʉ������a�Ƥ�q�Z���qr6OAl�N��ʻ�|>��#��a�.E8'���g	_W��*$���b�"i��9X󫴙U��IhV�]d@I�zz�'hS������J͞�KZc������'��)߉x��5�T_� �f�5�����2�a��7N$X���1ƪ�_u��;���D˩�-���@*�l<����=Mx��������/uvH2�2t��a�u����޷d��<��,��!��Q���Y��m��(M��b֒B���Mz1�k]㣯�~^��H��kF�o��a�ʠYʃ�{Ϩ�N�˨
�c�9����5H�����qg�P�v�okA�r�Eq�h�S��:�O'v�i%2��C �{�{X�&������DM3[���9nK1���S�M(&�v�1Uԯ��g'�7I�N��~1,Xw��G)���L,D�bpr���N]=����oS��`������� ī.63���U�	�lQ+���y���oo�tsB���?���!�����D0�����<}l�^���v�y4��̊&.��չ�0��+�^����F�����5�+�o�+��|���c������_r� c|m����fMBU�����U����Dl�o���L�bqۭ��.�X#��ke��bx�u�t�Q�ㆌ����:�9B��*5�m��j@t_�37AS��db�d�_���Mϒ��-��2��B�G�LJ���h֟�}�a�+��D�Y=�jP��4L�Ļ�-B����i�~�Uz̆��0B��Aqp�\b{Ǿ�!�Q��<n� �R�2�pylS�}�j��%r�����K]Aӑ{�U�z!M��j(Ֆ�$����B0�q.�Pi�ç���^�]+�0�I�R9��X�x�ҁF���=Q�� pVEYݿ�U`m��$�`J�rN�1�5)ZvS�Jˋ�o��� �}��%^k�+I�L�A�@Ec�g6*���!@�п��mw:%bYCx 앉hpߌWD��hJR-$���c�"���^���L�+�zc�.1ń����Լ�VC�!�g�)��;�j�ˏ�se���r��^?O�e1H~��5P�@zW/:�+��-�3'��]���H6�B�A��;LAM��o�(�&�[9��mh�4���x�3Q�"�Z�T��H��/l�oÝ�'֯�	UV���)����8��e�9����\�1p�zKH߱����������u��؈T���{��� ���������־�z=�:��"zG�$H����i��t��+�X���=�=��^��VnWPֲ�B����.��������t�M���`���\�jˣ�����Q�0���������R���?��ɋlב^8��ܽLEvN�b�K��\�č�f�/�⁂|A��)��m("*����e�4%�>G8�"4h��5tX����y��?�a��n|��*'7BY�$n��j��{�����$���\H�a�8�,v�eo�k�WZ��*��U}E@c�&9��\�� ��'�{ϽZYX#<Q��s̔�FB7��B�1o����Y�m�gi�����.�x�+kg����=c{�߄��2�n+ї`�v;���sI�-�1�a�S4g���DSq(�15�)���K?~�OZ�0T�	����_gl)A��ԜO�PTf�?�9M��~_�{��gk
Zp�F��R��~� ��KǸ^�j}���3t����+L	{� 8M#��m��c����ᾄ(4��7i(VJᔬt('���R�u�XM�b�2�zⳜ�MVͷ(��J�#M�܅�#��E��������Xه���<]�����Z�ʹrWcw:s�����T- ����{M�Uv�ng{gb�*w��S��}����H�]�Dpg�lr'�ۆ����T��ǂ~���#b����.Ep/���Ï���\<���f�Ft%��U��E?��a��uΎ�"}/^d���y�p �5E�+H�+|DY���H����Q`��꤫Z�~��:���i�qٽ-����0ғ4,!��i>�������u�z�'z0j���;�Uw's���L�` Gw8H�>���i�B�aO����1V�y�U�YA��x�����!y���$a�¨4w�ɮ�°M�"���&@Bk~�8R-�_~KFԃ����h��g�>�Pc�SA
Q9� �[��.�g��|@�5�n�_o�k�Q�Q�#<Y`��wO0dY�ӕ%�<�l�K�	�V�j��=#���[bνg]�F��=�;��;37��W3C������W��mZ���S�G&�)_��+J�8��~'�:��0�!��XU�vd�.ry�~���H(3�k�؏]�ғ�D1n�b�;b��^��0ޞ�����Q5�g$�VI��S�;#�˭��o�]��]�7w����~?�K��d��V��ֱmQ���f��|S;�뉮��`+����������rh���=/�?����m �ṖlS_V��l�a,56�7��ioO�I֢��t�<��V�h��]�o�E�YX�OTjUE�{ա�& ��Q?�s:��ґ�JA��y1�������*>��2}Ds������׏8g6ԅ�\�'X��zDz���jeά��4�˻i��[��0��v,�N�u�y��Aq����> kf�0�""s!Q-�4�p�Z�3�b�C�`���Y�U�q埙+]A'��&�wR�(D��i�=N��[���?���Rl��KswX�Q��I���k
�>&U��
p)1�X��X��Рa��4��U�pF2�_ۃ���"5�`���x*�(Qf�_m�`�32'Tkg̈́�������K�x�)D4[!n�C��\������=-ߟv�NW��X9�����Hy�7i)w�)����lnZ>�_*�e_[��PCI��%m����>t#�	����U3C�I#a��B��P��w�6/Y�D9�]�B!� �l�mz7��l�k��9U�{�����@��O��*}Ι���*�T�}������2�E�������ϥ���V�l�O�O�˜����|�'���;���)E������_�o���'�����߻��\���6U�hQ�Gd��5���ʱBd��=F�ˬ�Y�-�eZ� ��I�';'��Dh���^Tڸ��A�ĿB�H4��\|7��F��1��ŋ/uE��aQ���-85/@%��<�>��R���]��=l����zv���2qa�����~�����W9),2m%��6ʗ�����Am�Ȼ���b��U�ڣM�'<k8�J��r��{GA���*��aIYEŝ{��N�W�
(w�9�d�א�4�P�q���(��;o�ؒ��wEl��M�:s�v���%���C���{�'��������	7[dF�9��/1U�aS��&G��H˴,=3�G�$g��I�x����dXR��Gd�ȥ�m �H����]��Nr��l���7/S�P������n�l�3��%Vn	mps+�)[��k��q:�o�_���?|:!����iL�0��*��}�F��_��ǹ�N��&IX��4j��h\?+,Ce�kT����F�uf�=m銧�������*�x������zK_�}D���`Z��|{0<����U��q�?��o�<�H\��}��!��3�R�eLCx���t��A�0�Kѹ�5��O���jۋO�&7��q�������daȅ��5����-![���(G⤚J.ֺӅ�z����=5X<P�g�Lk� ������^��Gt�0�v�.�)BaqkgsM��yUw�l��<��&�-��������}�G�I�trT���&�]��{Ხ��h�&+&(И�$��ʓ��
qI��iK�cZ�^���e��I���Q��3�΁a�!y*��Bc����Z�NU[]�\wJf�7�L�-5�w�S�ċ�i��T( ���� �kg9DI�UA\�1c���6R���jp!;�b�8�Ew��7Y^(��=�hKWT'���-�GϾپ"�o^��I�J`+�H�c9���k���ש���C�f@!������;��G�_������t�'͓O��G1c�İ��@条/uc���}��ڧ�����96�m� ���";�븝(P�#&����S���O�����,a�敏x�o���*\�o��'���	p��X����XsgSemJݾ��TL���ߍc�@���Eۜn�ݛ�u9Ö�O3D�]�������C�K���~Ku�C��z�oc��s�G��j�ᄋt��3Ʌ�x�#=.�,��r�W�q%������ҵ��5U�����:arMR48`��\ۃ�^E�ќ������Q����RIxف:��$}(�L{r���;L�����Ϸ����*�~��/
�ڂ7��D3m��o����à��%s��8�j�4��p��r��0Qy���<_n��*�V�Y�7��2�@�6ݖ��/�$�1G���$��!��� hejs�q�jZy#�����E�v(c����������m�x{��oYsn�Q���s��F}pWC�<1j��IM�(P�i� ��G(�xdT�g��
Š��=^�e�߱�2��AnF�w�C[;�jMs�5�̻R�N>�H+^S,�1P�)��K��K������	���he__"l�A(���*VP/�?��I��&ZP&�Vj
�FӀv��+��)K)�������P��[+�a�	5H�{�#�c� �\�\��Ṻ����7$�$e�7����(����uj�t�]�C��$7�n��h� �2/�%�4#�?�F�h��mY��P~�w-�!f��b��:���k��عm��W��.�6񩐐�Ϯw ݫd�C0�M[�N�i�eg\����������j}��X֔��i]�	#pbDYl��x�Av|�ꔱ��lӢw��,b���)=�/����?�����\�a�ؿ��ǁ<A%Tx�}�{?�q�:iΩ�}�&ꛓ��ӫ�5��HιWD�F���b6�*�<�5oV~�^�:?\i��46��YVu�K͙4�������Ǖ��T�u�����j��#�VϕU��4s��V�I�j9�< Bf��Q(�͎i�a��/�е�V�xs��A�[��z~*�{��y�B��� ���w�k�]pM���� KyB&�w~�e-B�K!�m���c�%]������<�c���A%�;9r��[sp�.Ƈ�ꨣ�!�����o�1�Q��\e`�Ok��n(k%�
��8��ZrV�Ҵ�44#tsD[�;�[.�A��̘o�;ykQ:�"�S37B�#^�i��h�6� O�G׌?)zӪ��K�8��'�_\��r���v~�1Vi.�?���9���$i3Sȕs�D�ͥ����[���Vv�ٚ�ѡ����y�2���LGg�QN��������.�C]�.I�X]�w-�N��B�Z�9�a�V�1��*>m�}�a�|���D�v�{ ���iT�H[��b�r伡8m>?濕�R��k�l�"k踟�ל�5�>���r�O�qG�]�
�.�X���Z��;?��aEm��X��JTŨ��6�ԡ����a�)�N�؎6�J��y,�UϜt���D�:��ӻ��?1����v'�O�z�NȶR�eI�؃�u��Lj��-0�4�,��1�0qTy�Blq1�.���f3�Q"�߇Q(�h�ː���}-��o���c��S��:q�]<�����R�����=�}[���z������Myo�s2Y�Q+xI	�k�.>a;���ʔ),(�J�H\wa���E�Cp!h�_u�{��5����X�:*[?if�M�Qw3�kXc~�z�� �(�9�8K<7)_�!�`C����4Җs�8сzW�9�v!�}U%HT(�7�;���[B�-ȯ7�G�>� ������NC>fd���j����p��#NL����������Դ���rd�K��w`"[/��Tv���I ��:?
m���gn��������q�x�n�*��,.�}i�F���h��g���  ���y��]��n��_(�gZO�R���� (�|1H��tE���En�����w_M����#��i���1�!S�Uc,hLύd��>Ӊc��]�u���_ˇH֞hbtZ�����.�'��F��wV��#�TU�X�1d�}]�ϸD�W,7cU�r����}�u�B|�hF��m�-Ӽ8@ `%<E�ȫ�x���:���8��/�v�(�2�ca����<�~�����r@,�8�oq��+��7Yem��J�bL���V�Mp>�k�B�%��D��߭�a��^fa/�Y�&s{��QN\
ê�9�.��4y�,�q7Y�������o��ͨ7|Eg�=�	�g:.�<v2�%(}�C���{3���\�����f���:[�|9��1�+ZS�Q&����?!'E.����g���I���t,IX-�eG���!�e��]���a|N7�������SIi��->�����a��3a��!v8	蓁+��-��Y�����j%y�a~'?7�Q!������0�:�e�j}�G��<c�/{D�	�&dN�կ#L�CEZ+gGݍ�����М�D���r饈Y�������ec�=����D�_(�H�œ��,��\� {1�2�EU+7��:vMoN�u������?����e�Rx�itG������2��/�G��>���#|jv���
;�7�G	њ\�d��w��7n�1-����dGu�_��'�Ւ�W���l�ۺb�=�e^P�( L�c��V�m��;��_v����iP�B���qf���X��4�p���<d�X�k���U�\}��6��r�ܮ`o]7l@{��׳���y9(˺=$M7쓸)Xqd�i���>��^�! ��I���QJ���΁|�$�����f����)UV�����J!�E�g��5��S��.����? �c��5k"g�I	��A�1�cy�6�0��Pe�!6ѿ��}w�vqYy��.h&E�W�򴵞��-���";^�^�H�i�+�6octa�ź;�����r^C�5!���do;���+]ʩ����Z���[�Oz%�1~�,�+��@��/�"�O$K��`���\�6��� �}�D;µ����[����-%�jzT�n!�[��d��
"��%loy�T'L�"	����4]d���G>e�ݹc���n҆e~9��r��w^��bu�-�J٤��%7�� �'C�����Y惾~��zs-�����Gx%U�%.4៞3t�{|�߳�I=������W-8������d���z���um�M��`~��\g�]������&��ô�ۖ4�.R�v��5\O�������d!L;#���z��й��}�y�j/e;4�򰐾_�mGA������ �%�B8��p4M��������Yy��ϛ�:n��d*]��Y�j���o�����$�i̠|�P��dO�b��eeq��I�Z4�[��5�E6�/c�츛I��6���}0�`7{E�Y�٢Q�d8s���F��i�#�1e��Ϥ`��HiW���A<x?��g�M�;�'=YY�:��2~ �na3�V��;�^�s���g��Ih�䣔WS�1/1k�)v��K����#w�f�R		������_݋�AC�RԒ$~P
�9?$Z�S(Um��ƈ
ХvF�B�}�w���K=�������)�r�+���	P5w�8�#p�[z�����W���7߉W�q¬j��(��I�u��X�P�0e��)���ͭU`� ��#��Ņ����Y��I��CN�<�}cN��~��9f���P�hk�W���`n��)��Jk ����~�M���dK�g�c����p�x�����3͒�P�&]*#zp]��l(�����}�1Yű٪�}��Ib1�p�$Uf/P�����I�t�\2��ؚSǼ$�%�gG�x�n?FZ�������M�}%<�n�G���u5{o�H�gD��I�.��1��a~]X:�![i�e��κ��N�f�4"�y��尟����*�u�����EjgצqծUm�ns��ɫ��<�1Q =uL�?ҋ�H�i3raE탫YV�����A�5��՗�6�+y�# \�x&�wP���sFM�LO�{��B��~&�-��K���*1M�4m��Q����#cZ3~A@J�9���[N�.Ȁ�C��\��$��o`�Q(���=`sc�O��٭	۞%䕴�"��c˵V�Zf�#Onx[ؑ���xL�<����_�;4g�U���}[3��D���I]�cr�{j�G��)�1g�!m"8v4g'�2�"��V���s��g�.����t�{�� z3����-����ޤ��|��q���TR��H��gߚ�l��Ggڣa�x�
>Y�1V�1�ij�]Ccp�S%�w�{�~��u�ϵ�߭���Lm����\��|	 j��	�ɖ���s�f�L�*�r�3˚?A�}��sنlilIl�����MG5l�����KOG�8�%�I���LY�w9�¤E��X��aT ���x��r��$@�)l��H�`Jwfwy'>I����Wފ�U`Di�?��7�M���I��P�'�z�C��&ޏeīp�����&D��B0��m,?����y��q�R0��S�fn�"Xl�Q# 9�&�⧩s���N����� ���CG��h�]7� ��/�Rd4Q��n=Dn0[e�Ǔ����!KIH�Gf�5s�y�Q5cPI�#�k�?�>�Ar�@��)'��ǥy��a-����B�p���_Q�Խ��5��׳��*v%f�[���3�"k��ͺ����ܔ�rK�ۯ)z5!d/C�Ǐ��]�1�3Ѣ�,��Web�9�Z�����H/j7�m��_���+��� Р>��]�[��s�\Cy�2�[� ������#	�]�;��K�������*���F�w�Ŀ/ϵ�oä8�� j�du��m����b|��y�:ڑLf�'��G����g�}ł�{n��
a��"�F����;X�ot�U�ʂ+��b�4ORv^A�g���|�Z;��͝��<E	�W��T�_h�-�[���_o��f@�����\��U��!hG	0dQU(�D�x���3�4�b�B���vZ4�K��3�'�O�ߺ����JhTЭF������ij�1�R��7_2��-������u;���CK��Z�-nd�@�<����n�ǉ�7I�3���]�uv��2Ev�a�G����޷<v����>,($�J��f^���րm�
�^bF�*M�t�k�ʣ`�\/-q��k�}ރ�E�aJ��Y;�t{`[�NW��
^�49�ҹ�F�}�ƝsqRa�UV��)og�C��Eb2�d��:��v-�Q%��oC���{n ���2��C_�U�>[�5 9���1K��Sk*&�y?�~�%"mů���gX��I-����X;Gڤx�����.�s���UNR��b��\'MS�l,�Ȩ3���}ļF.3'�<��	c�{+~op�*hS�����e����&�?�W�!��_I'0s����}=O_������No��(.&d��*��N%+�k	��������+Cof�<���\�(�7�֠3!���>��.�_��,������;2��p�mqUƸ�5+0o�=�¾�k�����u�����W�e��-x���t�o�l�M�����ۻ�^�tjX��@7R���=�sѵ	`dWI6�`���C��-W�	��$|G�lz�����*6�ґࣼw|���E=k�xP�	`L!dX��I������;|����BR�qaL�)�c��b��lT<�	���h��!�a��}���sSr����5�m]��	{��г+W \�(��$���s։qPNi�R��#^2�m�]I�l��x��Ӂ�ٯo��n�y��ݐ	�UQ�x�5�J�Zw���Y5�zSzF�i�B�T� ���6�kݴtI$��AR�ncT��6����f!1����wkOY��r��h�<W����9{-< �tj�"���^�#��\+eD{c�*�U,]��������CO$�!�Y��;�Lf�Q�D���).��	}O5�X1�1�Ħm�@�E�/�T���]�U�������640��?%X�V;��l�^Kz����l�ɼ���K�����Z����~� �;o��8'��	�L��N�?W��G]e���ݴ^�
�M�A������r��RnS�/uo���E����J��B���AM��4����+z���u#G��������gt�7��t��=d$��
pWa�s!��;��؞�U�밙�M�{=`y��\������թ����dÏ�w�o�AR�u�0Nڿ@�����XoL�|/Ȝ6���-��t=�/�������zѿm�	��`�	�N�%��$8�Z�4yԳ�fl�Ԥ
y	����eFn--�*���YĽh��!
������y$v��W4͏�X��u�e`��''�Z������E��#cs� ��G{���]�f�8i�{ �%Y�dbQyS�s]n�F�By�1`\����"��m�i)��={�xlg0����Õ=T��ߕN29*�n|��,;�r�s����=�D����1S��91�f )�GK�Z������b	��|_��LA^�_�?2P�Cq?V�~����P�O���
�p�F	����Np��Kxi��;D`���=�͊�+L��	kBq��#K�f��5���ᯆ�ES7�j��i5�奷(����E�u����S/Z�����'���(�����D#���|����eՔ�Gy�D��W�����e��?��tB;�+���cB�Wt:(��i�����G� �c��"M�a�_�NgE��F�C�:��`��������]�\IpX�Il��۷���L�}��Ku�Xh��Z|zb�*����/�������,��\����uu��,%%�wT�s�?��O��Y�߲�}�Z�I�&�!�75�H�5�Dj�yG�I⚉ �1����~H{+:u�i����A�Ͻ���#�4��W�`SB�=�q��{4u�F�8�@j"T.����U�u�s��쫿	�o� 8�0YN<�C"�iN�a�9���7V>��&��A�/�0���P�y���#�S��w�H�Փ�M�p����B�w?~A�%-8_�K��уe�J�������O;�c�IA[	9hg[)��.<(���R���\�S}obQCl���`N�O�E����%߻:�}�\]V� �k�#*�[�8�b�7���NpV;�	p��to3Ԣ�B���^.��֥�GM�z)��K����8Q�c'?X������m�,+���.����2k��<[3�&������)f�U�"�8X�����)C�"�O	9�hVQ�B,ag5`��V%}���*�\�)��C]޷/�Naw�b��9�]���WM���d�z3m"w�Wd�|d��g�ɱ
����]�A���e�:r9��.I�?������١l�l�	Y�neq��5Jp���O�"�����d�*��Rc�RWW�L�|E���X�͔T{�%ì����H_�W���5T��ޯJҢy"�m��hױ&>D�����������8Z���M'i�zuX<�A��e?�t��!,��0���,������yQYq'ͽ���f���"�Q@���֧d9PQ'����T �p��]2�^�7��R�=�&Q�=�~![@ۓ�u��ͣC���y;s���QP�I�~bk�
,>�g��ۅ�)"J|� :��ӰaH�D�;�p�3�_��X��T�5�D^���*�̅f�6G��3�)kλp�U������lK���)�!�kC}�[�̰�.����rW �	9�^��sD>H
��7����nc���Q���>�C��v�N�zC� ���.��*ܴ&�X#�1R�"��+�`P��Je���1A�AsLw�d/��/�ࡤ��� Et	�mKgG�]�n�ԡ��L�F��n�U����
�}�
��vgm�ey�ݮ%�66eѶVF�JيƐ��Ơ�]�lO����H��6#|��Z��F��M TE��a����_�	-�K��	���b�{L�qUPPohBc.d��������8���u�=Ɵ�ޖmZϕ��X�'Ld�u� �둹TK����ӿ�R��M��7�!ӊ�a�u�m�p�˕��-	,t@��<����)$��TC��M�8�kv4��2ਁa�͛��.���f����%,�/��%G֗�4��mt�m�[]���b����+�Mf�_k��⣛�y�5*��ER��[Ldae�wY�I�{;,eN���
�q�9ṁס�B��/�qm�pB_���>oW^���ԍE]ʂ��U:��vHz:%�nC|��{��Kݒ>������B[�݇9�;1��SF�J&��z������X�g��I:���j�X��G��W��ϻ��y���sNmq��ݧ7OTS���c3��������3�oMW�	�:b+YB#�e�`�B�j�`W���4?�+!M,����0N����}د������A:��W&��?ե���v�+ݯ�<W���G���a�!���۪���_�t=�ۂ��s��8`_���O�J��$�R˯�X���y�UaZ)�0 �o���y���΍J�uP���
5�e	�x�5�t���r�\�h���%rۖ�.�Y��j��p� �g7������!����dҹ��;��~�-���ZpG+b��{�v��C�MM������0O'=�P�
�L|�4�����aw�U����׆�R�B��Oq\/�ϛǪP����<Z[A���c�\*��!}���Z��r�>�P2�]-�{r֙�f��vh(�^L$Zϓ.��q��i����~\^mf�6W�I�Fu�bʧ�dpہ�(��G��Ih�Bz/�+n�UL�����{J�=͆�l5��SU>ϋ�b���b� ��X��'ik�"sI?!aA͢�c/�-6��򆺥!,B�IEw&HY����h�*W0�,�� H-������"�E^���+@rc�@��<�����(�,C
3�!�?r��;r%����ߓM���8�O�8�1���!b�@w�`/&_�����[��B���g6O�\��~�3
Y;8�����ðE��
��l������d9����Fo\�@{����o/='��	���ɿ���$h�e>Gݯyde[m���������f�-����Pu
�@���nPB�gq�]�'ɼ�`�|���z����&TG.�b������$�ty�������)\R=��'���SW�>�.��� -;�څ�0�����]M#O�`t<�\�Qˏ�t�"�����j�㖪;)R�G�+`'5��}�y��l%L1��w���7u����o*/�h�����im숋;0�Q�m%Dў8�N4�{�!����cy����B�nh��*�u�Y�0��C�N�g�g�O�$�:;�2���MK��`	e[�o�$�Z�����E,acN2����Y�l9�o����{���Y�*Q�a�s8L�F.�J��1[03�Z�"�Y,�iDcy���zx���gkvC�q�;=O7�����2�scn��L��;i�ts5�C՝7�?��Y��S]�(1���)l�>K�9��wdڜ��	��"�y�_S+�AyA�ԈyrP�͸?����R3K�ηg�&
F[�F$���s��9K�9�������N�(�+c5	�ok�#&���n�-N'���]C7Uk�����`�u(�%�+�u;O��N�_��E��	��!ͣ;�%#9����o��=�����[��r~�s���� Xί>1��7P�^9<W�M_�)���ӄ@D  n����M,P��Z�MgmF}���U�U������_���|]`��pS�|l��r=��g������3J�����bg祝��/4��p��G��\(�U�P �2U�%%��n�?�>�k'���7X}@D�$�U�\-N5���H�#Džn�4�+�dR)�����Ʒ�~��r:�i޷�E_H������~�4[A�;�c�x��%��u��H���j��)��AYUcfsg���]�
�" 3�P�|f��iiGa;�K�a7Vy6��(jA�I�ߋ*�����y�6W�.$2wƲ[�.�[M���1x%BW��~\��-�I�K�+����[�jU�������vc�H9Av�9�6�[�(.w��y��~2��-�o�B2Q^I��~R`)c�OѪ�?��%������iVˁ7�#�0[N����q�2�h̩�r;����?����3���}� �:�,�Y
��1TG�)�MX�78,6'z��X?�������b�.�zr�jߦ�_x3�ՕDJ���I��6t���rl�J!5b�Rފˆ�`W�=i(g�<�B(�@��'mP75U����]y,��I�w>j���E�<����`����R�m�V �R7�|�D��u���?��
��� ���	r�c6�)��?�wn���wټ��l?-2�I�n�M
35����MO����������B�y�-�;㇔�E>�tX��T�b[�gƬ��>ϙ�w������J�]y�fK$���A�cD_��d����P���C'�6z0�̶\VUe�*僠-�U;��Q�0��T,�(ޛaP�y.q�gד�>f��"��KQ����N����γ��6��*��A����']-Y��$�Rڿn�A�==:��[B>�+�@�Wp�>�y/�sc�Qk3�Iz�k}��>��v��)+�[y�acZ����p��2_�q�L�5����i�C*�C�f.�����3�j�k	����t��k��J'Km��)�X/!Z�TCXgHs,�g��)�֟�E?W�[b9 �'����H匁7U2���((�g�H��F�$>#ܱ�Qi�)?�C�}�������f��[:#�j�O�Aik;=R��n�`�C�<��wqiI/E���H�.�6  �똤m�a��X�'�/����� ����Ϋ�W�ݨ�}:p�q�&��������Q�0�1u��%�1�˴?�aq-�X��O_�}�Q��|v��b�^��E?��̒`_��ѤT�$b����ѻVL���0�U��h=݈d��Ӻ�����5�)�"���aXZj�[�|��'����0g����T�"�Э���.}���ԕH��71B��\]�1 u1����e�ЭV-��@�=<V��䩦���).���vo��2{�a�sG�M����w���,[m� ���*��2�m���tb}]˞F0.M�A�k�)��ַ*e^��3<�Թ�s�a���Y1�{�N�ȯ
��9������Ǐ<��q���~N��[A5o�u��yӚEX�/�Ӝ:_?vcN�%�#�CWB�{����-o���]��;G[P�9��1A��S!�{&3���]�ȯ�kUg�;=IUa^���X�T�GP����J���)I��N���X�e��S��X����ȼ�]�r�	3��"r�	Y�4+45F����ݛ�[ ��r��?h�!*�N�U��0)�JB�}s0�����@U��:%&��� @�Կ�+~��B����ל��ܤ���:�x��O�����XO��b_9c�
$|�Qz��z�������U���+�io_F"�4@��:��Jt˟T�>B�e�5�x��ItX��-�^������]��q�.��t�jG*A��{K7�D�����	dMJ���Ϲ��-��ѥװ@G�wК6q��&�9��(V�r��k�|=�N�P�+L�Đ��h��%��!ĳ��B���qW��:t�e�5�بm<������觗��&eE}�c,��2r@�W�k�B]�A�{M"3�����%�(���$^��鏙q�8Ui�6��u�^�8	�p'I���罶֟��͗^e��$
�}W����KUG����JR@G��m&5�-�S0����J��R� Ь���ickS��IZf�AH��c
��6>���!�!'�D���fw�`wY�(���JWh��7Wk��o�q-��*{�"l��^:����+�Cc%�ŋm3��'vԃH2C�a`!F��`�;M���W�z/M��'ؗ��fO��y1��1ĜvE@Rm�/a >� ؋�5A�q����3�6j�'�w�YK;s�������"Op?<_��o�������恤Т�W��\Lo��a'}5�	ܐ�D�t��_�7e�_�ݪ�����ҷ�@ϰN�w�	�����u�� �;������׿�x{D�7D��vP�/]4zD&�����G��)�V�����t������d�4=�V��"SW1��
*�;�b����B�&R�M�B#`o�`\x4l�J�ש=[�����E����R�2r�&������8.D��CL�ˌ�Rd�r��c��jD/v�@�#�+���m����lfÌHn%��8�ʦ4/Cw�ܱD�
�dy�2��?�n�=�*.�Y�����ӯ"��2Dg$l�$�d����g�3k�eV+�AvZe��-v{E�D�c)�A��������a�ً{v �Y���Qo�osJ�Fi��eC1V$�ϵZÇii_�3N\x�7�g�:i�;=J���Kk�2���n���Ǖ�;D�!sp���8ֈ�:�x䴐�S��1�^�)珡K�8M7R��7��	�K'��v�_�#A����>P�w?�s��F��ĥ
f3F?I���yegc�K�)��q��������+���	���g�#����Ȱ����ғ7�HѹӬ��(n��1�u���Ia�A���Z�n��<����X�#t�z���L�����Z��t�qፌ-��w��!���Zۊa�=�YP�W*2F���τ�`� I���/�M�^"�U��g�g4��i��p�Z�V[���q-�]�/PpN8+l9e��-���f��~���L����b�*�]j/a�?�+qo�bB�\����+��m��%����i(�?W�.�&����}�����F�ӗ��5L?BH�1_D �<����⟉�֫��!~�.:�2�iِ��WϿE�����4�97����z���|�u�n���j�Qɦ§�Uި$sBpC�5����� .b��P��5Oi���a��<V���\�JA�����;�gz�ys�����	��w=��Ɉ�M��%�_B�~w�-.T�K��v�ې��X-��a���Pc�MA� w9^��[���.�H���ny�#�5('o��FQyF���`jOW|��ڲJ%�g��3����V4���"G#��[�T��n�w�-�>��;e�����3����h4�բ��T���||G�gF)�����8�l'����R�Kߟ�WB�]b.�#���.�:ԍ3?����S��-���GL��X��8�=�s�ŭȚ����8�kg�8n��o[[ߔ�ϟ��Ғ]�v�D=�w��*ʯ�QƦ��M��ӝ=��J�mXV��M*�|�x�0�p��
��������ۯ,roι�$��?R�v�>�����l�p��$��׈W5=�í��xOXS�Iǌޚ���O����­�E�xX�UOT161�"=�Ug�MQ���&���jJH	�y;��IYψۼ�\��D���?˞��;]ng��Ԯ�'5�z��@�wBTe5���{�~��u�b�R0�H�,P}0�yI�fq"}���fK�")�Q R�7����S��uK<��b�m�|��s](^���tR���\�Q=��g[���f:`��2�9��wgs�,Q��II���kX �>M����)��Ƕ4��a~���1�^p�(_z��eV5�|]�ĸ�*G�2fIF�=3y��kD�3͋�����ܥc�K(�)˱�!�D�C3������n$7��=��W��9���i�H�C�7�Ă�0e�?�����3>>���{���C*�,,S������2<#:��*$����J����t��p��7��w�kn/ ?v�ʷ��+� ��B&L�m�|�Sf�������v4;r��d��㖺/ga}���l�ی
J�SVp�l�Ѭ��� �h�~X��a_�S�0Oc��r��l�8|��=���è�E�l��a&_yFl����?����1����U��h8w?db�%�u����0����;���)�TK7Z��w�'�������!��TA�YЈX��ir�;k��C,7p`ъ^w��L�u�X��c�� -?�@�h<�0q��O|�.�.ȣ�Gv��2n\a�9���@�m�}��a�,���ۜ��A����m�]`o��b8s�ac�M\�^k�ã�o ���N��ѹ�a���Y��{�-9N�3
/��9����W�����q��h�zU�6��oͬ`���ES�8�u�:�v~BD%��C2�n{)~������1�f�K[��9ڞ1�u�S�ؼ&n-�OR��3��1g���Ip+z�`��X� G�M���z�U
�����{N�����8���RS56��ȷė��~�3Ma\�6r	�a�+H���R׺xѸ�V	����B?#3�!ECy�дv0rDQ��}�8��L���������&�fb՛I��(�+S�ƍrN��%R�<����2�M��H*��Q�T�������:_���ؑ�!�F�HJ�w�����U����&
�o��[��Z��ܲ�ke��z��y�[eS�Rx��wt��i��l�������L�L�^��$j��ə�&�7c���n7J��
d��9��vp��]d-(�y��&�G���QV�A��C$�MX�ۦ�F=<ܗP�lhL2%m�B���3[�Kh��w=�UյB#�gqRA:��� 翩�v6<P^ڸtK��«�ȭ}�:�7Br�!^���]#/{(���ܬh-��(���$��2���wq���i��ʋ���^�*El��I� ��������&�������T��a��UBݴ�F1�Jc���5�S�q�S��%b� ˯��G̝k^<Iu�QAÓ�c��6y��򼏬!"�#��?w��AY�x��w��h���W��t�
̓-�Gυ3�"'�Q^(u~�"2+�- c`F@�&�������+�C���!"l�J*;(7�%i����V���{Of�01����@-1F/�_����/����`�H�P6��Z��]���-;�!�/���
�g�}�T�+���V_�Z��s����X�vTo��>o��'8��	�b������Ee��et��ݥ��l�r���mƽ�3y��])t�u@���6���$���{hrѓ#Iɲ��ő�j��z�c����G�p�ݿ�+5to���zf�ߟ>�=5�����nWrZĪ��$�V	���<س�i�a��MYV�`j*
\ӚF����Xjh��� �+� JtRP��!�o������(��L'���-+������z��e4�/�l������.Vm
��ݬ����%zZ[8���4�*	����%�yz� ��\�n���*�� Y�v ������q�MY�$�ڠ�+#�ñm�Ε�eQ��8iZ on�Hv3E"H�c���5Rs��DW��IB�{1��Y���Q��Ds�gZF�n|Jf1Q8����	�iz����ix� �g�Cŧ�0=E�ߦ)�2jgNn�wBzF;n�s����Ӭ2�5P]�z�S�Ĳ1�
�)b�pKaWrL"���b	����/�)_�J�A�O��~N�PvAx?ye��E�AP��E
���FZ��i?bB�3K):�+�������i.+}��	�)�⺿#��0�G'�c3�ᠨVhD7�����VX�(I�x5Xnuq
��D�^������X�`͙/F�lΕ#����MWB��Ib����/��ᨺ�ii��^B��%�9���c�T��W���'��0��6�b $g��jT?Mb���P�_g#�˺w����ǥ��ß���<V�]�ɇpIVl�������Uر�b��mC�4�b��C���/�B����n�}�\��|mǨ%[f̝d��?��~��"(�0�#}�|�ھ����v5��H�_�D{yj����������?�|��~��]:Fxiԉ��oֿ �ޡҔ1489��\W��(�[-�u�22I.�jS ��-�UY�s�v�pf�@�� )�Ej9��toGi�	�a1�ڃ)�V�Ta��A����A=��"?�y/ϳ���Qw<�j�dzQM� �����B��~��-�~�Kh�`�F�場���Q)�`�JcFބA�R�9�/[��.�{�I�t�!��B�oL�Q�c��ߗ`��O�G̭u��%���ǎS-OάVO�=.�#���[�*�	/v�(�_a+; �|����3e���I��p�\�O"׏�EG~n")��3�8�y'𼕅���2�=�����.��`��P�3z��z���$�f��/��ݺ��@p]$�� ���9���3C+gFU�Wv�ƔR{���U�X]�u��?�w��q�j ��0���U��x��8c*m�u��H=�|u	S��@��
K� �����4�ӣr
Y���?�����A��,l5Ԩ��}���F�5��a���O�����޵��8�ʫ�p����|Etr�X���T�)���cq�/�'��JS��O6�4K�J��uyzhN�C�U�w�DUQ`��a�9�z	�U�ϸC'z~4z�V���N�e�)
�Vٻ��4�tH0�,,���/jyd�9q����`;fZ��"��qQ���mt��y<�XE}aŘ=�h��Dd�A�v]#Ɂ�H�4RP˜�wX-=0p�[�!��������4����s�<Q���IpQMk3+q>��k���)�|�;���ea������CphU�_=^���5H�j*�fd�h�ih3TL�k0#�&���y5� ��K�"<)�*J!P��C���Kҝ���{��hxWQտ96+4�䚎H�Y7�va����Γ��V��?G>YZ&�G���"6Ce�4�ǐI���P�7*^#�y3d��7D�v���]���@q�2\~w'��/�����$�� ֛�a�m�=�N�.��)��}oAV�f����q= SEb}p�$�g��v�&���ه���'4��0�Ag��r��NμO�C�-#�f�|l@��q�����Eu�н�P(_���G��Z�q�x��4��HMU!�hh31Rd�z��0�c���h������V��U
Z�*L�r��']!ߦ�o�<'�T�x�c2r�����'ؕ>|7˯���k�g�u'.ᓯ���F��-�B2@�O<�;�Z��Il�Oj���-v���2� �a�3�� �(�r���K,���wӗRw'�>�m��ʒ�b����|�tM׎�kZ��LI���}c��� �a��=30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�ڜ4iy^�����i��]|$-�'��������f�j~tɛ��T��h�6]�X�_3;B�s����ݦf~��fcÌ>��K֯c���y��b����PW����ܦ"������T���
t��hRDj�Ŕ��V�2X�u�w�0��jH��w���vF��P� CO�2����E�DTr�B� ����8-�����-��
z"1Y��+(h��D�}1��2[+R��e�{_�r���UOQ��ʪNΊؙ��X�p�����\Ȝ"�;i8T��k�+B�פ���B0S)�^h�ᱍ��r&��������v���U��W>��"�?�~�L����� ;�wo5������s�>�cl#�6�P�8�o�$�u�U9L��D� 3p�]�<��Ie�W�]bA�+%���'�*5BA�@]��+����e��*l7��6?{�?a	:�Ǽ_9��L!!���Iˤ*�ZE���n�b��{oQ�nRIwۙ��,2�*��#��(�<�`��hHǄ�{���P^w �S|w�ɽ|�K�Q���脡�)�B��Ð�����?�Q�a�%s�#4�d��z+.�,֥(޴�h�S+|�'���58I��R�s+������}G�<��.���F݈8��]�����)��Œ�r[s�)���B�0h�ץ�)��������`[�������Pɤ��C�,b�.�}��B����(��1���p-�9�VMz�u ���:��~�lJ]��F仞�O�~�]�|���s�M
Kˀ��Zp���Fh#2+t�nXU�wf��p4�AgB�h��~M��#ꤟk�m�����'`Ņz]2��ґF���SH\۵��m��2�+�?���>�U&GN1������K.�_�T��'��T�Fu�P%GC��L�$O������ӫ!�w��JѓT�q9��`��'�k�}��
��p!�fz�j�"�r���42�����Γۤ��a߰tH1-����y}���M��w��T����.Y�-�ے�����lg�bG{�CA����h���|��զ����/7�0z"b'2���;tK}| ���]��������ʹ��~�@���!��J5�����fa�M5N�2�-JZ����w`$�8���L]O[B-��c�d�@Ӆ��8( ;Gko�p�R�A�c��>�j��#E�t �X=J�F~t�#pP��ΰ����a�2ʪ�e��}#=ձ��I�ܟ��o�������r��/�n��o{�%�$��E��Fj��i�7쨾	���gಏ��$��ɆX򶻏��[�~��,ߘ����8}6�����xBp�˳���>�~"w]cu��}�a��q؆ʙyDx����uP�R-ʝ�X�̥�?憤)�|�����j��p�	2~y;'��"B?jz�w#y�v�q�B�k u�2."���ĺDF���t���L�k�����q����ю��ϕ�Y�u�Z�	��g1��AM�@�V\��qpG�zYӡ�A9�+чb�\V)3-H*4��{�x�U��j�0@@n���V3N�`��n�jD!~`�hFN	�@L�e�4���H1��ݚ��e{�y�+��7����ޜ��s�uh�<4�YN���vɬ�n�K� ��_M���{��(9[9���xO��y���"�=s���7��N^e���Nm�r��}��H�,d���@�����s��&�NywI3��p`�^O:��Ź�I]Oț�� S��5���Y7u�H��������$�:���f�4um���x u;:�M�G,F�� O�С�����g�#�E��1s\���}I�O�%�T�4��%���?��)w�?�>
D\5���L��#�ɶ؆�ҾT).n�r��&z��{p�SRU��+�f�ȕ]	����ݱ0�a���2yUq�e���R|^�;b5�_���;j�ӐK���ݪ�S�	^���E/�5͍�&�8�;�j /,�l�|���y��zכ�#��/��		�H�~��xRY�/Ĝ�Yi8��V�rc52�G�'{>��U9��b\co����k9IlI�B������0ӵCO�D0x��64�k2	�b�'�$�||bE�%��07�xZ�g��|R
�8hi� ��+W_���RE�A�
������*���x��Z��{#�7��1�{6�^�n,j�M�����$��q|�=�p�e��,���!i,tո���˾�&���H��5:��R��H$�>k
��.~Jn��rL�ԯ74�ä�k7��������kqS�����3�4X���%8���G��:b]�r��K~)&@r�ѹ�:/�����5��r�T5�~�߇�H����:gE˟QO,L�_|�p0~��d��Zo��-���DD�O����ha�V"�82��ˤ91�6&����7`�Q=O���a~�M	3^Y[��Y<;��<�1\�f��Gc� ����H�����&�;�w��o�4�á�L���@�JV%�H�(�m�r�,�~�O#~�\�'�4���c�.���i���MT�]�����A�^]n�/ q��{� �л��M�
������ds�'#j�j'��؋C?�c��:	 ���4�MUT�'�*,, �ya��m�	S��74��D�F:��}�ߥ��J�l�v���O�uF���N�R@��ۅK�#�����s�*��ת&�1�q�F��$x����`�ʅ-�F���#�Px�2���-@�z�g��=5B4X#��`���z6�?�a���ϱ�D����B��S�D�T��3�@))��w$��ǻ�9`�6�_�d� g�&i���*6���A��u.o>�����WW9F�i}�Į-qM;?����9oC_�,D*�������%�o',F�P�1��X�lC��1ț�c�pשT�ZO��^P���u'��qyA�׬ŋ�����#� F��x,����<�յ�xw�C���x������[���I%��J�z������Iض�Gf��sU��`���Y����ЄhuI��^����6�Rm��t��1�"I'���6 ��h^��'C��p�H���9����zY�Cի�:�0���������Ņ�sO�gOF�y�;ݳ�J����ZJ�s`�/Nw�G��J;QW ��VqS�_����?�{��w�w$K�����l	�b�_�_d��d�B����<�K9�,���#"lS��=���;�G��~T{':A�9���~�/NJ��uhab�d�� Ƃ�@��W�� �pT� �/�c�S��A�e7�u$����	Ti.*2� ��ME���M�~zn�.[ c�D>��cο�a�U���H+�HD�rz��߸
��0�.+�bu��������ǽk��y@lv�XX���6bU��yxp�f�*E�6�.�3r����M{�B�s��#��{�e�|�s�.�f�o��@���_�6�b4�)��{tG0 �1�B*�7�U�= �\L0�Oe��W�����'�ۇ��8F��*�/�sJ�´������󫂿�CO�J��=W�Q�V�e�_�I��!��w|Rw\h�$G��Ñ��lЃ��-_`W�do�ڱ����@9�h��V��lOA@@�@����Þ��z��'���9�W[~��J�Y��^��|��~s�Z@r�r��� ǫk����_*E�D��e3b$}��Dk.�!� �͋E,���g��zj��[����@j�aԿ�!��4�D��H��z�Ʉ�4c�,�+$�<��4��a.;ǹq���S�yX� -��a�b����Ey�b�f��E2�.���^؉�I[��!�s�w>�K�{���|Y�'.�SI�$l@��_7�	�^?)�j{p� ����>Cw�~�U��[�أֈ�֭���
M�y����]?l����U���|1�'[��&&G�/&RC�����G}ٔ�/��&�1<4�F]��"/���4����>���	سgʻ�f<Nzc�!�ΐj����a� �vb$	o(�NS�Y�$RZ�{� r���5Q�{����n���e(~��K��I�h1�
5��-�f�Y���g�z�a��#�u�i�sp�Iw�J���+ͻ���������2"q��<�w IMlqJ	mʯ5k\G�����ؤ���J����0�R_>�p�(�DTq���2M��f�I���6�0_ɩ�|�_���q_����QC�UK��+K*�}LVJC�8��[��4"�/=X���j?�K���O}��M�\���%��]f�� XSf}�^!�L]IP����kf�;<%��� ���y������8���;߲��^�C�|�c{#l-g���e	�)�VQ��H٢�7���<	���\�C��}�fK4����	��H������*,�������,f�$�K<�x!%ܗ�����z�a?0��D��8�����ćkɍ����u�"X�}qRR��f�Ǝ�؍=�������Rk�
_1x)^�R�gj�n�[Q�E��`�,"����>�t�>$��s�ginlo�3���x�5A0e�t� �&p*E�>�K؇�Y/`e�A���j�CɈ�_������Ώ:l�����~A/��E�($Ƀ����~m̍",��� �6W�(b�M��G�O��1����cޛS�Î�E�<�Xs��ײ�4LPhۂ��h��|�7��3��������5��k#�%)�!<tt`&�x�-�hjŽ�܋�Ӂ
�In��OM��6o�͗8���d�S����{�J��+~���i����6��M�HL>g;�v��'18\$�WZ�K?�r�h�	]���dN,���F1"y�X�d��
��n��]a�-"���/�#�.\v�7h���N�TSOwD����D��ZDQ�pe\˕7�z<L�ȉ/[�Ȇ�)�l2��\�D�o��^˥֗]%���F�J����P7��LV�+��Eҫbh���쏵����:�}���F7�%���)�\�d�:+p)؊=����N���D�7=�0[�Sj�t���kRB��3o��no8�J�>��)ܖP=ן�� U?R`N�_�d��0e���@���8��k�Ҥ�|%�?�0Wyyx�o:jCw��'�Q#~�>�h�wZ��g9ey}4�q��K���	S�\T�V�ڬ`��n7o	7�*�` (�ES*K�wu����d	�-qX�nyÚ`����>��?:Q ���E�̛�u-��@�t�S�n%������=�s����� ���Tkw*i��d����G�!��`k�0I��S��^Td1;����_�Z 7`�/�ߊ�S�]���ux��XMd�Ln-n��`����c���Qn�[�s����L�-�]���m���P}��8�>s��7q�+���m1��H%k�5D��5s����W��Y�!���(��s_z�Ҫ�@|ϹEa��X�i�ӏn���O\�b>&�gk�b��2'�@1`�:�nn��pS燀�J������i��i�@��H��.�����$�֙�"��Φ�	yZCe`���"�J�Ǖ��Z}�-g���fw:o��q�o �"��ۇn�D4�'��g�|���/�o<��t����״� 6$�I1��
=To|�R�!�(���18h֪dE7�V�I�p�i~���ƽ#Z�L$�j�־1ƻ�Ƅ�����0����Wzz#k<���&�u�' 4X�z����>���0]�U��,�>!+慊��k�g;����H��Oλ��p=�XnH�Rͯ�ԡ����;Z`j�ܑ�\*'���7ܳ�-)�%�hV�K�^<�r%��?���wv+�-U @X>Ff6����������c��������7�i>B,�#�1P�io�o���� 9<:��u�q����g�0��e�Z�N��<O@�ғB*�4[���7�� Ӿ(e�eV*y7��P6p��?����ܯE�"'WO��!D��(>L�f�m��?�D
l������]��@��a��L����TP�<!�>G��QU�i\��`^	�%�9�j@���h!�]�V�5�^��g'����׷ߡ ������;�`�xժEʫ�y����NlQ�� ���%L�O��񧜪Z�W�;�g��E���`��ڤ���ǧc�(�ցZ9%�g)�l�|P��մ� i�����js����A�8�ۜ�	B�洽��Yw,F��%����NoQh1���ƫy�S��t��Y�[F�\�������i� ���?B�hťm	U�*[�����Y�BSl1Y15��2võ�hK屍�������Y�Q��Y��֔5�[�Fp���k)dU�ؐ	]��TuY'�|��PAVs�?�;`�=��F��J��aE���W�I醖X�F�s5��ۧ������v�{3�q��|��ʿ"�����"z�4T[w.��{tt��`���-�,YX���9Hۡvz]Tv�=9�g'+��}�߄��}��t�x�����X����Ձbl1��yO�of��1EM5�.1Z�9����/��s�]����{B4�|t:.�����@��_����Y��)mX{+�% ���͹�یY�U��ǖsˈ�X��Rųny� ���@��׸!U�J�'VΌ&�m�/�C u���[�*,W�7z�����q(��>��!L<m��"m��w,6���6�6��(��M �� ����A�+cT~����N�;����M�W�A*P^ut�A�.�t���m��3��o܇�D�ey��>]�"�!��`��ʩc��j�A��A�Ӂ�UJn�+[M�}66%`ܗ��p��n���:{��T���^����(t6��$�A�H���g1����Q�1��$����A�vս����]��l�Z��ǖҵ��"��������dz1��#i]��"�g�/�~'.�'�7SH����L{O�����u��w�D��eҒ�78d�<BH���v=��'b�M}��d/D�vG�Ԩ.���ɵ��|� ����=��(V��2��.Rb����d��^��\��������� ���I���u�>r]p=i!M��"g��!-_��ck�=ЊH�鿚�R��3��Ť���@ؗ�����rH���, K��R�)p�տmd���[�ݬ�Cnͮ?���N��}�H_�0�0y��	:`�M��23Q�ߑ>��m�LE}g�K.y�8#�g��K�_�ʊ+�SûT�<�x����m �7v�`xW�g��S`���m�ǥ��di�-���no�`v�O�E�>�QQ�Q�O���t��Uq�-"��j�,�$���*a�Ƭ�i����f�.�9�M3km�	VX5���{6��b*Y�<�]O��$�Z!>��-�͙ަ��w�[
�n|d��Y����&J����o2�g�Ȃü�8<n3��S�+���Ƌ�@lzȏ�ik�i��m�@,�����wKܕ��;�!S��u.��1Z�Z����t4"o.�6YǕ��Z6�gf���o'����"q����t4#���q|%ry���o��tU���_�/ ���I���
��|ʍ!rw?������2`N7p�"I�����t�1��37�#�C�$	��F5��$;u���{]�03����!#�ŋ�Z��u3_4�h��!��>Dl�0�k�U�E;´j!��#�R�nk��S�l���ߓ�c���C�����X�w����.a�h�,;�.8�d1亢�}�%�;��)I�h�?���a
r��^��i���v�OHU��>Α��x(ܱ����^���=0:U�k�Ҍ��/>�_U#��P��o%V@�A!9ĿQ�d/��xS�v����ae�����ؘ�$�ZD�*�,�9�A�9I�F�xe:��*�ok7+��6�@?:���d�=�nW׍�o<�D'@L6m�U�?�| D�n�6g��n"��������L>���
����q��Q$�ٰ��(#+��^��#�fj���dJW���H��璋u<踂��?�� v������EJ�x�ER��'�\��٤ �X%��g���,�/�@Zi�.;w��w�N�t��b����ާ�Ɣ(C6Z��!��NlC��,�3 �Ռ�1�@l��XQ3�ɢc8o�M���B��E߰Y�$�FF�/%u(�U]�o�d�� w*�3�qS�n�xZ�[���\|&%!m��En� `]�?��0hM�"	�Â[�����խ��Xl�e�5"CvK�h���C����Y��:��5%Ş���o
�.�|}9���r�� �'x�����sY�^Ï=	�"J���a͛)�����L��*����c� �7��>�v@7U�1|�y�.F��gN:ŷ�ç�3Ă�v��[��-�����ĬWДk#q;��X�Ht�fY����W��-����N�_�b���l�m*@'�(lÝBh\b���o!��n�_�w�|��Om�*h���p��<���]���$���w���|5%��@���	Q�i	+����)8����#�!4ޛ�O?�TQ[e��m&#7M����y+���,�9��7��6Tz�j�/a8L�Wٵ�Q+����Ѱ}�2�<zW-�l�F�i�8�=]�����)�t��S1�s��S�D���;�ר�d�)Fvߟ1`~�Òc�g��Q�S�9C.���1�R��߬���KV1$FLp�J�Y�|)�.�X�6�/>���
+sx���\��4FH?�+T��X5VnwF�P@cAG�ӓHt^M��|]��vm�y)�a����e�h2zUK�&�+�3$}ە*mjq�2��\?}��>���G.u���w��+�F_���Ht��7sT�]�u�x�G#L��W��|���[!ċ��*a�T�� ����
�K8���gu��*!�֮fZ����r��P��B��r��kHg��H��5%ߐ�A�|P��vh�YǢ���M�)<�.7�44��b��-҃ٚs$��L�Jb'�qC�ج��ns�զ٧�Ԧ�x߯��0�yDb.���K�t+�L �`�=qT�����'u�����(@� ��GTJ���}�aҕ�Nzv�-*���`w�y���,�["����ъc�2�d��)�n��䫷(�NsGK�Rp���I�c��G�Jq?���t��=*��~T��p��4������a�DNʊ��U�=���`����7�aR��f���R�\/�&���"�{rU�$�)wE��d&)�/Ci�So��������o��$G�f�!��$�x[~��}�xfD��6o��ñ��BP��˓����~S\cUߐ]A��uA��f�cy$����;�Pi"�*�8�E��fT;�\X�����j�S��)2^6�VPjZsSw�v�y�"ۣ U�'2�F�׼D&~0�T��,(O���<�U���l�n+p�m�Y�I/:� ��^h1k�l-���6���QI�GqЅY�Uk�!i�+��axm˞N�ڿn�YS��lHv���cK��>�/�"�D;��� nb|C��n��*���hU��-b���oclIn7��w`�\�QC�*�$,���<���dK���w�Ww���|7݊ɂ��BϷQ�݇k��5)���[.I�#���ݸT?|1�Qإ��8Y#yxF�\�+��,��u�y�Wø�M�,�1�'8����7�w+L����/*}�P6<�=v�#F���8��]n�Sʕ-�)�����q�s*T����լ���m'֫���a�`��쒥��Z�J��hC0F��s2��ݽ�n��MZ?1f��p����Szud��=j���
~,]"��F���+N�b?����� 5
0O�l���"�F-��+��XZZ�wz7����ALu������f�a��,�m��q�D����Iq�j�2���k�����m�$2�n�?�dt>��vGӭ'��%��	_3?>�K̫�TS�u���G��LԆx���O�RS�!��V��;T�������m�1Őo��i]�!�*fds�g�r̯����i�7��P}[�i����7��U�M�n�ЂJ��Sƀ�0�Mmsu}���Y��wS�s9�-��u������b�4C{�������ŧI�F�����0-��b졑�{<�tP�K�@��O�ܠ*��3����}��@��5�&��Jڞܼ<�a�uNW'-o��#`wu�l�=�6��[�����c/�d�J��!/�i�(OIG�pT��œ�c����P$��ttez{=O��~��pb���4�a(�,�o䕫K�Z=�/�%��!�u�������n�7�r/4U��"6{79p$b�ME���1ni�Z7�#����O�4�q$���k�
�@�0���~�=������U�64m5�:�BUQF�8���4F�~�Wc�]@��?�:��˱�y)H��q�YP����˦ܽ������+�����}j[d�.�i2Cpx�Վ�'��j -whJ�v�k��� �#�2���\)DK{���>��쭥�tt]6�i��S�4�9Y�A�v}���W1p�I�^M�{o�6�&G��Y������#+�h�A��3��}4۰9�ZC�˺��o�Cի.@�L���?,3Ӷ߸<�΅/�rD�6D�-�N�;�@�(�e��Ҥ��1�>e��9�{<�R�%�҉?��Wށ���%�h�Ah�����X��DKl0N�0d�2G?獤S�M��9g#�x�d3�~!v�9�B��Ù��9��<;e��N2G�^���MMr	T�����@��z8��*PN> �3e�`�,�ߚ��
QIB}���K ;����Y���m`u�KD��"֨�����|:^����:���\DAuG�:d�6GGy�F�v�O�o�ƿ�/�g��*Ƴ.?\@K�}.�O�>T���S�थ`)|�K����\z m�l�D,y�H����{7I�)3�n�*��d�tzj��5xT���ZO��	3ȚiZ�Yq�¡��y��/]����U6�2g`݄��a����5�e1��<$�!j],K��ݯ~���6��PϮA/����8=�j�T��uJ�|��la�zĿW�嚬Է���*�D	��H�[��X�R�����iiC�V&�E5WFuy7�����j֝c�Rn�}�k�XTln��U����0���OD��x	�"��k�����&ɽ��|��E��9�Ֆvx��t��Y

!�i����E׳�`�E���
i
��}��-<��Y��@�7^L���F���,�)Mw��z·$�n�qAm|�����JS�� �,��������w���Ղ����7��Mw�>�J�s�hJSI����2��5���g�k��������T��끯AUӸ�(X�"?%�������?��d�.^���r*ɇ����:�D�^@V�:�Ir��z]��~s�;���ҵ�:,���)XL�#�8
�a'����SOÌǖ%���-�a��"�
� =x9:x&9�E��o��AO`�a��n��<3�?��oX;�</<�-�+Z0Ӭ�3 ��yi�&H������;J� ��0���L ݲE��V�h�H.��m�{ڣ!9�*a�g�\�>+�(
J�-���DX��G5 ��p`񥢇���z����S��%�ݝ��������=oAX���[l���͊���fw���\�j�m"��V�d���V9�(��E�}�B���Z����h��T�V?jc;-�h0���UJ�O0kQ(�٣K�7(ù.��̴h��}��:��D���Yq�V�B�[����y
K����}�j�B8�O�E�N��<WQ���^�I
S��o����ݻ�Hd�1���iWVm�\$u��@����1�����u*dߥ�	Ͼ1��/��t��F9"�q1>�v;pR�=���kD&��K���7 ���-W��M8Ga��$�?�f'�E5�������K�%3�Z�D�&�#�����R���3���������З�i��Aw���7 ��0Rc o�ЉKdC�V���)o��|˰�������0ȱ�y	�:������Qz�>����[��g��y��+���m���=G�.���jC�0:�?O�[쒭��V4�4c��U��'P;,X�y�sڸN��a�L�c�4���ٞw��Ց��������8��p٠Fsd��7R�`���8�{�Z�-�s%,A�/�,���=���ŉ|e��&�#`n�-U�ˡ�qT���?����c�z ��ٕ��B��H#�wn���hz�	��a&�Pmh��=LN�BL����ͺT(���h���I�(=��YYy����9� �E\i�#�*��'�lSA�.�6�������W�]i��8��`N;����^iC�akD�����
�eF}	�'�&PD��ɂC�v������TA�_�&^m��P2�0u�9�Ɂ=Al�c�/���f(�`�X�l�Ў��T=��-�x�0����+�Y��-��[K��K%_��Ҹ{�40�I0]���x���i�(��T��녖(�	u��^��Y�Ѫ��t`�f5"�\N� ��S�^'J�C�p:�֏���T�YUQʫ�?0R�6��CӼٖ��L��ƿ���M�e#J�,V����Cz������J���WX-V�E_/P����oӉ�w8!�$�n��m	la+�q�O_��ydK���~���O9)��2[l�8�����4�ݟ�����'���9�c~�>�D{�ͭY��eߡ��T?�6M"�g2��;� #�(�i�L��� xe��@$���a��.�� ��E̲lyi{z�[xD	�J]�=���O������Ǡ��H�tOz>i�đ��l�+ ��@8d�=������ћ�g<�X�����yb�{�rB	y��)f;�-Ej].���:q����\a7sU���i�{�e*|5.�ܚ���@9�_.���)�J�{�i _v�͚h��ZP�U�=����`	�t�~fy��m� ���t�U
�X�h'��G&B�/�����l�BGY�Z��S}���<�J(]z�9/ߟ�4��0�*8��S	4t�ʗW<��x��S����y���.��n��R�8	˄xN/{��twZv���|?]�������{�13��_�͇��������k�M��'=g��I�3aDǈ�3�%k������[|�9FE��G^x��R����
9�i�G�f1��fE�{b
�S���'��E�#��n��X�7vS�z��3,�-zM�C��,�$�zqY����<q�� o��yW,�$r������X�������O�[�e��>(��ˋ��Jk b�4x������k�8*��u7��������ǐ5�� X�o%�(���W�N�/�*�Fª&h�rB�.���v:�&v��R��r�`�u�~��F�6��Z�:D/ߟ�t�L�42�-��&�������kI+��ӌ�,v�.a,<*"�z�i�9.�&Q5�ܳn�UOxe�a����
\P3�"��O�;�f�<Ú��Cj���2 �.:���H�P����y;bz���#����0L��]�eV�9$HF��m�ڻ{9�Ƕ��e�Vn*@���E�\��_D���kpx&�l��]��6�S�������]�ﴇ��U��Apl���0��� �KC��"ء��Ԏ�:6m:_sV�l��bk�@]�^�Z2��Қ��	RQVW
�;E��hH!]��w�g1Q@]�cE)(�NJ��PZ��8}�n7��-����n��B�Eơ��
c�t릔}��BP�O�a�N�l+Wi'o�vq\
ko�a��û�ٱd54Å�2Wn��\<ҩ�#@���h1_A�ߞud��T	���#q#�j�^��Z-1Vv�~j�$�H/\p���ľ�g��5���E���ej"_�E�$�	�!r�y��]LY�C�u�&����3F=;���k	:�Sr�R�Sg��jJ����ڷ{���Xl��I�@��vr��}�w!0��v�#%����y�`ſ����ĒXYG�JP�����:Z*��̎v6qk��^5yx=Gt�&j#����Ι���QO�k�_�|1�sU�at�Κ&�" ��8�2~W�]���3�!y	ks��������l���uMf������6�w� ���q0�U�yݻ�c�M�M��_��|�}��'\�����Q5a?�<����M��g�4��Um_'1Kk,Y�y��4���J��z��<�4�P�_�uƶ�������y�
�F�y>����RY��۾M�|��1��sf�_����
��蝿ʉ=+���`��-.���Y����7�裏U$��z,�ٖ�}B��#8L��UJz��ZZ�z_�}�$��Bm�&�S�T��L�B^������z��:O������+p  |�i?"1*�]� BA�~~.�}��1W�f[i6��c;8Ì����C���D����15ۦ��ީ'�zP� ��q��C�_s���ו隔T�̝�-^�@�P���u@�⪻pAm��Pٔ�H`8s�o��Kd�q��p���kx���������E[�Su���%�¼�����5��IQ��3��,�K������٩���	�u�ϥ^,�5��������գ���"b"��ʬ��%^H�CW�Sp���oc踜��YH2����0S^w�O)�Ʌ���@BƸr��̌�J�L
����d���? �5J�W��+V�i_���?����wy�"$hG��<�lȍ2~�_��dL�{�4<��0��9��y��q�lL��e���G�ݠ^��1�'���9Q��~{F#G<R�����������4�w1z�Ȇ��I4� ��I�*���U��!f�e�P$#;g���$.�� ���E�_;�Mmj=�z��[�����X���՛��ܾn�ǁ��H���z_�Q���K +�����si��L���c���?z�`�X�E
�W*)b.�V��\y���fǆE�.3�[�{�ԡ�����s��*{įZ|6�.#�@f��_�̫�[��)��t{��1 `maͻ?U��sUH���5���(�52G�8y�0���hI��~Uk{��EN'X'�&���/c�ʰ��/�:;YG��x�>_���<1�];϶/�-�4�B:�K�H�!��	�
����<Kt5�Z����-��^�މ	��"C	,��N��(��Z7��]on���D��.{b�s�W�N���b|v��eN�.�Fh57�����=.`��Rn��$d ႰH��&3�J>��+�⦽H���c�}�/�����!?*�+J��ͯR_�\pR��D��	���^���^�/5.�~�(��qB�2sɌ��nQIJ�w6�3<,���g_vkq����%�C�
�³3VKg��L3:U���'�xK���/y� X�h��FK yN�,��"f�\��}%� f�q�XP&V}^M�CI-�����*0�%���]�m�vN����F�uO���m�AuL{z��9�c�˜ m-n������Q"�e��V��_WԚ=�g
��N]c��-�}���f���eH��~������oe*�8���r���+]f).KY@�x�q���|����aܟH���8���~ݠĤa2�x�T�l���-��.SR�����U���h�S�'R��_.B�^`\g�~�v@Hm�{��,�9Q�*J�t������Lg��lLh<�5���Rs�A��xޅt�$m�
���(��΀�/}��A<�Q����r���;����,��B�����;��x\(��� B�S��*mI�0,�߾��q6_��(_��MGb뺌���M���c�,���C���W�UK��t�^�H�PEE΂e��c���3�_m�΃���Z��E#���!�/?`C�����j"$�܈Z��m�n�H*M�;�6���U�ʩ!�H�Y�W{�)��<8�#��v��6`�j�]H	��g�U��.D1�g҃��J(i�Մ�1���]spw���m��T���"��}��W��+z�ˋ
]%y"�%�/�	!.��7Z����I���FO�p�y����<DNw�e���7?��<)�9��$;ȣ�X���<WD�d��
��Ԑ���Ǡ��%wa�V\�W�B�b|	��"�l���#������F=6ς�s�1������EGp�2=0TJ���
Ř�6��-���D�O	���R�"l3����+@?�����ږ����� 2��R�
�|��do���>�=0��Քݟ������(�
0t��y5��:�EO��ucQ���>&*�TC��gV��y<���Ι�K��ʱ�S&T��[W� �:��{7�Fp`�HO��@Sg��T��KA�d&?-.J=n���`������^�Q��g���DC*��"�_��Za�|����T9=uF��G.h�L�ʓ��P���8�!O~���T�H�X�X��J>Ŷy}���f!~$SfE��M`xrr>���2�]�&�6R0��2�]�W�{~�3tϩvW��d����LMSΫ#m�տ7����Y��-}�6�~����ymb���C!V�b�C��ֵ�/�6��O��gG0S�<b���!��t��,��7���݂G(���\����co@)0R��[nJ *B�"�a}bN�ع-��jv��w³��|W�n?[mW��~�c�o-d$������b(k�G6\p:��ksc� 赊���t��=���~?��pHp_�Y�E���aN��U鞫�p�=@>K+���O�ol D�ъ��\/�<��{��{]��$H_E/�I1��W�Ci�k��ɲ,�92��Z��$�����������`J~��lߣr	�8>c6Zb�����B�'&˞M��Z^�~͠�c�א�-��`��ر�Iy�d���uDPԍ��n�c����Q��ا�7���%j���Th!2)�$2�����jEg�wNvYv��-˖ ��x2ټ���eD�{��?Ƨ�w�v�K�U� 5�-���9���`�YW�%J���1�8(�������G��aY>	Ş�^+�u���	;3mr4m��@��`i*�ջ=�
k@���� �39�ȸbp҅��D,�0�E"N�`s@w�
eb�a�
�[1ˆC�l��{��KD�ү*&����'\\�^�hP��˜���.�V��K����:F������sg�9M|xZھ��Kp�_%��hH򙊲3�9*pe�E�N&*�Fw��}�/��k�+D_�n����N$er3�f�`3cj�,����I�o�
� a����D�d��u5�����F���O͎�C:������ Q��҉ux��:��G-��F<guO u���q�&)g�WFlr׳T�;\&E�}�FO}��T*���{�J�k)�ι�	�\`��o��=��nǑ��۠ݨ�)�;�n�%�J��zȗ[�f�XM�w�#�q��� �t���N����NLMJ��S�U��L�����)�f
=5+�֢�_s2UjC��K��hܢ��a���`�����D8+��j�o��§|�+f�~�ĥu��@���v暼P�	Ă�H��>�O��R$�L��M
i�cLV��5}(�_^p%�����@�ÝUc�|��L�4k$��l�u�;���0>~�Ojqx�j���k�7��$��P}|%>�E)����x�ɝ7L�
��Ti��i�����6�E#��
���9%�GB�da��S��&F�7h�掀�)@,�k�M;��o$�.Jq'2V�{K��,ᱺ�c�,�P�ч�������膪N��݀���>6��Y�jJ�S?�]������n8#kB����1���C���ⷁU���TzX�4�%��)�+߭�ǚ�=������r�4���:�!��խ�q�r��C�e~]���&��Sz:J�\��LL;��;y���7�i9��Ƅ�����~��2�az�}"�<��(�9��H&� #���eLtO6a�m����3������;��<���O��R�� 	X�4�H��z�Y��;�A(���(�n�	L����o�V���HwXm��_�	�9��(�M���H�����S�X�*\8�����p�3��m%援!�RS��"��'R&}�����cA>	��l��7�|�] ��vW�`�>�й�mHȆV��5��F�Ɏ��k ��(TF���� �2��V%�4;�D�h�,�Ɍ"�5LJQ�/����M(���i��y�} ���B5������ B� ���w
1 F�4�}�`�ƭ�(�ry;�b��x���Y\<��	�6E4�n���4[�����e�	M��N��`�v�AZ��������w�����{	P���Ǐ����<U�$2����h��5��<�^���&�Q�)��X�Q�:��TJ�+�xӽin��(��2�Y��U���Jg|w�Sf_\%W�6ӤQ=�hD{��H����_��(�}qc\I2�E}�SsQI�:x6��E��r��&�__Rq�ɶ3S�C���4��K��L����P�y�[{�/���X;(��S2K�;�����Up\���%�+�f+�X���}߰�*�I�,6���ѓ+l%�hQ��v�ז�<F��4�����"�|'V�Z=�c�~��,-����C���`�Q�Ő�t�ـ5��~BCk	ױϓ��!4�}��%ffJ���^���h��+&*!`a���c��7�f
��KZ@�x�q�T���"wUa]��";�8|��_�Tĥ�`��MQέ]�����7dRtQ��dTQ6R��J��t0R	),_�pw^�V�gHY�7߯N=�D�, �e�ka�t ����g]�l83�``�S7�AH����t��0D�G#����a��/~�~A]˂{}y˹�����JuJ��&�4�1aϯcNП-g����wmh:�5����[4��И	c'�d�Zv�0m�a�(��FGP�pLw����cx�6����nt]�=G8~�BpZ1ŕ��cz�a �9�g�B�C��=�����n�������<��/H�/,�,�7�{/�$Z�xE�A����)^Ai�I3�S���2�,Ӗ$ܯ��c+�8;R��v~�s���Dk��Z�6,��]BM���0c]�,&~�b�c�ǐz�p�2 ���L�y!B��i�P���"]ܵPw���7�#�1ع����jS�&��2;?����k~j,Dw`Տv�U �6� �k2�TI�TOlDC`��=���\���l����(�Ko6,-zY����r]��H71h��w��sE\�.�G�&Y��)��h\+���9�3�.M4�`��R�˲���g��͗�@�����	�3˿̸4]�'�D~<���YN���@��e���Ҝ6�1�޷�~؉{4E��b�ҁ���O�yɻ��h�Yw����NH��RKd���(7*yn�i�E#�9_��x���vNK�1z��z7��܃���%Ne���N*Nu�Vp'�E�@�W�}��b����@��dN6%3��`�IL�VK�X�I:����A 3�t��PϬ�C/u���V��Ƞ(��5:V����2O��T��u
T :\2#G?�OF� �O�8�о��� g�I���*�&c�\8�}&�O��T��^������)t}��ۈ�\r����<���@a綕��/��)+\n�>w�\7%zb�A�	Wp�@������7�ȒV�Q����Q�����;��Q�U.�__��|��dIx{�5}Gɢ]���9jUCLK�
�ݧީ��ޯ�Kf�����#/8��j���m�|�BYy�ķ��~!��|�"&	��H��0��%'R�>�ٔ�i��VV�5O�q޾w	����/֕�c����?�k�Ynlf�AM���0м~O<+�x�'6'k�o9��_�ٴ|w$JE��d��jx�;A��a
�Hi�����T��N�E���
aV9�H*9�%�栫��8��7V���x#m��f�,�lJMo^�r��$�n�q9l��Ǜ���꺀<P,�C����o-���E��z��//S�E��>rn�k�JK����j%��%ۆ�Vkk��Θ}e���~ਹ$��K�Ӱ7yXΊ�%�
p��=�7$��R�&���r"�-�֢T:�#�V���2@Wr��7U;�~kz���t�:$>���_�L�{z��?�t��Q�K ���ft�e��)ac;"{!�����9$�&1̻�&��w$�OX�a{�@��>K3�By�gj;���<��>�#HӤ�C �}a��H�o��;B����V,��N}L��=xV��HH&�m�ͅڛ�9}�1�_PC�6�� W��%���<���?���wpXC���w�����S�H��Հ%x���~��5��AP����ٵ��7G��6���3��T��b�mV�{���L=� b=W�:���%��Q����_V7��;%}h(H5��!T�G{�Q A��C�y(����{,�`�%}�u���ϰ���NhB��/��!�
Cz�}}�B0��O���N�g.WI~��V�	
K�io�̖��6��|}d3���qWN��\�K�����c�1���!�d�Е	�HH����\~�>  ��,16��v�^�JeF���<g{��𾺖1��\�%T��E��?|(�a@��w�Ylo]�#9��嗼h&w��u��=^���G�	�r�A�SG���JqX���^�[�8S����\@�Nr��V�W�"��}B#���*��@�̿w_��r�'@�Po�mZ
}��n��qK�g^�!='��&J�܇qX{����1�Ek�^��\�s5��t��c&��v$v8�� W`�����!Y�.s��2�g�����Ȅ��[M�찎y�ր�MߥWc����q^��YF��wn�M��t���>]bw'<�9���|�1D??p' ��;닷��4��UMa�',9�)y��#�o�����?4v���?�lƖ�ҥՐ���ѡ�Yg��ɜF�\.Ӹ�R9�9۞�D�\'���sF)&�px���ZV�}�������`���-#D�9Y>��������胎��z�b��v�mB�(�#�õ5�az�t��:9m��4��]���BM7���}�Tic����!�sj,��F0�of1�Z$ ��%i��*�	F��2A���.�T���(��W�Q�i�W��>P;B��Y\Cx��Dc|��+ۆy���<'�LP���Q�C�����(���i{Tbw^�^�#}P�Mu ��2�AMX�0�L�(��S�����Qh��j����x�J	��^�o�n�[��5s��%��1��ː���I1$���~��}\��{��c��x;�����u�^9��z�����i8��k�"B�~���,��`�^(�C7�tp{�яO�w�|�BY��ژ�03���]���6��6�� eZ�R��ݬ�J�>��LtD��
]���)J�]W�4�Vj��_�W��޲ԅ�wY��$�n����l�?�_}2�d,߯��q�"%9j����4�l,>��`K���}݀J����f'�8G91�Y~[�';��nt�{(0��=�ۣ�W|�ب-^�)�� �¦�
t�|l��Y�e��x$f�L%�I�yCr	"����.��Kj�v��7;�eK*��^7|��6iA�?˔$�����d�W�^a/^S�u�4Le-�m�6�?8�*DCpt����_TR�s�6�L�p��{�T�U���wt��)P�]<�@^��N�i��j����[(��7<����f0���c��p�I �U��T��\Wx�T;E#l�*d�m��
�� e��%\��hi��D�Z:�;hK�͈/���}��X0��C��|ۯ(���Z�T��,�lT�H�����[���קс��	��`�8`H���zB�+���Yp-�F�\#cF6[�8�{��4�E����(�]*Gu��pY�?j�7c�l`�tbf�m��t���=�~~p�pg�R�XA�ǒ�a�@���._z\���ޔ_��	ޮ��s �0�a+1���͠8��m ��s�'w����\��O�i�R������D�.��h���RW�_�c?^���g�G�腟^\^�O,�r�˹�+t.�t���g�Bl[f��$X��!1@A�{L�t Di!��i��7t��o!\/L��A�)�V�W���K���l��h������x\������#z(����o5�2���@m8�",����l6�6�`�(���M�$���k�QZ���zc�f��/��1���f����w��PT^�������┣�3|h��=�����q�t�����!��Z`�-��{�j�K��8����nn"zM֒�6�ٗ$������>B{bBP�c΃R�p��Ӗ6O��9�,H��g'�V�OF1$m��Èn7�7�s���T.1]"-�P`ِ}�0�2nE"�Z���Z�0��Z��]�"|��/\�.H�!7��3����&)OcCF�(�ԛ�o�D��ieH`�7n�:<8K����>�r���]���$D_���J���<w��Ԟ��<�l��& V������bT�-����{�����i���&^�ژ��B��H���tpdp��=��l��G�H#Wk���?c0�~����R�ҋ3[��ڧ
�6 X�c-�<�Y�
�e Az!R~9|�K��d�:QN��>��$q���Ѥ�����0C9�y䇝:V�V�6�^QG'>UO�c�g%~vy�q�]T�Kq�� �HSU�3T�6�F�,�	0��WB7l `.T=�6�S��"�cl�:l�d���-���ne��`,	����o�)'Q�.���2����l-X5�`>���0��� ��Z�_��iz��$~̃�kc��W�5q�x����m�Y�N�����1��P��~u�C��T�Q�Gn�;�M�� �&@���C2i)���,��o�n��dS����!ޟ6.�E�i���'t�@"V��@��-}�����#�+���MZ�Ĺ���"%��Q��E�{Z�#�g��>fu֍o]��� "ň>�l�4Y����|�t�-mqo���tK&�_ 4��I�y�
��|5#�!��H�(����#7��I�1����	@�����#x�$�����N�����M%�q�0�7E�U��#)б�P2�u��04VϺ�W��>:HO0��cU�����9!�����k�h������QF���ιo�.��X�]��;�󓜞��;�6`�8=Z��׳��1�)ɺ�hT��Gr��2�\C����v��U~Å>�Y��槱�;��TЃOŘ�C'���匵�>�}#���PK�o ��I�9:�x��=��M��,2��.Le=�k��\�zm���y�*Dڥ�/���[�Ӽ�ep��*�e	7�;�6n��?p@�Z�1�ˍ�WM��TT7�:��L�@dm���?��D�����w��N��Q����L���?��J���~w��|=gk�aO�^������ij��#�۶��s	_��8��X�5D� ,�С�s��{\x�H5E��wD�͒�
ψr ��%�ʒ���%�7Z�;�ͭ΍�j@�U���F�!��(9��Zw��e�\ly�'K��.��iT�v �Nl��8倲����B�����CXYu YF|UC%k�#-uoO+#�V��)�-S�����k|[�\rm�גc�J� ��]?���h��	S�[�̣�{��SY�l/X�5X�vAl�h�k��9�F��Y�T��R壍�5[ܘ��Ĭ��'��C����IH�'�N���sO2�y�Y=N�������a���U*�DD��T�sd���OI�mq9��s�v�
bקƫ�P.<�J��i:;M��:�xӅv��k[�Kۈ��
����J��q��MÎ.6Hj]�1F�W'���8��#�Lи�ն�b�"�b��*�������x��b�O�o�g�n+7�w�B"�E�r*����Z�<��up�x;U�kw�k�|+H���s�6��Q2�_�\�Z)����>���Q�j?p��Q�1���I#�F���}+'G,�!��~ì8:�tG%ݫ8���+�+�!G�ȶ#}:�`<�Q�3�mFv�,8X�]b�[�	ښ)��k�	�s��d.��A��^�!֟�����`t�ݒ���N93���`C$���癯�3���#=�A��1���p�O���zia'�?��~�]�]�Fϵ��x��{���SM�,�
$���4��OZ��c^*��{�-B�Ώ���_���b~� �c�o��*������sB�y����PV_k|p��eT��\���O�i����K�j��֛32�<}47-�ϔ�jǋ�w+v�a�o�? B#?2�O��'D�9���L�9�M�
0��������&�@vY���2����~10WzY�#]���'FG��Y����؈+�j���!3Z�74�(8��h�bw��}�p@[�]��3{F�����p�D.`�2��NVo�@9яedU��L(�1Mn�.�{����Z�1����'��)�<���h�1���c���׬�L�K���\��Tx�5g����s90�x\�&�A��Y��*���چ{'�eR�N�{�T(��K^�' �-D�F�ɛC�Ӝ��MN�\+3�V�`uS@�������I��L5� �;����f�auw�h�HF��x�8͐�A:+>�3`y�{���u���:�G�9F>L�OB�~�n�fbfg����³ֲ�\�3�}�mO�?:T��z��P��L7s)$G�ꋈ�\"q�������G�E���)�ՈnC����zSQ��Q ���9�v�s�C�B���]�z#o���[�Z�Q	�U�Y�j�,��t�(��5-��/� �I�j�gK�d�Wh�V�x��Y���S�8�ojm|���|3N�	�q�g0��B�3��YҼ��	�ΙH�sI��NR�^ĉ�O�2�Z�6���JD�ŏ������<�Ds5Ϛ�I�j{���|��.��6�a@�^_�-���)��{��� ?fa�zTT�:�TU�������@��T�FF[�yo�����ø��U�ʙ8��'�R&�y�/b�簊�����G9
���w��C2<p�P]Zv/��c4��ҁ
�����	xq�wר<�=���K����~��ZҖ����2�w	�h�N��TcZV���\���ے�q�{��K��T�ǭ�1��@�´e�-�Gh�85���"����Ȱ�6=��/[E1邯
��5�J���+�خ��`����Y�n�Z��W+��rl	&JE^����\�(��T�/������М��=�$(aY6q���2Ҁդ1�Ii��6�{���U_���q@��Q��C�|����Kf�JL���tqw��]p��/�h�X���&J�KH�'A��.,\{�'%"��fI�@X�6�}}e��;�I����@��?b%������-��ڸ��t�����<� ����ĸnc7.�_ -#���߳�0(Q�s��q����x皜��I��m����J}ٚfD�ǳ�E����㻓*�����x����f�qK��x]�D�r�P� =a�"泀��8���=��C\
��
,��Ƶ�^��9`�RҍG����h�y����X)R'�L_m��^=�g���U��,s�I�,^�ˉFt�=���ZUg�',l+|���'�����Al��t�{,�R����Z�?��/FwA����&��S�8���ɨp����o}�H�#ີb�|A/(X���?ߨR>�e�m?�,|���<��6�NS(���Mf�����Pi�ڂǺc�p�������vǔ�Ɠ��G^�P$� ��\���s�E3L�q����l�D��!x�+`��i_~j��R��PӁ��5n�ŴM�X�6����e������l�{2*���D2�"Q�Uiz6�	�LH�s�g������1�f��tUd��CO�$H�]�rE� .��Mi���R"�w��������*zj]�6�"Lg�/,w�.1<7Yz��b"�����O3�����:�~�	D��e��7><<!։kh`�BJ�׸"қ0�D/���~c��g���6<��3��<����V��_す%b$�N����K���}�9�2�ŊP����Vڤ��H�D<�p�!=�N�<���
�S�l�ź�N����R~�x3+O�Ū�j�~��3e���П�� `,RN��`Wd�	!���|F���r럧H����&��4�0��y�+�:&��[dQ��>%[�3�R�@{g���y�-��-BLKA����JfS%�T�������9ps�=7<�f`����:Sf5��3?�
L(dš�-� rn5s�`�P4��Ͷ�W�VQ�$���⛛�� -(�]�0���H��p2�̦��/��9�t���S��k3��>�5Aw)�փ��Y����SG��X�� �YNл�7.��?��!�n�[��*����&�J�pm2�ꃻ�n׼���n�ͭS��_��E"����s�i�2����@�[� ̽�ؕ����U���#�w��Z����b��"��|ۦ�­Z�a^g���fE�~o-�-�9�"��Ǉ<X�4)�.ӵu|�<��.�oʅ�t����E� ��I���
��F|�P!�x`�5�Mbָ#�7���I�eَbu�H��yr#��$���� �jU�)mA!�0�ob�%��#�;�� |u�B�4&i��'�&>
�0k��U��Uº9�!yE����k�҂�r���n��o�ΉA-����X�'�`D5�t-֜nb;�$����*:W׃�i�$�)�ʋh$�z��\�reW��,�9��}iv�]_UN��>T9����C��O��$�Ƀ�v���qZ��V>P-B#[4�P�Lo�}_��a%9
�ًj�C��������Ae�P���n�JUk��[�*�_�����+S<ӌ�e@>�*Pc}7���6>>d?@,��*�=W��$�)�
��L��:m�8�?��NDX; ����д8�u�گ��L�pM�P�����6�����_<N7%1C^W���uj⿪�j�������C�ڋ�&�����) ��/�^e5�K�x��E��ZG�.�b����� ��p%�q�������#�Z���;�Cf�}2Z�:ߘ���z�b^N��P�(	�ZGć�5�xlIT��L�������x�F����i�O�_8�JӁ��Bjt��{"YERjFL�z%;�H��6o��&�\��A�S���ҾmJ[�Kn\B#@�p�h flE?��hhӥX	#�u[��X�KIl�#��l���5(�vZ�hYk�����sGY\���"��]��5+ n���*��@�A��t�W��b(z'������os��I�1=O�wP�U�/aS��%�w��F���-C|��a��=���Y9WvƊ�w@��ơ.�һ��:/eí6��Hivz	I[̕b��u{�� `�86qW��^�H:�_�P�'A^�]����t�Ј����8�b�s��2�*��Yn⟝H��b_�o��n���w��M� *�y;���<�����⻄Hc�;)�w��s|����OQ�Q�%/���*+)~���j����!N?@7Qa�k����#��t�ǣ�+�B,�� ޽Ml�|b��p؀��8�?���+��-����}
�)<�K��uFF�;8(��]2)���u8)y����3s�g�ʙ�z�.٘�o�)ߥg:`D����X�����Y]vC�ܷ췡��5�߲_����1�;pV���_V]z9��K���~pi�]�kfF�
�xIT�����A����
�k��������Fqo�+���X�4DwϜ@��\*AY~�1�tg��hD��QGm��1�7���.M�2cّ/r�\���ޮm��2D�~?&�>T��G�����Te�_�l*?2>��NzT�E�udU�Gy�L��������!-�\���TI~�v��Y��Td̮(/!!\r�f���8r�'���?�������l�->��;*t�Fo�/.��~��Bȷ��-�M��A�՝� ;��f-�D9�\�'�U��bP�'C?�!�@��^���������m0�b0?�?�{t����e����ݠ(ݯճ����\�#�@Gp��j�RJ�鮼���a���Nc۸-3J��cw9@剁��ε��[ˈ�ڜv�csp�d��(��-��(IYG�V�p�W����c���SeO�,6t)о=��n~��Vp��[�w���ăa�1rʳ����i=B���
ef-mPJ'�o��{��/����Y8 {��$�=EMO����Ji�R��f
�j-��	�$(�o�/"`���*��3�~����d��t(6�S/�Z��n��%F���ֻ�v��(�4�*��\���%�vf�XX>}ffk�Y�I5`߲���2��%��x�e[��~��Ò��}Ԁ �^�I�]�_�Avc��(��-�����yB�Q*�~�����geؚEo��ƱV�����}�f����Z����Q���8*�qó�����	f1nKa�)x�'�a��ɪQa�`�����8��}�a Ĭf���b��tZ�'u��"w�RہC���)]�1���w�[)�Rб�_6�^h-�g� ��~s�uZ2v,����2�t����#�g�9lT#S�=�}�Z�A�A���t���������0dΈ��/��vAD�x�ϡ�c�9Ҁ2����n�����Cj��%��(!�}�(38[j��W�mQv�,����26g-�(gQ�MO�i��kk��N�+�c�h������/��]Kj�|�)�P!1PM�]�)>�#�����63����>����M�/�
�!!�{"`K�����j*S�ܐ/���~n�z(MϮ�6��9�]�w�)���a��{��J����+�	�~�H6h_�r�sH��g����Nm1݈��<0�Ռ�{��~d]{vʞɢ!�s���2�"��t��b��3�˓		]&�U"�t/�9Y.M�7b����`��O�������'�mDV/�ew�7G��<1􎉴�3ȫ�`'��DpRD����LB���Q��"�Ϥ�������Vd�%�J��bE���l�t��+�⃢�,�N�ϊ)��w�p�M��p@=8h9��C�Š�:���5z��4�W~�B�RǾ3��r�3����!���}���e��v� :��R�.V��^dwUf�ئ�EX��}c������#���70|��y=p;:�Ա���Q��>.�r\@g^hByD뺾ְK
��ʹS.%�T�'_���BC���o7���`�Ȳ�>So���\�S��d.�-6�n�q`���t<��`�eQ���T��K�-�"���Ւ�s���Yz��녈X�K����ݲ���49kܤ��f`5*�u�T��Y�u�����r�� ����0ݦ�vI�J)�n�x�φ���yx
&��Q�9�T2ֽ^�מ��֨n$�SS̀R��i�����i�޶� )�@�{ߏ��&`��;��֐O��ĸ/�`.Z� ˹��">H�Ε���Zt1�g[��f.&�o6��浘"��ڇ��04���^�\|t�Ý�eCoә�tD1G�.�� mZ�IH��
4�<|��!���!�T��b���7ԳI�Y���7Ԛb�#��$�����u�ӊ'���T60f����#;>�I��u�'�4��]���>�b]0405U�����1!�>�!9�k5����w��~ԟϲ�`�r�����X�'N���>��m
��O;Q#^䳳��׌�3�*O�)�Zxh����u#r�-��G����v�@�Uw-�>���'�U�4�7���!��R"_��z6	�     �  �    �*  76  �A  8M  �X  Bd  �o  /z  ��  ܍  ��    �  e�  ��  �  N�  ��  0�  w�  ��  4�  ��  �  \�  ��  ��  � � �  ! �' �. {7 H? �E �K R S  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع������?i	�}�,$Pt��-<�AZ�~!���q�`��T��qq
���&@�Wڱ�ȓW�D�˵��73I��Q�(V�@�ȓn`�x҉@*L<Vd���!i��X�ȓ�Z��c��&�%���d.2!�ȓA$��E�°Ȑ���{�f��ȓ;��a��:D#��B'��7V̄ȓc�l�ᇏ��a�(�q,H:Y�4���/�@�GN�X��c
�����'9�~g�w~�iK��\-X0�B��y���z��H[?ʨ�jSA��yrN�{�"�@�%�\���yR�&t�mk2dU�ATR�L�yR�*zA	�#)���G����yρ�#I �b�p���J� ��yR 1
(*|�`j!a��Ǌ
$�yrM�{ 4��lѿH,,��6EȾ��=��yR(ʄ �hTz'�P�L:!���	;�y"�  +�:�x��RB���ŝ��'�ў�O�lp���ޠ#P����w�F,�
�'�:)�Ƈ�#)X��mT<�ȕY
�'�(d�Ћ��~c�S�(?1$ �	�'��5B�(��J��T�7��A;��x����i���@̕��"���B��y"ˈ�yl.,[7b[��\\)s%�y�b�7U�Wn�1����� �yl=?~"��)��8I۱�B��y
� n�Y��P�n���� Mv-%H>�S��y��L$_r!Ӑ���mWpPh�aL��ybᝑ,+��J�G\�h�̉f��y��']�qY��.�2�JUDЃ�P�'M �a�jВ�F��7�˝Db9��'��j�
�[�t� $[�l��d"�'�0�DJ"M�n����ƣf����'\튦��:�B}V�	�+�@��'��t(4!�oL�c��.҆q
�'�Hpq�	�:��1�S�?P�|��'n�L0b��2�����L�!�'4(D�F,�|� ��`m8L��Ic�'��,��i�x�$�0D]5K���yr�'9��h�L'@�X(��`���>9��'ԛFD�5,�Mۆk�"%���E�S��y�ɞA��i��]�Evbeѱ���0<���	�bP�d��3g���K�$�&g�B�	}��+$	���٣�!\6?��'�ў�?��t��3Eθ��F�5"9J�	"D�P!� �tp�"��	X�J��A�>�	E؞��`��#ڲ$��숅nZ6��;\Ovc��Rv�+�.��Fn�l�u��5D��A��Q�H�T@�&�Z>��xȖ�>�PT���O��tX���6|�D2��ز'�
���'�t�%�4{޼��a&X�#~���}r!%LO.�r���ebE#M]:
)aDO����ֿxv.A�s�0>��)JdF_�<A1�H  j@��.x��I�(�e�Ij��ɸO��6qq.���r�ab�E�?�!�\?��p!�Ⱥ^���0W��<�!�dT�r.�����5�D��j��OE!�DE=l�J�nZ�7��D���B�z;�'qў�>e�Ԭ���]QeL�6�,�h�a;<O�Io@�W��$8L���iZ%[+j���C}�=(�f��(Vz�oͶl��<Y��9�ŞA~"��e��$�T[�2!���T�����l�6i�G����Y�=��6��ē(�z�%���3S�,=3�͆ȓ-��0 l�Rd�:�o(,O"`n�|(<�c�s4�`����&v�tJ���d�<���H3�,A��O�e��P#�`�<�"���thEʂ���P�T�16��R�<��hM�2ؚPP�$�E�i�L�<yb%[�LB$��F��:��<�\H�<�0ի;�⁚�%�|��1�sf�_�<�f�D��A�F�.S�͐�h�s�<��*�U
�����%haT�!	�m�<��ͽ'�X #0���Y3��Y_�<!S��Ge��:�"9O�
��Hc�<�4^2g{lu��l�5Ǒ�S\�<YfK��\(Pf�U `��LA<y��HN`���,�mBAQ3n�$2'�|�ȓZ1 ���zݤ|K4 �m�r=��	h�'��|�N�z9��&��00���	�'��i�k�/6���R�� \E�E�H��n�y���O܌�m�2=0��D�gt�Y�'�T�b��V"��&nDP��(��'�	*Bl��^��CV\$H�����'�|��'J�Aq��@V��i��m4D�[��GL�ijs�5v��ܐ�.D�����`��L�F�,x<�($o6D���V&�q���JT!�,u@֮3D��_Md-� $�2D4D�Ë��yRN��:=ydd������N2�y
� i:�LX(S��ٰ-�$=�$\�t"O:Er�S/M��BD�͟M�B���"O0M�e�<4c��S��p��$"O�m��� �}f@��a��j���"O�!�Ł:����JY3/H<�K�"O6ԫ�M�f��y���F;z%H��C"Ox����a��⤌X�w���"O�d�rkA%��!مM�,��x�"OT��C�g�����Fّ�"O��b�#Eyf��,ڗT[y b"O��fY L&�|P�aP$VE�%�Q"O8��t
��l<�9AF!X�k�H0�"O�`�T6zs�t�o�b��P"Oz���쒁kݠ�3�΍P����e"O�(1�3F��!S�.�t�Ĉ��"O��3��1UR*��qm�)��h@�"O������iKVl���'��7"O��Y�J��Qi8P�C9��"O�����Z�q�Qi޺]���%"O�)�ϗ�s��vE͊;F|��q*O#�+�)��-+��?r�||`�'D �F�ɴ �H�i��,yv���'Y�*0M���cf�i|����'�<�+�lR� ����3n�$q�(Q�'b�Ӆl�D�	v.X��8%��'&^�K����M�"ʳ	����'l��P� �S��@M�3�����'�ک����'<|]@�/�!q }0
�'���3��Y�B��Q�1J�
!p�'P<�H���B�$ٺ�\�3��"�'���0�E�O�$�A�)ܺbN�	�'i)��nR+A�8ۓn�|� ���'88ઃ�)�TU��
_=y�XQ�'��͛a+
k�f삤�^?��)
�'H@l�&�35�Rݣ��T�*H�	�'�`�Ӷ��\����ҩR�E�� s�'.���rǔ
/���78�M��'�f�����8���3�6�<���'� 
FIaH<8�a��8��'����E�T����S(,$�	�'���
� �����I�Ť�X	�'5jy��oC�%� �Y0@^;?Ȉ"	�'d6d!瓇>��:�C�*� �(�'�����^��#��~���'[n�YƌݷkR���H+����'8��pG,	}j��B�"�P��'n���W���|��@P� ��'^j )�X�W0ٛA����Y�'$�,�ΈLܔ� �m�<c
�'2�!�ז�Lj�L��}
���'Z=X���(��MZ�b�vWX}��'���i'j�~C��0F�k&���'�h� 7jEz�&h8�I�0kC�Y8�'�J�X�J��%L0��G��<�y�'4��S���/b���x��� Vѡ
�'�fe;����8Sr����	Ʈ�9
�'������z3���VJ�i����	�'A�-��蓸g�2⥥L�b�"xr
�'�0�`i��%�4,+e�Q�\g�ܑ	�'߈�*�G%%��z�iUZ��c�'�(Y�vgS27 ��R���'@�|b5��o���r���M����'v�� �G3P3��s�K�E�����'\���tς�X��ap�[�;�|����� rA�f�Z�)�ڍZf 	��ɪ�"O��Q�.�p���� Ҵ�:�"OZ��a�?������I�\0�0"O�����9+v��.҇6�HԳ�"Ol��2�Y�QRh�J��w}
��a�'���'���'�"�'!��'��'����V��c�@#E��yN�AU�'$R�'���'hR�'���'br�'*d���'_�F����%?u�xT�'NR�'��'���'���'��'@�������'a�urJM=/�����'���'�r�'��' b�'�r�'�>��w(�����V�!*d��'���'eb�'���'���'�2�'�zU���ʐL��`����c��%Б�'���'(��'bb�'�R�'���'��K2ĕ�hA�	W���3r�'_�'&��'[r�'>��'���'#�|(w�E�8ND��1dڌn?�)a�' ��'w��'1��'|"�'��'`(
0hN\ep)�*�c�y�u�'���'�r�'1R�'���'���'^r=(��_��$JB��+^�t(��'B�'���'�r�'�"�'�R�'LZ�;Sm[���҇�#blU0�'��'#��'���'���'f��'�켙�B�����B�;�`���'�b�'5��'���'���'�r�'�EAw�Z�Q�\5 �#�1n��'Xr�'F��'���'t"|�\��O4��,Y�p׍L�<�a`���Ay��'�)�3?Qr�ik�J!o�'j����iڕ[��7"^0��d���?��<�t�j@Z %8�*�JR�����:�?���O�4�i�4��$j>���'���/!��%��ʉ7mގ����T��bc���	Sy�퓨h4�J�@�q�X�T��%bP��4{���<����z���wM@�I�枉Y'���3i������O���X}���3X�F1OڌxG��q�T����?~�P2q?O�	5�?I�g(��|b��
�K�ŬX��8���[�������;�����僃�!�	2rV���"9O0��	Eꋓ}C�%�?!�^���	韌���DM�4��ѣf�Qh�:ܸ���mo�	��\)�	^ڲc>]!��'۲���0#�f���@@ [G�Y�C$G:[���' �	��"~Γ�%�Z"_bZ�q���x�Rtz�y�s�4F>d�'y�6�8�i>)p` H g^.����VN tw���ȟ���<em�}~�6���� ӛ�d��,���P�#2骢I:�$�<ͧ�?q���?	���?ѶcͿ?T�8�mI<]abeȴ�+��d����#��I���&?�	�K��i�!\*R�xS�e�28,� �OR�n���M;6�x���R**S�	ф�J 07�Ïtd��0��-4���D s�:�jGeI3��f�	;��
�	7li����Cnkַq����	���I�(�i>Y�'��7MQ�m��D1%{�	�˱k�� `�ѸK��Đڦe�?a�W����ӟ,3޴K��5b�%I zlQ���Z�(EF��M�On5آc����4�w�N%��J�Zv�!R��"a���'��'6"�'���'j񟞡� ��'�|�*�Bξ/������O����Ox,oڊ~�������4��l7=�cd�5��D A���V�xBdb�Elz>QS@L���'�nLxR�����]Ƞ*N,��(T+h�\��I���'��i>1������x��~��=B�M�ls�����$�'��7(T����O��|r�X�,G^��Ȼ���J��'K��E���sӢ%�򧲅	.k�X��3ٌYz`$/�0����f�2^���t�� +đ|
'(2<y��� @l�hyVC�����'���'���T����4xȈ�뚂�L�b)�����դÀ�?a��h����d�e}��i�L(qv
B�hbui�JS�\|�M����Ҧa�4U��A��4����(%PyQ�����'L��$�O,Q^f��Jb��Ay��''��'$�'�BR>�0�ĩ8Ȗѣ�h T�ެhW@]��M�u/���?1��?!K~"��P���w8Q�`�JӖ����7x��j��pӌ�nڶ��S�' ��ݴ�yb�� W�*EЍ+���z�B��y�!��bM����,�'I�i>��	�T� �	�e$��AÂd޽�I������L�'�&7m@�>K
���O��D2)�h����!SW�<SՏ@�e���8�O(�o(�M�Ҝx�2v���P��0B�&-��x>ޜI!�B.3�1��q�6�b��0n%��	ťOJ���&l]�v}4��O���O��$4�'�?�v��-�X�I�)Ky�r�Q�?aұi�>,9U�'��rӌ���;�h Qh-D�䜡��>�扶�M���io�6���z�66?Qc�2q���V�PP����F��w ��3�iM>�/O�	�O*���O�d�O�dyr��B�+u�	�O� Sv��4��$��h�eX�<�����&?9��9p �8��U�(�b���-s�����O@�n��M�E�x����<hF�P���U�!�G�+X��$��7��$P���%�j���O��e�X��1��)�=��g�@r���?9���?���|�(Or!m��|�%�IU�6�ag�kb�%��w���)�M��b�>Y#�i�n6��1�𡛄#�k�N��:���G�FEoL~RN�7(`��i�'��� ��:p�]"u�mZ���>�HY@�3O����O:�$�O��d�OF�?p�B
�ҡӦ`E-sC򬲄����������޴'���'�?��i��'�퓲��:����U�H�gT>���+0�RѦ����|��m^��M{�O`#�^�Z-�V\7�� �U�;cԩ��iUO���|���?�]}��
Q/�.r���I�� �����?A-O�n�uvN!�'��T>qPS�ݐWr����J�5
HD�i>?y�V���	o�S�t�D(,�u��J��p]K@�["}�N\"�mV�$�TU���Xm"dG�A|D��+C���@�_ބ��	���Iݟ�)�SMy" b��I�AO�zu�����I���djG�y����O�To�V�r��	ʦuh�$Y�n~dtڄ�J+kܞ�3�S�MKƽi�H!(�i���2n$d$���O��'&D��ˑBF+m"�+���}�8����O����OZ���O*��|E��5<�q	�l�8"��j���1w���Q�."�'2���'�7=��d��ᑁv�A�K��6�М���O^�b>u�fV��}̓
�t�H$*�N���r�^("�z<�D�^�����O�jH>�,O�$�O���*$�F�E�E
�n���O����O&��<���i�Ⱬ�'r2�'�ܰ
�GA�4���B
#I���d�g}��'b*�$	f�
8 �W�}�"Y��mM�-�ɮb�d5`r�]�<^Bc>ip"�'[B!�ɯgg�*p"��{�l<�������I����I�<�I}�O�҉�6Q-�L��P/V�d�fe�w���kӒ���O����Ӧ��?�;%Ft��ɕ0�x�p�`�2H�vl��?��4S	��k�@y�����JJ�j<�ĢK�*��PѴ���l��0Ks!K!x��Q'�<�����'�2�'���'�j�D$��qЄ0 �dT���:�]�p�۴_L| ��?A�����?�Eيk����j��'$h,��e�"I�Iݟ���>��ŞL�)G��7�8�1/]�Q� Pk�Bd�'��i��aڟ��|�Q����(Kn��%+�I�y�E'�����������ny�Bt�\8ف%�O4A�uk��CX,9�d\�_�B\�Ug�Oj�mZe��_~��П�ɤ�M�6f��ea�a��4`���H`�R�ƕs�4��D�	}s��a����O��"C9��y��^)rl�`�H(�y��'8B�'��'2�I��-�<�q�m]x%{W*�",�R�$�O��$^��%�g@|>a�I�M�O>�c��Ƥ"�N�i �4�1#�.3�'"���Da��V0�֚�X�1D�(ZI�c�۠CP��B��������?�M�O~���:O���|����?���:x�@�g�H�C"6���#Aj�H��<Yr�,O09o��5�����p��t��)�"%!s)U� ��]pBcC��y��'�T��?��������'6́ᕬ%~����
��4�#�^B����
0��$䟪����b&ڒO�ef�Z�=�ĭ�!F�-,@XF��O�d�OB���O1���]雦��Y�ru�q�Z����;���26Z�L�U�'E��{�x��j�O4�D�o��A��6�F��$M4���ݦ�+ԇ^�)�'��H	ƀ��?���Jt�����9m��o��I�1OH��?	��?���?���򉌸[��8U��$\6�bd��=PHoڑ&����	ǟ0��[�Sǟ49����g�hZ\1{�ե�����%p��i��O���O���� 7J�&2O�\�4��b��Q��"Q�S[���$8O&���ɞ�?�e=�D�<�'�?i'V�V<90���`��)���R��?��?����٦	!��D��@�����0׫�]�9e��;+BZBG]O�X�	�Ms�i�O���t�iզDgO��N�S4��X���*F5��&擁-����X�5��b��JcH�]�dQ���������IٟtF��'>��ڥ̚),R�`xdkX:,a��X�v�|Ӥ���O������?�;)�n��*_�"��F�8IN�ϓ��VBaӴmڟ-v�l�}~���p	���S� �t���6�ґ�Zf�b�q��|�U������ݟ��	��h��_�W~����L";���S*\^y�h���u�<�����'�?�էʹ�*-p(��%/ܸf(�6n��۟,�?�|BViϻ�i)�I�8�����Z�D�sL���$
k�H`���C숒OB�u!��� Gӎ4�LM �M��H�6�j���?����?	��|�)O��oZ	&/x��I�U���`	f�,�B���9J��	��M����>Y���ڑ$��͚��OV�����	��P�t������B�߷"L�d��Q��ߙ��Z	m�1H� �(i:�x��|����ǟT�Iß@��͟����!0u$��Dg&%�|a��-�?��?!P�i\�a��OaB�l� �O����	q�r��=.Z�|��
�J����P���?� �Ŧ���?����z3���_�Mo<�+�JO C�O�%�L>/O���O �d�O�ɶ��&q�DS!�U>N�l�c`��O���<ѷ�i��R��'Rr�'��ӕD:MJ���1XE.|�`�Q��p�&��I��M���i�VO�S�װ!��N�_�6��p�
�R��a��ۿMR��u�5?ͧq(���S+��8�byIg`sz�*Tء&�۟$���\��՟b>��'<\7m�xx`�۳�	
��8��A�����"���O���]�)�?!�X���	���lx �}@Z=2��S�H0�'2*و��i(���77�i�W�O^<u��� ����G�}�yY3��x2$��7O~ʓ�?���?Y��?�����	�%7:d�l?-o�{F��@ʨ�m�r����I������?!�O���yG�:3��Prf<7n)!4���I��6m�Ҧ�ѩO��4���i�>e���J��8"{Vh��𞌒���gN��I�p~�
p�'��&�������'`�tYІB�Y���PB��&28BaX��'pb�'	R�� �4eS�,Q���?���0�l݃d��<,�5:�@;�p�C��/�>�F�i9\6��C�	�
�u��.0��XwAA$���^`�БBeN�q
2��|zr��O&����ivy���3�l!�ˊ
�*s��?����?A(O>U�I�EY���nCp�\����]eD�����M�$+E�?��[����4�VP����*PaL-���F#�l23;O��n�	�Msd�iT\ H��i���"+F���O�����B�5mb�iP`�&z.��L�n��gy�OfB�'�B�'��8��h�(;b������xv�ɱ�MÖe�?�?����?	L~���K��v��?�KP�ֽs��-� X���شdǛ�0��ɐ5,�6�8Q�� ��,�Zg0M��a 6�l���O�`B�� ��?91�'�D�<Y�gI|gPk'�U%����k���?a���?����?�'���䦍A�e�˟�6��p}��:ǁ:ٖ`��v�,��4��'����?,O���CN�j� �r��25Qg +;B6ml���	�&���a�OЪ-�'��t�w��,KF�O>��H�w�!��'`"�'�R�'��'V�8mpb�ʍs��	�bP���5�O����O��m�}�$p�'��6�9���|�.�JGK*C´����%H�1O����<Ɂl]�M��O��zF���1a6�bt�ՃHƸi�H���a0��D�ʓO���?���?���1�4I�b��-0�YQ��TN.�9��?)O��mڏ3�&��	ɟ���F����$��D�EC1"��t1cD����W^}b�'h�O�S6P�}��,=����
$`U�Q�:�"a/�]y�O���ɼ>1Ov���Inv�ѣN��l&��2�'�2�'�r�����'d]�Zܴ5�*����qK�����mKF�01&T�?�k��''�I��d�ON�d�V��Q�����5VX`r�%'�$�$�O�=@s�j���ԟX���=n���}y2��,5�f���V�y�����F=�y�[���	쟨��������O�\���OSMa|l�#!S���=�S�s��q�I�O(�d�O|��,�D��]�LI�7�T�J7��P��?ڲ�ɩߴ�����OA��%:��>OXl��F�l��Bc�ޜc ���>Oj��/���?i� "���<ͧ�?a���S�P��%��yU�8Y��M3�?A��?�����򦹻�͉��@�iYnZ/Y�X��ݞ2x$����0*�6��?IrT����٦�H<�WEđ'��(iƬ�#K��qd��l~���9G���sA�P���O����Ʌ�b�2'e�] �L	2���$M�{["�'��'}�S؟���&+\���wDV�5��Ȉ�ݟH3۴�2���?�7�i��O��?w8��C�=&��H�����OP�D��������'��0Ɨ�?�����i���\%�ڡB��9
��'��i>���ɟl�IП����bX8�@���1�n`�G��NՔ'�6 ������O@��5��4C���������`T[� ��Ke}��'C�&5��IW s�i��C�ݥ�
<"P����ޡUwPi�Ø��jC��B�B��v��xy�!�y�\���B��H	�8#��'1�'��O��	��M벫A��?��$�(*�2�1��`p򔹆���?���i2�O�p�'��6�^ڦ}i�4j�0|���O��j֝t�,\�Aą2�Ms�O��cr��z��t�w��s�M^?�՘aHK�Bh�E��'���'�b�'b�'��`�ьҹz�ʝ�cѹsW�!Pq`�O&�$�O�]o�ze�䟼�ݴ��V��1�0z�� j�4�� ��xR�'��O��\z�i��ɫD�r��6gƅD���Rn�)���0E)_�jt�dO�	Ny�O���'ժ?�V���T�$!(�`�R�'剐�M�@㓟�?���?a(��8����O
;�Oچ���'��<��O8�d3�)Z$F�A�jx@��]	Gz��4kB/Eb����k��M+O�	��?q7i%�DI"(9hѩ3�j#�I ţ�7�����O����O����<1��i��u��F ;؁�Ђ�<�*f��
j��'��7�=��	���צA`� �8 ������8f��*3c�MS'�iJZ�6�id��;�Ԛ`�O��'*�R�˕ʝ�}��pKPi�.lTvE����O0���O��d�O���|D��o���c$�4.����ժg��ʳ|ur�'���D�'}V7=�̡�nʡy��I�0C�ɩQ��O��b>M��-�צ�̓"�v�KA�L�1�r�b��3T�0�Ԣ$Y3��O@�xI>I+O\���O��r�`�5q�y����s���B�B�O����O:�D�<1��iX!Y��'4��'���y���&�n�J�o�69I �Y��d�@}��'kb/>�U&Y�"c DA��,a����:��I�4IB���F_�u5b>����'0��I�Jy~�Cb/�AG �g'��66:��	���	���P�O����ܴ�ҍ��Al�,��,՟ R�k���!$��O��$���?�;)� �P'��P��!U�:{@D��?	�VG�6b�! ћ���:b�8!�T�&� �li��ae�9��Ŏ�!��Qq��,���<ͧ�?���?	��?�_�ERT��U	Ôl�д��K����D^馵)g�Mן��	���&?��ɴT����U'��	�Rp8WCP�v�FdѭO���O��'�b>�j1Ɨ�l@0�
̂/>4�#Qg��RZ:8� 0?G�Ě+�����������6��`a�[�_r\��7,<���O����OR�4��˓-'���
4B)ˤǠ!{�j�&J:41��߶	�bdx�X�0��O���<!d��9A!5;�/ɧ`]D��"�Y�d;ش���+����'A͞���.�{���ٓ'Ѐ}q^t�JA�e���O(�d�O>���O���3�S�!�^�3��ħn��l>@�6�����P�I��Mc"���|��
8��|��ղ��Y���	�|di�j�G�X�O~�Dr��) ?�"6�4?I�j�qj�;!M�0}���c�Tv�vZ1�O��O>q)O���Ov���O`�thX�i!bd`�._�/��Z���O��D�<a`�iW��2��'f"�'G�S(2D��uA��E��HW'��_ 2�
���ş��?�O�������"A��0�y����_���H
�8��i>�r�''��'�8)5R'Ei� Q�J:9���kւߟt��ޟl���b>}�'*7M-�j�+��eu4���tt!iSo�O��������?�T\�h�	 0D~�13"�.߾#g���]^Ā����M�,���M��Oɓ���JJ?����JGpxW�ǰ����(j���'���'/b�'B2�'���Q�vy���Y����r򤜃u�|l��4kO�5����?����'�?!���y'��CG(xefև �n4BI���r�'ndO1�28i��e�:�	�e�$,�sC$z�Հ�)vK�P�	�9m0"��'�b�%������'�,�3k��(0�)uL]X%� �'���'��P���۴e�����?I�3�l	H��
}<�A�C-w��Ah�Bf�>I��iv�6-�e�Q��q�%NΗ�P	yFcݵu���-/��En��.�h��|u��O|�������rb�����$�����?a���?���h���Ľ;J +BC� $49��a.AX�����iq�D�(�I+�Mc��w�X�C�R�VA,�(�ʶL��r�'��'��6-ގ6��6�:?�GeQ,YJ�i�}�@D8���gֈ��Q��I�O>�(O���O4���O��D�O��s���F,3��Ļ [$�#��`yr�nӶ�(0	�O���O���
�dD�J@f�(CC�00�P��ա� R��'���'5O�I�O����+h3.X���,@����Њ��Nc��)&b�5\I��A�ƨ��'��D%���'�ĘK]�vpaV���,E��V#���?y��?1���?ͧ��DEݦ� r�O��"f��`���!� ��YM��@L�Ē�4��';���?9��Xƛ�;��K�%�/V�8�M�Wb@��ӹi��O&I@�̍�����@���ߝ鵋�{�������n�����q�t�	ğ@�	՟��I؟��j񥑠D����q �9��?���?9ųi�`h�O ��i�^�O�`�߼^�]��#d�6�xg/QJ�I��lz>����^ʦ��'�V�`6��d�^��|��	n*l�V��ן��2�|r\��S������K�)fHF�:�O�8d�U�fÚ�d�I~y��|�l���J�O���O�ʧo$-i��ywJ�ˇ5zC|5�'x���?���Rꉧ��4*޸M)6ɴy�dY���)8I#�M�e�M����2/Z�g��)6Y�F��2�T�t6(�	ʟ�������)�`y���
�mJ�^�8A�p�+W=: �&�SNР���O��nE�*��Iߟ�00��~��\��⃳�n���D������4�"�ش���ǿn[�Qx����S�m��@�K�8fv4 K!CQ
(���Hy��'��'q��'��P>U����:�¨Q�@�*k�
�K0KY6�M��A���s���?����
����4�>�x��=�d=;u/{s�$�C��O\�D�s}�����'��t����&5O��Sqi�H�TR�l�8^��=O !Zf�å�?���5���<�'�?٥�TN����&I�BZ쐰��R��?����?)����R�E�d ���I��P�J��G&�KvƝ��Лs)W�?`�	ȟ o���ē#�f`C)�����@�Wzl��'"ZE�q��?��䰈�����ذ`�'0��0���"SX���@�,fX� ��'���'��'"�>��	
1�z�n�F�y����4�	� �Ҍ�I=�M+HW�?I�Qq���4��}���X>�hH5Hʢk%�0�>O���O�$n����m�b~�%ѡF��?2�B�"o!��cS抆��AǑ|rV���Ɵ���՟��I˟D�e��	���ɡ���5bUAyp�f��.�O ��Ol����
9�D�ԨW�c� ����%v���'��'(O1��y����\X�I�ǌx$�QtMзNͲ��垟D2��Z�n���]b�ey/�h[#l.4�fM���02�'��'#�O*�I��M��'D��?	����%e�18F�M�6n��Vh���?if�i��O���'M�6m᦭��4�>��s#	�t�`{BV<3�P�Fߵ�M�Oʄ�B�%�2����w���� 
�J��x*ν?*�Ù'B�'���'�R�'��1Jb�-/�UJ�
(
cX-	���O��$�O�@n���ߟ 0�4��oz�����(:4)��HL�T;���Ж|��':��O���!�i<���7��� z�JD	$�|!	���O�*fh!�?ib�7�Ĳ<�'�?����?�Q���0ԛ�MY�lӘI	s�_ �?����զ�i�ɟD������OZN�9�gN��	-f��B�O� �'����?��D&B {��IuM�&�z�H׌ЏJR"��h�TҘM�����R�\c��|��'ƨ]�B�#\ �x5���k���'���'���4Q�P�ڴo�xH�)ub܊%��$���4���?��hC���DT}r�'�FX���n��Eƛ!�Ɖ��T�xK����' �1!A���?]X�<"ӧ�x�TS֞k@X�H�u�<�'z�'���'���'a��$%̆��G@�o�,M��'C?o+"}�۴%�~����?������?�Ӽ�y��؊v+���W`�8F�T	��׃F8��'4O1���Je�`�v�	!A��-|�J�䎣T��E��,}����G�L�IT�	oy�O�r�3Q�BX���\�6D�Y�(Tt���'R�'��	��M���?)���?���e[e�����n`�"ש�6��'n��?��B�U	l��И��]�8=�p��h���߻{q�XۤW��$?���'R�����-؞mr���;V����PUUd�	����Iꟸ�����1A!�$
�X�p���NXe�$Hݦ��Uh�ӟ��I��M[��w!�"��^�}��ۊ'�F\(�'}rX�{�GK���'ٰuxr,��?"�C	D�̽�t��.1�h	��ͫ"t�'�Iݟl�	�����(��:a�T��D`�8<��p��
y|�̖'��6��K�R�D�O��d=�	�O\ �AŖ�1M*�1eR�Tac��F}Rl�em����Ş]�d�H�I
Z�M;�ͦ�<�C�cC���X�'>X���ǟH���|�S�(�6�,Hl�h�ɝ�[}����������,�	����hyr(c�ȁ�d��O�����V�F&F��N��Vo��,�OnHn�j��^����� �'�Bd�7j٤]Ѡ����C�}��e���Z>�֐��
#�W���diWf�S���Cw�ԥ~((���^h|�:�j�X�Iɟ��I៤�I�d���L�JAۂGM�3���G�Ő�?���?93�iHl��O�mm�ʒO�}srDI"@��5��� d�Hp	ՂYw�	ȟ��i>��	Ѧ��'Ǿy8rH˦,��A���V4[r8��K���x�I%h��'��i>i��ӟH�	#>�,8�͗�U�p�[c/Ml>p��ßĖ'	�7�_ a���O��D�|ʦ�_��Q:�BN5q#�\�P�VB~�
�>����?9�xʟ��B.��J6��k�Ǐ�KI�� ��>�rpR���8!��i>����'M��%�(��a�q)BH8��L=~K�tÔ���l�	ϟ ���b>i�'��6M[�Fj(�
E��'lK4x�hF������O����Ǧ��?q�P��nZ /�Y����\�pT*��?*�H�4oқ���+85����t�f��]���~Ҁ��(z6�,AA�U�j���g��<�/O����Op���O�d�O �'#`�tAB��+U��䳠�k�tdS �i�"�p�Z�p��S�şt9����U+�Bg���g<a*��_�9��V�l�0�%�b>Q�&�ڦ��2�H�
�]G�9�Wf��<�vx�f�0Ed�Or	�K>-O�	�O:	b$�ڋ��5i�/_�Uوв���O��D�O��$�<!��i�~L�g�'b�'q"L�hʀ"h ��7��hHjb�Dd}��'��E/��#�*��I� =�4�K<<i�I8A*��D@0x}�c>I��'x���I4}b@��妜�]k��˚�/3���Iʟ\��ڟ��	`�O�R�9/6�H��Y+o��k��H�W��fu�����M�O���˦��?ͻ<�%0�ŕ�@�L �$d3< >��?	��L@�O̩#ڛ���h���t(�6���@�%ѝh�>󥊗�^aU$������'T��'���'�J��A�p3�
	�7$0��a
98���9�M�s�J6�?A���?��tӼF~��ۣ����jxh�i
%-���f�f�$E%�b>��������a�-Y"T�@��cH�h0Dݳ��<?!g�X�n��޹����dH�!xV��уA���X��
=^;��$�O\���O��4�:�1�VON9@ҭ[���A��F��w.fh����)�� |�����O��l�.�M���i�F��2��	T�<`JtF��z�� *'�*v�摟�3��8Pf�������-1�
<"�����R,��p�G2O2��Oj�d�O��$�O��?-��⋀_<* ���4��#�K��Iß��ڴ;­�'�?a4�in�'r�x����}�L�ٴ��i�����+�d����۴�b�b���Mk�'zrGK!| H��9M��YZ�LX9.��a��@埴�T�|�Q�����8��ɟlA�U�s�6X˶�Ѿ�4�D�Ɵ��	dyhzӬD��j�O(��O�˧)qH��2���I6���4gY�MK���'J꓍?��ʟ�PRW��i�����K˛Eo
�Z�O	%nUJ�a�m��^$��|Z�'�Op1�J>�aP�t�����=]�����?Q���?����?�|�,O��l�Lm9â�g���kAF0rq�@CP�����MÊ���>�ձi��p	�lRz��q���,	"~ER�.mӎEnZ��Yni~",�:c���Sn��V�j|R��e%��J�eɸ:�<!���?A��?1���?�+���	� �X/|i�2�ؠ!~�	��ӦA���E����8�r"��y��<��(@�2e�X��3�$K;6͂���M<ͧ���'#�H�Q�4�y
� ��+#+� Br��+�MY�=O�� ��?��>���<�'�?�"G�x��܉c���qs�=�
[��?!���?��������f����	ƟTy3M�#���f@R�9h��W�B^���Mt�iiLO@ ;�?Ao�KT]3ƭ"���$#&�^�"��$Y�)�#�B�Iȟ��R��E��*R�<�%�n�����㟤��Ο�G�D�'~(����s�P����:���PQ�'�6큲F�x��O�nZE�Ӽ�3�P%�%�Y�Z`̝{�, ��v�6�Mt�i��6�5̾7m$?QצJ����Q%P"�ZӤ�5Qƍ+�B��b�M>9(O��O���O����O&c��ݺNx{��3�ܫ"N�<�g�iHr���'OB�'��ONR$^5��0��D�t��C����?��v҉��OUN\�
ȘN6I1�l%f-1{t-��h~��Y�O\ ��hX5u�
��0%O�2v�*�+��x�P�+�	O�|X3%�v5�ت���/	��p��Ȍ#z1�"��d��2��<6�4cA08��t��k��cj ��܋-/.Tt��lh>) ��קj��=�N�-Pj�1Vg�<���8+�L葆��G�	r���Z�S�JW�!�p1HI?��i ����R�-Iנ ������JπxHV�։NyB�1�ND%!�(��7���n�F�T�)���(���7%��!1r�o��&U��y��@�2+ܤQ�2)9����U�bz8�rQ
�n, ��/ʇ�MkS��;z���)�$�B{pF[�,��'2�|BV�t���>q����r�HH�6�X���8���N}"�'���'�	�(���J|���];���sdTY�v�#"B65�f�'V�'��,B,�O61�1nJ	]�����U�jZ����i ��'0剽}��lO|����0C`Y��X�|�xԠc�O f�'��8j,�"<�O]<e���\�_��E���1^kF�8�4��Ğ>_6�n�����Ol�io~r�#VT�|�P�K-t8����@��Mk,O~�+f�)�ӳxÐ��ǉ�
F=B1�pm� sJR6mŒ)���lZȟX��ӟ���#�ē�?Y�,Dq��j��Au�(ԃ��G^��Ӟ�O>��	�8 �3,(q�!%2�2�+޴�?	��?At�&ƱO�ġ��(a�4�M��̅}�(��5�	�`�Xb�P��ʟ��I�9�8k��܆+ ��@/�;\R��jݴ�?��"2�'���'D�^��+0Q�-�Pk�]��Yj��z�,�I딈�<q���?����$�@� �ӱP��Ÿ*D�0$�Z�nа'���I՟�'���'���b�M�r�\�ـ��3b� �3"��Ș'�b�'�rX���2�2�����Ll�۷��O>8�"�"���O8��5�$�<�V�E}"��(7J ����->~�;�����OJ���O�ʓPS�Y��$�M�*r��N����ȃ�>��6m�O��O
˓;���>�e�أU��uI�Ј�$l�ۦ��	؟��'��;ӂ1���Or���#z�]����!:r�4@�d
!���&�T��$ʑ�*�l[�ah�c�'�6��<���rЛ��~��j1��l���u���O.-���j�@B�I�%��{t �8f8 �6[%ǖ6ОC�����O,���O����ON�D�|
���6���J�5~���3C��;/m"<�|j���``�������Ɇk���a�iM��'�b+�w'�N�t�'7���g��:�`��D��?~8`�Gx2�8���O��$�O��BW!�f>F���"���F�J�q���\��I�@���D�d$�`��{S��*]*��F(��
%�e&����c/?����?)��?��O�T�3�]u���5�ϔ8��d�:����O��$�OH�O������KI3Dz�%� Ă�.]d�	��nӆԒq����I��|��^yR�� 7���)%�0��biǠ�\� ��,�C�i���ڟ�$�\��ڟ�H��ܟ8SG֣c@��"�i�9-��d!��b������֟��'�@��%-�~z�Gǐ���˧�$�p��5^N����i|��|��'}��<qO�$�D�ÐPOx��@Dь&��9�t�i�B�'�	�A���9��&���OH��9>��KΈl2l�0/�4���$�`�	�0�b�=��TC� @��K�EV+,��k�JW3�M,O�ȡ�m�����៨�I�?�k�Ok	�U%�|���ML�`@�!<����'��!N7�O^�>Y�4j'�|��$�4D��p2F	m�V� �AϦE�	�T���?�O*�I�ЕEA0,��<�U��!��b�i��HK��$7�ן<��d���(�����W	�ZlD��M[��?Q���r���Z���'���O$�����y_�����V�#5�x���D�,y�x�O���O����'r~+�
�w�8EkUm��r���C�i4r��he�듶���O��Ok�'7�M!S���|hah�0'Z�	O��<$�x�	ɟT�	Kyb�95H$��r!ЍD��aXw	��Z��pP(�>�/ON�d4���OL��:5�<(s N#L{ǡْ����� ,���O����O�ʓzo≲�2��pQ$��'��D�E��)<��
Q�i+�	ǟ�%�8�Iǟ�B��I?A ��BӀr���|~)�h^{}�'��'��	S��x������~f.HI���3]��x�^#z�m���&������g/�S�d���� 3V&�k���N n�m��P�IBy��ld�꧆?9���bu� �dqS�Q��l�c���8��U��I���ɸ�
����<�6����+L�"��ZB�X��8AW&֩�Mc.OU�R����M�	��	�?1A�Ok�I!t�x%���{pI�Rk��?:���'��cƤ[�O��>S����Y+r@+�)]2"  ��e�i�t5�%˒Φ=�Iȟ����?��I<ͧ?�!��K���	{QĔ�d���ivASc�'��'���O(�s���ɞ_�d�3A��>�୳����+� 4��4�?����?QTJP�������'&��ߣh(�X#w��, ���q�+����'��ɂG�.٨���$�Ob���O��@%]�}�~����#a0��!��������3"&�4`L<ͧ�?qH>��U�(-���YI�,⅊Dmr���'N�c��'��I�`���ė'$�	B����=�E$�2������E ܖOh���O��Oj��@��@^�a�n�@D�G���V�K��?AO>I������O��@�?����pT̘xRᆅ���H�bs�*�$�O�� �I՟Bs�52Ԏ7�=�dpFM
�r-(-iA��o#������Ɵ|�'pLXH��%�òD+Xx)C���]�8l�a��^�tl۟<%�L�'_Tj'�'N�q��\��DK���<Tb�-/ܽl�ݟ��IZy�۩Q��������k�G'\M�1��v��1	@�TE��T���	͟�@�@�؟x$?��s�=KǤ�����Rb��_	`58�o�>��;�:�B��?���?1�������qU�S2���S���s����U�i���'�-��!ȃ����O���$JL�r�eL"�Q��4Dg̍���i���'���O<PO�)G%9��i`���^�H�g�Ā4��lZ����I�������E�tR>�J�F!!�o�;a�2�E�A
H��l�����I��ҭVCyʟ~�'��@���K�t�`N\
bN���vG3�	�+1.@j����'����S�2�˴���q��OE<(��'i��z"^��@��P⟜2�@�a��'N��������)���ZR_l�#����������zy�H��^�(hbZ3ʊ9c�)�����"��O��'�$�<�Pb�?8Z	FLP�e3��q�爿LF|����䓙?	(O�����Ӗ��HG*/Q�*\@��U><6�<	�R�'��(
�f�"޴y�N��w���`�Z4�Ww��,�'}r�'��U�0V([1��'/T���J^8����G�V�XX|���i2�|W� Ґ#X��h�����#�T٨ieo٭;�|�ķiR��'��G�~t
J|�������}kFo��r���a�ñBt�%���'R
b��'��O�������5/e���m
Y|��ʯO6�d�HR��$�Of��O�	�<�;Q��XX�&�c�I
ጆ�".l�П �I$c�-K�+:�)��P�)���=o�. Pg�Z��7 
d�|lZ���I�� ��&��$�<I�%Q2
� ��jƱWeL�� ��~�V��?�y��'��E���?9Aj�'{��#w$��=X��x�gB'k	���'���'����B�>!/O������SĆ�~�Y�g��.P��-��|Ӏ�d�<a�$��<�O���']B�F9�z-���՝��\���R�Plx6��Od�� R}rV�L��Zyb��5F��B�t�[����*0�!2�)�,����<fJ�D�Ob���O����O�>�|%ѥ˝�A��1%S�)�|�թ!���LyR�'Q�̟H�	��\Y  ��p� ��T�E�g�Ә�>�I@y��'0��' �I�f�8-��Oj��:��A
����ώ�w�|u8�4���O�˓�?����?�rƊ�<�u*U-4Y��C(J	Ԁ��N�=���'?@��r�'��W���`���i�Ok��"*���7!Q4w�&����A�W�F�'��ǟ��IɟȺqes�\�'ڪ���%���i��3o~E�3� d��'[剐ђ�R������O�iI�5J�ScJKhLJ9��
�C�~!�'[B�')�=�y�U>�	o�t�T��~��H˖un���Y����'(��z��g�����O|���N�ԧugO��2���r��Pa��CL��}��ğtb&`j��%�,�}B6�"@��he[seOȦY�S0�M���?����1P���'��C�
^�:,bLB/ZB�
2�cӞ�˶?O���<����'N�8J�i�i�|��	2�@�
��6-�O2���O�4�Aa_}Y���	J?aa��t�X�dP��u�D�C妥��Py�#��yʟt���O����Q8qI�,[�#$9x���!l��mZ�DRe�����$�<������OkI�Jhx��b��Y�����F�|%�I� �|�	֟����<�	��d�'�����;C2))��/N���X�m�)WN���d�O���?���?92�� ���`�/�<X�*��3�X���$�O����Ov�4�P�x�:�,� Ac3-��!�Gϊ-6�Je�v�i,�����'-��'�B� :�y��ƨk��Y@��1����.��3�6-�OZ���ON�D�<�%�R�:���Ο�ث>_��l��4�JU��Ҕ�i>"]�P�����ɖHO��I�d��i��H�"�
,!D�! � �l(mӟ���Hyr�� {��맕?���r#�R8ǰ�����0Ar�0Є)Z8��I����t8�*e�\&���'Iݞ�[�.W�<���f�A�$Z�m�sy҆ʤK��6��O���OJ�ID]}Zw1��p�B�u��-T�蘉���צ�	şd��fz�<����$�S�L���'��F�&�0���-=�6�ˮ_R	l��T�	ϟT�S�����<��� ����뉸Pj�ɸFMOYV��Ȧ�i�"���'�[�|��t��p���J�<�,�����2�x\	�i-�'T��Z+�Z듼��O���#w�*���o�31nHԀԅPPF7�5�����?]��Ꟑ�I�
�,	�b�T?N�H��(R?&q�ܴ�?Q�ɍ	a��	Uy��'��I՟��U%�Q�����mА��S��{^b��?a��?	���9O��SwW�a���k�\�� �T�ʸ�'��ٟؕ'���'g�BC�q1иi�(W�) �=�RHL����'�"�'���'�s�L;E ����jC ���"0{�D%��/��M�(OB�D�<���?��nA�@`P�˚�A�n$RAę�5i�q���iR� 2;|�'�	���;��>�$A�[�����MX�s��uk0��`���n�ƟD�']��'�mع�y��'I��ä�^�r���w�ZpZ�E�H��F�'W�^� "�DR�����OT���b�۲��1�v`cF4vꉠ�k_}��'�B�'^X��'<�X����l�~��q����V�<^��n�OyB�Q#��7-�Ol���OX�I|}Zw[@�:ƣ�O�9 ��,���۴�?y�C��!̓�?)�ha��i��Tg�%P���F �bY�h2�"�M3t�Ҽ=ݛ6�'���'��4Ȼ>�,O^���ƷC�6�'I0$|��� �֦M�A
z�8�	tyr�I�O2|�䔊m6����J�4L,|�HV�H�����ڟX��+!��O<����?y�'B1`c� c���h�#�/���Iݴ��	�J�������'D"�'dڗJ��9+� SWC�<*vH� ��q�Z�d�U�'����֟p'��)\B@����V�U��u��dD�+f��N�������OB���O����q��G���H�j���e�,i�B�Pb~�Od��:�D�Of�k�*U#'H�����'h��j����P��<y���?a���DS�s���̧l�t���.d�>|JRd�+2���'2��'S�'3��'�����O���ݟ=�,,��9s0|  P������I@y��%{d�������&"^8ԣĎ�#` 8��@	����ICy�'KB�'�4���'�
���p�bէOU�NWG��l��L��Uy����tF�|�d�����><ɲ�L�
s�l��I�?�'b�' N���'\�'<�	 �&�(�6�C�Һ�3!�ӵ��3���M����mZ�����O��)�\~b��.C�R�3�ӸU ��33K��M����?�Bb���?O>���\�$�ey��_
�4�YS��MvI {L��'kR�'����)���$F�`�� �p⥐�+�a��4d2�Γ�䓠�OB!�3>�����V�P�Ȥ1�F�A��7-�O6��O"0I!(	|�I���	V?yQ�2pM��;1aLiI@����u�VT�@�L>)��?���~���/Y8z`̻B%U6(,��G�i�Ty��Ox���O|�Ok�݁W|
�Y���lB��� 	.E�	�o��`��Iy��'{�'&��-Q_��Bf�123�(�mi�M;x�>y��䓘?q���͐��KX:�{Rn�Q�*}ѵ��<�,OH���O���<�bj�)��鎈o���	VdZ���9��Ƙdԉ'T�|�'U�낱�y�ބ746ɠ��T*r� X&��+x��?����?1(O��V�^�S�Mz,���A/Kޜe�3n�`���b�4�hO˓�?9I�BW�0	���#E͡w����cu����O�ʓy8إk����'K�\c�<y�
װKCz,�u�^�RB��X�}U����|�Ӻ�f	��-�q�'S.n�͈�T���	�@Z�ɜ����	�,�	�?�5�o�	��)���Z�ܜ��N���M{����	��jya�a�=i��i��Ȩ+���)ղi�dq�7Mm�l���OH����6��'V���"09�@L't�ఒd H1�)�ش�?����3�d�O��	��~)�ѮV&U
 �Di��5�����I	�*��	���O�O2\�*ɛ
��嚂�mT����z�'B����$�O
�D�+D�N��W�v�B0�[ 5Txo����ҫ�?��D�<�����d�OklX6f��JG�+g��ٓO�?w��x6��?A���?I����DOe���۰ꕍ-��I�L�4.YJdVz}�_����hy��'�r�'���
���2@z*�����]�6m�s��y��'(��'�'x�I7F���Z�O�Lt!�A�Љ)B O�/��i�4��d�O4ʓ�?Q��?�a#x��dݹ"�� �T%�
"fv������$�O���Oz�0�@vT?����"D6�r���D��.�N�$iٴ�?Y)O���O���̓Y%1��6$ѕ-�"51a���R�����M��?i/O ��V�d�'���OG�Pr3j"I88�( �:�9�J�>����?��J�0��?����r�s����JEI��~��0��-��@!�4���\1d�o�Ɵ��	�����<����$y�%��6�٧��{��dBR�i.b�'s�z�'A�I�dx��}�Â�2��t���ޅ*���@�ӦhG0�M����?�����Y�T�'.�MS�d�Q��-���YC�l�^��Q;O��$�<I����'�����5p�d2��K�[�*�!jӤ��O��ĕ�J��I�'p�����2�$�a�N���l٠/C"#�UnZE�|h��)b���?a��	|N8�U�ϕo�0��c��35���� �i�r��6|��꓊���O"��?�q�? �H{��h��S�"M�:3�i#cW��*��u���Iٟ�������]yrd_+I���%I�P�0XhReJ�	����E�>a-O���<i��?���/� y�͒��X)e��=e-�{�C��<y)O����O �ĥ<�A�#;�I��d$���M!)�xH ���B,�VR����}yB�'�"�'���q�O��j��):�vᰁ	��X�e)DW�4��؟��	ay�%���6�'�?a�H5x�TU�f	M����i���;|g��'��	���	�L��p��'o�db$���K?~H`e���T�Щ��d��9�'�	>7��z��>�D�O �I3o�� ��;�`TˀD{�U�'"�'YN���y2�|�ݟ��VkQ;"����t�	^
U���i�R�'���b��'�r�'@�O��i�%(Wg�K.���?$�H�c�Lf�����O���a�IJܧe�IӦ]�cf�$���׊^����	�S&&M�EaC� =�����R��!am�!���1���WS!�dY�K���;��ÿ}k@u���۸k���T��{��V,.T�]'���_��{ �ƱaS0�B�ܲ��	Y�.�%5������>[PP[��]6BQ�2L�DsҸŀ�c&���U&�/�T�u��0G+,���<Vyʭr� S�7�asG�^�X��t���{���P�L�Hw���O>���O��?�����$��&�̜@G�)mz��G�M�0���)q��C2��1�[�Mc�yr��l5#��ޠ>_��҈��]h2`\�Uz�9�Ì��yB \;%%�����9��Xu*�C�� i��?9��$(�ɻg֙�G�ʝt~	��EY,�$B�'sXR�"L�*^���;0�N���';*6��O~˓Y�<t�QY?-��< ̖5�%L�a��`{S�ѳrc��I��T��FO�|���|jT����JP�.B0�:�4�	�!����<���ܝZ�~���00��ĂSB�>c?���րI��H`��,�Ѣ��2:�Έp?O��D�'�Q�\v�	�#��<cpJ_�Sݸġp# �w��Ū 90z��wk��2��I��>��hO��Gצc��5~�I��,9:���3�V�8�'R�I9k|����Ofʧ-�|ق�-�>	��V�H@�0���9R�S���?�Ek	9;L�Y�@����	k���I�|��)D$B1TH���!&0R�94�P��A(x%�ӂ�8������O��*��2����\��\Hv$��BenQs3�S"x�L��@���pF���'S���'�X�%��!�2�Z
|C4�k�'(��Y�/�;x0�y��V�li�13&�i>���䑫L f�Q�È�V@jYS���l�̟��	���S�ҙd@���ӟT�I���]V�x�p��83�Z��fC"0`h�Q�+N 6�ɣ,��=p@	"�3��V0o�글Ԍ@%"�i	f���Rt�������D�+I�,���L>y���u5���*�	D.�q �צ�?��OR4ړ����I�60
�����d����ZWvB�	a
�<Jw
�~����&���g���S��' ���w$�<�.�PS��̐C��~d0P�'�'�Bqݹ�I�̧g?"�q�-�+o���R��׀q7��#Ӂ�B<IV��<��m��l�2��)�@�?u����?��A�υ/?�J4�5斬l�*��ڟ���	�I�>U2Qe��RGd�@�N˶TY*C�	�W�Zӥ:Q�N���ɼ`��b���4���Xh�Q?A�I�B���!!�i���Ԉl��	ߟ��UE�ҟ����|R�Uj;T���k��[��D^�h�!���0��F�k�x�a��C���p7L�(ߌ�	�^�l�:5ě�I����j�3$���o��'��% ���f#L1.譻�d�-+B�b���}�F�P&��N1�er`�]�d�B�I2�M5�_�
�H�W�\*= XM� C���?�*O�hƫB̦��	Ο�OH�q���'��ɂ��2�`ر�R�adx=Cw�',���'��u D�ٳB����5O�SY�$M��eBփ���>�GF����ɻ@$� ��A�4m���]��M㄂J&5B&�'Iz-�����g����D,�����O>�C�')���ę��	�w��=;�j�������'���'�.5��b�Y���!.e��i>����Ό2��$�A���HAz��Z�h���lZٟ@��쟤@`J�	�����̟��IΟ杏/���d �B&dB<����<QPi�&/���iU��ˡ��'jڡ)����qOT�X��C�0<iDėI�8P@n{�}���L��?a�O8�����?)���?��d�l�X���荭;��(&����x,S�	�|�0�Yp"TaGJ���IB���i�<I3	�c���釪R3Td��S�$$��2�I �?!��?��c���O�Dn>)�`Z���ų��˄xPt�e��9�~%�"��%�v����nx�h�ȎL�Z���@�;x��9Pe�U�-�2�wL�7G�=⤮QZx��ẅ�'*��h�L�Mu���ā$�����O���,��T�g�? "]�ԀP�"�P���EK�<ބ��"O6�ۃ�]��x0�� s�,���@ߦ��	sy�f��6��Or����Ⱦ�{Р��o0��1D+J�6����O��I��O��D�O��:#�T�c`8 '=O��O&��$�#�����Wi�k�x���Z��5�=v�ܬ���.Z��	�b̌�l@����f�	��к�bg�������!޴�?���ǘ!��]�`�K{0](�Hٝ���O���Sy�?���(�h�<��OCf�QW�,��R۴R��]�I/e�Ȕ�BKO6V^�!�i��O
�$(ړ4�x�/*�� �*ɍ =��S�R(��lJ��f\ �/S���ʓ }���C�A`V��Vb�:$B�I80�����C
�\}�C3A"+�C��$$�:� �MKAO	���( άC�ɡ[�������0��kB�W�WvC�	�vJz�Җ��.��X�,Xc�C�	�S`!ɕg�
(�Q��@R;�*C�	�`'� �'yѠ���Q��B�BW�@�Dn�z�hX�A@�>��B�IZJq����}@�R����ĚB�	�A ��r��0�p�bt���}�tB�	�8aa33���
�`�c���E�dB��3n�X���ǁi�X`q��4.��B�	�Fg�	�1�?#\`-(E�;phB�I"�h��?��:6�<Q�8B�!h�\�8�]�QyWf��\w�C�	>:��}(� !�����$f��C�	2����,,vЪ�h��5��C�  o�1`S!�GL�؀7[8C�I4[ւe:d#ުgΐ�D��&� C�ɨ]���;!��9=��Ӥl�̴C�	����J��P۸-�2��&h�C�	=WGJ�y���98Nx�Z��N�)?NB�J��!Kpm��A�=�hB�I�(���d�ܪ�OR1p�XB�I&A��ɉ�.��$p��S�i�2B䉑,������O��90?=R�B�ɭ2~:��5a��p��)��nާI ��>)篓�6���{k�|���α�HUwɃ!��5�j�P�"O�a��Ė��͛n� �8O\�bEdYk_���"�X*�`
��)	���P��D��B�҄�&~o!���C��\�U���p4r�A*�<L�9 cߥ��I
C+WQ$B�ǜ?#<���_7x1�š&!�2O�8���n���h��~��k��
�rq��*q�ªqx�X�Hԙv��+�	�R��|��t���k�jG�9L\��`�&A2pP�������I�t���2�V�
�(��+���8�<	rϗ;5dv�٢b�g���W"OXY��R�6	!�V����ē!�N`b�d�T�j�E@ё�H=&�V�&)C���H�t`��!j�*�$B���>h[az2kv�	�`��y��M��E�AU�7���ٔ�ƥ.ހ|Ґ�OP�z#�yh]�N?㟐�A/�t���D5�sީ�1O1��߫�X���0�*������?s^�#f*��?�7MI�TTU2��6�H��
�8k�%�#�`k�mB�P����'>" �N|*��p|˓i;H����	9B�T����M��ɳj���@)O4e���C�0�<MR�
�9*��bHR,S(TI���&���(Ww�H�=%>�B�]/.�ؐ吪�U�Q���'�����R}�CC�G�J���|��-Wlj���6f�6�����n\r�Ê{�L �g}���~bb����;؎���� �,f�ت�&�>����bx�)�SԼ��ӟ�R�{�
U�X��Ai��q��IN�0�}�oD,Q�z�8mW����̑'5�V��l��	1C���I�Z:^6-�)3Px�"*O.T��b LG���R�L�7�zv�'-����m}R��*]�����	[�`��c�P}���5�Y�)� ��4,p���?�)�I�9ƀApï�}���C��&��O��Sd������y�ъ��&�;ضy��(0�ȘH6�!}Ⴘ�����^������=��pS�D�jUй�sk��1x��sO�C}��_>��S�'�y7@��XgB�:8$��T&I��M��_TkL��� � s���$N�u����&8z�yB�'�ybd^e�'�8� O_\y��4\��Õ*K�^#��9BJV���=���'�t�o�Na���v�%*6mnn��>Y�K��:��"6�֠I�[S�C%`���p$Ds���(�l-ʧ&D��� W�D�P�Pc,X�uȬ�QLε%�pDH����r���d��N���?9�T�CbC�\� ���UZ�$ԦH��C�ȉpX1���ݒ%gBycG��`PnIӦ��8�N7�\/lH|��a������ܥ-bp�j��˄K�,�¡�(�|���>�`	�F�:���58F���m�Ey�M/9�< ���Z9�� Q�Ͼ�0>�d��nv���{Qԡ��fD<+�����E�w�p��M�}�Fű�`
��X�{� �y���S�m��4a���T~h@�.�)Mgx��I�N�4!Y�脆s��m��&ûS�$�X"�ռAPNHۆ-� �2�9A2�	��H��I,T�zY��⎕Ȇ\r@����b�\pH��Ht��@���j�Q>�#�E�J8B�p�L> Ȩ�b�v�+�:
�B����l�M�4��6���%�G#K�X�"'˔s��i��OXP����	�/bz5�'����	NW�.����S*b䉙�'���!p��6g"6u�E!��SVd�iR`�:B��mq"jC��9aMF�f�qO��O��P{D'U�L����VK	J�VѲ	ӓ�\Q���6+h�"���#$��i��O���
��+4B��DJ_���'�l"}�'
(y3�k�<j�[w�d�Ŧ&�/��e����"
^��ӻ{��Y�`N0Ĥu�W�N���7m_�}��
�8(�U�$@z��ٵ�� �@m���M5��#!�;��)�9O�4��<Y2�ۖ?��8QgY�0dA�J[z<Y6�˶)%r�P��Y-7���K�$R"3e��uMj�s$N
��TY����z�m�O�Y#��ÊSO�d���8�^�j�;O>�:�^�	 ��7���t��B�˫i����)�>B�2=��C�fڌ�ɠ������?�b�����=��I8-��xP*���ЈH'��O 9�m
��If� 3�Бc�*`�O�{�H�q��&�v�M%L���㉭K�05+C�x������R6Jys�닯G� �I )����U�߉'���a�x�B�<�\1��@:kL���D��9i��\
��l�'�f�XP(�f�`I���T��'ܠP�U��2�"i�bN�l�|�ʨO`�H�MS2�	4*2*��W.Lm���ӄE������&�.�{���)�.erf�b��k���Z\����B'6���韱O����'4�h:�Q@�vU ��ɍB�}p�'��cN7��;&��7G��i8��$�n��yQ�L�)UT"7��F�]��UN�OJ��ΟHMk�(��@�8����ͷ}/¬�%
�DOF4 0*��X}��.܊��<!4"�1\yX|�5ɝp�2�3@`7R6��c'	�F�'��A��o���e�e��.N���IM<� ��E��R+���2�Z�6�`��.*��E|�M������6�J�v`�
�M��yҊH%.p������I�7菓n�T� �@xpP��o�$\�ҊXn������?0H�3���.-B�Â.
�h�F���>#ܜPcI۝�y���.�j9�7��)u��+A�Ӣ�Ox�P��7BP�h��©u:����d�O�x i�8@��Y��*�y�T�	>c!̬�fA�.���sgjY}��1��
)����ܢ.���a ��)��\CD�( ��el�G����e�DxA�ϓXǶ���m�5$�]�e(��
�.�HP�E�ma��Dz2�x�.�3K[�GW�I�a���hpeW���h�v�کC�N4{������k�:-W.P9q@©&���@�r��`�G�㮍��,@�el��D�q�XQ2�Ҙ)��d�'�)��h̕Q��ʴ��|h5@�x\�9e͑k�l�y��9��ϓ����V�g<�ԣQS�\�G|"lF�l�Fj�υR1X�����y"fD�Fj�]+�� �.�B"dV���O�j�Vܰ���
y�����މֈO��Bǂ�OX��O<���(I(<Ś`�@HA8ѹ�/� JH���=��]�='r�)���8�Iɤ�����ٴe:,rt�'�2h��|�'����	�r��R
-C�E���=1�-"��J>a=��hF&ʕ��EW�THݴ-<Lk���=��� F'@P�UX��'�6mǖ�~M�O<Mi��?�N���L���b4��v��� D�I�	�!@�I��J��	���T?IԉV��l=@/�.i�L��Sd%�$�������Ŵ>��,�&��O�Y�揠b�1��#m5��-?q�'�4� 8��	("���Qs� ��Xm�!]��PJ'ar��h��"A�����E8��Q�wZ`��π��y���(-�m�-�ߛ�Fh�df��7����?����)�w��=��Z%-�~��߷rnaxR���]V*h�>q $H�`�� ���
�9I����>l�����D����S��M��$CX(c���'~�|cd�h�ɫ��!����)r]X���i��b����b��)b�	�T���6c�N�b��cO6d�HQ���X0F�-k��Gxi�X�'Z]h擑g��):�S�i]6|�uƏm<�P�#��C�0���شs^�Ӥaݍ$J2����00��ЂedʙI��hд�V2e��π 
1�G�E\����@�E& `���"OHh��]]���ǩV�!'��	�i�޹	�c��<y8�H1��y?E�ܴ}ô}��A߱e���SӞJ��(�ȓS�e�cά|���R��>{�:��Of�q�̄6&���D��|Fy��4��U�%��3�E��K��0?�!�$p-8�����Hqk4��D���A̘�?Ji�%�O����[��N�R�Ɣў�y��	�"1�X�w����2��V*;�
�1�tL8��˧3XX�@!�X�<9�֜��N�k5t���E��<9$�H�h���RK׋:��<��ӣt�52�A��pd��4fdB䉝y��<i��N�3�lI��9R�p�ۓ�m��;g��6%�N�!�&Fxb����ZUm�9�0�Pg�N)�0?1Q�$7�\�+O������|j�{�  A}^��v��K��� ͕%>�`��-�;,Ɯ��D�>�1����@/.c��:͉q�Dg��d���9#���l�Q����yr-Br�$�H�� wOʁ(�N��y�A�*p��Vc�\�ç"�
���`�#m��!AF��&ֶԇȓ^%9�pD���h=��8�<���*��<y��ƃ8��!u��{���d�14��� �Zh����a~bŞ�3㌠K�@�N�,t��6����ʧd�����0�0?�@�#<sP��C�;�Z��_n�'W�y�o
=7ziCvh����-�h�r@�Ӥu%�S�ł��!��J�y ��S��_�UIT�C<��YULp��O�E(�s1�O�x�Z���y9��s (B�~;�'ʄ<�c�¬ �(|Qf��KUdUzI�P��.�:S�Ʉ�ɫ�`QS��Z(WW��b���3q�B�b� =
��@�.�pa@A�� j�C�ɵcM L(�(��W�1�Fb�}V�C�	�P4���Õ�A���0t �>G/�C��.��T:Vk�|.�	0�	�dB�ɣF{��tƖ?� ,�c��'�^B�L���qR�^�}�t�1�@�}6B䉸2@x��vO4@���E��j��k����j��O?������)%�~#HD�A)��+�!򤄖"	��
��֨W�,�Z�)����DW��V���I0T���t|X����U5���Su,�`�0O�ц��}��+D��xX�`h�"O�Œdl�k�8�hy9�A剒�������,3>���P�ˢd�� �ƍX.�B�	�c��S���s���u� ��x�.A819x�"~��
��sTA�`ǰl
�(�C�fB�Ɍb��}����0�z8�t�؞=�D�		��YV�'op��&�[�v�RY�'aދG1��S�}'吲Nt�"��c1��ۥd�O�8t�m D�8
 o/[kV�;�0���m9�ԆJ�o#�'9�J`�◂w�P��X!@;�I��u�ƥ��o(L\����L\oںP��-B�}���i����CD��rpJ��Q�:m�8#�'�J`yt�ƫg���2��/Ƥ��'Y"8��"� �.,�qLЀ<d���'�줊U�\�J�N4���B�Jx:hc�'��Ph�+D�1p��FGB�D��,��'Z�$��r>���<ʭ��'�Z��ǆq�2Q�B�3/�� �'�l S,�q��d;!�^)���'Y�р$Қ[�.�IG��=)B���
�'BfhɑC� .1��Y5u��s	�'#��P�+)� �����4>Ut<��'*>US�*��q@&�r�$��?�LHj�'!j��C�5����Y�2fa��'��0i�C7�2\�ϊ���$r�'E�J�DՐ:VС�!�?��C�'̺a�T
�~� ���ޝ	����'"N1�A&M{��������-���� �����֏}�Vɻ���Z�ԁe"O�mQ�$�:T��d
�A�D�"O�a2tꂋ=l|�+� �oI<(�e"O�=�2S��*BAߜ-K`�I'"O�ͰnǞ�LX#���a�.!-�yBnyϮ8��-�o`�U҃i[��y��$��)`bb�h������yBD��q:�$�1)V�)�~���=�y��_U�Ph�U�v�@��qŘ�y�J�, �lQ�'��d��+�!C��y"�c�PM`�I�]|�p*1ǐ"�y"=b�"���]�>�A-��yb]�N��Y��g�Ƽ���ի�yB�,��Q��e��K NO2�yB�֎_tK�s��UP�OYeb��ȓ=�.���L�gX�XtH��)����ȓ2��rɍ�Y��5)��H=n9B݆ȓFF�eQС\hؾd��&�7M[$<�ȓp��X���z�`��Չ�d؆�[��LzB��X~�iqm��~�> ��J��h����&^܀y2�nX.��ȓfH��I.HXb�: �29-�	��^ʹ���M�0�l@g��[��ȓ&��y��V��£"F(6{t1�ȓ	� )3�
,��EQ�H��H���r, �ೌՠv�ᣠBK�̆ȓ �:��O*Z1�%a3E�M��݅�~P~�[ҬU�"���Tg4>�
���*�|MJ@%�+:\Qモ�:WX���{`L�3BOX�?a�u�1^=8����ȓ&��!��՟��5z�	]�!���ȓ?9�+�!�*w��xT������ ��Q�"�-�q�W��)���B��� $Q�<PLL��(��ȓ8�,�����7|N �ec-qS� ��m�^�*OE���3Ԣ�/%�؝�ȓ���8��45��1��aF77����q���	�I�wx���ꁻh�ȓ�������a�Ŏ��x�ȓI.LaW�$/��� ��~�\���z� ��Ħ�epNx��'�����L�𒥎_�mOֈ3b�e`*�ȓ?6H ��H�~�R<��gN*By�ȓ>	^���΂=b,@3�Y�e�ȓ&�1�ScA-t\T��&����ȓU��m�,�%cٮ��Q`V�w�b���D�	�@���F�d�aNʥ��A��rWbC�	�VEC���=�	�ȓ-I�{f�A�b[	�2̓!cb����Bv
��d,^� T�Ac�oJ�_%@)�ȓ%�z���J�Y�b`��]�J���P�D��#�D�H;^���4���ȓO��ڴ��%#�l p�>Ov��ȓ> )$I¡�й��l��ÂQ��a$��(�^�|���A�8y�ΐ��4���J�Ά+#��	"��;A9nA��	|ꧠ��kv�pXf�]�m���J���1  7��B�	z����ȓ]��D����+�x��f��S�t���*ڬx�`��%	�����xrC�	� �:m�-�9w�����$C��B��>a�ls��(ɾI{� Z�J֖C�	S����Z�U>��)�B�h��C�I �"�qF�Z7D�횲o��JNB�)� I�L��vl�l:'�Qz"QPq"O��@E�#i�2,��XUgZܺ%"O�EY��T�q�r�;am�=�m�2"O� Pdc��r���´Mی`4LEB�"O��4�q\l���V|�c"O���&aY�:<�����N�����'��O0�SY�)v����ҋ\��Ta�"O�HE��"y�T��/M��т"Oбj���4_I8`�GI:�h�9�"O.���-�#���i1f�}X`t�"O����-T%P���%�a6��"O H��Tb_��f�	�P����'"O��s�E؎j1Ԝ)"BV=\ȸ�4"O��!� Ȧ6{�8�F�S�F���"O�ThB#O+l�PH�w��� �hY�"O
{ǎN�Dd�d���_�@�1"O��egX�S�6)aW"����""Opd2��\( ��@�d��F��̹�"O.��WD@6S��h{�D6:�� "O&��L4�M��E!���"O@0�k����\C���BkBHR�"O�餫]�x�J��"3WZ���O2�՝z���{G�"����L�yd!�˲w����+;�����O;wU!���D^�P�H�O���@m�N�!�ē�VT��mP�R� ��+���'�8yy��ۛ!���"釟�*0��'��e�B��P�`�Cͱ1Pl��	�'�Dy���]�-�9��"G:*�@���'�]��Gy���Ɠ�,>a�'�&��o�o���тI��*	�'���R#`
�0*�ڦB.v�� ��'OP�a�N%y����c @ ��'zz](��Ih��1�k4'�vX��'�ƍcu�\#�E��J�	=���"O0D9a�G��q1*P�e����T|�<9���5[�d�ۓx�XRM	y�<�)�).�U�cГ4���lV}�$)�S�'~N��!T����0��}��L��'\�,�Le���F�J.�(̈́ȓ1�����-Il8���J�*نȓG�����h6��thX	Yx �<Y�$1��p`.A'..��)���
>:p���c�*5k�gGv_|QA��0c���ȓ@��vm\�bH�@�����+UdEzr�'J� C��*t̔AB�҅v~MX�'��[��#F5YL��A���%$���q�ָ_�SgdȌ2[&��/(D��b�Iy�=#�O�\?�fo;D�4����X�TC��A:2���!�j7D�Ȁt`3A�#�`@9o���5D��!�L�S��<{a���Bb��4�5D� rԤV���˶��(`[ �p�1D�PJ��S�K�i���PDy��#��w؞<�$�S�,�a�3A	>���� LO���KR*�#sx	1)�hC�H`D!D� y�O+ �\�U�8Ja∃��=D�P9�oM^b͓ak�(T1�0 ��6D���!�P��$���Y81�����7D� ����w�,�ǌW�,-:UYD(D� q��	s�摸�Z�B��`�&D��밬�

��t�%	�Q����c&D�9G���}�� ���U�"��H�
&D�`�@���B�[�"��D�ґ�B�1D�� 
�
�'"rS�Uc	�226�K�"O$Dr��Z>`Ռ���];�MYW"O�$y"ME�<K�ěR'�$M+��[P"O���va +�n��u��R�X��"Oj9�C,�1�Xp��ɨ>�I��"O��jr�Eq\�;)�h4��"Ov4����:Pp�եL&Fΐ�Yf"O�96l�2eo:�a�b
H�ĝ�V"O�pY1N�^���Ϸ1Ȝ�6"O�I!�hD�&i�dI���
F `�"O�a�F�C�Lz��hML�{��Z"O`,04C��	;2����qZ`�ئ"O�|�У��\���ڂ5ODH�D"O�mC�Ȕ%��#��5)�R��'��Ol�����0�Pe{�#Ɠ@ Xͣu"O9qgU�gV�8�3��+�@|r�"O�Ԙ�D�e�x�d��Q��X�2"O�����62�L�s�C��M�� "O��Hn�?\�h)��X�	�
%��"O����GZ�}�>�`&�O?t��"Oi�Ǝ�4��(�τ�+pT���"O"��e��m�v1�S��lo�AP�"O�m3���l��2ƫW�|��B"O(I�Al�3"Xh��%ݪ)�"OB�H�7!�af��	��m�q"OF��g��=mQ�%�/Z��E��"O������*|fչQ뎬#��R"O(��7)����ݑ��Yv�K���y��͂2�F8���	�T`T�F�J'�y� ˆy��txO���ał���y⅄�RK�L #GPF�	J����y���%b�sDl
"C~�A��h�!�y�'��ǔ�Ʉ͖;12���l�;�yR`�s��!��5��@!���y"fģ*~��u�S'I��Mۦ�3�y�%S1f �P�Ê�D4r0fÀ&�yB�V�Z�ޠ�eh�g�fa9�e��y�ÞO�Z�%ȒP�Ԣw㎦�y��I�g�I���E�z�6gF�yaN`z����WPp�I�v�+�yB�X�L�r�r0Ð�R+��p���(�yR�Y[���f���F��-�y�NE#7o�a����
h�X����y"�V(�4eC5�ؠu��|�$l��y�O���||�3a��o�{d���yb��z��Z֍`q�E���!�y�eC{:�i�$�l��ʒ)N��y��N'S��YAB�	z�*@��F>�yR㐸mڂ�"1�n���B"�2�y���pVjqtƀe�4��ԅ��yRn��ck�	bZ�g�����/Ҧ�yb�^E�����=S�0�N
�y��њ��m@7F�v~����/��y���4���1��hX4
���y�f $I�� sW��qN�i���y�E����j�(v�E@�E�"B�C�	4z1��QG*�;��i薄 3�@C�	%�P�9��H������S�uaC�	03:��BV8`��}H �R�/��B��/O4Ε�����)8�*C&i�^C�	�A@�ơB�.�h�g(͞t+�C�	<a��ު.��e�&���A]XC�	�BK`�p���/V���j�&mB�ɐ!hr̚�Cf��-@�D�	~9�B�)� R|�&��3Dp�Hv�$t��"�"O�1+��G�T�:$	p���<f X�"O�·ĒXe��:�&F���(�"OpA��΍6�@����Efb�u��"O�qcem%c@jА�OI./�v���"O�`�`NC,u,ı�.�) �FKr"O�$�D�M+�|�	�_�y�J2"OX�9"��7��,��ي8��kv"O�-Y�������5mY>��0��"O�򅊈��=ۂ��l�X�#5"O ��c�2�d̘ �K�\�t�6"O�m��gJ�U�^��I�Y��$y"O�)��/��:a�x�h��
Xq"Oę�0��4�6á��"��se"O����Cǘ/����K<D�R�"O��
�C_�rúA;�ɓ5h��"O��Q!kY��"����WO�6U��"O��h߱m����@`Ŵ3��IR"O�Yʢ�ޮ(�D8�͝)�^Ȑ�"O(���[�$4�F"Q�D�;�"O)I�/?�P 3A@�(���z�"O�p����2&�,�f��Pv*I�!"O�a�C.�SW�ra�M�uD��"O�}Rr�ިd��ɻ�o�o^l��"O�]:���Vh�Ť����)�"OD��aˍ�X�(#D0B�<EA"O���'8>B�8�������3"Oʌc�h�-4�BmH�с�ڐsS"O���P*$`�ܐ�]�	��Q�B"O<��3c�������b0"���ss"O �y�)d�y��͠��!��"O��B�I�0	�\Y�G*���<$p"On��W���P�w��y��"OF��ө�.����w�
�6�zx!D"OL���U��͂��U�Y��S�"O�Հ��ʝ
�z�3�jİ!�T-"�"O�P�$P|�c*��N���"O�|$N�>7ܴ���G�:�>�0�"O��3c�"�d���)�x�#"O��k��@�z$�N��8-�)�"O"%�b�?����V��/$���"O<�i$c>���@ F�$���i@"O.�K@��C�� R���Eȉ�0"O��Q��ġ^5��2r�i���VO�!��� QZ�� A�=�0�Y���5�!�$�=d'T�
^���e�@�	�!�d�_rD}�'��zڵI�`��Z�!�9N�e� &�DZ}� �Q��!�d�� ����"Q#9oZ)��� K�!�dN>U<��ޗ�>��&�%V�!�
(%��3�!BI�08Kb$��~�!�P�P<�m��K�'n��@�h��/�!�DG�7�L��b9].���U�aQ!�0j,��d�lt�ĩ�A$<!���T�6�-_18b�٭JV!�dT7h}�IA�j�7N�1�LxE!�D$%#�4F�:�P��d�΋&�!�d�"@8{� �,h�|��lFes!�P���h��;����k�l!�է�`�� ,��g�ɮad!��W�+I&����A�>���9`i�=d!�� 7��������ؒ'��/�!��_
@�� ��:�b`��&�!�$�1r���C��7R�(c���1�!�� ��q��h>~�㆟<i���Zf"O:�b�c�D��Y$�ӥh��ɢ�"O��� ��_�b�Sp�PF�R4x�"O�Lr�ɚ�BMp��ikF�i�"On)�n��m��]���M3cw���"O�}��+������*I,�	"O�4���N:K�d���j@1C����"O$��3>��;@h��e�B"O��XP+S>fg����Z�O\�aR"O,��vO�zMі��.���1�"O\�!���0Ѻ��6��@���r"O8� �ŋe�. �у�Q"O 8�W��7%3F���)f� s�"O����+X"Tn��6��#=�"��D"O�HRG�}v�� �K������"O�cĴd��6�C(^;�A��N՘�y"�UR6�Qӆ�]L�D��a��yb�T?j��z��I�?"�ܺ����yRΐ�&��aH1�U8؎ԩ�h߽�y����L�� �����(v��kS
�y�'_�eyـ�Nщq�RE��̦�y�H�&w�xA�(��xKp�CHH�y������8���u@j�@����yR�W$kǜ���ˎ�p��Th0�޹�y��7r�0;em:f����G���y"�	;H��KI�+\XɁ�BH��y⊚�+!�lÆ �j�f�0����y�"��h�7��h\���c7�y"���|�q��T	`0������y��*8�\1�T	��TY�h�ǧ��y�MLhlh\��nџ{���Sg`��y�B��.���ܕ}F}rF����y��prqSQL[�t�����y�łnd\���۽lq�骇ə��y҅�L�̈�5'L1�"��Vb؂�y2���mڸ���Ϧ@q\�P�̅��yk�%�R�x7Kg,I!3IB4�y2��#c߰h1�Ju�hY b�y�-k�� *�܍h��A���y�Q� 0������__�M�$MϤ�y���*+�-��'ʟ]C`��2�yRa��FBrP ң��*�M�V��yR��$J5��T�Ta�@R6A?�yr�ͦ6Қ����<E��-&�D�y�J�FV�a��D
�82L���X��y2��{��x�`OR+L쑁�	 �y�/��L9jS�BL*pt��X����U�r��#_�j����2͐=�X��ȓ}1�IA�k��kE/�>n�r��ȓ0���R���X�P��0��9�ް��"9�ɑ��66��1��+
�G�H��pCjū�Þ�e_���%��G�h��_a�L�Eg�خ]���Y���� (�J]$'[�z4����`���Y�p�`D)}�0z�E_l(�لȓWxrm��Fڊ^>p2�*ބ%<����B��HPC)��ȹ�F�Bb��ȓ'�" r���� ��2FP'iT�̈́ȓCr�sd"U.3�"�HV#(H��nM�M+�Z,<dR�g�.�m�ȓa(e�aJ��l�I��&�@8�ȓ`�l��ׂ��o�\�Q��B�qnU�ȓ%4e�g��>)R=���_�Z��5��n��$i /�6��}�q�O�Q����S�? h�b0�T*�(�34���1��)��"O0�2;F�,��-��G�b�"O�D�l+)Xq�A��|��;�"O�I�������!@�&�&��"O�MR��	(f��Ty�M��{�ٷ"O����&I�\@�.S�{�� �p"O` ���=^���r��/)����7"O��`fФv �S��	�(
S"O&��2nŢCd������!9Ml!�E"O9ç#?�`��Q��3+Xic�"Ot��A	N�U\C�  ���"O��q���"/�)Q��$�@-��"O�d�u�Λ ���&�^�=��\�"Oz��˂6auR܃�� ��;p"OJ��ՁA>80�lP��Ƕ˲� g"O����L��WY֙1vB���mj�"O<�tiB�1E�ȡ��Ye�Hy'�|��)�Ӳ�=��ȒbD8�+��х
��B�	0d���HN�X��3)Q�hq�B�I��v�zP�W�|���$��62C䉛a��T��鍖a���A¦5�B�I�\CJ)ч�?�<SE�3z��B�ik���ኞ�#�T�`���he�B�I�I�z�b���`O2�F�Ѭok�ʓ�?����?I
ç$�le#wh�O$�i%��;�h��ȓB����9=2I"c�d̅�b�J���g_:Ob��9V�ü hZ��p�j�ÕI��hҘa���A�����eh� GF�"R����HͩP[|�ȓ^�n�q-�q>X�B��Sk$D���w	��{�*PA���\��#D���.�j��,��@�^��D/?D����5+��0�L.ؼ@�<D�p���Ǩ9l�]i�ӀT����;D��h �J�L��uF:s���%:D�P[��ˆ��A� F��J�V�AS�8D�4�Q'��V�9̶r�N\"c�6D��{��K2,��%�&��p��3D�� �ȇ>"��d��E�����g'D�/�g�r���@W�ģQO$D�������]�W	�X|��"�#D�TY�I�&k���nA �Jċ� D�\j���c�Fd�r :�L�X�N?D��J��:e�&}H���\2Q�UG0D��Y��%�~���o�&O��k�E�<I���S3~�1���5���ϋ�a��B䉺4�hH U�ִ2��2��|��B�(}�n��QMۊJ��qB�}\dC�I\[��ygBS�ҙj�.�B��C�	=
��@�Pf�Kft�3��(N��B䉈*����o]��	��V%d?jB�ɫ< �9C���w�8t���o~NB��8��BAM�|���U��+HB�%/�̱�eGG+���0�C�����d/?�7�ɘڈ�Х�Q�=`ΔL�<�E n ��+��y�N�CDA�<I�	C 8shy:���L@ �/�S�<QU�νr�z%!ˊ�o������L���G{����'��P��:?��u!U�t�|���>��}�$��'��5���oِ��C�	%<�m)�k�2lw�m���2@C��=���%`�y���A�FC���<�-, �1��U�U=2a�B�.D�83Agۙ����U��p��9D�� �Ӧ

�@���C�(@�)�v�٦�'��'ߎ�Zd���NB4���O�<�:���\��E{��I��3zڄ1���JrЭA�D�h�!��V�1�J�Ndf��dʬM�!�Ė�oJ��sQM��R�ReR�`[;b�!�]m�6�r��2�j\8����bI!���/5:]`����=������ P!���֡�E��!%��clv7!�$S�E��1[E`�',o�L��Q�(!�'Dў�>�����R}�hH5(�=d���#D��Y&ៜR��-(ѡݭ�.�+��,D��9�m�s�.8��ǆ���!0�(D�h 4 ��*]s'E��
�
@��%D�P3$�3~ީqD�W0M:Y�U�$D�0�#�%P�f��kX$xIeL ��_�'	��3����U��%F�>��C䉉+g����g;^Ȑ�H�Ln���hOQ>-��k�1%nňD)��K%֠+��<D�@�ƕV*�!!���#��`I��8D�4;r�c~�ڴnD(s�8!�)D�@�2�F#<�bɠWR�e�r*�Oh�&���%Y!�RX&��,7b���u�����ɽh$D��3��E����wpB�	�{fՋ��8�ލF��2\���3�S�O�@����:%�EȦG� �+P"O\�[���d&�3tB�,&�F�Pc"O�u0�j7HR�*��T1�t�s"Oz`��N� q0��K���p�`�"O�0�NIaRDE���^�"�К��'��Id�)�'v���!(S�L�hXEF�5wҕ#�'�\cC�X�x����v��"X��!�-O��=E���`�L�9���;c(b�x$�S�y�Fգ��ؘU%�kH�[�`��y�k�j���	�H�z�s����yr&P5q:B�i�*N�}�6�Q���yreX&?Rj�ҷnJ�p���8�*��<��dx�x0�4*C;'��j���R�!�䋕}���cgѸN��U[Q�0�!�d��*��$@C3�:�j����It!��	Vz��q�iE�B�`�z��Ѕ��X���BY�Lؘ�	�e�f5��}���(��
 +�
0
a[\��t��7��M�"LQ�Y��H�`�.x�u���z�/'�����]|� 	��r�A�ȓ
+ȕ���]9F$I�#%�Zͅ�n�����@D�"���e�p]��C=��b	V�2r�O0+R���
�CG(ɂ65�}:����g�D���o�������&��*�k�0-6Մ�)p\ѰoS65�ȌrG*��K,�$��?��?q�OڅёkJ�L &�p蝤�t��"Od�Q���:���H�EM:��i±"OX(0�KK�y���	���1"����"O��2b_��jh��!\j�5�s"Op���Iтe��Bv��g(�:%"Oxl���)oa@l��.�R񠠻`"O�:��@ v\�ٺ�m���"O��S�AO=��l��!�>���"Ox��`V�M�q��<c{n�@2"OuHR#��)nP�(r��*l�n]��"O��A,�;%��K�ĳI���	�"O^������CpP�أmܲ9�$�"O�(A���M�vAbM� ?MzAs�"O�؆"�'Ojp:A�L�g:J[`�'��'V� ��!s��5l` ���ՠ7?h�"��$-�S�I6.=��#�%�v��@Ӟ<�!�d��T�*Ԉ2�]�s�ꠏ�]�!�N�>���+u聵nƄ2�l�n�!��#U�b�Iѫ��Y�T)�i�4k�!�d��M8hr5�{�� 1��L��}�8��8U���G���fW 2�O������̋�4�N�ʎ8�	&�@�	[�Sܧ?�D@)#B�2p����	�S�4��S�<���W;~}`�����s-�5��)���t`��2qK�O�لȓ"���p-����y3 ͕i��i��U��%*BDC�DD�D�� �S*����n��h�~f�#1B�~�8-��x�nՑ m]�"�
�kT.�-KP���I���Vc�q:��2�*ڽ`8h���f�^�i�4��
&�� H9��ȓ&x�<J�E�U08�)����F�&���G��r�j�� ��[�d�4F�ƨ�ȓqfс -͚v,p���a��Y�ȓi�H��6B�?m�pq���PDu��#@����W:2�^�ˤ$\�_°�ȓRά��3$Ո6�����+�$(@�ԇȓ0��]�W��/��(HƧչ%Ӟćȓy�D��J�i��UAUj2@WX���[��e�v��o�):����g�,*�e c�ļP���8�{!�D��o�p�	c��6�Ze+%d܅{�!���5-�\Aua�:n����%րG�!�ǡ9��)�M���:�EM�u$!���q�`S��0�����m�	J!��Ă�	�K�I��<k#,�f!!�$�4Q�8qB�	S�Li�!,��!�Ą�:V����@�0x��� ��!�Ă�Z�04��C\��x-
GЄA�!����׆Ùp5~]`bg�?.-��'��0g��r(�Q��,Q�Iy�'��P)���L��C2��8w`r�'"��B�
�DlY!�D�i.r��	�'漌P�և6�V��ذ.��5@0"OL�����f�Q4a"�A�w"O��C�E�o]�\���XYL��R"Or�##�#��i�!�/|D"�1"O���5�%P�a�f�v��"O��&	�d��m�1 �4rgI6D��17	Ɂ��Ó�ބ>ʐ"�1D�\su"Xno:`
�M�FȞLSv:D�@���@�5ȓ�4Ƭ=z@#ړ�0|���L��xq@*��i�|HC7lW}�<��F�3QT�!� L�$��"��|�<y$n�0)��xS#o�
I�X��O�Q�<ѧi�� ��txD�0'K�J�<��O��w�X b"/W�R���q��I�<a���4W��AV%�$0,� �ňp�<��]d�@"�4�Ј��^j�'�a���|��릍T�Q�Rܱ�쒱�y���6��� �Ì�LN�耋£�y�#�$yBL��Q�RI��=���E-�y�(β#=�@��^tR�3�D�y2�8��ءThNo���R#�y��"�*��r�
d�����d&�y��	ǰ@��dݑde ���y�lŞF� IJ���7T*(:��ybAH2/��N�<�6��E'Y��y
� $	⎫X(N�B���&�R�R��'	ў"~1�$5����p"ȟ�X�JtK÷�yr�j@��@Yx�h���"�yBոZy����B?���y�-��y6E�P���
�+x�X�!����y��Y�`ݬ�v�k�hQ1!!S��yr�F�{��Q;.֛V%X���7�y�k�"����p�+N��1A�3�y�е*�A��^?L�J�CF��y��ɋR&����"5T��(�B��yF
�2rh�`D�:C�Ɛ���[��y��T��T�l�>�2����y〛E�=���ًaйز�	�yR��,!��]H�坰ak���MF�y��= ���K�&_��	�6\�y��JV+Pfi^�X�)2vG�=�y�#� w�p�����Ř�i�"�ybE�Dђ���)P33�;EM8D�8J���\�~�tdϜt�!�P,D��z�AP�NA \Qj�	h�r�*D�X�`ҾD��>(�&��K(D�8�a!ͷ:�:d��o�%�QSa*D�d@���%/��S�H�A̚U@� (D� p%d�+O� R�7<]D��6+&D�X�@G�nMx\��
Ѩi�pP���/D��؀��RM�<�&N����Agm-D�|r��վJ%�E�qn��j��=x�*D��h��L�n�2�M�L����<D���M� =�ᒷjBq��:��6D� ɂj�cN��R��"�b͢��(D���I�aG����0B5��X�J%D�t2Q�P��0��\��ٰ.D�(&��3t�幂ֺv�x2,.D�|���+~D��k���0<�t��+D�����:ђ-2���*}KBLx'L(D���8R�X�+��{�*DJ4
9D�i$�Z�$����?r�فE$D����G�*��� !0�04�6!&D�|�5�sh��bVE�$z�'D�|����?�:�k�%����J#D��V��2L`�`3k�2&���g&%D�P�2�D�!H2�Ʉf�8��b"D��zVԏ>��B�㌿_���6L+D�$��)����ݯ[�<QŁ(D�����E|V S�*���I!�0D����L��2�aP���f�B��<~w,钓F� C�z�HV�Dv�B�	�yf=rEe,X$�!Q�ƾT(�B�I�"�(��� bݾ@A��%M�B�		qAjq�W�B2vzaS�GO�8C�  ���xpn]�.�P���k
�7�C�	� �ޑ(��ߟ.�8s�F*Z�C䉾WD��"l��B�ʀ��d�6��B�I���:�EĶ-�~�"A��"O��tDlqD��(�y�"OnYZ�������?K����"Op�K��u�%��/CR�9R"Op�%��0oҝ���6w3.əu"O��+1-�.1��x#
5_Ȥ���"O�aC)�j�ZA�K\d�,h��"O�Y�u�Z,l&���)�#��H�"O$@+�O�.�btu(�:�:��"O\�H"04m����gW�����"O9�� �Pt�F�f�e�"O� ΅��L<n]�=��%�Z8��"O�i�"M��������ND�{�"O2U8 ���[�L,p&dŤ^/���c�<!2&[��3�H�v�B�\�<�
ί�0e�O�5~DX1sfTY�<�1Nծ/��Ts�@	�n�Z4���
]�<�3`�>7<d D ��f�h��d�A�<�ĕ1
XB�#T.K:`[�FYr�<1��H�D��
�'@��c��k�<�,��}$^	{�HǤw9���k�<aP-�+6��%�8#r%�v��Rx��Exr@ɠ~8�È�F ]��T��y�ؚH̺pzSd�
V�����"֢�y" G�`T�PI�)�;'^���5�yrJ	�1�i��[�����მ�y���F�^����!��d��S��y��,V��e�^�	cn�z�!�>�y���f��Q�HJ�u�r�&���y�N�LH�3�&Z,cYy��K2�y"i��bJ��i�Q|��۷���y�.Q;|`�� �'��ta�``͟�y�`P�c@̻�h�iT�+@�_��y��Q�H]�`.�9k�(�������y�XoI��F�U��y(��ɽ�ydI�W��Iy3�O�H�����yҨ݀]�<��S�U�U;V�S<�y'�bp�aP����Ƙ��y2JU3:M+�C��hP�Kʷ�y2�]�`�n0���̸� `�-�yR�-� ��B잶$�2����:�y���4�p���f�~�t�M¾�yrON",Վ��O͋QT�I�l���hO4���B7����8�L��G�=q�!�`��`���Р�;�!�d���>��S"N�@�!��=>���0���/d.��{E��<!�!�$�p����;UA>(Z�F�4Xk!��>a�m)���A1��rgg��a�!�$@���C�9A���X��J�(!��R��)�D�ڏO�T��n1	!�DC�{<xؔ��e�4q�5��!�d�.._,zt�A<倄y���!�!���p&��2���͂<�FL?(�!�d�1O�X��񊖑%�C�M��!���p� ���`m�ͣ�	7/�!�D�{j�}A��xd��z3��f�!�$�-*�R�1�A�tQ$i����!�!��
4�l2�U�B���>A�!"O�2��������/r����"O"�Cp`ZW����-�a���("Of�2��
&�(��GAY�(:j�""O���χ/2nk���3>���"O8��櫆�d���"Tb*zȲ�J�"OxTz��J#gَ4ʓ��o����B"O��h�
�%v��9���^=�h�p"O<�UMV= �w/A�g$�!��"O�%��,���� �Ѱ@dD��"O橢3-�@��P��ʴI�lЅ"O&��qЮObbԒ�?S��2�"OB���'���jT8*��I�"OH����>)0�+W� G�C"O� )&�R1a�"K)'�R9QS"Orx{�h�h:����c��z�"O�sJ��#�>U2��$�J`�7"O� �Z�ڰX��pKs̖
V`���"O�۰��A���r��&��A"O�e�r�SJ �ء`�1��m��"O��10Z�8���Q(�2�"OX�3ab$W��t��E�e��q�"Of�kCO�x��| b˘�
r�;e"O
U��C�a�H�(bjo��R"Ovub��?$)!��6f��3V"OĄ�nBq�VE��hSFY!1"O��{!#U*���a�
D�l-�Ԙt"O y�o�
S����)_C
vL�"O*m��N�##�z���m�/I�ӓ�O@��W"r������\*"��m��"Ox8BF�ʘ>߄��v�F#!�&�z7"Ot�Au,�%P=,�i��(�N0�R"O�tA�B�*��P�A�8 �P�P�"O�� M�#�\�3�C(���{D"O4��߈_�N��%b�	_r���"OZ8�b�U��k!!ʳSTѨ6��Iy���ӏN\��k�@�=���:�����)�'.���0� �q3�}� H)/� ���'%��!���7�����rz.��']��ě�j���TiG=iF����'ZxX%�R?!�1h� O�ZߓŘ'Da�� �l	X1J��OMdq	�'��Sa���z���
7H+\h~"��d�O��$5§L'�LH�E��`��q�	5[0�	�'lў�|bV%^
�LHY�P�-k�ƥ��<Q$��_EZ�XZ�X�`��j��0�ȓ[.��B�Z2tb��K"c�5!�(̅�9���Zs�K�}���)s*L�6�b��ȓa���E�',�>���� F1���ȓ$�jP�D"��J�H�q� �rTp���8y~|K�"��N�n0C��&O�L���I7�`U�	c�̌�B6���2νa�?u'ne2�HY!Q�j5��/�A�V@L�{5�����
m��(��`5�p���v@@�FLK�1��Q���H��Q�m 4؛��
��H���F~b_1!(B0��ö"�X=�M���yrl�!/lY�����y�����y�(uzV�!s"�;�8i�ό�y�L�}�>5Ƞ,�MP��X�!S<�y��G1a+U+f��,L�,L�@�?�y��Ʀ̩�d���NӨ� �yr�_�.�SL���ZC��y��2e;F�[s��[���"@���hO���ɘ�3����AX4�@�{w@�)(�ўȆ��;h�����L{S�|{t�SO�C��?�e��"��a9.�(���/��B��x
X-J�|������5��B�:x��)��I�b���	�	ژ~�B�I2|��z��B�J̙b�V:1XB�I$HĠ����q�F4�4JԐ:hN�=ç�]���;+�X@x�o�eu�$�ȓ'�80$Ǵb�q�c��@!,<�ȓ���IȐ �b}b��uN���ȓ� Հ�(�� 
���R���S�z���E�VC��<�٠�^!�n��]�}8A/طs�hX[FL��C�
��ȓ��"�ʀi�,�+B�˛{(HGR�S"W;81)��D2��}+�#3��9ړԈO�����:3��0h���E"E1�"O�l 2�d��%Е�V�aʜ8ʳ"O� ���eÃ��TѴ쏛<K���"O��òBͫYK� %.�$֨�ˑ"O�A�CJ����B�e���A�"Ox�s`j9���*��Z,%��)b&"O��X�N���Z>�n�"�O�D��'�BY����(O�A9��.�8	%���F� ���'1O̍��C*9�$���ɋ7v��+�"O*b��M�v=@Ih�D�7j��3�"O*����B����
֗n�(�T"O�xc֣ץ@�>@�S	5�d��"Oi�lE�~V=��h�����ʆ"O��(dhG�uL�y�MV�_h$��"O��c�bݥ,�.�����. �r�' ���$��3b@����V��� T��`��̳Q��1A*�4��@
�"Ov<y�aŉ\e��As*M`�D���"O&)��#M�-r��qK+z�l2�'J剞l�r�"�)ˢ&�~�"�h�R�u����A����
w$(��#��k��H�ȓP�@pBD�*�b�qwcяIsBЄȓ}��,1�EF/������%0� ��ȓpءQ�R N��z��"0(��ȓ!��-����"{:>\�U'�:< �ȓ(��ժ�@�@0E#E�KO.y��W���;SZ PＩ{!�&`X��ȓW���B�JM�hj�E�����k���h����VB.���!\?72�`�֊0�!��Փa���0�:/h)��/G�!��TAQB��p�
��B&��!�G�,7���� �Y�a��eۼw�!�D��f+<���X�Bq���T�V>L,!򄄋B5��A�nQ
 E�(�!���<Jf����G-kW���D&ׄ@�ў ��	8Q��q�Ɛ8�JA��Lgn�C�I�E/z����=DQF�Z2B��@��B��<&��ᢖ�Kn-:��*6j:�B�	���PСcX!Z��%A���r��B�IOԝ���p�X�D�+3�^C��/%
�|�W	ҙ>ɢUr�Hch�(�S�OPL�x#g�Fޱ��.��&�<�Q���?LO�@2��� ���3�\8U"O�����
V]D��硞�6Ф""O�a��-ϣ(e�yy4�˗k&��#a"O"��������2HOR{tT�"O����A>	@FN�En��[�"O����ЏpN$A��;v��䈅"O� *��S�HY�@��-3�\lPr"O�X�B��7��E�s������:�"O�kX�k��H;�]F�B�)"Or���C;]�*���T�\�!P"OV�bC�(b$�T��(șK`y��"O��b`�N�^�0aBܢaG��"O��gF^�#�(�B� u4�|�5"O��k�l��M+�J���i$�i�1"O���ݺa����Sjѷ{���w"O��9Iۈ9�@9�6��!DnN0·"O|YQ"JD|w�y �2Ym��s�"O����M�EK�x�ؒJOfl�v"ON���C_Eg��B��@wE���A"Or��hK��^�
���$1�6��'�!��"z�sD��06g>\�'#FB�!�#���HK<JW������"D-!�E�h6(䢉�;d�Tb�!�dM�F��}+�,�#$����a�6[!�� ,zW�-;pE�@�f6zq�A"O��I3�Fp^t0�m�Ϟ� @O����P&[��amX�NL`�`%9D�tʂH�qj}�u�Ü&U��Pb'<��џhG�$;Ot��>c_~���cΪ-k:y2�"O؜Cc���u��T]]$���"O4�WA����z�G�]:�X�!"O.�*��ˋ�p�㔠��+p�"O�ɳ��&j�J�[U ��OfL�$"O6Ѩ�Ȋ�����ڶ"����"Oz�[a̤/��I�EN	�j ����'D�'I��=�\	��@"���cĄGCT�ȓ���;���U��Id�=m�P��ȓ,Fp�i�,��Q⤟9Sz�ȓ�����{,������^ ��=j��"�5?p8xW�T�a��	R<@b��`�dA#U��g��m��O�Th!�ȱ�Ly�A�:����?a���~JDk�RL�	H$/�0Y���	P�<yD��9V���㐈ܽ2S�� Ҏ�U�<�%�(�dT��*��pd ��BCg�<Au��58���R)
8L����h]�<IG熭'X���U��7,J�Ei&��t�<���
wZ�����4���{��f�<��.��а�.1?v	��Wf�<Q �I:,���1���@Z9� �Wb�<q�/�2OK*(k���1>t����_�<y2A�$6A�d��$��a�Gȑb�<Y��Ƒ=7؈��/8����gA�\�<92g��B�T|cI�6gό��U)�~�<�BȬԂt��ڱV^h7���ȓW�r�p��x���5�~�$'�,�I[�Sܧ#�Tʡ�vf�-�s�A�Dv|��ȓt1�lr��U�6�<<S��/ =���ȓZXC���0i����*2}�0��1YB!5oW�wʸ�I$�����y��=�X$�C�;7�pQ��L�e̽�ȓV�n%	�c��l��9i��49C�5�ȓ%���	�,H�$�H��/�(HG{��O���A�I�wZ�8���4F��0X�'/��G�H�Uix�"ŝf�p*�'u<���\�%��A� �^�f��'@3bj����s�ˈkV*�(�'�f�9
K+II�ȳ�E��^0n$*�'�,�CV��/7H�]@�[�P�X�'!�Qy��@p�p�!�D�1$�R�'1�#,�j
��LQ�&ؕ��'��!#W��2ǐ�@��~�a�'q���s	Ĺ ���1��Ǖbi\,�	�'�i���
2(Y')�2����'��y��(ҍ^Ѷ)G�Ÿ�{�'��أt���*�Nl�!Q���dz�'����B�j{�H���h6(YK>�	�@5V�JR���H�gS>8h-�ȓF<T��"��x �11KĹz+�X��`�^�٦�(z��xW�h����	S��puN�'#��ڤ��Jar@�ȓp�T�;�֘Q�xE�˖�2���.�0���:�v�H&윋E��ȓq,����ՑQ�`�� ��4�n̠1��6>�P�Q��L�I𘅄ȓ��YQ+���9��O"t�2��s�h	��9a���ӎ��o����a	�H0%d��s�Qp+���p��S�? f|�A͓;�ޙ�� ] 
�I��"O"�ba�E$3R�@�B��!]�T�S"O�T�����7�6����?of�)�"Oƅ��+V��xsu�O�(�@"O����K�	Z�@�V����D"O F"�;X�J�z�BN�l�<��"Of���ʞ|ɦ1z ���8YC"O��{1GW0w��ۂ�ա��q"O^Q�6�͵r�
H����>�Xf"OT�+�oZ(xttĩ���5�(+"O`��!�o�浣�@�%�nas�"Oh��2囝�L 5BT�K�l�'"Ozu��&نL���xT��.2��9�'"O~EQ'˕��`��Ď�.��h`C"O�M�j��0����)YC���"O�+B�")(>�+��
<�4���'!���9�2es�-�:!����6Jf �'�ў�>��DQa��9�4�W|r!�ro/D�Dk7aƺ?:�)7mֺQ�D10q.!D�4���54����W#x���A�>D�|oĞ�v���H��%�t�7D�`��4ft�a��wAfd��;�O��	�i��
&	*+�����"DU1���0?y�-W�}��iKq.�7Z�J��w�Yj�<B�_�	����G���б�OB�<	2&I]g�`9��l�6ax��@�<��#
�[�8q��qAp��
t�<�7Ɋ�/���k��<yS��F�<��Q)�<9K�G�
l1�8c�x����ɈR��mZ�����]XG�&;�ͅ�~����%�ߍv൨a#�<nh ,��o�:�j_�k��������ȓVybЩ7�ٍ<���b희�6�ȓ3�}���E�p�4����+5B,���V@A�M�K�&4��)\b����x>�x�@� <�.���f�0��l��f.%s���\��)��U� �獟9��Z7�&��-��8�<�$^6\ɒ1�_�j�6�ȓi�h�d�Lw�KC���qX)�ȓ_�P��n�OOI*���I��ȇ�\�,S� O�9��
>&G���k=<��H�B�&���͔7x����1vD4X����D�:#�q��
׀%Q�ʜ/NA��ɳŇ�W�j�ȓ�֍Ф��,��]�gA5W�$H�ȓ!�4<�rn�*o�
��6Q)���v��dO�z~�m���{�⭅ȓ?�҈q���>du2 J�{�]�ȓVyfe{���(+�,���Z0V�E�ȓX�hbя��v����Ζ= �Q��z�Z���n$ޜ���Pg��ȓ|���b	#PI���JM���ȓ����Sċ,����a��K/�$��\�����H�w������G��FD��FiLC��DE����oT1_�J��ȓk���I3����6�	�i�1���ȓ�e�5D�,C�iI6�HW,�ȓMQRl� E�,t"}igA+B�u��]@ ����+8�TŐ�WE�p���e�u8`��-j^x �lW�{�����I���y��IDPto
&}���@���N�%-�( h�f�:"*@��^z�z@���Q�d�{�)B9f�@���S�? �i����:MDp�An��}�2��"OČ�V' ^�D��TâЖ�T"O.I���`�d�IO%M�jQh�"O
-f��vD��A�H��p�Z"OLȷbތ.8����_�'��{�"O���Â?]���2ׂ�S�4ib�"O����϶80\9FO��4����0"OXm9�I#Qkh�@��_(~��:�"O�M���~�|�s�)����"O|P�4���ND�!@�rnhU["O�}��쎲D��@�hU�-5���"OT�rCBӯZ�
D1T�ڗ? �c"OLm0n��o�h-sr
9bz)�"O���`�<KΘ�)OS0'If� �"O���@�m��M>~�!��"OXA��L�=l�H0
e��k� p"O�������^A@LP+�T)�"OE#1�C�(�Q[Ġ#hR��$"O�\鰧�Vx�p#	�q>P#"O�<�2͘-v8(!�ԣ=2���T"O��:@�& ˑ%Ո$r�"O4��4��d����ޅF��A�7"OI�Q�֭�>��A-�1k�"O$1a���8r0 P�K�G���`�"O&���M>m��E��/� ��S"O�T(��ҍ*���NQ�H�*O<�;�.U2,I�oڸ#�F���'�c7e��:�ic���'B�E�wm�`��ip�^c2�e��'��Dc�� T�v3�)���
�'�>EHlQXI9����|��Y	�'ކ�R
+�$�a�B�"�x0��'*�`�AC�V� Q��R�`J�8	�'�@л�A	� ��l�j&~|��'d���,�3�����@=c�d��'wNDX�ېx@�PfI�[JfT:�'Y����­;o��$�,_5��"�'���7y@��E��^۬h��'_hٺ��V]"`�
�.,���k�'�jHɵ�ٮ^n"�W�X�P<ܥ��'J��wD��kvr$z��Lj���'�Ȅc��/E�d�Q�I��`�'&��+�.D�a��Uc��R!Hp�	�'��A�c�5Tkr��E�-:�� �'J�Df�"4��aI11lIp	�'lRXst��R�H�V�M(v�4y�'��=rq�F�
���84.G/&����'���wJ[6V��Bn
����Z	�'[�0zb�4q��$:���Ea�'��hy�샵5l�	�@V�X��'a���1ʌsgԈ���h�"��M(�E3W����/S�i �T�"OL\@Ah��W͒��1$��F��D"OƵz�,~�.�6��5��L��"O`�5���<:����KY1Z�4�zW"O�t�eF�8~����L7&]D�P6"O�X[��R�E��Y �Y.���b#"OZ�)gA@;y��PUH�*����U"O��aA�2{���8��P��t�5"OA�פ��:�Xyb�F��y��"O\9a�*�,q�N�ԌE̂���"OHc���#jD ��.J�~��mڃ"O�p�%���|$���Y�*Ę��"O�I���X+)������2a�"O� � �LRS�:x�� �~lbc"O`�1��ռB^b%Cc&ҢO��1@"O������9^8�!�$��`�\a�"O�Bf/�K$�	�Ý.jPq�"O���c`�K���)�"j��P��"O�����BJ���1��'
�li�g"O�T�pfH�<쥙�O�p����"O����\��2aDҿ�����"OR��
�<���s�(���4ѡ"O���˄�%24�T�C-8y��B�"O<E �k�%�JS�?fRP+�"O��z�Õ"X�]�r��WL(��@"OUA��%>�|Q��(S8����"OH���GJ2yʈ��~n�"O ��e]�8�T��k� }4h#�"O@5��'�U���PF˘)t�1b�"O����֯T!Z�K։ �D�e�"O2h֡�A�3i8`L�<�a"O�E��mE7�mH�W�%Lڥ�B"O���fCو_.~��G��3�(�"O�]b%��S��0�ݪ(�|�a"O��pMʱ���#d�Q�x:�*A"O�D����M�t��N���4"O�@*C�͠r������08�Y�u"O4��C!
	�����W�N�����"O���U腑�pR�΄q��\y#"O&��`��{�+�*��Y� X�q"O�Bs��Qox�� *ƨy�X] P"O���G�@
u��f��<���K�"O��Aq`��6r6P����-;�x���"O�pۤ��:�X�wEV-.Тp��"O���7����Κ?��� �"O��Q�P�g"�u���[PS�"O�A��'�<���ƕ/��@I�"O�=��O�^�%��;�L�A�"O�<9q�Y20h�� -Ir�M  "O�y����0���󌞁Q��y�"O�u�ׅ7eM`�3��2�.�q5"O:���N�6m�m{�g�'$�Te��"OZ�����M��dӈ) �@�"O�9s��_`����K�e�tA�"O8y: +�=`��S3�\�����"O�8a�H?q ֡�"�Y?TX�#"O����lU�sv���eʓ{\���"O ��l��IgBdX�D�HXH�"O���[�r��Qc�X�D��T�"O���QES5 �9�2/�m��B"O�U����" D��7-B�'�1��"OfH*Ն�Q��T3@��[]ΥX�'�2#�J@�gR�ܫb$ާz*1��'�e����g�N���
̝lȌ���',)ȗ/�&ѼU�'����=8
�'��13�ܓ4�TL�q�އĲh	�'���[COX�V����L�|r�!*�'Gv�A��@��1E��>��a�'�t�Xw΍4wP�(ǟ�1L��K	�'a�I�D�E�D����&`y�%��'N�Lcnڲ:Þѡ����X\>T�	�'�����+?ޅ� �Q4VT&)A	�']�y���}�^��AD�\`�b	�'�4��	�nu�O�X�f�K	�'m����ߙ-b�i�T,Y�f��\	�'
r���A�Z�4�3,ln:p�'nvdct��<W�Q�`J�`
�z
��� ƨb�腩)-�	�%L���ex�\x�Q�LR�)b��8�@CW%>�O�˓Pz�[#A�D.��D�
���;�'78庑+(7�����J����Y�O�lh��(��0�􀑀��'+�OFt�0i��>�~$a��L�ᠹ�b"O��b ������ō��ĝ`g�'�V��'����j�޴�"���]kD!�W�&�S��?!��B�m�
(۬M)���z�'Dўʧhܭx�l ?Dp�3R,ѩ��Ȇȓ.��+ &Ғ�����BDZ�����OP�Ol�g�'Z���v�:��d�!�><����9�'D�t4ᐄ���"s�ل@fT��'L��^X���'n�\q(�)� 2��5��*Q�F$�m�����T>�sO~�'̝N���1���:��=b&OP>x��#=E���(��H��9��܅V�H�Gyb����G��Ӻ���B0hh!q�LTZ$0ĥr�<�V%��<`z`�	%+�kSjZ韜�?����O �q֯�"G�����+NP@D0"Ol�Rr�+]������F82X<A��l���i��Nv�(��B�O�v �5�5+�!�ό��#eBϛj��%��d�4�!�t�l�Fc�B� ���1�!���%k4��!�mܨW�����Ҳm�!�d	�8�zp��͹'�,��3.�7t�!�G:ab��{îۨo��`N0�!�d�i�,Y@H��t&���K��!�d)h�4�	�?b�R�kTK;<w!�d�&?�&=X�ʔ����8r�Bi`!�d�17G��z�gGDij ���ʈ
U!��=(�цު`v�)��8)>!�dB�d��ٖ�ND��	�zQ���)��Y@$�ܧ(KvQ���R�g���=D���5�Ժ2>��� Ю ��l ��>�
�U�J��qkM=HѐEdg���$��D��Tዖ]�������!AT�)��$S'��e�-jO�[4��B�k%D����J�
}<��Rb�<��,��6D�쑧����h��AJ�Q�0���h&D�Ti��ՠe3h|��F	7Ur���"D�d��Ew���h �C#���S�j&D�@�XmYn�ks�Z���	(Ι�yB��++����K
�`���i=�y�Å$u_*z�
�{�"�$�(�y�N�k� ����|�dx�4�J�y2�Ǒ���h��ԭ}`�]+A�[��y��$F�5���L@�I*r��HO
�=��-��s�ݼ7���TA(M��|x�'|X��T��B[�j ��7�Iz���X�j����#�I�U�Y��XY3"O��"�bS�A��j��I�c^v�pd"O��J��V�Y��8�B:4UtpS"O�4�q�ǽ{Td[�#F(0�'��kx�\ƃ �f�`��S�2�N��%�3\O�b�hY�B�n���ӗF��^�V}��I3D���`�:r�js�H�~�6�@ �1D�t��#�c��	�K��k�,��� 1D��B�^ 0�.D��B&[��"=�ǓE
�Y���a�N�S7 S9�Ņ�}P*᣶//�.�����t=��m��]GQ��Ï�d� �x�{֋v�[g`��Ma|��|���:�(�]4�,���K>��4�Od�2�Q�f��p�k_!A"���'�� �4��@Ӣ��[�\�l�R�)��� ��C%��pEA�O�`� "O0�j�Ί�ӀBr�)kw"O�%ȷDN�Y��Y�a��#�F�����%���	ˉ>.��A��I�7�Ƽqpe΁�a}�>1���,PB���ѨӰA��"j�<A��T�Y��a�-.����͔e�<qF��0𨡔��1Q��� !Pw�'\I�ቑ_E
�a�"�Fx|MCr���r�.C�I� �!��}�v�4���ZR6�t<��lr���
'h��r��a)�$0?!K<�O��O`<�-�(y��0�v�V :��Q*O PË�ܼL��Pb�(O����\�2����oI�HE<�X�J�i�!��;t}�a��(��y�~����V�!�J	pF�D�Xt�q����PIqO����Q��"�`[�tZ���%�L�nG��nӜ����%���y�?�2�����(\O"�@�\ 	�'f�!�L�0�"O\ i��
Pn��c����K�Z���Z�h̓�ا(�v��!NO8����#%�>�8�"Ot]�C�9l���!$��	)���d��}����Ć�3��X�j�	G�P��Eoĺ5f!�$Q�O��]�A.����USb�[�x�!�D
�;�<�N �x��W�))}az"�dP;0<2=r�HT��2|�t��G?!�DM$2��	Z�l�M�B���A !���x�&��⥗�����	U�;:!�$T?�J��&�ߌ@d��B�3�HO$��d�jp���<
Q:I�#a�%rX!�D:nw��jGǐ�	-b0bg��EG�E	c؟��ML4"ȥч�R9,�U�'�O &��8���8V�j�[�%�@L����!D����EŜh�@����p��dɁf:D���2��&r������A��H0�e8D�t˧E~|��E#}���	9D�dӔ-�4LPn�1+�hff��TB8�Ih/�#<�|2�V�2��(�"K��Dz�$��<Q�'O"0)�8x�3A^ 突Jߴ�y�A�<���h��џ�Oz��q�P�*��5f҉;��p�"O�}2Ţ@>*�(=�p�Z>!|l)"C�ѧ��_l�FxJ|��/E6{��٫��Lwd&Yf��\���>i������@�Ӎ6B�p���hO?��c�ę�U�t'B`�Sf��;4C�0`�t�/�l�Y{�*D ?�0�D���?a&��({@��S �*�Z܈���{�_���O[����eH/=|�`y���H[╙	�'��K�nϦ ���+1�^k�.��'�az��' �0p��bQ�?|����*�0=����g��ӏ�7
�.���Kcπ̆ȓ 8��#!ن��A ��Rq�Gx��)Z�gk����c��0 �$d�<���5��Z�ѧh��*.ߟ�G{��	�%bZ�Z��2k �DA4Nr�������ѡ�#b���$�H�.U+�F�<i	�$d4�c�e�P~>����&)�~�F{��OȀ�)����$���F1FGT��'@����B8- ��d��@b
T���HO$$�e�@�C�P2�e�V��5"O��b���6�X�c��?)�.��t�Px�x`�����AnH�-�K��_J�}Җ�8�f�I�B]9KfF¾<�x�B�'D�(��'�\�&��d���PĔ�r�)#D�����X����#"dl����.D� ��%կNÌ��t��85S���P,ғ�M+���H�� ��S1OV�|i�X{(���!@B"O�!��-4B�x���(:��Uq��iꛖ�)��](R�X; ݮ� V�ʚLVڤ�':D��dG/��@���� ���,7D�� /O��$���Hmd��y��!D��⠂�3T*�X�Pe�&nA�Љ��*D�Њ��G(r�z�ӱ��4�� �D�&D�ܺ�j/�Ƒ#a� ^QL�yb&$D��A�e��=HlP���1�ص��"D��dL$]��S`�z�ȩ���>D��(p�� oh��g�F�+ U�/'D�!� @*A�������p���E$D�3� �#mX(�q	��|�Ä"D�43��í_����A�A�V��\bu�4D�p!���!5�* ��)����K2D�<��`�0N�I aB���=��
0D����E��<�z�������n(D���)�J��`�F
GQ�)((D�<iV��6;���
U=�Xݑ�`)D��SBd_�{�R���O�=v���h'D��y���W$��E���{���VC!D�ȊNO� M�-�e�w�v��)D���7(@�jL���#"ZHc��� �&D�(� @���{��~�PH��B7D� ���P���X
0ů1�]���9D��#�kJ�D�q��l�0q�~��<D����*R�l���OW0@��/:D�T�(�$~6� �l�|����9D�ha��U�$ȕ���6U�$J�j7D��Yk�$%D@����T3_ <`�6D�H�4�v��!��R'zA``?D�,A,�c�^Pkf�M:AHtФ�<D�D0t�"~� �ɞ@y��6�.D��iveU`DtHY�H/���*D�p�񂄎YY�D�kDs̀%�,;D��@fLNj�$ab��6�� ;�I1�8����#n؈�TF��q.�c� �P��V�Z���U&��x�n6D�X觍P	����敍C���)��!D����jڊ4>.\�IL#a��*f�;D��EL�?FTt��	x�t��FE5D�PQ�LT��`]�G�B�,)��!D�p�W��,\��vcS
V'��Cw�(D��x�h��ZDJ)�f�r�˒B)D�i 
G?D��% ��'I:p�%�2D�\��
+|�!����k�Y��*/D���Q��D@�'جvP�Aq+*D��av	�&��1F�������(D�S���0-���Q��0o�viX��'D��!.U!���&U �T�qc!D�8��ϑw H� @��cҥ���2D�2�f� K�Hl`4��Y��(uK,D��$aM�J�I�4Ʉ��p��i*D�(B��֊83F!X�ᗦ X�P�+D���vē�A��x��5Tp���c$D��c���7��PZ�㜺/Nj �) D� bQa_�s"�cP�X�3^�iI!m D�P�$�JP)lh�P�y��)Ӷ !D��kSCů4v�,�/׿ j��r.?D�� ��Ҡ'a�3�
I�t��ӳ�<D��q
τo�<d+�� q��٢�m6D����P?�P�2��-M�<�@B7D�;2@�3G[� ��5T�FqT�7D��ҪW�8��� 2�E�:�ӱ�4D�Dڒ��<�j$C��F"� �%�5D�� ҉����n{g(^�m�R�(T"OM�`��(Sz�ez���b�D�:q"OjA�b�,�V�9���q��Q�'up(�@�I�2)V�b�F�nh��Z�'�*��#�D�a��	:����W�^���'j�M�gCH�K��[�)�	F[�(�'���h��A�W�} �T/�8��'�RǉY�L�`(��߾lB���')�TS��e�T�iFN[Ί�6�*LO^�"��6��I X"�!#�܋X�T	�� ��6M�$>g���$�e�TDRgC��ցÖnX!��'�ґ���X ��M �;�m=**֔Z[\� �
�&T�-��j�]�<qS�¤!^�c-�R�\}�����4&D��OJ��-���O��h[��`���@k��H��%"�i��=�?$�غ�&}l�l��Ϝ"��F��$��U�gH�8����J1,��	2U�$,�r��.0(؉2i�%'p��T^(x`г����$	�&��Q�H�r�@�"��͇�M�TA�[1l��DN=S7��:@�~��Q�FE�2�'����m��`,��'�%�7��U��j��$�����L��!cB˚��y�>%fJ�f@шB�9�b`{��{B�x�����p	��p3H���!cB�  qR$��<$��(���S/��q�j�W
��)Ʋ߮-I5��6�}l��qꮴFLT�6����B_��<ygl� a4IyŰ<� k]=H��P��@qa�ܰ�k��<a`�X�m� c�58�n,YǎLc�:ivp����D�?��2��0[����h�d�*�`.D�����era��B�n(���)-��ĦO�� 0fMX�g�I����RƬ�d6p�p!�N�l��B�I:d�v��.D�rp����+�{o�uQF·c�FЇ���S\č 2EҼ%2a0�ኀW���D^�4��H�PAgJTdM����Q�	͔\A��'D���AG�-t�ґ�V�ΡYNd�G�#D��x�*�/Q԰s��#J��j D�P�FGԭn�<%ۢ�	G�Z1Id�5D��c�\3F%���FC݇�r-V�'D�Zd�R�I�|���o�: K"D���P��'aOH��c[�+���1�"D�,;�Mc6��-�,�z���#D���0A�B�|�ɠ�\�.c�"D�@���l�J��JE#����1/4}B�
:G�Ň�	B+�,0@�ůM3*����F��ē�G�8��ϋF[��C啹v�:l�P��5�ܵ`�'���ـd�1�0� �޾ku��	����a�����䐰�4����f��f�v���%�w�Q�g&�y�l��zJ�'z�+Ё$N�R��� �lJ�Ag�8���� C~:�W6��ˆϔ�W��U��(�0������:�b,�ǡЎ}��!L٤J�H�K�-�g�`ŘU�Є����M��O�D�P����b�  ",��>����"��
� �l�5�q�D�Lx���E��R����3I��hAN����ڤ=�`�+�
9�aBE��z0CV.�d�p�V !U���d�XE�K� ��)� uT�A�f2P��4�мk,��_�xZ�ˈ5�P����f��hzE�Z�M��e��a�5qBbACF֜�:��
߆�qK��7uj|ũ���N��q�1�d���E�&�~��=m&T袭K?[��d��Z���O��`��
�+�`-ʚ'��ܰ��+yV�&OQ<����ʜ �X8b�J���q�����y���YRhĲr/����x�^+.��Yk�H�kf��y����-�!D���9��ȯ;d�����d	75I����nX7h�����Z�h���3i0�U�FL��p?i���-a}����
�l��t�7+d��0�U�PO�/�(e��lΰTZL}!�Q��~-��w8$��#%%i��U�QǗ4r��S
�$=*�l�Ҋ,�F�ۤ�� �P8�gQ�i�8��RIU=KV8
��!x��&+S/�Bc>������)Q�H���1���Z��GBJ�$A�6�
��FH�Ӽr�:�ʇ�]�'��䎊'K��37��.~nȱ+�!\G弼1��z�IG}2�ز@2�I���%l3�������R�r2�F�!XD��O�TI�)C���Q"g�Ea���^��yr` �={�P��I�5L�,���'�b-B�nߢF���B��,����x�%e�� ��r	f.��B��BU�&����� Xh�p"��!�>9�*��<����'.Rt� ��2M~�|�th�,Hf=�/6D4 (��
�M��¤��2�fdCTC@2L���Zi`�iN��r�u,E2.<ax"�@�Mq�OV��7��
��;�C�}�� 2�L�O������p9�-�G�#A�V�?a��Z�Z4�s��� 8��r�oYj8�l�T�Ѯ�d��J�>g�R�F)�e��%
7�'(�D`�j��Z�H�<�Ozp�G*�V�b���է9�Pi'����GC�*Mw.��0��o�@5{�
�,|1�c>q�H�7]�6|�F�Yu��k�-D��r'H���k�
�Z�,y��˟ w��� IO;7�&mA������"eII<����:�ޝ*`�
֤h�	W��x���I8zi:��X)�����A2�F�H��ߘJ�,L��N�)�'�Լ��K�Y���a@�dP��C���߮N~A��ƃ���' >^���d20#��\�����.��B94�$(��:�8$�'��L��@Y1�6�OQ>�㟞pe<��(r}�)��2D���3��&��\HǨ
������;��ɱ�A�Ck�^�3�I�a�����$�4B掝���e����M�b�������.*��6M�h\f�T�,}�����o�<���J'�xB̗';Q�,SR<��A����O�L�Ҭ�98hD@�4/jQ�kS����RA��#E1�ܛ7�B!M�h�R���i<���9Df�y\��Zeg̼�T�G,����JN�?��M[;Aa�!D�z̧`*� �poC8��
 ����Ԇȓ4b���'J��u��a��'H�Γ�M��H��-܁IPmܧ���j�����%�!H���a	W]�9��Hҩ{v���elnT���!����'����6��I&-�1����Nw>�EGCW���	)K��q%��$�d9��N��gC�-@�'4e��d�6�x�O�Y^�'͛�b+��C1B,�f��0��� s�q���a����U����`k�	zH�E v"O�a ҪC�# 1���!-�R�Z�y@�?T=�b�"}�l˕gi�!��I32�@���k�}�<	�h	�
x��	\�O�Ɣ� M�|�<	� ��d��� /W`@tsPOBL�n�A�1�;j�h����^�4�9%��9����Ĝj:!�d�t!�R�W��"LaW+	2@"N`G�#@t�8�����Y��Dj��h#TI�)�BZj5�@� D������3�R�Q���:U����_;(�E��U#4d�3�Y���<9��׻Xܐp�@�>Ċ�rC�u��Xa�O��gN��ҭ��[������?�*��c� 1�����H<�WפM��̺CI ������Sm�FwX�')�>y�>]�t����O��e��L
�q�<a���T�(�'0y��K�&�=bq&��Ҁ��R���lB/P�bV�dM��(��I?v�Rl����<AN:\�G�4?��C�I�s+\b�'"�t]���ԑd"��ء�#&bHB"�OgV-V��NX�0u�Jr�I�;Z�X��P�'A48QTh}98竝	z�0�� s�NL��J���	�$�-:��0wO>���D48�Չ���`a�cP�D0�ֿ+`H����O�L�,q8a�Nst���P�󈖵��q���+�H��$"O�8�!�w¾s���	x��hˢ�IXwL[1%�� �,O��O���Oj� eBI�.9�12q�΍c�m:��'�`�p�3�mQ���Έq���?� AZt��E��̘7a�azZ1wl䂷bY$Ug��B/����O�ȉ1��c�Z��O|���ؼ����#��)��� �I�<���}��8Ѣ$�&G� ��M\Ey��K�}Ђ,���v��%wE*�Q�c�\�f���"E=U��B�I�|
�i�(����{�e@;tR�d�O��BJ�s�%?㞴Jeԟ���:�O
�L���B$+�O��be�T8 X��	6,� ����T�>�֙;�%O�?�%�.p��4b�������e�u�'���s 	��:<$>U�N���e�e�1d^��!�	2D�(h�#����ȉ�e,�`�<q�o�!!F����%8}���<Xt�(��aѕ:9��p�gS(I�!��Ϗ�H�*��[�p)+����O��A��58\���qO$-�� 
n}y�.��at�9 v�'%.1�7� jґ��	d�dq�w&��!i�y�!�#�T���I�Y���N[�)Q������ p��?)7�9hG�d��&��E�r!X�	Ҫ`YLe��e�~C!�� k6,A�fNX�~OʉJ	�7S��9`��!W�)$��S�O�����R=y5����y܊�
�'9�� ���h<�Sd�"d�
��|B$��f� ���yRޡlݰ4:� A�����Px�жi�-酯ͩH��܋W+XYF�[�ƚR<���E�dH�yA��>����І�y�<�d���l���@V� R�@p�<Y�l�3,��i+�&yHz��V�V�<�a���9�`�R�-�ݚ��U�<U�T�?l|�H�FA� s$I�L�<�U�C
e�8ۅ-�y�R�
�@�<Qg���X,����a��Qz���|�<A4�.1md�)�I_�]��;B�U�<yS%�k*a�`�b�r����OZ�<�v	��!��)Ru�CJg>����m�<����J"�Ւ&�AB5�Ko�<Y�+W�'l��b�_�|�����a�h�<�I�1u�X �꟡x�h���j�<�u
ؘw]Ȑ:��P��,Ͳ���L�<�C�F�h<��`�N;* ����I�<�a�[::J�]h!��&3
�K�_K�<a&��_!~Hi'V�4"dq�PA�<�C�BF1�m���cC"Y�%�|�<Ap�$�����l�!�e%�)�!�D��+��8�)�{� h��O�5�!��V�w%^g.]J����Ь�!򤞷(Ș�:�F6Q�L�i�V!��W9?.xl9�"9$"J���i�@k!���t$�1Zw�� 
9.8s��JZR!�K�l	87��
��
S$jG!��>H�����@[`�T(�0��O5!�$����� ����z!��i|d�K%ƚ����ۚ!�,GJ����$b�t��z!�dY�~������.S��	�)�,^�!�"\����O �p]!��$l!�*y6���(�f}�\�å�4X!��Ǔo�A��őh�"ӂ\�5!��3t�A��OHnM!�Q� =!�$ڀ���P�m�:K�aj�e�5�!�d(|^��(2��"�J���a�!�TfR����w���0C�!�D��`x�ɇ;]���Sm��M�!�@(9NФ\��� �c�_�=4!��ϭ)�	��ۦ1������ќz!�$שƈi�T��c�f�Sl�,!�dUL<\�� �"�T�B�[�A�!��a���6A�Y�99�J.9u!�d
�fK^�5�CS���h�FX{d!�D�Z�QZ�j�1�N��e�\�!�р/��H��a����d�S�!�d��DѬy���
98�T@8�eկ`�!��d+�hI�A�:W� !��]	d!�d���� BS�X�d9�h��BA%1T!�$E�F^�%��t*̴�����o�!�.kD|s��E�T*�����M�#�!��Ml�H�d���8��u��s�!��p4!�0�ƭ˅-ڭ�!�d�!������'���Jq�O��!�D�+{Ҋiz���:hH�YP��M�!�P�Z���W:CeP����\�$�!�� �3�"T#�X�q����S~�A�"O��쇋J<���Q�S	cY�!��"O�x�#G9��� ˨SH�y��"O�q��(�ߐ� ܳy��ŘV"O�tjbW1~l!r�M̜~�`���"O�e�u�X �����X��%�7"O ��GJL$V��)B��R{���F"O6��&AzmDh��1h�d5��"O�a`B
Q��Ў��dh�"O����b[�A�Z��5lF�3c�u@�"O�����5�`|#«Uh��"ODe
��Z4o�F�2J�P��k�"OH���+X����qJ8Lxɖ�'�\�(H�G��V�v��ڕL	�wx*]�`L�:!!�D���O���m�jX��'��}�W�X~�a���ϰh�!�d➴e�ʈ O��y2�}��9�����C�y)bj�68T�}�י>�rdT�nw���'7n�C`G�3>�-�RNV�]����'�L�f�
PhݳE���c��0
@5,k��`V}x�D"�ۗ6H(����*<�+A!,O�DZ�i�^l�/O )�Y�@�*e�Cj�Ԩ��"O�l�!U��lU�V(�Ĉ��x
Ĭ\*�AW�[U�Oܨ:G�֢py�A1f��: ꨡ�'��PӠh�D�25�[2+&>�eδ��eSBT����x�eµeZ���	�0q�����т֐xR�Y�K�����`��F��ma���5L�~��띎\���	�+I"1�f(!.�RK�9{�����HD�{�D�5��D�-�F!�TJ��?�f8i��ʑZ!��;2���&̈́���Დ( �$ԉ';
̓�g�O��E�4MT+G},Ģ����@-��P�OC��y���?+�`�q�b̑Eˢ �����(���R�>IV'�V���']�S�
Yx�16n6D%��S	�'�^ �b� (��ԛ�\�*�bU��^$��"�'�h)@�L�9<V�aBuNԄ?�`��ӓ+�4�*J"}��ů8���s!�S%�\������y���z\Ɣ7��G�D��y�k��-M��ō����h'-E��y©�I�^\��)AXd��$/�y򉝾Csre���@� ��!��*P�yr��$]��`G��9#hR5#���y�%dd��1��L��tI��y'��6O~%Ph5�0�cĥ�yB猕���x�Pm"����y�
�{���p7Ϝ�LNl���i��y��ύ��r%c�D�h���E^�yI�K����H�9K`-�����y��T�)HLx�Ă_3:�$k��G��y��Ʃr$��8��G�+/� ����6�yNо���ʷaƛ���I�]�y�$ޔ[&��w��(C�b�����y�o�)B梨�'��4s\Ȓ�DW�y�#V�G7D��D��*1@����V���ɟ0Vf�����Qkriꅧ�&^���24f]��!���Q	����NQ	�d��L���"�Of��G�Ҝ�1�1O0m���Ωc�f�s��	&��)'�'�4y��$X�n��i�@F	���k�u��چL�V؟����
`3��t��-�Xu87A/�/��( ��;Mx���͘ӎG����iՕ#��ܺ�"OBL2u�ߐ�hY�0��*��|�vT��i~�(ґ>E��SM���t��R�BSjR+�y�#�&s��q"�Zr9j�zH�p?��'�x��5����ϸ'� 0�w�_�L����F`�-�И��o�.�f�y �������S�J��l��bgnt�W`:�O�A�e�1051��i�P3�e���	�5���(d(ʦ,�π \p(p�X�V�vQ��0D�ӗ"O^�9I�P٫��%D�	�_�P`4oƍ�  5�>E���̀D��0y�/	H�dg�y�9;�8���<z�h�gLǝp��'{�x�7�ǜ�Ϙ'Ո�9g���Q�B�f	G�g���'EҔ�eI[�+�@R!D����$𢄍-�I2/�"4[���G�M�@�@� D��RrHW%~(Z�07j^�^%��f!D��
*��XƵ�S*�,�P=[�?O`]���)Ԙ',N$Bp��2�v�{Ua��W��`�'�<���mS%`�.	Ĉ�E2 ��O`UB(Q*X��O>C�^*s��EC�/[�B:�r�8D����ԡS�&|���x�� x��ӯ���31���y��[f�3�	PJ���4�������=)����?�Ŕk� ��j��#�A�d�P-q�|QäN+����䌠EZ�$�0 �&�@%.�3�џ`!�Ãz�l�+%��D���!"����bԻhS�ppЭB��yGJ�(@�=���iS��X�lͲ��D�Cx�qᢃ]���)�'}����^+F�y���~����2��#ׄ��[���[��R�
��x	��>��bC�Hzu�J~�=�cAGlv��p�Q�( �ACw�M��؀A��r��T�ci�b��	�4珴U��x�nδ=�rj��Hq�D{�k1OP!�дSd�Z!�	^�n����	,C�Bu�ժ�q&�V���d/�����b9ia�@�+�-��JI����'\T�G�;8�D"�T�8,����Orԩ���DsZ��A�/�|���gFK�1�~�b�/�=�x<C�N�MQܼ(�"O��B.���A����8@���%8O*��u�4��C���~�}z!G(?ق�Z����C������b��H�<���L�AnRE͜"l�ʝ�2$�m~j�@�ʹC�%�#�0<�Ԭ�!��p��p���y��a��4�����c���Y���'jr�5���]:׀P��v�(B�ɇ%�`x����kg�X�Hp�>I���T�vĐV�)�J���6+_wm�Uѥ�٬u�!�$[�q�8�2D��AL1�$�Q�1��I 
 B��!�)ҧ6	RU���Ş�⁈P ��g��a��xV4p4�N�?�.����7-J�8�ȓW�<p��"M��0��܅M@\��?��I+0�\q�@����������),���i�U�>z�p�"O���i@�sUP�!��K%~�J��g%���@����?�H��	f����M�t0�4IV�u�NB�	�+�f5���?�bԚ�F�9,�nQ���",�"h�ˆ,iN��
˓%����ص�x-͘�G恆�	=\��mc��P�}��<�CN�\�����Iѕ��A�v�J+E����MCF��B-��*������9c&$��=Q $3rA"��_l��@Q����Q�%8�0x�KX�Frd��&�y�L֖E>Z�1c��2IT���ⓕ�|Q9DC�U?�`��O:M��Y��J-�1[�E �
H?Vl�$�9� ���FO���C.�a�u8�k^
@j��t/
:���f^�6�쭄�		P��1�шL���A�F�"[����Da��Pd�0��Ҡͅ�F�(��w猕}-��@7�\�;������OH<�Toi-FaQ�A�Y^NX�'[ly�M�he	1�o�&�k3���R]��~�� L=�d��b�(!1�c�m�<�m�&ҍ��HW+'��16��^լeJ���^�|�Zҁ�f)z$?�RJ>��eH:P8�������8*���B��$��%I9D�>[$�@P����eI�s�t #4�1G l�m�<_�PD��	iHR08SG9l0�l3�ɏ5�v�?Y� �[���8�iW�W�l�ZWkJ�,m�D��1#�B�I�W<�D E=o~ވZ��3l�������}�ҧ(�ܤ�7b�4�@��w�L�8�𤢶"O.��,�% �@�z���9'�@d�Cl�]�$A,pF����G8���X�fJ�k\Ol���*� 	����a�d@-�#?�~ ��?+��]+��7��8���$Z��� �%�a� ���<i�?�s��:�h#�)"��ۑi�|B��;�=���Q�!�� � cD$;]<!*6$܎ ](t�uZ�|���ٓv7�h��>E�DdM?R����$��z����yb�I�
9Xa�����ʌ����	��')����{�ϸ'@�C�k�.�J�q4+�	�b��pE�#`cW��ViD�nnr�	7�/h:n-��+%�O4zrE�.:b�`�˒=g��۲�IK���1#iI/I�O�@�Rh�)������N	��	�'阄��&�W�B$�M�FP���+O0T�3�Q�5KI�J��|*�n����]�A�/Ț�A�gL�<�E�E4TxT� ��+1d��fØ���1l��6CK�g�V�\:B��	cӒ���.�-���+]*����Q:�\52@Ȝl�������K�C��m��HR6�l��cb	0M��C�	�6Ŋ��B��B0Ε�e��C�	�lH�S���r�Lh@��$0΀C�	������:���Dc�O��C��W�0h�hN�|�zIP��$�C䉳,w���3dٶz`���* DΈC�ɧ/�2	ڲk��D���E�$�nC䉦(���k��9�b��S��j�BC�	�2G��ЁM�D����1�ؚ)�&C�I(��M�2y��;W!��c��C�	B(�{���3��`�WV�V��B�	�?'�y�5f�A$�0s�צ�B�	�zy�JP�H�v�F�*��O��C�I�P`���5ifh��*� NƮC��4RP��#憇�8J�T)ޞ�fC䉆K��m���F�`l;�eS�0fC䉙j�T:�*�>e|�٫���tC�ɐ~D�#ufE�SԜ��&2��C�I�oz���#� ��Pv'�9�C�I<��t[�ۗ3���eI�m|C��1k/�DI`集(}Ms�	\`C�&f2ek"*T&v�=�U� �,BC�ɛ>Kj�P��.�bϺA	
�i�"OBĂV�,<� ��w�'u��MU"O<,`g#�-��5�g,O�L���"O>�(GH"y��xsg�?J��d��"OV9Ơ��s�d4���tJYȇ"O|�寞�^=q��W$�W"O>�ô
�
Q��ѽ"7ƹ9�"O�]�v �9��c�V8Iy�"O�{�פz�\�ه�!Z��2"O��Q�RafؔiQ�/�����*(���&A���S�GJ��ɄAu\Hs��I9D�P��^�|�s��4�z��	�D��jh�c�'^����%CFRR�B��2CY�Xꅑ>�I�d��X�ç N�h�⇩#=pAy�A4|���<q�+�����O-&��BӁB��рh[�.%�U�Ot=�!1�)§C�ҵ�u�M�RGL�RrO�+x;�͓[�� #���)��zcD���^4f��(�1�!*'���'f�* �Ak暟��ӱ<g��RoӉ!��� �m��/:�c曱*����^>��)�3%bҍ�Q��,i�+�;]��=[2��$P´i�v��}�S�$님G� �"95\(��T���H��$�>[)󤒙N����$[�b>�I�]2N� �,��&�����d������<a"��\��S�O� ��AK��؁f�%�����'[��ԟ�T�T�иz�$�r$��5��/v�p�vH��ا���C�eԈ�1���I$'+�TҔH߹��'�6!����<8�V
2Z��ya�<��ʓ(����9
f���4H�~J�'\l��r��T�������3Y�����)f������	e�>������}(�;4�}��iBFV�W�֜ї� �$v������Z
���(Vj����K�n�y�*a�I����2����0|�%.��-S�O�;!r޵��d�wy�l��E��qǖ|���Ef���A�M��	�TB�N�>2�b_��M���|���5٤�@Tc۽��������Uˀm��D4�'�a�� �������0�|7�-f�� ��9O�'
d����qO�'G���*�5�@�qd��&:�х�Bn�&�U�L"&ԇ�Va�ȓ.��+�;H�*�*'�r��ȓ=Q���!�^��Y��
-P�ąȓ���dT�E7���IO=����"U��"�f��g:te�a�ZmBd�ȓ}��4	�&+�t��B�E�T`�y�ȓ
���	��D@��J��(��B]�<�OH�.�,�c�'׭Ss��4�B�<Y5��o��t�.,p*��$BB�<�v�9�U���7L��G�Z!�Q�l@0l�t$ޮL�J) ���o�!�$Z-\tpؑ���
@I=:�!�6�@l�Q�H�ڍc�!�ܶXJA�F�z�>\q�+G�!��K�5�kL�<���3 �!��;�h�����;�p��UNW'�!���!le��Ѡ�
�6�D�Pv���fh!��AH��J5�O�p��u���!�$\�I&0�tLK'�x��#H��B_!�dK�q6F�p�N�Y+���=	l!�L
���'JS$}|\	3%O!M2!��?�>1G�ro�#uD��!�_�F9I��Bݡc��'#Y�m�!�D/o�����*C�nV�E�W��.W�!�N5!<�Qðl(څ�غf�!�I$Bi�a�B�$~z��@�K�!��]6�[��=V � �c d�!���%� ���٧R��d�A�rZ!�$��	z���`�B%d��T�a 'l4!�6-���㊚l�d��j19�!��!�P��VEB.,�@�K�Z0.w!�D^x���
D	J��퓰Dze!��ݤ
dP*ǁ1*���YFE��wW!��k���h��\�� �["̯�!�d�K���I��,�a�X8=L!�$���0)�"dب���Z�A�0!�S^�\����ڞX"��ٲOI!�@�5S�q!䁕�7�B(ʲ$�:5�!��8��ӂ@��>���q����>�!�$�spZ�S��:�LikX"c?!�$M�l��dE�=Okb(a���<<!�N!k�����a�G�J`ZsI߸*�!�D�t�p���>jAPm�6�J+m�!���X}���N� $�0�z~!��xW��2�Gβ=�
�b4͍�lL!�I7[tP�"�7Pv5�l2DN!��O X��l�%&kJ!���L�-!�ď�":��#�Ɲs��0�̘/(c!򤉥�H�c���1�pQ� ��wd!��P�Tx��̓�Z���S"�H!�$�5:_t�;cĒ?f��ٱ��I�2�!��I��ޑ���_���G2�!���V������FkĜ�k�H�'_!�D�2��yr��#���#H��xE!�D;�J��
I�bt�I:EGD2r:!��_�ڐ�TM+cs�͡7�Ή6!�H>x�͚t}�0��B�ێW!��TbB�Әs����W
[�&!��Q`d�
�h�)'��t[k��*%!�d�&��CF �� ��
�3"!��3	I&g&��f�z�
BH��6!��E�	�f�2��5(�D �FFK�dP!�� "�c@ȟ6%��A�
F�4h"���"O>���-]Ժ`�0(�6h���[�"Oޘ3a �&~^Q���@�i%�:B"Ol�K��\�l3����G�`�R""OJ��ć��f�JM3\���KW"O^��B�
 � S�M��)��"O|9��N��oh�H�$��<j��Rg"OZdb��M�b��H�B�b�Q"O��[�)rSTi�@��BO+�O?D�d��i�0nn�� NM\	4�E�;D����2���D�J-| ��SQ ;D���X�	�,=J��F&���g8D�$C�NDp�����5o�p��m5T�l�􀚳��c�I�i��a��"O��ѓd˼G7Nԓ�c@�t�Ԑ{q"O��K�'I��\ss�ԸYu����"O�"��κ��g�I)h�A�v"O�h��<H�ʀʃH�G��<h`"O�A�t��q����ҦD�W���pr"O�9��(�l2̈���	�`$�E"O~P���$�(\
7�k�u�"O�����cx0��G�$n �}��"O�D�BW�
�0u���[�����"O���ō��i� �3�\��"O�P���!J�q���`��y�"OX��T���+�0�4()%�Lpq�"O���+=E�PIW%H�l-�DS"Od�0���V�f��IY�G+h!��"O>����� I��  �jֱrp��"O�Kj�;sO�!��o@*-���"OHA�֭ӭP�4c��!8,Z}Z�"O�;�͝0$��ع5�8&���"O�h��M7K�vQq���@��17"OL}�� �-F�+�✢?����"O��"��}�%{V��G�ΐ��"O\���.f$d(�ЏC�,Ţ� "O�}Ӈ,X�L5����Z� ��Di�"O���"�	�݋p ��2�6"O��P@�B  d����X���h!"O� ��ۉa�����Z��dyل"O����[�,�@emM�	"��"O�d��m�L��Qx��˼-���"O6	�s�єQ�b��bD�1Tw�M�"OV��b�"���9#c٥=n�Z2"OD�;#a�"lȥӒ��#*�iI�"Oh����<2�`� ���0xT��D"O0�ÇJi��=�DD۝cl��Ic"O��2g�Y?���@!>T"��"O6��d�ɵ%�J��!-���(&"O�P��K�c �� ,98�*�("O�D�`��Kz�$s��3l�hي�"O
iq�G�V$|Ļ�.�z�n���"O��	p�,fl"��V�0Yy��2"O�4[ss��Ȩ" a�x"OH ;�,=X��ـlGH�9;�"O �Rn�%kiB�C��GA�dW"ONX;�KLv���B��d;&T�B"OlDhF��(^����Q�2"Bx�"Oh�D #L�4!�e���\z��"O�����{� i�^,U`2�P�"O��Cm�>{��Sg`�3W�i��"O�5x6	��hh��Y��O���"O�K�eU�c&ظ�F�ʦI(�\�"O6��A�w~n��P暷x< �U"O� ���
ܗuAh�ѶB��z?F1A�"O�!6���r���ӧZ|�0q�u"O�� t�Ă�	'�W�>��p�"O�`�%�+7�ѩ&J��q"O���k�?'z��.��$K�"O`���46h`A���X�C�"O,��@��(����ьM� �Y�"O�%�#K�CX�	$L�9Q��챀"Ox�c��D��bPHF3B[v���"OI0���v8��ZI���9��T�<�'�_���:��  ���J
R�<с��D�q1ȏm���R�K�<IУH1,� �I����0�	P��a�<��@-[�T��1���&u)3�`�<93 ������'�V|!�g^�<i5�M %ڌA*	3��XAh�S�<�c�\�NoT��@,[#�����Z�<q���$=[�����Ћ.�l��T�<��D�Jώ� ��C���񣤚E�<!�A Z�h���ۅ_i�(!�m�\�<q4�@"KY`�`�lo� �e�M�<!�^>9�z0��<T�TRQ�<ن�ˌ6�l���ϊy���q�@J�<I�hV�*;�e�v�τS5��j�mo�<ULG#WĂ�� �x�FD��n�<IǬؼ~`J�C��K�App�@LTm�<9G��<H�bk
"ttra`���R�<I�)��=�Le��mךh}�Ț��N�<Q�HZ�6#n��e�g���F�b�<�aiH�+NpѸ��Q����᫈[�<aqo"R:����,!Z�� ��	a�<1��y��`1'O!S���k�Y�<9c���$@<$�C��!Pd!���R�<���H$�@#���_�݊��K�<�D��,ֺ���(�$�}��O�<��%șM����Kь"+ܽ�wK��<���_)kv��$'��c �����s�<2!�/qް�cvLHr)ьHu�<���VE�j�;�l�xk\���mBo�<�%�R���E��E<M�$ʕ(�R�<���׉}M�jr���x����GJQ�<9��ׄc�R�sB/�X�jd&f�<�˟�?���9�	խI��p�!Ub�<�U(�0J0�%�(T\b�DS�<���K!
{���	??u:4"�"�z�<��OW�C$�Zt;w<�=1Bn�v�<	�� ;�@�ꦆM;UQ�����Yr�<Q�A��$ٰ�9qc@��t��pAB�I�}a����.C�I�]����Yj�C��2w80h��`T�ڕ��{��p�',X$j`L�E5�@�U햗o�N �	�'�ڬ:f	L�͊�Q�Вmz�	�'�t1�RkU�d�����.;`����'�@ ��eT%g+�)*�O�"]�����'�*�j�ł�l@@���	`���
�'Ԕ��d�qb(9AD�ӒS0����'#�Bf/N+4[\@J3���ș��'�0��dДH�����	\�ܔ9��'PR����ǯh�,���������0�y�K�5��$� A��eL԰�y��%q� ��lC�g��5b�<�y" ��D&t�{ �b}�$����y�@βk�bB��DmJ!ى�y҉�3Eap��aȜ������_>�y
� �XHv+G� DJe �*N�ŋ�"O���q�=Ok�Ё��]�fc^�rS"O��9C�_������
�gVP�w"O�Ii G�Z/dl�`��39Z��"Od�0�GR%�%��?_��4�F"Op�n^"(���+AE��A��!�"O�� r���4��1���զ�+%�y��'\5c׫�'bj�p���y"�5d�ÏN�	SV�)����yr��@ @  � ������4�Ms�:(�Fs&�MG�O�=Ғ�_��E{�,@�v��Pi�"x��b1�4W� 0cG.MF(Q?9ڂ��i��_qYp(��m��'2.��,Oaɱ�7	+�̰�s�0�t"R&�$�y���kTr�;D�T�¥�'4�`ic!ӣ��0���4D�T(U �;ҪX���>Ā�#��4D��Z2��z�ԉR�o����{tL1D���℆z0i�!���*��tq�	;D�HC�H��
ѲxI�.�f�LxS>D�Dx��Q.��-[����C?D���p�W� ��'�Aey�����=D�P{2��k{>|�`Ք�X��=D�@{OG~d�d�2�� ���:D��Qd���^�@z��6X���p�-D���Gω8�Mc�T�Nj�Pd�7D��X���%3����nT�d���t�1D��x��� �}�@��O}�L�F�4D���G�k�0�hrJ��C�N�;��$D���'�\#�6Z0��'"D�|��!ˎz(F@֍A,t��k�!�y2�O�R��Vy�����M�8�y�m\���|bǂЏhRR��/��yb��	7gh���H[]��
�J2�y�`���P-�TX%㗆�y���5���R����xL�H�3�ׅ�y2+L�}��Q����j�p�������y���.&	�IX�
\h}N�R�,�yrF	�j��u`4C���y�`��䮴9B���C>!Y2C�:�y�C�]���Y�.G��98�e�0�y��8M���HWP�t}{�
��y"d\�s���2����]�� 1eA��y�Ȉ�*����P�T��e�  �y���z���HJ�y��Ņ�y��[X��O
	) y�E#�y�Ǖ� *��Ug�Y����B��y¢3����P��Q��H��y
� ��P��N�R<��P��Y�ltm�R"OB���A+=�e[G�T=n´�"O ثaJE		�L����@b��q�"O^��p�ٛ�H�[B��#k�7�$D����T$'Ѽ�p��Y7L���-D�����T&X�ҥV'/���!�*D�l ��*	�Ȅ����\F�!;tc)D���� ,P�a��� G�b��(D� �h��,��l�Vjԁ{�dg,D�\GNɗ)A��@�F�<�ҹh3�)D�TP�@��@��ŕ�b����3D�`�bLH�|&vx`�f�P�R�CE0D�HK�Ý�GĽ�1�ؚdB��AL.D�
���!a�
�k��sJ��B�ɭG�����@�+䰭��`ʄ|i(B�I	V0ب[0�[6��xr	�n��C䉓,�0"0�]H���H��	��C䉍B���ݮH�d���y��B��V�8Li�N�$_q�%B� D�J�B�	'H���#���h��1y�]\"�B�I�jp��R�����"�ڭ5g�B�	8q&;��^�������Q�$B�ɄJ
<�H��L��$3���C�I�\:��/�18�<�r�Ĳ!l C�I-?�ndx�(Q,-ltX��BB�,B��D�vp�#f�4Ԋ,p��C��KT�0�� 7ۆ�sR�-mg�C�	/Ft�Rg��4��jPf0@l�C��)_����!��|aI� �#2��B�I�)
��C���`��c�6�B�I#>|@�p��_c��#F �4\�B���JG�ӵbv���bP�z��x�
�'?Nl�G�نh� �J4�#���	�'O����8���SO G>*���'��s�h�yJ��sS�1;i�}"�'H>d��C��?�p�
�} ��'�	Sr��\�6���*e>��	�'�������Q��ʤ&��m��'`D`:a�M�Z�,CA�C P=J���'3b�KF�M8A(�Q���0I�fu��'�Ԅ
��4#�D
Ǝάl_:��'��$B���=o�T��+ aR�i�'jR�1AI�#�\���X�Y�'��uC�!�[d�-���@�V�Z���'�t80eBW<�@��S�M��M#�'�m	��?,���6C֥Bs�x��'u:4sңA�/t���M�>�j���'N�sAK+1�ix5$�(��$�
�'���i�J:*����E[���݁�'�٫#���d�@�b�4m0,��'��9���	�0���1A㕑vt`��'�ty6��]a��2gDߟj�A
�'~��*�Յ\�[���aw�!��&��Sc�8?%ܰ��m�PV���r��h��M师uʜ�X� a��st` À雼"�t*��/T&���Z�fd�#kB)}v��)�g �DZ�q��lRv r e�|���Q���ȓ�^����+1}���"cN6CwzŇ�&&@8��c�j�P��.g�I��|�<��n�Dp��T�����ȓ}�p�2�S�Y+bqP��$�ȓvj�E���_�Q���"��1�ȓ~d,	��T�12=�C���#p`���S�? ��	T�ե �vh��� P��r"O�l�t�/��Qbjٔ�(xU"O��s@.� 0�H�1�(��g��J"O��3"�7�]X6ϱB�F�3F"O@l�jY"5˲1#�Asy��"Otۡ.4T�s�J}���"O�����(���k�6��"O,P�Ձ8@_�� �\�f���D"O�m�� �&�� �3Q8#e���"ODh���&�hՁC 1����"O��J����[!V-�� \#��+B"O��k��L�M@�Y`.�&E�Pe"O���RmS��Г���,�c"O]���%|V�<��b�N�8�"O~0��/L)�t�pp�ŗu�d`�"O��S퉧{����f�^<-��+�"O0�B�J�x=���JV�B����"O���JhP����5v��1�"O� �5BF�2=��H��k���"O~Iڡ�s����-�3tߦ��"OF�;G���.�l��w�_";����"Oi�14z`f݁�DU�D���:�"OH�BG�T�/\��W�F���w"O,�CZ�j9 �8�˃�l,H�"O��@}���� ޴P�(�7"O�}���4Q�8v��o��U	C"O���&@�#]x rh@��8�H"O�1�D�m,�@1� ���]@V"Oj$PEB�1��p���<{�eS`"OP@���b��!pÈK8x��5;�'y� ��0�+�τJ.��'��t�R�ɼCb�(I���;<�v���'�t0R�)"ul�Z����4� �R�'�4��c���.�`�^9�j`�	�'��[!o������6!#�'�Z@R�M,5���beHˇT��R�'�T�0g%IE��Бt���V؎��	�'Ԋ�S�ƀ{lV�@t�G;N�*�'z�)��fڋl���@朚7	����'K�Tz��_�T�$)	�X>6�TH��'�����o�*T9�	j&����5��'q���Cͦ<+Α!}���b�'�ja�Tϗ�Y�bԆB v �qK�'�Τ pc
����R�w�b�9�'�:%�֮�Rs$(�a�qP晇�_��TK�E��|�@B�]|�$�ȓb�ЩhR! =e��b��5bC�8@��,�ЮO?2�$=�v��5(��C�;h�8�f��<I��,%)�>_�C��9Waxlz��R�HΕ�v��"O�=	v� �i�r���-��'�p��"O�1R����X�6�R(�"O U�e�0E��QJ���'���"O����嗎t��LᑊȖ7�8�)"O�]� ʛ��c�鉍tsN<�E"O��A��zO�S�ǃAX���f"O���p*�"q�j��B��6AF��"O��*�E��m���EO1*5:�!"Ot56m���Q�.  x�yt"O������ `V\[@,�"O@�����UR�hc��@jա�"O����e�0B�v����E�5���5"O�PH#-M�)�<��*���B,��"O����Ye��a�&��Lq:s"O� ���h��z� ��"��9wR�i["O��:�J¶������!t7hp��"O���	�<�v bd�Ȃk���"O^�˃��yt䈦d̓O���0�"O���Sk�0m�4�n�U�4�� "O��Yѡ޸@{.��g��1(�@a�"O
�����>W`����Y���0"O^��q��Yh�����8�ŀO�<��b�4ʰH�j�*O�����]P�<	D!J�2"��aMϤj�����`JI�<1F�ܮ�D��fQ#d�����}�<! �)QiV��dZ�`�@(��gP}�<٤�O���I���!���@0�_�<�&o˚X�b��rYC�ƨ `�<�#l��n��O5??hp�BY�<��L,gļ`��N1`��U���L�<Q�;6��<��ٸ�6��n[E�<�	F�x�z2ٛ:���`E�<!�Kұ���a��1;���ȜG�<qr��Y?�U�����i��\@�<qE���uPG�ǥ&�)��dTF�<� = o� 3#QI^J<�ȓ1�nyx��v�B��N�:^`��L����v ��g�Ή�3�F�,�%��W�P�3'g���J�D��>MjȆȓW%.[�l��`9<��u�M耆ȓn�A��aŞ�9���y#r�ȓK^�	��˶u�����JJ�ZE���ȓM˪��&��.�������lzn�ȓst�0{�	T�c��a�I!��%�ȓjm�Ĳ2`��k�x���Z�[j,8�ȓL��H�d�ߚ6������ۙL�nȇ�Iy�FK�1Szh�q%�2ڬ�ȓQ"i@�J�
�2�x��ʖJ����ȓ����s��..��2#�_�{Ld���/Y���	C�PЪ�m�"�4 ��8�\�� @�?+��d�dBG�"9H�z�;D��1��P�c��U�E=%<�1�9D�����E�+��X&��L:D�pX�n����a���9���q�*D�,��A�0����Ԯm���#)D�y���
6���H�w�`4��O%D��* �N���Ҥ-|�6��ҥ!D�h�1��?��H1��
�N�$�8u3D�T��̒NzƸQ_�$�T4W��C�I=[�x-5�։j"�=z���p"O�8R�ͼ
J��L7(��"Op�*�F	T��u��悖$:��"�"O�;�E�N4ά��/�O�F�G"O�!�#�V�&9vL����&m�hb�"O`��@&E=*Q҂c�b���Z&"O� \%�c��*"�%�a4>�@e+�"O�I���p����p�jL�g"O�0��._�;���礐�$.�y�"O��7˘J�m�D��J6��""O�L�h΁���7�7?|�"�"O�b&�wP����� 8�DY�"OV<Ɇ�\5`����P���r1"O��THݵj����Ј3�N��"O^-;�G�&�<��û&��!��"Oac�oG�J���&�
|�:�k�"O�mÁNY)Q �H�\ 3�2e�"OP%ipg
q���2$ڕW��=A"O�@A���8Ed	VC�f�}J�"O�AQp���#�СT%qH<S�"OrS�T��6����TZb	;�"O����֙_���y��1I����"O�|��5�6�h&	�,3�a)P"O�(r�@As��`��Q)�Y��"OJ��BdZ�7Z�L��o��>��0�"O�l�%�:t��9���ƀ`�f�#"O���ƣԍB�0��Եa�:��v"Ot,@w�O�L�$I	��
$�dL�@"O�zԫK�[f�����B�_�~��"O����i9L��0z&��,���Kq"OP}�+	�` ]`�O�&H�t��"O4)ɱ�֓*^�	����j+>�au"O�x�ՎTBT�s4�޺o8`q"O���Β�d�����#48"�z"OT#b]1L�^�����/d2@���"O�!�!� ���k��QRn�B�"Or�
�Nʖ>���o�&�Q�"O�%B�!S@��A��a)+�a �"O�� ��9��l���T�OR-��"O�%!�!��T�*幕���oZ��SS"O�Pᦩ�|"Hi�A�.�`D�W"O��q3�V����U���r�=�5"O��RN�m������'mEP�S�"O��`�W�S�A���R,�吳"O$���G0.�n� 1f�4v���"O�i�wE�>��b;<����V"O��;��ˊt��W�#~b�:w"O�2�(T�s�P s�E�5z:Ĺ6"O�� ®�L|�,WG��Փ�"O���G   ��     �  B  �  m*  �5  yA  	M  �X  ~d  7n  �w  ��  ͋  g�  ��  �  o�  ��  ��  b�  ��  '�  ��  ��  '�  k�  ��   �  B�  ��    �
 � � �" �* z1 (: B J OP �V oZ  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p���hO�>U2��F1C4ӡ%B�>��eW�%D�����9]����"8�
mS�#D�th���*��6��4��$#D�\��2~F��u
�!.���sA D����ýe������[�<�����?D�@�w%��&�f�SS%D��8a!�(D�HY&N�1V�ȥ���V&D�A�`!�	�#��yr�C>s|D劥o^2;#y�Qk��Px�K�{�T�:���(8��+�#$����>iS�'lO�m���KTѐsF�W�ճ��'�铤�$ũN���rć:5�@3"��)rm!�P-s�h3eH�r�xb⪙�j�!�䈾�Bl�*ݎzp��a2c�1Y�!��8$�N9�%�D#f?��
�#��y�!�$R*l���2�Ɵ�1���8cǈV!���+ D�
�dV�e"⼐Fip!�$�8p�,�7�֐:$��`H�;�!��vM��­�@�0��/Et!�ĚYゼY@!҃&���K�f��l�!�� ,.�T�%rd$�4�]<~!�䛱���kah�f\삑�M<+`!���8�e��2G,%s�FS�gI!�� ~��d�)b4��ci��.�2�"O�a�L�I��=@Dg�0��TP"O�1���F�nؘA�5^�
���*O��(�NB4)�xt�θNy�:	��Ms�O�ݒ��hҊ�Q Ў!�ZM�"O�������@K�ux6Q���{�O˦�l�+E�x�Q�đ2 Na�	�'٬D9e��91��p�X$>��a��'�б�Q����i�&D ;? $��'͢\"�b�^�@!`�A70uش�~"�Pc8�@SD�?(31���T�j	���?\OB���$�`s8�Xt�����I�f�!�D_�)��#��R8�$=[���F��'Mў�>]@EÜ� ��9z#Ï1�̐ .?D�X�h�%;��hK�ɚk���F D�*$J�)" � I�3*�q'�9D�L��l�K�d<�7�1<�5xү3D��q3O��%pafӀ)R��p�/D���f��J������Ib"���-D�L� R.أ#�	�D�*u�7@+D��8R&R�2���B*^,�Tk�k5D���3
L0�,��f�1(��xC��t��=E�ܴe����Q�0�Z�(�N˖|���ȓ[��}(�h�0"��_�Y �0��j��s&�O @�B�I���@p�P���F~���`F��%�^�7��H�ӳ�y��9P�����:Dql9�F���y��N�'�4[�IE�%ߘ��E�̥�y" h�^�ڇ��5�-�'�yR	 ����P�S?`*y�����ySc8P�{��`���'��y"�U�S$�R�$b��z�K&�y��X�rm��"��\}&�I� +�y�)>1��E���O�H���؟Ǹ'�ў���a"QF�D�A$���;�"O����7��<�2��5c,dts�~����BAH�8�YPg�rhR����y�$�ޘcF�U�n���^��?qQ)=�ONa����ph6��F좱pe"O�e�/���Ukֶc�I��"O���茰+�j|����vp�d4�S��z��X�W {E4�(�&�DhC��2z��iH4�l%��7|�\C�	l��2�利@��MR���z'HC�I�)r�(z���$㠝c��+�FC�	�L��<�����Wl-s�D�$2C�I�]��%��� �X!�BE��ybgH�(�L�g�� �&�Prm����d*�S�O�<��� ({��Ar&�T
#��t`
�'�<M2�g��h5�����	�'�0`!�(��&��`ժ���� 	�'%���7�L�RE�Q$FB��"�'��h�Wl�B��	�qO�+K��ea�'O��Ȱ�H�j"�y��W�>��z���'*fՉ�Q*y������gӄq�'6Ȍa��5��Y2nϤTTh�8��Dp�ޣ}�qb��T�6(��Ob��u.P^�<a!��Vp��ᨕIF��S�GbK$P��O?��B��*h�w�ۿm U�6(Y!�\s����?s��!��$�����>��M�+�����*@�Rm�#�e�<�b�5q�������1�|0'"O4t�2�մer2�/�(i���"O������<4}B���M��!C����2<O� ʅ���^#7
��bQ��];bOx�����&PP�,[��=��( �� $���`8��2����7Z�����>+��;W�=�O��A�'^�}��(�d�X7��<wR�52��HO���&��&X+�c"�r��$I�"OJ��`S�l�1O�
���W<O��=E�t�܉k�Z(ˉX��0Bd	�:�y�: +d��)ɰ\�`�� )T���Cݟ̇���	7G�I�<}���������<IR.��h1����%"�&���n�p�<�u��0Am���4�D�e���yĊ�e�<�W�J�I%�a���
BRV�١AF_�<aTE�TԤ)���=0�U!7�x�F{��逯L`�!#$�˯[�&e��	�"|�B�	j��e��޳�-SET��ɧI��I��~��hO����Ǆ�$L�rs�<8oڅX�'�d��'�4��b�d0Q.Y�f��n�W������m� `�z�nZydN�V��0=A7�%��$o��<Rŕ�,��K�肍M��듚p?���	c����e�E�mhb`а��}X�ԦO�<q��ѷa�pz�X�L���"O<p��C�	R���y�-*g�|B�'��O�c���Tyƚ����Z4�����0D�x#� ��@�:��������d1D��!�[����g��r%p%��/D�� ����7x���ʕ3Y����&-�	��Q��O��좷��'>i�`��o"��	�'
�A4i_�f�\ѓiD�3L�ّ�A,ʓ�h�����t��|f)*>z���t+�m�!�:�1gI�>} e����)�Op��r옺i��h�&ԠXw
"O�p�A/EJ��E&��Wg�-i"O8���R A�	&e��d?N$	0"O��C	qȜ8p�!1`�V"OlUAR �;I����.	�(h��"O6�$�ܻZqd8S4�L(��e�F"Oڥ"`��?bH����t�(5�s"Oй�&ǝ5n$�`vkA�"O2�Q�!�Z�|�o>1���"O� �r�E�1ಸ��͔�/�1�"O`,b�m؜��H�&��8�`��|M��jȞU�ƍ���Ǿ^o�8�ȓRBL�j��@>A>qKv�N�pńȓP�0Z��E�
C�s��!9����ȓ�Tڰ�š<����s�T7R���ȓ-ъ�J0�O,B4^�#�a0|�ڴ�ȓ5� �+�!;ЌS0e��Smf���G�\���
U���dO��&�h%�ȓS�Pe�4DTJ�Ve����*p��m�ȓa@�����[��q��G)�,��ȓSIl��+m{B�ѳ���H
�ԇȓm*�U�#�>;�`p��S�y(�������Q@M��}��-S%ƻ'*Ra�ȓt8����������P�>� ����@�A�A�7#O�S7D��+	���JR᳢G@q`�[��\B��ȓR��;�n�iP��J�:{ņ�?x$I�6	E���L�ES�2.���ȓk�`��3Oĉ�7G�p�4Q�ȓlA���Mլ9�ɳB���$4l��l�*��T B�Rf�P�̇+D�$Ņȓ[z�akFk�7tv��C޲C4|�ȓZ��5��^;d��;A��+��|�ȓ���G��%Lժ���[vhɅ�S�? ,�T��5M�<���"8=�"O���Aٓ8.�ᡧ�7B ���"O�%�X�F�+��B�/�F"O�T� �/f��\u`�89��Q"O��(q��uJ~�	6k��&���0�'�B�'U��'�R�'�b�'���'arP�$@�[��9�,�95����'C��''�'�2�'NB�'���'��lX7F����ȣ��ͷn��H��'+��'���'�R�'���'���'�ik��4+*��'C�|/8DF�'���'���'�r�'���'%��'�t��I��[���LV�+-�?A���?q��?q��?!��?y���?q��ؽ�����K�MX�O'�?Q���?����?����?����?)��?���N���p$̂�s�:��D���?����?����?����?����?q���?�B��*�~�i��Z+Z�Ő�����?9��?A��?����?9���?!���?�S�F�)�d9�C�ab��A�����?����?q��?���?1���?���?�0E��g��A�Q]0,-p̙q�� �?9���?����?A���?��?���?��!3,KHI�4��/M.������4�?9���?	��?���?A��?���?I��=�X���R�;rr�$E���?y���?a���?q��?����?����?	P��)n��LS�ĕ5>F���6)E��?���?9��?A��?���aG�6�'n�x.�3��|��p��@�-8���?�*O1��	��M�#�?q������¦Fr��,/`,4��'�6m0�i>�	��p�v��.E����w��`Ǐ�����-��5$���';��đ>�R�ӂdY��N��Tf̓�?�*Oj�}�0�^.8�����֘{78�R7m̋H��$�'��'�Hnz�5�Т_v�x�ĉe�n����Bӟ��I�<A�O1�����<1.� ��Y���ؑ���<��'^��D��hO���O֡� Aհ_���xZ9��2uʑ�<Y-OX�O.aoZ�,2b�4A�DZָ�b�뜂&S^Bo S��Z �Iݟ����<�O�4c@o��d�lS�_�W�d\ ��	�6�>��P�>�'Tl������dTC���i��
����]
�,i!Z���'��9O��Ђ/�?X�ań�.�Xh�:O��m?Ϛ�3|�V�4�8B�` �j���H aDc��R�9O���Ol���2�6�Ot���J� Ҹ;��I�&˔n!Z�(�B��}�"�OX�S�g̓W�� S�
*��r]
,n(�'h�7͟Z(��D�O��D*�Sxê�q`l�8#�jyxG&�	 �H��ODm���MC0�x��d.Ёx
z�h˕��\�f!P�:�p�B)A�7�剄@��R�u��|BR�T�e�O�m��}K�/D�
jK	�*Da|�a�}V$�O�t���^�l}v�k���9|�Tu�p��O��lZN�u���pnZ�M�It�4���Wt�L](��H9XZ�K>��R�1��^�S�ߙxr�	g�V�"P`#	�0��Oe�����3g^���W�=F��peC�TRj(��ϟp�	�M��AM�dBg�t�O4����՛@2DmJ�+�
'
�:�!#�$�O��4���3�''���4=b�G	�Y�����k�iM�A�"�P#|��IO��Py��d�/Rʦ�:�A��pd	%�� N��,�ܴ9	X,���?�����	T l�
l(#�
$1n����l�62������d�O��� ��?p͚���-Z�͊'+vi[����YP*�ş�����D�i?QI>!g�S\:�\��FU�C"�L�1�?I���?����?�|J.O�5mZ�[��DC.0A�IGA��@$ND_܆�$�Oڍn�F�/��I�M�N9M�ea@AE�S�d�	O�i�Ȅ��%3��œ@X^\0�'w���B�N�2�c��H-HјV��	ܼ����D�Ol���O��$�O��D�|�D(��r#.���̕c���u�ˎT��V�G P�I�t&?5�	�Mϻt3�E�ǋ�^x���Y�1��H"�i��6-�g�)�}���'������ wP ��ֆK���ٙ'L�A��&C?�N>q+O��C���Щl�6�i �O@�̄�I1�MK�d�?����?!Sb�"7��+�蘔)�.��@?��'� ��?)���J<�s��[�x�0�ȇm��)�'6������1C�t�E?���v��ْd�E1=�����������?���?���h�����|��ֆ�+��`�'eŦ]���d��e��۟��	��Mc���4���Y�Zφ�j��� AV��g��q�d�5�4A�����?X�Iퟴ���\�P	��B>9�,�W#T�x���ȓl�)a��O����O��xcaE�7�|K�-�JiP��0&i�n�r�'""�I[�p�P�����l	�@Ґ�'%�6�Ц��I<�|b��<ک:� 1wڄEJ�>,������/{��@��'&�'A�	<��T���*7.����N�f��ݟ��	ϟ�i>��' V7���F2v���C�pc�$F�&h��
E�g2��d_���?A�]���	�0sشp��U�7$��]����Ŋ�Q����d�,��Q0��w�����>��=� 4�y��^�d��Rd�T�{�2�+`4O���ć�K���+�gT 9@C+-�t��O,�DU��)�a�3B��i��'3�Ы��wP`���ܨB�Jt�(�d���� ��|�G�)��Ax�s�l�2T�:��,�z���O:I��ӟ�����O����O�dКk7���T�`i���w�W�\��O˓)��AC"C��'��V>uQ4HC<uhe��bݪ(3 �-?Q7^�����CO>��?M+��Ohf��wb	,k�v�x�eL�b�̓0���"��*��O�.6�D"Zz2��@�},��SC�Z�P���O����O��I�<q0�iC�pbQ�x�U�e	O,-�m�5vR�'.r6�$�I'���b�P���l��=޲C �0o�� F+�ڦ��ݴC��1�(OP��ޚk����	�0{�b7�=����r��O���	hy2�'92�'���'n�U>�Q���%f�8)�N�)*f�œd�ې�?�� ӟ��I���%?�����M�;rߌ�bgd�fL��צBTD#��'u��1���tꖎ{��I�1&��F�΃q����աbgt�� j�� �'X'���'�r�'��l�!�T�4⣣K��Mˆ��O����O�$�<���i ���'���'4.��k�=+h�{���;S�D ��F}��'�"�|r�\/D�*%�qZ�
��DT"0
8��f?�4�H<��'��NײO�a��L	�V�����l�"�'���'t��S�����'�0s 6@�&�6/|Xزg	�ޟ���4hb�����?��i��O�� ]Yܙ���Y<I�2�@ڄW����O�7-�A��ÝF�@���O���խ�.T>��q�)YO��!�Z͟��'C�i>�Iȟ���ϟ8�I23�(B��8~�bM`����Q�ba�'��7m�'z�"���O���<���OD��d��YЄ�tO���D�*Bx}��'B�g2��!j�����e�Z6���n���(�1�J]���	4-[��3��u��|P�P���="���'\�0lni� Hɟ��ɟ �	���pyBKo������O,��W�#Nm�'mD	O
����O~<o�A�F��������ğL��g�&"�ht�S�ը��̚$�*>O��'�bo�<k&��`���� ��/ N9���-%�9��;>����O��d�O*���O
��,��@�R�	�p؄Z aH�#q ��	џ���&�M��C�|*��!z�֙|"A�_������^�&��1
g2@O�o/�M[�����,O �����$��ԭYA��x�v*üZi:��5E�+�?�h'�$�<����?!���?��I͸�	���J'�@����)�?����d����#v@\Ο��ßt�S�?�V��QI��H ��<@��1?�#]�<b�4cܛ64�4���ɒW�v@��	(4��Z2#@�,���V�L�M#���ch�<Y�'"�.����O��C�ǝ@r��[�l�&a�(�ON���O���O1�(�*]���U�l��Pa����v5B�B�:0��f�'��E�X⟤ۭO��oږ�B� 6+_%��U`�gE?:��ts�48ƛV��\$��柌0F��$��dfEoy�Nٜy�Y�s!�nQ��x���&�y�]�@��şp�	���ӟ�OO4T��+�&a��}�f� fy��1'`�,U86L�On���O����D�Ц�*2��(!O.g�j��$C�K\b�)۴{$���9�4���i�����d�<A6f�'BK���� �I� \�0�	�%"l����']$'���'�b�'Զ����Y�]`�T5i�~4V�@�'#B�'�rQ�|��4C����?�����)��/�4*&�I�4����H>y��Z��I�M�i�FO����F�N%�ƨ�8����8O�Q��4Aa���O˓���<�I�q9��rC�¸i��(p�@�,[��\�����ʟP�It��y�&�=Oն�1�ɓ8�,��d��`�h���O�$즥'��s����]�o8��w�J
oT�*vOf����43����{ӆ�y@4���7N�0��'T�}�c��FG�q�"�M5<�TRd�9�d�<q���?y��?����?D�Mo��(�I�t�}�Q	J���$�঱�'ŃLyr�'���^>q��H��IR��K����+"����OXn#�M[��x�O���O��a�g��1�&�[���1;SNöm�RU�<"��L����#���<YAZ�{��piEzH�!)��=�?����?	��?ͧ���ԦA�C����s��I��P��Ô|J`Ѝ��H�޴�?�J>	3Y�H�	֟���15({P���0�����:I��D� y��'�$�[�l�E�+O��I�Ԣ�%P$,��qH��+�(p�78O��$�O��d�O��d�O�?tm]�R��J-+���������ٟ(j�4ydyϧ�?���i��'����S�m܄��h��ƞ|��'���'���X�^�0�'40��b�O&[�n,Hf�&h%�Ɋ'"�-�~�|�\����������� ����?�;Q�/N��ek�����	~yreu���!p%�O����O��'+M�=�c�
��ل{�(9�'����?������|���_���A&�f�@����q\1���4���O���M��D$��S񆁠s?���b�Σy�Ib�A��D�Iԟ��I��b>��'�b6-հyT|H�4��[
�/A�>����SE�<�զ�?a�[���I"0�4��B�6$�
0۾e��t��ȟB��ny�П������?͖�� �J+��R�M�싽;vL�x17O���?A���?Q��?����	A�ߒT�$,�a���JgfW)?^h�nZ'�U�I՟��I@�՟  ����3�"Z5�|�B�(�CJ�?������|���?��&��
�(C��b�Ꭺ&��$y�b&.�d�*��z�'��'x�����I(��h��DU�|c2=0Q���T\ @�Iݟ0�	ȟt�'IN7��D�D�O��$H���0���!��<��� 
�xH�O���O��O���&^�e���[ÇQ�~$�-PĞ��鷃O;�tZ �>ͧw:�����Č�~�JDy��gyt-��?v����O �d�O ��.�'�?�'��:�t��-g�8��2�G0�?Y�i�� h��'_�dhӒ���q�:@P�a��LH��L+�~�	��`��ş�p��D�I�t����O�:�`-���N�[�h�`�ny�O�R�'���'�RJ��y�~�a�Ԧ<0�T��.l�剆�M#����?���?QI~�� @�T �Ϟ
g�"���[�5�tq�P�������%��Sޟ��	��nXP�J/BN��We�3�ZM�PJ�
��Yg��
��O�7��<1�ΕT?��q1��/|@����ׄ�?����?���?ͧ��$�֦��qLȟ �iP�5�Pё�Q�����Sҟ�P�4��'��ꓦ?1���?)DJ��h��p���2.��CG?+%�M�(O���Y�"�z�'���?�]"L(,	�ًkV�b�䍈#H�ҟ$�I���柰�IO�')ҩ�"���`�RЈ�U]X����?�����& ޜ��I��$��:F�<^ ���S�p�xb��h�I՟��I���Lny��'�����ӳp׆(�U/Y�F�(@��kʄ7n2)�	�[��'l�i>��	��\�ɰy9,}�oX<}�8�4%	U��l�	�T�'b7mP�3�N��O��d�|rs��<Y�T�g*��!�4�H�a�O~��>I��?��xʟ�(��A�0R�2�8�.[9x����"1�dP�����i>m����u��|�M�~l|�!�Y^�����U�1��'��',��Z��۴j�X��s/�7@��:p��-5*�+SHΊ�?)��_�����i}R�'��9H@Z�����A��^N�"7�'?�7��%g���?Y -C�|}T��,}r�ӱo��y�s���L�
�P�yb[�H��ȟ��	���	ȟ �O�te�V�:�^E�!��?I3I�/tӲ�"Q��<�����?T��y�%w���ibm�
0T�ك�G�R���'ޒO�I�O���ʀQM��2�>��U�)t�l5��ĕG�ϓ^�����o�OV�yL>�/O��O6E�F�Xp˶�$I�Z{�1�J�O��D�O��Ŀ<A��i. q���'��'��㳧ߙ3w�2�Z.�����ĆC}��'�b�:��σ7�hal�2tp�gx���Ox(�'D>�p�O���Ӎ9Zw2�AK~��Ʈذ,���ä,�7I���'���'�"�S����a�T rjP�E�(|c^)��OʟԪ�4Z����?��i��O��;/���ȇ�
h9P*�z\�o��l�1�M[恏����O�R��:�����E�`��[dIsQ(���UK>Q,O��Op���O��d�O",����x��X6��_� ;q(�<�g�i,�4�'8"�'��@�"b�}�Q�C.˜.!�{e�\D}��'�2�|�Ou��'���ÈؗEے��%jRj1�A���V8*��U�Of�d�-�?�;�䓶�d5a��6�W�o�t�(Ѝِh>D���O(�d�O��4��ʓO0�v&ƣ�R
A�3�B�h%HƵg)~��b��� l���
)O|�Dt�^)lڒ[B6Nq�}8�Č� ��J�m�S�I� ��}) �O$q���.�i'���ᣏ�:MP �bV�r����O`���O���O��)��?qT�7��D����ԏ՟y��e��ԟ�	2�M��*�|���<ț�|��&)8�a����%����l̢Y��O��o��Mϧ"��!M>�u��0��S�nZ����Պ�#h\Q2���O�%�J>*O�⟨��\4c,E#q �lgF�x5`>����U
r�"�'�2S>	`�EO2��惀 5b$ 5�=?1$X� ����('��'��A�"E�����6,j*�낺�dq�����4�FԂ�' �'5XL��S�D� ���c`�q:�'*�'����O��I��Mۗ�Q�;�.yU��-�*u:�n	�U ���?��i�ɧ�4�>Y��*Tf
`�z��1�
 @F� Y���y2��
��Ӻ3��ٹ���\���D��~���(�֫@v ��os�T�'���'Ub�'��'�������N�i�$�*O�b4R��Wf60������o�S�8"������Ir��Q��,�h`��@��?�����|���?1������$��\`=K�l�0C ]�"��:L0�dֳC�b�'e�'��	ٟ���r�x؁"��q0<l��� `���ԟ�����Ȕ'n�6-\��d�O����<i��[��$�U��j�5|LN�`��O����O�O^�� ��A�Pr�M�
���P����L]�.�����y�1.����O���B�#�6�J�Ĕ�LF$�p��Ob�d�O��D�O,�}���0���Td�ȡc���J�h��[ʛ$�;��Ŷi��O��X�B$�'(���yRA��$5��$�O��D�O��!H�<I�k���H$��v�� ��@��T9�^E�Ď� GD���.�$�<ͧ�?����?����?�"�Z/|�y�4E��tp��k����$Ҧ�B�@џ��I��l&?���9'�̨�*�.�\��V�I�y<T��O����O�O���O��䙐4���)E��D+�"�xd����/�O��P>���K���$�ԕ'�(���C8������4���ar�'Z"�'Br���tW���۴m�p4��`:�{ Ϛ<eVX`"GcO�~�+��ܚݴ��'���?��e8��\57�ءx��ՍR���`b�����|Rb�
�A�SK�'��{#h�f~�P���I#?ӄ�i�j��<i���?a��?���?����ٝ)���J�֣�e�r�ݎ/�"�'��#~�>d���<Y�i?�'�b�Hq�[�"��`E���`����|B�'R�'D�*�^�8�'&)|]�pΐ�J�lsԣП,D0RR��%�~ґ|[�p�I�D�I埀��Rx�<�`@A\?�9�M��t�	my"x�v�d)�On��O��''�N �Gџ@���`�� �J�`�'2�듊?q�����|��\��A��R�6�`҄T3~|P���Ñ.��L�����������'M�'c(I��)����� Oh *!z��'��'B�O$�ɗ�M�(KDȔ�ՎM�l�dY�M	�Q1܅����?AW�i�ɧ�D��>�ir��R�P�?�VTi��O:"�|�)��p�zn	Sح�'�2�І?�TD�'��̕���[`NC:O���⃋/[L�D�<q��?���?A��?q(���1��(<fb9j��]�0 U��\ަ���l���I�H'?���M�; A$5w��¯�I*�����?	K>�|
��E���ĉ�nMj`LP�U�D u��>7.�֤5�@�j�'G�'��i>��I�O��S+]�;�1p1`^4]x��	���ʟ̗'��7m
�@�\��?V��"g욐hՠ�`�+���.���?	�T��hߴ&��� ��*:���`'��(9N(8��D�W�IQ�r�*�噠j�0�%?�2r��u��'e�R\tZ 5(���)���y��'�"�'���'I�>��I�~x�qJ�#�2qoD`��&��y�I(�M�)ƈ�?I�3���4���S'�/'O�US��Ҕ��<J�5O����OpEm>K<0�'$�)JX^1��:���b�#֭?�r���	�O�D+�|�W��ǟ��Iן(���x�I	d��82�߁7n
̓W�cy"�oӞ<�G��O���O���d������ƾ �� q�'T9Mi ��'�7�JЦ�"O<�'�*�'"(8dSte�[�I��Ǩ�W,D��?�/OphؖC��~b�|�^�8!�ǘ#"G4X2�Ӫ���w�ڟ��	ş<�I���jy2�b����N�O��Fgӻ8�*�pf(?bƴ3=OB�n�D�I��I��MŲi� 6�ߕQ��!@vC�		���qƈ� u%�P�*�<1�Lp� g�?�'����wj�Hq�P�l�{DJߩZ�}�'��'���'2�'���䁤��1~F���-Nd̑p���O8�D�Oʽn������'�\7�<�$
��(�d���2���a��P�T'��mZ)�M��'(1���*O���
�jϨlY3��$j�����Y����/���~R�|�T����ܟ��Iڟ`C�$��-�� �0gÌd�����Dy��hӤ�҆C�O,�D�O�' �q���� nQrܫ���(_G�y�'o ��?	�4�ɧ���|0p���mS��ɞ�&�FQ�8u���[���p�>�Č<	gDe��\k_Ft31�
�+����O����O���i�<ђ�i��a򉞤tǾ�c�͒&���i� ��&�B�'�R6M>�����Ħ��s/=*����E�
�TARRk�2�M�W�iw���0�|"���4ڬd�'���@4Pak�.��7.������t��<����?)���?����?a(�.� �K��	�F9� b/W�����lE˦	�Q��iy��'�O�R�w��n�Rtɸ���dn�P�Q��xͦdn���M+`�x����*I��	�x�F pG�G[�)�����I��ps��O��O���?��AB<��⏬c�ԁ��_x�a���?1��?�.O��l�E0�@�':�-ϝ*(�xFEM�I^����"��'�$�>Qc�i�6�K�pФ�EF�
 I6�(�ȑ7 b.�@mh�J
8>@�\2I~��j�O���O���F׾R�9���J�a���8��O2���O��D�OҢ}λ}���+^Z�9��5,Ҙ`Jwa������4�������?���i�ɧ��w�Z���iKL��K�m��X�5�'x�6M���eܴ"f�HK>�&�U#ʈ�i&A��a��`�����4J���^�YN>�,O���Ol��OL��O���V$S�q�X�X��<� �i�l�OB���"��T� ��s����̙q^�U�#l}��'���|�O1��' �	k�Ô� ��,��`	�.bv�U�6Q�'avm5&w?9M>1+O���H�P~biK�Ŗ�!.t��PJ�O�d�O$��O�ɤ<qջi�M"%�'|�i���&C8H��)�#%����t�'�,7&�4��\�'���'Bn�$�r���<��eQ�x�X�0�|�eј딹����'r�"��0E�:
.���q$�8e�е�I	�O|���k�<��[A�찙�G�0�	!�'�6q���K�/̸:��!#0�Af��@d������-�l���rzf�r��S�<aX��C�ί82Z=�G�5?��ǘ�]w�HsG�=[��ژAN�eٱf�3}p� X�D�O��]�%�]�_����f�4�ߒUf��3c�%р ��Su�@�,��A{W�-.Ş��B
=["4h���a��B�o�57`� ��G�0͠����':��	�� ��oO�TkvcH�Cd��C�9����i���'aB�>T�����O��Ɉ*,2H)7��z�D�p��LNxc��1ӦS�	���	�ȰN�|x���HW�<VP�!���M���%5 슥W�<�'�"�|ZcDX��'����O]$	4���O^�8%��O�˓�?���?y/O��!�ǎU�u��o��r�@E8D \3���'�	�P'���I��@v��:/���F�@��5q�-�(�$�����x�IKy��4KF�S�>Q��ҵ-�W;6���A8)&6��<�����?���?���'!��W��E�&�!Т̙�@�"�O�d�O����<��Č�E�� �G-�5�P�@GDˎ|��dP���Ms�����?y�
� 5Љ{B� %�>�S �ڙC�<1�W��M���?1+O1q�]R�$�'���O �Hl�l2l�!��ͼkq�qq�&-���O��H�
�㟨��3p���%=A.L��خ}>�nZAyr��p7-�O���ON���n}Zc
�}
Q�]��V���]S�LE��4�?��y��(������:;��T/M&}ؖ}�E��//țf�\�7-�Ov���O���R}}�[��%I�u�Q�e!�?u�rH�j�M��K'��'T��������bdW
h�&�L&c�>�l���I͟��$���D�<1��~�c��y�	k�g

v�T!�0	Y���'�D�Xd�|��'�b�'��u��hԹPT4�h%d[�z?v��(l����U�a�'��I���&��؇#6��PAK9���ZPh�=Ȭ�A�yq����d�Ox�d�OʓA]����1F �
� B%
$�1�&gJ/U�	ay��'��'��'ި��F�r#�Q  �F0L�x��J�sh�' �'9"R�@�ˉ����C�!�
��'�
u|�z!���M�/OR��4�D�OP�Ē�8��0�޸s�BN��ҡH�����ꓖ?����?�-On=B"��z�S�7�����SX�س��0G��ٴ�?�I>*O��S��O��O6rl�F�'F�
�IRM�}���4�?���dó+8�@'>����?�؆p}����b2|Ollq�^CRH6��<q���?�qk	��?	H~����aπ	��!@WMD�=G��{@�����'��i0r�}���O��O���gޤ�ɱʣm-��H��E1Pp�l�Ty�͋�&Rb'�i<��iy�Ȃjԕo��$_�V3�5I�4S���2ǽi�B�'I��O�O��G�9�0�6��91/��	c���t���nZ>3v���ٟ���ߟ��S��R>Ya���N�� �#�����hۛ�M#��?y�Lبis+O�Sv��ma(�e�̆:
j0�C��H��m�<)Em�7C�Ow"�'\�-�a@��V&F���E�� 8��7��OH-��(N@�i>���ܟ��'�)���%�v�`f$єpm:-���t�<�$_�k����<ͧ�?�*O���8�d�b��=�Di��.��b�o�<���?Ɉ�'b�i��(��ˌ	`uѕ$�=D ؠ��P��d�O����OTʓh�,%B�6��Ly׏\n�}��@'PRF0PtS���	�����by��'��! �" ��s޼,�U�N�$x%eH0IN���?9�����O�s҉�|���h^L*u-�&Q6��C��bU�БB�i��O����O�rB��9��'m.��EC�A�>��B�
-X���4�?�����D��&>����?��	xqv�# N�0ia�-v��#X7�<��?I�E���?IN~���C6[��^Muf�o%�hJ��Qަe�'�B�"(sӒ��O���Oh4�A9��gB��`A�S&@':7UoZ��I�t@T��ɫ��'�(����>v��1���X�m�>4cT 
9�M!�9?����'�r�'��d�2�4�k��YP�!1�ω�e�|12G�H�DK��'k�'��X������N�2�A�����RQ4��yo��8���@���Ҍ���|����?�vLU����4��Ri��!B��Wś��'�B�'I�	3��~�'��'�*J I�pk��	)^�"��A�i�F�$N�S��5%��̟���{yJ��,����$�F]�W��%t6��O��9]��|��'��\�XX�(�	`�\�{#"��Ԁ�?~� �I<���?Q������O~��QBv�� ���I������ӡR�E�G'�ONʓ�?����?1)O
�!v��|�e�]�K�FX��+��s�9Y�fBD}r�'(�'�ɟ����9 "��ie\H��G�l����B0Z�؜��*�>i��?Q.Op��:ns��'�?�ҐM�i�D�E$1-I"fJ������O~�@6"�:I�xR�[8�NP�p������C�M����?�+O���-�D�S�� �s�	[a╕zzݰ,C�N���17�!�$�<�C%	�?�J~��O����B
I�0�ֱ0)^0��O2�DO����D�O����O��)�<�;l�
<3�ʑwRtJ��lRTIo��D���N�D�u�5�)��|G�d�A�F� �̠x�I)U�7��%\<��l�h�����S����|*��+�s"�	aa����,D)r̛&O[*{`��'��IN�4\�x����tC��8�b0k��K Q0"��ݴ�?I���?IT
n���xy��'�����eJ�h�A�5(�rU�wn�&Uۛ&�'��'׆���)�O���O�)��cת��2��N�%|q��o����	w�<r�O�˓�?�,O����� DQÊ����p{#f^�-���a�i����y2�'!2�'F��'R� x�.����>Af��A�ԅl��E���°���<������O,�$�O]i6i�)���aj����lP*6���OB���O0�D�O�ʓ^��[�:�v�b��&+k���ab
Ѻ �iU�֟��'Tr�'[�'��yb��1�Y(e�8.�����W�V��7��O�D�Ot�d�<�6�Cc������<�:�I��1X��%5����7��O���?����?IwF@�<!���~⁘����!ȒO���r�A��MC��?Q*O��2T̑D��'y2�Ov"� �aš@˪���4�v��!"�>Q���?��v����Om�IH�QjK�V�J�mǉag� S�i̦i�'j�P2�oy�(�D�OT�D� קu��P&a�ƠCf�ӚW�,y���M����?�F���<	���-�ӟbr�� HW�V�y�rE�5QX6��<J�n���p�	ԟ��S7���<ɒI��8��ńL��i����֏C�y��'l��O���?��Гr����a�Ǚ}ۨ�CFbR�9 ���'8��'��#�h�>�)OB���4pg�Np�,�����yd�2�`����<���<�O��'�r��9j>��s�]�B4֭jc�v��7��O~��D�z}�[�x��wy���5��E
1�~�����gc�K��,����T,���@�Iٟ��	|y�k�hdr���O�0Y
�I��E���F�>�.O ��<����?	��S�!�����Q���ly�H�<)��?A��?i���$˪pF�1�'F�œ6g���ة��B�6v���lZ{y��'��	��(�	��@CM{���WÁ?RӨTã��211�Q'X��M���?���?!+Oz�hrjDX���'�H}٤�C��Ai��N�^���O`��d�<a���?Q��&S�@̓��i���j��B%��t:���+x�^�r�4�?A���L�в8�O���'���ɁD�R�RuGS� ����4�~��?����?�����<�K>Q�O�	HU.ř9��G*��o)0ݴ��č�y�HqoƟ,��ٟ�������Z@B�k�v��l0&_6v�z��i���'l�@ �'��'q�X�k��)����g$)�v�j��i3����Os���D�O��d��I�OX���O��"WMV!��;���>�h$��n�˦�A����p��͟ s�������^�]�^IӐ �8-~Ъ�4T�n�����ϟ�pT�
 ��$�<1���~����ov�y��. �@i����Ms���dɢ:�?	��؟���o�D�������3�D'CzX�"�4�?���A��ky�'��֘)f}�)�5��I��iЁ~���F�����?����?!��?�,OԼ{!���֤��R���	���b��>�,O����<���?���2��"`%ܰRn�)����QX�dꄦ��<!-O4���O`��������|���ʛ�j��?
	�౱�Aئ}�'>bV�x��ٟ��I�`~��I�76�-j5�<�p�g�4��0[�4�?I���?�����W
���O�Zc���$�
�3�~uv���@���hٴ�?9)ON�D�O��d�b����Op�Ċ������.��r�pcw���dZ*�n���|�ICyBl�K�h꧂?���"r�J(�H�ʰ�
T!�iـ$	*6�	Ɵ���Ɵ(���z�@�'��֟\�cUR)�@2�NW3zARb3�i��Ʌ[�=ڴ�?)���?���[A�i�A{�A9O�$rp&\�>)(��Gu����O�0OΠ��yB�	�t���	���%���
�j�����%2��6��OR���Ob�i^}R�@S��L�1S��C��E鹄�	��M�ah�@~�W���R��vc ����#�� b#O�C�^����i���'M�ҭ�������Op�I�	�����H ��6��S�$�6��O˓w��S���'ur�'�� 0W��4H�r��7�a4jx����(\~��'���۟��'�Zc��a(�'�
N�x�k��?ɲ��ON5:O��d�OB���Ox��<��	ǐZ @dE�Z��@��Vo�iBQ���'��U�����4���6O��@�1`�j�nQb�:�
`�c��I����	���	qy��2NR����p"�Fr��)Ë&?�7M�<Q����d�O��d�O�ыR7Obi��V�F�\��B �d(\Ij7����	ԟ�������'�S�n�~2��+��m��L�1U��p�7a��9�	QyB�'��'AD�'G�s���P�'����@ ��&z[�9�@�i#r�'	��d7n�����O��IC�p�K7#�;�����F.syR��' ��'cr�������#�0�y4��+A�$Z&7��(nZFy2h67�O"���O��)f}Zw�B,�K��vü!X��Y6=S��i�4�?���S���ϓ�䓅�O��0���p`�g�N�4���۴&|��Xưi���'���O3b�� �!(T���Ͻz��}+�'��MKD�<�O>)����'ц�Eē�\}�1�f�	�Iz\x��m~����On�DM:�H��>Y���~B-_�[X6��֛7��cI8�M�J>q���?�*O��d�O����TmZ��D�D,Lh�C.:h��io�I	5xO���OH�Okl�?��e�'+�-���2��?��I�4�i�	ay��'���'���r��HZ�m�/�luva� <��Z&�����?����䓟?��=6Fd���)/1����q�*�2�䓊?����?�*O���@��|
���%(��`��5ne��L�h}b�'�|r�'��h��$� ZuX��ՍO��Z��%i�x�qY�d��ҟ4�INyr�S���t���ЁF����a�}�Bm�Wn�ߦ��	t��	�����i�$A<���2�ݷI�x4���qu�f�'"Y�������'�?)�'�d[� �	,�����Px+���f�xR�'���߮�y�|�ݟ�,K��7"P�B��M%j2��i(�8�v�0ٴXJ�П8�����ÑzdJ}���B�@����&�G,(7�F�'��%��yb�|�iV�J��pI�CR9i� �F�(8��( �.jp6�O���O��I�N�I���B�n�z$�[%"�d�XŴi.\<��'��'�Z�$E�֮5��oW:-����E�8m����	�����-��'�R�Ov�ꖤG\�  & 9eX��ӳi��'���b5�'�i�O��D�O��'&U�8Ј����G�F#"�Ǧ��	#q�:���}��'�ɧ5F�Z�J�q��/{��,٦�Ǯ��$�2+��ĩ<����?�����$� P��J�>Am:�a�50���1��j�I����Iy�	�����<ruC�%���w�99���r�v�@�'�"�'�Y�0�1�$��$��5U��"/\����C�����?�O>����?�ъٯ�?���B$9<IC�л_��Pr%�+�I�\�Iß\�'`�,sw% �i��F��P��$̠|��@�bJ�?A�doD�'�g)m�B�'N�$ْLЙ��F�e�*՚��$13���'�\��fHI��ħ�?���ö���`rDE�k�5�\0bǧE쓗?)C�ߔ�?����T?�%y����h:�>e!G��>���rA���ʟ��I�?���u�]�Bm]�MIq)G-� �4�?��Lݸ�Q��l�S�q$�M�LմN����B��M|�o������4�?���?���OӉ'��m
�j"���/�#���6Ɂij�7��������	�9�v�ݍ{�04q�f�ZP� RG�i�b�'JR'��DnO����O��;��M�fg�	�i�^]0c�ЊFJ0����ܟ�ۆa�A�T�I$*Z�v�&]��P��M���X�D�,O��O��|�iP�N�T�!�NYe-X��.q2�:q���v/�z~��'#��'��I�V���*�ڶYF*Lywd�$J��m�4+�����O>�d�O��D;�ɹ
�6dy���VT������@�D5@���S����T�	؟��I蟈` F�C��O+y�F�q)�e��}��'Wݦ��'��|"�'��E`
6�=\ Z��f
ܞ]L���&��$n����|�I�� �'����3�~��\ ؐ0r`�3N�x���9*k0u�s�i'RW�T��ܟ��I3D��Iן��I�� ��!z1�i�`N��]X��M#���?�(Od)���H��'{��OB�A�*iT���OA�a�	�%�>A��?���V����9O��ӵ9{,9߻D��}�%W�6M�<��-W����'r�'��d�>�;jP&xC�L�}�d�!�"^}��o�ğ���u���	|�Il�'G�������E�,�AR�2g��n|Az#�4�?���?���g��dyR��!I�P��$fʜрӫC�xl7m�%���9��3�SП�Bd�v����_�a��iB���MK��?��i池�_���'�r�O��	Q���
�����HA�Sp�"&�i'�'ϸ��S�T�'�2�' 
%�B��]i!�/t:H�b�
b���D��g��i�'���ڟ�'�Zc������w�H���47ڒ�!�O��h>O���?����� �e	$��+u7���iT%!� !��<��Ify�'j�	��	П�ap��-f:���ڗHrƜ���
e5��	Yy��'��'e��'϶�1�ҟ�y�wi��*�&�X���7-���E�i�r�'���|b�'���\��ݴ���3�i�P�z���&H{8��'�R�'U�Y���/0����O����	�Tt"1�Ye$��`��@��?����'��x�&�$]�d_�����Dku8L�t���Ax�F�'�r�'�"��l���'��'�����(Ⱥ��W����@
���(��Ob���OҬ
�(a1O��;�Є���LaK:tH��	�Q�6-�<ɤ�*XO�f�'���'����>��u�f̩PhÑ(p���皍m�To�̟h�I�nט�ԟ�����0�}
���� �ڜ w��>r��8AU�y�`��/�M���?I��:rR�X�'7�������@z ���
%eh|�tӢ�<Ov���<y����'�4f녺K�H�G���r�2���&u���d�O��_v.��'K�I���;��Qi��XA�ă���rc�4n����'�x�����)�O����O�Q��#Ρ?WVx*�
4r�Lh�&JEަ���a򐠚�OD��?�-OF��Ƅ	�n]�Mu>�B���5hXpek4V���oy�\�	���	ß���uy����^��d33(��Z�~p15A
>��%g�>�.O��$�<���?��"8L��[2.j���Պa_��٥�L�<�OB�8 F�
I̠��ooj	;����BlV�:��x�	�;�U���+9|(��O�-���"]͂��U���������K
K��q��n��@4��l��k7T��l0�.���H�_�(J�+ؓH��:��י��	�D��j��m)NQ�5ŔMx3M�?7|�e-׍t�<���ڃ9�<�Q����4��� � 8�4�
#"�].���SJ�X2�P"�j��1N2i@��� �PY&�E:��{�N;dM'�"��A�E��p���m�X`R�'N��q��
����W �j�r�X�.�� `ts�L�-%Z3�� �z}Y��>����n�I˱D^^�D����T	*�CC�~2��ƚE�P��Q�Ӷ.��p�t�D��m}R�'4�>��>	|k�$�J:�"�F��=��C�	�]t��Af�	�����R�r�h��$p�'�V@��`:�6�X;�*��ei�>���?I�BS�>��pQ��?����?ͻ �����H�} e��ѿ�@z��:X�F����&P�g��83� ��Aj�7HC<Ds$̀v�1��.����:���|�� �~�%fX3=�BH��Z8}�����O�	=ړR���vbZ�<��	tEW:7?���ȓ*K�Ĳ2��4Rc�NQ�;����'��#=�On�ɶ�*�zs�۬2�Q.SZ�Y!w�*Q���Iڟ ��џ�z_w���' ��b��C[�[��Q'�]"{6|�8��K%JQxe�׏݄A,��ā>p�D���C�-��
�cD� XJ�g�{��t� K�24W���{}֍Is�]6�V�8�]�=`(���'�r�	}���Y��bT?d�5�WN	'�8�ȓ�� ��=)�b��ë��h���<)4T�Ԕ'd�x�HhӮ���O�<��t_����AN��Da�`%�O��d�����O��B0�m�_�"6	BW�n�4�;��B����$T�'�lc������8Y:��1��9�E?O 0�4�'�rT��" ��oDP�`��,�k��~���	ş��?E��a�[�*I� \1�qrwJE�xR�~Ӣ,h��_6�@x�$��*%�AJQ9O��?T��Q�|�IO�4gŷJA�(қo�@�DH�V0��I��I���'P$ȖEV�D��٦� [���T>��OH�@!���",U���T[R�r��H�b�í��}s��F��/�Myt#Q A�"h{%�����ɛA�P��O��}���X��p��ؕ��]�%�O�S��d�ȓ@
T��"F�����oֺ8� 0����HO�<S��&0��� �<8�@�Ӧ��I�|��.~�yR�
����	ğl�i��C�LX�
B�K'` �]dFc`7>�\c2�	 Mk���I(����|&��1"g�=D"���Q@�.V�de�O		>I��� l��Z�[?{�X�>�O�)H�� �`��oǬ?�"�#�?�	�=�*���|��ī9�,`�Z�q&��`�`���y"���e��	@%�,�9�V�������8�t��cM�Y�JVW��\�^7Af��$�O��D�O��dB޺S���?Q�O�������=2�:i��j'	@9���O}�|��Щ:[˸�3�}Ѵ���I��m�L���X�*���qB�X����p�M	�$E�q�A�@A�p�'%��6�"ؘ���-%�����m�e���$!�O�!�X+y�6DhCJ������"OF�Z�ĵd���(ЭQ������R�*�PÓ�i���'���e^2~^����.�#0d�����'NbڑM���'<�	*O�j7M<��V|"<��'�1a��}p"j �_i�x���Y��O�A�W�Ǎ^��a����F���"u�'6x�����?���?iwkʱUD�p@�,��I["�W����Ob�"|z��T9T�q���A�p��B�n<�`�i:p���F�a����Д
�-c�'��+kP�ش�?�����[ �`�$�#D��+��F4� @�O�&ky����ONX:��O�b��g~�r!���c �j(f�������	�C��"<�*tnW��@* ���dF(��'�S��@.c������~ԉxu��b��T���ɯB!�$.l�~8C�^�b #̘6.axd?ғ��%��ףiʐy
0ş�j�YгiX2�'1bA"-x�H��'��'�w�J���âS��a#�
c�-��
U��yV�en`��%"&X��ǝ���'Tr��ϓ8?�`��(S65[������5��yr$���?�}&���1B�w�LE@v�#	�hX�0�<D��&U?,V	Ѓ�@�^�[#�4?���i>}$�T���@�r�P���o8$s��/.k0� �@����I柼���u��'�?�6��B��8D�����՜y �xk㄁TN4���'�O���r�*s�p��'.ؕ����QcL$�'�pA̡�A'QTX��hF)б�B��&?]8'��u�
��,�O�iSPOB��15��	�����'w�'B4�BO��n����l��]~���yB�p���OꄹaJFA���'��P��DO+>���I�,Ȏe<��3P�'_2��D��'��)�3�r�K��ĆMYNz��`�p� � ��m�(�	AD4N�jP��'p�7�Y�&�x��Rk%kV�� ��������wB����#$�'C����?�)O^���C�;�� ����m�|[6��O����68ƅ;l�*)��qr��+H��G{�O�7�D�#��Уu�ݵv#V(2��"0N��<�f�Ʈ}@�&�'	�]>u�1�ʟxX��=5�"caD��ȩk��ğX���w����z�S��Oڐy�%])*OpAi���[~�)3�>��ȍN���O�� R/[���eNoo�٫N� �j�ON��O��� �ӓ��1���&�h���p�c�X��ex�hK�Ď�Y�,Hu,�}����<O�1Ez"Iӧ]���Fcý+rp�w��^�66��O��D�O.�K�4�����O$���O�N�y����˹e9�L�*�2$��@����v�h��4
�uSF"�F�g�I�0 ���B���f��s-9`?�: �=D-���i9p�l�h�g�I4n'���E,��Oǘ��UhV�i���<�hV̟�>�OȜ�Ѩ�+q�bU@�d�<|��t"Olp� ��dG$�K'Cˌ�F�w���Y����~?^� �l\ �N,�f�+sH��A��Ň 8�a������ݟ�^wS�'���]�!"LQ�Cn1:��l�r.���aO�퉐��M��� Y�)��(���!�d�M�N��B���jS�,+ᡎa��y�'���-��C�Y��suB�y�o0E�����ѡ8p :V�[���'ǎc���!�O0�Ms��?--4*\[R&�:;&�)�a�A"�����,��\����|b���+{����b�ȹ6sb�HѤW��#G�Xr���"���9 l��d�"T-+�4q	h���F��<.��hi*9��@�-ڕ=u�m@�%5OF���'@�'*IC��	@�bSń*tq���'>,+тL61�kbLǰ�|��'��7�+|<�,�cݤ-�aj�"��u�1OV4�t��ʦQ�I˟h�OQTp T�'L8�S��l3�Q�w�ݪ�����'�2"�.MCb�T>�9iX���̏�2����"oF 7zrȥO8Q��)���Q(�)�N�=E����#�_#.t�'�����Θ��O�.��cZ	��Ҷ,͡q$�'�Ƶ��nI?1R�%�Q�@|��A
�
����KUA�k��X���٘/ΈtK���?�MS��?��e�q˖B��?����?��Ӽb�Y�S��[f匤y2 @Ǐ)��'>� ϓi� �ӶT�܉`�	�Tm�=��	^x������+�f���d�p��m:S �G�s��}�)�3����c=�(��/�(�  �ߥZ!�$8k��DA+ׇ)�D�ؒnY&2
���HO>qj��À;�� ƃ��a���^.Y|x��Ο|�	Ο4��q�$�'X��C�/\R@�e��!1��Ų�A�:u�x�Ɇ�)�O�&h�#!��3Sh[\:�T;7��i�<��r�ݡ�l���'�^}!��!��=bh��3� ��	1�?�2�id7��Oʓ�?ы� ,�0���QU<�a�Z��Oʣ=�O۾�P�F]�e���_�T8�����|�i،T�7��<���	�A���O��7i����0+T��͘w�R��z�D�Or@��	�O6���O���C�K�C��O���0䘘t)f88)�K~\h"s�'&9���V,sal98������'ǊPv9P�C6j�d��Q8�D�� �O���W˦Q�I.aE�l���Y�F6��En��_�<��'����SJ�����Y8?T�x��]�-�T����O$�n�:" d�Z�L�4��`A��G�j8ڴ��d'@,8n������b�D�R�[�t�k�oD
0�l3iͳZ(��'�� 9R�'�1O�3?FթZBR�g雁E�Z}�CmZg�d��2���?59�� �
�h4��:w��I3n/}�Ĺ�?a���?�����OT�qi�OV�Nt:)H���.(,�ˈy2�';�y�h��\1�^΢�E�՛�J��ቆ�HO��I<%[��ht�+�����Z�e����@���I�h�)� �՟�����8�����r5L�a��F!� ,L���k���)D�0�)�l�g�	�Y��M�톫"��5(�*yV=!N>�B̒Cv��>�O����lԍS���j_���'7�����,O<��=��F�N�uŶ�ʴ-�-aTC�W+jq�Kϲ^V�����������?I�'���c���>( J��$�[$K6dr�@�G����'��'�x�	�I��<���D�� �奇;T.�Hk�b��1��XQɓ�e~���ũ@A�3 m�/'� ���S�]���1�C�7캵SF��f��X��h��p��"u�N�HH�a�D#<a3�7� �����W�t�ʳ���z�D��Dg�O��DW릱��iy��'�����Q<�Y�'J4 @ׇ��8�)
��H�h��h+�'w��#]�,�&��_��H�y��;�,X0ņb�P�dTL}"[>�2��)�M����?)$+��.�n1���Lui��c��H��?i�P851���?i�.춵aS�i��'⢱�ק���ڤK#*Еm]J�zǓO��4B�� �P-|���O��X&
�%� \X���jʌ-'�'�Z������f)pӚ�DL�!zh�U���s$3��!>�ʓ�?����4�'+��ED�P�j�Ȳ�Yޮ��	�'Ԯ68i48�E B9���qs*�	520�o�[y"�]�{eNБ!�'ARS>!(&HF� z��� 6�
�F;�\����^㟰�	%I�)�,ؤO8����0t|૭���'I!f%�$|1���KJ���O��rRL�3B�A�2o
5v���B�(��Md��gdK6V�����<V�'����l#���'w����'>�z1�u��if�H�eت��'���'p��'&� @��ҽ�Vg=R��a�=O��FzR��%UН��&�3o�@���C�p�z6��OR���O�=��I�SJ��d�O�D�O��;|Ϟea�Z�1e�P	�� �l%�s�yrB�_�ʏ�D��<
J\R��	6&��g��.!�Zc���J�& �q��'*�Xj��ÎG�*�
�!�ͅ�:G��'��aZ�:�)�<1��7�;�)�,-@bJS��b
�'�U��.��}��Y ��2��p�O$�GzB�AZ?�*O�4ш�D6��"��Ҽ��J�ݢ9F��O����Od�$�պ����?)���̒B#(Ť%��B5)'*pC�'���<��+p�1PÌ�N
�0��R�~��A�4S�8{���g��uR/�E���b�=(�l�cڂ5ڊ,�Lɭj�,�$�O�	lџ0�'���D���|�tjW�L�n	ī'd��*�ODyХ/�z5���������6,4��^��j�l�Ky"�M�1�םퟬ�ɶ;V�2���>lg8��*T�n�����	������|�b&����z�*]^�Ԥ�4J�d����Rr �C�#*h�	��6\�����؁o�b$�F�����Q�I)	,4�P���]p�4���:O ���'���'��ҳj�Ё�A`DR�&�8��T5L��ß �?E���O�LM#s�_�G���-�xR/p������()��1�᪖�Fk�s<O,�R�Ցb�i��'��S:/W���	�@��� W8E��!_R�
T�I؟��wgިB:v=��)ML~*�@ʧ3tހ����PYb&k��(�bQ�O~����*V>�ŢA���r�"}�U��� �|LXC�$]���2g�Jl�Ĉ;H�"�'��'o�Dly�bI���Tԡ��o������O&��8B�$CG�U�}�h�j`ߦ�ax��&ғiq�Qp��Un(�%"3�F�-@�\�'V�}R,]	g�2,�WF]�/�ثMN�y�m�dL�f�� 8Ā	ǎ_�yBKBJ��%�3���[���3�C0�yb��}&��zO��|�d��R��y��Ғ^�(��"��� ����y �)>�I�5-Cy�qF�=�y2���]��uB�oW�Nf~������y�d�b��ҝK�r8��k�<�e��(A�ਇ�!� i2F^u�<IT��L��u�R'w���cǞu�<�@�N�ꕁ��H:���P�Yi�<��  B���9tA��J�~�<i��ڪg|�ӆ�����a�x�<�SA=w ���s�߁~��s k�<�udJ�Gt��1SA��P�$��r�M�<1!]�&����`J_	"`�-
��F�<iP�ӟh6��.���x���@�<�c��	��M����%0�(QI�o�F�<qKοyDUi�-آ-8�@���w�<��պA�H`�r!�a<]����r�<Y"��4V�} �L��8�*ݠF�X�<�"G 0{+�P�$%B�Z�������N�<)D=Q�\�Go�
{N  K��u�<�"�\�q$J�䔂^՜�Z�L�<Qp��=�^��d�N����W��M�<iGN�9=���(T�0L���I�<� N��E!A�6T��/Ir�y�"O�lÇ�D&�xi�Q�ǙX�T	�"O"}�����r�D$�J�'�x� 7-�j:9�'>�����O�Ϙ'*�@4�U�3<~��e�M�/L=Q��g�T��@ҊH�.�rբ�7��"��1'g$����zxs�&[ʠq.�6/m�t86�Ś#��G~R��0a�xk��Ñy����ן~ ��؆�H��L�h��
�"O�8�B瓔M�r ��cI�(1N�!1�O�m���_��E�q��Y�]G��%P%��f��ՎlI�*1�yb���"�`���G�x�<�kT��".�Hh�8`��S��u�-�媘�&�p�э���Lyp�:�㝑2 ƀ��v�azr�Ɍ� #��Q���dȥ��4���� ��u`�K1�V:�L�5}�RiKU�'�2]H&�_i"�	5n ��x���y�n��hỗ/҇`j�*Z�caɴ��?q�$�K%<؉P]�R�d�I�H�)�y2�6�� s�F�.�S2/V	2{ � í2�h2�.B e{r�b7�-vT�O�r�`�w��Lan�k����F�.�
�'�20�I[=l��hjw
��'D �X#!;��r��r/�{D��U�"�7IZ?h��b�����M�����ewV�#��0LO�UI@��?��税� hP�� � "Ϣt�փۖH�.��s�0j��!�$Z�*��l�דT����&hA��"F�ǡ|^���<aƆƣxV��i������`������عBԸ��u�Й��=JF/T)��ywA�U�<g�>�ژaӠl�H,�5xF`����+R���0��"zAo�~��O�����wFp���Ev�M����O�DY0
�'b��B�έn�`Xاj�6+�U�J�>h����� ��"Fh�D-D%/j�ϯj�px�=�qB�{D��ՂȈl��9z!kAO���*�dE4`���5���w��M�@O�k�\([R0�43Kє!�t�pǕ�eՀP��'��l��j� ^�f��42 (H�y��0:�I�x#��
䩙�ֺ�J'�����;�x4���{����Φ=�C�I��l��vy��eOB�D��S$�A?���R0 ��M�f9�#2�Z�8	����'b*����n����(�%ޜ�s���t���+9܌��AK�?���|皕h�q8���!��1;�`<���X�R4�Qc�8b���38o��*A15����'��{���3M�8��@�[nP1�%�G ��'�4�H�@b��7�F�~�Ad�Z	���D�>zm����F[���k���-D��2O���q ���:!�I�������ɩӮ���MоYW�tsm�~M
����K�(�͛u�]'qW�i�Ӭ��_S����E��9�qOz�i��E�#�:��`�X�B\J`�Ǧ��F�^;ƦӉ�p>arfԽl!��p�� w5ԈpOf�F���*��L��,2QO%�3������m�Nĳ{����ҡ 3>��2|Os`#�<�:M�FT�&o�X� ���J
�"�H�1�ax�Κ$ ŜUP�� �R��� "A�w�r���?$�h�k�m�&�$�G��� ��Q	(�6�b�D�d�P(J$�P.U����]��@�g�H�Oq:hiv�<)m�b->�뤭�= j5�1OD�'��qħ^6�xH��U\|���]Ct�E��')X����^�<���s��NE��yH�y2�D�NUPa��Ό0N�& �wJsN��P6Om�	��	;&���! `��kd:)������aF?F���®��MS6j�ߺ�O*C����Zc}ܰ��eB�w��,#t�9&p>�;�'��c ƵG
XA�AY�T�T���b���~b֕�X@�II�|��.q�|��ʒ�r�����H2uMVAS�y��h{e,��f+�(	�#� xAcЅO����!;Q�8� tY���"�  4lD\�@��x@aԍ_���'(�P�@D)I��PX��3��y��sB���R(E�D��	���'����,��:Q���v�ɐ^(ljSg��~M�9�M�/'�{"oK%,?�I��ݗQ�r��FOY<9r�U��+�@�|��9��'#`䔧��c�� DY�!�#��c���C(<�T���sR��p�aK�&��EЅ˚*2�#<QA^����-A3_"��a���0PuF�t� �ƍ�4�U���%�)��.$���t�Z,(h�-C3EQF� x�e*$ @�H��zt\ݲ��!}���}u蹸a��#���@��$��'dTX�]�h��u�*[�1F#�O���v%E�"�b�0B`��J+8���'_Bdi򘟼*Ճ��(8�Hr��W��D٘#BӋ�X���7�|���V�my@�f��/#Dq�"��-aj�ے��!F�Y�6�'���0��OqP�Z挍++TQښ�y��GeB��@V�ytt�ڷ�V�*�!��7�l=wl�j��pY�O�7Chh(5�Ǳ5O6X�Rf�Qt4�9����V��t�'m�q[�G�w�hi*�O�B$�O�u��1�C�T�U����I������P?'�h�d�'IH �ELh��E
穑���g[R�T��N柨QЭ�Ey�1�M<�=�Rd����v�ԻJv�]�6��U~"��3���DeZ	k܊�0��
��M#���=5��Z�n�eS�������G�ŚO����6�M!�zx�D��==�a|�J�e���#ŗ�
���r�.-�(R2�^�|�|��ϓ�y� U��Q 0�
�H1"����HQOT��Z�9a�4hcZl�Z��v��H��2�'�5jkJ5,Z��r��`!�Rb^8^#2��[��Г��2U(f�Er�ؘ
�n��H_:bJT��1�����c$ұ7|z��邟h�(rT��	}���X��E��M��jN�]�#���Dy2m3<�p!fiB�����õ�����tr���t��4�2�� ���}���K�i�J�&�VX�$3oo���i�&*$m���:<8���r�@��b	�shJ�G��`�SFq�O�����>H����D�z⚯o�8�����������t�.}���V�yv=�=��F�^�v<�0OlPK���7K����8�% �E3���Pk��WZҠ�%��U�'D���NS�=�^hK��x��$=6��e���;"~Ͳ��W�]˲�a'�Mv?�`��?���|�<�Q���h��)�Dٳ\ff�tn�L���'9�d�l�3}��3�vU+�K�no��	F�D�D�Z�@�dG�?$����M~���]�BVz�f< \���R��69��7�:���<��H��v�� ���Tw?�ӥ`�u@ᢕ,1[hё���M2�$3��,Od���H��ܸ'�ȅ��!z98�C�MP<�ez�)H�H�����tX��g)���?ex�w�2%!'g�X���s�P;4x�J�O�L��������T�ߩJ��&䇡Hr���у|?ϐa�E����u��Q��Z�;yx�ܪ1n׉��@��a;�ɩWF�A���|2f�|�rcY�[�t����Cj��ap��f���DǏ�x�;�N=lO�N˰gf����e
�����$솃��yJ>� 䖣B'�d�I;hۦ�)u"�Ο�'o4����(X'E�����E��R J3�	697�^h7�� �(���o��%rV��흋P�.��gU�yz�Y&oE,\޸
�ү>�V��S��y�h�5~��Qcs�>+
���j ^vXᓄ6�n�㷪�;)(F ���e�D3y�,0b�ݳcMp���#
�?����"c�<9���<��ם�SMў�9���&��01���<)��y�@�q�{�虼�?i6f3���Ӽ#BG�.qK�u�ӎ˿)��$㊜b�D��,J��hO���gZy��� c=��Ѹ� �C��,�ݖN�����'F1x��ڲ�l�O�1`��#��*H*6�n	d"V��J�cE�U2�؀У	Rh�r ؁ҧB� �b+4�D^dc��J~��}$pB��_\��0��"��$�+IB&]s�r��"�T?	��� l�UZ 9O�չ"L�IB��5l��`�H�kB�p�  DzhQ��f�"r�O�-�ED��Q;�b\�r�8�(Ѓ��e��?Y��jL�28�*ԋ�B����s& hT���e� Dvr<�5��	=o��T�I���yc��!Q��Z�`P<�B�)E�?8��(���e�"=��8�Ȅ�W�.?��nѰU{�M�UDޝ~�̍pbϓ�2�'����ۦ�9�iʂ!+����$'h��kנ�*c*��#)�	�j�*��+��1jMp��Y�6ZA궦#?A�i\�DT0ūҀ���4F�k~�V�qODUrA�âF����0N�4�z���V�!r��Q#*���iX����ja�G�4��c�8{���?˟����C[}�< qd�R�#O&�p��|b�B�c�&�r�+����Dӣ�2��'�Ƥ�!
D��Fx��֗/x��� e\
��'��>�I�՘Ł��E� d� ۥb���xT�I<Z\u
D���qO�Ӑq�2qϻ���$+w쉷M
�F�h�����O���{��}��6b>(4��E�YfH�ӌ��y�1OH�ׄ��9�a!�R��t8����\oA,}��jӕ2�^(��΅�Q��y�bõrS^)��ƕ�u���,G� ��EpjU�gLؽ#/�$U�rU��O$'!V�{�b��IP���?���`	�x�D�$,h4Li'Kݡ^<��螧T�I��FӴ62����$ˍEQ �p��F�7��t�al�+���Z�DWAj��>�Ą���&�u�'bJĊG�N9-�\����0xj�#�T�8���&�U)/�.��=�O��� P?��YK���-6�䋃M��O�^�"a���d���`w�L�xXy���Rf���O��PS�k�*\_Ȳ� G#(����/�I-c�����u8f���M�+�rc�<�E��l@&�pB���q�z4 b`ΓQ��l�<ӣW#`����9#P�;��F�`��(��Oߒĭ�9���+R�n�
�A�"*z�,K 薼S~�xR#��>dV�Y�GQ�}��(���0d(���5����/�)�'(rpd 'jV*�=i��Ζ&�:e�㉊��e��zۚ��	�O�8�(�Ν���Y/;�ڙ;qI^����e�̉]����{*�j�1s�b�����]4��p�@��F�\pȷ�!}�=x���gQ#�޹E��F6�l�ÅD�*=�މB��zi1OވF��:��aa��V�t��w�ĜN� J3,C�Pɦ��	F�y���� ��tC�$�'���A(��dJ"ɔx,�h��bX��E([
R*���gy&�B.��z�Z���(U�"��ys��'��` o:_�1�I�)���GS2Bx��a���1S�@�Ƃ��4$!����y2AK�v�V�9$��+E]X3W i�铗�' F�{���+�X1S
6�y�ρ�`IV�+C�����97)�UV�$e��6��H�'g��]*i$,�ƅ��1*�kW:g�d�DàjT�A���F:v�qRGF�?-�&��'j�$�3u"���tt "��|$���#����%EW'��	'�?� ���J��� 䲀O�H]�͸v!�p*QOp$L��Mʬ+��I��A��� O�T�S+r2"���	G,	���sF�ޝ!���I�=pŐ� X'$�S�?Kd�)žith�R7�+!q�9Qt�8)F}"G�5CN�/�3E��郗j���Ϙ'αؑJC�;J�1U�ì' ưX�O�Aa$�Ƨ�@�c5��;3BI�=Y���]qΡC��l]&%�,�v���Z���@��mBH"qF}R��yg%�B$���kX�6���&)	ֲ�"4AC;��c�l�T���!��-�'D�$�-{b���dS��|�y����#>�aG�Au�m�j#�S�u�������Ov�p ��ϔ�'��H"��(+�f����|�uH�~]�"R��<���<���5>�"d{��3}��I�<>c��c��)YH�k#ɉ\��ϡvn�{����	Ь����-��鉠!�4��g�L��IS��<)��
r����b�#۬e*B"�b�������Ğ�,��٢�	�4{��CvW!�D<M����p �+x��T��F!�$I8|ڄ�[=&�|`:�%R9K=!�d^�%M@lkW�A&L�y@1CL�E�!�č�3�֕�K[�0�+�G� %%!�H�F-hD���y�8bU�B5);!�dI/lX��X��ıyjt xI �!�D͊њ�ҧ%�sc���! �!��
 �Iz�MN����i���MY!�0sY �ф� �z�@�b�ƞd7!��d��X�(�!U%���R�Bg�!���0����� �.\""�ԁr��C䉠>���3%�W�F���e�?VFC��(_ƹҧ���v�t�#Q�˧��B�ɯH�zY�'�ץFVJ�b֝��B�I2jݦ5!pJ	%&I�H��һ��B�@�NVR�@ L0㣞$��=��'u��M�;P�'fG;�H�'r�k���|�1	�Z�2�yr����$y4L��afe���>�y�ϚWS��7#& �:��1�yo�$:�R|�Z-!� ����yN?i�<��(\�D�nH�f(X�y�'�2��i{`"�9�� �T��yB�͜e�,Y#Ç�$�pq�b��yb(�Q4�Ԉ^��Xly1���y2)�(K�fG���D��s-�y��
�]y\e��!��h��T=�y�`�*j7����l�j��e��y ���Ȩ����^�dA���y���0P4uC#�� VIЃ�D5�yB^�N�F���@�p���iC��y�$��O�L��E�Μc�y�s	�yүD�dļ!�dj��X���S��L�y��=�����|��$�B 	��y�dN/f摸e��:{�q�򭑭�y2DT�,�R蛺)'��� L��y��YR�*�H�"�v8���4�yr��	�F���K�o� Us�̖�y���U�h��O��|�\��R@���y��	�&v����\�r4����Z=�y2I��o(杀��"m�ƙH�چ�y��
�`��q��bܘQ8��	�y�Q��1"O��H�%�����y2(L�X|��JBC9N�����mė�yR"���V���_[��$̎�ybO�eޔ�5j�&(sR���S��y2�Y�R��:BM� �d�Kt���yba�V� �"p�ˬGҰ�j��J��y"�M2B� ��@��iA�H����/�y��Ɉ0����3���54`Q��P#�y�%*��t��Y$��)��͈�y
� D���B�Kz����p�T;r"O�Z&�0-���P鞗o�,��"O }���}��� ��Q����W"O�\�q��(D�����w��E"Oʠ�䯗�� �#7!DV���"O�Y�s�W�Nfh�����>*&"O%����q{��S���$D8h�6"O�ա�����e ʕ8#B`R�"O`���#2)�}k�,v��cA"O$q��*li2�K'lh�\����y�n�2f����%@m�9@�П�y"��d�����$�pTcB ���y�@V�.$xh�Y�s�J����yRH�;��e0!�;3�}C����y�J�'
	Н�!G�@r���D��y��o�ڳ��"1��1��(���y��=qL�c0�_%�>��@$��yr�Ɣ�^�hdȜ#����e�&�y"�/+X,io�p�t��H@��yҫF�9�q�Ҿ~u���	�!�yR�H�g$�C��R�w���dg��y#�?�|L�V���&!9
����yR��	i�tS���6zB���Ǖ��yB` /ZS��)%�ě1�1���4�y��9KIҥ�'��<$5ڽ�����y�� �Ʊ���Ѿs��bDE��yBe֯*0�%Y��\(�u!���y	�*[�֡�D��#N6��9b� �~b�)ڧtZ�`�E�"�Iҵ)��~�P��=9������A�NDf��3M�3�+!%����R�t�8}i���|.=��Ɩ-!�d��� ӃǍSQZ��A�@8!�QPd��P`��S�PKR#n!�D�;B,�LǪG� ���U�!��=��Ȁ�[(������q�!��-�ASbə4������;�!�D�~����u)(�ڤ��a��!�DR�d�̌ "��x��#�b��!��.�N�RH�R�����L��!�$v�i��MH�;�@ȑ�O�	m�!��3d
.��߽|��H�CC�B�!�D�8a����׬�Ш:em�,F�!�D�C#���e ˶c�p 6�[�Z�!�$+f�����3|�G�8
��*�S�OZ|�1��t>��n�D#Fy�
�'�m�T�9S�<��敕D��̳
�'�N h����{-2E���8*c
�'*�`cM��G�zd�G��2&��S
�'݀�c��)D	�	@�2ŀ���$+�r��(�x�9��E�(,(AQ""O:I�3��0�F\��₈{��F"O�˰���c�4��p�v�
 "O�����L|
��1�8X�P�"O�����2A����M;���Ж�M����ú>]�0�U'@�lN���$D���'GR�݂���R�t����'�d3�Sܧl���M�P�,�bΕ�|�XL�ȓah8{�H
k���S"L�����ȓt����p�ƥ��I�D솴e����<�* {�팈��x1�@������X��0iT+�R�:Ԯ�0( .q��	�I֨#<I���]��I6�űM��В5��_�<)�bص#@x�HS/YIx���	UyB<w���Ӟ|��)�Xo|�9�BR5F��Icҩ.I�!�� �� S�[%:͊�2�iĢ1�
�zF�d�z���C�G� Q�N�����D��UG�+D��)�(��ؽ��Y�mz� G�.D�P87��&��M��-�0m�k"c.D��HU�N+b�D�	�Ɨi ढ1m0D�,A�с;~�j6�%4w��f*OZ�i��R鄘sc�0/���t"O�)z���Q#�t�&��&�q��"OTLɆ'7B`~	砗(WiAu"O�yI炙ȩ5b�w$iAG"O��x�h��C�K��A�$*�"OR�R���-&��ka!�!�R���"O�m;j_9�܄����-?�<ĒB"O��g�$
�f���F�-x� ���"OV�c�jD�y���s"����@&"O�DC�l^�/R,!�%"۱8��Qr�"OL���~�T�aR��1,�����'#!��%J�ҹ)U,Y &�hi��	�!��	�AT��l�3	�n����v�!�D��0H(�S�G?,��ۑ��Nz!�77h��ǬR�N�~:�B(�!���$&��+��yY�a�Y�s!��^%X� ��S5x�`p����V!��*A�R���Rp$�x�C8)F!���1#
���`y���(��ךW�dB�I/Q�~���fՈ�¸ʶK�(�NB��0w��$ N��h���ϐ|����hO�>)0Sd_8e>2a
ɺw��Xe@.�O����5�M;y?��h�A�7m��ȓ=��9�?|�2���ȓ|�p)R�f�(\����M���JX�hC:�����ǁQe���x���hp�����k�M�1��Ia̓=9P@��6|�t`ۡL�)z܆�V3R�fж�*@���ӄ	�����ܛ�S�a� �z�J�Mn̔�ȓgV��	�-!��vAۊ���Ol�=�������`�B�5(v#�]�<Y&P�v���	aę=1�Vū��]�<�%$ɫ�də�K���rY{#���<�*���L]�u�ڿTtNȋuIU@�'��?��yz}3G��OފU[�>D��"SD�h'~e)�.^*4�hU��C���F{���_=s��QCu�U:"8��S�[�lN!�$���֐p
H�k��xc�Ӑ$!�$N��=
��@$p1ˤ��z��	h��H����-
��y��n7�!�v"O��rPi�xr,I�l( $�"O�X#2��<����	.0�#"OHM�fՠD� +�B �=�L��"O�6�N�&��;��Y>Ӑ�"O܅i %	{~�C5l�JWPC"OPʗ/Ɯ3'*����M�sT�Љ�"On!c�`��pHx����ZS(�b`"O�#%���d/��m4LJ�H!�"O�MҡI^?���0F���N8�&"O��{4C�h�8��=��"O@,��-��N-�DIH�X���S�"O��b �Ԋ  �T�a�ƹb���N�<I��_,��x���R24���b��K�<1�}hB�#���9/R�Җ�_P�<@��>���@��;I����kQ�<����#�����X�3� �O�<��ʛ�Z�����Ψ��Pw�d�<� m��j�:a>&	ۓ�c!ƍ�"Odth�/3�P��A+܁3
�ػS"O�̒2̅�Jr�Ջ�»2�B��"O&H�A�9%�B��
	w -��"O�HFȏ	 ��8&�Z��A`�	F���i��1� DҲ�!�����	 ]�!�dǋn�Ҁc���8A�~b4a��"O`���+@6�u�cD�ߒ�K��y����^��S@E(!*���'���yb�]�"�d�'+��r�y�Wo��yb�GP��DcQ�4���b�-�y��\e�ᙦ'ŗ~=0�I"���y�΂�z[��Ҁ�$qU �k!E���yB���.�Y��탻j�:]Y���y2č ����rW	�<�A���y�F�\��<xw�ðG!���B��y�R�إS&��Ȑ�A���yr'= :���I[;|�b��yB W0R� Kb.M�)��!�GH�y�JIDz14A��~T�ȃ�y�H�6��}
g)Y)�s�F���yb�Nb�|b@v8`���ylFL��H�V�6��`'�,�y�W��*d(s  [��AW(�y���&���"j���zqB��̞�yr"�
SG`��#��f�8TLI`�<1�oqP��`��ˁR�f�iv	�M�<�``��3}@��f��@��R��M_�<aB�ya7�s`�i"CH�AJ���2��t��;|�[�mޅ>ȓ_��<�3$�5$�p�YL��~��T�ȓ�4d8��T��Ixģӽ��m��\���J��''�r ���:@�hD��JB�$̭ k�4�(ŵzhZ �ȓD��x��b��[�
dC��ȓc���H�p/ZQ�ABY ά�ȓf�,`[�@�6WU& �6͹-|�!�ȓJ���q硆"&δu:&d��V�Đ��F a�Cc�,A�6�`�Δ�$5<�ȓ?�V���n�1�$	�	����C��A9���h�VY���S�+�̤�ȓ'��m(�Nަc�&���A�[�L�����ـ6D*hsj�27�DTK�AZb�<I����6a5�[2��]�,�v�<�U-Ørb�����Y�8 !	�^�<����M!������+S�U�%Z�<i�e3$��ts�A[)��4�HZX�<q�a��J�*p�c��%��:eόi�<Y�ˇ:p�aB�L�!Є���M�j�<��hX��n�*�E�a�ޜ*lD|�<� %�f$jj��__��{��\�<�!�.~ap�k��Vp��j�Y�<1$fU�^I�e���Y�p�v��'DM�<م�O�z��ǀ7n�����E�<P���(ǆi�&��4��1�� �C�<qԥ|����̖!fw���$Rv�<�A��2�x��h�c�����X�<�`��(���P�E1XB�)��c�X�<�i�7�<��a‸{HдeWT�<�E�1�}2��_����V�O�<a�lGt�X�ŕ	+�XT�@/�G�<IaǲT�ȸ���C:ӂ
���E�<��I�OO����%AzX��P~�<��C�ۂ�(�%��#��mIT�{�<� .� �+���he��WKS�X+'"Ox1��KIn ���!*�',B�!qS"O��*�+��g�X��G6++�-b�"O0��⊌$�=�d���iA"Ol[��?VXb���&�$66��2"O�A�mQ�]�)M�m��B �>�!�d=>Z�qN�2~��py�Z?}\!�D�#�`��Rl��B�����C+\P!�d�.qZ0��HE�[�@pj�V�?6!��J�?����&��%�Xy$�L�.*!�$W�∹3A(+��9��ܦ !�$Q
A|��p��&!���c�Ǆ!��֚Q;E.�B����!Y#!�D��K�Ɗ@���@,Y!���0d��ؐ��R�4��xH��U"�!�Ӕߢ�ƅ�Rt�r@E�.-w!�䆹W�@4��e�zM
Up*�`l!�$�~9�������b/\i�j[$yh!��ѹW��X�D. @#�i2iQ#K!�d�@*M�&�P>-��Q�NW 
1!�$��V�X�k�o�<b����ؙ'!�Dϭ����k�$�t�v�	!�d��6�Ѐ I�f��<�iV�%*!�Ċ�S�4YҡŀM�Duا(��R�!��[�8Y�ɖC��i��@0g薵&M!���VONA��8t��P�u爡qC!�$Z1,���@kmb���+5!�Dܗ[�|Uh��#O���/xO!��F�Q�rD�ud˵e� ��ƦFD!��]y")Q�-
�%|h(H�ʈ�3=!�\�Y��h�턮;g>U�Dǐ�!򤚼0x����j]#+�\!�ǙMe!�V�bz�uˀ�¬}8���Gғf5!�DV�\�@lS���"��E$��"�!�D[m��p��ίJ��IjD,R#4�!�D�J{r��LYP��}Q���!��T>)���:����X5!�d��VNQ��K�' $	"j��z�!��K5F`0!m'f�8�wBM'!��A�t`Y��;b`jq�۶�!�D�j��!�'�N�(����!�8Gh̙�l]�p�ʙ1��œ1�!��>AS�8`�:h�blxu�9	�!�$���H��]>'�С҅��!�bݎ��&��(c��E�n!��/^�Y��!��;$+h�!��L���� �	�88	����,�!�D��/H�,�-8zp��JD�o�!�䈕��0�$�B�%��X�S<u�!�ǞIQ�M�����'aD�Pn,|�!��X���f�ݟ+X�چ�џM�!��1�)����BK J�F�c�"OD}+�4$BHCq!�8�h��1"Ol�9f@ϲ��ԩ�@ r��A"O
��'�8|�H����J�h�"OȄ/��80�E�Zv��o0�!��	�(��9"�ӭ$0*�$��O�!�Q�Lxt��fG�s�|"CMY a�!��|{�s�@E�a�vI����p�!򤋞
Ș� Ö(2��t�7�^	�!�[�j�h���	o,V�� ��,:!�dD-� ��J�	 q���r�!���:+TTK�O�Y�`ɰ�M�S�!���|5LHdO�#�&$Y���!�� ����q�ظV	Z�N����t"O��*�&�	7V�T�EW�i "O�=X��� '��E�ӊ�O�Șt"Oօ�U��lf�)5�X9z�d�u"O�h�*��'v��[L�L��Ȁ�"O���c�M� `^@�sDɉm j	iV"O~\)�(M�<a�r�b�`���"OXc�w:�$�c����y�"O,d��`V?1!�	�BP�[T2	%"O�h�dY�dhʡ�� ǹ=���	�'I�%q'E�,���� @A�',h�Q�l�h�"u!�yx�"�'�d�¥ꉴE2iP��`��
�'���bC��$ h:`%���	�'��h�@t�-���V�h��'� �� �_�h!uŖ:#����'i$�P&:����Q9�<��
�'�T����.�PC�!a���
�'g�|����|Xp\�C�Y�J(֠�'A{Ã/mj�Q6�<�� �'ڗ��q��� 8%,R
�'�]`e�]";E\��B9-�"�	�'�$Ԑ!�W���h�--j�,��'x���w�I�XfȁY�+��T�r�'ٺ]�2�]�[f��a �7V �"�'��SȖ�G��t!�POA "�'�da�B��(��Qg�"D���
�'rbx�q�	`ܦ���<���
�'������#�)��)�.1��'
�4��	F1�p8sFG&�K�'��TH��Ư7���s
U<�Z��'�ν!��tt���mY .�L���'54`mX+�����6r�> ��'\��Q��,30L��%ߊl� q�'��!�D�F�Ja�H��W�/5Li��'�l��Y86$<3�D�-/^��	�'�2YK���|���f�s�&H��'#l�$%Ό,�8`FLÇ6ZE��'�>����W�Q������,yJ� ����Op��0§�
�ۣDZ:<|��
Г6�T�'�2�'P���O|�J%�u����"j������.28HC䉺E�R�͗]7�(�GeD�BC�I==Bpiu��	���Q/�	,�(C�	�9&�z�@ӊ͌ �F-��}"C�ɜ=ٺ=bq�Nt��OǴ)��B䉮a��h9R-��R����'��l��?A��iO�B`�c�b]<���"I$E�S�h&��gܓe�F�PT,�P��X���	9�ȓd�m��
�GƠ���5�Ň�8��%�g��#ae� F.�&kyR0�ȓE�>��JU$8���M�O�xT�ȓ�=�fÓ >̱2��rWb��ȓV���8E��G���Y��jJ���T�����؞�i�@\<"EL��?�ӓ^^��5��5�
-q��ȓ\� Ȑq@� x	p���>���ȓ`:���Ț '�\� BJ/M,��bu�pv�Q�3�h��4G�)��(�ȓ���RE�Y�8<3�l�4����>�l���H7�DQ+c-��PӤ��FL���"�Ё�Z���<�'����Э�0@�0h)���)`�C�ɮZ\"�[���7�b�1��[x TC�	�	!	��d�>�)Q�k�tC�)� dX���ȹV$A�q�ʶ�̲�"O�|���YT= ������ʵ"O�`��G�_��)�C�/����f"O2}��j�uN��d��={�4�C"OT�[���`
�[�Ⰼ�Q�^J�<�!�]mAP���WrNS�TE�<��oՕ;
v}(�/�e4�]����|�<�w�.{��L�%��<H���s�d�p�<Y�e�\��9�d��?lV|k���m�<�A��k�z�CF����n,#e �O���,��@>y��%F4?J�=�"��Y�h�"E1D��*穕/L���k1�[13���P5D��P[���0,�4[U�HQa�0z�,C��/n�@X�\�{̼��C�.O�B�I&���(��t]�M!�,5�B䉃|R,�pn��!�Y����ra�C��	9�����O� #�œŮڙ'^⟬�	D>e�`�z��D�Dم=m�\ۀ.1D�4³�R���E�w�ظ�ĲRD$D��I�J��(򖨪��*2D PQl!D�$�u�� eU�2\���
���y"�2v^�Ԡ$��O~5+�J��yR���%v��X�H?2��HEj�2�y�GG�6��qCNY��q�gDP���hOq�lI�!D� U|� ��e���C�"O�dpQ
@p:�X���G+P�-"3"O$"�+�\
DF�0���X�"O�UB��X�R��ɂ�D��]��<��"Ol) �l�)f����������X�"Of�c�J�1'¬�T�Z	
�~� c"OR�����бo�Ќ��Y�xD{��N�R����Bo�L���9��]�!��>Q����Մ��fy섂�KڂZ!��S���:ce�qL�A�j��!�$� V��ѐ�Ί#$:"�7��7!�$�1d��VC��<�����U�Q!� k��``N���
y��־�!�D�g�.Ӏ+�)"�`��A�P+�2�)�'E]0����@�j�,�#�%Q����'2��⥝�'��ccOW+6!X���'U�K7�0=B�$C9����'�TMec�X��9� �95�v�!�'TV ��e�0b���۳d�+.�����'�r,a�"Jb@H�83	Y�z���'|��.@�T��D�c8n��'���+s���W����U�9#&�
�'�z�IQ�Y�r���3���7�zi�'/��W!U�v�PLE꜁k�� A�'`L�HA���>d���#{F�l��'�	2e�g�5�H4��GaU��y̋&/���hH�Bj�Y�����yr��6N�F I��Ǩ?�I�G��?���'J��i�^}�� 5Z���t!\k�<A�D< O�-#Rjͫue^��7D�c�<9�����n�*�o�L���&g�G�<Y3��2[�8�	�5P}NdZ�A�<��B�q��tG(c{"xB  {�<���A���	�,�����%�x�<Q�  �-�$������r�(��q�<����bl�xp���9��4��E�n�<3�Ͽ�J�2��-C�����j�<qe����!׭5jK�bK	f�<�"��;4j���¸iJ��V��V�<�䪙x�Hu��1��ݺ�.T\�<� ��" FP�9�Ty�5l��w�b@ Q"O&��$�� �YzKF�(��)y�"O�|��Oլ��Lq������Q"O�$22�ݭn����� г/D��J"O@಄�>�<pzr��?"��t"!"O.��P�̅#
����ŋ:�R�a�"On�k1c�0hOh�rg�<(��(1"O�� ��V`��&�\��"O���dl0%ۗNu6�iY!"O��h�0o�,+��ӏ ���"O��"�L�#h"��K̠X��YV"O�5c�PE��H{j^/Y�Hc�"O�pxl[u�dhPF�Q�*Ժ�"O|,R���o�4���G�����"O�u�D��-�@-	UB;8h��A"O�`Z�aEK
��D���3�
r���O���2���"!o��5v�1���ص�N���%��i88����N\��m��P��Ș��53\
�����X��!��y�t�D�֛	�B�R��*)q�-��:j8��ƀ�<d�d
�.'zj�l��'���Q�K�2M����j3r��JP�!��h��D�93�oO�d��0�?�-O#~��XK����	t������H�<Ib��Eh�Q����B$4���j�<�צ�y©��͇�l�jۤ�EQ�<�ȃ1B���u*�1��ݪqL�X�<9� \$Ei0�y8�z���V�<�T'W�>
ʵ���B/lI9QGJ~�<�C�U
����A�M�z��$�TO���?���ň�b��cO	�T�A�'KE;�&��"O�i�D��
.������[�]��Ma�"O�$ѵ�̥d����H�A����"O�-���Ȁs�J�s2�89j�"O�!ff��.���EC
Eiy��"OΌ�U#I�_���C�֒C3teA�"OV�J�"�"%��<[Ċз	-�`f"OR8T�6Ÿ�Z ��2�P� "O�Ak��K�|A�D���R�D@!�"Oܜ���܉���Cd�$�g"O�H����(u�\�s�E�vn	��"O��ë]����b��N��Ʌ"O�%-R)%=H%���@Y���;�"O�9�qN)q�9Pˋ'0l�aA"O� �%�2�-Ѕ�];�N�U�|R�'�az"'�,ph�V�����p����yҤ�$/VP�Q��&�|+����y�-�I�d[�E({�YY'�;�yR�J�{������ku6]oJ��y�g�JN���s!ɏ]n��S�	ŵ�y���25V�1�B� \NZeb�-�y�AX�4tZ\p%��#D�ROF�䓥0>	D�7���Qև�c�x|�uJ{�<W!�{j�)v��	o`���'Xs�<��'?i�!�4+�-	P�@ K
{�<Q'�v	��(S�|w�(H�u�<�se��D��p� [������J�<i���:̜D�A@Rlơ��A�<Q C�kG��P�gV=Byv��`�	~�<�4IהX���Ygė6k�B=c��{�<iH��	&����C�6F)�y���t�<���I�X��h��m�R�ҐH!+ Z�<qA�+K��X�Nź��a((�q�<a�Yƒ�w�
�bڌ��Uw�<� ���	\y���z��g�2%��"O0"�d�n	���GMkJ��v"O0Aڂ(f�ɲ��>DёR"OF�DE�6u&hS��R�Ftb)yw"O��c�/Q� ���k,L-
�q�c"O�H���!���Q�/�����"O��X��
�>�*M1ʃ)��S�"O��8 �0/T�J��E7t�Hp7P�,��ɴ]�J�Ƈ4�l�сF!��C�ɉYU��{����pe	c��C�I�O���XbH"AX�W�.6^zC���,��� ڼu9�����̄.��B�I�6��qq`��#d�9`l�,_��B�ɂd���c���OT�����"Y)����g�(*�����ćU�%�h��8D�,ʄm�-�:���KR�2�` ��5D������2S#2l)u+R/]���hp�&D�\���{<q�&!\�?3����$D���hG<얥&�@Y��$D���  �w(��#,V��(6 !D����M��e�`�q@�, ���
?D����?k�l�!6I�-�ހ�/D����)<(Ķ ;�KH�}�l���.D�X&�ٔP����c�)
�����-D�<;a�2բ|�oF�R|xz��*D���U���	yn�H (EBh��b@,D����Q�U$���- �A=�}Jm4D�<Ah�4i�~,��X�Z-���&�O��d�i�B�L��@����R&�	�ȓA��0��N_8]X0�;�C�,��ԄȓNDzz��C58q$�;p�~U��+�Z(є�?$��(��7hm*U�ȓit䉻v���Qx�����X5���ȓ
�]��,B�+��3E��2cؐ�ȓ:RƸ�4o�l�Y��g�� �����I����I�<�6���p��(hf��We�B��I�<��L�$����g���W��l"�E]�<1U�ڔ~c�݁�n�&R��Ѣ.�\�<)�a�V�&0�Ԉ�1o)�I9��m�<�EgK2p/�����2A��!��u�<!�CWd��L��'�08����&�q�<��Z���pht�N$j�b�B	�Ex���'��Pő�:X����gO.Z�^ #�'{Z���ǉ��(������W<$��'X�y�tCD��\Rd�I�b��'���蟶9��T)�([�x���'Le�e�RD�PX�cC�Ԩ�'2�����t�U�GJ��R���'4D I�A�a*�X�%�$E�Ɲ��L�H���KP��z��W!d��݇ȓ�xq�s��ee�ݐW HqX$��:�X�2�#�~$�V���{b�Є��.� �,���S �	�t@��U����h�Ly�mS�h�`�ȓb�EJ�&�U<��=��ȓ	C�=
��I�v�*'�@�����ȓ�Tإ��u�TM�@�d& |�����c��	k����W��z���$��,a�R�n�"m�v��H����Z&�;'W�d��ʔN&M�JЕ'�a~�Iϛw����O?`ϖi�c昚�y�g�3e,à\�OjL��3d�?�yr�Y��lk�A:���q�@��y�-\'A& ��b��2�b\y��E	��d�Oj⟢|� Ɓ��d/y�@�RԤ�-�,*�"ONR@��,4�3��CY{�	�""O��cT!>�arD��Ef��"O� �� ��%���`,�o�����"O����@1NڒD�kg�`�X"O�x���+)V��L.`�\�R�"O���S��2))�	�> � x��D>ړ��D�3xX��ڄt���yA F�Y4!�>桠�
�W��p��ˎf!�d�^n�k�&�?U�j�Т� �.���'�a~��J)C��أ&�� E<�+V؁�yBc�%f�ډ���K�S?40q��ݷ�y�չ&�
<`T���PӞ1걉��yb(@�1���`)]�EL �с�A��hO*��I��~�5	��	������!�d�
8�K0�D�cLa�v���!��8d��L`r��.�^9�p&��!�D��L��֪M�v�.T�4��+]~!�M�!���RQ�Eln���eC�/�!��D��8"�i̝Wax�@�ݸ
n!��[�_�	i��K�riq�8 �Ox�=���
5���v�d�mX�@�VxA "O���2�������b'.�ȷ"O`U{��OB�E�F\��R"Od��¢�8�U�-Q���ʇ"O�-�Հ�%
��d���VF���"OYZw�Ƚ&��#�f�*T��I�"OD�����L�qY���_�D�#"O�s��Q�<��l�7P3`Ⱝ��"Od�q�O1.2-�W�-OB>��G"O�}�g �)����_%z�c�"O愻$i*aP�¡N�!rb��"O"���F��>Jb�rB>8S�la�"Ox�ke���U��p�a��w�8�"O�q�<#VV*�O���y�"ObX�G�E�2x���Ņ-�`a�a"O�V����������o�` �"O�XfNԸa�X5 ��.��Ы�"O���+~,����n�1a����"O�IQ��>K~d�Rc�L��Tz"OX �@�0 H���ޜU�r�C�"O"�xw�C�-˶���6�4%��"O�(S��AD2Re�ٽd��0�"O��A"]�h�� 9��)FBE�"O�!�nS�9	��B���8�my�"O���+�zh�#�oTA H)k&"O�S3���=��������C
2��"Oƭr2�٬'/h�p%�#e�� ��"Op4�@/�-[���A��%Ҝ�
�"O�S�R���a��D�1"OгũW� ��|:��σD��h��"O��Yd�����w��0�.��"Ot�;�Ǉ�1�
̀���?Y����B"O���FA)栰PL�Ny��&"O숑d�!w$��q`X�5[$���"O���U(۹l7�0&m�}<�Ix�"O��rf��,�OKֱ�r"O��p���Lq�3���f5�tXV"O��rc�l۲	r �C�Y2lQ8�"O*�[�o�s YKi�0"2mJ"O\�ȴ�
��@��f��>�#7"O�Z���+e&"I���
����v"O$���n�<1Q�1Q��Xjt"O�*�g��t�f	;�#�<w@@�d"O� Q��g�V�� ��A_�qY�"OF,��Aڲx����g�*+"�x�"O��9惞:��P1��@��^��"O>03f+�*m`B}��Ř��D7� D����W/����H�"?l�I�m"D�4cU��8H5�C�XÚk-D���2녫b.���@N�;W���ɴ�*D�P��E��y;D.�9rFIե(D�����ptj��]��%ʜ�#!�dԺk~ )�@�·dFN�HQAQ=}�!�I����A��92J0ء@I�-�!�d�o���W�ǿo� ʗJ��!�$D2J�*)F����R��!�K�4�f����W�=�f�r�	�!�D	�F)���	�w���8�LD/n�!򄜶�n-�W�G�G��D`r�˱�!��Ly@.���JX'Wm�(�Q�[l!��"�R�dؠQ\��;b�]�!��@j��@�L^!ONH��5�Y�[{!�(	���%4���� {�!�M�F�xQBCމu�n1��x]!�ĔJ��h�#:���#�V'Z1!�dM�kҌ��.L3_��-`�&�#!��?�P��D�c���Q�E &!�1��+Zo�n�бNR�!��>�:1P��Ύ&R��Q�l�-�!�D�(���4��'.�m�Pl��X�!��s�p�D��L)80�Ʀ�!򤛲U*.�"�.u��x���=MX�C�I1.$�أt�@	aw�5cBØ�_��C�Ii|�=j��Ԍ<�!�'"�?�C�I�E����u�x���߲V��C�I�u �yQa&�|�F�����1U�B䉫!_���.qL��Ǉ�dxrB䉊H�
t�E��<e:حkV@�>�lB䉌O�.�
��XS~ĽK���oJ�C�	5rȍx7 P��^]sc�˷Nr�C�-c2J��I�B�2�Y� �&^�tC�I�='b������N�X�Z����q�RC䉙\���&	N�$J]ʑ� &2fC�I}*B1�#�D��x��BU�JjB��
zT��%��[�P��"O�RN�2?��$�%�7mD���"O��s�jֆt�Y�'�E�j��b"O� +�
���`��@
�&hXM:�"Ob�0aL�-���ToT�R*t��"O�A�Ҋy$�`QTI�~b\�w"O2i#���B���(�G�>B�]R�"OJ��_�2�p 4FK�uX���"O�!�P�ZR�=q��R��y�g"O�9��	�t�����!z�l�؆"O�|�s�]�|V�G:N�
��"O�p`�IY�}R鐧�A���$"O��0J�:o��a�GVi���2"O� ��jS�+Č������`��As"O@�Ґ$B7b)�5�0���'���*2�'�'�B��>!a�X�<(�0�Y�1~<2E
�x�<�SF��j��Q��2���#�u�<��	&yx@��(Գ+O����V�<yf
��|�,�EN�/�@!�mSO�<��!K:v��erC���[�x��E��D�<��J�y��R�٩-�\���
@�<�J*wr=P!J�;�v)��~�<Qs�Xf�}�Ɂ;U+<񨇅�y�<� ��+Tc
������m �=���s"O\�8t��9=�ᰱ&�,<&P�k�"O�qq�ZB���AS�=�$"O�5B�,�S�~teɌ*.؄��"O|�����:S�5�v�K���2"Oh4롊@�Lj%H�r��3"Ot9H$�ˤ$δ`
Pi�/L��څ"O�8�'����D�"�K'�( �Q"O����!]7�QÇI�R�"O�)2�Ĝ�^��5���&K
�ٓ"O�бc�����F�_`����"O&��BÏ�g��u�Ȑ�A6%��"O���5��1���皱w����"O^�sCoY�Yz��YUg��HFY�"Oj��f��a�f�a��Q,�!�"OX��"ْ|�� ���*G;ؐ1�"O.9�ǖ�p�ū0��0���"Or)	5-G�tMq�%��G"O.�;5̞J�"���ܠ)i�"OԽSĭ�=<�����X (�6"OT%��d�CV�S�쌸j�= �"O&���Ϙ[1���j��y����"O�|Ҁ�h��*�X���
%"O��Ti���T����[�A t"O>���_T� G,�&��II%"O|�ja䁐j ���ʇ�D�j	y�"O��2F�ֆg�Ȥx2G�0�(�Q"O��AF���_f�ak�*4EJ�!�"O(,�*:&�D��P:
�@X$"Or�+����#M"�8vcAI�zEr"O̴8�O$P������1]��Rw"OtU2i��ZR�D���A}�zD�"O��ҋH�[��:��T�Hqc�"O�qPP��=>ߘ@A��)�N	��"O�t"F'O#w��[E��y��D�3"O���DҤSB�i&.�dv���"O,q�
�*-j񀃂CYj�q��"O���T� `b6�[�yp��ۓ"Ov�"V)��.p�5Z�Ŗa!zb"O`ui#\{&�k㪈�bRR��"O���cDJ�^��#�g�3@E���"O֔[w�=ԁ*cF��WAưK�"O�ЛhW-�e�d>6�D�'"OХYPV"\y��r霅"��B�"O��TeF@�\H���Ão?���""O����@�"9&DrV�3
���&"O�Y�Ӌ�^�P�����&в5rR"Oެ��+�,5V`C4�)�d� �"O4!�M (�j��/P<�8���"O�A	uF	�y�x�2,�"n����q"OR����@�X�	S� ��\��"Ob�zV�I_V��������7"O6�� �$eEV����J�^� "O
��C
�Fp�`�Mӓv�p|y@"O��ѐ@�Y'�Չ��Q�KEr!��"OʙӲcZ49|�T��K6_�%R�"O�țB��*R���pNI[Z|1�"O$J2m=X�4I��qR�T�p"OD��4�ɹ��E�m�6:H�� "Oȩ�6�B��|i���J�2��0"O���"N�ܔ�eB�)HՒ��V"O�9�%N�J���c��9�f}i�"O�$3ǅU�c���p��	/�.g"O�a�G����9HT�#j���&"O� F0�m�i.�h��_T�@aI�"O�tP�C�ď�A�Y�e"O��b�.J�=��+a䛡5qP""O,,R�J��-����0K1��b&"O0� ���Gr=���m��PX�"O� Cs���;pd���Y|@D�#"O.�c�%{�xaS5�� �U��"O�Ē�,�Mv���!$A��"O|D��,i+ !��w�ڨE"O5��$[�+䦑*ԏ$d?���"O���@B$+��Mx��@�A��� "O���H&?�05� �(8+F��"On��D�ǥB'@����:z�H�"OHZ�E�m�HX�H��Q�	��"O�fG9	��9�F�=.���"O�Eu�G,Az
�d�@/��0�"O�E��lQ 4�N"� �`��"O�I�G4B�<��!մ���"Ot�Д/U-$��]Ɂ!�:~$"Ov%: 	M�|�x�!���**�J!p"O�𠲨�q�����7�8 �p"O0HǮN =��b��պ
�v�"OZ%{T,՛5(��rƄ�@k�T��"O� ׏�!z��c%�A>���"O��B�a�(l[t=�ă-(2�Tau"O���� ~ִ;�Y�!�zR"OV�X0%��ab�-9�]8;/����"Oδ�T�5 �jG��HoJͣw"O.0��#u^�dn�"md|�q�"O���u�_�BUR����	|X�0"O�%�n! �u�q�%hV0Ա6"O49S`Ç�	�&��_C4X�"O疴�B��IװZY�a�"O^�S��2-�Xq0��H�=�%"O� �g�X!Ct���65�Zt"O�1g�-�4�� ��.(�"O�x�ĦC���
Jt��%"Ob-�$I�3TJX(p�I���C�"O�D#�# �*Q�G$��t�"O ���	;v@-Pn�����"O���edǣW���Ҍ�E��B�"O�!��ںH�ܳU�'"�m�"O��!"M�p�pykSǮD-�U"O
0�4�{�Bo�L�"O�Q8 ��	0���j�m_�A�b�H"O��X�W� '���$7M(�"O�i�0g�&@#e�ˢV�+"O~Y�0�W��)�U���|��=�A�|"�'g���1�%'��	�ΕMff1�	�':���qȕ&F:����:V�$�k	�'KP�7䆪Ob�4���0R��]��'��SSL��rN0'��K�.�R
�'s�ى5��(s�<��Aqx$�	�'���� �*.p�]rT.�7C�5 �'r���r���@Ϻ�#�/�?���K>�
�c��ܣ�K֎��FEY�[ ��3>��U�ݽ����̀) ���ȓ`��I��1m�j�"B�?u�J��ȓe=�-�$�?*�Mqf�>>��!��p��Y��#<U4���ȱ� ��W���b�<]Ԅi���)U,���Ed���d�Z��yi��ܧ�d �ȓ���Z�@�q?:$�DdԊm��(�ȓ\�" v��c���@�炬r2���S�? "�P�'Y������#Ϛ=��Ī�"O�	��ْ���RF�K�/C��t"O:UZfm��n08�� �v6���s"O�B0�K6�٠�^4"�3�"O�pG�W�Q���+Q���I5��"O�����;"����KׅxX$2�"OȽ�#@әH�N�P��]k�Yk "O�3h�(0hY ���<<�qzV"OB��&n�'�rdQ4aW�h��d"O8�@�-a`�Ж��5-"@|ك"O�ap�H�7���vN� �U+�"OJ�3v�?42�ӊ�\�4��"O��P����a�ԧ	vø�r'"O�}Sw�F�x*�@� T�"w"O������:��1aۀ[R�e�"O��b���8�� ��^)6���"O�(�5��Z]2e�uo[z�@"�"O���u,A+.\������Ig`u1�'���q0�-�.ē�7 ƌ���	3D�(���9?��&�ۜ �e�1�1D��C��F4?�%$�s�1S���	�y�&M�.>�@XA�K�RD�rv�1�y2Ak �u��'\�N��@�B�Ɖ�y��I'B��kH�AT�ٳ!"�y���+@��X�k�&=�h�Cϐ��x¡]7Rp7�N:d
�Ea��&�!�&N�TPVa�� �)ai*`�!�DH7T�݋��X?�48�h��{\!�$D�f��)0P!�?m�<��)9A2!�NBw�#e�׏Bp�xҳ�SF&!��t�J��%kX�4Z֕!)��!�� �{�<�g��::jh���x���1Oj�P��O2v���I�o�0��"Ol�A�&�8{bp(�(,B�)(�"O"t끅��(���bK%K� ��R"O�|#��S![��@Xfg�@�N��"O���D
4(��`�����k��3"Ox�l� �qf#ة	�Ԥ��"OF,b���⎽��"��u
"O��JE��2�@�	ʦhQt"O0�����k9А�ԏK1.���"O>���Ρ�	��OE��m�"OKF�>���3�E�d
��K �L6�yR�Ɋ^^^�K�e�]��%
��y�a��xS�nR�b�3�cK��y�؉�TCw�}�2������y��V8bNw����_ �y­��l,�g�oi *!�L#�y��O�R�����jG�Pjp��ʁ�y�D�t��H6GR6��A�W'�y2�˕~��"���'��ţѥ9�yb
ڼg���X�
�	B�۠Dߎ�y䖌?*p4���ܜ_z��`�!�y�W�9����u'�+4V�� �@�y�%�0� �0ŏ�niq��U�y�4	���)q��H��,rɕ�y2�� ]���aJX�m=�q�v�C��y�՚Kb�|q��/\A�( ����H�<9��`����Ջ]D.�ȓreva��� �h�2���)Ȝ��6����Z6j��f�w`X��ȓ����`#.���Ĝt�8���iVʕ3D�ԖX+1� E��d�ȓn��U@��K� �G�G�����S�? �);s�ىR�FU��h��	%�Qȁ"O���iJ(ZX�$+�ߧf�!R�"OF�Q��z)N�[�k^�s�VQ��"O�Y�#�̋@_��j��
>a��b"OF��@��W�,Cb
Ee�����"OșdF.��<BlS1^�N�t"OܠPs%W:xh�%!�l� ��c�"OR�` �Z
	�H�s�I��r�,�I�"ORՒ ��k#��ZT#�^pbذ�"O �`]���yyС�:j ���"O�1��@	+l�@g��b����"OYW�O�R��yG�� �D�*C"O��� W�JB�����ԕQ���3v"O�p���)X�%J� P .�X��"O
L`�K&J�
ШP/Q'��j "Ox�U��1pT�MX�/W�&�F��"O�-���ݼ4P,�D��mwT8B�"O��ǫ�E� Ô ��[P�X"OH!�vj�36�b ��(ƩkCBI��"Ot�%̘�9s��²g�+jasA"O����^,sZ��� ���d"O���P._�fgi����H��"Otʂ��f��p��S:/e�&"O�-;��[�n�|�C��l��1��"O�8�"#\�m�ހ�oE�v�t���"O`����F�p�C��C����"O�1�j��������\N��)f"O�Y�cK!,=�e���\��}I%"O�`@�_h0`+w��Y����Q"O��ض�؇Q�D�чF�s� ܪu"Ol);&�� /��5)�̞���"O�m�%fL}��Gk�- R��"O��H���i(6	 ��O�<��1w"O�±�\1o��ɸ������`Q"O
F���w ���f�4���s "O2q��#Ǝh��I�4c�Fd�Ҕ"O������nX��9EKW�xӲHJ�"OX�U�Ӹs�b)`
�Ϩ�0P"O昂�e#6e��3cT*_�م"O��3�IF�F�T���Ѝi<|d�%"O��� ���U��4��"Q"
#P"O��F�c�����f�B�X�"O�-9��Q-aFH��l�J�:$ g"O�l����HHBv�օK֌�05"OE�����h���Sv��j�\̨�"O�Z���4�fu��/��\c�"OTU P�'������ Z�6x�t"O�9��9+���ňBKL}*�"OⰂ��+�1�3:�3�'���EF����,�P�(>�<��'�u:W�ȏmc�Р)X�;^4�[�'�F�SA��S�)s�!�=5��ɚ	�'xj�A�^�h�u�;+�4��	�'&�����+�$�H&e�>L���"�'ʄ�d�Դm�Xha�LB�Iun�x�'����K�~=�Y���A+^)�	�'�R�!Pj��5�ޘ*���:.�J���'+��o�Q�[�|TKa��U��'/���!�E�!�ry�'�Dd���'"��a�L�Vic�/� ,�|�
�'�.�T�UnUr����9�	�'�̫� R�r}��uGHuC	�'����d^�F̩��I/g'�ث�'���B�+82��X�)��Y�@�8��� �|�+JT}����٠m�င"OH�X�F�9�vMk��Ro�x�`"ON0	Ł�� ^��#DB|�|��"O֡����@���C+�:�Ӥ"O���c̥E�Z�׆Y'."O�`!��h]���2�\#"���V"O�ـ&/,I�M���,X*��a"O8�f�ɖ5�r9ZE	J+ބ��"O����0��gƟ<;����B"O>��. �ri"0����h��"O�9 ,��'���"c��8؈��D"O<�C���% �D��s���,�$�`�"O��KA��c���QE"�=	P��"O�Yr�oE��s!�J�
Yiu"Oy���X)oj� �7!�mި�Q"O��y�J�E��F"�o;�98f"OjX��f��U��k�斋 ��	�"O�����
c��J�.p8�"O�@CE�Q���@5�Q'89#$"O�9�u�V�+6�Xۥe�?i�!)"O����l��T����ì7�����"O�H�$I���y;&�����s"O���ă5�֘"@���v�r"Oށ�d.]�x=�D���!7��z�"O�l�ԗ.�2ԑV+��>�X@�@"O��X�*N-;3�k kB���:b"O����a?F�����D\Q�"O0���3uO,���.�Eh�"OT�5"�4&�dL�6G�w�Y��"OI�+\�ѷ ݣ0�
�i"O��3iD��IpT�N`n� jt"O�x%��[����Tm�.Y�"�"O�y�$�J3�T��NwT�i�"O4ɠ����LL�	V�*fj8I9�"O����xӨ�YCG>��� �	1D���g�Q�as�U2C�!_���"��<D���"�G�/y"�9ϕ=�t��ą5D�iF�6yjĳC�)Z�r�j4D��B�A��J�!I"K��E�α�4D�@��`A0I���`��Fm��%�d<D� � J߮*�ȸc�����i��9D��:�nC�~m��w��71oؑ�b7D��A�4��1F�Bs�U:sG3D�P�4mٻcì$�2'U�d��jq4D�4ɡ��)}�B�f�my��xw�0D�@���? ��\��E�'*p@ Hg�4D����BB��^�a1*A�B�>�2â%D�
G�ݫs�N��_9�8�K�o1D�8�p��zY�T�^)��Đ��-D��#��ӷ3�4���!��p�s�+D�D;�ʷ7͌My�΃-?h�,/D�hxv��<}P�ܩ�L9� �kD�,D�Љ�b��I�Ƙ�PF����U�D D����oU�)�T[�DI�E��UR��(D�`�¡H_�Xz�b�2p�\�J��<D�@Q2b�'��q)AJ��~  ��j;D�$���'.��1�u"��F �1%/8D�8[�
\f��ؔ B''��ca�5D��!�ʍ')�6\��!�N�Jp��I/D�TI��a��iP�D��>�:��(D�x�ꈿJ̀J�<Sg�X'�$D���an�)#��fG8.=*�s�"#D�Ђ�\q��蕦32�&��6D���	M�j#BmЦ��}_^���(D�� ��Y�A#n������GP8�a"O�)bQ�E01���j�CN~��Q"O%ꇋQ68�^̉�a^5i�� �"O���W�he�B�P	o��ܹB"O�5Sq��9R���H%����<D� +��L��t��ѧp�P��<D��s4sV]��O]0*�����&7D�`�1��1BN\�G\)&����J*D��8eFM<-ab-+�NZ�2�d!�)D��ūW�^�eGbR�l\,�;1�&D���c�	f (Q�5"�_j��� D���b ��&���r��0|Fc�"D�l{� %A���R3��#�J��>D�$
�hO�`��2�@��s������/D� ��85�PT҄拣L�ȉ8g&)D�����H�z>�)�/�4bU�A�'D�|Sb�:2�%��2P(4H!D����G��\f�L���0���4�,D�$�`�N `n�(T)F�*��̢��<D��y�%Q�(�9�G�sa.�q�<D��9�!դl�=x2Ƈ< ��k:D�$8�GB�\�ȼB�*
a޴�4D�i��Y��6N�o��@@�%D��C0J��=� �c��cN�QN!D�$I�$͇6>��3$R�/<R��#!D��Zplө�6�$�ĭ%�hQ�w+!D��c0$�>ɔ19vLC�3j���t!D�|@W��n�RM���b�(0 �=D�$��i�l�h43K#�q��<D��4�n(�UY)R� dx��>D�p�4(	��lx���Z���ҡ�;D�d!�-�d�L�����B�P!�7D��R1� �����?da�qs׀;LOH�@�7��34�XQ��A��sF���v�;D�L�A��)�  ���@�"��m�!'�IF���ON��XV�N.\�*��W�P!��'ŢMX����zd� ;��N�z��M�
�'��]��/p|d�A6���\_�,��'	T���Y�IdA&Є[�(�c�y��)�ӑF:���CZ�F=TX��M�-q C�I�k?$`�	K�LP�8��)9��C�	�IE�9�qL�|:lY��lC�ɸR�࣢G��e���{"�Y9�pC�ɭ�pYqU)�.�m���2Zd��'(1O?�	?gr�2�H���9����Y�JC�	�m�j��T�'S��UT$Ԙ�<�Ip��໔ϋ TTB5�
�;]��� 1D�T1�o	�t��؃��g���e:ʓi�xˎ�=���9��� K������y��]*v"�M�|�Y�с�
E��i�|FlA��&�1e�֙Hg�"��	I���,�ɯm�-�Ӄ�@����󄁹b��B�	 /�Q:�c��բ$��W|���u؟�i�����=�1�����)5�'D�(V�j�Hw��,Yt\�P`(D���U�^3��}PA/U	v�ڰ$&ʓ�hO�&Z�����X�X� (#��RB�	/\\�Aj�
Z$D6�Cb�ϭS�����.�DJ�L�
 D�92� ���u�!�R�ԤI�+"]:��4:�B"�}�'����+�!�&��'a��%�x�� �)D��(���~B4ق$��zl��E�&D�abΝ �|l���J�QMh�&�/D�8� �_.���֕7�F<yv,-D�� ���2դ��!��t�"%i�"O�!C
�[�.�z4*B��
<$"O�[�aԾ'�d)׈*qX^�8��'�(�<Ad���sp�P��	?|��8�HF�<	�8z���@��$(����JM~'?�S�O[6�	�A�^�r�ƋD�1��H��)��<��Ʊ�΁�C�K:sn^ ��RB�<q�ᔚ�^�Q�+W�I�A��ʔ�<�
��,$8�Z@.���bcم�FX�$�O�3R�K�)}�5�%E§Z��@��'��'�i�v����`�`cW)F� q���'�S���C9K��Yy�E��|7�Уa�X��OF���k�-�d��fj�@�|�q�DyX� �O��9U΁�0^j����p����7"O�%��ގ+��	��NNF�4%I�O&Ͱ$/� Fn�8���70�yy��#}"�'������,D��݈��++�X���O������}�j'�� / �CP�D?C�a~U����ꏩ\+^:�H F�Z��v�>�
��P(&$��7��dB�"
���g	�p����'l$��'���
H���ӮeH&��[�PE �[4w;0�ȓTAf("V���/j8`���f���'�a~��>mP������qT��а=9�{r��_�i#��ݰ,[���D�	��y�b��+@p���0k�y�G�D���'���FyJ~UC�0`c���R�����`9&�UV�' �O��'źl��"G���@���WB1Dy��Q�ܪ��%���`Bǀ2Yݔ���g���?i���CRU���
Ul�i7�X8,�V
Oޅ���?#�V-#Ü	Щ�|2�)�Ss �LIe�j( ��z���'&n����|m��:�,J�}, hs�y"�'�,ѺצT�t��E	{��k
�'��X��1�v4��ũ:N��	�'�>��6�L'h�~PZ�C��5�ޡ��'0��@"Q|�4{Ҡ֟*8%��'������YX�P���ة�	�'A�Q�#�.<[�0��w;d`	�'�`�
љdxȅx���Eb�{�o�'<�'�� ��N�"8�
�K)"��
�'�D�(�#�#y�(�_�Hٖ�u"O���e9>���ҧ3*\IJc���'�ў��,!A�<F�
ё%���T�RX8"O<1���x�&@s�Q<Q�T=3"O�ݪ��-3[jX��F!z�޹C3"O4p�2��7 *a��F0e(���"O�h�q�S�0%KkL6y���"Ox�)�b�1V���P�I�;θk��$8|ODZ�(ג(cؙ�È.Hn���"OM�5�οc�\a:#h��+�yqP�'�	D
4��a-��%�Ш��iN�*����q���qJ�5��{��]�g�ȻM>�������|����0$� � (ɳ"O�i�'��*3�`1C�X,m�*�PA�6�SⓥS"�d�a��Q(��Q#k u�jB䉰 �>�u�SM��yc�n<�C�}"�i5>�C@��V��9J�M[tM�o)����f?i�� |��<��ů?���Q��M[�z�Z�RK�4Di�Ӹx���_�O�h[�j�p?��j�d����,�١FN�e����!D���'͈�-pʥ�QbȦ���C�=,O����Is�
W���Hءe̼8�p5�M<�O�Ϙ'�����%X���kg%��7��MQ���1�g�? ���`��:d�� pQ�R�a��٩�:O����� �慪e�>����&+�44y���$>�ĝ2$�+ٽ-�2��K�[D�~P�d�fعl|X�s���'�L=���*}��'�6�S3V� � ��]۩OVc��D�T���lU�U����8�#�eΞ�yR�T�s[>��eC�-��)���'�ў�	�䂔��y�B۠_��"G"ON}�!�Ʊ?����4��*^0���	g8��A��\��$�!ԩ�Ah�c3D��ذ'
�p1�y:��71��9�2�(�	a�'�N���'֒�܀s�Q6=��,P�'�EyZw(�'~��P3��!�S��km3G�!����`�v��I�r��w.E�l��I.�yR�/ғV�Pa���(ƈD��-WO\$�ȓ$4&��#��$r�V��)W#�6}�O�=�bE��(�Gb�C�АbJ^H�<��:`�Xh3���		���)�o�Fܓ���hO�%;F��2����L/x�O��Z�b9�X��.�E�"����6`�!�D�51I�SFD̢m��LPw����'��'��?I�Dd�"�bAJC��)&�aT�.D����d��b��AwANh �G�O�7�<�S�'��^!+d�2�C[�xp�uΕ r�!���`��0U�?�jq�U5=��o-�|�DؖtoH<�a��)#�y� hӶ�0?�,O��1@�Z���X�.A�W6!��"O���-�;+����gKD2(��+�"O�� �'l�}k��N.
�f0" "O8���LUdy��̐t�"O���&C6��5��J��b�I��"O�s��T�y�9s ��e(���"O��sASB>4�!��S1C� ��s"OT(gl��\� `¥�7�Q��"O`L)2�/aH��Eg�&���"Od!�W�s�Q��E�	w,}�t"O�e��Q7)����پ���!�Ó\uԩ�fɑ�)+�Y �ժ!9!�$���p�I�`O������˿3!��=��@R�J��߀{�,��<!�K
{6V���-�*�}SҊ��&!�$�CJ�k�	I�P�0�)���q!�ѹ+&�	ԠE&D�
�:D�`!��ϫ	�����#5.ʒ���<U!�$���֌�@�E)t�.�ʆ*k!��;y��H�R����ZL;׎4cb!�-p�qu� �<�ܥqQ(�7jI!�d
`�L�����$�28�pD(:!�DZ9:�8p�!��{��t��E!�dA�Ww��J3C�1O�Xc1�	�p�!���;8�����;]d^����D�0�!�dŪM�p� �&��uKv���
�9.�!��N	P����/eI|��)ġR:!��@v�LBf��n�\�q��<_�!�dP�`Dp��Ð_� Չũ��!�D�7ij��)��A�PD�v��?�!��'>�[�D��S�� �Vh�>W�!�d�9=�M�#H��w�T4҄M�2�!��	1Rk�5���	PE�����H�!��9��)���i;�t+u�	1D�!�d��Cdlu�B��>u�V�7�!�$Wp�dʥN#�
�Q��%J/!�H�Ʋ�����l�FY(�g��9�!��R;êm*͎� �Zh�F��i�!�� 4���&:rVѹ�LT�!jp��"O0�`�䕃l&��+˄�s�N��P蒌AF@��J9%�R�A�'�&�PnU��"�5a�.�@��'�*��4[����eQ�����'Ȁ�#�
ϫ�N-�U H�}U��[�'h�Q��ނ\��6���jy����'���"��5C������:g��9��'�1�V��&��!�^�g�T��'&�������9qV=i�ԜZC�I#��"��^|!@�̀��C�	;3S���F�A�%��1m�� q�C�xo�$�GW�:�=s2/� 0�^C�ɞSY��s-J�NΑ����7�C��0����BtI�hh�NI�*C�ɒN�0eqehAL�Lp��:*C�	}�ܐ���˨:�oʔz�C�I�s�b1됎��8�$�¡L��C䉿Mf��� ).p�؅�BڈB䉯(\P�,I�d���P��(	�B�Ɏ����Ǚ�0:��J7�X�	/�B�I���Ī&D��c��ʦ�ܮY^RB�I0���2C�=Cf��#�e�(.��C�	2�x�g�ʚJ��'F�8��C�8��Ei��ܤcq�2�K�	ntB�I�d>B)y�j�h� ��d�/�C��&8v��1eT01�Ԡ��'��Ms B�IZ�a�&� �`��NB�I�p�j�1GM6og�l��`� !�$߼pݐű$�֢5|�i���fe!��'Rc�)(��3|
����Z�W!���7<�� 5+	P9K���!�DM�i�x���W�,�|���ϋ6/��~���5��q�!dF�OS8�9C�.s�T=Xe��u�<IA��4PTL$+n�=�E�S��Z�'jV�rmԕ���~��L��p���m.N���Ya	�W�<1�������+kRl��b�#.Lȑ*\_z����Y?E���[��@�,#[@U�ҌD�i�Ʉȓn�HA���H�q�dh���.Ԕ��:��8���'I:���� ͉��O��(�-��O|0*`�C�S=�H��'��1�
��N���u�hY�Cʌ	B�M��oXI�'+�Ȩ@`V.t �lK�"�#��I�r��"�Z��с��X�H���\�Ӑ8$�u�S���M��a*��B�I[~X\:#		K�t����葵G�7�����J�&U���+�g?1��x(��s+�':�p��L�<��%�$Bm I+#k�
\"���B XZ�D:��R�6�����a+,,��;��O�|#�o2k�*�!A!\76c��'24 ��dg�ę��޼�rE.ƥK��]+e� =?���Q�ȠV��~��PxfHa@l�u���C��4��'��1�p��J Z�����r����>�8�Æ�E*'�NKA�Z�G��B��?=��ZqT2�A�5�� _U���à)\iQ�N��\4��UE,�'�~�o	�	BN��㜠G-T�Z�n���=���X���]�ȁ�7�G�{���U�	:������(~�v4�W^���c/�̺+���ã�؉q����]�eA��D5sKqO��s7ڸ'�]�qq'�ŷvG"bA)��4V<QK��8?���q�)� 9x3E�5�p?�򈇇}��xz3`��uӃm�#*�v`���<���7d���Q^,"���Q�n��hs�8�Ī�"Ϫ0���Y@��0p���SG"O��{do[=Q�����b���ŝ?F���u��<I0E`f�
)]��K�/�?T���˟�D�4u:����$ljݐJ�~;azrb�3�vx�r�?i`�u�jd0��K�̬{������A) Z�t�`��Ե5�ϨO��Rb�
�HEZ6��-ߜ�{���E.Մ�d����	�_�-q�h�5YF�z�n�S��1;S)i�9+�G�U쀉��	�$��DBR��1�
d�5ə#xX�)&��F1��"�$JM �����?a4��B�4J��}����<Y�
=��cRk�<�wf�6x��,�vн`,���n̸yb@�׉�o��� �Rk?�@�>OHh�'���S�? �)"�d��3CoK�f�d�I��'񈍑�Ř2B�Ҡ���2�a5�6�� JZ!s����'�`��3��h����	0�<��ФI�z(vu���['���\¢ʒ]�,��z�+X�0�>�@�'���vg�;V	�e���9D��R��Jnʰb0fU�%��A�IW,dJ���=ф�<�`LS�[��Ijâ�3X��8�5D��H�)�)w0� �Dʂ;=>�9��'�K��W}B�P;��9C��CO�<9e��1�d���:f����@��H�<)6�,lhP^ؔS��/`c�!��b���+sC�UY��XKA$;#FA��p9��%�B9�Ó@�'@N��ȓ@�|m;uH��|���#7��2������R�`q��j�x��	��,2Uy�#%�
ap `�!�YÊ{"���c�� uX` �ޟH!wI�;IQ��P�ᖩR�D��)D��C���:�>i3w�,�us�q�ܼ�G�&o��7��9a� [��5:��S�S9i�ȵ��_�-��A#������DK�o�T���C#�ybOK�����G�� ��{�+[��|;���~�ʓA``�|�'���6bʠS^*!B�χ
�yX�{�gC�(�"T�Ht�O�p8r ̞v0�a��a�e��NǢd��١ǀ��t��d�O�iP(ׇ0���ٕ�"���O��09��O�lj��V�mf��T�i'lz��F�4H���F�����y�'���:#��*�@��-�VSB�-p:z��� ]��R�T3#���:��<%?5��l�6Z&q`��¸	�t����=\O%����(���q�'" 1�$�6wW�ٛ����{Z�y�B��D�IC7��<�r$9�gy�_��8�T��33�Jt�'�����''2��@�Mt���D�DJþ,� 1���+~,p�1d�\;�6�� Γp����"7lOtac'���t��U��n��'f�	s�׷u���[�߅z��d���'{�^,R2&�3`v����S�T�	`$
e�T�� � X!�Đ�B>}1j�67�ZŢ�nC�"�F��&-&L�æF*Z��a�t�!V�8�O�i�O_����j�#-R$)��Ϥc���3�2��D*I�pX���EE��IبD���4+���9F_0vV�B��!X�ԲS�_�h�qFBC�^�=�3�/��4��7�����%�܇y��LI�@!$ވC�	�Ѵݠ�I�)8�$��T�+�z���y�\��ӫ���)�'m�.%���a� �r�A��6��dJ�'g���	�
����ï�&�tC-O,�{3�μp�h˓0�~�C�k��Nd	����'ꖡ��ɭL`��	%킑j��V�?�H�&�	d�ʉ��NX3����SO��sꛭ �*�r�A'(���*Q�x򂃋LU�ţE��9kZU��X$��O�ԍ$���0����,[����	�'s�|�fo�"}��=R�B�c��TgK�i�1�'H\�� ,�.�¸O�'k���(͖[7�W�.E�.�3B�,�<�sc��rr�-F���o�8O��A��ߟ(O���@d��<�����8���HB�p_69�R�ZAA��"qh�c|����	h5y�� Kd���K\�LOڤ�S�@���(
QE:�C֛��Q�����z�D�@T �b���H�D�!�4��ɧ}� h�Ֆj�>�ڢ�S�?VP0��dm��ɔ�o�RH�gA3D�t6�C�	`�/�FL�wC�(-y���>���WV�d!�k�.
dqO�n
�)ڬQ�n�;�j��c ��S����n�v!����A����O9jN��*B.��תE	���q�jҶ(D�D�M�Ffh��I�w�����6�p<��M�9$��!��.?9r�Ƞf�Dh���Nv�D����R~B��>��x��4\��dc:���H�e	�8NO�œ�ċr�O�ӆ#�mZ#3���C�T]©"C�1	LxB䉕	�r�ڂ�	���8g��#L�JP��{b��&d'��vј�a0+��l���@19���ȓ�J4�6�ޟB�����N����'�F�����yWl�b6����@9����'q�����<To*��UďE@jP	�'��Z�՚$;�p��dC�9V��y�y��)�J�%��Dߠca�haJ�	�C�	JZ�(Q����L���Uƅ|#<�ϓ��]��F�$7�T �h\Z����S�? B�Pvnڽe��˔ �k���@b	$4����=>�2D�u�U�iz!F!$LO���r�� ����'�QS��� D�����Q\n=S£B.^����T$4D��K�Á=g$&����D��DO5D�LPT��u�Yp5j�'Y\(�b�>D�D▩^ w���6��0�p�B9D���u� j�ʇ�͇o��Y"*=D�p�L�M���wI	48���S&8�O�	���~��Ɇσ�f�@1'£X ��'�EhS9e�j� �#3>�iN>�#�~¬@�@��9�D�|��J�4dA‒=�d0:W��/�$��	a��u���>S� ���9�$=*����!�"�LKpt�s�c���� �<D���5f�=��c2�"ԣ�+K��O��`C����O�@أ���lx)@"ȧ`ͤU��O�����ŒJɖY� ��yq��!�@>�4��m�!�SvNi�A�H�n��0�t_���êqA�'�e E��F��'Ѥ~�.���J��E�6��HMw�H5:e�P�&��QQ��C�,��LY��4}��i��|���K��^'��\2��Q2�V�\�R,�'�3J�����cPꙠ�OŒ\|:5���4+ĳL�T|h���8���%
���Q�P� HB�@���Od�e'#l�P	��	�'�^�c��L�s��#��K���,ľn��Q?���X�x*֌!@��xH��Bg/"������E�
ܱD:8qb�>1b�����(vv���$�';�L� �+ĸ1��,�e��.5F"a��8OF�#Ӊ
]<��BC��'<�R�P��y�ԟ��j&��||�Q��>$�����,d�i���F�7l�D��"1��
�n�R"���A�$�N�=Zq9�/�)zB��F�ŀ�@ӧ��Dx`�Z�J�I���Mh8@�∥�\r�>`4�tj�1O8�1��§p�(�k���l\):��m𕌂���ɵe���W3	~Vp"��חа<%E]�� �p�Ax�y�� �<!����`�A�$xɦ�J!�o´I��u�
;v��z�ɇJ԰BI
�VoB]���>�OFM�b�_�2�m���8IP�-x���;?�Xh�-��~B-�gr����i�m��A�9HQɧ��ʟ2��y��E66\���AF���O�!�Y�_^�ih�O��H���F6%y��V���JU�"TDy`�'��xu�Ii�S�O��	�X�;�1�t,�%5G&X0�O����/�a�.�O�>��s⒂'����OϘi�l��)1D��y����)�y$JT�V�G�.��U�R�˓
g:��`��~8��C�E[
B>��ȓF=� ņ�F�>�[e*L�Z��ȓ~xA,D�!%D��!�6�T��ȓH������N����T� �T��чȓSY���a0W���P"��%��+X8��l�S~d#B�нB+�!�ȓPvN��O�&��ђ��	?-FH��	���+4��->�d�:p��9Xh�ȓA���ȉ��cP,F�_�,���x�#ef�^��'Ɯ.r�0��*}d��;?}�գ�@�f��h��I��+��S}�J�;�H�`�(�ȓh�Di��F��=�a�
|I�ЅȓqW� ���	���UxD�B&(��ȓ:��p�W'Yc������%���A�U(��M�1�`Q!��& B剪;n�$!���2=Jؙ�,��l>D�؃����{���"��Dq-�1;�?D�X�d��Z��d{d"!z=i�H)D�$"��ǚ<�X����U�52����;D�������4xG�9�J�@�ȗs�<���#oߌ��*�ilpyPcBD�<cn�)c�����[)o�>�3�+�H�<�5La�ͫ�Q!
jl�I K�<�c��26qpb+W����Б�FG�<!�g֜N��f�ܙd�	P4	OA�<)����\�Ru!O�1�8�+P�@G�<�o�t|3'�Z}Z�I�u�F�<�%s���ʑ�(Wx$�2��z�<Qï�
�����JH&�����
r�<� �p��2��p�f�:K��M�"O,�1@��P��s��K��ҡ��"Ol��N�o��t�s�!|��b"O��R�AX)f�ؕq!
%��"O
yK�Z*L!F%27;_�2�"O�m�2́)h�hbi�	�j��A"O\�����,�@�]1Ko(�(�"Od��.�Y�֌ �eD�uAd���"O����+��Pw$�&OW�0)`"O�-��G?%y�L�`c�:A4��"O��%O�}=@�C�!0�a(�"OX�S$H�25�`��"�)(ȡ�"O����%� ��U���k��"O���6�aO�h#�[�M&��!"O�T���_-)DxD�Ԭ�!%n�*�"O�ju�W�mKE� #څ����yR��.0oyR%W,'�:��ꃤ�yb >(/�JF,/Xnij6O���y���}6� ����w��&���y�%�)� l�b��)�ċ��ɢ�y�1]��C.A�O�t�%��8�yr�ʫI����k���Q�@[�yB" jDޱ��tݲ�U� ?�y"'Д8Q�2F��n��DY�%��y��E�&4�aJG ^�)"�H�^8�yR�ٿS�&5!c�%�8��2�y"ɖ�~\��@i��x�+�)�y���5�V���۝| @���O�yBɏ+&�ԋ2O��v�,l�K�yR�ԑ޴�x���r0佚�d)�y2掼nR"����]x��2�A�7�yb)�L� l��̋9�D���C�yRgɀ=��<1	"Q���yb�/n�h��%%�l `��y�π�y�r�7'D�y,�ා�2�y���4鰁%Jެsxʝ $�y��E��,B�B�4Y���:LI�y2�Sbd(aR3M/]��i2�o��y���	Y�2�3�à �fpI��9�y���=w-Ra�i�Bm�!-�"�yJ��F[p���ԅc��U�`g��y".��)M2� �ҟc¹�0-P��y�[4����C�g����铏�y�k\�;�|�@�
�
���ؤH� �y���*��10��U�t��8˳e�y�D��:Qbad���z?
!C����ybK�$h���VM֏h���X���y��	K�@9�i�4l���#t!��yo �CFT�2�$E"�����y��(tnpM�ѷ"���R���
�y�,G��ٛ@Z%V���J���yҪ�� �\�V�Y�<99��Q��y-��D:��CN�9�0���yH�l��LN��$=Y$C�2�yr�W�;UѰ��t�H��s�@��=�N��;|�W���N�n4D3�͖��X��	��c��!9>���L�2�6��=iDHtZ@؍���B����M�1x�ȃ�	]!���9wK6�H#I�x:�
t��XyP�K�����	��"|�'2��)�$ׂ5NL� TY ̌0�'�0ژu��� ���$�0}U�� %�����@x8�TY�kU<�:���	O3���&�6LO�L�$'����Y��'�)RЬ ���D�0j0�P��'�4%e�b��<��g����y¤�
b�ꅳ���p�π �I���'+�z�Ç���:��"O"��*��S� %h&��6K�(�0��O�\\+M�X26!?�g~��˰��M��ʠs��;�fʉ�y"j�!*18�f���,}��J:L��ePrᓁ7mα��IN�p�R��}��2� �%|x���D�	<KT�c�B���~2���q�0�S��Ҏd�H=`��С�ya�0W����C��P&��A������'Nְ�m�	��?�:��:��)
E��E�޸��j/D�X��,��I���
E�C��(3_�X�="�>�#Wa!�A%���yI:D�gM
a�<���9��E��K�s~8m3�]i�<I�ر\�z�*��7`t��Zg@�k�<���_m�N}p�A�&�@�;���I�<a�D��2��u�۸X�:��^�<F��<2��)������P�Z��B��z��)1 �Ц���x!��
%�B�	�w�h0���M�#�����%�;`�~���*��+�)+�Odq+�DXTB%��C�?b��Yc���s3H��=�O|���Ⱦ`��MC�o�O��y��"Fc����Z1ex�4�b"O��Fj���jL����Y
��c�i�L]��bV�Hs��(փC��D�#�ڨJ��)�	�$*��2c�lH�I���z�`[�z�H�˲-��<A�HЉrOؙ��K� #�r�ˤA�1@��xW����	�Q>�n���Zfj�0d�("�.C2��H�=q���rt�P�t4�'��l�"�@����-��زp�'y,���$Ș�a{�3?a D��.�8O��i�,�V�X ��� %��ɠf��-2�AW'��G�Z9�4Em��X��۶tg�|hm�{60��ȓ�~}j$��
����0 pm��h�I�C>@�� �L��}P�L��`}�S���~�1R��������ҧl��H�'��(�4��-9	�R��4���Y�$,�"��="D�aU.�4��Y��0��<A�#Į*w� h�l��?��0���W�@j�T�ժ
�%r#~��oF!<�H}Bre�1Z�%p�L�h�b �3o�'P����'w2��d�!5D��H��-��U��C�MO\�qĜ�~��D�P�h�b�aa�'��}aB+�!B�E5�[0�&�8�'���q�@�b�x���+K+%m�!C�4��-0I>�d��%U7ǔ�)dMc�	��T�+
��$i��_�FD3����{k�{�(�4b:��F��(���B�C�F]���%N+&��b@mH<9rm�o ����0rj@�+w��_�'}�D���`(5�~Z�
W�pw�U)�\$�����X�<)t�ô-��X��C�\�2-�R���D��k�.�⥚>E�4-�0_��i���-7�����%ϐ�!�J��e��苄?��]����7��$��
u")�V'���<	B�F�x@�$B���R�]x��h`O$C���"���6<4�x�H!mY[��X�f���їȁUn!�dQ�t����s�ҍ|.K4 ��y�'��L2��@%8�<Z�ޖwt�A���d��=%p�A�CEV���ʦ���y2� p�)а�fA�6a���U��p�1��"F#.h;��+ܸO�' <8�va��'v��`�U�g ���'�q��<T_H$��3u�8�Rr��9hz���Ĳ :�({�����<� 
��[�.5��#V(і�j��{8����
�^� Xs֪��c�:��3f �|��y�2��	�ň�?�!�Ė
Hf��t-.y漈��\�	Y����#�>���қ���!�E�f8(�����!�;
_*�`C���=�rq�e �>��Е>��J L��>�O��b�'!���S�ٖoIb�;�
O�U���^�G[&l��Q�R�6�J�샵k���(4��'�0?*����k��1�
��D��v8�L:�o��e��:𓟔��L�R 8U{P-��{N�p�*O�����AO���R$�/ �Ǖx"�H�4Z
(F�|��d�ߗq���0lK#$�(pN-�yŔ�L&��B����v������$�DL�g�D��z|DM��KM�:֍îY�!��:F��t��,�Y����P�>�!�
*1I�5C��?.b��m�!��̄s|�UG�3z�f� ��0�!�� zM�r�
�����Ƙe2Lk'"O��S&l4;�б���	*�5��"O`��[�Q��́1CT8s���"O.8 tD�	�vH2�HlbD�"O�t��VEӺ�SF�'dN8�"O.�)�h��M��P�#kM�$]zD��"OA�cC+-9b5J�*�* ���"O|H*�E�<
p"_�]u`)Ic"O��L�r�FE���dPl�U"OP5IbCV"r¬�P�C@pP��"O��R1��5�t�u��v�j�I�"O��b�Z�����S^����R"Ot�k5,;v��rF��o�Ԕb$�'����*��x/��2g�yI����O���{�	��j�WN���ٗ2�
\E}2.�!)��a��i�9,��)�9�Cr��TX!�D2k+Z����Lp�"�T�2H�	<�l`k�7��)��3J0)��Q�Hؤ<���  �2�U��!
%!�PΔ��(S
{E��A��V�ɦ�4#f�!�2��Aj�3?�i&���>cG� ��,Q= ��{��-L\�?�#�E�:�[���l�Z���(6c	+7j��U�!HR� �E��c6��J�`��\�S�O1ƹA��]�w����@@�b����]��U�/���pk�D�i�*klv�>�r�N;Y�|���ڱ �Xy'n�<�%��1o�f��"�=,O����Y`.�e�1S6�يT4O4���f�X�Z�۬ID�'�F�jF6Z���[��K�v 䨀*�h�"5sfm0�P z�1�\ *@�� ��(�%�%/E#�G�H"�:RHk� y�"Q�6d��`�, ����^����?��*J�<t�+䨘�n�\x���<�{��|��'�3A���i�_ (�gj2N1h�s `�0�4�{��B�0�=�4�ƺ.jC����)�'	H��5�L�rb���闩KB��'d�y���D?K�F%̓ ��J�fX:�T�>����(L�����ٯC&ȕ��Ƣ<�S�Ra��*/,OBi�S�_��EK�G�}:Z��!0O�����5�n��g� �il��Hw�F�38��P^���Y����[�|���F#"ܽC�&НP�����	Ň��l2�ǟ0X�����h ���}8��m�����BI�G�i>�X�ŤM���q��C�4V�`*��!�5ZZT℩ܟ{>�DT�Ѣb
%(G�!�F�F8<�Z����S���Ij�l�����S[B��"Pa@t����-�2�
2����]���S�O	�0 E�b���"AE�yf��1�'v�ECv��J[�A���r]���N>�šs_���dB7`�������{�蚃A~!�$�(2�D�R���^�,��uA1k�!�D'7=pTKr�����A
�W�!�$�{�tZ� %aɂ@B�V�!�	�"%�wOZ/�0�o��!��6cSB�QA�_6f��Q4��6�!�dE8H{t9��T>a����햤�!��7O�6p���	qgDh�K9:�!����(��&WR�����Y:G�!��a=,�� ص6w��#�#�yM!�DL%�����C�xt��2$��'#!�ė<g�l7� �G3��XP㗘o)!����(�P�H��8���b(�0d!��O0(FA����2:���S�A��!��P�8�B@'�u̔��Ꮛ;�!��?y�Ȭ�$kĉ ���RV �e�!���<{F@�buC�� ���`!'�!�d�L2ޑ;��[�4��� ��S�hq!�51j�P7劔H(����@�
l!�d��P}�E��
�qR��C�N��!�D��2�2��4�Q�	$I��nH3/�!�ϖ}���h���#4�������N�!������bo^S,0Tr[\�!�DE �p��J.>A1w��!�!�$��K,�$qw�y�i���+i�!��Fg>�Y�ׇ.L��LS!�!�� ��dsK�9��F�%h�$�"�"O�󀝶K�L����,���C"Oj���)F�;�Ta�O��v�P1"O�1B�g![��U9Pm�{��л�"O�q�6`"*�X<J��L�h�:<�"O4���.���˧צ\�)�"O��i��Ƌa�@0��HI��.���"O �p��"w�.@�Ԫ$��"O@�1�kL�Je�A��A$�"mc0"OV�b��w\mi�#��
'"�9$D��lA<<����a)Z$Q"p�;Pb�0{��O�SU����2(U�Ah2����4L$ Y՚>�Ƀ�!i�L�|M~�iLeRr��ӏ�-M�.��� RB��_�[��YH��A$�0|b���T |����&Ul�j��|?	�C��6�:p�6}��� �5	Z�iA)��,���J��+<�S��U�@���>E�t�J��S+��Q�d҄ș%1F��j�$>� <�M����.6Mp5�ᓬL-dD����=�����#!9����b$M�-�JK�8�C�~z��)ϵ�n� �J����Q��%8�X���R�V�q��]�>+bDP�S?�F��ɜ[����R*
 IZt�	�I@��?��

�,����e@��)�GҜ-{�L�\%x�	���X�Xp4�2�}�E��p���"�f�[6�K4xB"l���Ǩx�A�>e��@�7�V?1V���L�$��@�"�lT�MNR���P�@��� ԭb�D����t@�~�	&�I�|��)FT|���umn)�1_�4���/txY�۴R�a@�J?֝ݟT�l�a��}��JV/s��!@�J~Ӕ�)!��`j� e��]I�O��Sm��T��	��լx@>�O<AJ�+Y��xn�:�PG��)h�*Tk@�@6>�"@�� l0�	� ���i��Ȏ���d��B��4,�j�N�gBҊ��	�nԛ<�?O��AH�<t��wl_�)o�Z\�|��h~�a��F�"D�E'��t�>ɍ����D�<+�(z��%O���k�����0>��fķGpe9��A�0�,�`i0.kDx�a��+� ��C��S���`E��j=:E%2�ɚA�LU��S�w��eZc��;���bP
F(�O��'� ��Hv˧V�$��o&b$V�V #����F��8;Jr�'�l:���l�����>﨟輨�.۾4�J��b��6i>B7�'��CÍ�*,�ʤa�Ɠ�t"a���ֵ
��t٣�M�h��y�Ҋ����h��}�
�Jf�qP��ˁB�xS6͇�D1xu��?N~Lb��؊lZ����)�d���ujJ(�A2)lZ}�ۍo2Ɇ�����r�˖���P�AS�6u��Lj�
�dV�Wy����
?�D��ȓ^��)c����LW�T8+��C�fD��`q�I��O$�P���	;>/&���OD�@�-�8��d�7�2%��]z����&`M��PîB�Tơ���e+��H �0�kG�!��Ćȓ]��'�7l��Ҷ��gt���>�\�':SeL�F��?^z��ȓUa����Ί�p�H�fE
��@`�ȓ�H�SSi�zP� �P::���C�^�CtH�M�����A]2.8.Y�ȓ���'�ӭz'&X�cҵQ�J9�ȓ \�}��Gεw�ACA�\�p�ȓu#jm!#�1v��DCƇFK(�ȓ	���{Q�Z�3�`4�p��o�,��ȓ]���Al %ˁ#J�%.���p���cI):�n���"R3�d�ȓ���0�ˋ�t�Υ�t%��-��b��]8q��XDpS$�]	�͆�L� '��p�������Xc"��ȓc��,�"�ޞ+�<I1$��,ex��ȓ�e�a�FH}����fV�]jņȓ"�H'�J�Jf���uL�:F����X���)��#(�!�"GW< �&̈́ȓ3��\*�k.���� xp��S�? (�#`:6���ِHƌ.�ͪ"O��vE��A��QBBH@0��i�b"O`�[��PP��eSe�*���d"ON{���a~,H�W�+jd�i�"O�av�)=��V��-�BIx�"Ov5����a��*��w�����"O��a� �`=(���	�.[3�y���r����c	H4�l����y¢�'`��
�ʝt˨1ᓉ��y��@�������aI�U�r�T>�yd��L��H��� B��8Â�̖�y�'[��D��ʒIU�8C��yr�סp^��d�A�@�$��a����y�j��7BPh1��7h�ݛ!l_��yR�҇!�8�0��_�,a�9@鏁�y"^!8�tX�G)���,(�Pn�0�y���IHbY�T�D&z�vؐu�M��yb91�\[�b��ZD�o
�y��>`
Ⱥ����"�L�Ys�ʊ�y��</�Չ�E	.n<pg���y�&r�� A'ȸ_�$�	U�H��y�3s�1��	͔,Y�<����3�y�tb��!�������/]��y2� ��l��	��n�n�94� �yr�}�B�1���f\Ą�I��yrǤdL���K�O8�))`����y��P�鰤��HB'L�h	ڒ.@��y�g��g9X�pK�:���/W�y"*Z" s@X;@�RW-E"�y�OL�p��{��Iw���y��	G�&N�z��|���_+�y2B�h�r�3��=��2&���y�'M�>�2I`�O�3;��P�Iȭ�y�޹Jf
�x�䈧%@���Vg�,�yrj���s�J}�)�����y҄��7��1�!�;�@� Dᘰ�y2�M�D���0M�70�E@���yR���Rd(J�+إ�u.�$�y��K��<� P(T�o+�Up5Ȃ��y�"�k�F9Jq�C�c?j$)ƦO��y��!�viI�⁻*�2�զ���yB���`�|xҠ+hH	E%���yb��{>��H�ۺo3�m��*�yB�o9Ry�cM�9j�H�C!���yB�@_u�U���aݮ��B��y�6x��`�LU�x\	abD�*�yRhӆf2���eӺ6g����dҥ�y�X;����BC#,�(!���\.�y�8m�������e�֬܈�y��:��A���t4����y��O"�R
� �-`�N5�A����y"M�*R�8�x ��
D�Q�1)E!�y�Cբrj��6�Rx��(��y�`%2]�����(�$�I�K�'�y�mN��������Z�qa'J,�yb�6�|s�DX�0��s�̏�y��ܮKN�	@�1�6U:�bP�y�J�^��'�8?�jXB���yҏXK6��(�hC=n�x�Æ�7�y�L%M+�;�/�Z� H �́��yr�It�.� �ũW2���*й�y��\����MKU :�������y��څEl<C&�E#}J��'̔��y�	�R��%��'S8xܔy��	��y
� $b���X��k��[9�ִ1�"O>�iP\A�5k�C-\n�a��"O�R�e��h��䡕���t\��1"O��;P�؎zMĝ�6(K�H �d� "O]�3l��&�zI��ң"O�kS���+|��s���4)��"O��rf'�'LBtɂcfR��U�&"O��(� U�C�Tu�S	��
�"O�qSV�����W��~����"O�����8�P,�6�	��9�"O������%���g���*�I5"O`�4�G���٠�bD�w���5"O�}�5�ٶ[L��y2�)�y�"O��"ca��2l9vaӼ)V)�W"O~���M&R?.����T�z�"OfH)W)N�S��d D������"OU�2%C vm̅����%�^��"OɛN�5H4��3�]�TAn�w"O +r��PJ؅�b�ݭ1�42s"O�q
�扝w;K嫐��Z�"O�`�V�Ӏ7�d�4���*�dL"O�u!��Xh��aM�G��`"Od�B�">
Za�j��b;V���"O�E���  Dz�oL+N4�u�"O*����.'�:���Ͼ3���""Op=��� �9"�m�JR�$C"O���`��b[�,�
K'h�Q6"O:h�U
��W��$�P�̴ 9\�@"O�<����¥�T��RP��S�"O�U�E�Z/T�M�Pb@�5����"O8�"�n��`bZ�q�BX�`9��"O4=�0▐V)2$c���p�8�s"O�d:�BƸw^
���]6[Vvݐc"O�\� ��S ,��E�+p���"O�[�c߄)}Ȩ��c��X0�"O\U��[��	�bB[�8�=X"OP���bOزE�G}ܝӣ"O�����������%΀�}oVB�"Oh<�Eo�$�@��*�3r_(\�5"O$��r C>����@	 
�x�P"O�4`�Jͤd�ء���6�@G"O��``��)A��B7��k5�(�"O��x�ǅ��2ex�L��w����"O^���Z�T�ܤaQ�V�uV��c�"OD��bH�}�r�P1��j=T��P"O�A�ի�1�riQgFC�uG:�"�"O�Ir�lF 1��d�
C+!��i�"O���+ X1������b"O��l����ɶ)U)%�
i�5"OR!g��0:H@�
Ȭo��D�Q"Obe��섳�����]�wκe:u"OT���#�*Yv�����N��x�"Od��gݨ�l}HA��<q��Cq"O�Dz�E!fY���fd��k��y�$"O`�җD��<�\0��ɽd���b�"OHɉ'f
3���t�̡in�� �"O|����׽9��[�ɓ.[�Xp%"O6��F#V<I�j\ң'�/@Wt���"O
�+CK�F%�PF�]�8YS"O���� ��q�"yq(7~Q+�"O����P���F/$�yV"OZ�r��J)&����&��7��D+E"O������|e�4y��pwAk�"O�#�_T�q���˯FEu�Q"O� ��k���qh)����04QXd"Ot5
W	M�(��q�[,#��H1"O�9��є&�vh�&�pe�t�"OTxf�:��	�� 9J��Q"Ox�)A͏�y�赩����"7��W"O� A��Y��
ҋ_	��R�"OV9@,B~���sT�N.��	�"O�ų���:F�1�D!��!��"O �A��̈A
������Q"O�|8��J�i�p�!��O=	�N!Z�"O�RpEPvA`���(*l�܉�"O�=���k�P��凗)>�-�"OrqRf��+: 4����08�iD"O��,M�i��+U
&��6C���y���$j��	��Ӆ*D\1'��y��ռ
EP�R�'l���5��(�y�7f�H�2큼m60��,��yb�^8VVb�b)�0d |�	�b
��y���̚%��Ƹ���O� �y�(�eL�	���Ѩ�3�Q�yB�M�L	�)RL�< h�"��y"�x\��0%�!a>e�!!G��y�̎+�n��c��щ��yRP���H��bW�I��ba�-�yb��ZZ�C0+*FKJ �E�:�yb��6hW��C�DJG1���c#��yr,�:�h�c�B-P$!���8�yb	�*2D�7 ��At �����y���";gT�X#�_�c2��� g�2�y")F:Uľ(P!(�_��R���yҩN�7x<�bo��Q{��( g��yR�N��x�A X+�d�I�,S�y�m�Pز�k��`���X��y�Ό�1&�`j�g��+	��RW�M$�yrD��zNR��!�FaA��yҮ����ӥ��򩂀O�.�y"�C�>���
�$�����,�ybo� ������R���Rb埂�yR�?�Թ2�E�8S���f
G��y�HG    ��   �  i  �    �*  �6  UB  �H  �Q  X  J^  �d  �j  q  Zw  �}  ��  _�  א  1�  s�  ��  ��  <�  �  ��  ?�  ��  ��  �  ��  �  L�  ��  ��  ��   ^   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.�T�DxB�'��PnS�8�2 �f6Q��$��'#j��G  �?�	{7�>� %k�'A�)0�˲e!>�i���%��ə��(Oz�J��_�c�q7(�4GW�ȱ"Oр�Hr�́a6-�E�	f��E{��i�dI�hSm�?�4��Ń�	O!�?�[5)ɂPɌIP��vY!�D+q#b��@^����A�芢
I!�� ���2iR�7�`���R�/PFxe"OP���]���A(�1�4AV"OPձW
�=~�����T�Z�[c"ON!)�fi�	5 �H�4 ��d,�S��:6T�����x�d@�PoxB䉆��i�7�Ʌ4�0�sl."J�"=IǓ�VUP�͎
#nDc���0���ȓu���Т�1�Рxԋ��B�J�<�指�$Ҏ�3�Kh|Y��B�<)��ݧ|@�����E�D��v�<��胹����g��>6X]tg^n�<a�B��m����w)�C�ɟ��b/��C��Y(�r4b�O�����7� ���I��&�PU8�.�x�!�F�3@(�Q�K?<�X�pG+1��	@��̫7�\�Mİ��nW�_UTyKa
-������~¶��k�%^��L �f K"1m�O(<���S��3F��e�h`WGK?i����n�NQ��N��a����$�@=c�C�	�EP
���cJ�z�̀�C��_;J���<��'����O�3�I9Hj)�.@P��5��8<�DC�	� �y�cbN*B�{����M�C�	o�������9��%Bm��Z%�>��)�#Q�����g�^,ц��[!�Q/�$�p1��6a���F���!��1&�̉�"��'�zDBcFM�	!��H��Q��Q�qc�;�$�%7c�'�a|�O$�4��&�Et�2�	/�y�F\�r8bf��st�4�p. �y�G�2:Ѯ�15�a�2,@�I��y!U�p�n��7��3Zcb@c2ب�y�K��*��U�N�`V<������'�ў��ȍ�E�Z(
��2�Pc"O���R(�/(�z���_�{��hB��0L��x��;Y�ȍH�*W��4����y�GO1�DՃ ��2�j�# 3�y"GL5~X�"�<��H��yR%�|����!5��H�숝�y�埕t�\�ƥ�GfU!���y�&֗���9 �O+D'��R�b�y��<s�|y�T
E�?���rʔ0�y���lV(-����%ېP���	�y�f<V��v�T#�����2�y�윖t}HI��/0_|l�e���y2'   ^"���*E#h�RqoI��y� �60 ijQ�>�>���H�yB%�s��h�V���=�V�Rd���y�G�7<0��!�mS(*B�PDB^��y���xQ�D����a��Q�y���9P�Z�����ty�F��y�M�'e�\���R"����w���y2�.+��LyV��~�@`�!B��y�b�2���zb�3.qj���)��y�C�=F�o�#S88Y6�Ƴ�yRE�t/�@��<U@����U�yr�٩,HY9�#I4W ֨�d�ݰ�yrB��Cl��uiO,{����ʑ�yܑ*vp3%'��K��P���	i�fO@LD��0��ƛA(��ȓl���ce�}�ZP pʘ1q�Q�ȓ4 xI���c�,��D���A�ȓ *�m�(�� ���
66m�ԇȓAW^�2e���5A=a!�� ���J��!���l��������S�? H�ق��"c�����s��!�"O
����M��HP�� +t���1"Ot��c��'O��	�B � ��kg"Oa�4G��T���dI�$2�2�"Ol��Q)sN�c����'#�-�t"O k���,b&��5<��t"O���T�#$?bl�g��1��� 6"O� �pa¼�0|Sp��03��Y"O"����|�����V�	���%"O.P�b�ۯ/v�����k��c!�ڂ/ov�AFl����I��+@�6�!��u��x��d.ƘUʏ� �!�dW!=~ �����]%0�(��:�!��C�j�C$)Pa�G	�1�!�D��w�6���p���(���C䉆��x���X�	�ε�b�EV��C�ɷ<}��;0EL�j�	I3(ޗW�C�	�|���v��g��-���APC�ɭ\���C�͊�4����˸ PXB�I�(u"���dDP_|��R�ɋJ&�C䉊5���*���T�DmKJD|� B�I�t�xMz&��8�.ٺ�IA��^C䉡/�n�.6d%*e�@> }���sSD3¥�O�q�/	=z����ȓp�\I�E�P\�сN7n�� �ȓ4�zPP� ,"�|����.]�(��V��VE�$��2�%
!}��`�ȓ�2�36g�"v,��*		W����t-jv�1�2����񎔇ȓk��
�eׂ5�����J��X��Yv���N�w�
���Z�;{X�ȓg�Zx�5�N3�f���#L�%����#�����J�J�b�{�K�3g8���Bq��t�	�=�N|k�H$fK�H�ȓ
�B�Ba�D5r�(e٠$�B��ȓ\}L��Q
K�G^��Xp��#��$���8-Q��جJ��U�¢n'�y��`��@�#�^!v$�7e��(&���K�ɚc� �N\;g,�<a�$����,��Ǡb\�ď��s.���S�u��O��^��=����?q]�݆�!.���U���җ<:U�Іȓ�6���	���R���;y��L���������h��e�tQ�ȓS�H�2�c��Y�!`Za��)�ȓ���)�I4�"7ɔ #��Ԇȓs�~�#�/a��┘U�|�ȓO����Ȓ��)c��>Y.�ȓO��|��]��`q��5�de��k��x��LāG1�LI n�Gp�X��\�V5kd�L�6�:©ݾ='����\�T�؁ŃO��P�$�Y�?�Lx�ȓ���ů�*~Pek�f�6;�D��ȓ1����`^�zt�	[u��(�>��,3,=i�ą�\�*���-�=��G(a�7�ݑ+���2M 0��!�ȓJv���I;�q �ϗ9kx]�ȓ�4hr�"=C��A�Iʑ=͆��N�|�H�j�hD>�����^��ȓ5��{���1(��v�˪d)�ȓ�Pm eƇ���T'$i����y(�13��3\uT�iĤI H��X�ȓp�<E�V�-�0A�MtK6��ȓ�6�A+�T���KW�ü=�~���S�? P�k%H1�輣�+C�B��"OV���U)%�"EhD�Ow�l�'"O����OB�UVE���!�|Q�w"OD%Z��l���&�:k�<tH�"O���0k�����aH ������'���ٟ����	韨�����I,tvɲ�NE�E����'�|�I�`��۟��	柠����	ɟT�ɨ =���V�Î[�`�Ƈ�*N-vd�I֟�	ҟ`��֟���ǟ����X�ɕ#ﴠ�w �4#p��螄p}��ݟ8�	��P���$�I����Iğ���_�
 �t�M!���b�G��]O���I����	���	ϟ�����P��ߟ|��9}B��a7�Q�l$X�����z��$��L���\���8�	����	��I�0P�ea
1� z&�T<}8���ڟ������	럸�����������I�PA�q�ӧa��]+jD,�������	� �����I�������I3�$AQ���-B�m;�W�8 �9���,�	ȟ�I��	П����I(c3�qS��^�B�@��W*�=_'(�����	����������I����I�)u�T)vB<";��fLħ.+RT��ڟ4�Iǟh��䟼���@�I�|�	�w��)�Ɏ6(��1�M�ff���	ן��ş����d�	�h��ϟ���	V���6f��(�,@+12>�	Ο���ן��I����ڟl"ٴ�?9�}D�K�n H� �ON�-�QWT��	y���O,�n%�^L���ܮ*����EK�0�RP�"�%?���i��O�9O����-t<���C$m����EL�d�O�$r�r����$��$�O_�h���4j���RɀF�b0�yB�'��V�O������^�q$V]*B=h_�1A�l�f�s#��4�Ӟ�M�;U�"M����-V0���L* ��P��?љ'-�)��8'y ilZ�<��!�=�e�APht��d��<��'�$A��hO�)�O��Ѣ�АsaZ���v-���0O˓��ji�&�2Ę'������fڶ����"${<�����e}��'��=O,�)9�<���Єum�u�Q��Ar�$�'���,p��,���#��(5�'�F��7gş ��=��L؍cT���]�<�'U��9O�Til�*�~����Y;��q�:O@�l�!x�x�=_��4�F|	�"R.r�����X��-A7O���O��D�>Y~6�(?��O�B�	��|<� ���f���``�[�3}\qI>i(O���O����O��D�O��G� ���[r艎K�~��pį<�0�iG��;�[����S�ߟ�qGJX����Aȓ�c�4�jQ��DLΦ0�4g=�����O��t���<siZ�CZM�d��=8&И�iB����ZX���1BL?�I���R�a1��icr�k�b�=a�d����؟�����@�	՟�SOy"}��	g%�O�a��d5���A��9v>]Y�$�O�yoW�{��	�M�R�i�47��J>�!OE�v���� _
�)C'`�6物9U���̋#���B�<�+H�����VQ8l8!/�6g��1A!�U����Ɵ���֟��Iџ��	s��%�j]#��Z3X��P�Lު6	��y*Oz�����4m>��	��M�M>Y6iAD>*�k�Tx�.�d��'J�6���i��(} �l��<��f�A9��K�5�*�A�^�-����臬rO��D������O���O���6�:����$�A��		�~���OF˓r���PA2���ЖO��� ��P�XsF܀�oD3o޾���O���'~�6�Ҧ� L<�'�Z!'�*?���y��[�1�H�`C�?r��Z%Fݓ�M�R���S�1��D,��ol�J�G}&�Y��1>mV���O��$�O����<�&�i����ƀI04 ��
�U�~(�R�.�&m�'D7m%����$�ަիF(��M~mGte����	��M��i�u���i���O�`b���R�o/?C��4T"���ڻ��-	��|�@�'���'bb�'��'Q哚o�� `�`RV!�9����4���4|9�H:��?�����<����y�R�^d~Y
�Oڔ%�F�:�ʐ8�(7����N<ͧ�r�'%�f b�4�yB.Dh�u������gj�Γ{�����On��K>�,O��d�O��qSa�y��P�����򄬩���O���O��D�<1T�i@�B �'X�'��t1�QN�|1�Ϸu���s��$�^}2�q� �n����]B�)R9�Q�����J�Γ�?IC�
o��Sp�4���
�a��R�F��$m�"x�)֙c3�����N�d�O4��O���2����*�V	XTJ��P�L�*I�vL��?�7�iو���Y�d8�4���y-�K�)�5KJ3Wߪq�ACP/�y��q��LmZ#�M���M��'s����-��'j��<�u�ʁ0M�p�M�-��L>�+O8�$�O��d�O\���O�0	�EȚ'�S�i�I%�h����<���iw~9#A�'T��'���y�C׭���'����yFJ�.n`��?Y�4S8ɧB���br�D<	�c��sօXKE�NP C1AК��A�Q�xQQ��Fk��O|˓˜L��`��U���"fCY�}.��j���?Q��?���|�,O`ql�Y�z=�I4)�x]�w@eY�����4lK�;O|�og�M��	��do�4�Mۢ�s(=f��0��5��y�|L��4�y�B��V�������?mz�8O����he�=� ���^��Ea�M ��8Ѡ:O��d�O����OL�d�O��?��-[+l&�+g�
�\�H���-�Jy��'3&7M A����M�����^�n��$Q���!dW�;�h�~y�'��o$�M���*cI��4�yZw���G��e�H�B�@9l2Y�g!�!Y�x���'�&�|�.O^���O����O���!˦j�n-	�=I�]�Aj�O��d�<�ջi�dh���'��'��>U�|��� Q�i���I���n7��S�ꇱY��P[WCB�u�2X��+�z�~P��H�
em�&ȵ<ͧJ�\��y�ɢk��y��� �Iy�N*�t�	��h��ݟ��)�Qy��Ӭ0��&~�HI�cnG�

�I8CË�a������DF|}�ak�l!@��P�>�J�C����3�A�֦9�ش4k�iߴ�y��'�,�f�Us�,OT	��f � ������5��?Oʓ�?I���?	���?����) ���}�7��շ���m�Y��ij�&�'�2�'��y��l��&4XdрS�8�˄�X'3�mn+�MӴ�x�O���O̬*�it�Č�6�2HXW�T�.����D>>󤃄85ڴy�o�ؒO�ʓ�?	��S���r�.�'E@wc�����?9��?q.OvhnڛFv@�I� �I�	C�5�5��&�%��h��w��I�?�T^���ݴ}���"�>��������'�<�I�"���O(�V(��h��Qͽ<Y�'7���H��?)%,K+Q�$ec�6p`��e�E��?	���?y��?1��i�O&����0o#ȸ�׋M=&�2u\0�$���q���Zyr�d����,=l+A�r�P�1�m�,T=b��ɦ�1ߴ#'����b��=On��Ή�T���O��u؆���]r4�9E��;I\�qs�|rR���	��X��Ο������wg�3��3�T;`�N
$dUyr)i�J��p��O����O��?�R��	�P�Ԑ��%�/?�@�V%���T����4cՉ����O���Z�):>�P���)z0@�&O�(:��Z��E�=xbO�y�Sy��W�.����6f�_�X1�,\�&F��'F��'��O����Mˠ���?��!����Ʃݩ"�����?Ɂ�i��O:��'�¾i�26�$(�ҭI4V�5�l�#�ݣg-��Qw�x�4�	ٟ{d�JZ�dh�~yB�O��
�0�,`��K�\6l`A3E�%�y2�'�2�'L��'���iJ�Y�m Sa��B�N��V@s&����O��䦩�t��Ty�"d��O"];Q�צ�c*R�+�|�XbRu�I<�M�ǳi�����s|��<O���ҵ^��4�6I	�|`�h"*��q"����?�&��<����?y���?Af�^B��A�DW$N:vD�����?�����dXЦuh��쟼�I�`��?���	�=�u"� �I
�!�a"'?��X���ٴ`q�F�%�4��I�;U�A��c��s�n(0��88��G%=
�HCǪ�<��''���+��L:T�2@N��F�F���u��T��?���?��Ş��DĦe0�R�Jo�lV�.+���V�I�,��'��6m7��-��$��is�"��Nh!��)�5h��r�թ�MK�iV�x�e�i��D�O�|D������<1��D�e��3��O�s�꼓4��<y.O����O��d�O��D�O@˧.�TS�*!_���%l�1tHdx��i:p )��'���'W��yr�o���]��CW�S�+F���#{N|m��M�t�x�Ou���O��}�Ѽid�Ĉ=�1�nC"bTڸ`W�~,�d3�(��t%�O
ʓ�?I�WE2�����t���"W�QފI@��?����?),O��oZ$kBܗ'��!��u��u$�$y�u�6J^��O�'��i{�O�apR�˦UHe��@Ct�S=O�$Q�bT99�'�:�@˓����O��Z��%�A�>��L���1u�� '�������㟀�Iş�G�T�'�<��n#
m�ݛ���,!�I��'��6�DS��˓` ���4�P����ݰo� �d�Tk@���8O�o��Ms4�i��ƹi6��O@�`Ҍ���Ŗ2	�m�$N�)�Ht�"�)@���O@��?���?����?a���X�a���^.��	�OibT�)O��m��i�u��͟���A�s�x�1ߧN݈HTO�E0�Ǘ����̦AIݴ	������O;��#[L����+A6(-��٣�Z|F���Y:�� *j�e�'p��&���'`yP��Z�X����@�U��`S��'V�'������W�`r�4a��,Q��s@0�j�.�'2�b,�j������'��'��k����~��	mZR��0���9!�v4��厏]�b�sG)�Φ�͓�?�+�!���釅���䟸��N�R
,J���H�}�7���e'��O����O�i\��'��hy���zv$ȕ�^�.���"�O��d�OB�n��6@��'�6�4�Ď0*^V��u&�Ȳ��$��'��شZ�6�O1Vp*�iO��O�3䥁=�v�hՍP�nn�%�(J,ܣ�'��'�	�t����	<�֝���&m��T��b��p�I����'d\6m�&�E�'���'1�S�?.0ɘ��>n�f �� A�mX�o��I��M�ѷi0�O�	���y�@''�:Ǉ�\��A�5�3٢@i�- t����C��O�UhL>�0j��i^��i��_(Ҧ@������?9��?y��?�|�+O�$nZ)}T�):�/��lahZ�/��9Úcyboe�h�H�Or�nZp��@�ah��c��P�[�����4E6�&O&�v;O��Ē*s�8�Oq�)� ����%�4ֈ%�0��?��\��;OJ˓�?q���?����?)���?iMI�|�:�Vj6��2խ��Fl�E/9a���.O�ܦc>�`�4�?a1.^'Mv�C�@��i28`�"[6⛦c�<$���?M�S`�d-l�<�d�<o���B�.̽	}�����<�V
�/J����H
�����Ov���/��E2�K��Vyps!�.$���D�O��$�O��H��&HҨl���'����o�Ayw�BiE( Շ�^[�O���'S7�Ŧ�H<i���0��e�H�%JЋ6K��<���W���0pa'u��M;(OR�ӄ�?�7��O�I�3��/�Ҹ��b� #�Ƅ"�N�O����O����O��}
��w^p���P f����E�5o`��!ۛ���	W���2�M[��w��0Ư�>�9#ժP%Xp �'\�7M��:�4v�I��4��$�!������jp���/��Րg��
+��"��/�$�<���?���?��?�b�\�lp�pB��,9��Ӗ��$Iæ1��BIџ�I�L�SG��'����?x�F�*� ��0yk���>�%�i+�7��f�i>����?ɪ�A^<����5���Ť{�R���LayR�ߪ�����2��'���$F����D��Q���Ba퇗1z��	ٟ�����i>=�'�6-�#�"�$ݓm�
E1���̚����e�?AfX���	���cڴD�&�#&�˥5i�h���X�v�1�۠�M�'6t4+U�%d�8�'L܆K%�O�4ט� F��tO�VPI���r�f�	ϟ��IɟD�I�����s����AQmR s��� ��C��)���?Q�Z4�v��e3剰�M�M>�".L�l���+5�qk� "M��)��'b�6����ӭM��oZD~REܾ
������V�s
��[>�I�����!P�|�^��	⟰�	�x�U�H�fji�0cK�u�"x;!�Zڟ��Izy¨a�ҡ�b��O����O�˧4�Ҽ�2�-<.��#�X� `��'l����{Ӵ%����?��HI"F��ru`�$	a�Y룪ѭq���U�=W�e�'�������&�|R�
�J^����%*�Բf�@+M�'���'����_��۴m�5�R� ��aL6��q��?1��k���d�F}��hӬ�1��7�	��e	�&�<X�L���޴D���ش�yb�'뺽*����?	�EU�4kv��4~��X���YV��``|�@�'��'���'B�'哈U��KRcX�x���	2ǈ� A��Yش}����?����䧽?Ѵ��yg�K�q�n�C'�G�:G0=�Q��,;�6mKͦ�I<ͧ����)&A�۴�y��G;=vȘÅD�71Ѽ4Y���-�y�̛\j<P��� �'k�Iȟ�	�W�)�b*��y�� �Z"�%��՟�IןĔ'R6���zV����O �d��XA�p@�Zj�"ǀj�lوr�<����Ms��x!�a�Z���m � �!P�@� �y��'�H
۩Mi��*�<����F�	ğ4)���B� �H�aĩx��D�&ߟT�Iğx�	���E���'��PRW�Ʋ�А0� ;2�	+��'�<6�\�_b˓hh�v�4��x�h�g�������"����O�7�E˦I�ߴ�^M��4�y��'��i����?�
d�9BZ4Q�#H�|@H����΄G=�'B�	ϟP��ßP�	۟���1vQ�i�aD	+t#�`5��-��ԗ'��7�4f���O��d5���O|�����a��".�q �$ �G�\}�n�b�l����|*����EL�S��l��+��P�
� ݂,{��wO������0
�����6���O�ʓ^���a�� 
w�E �.��7޵)��?!��?���|�+O\o�U����ɾ�^�ᑍu��e�7e֫D����	�M{��>�g�i7m�ɦ�@��]y��re�`w"� G+Է�,�l�<y��:�z���h����/O������=y��A?W'^(8�c��&���Jt>O���O���O����O>�?��G �'`��	Ck����A�bJ�Οx��ß��4~���)OL�ml��� ��V&�Aī��c��P(I>Q�4ś�OXYt�ih���O �0T�˥,�3r�ؑqK<�0U�ņi�L���$��O���?����?���xt<���x'`�Dʳh�4	���?).O�mZ7Lfl���<��B��8��p5��7f�@٥�����{}��~���l�5���|"��H����s��,	�8�*҄ũ}cE��	!�l�bjR������F���N���O��4�؏}EΩ*L��9����e��O���O���O1��˓,��&�I��r-X����St�s�d��_�%���'҅pӎ��q�O�AoZ<��Y��"��Z��P���W�&�,�A�4_��V�M��'1")V(xab���1^��I�=N��Ӻ%`���3�6�IHy��'r�'7��'�RU>��+s5R�h�%M"Mb����M#��¢�?Y��?�K~Γ[&��w�N��f��]�궧 
=	�@Ӄ�d��1l�����|2�'�ZD䕗�M��'��%A��֚5�,9�j<Q��ؚ'Kl�Z��S?�H>�(O2�d�O���)A�}����G*֕d���'��O"�d�OR�ľ<r�i�t�*��'���'�N�C�"%_~�;d�כZ�*ͫ��D�g}�HzӼ!n%�ēQh�H!�ȅO��0��'�;e���͓�?��_��fa
Ԉ��������iD�D�4@Z�ЀJY�
qx'�֜n����O����O^�d*ڧ�?�Ō;l������N��I��o��?IT�i��I�Y�d��4���y�CG�d���ӧG.H�X5H����yB��Ox6��립��k�ܦy͓�?Y��R�:]��	�M�? ��B�5%�.�@A��P	�y�F�9���<i���?1��?Q���?a�ē(X=���~�:@��X���D�Ħq��$Jhy��'K��e�W��C��]��%�536PT���tyb�'֛��:��O��$�OkҰB��[FH`���V�= ̳Mþq(gU�H�V������*��)-�uГ�IX�P�;��O�=��O\�9m��8$�H�s��ܢ�1D�lx�� $0]Ft�##گ�D����;�	�y��l�	�Lj�����G0W'T�8�j�1��`��K
�nk����e
C 8�di�	���H�'Z�E�RW�٧��3�P�5�U�;1v�A���w�&�ѳ� Ԃ-�@̇-,*H���'�\�a����T�"b�!%]���\�.���c���L��1�Q<�Rxl��Z��r��^��ڱ �!خ�Y�O����O��O����OUʴ��ON9	Bk�2F�m��Eьc5�A�q}��'��'.�*+���I|�CΆ^��̨�CL1|/������iכ��'��'���'����'�� �*9���W��hg@H�m�x�IAy2�OC}���d�
9��HJ��EҲ@́[�&E��Xt��؟H��>�`A�	`�Ip���ǌ�� b���v�l)D�զ��'�T�J�!i�\��?��'sJ�i�%�v��?h���c@N�k�Ҹ#A�r�,���OlI���O��$�O��?��T���:Q���&JМ��DL�~�D6-�&F�nZڟ�	�Ӗ����<I�'��N@*���? :�=����>R
�f(N0xW�'}��'��Oq"�'��F�\33���p��	
E%�=JRE ���	П4�ɸ ��ۯO�ʓ�?I�'�
]p�R>'¤��A�En�3�4�?����?�cBX�~��������۟H��I��	��F64���JR*�dK"o��*%�Ҧ�ē�?�����{�EEX������0Cv�@0�Uo}��Ѓo�[���	��t%?�0��A6�ZE���f�Y-�(Qj���}"�'0�'x2�'*f��%Ҁ=4��j�F��c�]JB]���I���Iuy��˽:>��U�~��ӎљ
Ш���LOK����?�����?���k��K��W?��Hbf��ԃ�㎎ah�u�gR���������~y��Bzx��?Ab&�'e�`�F� 0b��p�S�,���'�	ş`�'�f"�P>]�I�ϸ��s L>,P, � D�'����4�?a���?	���t��W?�	؟\��;>�$`R�jL�C����GI_/t.�9�O���<�@-���	�Ol���?!0F�V�WnR٨1@�CTx@�сs�J���OX�`��Ϧ��'lr�Ox��k$Ǳp�<��"ͭk\-x�#U���Iß`Q5K��I˟t�	Z�cr�C���e*L!i�-\+:�)�4s��Z��i`B�'f�OÖO�)�A��)"�ֺ~�V)�����mڥ)gzh��������h�m��W>���Nj�pił�%{J����ż�M��?�3�ཐ/O��I���# b��``�� =4���#��L�O�������./jQ�J�&I<���+�M�l�H���Gy��~��B�?���Xŀ��aQ�@5w�7��On@����ܟ��'v�C�P~D�!^�C��e� 6F��m�W�D�	����?)��?1��[(Z�$��G��l҄�V)g�4�ۈ�')��h����s"�_6S<�䒧�ϡ�6�������ڟ��?Y��?A���]}򊕘h�>��PbY�>@@%{�Oŧ�ē�?�/O��ŧ4��ʧ�?y�U��p	V�״ k�x���"2��F���O���ւ*� �O� s'��K|��*q,qi�#��I㟀�'` �bc(���O���Ƽ�#Lx�8ę��N�k�=`��x"Y�� #�ӟl'?=�'d�LJ�J�&`भ�7�$ �bL�'#"�U/y�R�'y��'��Z���07�n�S��N;�(x��P�<�`7��O���G�\��b?ɐw�1,�!0�=)8�ȉ'IxӚq3�P���IΟX�I�?��N<�'J݂���_�W't�SCڭN\4����i8H�'P��'R�O��s������+d�̴��h�
_����rΟ�&z0��'�ʼ�2y`0���b� _�ݙ��Fv"
���3W�lx)D������6e5'I�uJ��T�@����vo��2��9K���ŉ���м��g�)�OO/'L�+�䝱?)�l�숎,A��Q2C��Te��[�a���hS�_3<h�皿+� ��.�7������,�5y�#�y0�	�"�0��	ޟD�	ڟ`���ɟ��I�|��dЍ?Sp$���� p��#��\�d�ް��ݟ��%�Q�\�Bp��DV�N�X�f�JQm�����PXt1c��~\��bG@8n����Ǔ<�u�	��M�G�4<�M�0��<V���DbҼby���dZ^��yB�(���n�y_��"�y�b٪@"t2fa�<6��f��y��>9+O6HC�d���M�Iߟ��O�
p�CD�:e�MkƇܥps��▊B�2��'2��_�� �[C�24`�kT�K�$��O�jY��܁t�vi��� �lo�4Î�D�]���Yb
=�6c��;iT�'!NB���)X6ɂš�	@�HGy�a���?���䧡?9b�rV8�y��KL���r����?����9O0��6k@$^АYsV-<(S$`�'�O~]�)�|T��*�?q4�#�<ON�[�Mզ	�I��<�O�X5�'���'��d�Ȇ�d>�٥,�"����H�=�l H��{�^�ԧ��'��O� ����ԭ$ܜ�3�L3E>܃&K[)���:�/�&#��J�O?�H�$R *�q�x��5�	����i"��OZb�"~�	*hu�l�g��}<��,&C�5J��H�����1.}����v�2"<�$�)*G!OV=�+*�����K�<ivG�Q�|DK�G"J�����`�<1�HXc�ԑr2큞8����Y_�<��fW���������kB*��\�<���ڂ4�!�D�iB����D�W�<qfd9qH��R�P��=�F!�L�<��:�P�Gg��S���`��G�<a�G�J� XA@�^�^A����G�<�V$�8iF8u���GCT�`#$�]h�<�GOO?��< �J
�\V +��a�<1��ۀX� @:�.۴e������`�<�6�ҟLt�k#�
e��X`�r�<)DLK0[Q�=�qB�{�RdrQ��j�<�^XS �D-fuz����>u�h�ȓa���z�Ʈ+���	��&\lΡ��u^�d�S�ͧ>6� �Ӌ��~p��0_��*�Eǲe��p��]�5����%��F�3F,^�]¹�ȓ(��cE��,)����1�B':��ȓ'�
)Y�%ٯnL��PB�~$�ȓ�U`�.��<����8�"O�q�F/�X��)P�T�����"O,��Ӄ��F��I�&Ne��9��"O��â˘,<��waA�i����"O���"ۍ	��̉A'�XJ��h�"O �,E���i`�"5y(�i���y�aJ& �� ��`�3% �Cdc��y��W��ճ�>~��E��y�"ݏj2J��0ꋦfFN%�b���yr�'Z3ZQ�gƣfK�@rE �yr��3{�(�JT
�Z�����y��ɑ{�H�{��E�Q�=��ԙ�yg�0H��Òk6D�$��3a���yR�)H�HsS�^�5����w�ؓ�yBf��v<��V#L�`�lI��O�yRN�AK8�����Q=bܺ7mT��yBgR
$p�XQ�fF�P&��ö����y�eŖ�R��s`X-=�0Yj&�R�yi�J��4�P$Ω+'��K! �yb�&���(Z���Ӂ����y����mx�t�%�PC���F]��yH�8�84�-��ҽ��c��y�
�zx+�.�-?F��#f�y"jK8�x���	�2�y�֎�y���w\p�E-ājy
�Z�L� �y@^�6x���"�4��������y��ԑp���Q��%e�@�J�y2�W����-�T�\�3�kD:�yR�A�\}B��3M-�ݙ���y�e��	�g�I�H"���Pl���y��0V��)Qh��>ּ �"��yr���$N=A5ِ0Z:��r�K!�yB"�75P�ȴ��!�@4�2`�7�ybW�W3�u��n�R��R/��'F(SR�2S8ҽD��-�Lx�z���3*�����y�n�)��"� ������k5yl����B��	�]T�"|�'���"o�?�rq��A�  Te��'Ѹ���� �)�ȟ�����Q���uP�1�{��0�>�!���B�AYvIP��p=񷌀�Ж\P.F؟D����Ĉz%.�9-�����.(D�� \�0���<����@�F2
b�S���VD�b�Q��E)i.�}��l���(!$&����d��	XC�<�3��0h�F�"dI�Ϯi��g��~s��rc��򄞾%
>�snm"e�ܙYv�͛�`�Ʈ,�ȓ,Df����ވG��)@'� ���Bl�<L;�z��"��='I '2a�DÞ[I��FG�gX��9օ�`�)+>�� �C���&l�A�N&�y"�]00��ގf��<+�ֺ�HO�\ ����h�V�SR��C���3��B6ȣ�"O����y�~��K]�q��ȁP�iS"��%'�o�S��M����Tas"X�i^�qS��h�<�c&�!WlQ���ܼFx�D��Pv��}���i��Q���V`OR]QC�
��z��R� lOh\C�hI��J'�АRi���/С	A�(�B�Ԧ[%�Y)I��S
�.�$d+j��_�f�hDO)�~T�>QEB�_պ]���P�5�~�����'�j��	:S�t�� ���M�x��	�'�L���t�vT�0�x�\%Kp��$X<BsfW�N���	bӼ`@��Y�)I����^>�$���"�;&R�{Q��[؟8y�CO�P���+e�G�"`��Ytd���1�4P���	R ��Q�k� qf0 S�F�@��!ӷ�8��է'{�Y�S͹��0���QmQ�|x�o��y5Н�����A��ю�O^؈���{��8`��Kݺ�`앭��'�.��)7�J���<i��P�vi""N
j�0�NSW?i��X3Q�9RT#�95��Rs�H?��̙�:�L��ҩ��S���K��!�� �n��>}�Pڒ�&4���&,G:)..�!��b�~�#�DE�(Br����z?A��jZE�/�$wWP���A��s�:���"P�ADj���o_�_�����'=�m cL
(M",H�(�<V8�D:A-�8#L�@q� ʒD��b�gE�3TB�1�$G�"-J� ���E8M>����=h/�R�e�u�S�_v�'�݁���e�*IRb`@7|��d��0�Z�� �X9P^$���M�%�$7�E8kR
� �Iʋ=�XQϓ"���+D��.8���G�2��'�z��q�ɷ�Z�+��H�/��|�O>��צT�'
}f���wdT�1�N�)Uʠ�C�:�JB�ɎN�<L3b� ݢ�{��"q���`��cV�	��%�[?�1b_�&��t�)����g͌f�����:#`drc�x�<Q�I�D��E��;�޹��dE�!K�lٲH����72�I��D��[�)��p�Ç�	���1QF�_v쑆�	t�ʩ��Þ���f�Y�8��_2;w���*A�;6����+)4��S�ăC� U�X�p�O� )�	�{�Rizq�4�']��
���_�f!j�l���q�Z�!P M�j��2 ��l�MlZ+{�
�+R��s�h5*��֒g̾|�e�n#6�I`"O���)Ki�=���&����^�H�T�ɸ05�{B�P�"IV�R�z���K��G�>��(��v\��$F�D?PcW��@�CF@֚a9!�Jr=�=;�]}0)�Ta^:*ב�P�R-�^K�>�t@
9D<�ȅ�T�[�9�);D���sI*P�2�ҤӦi�j�r`�e�.hA�E��������چaD��suo�*-\x-��cV;�y�kM9^L���hrI��Ί���d�x�D��-+B!��F]�V�`	1���Y��u��I9G2n���'$n���@�2�0�aX/.'Θ�'
A�2dA�=y\��#-��r���2��䅩L y��	$?EjH(3�3I��PN�rg!� n2ܱ`�N��ꐓ_���]�{�LX�=E�ܴh�&�ց׌#s|`�%N՝*?�����كN�x_|���ޱ*��(�'<�|���'����׫wO�m�1D�c�����'L2ء��o�l���)��S�'Y�!ÑdP<�$����wm��y��Ip�%;�Q█b`��!�yҮ7�D���J9L� q;��,�y�\LLEZ���K*�pL�/�y�ĈA��rԩ��N@���f)�y�˶Jtd ��M;I��10#0�yR�H&B�&�)��>�^�4�y�]<�
��a��f9`���޳�y
� �(yta�Ml���L#l�m��"O@�ѲaB7AR��BCI]�¡�"O���7Μ7����+խ�t�2V"O�y�.�A3` ۖL���݋s"O,�����	(q�ņ�Ȍ9"OH}z�A����h+�� |�8��"O��`ή1���Y�d�Z� tP�"O�\۳��e̼P��@ج��A��"O��g!��9�RAW��� ��1�"O�����"bBh	�-�
u��a��"Of����� �/a�Nm�"O@d�ꚝm�H0ӥ䋸%z\h��"OVH	T��.'w���D �JF6�Q"ORܢQU�H� �H8���"Oh@��ү~�*%&�-!R���"O��W̋�,o6�Y�,��	d"Ol(�/��Z�tIժL�H�=��"O�ݓ�䔡O+\�D�� �$��y� �����[�6>.8(�KG�yR03��$*����'��[�	ޡ�y⢜�s�`*-���n�0Č,�y���xEK���J̘Ӧ���y"'��w�T���)�$����<�yr��*K�\�H�2i)"o�:�y�ʭN�*���<R)�L]&�y���m�R���>�P��h��y����_> �Y�V
�(чل�y��CKl$I4!�~���4�y<a�y�&�&8�9����y���'���QK(`����U��y"�޵��m����/h^�tٶh[��y�-�|�6�KW늓*�p��P&���yb���Q� ��-��R���'�y䆹-B�yӐ�M .r�(d԰�yG_+6����G��~9 
$�C��y���:c��NH>he���y�f��#�Ip�m�,����y�B��VMīW�C�f�aÀ���yR�$ֈ� K��;ʞD�RB�9�y�n	�ʬr���!=*�#�(_��y"�L�\�`�A�$�fU�D���y��
7(���BQ+{�zQ��:�y�H��[]����]��Xk�=�y�ǀ� ���P'[?$��� q�Q�y�C@+	�5��K-kMZ5�͟%�y2!����)��K�K~������y�&�JV���B]���q����yZP� �D��t!"T)���"C�Ɂb9��xS	G��ݣ�v�$C��64����Λm����s�f��C�I�R�rm{pN�W&��ifi�	<"C�	� �P@�g�D+1`ŋ4�{UC䉦P��С���DYn�?V;�C�	�x��I	6�� TI�u�P�~èC�	#Z��a�M�H7��� ǟ:z��C�f�E:�+�L�!I�_QC�C�	�r �L�`�X<�,(�C��7:82���@�.�F����6zC�I=X�hF@�*h��6�V�j{2C䉍`d怣PjJ�)����G�7^C�I�t�� b©F#�i%F�O��C�I���c��.����DY+ǂC䉋]
�bD�Ǧ[�~Io�3Sw���ȓdl]��&�<&�yg��6f�H��S�? �C�mH�B��{��q"OI��`T�2��Lp�"O�a�'�� �r�ل@�T�V�S$"O�����B��
E^� �"O��ឥ_A`a���P��<��"O�Q"_�M�!����:�&��"Oҩ	g��J�05�P/��h�"O�TU�ا$H�:���l�ĵ��"O�����о3��ſw�\D�"O8Ա�hK5�
�&��L����"O>:w�J�sXr�EɧcX-�"O���eoL�:Pes��Te�C�"O~X����!l�촩f��;F��g"Ot�+�N
�HRm ����Y80Xҗ"O�!�"�O*���sr�R,Na��"OݓTK�BT����˜ �A3�"O>��QKP;<4,��ᒖ�X�"Oh���ÒH/ ��P ��v<ͺ�"O΅X�A�s/.��#NJ�2H���"O�����a<r�,W�5��c"OH��䎣|�(�;�I��0Jh�"O2�j�,_<A�z00�G	cW��p"OH��e�9]ʄ��V��[4R ;�"O�(Ś�eV4�(�Ћ#�Ft��"O�t���*0VY��蕤ɘ �b"O(����҇nl>����X�b�T��"O��(û)|.\	�,��	�j0��"O��A�腰L{�D)UkQ�`�c�"Ol��*�3
��`�	E�T`��"O��SGB�ma��S�G%�U%"O`�X���KP@�����/0x��G"O���p�J�@��FB�]v�"O����dޥ7��ᅌW�ez
�@"OR�el��d`�X�ą(uU�t"O�逕杵t�Nl�"�6qY�s�"Ov��p��r�vpd.ƄlV�] �"Of5�O���}��.�9��"O�{���~�Tl�����q�"O��Wj�/4u8�B��b�K7"O����Ȫ��y�S�g����'"OI��U�n6&� �=u����s"O�)1�ω'A��I���^�0ؓ�"O��Y�d��]{��rn�	�`i�"OVt*�ˋ*�P�mW�Q
�� �"O�s񣃒b/�Ål��Sb�q�"O�����n���Q�LlAn�V"O E�udԞ~2ȀG�w"$D`�"O�����<q�xcDmXsx(�"O�01���6���d��lb�Cw"O�(�#�"e T�`oY7EX��r�"O^����ҖBRHre�I.�0h��"OL���8����E��tk^iKu"O&��Ƈp�m҃�
����"OЁ�p<]l�ԓG��f��9�"O�J� ԟ4��[A�"~ŔXA�"OV�Ar��=;�U��1W
�͋U"O�x�����r̆!���;Ljd��"O��e�	<���AAŸP��E��"O��ۺG���q���6�B�8d"O�$r@�ѻ^��`��Fz�
#"O$�"ed�-~��bD���d~��"OΈC��\ jnh�C'ׁ;��u��"O��V��(i:-��ƀ�|%���`"O��c��O/c��r��;j��Bw"O� *�j�E)��xDS**�ٓ"O�\k��30+�Z��W��h��"Ob ����
ir��Y�6���"O�P��g�*^<�D�=P�p� R"ON�і�߱LAZ�ȕ:\s��y�"O8}EK�U�M(Gk��"O>��6㝸'.�V��HS�H�"Oꀀ�kUM�ipb�rƝC""OX4��r���i�b�(NS�� 	�'�p�� �ʦJ�$Ո���:W[Ą)�'���[�ˎ���1�B�NU�Ir�'p,����_�hse�M�K��@*�'������Q\ ���сm�����'V�i�#�w/��0�L%̴���'bd�aĝ�c�R����Ŏ �U�
�'_�4Yf�o ޥ����.%�e��'���nT�*f`( �� sJ��;�'�aᦩ�� fm���d�✈�'Vt����);�j�H�%����'M�U��a�'.���&iS��4)��'E�H�GHh�q��J���6Eh�'�@s5�ҿ%� ��&N�uZ����'���$�	BJ5Q�h�'�l��'�1c��;�i�V��Cn�ӓ��'��(7C�0:�jٸe�6\!Y
�'�.9�F�,Np���&���P�'�h$�a$CFl�l�7J]�u��(��'���	���$>�B$��,>����	�'������`���N_�NXy�	�'w쐰S�BBԀ��o�.����O�왕��`�$_'uFn���"O��qR́1=.�84dY�\��z�"O��K%5Dv<�EH���� R"O �B���?<ÄHH���v3�=�4"O����$ޮ
�	���Iq24�#�"O�T���S;?��E[ŀM/w0�l�d"O��h�� ������4J�J�"O����<F��ER���]f��"O��u)�%!vq)��F����!"OJ 4HܕC��@(4/H/I�@%��"O8h�6�׉0�(�0�N��y���� "O���΄�N�{f$��B�XX�b"Oި` �u3<pCp�F
�0�a#"O.X�U��(͈�`?
h2���>A
�CPbE��f���e�F��A�r݆ȓ07r�A�)�]���Y�*�	�"\�ȓ'�����	p�)�MJW�V|�ȓ=��uaU��t�#��9��1��;k��GE��H�\���x^Ty��b��Rf��(��u�k`~���7@�,Sd[7������?t��(��P;!a �ǚU�.yDÔ�BF�� ������)���ĉ�t��WRv@gŃ��d{BeQ�'�-�ȓb�KE@���֪q_���y�@�NΈ�!���S�`h���Í�y��ʠ<�
�p�J�A�4����y�F�:/�^\h�ئ©@K/�y��Z�{����@j�|l���yb' N�E��{Ҕ����:�PyR�	&S���R�dn�pƧ\A�<I����!0��?g���XƊt�<�P�L01E��xR��V�����Hr�<i���+��r�KQ�{Zn�"�h�m�<� Zu��� m|�5�ԃ$3��\(�"O��G�� ��]���4^��=��"OM��*K<
x��aU�S�Tq�s"O��C�.(�V�Q�+�����"O���E�z��x!`Ȉ1�t��"OH`
��us��3��tm�� 5"Oqj%Jڛt�l�)�*R�{:�䣧"O�]yw'�":!�\d��/.Yb}�"O�2�->dz�i�4b�l�"OHY7 }�Rm`i�"�����"O�0RG\�Y Z͐�CBJ�m��"O��؅V�yr �r�8;+ᚒ"O<��`]M��` ݫ%^� "O��s6AS ���r��	:�1"O1�E(ѐ�2��$d4��s�"O*��3(ڒ^�B�x��q��_��y¥���L����i|�P�͉�y2
 f�%� ��X�$s�� �yD��(�
pxą
:�X��Y��yR	��*��p
�c[�	�<���yR�)8��1T���+�0%Z�,E�y�(S.ϤdP�'O<veH����]�yb���B ��8�ɀ+qh�� ����yR&U�a�p,˷�͸Ln\/�y�.֎K��b�h1Nؠ#tmԳ�y�."�u��'T�!E�a��5�y�B �QE0��Ą1!��@�;�yBkL<"Җy��F�rT��G���y��Z']���2)����#���y���)���󀀿�D�(�n֝�y�E�J��i�������Y�y� б��(�uC�$�Duy��	��yr���D-a��єLz�ݲ�#(�y�JɎH^,\X!��<��<+����y�EN�3��/Q�-:������4�y��1����dF�3$�}1�<�y�(�]�0�j͡`Z�H35�I �y��)K��U��,Yb�b���y���b�˴��O"�ġ���1�y�	�3C����Ą�J�%�R�Ȱ�y�+�A�<�����::��)ǀ�
�y��̝i�̜�&U�H�����\��y���B��QR���o�؉X E���ybŉ'�
���� 'dĺP����yr��6¼�뇁עW�V(H�a��y"C7By���q��6Y��uK��Ņ�y�S�7�V`Y��A�LISw@I?�y���@1��ȁ�69�	P�HT2�y����Ґ{�eL�vE�?�y"K�_��Y�CK���rqp ����y��S;�~�Pte��w���2�-�
�y��YO���k��R�D� ��&O��yr��{߈  �nR2;?��)����y�Vj��Y�k�3����mĤ�yr`]�a�4��< t 2��y��E�$$�w`�&���I�yҥ	.\�����z�tT���yi�@�S!L��'uܝ��F��yREس�p:JV����I���y2B�m����'�4���$���yr��0/ �{O�j-�8#��9�y" �!n�Q�I�*hT��!��R�y��|����,�M��DjX��y��f
�۳�O�O|�وt� >�y
� ���3'���i�&Zt�$ v"O�m;E`�0g���P�=:��("�"O4�*��d�^���ăRS
�E"OD<�.��8��a�Lt0��T�<AЎD(~.Ź�3@ ��
�Q�<qdnթ�!z0H
/W!������V�<qR�;P����l�g�<A4(G6n�|c�Gӓ�j�u��l�<q%hș��-��ܦ��EQ�Qs�<a�K�Eh��Z�&��k"����W�<����Q�a��D
Q�1d��J�<��c7ms:�K$�("�,1B�JE�<1�"J9*q��j�#(&B�H�l�G�<���6D�48�vjRIܒ���#NF�<a�N��Lsd�H���:h`pQ+��<iE�b���a�lN��K�b�f�<��n��D~Z�(��ŵR�"��A�a�<��-q7&a�DW�d����g�w�<���U�j��B�6�4��F�h�<aT,�W���q�E��5����y�<y��Vn|JE@$iȹj�V����x�<a�-Q?=��k�B�?�,)�d�w�<����(؆���*X<1%N\��l�<I��FTn�XzdJ�8�l�p�@@�<I��Z�JlXI^�b�p�}�<���K/B
�yF�M�,^�u�uÝO�<A�ɛ�LXūQAlJv}�7JXJ�<Y�#j��RPpC��A��G�<ARaD�lQV�!aT�M&�t"�`HE�<�b蓘o\D�+��T��"�&�C�<��[=gˈ�儒35>�f�x�<Y���>*�q�c�':�{�ii�<�tǖ�{(�h;���A���ӭ b�<�6 
 T��@������@m�a�<�4�ɱX����2DԐzf/a�<�.���i���ܞ:d��PG�[�<�᥈>�V�Dg�0���7/�\�<Ia��=;�����\T	��0�(�|�<��֥^)�R��$�؀��Oy�<y#�^*z���d��D88PT��u�<Yuf�8 "l i����$0x��G�<9���n��A�J�8`���^�<�r���=<6�@�B�6d�	�mFW�<Y��-7����˻`�ʉ��]O�<!�� 0Q�U��M�8;f��b��L�<)&$�=�z�ۇ�*u2^4c`#LF�<i�B�q����-K��D äh�D�<i����7g�x�%,׉_����G@�<���۶/Ct��B́�ZQ�Q�7�GW�<	�L*k��m�F/�e��)P�T�<��ӎ�v�aq���Ƭq �v�<!��N�=�����79Φl�.J�<Y�)1����[�y��!QWH�<Q�LG�pM�q�(D�N�_�<��C��J�L�9cNˢ)<����r�<RMF�w������Z�Z��W��r�<�pkE����Lː�BDڥ�Z�<Y6� �<_�����=J�u ��YT�<A�,�� ��P��@Z!"�����eR{�<�!!�`�D��S!�r�<l�d��y�<�ҍ�_r�6��z�ިAF�a�<��l�u�ș�-ōM�E��O�h�<��쐾o=�4� H���S	�M�<�d�6*��H1셅�,�̈́`�<� 0L���ЗZ5��C@C8$�h��"Ou��D��T� ����4��Æ�^�<၌�J�nq`UG�>����_�<A���Ŵ�b �Đ<�*(e�W�<���	z�Yr�-�5h1��h�V�<q再/0P5�G�	X�4q�3��g�<���AϤ����Y��т�f�c�<�q-@�J9{Po��7�����k�<�4/�<CJ�A�a[�n�X���&�g�<����w�nI�CO�IL�*W,	L�<�$KB,H@�D�]4'U��Ba�<Ƀ��97jʰ`%ШTl�B,_H�<�����d��x��$��1��Yy�<)wh)0z�4����	B!ڴ	�)�o�<!r�[c�mR�K�;�ai�"�S�<�2(S%L�KӮ2��w��V�<V�ͫq �)@�N�d�����CH�<ye$Rx�Uk��
8 Z�Hd*Y�<A
oa�/��q����T�A�$q���{ȴ�I�$ˎ���KV�X�n�.M��iֵ𐄐�GJ��7��5U���ȓS;M���I�lTL;��� �:���-�T�PR!;n?����l,K<�,�ȓ\��=IR�^$sF��Wj��LVL�� ��(R戠��q"Š5�q��J\�ej2-�:d��OɁ	�ԇȓjr�(r�%�=�Z򇋇{�H�ȓD��l	�B�0>�ة��L���NL����u�Ѕ�G�, <�������q�R'4� 1	ƫU+0t�-��"�8 ��)9 �u�!��Eb�'>�@��F�S�H��Q@I^|���
�'���Jʝ~�
 a��?hFp`�'P�E�1%�7.F�[�œ9�E�'D6��ec�?\
����K�)�����'!.!j��]'M��Mۧ5
Vp�
�'�(��ѫ� 3�> a4��=6``a
�'��;���}(���ˌDy�ٸ	�'fn�	�&�y"8�JQ+�>�ʘ�	�'3��"��4d\H����ȓP%�-JBER�E���rGE@����]�R�b�"K"�\س�ļM�,܆ȓ"q���Ð(8�u�V��!1�e�ȓ{��u�����T����H氅�}�����żrt��B7>������d�Έ�j�i��]'Fn�ȓd����KN�����iZ�]sH��+��B�,b�@���8���ȓL�@��#!�b0���7h<���\y���A4�����2g@HI��#]��#ϗ.�8��A�(bx���}�����!�9;�%��F��m�H	�ȓ/�ZlRT�ѲZz���C�?���ȓSV`�q�%B�aԈ��EJN�%j��Fh��O���'�P,<��]�ȓ�ؔK��4�D�ӕ�̦|Z�Ԅ��j)�a���	��i�"���h|M���Ԓ!W~A�1��Z�@`�ȓ�(�Yb����T��ȷ_�t`�����cG*G])�C޻E�@8�ȓR(pP]y��(cQT�2ئ$��"O �Ic�I�e�Mh�!�!M�ʹ�f"Oذ�6W�����֋3{�d��\�<A�KJ�3�hi@(�]���J���B�<� n�#e�J#:�^ �i�w��5q�"O��I�`.���w����䐓"O1�m\�cޢ�1'_1d��dQ%"O�Lk�'�59:45jwK@m�"O2����r$���f�� f�h`�"O�9)rN�c�(�:p� {ʥ��"O�a�!�4��šp%�"+`���"Ob��C��Xa���s�7�b���'�(��!�5�Xa`0%T+�J���'��e���#�x�K�Qh���'��+�`�i��2ք��'�|��ubZvA�tX��A!��\��'�`["��xt��D	�ܚ��'f,�ch�7@m�V�(�bT��+��= ��G'H�mA4�	�ȓz�����-ѷ9\2���&����|��@a��>-Tj��w(���i���CX1�Z@��o��@���ȓB="M�s�'&$��`&$�%����ȓI{�@���$�]PC��ä���%��"lڽ1���Ɔ�P^Շȓ,�1!g"̺[�&h� �"O��ȓ>R��W��$r�BA���%#�4H��!�8Ê:v�@��Ս^Ϯ�ȓ2É�Z^��Wg5��a��v,�!!�u��v&�>:��ȓ@����P�ȕ:�~�2��G:p#̵��*�Z`{���W�$��+�4z�"��r���Ru`Fk[xDBh9=�Їȓ3�R4�FBǺ�E��gӴc��̇� 1������7R�5lU%F0���l��̰��@$�"��$`�����oQ�q�d����!uE������D�d����l�j��3 �3e�LՅȓ�2P�u`�	t�|9�)̭iKȘ�ȓ �<�d�^������,(>���e�s�+�1S�Xq�C�)�Ć�QX�Qr�7S��0�B��B����ȓfR �f�W-3ޘ 1�T�=��ԄȓpŊ�0���Z� ��<l��̄ȓh��<XB�5�]2�H�Y9��ȓ,r*i�ghly��] 1�,d���� X�>pH���ǿT������{�,$"!ZR��;/�r=�ȓ��0�K�^�NL3�(ǾM�p��ȓ+_�����i�t��a\?|�m�����B��P�pd:� ��v��نȓ"_�u#��Q�F��\�;�R��	v�������.���� �L]d4�-�;D�}��<D�p�H�eR]B��K';	8�q��/D�P����'ZR�����\7I0����+D�4R���xpnEX�+V�m�9��)$D�D�򢔀4t�
�\� Ai4-/D�lc��LE.��fO^�3�����,D�`�V$'pd+��9,E��Q�?D��D,P�
�ɫ6B*
t� C#c?D���獢1�mф�@,^����<D� �4C�/6��� C߽#�:���9D����LØ2��g&_FP��+D�d�0%��O"�Q�°$�N��D*D����U+&�@�+�ø+D�z�h2D��@!#E	\��9h����D��i�O@�=E���&&K�0�B)��\4�e�R�,n!���[��z#� �y�Æ!;P!�� ��Y�~�<uǚ4pY^��"OtX�V��
7ܞ�a�����"OE(҆�-��Q���ļF}JT�e"O��#�R�3�n�"6|��
�"O�H8�����Xx�MHSqfi[��d�O���Oj�;w��J���HE
^�*��)��'�f���o��'R�;Uo��z���'���vNȝM�f`�A�ϝw>l�B�'��ҍ�~@����}'���'��ybEAV�0���*�v�r��'l�lR���<E<��۠=F�8�'�l1���I���H�� ȄʓB���`u��u�fZ2)�A��ȓ� )�S_ N?2(��н]�bH�ȓ.��-��
Y�*�hѓ"U�I��`��w)��
'.ƕDڬ	�#��}�X\��e��c��ͣ~�$|pփ�)C�����!��!�Q�ld8�b�*H��'����ԔȠ�ϔr< ��"�4؉�EK�"�I��T�Q�Xi��:��o��8�ұ$%�@���v��%�@�L�~�J�z�W5�F���G�Z8�ǩ��_r�
҅	'o�9�ȓy�ع��,q��)�ACT�Н��FN^��$����Kw'�G�ńȓzLnMI���-+���E�T�9�*��ȓ+/ u+A�L�_�̱�MƎ%,B��(�����#ƫLR�1�JF
6�0y�ȓh�ɒCU�3��pѠcɜt|d�ȓ-���!��T�P:|�6��(��`�ȓ����݊a�RZ�KYT�d��ȓ5�d*D�H^d��ɲ�#F�rp��/��Mң���X,yA�X�F�h��!���Gɋ&r@��x!"\08a*Y��af������<Ft�H�c�*nN��ȓR���E�4%Cf ���>K�4���3&hy���	�c���ӀO�;gH���ȓo�X�9S�БOs���զ�7s�4�ȓ�*PbG���OCL ��O�/O�>��[8���5�b ���.t�61�ȓ?N8=�P�S4(�ڔ)���&)� ��-�09�`/R�Zd��OH�Rt�Ȅȓ3�P�Q�`��n[�$r4GҊw��l��V͖�9���%(�pm�.R@���ȓ�(���۳_fB�i�CX�ZR���i�����טPÎU��<�Ե��/֩�Vb��6e԰i2jF�%���,��+0'�'wV&��t��P �8�� >%9��ɿ/�0��M��5�ȓT8��r��';��p���cq�]���r\�`�_1I@H��I܁p��ȓCӰ��rLI;F*�s�&A?yVv=�ȓ�⭃�K%P�Fh3H��(�ȓC�|��$��!h�-��dQoR�!�?9���0|
֠R	3����G.!�H!���d�<����K� x�4Ę�r�DXaHa�<��	1o�4	1�b��*�[�<I�쎀e8�m�T"D�F^bh�L�<1A@�1)����#u���(7�P�<y�*�^������S�
�8��[W�<i����>�|��X�u������m�<��%\�J!�Th�"��� ����g�<��ģ,�, ��l�	2@ +w�]e�<�Ύ�kT�(F�ֶW����BCEd�<� ���ĕ!%@�h��J�q"O pAPf�o�J��P�!s��0��"O�ݻQ	�e����m�x�c"O2P�[6~-6��cϜ-O�� x��$�O���IB�+�
� ƕ�v� �X�aȋqў���I�+(6Qi�E	�:ؙ�l­w]B�IX�D�KEN̋} ��P�E�1"2C�	�K\1�rO��hXN���l�<47C�ɪEEr8�ǃҋq�,* �R�B�ɷ^k���$K*d���J_����$h�P��f�.1 4��$D�)�t��'&)D�(�f=R�|��%��g�(�4n(D���t�:WF,�aw.^�
$�(�E!"D���r�TyG��`�%юyK~@h�B>D��	h����Q5R��K D��2�J/��aJ�P.t�t��g�0D��!�I7s��PǪ1Kz��/.4�x��Z3(�$��9	�����ψ|y��'��83�.i��a�FĔD�FHH>I�
tC�O�z�V�ZP�òY��X�ȓjɖ��p�O�D�4-Rd̗�~ނD���"�z���vp!:A�"Fв$��AIEK��kr�ꏢG�Ω�ȓO�f����?����MJ�!-�=�ȓB���)Q�+B�Eт�	�hh��7<�h��C�>���!$��bٕ'�a~b J(�4�^�����%�K��yb�E�'����,�X��� �!Ƅ�y��FD\q�߃}z�A�'�5�y��Υ���G�6f�\]b#�'�y2�~n��;)U2�� R��5��x�V?z�� �#Z$�("F�V w!򤚧zh`a[�j�-%V�E��MS!�$O"S���e�*h��%`TJZ?!򄞂<6{���8}N��FI>X%!�E�m��L+�  �(�V����A�!�d�-!`T��V�=/ڬ�1��
�!�dD�l2�����X-�\J��n�!�Ę<Z��}����;��S@����!�H�xX��)'�_^*�k�B]>�'a|�!�2�	�B���ta���C�y��firAk�,Y4��`V�3A�����2U���ȈDp��#��2<(�%�ȓV �@e|o2e�b�+NZ����}K����:b0�;���*"݆�Bs��2�2�b���lI?��5E{2�'}Hq���"ŜQB�&ɶ&錐i
�'�r�Y��u9�	Bo�H@��	�'h@�5��7\��A2��F_��I�'�6������^)80�7C�<KHb)a�'�L�G�Cz���V�š7���P�'$b��ˋ*k�"!3����0�ȓ�(���̔�_���Pk@�6!�M���g~"�E0��]����8G2\������y�#��^dɁ�P�A��qS�;�y2���J5(i�H�#���y��č�y2ⓞ)V��3��Уl}̵{D���y���g�\��]�9�S�^�y2�L90���YS��]�b�s�I�!�y� P�f��$IfU�0�7�y��2n$f��*	�����ꘕ�y��N�4U^����*����V�y�e
)W��!*2+$�L
w��5�y2�K$Fh��R�#'�𐖠��y
� <�i�f	�����S��}�"O�ʅ�^\Y ��BjR��ܸ��"Of�1GO��V3*�0G��-t+����"O����l١�(H��Z��"O<āGA�$Қd��C�h��"O�=0�G�x��A�U�Ț��Q�"O�l9��'E��P��n�L��졤"O6�I��);�O�	ƌ��"Oz�ە@O薌I mηP���E"O&H	�
<u� =�a��$4�؁y�"OL��u��>�n
����HC�'��Q��Y�lA&C#�T�C�'����	�+�<h� �ن�p�J�'8�"V��',|���k��?�Y��'�p�iVn��3#�U��c�;}@�r�'�$���ʠDSB,3��i{	�'jN�̏-;9��0�mK((qx$q(O��OZ�}��0�����,h�V	�0�
� �vm��~R>�C�֘[�n��%�E�5��i�ȓ��WH 5���x��4 7 L�ȓb�p�kaF�W~�`A�%6�ؠ�ȓ^�zYi�P�.��$��F9W߈X�ȓ�r�t��Q}¬�U���ȓ@�D��'�S&4�TMIV�ͅy�����|����z��# �|�@IAL�
�<�3�8D�0C�;>�:���� 3LLu"��!D��R��%CW�y�aO�"g��)�&%D���F 9ig����М�,u"��?D�\���ڷF��PY�G�%n�b99+?D�dK��!`�S�MO�3�P�<��Vy��58fFE�2�ҒUݲ���(	�˓���h��d����%�ʎvevP���K3�!�&!�T�� ���Qba괧�&�!���K�>�[�ށ�l�b��R�!򄖉}vޠU�3>�p 
�e�2k�!��R����d-N�5δ��E_:Kp!�$�q'.��E��� �T<c%�H~4�O����|
�O7�H�gl����Okux1�	�'*H|� Ɛ�j(�%�>s��A"
�'8�q�������T���d����	�'qt��e�\�N��Q���Z	�'�������z�3�o P���'�
D+���Xn�a�PH�y��er�'14��G�^;\N��w�FgD��[��'����|:P���<AހI��>'#�0�t�YV�<���4f��kd˼Q��¡)�{�<����96pMb'�ܶ�J��db�a�<��c�gb��(1-b���֍a�<���
�%� �It�S�|{�$Z���E�<���I�Lø�1��V!:�)��\�<a��^+Y��W�&XZ�Ы���X����$2�
S4�'	�*IwA�A)�v����L�H9���ߍ~Tb��v�4I����족�˙',�e��/Hz�u�ȓiU*y����P�b��,��v;Q$/r�A+�.5Qsv��v�`-�2L��1xz��f��<{j	�ȓPa�� @�	<؂�
f/5Hp6��wwr��-� �N�ʑ�J Dx��	{~r/��FF��.֬z�b,�Eg���y��� *)R�["Z�m�}�u��yb�޻#�L5���ߢ<�"���Ԅ�y�h�)��X9 �K	0�@ѣ�T��y�@�L���K+��<��^��y
� T���D]D=�� �r��D"O�r���:R
�q�N�O�8EQ'�P���pO״�8��ݫZVP(U�"D���#@�=5"��P�`	t�*��Ӌ%D���3�I�yn���#�9v�u�1D��x��ޑO� |�F�\�Wn$��e�;D�Xx���'_[�y�CN�q��AIt�.D�,y��L+XB=#�M־�� pv�,D�p�ć&-������T��`�!+D�|�W�S�(��,�rL�+�\\AF*6D��`�D.\��4��H��I���a�9D�\I@e	�B��z5��n��D`F�7D�<R�n]4䜌���D �Ԍ��+D��R����d2Pܨ���#�b��7 &D�䨆�E_E���~R��ĥ$D�XQ�
Y�V�l���I����O�OC��<^�:PR4k�*�@�
\abLʓ�?��_�l�i��J�6�bF�J6s�����;-Dp �kL<6H@�鰦P3v[��ȓ`�|%�E/\���m-X��9�ȓ~��ɢ��Fa�LA ��"\�Ru��%5�łBJ�V<�F(	H�.5�Ɠ|6L��*��n$BD��z9�X�-O���΄k̥��&,�)��r���d��@��g�P��m�4�PCY��j>D��0j��m��p�Z�~�t��i<D��ئM�q�H��$��`)ҥ��.D�� Eǫb�\�.�!�E��c&D�)3Ï7�tA9��x���P�P����
|�i�E� ��`Ѝ��/�B��ȓlt��ࡗ0Wit$z���>K����?����hY ��>ju���|�x��ȓD�t� �N����(c���P��Մȓ%�x��$Vy�4¤h[�e~ƀ��ON��s��ܿ4���)ѦC���d��9\*E� b͌Z�,�	�G�*3$���;2Hy���Ѻ>�lX8�m�K��<�ȓb��h�F�!M�`��fL;I$^��ȓ�T8��M�NV�����P�x,Ԑ�ȓ���b��8��t#S�l\|(��nވ�G*��.���#!S�i��V�qr
ز�L�@�&�n��ȓw��!��C�":瘈�g�U	��ȓ&6����� Z���t��+���2A̽����%�p���<s��J0,`#  W.:� ���$ȦspD��tY��"<�&����8t4��)Z�L�����35���k*l�&u��8bPia(߂?1�ET�/���ȓ)�]Y��CQ��bǂ�@�f��ȓ-ty���¶ckZeK�(6X�l��B-�A�R�Ń} ��f�浆�b�����V�zAƠ��(��9����P�c!�( �<�p�®E����!����J��~R�*E��O5��ȓ?��bQ�ԌZ�푫l}�	��=D�d�"יTg���O<n㸑�Ԇ<D�Tz�G���1:��M#<�X� D�� �J�U�݊0e^�{�6���@3D����НK����U^4,�;D��zTĐ�?�y��[M]���p�<D����fG,F�i���x���:D����@_ �4�����<���,D�T���̃ ��R2*S�z�����'D�� \5b�gZ,��H�!��W��X&"O��jq��kײx	Ȍ<�Eb"O��aW�؈��\
'���`E!�"O���`�kE�Ih�+��f�ni�"O0��&H���B8�d��H�@T�%"O�Y*gؗA_N�[��#q�(��"O��b� �1��3��;����"Oʽkw���4R�J� �F&�"O�M�f��bӾ���	=$#f�:�"O"�A�38�С��)��0����"O =�W@!~)�acwȌ0Q��
�"O  �e�.|�LqP�G�n}ހ�"OĜ�p�[�&���K�M��ڜe"O�`Q�i���R޶	up"Ol��7�H>4��D��ܦP��qxV*O,h����n�ؓBX�[����'K�0P�� �% 2J�K�^)0�3
�'�!���:��@�$O�L���A�'�\EH����x@ C���{��a�'�=�7ˇ5�V�*7�ԅ!E��'��h�ӧ�1A�����o��ɒ8�
�'��0��K8��pHV��&Җ��'�fi��8pB��u�N���9��'Uz����+&�����c<�����'��l+���g`�(Ί�}�`�
�'�� 1K�洂�'� z�j��''�<�vn� l���e
V�>��9#�',�Q5鏕KA�c�[�3��l{�'�r�YG��N���k�ȇ0��
�'�M�$c��7]�(��7��i;
�'ؚ�P�ٌ
z���Bҿ�0y��'b.U`���@���N&u�K�'�r��a�Q�n!�E�į@$���"O�� ��Hq��d AP�F��""O�@�ZR`��8��Im�� r"O�p���E�f�z���N9vɠqx6"O��؃E�Dj"u�U�����"O���GcX��u��&؀|�����"O��0���!�Ba�䐫+|x�!�"O�����Py����7�E�x�FY�W"OV����x)�!�!{��[�"O���W���-� ��0����@I0"O�,��*ޭ*�)�Yp���"Or�Av�?�8��l�-�j��"O���/F�e����V',���.�!��	��hc��.h �� �ϑ?2�!���FC��"�Nꄝ�A��~!�D��tE�,ƥ�;u��aVMV0,i!�d!ݴ�ㄨ~�$�� ��vq!�$a�l%�foR$a���c#$�>5!�Ę�@�\�� �S�>��DIO��!�$B�pU0���g�rYR�']4B�!��-
�x���k���AL�4�!�$2X7����ÓXʰ]��do�!�DF�tT�"��\R��p䋋!�$Q's3�!�hY�RV"�#��Ppg!�C� _�yjflN��񁓠S�-Z!�$~�"H6K�8I'V�!v���A!���0t�z��-�>'�U�r�Z�9'!��DQ��e�G!2�~$8���!�ė�5;A�#�a����!t�!�d^��R��J�NҀ�U��'�!�7k�
1���N�Y�amG�r�!�	��&�9�L�m+������!�� ����APT�,b"D�ar��S"O\�
w��=+ؼ�@@Ǥ8�Y��"O
T�d*�3L��9Ơ�[o�	�'"OP]�q�Yw�l�UF�u˄b�"O&��3 �<�ly+�D�_��P%"O�)��,� C����PW�Yl*ȑF"Ob���")4G��;��zb�"Ol��r	[^u�À]|�: a�"O�ڠ� �{v���Z�{���"O�p�q���������C�"OL��Z3�RܪԢS�Hֈh�"O"����2����'�b*P�� "O�*Q�.w�DY��f�.I�=�"O�{�䁚0A�2�f4<кm "O��be\�4��kA��:�N��$"O�E�C\Khp��@��z�n�g"OI�'�\"��q�" �p�r��"O�<"����5H���-���H%"OPdud��
$�Qɀ�˵>�j4I�"O �3�HЬO1t�a��1m`NT��"O8`ꡈZ,0G
(e�$S.�(�"O�𑬁J�t!oD�"CP��A"O�qREʴc/0�nV���.!�dг<U�eB���F�b�͌�Ar!��4�L��É&�R�X2J	�4t!�dP������#�l�&�"?n!��Û:�:� Њ��z���ɶG�!�ʶ#������9�Nݪ��W�J�!�d+�J, �dG�?�����9�!�dڍ]������#5�I�|ќC�I"�����ŉg�Z�A�41ΞC�ɽ"H���i�-PFDxD,��yP�C�<T���c!�̀<�D Z��̨u8JB�I;x?�Y�K�;m���g�~} B�I%d�x��_9Y�������,B�ɯ�ua��	y��qXE䋳R��C�	U��M���LI]�1�E�՚5�C䉪wU�x�&�M�	%�� �m�(#M�B�	8�t�5(F��X-]P�B�L��K��	.Ek�y
���9d��B�F4�	F�42|��1�jB��,th���z����^�KDB�I\��T�h {��ȆB�I�lݪ�+�-�(b�.�B�C�>��C�	+-�ʩ�Ն�d��8�PkT|��C�ɚ4!����P������L�<B�#E�Q�%]�NR�q"a�1o�B�	�^�HC3������Y�W�p�
�'"���[b��h�こ�L�RU�
�'�6b�![�?��`c�o�(}`
�'�ؐ�tgY�`R��˂�:gI��'��R$�=,���Ɨ4:����'�H���Δ_����"Õ%g}1
�'.l�3BƆ�.�v���l�P�*P3	�'b%�aR�y��i@>'�1��'y���sD4)aLa��QQ0pZ
�'U��R��6c������)�'����4�_�.F�asA��-@{�y�'�����RA]�0��j�6�P�J�'<����X?m���uHU�𲈘�'s<��_�$�z�c�
(��'6j�X���	��d��|�~��'��I�C$[�j I4�;?��k	�'��mȤK]?D|8�� &������� $�F�&� ����p7���c"Ox���|C�\�#�Z p��e"O���1NO�,L��Џ!���"O6D"�ƿw"�A�t`��-�!�s"O�ڰ��IPB�ޤR�`hw���yB�<����i�}��|��K�y zIr��D�ܼy�A+�䓶�y2��bY�!������F,�y�'�<.R��ˑa�,
�R%*����y����d��P��4�����G܁�y"j,1���6��*2�2����ԅ�yR(@6�^��d΋�3:�ٻ��O2�y�H�sP($jsl�#�2���e�yr��/{ )����!v�8�a&X��y�K��N�LMP�΂��	8dJ��y���0:�u�P�E,	o@�ϙ�y���6��2��(w]`Px�R�yR�&����Իpx	��!�y����1�Jv����1���y���y�v�9P/	��\<2�*�3�y�c��x�0�D�ا'��p������y  n��p�SZ#:�$��	R��y�D�&<��qɇ`
�P�V��)�y2.5�ś�G���h�㛵�y���,&"X���ҹK�-ڤ��yb+M�e�j��emw�ޥT�� �y2��rȤq" D4m��v�R6�yƃ�?��8���7���p$�y@�sV ɷ�"6���qť��y��]�v� �!����3���;�F�2�y����m� O����ˤ���yr��i����)
#*�&�Db_6�y�
J53�̸�b�&4����ȅ�y�Mߖ2�L���Z'O��9��]>�y"fX!¡��Τ��Ȣ��yrK��IZIzw�:��l�bJ��yn�@�I`��{�l	�c��y"kC�	a����\VU�vJR��yb�%AY���3N�조ࠋ��y)$���I�<�������yb�D )Լ���������#�yb�u�ƅ�'pq��E�y®�6�tzt�+��� ���y�$A��Y��I�|t�u��bX#�y�d�2 �R�FP�pN��xv%�1�yb�V�o�h�&�e��� K�y¨J��ġ�N?aI�]pS��yR�;A45�J�.��H��E��yB#�u�xpG��[` {�n�"�y�3a�:AY�C��y&�)�	�y��ߖ5����&a�����SsϚ�Py�
�T�#���J?@Z�ώV�<A�Cӊ_Ȩ���<�l�f S�<Aw*�'��C�B
_�i�T�GZ�<��	+,���xRe�2[�j帆��n�<1�Dk�V���o�+���`&Âi�<����*������'t%�� ���N�<�P�^z 4j�l��>?"ٳ�L�L�<y$��H33�Ě
K��1G�@�<�s�ɻBa�3հ!G���%�Js�<1C` 3>&@Bb�ߑg�ج��Gt�<9dKI2)�B	���P������m�<��ǌ=ҡ���D���ف�h�<aD$���B��Q;y�L9�&Qe�<� L�3��֢R���%Η�
IDE؅"O�m8p�N�<8��l��@��Q�"O��2U"Ѥ	|�ja&�T�~��c"O�򓇙�Im|b��w� "O��V��˄�0t*_2|�*��"O9��m��ZEkħF��"O�8�6�ƷJc$���L�D�N�	�"O���E�^jr��&�L��,+!"O��sՎ�q�܄(c �[�N�0�"OZQ��iT�����l�
�zW"O�-Y��9
�&IU��'Q��8�u"O� �Ů�d�[���2ܼ*�"OR��d+ݐ-R�ݲ�o��e�r%��"O��	e�׆\�Pq�`E�-�j�:D"O����e��d�t�p��Ђd2P=�2"O�ZW�P[�j�H�)S�Z.1H#"O���2혇�XE9Ї������"O ����F.���>T�N�yt"Or 9BOS�7�H �D�gODm��"OB4!�F�ґ��B8`>ʹ�s"O�X1�Ŏ�$� �JD��|�`B"O�1�U����f	�:R�`�G"O$�[pkȕFLFHq� 9��5"O���e-�M�,�zfCH�K�8�"O�]a��D/j���DN�+�dՉp"O.���
c��#�⚣2|nثS"Oh��pG,<���7Bd؆7�&D���G�V
��Z�LX���ŉ&D�h�ǧ�P��rT��G�\5�N#D�pQ¢�J�� � ���i�$"D��)�$�2,��9A��M\Ҵj!D��uj�*��؃�ɑ�jH�V�)D��&��>64�HD�.;ht	f�,D��ą6Kn킓�ěl��H7�)D���L��Ҡ��3-X^���!D�@ e߇��Baf�
I���0( D��Q��A�<�+�j�9�q��+D���.R�}ɲ�Q�
H��|�6"$D����9��׀�8W����*"D��ba��+�M���8D�|b'�-D�ԑGc�H�h�X4�7V�q��-D���sR9v��ԁ�`Q*kV�ԈS`*D��P���	X�5�'P4
z��J0&+D���#!Wy؞H�!�_j���'D�8	Aa� E����HL� �P��&�&D���gBf=�P+�.��%������0D�@�w/�>O�a��D#tb�9���0D����P6�T��g�]*j'�d�G�-D�@���\�*��K�k,X�!�i-D�Tf���|��e�4]�py�%D��n��m놵�P̙�GN�b&A#D��@���:UM���T$�2R�� D� X�c#iB��Yf#O;�
���I>D�\�#fS�/�b��F�8򶀙�'>D��H�@ע;�H�qFE�j��ؒJ?D��@V��]A��[1���r��(8�d>D��(���N4��(����,���׮?D���&b��Ea0,�㥚 +��q`�=D�عdMۛV6�� T�>r���EN=D�@[*ǜg� �I�K�fR*m��.:D��B0�V3��h�$�MO�`�,8D�� �#�6
P8x�j��|���0�6D��h7c��5�F�H���L�F���B4D�|3S,�"|`� �D����$7D�� �l s�3�)����za|�XP"O�� �AJ.#>��cd\C��0�"OZ�&�Љ�IZ1��.s9�=�e"O4�8a'V�v�Z��ŭѠ`%
I�0"O^$�%�Q5n��騶��:F,6M�p"O�Y����.5e�5�������"O�m�f���
��j4bf"O�0��H��d��$��l��T#�"O|�z�B��W<a
�dߔNE2�"O� ��'�#?�0�I��=���{�"Of��"S&㎙ѓGA���[4"O�p���F�lL0�Z$�T�gB��SD*O�1�J�6B��h�\��TmC	�'����o>en���M���M�	�'�՚���P/D�ITc�
�����'��LA㤉 �v]Q����xI�	�'v����H`�c�E49��S	�'r�p�b�A
pyF��� �H�!	�'��@%I��q�E��	ML��'\�	����1��t���3l��'��aP�ڹu�u�4�ъ}%��:�'t�-p�ɔ�<�|�n�M�r���'J�8���iz�$���\9���'��tXF�=�А�6k��5;�<�	�'��D qH� D�pt�f$My^� 	�'D��A��-@�}a�c�.E��,��'�|�(��OHL8TK*�\�B�'���8/Aqzļ!�g�-/j��	�'�l�����-V���4>�`�y	�'�H;��:4�H*�P�:hq�'c.@P���]¨������`�,t�
�'t��*��F>?�!gnQ��j�
�'�F��&
�)ف�@]Y�@h
�'֘񐎓7jԠ�-I�]O�]��'/p��`���krmTaj�A�'�H܁ө 6pA��a�I�2���'tx��S
7Z�Y�pk!� i�'ڤbv#ݨSܨ�B�����lQ�'\xQ륉��/�$1�RDΕ|40���'`���2�O�+x�IKrdO�c7�%��'Gt�J�'mrf q��V��<�']\��#���9�a㐿�\���'�h)k��X2,��0ao�v��A��'�P��D�U���KA j��=a�'�:l�T���Y��03�Փi�Qs�'D�9�r�ݘdB�P�NZ�/��(I�'�,PA ��!^�Z�Q�L#.�l��'=�H�,S Q"n�HRA%-���
�'���¤ �;�H��dȮ(��@�
�'�-���L�h�x���A%$0L��'�D��&��'�%�O/�x{�'�D��ĕ�9s��[�iH��RU�
�'}� (��G��aJ����9
�'_PX���U_:Mr�ɔ��i	�'���N�$�q��	*G� �'ւꕏ�=jA|�b��F�#�X�'�(p�Ë�'�XcP˅�+��I�'�N��C#N�.��;n�'��9c
�'*V-�D �vY�A�Ҫ-Y�5�	�'�F\35�� ڢs� ���%��'h���4,%�(�H33�`��'~6lke��+$��pt��W��Q�
�'f%� K2aG�ir��D��
�'�1�L�E�D�) [�Er	��� $D9R���^����cd��H�K�"Ob����V�b|�P��l�^L+�"Op�q�*t�~�p��[�X�����"O ���d�(< ��@�Ə7��"O*@ b��f
�5k�e�:"�C�"Oм	�E�h�X�d��r���@"Os���"[֡j�?Pь0�U"O\�����$ie�F�W3H�F���"Oޜ���=���Xя�2u��`�"O�hQ�B��m���`�K�v�pu"O4&l��y��T9�8~c���"OF�Я�%���K�lL�]_�"O�]�&K7Y�%���&Qhj��A"O����p肶�J^��5"�"O�XZ5lW:sT�ö���	���r�"O�@ NB����C��4�=z"O���ȇ%S8��j3&�75|�(�"O�!F���#s�	��'�3��V"OKB/l����Ť��A�N|���C	�y"�K#�Z,H���=Z�t;vLS
�y"�E��vȩw��0�,��#�y��4;#���!&è�j!ZBOC��y2'M�|��D�A��pp�NP��y��N'̙��W�4����,F.�y҂גt2�K-t��o,�y�$O.��I��GW u-��ꂨ���y�+Ғ2�p��R�یv�J$XŠD��yRHqQfE�RAP��9�CNH��y2�߉T���CK��J��FS��y��P�u�� ƌS>��QT	�7�y"�+D�@�JV�H�j�@�B̈́�yr �@9�F�O�dX�y�	ͽ�y��QA�4���Y�[�\m�wO��y�d"��K&��/T��12����yb�N.l��ty���9�@�i� ��y��>Z�y�N#Y$=��Z��y�Gpa�J�A	�Q3���0�����'��dEGP�(�s�ٶ%�ȉ�'R�܋��.G�&e�EVlk��K	�'1�d[6h�zb@X�A�*f��<��'������(2us'M�9[lʄ�
�'%�<���4aꈙá��`���	�'X�H�!��1_	&XB�j�_c2�R	�'�z\�-��։ipN&Q2�uI�'i���$�n����<J��<�'@밉P�}�d��sĒ B�v ��'f�Ʌ�K%	k�!S`E5f�Qb�'��E"�A���6���](bEZ4X�'�� �)
5d&��{�LP=h+ ��
�' ���&�[�ΘkQ�20\q��'�*@�ۡ;��uh�C?�����'��(㠜��|�"�δ]a X��'�\�qj�< �"lY�ט��'�z5�A�0��*�W�x��
�'$��!��A�/��d���.�x���'F���qd�$W�,�֏N}kt��
�'�X���e\�1T����'�����'�
lva�Gv�@�@3�:�	�'�,d��*[6���!0x�n1�ʓRH���uØ1���$b9?�Ĉ��H	�u�%�:n딴ZfB۹S�Bx�ȓj6���b,N�|�£oV�T����DVN�x�bH@C���n��H��D�ȓn�Tz��D�m� !��=����S�? @ pBa��IB �ajM���52�"Oj�J��!�R���h�5̢M�"Of�P��q��S��N�@��15"O�$@I c���3���>Ԫ�"Oʙb��O,W�	�*]m���"O���a�"C]�H`wV���qa"O}"v�� 1���sa�E��@��P"O�)s�O�e�:i[�
 !q��"O�w˝$Lo��롄G�un���4"O �Zp�2�`�գ��S1V]���Q@�<��M�2eZ�z���[���U
%]��	O�)�?��b��X����j:�PAc�<!D�L�m���a��LFʌ,a�F�C�<�)^�B^x���WP�\8eC�|�<��bҭ&�n��F"����c�y�<y�+�:�ly��/�\��� &��\�<��@��g���
1?�| �e�Y�<�Eg�>��w�V�Y�`�U�<�����D\����� W�����H�<A- ko�4�G�� m$���	P�<���
v��-�P�K�K)-���f�<�E_(X{D)��8�`8�w��m�<!pN�;�ʗ�#�~�A#`m��X�>�f��>~�(��� 5�����)�D�<i���A�T䛧�H<_\	�'�Z~�'�?u�q ��;\���>](���(D��8#R	n��|��4#�:�>���"�0� Ƅ8P����^#V���ȓs0p���%'�J�#/Ou44D��:�jՈD����d�c/X,��4E{b�'�� ���v����!C?']$+
�'X<@2�j�#�n<At�0 �E��'�F�G٤�p�:��#%z�=R�'�.����G�4�TM[��đr�u�
�'Q��B2G�0lZey���&J���'�
0h��ٓf�����aT\"u�H�,��IC�xT����}q(]e�@L,�C�	9R� b��D�G�1 v�D/CC�I�}<: �aΊ�p4u:��ś0H8c����ɐ(|�4�q�Q11gh���	7�C䉬[��]�aN�6c�Zٙ$G(��C�ɻJD]`w��~8�ڴep�d"Oؙ��F�0��
�J��*iY�<����=��,(x�0�K��7�(t��^�<�Ph_�Q{6؁v �	a� ����V�<�r�\�ju��e"�_����-�x�<��o�N�Ը�b�?u��Y��	t�'�?%���)I��M��o�2H��R��7D�P����=@ 岴	��1���2�A1D�@@�K�TVH�����{B`$D�(XS��`8�������E(�=D����H����qS�L�M��ݰU�-�O,�I,Ph�P����6(%��2�bWv�v#=�'��>IBt�=C���酦�n�`�)�O��'ޞ#!E��-�L�(bPc��J
�'�(���C \�A�
K�0l�*O�"=a��5g5~!q�L>��r��@�0C!�D�-3�����cŊ��1Ԥ7<Lў�P��K�M
"�tQ���W:^�b�"OJ���A�ܨ� Z>:�a
P��z�OY�R�X	p1W�.l�(h�'�6��1�E�$�����kK�a��%�'�@�a@�2��A��gָ�^x��'�@�Z�Bž�8Y���0?����� �I��%[q��*�ʇ�H٨��"O���ːf=����G&8J��"O���1��/�"�+�ɜ�>y6,��"O��c�P�Hy"Ƞ�*��8a:�"O��zҢ��u��5�
�R��!�:O@�=E�dI��WJ*�s�l	�d�0m
@��yb�ԴP-ܝ���NmY�A)���y2kT��D{g�?b����p��5�y��ܧ8���pg�Y���P`Eگ�y�⛈�2�౪؍PR�pp( �yr͐��d;D�.CR渒P`'�yr��1p�T�Ö��2@� m˗FD"�y����Yi<a��%3}C��:�y�'�M�1R�KĐ��L�R�yb$��������x2�wLG�yrnI���J�E��aNQ�&E��y�%�\ҔQQDS�^DI�a�Q��y�7l�U���T�aF���pM���y""��(���3��5H����@4�yrfA W�F�2���X�N܁�@��y��_�	���tFK�ebl�p!!F��y�ELhml0B�nͧF��؛PR�y�B�m.IZ�+��=�D�6(U�y���*�Z���+��4+��%i�4�yR.v�� l�&3@4���F��y�H6X4�i� *��Յ�y5L�b1��0�xk��Ǚ�yRD��~$b"$DC�l|�:��\��y��/	�܍�S,U&]��������y"OǜC�\8������P����yR ���K� �>3H �� �y"���2:6����C�#9��r&^�y�BV� j�E*@�[�6kvF���'5.t*��Y�$�-`F�+\��y��'��͑S���g���'`�L���(�'�H:��(GZ�1;���<�<��'�؈�h�� � 
$�A/EU���'E~�����1��`�*����'e�9Q�Α4z޸�VLO�$ê�'~p���ς
��ӕ�$n��	�'�dkAZ�8`�M)��V.�,�Z�'�L�qa-�t�j�r(S)��<��'���Ѥi_�$��`2�<I���#�'l��{�X
7#�-p���?�l2	�'Nlآbu�h9�Ƙ<���y�'r�}�2�L�æ��,�+,Wn���'{�y@e*�G'���ƥ[0$D���'#JM��,ޘR�,�8�dYs�8C�'�>Uq�0@��F�s�((8Q�m!�'W�ŉ�ڨ�@��Lϓ5z(P	�'�А���:!hF�Y�.��,��'@\ݨ���<t�B'� $�<X�'$�<�5&	�#j� ���s�<Qh�'O����]�x�8���N� �`���'G ��aG߃t�i��V� ˒���'�<�#��A�	}�Z��ي��tq�'H>\�UDN'%�(�v�]5xj����'��بp�J�s��`���\t��p[�'���O^H>,	a�Èw��	�'��#�X+�$)��-�0�X�	�'���ˢ��798`kL�%;�Q(�'���òˋ5E��!Z#�� 2����'h�����5Z�U�+���`��'IvA�cM�9~p �`)ڜ6|L���� �!:��@�7H �4��	h��"OdXB@��N�X`�0��J��݉!"O��J�-$n�¨S�៮h��@�"O�ݘpk�P����E���"O���c@�w���P'�S:f"��"O��8�+JF#���5�/h��z�"O�E���E[t�8B� ۱*��� �"O�0�Y�y��]	dbƧz��D�"Ot���%O�JDH��c,� "O<� ��T�h'Z���f�<U����"O,<x�c�# ��5pƜ�|FPd"O���$ 0�С���'xY��"O�a�eJ0L�`(Qe�ޢB`�V"ODЂ�A�y�F�©���l°"O�q�r	�'�05Cc�F�!��I�W"O��Z����� �h��JN��y"A�'z����U�f��}�����yB�+YbY���ϕe���Y��� �y2j_@�hf��g�Q�î�;�y���}�nK T�S�V���,��yҪ�������F@�P�`�!�y�Sl?������g|������'�yb`J����J����O�\���L� �yb(ˎ@�9�#@�B�b��E���yR(��9?ꈡ'��3;������y�Yd�%� Ђ;a�l��m7�yB˘�A��7KP,7I�T�����y���+9v�����+��0B0��y�&F�tb��	Th�VU(�B�O���y"L���I��o˳L;pࡃ��y�:]�q�CX>y�H�z b��y�kޚ��I7`K�x���h��A��yB��#��p�ړ�-�ge;i���`�M��0?ɵ��w��h���N�5@ihqC�r�<a��	o�t���-=B����j�[�<a�-�	�(Y����6����DKl�<�F��Q�B pT꟠��y�m�<�REW�P�@,�G �!#�N�0G&Md�<1D M.��R�[�o� ���c�<) ��S�U����0`�|�R��Z�<�E� F����\2��U�#�Q�<���){`��G/ݯ-�Z�Hu�<1��)G�8��uj��W��Mbd'�o�<a1C&oh�0�`��nE\�Z�fCe�<�eAB2+m"�����'Z��a�z�<A�n��,AȪ�'B�i;Z�֥U]�< ���/߀��g�E_
#%mLg�<i��	�L�f�A%��m��=��ȚH�<�Vd �1ؐ%Z	L�X"��D�<y�I�J�T!!J\�:�@]�GA�<�՗��\��8R��j��K�<�ը�Nutt�"�8� �q0� ^�<�@J�$�xe+��YoܠYe�c�<��f2s�x� �� �c���1�KZ�<y�eN#n>�C�Hv�\�Q�I]�<�R/Q-D>b���WQ�6|�f'w�<�3��#>���`T+~� ݀a$^s�<!D ۙ(&P�"�\.:��aYD��g�<�K�3Eǐ��dl�Z��Ѐ�j{�<iCP*dM�e	�ɝU"�}BC�j�<�g�Y��\*E��2��"�%T�D���ƲM�fT��`�LZ�YQ�2D�����Q�{Ĉ�Ivx��7�.D�<����eْ�����|�\"�f/D�� �t{���4lxw�(�,� Q"O~2�O�@N8��O3T{�D��"O�aY&cݮς�;���)hQ(�"O
HU`�kî�� -ú,D2H�C"O��BW�@�qR �1���9@�5є"O���B/�6�
�)�yF<��"Op0�5�F3E�R�K�ОB��ɰP"Ov`
S�S���Iʗ'�?ky��"O� rc��"�6,�����f���"O�4+��B�Sy&�"F ��]�����"O�`!�aû*B 9�O;k���2�"O��ńG�*7�{R�N�n�(�B"O�\�F��8!ƍ�A�� (`���"O�$���J`��i$B9J"O eG�<w:d��O��`���"O��R�K���eX��J?��ܒ�"O:Lũ^�M�=�F����"OP�����Xul���ڛ@�x�5"O$511��\�tU�2E�O
 A�"Ob1�!7D�Ȱ"���)#"O��8��X�X<"��D��-�F�W"O�!�3�F]E!���1v��5*2"O�9"!�O)���A`��uҜ��"O8A�-M�k�1���k96�"O�j�1S�x�NG�/p��"O��I��H5���с���)��'��P�G�a�S�O�P̛�O��vo���1dK�`Z~��a"OX�b lA �����cV-2�Ĳ��O���>�ny�	�*�f	�d0%h���㇃&�l�E}�IJT�	=|>d�I(�`YcT	"�~Q�w�N�6`��ЁL "E1!�TD<`!��)"]����dR��� �Ԃ��:�X[҂VA62�4ZR1������Ǜ2AK��G\��́]I!���m�(�"��x����~+�,���ۀQ.��ߴy���? �BO�z����O�@�&94�v��&坴2���"��$�O���EV�_#�� ȏ�F�dp�dF�
dÎ��1'!a��y��FMa� ���vz��'�D�@k� �`�5f��Z�l<��P�E����w`��M�!���z9�QH^4U� !��Y:=�����'�DŐ��\`��C�ɵo����`�-	��S �7H��jk��d`�)��CE�K�u�Af�+K�(�`Y|��<�
�p��K16�@�Ѭ͉ �3�"O�|K�K.r�dm� �҉, �T���50��j�W&�2��2"�%X��4�K�p�jM���S( ��x�A 9?�=�V�M0�^���I�F�ੑ��\	5��m#�B��������>zF��p�](©��J$`��c���uY��	�lj$����:A��!�b�;f7�c���.Y~���Q��)�]��
Z����ˁ��`�QC*�o�(�v	��A�"݋f�֟4����I�D�W��.d�4"�aP�~�d|�0dN{;@�B��A�@��M��E�l�'կe������+��� �n��"E��^Dt	(qDGw�'��@铨��l���,����"����P�v�۟,�|�3���C
`ם�"��Fg�-�T��Z�h��&<s����w`�Eu�l"UEa�����yqO���ɡ�U�T:�ɐ�K�oX�Ѷ(,b�~a�����q���Зf��i�4�z������ɱe����g��*C	4��AD���T�D�QlC�&ds�^���7m�
=�uP$��mΆ��@ҖW�I�Pf΅��(��耩k,a��G Za{�Kp��(�"ѤyXǏL�2���Q�6�t�x�{����FO9\�X�Ѧ��@�A������;`�F�H2���:C��)g��Z��F|2\
C�D�TK� �uC�eO P`���	M��" �sU�<B��ʟ��\w��{�ܔ8�X�y��>q �ݘx0!�F��2�đ���<�W��#l���;��h ��6%� 4
7F�=qeL�C@':VEpf Ԓ��6�L�|��g�+
�
�J��'>F�;[Ԗ�ȅn�5w���խI�D
i�$����:4P�K���<��B��eKB�xe"��$`�`�`�nJ�TB$#��_H<�p�X*J�a;�l�8m�qʒ��b�_�$��S��p�gLU	$��.eͻ|��:Bn�!n^�˦.	�%�l���%N��G��Y�`A�� ONj�n�	^��t��k�.n�h�'�6�� C�b�e�&9���h,H����R&�ȸ��I	Y�L�C䗛R�6er&
�%�μ�ߔ=�61���g�!��U
|m�%�p���DkSD��Ola
�H�)$� Њ2�3� � �%�*X���#�! ��͓�"O���d�D�]���#���35��X��Z?J�B����I9��d9�g?ٗ� G<�z�{��('O�U�<q�]�N�Liq�F�K��	u/���?����AdX���[R�*�p��j"&h�㤝#�� 7�Z�&:a|b@�8(Ҹ!�Q�M��q��+�~���ʇ�	'.b���q�ѧM���Lek��ضC�Y�����H��(O��9�,go����ޑ٘O�j�!⟝j?��q�dI�X,�2	�'9��s�B@>=�Ҩ���n��0z��( ��KM�xӧ���aG�b�F$b���E��q�A	"D� !⊂!����)G�"D��"}2����A�鉉h�� �uh��h&����B�|�C�$����O�<,��AJ0G7�C�I�L:`0�!עd�����2c��C䉔W#����a��@�c�Q�C�ɸF�>)��̴X��\KqA�8]�C�ɞ4�������M��Xx�IP�2��B�I t�<�9#���P9���4%�9u�C�ɦpo�D�V(�&�����I1:�B�I0v9�i�V�?7��4���	�mO�B�	\u�%�%��>Mv����>L�C�	������h10L���ǂc�C�	�p��؈��	�ӃEPۤC�	T,�]�Q&$W��%���Q��C䉱Rm�Qb`�
1���2��+.�C�	�*4c�Y6�����!�>*�B�I��\��݊1��̘'��_޲B�Io+|1�a��b�̬P�c� -ԂB�	%��Ш&OBF{�D:�a�I�PC�	�jP�#V�X��$�ӏXwKtB䉅.����n�#��qP��*�B�I/i�u8!�]Tȸ@�cۮ0V�C�	 v��`s��<"+�]�sFU-w�C�ɴ���S��4�pm�Ӭ	dC�	 ��ʀ�׸G�^�b3.N�OA�C�I9ĆT��#�R����}n�C�	�n�(��Uj5�\Ej��W�g� B䉀<7�zU&W�GO���K�Q["B�	�<!>��#��84�eP�d�4B�I0�dE,�!l�t�i��7��B䉳)S&��D�G ~��0*�>)�B�I?g�:������5Bqx�g_�ٲB�I�#�rhkq/&n��JBn�'m�\C�ɑ�B�a�X8M����ca��"�(C�	i��	82c�K����F�+�C䉜��u�Q�	�b ���䇓��C�	�|OZ[!%�=�$�ۦL��}��C��6��	��.�;*�w�0>N�C�	!VY�����GG>���M7(��B䉊<>6�@��O���m�� �:2�$B�,j�j�R��F�D�hj䌷?\��D�.6j� (�OB�N4� dE�aW!�d�G��颖&ģ��[��]�!�]/DS��ȖLL��Fс`ˡHw!�D�5,7�QVL����@����!�֐y�PH`C�H�`�\�A��k�!�e+�<*�p��L*5��@�!���8`-��/F��쵙�#1!�$Y�m/�h�W�'�n� �Q��!��� CU�d0vQ�)��A7M�j�!򤑻h��5� �;+?V	��@;y�!�Ԏ.�@�ŋD�f�J��
j!�d״l8!��*���"q�Nz!�$��tB�y'@� �Y�~!�� �x�@4it$\Z���C��P��"O�uce�T;iN�9s�eյ ��'"O��82#�	K�~t���P�)�"Ot���ŭ���c���L�
�"O���aB�W�	aw5�]*2"O�u1���I�d��4 �7�ڌZ"O�l�fOG� Y�1��A�
?Ѳ��p"O�d��j�;n�)s)�(q��K�"O@�#�W�Q����^>�b=;`"O���tę'ir�es�:0�>-��"O
��ѫ�&s��8�G�[�´S"O.��̛$c(u�"E+3�`5`�"Oް�%��E��J��P.�7"Oܤ"7@.2�"9 ��/C��7"O�L�wΜ:�ٹ�d@.g0���5"O�D ��S�[g���wC�%A)l�; "O�T�&MX��Q7�J�EL��"O����$�1m�+*$&1�\QG�~�<�bK�+��P�5eU=?�1��t�<1$"U��zs���J`��PC�k�<Q�'�	3zB� "��1'B][��3D�� �O��������J=�G0D���7h�$j����(�O�<5���/D�X��`3./�	��&I�/�)�r@ D����U�me����X�frrx+a�>D�4�g�ڿptdI1Mݩ"n���+?D�t[U�&w88�P�[�R�r��/D���wB�+W=*��H̽7Ur��9D�L��ގt�ŉ�
�&�`���1D�@��K�j�@����?ht���("D��9��F�1�p��&�=�|��n.D��X��`b>dI����b=����(D���&�8IF��g	�t��ru +D�8��"��b�"���-���1�)D�@1e�h�����M�8��F�3D�l�&�U~�b-k����dճ��.D�lC�IE��xT��![bO�)SA�(D�<�!)� =|DH!�d�!O�ƅ�bb=D�D�S��&Hb�9jқ{�B$[��:D�jW͞�H�T��`�R�d���t%2D��𒁒#W16����kT��E�4D��$`��e�#ច3�$�À$D�����m��A�I�m�� �"D��[5�� =/��c��ض[/���I%D� SM�C���PQD�6'�p�r-D��K$I�j[��.1�&�(C��
4C!����d ��e��~j��
�Iܫ)C!�ٻNO�ԩUoځE�X��t)!���9­�V#�(��9�m��7!���>O (��ц]�Bz�C��׏=`!�
,���p���bǄ���I&@r!���w�P�o�q�2�1�@�#_!���6\��+�3I��@���&J!�$�f�X�P�`���S�hJ!�đ2,`J����BM�ZXB�g�!T!��
��H-Q"��bؔ�БE�*4.!�J�`��$��l�3�N�)���Y!򄁽o�&�+�H�H���@��#c�!򄒳4S�$����q�*l�UfR$ j!��fu:E�D*`���f#��E�!���Y�%L�\�D;�b��_�!��1a�F�R� Q���J�O�A�!�A�lr���4`TBw�*�gM`!�DM(�4��ūN	h�3\!�� ����G)?B5�F���+��#"O �cgV��м�p��j��\��"O��@G�@�@A�o]M��r"Oƴ��Ũ]�"Xh���<-'�yav"O�qA�W	F�0:%��	Q&ò"O�� �Ŗ1h��iku/������"Ox�� �_� p����� E���F"O"Q��i1��<��J(c�&d0�"O�E�W��8��/+�8ˆ"Op��S�E��:'�pJq
F"O��`�aA"F�����jZ Y}D��"O��0Ğ}�� b0�FO����"O%��L�6X�ʩx�ㄇ2��,	C"O��:'�?�h��њq���`�"ORq�QF������Sȃ�N�"�w"O��1�mΑP��)P�� >h���"O��s� �`�����E��"O8L���;%�b�Y�%ހ���"O�������$I��E��}�2��"O�, p'
]��R��	1�ڭ�"O��*�,C��$#m�025"Ot�vf�����,�)�$-�`"O�|���+i<��jły�"@G"Oh��#��<�%[B(�1:��}��"O���v)ȓ )lQ �gB4,xz!6"O�@�`@ΑD%�6Ǘ+�x��"OR�[���h�p)�E�90�0�{D"O��$&�o3&@  � =L��"Ov�I���W��E)�OKN��9P"Op�����:2B��"�]�;���u"OlZu�^�P�}��X/*I�"O4pA3���(Ы��d�=�U"O����D��r�n$H��A ���i"O�����Q�`��S��t��"O��c%S�p@�3�	Z�vy��"O�m�-�m��Qg��;	q@"OT�P��7��U�2��k�̐�$"O�v�ۑ]d���gԸ\4��U"O��!�أ!�T0�E��]����"OP�䙈uP��# �� ;=�U�w"O�5Q荙�^��Ղ^9Z;��Ң"O~�4 �,,�L�I��2"Oxiu��=~3|�cΞ0;� �"O��)��^
������ >"e.��"OL piУ��<` �O
"B����"O��+7+�F�<���͒�pNBE��"O����x��,��J�1)��0�"O&�Aa�)�����J̻L�h1"O�M�w��:X`��d��<6|��"O�s҄�:5 �B�.4�䱘�"O"M���#��yc��O�f( "O�$s��@>T�0Z�c4[���Bw"O��Y�`�,-8�`b�-h�^}�"O8��8=��ᢌ�_[rMB%"O�P��`��*'�%� �ǉOM&��"O���&����EۚV:Q��"O��##F�U����aM�;�rq@�"Ot(���sL���<��-��"O�}r�����`���&��%YU"ON�[��cD$#Vb��Da0h��"O���5�ʁ$�)��B��C�����"O���RI�hXN1!A�ҫ	�
3"O E��E�S������g'�,�P"O��(6���7�ʔ���R� `���"O� ���Bس1݆���Օt�,���"Or��E��5��%��Ż�"O������(A�gjI�O�P��"O>�"����cƊ2$4��"O �J�V�wU�H�.� �Ț�"OZ4���R&��f��O�#�"O(�� ��A*B��� p8t�r"ON�ё�0T�,�R�Y�d����"O"Aᢍ��U�V1 wI�n��G"Oz�����H4��!�h��Vi~!�"O�0�@WK���S��(ED7"O~���4rw�-âM��H@j�b"O�@8�	��H��͘�/��Ka"O�i��E� �e�wPD x�"Oрb��/����J&j`SA"O��'��(Y��X �G�T\���V"O.�0�Q7��h�	�15���"O��b�.�L@8�C#>&���"OfԠ�*��IJ,� fE&0b�yg"O<tk3��>4��"#	h԰ې"O�P�$���-�@jf-�}>�s"O�4�+��R����A-^;���"O�41��s���ɀ���_&8P�F"O41��wG�p�c
`����"O,��Ƥ�Ada9ǣ�) 
th�S"O���c�Ae \("!ĺ\��"O�q�ă�4�ԢU���b�,%2�"O4���h`�MK�l�:��A.�yr���i8�o�[��A����y��3rq�S�	��M�`!T�_��y�iT�{�x���i��K4.C��y�,�2w��87TX��r��ȶ�y��qx�cVp�"c
��y�gS/wі�Hi�Kc֙3vG�yB�RD<t(��ډi���⩌7�yB�:5<�<ѷΌ�{r|ݢ/ϱ�y�,�v!�p�AE�ioP���$�y�����߉\���s�+�jfh��`����J��f   �?ɸy�ȓ{�~���l���Z��剓!���ȓ~Z���F�)DԶq{�_	[��ȓ-�Ό��ҴEt5�'@W�Y�ȓk*�8a&B�3�����D�{V4��jz��giַͶ�p�An�A�ȓW?^�:֦T)w�����6B{N\�ȓ2�t�@�Ț6|؂2��j%zL�ȓC�H)��k[/��K)8�)�� W��@�G�z��J�
� mȅ��*���tb
$[���
�.e�a�ȓEH��k4� �\:uO֍H��i�ȓl�d�Rj )zp�2h2[�Q�ȓ�.���l� xN$Uy��� �V0�ȓ?�A fb�	8���b�@_F̇ȓ�J���	lB��3c^�}r	��
�H����Rt���FG5(A�����E����%VR�s�E1���ȓ��q�S�II�ʁ��i�)=����{�hs��P&V`�˃�B�PX�U�ȓ���Tk�:b���Q�A�x��ȓ P���"���F�1۶��`F����IR�|Y�����r㩁�x�bІȓ \�(���Ӡ�~"u(�%l��m�ȓ+IT\J�#Ȧ|�9�aS�<V���ȓ3����j�8&���!bm��cm�P��S�? D�&h�&���� �Y/T�w"O�0���D�@1�4`�#7*i��"O䀲jG���@bo�2��s"OL��Ba�,{:ܡ5Ė�~>�I�s"O�L񦣛�^���9�39>��W"O����3(D,$ Kӧ%z��v"O���Y�VP5�ʬY��Z`"O�]�rn�Iۀ�����$
��f"O���1�ݢ"S���,N(t+d͊�"O�ų ��)��T�����`*x�4"O�CIM��V4��#*Dv9��"O��Ibo�)X�tZ#�·a>���"ODP��LH�h� L#�ɋ�S�Z��"O tإ
�
m����Ǉ2u$;�"O脐��=LԹ�ɢ'���B�"O������,Ȧ��
�*g���K�"O��	'i&mVu�D	���5ӆ"ODXJ�+����;�fЦG�4 �"Ohp����Ӡ��e��o�\��"O�u�3�\�*أ���z]��
&"OqQ �,. u���I�P)
"O���Ԩ�6}>9�sϑM��-�"O��(��Ru~��CD�<�I�"O���R��l?��+#�/9�jܘ!"O�� b� v�,�©��eٌ�@g"OfE��'%���au��� Ƙx:�"O4����p�
&]�q@ ��"O��S4oZ*=�|U�f�-RƌK�"OHd�g�]DN�
B<7\Q�"Ob$!6c��^�@4��Z� `���"O��R4B��Q&��֤	�}�t"O$p`#hE�R����mH��6+ "Of��P�&| �O�62x�Z�"O ��^_���`��<Z�L��"O,�ڥ�W<�2���%U��3"O���s���>��#lZ�i�"O���ӤL	��+P��-V����"O�sP-ԊG	։q����O�<P(�"O0�+�N�lF�(���1v�b-)�"O qr��/?����Eй�b`�"O���20gK����R&mn�I1�/��<F�''
8��D�2H1��@BDY<��3�'X�8�@�U��ē!H%,����'��-� m7Ux�+!	� <D��'p0�*
�c�*Q��=�jI>��ν��<�}��m\>@}�rG���]�~hqr��Gyb�]�v�t)�y��)]�d���B+�:���μf��ɷ>l����.�)�,vZ�"֋ .R��AeN�X2��r�Ũb�
�*��T��)��� ��)p�m�qv#C�lRl��q�Ȕ8���6Q�<���v*���Z�"�0���IE������#<ب�"b+���`YdoX<[�<ʓ�Oc~�������mV2R��m�&�Ǹa�R$���Ͻm�d!+����0|b�I
�k�Me�N�uv��:ZR|��4%5����q��;{H-"����~�K|�uJY�P��Ͳn4}�X�֎˕Z���U,����S��M�;j6�Pt	^�1َ�I��٩t=�$i�F3�	�0|2�K�MlY�׎]{f�J�B�Q��P�X�J|j%N��l3�Da�м��D�P��	2ê��?�~��f�,1�U(���:^�2H��TV�<9��=A7��hS����H�{P�BR�<��,ܭl���3%�}�!�Wn�r�<�.ՓO|���&B[n<HU��n�<�r`��	u�0+ �Z�~�v��C��l�<��Q/b��
3鄷#z��3���e�'~ay�*�Hx<��MՋeB������y�F7&,� ��'����FL5�y
� ����$�T=k�iV�y��Mb�"O��1C��7( ���0(���"O	��"�9:��]��m�6$�	�@"ON�)�'6���(�i�'n��0�v"Öq��^z�l�	H�<@����d"ONm���ߓ{��q,J�|d�Q�"O�� �,�#`FH��̗vY�b�"O���S�ƞDj~��ɍ-s<���"O���c���	������y0�Ub"O�TI��U)1XP��9x�@1"Oȸz�Y(�2��)��5Be"O�]b.mjn0ڳmL�0K�H�"ON�
ce�@z2�C��,T/ܬ2�"O� P�'G�8�4"xJ,{"O2y��s/��Jo��&���'"O �q��N>P��MC�" ����"O�Pk��%���P��e��H7"OL�0�(]��9R����E��"O �҉ZU�����
�%
�}��"O
��AEߤ>����
-M�|"OD@��gӼp�¬��J4z��bF"O,��6 ��t|�أ���Hx9K""OB�@��}�^Q8j4��B"O�Lk2���\�s0g],+`P�{�"OV8�քS� ��P��8PL�(�"O�UYUb��U~Ri��'���Q�"O�)P�Z
7�P�M:l͞�8�"ON%q@�"/��J5�>�A)�"O����hM�C��XX����_Fl
�"O�1C�]�S	b�c��B#��K$"O<܉6�B cr@A CdB%�
m�e"O��؂Kώ�6l�K���|5"O�q����_p�(�2a_����36"O:0�5䉻i;>�ɤ"')���q�"OpK���8�D����GQ��yТ"OȐJU B��I`#��|T�"OtL�� ߏt9Z9I�O�D}A�"OL�ySG�&8���q��|�䲄"O�<X$N��]�t�igʀ�{�L���"O�$Y �ØR#`I ʙ�;~x])�"O�5���-�� !B�%>�I��"O��� >:���Q�m�|�uzF"O"�x3,c�P3ƥT��;f"O([�DU�@NA��g��\����"OP�C���<ʄ���L>@m�Ts!"O�qY"�ߕ#"V��ܼP\��`"O����+ S�TpWʝ9.바��"OhE �+ѦZW��(P|�*h�R"O��eRP�=��7�hI!�"O cC��%#�B���eڼ5�����"O,�(�=G��� ���L�(@H�"O�$�2d�h�4dw�r{̅:�"O�x��O�t]�
��* ��y��_=�89QʔS�ڐ� ��yB�K<F ��ʧ*�2OKZ��rͲ�y�m2Yih#)� I��9b`ݶ�y�J<��0�:qb��a�@��y	��k�0��a��,`���Ja���y2F~�F�p���S��AY`�վ�yr�L��� d��a1��q�ӽ�yˢ&u�����C/`�P$� $E��yR�Tbj�!��T0ڄ��,�$�yҭ�P�Y��c�%QP���s�O��y���=8��;��	�8BY0�}�<� <���׊q������JFp4�c"O�,���ŷs�ވ�����3.�5ap*O���e�9Ea�
��\`�'"�����&M���ˌE�@�C�'� ��!Q<r�� Hg��9.m+
�'�p�����7�^�&�?*ݖ`Y�'��=����-ub�	�#�z�����'m�Y��A�k���E��xO-��'8�$qJ���t�vl�4_bΩY�'�J�0�Ł��aBG�W��m`�'dp��FK��Q���H�>�E�'  4����>��Y��(:,\���'�z)1�cȧ��*UJޡ!/Li��'�E�'�§j���HD�^�J2Ʃ��'�fٹS	��,�æ�xa��{�'I�m�u��6����E�o�p+�'\X�7ɇ�ow�9*���`��AS�'�h�K��4���F�A_�d���'rh��.��x���LC%V}8��'�8� �Kګ��!P��G�M����'�REHq �/4P��gX�L��L
�'rn�`oV�ܳ@��H��
�'���b7�ٹ#U�g L�9�|��	�'6���KBt|}p��2��	�
�'�8m�sKB(���4�69N�z�'����1�E�MRp���3�(9�'��d�V��M���E;�}�	�'�N}��
�l^�Y�GL+ Q�t��'�.y��G61u���	�1u��1�'�`P!�R�l�L� �o��k����'i�h��ɍ,�~3�/ݖa�@��'�ny�E�H5*�@fk�l�����'�B�y���5b�K6�ːz���;	�'K��q�jNx����]G��q��'O>!B�l
�M����"��<��`2�'W|���/����5�ʑ4	�(�
�'h<|q&¥@�� Vk�#�f��'�J4��Ǉ*_��3���*`��'tlQ U��-��Lha�1�N�2�'ld�I `ԫ\��S�iY�_�����'� m#d�݊�b��g�5H�p���'W�|��$Ō`]n���I���'S���ǧ ��cM:q� :�'ʦ�qn�3Tea@��
0��)"�'�n=+uL�;#/��bJ�$ݺ��
�'����qe
Or�0���L���ȓS�<��`D�/t�1t��C�Z��ȓK����&\ ���Q�@e�x��X\I:+��s���AQC�=����K�>���C^~x�ۂ蜝}Kꠇ�[C*Sh�� ��X� �K��x�ȓ9O�IRp�2qV�%{�A� 40��L(Jxg��j~lx;eNb;�y��y�0�t�%�P�kE�F�|���ȓm;D���>8�r5�1�O15Be�ȓ��<��bD�o�^�SP�4~.�Y��eH����X �Qs3�-� ��M�r�-�I���� �*�z��$���a�郯9����XBT�A��5�n�EE�'*XD�@'�3������f0I��2/"Y��/Gmp���'G�<Hb�͘^^3#��1I$ʕ�����2�X��X��$��1E��I�ȓS�ư+2a�� ��oC���S�? u�A�ħ+� KO�_j�Z"O�IYB�ߢl<��Dt��tY�"O8�	3�¹h��z�.�.9��]b3"Oz �6A�H]�b�,�ɒ�"O�ظ�n��,ش��Eg��V^�"O����`�3�p�2�(�Vيc"O2H�S`�a��f�LP��e"O�	���e
�� �+�%b��d(!�$��&�Dd���~�:��T�U�R%!�.Ex���֎�'�,���2!�
.u (�#�>R��`P��I2ko!�ބW��\�AѠ��}0��֎!��D�~	,4�������r����P�!�ߓ�n����$u�3��ي?�!�w��Mp����>�* ��� (�!�D�	\w��@f'�=�X�� �!���,�t�B�'�ܽv
�h�!��E:�ج[V�g�M�T�R4�!��T!8��m�r��m��U�7�E�g�!�׉�DI�]�}��(6��Q�!�$�Ixy���t�Z�j�1F�!�%\�f�a�Q�y׊z��L5t�!�DU�0�t�QT��7<]����A$�!�D�H����Лf2̲Sל"�!�d��^�4�6EIv0�7ki*!�$1I"�A�F8F�Ī"-��8!�d��&tv��WgM/E��Ȧ�Py�ءa?�)�M��'&y*d�ڮ�yrf�
���DF�l8�֒�y�B[9viM����H�r��:�y���r�ة8B��6QE�k�E�y������Іޡ2� ��� �yR(�)o�UH���h��@���y�i�-@�(
�*	�j���3C�y�����҃��2��pi ��,�y��K6y�(!t1>�'	���y"V�8|	�S�� �@�뀍�y�<8;�q�Dqm;&��d�!�ߜR�~ٲ���%M�*�'@'�!��5G3^E�G�%�n  �hB�	�!�$֘�ȡ��d��B��mI�Y�!�dJ�!.4��+�?��(;u��SX!���Q��
0��+�����;F!�D�yw�E��̊�yl��H��!�P3slZ��«V -s�e�JJ;S�!�$�:��CS�N�ȤٳC��>�!��:wݎ�*����_HU���sx!򄄯{�����^'BR��%��Qj!�<L�
�+�n)G�(�k��p�!�d�*0GB�{��O�cj�P���6QO!�\�=�6d�C�r�"Q��aV8R�!���X�. �e���X�r�A�&�5!�$�O;^�s�m 5S���9���!�D��2HB��A�_M��; n32!��˰EK�T��ϫ.� �I�ķ	!򄊵I�D�C,�	��b!����!�DL�6���W#��*`��F�U�!�^&V��*�
��]�U` �.L�!�ҏf�fDcK�lYfx�n F!�DA#��%�V@��x��V!��X)
�jIJ'g��?0d�F+��!�䎙�]�CkW�	&h������!�J�+��h��_v��*��E�XV!�DB� ���^)2
_(��"O� �Q�N�r�% C>��`@�"O�t�Ώ{'R]�ph�FHXe��"O�t�$���u���Y���}�"O���A��	g~a�Qχ�"��@
�"O�}`��g�mIԤ�.b�e9�"O�qC#�5�]�2ꆾ�M��8D�|2�
   ��   �  ?  �  r  �)  �4  @  �J  V  �a  �l  �w  ��  0�  a�    �  U�  ��  �  *�  ��  ��  D�  ��  �  ��  �  c�  ��  ��  =�  � � ; - C% �, 4  > F �L �R Y [  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+��6-\�c
�<4�d5h��'�B�'���'	�'/�'�B�'���k'�M�=��Y�A�D�S��܃��'���'�b�'���'�"�'�b�'�t�"���#H( �TQ)G��ڟ���ğl�Iԟ��I˟d���x�	؟�QH��&
ga%@B�Z��[�$���<�I�	ӟD���������5i /;N`��M`�
$��J��	���	�������ß���4��$04��)�¢�6���N��|��埬��������p��ٟ�����D{ ��n��0��/�'j��: *]�l�I̟����8��ן��I꟔����T9���Y�`��DI ªK���韴��ퟨ����	ڟ���ٟ$�I럌aF��sk��C�cV��p��ɟ��I����I����I��(�����I˟�������H���-�^�rA��Ɵ���ɟ����p�Iٟ��I蟀�Iğ�yD� XCbE#!�0�� �����Iϟ��	͟�	�������������Ɍ|��Q�C�%����A��)n ���	؟�Iʟ��	�����㟐�	������Pӧᑘ �􁣃�ȴ1������|���X�	����	��|�۴�?���4_J�2���7[��R�Z"Y�VH��U�h�	Qy���O�Tn�9g*�Qq4��d@9�L��|�X|{��>?Q����'N���ĳe�����(P����m$es�KB���	
E���m�f~�7�R1�[�iR�5j�P�1a�	/^�\y�h�Z1O��D�<Q��IL ;�S��NA��@ס�$G���lړ��c�����Ӽ���:�⡛�.A�mS~��b���?A��yU�b>A���֦��QDp���I��>*��a`F�\����y��Od����4�F���lg�C� �~e��]�h:�ı<�M>��iR� q�y�;s�[�8>'�M[���=X�O0ʓ�?���y�Z�$�A��;!2���P��HQ��,?!�r�h���.�[�'r�j���?�a��(��A^-s��}`#���D�<i�S��y"�l�$���'��M�v,�@d́�y�Kdӈ�;������n��|2t�>s=���K��	xp��<���?� R	ܴ���q>�1��Ct`���OZ�%@� YV�;�9@%&���<�'�?)��?���?�s��'���I"*��#dP�����ď�}�qy��'C�p�9���A D�+�v�0�S���<a������O��{�ڢR��Y���Jbe@�@#I�9b�U�8��� h����D��Ay2��Sr�� �-�hI����'��'��O�	&�MQh�?�?ٴ/�#��!��"+�`�O=�?q���'J�۟���䟐K��^?��L��&�5����1m[9.Z�o�Y~Bǹm�P���p�'�#Pc�Rr|0��S%�!�s��<���?)���?9���?)��T���p�'�J.%�t|QQbʷ��A�����I�M�$@Pv���'h�'>�r#��W`}��$YT���|�'9�O�a`ӵi�I�O��ĩ�%�N0�7-�3O���Ecj���8���<!���?���?���۷,���Y��K:^sv�Y��?q���$��]��ӟ8����O�Q�u�� z�eD5!恙�O�˓�?�����S��#�*/�f��R�ֈny��r��D� <���B�J�*nn���O�i��?A/�DG�i���HW�:�6��1��)DH���OL�D�O4��ɰ<i��i;�5��iڂg�&X
�A�P���!�܇���ݟ��?�(O���|�&9P��B��$<Bꂣ��Dz T�ش��D�^�8l��'"���Z;�U�1��m��"��"*�0����O����O4�D�O����|��F�$$bx��c���a(Ǐ�d_�,Ęqv��'�ҟ���'��w<��EdO�T�(�sˋ��,�R��'��|�������6<O<B��#c�����8r�p�;O�=�1�?�?qW?���<�'�?�`�F�J��T�ǂ2Q�0����?���?I����ɦ��F�ʟ���ן��� D$ND��	�$Rz��))a.�K���$�O���!��]	V�@󡂛J�h��*I�x��	7�� �ӑ$��c>1�@�'������hWHĳ��Ռi��@� 	нP��x���,��ǟ<�Iz�O����e� 1Bbh�1��D���v���2 f�O
�D�O���]/,5�@���ue�$*�i��hb�I�������˒ܦ}�'�
x��� [�W��o���WC�� )��'�'�䓢���O����O��d�O.�$"IblSf�־\\��g#^r8�A˛F��6>o��'����'4��sq�E&�@��D�%I�| U�P�	���&�b>�ّ�Mq �b�I�V%l�����O��d���~yR�)M8��	���'O�ɴ�P���ջ*�5I�/��1���	ٟ4��ן �i>	�'h�7"yG��DN-s�Lѕ�ňM�X�K�������OV�`�'���'{B'	�E��AcH�6^��-��ʂ n��B�ia�	�*%�Ar����� �H��P�h��k�$/lT�(�8O��D�O����O��d�O�?=q�JfLq����"���b����������42_(y�'�?�����dV ��:"��YU��I��5�<Y����)ͬ6m.?Ifń JO�-P��$ԺA��6&x�Ԥ�OrP	H>�,O �d�O����Op�9�JԻ^�� ���-��0#�C�Or��<�ÿiZ@`a��'q��'K�S����2�_w��u2f�܉M�����O��d9��?MQ�U�v�7$�l�=	Pm��X�(�}I���|
A�O�@�J>颠�rT������-&����4����?����?q��?�|�*O��lڌ?i衡ՍG-6jQh�+~�ڳ�۟���ޟl�?�(O&�Đض�b&�B�N4�i⭚5�Lʓ}b�qܴ��D�)}�>���'$�:˓n���D&�&�~4Q�CL3$��%���d�O6��O��$�Op���|ڔD�X*L�#�^�,��,+�$VY���	��'�����'��w�B���ӣP�����>LD���3�'
��|��D��RQ�7OF��U���1�~�%!�P�X��a5O
��Ά��?Y��%��<�'�?�ǂ�'�:��Y�As��!�j+�?9���?Q���
�u�������	��P��
A�a��c��U}��ӡ�TD���$�O��D,�d��<a���T��1z������ɷcf���R�Ǧ��O~��%������z�6}��N�iq��Q��PF&����d�	�����_�Ob"��-vl�u㢨�2%��]��b;���Ӕx��d�OX���O�����!���`jH�9R%E0o��	ҟ��I؟�R��æ��'`��I�!��?�C"-�40�'��-5�HtZ nZ�H0�'��i>-�I�������P��2�%)�� �w�<�Q�D(@[L�'[R6��q'J��O��-��3p�>� D�ˆ^�t}���P�c($��'���'�ɧ�OZ�|�P�'͖Iڢ荸U��yt�'p�0y0RX��rG�	-�B�s��Hy2"�>j��J�%J�t<s��D10�'�'D�OZ�)�McFS�?�Ԅ��k�s�nJ�n:v%It,���?����'��Iߟ���䟔xQ�&'+&�l�p�j�Ȟlx���i��"{>8�p�O-q�B�.Cn�䨳"$���ِ�W?!�d�O����OD���O���;�S�������l%R#KO�c���ϟt��.�M+�	�|���?�M>�@��w��4�b�&:�x��C뙶���?���|��	��M��O���=D�J['K{=�n4z�^�Zc��O�u�N>y+O���O��D�O"@��U~Fx��#2���P��Of�$�<I��iR<@q�'��'�������D�9c��Y��F]�Hc���$�O�%��?E��o��,�!�c�z����o�H����M5�1����KSʟ�V�|2�J�.��S�M�`&���a�n�b�'�B�'_��4Q��;ݴ9X�rR���;��עޯ%%���e� ���O���'������hx�Ä6M�Q�E@"p~�	�vlPl�m~���g4H|�S�_�I�X��qUBQ;aZ*�顥K�G���	[y��'.�'{��'x��?�@EĎW޵�P���xU�0��m�Ħ�p�����p��ܟ�%?�Iǟ杜=��`�JN�e�T x�L�2k����l�Ş����ش�y"NS.-�N�"� �a���M˵�y��T&"�d�Ɉ ��'����I
6>\aX5(�f���IG��8UTJ��I�����ٟЗ'267m	�a�����Of�DS1�Ե3C߯N��y(�(1� �4�'J��'��'�l�J$MB�2� ��AI�;�����Odp��µY\��	O>�i@5�?Yo�Oz  5�O3<+� "D�D�؅��Oh�$�OR���O�}���j�tP�>w�p�P2@��"�����]ћfl	H�I���?�;,\LH8�R� }��L�?��	ϓ�?!���?��@��M��Or$�cM��b!�A�3<�]Zb�Wd�I5' H��Ob��|
���?I���?��Z���BMڄX����g�S␸
(OWc���I�E�O���Of���D��0d��\3
��l�$^�];�ʓ�?a���DȖ^�8�"&	�0�r0I3���D�2���-*� z\=��'N��%�,�'^8p�&�"Y�����* 6\S��'I��'�R���W�p�ߴ ���Q:ೡ�V(Z_�Y��
�0q� i���?���S�P�	�<�	�Fr�ZL�1�,iX��˓P���1��ᦥ�'MBQs���?�Ӕ���w� �AW�~8�B��٘)���'��'/��'>��'K����W4;�P�!0��T7����Ox���O��n�b|�'��|�e��ژȂ�1�TAӰ�N]�',����Ԋҁ):����lY ��9Rh���OݰT�d�F@5Is�+��'��	'�̗����'�B�'6NLbU��0�� H�u�h�3�'b�^� �ڴc��
��?���M�m|���s(����CE<@�	Ky��'���|ʟdt�f��H\����u8���eaF�s��h�f��_��i>!ل�'��%��d�� F�MZr �o��\��o�����	���	˟b>�'�N7Mٮg�H�12�5uZ����GçW�@16��OL�D�O&���'&b�[<)�F��� 	f�M����'vR�'4�� #�i~�	�^4Hr�� T|�f�C�d�$Љa�C�	h����;O<ʓ�?	��?a��?i����)M:B�R|�d�Q<w|��!D�,��doZ�|��8�',2���O��4�.4I��ϟ5z�p�'G=^�����O��O1�r��c�
��(��;׌ ��B���V��	�s��0�'A�D'����d�'͠�Vh1��P1(�(� �Q��'���'��Z��ٴTJ�����?��|��h�g�Z�k�[�'Ӛ*�ؐ��W�������%��Q��ͮ��lZT'�/J�r���j8?ɴ�E,&�ViQā�2��,�X�ĕ��?1�L\�TKH�K�NJ�bUh��#c�	�?����?���?��)�OD�	��@<D0tP���`#���Oho�:H��'F�4�lP��e�����Y�E� �D僇2O&���OR��	�-s"6-*?Y�)�0[���IG�-é�.GԚX����(t��dxL>�/O�i�OT���O����OT�Td��X�Ҽq��E�'��a"��<��i����T�'��'l�O2�-j���K4D�{�����D������t��S�)��yL{�Ī�D��q��Z��������/O�
�� �~��|�_�S�i6G��)z�kY&y��|�������I�(�	ϟ�Ssy�Kxӈ���O:)�B	"'縥K��X,�P q��O��:��Xyb�'r�'7 )�߈;t"�@\�[�����J�K��旟��v��@@Q>��]7C�j(��̠	HT١w��;e����X��ӟH�I��x��n�'>�>aE.;OlQ��ş�Ql����?��k��nK���t�'\2�|��)1���(�Fl��Ѧ�E�S�'������D
�F��F���
)6��+�l@=g��5c�۟oظ-)0B
���sv�|"R����ߟ$��Ɵ�Z �^m��[��K:
+�h3h]�����ly�nj�R��R��Oh���O��'1����W_�ja��l�jJV��'��	՟���q�)�A��V�q�L���I{����$�#6{�P���4MD˟�XA�|�-��3����gJH�0�x��@�8`�"�'���' ��tV����4TĤEp�@�'�J�C�mb��}�����O���'X�@��Y	��p�nI��KH���z��=o�V~���`7�T�ӵ)��I�E"��iQ�	�so���cj��#$�IXy��'d��'{B�'q"U>�Z�(����Z��V7�\�C�A��Mce���?����?�M~���?ͻE.lD�c����rb�Z�Y��?QI>�|�0���M{�'n�	x�LG�s)X��ő �(�(�'�t�8W��A?�L>1)O�	�O@}�rΛ�#���EɈ1N�*a����O��$�O���<9�iY�V�P�ɼ[���%͕�5�Ѻ��-Jo���?�.O���.��*�4XhslC�p���C%쉋eĴ�
�<qe� ˂M�I~2EA�O�M��}��h���H�/v<��G	P�EA��?i���?���h���d�}J��iW?=� ;KӎlPP�d�æ��0���`���H�?ͻ�H�NTv|lՍE�G_j�ϓ�?A���?��`
 �MC�OTuP �����R�Q:lyKW��4>lBW��+l��'�i>��	؟�	ğ��I/p������
�`B�%�δ�'�f6�PC�d�D�O��$=�	�O,�Q#�9O`J�&�
�"��E�<�������O�24�oʛo'̡�fO��_
�)x"\ʦ���V�, ��#1��ƚI�byr����0��K�[ʾ)s�R�b�'���'d�O�剺�M#�KH)�?�B��Cd���ı#it�{3bC�<y���'�����I��0$�:K �]�����)37JQ,{�doZz~���8EY���䧂���Kn�e�B@��r��`��<���?����?����?A������ф���9�ǚ� C��'db�~�v��  �<a����a�$� (Li���ɹI��!0N>����?ͧ@���ش���7a��)E'�+spL�5��y� j���?�2''�d�<�'�?����?	��.W�Zl�	�8a���A�O��?�������e��@W��	ߟȔOC��	���mRlZ!��taȴ��O�ʓ�?����S�4'.�Ё��h́_��d ��/r2 ��,ʌd��4��O�I��?9`K0��ݡ؅JЅO;<P��[b��������O����O��I�<�v�i*��=1�:l@�F�):�J�peB%O$2�'���<1��hZ�A^��X��m�Ͳ,O�����b���exP�E�ҡ�,Oѻ��ك^��<��0�j5�G:O���?���?9��?������:5
�iV`UUˈ����g� `oZ?(���'���T�'��w�2�HT�#n�*Y��a9#n�[�'5�|�����[�&6O>8��H�9$�@|#3#]�&Ԃ�4OF�CP�7�~��|BS�l�I՟��� ��j3�Ta�lF��ba�ϟp�	ş��	Jy��|�$��OX���O�8��@�*��x��D	�6.�h � ��yyr�'��O�X�54ޅ���SY��� V���`�� ��-�Q��N����ܟ�i�iR?[q�$jņ�
N�Lx5��ɟ0�	��<��ПE��'�n�r���>)��� �-"lh�c�']\7-J�f���O>�$+�i��2�����c�̜]β	r�+m����˟��ɒ&� o�o~�g�l�^��g�? rPc�6L�Ў]�z���2@F ���<�'�?��?���?��eP�5L��ʶ㔺 ��ڶć����¦U;P�T�����ٟH'?牼3vЬ���������nӐ~�Y�'�B�'Gɧ�O�0�"nؤ-h�;C"ی@��Gچe�O�	�2���?��%���< F԰6��8���L����8�?��?���?�'��� ��!�e���TH��� �&���o�*��9��ş��IZ������O\���O��R�O�cb����5k�@=�FNR#E�6m-?�,�(�������'��s"@N&�`@#V�Z���1��<i���?!���?���?��D��R���{%bB-�lm�%M��')��p����F2�$���OܓOt�O_�Sf��C)�q��D�R�$�OJ�T,���ٴ��d���Q�����z%���F;IC�U�CF��?a��>�ĸ<����?����?�u�s<zs�Ѭ"�2D��]��?�����d��}r������	ҟx�O:(��V�O���GM�sq��O�˓�?���S�dJ�pr�P�O#pȔ�#ĝ	^�$�;����JX��S�/��(]r�I=��� ��!d��f��rv�����4�I�|�)�Sly"�g�H�8�@zjh�B�˂9����5W ���Of�d:��Uy��'z�%��K�g��u(�U�aС�'���=L���������Y(nq�,DPJG�m	W� �4�v=O�˓�?Q���?���?����	��vc�h�&Df&0)�EX6Ξ8lZ�i���I�<�	_��柘�i�	�2o�*]��Z�A?�H�1$���(�	o�)�=t�Em�<	c�;��$���s�\��F��<��U*KP�dȥ����D�Ob���VtC�Ǡ�r\��������O��$�O^�5���Ej��'z"T�x#���6a,R�2����
<W��O�˓�?�����$0��0�V=[�4X
�A�X~0��'�zѰ���%��f�H��~�' `4h�H��9TkQ�#x|2!�'b��'���'2�>��+v��9C��"zNX(V�H�,�֌�	?�Mp+���?����?ɏ�w��A���>pd�Q Ѫ�G�Vm[�'�B�'�d�@˛�����Q?U�����^�̸:��̊-��9q��M���&�,���d�'l2�'�b�'bDY�s��:S��	��>1�y�bR����4HfN�i��?Y��䧒?���$NaH|[�Z�fd����nҐ��d�OZ��#��)l�����DÞE#<��O��U�܀7��G��<w�D�A�':�l$�P�'lF9��Y\���@g�җj�r�zt�'OB�'2���$W��8ݴy}�9z��rxIwm\U�Ȅ��/v<zI@���?q�R^�d�	۟ �Ʉ?j:��T�g��!�Q�W�e.�������'��������?Q�}��;�@h�	�CL�	#)�1`�D��?����?����?����O��}Q�`YM����g�(W�l'�'	�'F7�ܙ#��˓�?aJ>�vG'V�@�����R�"�ݳ���?���|�4O��M��O��BӉ��h[��KQn\�y���U� .-(ܠ���ēO ��|z���?���|h��
T� �V4"��B҈�`��?�+Of�o� L6Y�	ݟ���`��,��hg���.�z���@4��D�<����?�L>�O��-I
>WAfؑRjF7���X�t��r%`�-��i>ݢ�'v��&�H2��%$=4�q�m�:�rL '������ȟ��Iɟb>�'�,7��|����X�E@��pCL
��	��Ρ<)���'���ş��`�P�r���q�A�<T�b�
�����,�I�1B��nN~Zw�ԍa��O�b�'��5�ׁ��	��#IP�
^69��'��䟬�I蟴��ҟ��IC��!�-��˗�$�n�/E3��A��i��§�'���'�O�"��y'�T�Z-�aF��xTy`cK�?"��'nɧ�O�Tp1�iv��)��\�P	�>!|��f��8e�D��z���h�j�O~��|��C�l��-��,��B�2-���B��?����?�+O:�oZ�
����	ݟ���9�&X�g��4k=x)s �I t��A�?)/O��d�O��OIj�MM�D�~��V�˵:�dsv���:e��f<��l�C�'�~����8�E)݌W *Pa���:K���������Iџp����8F���'+�ʆK�)$*D�N�>��r�'��6��G0����O���=�i�I��Ď*t(���� #V4@P��k�(�I��,��1��Tn�_~�Ȉ���;����V�U�2\�O�~�I��|_����T�����I�%k�~r,��HB�:��Q��fPKy��qӪu�f��OT���O����4A���M$#B(\�)V�<���?QM>�|Rf��4/�����8�:P� �)*�B��0*I~BA�1SD(���0��'@剫A[`� ��͍)( �H�j�;	�4��Iϟ���ݟ��i>��'A�7��~T�D�;r�6�X��Y�v!l�I��[���D�O��X�'v���y7C�n�>�*T�*���y��2N8K�i���86UȜ�V�O�
�'?���L�<� �J���0�Q��-~��͟��	ǟ��I��D��@��y��bP����rn
�aN����?��3כ6�ȎW��Iݟ�%��������\���NB	"h(1e�I�Iџ��i>�j!�ڦm�' l�j
� �ta�F�4�;r�֊R�N��H��?1�l3�d�<�'�?����?�2�K�rR��"��zSvtK!I(�?�����ă覡�#�_����	����O̤1s��}�*�9a�W�>Mt`�O`˓�?a����S�d�N1Z��]c�d��jic�`
384�T�G�hƘp�O�)̴�?a� 8��2�d�A�jJ-�rϥy|j�$�O&�d�O���	�<�ƵiI��	p��m�(�%����"�� ���'4"��<	��Z)h�yC�JB' aQ���z������?q狅�M3�O��AH%.������K:w B4��造0�Qq׹���<���?����?1���?�/����A%�
0#�\�У�:�ء��\�EXcAߟ�	џH'?�	˟�6_��E �"p\�=+��̝�h`�	��$&�b>awD�Φ�̓-|�X�KO	�d#���{~8�̓h:�H�����&�(�'��'�jhR��M h�H���m��9��'���'�S����4@�ɡ��?	��%` ��%�0�pg#�2�
�"R����j��\%Ѝ�6mG�]!8�����	�(�'�B�إc:t]�EX��D#^��PX��'MY����[v4�!��� *��C��'e2�'��'q�>-���1R�tSΆ�m�N���F�]t"��Ɋ�M��������OT��]�\e�e���Ed2	�GX�U`��Iޟt��џ`8�����uGBX�Tg����>H��P��"�A�0'U�J���&�X�'���'tb�'���'-~��K�5�`��S;��)Z�P���41�6�����?���䧄?�j�4 ��p�!E�_J)H�+����O��d9����\L�g��?y*���
�3W�MI�o��l�'�����LJs?�H>A.O2���ʒ>7wT(`�ȍ�@������O����OP�$�O�	�<� �i�bx���'�~}p�g�.m������K�w��#��'r���<���?ͻ@$R�����sa��x��
??\��M�&�M�Op����	�r��5������	�!A�Q����!���� �B8O��O<�D�OP���O��?�`�皗o�����PR�/� \����ן(���M[�/��|���?�K>��f<$<���l�� ��%µ���?���|�
T��M�O4�9���:O@=��L%Q��a�͗��M��?QȒO���|���?��"gZ�3PK�.-��9�h*<�����?I+O20l�F��Y��ڟ���J��A�-UHtk���Ժu;��M����<q��?J>�O��pqN�h=rM� �S�P8�x�,ߊ���i�i>E#��O&�O�9;�b�Pt^��C���ɡ�-�OJ�d�O
��O1�|�u��fCޱ&�``���й ��+��k�mc2Y����n�����O�%��I��+J-:��՚:�6�[�O���	!G��7�1?!�� �X�D��/�� ё[�a���拄>3�V�ʚ']���H�	џ���ʟ@��m��
έu�J���E�fvdɊZ����	h�b���!�O����OF������O��"\P*�Z�M	z���"�w�����OڒO1�(���	l�2�I�>)�`�C��&R�0���$�+���I�?��0*�OғO��?	�|��ȘF��'�H|�u��h�PX���?���?1/O��l�r6������ ���B�R����5Uq�(��2��5�?/O���*�	�Bb��!r�����_���B&\��w��:�Z��J~�W)�OP�o�i���s���3Ɛ
0$�D:
�'&$d
s�	�츇k��p�=��'I�6-��&�z��?��wy��)���9k�q��$o��)�'��'�c�=.�ƒ�L���#eB�	ӹ=�FlH��K#	Y6�r�'39��O>���O�):'^�i��miFo�,\�@9T���[۴��)S(O��9��9Y{����L�W�M8cJ�?�p	�'�2�'ɧ�OB�{��r�P��T�] ?�\���h,X�uiGY��sQ��hr�]w�	fy��� N����GT7��ř�մ�0>�t�i�BQ���'��]qP�G2y��c��	,z��',���<��?	�XsjI�σ�}TaIDϽ;��VhϠ�M��O�l�1�T��`o6����V���=1X2X��M�9 �*H �3OX��� (%x�g
�4��d+GVq8J��?a��i��P�ɟ���(�ćB��	I&@��k��@�v(��h)x�O�$�O�;^I�6�7?��&L��
 e�xh*�-����@P�.���%�0�'d�O����Ƈ�=�~�Ӆ�߄�h�j%�� �M; hԛ��d�Oz�'X�ZC��?�:��J/:/X��'a�	͟��IP�)����c@)�cd�������>���V��M�3T���,x��D!�dH�����á�1M=�U)w�ˎz(!��Nۦm(3BS�pu��#Ӆ�y��Đ���6d6�'�����<��" �D0�Y�9mn	
⊱#���+���?a�h��M{�O�R�3o`������J$NP�*�� 7z���Fks��d�<����?!���?����?�)�¨{��̕z����%�K8%�����ʊ����rn�yyR�'i�4�4���"am�{�b��]8�yp*�O��b>)� k�ᦥ�S�? �@C�˝+��1�H߱H��l�9O��	�H���?�d�%�$�<a���?q���X*�$�@�ՓRI^�ڇH��?���?q���Ʀ)
�ˉ⟤��՟<BD�n�z@i�D��n)��T �a�����O���[ K�Th6P�2��&�6!�sM#?��X�i�Gڄ��'k����?�VeQ�7$��g��S�r��D��?����?����?I��	�O|���'�� ,�	�-BQV�Ī�O�IoZ������h��w�Ӽ�PoT�[��!�&V�)�4�yE��<����$�)��6�6?�≕�R����T�&� 0%IU~8�B�G��Ѕ#H>Y.O
���O~��O���O���Q��2@_�%��Iي(C�3�̩<y��iN\��'I��'���y� ��^k��l�n�ՠP�ærh�I����?�|���[����h@�\5>~�ГWI�sP��蒸��'�*��N
ڟ<[��|�^�q'&C�o�l����va2C�D۟t��ӟ��I��sybgӺ��u�O
�%�+%���i�?�z$����O>�D8��^y2�'��	
05�1�uo�3'MM�4HқO��z��W�I�'n>��&B�?��d����w
��c`#Ȩv��x��$Ž6�)��'7r�'gb�'%�'��t�0c�C�pD�7���!m`���O����Of�mP-@<�'\��|r��?-�>t`͜�rdAcƩx��'Lb������Y�������J�0�D���.���Xj�(�'F�'������'s�'6`�a��_@b��)�4�)f�'#BW����4O�J���?������Vl-�W��
6MˁA1��IHy��'/r�|ʟ"	�d�ͽ*�`��nV'Y�6��cc��aF��{��|��i>k��'���&�`I��٦!1��b�᜽$�8u�4B�ß��I��@�	˟b>��'o26��x �	#�n�c�K�>ƼM�@"���I�� �?�-O��D�^|��˅OX&?t�E
4��P&��Ob�p�`p�4�=��᳆i��O�t��	�w� V�ܵD���'��	ɟT��ʟ<�����	^��o˫"y�PD�³m=��4M��%[۴L:��?�����O��w ��U@���$��c�B&8�Ȳ��'e��|����s��=OVH㗤�4������&+�X�R<O�MS��)�?�� �$�<ͧ�?1F�¶gf�8q刞%�z`P��,�?9���?�����զm��a�ƟP�����s.�/� �� � �5a�E�c�S����d�O �7�D�;�04��,0Q��H
U�ѩy,�	,`�>u%��S�Jb>]S�'�J��ɡ-(�911�E�q�x��O�RP��ܟh��ß��n�O����?RXa�^����A�L�* " c� ��&��O���O��]vo���-ӹf�R���gS�Q���ޟ��	�t1�k�ߦ��'�>9٤J�?���i��p���*�X���#+��3��'��i>��	��4�����I�2\�#���~�L���J�J�� �'��7M|T˓�?)N~J���8d���\f� �0�&7��*O���OؒO1��Mq#��+:=4i�Ч!a���y!��_6��tyrE�y:���䓁�L����P�ͦ��� ��,>A����OR�$�O �4�&�W_���� `���/|b��eh#%H�|�6��B�'��O���?��?yP�тK�^��U��7��l��Ci��-�ߴ��$��.56�X�O��O	ǍݒJ��]�Ɔ��^Eb�MI��y��'v�'���'����'�����B"�X�g�J�_h��$�O��$�٦��,m>��IƟL%�hLT�c~f��A�t�S��IA�IΟ�i>!������'��o@�C`�-����m��ȩ��ˠL�d�������O���O��çu�N�x�ºG������אJ8����O�ʓEs��T�j �	џ�O���$DU���uk�c��P��	�'I�Z�D���,%��'0�^L w��M�T��%!��\��
#��a��t�ߴ��i>A��Ot�O��#�����R?B�Kh�O(�d�O��d�O1�f˓?��f�C7O<��Tg/���/U9�F����'~b�'�ɧ�4W�X�	�w��+�.1_�h9�FE8I������`�ͦ��'�ʭ��a�)O�5�1�I|���3� ��=Ya<O�ʓ�?����?i��?�������5i2��AKɋH�L�H�Ir� �o�'�`=�'�����'��w��u��N�aٌ�J%e�_��U���'��|���M�mӛ�?O�L�p�ɣ\]D���@$K���S>O�<�ׅ�~B�|�Q���ڟ��ǎZ�J��MCn��q�ꬣF
�ٟ���� ��ky��t�\�3���O^�D�O�ӑ��_ �-�V�oc�9���,�d�Ov˓�?�����M*�p�W�ETpB���QMNE�'���d,�&̚��6��dm�韜¦�'��b&�N�ׄ�A$h�s<�[S�'�2�'�r�'T�>�]*=���؅)��~�a`� 2}����I��MSB/�2�?��?AH>I�Ӽ���a�E���~�����A�<��?���)��!�ٴ���S��H@)p�@1I�┊�i�c~��v�J�����O`���O��D�O���0���p��P0�]�Č�
Xʼ˓%^���f9�ӟ�%?U�I����B҈��/�>C�"�`��'�2�'�ɧ�O �1� n}PGD�tVZI���x��e�W�x��'F��z$|?I>�.Oh%�N�~�J�ʂ��F�i0���O.�d�O<���O�)�<Iq�i�J@q�'��I`�%0�Hm�J��r0j����'�ҟ|�O��	�@�	��S���w���b��yfhL8Q�_EU�(nt~"�D��'����3��<`���hqa_�=���K�<	���?����?���?Y�����BB�!�AN`&�FX�yN2�'��nӰ,S&?�����O"�O����QX���lڌc�^a�H(�d�O��4�~��5�qӐ�Ӻ�䧖�|}��"�M9k��9����x�N���(bN�OB��?A��?Q��uʔU � J��h*r,�.4d�����?	.O�l�z�(8���$�	V���	R��ևZ�?i}������$�<Q��?�H>�O�>�;����dMZ�A�q8��bt쓬C�8�� �ib���|rԩ��d$��a��6'����^�$��jb+�̟<��ҟH�	��b>�'H�6�0�܁�$�)J|9��P�qe\ �m�<����'��۟�kD`��N�f�ץ+t�=qF�����I�>$�mt~R�S��e����ā*G�nm� ����ɚs,��$�<����?����?A���?	,�*xXX1� @�g����|�5@�˦�2@Zş4�	ޟx$?�	ğ�<n?��Q�)�n�@1I�@M�2���ϟD%�b>�BG ƦA�N�Y�3$P46lH���*� ]�'}���h?�O>�+O��d�OFHA�Իm?��xUb�,SDi�m�O��$�O����<���i��d#��'�r�'PL+C�U%9�"d�sˌ����V�d�<!��?�M>)U"X�+n(���8��,a�g�W~"�ӭ7C�����iVړ��ta�'��H��	�n͡'�M(��!��'�R�'&R�S�X�΀��^Yx5.	����A�֟���47�*!�-Od��$�i��#�O�"^:��*�SIഛ�p����ɟ��ɳG�n�t~��T8����'Z��B7��c�Fy�M#Gb�*K>q+O��d�O:���O����O4��E�v68I��#>���p�*OV�lZ4`���ԟ��	d�s� )��^�U�z9�Pg��)���Ky��'*R�|��@�[<���XL�i��[-	�k��C"����Z8,0��A���O:ʓ[�z�`M��D�n�����CG�4����?���?���|b*O}m�0[��ɩK��07ON8J;~!���,��Iڟ��?i(O�D�OF��K2=n>��D�	>�r�P��[79r�yp�l�z�nݐ�P���8�>y�u@.�M�#�ص��!��9p����4Ʀ�A�\(,�`�f:�Э!��߻ �Ea�3d��p�`��s:��蟚�@�Au�1RӋ7�x���,KY�ܰ�aH��7�~%PR��ߘ'�|-H�ޫ.
�!�P!R^�.)W'+T���
�A�9zU�tj�/kI�A���ۡ:2��[�"U B�~�R�%!@�b��`Dً=r,!t�%Z>��Ԡ��y��͈���Hۂ�¤ �4[1��z�K܁����
+F�=SU��+J��!R爇(����
tn�Y���3Eޛ��'w��'j��x&��>�+O��$��(��+	'�^�kā�0q�@"{�ޓO����Ev�˟���ǟ�
瀘�F&*��bW!/G�A�1�M��M;��#�.�j�U�0�'��|ZcT���I@- �TY�b�#V��1�O�,���O.ʓ�?I���?�(O�����Îtb�S�(h�(4�ВHn ��'������&�4���������J
�7I�,R���Cg�c�b�X�I����Iy��_Q<p�<%���!gӯ6.�0�!��6-�<y���䓹?q�H����'�v��TI�S���Ý��`�O����OH�Ġ<��"ԀV4������4ʘ))�l���[>�ܱ�iĬ�M;����?1��v�������I�EV2��t�؆Af�9��#ܪq827��O��<�"_��؟��	bj �D[f��S㛶h���sm`����	 L�N��?A�OO�}y��.h�x�F�ʢ@�VL��4��Ā�T�n��h�I��yZc��5�@���Dh�](���O��YS�4�?y�L;��B��&V������f�{Ei�`m��ŕ�0�46��OV��Od��HF}�Z��0�fܣ"M��o��D�S�T��M�c�O���'����Yh�dip��ܨ���>�tHmZ��`�I�����锼����<����~¯U,GF�'���� D�P�+�M;O>y�ˍR4�OfR�'�ˑ
]H=�f���!��A�O/Tr7��O<T�#��|}U�|��G�i��q���P?L���=7k�|���>��M����?����?Q+O�����q��A�%M�o����d�˅;��,$���Iǟ%����u��;\RPh�s��ia���M������OH���Op�a��ĺV6���h�BT;L�8� q�VoT�T��U�h�	؟t'�l�����'�^x�R�'(~�<�m˜<b������>����?)�����ܬRr`%>Q��C�<���@�D�#���b�և�MK�����4����1�Ġ�-�u�q�#�<�rE�@<�M����?i,Oֈ�K����s��9�o�>����P�?���w�)�d�<���?AO~�Ӻ{w�΀[�r�!�
��\+����
RY}��'��R�'���'=��O��i�A� *�3A2ԭX�Aѻ�^��1Dh�B�d�<Y�Pq���'׮u � �wN *��
*(0�l�� u��͟��'���U��'k� L���g	N��R��T�@U�İ�m;�Ş�?ƈ�� �<�d-�'��#�c9��'���'�ĵ��B'�4�\�����i�eZ�RXl�;���,%��vk���$+�dV��O:�$��Ș�# �W"e5'˽}+��(�{�h��%B������s��f�h� Q��Y�6Nҙ{^��j�x"�C����O����O�˓J�ls%�!��Y)�@3&6����6#��'M��'E�'L�i��C׏�A���(��N�~�ۇ�aӢ�ĳ<���?Y����K�z��9̧�`YA��6M���k�߀1�J��'|�'��'}�i>-��
,����$�.�
B��q~��O���O8���<��MD�!B�Ov�p�q��
0�ƍ�Vk�,z̥s�av���$;�d�<ͧ�?�I?����G�>�Z�H�� b�J��tӘ�$�O˓ y\a�e���'��\c�2AgFN1"Z�9C̈�(X+H<+O����OГ���؊�Ț$K��F4j��1Pбi��_.�i�ߴ'�Sҟ�������=9(L�����R2�I�\�O0�6W���I��ЂI|2M~n�Z4f����1)�00���4��6���F	����������pyʟj̠v�;8�(�܃����`]K}b˟&�O>	c�$��H0ǉɟ�X����U��M;��?1�R5���/O�Sy����0�@U���.'�H��D�Z(��tFx��3���OB���O�����F��0x��bٵ1�^u���T���	0 |T��N<�'�?I>�;�������-gg^�1d��.���&��	g�I��\�'�b(^�Z���r�ߙd�؈y�F^��怣UZ�p�	؟�?	��~��@�"l�!��U�|CB���!׍�Ms�k�K~2�'r��'I�I6p}�OU�8 `O�8(����ME+$.<q�Ov���O\�Ot��|
���p��F7?T�Q�T-XI�x��S���	ܟ���eyb�	"�l�rjQ(O	@MW���pB��ɦ���h�IVy�Ojr�~z�h��rTY��	�/d�!� �Ȧy��؟8�'��Q�)���O����h�AT���Mz4)Ɯ[
�0�x�X�L���H$?�iݥQ2���YаQYv(Q}0P@w�>���'��K���?I���?9�'�����VK�s�TP���.p��(�Ѷi�r^�|���.�Sⓛ(R���J͈)Q��"7
�06��xp�m�ٟ��I̟4�S>��d�<a��ˇp�T �ᏼb5�$����%�V����yB�'0�x���?�H�}���K�i9Q�r {+�Nz�6�'�2�'���W&�>I,Ol�Į���F�s�����P��L|+�ϫ>�-O.�擟�şX�����P�V`ee�K�F����>�M��0���sWY�ȗ'�_���i��Z'��V4�����(+4�>����<.O��$�Oz��4Q�2��2��L)�Ó&W���k��*2
!�'��ϟX�'���'?��
�I�F��2M��=�Nqp��R�'�2�'��'�r_�L1a���D@-�4Ad˫t�"����T��M�-O����<���?y��&<��\2��谦��dT��YC΄�[E~��W����ן,��_y�7��맺?��	N�\br�#9�;0�7p���'_�����	�� jd�1�sӤ��e�L�s�ޑ˵�8<��xز�i���'��.x\|X)��`�$�O�ɕ1k�"����Â�Qs�ÂI�m}��'�B�'��#�'�_�D�'D��l7�Գ'��x���_z�PlZ^yA�7!�7��O����O�)s}Zw��8x!ظ~������[#�jش�?�e�R`͓R�s��}���I+�e���"LTt±�A��q�7d��M����?i��R�Y���'uZ�6����
��ɇFLd�rv�wӺm:�6O|�O��?���c|��C�p9����-O-V�!�ݴ�?���?ip�2��	Ly��'#�d�suh��
:ϔ���Ʒ7��I|yr��)��4�:��O���\284�)�%j>T`�O�WZn�Ɵi�b�9����<����OkL\�"H��A�H�<0D�S.�p��I:|�Z�ޟ��	ߟ$��ȟ�'���!1�J7t��5)�?;��P5�������D�Op��?����?�ԩ�r�k��E,�*4۶��fj����?Q��?i���?I/O@��D�|����'L���f�
�̈`k�Ԧٖ'�T������0�	4xh��	-f��!�M� T`�:��x�ٴ�?����?�����D��!m��O�Zc�X�I�����F4Fd��4�?�+O���O���2bw��|n�!PR����#�#>LI�`!��\�Z6�O
���<�GZ(]���џ\�	�?	Q6�R�k&�")�4&�1Q����$�O���O��;OR�'�?��Or�!��d�5j��P�2E;�2}�ߴ�򤖚.3\�lZ�����4��5����&��Ι�e���ъ����U���'���^&��Ļ<��DIU�6BT1���1"z�P�p�W�M�gEK���'\B�'@��ƴ>�*OB��ׯ� T ,AA�T�/s��J4��٦9q�B"?�.O�?��I�h�h5�W�Cx�)A��5M��9��4�?1���?����;{��ISy��'��d�#m�����>�	��B�՛�|2+���yʟ��O6�d[�CU�1�gK�&��P�I���bel�㟌���/��$�<�����Ok� X�٢��$�P�(�/����i�ɝ��yb�'�"�'�2�'W�ɠh*p��!��z�D�xìԜ:�(|�A"���D�<�����d�O����O��Vb+^ȉ�/�
<	"Oه,)�D�O����O��$�O�˓nt���1�( �u���	�f��Y9��,+R�i�������'�"�'��E]��y�-�$L� ��	�<E:#��UM�7M�O����O����<����	7��O�$���AҨF}�;�(S&H�u�1�s����-�D�O��$M�a�d#}�9cEv��cHNAy�Y�ҭI��M���?A(O�5C��Aq�ğ���=c�e��ΟR6�(��&�$�jI�N<Y��?	"o�&�?�K>��O�|�p$��;
�x�A��e �H��4��d\�6��%o������O��I�r~R߮X��ܛ�ѣ(�����L+�M���?�&m���?YM>q��4D��v/ڸ��i�q �1�����M�P��Z�F�'���'����"�ɺv���{����}��(.�d���41�,5�����O���Y56�C�a���萧��;o�6��O8���O�(d�S쓑?1�'�
����H�)���!£�7�|-�޴��Z�m�S��'���'���	�f�">�|��c�1��y����#z���>9�������lӶv��aǣrѣqHl}�o���'���'"X��d�
5T�0�LX0��w�W�G�HKK<!��?N>)���?����03u�t����{k� q�Mܓ}\0�<Y���?)�����¡}N���'uJjܨF�	6�H03d6>*�T�'*R�'��'+B�'�Z5��'6n�J�QO��]��fG��8�hs��>����?����@%Gu
�$>yAtH��Z#�yr����B�E;/w�)�ڴ�?yL>Y��?�vj[,�?YO�p���*jg���g�ށ!T��!�OjӼ���ONʓݠ�8ԓ��'�����5c�=���V����r�0Z4O ���O��8O��O���<~!.�$g+2n��G�ik$7�<���>	&��E�~���RW������	-�3vM�����|�b���O�,y���O��O��>M �
ݨ\�Έi��4(.�m	�|Ӑ�y��٦���˟��	�?q;�}�
��1�z���ήa�a gJ�)\6��,��$"��>��˟�����}Fh!+c�P,a�0K��)�Mk���?��r�,����x�'���O���/�:|a3�(�,d*ֶiY�'�He2G�-�)�O����O��BR���ik����?4UzU��M�	1T0���}R�'4ɧ5V"�p�����;���O ��$�1j��D�<����?)���P��ꝪaK�^	J� *��+AT��V��O��$�OV�d�O�OT�D���i�Gўaęb5'�.Ը���Me��!ĝ������@�	XyB_�Y1R�S�(�� ���іmz��jN�Y��?���?��(^.��)��y��!����z_�x)'��!��I�t�	��4��P#�E�}���'�P��N�[>���I�,����G {���%���O˓c���&�����i����&��,��� �{Ӝ�d�O��4#l	d����'������`���BNO��\0���&ɰO&�D�O((��r�4��-Z���x���O��5�'�>�ȃ,t�p�O���O0D�%*&�ӡ���� ���r�<n��p����"<ي��MV�"lh��%/+��U�LԵ�M��
|���'�B�'���/���O�����=x$�YX�-\ ��7K�⦕�q�!�S�O���
�xҥ(�U�^�2A�őg�7��O�$�O�A[��a��?��'d,Q��h�xL���A?7$�j�}�$����'��'��DE2���i�n�f�8��?H�D6��O�U�L�	����	\�i�JCg�^/���$ @�j�걣��>	#�u��?Y��?9.O8���n%\%Pe)�",o��ۀ X���$�(�	蟔%�,�I�p���#6��=�-R�gfDIa�`%2) c�L����i�lڟ �o�eG,ρM`e�5��t��Ԧ��'�r�|�'��ɤVv6��}�ؑPl�b�0���%^E�I˟L��ڟ��'��u��"�ɟ;A`B(=o�P���%M'z�LoZڟ�Ij��xt���~�q-_a�L٢��I���$����������آ��~�4�'��O�"d	�	W�RxHb��4�b��6���O �0G�GxZw�r���	{$h�Q"Q1o�>0ݴ��D����to�
����O���w~RJ�C%|��j�p���&aդ�M���?�׆z�'xq�ƥ����6R9�@��> ��}Hg�iwXA�4�f�n�$�O������?���(�6$� | Xl ���u*^u�۴ �pDx����O��ӷa�q���u���s�qxb�צ�	ԟ8�ɀpc@,�J<a��?��'� k�
@ rX�=p�b͌HH@Ȫ�}Ҥ����'Nr�'�r��7n߆%CD����@i��XE���j���h��?!,Oj��?��۰K��	��'k��������D�$�8�v`<?����?i�����<^���Ɖ�.'�Ҍ�G�j|�����{�	ϟd�I��?�R��:<dZ��G��3����B�Y�\a�<����?���?1��C�
���O0@�k&.�2VA��iw^q��KTͦ����4��o���0�']�=��t�? �|��'�<1%kGܠ��GY�<��ßЕ'7��3d/�'�2CO�
D��aR:��0���N�6��O̓O���<	�i�s�4B�^qI�� ݘ؁ ��D�6-�O���<��[!1��O�B�O�^)�ġ�--�B�sJ�Q�ȐSG#���O�������'g�Rd#�c̟(��!��:E�lJy���'��7��J�t�'���d=?��gD�C Uh�W%x�X�y�%Nᦉ�I�|�5�3ݸOs�%���O�e߾�c���=���9�4]p����?���?A���?Y���)I,>��1XpΊ�G�z�����#_"�$�'�R����I�O�1XcA �:���WW*���DEΦU�	㟬�I�G��H�I<ͧ�?	�*d<�YD&�!d8��R�ݯ��= F�ć�)1O����O&�D� Y$�#�úY��|aƯ[�W�l�mğ�8@D�ޟp������OԒO&�"v��%�Z�i5��U��P��m��8VU���?y���?.O���R�9b,���"������(����>�����?��GS�%�Ge�.��u�%�̲[,𹕫�f̓�?����?�*O������|�㢀�~��<��_�}@yH�-\A}r�'�"�|b�'�¡�8��Ć;�dE�2�^
WH�Y�����	ԟp�	ߟ���ݟ$x3 �E�t�'u�jM��J���Z�ՂgLTYcA&v�`��7���Ob�wS��$��r�� C&��]���T
��r��$�O��wK�=A�]?��I쟘��ovd8b`�8��0�v��~�ZM�۴��'P�"}�'}�T��
7�TH��I }b�%8�4�?I��E�,1I���?���?����?���TܵO��4�Ǉ#��ˢ��զ���[yB���O�O��Q#䏒]��9 ���v3�D��
?�6���0>��勦#)8��Ā�8��$��o�K�<�e�+#*��y&�ޒ7\��H+�(8N�bc��i&�}�g߃2�J� C`�!7�	9��ٜ+d�m��)�<M�� �/6Tx*3J�,
R ��<: Z��<��y`b� �W�8�a""�;�j�I�02"��e
�(6j����=�tG��c�8ga�=3�����!�?Y��?���=&�.�O��z>�Ue��"�$����"�gL��(�#�0R ����՗T ���d�&�0��R�	T��8C��? �l�kbn�<Z�(ZB���d�tY45It�9�x���d��0K�
�xc��d�Q
�����	C�'
�O�uB7�F9,�r92��d�q�"O��1�C��n0���*c(�ȡ���U�	uy�oɠV��?�l�`�b��ġG��<�����?����5���?i�O��M�d�T.�|ٹׅˤQ��q!���Y�����8�|�H���y8�PQe��->�0�*D��,a��� $tf<��N/J!f� ��Ѡ8�x��[;�?	����D^�{�T�!���8e /A�]��yR�'Լ0u�)S$mb��L�FiJ����+��|�W�iT�[�  S��H�0!֪j��0�'��uK~�9��|�����Ia� ��V��w@^�)�lH�b�	B��0���?")��)�P�/lm0�����|����#s�~Uq��;��L0 ���$L22�9����[r�%0���O"0��]���)�QaT�b�A�@Y���B3��.���	ɟ�D���'��JA%��O�� �G�j���'�>-Xdh��s��J�ub���3�i>�����$~9hmr¬Q(���f�*\i�AlZ���	��Q�ɗfr��I៤�I՟�]"v5�em^�Hs{d��,qz�cb�i��ɷ,�j���1�3��ƿ?��-�w��89�1J�_$&�d���P9����N��q1��L>A��J9Ɣ8K��Yp���h4�?��O�)�����	.�^<�҉S�I���� B�=DrC䉐r�N(�b�#"�lH��I��jp��8�����ğL�'���8t�݅fH�h��[�\�69�k�l�~ma��'���'�R�m��I����'ZahM�4� �	jె��
�8	W��HmĐ��B�\��W%	`H��r���f�f��$���U�#aP#?�2���Iw$XJ�'2�9e�Q6
���m��4���uQ4����.Nى��^������(�DG>v�~�pfMA�y�Q2F.ƕe�1O�mL��?S�Q������N@HVES�v�((�Vj�)�����O��P�O��`>Qu�;�찑����\mZ&r� �D��"q�H��PJ�'M,���ؽC�#�-O�u��� 3fd����%Q�"8q��
P)��i�!�'x����?�,Op-��X�%�l����d~ ����D�O��d@�>�6��C�)u��dkc)�	L!���¦!�V ڊf���	�������%G�ܕ'f��QT.lӆ�d�O�ʧo2 ���D�|(�A�X7N6F(�� ���?�Sc�}0qB	v�|�����)�|�) �Z��7-ױtZ�	��D�P����U��4ZeEǞ羘x��Y��M3��'��	�*M>�ѡ��U�
#1�`;�I[�S�'	¤#a�ʲ@���ksE�+�����S�? �YY�-����,��^}�,�A�6��|�S�I���I�)�!����R�{|��Aܴ�?���?鰆� ۠�����?����?ͻK޶5����t�=!S:+�鳌y"&�!��<��͒T,<舵��k��:�e�@�Ak���I>@����Ȫ��`��w�	�<! ���>�O��A��c�@aHt� v���"O4l�ccF�WVQBq��/B���" ��PY��4�X�O�q����:.��}�̈́~"FŃ@eX�F|<(���O����O����Z�t�'��I;2z&lK��q��0b��b�IY��RBת(E*ͱ�j�?:���ã{8t�'!(ͩևM�x� ��#@�������,�?����?�����$�O����D>xlzRjC�f4!Y�H1D� ��fš!�<KqN�E��yq�2����<aqMR�����'£]�+Ǌ�b���^5Yb��r r�'ֆ��A�'-�'�,\���E�:��O.9(F�%md�B��/	�X���'׬ ����z&i�K|�!H�o@�36CsD�V�D����c�џ��Ov�D����I�䊕��şo^��b�����'xb��ӷN�p�;g�(|R�h�nW
K����D�O@�\��0�(ނY�����	@R�\m��.z��=Q��$R<
�T�R"'��b��P>m!��$�$��2�����,g!�$�_� �*��Tl�m�`J'z+!��*(+�0��C�}�^XA�)���!��$I��#6$ l:V�1�i �!� /�n��R	ӰP�!�5հ,�!���X��p�'ƈ6��ѷj�	Z�!�$ʺmդ`�2�
B�Qʅ��!�!�-�+ҋI�N��"	*�!�$Ҝ���`gBc�r��e͖�L�!�䄫Y���$��'�d�è!l!�wf(��m� xy ����ٱu:!��C�[_v�����[m�ht!�dA�ب�c�Q�aX��R�E�W!��/dQ���G�/HNQ&d�j!���v��zQc�9�8dC�d�]�!�$F1x8����!q��AAv�֋B�!�d��< �I$�3k�貄`>w�!�Č,��a(#�XLĐ�.�!򄖀D���)+Dܬyv�K�1�!�Dy�m!2M��l0���2$��!�$\Zu�ĳ#�#�d��L��H�!�d��[ ���B�l�\���V�!�D��9�D�C�H��0D<ڑ%�|�!򤆅?��A���,��`CԢ�!�N�W!�)�7B�.5���cΎB�!�d�2n�Y����4�1@���P�!�O�-�����gX�2�=Z�'˵�!�$Z��Ų�EO���R�^�!�W�{�{���PK~1�Ă"}�{2�VF<�`R��OD�(�E�g1�l�q�N7L�YZB"O*���J?�v�b6�V&<4�T{�����ng�u�����H�dAR�iˢl���j6J��$"O��0�͞B�bĉ�+G&n��#�ɜK��i�-G^�D'�g?QSF
*{�DЇ"F.�YP`KI�<A�Q�vb]*a�Н7�Z�*�@�۟x�'קn�9��'�J��OA�c�X9ٓg�O�:rߓ9qv��R"3�Z7��_��pz�g	 X�,2Eh��.�!��̸k���x��>e=�e��
9n��O,|aG�ٛu�ڝ��Ɇ&Zߴ)ʗG��B|!�c�i�!�dq��em� v�n��f�� R����HO>�7��>*U2��.��颐4D�\2�l�')
�� �D >��m���.D�L#E�I @�t�ea�(���R�,D���BAM�U�����/�x���!,D�� ��A�M,1I�!���Q�"O��R��
�Q�m�!B��t(a"O���ݨW�d��,٪R�l�E"O&=�ƠWHрH�኉(wa�Cc"OT����$�$����(w�JA��"O��+�j��J�h0)P��67�]��"Oiԥ�+$���aHN��p�w"O����)T
��-�4)�5*�;
�'k��!mƁɰH̗o���	�'�&5qp�޲K����Ҩܷg�\i�
�'���`��\>�:ҍ��Y�ژB	�'���W�x���&f��9�'3��B��S)V�,�D�V�Gpلʓq��,Z�i[�b���#�$�*����ȓK��VZ�4�"���T�[�VL��z��3w+�/�<)c��IsȽ��vp�0���/y���$c�:¼��c��\�@�܌-r� h��̛m,L��N'��*�Gċh|z��G�u�^��ȓ;B��_��*�� hPXJ�ȓY򄀒��/RUZt��m�~�<��^:��ķ]�R�QT\D��ȓG�03��ҽ(Et48v	I�NbԄ�gyH�qƤ	��,L��SL�DP��HAn�bI� [��,*P�4vr��ȓ�j�x�i�'\뺡z��@.���Q�
Q�?�P2��́Q��ȓ]���gI�R�~9R�L;v�i�ȓ{B����H��W! t��B�\̅�S�R`�=!u��XېT�d�/�2!hSA]V�<���M��(�Sҿg*���4�AP�	�{GDa�?�~��ʇv�x�`�͔�,��x9U�]G�<IqA�S���́>$-�ʞ�t�� �6ɒq�Y�E��<h|��}&��3u�&	�}3�'܌y`��p��8��1��(yh�\�F��z�x	�(�9�j��
ե�졪����0K���p���@}�<�O�~��	���Z��J	NI��@n��c�Ͳ&�ڙ[�Fڗ7�r ��I��'P��{6C�p�hQH�!{V��9�ō�c;�'^�>�DW���ͣB ��f�j\ ЄLl��I>�Ի��t�ȩ0L ����҈�ī������� I�j�ڦlϸ�~�ħImi
��'��Q��J%k�0!au���ؙ���7fdP�"v���rǃ����'WH�2G���l��7͈'t�82��>Jf��W��~B�Ec^PX9V�)u���GE^�5�e ��Q�Uޙ��˔�d��W�A6 %�y��}��'-�.x�0m!Pn�'a��d�$#ٗcp">���m�Jl�" �LP��� ><0�`����501�ɂ�0%؞	��[���yC�c�(��'��>����s~��[�=���)	>����OJ�v�	p��M.cilmb"jܬ?�vY:���O�%�d����l{���샓;g�	�D���=lOܙ
��N�~����O�x��
2ǅ�P�lբ䏚;�|ԉ�쇜@��'U��'�T��KϤ2�Xe��ݯ�43� 4�T��CW%�@zu�[�C���U>S�\%R4\�7�<d�7�X
P}���ɇ[Z���n�?sX	��AKPOX�?ᖢǚ-?L<c#D7M��<b��&N��E"_�N+�f&v�PW̚h�<9УU�x�7�ȝn���[~�g��{�\# �I�W���I�����<ؙW��@����v̙�m��`b"O�hj�вQ�����*;t��D���F��,s�韬`�K��-�q��'r����g��,95�R�Z�y��'}�)�6ǖ+^-�bD@ʺo���hq���+����.�&�$��
ۓX��Y�Eǜ'>�X�䆓�s��%��	�),Tp��ى&|牅"�Q���_�l�25X�C���C��F�Y�C�z�Q	��!zw.b���D�νK��~A�	:=�Ly��[8A����.����S�'3b�1Dd��K�m)3����@ϓC�Mi��%�$�/\��A�J�t m��!<2C!�d��<Z��.ZT�Wg�B��'\
�K�g�T�S�'rK<]���)
3���%���$��S�? ����W	�ؒ��Ur�������=[l����L�@K���V�B�[8a�h��!D�x�4Ꞅ���4b���HR�쿟4����4�t��g�@�O�%�̒C��C�I+�p@y4KF4>�T])���q��C�I�a����\9I�F���aĆ<5�C䉏6ֈ�hÊ	2il�@1�pB�Xkx�zO�.��	�L՞B�	,q�΁����0�΀B �j�p�RY���� �M�6	&������B�a㍚�R�S���p?�,��R�� �=3�a
.žc�Nu�2)/dR�s�'���)�G�;K�Xp�&R���C���K�pԉ�D���A���	Ҡ�,WqTq`�a��Ub`"Ol1�6�԰=�;enA�Nk��C$�O��h�+wTS� �0|r/��D�j�AEO4)�苰��{�<�WKV-��yPҤĳ�t�k"$@�y�t˓��M��������'�9z��i*�����$H���'"O�U��	�o��@���M�¦L	S�\�HɌP���P�v�����a�A�A	P53��� l<8!��O�L��֧�����s�f���"O*�x��L
Cla��NŨC3r���"O6Y�u��pn�%�g��nD��f"O��� D�'�}��$R*���"O�9Pv�
�a(��=g�0���"OTH2 M�Z�&�C
=�U"�"O�����^�R@(�Q�uƈUC"OD%j5�M�]��[�,�#���"O�-sv"�#A��U�d��.W�c'"O �Z��ŎP����
�U"O4y��[�~�4�����|:l"Oi���(c��i�2*�'(T��4G�V���$��#a�R�3
�''dir$/˖t4����8L�����'�B\�ulPj��tYB���H��I�'�Y@&!ֱD�>��!m�S�*|@�'c�1#J��n�� �E�M�DP�
�'Q�-j�L�$\lf�A�%DKF"�'�,�
A�M?��В�.I�F�p�'f��a��p����/�%o���
�'p� $��{NȔQ�C����u
�'Xp�c��6�L	d*��z��2	�'�6D1f�+8ޤ��sI+n�8��'gp�ZK� up��
'1 ����'�T �⣞�MM�� ��?%ƭ�Ǔ~j&AG�V�T�X7��5 ���`d��}y|�(Ҁ�J�)#Ih<ٳ�Z1:vN"`	o����f�Yw��*֞�3�͋�js�|k���+F<c?��,J H-�H�Cf
/!�u�a?D�l�F/��Dsy�W
^:j5�}y��ܴo��)
�G��x������ؕ��>q'���G�G�OXJ���-$���<��cBC�Nv�ɳ��� �Z�P�AAn�1�䇟>?!ZI@������	� 3��@"T�Q���� ��^k��D�L�$H���A>3�� ��`�2������^�.����¸�)h�O���E\?Ԡ�jj�pq���I�?��0�֍ =��`���B�0��ȃ�X�
Ԃ��c"O�|�qn�~)�k�υ3�`����'��͡�P���|�O?�s���uP���h�|���ހ�y2�J����h��ȔW��
u�O���&[N�C�+շ��<���±(��x��Ǩ [�i�aB�\���,zrH��I�CJ�c�@E�$��R�\Z�$�� V�Y�ȋ�^/��a���`ڌ0��w"(]A�@ka¯�vG �	�$AX�<���
9<Ձ%VU9h��mR�<�d���_Ԅ�E`�<��]����P�<��ʘ6<(S ��7J�P�A���H�<� �� �6�y��� cH ��"O:e7K�9tI+��OA}4�4"O�� ECWq�$��+��*���"O��o�Q�k�
s�*�b�"O�%�ī�vi�h�E��� ����"O��FS�U<������qr�$�"O�rcfнW�f��锰3dXZ"Ob�ITE�;,aI�h�!1Az%@V"Ox��C��Nh�m�愥[\l��"O��#��%e����
�O�2U!"O� �&���,�h)j�IɄ~��|4"O��;`��a|8�Y&H��xh2���"O�+�K�2r�jH�禐��d�"O|�1w���Tf��%��q�s"O�#5H�7ݾ��V��<��̰�"O$m��|`��K�D^=ju�d�"O>���S�pF����#�sW���C"O���,�'>�
�6��($��"O�
pG< ��tC�9K2��"O� g�3?�P��Ȕ�"��z�"O�}㤤�4)���u�
�P�"O,�KS#Հ �m�U@vw܍:�"O��!� �j�S�-׀vcڕx�"OJ�(�$�l�ع2�lR(Vf`�E"O֔� �?��8�lT�5H���"OFq 6��7N��s�4��k�"O�@��ք6�$�IE�0(�P�"O:�bUυ,y�����)��H/���"O��S ςފ4*��F,jMɇ"O��[ ��Y���P�)�>1hx�d"O�x����2{~Vi �(H-����"OLh�@I"��qZ�g`p�{�"O������6"�f,��ĝH�i3R"O �;��M��C�đ�@(��"O"�q2�]< ��UC������"O	k�N�n��  � 6�`��f"O��"\��2��D{�"O�����O
9x�\)q!��"O*X�LFR��OO���X�D"O���r�]�1j�Y�ڇN�4=3�"O��c�'�A���rp`�q�&I�4"O��*�+ȓh�\�	EE��|x�	�"O�8�T\/ozxHs�	�!�(�r"OziɃ*��~5H�zL5�eX�"O��x`�7m.���	�F%8"�"Ot�uDN)��`j�@,'���"O6qkY
9���@CƵ���Y�<!�ޡ�x|��K\^���y4�MJ�<I���	�a8���I�F(���l�<)C��.�D����$����h^S�<	�FáS�8y�C�͡��ìPO�<�G�֑�
�bueJ�Gj�4���c�<i����`7 ��!4J����&"Q_�<Iw�A1��R��*��,�c
S�<6떲v�t�p'O�I�m@�BW�<�Vܢ&���1JN�a2$�V��I�<�V�I�Z���@A�'F6�i��A�<�/
z��2Y�DxV�z�<y��N����qnM+Y� ,���u�<a�	D>0��pǢ��ʹ��$e�h�<�KC�)�2m����"H֢�G�Ny�<!/�<!��Ia3"&���l_�P�!�D�0f�(�Gk�>1 �̓��߭a�!�܇8�P���ߔ.d�P�_�f�!�� ��ـ�5%B\��Èvװ��"O�ca΋Q68�����|,�P"ODP��,��� {��,[a"O,Q7a�h�p���&9��"O�=�F��FK|z#��?��@r"O(5��M�yT�ˊ:z�z��d"O~���˺`�Π��
D=�Ș"�"O�0��L&ok��آ냜xw@)E"O�����X��HP�\Gݸ�"O�E�R	 P�J<RP�H�%1�m��"O��jGL�S/l����	��-��"OZ�1��9�>۶�nT��"O���N�6�x|�0�ց3��l2�"OΡAO��=N���&ǚO�z"O�]z*B�,3��ʹ{0�p	!"O��2����6��Þ>-��"O��(�fZ9��8���">���"O�a��M�>{�(eĪ��:�D5�"O���'��[�$$�QD�d�"O�d���&�:x�-�B�A1�"OV����<GB���5�P�"OJ�
�^9�L訢`�7J3���"O�r1o�9l�~��oؗ,4��Q"O�PZ�^�Q��Q�,��B���1�"O,��#;��hSs�ڞ|ܐ�"O�����L-|����m���D�]"!�V�7��,RhU�5[FL�1!�$ �5I�2���h �� 0�N/
!�D�8$���(7@F+w�\4���ޕ !��	����˜�yӬ�� �m�!�D'x��Ҡn��:����'
 	a|R�|B�\+6��a%�?%���K)�y��l};�'\��LD��y�(�2:/B��UeA���)B���4�y�F3l�&pj�`���@UӐaY>�y���B��̦%πi�Æ��y��"U(l����6.�`�G���yb���]Ԧ���(=�-[&ƀ��y2"G�&�0XZQ�H�B�x�	ָ�y�mݿ"Ob���>@�"��$n�+�y�J�,s~8M
���l�����U��y�i�^�L��Ab'R�p.K �y�+ʠjv��0ˈ��H�{����y�H͈'j��$��%(2 m�6�y���T6v�v	��`<Xw���yr�#Z�	�u
�A�< 7�P+�y�ǉ#j��q���	�V]ȖI��y�L�� 2�L�aLQ:�vqQfNE	�y��D�A�H��앣~�X��t�݆�yB��F��u��P })��i���y�MJ�DmL��N�r9X����L�yb̛.&X�2cpJ�sw&ة�ybǉ)]�L{�5_��rG���y�F57,h��a2U��ܺр���y�����J�JA��!��y�
Qk4�
"j��rC���!E Ѹ'�a{�k��C��EB��O�BhO74��(Z�'m�4K�*��`v�*7j�/z�A��4�PxrU%(>�u�!jR;���r�Ƴ�y�脺C�dh��ɭ/�Eb�M �yү��I��YFɟz�����LW��y��"�M��I�w�8�C����y2!��7�̛��8u�8hj3hѤ��x2H�z��פG#&��) ���/I�p�h��� �I�0�.X s� X=z�z$�'��Oj���1D��% ���L6攚�"O4�yAT=3�(�rCE_?MY��0�S�S����E�6M����3`�/y�B�I/K�P��ؒ\Px1����B�	�[<�[um�X���Zɉ,A��B�\�PjN�~c��spF�C �B�If��F��	i�P�Ö
JJ@$C�)?2�yW��l�4���I�
<C�I'P�~����/~���Yl,C�	� �qS��"N����M�
C��9ʹ1!��ftb�g�F�$C�Iv��}���7��d��cJS�>B�Ɉpk�L���3٠�ADhվ~rB�	�nV2�Ê+\�r$���nG�C��0��Azãԑ/�T@giA�88C�ɑ&9��)C��:2�"w �%UpC�I�L3�0�%"`�(TCa�0��B�	!nyv ��2tO��`JW
��C��P�I����-��I�� 1 ��C�	���·�E|p#��Y���C�I�O'f��T	�|�4Lyӏ%WfC䉍�����[��u�էU5,�0C�I�cQ�����09�r(�t)��ZUC�	2RK��+Uj�p�१�+c�B�	�b{��A��$Ե�GC^�y��E�F��A�ǃˀ-��I��g�y�]�r��qb��ޟ(���f.���y"#ǥp :!a*Ϯ�.=Q�P��y�FM/?� $��;A ���s�ؙ�y��7��i"�̽C[� B�y��]�3�[A��k��=CeY�y�."�LS���V�Zű�C���y�&�-N' �`e�F2"_DT���y�CV;3�k���2x2p��N#�y�.����S.�	/�iJ�f�(�y#̐�nU�ٲsCZ=��϶�y�k_d=c6��:Z:.��6G�,�y��Ȅ>`�8#1��"=��í6�y�kpIxG/��^" 	�
μ�y��_~�@Q��� �<Zq�珍 �y�	�r��8#�
"�&��p\��yB�-Uox�0��܄!�.�1 F#�yB@��nt�]22`���@��L��y��5ֶ<�6���7�|ؒ�I��yrĄ\�m��E�*�H,+���y�G��Q%X�ZV�?"�d��E��yB-�6c�N����a���X�yr��`|P��k�6���i�0�yBC�?N� �ٞE�=�Cɽ�y�ȉ;���&��ApaHF<�yR�٣0�Q� �J4~mN)��L$�yRIM�zcFy �kV�eb��t�N?�yR�R��l�Ąd��A� �A2�y���J�ݨC��$^ �����y�*R/f-2���W����H*�yB$H<t��(��Z7U�t���2�hO���I=7($E��eB�i��)�	t!�Ĉ }w�Dk�������l���	`x�hT*Oovl%�V4fkfɘ�8D��h�	�	z�"r��[V,��E6D�@�A��j�n��B��o�,L�V8D��0���Ѐ�)vfзnY@$��/:D���&P>ar��S��3t'.\C�8D�� B����/HV�م��h�ƽ�1"O̕�4���cu��hҶ�d!��"O:�i�m_K��� �O�"V�j�"O� cv�šc��k$_6���"O�����{X��]6 <@��"O����޾sR2	aeUH�t8�"O�)��H����l��y�"Oj���޲z�.9I5*L-X����"OJԪ�F!d�� ����		�)!�ĉ�OJ��������)�IѮ(�!�d #]F��!�`��'���K��K$@�!��( 2�1���p
���X�j!���;Gb\���GZ��Y�,�2"!�$�!:�����M��jx��E�aI!�� �l���J�~.�x�'˲07!�ę5J�.L ��6J^i�d�,�!�Ĝ=Fx5`�ʓ�`��+�a�!�DNi�^p[R��(��R����!�D_�<������J.9�Փ�.ϔ@�!��)^8�KrK�ձq�{!�dʎc�<(;��Bn� )� ̝�A<!�dʚn� ���"}�ƙ�%H�1�Py��5�Q��i�64Y�%c
�0�ye@tJB�pU��=w�<�R«1�y�G\T�M0��ݼy��B�C��y�I�&'vX ���y'~�YB(��yB��P����2�HHR`�o_��yR�	�.�%զq���"7i�yb� ��ycG�f~��VF@��yb-��kO��`a@�+jm��څ�yR/	�s�(��m�<%z��� ���y"K�oDq��ن$�B��\��yҦ�>/�Ivd�!��|�m���y�!�	N�2�>����ԃM2�yb�4�����+e/��#�j� �y�eS�z�xї��Yx��qs^.�y҃���`w�:TQXU×FB�yb�&
h��7�L�44
D��#ϟ�y�ˎ��L���!(����$ʂ��yҫ�,q��, 5B�<�Z(�d�'�yB��>�捰��,[el��b+���y2_|#��;��E���$���7�y���P�4�` ��`x	jq���y�o�e���P#�_�"]��mQ��yB�6�.e0�b6,fְ�P�B;�yB���GI`�h�3+���fn��yB�Paޙ���M,ne��+�'�� �%���Q*��-c��p"
�'�H���ҬD6�A�2G��d�x	�'M���Q%d� ,���oz�]H�'�T�w��IU\�1�]l����'llu@���ܪMb�14�
�'�ڕ�CAI���x�Q��n���
�'׼{�%-Co�X���ߪr��tR�'���!D�GfHes���f���
�'th|Ya�^4]��P��OD-0����
�'Z�i�!��:`����R�2��u�	�'���Y��-%$v�� ��.�
���'b�hrˊ�M��LFs�v���'���SǤ�6\�Z� J�v�<(��'oZ�1T�~S�!ڵƛ6=�r���'*��QjQe��չ��< $�!�'��E҅&�HL�<p���$D�N��'l�Y��a�":�F��� 7��m���� :Lj�k
-N���FBeڡ��"O����ӊ ��Z��ZVxer"O~�7#}�n ����;N���"O*h��R��s�F
+  ĉ�"OD�pĄ�d6 djQƶq#�as2"O���eDR�R�`��%�`���*Op)��c�Љ2BEتwB�1r�'h�� ZZ����o�\��'��$�P��5�i�1Y���z�'*�x�X=�,	���
�n<r�'ZM�@Ok5� )�#w	n, �'��x��HR�9+�q
�s�'h�eyvF�@[��{���b*8��'3�����B��I�E�ġTn����'�2!0w@a��R.F�b�����'�l	�N����U�R%ĝhF���'��d�2fF$���r�<8�4��'��I���>����AH��.f�{�'zRH+ah�><M���c�.٠l��'���xo˗ �:�3���1^��j�'*r���A�x�Y���L�x�B�Z�'�Ҩ�Ǌ�9����a�	�u�@��'s=;���pA^[q��g��yy�'�Ȕ�6E<2���0	�fk�'�a�K�#AY��(��݂`Z����'L�p��KZ��Ga�"J
�'?����"��I�d`
�@���'?,����n�Ȫ��ͣ���'D!5bP���m��^�nDc�'h9���UB�-9V'�q�i1	�'`z�:wf�#d��O3p����'.v�z�B�.w���C��ry�#�'b ��nN�(�����W0:Bz��'�t���	9h���@�"D<< ��'^��k�8=w�Ȣ� 1�Du��'V�l�6%6-�8y�'��7,`J�'�)㠣�:�`�i�� ��%K�'�p-�`Cԗ7Ժ�[t��4�z<	�';�)�E枿��zC�فs�ā	�'U�A��8XB9�.W!!�<�p�'���j0�	/3��[�F
&�@�Z	�'�I�ː��*;2`Ѓ| f���'�$����=�z`SA�N�r���*�'�Pe�%{Ġ��W�	�'-b�'����QŎ�W��X�'��<H�I
�a�@@���I��0��',�YF�>��D9��=n01�'>����=�J}���� ;*��'�q{���\�(��	J�/�����'�f��:N�\ju&���}��'�zѴo;V���1��]cvq��'>T�w�K�b�� R �dlK�'�^I��̍�����diܔbR0��
�'8$ě��ͩbd~��k�$Q�<�
�'E��pݮ	+O:�^(st�%D��0����T\r|`��'f�H��'D�4X'fO��8���>M_*8�D�0D�Dq��4A�D13,�2((9�L0D�`�7��	�^���.^9,�	��-D���� ��U�ܜ{��^x�2�&+D�좁��~1�@�*Y����(D����AܜbĖ�ñ
� v�İ�#(D���C��$���% ��L<�Qf!D���M�!7sBE�d��S�N�w!�� ���IZ�S��`�(�"O�-�s"�]ǲ=*�CDz���*�"O��p@�B!F�"1rPC\�{L$�1"OĺCa-�~���B� l���"O����/�=;��v�Aq�h �"O�̃aO� �Dq3,܇n��,aR"OL)XF��1L�ڬ�0��9}y&K�"O<[�↿9����%�ݦi�ܛ"O�h�o@�)��saF�,����"OXx!���L���F4�\x��"Oh`6��]�D�p��{|M{�"O���6�Z;DDp쑠�rFi��"O ��rf�.�����!�-1�d�w"O�M�n_2���%�4a���"O�t�K���^9���Q�{T@�"Ov�
�W�zw�H�Ǆ�A^b�Q"O\����X�AX��fG�3zL�g"O���RNY�v-"��C�_���� 1"O\������DҘ�̖m�B��"O���0��Uʑ�5����]��"O��Z�ʌ;>¬Q��3�����|��'ݪ!0���&>�(C�I�"Y��	�'7�CCͳkj��H��T���'Hb��4Ãw��*�KϽn2���
�'�8ʱ·Z[j�ȷ�ƥQQN��
�'I�5�&B pH����ܾ]:n�
�'��9���t^09qWk��%d|t 
�'�����ɇ�,���I��
�3X�u����'�2���, x]����ao�qH
�'�Ru8���3�����ρ!F�Hk	�'߈� �@G\�8����z.j0k
�'ж��B�D����Tʋ A�L�	�'�.5��� 5����6�L#:�hЫ�'� q��Su�� �hX3Y*��'#���c��=
b�8"�܏+�.�!*ON���m��T葎_&�a��f�#;!�Dܘf�r|@�'�H��E;+�!�1o+�8���ļp�Q�cJ#QI!�@�y����5/:�ib�	L�!��JRd�sɕ�T,:]�]��!�K�,�:���+]6���!G�J�!�d
��,�0�b� Hߴ�V���!�d ��[qB��g��
�UM~!�Ė1��i�p��3��CJ�>_!�Z q�LQ�I�'/s������R!���v�)��GޭT��!gI��]�!���>���	��$[d6t�5�.3w!�
�}�v]�B,��oa�쐶�I�+I�y��I�?p�a�+I�5��`�TL��v8:˓�0?a��@���䁌fh����n�<��W5S��`ô(�0�s�<)ï�;`�t�P��Ǌ��u#�C�<�w�� u;V���cF^����A�<��G�iM<�"͋<@� x1��x�<1�n7�� v&��S�)�$�_�<��H�&�� ��͝n����iS�<�!�й�%/�7�F��r%�Z�<Y�	ӭ�F<��.ҙ�z- �l�Z�<Q
�B�Z���j�$d蝘aKQ�<�t�P�*�5���@�u�P��R��I�<���!<0����]�B��e����}�<�e�B���5��^�%�ڈb��	ҟxD{�����F�DIAY��HP@\�[(�E0�"O�LP7���RPcPN�<[ʕJT"O� @�i��R��馍�;:�r���"O���ő|H4����+g�~�#�"OB9QaQ�bw�`K�`
�$�$�"OR\�$&D�U7�sM�?���Sq"O|
 ��>҄u�뗯�TM@��'ў"~���fC�] ŮP
f����$ ��yb
�d���xݦQ��qĂ��yR �ϴe���D;F���o���y���7S����bH��zj` ��yr���E�lq*Ai�/��݉��H��y�'��^���ص��%|-�0�e/�yre�&y��Z�^
K��Q� ����yri��)��"���0���4���yң�,��(�k�-->�j�
��y�ö��<���ZD������y��S�_�t=3�k�>=�$���mK9�y���&����!SR�J�GN�y�KA�pY���H���޼q���yR��=[o���ƀ,�潀�T�hOp��Dc�̵�P%@JxqOƔ9!!���v<)��Ku��u �T�-!�$F�O�i�N~�.��Ƒ!�$�:2�3�Á�B�N����*!�D�'̂0
�` �%�|�p�&���!�hT�dyV�?8���R��B�~!�D�56��A ^�Z��-q%�� !� 7ՀT�Ug[��xI31��8t�!�ʑk�.����>`�-+�c�^�!��P�@��/H� 0;S��'R�!�$����ϋb	�A!2��>��|�P"ONp�D�Yl^��0-��d%
a"O�8j�B�*�9��é!ʨ�2�O<�(f�Ub���c��c�hr "�<����)05�p��zc�I����:f��B�	�FY��'i[�)�<��" Q^tB�I�qЮm�e��9�d݋qO^�~�<B�	)Jf�(2*��+��,��
�')�hC�	�4i��QC:y�,�1RLۘRC��f�t�rK�	�
�C��3c0C�
 Ԉ��7ƒ�1,� ˀ
đI����g��8� �5�` "��
������-D�d��KV�[�͖60ti�"J7D����lJ�~ب�%Ӿ(`]��(D�<0Q��T!<̃�O�.EkV���$D��$9c�x����$� y�5D D�8"t�I8<Q�&�M�d_�lH�n!D�[C�܅"�<L
4�E3C��(R�!D��2ЮY�*U{C#Ft�*�Р�9D�����	4r���a�� "�X��8D����GP�Q���JpMφA<�1�c"7D���1��#U��C!�K�#�� 0a3D�T��ÿQ�* ��+Id��PW�/D���&Ĭt�h!j�&?+�4���n-D�DA�ǳ/f� ��E�[-��j�O�=E���ٱ��l0`���	,���5(��=��Ie�� ��a����I+�c	#	Q*ؑ�1D���c����iCE%�8Pй)��0D��2�D�#�"]��<tِ)�2�+D��&���h���\�)j��q@&$D�б�	�fB�F�ڵ!��QF?D�x���Z?D�0B�[([�Z�#��)D�"Q&ǄU�f|�c��=*\�R�!D��ȰA:8��;3i�>��l`�=D�!"B�=<h:6%�#�N����?D�� � 'B�lZ �7�*1�c"O2���fF��n���"��"O>�"�Ù+�D=P���䨐92OJ��$��	���D�Т[w���'H#D�\jt�W�{l��F�M� R ��$�!D��1BX�����8�	�p�*D�@cԂ�"A�X;�6d�M)��,D���4�TULh1
%�����e�7D�H��!N��Ł�lR�v�R�5D�@�#��p��t9�#��yj�
�2�����@icwg�0Jf��`-�Rݺ���3LON���~ЭЁ��s��	�"OZ��W�ݧd�D� a���Vʴ�$"OV��Ff��m�� A�Q&lQ��+e"O��*0h��+�j$p�,F�8ā��"O�]a���i.LB��V�
`(�"Ob��4B��J�D�k��,j����'�� ��&<E�ި�'�0~Ė�9A�)D�|�gơi/z��jͬ*n]xpi(D�\A��ɝ)�ݳ�oI�BLq(��'D�4 r�ޅt\�щ��3DF--!��*�FiAg��<�����KֹK�!�$���R 9�	
$?<�R���K�!�$Cz�Yh�0�B�9-ܙ� �	V�O��Di!N��1�ty a���A(�M�����hO�')��ԛ���=G�ʉ�7ƅD F��ȓo���BN�SfE�e!�!9�Q�ȓ��񚤍ɬU� �(� �K���ȓW��pc4��	U�h�@����uv�y����"@
��q�T�c�z9��i�K�<�c�$W�L�׃��@x��_Eh<��aӵ��`"���.�Ň��y�����+4K�<�L�g�/�y��ޯH审�d&�7یMʦ�C-�ybD�,������0VB��Ƌ���yB�A���z�f��]����B�ӕ�y��P`m�����jg�A2j��y�AڠR�г���]:�1���Ө�y2�]�pJ�`��.��?�B�h��\��hO@�����}��(�O�*E�-+v�:�!�A�L��-yUI�gȌ��X�O!�$��j�yvIK6XZ�b'�\5^!�DQ*|3���$��Q~Q�̎sV!򄀓R�l,bӢ�d3�m��Rj�!�d�=1@�!q&�D��	@ˎO!�R0;��R����v�D9`�ErP�0$�"~�P@WN,b(��%�N2�P�\�y�*T�|�zEYD��	�.��y"��d���s�m���0���&��y��B�d^����³L� ��Q�Ǳ�yR`Ӱ/\��w�]�I� ,�D��Py�!�D�襢�R$'���Nl�<��I�4:Z����̤N.�ٸ����<�����(��GȈi�B�'��(ڲ,��-���Z��L�'6)�d�i����ȓ'z�u)Q��TI���J�*(��VO�;��W)mN>0&f�$�E�ȓD�:��'�wD9x�"#zrt��u�Tm���y���t/C�A?��ʓ<���� ��xh�JHN�hC�	�yb�a��d�"Pæ�yң�[Rf�D?�L[�/	-ml�|���,+(PڕM8D���A�E�����^�O>Z���K5D��r�2L��DP�I]S�2�I�h1D�� ������z�} R͙7!	�Ps"Ot�ccl��5�H�0�U9~��H)�"OH$�%��N�\y禔#G\���"O�b��ˑ,Q��À�C�-;�E� "O�m����;,��a�Fٌ
 Z��""O�4�u��Hǔ�єC��(�n]��Y>�X�'�E��U��,Ñ"����:D���$���|��y1O��]수 6D��Xw�=c��5�"gH2g�l][��3D�dHX�'2�t 4C�q	`��2a2D�8r����{1nQi�Z��QȖ�2D�\���[�P9,ت#�=/t��/D�h��aA�s�p��'+�s|�Ѫ1D����
�+AA5�7��3]�*���g.D�(��B4[ tJ��!#wd�)��+D�쩑I�,�x���j܌Y�<�r�)D�����R�>k��e��W� C��(�$9�O�Q��IP�K�}�tJbS�@z�@$D�D!U�u.�cO�T�؀��'D�P1B��q��eC��>|�Ԫ�,9D���ƍV%β⢯� j��8�,D�XP#��6N�4��[��Q��@4�y���6:쀀��¨cP�a����y��!Kb@��� T,�ɠ����y�IA�u��i�j�G��!� �+�yB�_(�ޡ����<���
���;�y�'j�v�+ �/����e���y�K��2����T�O1y����O���y�̭ل��2��H�D�b��yb/^�YdU�Z�F�P�1Gԩ�y����)Y���s��A0�๧AL%�yr��t��t�1/ۉ=U�5 ո�y�ג^����.rft+%��y��,"�@��R��e!ϖ�y�J3:T��ׅ�Q��TF�¹�y�`H�'�y{Չ�P��P�n�(�yb��.)�]�wD����5��� 8��>��OR0[geǤy���hßT��VR��'�ɧ(�B=��J���3%l٦v)<-Y�"OXU
�m�:8�0E,�;6]0"O�,�b�� R>�@t�G�P�fMj�Or���\�Jb�1n�%L~�Cd2D��# %Z�,�&t����r��l�Eb.D�pC&(�8o�2!�7�p=���f7|O>b���Wc��l��l�(+�hy��4D� �1#�@�~�`1d�	X�*�
�C(D�H!䝗���@ ��@��{�G%D����J[(	�,@��^�d�} צ"<O�ʓ����Hl~���C���JQȲv�!��¤4�0hY�dG�h$!�kڼA�!�$��]ib%���N%cJl�0k�6J�!�Z/|;d���ׯD7�mblĜ�!�
�UB�h��_�3���p�!�dS6��TY�D�97�d��!n�!�$�'���c#�)o�,@�s*C�P�ў�F�Ԏ�F�(�C���/x����&��8t'!�G�n��閔I����ҽi"!����-S4��C*̔+��˄�Z5!� ])�ia��O�R���d>^P��'�z}�� Q=��iI*êe��11�'ff8"��ݍ)�xi���Nk���'Ⱥd I070@PE��?{+��я�d5����H6C`"<�1�-��Q8� D�T��!
�$�:5;�֗Z��2�0D�� X�ɀX4\Z�ȗ`L,'Xh�C��'Z1O���F� m�H��[8T.^�i��';�I;Bب@���,(J��$���@C�	1 �<b".MVԅ�E�^� �C�	��|H%*�$+�H+�����B�>J�F��q�
� ~��w}��C�I�z��TAL;1�ԉ��V qԮC�	p��=p5�'t�|V�G�RM�v"O�@��뛹~���J������RR�\��	<{0N��p��L=fHK�K�pB�	�%��U��@�+(.<{Wl�+ݖB�5p���VĞ/�� kHmXB䉭^f8��$��Ԍ-�EH��(B�ɬ;thc��ݭo�YC��ǚg�XB�Ij� Ua�e���j�[E����%ru�a�0/U T�k��� ��u��Iv�dpx�h3�F�N`X�gKJ}�Xh�ȓ#ʎYq���>��Y�e��g����4��d�,3.@�D`�92]�T(�'��A��hY=f����Ȝs[��s�'AF���H~�\�)@C�=r�M8�'���*��P3a��`"d�1&R	ߓ��'���P�A�-^H8H�F����pܛ�'�Ru�u�U9lfYK�o������'6�N�:uP|�C ;i�x�(ߓȘ'I���(Ҿ0Z�=;'	�8���2�'�0�vb��0���'�=B�՘�']N��4$6S�V���*G	3U�<�
�'��U��gӓl��hx���w�-�	�'����	 @�v�� �����'���S(ؠY,�DV�q�~�:�'�6m�&]��	�K܍c�2X���y��
0'D��8T`�9@;��X��N+���0>�S�O�5
N4A�ͦM8�*d�X�<����)z$�'
A"	vq�U�V�<��ևc�Ųu�ŝOں,[3�VIx���'�|�;��܉>�ֵ+��%,~x��'��)KΌ�MH\<8�"�4� d��'�qR��_8'#���a5\֌�'���qMƭw��� J�����'0�q``eYTF�qB@O�_�h���'E ``�`Z�R�戠���Y���
�'���T�(u�}a�nAN�,�b
ϓ�O��aG�U�%�,0�H89�,�"O�9�e ��P�i���2�����"Od��Lę>fJ!kd,^	f4���d"O|	"k�4�
a�C�ܮy2��K�"O�|C�O�F�Y�u��1*��;�"OHQ���կsWּ	SG
E�i3�"OF��қn����&ƕq�"O��r�/�)����0�
 ��c�"O֍YuFK�G���L@�ڤ ��"Oj0s`��i��*_(n�l0AOn�!��|�|%@׌Հ4F%�D'D����Y��f�n��l<\��@K�<��nQyUś��Ap,�2�ǍI�<	�mµ'O�a��+�-�XQ�፟D�<�䃄�<C�ˆk=���1uy�)§=����0��z� ����U���)�'?�u��,\�.��U
}�4�3�'+���b��3Z���[Q� �qT����'��%Cv�DPz�#CM�U�����'��ܱS��ڊy�!a CҢ��ʓWF� ��Вi��D�^˦�F��3� ����?��2��>����'��	�T� ��堜0p ���]�RB�ɸ!����N�9[���XD�;oPB�ɐ8o�IP�LE�0F��!F�T�.gB�=��?q���U$$�eꍍq��9iv��_~!�dr5����+P�jI��zq
-l@!�?ܘ*���/��%��&!���5��]2ŉXteB���8�!�ȰA?�ڵ��pR`��'E�l�!�$:� ,��� @NV\�w��A2!��:I�0�Ca��v�eZY�Jm��'	��#&l��2�b��.�g��P�'�BDk��ؾ6���(g(�t
�' J���o�n�f�p�^&`�4E�	�'kx,ĥ�7ͺLHG��VD�	�ܘ'�FU�GbE3ks�UZ���?&H��'qH HVdW6d���
� ����D �'�`�;G�ŏ!�U�P�.7��@	�'��=ʤ�D�_�6�����$�6eH�'B<�g
�{��j��N�c��ԇȓy?��IwĜ&x6Q*�ŁW�����2o 	i�eO%u��{Gŋ	2Lq�ȓt�S��մj>�]��"����'�ў�|"�FթU��h��Ί�
���sh�|�<Y��X�h
 ���J��|��*
N�'qa�$䕘1�fiJ�+4ɦ�	U��-�y�O�f=�x�E�.~<`ᴪ͎�y����-�<`� �+ي�ł��hO��.�#�$1 %��87[`��V���*@��ȓ����вmL����j޴B�Z0��=��x"�)�3"�b�:W(�*�����s�j��fF�v3X�J#�A�8z�8'�PF{�����*ɔd�E3:2)Rb	���yҎT�����!A)5��
ra�%�y�O `!���c��{�LQ��!ӏ�y�� N�yC��)2|T�!	����+�S�O7�9'��&f���Yg�һ<�<)�ϓ�O��A�
�&ǯ��4=���|b�'�\0ʥ�E�V��+%�PI
PN>�L>���$�	J&6ai`FX:n�6My��{jC�	(l� Y�R�ݝX�|Pq�_(E�PC�I8�|�e�\�Gd*0H���W�LC�I�;\��q¨�t
^���D�_g(C�I�V��d�&� \�P��<�C�	{Dt� �[��݂'��{�B�I�X�:�h�,Ȕ]��0�@<%��B�	�(ޤL�ֿm��`c�J�RC�	�I��`S!M*'��
�.{A�B��@�H�I�'>|Ჽb�/ߪ��C�I�
�t��<j�� �(�kcVC�I�R�~��G&N�9�|�s7 �$7�C�>}ˢ�� [Z�*��ϿP���$/?�'I4̖�c!�
<"��y@$�Z�<�FKg�NT��j�=E���*�Ȋj�<���
�d *�b���2B8
G��M�<ђ̀�yD�&����j0'\`�<Ya�'kn����"b;(����؟���V��?����N�<A��dVf��Љ��/]Q^ey
�'�>h�&��.b蔒�ƴdL��H
�'9�����>�3ł"^����'[�S�,G� �D�k4�ؠX��`��'��0W�<��A�dH��C`̵)�'U�H�f&\�B蚴�H�Q����'����7�N�@��௄�Oe���N>�K>�,O"b>� <�p)@J�}8f�K� �Fа�"O��W'vm�1o�ThUJ "OX�H��k��H��?LK�� q�'��� ��!�,u;��9��B�1D��0���jz%���d��D�,D�xZ�#H.<m�N�e�O�B�I���1���
�ڜ2T̒�E�>�?1��?��4�V�gͦ����$)��,*�f
1�y��Ӓ*9v�{v�J-�f�����yR+�)el����΂Q���yD)[���'�ў�O��H���S�1����F��Q�''�dCD��Skdy����aޤ�
�'pQ���>)��ģc��J��=P�'P��(�5��H d/)Y�ĳ�'\� �h(6� �����RՂ�X��x�,ӽE��J'��{� m������y������� 
s|��^{�<av$؊6��АLܶ?��(2\_�<Y�KF/A��W��wQ��q�[_�<��
>X����W0	�J�ҁkLt�<1�I�(b�\ ��,-mm�"b�g�<y�h� ��]�j�o@� b7ɚY�<Y&Ƃ)&$�cV�_ d�@#�-�Y�<�KW(~���G�[�B����Y�<�o�#Z-"�.�1&L���Q_�<є*�0P�5���)E�}yB��W�<�ύ''���*Ϙ��.o�<��Z_%^@P���6�	�LTF�<q�-џ����`�TTL*a��V�<A"��u�����)^�7~��a�@^S�<i�ɇ:e\>A ��A�[�`��B�x�<a&�2�n��2'�ak$�'YH�<���	I<t��B3��S�^�<�#� M�BeFJ3[���C�	L]�<��g��'��-9���-
��|��B�R�<)��'?8�[vnN53��xkT �J��a���O���)85�"����9dQ�4K	�'7jM��@�<[�z��u@��\��`C��d O�X(���F�}j�*[�.���"O�����U4F��(�H��v�#�"O�qj��ջQ ��b�g�
�D�p"O^H��
@�.'����Lu8 �6"O�,��R~��R'O��9�d*LO���lE�2v����d�,iO�9#�"O��/H	4�|�2ԅ�.e�� "Oн�&f�V�`�j�0Y���A"O����P�d8a#�+�1~9%�"OH��h��YY��%\ �"OdP�]�n���Ģա
��W"O�Lb�.��4 �)�D�܃	���D"O�cI�3C�:Y��*�dȬ���"O��"^]�4 �JLS�ȹ�b"O>��/�-S�f��4I�+N؜�+�"O�I�"�CV��m`bA�"OB-�G�D l�!��J�h�"OZ��a�Q�A�<���m�	��݀�"O��붌0s�$0�g��7j�Z��"OJ@q�R
/T&ģ��uJrT�DD{��)N�i;f���g��ԵB��-H!���.�����:P$8��	�d(!�D��jJn�2��f�4��a��V�!�$
�#@���͛w���I�ǘ4F!��
e��u�qF�#�PԂAf��:B!�$B�U������)��H����[.!�� �)�W�+pYx!��6A��a"O�A��G��?��$�f��%=@1�"O�3��K����SE̴9
	3"OJ}�!nBm:��{���F�*D��È>�Г�$Ǫ��=K�(D�誡�R�[�	�����A���%D�|2!X#N��1t�K8'ɲ� #�d"�S�'xX�*Ѧ�e9��t@��v<9h�.P�h�X��;`�*�8T��@!
�6��h 䛔Q5C�f9D�HZ �A�=̖�0���'C��2��,D�d����U�<� �L� Yx`%+D�`�U�4.�$|Y��޹���B*D�(5O�Z�̨�cX�M�eZ�E)D��� ��"�`�u�Y%
q��(�&(D���,(��<��*
e��T`&ͺ�y"��Ȝ�2�m�g�$U�����y�n�%Yre�f��Y���t�4�y"JF(�0�Z5Q�[��(���y�k��7�D��D_�M�
T;�	�y���5w-Z$x���F�\(0S*�y�C�WK�y��f�>8�%�w�����O��=�}RAM�r)�}Xg�]&Q��HA�����II���O�����'i���PG�(=F�a�b"OL�jҩ���4��WK�a;
иS"O4�3���L}V���:0�y��"Oa��o�/t��ɫ��1r�֕	"O�.؄(C��� �:J�<�`�"Of�B���E|�P��O����(�"ON�9A��,,�d�� H�/S�1q�"O��
��Z r[x@vS��Q�"O�dɳ�Ƃ6��B���l��2"O��ƈ��n��Q���bq�&"O�6��l7���TfKD!6��g,D�~"�+T���jI��ɖ.�	A|T��d/?QC$��+ﮡ�Eԍq�;��B�<)2�Ԏ@2@�3u��	+��mW�UA�<�؃�,Y�n�/[�H���{�<���?_�8X��'�}%��X�FO�<����3`Ĺ�u��H�x��UH�<q ̘�>���(޼�l<�w��Z�<!�����ժ�I��=�.����B�<a���:{������R���%C{���0=�B�ы�$U�l��P�&�q�<�f�04�9�rd�^|2yi�V�<qDH]8xF:�7e>#~ܢׁ�O�<	WO�(X�9>'�dbPL�<�!j�(��)�,@4Y"����K�<�&UaӾ���BŚ&t���.Jh<��&|s6�SG�\�9�l����Dpm!�D7}�}�w�B�X���x�	�Tў��S�]G�y+��
�|����L�b��C�I�Qs2����[#>Q���r�K�xChB�ɱmyn����� ^��ɕ�\�:y�B�I�)m�� ��P�i݆|S���4v�C�ɠ~��d!> [�LA��J-:5�C�Iw'B�3�"C ��;���(XB�ɨj�4��FI�7���p�mƽd��B��=1�D�#��`E�s�B�s��B�I�/��r��Ю4��;6���FB�ɧ:���C�a�I�*��7\@B�I�]$�T�dƏ�f�C�凜
�B�I)мa�nԶ9 TR��B�10B�I9{�}��9N��3B��B�)� �ɓ#�bɜ��fY�\�.1����O\��$�"�v�BCƯM��I��P�#�!�$
��2)a���<I�t���4=!���9 Z�*0i��-؈D1�<b�!��3B���c�.�^�Qb��K:6�!�W/Z*T�:��N{=H]���?�!���&FTB/I6|0h��s�*=!�	?��ܢ�d u�nL+�%V�$,�'�ў��<i�cC �����i��߆P�!�d�(.���Q��L�fM�Xb4$��(�!�ĔM�f��p�ɿ0�D5� �ھNW!��3J��!��zè9Pv)��"�!��Q"AE�U2E�N�P���C�b̹�!�$�6EZ�$YC��0Oa�9�AG]�!���'��J��R�y5�,��"^�Z��O����!SE�ٴ� �|�:�f�G�!�dL�<a~��։9Rv��02�T�6�!���h�	���Ɲ s���b$�5}�!���-�lU�����Gp��1� H�!�S @�x"S'��W�رka�:YR!�$Zq
�8	FFF2w�riA 
ډQ@!�# J����[�;JX��qG��!�%�z<���a�dXE��q�!������ڲ�I�U�Q[g� y{!�Ⱥ~�6����H�T�y�ФE�!��!�1�g�B�@��Sb�w�!�d 5q$��i�����b-AwźR!�1V�*��嬊6g�r-밥��:!���r���
�l�tY��nI�]�O8��� f�Q;C��@�����I[!�D��/�V�ڡψY��T G��s�!��� ��򎃣	s��5��
�!�Qb�8
k�T�1�T�%�!�̖Hk�1�e���}Z��В+��T0!�K�t0���bO�DdJ �1%��|�!�$؆S��i��_�(P���Bc�{�!�T����f��*)9���r!�*G�!�D�mT�\�4͙<!1BH��:�!�$���a�A%ɳ$����44�!��܇W��H�1o3 �4	�ֺ}#!��	!�p#4'��Fp����)�}2Y��(��@�w�e˳&�U\xB���~�<� � ʪ0Igc� r%F<�T}���0=if)��:Ҟ��$���M"����a�<ie@�n��YX�ٰb�dy�č�T�<�T✰ݬu�#��2�Zy�RLM�<YSË}�Nȩ����h���Ks#�r�<Y[�Ƭ� �	�N�I�B׷P��B����4�E�H�Z�5�SE}�B�I<B�0},M^"S��b�ɛ�j�!�M�5�)j��� r����L�8u!�$׉@~�1�T>g�!��͚�Nt!�5R��)�pH@�h�taWc� X!��AF�Z��ѽxD�;�h��!����I����|^�0rK�Rp!�$U�`R��BZ�lh�L�3�!�A�|�X`&��
|<Z��'e�J�!�$ɪ����E�6Ǽh���sQ!�$���f U�a�n�{��(!��{	�Ѳ���N�>ʒ�.!��B4l��QA�-ՊTxL�u ڹ]!�$��On�#eF(xXbѓ�@@�!��]�;��)�O�svBCC�L�!���;\�1�w�� b� ���N�!�� M���H�cSXh���sl�d#"O���P)%�V�#��CNRj`��"O)K ��?�r�8sD��p���U"Ol��0��(�С�A���K`�0Q"O�ܺ6㏦Fܢ�#�'YN� �d"O����R/
-,�� �:򔰋4"O*d�m�V#��p� �t�ܐ�"O� �"�
].*<�sFΤS%h�:r"O�EජM�*r��-��K6��{�<�&��>x�P0jS��zzpP�S{�<Q�K��z`LH)P�:��t1W��Q�<�"O��lkF�[:db�'9:��	�'��%���U�S/���cZ-�=�	�'�����E�S��� &. `���'�H3�僣X��Q"�!�A�B�#�'�`�c���{B\u	VX�,��8��'��k�J�]�����&���'ڄ�B�F�X9��'�#� �I�'��a#�
"w�h�S� �����'��h8�� �6Ն���Ħ#��Ź�'���X�Mʦ$1��� q�r�'h�-h�D^������ؿU�=P�'��]��m׽:�6���ED�^�<�'>�M��E	 (�@� Q��(�Z��'�TT�W&P���(b�m �j��R�'� ��a�>��CG8,6�AK�''\0� �9⣒6����'���!��Cx�QA*ݛW�Y�'I��c`JHH}�x�nǞ��1	�'��@�iC�<T�밃M	0�C	�'oqK���6[�hS��X7�t�H�'���Aɑ9>�-�����Y�'�$��������;��P�����'�8S�$�O���{����uBxJ�'G�m�j� ��ޯ8�`���'m>h1Cb޽K/DуQ�ߨEX����'`���Ŕ/i"�	��E��u���'[�� ���+t�A��qBxղ�'tI4
		:��5�d+тe%�p �')�P�1��<�6���d;\`�'��rC��8|^B��E/_}�Ȼ�'C蝱�+T���`�B#m�X3�'�� A4l��8=Q*@㘣]a����'`�F�=����$���X�he��'���(/4ej���"^�d<��'ER� �聬$��\Ti�YK�])�'z4�p��/�P5�s�s��ail�<!�!t���&D�>NB� �)�!�ą=/ ����[�FVL���4�!��T*��Q��\)N8lar/��>o!򄌵H����+͈1D|�3^!��W:m����.Z�C�d$3q�R�!򄏽i��S@2I��Bnœlz!�$W8{�pia�ܨe��"��_!�đ�^�m"7gEX�D8���6g�!�Hq�Y�Ǭ�T�~�K���`<��_/��q5 �w�FL�a]R�Z݆�4��� ��7X�F���Ǔa��Ɇ�J�H��IN�^�Y�c韑^J�@��J��4�/הZ� d�j_�L�ȓ@ሀY7�%D��B��Dfx��ȓ3�M��N^�	Z|���Z ,���c��)���<sz��$al`dP�ȓ@�Z���Gƫ\�^uYo��nyn��S�? �� !���\J��K���S��pAc"Ox���\���Ӡ�3D2"O2jӊ6J�z�-I�m��z�"O^}+lN?'R��W��'�����"OYC����e�<-�*2����"OD%�e�P7yɚy��AF�uvd`�0"Oh��4(F~�$l�FbDko�P�"O��y��\�a�F��ժڤv^�D �"O�eS#�#%���ag)N[qX�+�"O�Ф��
��\bozϽ3���ȓo$�fDܚs��UǈU�ȓ�v0�rKR�M�x���ˊg, ��m�6E!a�60���b�8��{�R�w6rj��@M�����ȓ:�.PP��E��x'V}�����x�|@��ݶr������ i�Zфȓ=T��UӼ^�|P�4�#M**!�ȓ9���E��G�XI˗�Yl,5��/Q>��v<%;���Y�>`��d��8 Eo�3@B�r �	�(=��ȓl�|�:�fҴ$c^,a�M��0��8�ȓf�hA��&.��ࠗ�S�a�5��j�$"�H#Cv�� �۱B�$���V�Z�pc�$0�p�n/!=и��ul���(fSt9��G�v6�ȓu� ��M�8]d���a��/�ha��.�p9(v��)w���`��Z�ZQ��6�F���L����$�]:RȒ��ȓC<��ψ$'��8�כgB��ȓthv�[ BϒS� ���l��W�H �ȓZ0�A�D��p3�-�-3�6��UZ��&MH
{( ��*R�L�؇ȓ"T�$!D@	�7v���IY/A^x���?\CVEM�38(�Bq�E�[N����,zr�BӤ��j/p���V�G�B�	6h�u�o��V ��D�f�hC�,2����ɉ+�r��G�-#(�C�ɱE�@R�����Kf����C�I�E��°	[�C�E���L�w��B�I�����!GN3��-��ㄓU�vC�I�g������({?2� F���C�IHa��
צ��2�B��0�
#EV�C�əI��T����0����;�C�ɷn��Lj�R� �:��ڒ8QjB䉃[�,L�d�9G6��'K��ZB�I�`�(Т.Y.'�=p��X;rC�ɼw��b2D��Sq�:b��B䉀Y����e�I��̉�v��B�	@"���S	|nXɃ`ϸs��B䉙�	p!I�UN�Q�����B䉄 Ր3B�|d8��w#\ʤB䉛;dz��ć�Gd2gi�_�zB�I�k�<��	مp�8l �ؓ]�4C�	�l�KWJ��D-@��1=^!�d�(��4n"1���1��\Z!�D�8w7Z��q�¹�e0���d=!�((���c�0,�B�A�U,�Py��SbD�U�gθ�%L���y2�0xJJyy���*/����&ڥ�y� ��k@ ��A8O��y�L3�yr@�]n(��?2�(��'���yR'E0��M���-ب��DMց�yR��1Lr�zfaY���q���V��y"���� 3gm�	�\��-��y
� ���d��uѺ�2aK� ^�	�E"O��UfR+@L�x���;n��"Ox$qOJxp*F��[d|�Zb"OH�1Q�فm���`Ѩ]�j��e"O�ۢJ�qArEA�EH�`���"OBd�WEV�����E��Z�P"O��B%�ŇT'�9�$�����"OB�1��ĈM�&��p�M��`��"O޽�����{<Դj'ヂe�]��'���'�<ӓ/��N��J�U�xx�	�'�>Р �j�d`Yf�ՓnK�5*�����D�da̛{ZRLY��-�H�Ɔ�%�y���F'8��$�)O9��Qբ��M��#�S��M���N�",<��"��e^��	�f�C�<I�X+;��9Y���Xǒ�	Q�D�<	�'��|�ەJ��	��ڠ��tJ��_
�yb ���<�`!傔��möˆ��y2�߫y����#IS��33Lޝ��O#J�k͊V^�P$��g9�a	��^d�<Y�o�	�ܸs�!pR�с��b�<i���;�MSE�@�-N⬲r�@a�<�n_  4���S� �P� �JB��Y�<�b�0ZRea@"�b܉�	QO�<�r�����,�t[�,�fF�G�<�Djΐ1�r������h^2a�!�Z�<���ܤAi��[r�ͼy�Za���
Z�<�g�(A���#R@��`lZ�<ABG�r��Ы<( l{`dBW�<�/܍_Jh�ؒ��	#�1�SG,D��y��.y�U�ң�*T2l�b(D�(bǫN\����bI�W<Y`�&%D�`0qJƲ+��UY���`��%A�<�����%��%�$�n�[ ���lB�+_��LJ��%�>$�b�V�]TB�	�O�P�a�1j>>�Y�'Q:�\B�&�ԼB ާ�<p`��O6��C䉣f���p���;}Hd�V��/&B�I":�8R�9^����&�9>B��/m��$C�Cܸqd��'H�R#b��G{���掙C��KAYFr:��A�I��y"�C4W+%�/S�9��.
�<B�I/-�Qu�N!E��k��.,^�C䉑�d� �aR1i´��$�3z�B�-��T2�'�2<`f�g`�3m_�B�I3~��D��H����$JOp�$C�ɄVQ�*��6�q��4�,B��%�8и 	ր;�rܡ%`��B�	or���'C/o-���b�͋�b�ȅ� ��1<6@��5c׵m��C�1]x�������X�L�%N��C�o�|	�kA��C���aEvC�IzY��
�l�{t��	C�\�~B䉕t��U�D�	�n���o�hPT�'aў�?�1����$���S<?ʞ���L%D�*��E���Ye✠m��@P�a'D�����K7:nx!	�H��I�j	k �8D�̸Vm[�G`�t�u%��'�Z�xf7LO.㟤�6l9`L ��$,D�q��2D��hnWBZ�a9�
ɶ+� ��k/ғFO��ը�:�b�{��_�z�;��Z�'�ў�'KŨ��t�
���!�U�>���'gў"}�'��yJ�8�A�[~��r�W�'��x���/Q�Ѡ��HmԥsG@����� 5��>!Հ��n����ϝB�t�S��y�'XQ��S�? ���K��4m�p0�T��z 2�"O2I��(;X���l��B�)�U��}���Ƀ+wAvq����0��I/L4b� E{J|
dV|�ʡ��&@%��]�a�_�!�E/>j��G�A���8mʩ!��#<���!����
�	�@Z9�b}H�&V�[!��_:0�`�ӯ��`AfS\�Q�T��əQ�,݋��w�5�7���B�ɪ!b9�dg�
:|� e���c����и'&�'L�A�1*ߪM�`(B��� k�z��D�Y�O�x4�W#��1(�FѰò�Ҍ�DH<�a�ȧQ�x3c@�Jol����fy�X���<	��,��I^�M���|l��E���C�ɞ,��F�F2C���bG�ŽAdʓOn�b����ԎBC@J1s�J �-�� j��x2��3C躡+�:�U��R�$���d*,O�Ȃ�
I�J�Tq�J��&� ��'(���Ir��Zg!�xx~́�iB-��=�	�a�T�G���
�<��l
B�8=�=yܴ ��c��)�|*�
�Jf:Y:�(ҭ"NJ�Qp+Jq�<�"@�	�P����Q&y#P���'^d#=��	 1
�dpX{h"!{4�Ҙq�x0��D�>��8��)\�}��K�|�X�0C�	�lm�C��-O+�`@qW�:��8{9��I_}�*?��� |�X���+hO���g�%,JP���<O�I�*G�{-C!.�XC��p��'`Q�d�fލ����Z�]Sf�K��1D�l
ƙ�LCLpzp,��^�:8���$D���f��if$��w���e�.`qTn"D��Yl�c�<�8%	�B��}��B T��	Ԏ�(gbN�S� ����>A�����&deɠ�X,�����ST!�d� � $�FM����� Y��'�R��'��8��	p0(a@�
 ~�:5��K�=ђ�8�''"�
���0Ǆ���,�1Qa�4�'�6ܳ4d�R�3�JM�r
�y���MH����T�\��+�,J�f~�$���8D�`a\�v`ӴK-1S�M���2D�PP��Ӣ���y�L��
_8-��m>�d4�O����B�z�r鎆D���D�_���)�=h�q��g��?O�����1D�P"�$w��UI�H����W�0D���c��1h�S5쟩[c��ЧN/D�$�s��HVC���27�P�0�?D��#ѭB�:����/^�Lh�+D���kB>l}H�el�A#��3D�*D�x�b�<8�,Aᣧ�o��P�%@#D����������˫n��8ր D��(�j1 0c�$u �>���<�Ǔ:��8ۥ�����I$-�k`�������nZ>�D��l�;v�dq���$v�B��cd�y���?_
��2�2ɾ"?1�����R�m��Z�p���91"O �C��IuV��7g��]�"�'�1O�Y���H���pd�T�<�Z�a"O>�8�J�2;��p	�,Z5y�mP��i�ў"~nZ�;�,iD��tr؀E�]�2B�<G[jȹ���0�B��\�KEB�ɤҊ-FL�m�) �X��C�1_c�L:#M?NP�� 3�`m�7�<�������0�̤5�&� �8��V}�R�|�}
��ԣ��Cӥ��
3NEp�F�p�<�������
�|<�!x��TC�ӂ�)��(*~��*p��41%v(ʇ��aC�)� �Tq�1����N�x�V���"O����5��0˦�ҷ!��=00"O*��Bk��/p�,� �*�O����=���I/�:�(��W�`�|I��FLX��Z Z���u�ORWouf��9�Hۃ]�t�a"O��2�H���� HM0e�B,�a���+�(O�Ov.�v�J�mW�@3�fV!���x�'���3�_	x����dEa�'��]��ƃ%�$t��E�q4<��'R�)�a��1�x�P̞
9���{R�'e(���'Y�]�bU;� <+���'m �J���T��y�& .L��'#L�T��3�VY�h�. `k�'ў"~��&Ϫ����� uH�����x�<1S�R�jD@����Rb(26e^�<�c���5`T�ߴj�iKK\�<gj��[�
��ݴ.�d�q��KY�<)�ސ7�Pz��G����A2��@�<�ᧁ�O^^D�!��Y��I�JC�<�4�	��U�ʜ#�D2Ѭ�h�<Y��L�g�\AF'U/ʨ�Ȓ��Y�<��% �v��uE��h����k�<�V �^���*��'l0��R��g�<	͙2&Ci�/R;P��LY�ŀc�<��"	����s�%���t��n�a�<�7�]��zM�EÎ�x����`�<"j�y� Ps \�%��%�AŔ]�<'K�g��	�d%8�C��V�<	f��`�I���U,u������
G�<Q��Z�F<[��z`��cl�A�<Qco�u���[�fϏS�����{�<)� +�h��އ)zd���u�<�I�a�T���!f��
k�<Q�-�04�b�H�Ś7����l�<��W&5�%Qt�r�z�`t�<�Q�Xx���p���:��GF�m�<�S-^(f�x���Ȋa��<[�N�e�<��������hDN�	
Yȍ*a�V�<qP-�ak�AЅa17
�:�ǅZ�<��P*����A�@ µ �L�< �l�q�t�^ ^l��/@S�<!�*��h��ˋ�N`8���R�<y�o�"9��<!B��o��	��w�<��J�/�@L�!O�?��PKZp�<�jJ�Q�6H`�΋=����S�<fN6'��hpE�/av�3�oS�<)��՜6N�i	�J�z%��ˇJ�}*�(`"+F	EB��Y�J=�<���9�ұ�bTuΚ�B��E�<I�,C>"XH�Ȳ��=�tI���B�<�d�S>�(��F�SF�icG�|�<QG A�0��HU�G&p�.кF��|�<I�D�6&�:0g^(9��;�,{�<	U/ۢ�Ȑ eX�wKlx���\�<�u�M2rR���BN-	�⡙W�Y�<�A4�x�U��#T�D,�!��B�<��ؓ|3W�ԛ�Z�X�.f�<qt�Z�(~�	C��@�?����a_`�<	+�[z�����l��@�T�<����{]�uʀ�ҙ[H@��#M�<��&��H8Y�şaT������c�<�H btP<���˳6e�ܺp�T\�<��. -FHw/ׯ|��P��,MZ�<���.S�T�'E�+`�JҋUo�<q#m3'�tՒ�/ʡV�Lyۖ�_s�<� |��T
Q	�xi����T�&"O���I��I�T�P��j�����"O�qS��ޠ]��| �N�4c���xr"OZ1�FЅk��a
7Yl��aÖ"Oܨ��\�V�L�ڴ�F�8�4�:��'o��x%���L�a|Z	��у/��P!UK�O����D�h�j�	�����?Ѡ��!_��}B��ğ;1d1�H�r�<q�d�b��e���՛x�ĩ[��Dܓd��5��B�$Ut�����1@��f�F�(^H=��?k!�D�!"�a�d�M,2N��鱭@>Q\0r�,�$L@�̖'�LiE�,Oj]�!���|�'��l a+�"O�t�G��?�B���>Gv�@ۤ�ʗz�9�ӪźY�D��	�3�B͈� Ԏ]T�b�
�{����$W�V��}Ȳc�(o�6-��r�r�X%dt�J!����,m�!�$�=���PE�DN�S>y�qO��9!���We���Gl'ҧ\� B�(�|�{�*�o9�ЇȓF�p��G8���˰�]�L(tKV�x�@I��^�p�<y�OL�<mͣ'9W���|�<a��F<�z���^1':�a�1F�h��7N��i7�c��'�rQ�fJ�S�H?/bP��`�]0�G(���$��X�(�e�o��x��G͒R�!�$�9J��h��Z�]�e��
�O�ģwa�(r��#~J�S:*�L,3��Ҥe6�h�Ϛ}�<)2,׌P)Fi*@hR����$#�Q�<ae%|� �)�!WZ����XM�<��Ơ7��B$	ɆP� �c��K�<���@34��Ǯ�d��xq&�A�<�/	!^d��2J�"���(��T�<�� 2�.�h��mN<�h���P�<���R�wZ��Ӄ���U f�VY�<�#%�QJ�sg"ΓQ%�@�A�C�<�$�Г�̹Qa�J�t�d x�<A!튑_ar=(d�0r����p��]�<�-Ƿ^E,�c�OƲ@��Ir�R|�<��%��0T%A�&�-zHq4J�E�<�口�h���&�<�ty���Vh�<)'K��Fn�⬛�il�Cc�<0`�v�����H�z!{v�%��IN�,_
)s"�@E	�h��ȓuc����A�|kn����
H�h��IfV1 (�ntRL[2`�-�q��x�\({TNƈ(@��{f�ݤ#\���+�����MF�I�(�e�4wν�ȓR֠��5�4m��S#�5씁�ȓ��+R�J ơ;'"N
����;�dR��F5@
D�+U'؀-����ȓ�b�W�U�]˅ ƪ�]��$)9Qbk;U%\1���'l��ȓ>��]�wj[�w�"�J�@)7��t���⑚r��%6ܙ"A�O!����I�r�d !�O��D�>]�blc��%@Xt�e"O��X1NF�1���I%��8��P��$N`)}3#E��h�~b	Z:7�0m
&�hr'"O����MZ��$XF�[��U/X�iܬE��+�~Ҍ�-��bߖ� ����y�O4	�<@A�6c侴R�-�'��x���9j�D��P��7�<�E��gM�����8���RC*�^w��Y�D[�i�L�'���'$�N]�tb] �v��􍟛z�LY��	��~���m_y�@Mc��,%�����?|�t�� NN--(�",_�p��Y��`�<���͖	���KR+P�9�~����q��֠ipX� &aV�gr���b!WtH��	�������l͏1ǲ<�f��{�p�*P�޸����I�3Ġ�4��()7b����B%9������I{┺2C��	h&@�ӊ)�E�-5�|���D?d�)��ףd��G���Axeba��:�K"#`��6γy
�0A�N�H�P	A�-l��30�����d�� (z���,Oq?%��$���Lc��\�s��<X����b^џ�[�O/'�pU���	z��]a3ez�? |{���q�N�
S
�7BPqB��2A��8I��E�2���S�w:�9�~�'m�hE$WR�Y0rI)�RtA.OX]��A�&G�,�*�!�e�t)j�b>�)wd��_D�����6�"��B�T�sC*��� �*m�`SSl2LO`=��[�	zb@*fN�0�����n� -f��� '��i��x�)O���H��I��Ӝ~��Be?L�e�VgX*�����
38J|���G�<F�	���C�]H��9�)D�j"�A'���(��U�ڝe�V�ʖ�t���(X@���ؔ��4�r�eƿW�� b���r������N%[#��Q�j�����Y&\p��KX���0����0��)K�3�4��I�	wߐq�'��Ӳ��O*ܠE���ތ�"�h�v�zPZ��kc�J�,�E�u��+=z1ꇧ@�2�@�|�e�D�K" �a�)-���^?Q2�	�H�6PA��.LO:�������!Q�і{6��q��K"�8��
}�#
Dv1�e��J�Fs2��bSp"Pı�.�'��|�∉@ء��8�D0!�eZw��E�B75nA���D!X���g��\�$hk3A��[�H,�E;��|*��!^|�Ȩ��"{)�Уix�̰�o�#}5��cG�P��cH�lb�)�F�^W,AT��$:��C�$`�rA8�fB���4X�N�*�l�O�<@��Y%(�f\*&��Rn"<���T.�<5����G^��eJd��9�y2�1��h��%�v���G�_p�C��HG�>T��=��F��O@���I3W;*Q��/Y@dm�c"O�u�5��k%�0���6F.(JӸi�R�D�����|$;�)�#��`#J�3���$[�Pk朱�'��a�LȻ3�<a�SH/���c�',�t��M���!(c���J�x���'R���jƤ	ZE�bΙ08� ��'���ꆋ�t��rrDF�4ǂ �'Y`	���=ގ�H��%V�c	�'@} '�T�~*�y7�Q�b�5��'�*fJ Q��΅8dB4�&[+�?���4|�T�K>E�$�W�J��CE�)i�p��[��!�D�I ؈�4sS��B���W��	�	����R�)�y��H.m�ʕ�v�U}�b�pHɜ�p>�5,B�&t����ۍ],�s��S���<1��G<5�����B�9V\�~�L(8��SE K�׬u ���(O�Q�f�-2��c�Ҥ}ȟ��2��%VFt� a�.m�H��'�lAB%g�S�O����TK���(��G��#V܉��ݯN��(�;~�h%{��#~���0�8��� >�4qJ���T�x�	�*�p=���[9��y��ʶl��(�d�S�~��������@��4����V�'�� ٔ*�x���c �6�Ι�� Y-���R�J8�ثf�J8$��H0,��['F�X&��.�$k1&�Dص�
f����+�	�5N�ʧ<���;�L��&d�(��cHX7��GyRع8��kDL%n�� ���	_��Y; o�Vr�Ma��X�}h�럶�B�I�>E���D-p�Qb��H�O��I�B׺"�8���B�<@
` �ň��Q4��0�J�	mr!�_��~�GG�z\�}���K��x9RR�R��$k�({jTtR�j�'�(]+E�N3d�*��ǆE�q�B�g?��ޚ�ܥjA4I�x9v���i�}r@�ˌR�@��P�H��בb�I�$O�-F��ex��]4z����@�I���r��O�ٛ���d�'�c��.3�U�d��a�i1M��:Y$l��l���<a��!8\,d��'ldCU͔$k;�`��z¾�:�V/W�FA��C�}N�ťO����G����?��AM�&��6�H��`�*�H�\��d�:�h�>qpIL�DM��F�4s���*o]��/p�D�#�_}b��~l�k��'>�u���= D^13���5툩#K��J�
/Mg�{g�I�;c���hߴo����k�����!eZ�R�D��ȓc����F�f�����P2�8@F�N�$G"�|DK��L>Q�%��R��t,X*�hf�~(<�Bfá~yL�(ą�(�\jU�9�4�WG�QEX��[*�T�rp$�.�\M;� �
��x�JA���3UmPB~���a�΅:f�!�z��ǩ� �yb��0_ @`�E��5b��4��	�9	�S�[�h��K	n���~�� $��q�p�֢CS�	KF�u�<	`Ñ�`�um�Qk���� ��2�$FS�<�1���/r
 4�~�K�p�0��6Ch�a��
.,9���!4����m��5�B��Eغ{���'��:i��/��@�.)m�����'�p����c��0��+��f��%��h��풅�=3�d�C�*�E��ҡ�Y]P��F���)Id�J���=� �T���ٗM�����e[//,����;��M�ĬZ\_��Ғ���*�\���]*M$RSBO
K� 8P��c�!�䐜~c �7e$J����@Oٚ>��$9*8m�F^�x������>2L������7w�d�!�K����q��T.'@!��/�(�B�EE3���{��>D_�����C.SD$���q�����~z�C0��-X<�Qgңf-��	�5�h��DC��x�薠� m�6I�,�%/��q�,or$��I��h�"@��0=�ox���d�-ф�P�YD�' �M��&�jt��{$�/֐�(� X+kYP�F��*���`�dЎ���j�f/T��b������z�jA2V�62Bm�(���!�)���u�� �ιA-���b>�]&L��4�֋
�.�=H���f"OL���A�H8)�Pe# m�퀠M��[��PdҢQ�Rr�Y����O65�0��3M)�����
R�������4��{��;�Q�-Y�N.�Y�COT�%��%� E��x�ȱ��o^�@�k�
��W��'�'�(�b ��)�aJ�6|�����=�vl��&)��s&��o����!m��e�"�yB&Z���#R��Y��"O葉�h�w�M��$[���0��/ޘ}��\� �[}H�}��,MY�왙�(�Fܧ�y�)D�q&��㔟
��(u#���y�M �<��|*!f��v�[O���?��L�n�9 �*7lOf�@�B�Y�01�`��C��-���'��xTkX0J�n�l��D���*�ř!Cz-z�,T�&C�� Hn.B5�S�Q�\ !�Pۂ=���7��#p	�C��>����l�T� � �er�B��=D��'��:V��!�)_�g��T#�p�"�K�HXb�)��<锭ڟ@*L���$M!O�L���Q�<B� �+T�� �a��	��`�N?Q�J]�
���č�V��`�M�#����,O"!���6_�*�QW�1֌<�a��?S�!�$X�1I��So�4x�xٲ����!�D�'��Y`�i $��
�kY�!��<�-;���5
��ѡ@O2�!��R&XH���E
	��`2AMϸs�!�8zw��*��7�|X��,ɬG9!�� :��	�%
(]���䁞!�$L�,��!�d(Ɇo�P�hU�}!�W�JLb��s��/I^��Q/�(!�Ď�UJ����'K9�t�PK�$!���i��=�'�L�Q��1p�
�!�d�>���gGG��Hkf�G�s!�ˍ#E�u.�)��+S�+�'��Ż��R=T)�)�� 'B�K�'�8�pL4{Đ��K]�o��'T�� g�&"㾕��ړ�6A)�'��}�W�4J� B�5�n��'5��9�N���%X2㐊!�T��'W<�R'a�6����c׻(�����';
ǭ�9Hh�p�ϧ!�C�'��y��?lo�!c C1�VD;
�'t8�I��}��o�9���`�'�� ��_�¸�u��F��PA�'���:gj
�5��̻��K16[\���'tZ��L�8��h�U=pq�p�'Zs��F�:x�Si�0t� Y�'cz�c�� ��B����9�� �'�ld�$I�$s��Q�6-�fD�
�'�pɊ@B��]����+v���'�Ƅ�#��>���g�DQlM1�'yh\Q�E
�.��U@�����D��'�ѣ�D>C�����B��L��	�'�X�2�D"�,���%D;�I@�'�\��Q"�-�ʰ�b灹��1��'v�E�� �>���h3ŗ��|A1�'��XS�-Ɏ?` u�rM��|�:���'溸�U*O" ������āNp
��� J��bN�+D��CeG�+f>�"OD�#"��&h�<��tb�';Q�4�e"O��J��Y���{�]4MDft��"OZ�PD��n]"���`�)bM[ "O,���2XnH��ϝA��;&"Of�	�$^;xJR!�MU�5Q���"O�}xǅ��߾��#ػ#�E��"O��)b�"H0 ��+��-ƙ�f"Ob�I77�	I�I+JoD�*�'��aS��5�a|B�σ/�v�Y[��B��6䦱Pۓ;A�e��&�5h��D��(=�e{�"@>e+>��!�Fk!�ы~��h��%Z�(�G��pNqO
�C.��$�P�s�d;ҧQ|Z�(�E��,g܅�/WKN��_� e����>0^%t�7hX�(��N�$�a�#S�hi��<)��0"�
��v@��Z��iHb��J�<1tk��"��q��O�Z��ě���C��z��4:���U�'���!ɕ88�ҽ�0b��dŪדuj6�84�@._��!J�4�AY�����H1@g$�'M��]�ȓ��1��KA�;� 㩋5d̌�=�%��j^�5lY'�H��u:EBC�{�ꙸ��
aS6\xw"O>�H �R��	��;@f.�@�Ҏ�Xa�j`yB��L����%|���@�|��9���1!�$A-��
a��PX{6%#�`�ҋ�!!t��'I�u؞`@��K>J��0��K�j�,����<lOx!���$������@�)A"�3=�!�p	�!3ttȆ�l 1s�@ӷ/�9�P�]�!��P�?����"j���<F�6Y["L�3"��6��L�!�$'OeX � ���I����Y�!�D�H�`�c�'(zr�$�˥�!�$	;1l�@Pr�&3�-�0�׉\�!�pi���@+ݾ<�:��L7N�!��,\I��[@��=x
���BL�!�DZ<9��(B$R���_s!򄁸z��� �.�ib�Q���O�}L!��O�{3T���O��8A�=��Y�!��� ~�����j)n��D] w�!�d08�'dO�u�aJr,�\!�БZĲЋ�g�$rn����sC!�,ޙ��ʔ$�����gÚ!�!�䂴ulȘQu��/
�>l���6�!�dC� �Z��W�T��]k!gH"'!�D�+%���S�[�R��@'S�0+!�N[��i�E��O�Z�q�Ï!��6\�M��ǴsK�t��h]�A!�W� +|� B	[�M8v9��G�u!�B�DFU�3B8g��h��ۆ^!�$��hA�Ā�=%�d+r��E8!�dԽ�����7BW��X�*�q!�$�1�Tz��I�Ul���R��!��K#o�.�Q���`^�!��Ǵl�!���`>����.eAdz����!���,�B)"1ի	E��D˞8�!��I&0� ���혷(1���H�4�!�d�(,�L� ��+L��w
ӥl�!�$N(5�Lt+�!3�������!�D�t5J��pN2��B��k�!��F�틆��:X>J���*2n�!򄞘-�5�EF�L�l�A�Ɍ	q��{"��U�Ȑ �9OB���� (��j��َ~�`<b!"O=H�e_cmȤc��X�>� �����:�������h�����/&E2`r�ɉQ��8�"O�&��8fƝ;�Ww4�1�Ɋ bU��3&�yy��g����*K����B�
@�pU�Q(ȸ p����P�0�)��0�.V�P��W�	C��C G��,*�Q�M�r����� ʽ	���7s�� @@�X�0�.�)��<��ة2�$�	��~R�`��Ui
y���6@�p���L�����?c�\E�vm0�Oy3��0k���I�E--F��V@�WN���o��~"�L67��
�Y�xT�4�2�O���ϵ~p��0���a���~�ּ@�z�'�ʼ"��2����.����Mӽj�P��wa��;�v��w�FF�(�æ�T�z�јs�O�$"�u�gy��J�Iн�S&��CI��!C\��[�A�gH�?��Ɠw�ꌡ�0�9<B,�{��2��[2���h�*��c��"qX8@��P;&����dش�R\h�[
"�Th��LW95��E�I�D���p�Ķ}�j���~Ba�Q
m���*��P2jX1���S .��$���'M�tA�b(�O�$�,�/rr������&2�"-�1�*t��B�����?1��R0r�R�.rt����ɿ>��ԻB�I�!�v�N��E�&�2��q�џh�!��:4�5���'z�IB�(��n$�G̒����$�rPzT'F3��9�)�:��	��d,���-�d�nP��l��1�4TGN��'�<�AN��K�O�ݺ��ݣ|����������3�Ƣw����E�~r��"2��4]x��|`��]�P�JQ۷�!/Lv��e��<�j�xq�9���#X�b>⒄�	!]�lp��]�sKP�qC@��H1[P��1q��Bቹ$�H�Xb������g�xh
g�D�$��$�<��ܫ ��8�*�j+���|�����.�
y���Zjk��6�Hi؟9��e�8��@���?|v�����zY��cT��{(<�t�tC�*X6Kq�^R�'!�5�LU�'b���QP!d��+¡|��ʠ�B�	,b��a�ՎQ$����LW <B�	"7��[�+�=rN�B�(���C�ID؍�Ħ�#�(��`�+u�\C�	�#1V��c�r\zp �M'K�C�	f�P�P��?�T�3ץ�-s�C䉜'R¨[�J�<@Y�Ujv��B�I2TBhh*Ѝ�f�Up�cª^��B��!o�:mS'��zP�@�ku"O��$�K�>�>����Ӵ?�����"O���ի�G^�Ǘ�x�Z�a�"OVy	��k>�,����,;,89��'����M�|�ɧ����M7*��H�c`��~3�M?D�\ALմS٬H񧡔N�j��ñ>�F�ʾ��d�t <OJic�"9$�ད5��|;`�q��'G���U&M&Qݔ�X��_�T�� YK�-�̋fA�T��=YEO(�OQ�k�	!��}CR��-<భS��I:W]y�+B%��mk!�,=��Su]R}pW�U�a	<@e���ir��Uv7X��{��)��^Ut�b
� N7��H��4N�>���G/p�X8��C��G��\�4��n��?�Ҽ~�Ҩ�#�H'����4	c}��@�(�D�'��$�bGծKu	E)�Q숣�	̃,tP������V��)�p�:���O�!�%ϻ<��,ࢄ�1 D�a��>S�(��C"Q8�p>�����B��� )�ԥs�F���x���/1�@����\9"o.I�'`��Z#��vB�T�O�������^�� #0Tt�2�<Q����@hF�[��0s@��W��lѫ6�U���4=c�\:5ڮ��R��_6,��U�K�"~�I3&Z�Q����Ш�S�F� �P4k�嘤jVP|��M�8�vX���s��?�t T
��(yP���FQV�P �CB?�5�I�D����*%LOV��m&�Q��Ğ2��I�^��N��F�^�hI�]cj���m{���$�yGT��wm@(Th���憜'�#�9o��ū�8�O�ͻ$��1nmj��Q�D�T���H-#�U��#B�{!LQ?I�/
��@�@��^�
c�#+ʡ�!"��"Ƃ�y����*%F��p������( L��P���!F�,[� ��TN��Xh��\�D�<К��O���Q�>�+��=���>�$A%hX{G� 5uy�QرD۷3�1O�Yȑ[7����:����O���V���0� �A��V��C�4��0h h��DN��t�"C�6��e�̕$>��heA0}��Y*Lp,��j`�''7^Q ��k�B4�w��0/�
Q'n�jݠ�c�"O��CIA�qo��@�n�I�`���� �9��&�b隥�0�3�dɽi$��P��%yx)�$�8(A�𤞵b��������I#�2$YJ����"M�t		�EC��(�D�!2Bv��c����x�'ă%8V$ё�M~R�]�5���a� 46y�Q�e�yRۨ�s����J�#	���	+u,^%�{�R*�5yLZ��~BpM��G�T�˃��9�ԋ���n�<��
�N���Bᎂ���K�)8�B���,�<x�H�f����~
J�� �)aƝ��l0��;�H�1O�42���n��q�i�+Q�&�ab��#B�
E��!�l�*��$t���D@�l�Б�1 �L`M:�hF�[8�~2d����3�m�y�5h2'$?�e���G�~���'ڃ'q�I���'�� �2@GLM��V�ً�K,	l�p`N�������?��$��KHI�(h�  �x�Х�-�yb/�5Kaj�FY�2 y�P ��~r�O�5���q	��|,p��-Z�3��\E�$��H4�BAD�D�9�@ʜ�y�C��L��ە��8��I��BQ16;X��do��X���c���	$ 5SK?91r�V�K����N�a�,�	Q�1BA�~b,��_}6y2�E�75���y$.]��$hC��EQ�d{�
�A���
���B�����\�_,�!� �2#�D�o!ʓ��BܣY#���BU� �x�����}*������!\&��bCS�B]\�B�.#D����%��)�`���L�8q���0˺zZ�1�b��^�ք�G�,y���'� ,�b>睴n0͉p�R�lv��@3�1u��B�ɧcTZ�1�hj�+#�)q�|L:�)vrs��*-f�B��Ʀ�b�g#2��yҭ��S��Qŝ"qX�g�X��=�QGE�|<�Ua�ME Pݘ ꊉX׸ ���"whr�ѡQ����m˳-}v$zӓ\4T�gsS���-�0<[��?և��e�p�2V����X��CZ�c}��Y/���9Ѓ�pG̕���v����ы9D���aD]xX��#��-����T�L�y�w`ŋL3�a�2̋)�LɲA݄��O����%A�
i�TOz���1�!�D�>y�(�����^*F�r�N��
�b)�<��(���o؞�r��R/<,L-�%� &�Y��(|O~`�b�� ���bشWd��Q�[5A6�,����=ǀ%��
c��c%ƥ<
>]x�"��|�i�?��/�Nȴ�*ҧP �Cq/'\�
�\
e�%�ȓJ(t�$O�N�(ɔ�D?Nʄ����/I7�\I>E��'��i�AH,=x1Q�F!]�hM��'?���D��-�X�*Jix�8�'y�e9�(�R��`�ݱ?��P�urAT�;��:D�ث�	�#ႌ��Yv���B�8D�x�%.���V%�`��?T)cl4D�cKύ @���m�99�U��	)D��b�蚬ѪX� �E�ʙ��!'D�`i�k	 :~\)�7��;/&HA���&D��aਃ�5���)N���`��@(D�Գ�e�;Zn��ʂ�n`�v�)D� K�O�-XvTh�k��;L��3�%D�\��L�)*�Z�zU.�,k�VۗB6D���+��+"�q�
�f,>5��0D�P�Ä�0\x8ՀG\�k7}1��1D�`6dW����{���,��<�*D�����A�$�k�-��2�xIbc)D�4�w���14�K��V�=ӞĊ��8D�@�W�S`b��'d�נ䀤6D�Tr�ȃnp�cE�dШ<[6�5D�\�鑀Px�����T%"=�ܚf`0D������!$���3S�26f޸��-D�ȉ��AX)�m�0Nn��+D��$f��>�1t�ӐL�`5`��2D��e�����%C�Ռ}��W&/D��x�Y��Lju�Ъ?��pj9D�����T }��l@(Nh�Xq�H4D� ��C�S]��[���4��ؖo8�	�;���f�ف5-A%��<R��b����Ŋ�d~\�	�?������3D�dI4��&_| &� ~�d��R�6D��QBֆ8��6��4�6��6D��9�)�9;��y/D�e�hHS�g3D������z�Z)iP��� ?f��2D���a	7y��. �<[�B��?�!���<���s��|m��b0lݎo!�Ю"�t|�5�N�B���e
 �ON%Fx�nv�z��."��iRt��/�(��w��O��$!��??)��T�2�@�ARL?�� ��x�E�	K*��㨈[�ְ�w?O&�����	1����EH�<E�TGΛDg��x#���	�SJY(t�Ad��7��	Z����S(���sw��$,d;�C=7K<a��M�wZ�zo��g�T>-8�Lޱ`lX�Ʈ�(V�P���S��'�T���2�s��s�04���'JN���o�*a�(C "O��r#�-xit���ֿ%ͺ��"O���l��-{<h8��'\"80�p"O���0Y�S1� E�_ ��"O�a�V�2V�
I��MR�1Ʃ85"O�T�q�'�*GJ��%t� `�'ϦəC�0M��� xj���'E��s�*�|}>cĉB?~`����'b�q9ɛ��Tb��|��գ�'ð��A&�\������x��`{�'H8����b���T4_��|�
�'C�eX,�wK�H�DT�Q����
�'����'B"%�2|���W14�|�	�'�~���΅C7�i�R��%}��h	�'\���_�.�
�+��Y�]Z ��'�R�Ae��5d��tǀ�� ��U�'Qnت0
�S��Z�#�0|.H��'^�!����t(��*���y2⚯y���u���*�c���yB�ݙ[C4�!�A�+^6L�B�!�y�Nʧ@�*1����)�.	�s�ؚ�y�R�C
���,(�d9v`�y��,~h�#lZ�$\iUo�y ՐB���;/�
���t*P�y���uU%t/��Xf��wJ��y�D	,E}>��w��>��`D`Ӹ�yM�VO$es�4FZ^=1O��yNθWf�����'k�E����yBh�	&:1;`�S�"�1͘��y��-|L̈�QB-L�)9�͎��yrC�;: h!��u����'L@��y�`�b?�p�§#�Rб�Y��y��(.��[W��-_"h��gN��y�#��jte8g�*ܠ����yI�`�����J$V�(|w��yb��>���GC+J�Z�ef�x�<IuD�}o���B�!��9%�BE�<��GV,l�BU�1���ȡ�h�<�䥀R����r�ؒQ����P�Z�<1�����ȅS����"HM~�<q�ǋLȅ�gIT�(Ԡ8v��}�<�@�'������2� �GKA^�<9'�`)R]�DM
�Y���E�\�<�4��V[��r�eC8��D�W�<Y��p�!�m�lu�a�&�ES�<)u@[
�j$⵪ڽUD��0�H	D�<!bb�-Sp��PL:�@�&��T�<�1��,.�MhGd5m�0�3�T�<���,E'�X�A�0:���ٚz�<�!��9L�d�ROE�yz>���P�<��M�=1���S�
�5u�PU��M�<�gAʮ#t��J5�ʴy��M�%�MQ�<Q�B�A)�bѬN�k��X�<Y�G	�h����tH^&{a�آ"��x�<AD�]%W=VT��B��N�N�*e��v�<1c�6�� j����J�b�iE �s�<9U�7����n��_F-�3F�j�<AgG"_"�h ����t�i�<�nPrP���ÿ/��6(�l�<y���/����ed\�m,h�)���n�<� ��"GÓZ\b٨��E�	�d"Oj�"���|�h���{��%��"O��6�J�7^��C��(	t�˥"O��j���6aF�A��lY�+6D�"O��
gA��q��I�Q���4"O<��bA���t���V-6',���"O�y�`�@�����!ڴ��"OZ�	b	�_c@�5b�7f�̍��"OJIs� ���x)�/z�쩨'"O I��h�t؀� �H(�0f"O��r@��f)90���tX0�"Or��T��=!c6y��H�\�r"O�\2F��	UC��9ԃ��}����"O.��e]�9��-�$b��!��"O� 2 B�.�.��G��%u��R�"O|H#G�K�e&�Yv!�,o�aC"O�!wJB�R��J�E+n`���e"O^�B�(RK#�9 �{���"O�i���O�{"�"�[���(G"OaP�iS=`����R��qs~��c"O�#��S9D���i�D]�F^�]��"O��Qw�"wq�]��eC O^�`A"O*�����=T��p��/|5ʼ�"O��2���4nX>m��jW�.���"O�It$ڑ8��y�1��.�	"OT=0��F�'^��ko8]0	�"O��S�!zv���G�Lu"Ot`����OeZ���ʁ=�A�&"O���愘/�. ��^��(��"O� �'�k%��� �' ��8"O �����w��\Su&�+iA\�"O��h��:?p � �c�F��#"O�yТS�B�pІ�J�Vv��"O�M(1&�(
G�aA�@��IB���"O����A�(=���P��1A.�dQs"O���ugSG<t�R	�%*δ(�"On�7I�B���7��?B�3"OV�J�l� ;�8���\�n��yR�Ւ&�4�)�����8�w+؁�yB�C�xy"��W�$73"�3�!8�yc��*WeAccH�ѕ#E��yR��5f5dc�I�Y8VQ��K�y�G��0a�ir����` $1C���y&] �|XP�_4/����Hſ�yR�Ơ7��=����>Y��'��/�yR�4	�e�����9t����@ݒ�yO]�5�̅1�*H�Y��}�1���yb�
�sA(5I�OɩZ�Ua�͢�yb��1Vh�p��R�V�����l3�yҢ�U�B��,�,MN �MF�y�O[1m��yw@�q���N��yr���n)IB��e���+F#N��y���8)���+�W<\L+�@��y��(n4p�	دQ�0�dÂ��y���j^&yG�ԚCg@��f��y�'P QB�҆D�g��@3�M/�y"��nJ�A����+U%���҉�y�	8tAVёw�$S�"8��IV��yҊ�9�V��ȃ:HC�u� M#�y��T��`�D'�;|"�j I��y��I9�@����>[�9z��y���2!
�k2㝌Si�@0�yR�^sZ���蓱�\$�d��*�yb�S�k�����N��2���H���y
� zd4)Η&�x��u��p�LH�"OJK���/;Dz��Dδ4w(\�"O�u� 
#sq@<�`�~��Ⱥu"O�c���*AŸ$�#�7Q���&"O0x��I�+n��ta���{K(�%"Ox(�dX�d�KMW�81��Q"O�İ��Fy�mBFF�='t���Q"O�A�s�%\�RJ僪N��0"OD(�@���N���d���a��"Ol 3B��72�f�AqE�1"p0ц"O�h��Ʌf�|;a�� &�q��"OV;��;���1/��h�T���"O��d�I�s|H$� ��5@d,�v"O��ҦϜtD�p��L�N�T�C"Ob )�̈́;C$x��� Շ1�\X1"O8�y�i+v�1���V�x�"O8qRuo�A���׳,r�(t"OH�*��E6JOv|I��I��ܸ�"OF�P1���SvXp�JQX�Q"O<� ��G�'�4-���F��"O�Y!6/��i��q'�ږ;ԒȈ"Or�iP'�6Grt]J�j��;^;�"O"!�Cj�%�V���׋G�i�"O��"�ݜ6��1��A�J2-q"Oh83�W�X�h{q�̝!:��"O�s��CH�c�'�O���"O�X"��J���Aas�T�"�̍Y$"O
�w��;7��$:B쏄�N��"Op%�Ĺ0 �g�^���C���!��NQc<���rDp���>U�!���>�����V.x���G|�!��A��Z=�T�_A�:�m�3�!�䋌a��[�O
�!3X����R� !�dܧw�L�9�m��$ụ�C#�!�$VR����%��L���Dn@!�dN8I� l��ı�|5���)!��3yr�qd&:�La�&�7!�䏋n�����T=r�,�3��T!�C��ܱ�)Ͻ_Ȓ�0�d�!0�!��
M�0��h�	L�1U�V�{�!�D�s=X�"�䛡��{c@\�b�!�΀8h���]$
��Q�`�!�dA>���4��-稠C�aJ��!��q\����J�Z��W	S�!���\�pEÿL��\�1���!�d��Q=؈�tΛ<
�R���iU7Y�!�d_�\�^�S�� 
mܖ8Yv��!�!��@��y��Q�E�BP �܅!�$O<��Y{7g���������!���qh���h� +�T�1���F�!��L�<�(XI5ƚdx��2�!��fQn��׀��))%/̺fn!�M �`PK�J�/�Hy�cN�e<!���?,��*掤6�]�%��B�!�d�1<�2L�6�(�j�AԟI�!�D[�*�\[�	����U6)�!��L
\�t���0_K�E�����!�U�����v�#9�-� +�k�!��F�>�L�`o�,J�X����V�!��@�����3v���cƐd!��٤(�F���Yz�ݓ��Պ�ȓ*~�IK�enm�U�ÕD`(��ʓ^������)bj�D�l3{�^B䉶.�D1�7��+y�^��P��S B�)� Ph��m5QF�L��Ø�AbQC "O
�H"���I�P;���$0r���"O�Ph� A�uԸ:T��+,��E"Ob�Dl�-���Q1�G3:T�+1"O�(K	�UȐ���M��cWy�<!D��~�B��Æ�� �BP����t�<��DQ�@,�F	͠����AW�<9���y��5��2m���`�S�<	���b�`�0��P��B�%HC���ȓ!G4�ʀgF{�v��ůKn[�Ą�hUhpI�H��"����� e�Q�ȓ5~���� (,� ���Ȝn��L��V���+SF٣Q�@���y��U�ȓXZ���C��Trp�,׾d�ЇȓHH&)Re*�=|�BAP��>S����QI��S��Sid��Z��'��݆ȓN!�9"�(?j�LŀW�J-ly�Y�ȓ/ي��a��oQ�h�wo)L�T��q-P��&CM2�*y�bEO#\,��ȓp��x[���		���r�&�ƹ�ȓ.��  @�?�   �  �  ,  �  *+  �6  �B  �M  �Y  �d  �n  5v  ��  /�  q�  Ϙ  5�  y�  ��  �  ��  �  :�  ��  ��  %�  }�  ��  �  L�  �  ��  2 W � � �" �* �1 9 `? �E �G  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<���C����P��1�ޜ�F�Ai�K���3bH-D�x��U�Y@�L �2�3��??�
�"�^��"D�*N��UOB?U�E�ȓ0�v���,[�� ��T�Y����ȓp�s�MӶs��yU��9�z`�ȓaZ`�;׎R<g�����;UU
)��X��qaE��?F�d�$��]�ц�rBj���H?�dg�A�5潆�%�:��(�j�  ��I��ȓs��Iȟ&�������~_����@J�<�%��"@+'I�WưH#�'�����˗0oءh�hY-O�xm�
�'�x bi~����N	�/>��	��� �5	1�#!�����:(D�D"O��B� 0X����IR+9^���"Ol����yӂ(��'<x	Z����	�j��[�M�e5根b��O<C��K�����'�a��`���(
C�	Jmry;�	('�u�!�B��B�IR�����a� J݂ �F����B�"'ޖ�V��
yH�q'$ʷC����hO�>�R��L�%����)��x%��Z�a=D� j��K\L�B"�35T��:D��qc�gN�x�&+
�E�U"��6D�ػQE�2��B
-m���颭'D���c�57.E��\�Ĳ����'D�����G�:��#%�$rR��V,%D�0%!X�Zք�EL�~4J,�@�.���<q�.uR������0G�y���X�<�bJ�?c'hA���	�$������]�<��2m�~i�FHͧ_�\Y���p(<A޴Pd��J��?�0�_^�y�ȓI�i+AI>0�L��'�ƛl�����6�X�9���&[^2��� -��T��~t&���\�(4��C��?�N5��Sj�pZ���k����FG�\��@�ȓ{��؂4�J-$,فW"L���ȓl�8E��3zAA���2h�م��zy���w�r�.������R����y�b����9���p:)��%���O��G�4�03Nx�A2f� ��xPŎ��ybJA|��|3���p�ˣ����4�S�OVxDG^R�H���ʨ$R��	�'B�T���X�T4�qk�W��
�'a,Ƃ��j�	��C	���yR��G�4�8��
R�Ip��8�y��sV*�򢫜��*����!�yAW)W�pl�4�y@��(l����	�'8�MI�,�1�6)��l��X��'^��N]b}j�����/����'a��Z��°O��Y�F��`�N�І���2����g�%;Z̀!$C�h�b��F{"�'���%ph�bE��6'�:�ˆ�	�U�ȓ!JA����T�ai�7L<��>��'Uў�M`�jC�Ԏ\%���AÈL��C��:!��M���C
b���ۥ���(:vC䉸 �Xe)�ꔹov����^;wF#?Q��iD4n��|�&�·��S�Nե4�!�.$� �.`�
ik.�:���M��H�P�!eh��`X�sdiфq��[7"OƜمg>�d�(A5&Y�7"O�1��ǜ31�U!��TF�DX�"O:u�.��LP�q���>\`$�s"O�IZ�@ͧ9Y"ݣ1&��wO�B�"O��!b9L��T�d�N�����"O�c��/Z������&��|Z�"O���ר��6�ї����m) "O�m��I HK�H�#�ߴ?���C0�O�ʓ�hO�O$���6n��+��%i�*�X���N>Y���	?�"|�`�
@�����@)j�����	��!�Á+Vl�fm��%~���I�&���j���!fQ�V
�X0@C�*���Wm�=����'�HF*���ɐϘ'�>�sqa�D�҄i�'�K�ϓ��O����
Dq˺��3�^HԼJ�"O]Sף�J` �S���!���"O(��%��Q���k�6P��E"O� � Y���;+�t���\q����$�O�YEz�O`F��	PF�=����%Ĥ�'�)�ǣR��ؘz3��"!XҝJ�'�ў�}r��>	�ē�jzr��pGWj���>	�� 1�T%�BS�k��Q�"/�\�[&�=�O�|�Ê&W�~�۴�� �Y�y��)�Ӱt!aV��W�T酢]*H�d�$��(O?��H��D�����O3H�&L��m�i�'�y"�܀Q�Α���s�n��E]6�y��^^��PrA�=;�̐��ے�y��H�H�����U9AHQ� ���y��A\5�H)�ヅ,�:(���M�yb�?>�Tm`�n�QG,䘰��/�yrEʖy�h����!I��g�@��yr��PEv(ʵ�ڞ�vaC' ��(O,��D��4�&�sOc�d�F��!-��>)J�"��D�O=���ЌK8y<P����Dt��q��D��'|��@E?.2��
��!���	�E�➨x�o��HUJ!D��B٢t��
��P�}y2��ܦ�E~b��0b����6�L9�����֜�0>��xB�H&�* �$3�6�y�Md�!�wXpp+4��6@y�P揇����u��}BشC�4-CM�$Mt���o4L���=Ն�����D�� _�ST(��w1B��qh�p]��I%��"H��U<�m:�a�%��!`��
ک%����ɷ[���B�G�dP,3��;G��B�I6� F��
 ��'�5'�B�	";�z�r@�r��Q�fl�11��'!�"=��7��g���:u��2:�hYXC�\�<���GH��,G.r��<�BX�<��N �J��i�*xטx�`k�V�<�%��Fv(��ϱp�*vŒ&"O^D@�ȱ5$q	�K�"��2"O|�k�aɟ ������}%ք�q"O`4ZI�(��T���
�EY�"O���D��՚3�$(Rތ�e"O�<ӵ����
`��dA� TR!�7"O ��U��T�V4�E��pB\0�"O衺�I��h������=,�p��"O�W�5�q�����@|�a�ŨBZ�<�uaO�o�����'ؾ�F�S�<IA@%:$��p*�
dp>����Z�<����x�:q�G��e��0c+MU�<A3�jdK�	[�r�L����O�<dG��>��M��d��I�NHH�d
p�<��	no�tЁY�X��s��'T��Y������pé����	�#D���Ƅ"q<���M�:4-����!D����a�O�:�J��@��͓h!D�h���^+슐1�l��f�	l D���С��Lv4{T�]��y��N D��K���"�!rAͬ@��ua�c<D��*q ��j�̽cP�~_�(���8T�x	"FX/ZV���ݣg�R�"OйR6� jx��P
ԨH�~$��"O���!��=.&�"#J.q����%"ON�3@Ӹ!%|��P��,y���	"O���Bƛ.~��͠4N��"��R"OԽ�#O�x|)��1�ޙC`"O�MbJ�F�r�R�oƟl��a"O�t9A�
��	��d99��e"O0̓$���n�|������K�F�RQ"O<��"��c�D��"[W��!SG"O� p���	K�׼�6K�&?��%Q"O�����N�&`ڶO՚x�j��q"O�Y�tk������N��t�.���"O� ���p�x���˟ؖ���"O.���	�2<N�D�Z/2�6Y���'�2�'���'���'r�'�b�'�<��B�x �9�bG�#*Fy���'0��'\��'�R�'B�'��'>1�gd_�a椠���	^���1��'�B�'R��'fB�'7"�'���'�B!��!_�A���@��-̆}�Q�' b�'���'�R�'���'ub�'� ����K$L��ǜ5t�y��'Q"�'T��'���'�2�'2�'6����Ёp�i!��F�t���&�'4b�'N"�'���'�'V��'6i�qȈNCR������4E=���'���'6��';��'N�'pR�'�lش���A�H%&���hSJC��?����?9���?a�Ӛlן��ٟX��]$N0&l��F�Zt�"@N$���۟,�	���Iן��	��<�	۟��	���M̎*>Y��ʞ@F���Iܟ��Iӟ��	ڟ��I˟ �Iܟ��ɟa��a���ɁG�x�#�
�A�ʤ������Iٟ������I̟���ӟ��I�X0V�����R=����t�20�I���	�H������ޟd�Iǟ��/m`\S�꜑݂}�!<�N-�	���	�4�	��	���	�4�?Q�5S��[�-�&w��(3�CG�>��9['U�$�	Oy���O*�mZ�pU�h@l
)��!t�g�%A8?A3�i�O�9O���P�&ᰰ�ށ@:�pc�X������O���6�y�����D ���OLf��U�|1��+V�>�h��y��'��	�O[^PQUo��0
 �nG��p��abӚ���D+� �Mϻh��H��D�+����0�^?VX	���?�'��)��9
`�oZ�<уO�&t&ri*r��("��<!�'���dX�hO�i�O
�hҧ��F����R?v�(]0W7O����4����ǘ')x�Q"��	iN
�XD��mg\�у�IB}"�'?O�|�~���FRf�YR��?����'0�摕>TyK�����՟|K��'��0�fdG	�>�Kc��
���a%X�h�'���9Ot�1AƷpǆ����9���49O�o���
W�F�4����s�>D��ZA@7_�.\;�8ON���ON�d֫"�>7�5?Y�O��	�)C��i�5�p�Z�{�H�yp:L>Y*O�)�OF�D�Ob���Op��k�"Wl������lp ���<)B�i�A���'M��'�OL�`��~Mȹz�aZ�k9F�X��"x�\Û�i&�)�Q�XͲPg�HJ��E��:+��!e=p�T���_툽�HۊZ���;<�'�^�
����AU$UM�X�?C�L#���?����?!��|�,Oj�n<_2�A�I�3&h�&��Mz���1*�)&I����/�M{�i�>�F�i�6٦e�S���`��eW�I�r	9AL,_��o��<�!�S.#'Pɘ�'�3T0�xN?1���w����/S>m�p���'P��@�'���'���'���'���;F�T�hp<h9��6F����OB���O Ym�]��-�'1�6-3��Ō57��b�`	=k�.\�R��X�$�\��4JF��O�6�b�i��ɋ]n�Z��U�*"l Q�֐o�X�� ��T��"�Ty��b�h˓�?a���?�����k��:�e�o�pqI���?I.O0�oZ.r����	��Iv����HX�x��,Ȋ7�
c����d�Yy��'�e)�T>���A����E	�	�8���tJ�*M*T��+Ѕp5�P�'�6�]�N��Hwy�wt�:�iC�k�<�n�a5x�J��'�R�'���O���M�DmX�d��-x�M�V�U���{)�k��?��ia�O(X�'�P6�ų]�i`���@��03�M�M��8o���M������M��O�e������M�<��\�j�"�z ���J��y��އ<n�]�P�	̟��	��H�I� �O�\,�S�J%f8d����<R�p�0pLb�b��B�OT��O��V���Ǧ��-�zp�r✋�~Iг�%F�<��4NP���!��Ԃ(��7�m�`�C,Y�&3vQ�T�w� 0n�!eH�$��4A�� ��nM��Y�,��͟�@���)y�8�C�J9|~�!�@Ο$�I�(�	Dy��aӢjg��O&�d�OP�(DA�t�1�2��i� M��!5��/��D�֦9h�4_�'�]��N9MȪx3��N�[�&���O�UAg`D�~ӠM
Ca�<iF��Z���2����;첝��E�&c�l�S��`����O�D�OB�$(ڧ�?�r�z �ࡣ���¥r`�ӕ�?���iČ����'�`�f��]p�*���"@]�H�-Vc�扡�MS�i�z7l�6�#?���\�?��	Y�N��*l�mI����@(/b�%�.O�!m�LyR�'K"�'2�'�bLݟ;�4%�c��L��E�#��	��M��IC�����O��?�h �
��� �W�#L�a&����I��0ڴ>ω��O����0��2����~|:�`�^8
���`�W����
{���Lyҧs�X��8� ��p��YjU��O`�,����?���?��|�*O��l��N%��I�VG�!���G2z'�`r!Ȁ�r�
�	�M�2d�>���i^�7m���h�"��3�,y��RK�	�sa� bwĹnA~2(O�Q7^��S���!�u���� =kҠ��v���Yↇ�t��8O8���O0�D�OX���O��?m8��K�9���dKW�8�(�)a��ǟ���ϟ�kڴ*Q���O~7�>��$�ƌyeօ���[����PL&�d�	�<��s���oc~�B��h�sd�݆r�|��&�P�gL��Q�����D(Ǟ|�P����\�	şd�AO�{ ~�£��M�l�$D�����	jy��w�,%뵅�O\�d�O��'})(� !G�H˥F]�=Tm�'����?шʟ$ �S�YSHx;D�H�'�@m�k�&���G�7A���|�'�O�:J>�7�C h��P@F��P`j𢐵�?����?i��?�'`���N���D����k�V%�Y! �Z��2���a>����Пx��4���|�Q� o 5N�<�"ڮ%��I���|s^]K�4A9�V�ӓr�6<O �DXJ�D=���.��iوn��_b�5��m�)L�̀I:O���?����?9��?�����	^#���[rdK*h.T���5A�l�n�EɌ̲�"˟���?��쟜�I��M�;����BhK�h�ڔl̥`�f���'����=��O
�T�Oo�xu�ie���{��e�R���My��:1���! &%��]���O��|��4�t���i�}����c�)J��?����?�+OĔn�gT���ܟ�	�l��,���_���$';����?�P������x&�l〣T�P����� {�P�"� ?9r�ƇS%��Gh���T&��$�?�CY�O���
%/؆��T���?I���?����?y����O�0��ҟ; 9yf�,|�Xxyc)�O�m�Y�����˟�Yݴ���y�!�L&�(����J��В�yb�'��I!<�1m�d~��_�d�9��L�\�y�fŲ lؔ��cZ���|�W����ߟ��	ڟ��I����ҍ�0e�����$8P �HyRkxӴ����OB���O蓟D��ԿA&h���m8Yf�-�a�'�7OjO1��
���.`��Hs�(a�5JӡԄY���RF-�<y�hJ�Vr�5����䃇W؄	R�]�;�(�A�ݷ����O����O��4���eě��Nb.�;
�`�)�M.R�;b/L,6���rӸ�T��O��o�5�Mc��i'xĉg�7$ �d�ݗ�th�#Î+J��f������v�������TZ� ��ň��q�4a69ON�d�O����O����OD�?�`dK9NO���S�Ҕv�H `�����Iݟt���:��S��D�ڴ��j��qD+C�j�L*��I-l<�v�|��'m��"�<x �4��䚥lD��Ѭ� ��:h�Y[��gY��?Y�O9�D�<Y���?A��?qFo�!�Q����tʥ��Y��?����ć��
�ΐ͟���ʟ��OF~��pC
 ���`��T�D�8P��O�y�'-b:OFO���Y�b}����
�����.N"
�Np��,BQ�� ��Oy�Om���#v�'[�M�Q��Z��B
P5o�Z�'��'����O��I�MC2����q�!7iR��
>��� (O�@lZR��$7�	��M���4v�i"c��c�l�Pv���\�r�i#�$H�i=���;�4�)��O�l�'���+5����I9���wX��'P�	ԟ�����Iџ��H��ER0k̬CC�W=h��cP��*/\7m�wil�D�Or��+�i�O4�mz�!
�-: ����
+kTX���
�M�P�i�bO1��]['�n�(�*4����5@�ڄX�bD�&�*�ɻQ�*!��'8F�%�(���d�'���u�="T^ԁ�bˌ(l :��'�'7�S�t�ܴ4n�D����?����ݠ ��d#ԁ� e��2�r���>�1�i�D6M�T�	%e����j+2U[�H��5D:�W0�
�R�k�X�|����O�X��H���¡�y�����C:M�ti����?���?����h�"�D�x�V�rG�e��B�M�7m����������y�my���杁DGB	"q�T`��iQnK0 	�ȟ��'��ԁ��i��I�Ӷ,��OBBA	�C�h9��+�+���BǩIF�Iky��'�r�'���'���*p����d�n���c��4��	��?��Ο��I�T$?��ɐg�l����#mz�i��AT�f찰A�O�mo���?aN<�|*&B�=y{��$�b��R�gG�   4I�g���� �P�� JOʓ�4�0���8�j��Dc�S\�H���?1���?���|"(O�!l�A���ɶ1ۈ���;m��@G��"f��M��c�>A��i��Dl��;��g`K���(Ae�b*���e���%ڀ� T���J~Z����k I)X&��I�kr1��e�0������I�����֟�'?�[�
�-�|���ΨN�� �3`�  @ � �쟼�I#�M��GԀ�?���4��f�|�d 2��Z��"%Y l�E��b��x�M`ӂ�m��?u	A�Ц��?i���%�:)�U,��d�.�hg�C*P�q�B��Oz9@N>�*O�I�Oz���O�lXsQ�IxQ�s��,-�65W��O^�Ĵ<��i�����'�2�'�哊c�q9vg�^�>���Ȗj��.�����(�	��S����g(�K����82e��e��qp�+H���<b�O����?�b>���q�v�h��	#�S%�
�:���$�O����O���<��inh�ÊRv�� ��%�t�dH<9���'5~7�%�����VЦIR`Ӡ"��T/C4>�lJ6���?!ڴ%�Z�ڴ��$y�h���f��S�? �q�L^T��ƀP�F��Di�<O�˓�?���?����?)���ɍ#>rï�A��(�-�:xMP�mږ='���'��D�'6�7=�`i��G*�(nLwv�� F�O��b>�;�Nڦ��"[���A�
~���&��Oyp�ϓlvB�@�O��N>i)O���O��ـ'�wR��d�J]s��O*���OD��<�ƺiv��rB�'�"�'�V�zdn����Rg�3z�� ��|r�'��3����i��%�Xy3G$@���P���nj�U��$z��I�N(;�-\�
^����6 �O�h���E~0w��
\��EXT�M�pW�Q��?Y��?�����?���?)"f�6x��_)J}:���NZ�v��$�I,�M����?9��S`�f�|��yW��MJ
�!�F�p����U�ۈ�y��pӾ�lڡ�M�p�4�M��'r�[,����M`�4@p-Õ Vm���O�M���%�d���$�'��'�R�'���hT��.����"�Ҫ3�@���_����4i�L�)��?I���'�?���W�z�2m�Ь�6��pi��������Mc��iE�O1���K��Ǥ'.�d��)�6;;�P0s$Nm�@MR�����ș-��DQ�IYyb�À�Z,N�6<;��ηT'Hi���?��?���|*-Ot�lZ73�6�ɠ<�ꅂ���% �8!ˁm��pl@扠�M���
�>A��?Y��iΊ](�M
��и14�I�I3� a�Y'%I����������c���i��2�q�W5%��Uí_�&�]	V1Or���O���OD���O��?�U��	x���1��K�F������Q�4FX��!.O�qlY��h<�rA�"�pc"�_�Ɔ��I<��iz6=��p�"lqӆ�q3���(�:T4V�a�\�pA�C�<�6��W�����4�����O����PF*�� 4�x�z5��|,n�$�O$�y�v-�#�R�'0"[>5٣/Rl�����'�>�i4)"?	 _� �I㟄�N<�OB�A�p�ɚS���ɔJ^k�V�q��Զ�Y�@���4��e���0�P�O��Ȇ�Õ���f�(%��J�b�O�D�O��d�O1���B��D�+\邠!˛0 !�엂=ܾձr�'B�eӔ��X�O���2�Z����F�<����6nhʓJ�P!ش���cIx�a��:��ʓe��F#W�K5�8+bӨ��(����O���O���O8�D�|
�*Ʈ%�:��� �?���'�Q�s��6M��5=��'�"����'ފ7=�( �뚡69�%Z�d�j2�3��N��:���Ş�>!��4�y����tԸ���,�p����A_
�yb��~���	|P�'��Iԟ0���u�,@l8�ir�*d�nu��ǟL���x�'Y|6m�L��d�O"���=r�؁1N'bx
�:�C�W9d⟔��Oɦ��ܴF��'��  �A w2��`d,+ps��On8Y�h�Oʰ5H��)��?�l�O���P��=G����U0>�=9s��OR���O���Ọ}2��9wd]��
�o���a�l�����.��f�Q�;.��'\�6m+�i�]P4䏾M:�C��-�.d�Q���d��ʦ�:ٴ�d��4����	!��h��+@k%�U�"ڊI���~�}0DϘ�����4����O����O�G켠aQ�E���eAV �e��狍�2�'R����'���Ƨ^$�!�]�q���c���<���M;��|J~�E/W=I���ӨT1a76����H��T!�q�c�O�)�K>�+O�u�G�XS��_ k����O����O��d�O��<	շi��RP�'�\�	fᅰx�����4����'56�#�����$ͦ�Iڴ@��ƣ�j7�\y���`2(�X��:$h�봵i��Ib\���`�OCq�r�NYGq�(0�K>�<I�á_�U���O��$�O����O���-�	7������_�$��@%'�؜�	؟��Ɂ�M�E�@")O�dn@�I��f!1$���P-`��ȝ(_�ZI<���i��6=��5Zd�~��D) ��3I�����:��0C��ғ2�0��ܸ����4����OF����<�y�����@}h���T8
�d�O�˓D�V��pYR�'�2W>���H�6��Ф��O$�S�%?!4S����ƦbK>�Oi��Ri��#-4�n���d9֦�!)����1D5��4�h=��`^��O�pI��+|^\(���"���b��O�D�O����O1��˓`��#H�(m�!�J�B����f�ٰN��ԃ��'���mӄ��J�O�mZ?wkv����	�45"�#ya�Q�M끵i��s��i��I,�X�ؐ�O*�B�(rB(�!w�r����ܬj�B!Γ���O ���O���O���|*&,F�8�||`�N�Bƨ*��C�A��DYB�'�B�I�צ��y���	CK�/��Ix��]%�����?�J>%?M�wGަ�ϓs�H��)�1��8r&�]#I�r ϓN��B�O�5�N>I+O��$�O�	z�	ݔx#��H �Ԧkv�Qz�+�O\�D�O����<A��i���s�'���'�eS�n�13fU�®��w�U���}��'��$���C�p`$�ڃ P@$�t��B}�	�;�*$��7��<'?12��'�����B]:�1�ǁvK ���H���M��ʟX��͟���T�'x�6�0��-�ʘ@3o�	�H�N$ٜI��ϛ�ϝ*��'�Z7��O���?�;�����j]D�\	8Aaʺr�V5�K������Xl�'8ioZ�<A�έ�'/����� Di�tm��r���L�R �h2g4�ĭ<�'�?���?����?i��6"�Lz$K�Q��  ���?��$����!�����ӟ$&?���9^�昲䞧fb*��t���%۬O���&�)��LA��2�����Ӣ�
���g�j�'q`��Ä�ޟ,�ѐ|�T�����L�I�� T�j��H�$����X�I���Iܟ��Ly(}Ӳx�g��O��E�q����雇hd-09OHmZX��u��ߟ��I��Md�0M�Nx���ʡH|m���ġ��sߴ����>>�,���'��O��ĕ�9���G��!J�$ �2��.�y��'��'�b�'���	�_�r�0�� u0X�f'͍j~����O�����u��o>����M�J>Y0)TY(���E�k
��������'7�7O�d�Z2sh����$���������YBl��%5�d��E��H_M�	^yB�'C��'a2�Ԙkc.�+v*��-=��bdK���'��	��M6�5�?)��?i*��H�,�=zD�􎃭.2�2��H��O�l��?	L<�Ooja�d���m@w�цQ�v��d˄fP�n��i>�r2�'o�y'�LrF��w_6U�#�,jb}Ӡ-����	�l�I�b>%�'��7��D����m���h�E��P��Q��O0��L��m�?Q�]�p�I5b�>pyf�D�b$ )bBKE7�6U�'�p��ߴ����3p&���X*:ʓ�$�2�bI!��	SY������O���O��D�OP�Ŀ|�PF�$�f�����@8�I$)Y��fU�^PR�'��O��0�O'b�{���1R挹�#=h��k�"0:^8��,�i>��	ߟD� ��ݦU͓xgx$�waVI��Ó��:�v�ϓ}
��D��O��I>�,Ox�d�O�܂��(+��9u���6lX`q��O���O~��<��i��3��'8R�'�����@�:㌩	�NF7,Q��#��ďW}��'�O���C@�mF�dB��Ƿ_HL�HA����gY�u�|���IO��t���	ݟ�0'J��b_����W|�D��E�ǟD�Iџ����XD���'0,49����zx��sP=}��$���'�v6�y�d�$�O>�lf�Ӽ�G`ϥ�LPQ��$���ӑ���<yU�i� 6����+".�Φq�'
�!�G�?����Vj�1v�k.v�:g뛛K�'+�i>=�	�8�I�l�I�}æA�P�кhf���-�^Ԙ�'��7-�/R��Y1��O8�d���3a��O���R�had�� ��SA�Ԁ���	����'r�i/�O��Oa��������@�Ɲ07����ʳ[�.TpD _%��$�=��M���@*�O��)����D����D܏M��4���?����?Y��|b.O��mڄQs��	�%��T.�1� �o�p�
d�'�7� �	=��$P�����4J�c�6�JqC''��dJv�\"?+j0ɢ�ie�	�r������OIq�j��U�`��u�┿;�����3+O�D�O��$�O����O~��>�ӻP�J|�gc6���+�#'M<����`��<�M�q���|���=K�f�|2ဃ,S��˚�!� � �EM
�O�m�󩚧jhv6)?�p@Ws��$�O +���ϫ-s �W��O��J>�/O���O���OBi�u�سL�0���,L�i3�O����<iV�i�4ٲ]����`��+�)�&�	U�}R�u���,��D�qy�'țM2�T>���O�G�D!��!��][a��	<��-�0�^� ���|ⲁ�O�Q)L>�3�\ t�N�a��*O���
��0�?���?9��?�|�-Oh<nڿE<0��8nJ��� �"R쮝���������M�B&�<��4�9@��;�<���"�
^V�a`�ij7�D�9�7-$?P���4�,��:����{65���,Nؐ�
�e���yrP�d�	ş �	ҟ`���`�O�z�1����1��� ��L(,�O �� ��L���'��ݟ��I���9VʈHs#�&Blx
Q�4#�Ν���?)�Oj�������H�Qch���If�p0�jðs�L<�B<g�p扳1�6(#��'�.�&�$�'���'���*�!:"0�pR �V"�u� �'NB�Ԙz�"W� ��4zX0-���?q���8�d
�_u�Iӄժ���bI>a��$��	=�M�v�ih�Oh�P�`ʖ)'���j��3(ļ�!8O:�$� �F���d؋��I�?�P��'=���M�$��fDU:�*�!�T�$��ȟH��۟���W�O�*���^��e�&>�Z�9�M7,��mbӼh�ԇ�<	d�i��O��<-]j�Q)�ki&�jA� &��Or�I�@��˦Y�'�
@��?A�.� ���C�2Pv�30�N�a�ԫ�n��@��E:	O��lC�0�>p ��F&Ts��K�u�n4k�&Cq�0y�(B)tXB�����D񔈝�K��$#Ĥ��tmp�	b
U��m;�l
9Tg>m�ģ>��='�T�br�S)c1��M�98GF�R��.A1rG$f�L�#3��7� JB=KL��gO�7$6�WAƈ�)b�d�oiL�qͦGi�\i��90#^�Q�gã��<��G˞ PxI�ra�{AN��Ȩ[Q��*�v5\|���B3J�@mkw���+߮Y��ʘ$P ���OH�D�<���?)�k�4���Ӛ��ac,�9e�*���i�b�'��+W�:����O���)���'[ܠX��KF�b�N��43)�Y9���?!/O����</On�cd�E���f(�*C�l�2*������R`*�b�"|���.@��[��[b��h�r��7v�4D��i8�'T��C�o��'��S����{����2�P$k�,[�\�0m@��H�Z�ΐ'>��	ǟT�ɂ�� �a����,m��25m�E٦B�i��&ЅY��	��	�OH�Oa��)�;+��5�G��g�=�è�Y}c#`����OR��O���<��7TF�Tr#�
W�Ip��ntST���'�2�|��'��/��|���!#'@�AEQ,3�Q���|�'���'c�	�U�Δ �O��RfB�e}6$E��m ����4���O�O��$�ON��%�����k��[��Mr�Ӊk��8�K�>���?�����S>n��t�O��kث̉�RH �Y��1 D4U�7��OL�O���O�4�t��Oz5yQU�4����0�௎<Z�H� ��w����O�˓*��ɱ\?��	�t�S<d��kRB"�p��ޛ��tM<���?�#��'^�)�WN�(���O\>|8d y���Z������M���?!���BgP���=���R�A�*��tA��ďxI7��O^�V�zt���}�S ݒ�PP@KM�
�XM�E,NӦAS�fܢ�M���?���BQ���'ٖ�q�O�0Ҽi���[�$[N�rwm|ӄh�t�:�����?A��w�t��5��-	ct隑+�n&�f�'�2�'�0��A��>�-Ot�䦟`�!2G�"�@��H�-�4C'�a�ޙ�����3�Ҏ�ħ�?���?��m�/1-�$i^��`��!�BA��icR��8]܊ꓦ��O��Ok�]�E�*�zQ��H&V�Y�
��f]��*N�rb���I�@��Jy2h?1�p��ƽ 2:D�����nՖ��c�>�)O��$#�D�O���&@��|[�r:h�I��^t���-�D�O����OJ�-/�|�F2�X8�H�|��Ъ��8٬�#İi�	͟�$���I͟t���Sa?qcoD�^�q��P3O�VX�"�i}��'�r�'P�I�^ݢ�q����DD�k���sP�P�)��h!�Ǳ��yn����&�p�����!���ޟ��>�E�".���i�<~��hx�,�����쟨�'!�L�~r���?I�'� ,ЧY�m���Q3����x��'�$�@�O����i�.�c#�.���n#$.v6M�<���V�'�2�'���o�>��R�Dyc�ߎ&�U*��J�1��l�����	kb�A�?Y����P����sU��$>�hE�� �M���[�.����'�'l�T�5�4�X\P0Έk���T"�L��k����	؟(�	B�i>��'�2e�)*���������Dɱd��7��O6�D�O�s�x�i>���P?���B�EY�����hvE�@˦���w�	���9O��$�Ob��B
n@�8���	`<HD��XdmZȟ�Ȕ6���|�����Ӻ;� ��@���(ʀZ�9��OJ�Iߟ�'���'c\�DBŹeǂ�)~.j�۷%Q�*�$٨t��v���H���byZw�NQ!sAQ5OR��CH��Lx�4�?�/Of���O��$�<I��]�},��19�@��1"�����@Q(�����	n�vy�O��$G�3a[��C�(��e��aD�uf�ꓝ?Y��?9+O�L���u�ӘA�ZyᰯV )��T��Î']����4�?L>1.O�i�Of�O�j�5
�~�D�I�Ōњ!�l����<9�����-�����O���Ʈuӳ��K�\Q�V^�@LsԔx��'��I!b#<�;Ys�J7�8\X���p�@h�'b
�/�B�'��'��dY���E�*5�a-��5��iJ��27��O��7���GxJ|Ԇ-E]X�sc�6_��9��O��1�e�O����O"����$�S�ԏ�g5�L:E�<���*c䀚7A��E�Gx������L��+2)ZU�� I	Md,�nܟ��I��hg��Eyʟ��'�`(��]�h����CE	h�th��>R��O���'����5~�^�A@]�˒�!k.6�7-�Ox���c�R�i>��	H�i�K�&O�+ŊĢ�,ȟ;���@f�-�$�O���?	��?�.O.�C�͂�F�Rt�s�>�"����	�0��&�@��ß�'�D��u��-'�~ɀ�eY�4Y2,��M�������O0�$�O0ʓŔ��U:�*yH�Q?Q}���j U6�P��^���IƟ��	lyr�'��矐zf�@�; �Òb�z`�1�����O~�D�OB�J��G�}�ӊ;����"��0���*]��Z �ߴ�?�K>	.O�	�OX�OŬ�ٖ��	���Z�.�3xj�4�?	����0fW6a'>��	�?�ؾ9����`�`�U��R�?��Ol˓t�&�����'��tCη[�nL&l� F�T]Y4���M�.O�x�*�E��� �D��,�'2J%��a�4j���Hȟ������4�?��p�>��"��S�����s�ܴ>�*���gR�#M�Y��yV�nZW��(�	����T��ryʟ(�qq��x٢�&E�Gh`����-Ȗ+�+	�>c�"|:�P h�SE�lpx��	�d�v5�i0��'����/Z ����O��I<j��m���*�0��%��;0�7��OR�N���S�t�'��'��]!�]� D����-�x��x"�|����\�TL��'��I�Ԕ'�ZcK�Œ�$U3����@E�/�ΰx�4'�fY!3���<���?A���?�����$��T�Y��0�Nѐ�.�Of�ȱA�X}�Z�H�Ipy��' 2�'CD����G83�L��b!N�������d�O0���O���<	w��?t��� ^�05��*1jH��!i��4�нi��I֟��'�2�'X2N�y�j"Q�ꠐ�>K^��#ŁUw���?	���?�+O @�w��v���'��4���J/=��; h�:s��1sah���<)��?q��t��4͓��$*@�R���B�O�`}�ԧ�!&!^ ��c�O��$�<�jώ f�S����?�*��ޔ6Ϫ�"v�Y�^ņ��Ç��d�O����ODt�>OX��<��On��F_,@�p�ڕ	ˮ5�40�ش���˖NYԠmZ��4�	���������"퓃c�1'(
��ţ� fb�is��'Pp`j�'��'���F���74t���@�qs�ō�R��fi�N�6��O����Ol�	�V}�^�\�P����J<K� Jgt0��i���M[�o��<���$<���`����A�Yi��G:u�DԡנN��M��?A��jЩ'T�X�'�b�O$I��m�4|2�s��-Ua��؁�i��_�`c�c��'�?��?�ĭL:"�ry[�F\�v�X�sF���[�V�'�t��W�>�-O�Ġ<���s0�Il�uk�m�	0�@e1�@}���yR�'�R�'���'��ɓ&]�!ȒM2e��d/�:,b[,w��ӪO���?/O��D�O���J,$J +Մ<n( ��R
hE�6O����O^���O0�Ĭ<�� �.��	з���Ԉ�>�~캲M9P��6S�t�	Qy"�'���'��q��'4�#��/_h
(rOH�`x�nh���D�OF���O��4U�T?��i��K2���n���@�X���ۑ�g����<���?���f�y̓�?Q�B���$�ܿ7&�,�$�ÀL�����?1����!��O���'l��HP-1�f�k1�X1C�H��sض(\��?���?Y��I�<1-��d�?��3� ��F�
�U*pTl)��oӄ�<MZ�C�i��'���O�Ӻ��,P�n����D�Bff`��!ۦ��͟h�f	i����`yB�i�ZD,�s�R#S����Q�4�ք��rҘ6��Ov�$�O��I�S}2S�0"b��9�Y�sJĢl�qs���M{B�<,O�Eȓ�<���?��A�vi��c�G�j{�#�S)�M����?a�'��x�]���'/��OdYsA�������L���XaAt�i-�P�0Ksf��'�?���?yA�ݢ��x7��a�	��_~ϛ��'O�r���>�/O\�$�<������{�@�#s ۭoR�x�d%Xp}�.�:�yR�'�R�'���'d�	Lg����L77fM�O�?Pg~�Q0Fɶ��d�<����D�O��D�O�UR#��C&HIF,��2�Z KW��,���O�d��"���OZ�	�$l:F0������VT�eyt�	K�	�iW����'V��'�����y�e�+��c�݆(�F�g�>W��7��O�I �*�O*�D�<� ܫ/����t���Y(B� yW�@$J��1A.�M�����Op�$�O�|�2O��{���F"E��� )�eF��0G��?	����$�$�n��O��'A�􌄼(� H�N�*%Qa�nʴؾ��?Q��?��i��<aO>��O�@�uF�'�%�&��l���4��F#���l�� �Iߟ@�S�����D���K{&hr�AKw��� �i|2�'J�싚'�'�q�Ľ�@?��9(�EJ@
r�i���HR+x�Z���O��$�'��	��x;���(tm�`�X7y <A��4r�������O���;�t$�
:*�ր�aO-S8V6��Or���O���u
J}[����t?���!(����T�� %��Ve�q}]���V$%?ͧ�?I���?�p荤tD��/+`�q��� ����'�"tk�C�>I*Ov�d�<A���)H�s��3!�9F�
i�GI�`}�F˫�yX����̟�	`y(�=O��뗊A#?��-�m�R���s+�>�,O���<���?9��Q�ѡ1��N�r!���
/WD�2ŀ��<����?9���?������-��<�',��p�"��,0��,�7��"�ޝo\y�'N�IܟT�Iğ�hr�}���b-Ш����	ڡL��16�� �M��?���?(O���f���'�
����'��m���E�m��1�F~�����<	��?��%Ը��|nZ r�����ٸ7u�� �I�+;�n7��O����<)s�P9��ߟl�I�?㇫Ä�uꊯnX=W0�D�'��'�b��yR�|Bԟ���@��z�����n	55�dhxw�i剱O�i�ݴ�?���?1�'��i�}I�9n�x��/	�=Z�с&x���D�Oz���5O���y���7z��[�AUA�����J�����wP&6��O���O"�	D�I���'��>k�<�4̏! ���2Ƒ��M{��[�<	L>ُ���'¬P�F�g�>q�5�H'ɚ��pÛV�'�r�'1���q8�D�O��Ĳ���gHŭ_�>U�K�,y+�I��z��O~�I���u��$�	��RA%�?<��t�E��X�)�M��&�D��דx��'-|Zc�P� ��RV���d�t���i�O�ikRC�O�˓�?A��?�.O��pǥԊW���6�Ru��O��]]��$����ğ0%����ğ�#&#�g�� S��M�~�0��Y�l�V]��pyb�'��'��ɪsZ��ОOyjDC �P��X�q3���*2��&�D��l�	�@��9@[��+"��gm@��}��e�+e~��'b�'�R_�lB�&�	�ħ
�&�`3ݪkh�CI94p����i�|��'iM0���>y)�:;�����L�_� Deg�ꦡ��럘�'�Y�=�)�O�)�z�? ��p�,)�� qFφF�,q�x��'�U�eb�|�П`���a\�ݮM�`HV�'pH��i���9o���#ٴ6�ϟ��ӂ��ɡs�ѩ���>$�v5⅀\.!k�f�'��)�:K��|��	u�z݊Ҥ��"9B�i@�C�F)[��6��OR�d�O�iNS�៴o�u�b�1G�Y7-�D9�֡�v��Ve	;���|��I�O�U3T�QG~��C�;��0�aզ������I<_8���}��'��D��>N ����C�4m�W
Z(;�F�|ҌK Qv����O
��O :b�E�b�FZ�ż�l�<�(R��ē�?1������@�2\����G�c�x�Ch�Q}nB7�y�P�<�I���ICy���#EZQP�n��y�he{Q �tl[��5��O��=���n.6Q�g̭;��K3�sS�S�?(OR���O:�d�<�A��>CV��J!Yx�bؽz>�"DOZ"b7�����F{R[���I�����0�
�0��M��p=�e��OT���O���<�F�� 2R���р
�W���X�K�'�~�F�D��M�����Op��OY���i�xdjE呝�()q�A���Pش�?�����D��W=��OC�'Z���՛E�J��PG8�r�)�(LN��?����?1#G��<�,Oȸ�rF�?�"&���x��a!�S'ThJ6m�<��%I^��&�'h��'1�D��>��R� <��h�8A0�h����lZğ�����:�	"��9O��>QC��Ԇ$�p���e��-(�|�j����æY������I�?b�O��z���{�j؃�V|��%���i�b��'��	�><��*��]����*��29Xtm�3p�HDj�i���'���H�듲�$�O���=s�a5�ָth�C0.K ��6-�O$�>/ޥ�S���'o��'���c�V��d��:-LcR�w�x���r��4�'��	󟴕'�Zc�x �E̋K��tc�z���	�On�z�0OD��OH�d�O��d�<� /���h+���&J{�B1l�k/T���^�|�'��^�x�Iʟ���������E�7|+0쪠`]�Rx2�`0?���?I���?�.O��0�N�|����a		R�v,� ��'Kæٔ'��T�������ɺ��3�pu��E>"�0��*?Ԩ4[�ON���O����<I���o�O�P��>ׄ�H��޷Hf0�b�ja�����O2���Z�Gf��>��K� c����Y���ZtGC¦��I�4�'�r,Х% �I�O�I� .
��D�}�Q�aӧ#�8]o`y�_�,�Â#���4BV���Ȃp�$���G��Yo�jy(#(�27�u�D�'���@3?�����f�͈�,��\<��K�Ŧ9�'ut��P�4��'�4 W�RK]K�g��P6�p�شA�PU�W�i�r�'�2�O<,O:�d�5�,(��P-���G�Y*7�x�	0'`#<�3����*��@7`� �F��l;DqZEl�?ntପug�^��̠�'���J6��5i_NUQ�׈Ax��[���܂��#c�lt�1�1� �PaJ�v'�I��OD��A�B��)��6��)��j��%�V���cO�Z")S$JO�K�Ȅ���K/^��0Pn�%t	N-|$�D�!cS�M����%��W��db�L!.5Z�
�\�A���E�Y��Ū3O�L��� �[]��	�����՟�*���|B3�K�&ŲY�VV/� FlO!i��p17E�+��A��/ߺR������-�2�(��Oo�X�E-�&f"��:����!�Xq��?fF�,KlP�HO<��'{��'�\�+1H%/
�< ��^5�ў�F��U�s/���7���};)�0e�<�y�G!v2^9�F h{�Vy�W�_:�y�j�
�ľ<AD�ɢg��Sퟸ�O�U� F�1�~���
r쳆���>��'�!%Q!�1�b�J��Y�G5�-T�0��&�%5%��2@̟���<IcgW�c�p(�%F=D�0CL2��']8B4@��T�йh2�����K�'����?A�������Lu��f�7$\U�!W��y��'� �s���F�H-*�n�'<ʠC�O�=ͧ
�'��]�ԇ�(a*���<`౜'�*�Y2�r���D�O�˧dH*xK���?��E�l@�f��4F4�1��Xk.в���@�<; t�8䧑o*�2b>�$(�{�ѡB�ə#"�@o���E��0���	"���	8Ix�r3��w*L\����2-���ge��2�"I�r�'H�)��/���s	"��5C۽#V���NZ�L�!��29�6�R�A��|A������X�1O��dd�����'}.���IX"��hsA��>hDx]�F�'�B�O�n�5�F�'t��'b�v��	ٟ�˱��\�8��U���;����/���S��X�%RE�q��p<���0.�C�ЀA0�IG�TR?�R�V!�F���&"U��x`��F�p"��'q`�I �L8�~���?��hO@�7�Z��+��L��ӰD	;W[N̄ȓ-D���J��O�q3��9~�p'�i>���Ey�)R1UX7�\+��x��M!�DB#Avw��D�Od��m�P�p�O��D�O�L�qE>:��$N�zl|��"�L�3eݩR�|ăG˂}�0�A�? �Iɑ����a#'�[&����Ռ*](��$P-!�'�ⵏ����`��ܷH�(�Ҩ0���O���3�)�󯗏O?P��]��@���Q̓ig�Ex��$KŔ_hT����� �l���yr�v���$�<y��ڸI5���'�"Y>�5@ጴ�R�@'Pn����1O�l��ٟ����	��p3bLL�$��Τ�?�O���34��\P(����^ VT�����#��h2�j#x>�l343�錅O�I)Tg�&X�a#Q�uQ��jQg�O��}"d�K�E8袢���@C�P�<�3���!���:�*X~�@�1�I�pO<a��29:pr��=N�Z}�1��<yƉ$Up���'pbS>��1����	ӟ�fN�>�}JӤ�}� ��M�LJ
|:��P�4?@p�����<�O�1���L~0�wDU%�.�􉔓}�J�I����J$��"��t�9��ȘN�s����pΰ�n�`���`𢄐%��1�,K1�?���?Q������]UZT�[��B$k����y��'U�}b!ԗx�i� 83x�Y�鐽��'kr/��|���Y���)@�Z�nȉŀ�0,�����?q(R�F_`� ��?)��?�ո�����O�}�F6 (	ꥯ��c1l����O<�p�'+��4#�?�ea�2+]�En�c?1�OYx�t�J ?�ʄ����:N�&4��B���1T��O�����$\%��P�HH@N�S0!\5r!�$�3}�z��V�ɷ0�`�ˆ��,cd��Dz�O��'���R�i���K�F�(M���V/Q`Š���O����OL��8|N����O瓾f����O��h�ՉLC`,#`똽W�l����'��)�*O�e�	B�GR�2�CIO���c��'~4���?���,I�<,��팃d#��k�Iz�<��L�kV�a�n�'���T"x�<Y�(�%�R�Ӣ��[+�(�#H��<�����4}b�nڟ���Y�4!�LQp�Q���Ƽ2���P+��¤�'O"�'r�a�d
�l#��O�SW�DH{㥚�1,Q�"/N"��<IS�\W��2��T
i�QR	ù�����l��� _�dഴ��ЂE#Q�0x4�OD�}�'	99���X��)��I�<�sD��a��Bfl� }�0 �%P|��K<�2 $5��c�� $#6
�<Q�%�=����'�BT>�G�Xϟ8�	Ο�S���
�P�&j��8�u�cػ6n (�IX�S���W,
��$0�-@�Y@.h
��Zo�z��C	&�S��?T�K�b
p)�+��m��,�@@ϔAҴ��������bl��D�&x��g�%]����F��yra��: T<���\�U��0��M4�O@�EzʟtaӃ�F)J0�RP�Մ`RTI˶'�OP���%G�$i4e�O`���O*�D���ӼF��)��y�&t�I��Sc?1�H�ix�� �@7F��zCoG�����e��,��b<�O�L)�`Nv=Z�c��O0v�j��O,���'6�{�m�7AT<Q`n�E�ɢ�a7�yB5?,�Z�i&
�E��.���#=E�Tj  "7�@�H=�䕀gh���I�+�D�O����OD��p��O��Dv>��5��O�����=�v� f�
���J"^��|B�����v�P�ڙk�d�6
�v��|����?���W���"f\[�Ҁ��n>j����a_t���@� Q�Sf�V�}��ȓ'��U�O Sux��O7f��ϓ ��O�����¦��Iퟘ�OpJ�R�>��L���;00Fhه���^�B�'��
I�H������|�*P�|Ɯ��B�:+���Q&a�'&jĻ�ݜl�vq�шI�:^\��?�"F*�B�D��Am�@�I	�+� p�����x��4�?�*��ᅫ�d�* ��?�ڝ�'j�Ob�"~Γ#|���ؗe5�$sk�!/��=�<y��V���Iџt���:Cʉ������t�@��$��M����?�*�P(��(�Od���O���ӡ~n4���Ih(a)��� s�q��	l�t�S����'x)�6k͸g�xq����2�����ޯZ�DB��7<�)�矘�s��2���t	�8Q�PɅΐ�>6ZI��.�M�5�iV2��O��M�0M���꧂���<��9Ol��<�On����-�p����J�@�CQ�ɷ�HOh�[�'-���D��.�ӓO�#����:*j�O��+aA��+G|�d�OR���O�;�?1��FM\��e���!{����@Ǚv��)��ɰk��zqAL?jt��4�V�剽u�uzs�.,d��{��;���r�+=)��Q�A��&��d�r�?�Ў�� ��s�fԛ �HUP��Z�}H�����OR����O����O�Y�<��Wyr�^�EWt���]F��KZ��xb�'d,�cJ�YC��ap�\�o��B"�9��|�����MY�l�#+�,�U(`y�=�u��[r�$��ҟ(�����c@I����|b7ɕ"5�N��C+_e�� �@�F��́�� [ܔ5�R$�:�ay2��72���Z�wI<+5�03l����HL�C��$cE#e/���ј\�hf�ȝHӌ��h� �*E�<��d)tA�O����O����O����O����d�B=�)c�얲��8��A�W!�D�:%����aG�8��;bW�sh��R���	WyB`V�t�7�O��D�|��5nB`���߄�6}�#��/:�\����?���fiJ\����[#���S�[��7]>Y+UX�xpQ�V��A��9��!�E���V�չh7��0U�	w��z�Q.[�fR�q_��Gy҅<�?q2�i2�'��>RkNY�52��	��僨L���	�,�	��i>F{!%2�f �9lmt=He�X=�0>�T�x�־3��@�;_�r�2H���yR��.U�7��OT��|�3���?���?��X��Cp�$7��跠LQ�ZA�oD�8ɧ�)!��O�	��^h~�E����T���[�0����]�)�矼�S�G:�p�(P�\�~?,�x�-�=�zd�I�<��͟�E�����Z�D\���t�3BPYϓ�?��i��=[��E�9L,����"ΕEx�+<�S�T��5]ℍ[7�P Ix>��H� ���D�Er��2� 1]��	�D��4;!��Z�e�@ ��ss�H��ӏO�^B䉛FU���G�^���^?t^B�	/N=�L�ji��8�R�ئd��B�I�0R������aSf� �c��цC�IY��'e�>�R�����cSLC�I	^]�a��?MJ�(;��	FC䉂=�h�w�\��{�%͋^�C�ɏny���e��1�����M��B�I[�X�{�b�"��0St�
�q�B�	�mT� �	Xl�����\��B�	'6��0�2���K��������b�C�	e��0�EU���3ክw��C�I$P��R��Ą&�Rq{ժ
[��C�	}�E��@�u]�%�@�I�'�C�	!;ИS�I9��y	�C9zt$C��v�J}!��='��s�m��L}C�9f~r�`������%Be%��yTC��|�>1�7`Q�<Ӡ��C)�;y��B��x0,���\�2�9f	�)�B�ɨ6��ڄCD&D�\�J�ͅS�B�I/��m�8�6e�P�
)A�C�I�m��8��M�~��dj�*VU��C�	<H(` ���&A��A� �T��B�	�5bf���n5�)�vC�))ttB�	�M�.�b���DRbx R($z B䉡Ya���3%ץH6���F��P��C�v��ɠ�;7 v(BT�nB��0A���9%�C}�B�*u���B��[Zx �� ԓ/�Ү�!5n�B�	�@�h|8E�͛F��2wb>m�B䉡=�\8�v�ېE� Ҵ�V�(�B�S��\8��^"�D�Dd.��B�	I$(��/�}�����@�>
LC�I�zH���f������/D;D|PC�yUV�� M�6�
D!�0yTC�I���(�VZ��,!�c��� B�	�L�ҴI�rg^̹��GژB�������L�#�B�%�.#nB�:C^.zU
X�:�+�,ܮq�TB�V,�ȃM�Li0�R�dޮC�B�I�b�6�3�� ~,>�p2�X4��C�ɓ�N�OV<i�ݳ�ԥ	7r�'R�<�c��� D�('����жFV	 �P<h�"O�H���Q�Mx~=ӣ̆8`�f�9C�'�
Ś�'�� �3+�y8��;/CV+��b�3ud�y2�?|OHǦ{��9'��j�"�N��/F�!�9>��!Y�
O�Ȑ hC/�$H:��V��z���U�$r�ɦ��H�p���	��SM� �^Q�bj�7z!��",�L�K�dK'��u��IK8h� ��;O�UrN��yB��
#��wr�Us�/��BVb���6D��Pq�A���x�� k�f\rpm�O���Io� �bd�GW�x�`($y6��$�*��Dm���=�!"���y�hdlY(��˫[h����9�,@��Ȇe(<	D+ݣ� K�F' �, ���i�'4�Yz�'
�C� \mܧ=��%{���>�f�a��M�\�ȓ4K�TX�j@$�V\y��_;$}��'�d���&�_�S�O��XS@!H����A��sg#
�'W��i�M��pX����Q!(*B�C�y��Ah�Bԅ�I�}�8sqd+u:��c	�
'&O�u���"�)�)ߞ-���C��o�v@�F�I^���`��Px"'��$�2�P!
I@0��Γ,��'�A2��޳��d&	C�
�=a&+@�2�a�8O�\��pA�n؟h��DFnպ|�ӧ$`��BE��:#v�hU��7^K0|H��	��O>E�TΜ:x���h\?J���2�� ϨǪ�������'�`�)�, ?X|��lV3�����)z2�'�M!��˛����O~��f��90 ��Nn�
>O~y�dÉ#C✀K��� ��> ��3���C�&Vz�(i(#垽(hԊG&N��2��W`7�\��aX�΄'/�H��1O0�x�Ӓ7�<x�;i��!�&֟����hD��,j�D��-���KB��K��$#��U'�����(��W@H�;c�	~ |h�wǙ*)
B�n	5�`:��/Mv���(��|�4�D�%	�#h�j���"V�� ��oӐuk��'�>E�T*L�R��S�	IW?�'&��4�ጘ�-C8���;!��Mc����l���(v���f*&�l!r�O�U<�ǋ�;'~�
�3}��E	�9<���w�ד{)���&��ʧgwR�1��h��y 6 �2L�`ٻuN˞e�
��|g���e	80�"<����_�'�E���;MN�12��#d.��I��6e�(���'� q�-^�UX�(a��f'�)�����c7� �Y�R#�bl� %s��y�(\�1�2}�oW�?�Ӈ@1)�ǍͰCp���_�[�4�b˃ E�\��#�a��6�(@��?�S�
���Z���?Q��U�����3��<���`�)~��X�w$Ю`����G(&�)��ş�. �ޡ��DBqI����>$;�� 6�O�IF����rΟ�̹5n�C��Ւ7
ٻ\c���.Լc��yDN9#���1�@;)jB���O���
~�a"E��V0)0E���MS��_��p?S�T	~�d��v�$O���G�Op�H��I-/�a�(>��5��82j6�
�?�i��	 �C	m�����G�}�ĩ�A"%�O�)�F�.V���i@��A��&��-҃�� %/��$����5�O�C��ұ�OTԽ珞�W�Z�k�Lݬ.�H���	급9��c/:��������O����p�,*(��et��+��I~?Ae�4��)��Oy����V��rA�Rd¨Nr�ZQ��*�nt+�'&m�&�� ��U��!�6�����N9/���á�P<U���YW�"HDĔ�B�\��~b��G����QX���'�4� �y�[�p��A�A�:zAA-O��������
kB���#F5,�@U ��'��`{ ��w�p`�E�#uHX�d��8z���L$��V�E[��+C�O@� e�)��O����e$��Hhy���R�+� �
����x|���X/�	�$����OPv��҄O4���(gO�_>X�:m�J?���Wx����Ŋ�A���$Ż:�^�0�cɋ?|�P1۹p�R���+������ U���	������$ʶ}}�m�u�]cb��J� W�ׅ̖=��l�q�'0| ���Fl�ܠ��� M�	�'�?i���-`~|r�¤��?�i��A-3y]�Q����21}�8&j&�O������⡈��s��ey�O�.q* �5]��;�R�����P XVt�	�l/�h��i�!Gf� w��#���kr���'�P�T�Ԛy��E�ȏ���k���O��6��x�cY�1����d2f�a��'Kb�3�.P�d��0�˟���vf!E���Jq�?ߐEo��/.���S�� ��$���~6m!��H���ɜC{��Rp�H�W0��G���9�oE׎���b�x|22�؁y{p���
R���D��,K�f��h<+%0�{� ����g֋N	��S��'p����ȏ5P2����F'~�\5��d֠��'d,�1`Y�c��A����|T���%��Ok(��`��z�fN4z[1O��:QboӶ���(��!Tࢼ8Uj_�~�T6�2����Uv*j�/C�r�Jd�T#��zQ����B�2�%�Pӧ�^���P��� |���J�^�!1#Jj�k��^)=��(���8R��Uũ��F_�Џ�$�?(�a�J�g�A��b�5G��O<����b��s��%H��I���J);�i�i҇���_}h� �"R��
2!��=x�X�	˓Z�b"`J@9M���A&L�Kr�Yt����9��M9 J����!��e8q��/��C�\�֧�G�yG<�+L��5�2�b�B�Ȝ=1t
�"m����d�C1tdZ5̎�`�;���Z��>l��ȑ�f�h�bV�cM��BZ��	�yxڭ��@#T{��R*W,�ᘃ�ͺ9�	c�60Q��XC��b\�A����%���aa���DZ�Q`F��m ��'"��@����۠)�Շl��Pw��9u`\�Ծ��P��[��(��r쌣z�.Xh�I�:s�4�Ϙ�dզ�#!��
__�7m~����
�||��,\�2$$Q�I��	��u7 \jJ p��Y,O}����jE����á�'���bU�A"�]2_ؘ;t��6s�
`v!�(�$���#'
i2���FW��K����B��\
"z���5�� q�� ��3Kx�jt�#�yʵc4�8��]2�� ͺY���ȴx��d��X�pj��Z�.&Ţg"Ä%~.Rn���vhB:��I;d�Dh@�E1(�P4c$��jֵAD�&4z��*M�f��DՊ ���Ϣ0��ȂG�ّ;�`�Ӈ2y>p,���84���`y��!��7�<"�=��M�w�����]d����c~�B�HH�=�ɜ?6���x�+���*�?)U.��v�S�E��)�W�E�+!b��V�ɵ�(���N�V���8%H�Q��MW	,<�-P�Iމ�	��y���qP$��eȢ��?�i�m(�n%~�PQ3�%V:F;t�;��5��.a��c���m�	C�IB����	ܧe:
Tc�ɬ$�Ot��̦KF���`�:���DG�*� 9�����(�FC#����'
D��$��">�452F�~y�b"�d��|�OD��˝�N堝�S�ۑ=�i�P�'1���Pʹ|���g�&I�D����cǮI"P�I��<��¯��@�'���Ƨ�6H~axF	�?����Ё�+���ʉ�~�����G^�'ܮ�@0�g2����6�^H˄J@u?�hBN͒��ha��5|O�-[%`�%��L�0��z�N� Rr ���0���\�l+��[�s��	��ēd3���j�-!\��JT�nK:�D{2*�,d:f�ضM[(�v�ѯ˲�~2�X�(�h��"M�G;B� �ڮ{��d����h����t-�
�2?��\�d���▚r�d�*Fh��ҵD�),�n�+�CV�"f!�� ,�Sx�)AѭP̒�]	cqV�# ��Iܓx��B�'�>���m��Vء� \��x!rt�S�[��G}RH�=z����$����k�!�.1E�ۭgt���.)1�@M�X�'��B��*f�~��-��.pH�;�:�ȕ&�=F���xW�1�:��<yS�#qf:�������a@��o̓q�xЃ1A O�X�%`K_�����m Y�E�*S"�:��ݘ?�����(�,H��-�����	�{}���ӷ����M_���'"�;����×�������D]�?�z@�b��cp6		PI�$��5����iFjqy�o��D}�eCM�b����N�;u65�͇r!)�)�O��f��?��E�5��(���zg(p�uM�.����6% 2�#S�%2�����RA���Փt�H�A灉N-Q�l#l+^�P<K�4\����
�O:D#�����`dR0.B�P��dBn��R��SR�,A{D��M�1Ov���-QR,�WV�.J@���x2�����T/�:=4�!�P���'~:�Ҏ7_�����A*]�Yp⯓�om�p�Q��..�� �L1x���K<-�|E�B�N�`E��( ��ц�G�j����j��K5"�/.o�I�H��a,��D]1+?X� wl'C��Y���YN�.��~,�Y�$'�X�Ŋ�W΍h��R�"�L���,H1y1�'O.�(�����P� /�=X���V�c;�ī��A~f�)F��&VKqO���k�e5bم �>�I>�3)�Y�@�&n�G���3��w��n?7���xr�!�4/b�OX��OZ�lT,Ei��=?�Q���	*���
Y�Y��h,;��ԟ&�;ga�nuʙ0�@�|���1�hҝ3�&��R��)SA���	$�=����^IH��#��Rp�A��#zk��⑌Ԭ~r�\"��O�3��������*!h93K]���#�"O쉩G�U�:��q�H�=�H����:t��
]G����l����E��ا��`g[#9������H
u"�I!��~��EE�L@�T����CTE��	��J���b�A�,����5LE4�`��0��#ʓ, �U	��69��H6��d{څEx�d_�p�XA�A�3�r�9�d.�?�'t�$1�l�+�����=*tY�ȓܠ4Qa֭��%8;J��8�Z3u�f�xe�KL� ����ȮC\�>��?u@����:�X�@��5 "!�䏌L�Da�M�1��-�G�ҏX!�Y�u���7��%�z��E±Z$���4���2��A�S�����D�7�yb@̖},�m��� Q�ꑪC�E(�yR@�1 &Ű�UF���0��H��y
� �5���)~0D�ц�A3u��S"O��X�-ޛ<��۱"�"DW$Q�&"Op�ݸw��%�/�=jGZ�X"O��� ˉZ��IHTϑ�EH #�"O��D�N	?��A��.!Y��"O��j�c�l4��-�5V�ec�"O\H�&�߮e1�c�W�;䦉cQ"OI{eh[�{L�҆�(���"O���CO	� �����/�0i�Ÿ3"O+#Y^L�P���U`��D"O�Fl�$*�<0�@�
f����p"Ot5@�iߟnhK�AZ�
��Dk�"O�`)
{܁hԪ�� ��"O��@v� �H�ptɗ���} �"Of<��Ǌ�8�F (��X���S"O>�
Q�Ҟ �@	�c� 30j4��"O$A��	{<���G��%vC�"O��Bȇ&(��C�
;Gm���"O��*��E
an�t`�`�3b(�A�"O�h��&Ջ]�dKք�C��c"O��2��=��U��-ހ})Ĝ�Q"OB���!�3_J��K��F���"Op��3��G2��q�Üa-Z�"O�	ゆ]LW&��ၐ~.n��"O,3b�ؐJ��e�t�Q�_,ru@�"O9x+:�=��/ݱG�c&"O� ��"T:;�ڤ2�/�gҁA"O�2&ET,W'� ��olI�"OJ9�g�Է.~}3BGӌ|;��ۅ"OA����))2��cFA�e~�ѩ�"OIg��/���yǄ�Vj����"O<���i�+Z`�"��W�u�"O�go�k�n�+ԠCt&>Tx"O�����E�*��Q"�YXc"ON!�5F�(}��C���w�D�T"OL�1�fMN�h�#������"O�P`�KT�\��r��ąm�p�"OX���" �|�u���Y}{-�"O*��f�ұ4��!!6�KT� ɵ"O����È'2m��yP�	'r+9�"OX�j�ȗ?`�ɣam�$4�T�!"OtuzѬ�Zwr]k��S5�� qe"O�8�â$��A#A|�p�s "O��!bͣ�V=�G�ǵ�Pԉ�"OqBK�r#ʡ�挰X�N) �"O�X�"C��J�JP0�g28���"O��S4#��k\dp*e#�,-��#�'l���ߜS�p��N��k�%�	�'���iL1�j�k��N�xO��'���FتC�tJ�#m�qJ�'r `�d@Lq
4�� J�_H��'xT�ƂZ�[�jp! �(�)h�'u��Ѣ�
D�8H�Ʀ�)�t�	�'φ��t	�-ۢ�sl͛y���(�'� ������D���#�c�j2�U��'�tU%̆ Hb�iq�]�b�by�'���7�
!&�Ic1�_�i�
�'� l��Z��BσZA��'_r���Y,(la�An^�O�L���'��3�G�U�,q��L�A�*��'�`����&/�-�g��\	�ȓtʆ����դn^�U�X]�9�ȓ.zv��Wnr���`�U^�F���gE��OR	v辑��R�9(^���S�? V́'�-�@-�5ƌ7~�0:�"O`��Ao
f�(���_�u�"O�8Ap��+Ơ���l@�tm8�"O�x8�o��[��]-|T81�"O61��ώ���Q��='7�@a5"O�5�sA�D�f�s�HY7;6��7�'l!�XMh��p�ۄ~��	6c� �a|��'�d�����x5���I�鲒��?�!�*-AF�-\=�2U�a_�p�OҢ=�����%B@�}��A�ѩ�C
vl�"O���� ��a�����n��SBT@�'P�>�I1 ׈Y*C��-�6=(!�L�oNbB�I�9Q��'��5|2ݩr��Xb �	l��� BT���5ʓ�O\�`��!D�����Q�T�|�`�M$=�x�0�9D�P���˨.�L�F)��j��fA5D�؃aB��@-�݂FR#���(D�<+#K�#������0@��M�S�%D�`@8aZY8�
G�re��N"D�T�+�=SL��&.I���!� a*D�<c7�q#q��*/`e�(D�DsC��/_�����vu~Ti��&D���S+Y�V�`�H����c�!D����Ӂ=�,� ���C�}`A%D�l���Ͱ��!:ӀΛQ�r�Em#D���H��s�<A6�ʼc��9��"D�dsFf�	=��g别Ħ=��*$D�9��4G�e���Yz6t��c"D�Q �-�xx��ʃ���5zP?D�0�E�1*�
�ϟ6���Dk=D����L!)�X��7`XZ�E;D�H��M�K��D(�@�>h���8D�0Xb�П7*�����p$�!��8D���祇;_�� � �ӺK�DXAw�4D�X����:˨D��-_�;���&�/�D1�O����:;aq��G5P�[�"O�ɣT�R8�n ����::$b��"O�uP�J�9\{tg�24�j�Z�"OX��1T��}X�&����C�"O��c0���R�P��N�Er��ز"Oh@*�`U�l=����'_**�"O6x!�Z�6��3A�O��"O! piT7i�<�J�Ao`��9B"O�Y*% �0X|��C��
L��w"OR��� >RY3b��7`E4���"O8�(v�<mu����g?j9
�9�"Oĵ���ʣaX����`�8f�vx1E"O�乕bя"��3��ַZ� ��v"O�٣`A�r/j�r@��5Au���p"Op�;ҠT����"�2F�N���"O�M�AgT$q���Jv^H���@"O��o[����C�'���("O��yF�.�t���
$y�0�06��܄�	D.���a����Q��5D���DÿA��H��#��[��b��/D�8Xӆ	��L������R�#D�ਢ�Za\3��Hn΢�n D�)V��3F�Z�qqG	(4$���9D�ȂҮ؜R&P���ѱ#�aK�&%D�P���
��RTsB��e��A�#J#D��	'o.eoB8���Ǜo��c�"D�,�G�ĨW��(P�ƍ8r@Ãh D���'�b�,�����=���L2D��Ƃ��|�� q�Bչ�L#D�� j�"֣MW�n�;c���=�S "O�,��.�"\�����,�\��"O8��c�9fe9��Ño8��"O6�Y���E����5&K5i�h�HB�4�Sⓔt��(*5�Ɉl�v����E�B䉥%��0 Fl"u�^�-d�B�I+�t�r'�h��k5�ܢtw�C��	�h�3kʪG�銒�Z�}ọ=Y�G.���1���\B134Ά-��p$��F{��DJ��0j���	WM��R���y҇��u0�t���O��H{KX�y"@�8c��XQOڍrFv�$M�)�y����$l��LF�ZxJ��s���ybfT�h"��q�{^�l�	��y���*wh9C����^x@0�EI��ybE�1D��YS@�S��4��AR��y�o�9"
(�ve^�a�&$��G,�y�h�2'���6j�ST��L��yBj�h��PE�ׯL)��8�"N��yb_��ٻ�ɝ�BAB���>�y��>`_z��֫�;g�@�c����y�'�&h�u-^0,�DPӒ[7�y������
��zt�Ñ�G��y"�	7Q�!�%�yĨ���Y'�y�E�P�T��e�<���n��0>AO>A���j�� ,=����O�<&���t7�m0�-�z�Z��r�	�<!�}��d�X�D�l�������:����?��'պ�Id.�x���X����@�X�	�'�
�i����#��!đ7���'NV(��1�J�z@�}���S�'@*(�"��l��,QEC��t�Z�h
�'܈�!U�M�[�2ܪ��o?���'H,�!'\�~X�Ӡ�#mk�I�'Y$�%iP�~�dQC(g�`Qs�'��@-H�#�5Y�䈥5�j���'��lA�	�%3l���-���U[�'��e�ʴK�MRh�F���'t�0TE ����өo%��
�''D�*F������刎-v�
�'a21i�s�>E��N����k	�'���	�>:N$seL����X�'C`mJ���z� Ї#�	�j���'3�Y���\�@�l�O���'�X�!��)�v��f�Z�IC<��'*J��W�F�L�K!��M|�̫
�'���y%B:!ʩ�M!=�8	�'�d�#Z��q$�ؐ�;�'c�9`�\�^ ��n���p��
�'�L{C�L	m`��	��քJ���
�'�̵v��eN8Id��E��5�
�''�A�)�J(J�[2���B
Q �'Q̭"��>_��<��+�|��'4N��B�*!�X�A���z<PG�$�S��?����@���`PHވ}�ó( s�<9�H�'\���AQ�υoj\L��v�<) ̓!�� ��D�5�-��DMG����<1�ŏ	*1��cQ�2d��4��@�<�g�ܸ4�bc�"0 ��AE�<A��܁`K|@�r/�4H�%	V��C�<)��A�R�X5c��ښ_8�!�V��K�<�pjϖdw�L�F�Z!Q$y*��p�<0��w�d����G(+��U*��p�<q�E /�SGH� ^��ki�<� �՚��P���d�g@�S&��5"O�!��G�'�J���L#�6x�"O���FG#Yzy{V���?�ћ"O���IO86ؼ<4���=Ίe(U"O�uIr�]v�0JC-�6B�"O����Q��xx��i�w��"Ot�W�Ά`'J��(Ԋ\Ǥ���"O�5���sX9�G
�:X��"O����gt2>	����<����"O��
�lNB���K�LZ3t!"O\�X���T< ���45��"O�Y��d�'@[�P�hZ�m����"O ]���6H����� ��+b"O�
EČ�2S�ҡJ�:���"O��҂F7Jr� �KR�|�l�"O��ن� ���Q��
�o=&ᢗ"O�����I� ��$7�%�S"O�ŀS�ʺ�����c�c2��3d"O$�)�gH�&~�1���]'��#2"O:4�Q�C	x=�� �n
$f�J"O"%��(	`H�-�J��)�"O(�h�Ā	s�*,�%C�� ,�(Q"O��9�cZ��qA\�Ԑ�
""O���a5YH�#�@�A�P� "O��S���-��x�֮�)(e3e"O t�w�� a�|�J�M	(r.���w"OlщҨP�R&��s�lܒ|�ɋ"O���W��rt���܄t�r<R�"O�
���w_>�Q�R�D����"O���A�!r��Y�@D̠/�}�"O����@C2N�<)2�����%YD"O�Ƀ�e�0s�����\����5"OB������|̭��MƎm�f� "O�h;��J:_�-C���?�Bܣ�"OZ5╘yb6��,�>pi"�T"O�I�&C���L���Jr��{�"O�}��dI��*�@���H"Oʹ����`x�5�2�144��"O�h[��_L�p�
֤)j\D8�"O�-y$���1�b����k:\���"O��$X<��f]�)9�Yr"Oz	ӷ�����k'��"AQ3"O4�:S��'%T����I�(m�q"Ojm˃� 9Rw�lᦫӽ@��eY�"O��+�'zj͸������-��"OV���-A0���TL���6!f"O��q����q��Ё�ҠY�"O�ٓlۍw�h1�%�/���C"O��˒��wW蔺r���J�Z *P"O�U��x�r��4K�B��"O��B�&��((4$߶@���C�"O�¥_1S��	9We��r�! "O�i`���5X�(T��%LiB"Oꀓ�ƅu�R0kv�+)p&s�"O��Sw�]�Yn}I� ��3Rԝ��"O�C���~bֽЂ��%r2�|q�"OD�R(Ό"<�9 �4"Ot�����@mnb�O�~M��"O����T�.O��/�"����"O.��q�[|��΁4�II@"O\��	L!6��9`�(�.œ�"Oh��ǭ�R�D4��m�>���"O>H�6d�8#�v����s���ˆ"O�p��향t��kdB-fl�
#"O� �݊�(]	8�ʨk�"%F�ۂ"O�9��^��Q0G�	�	�I{D"O��$��Bl����ؘu���"Ox<i%�����2G� S��M �"O"-�b�X�?]��X��YN�xz "O098�,c: �넇A;+l̘�"Oִ��鎍p��Ib�C�J��w"O���2�U/���Ѣ�9��h��"O|u�A �;e>�}�����i�"ON�3۫s�p(�Fo���w"OF�f%�xw���pJD� ��\` "O���ș�hr�D!v�� �D��"Ol!��j�˖Ѣ�(
�\8�"O ���@35�:I3���T�2"O�=�F�'Q� {�GE�o�^X��"O��C1�'r�ΐ����L��%r�"O�U q������B%�Q)c-,�)�"OP���O9?_\S���q�H�"O�D�@�!+�U�r)"B���f"OT�iAGr��r��9	�Y�4"O���-N��4
PM^�Z}Z�"OB��%�8JX����L����}q�"O��ȷ�@�D�p�c ��xg��"�"OޑB�j��0�F�s��R�:R*9�"O�����#K��E ��8c���*f"O>$�@�V�|\"a��/�,N�f��"Ox1�fGB<`k̑A�.��srF]�4"O���`��j�NբW�Ta��S6"OHHk�F(�� s���bx�"O��%��h� �x��B����"O|]����e^�����,)�ji��"O��%���]9��X����S��t�5"O��!�c&@Q����L���"O�e�#R�i���[S�C����"O��)"�yJԕ����s�|p#�"Ol��@J�*�tP�E�P[Z�%"O,��!�[�BLF4@�h�	B�]!t"O�4£H�(�����W�n�$"O�	��Q����a�0
�u��O�<��3�2P��}fd��-Fq�<yv�E�0�Lyģ�%�QI���m�<ACb�'���T�D%S%��7��i�<A��^�M��Xs�.ҟl4PF�d�<���X� *VĜ>u�MrԌVu�<�4y�A�'��/w������x�<�f��PBd��D����� b.�v�<����)K�֤�Mɟ$UZ|"L�x�<A�D	'�����g.����dXo�<�D�58dj���� q�����(�c�<91���&	Q���"3�%�a�<��䖲e9�D�qÆIB`��u�g�<�gM�e!����]Ta�Ax��b�<I��цG
nU���T���Uci [�<�`k��.�$��Ą^N�ʱ�Kp�<�2�Vg]0lC���of��F�Tk�<QvLն:�IrD��!yx���P`�<i����5�0"��K= 8�C��U�<A ��J�ƥӝ_2�]c��S�<I�k؈/���a��#<�I�"iMN�<Y7+��bΐ��1&�^Y�k��_H�<Fg�:�`RdB�rU���G�<�@�O�"�f�30Ύ�S�2�*�n|�<��^snRa��e��^$=#��y�<��n��a�����:0t ����P�<� ����ܑD���1���E��8u"O���%��Ut�}�f#�*�rq�"O��S���5	����"z@L"v"On@�ᑅ/l�=Zf?#f� �"O��� Ǿ!��e��#�t����g"O���S,��h�=; �I`�Ht��"O�$`&	����4�Vb�<����c"O�y��埶pu�%�C��1��8��"O�����gX+"�!C��P�"OV���ȮK[阡EP�/"%3W"O*8�Si�=h����N(��0�"OX�)$,ڪPc�٪$��'&��̉�"O��#�B�qp��byx1��"O�̎�*qnӚ`�yq!b�Z�<Q���*���0���:_���b�q�<�V<�L2e�H�.Y��#D�,ᕤӛH�F���A &܊��$D�I!���Du1c�]�T#�M!D�D�qf��7,�,R�&\N��$U�*D��:Һ��h��VQ�Mr��T(!��@�s�|�$-�5y�u[�EL�C!���
}X��tG�Hp^MA��$!�^�t�8ʑ�ϵ3Y&`j֣��U�'ў�>U��g�)e��\��`�!-D���
�2�B:�&����#�?D�lp0HE��-"w��Ng
Ya,*D�P�b��~٠ܸЏ�'2�,B�E(D���ł�@߼���܆4�΀��+D���$�@�E�j-3���*�@y�c(D����,�����ءi�(h�˲<9���?�9�za�F%8�p��e���D��ȓ�L��J�'�V��`Ǉn>,��h�`I�5cD�t���p�ZIܼ��ȓ=^�+��h��ḇ���7-�х�Rp���E.2��{ ���ȓ&
�x��5�$�D��YkJ��ȓN}HD�ɟv��%���ĚQ�Y�ȓG�
��$Ӷi��b5��Y��ȓo�L��f�
4
��x���H�z��*��C�CP���SvN�c�
���r&J�h�A¿�`I����%� -����8�<q܀MG�	v)4���	_~b�ݿTԴ�tHP������\.�yr+ݴ�>���c����!�̄��yB����r��RBnpP��1���0>9gf+��x���g
>���d�r�<�����9�g� `֑�s�r�<���jd݁�,ѷK�H8y!�f�<���V��a#3�W8@�
��!J_b��x�u�ܱ�bΖG�}�"a��~��ȓ�v �E�2j8��i��8�(Ѕ�A����?���;ąX�X��%���IB��`ҁ�[it�d׺)
��g*.D���V�4���wB��p4��&D�$I7�M�=��hPW"R'Xmn\㥬%D�����<U%���ΫN4�B�I.�O��	^X����ֺt���a#
ܹQO�B�I`f�I֩RՠHz��.N��B�ɴl�e�@,Q�h��F�B�X�B����1ٰ)� ��|8����H��B�I=nx�i�o�A�~H��i]KڀB䉣��BՆ��9#�  �.ϔ>vpB�ɒ`��x�S	�W���ij��D.扷!܆i	�`K�k^P�0��_�(���;�� ���*�lє�`��ۃV�p��"Od�Tf<������4-�Q�"O���g�^3D��0����N)$m�"O^��fZ�L��]�q���z#��`"O`}�c�\��\���dP-,��x�"O��t/��������G���O��FŐ�=sf�RVn�[-�qĥ9D�(cc��=(�M`�܍V�t�C�6D�Ps`�t���a˛g@�A�&4D���i��9�V��� �(����'D�,�P�T�E7�7�����2D���`ˊ�� �3敯{��+@&6D���DS[�d��C��n^����'D�D�t
�1nF��E#��v�I�B+'D�,"aJ:1�T���mюI~U`F�$D�� ���K.���g�ҒkG\1-1��O:�=�O��Ũ�®Z^ ����~y�"O��+���F!�B���l�B�f"O��b\r�Yz�k� %��yC�@��y�aJ6�|�	4�K��r}�E$Y�y�o���9�@	'; ۴aR1�y"ލ����S"��"6�tj��yB���/�ZI�����0�R���/K �䓩hOq�`�K���v��0Q�Eʂa
ܳ"O
dx���,�v�����=`Z��"O�X[e� Հ�C�VG��H�"O�X�х�;�bT�6㐮�4���IS�O�衡FU��������c�����'�F<Z�g:?y���p枰o��-�)O���#�O>�p�g��.�"2����9��"O�4J�ߵ
j�����i���"O� C�׎d��\���5q5�%�E"O�肢�I0"u`�)���a�.��&"Ot ��+��#̐�S'�jЊq"�"O,�JQ��7Ԍ�BƐ(�4��OV%s%)ϋm��5c�=HN- ��O��d�O����oY�M�pGӷ ,��cXz�ń�5�p�घ�}�����	N&L�@<�ȓkjQ�wOü
��ѧ&pa�g�B�<�!	[�f�ج9P ��t�H��{�<1hD/QfT�V�E��L�(b�Ly�<鰏�s��"��p���%�[yB�|���'B~�ȓ�T�}H"�1��@ǈD�	ϟ��	�;��ئ�F2��0��o�tB�	*��"�Ĝ���C�A��>ղC�	�*D��4"Q{H�)���MrVB�	�=�T��˖V��$x�/|~B�2r��:�*BhŒ��G!��3�pB�ɽ8tn8��ć�,yh�95����B�+d;��� �>�pҡ˼flB��#������
i'6Ӏd�--|B���
��MΪ궭��ID�C�!��T�2��vN�%JDF߻mr�C�IW����qӘA�A�rk�2VB�	4���0�
�#u|��)�qc��=я��?��ƥP��u�7�(E+`l��7D�<��͗t�� ��=#4���2D�låQ.	��,q�CY�0�Ę�0D��C����0�'͘(�*�k�%<D�D��ċ0u$����֢NT�x�%M:D�TJGȂ�{��*P ��cۼ����+D���A'U.<���f�5[��j�,)D�<j�ˎnyf3cCoj����&D��P���6%��dPtoR�m�� �*1D�� ��9p_!&�:��㒘Ȑ\c'�|�)�ӵ�~d��kԣ"��򱂉�@ٞC�I�e�`�Z��u<ȋ6��;�!�$ُ���S#@[�P	Is��%�!�E�+�h����ưA��hX�������<1�ɘO���g	R�w�xDY3j
�l�`�'^(xT���+�X�g�F�̑�'g��b풶=�yqg�� ����'q\���B1[p����@H�qv���
�'5��k��>����N&eB����'��=H���J���F,37��S�'��%0��f��- 4�Cg8�����O��0h�Ő���e�	�"���t7x�QA̬��#q�Q�}S�C�I������L樠[��t�
C�I1oI��ca�� �1"���,6��B��D!�����]C��z�K q��B�	�`� �z2�1Uˊy�Vݤ)��C�	�C���-�<4(�1\>!3f�$&�S�O��	������@s��=��p�"O.P�CĭU[T��� ׮�̉#`"O$���ĒH���r�O?��)�V"O��9���o׾)�.B+.
:<��"Oҽ
ƪ��_X&��("��iS"Oޘ��J7uWl9��� |�$��"Odd{�B
w~��`��H�qdd��IH�O�%���M:f^t��-�hI�(@�'sj�1��b��+'X�S\��@�'{��[uu�j9���\Z���j�'r�|�V��s�x)Vg�V:!	�'�*PƯ\-$&��RK��X	�'��j�L�
/����r��8IF���'n����ԡI�4�#bΖ�0D4��' F�I$E�v%D�@�ܯ/.X���'�Rc� ����;�f��_��y�șXsx���+��=�8�z�)��y�h<`��j K�	hBLA��+O��y�b�oA�3� ڗt����Ɯ�y⡝�]*�	Qb�݋z>�d[&�yr��K�pe�⋬p�R434G
�y2.E�/�����![�e�2���,��yR!ök��{��Vv`9ڲeǅ�y�,N�P���B�-Lq��xe�L�y��I�J�d�a�X�`x��e��y2��q�����)�
ZIx����y��Hj�P
�O~@X �G��y",�+WRP&lE�EI��?��?�'A\����2�Hl�`j�hͺ@�'4��'''���Q�.��cDveQ�':Tp��hI$�V�"`_�Vz)1
�'� k2�0���� 9����	�'7�質��zU0D�$��%�4Y;	�'+ٳdi�xR\(S�o�G�he��'�j;ӯS.j���3�<��T1�'\���IB'Q� ��$,R�x��'��5��Y�i�a�1���@��7D�dhw�W$	Fhp�g�
|� ��i5D���l]�p�	���� ��T�P�%D�88��c�^�&Ǒ��SG�&D�P�c�0VZ��V�`���R2&D�(�֌�����F)�O�z���$D��;1&�Tj||�V�#JZ)�s�#D���a�@PC�4/N)K%'<D�\I��P�"
D��4�J�#XT}��);D�� ��+4�$ny"13��O�$��"Otⅅ.bz�����@�z)85"OZD�m�H� �Z��]*Uh�`�T"OF0�sK�w�@�փǨGf�8 "ON(c���~Q.�Q���X��re"Oz�D�e5�A8qo��~�nȣ�"O�=`�斎��x�HC>(��;�"Or����4Pp�0��в��Eq�"O���#9�̺�k�~�5��"O^-��-6װ��Q�m���"O��'�_�	�D���]0eb�"OT��I3kL����ُ>ޭ���'�^�)�'L����F�,}��-AT�����J
�'L�H2�	�3��J��Y�v��	�'����D�I��yYֆ]�=uxY��'* �̰K���ߚ/�|-��')~p����h���=�(���'�09�3?�P�j����.T�+�'
��Ir�P�sVH�1'�-��'�]J�攮�$��0 	*$�*�'��P�%F-r`7�"���"O�s���D
���:VaX���"O��r�U�A��n]|����
�'w��
�F��B��+eH�6�l��'|�5g;`���R7%C&ŸY��'Ղ@�% �;)�}�V
\�^���'�(l�&@�Q�0�-C��XMI
�'�����
E�8�zM�I�f4�;
�'��e� �78�Qk�@����`	�'��`b�9b�$�(b+R�*�(ms�'��m��D+/�ʴ{V�3R7q�
�'H�	���ц v¨���^)Q��#�'�ۀ�=/m����*���"OL1ڶ�͂sxd�䗥|t2�aG"O~�����}�7)ѝbI��AC"OX�a��7;��Ƃ��"�Vab�"O�4ǩ��W�X�8ga�r$�}B"O�!��HR:ߴ��@.�&Z �<��"O��DC�J2 Y��bS���J�"O�횔$�8�D:$��@�u+"O>�C�a�V�69r�hڛO�d�!c"O�9��lK'<� ;�&�%uj)��"O0E��o��>��MAdf�_�h��S"O�<E.�%�b���Bêz�&��q"O��B��Z��H��
�_Ypp E"O�J�C��q�q�~V,]���q>5�� �8 ������.ڠ@q�L!D�P�u�Ĉs4T}�v��
7�h0���!D��8�+R5p�X�����2(��B;D�<ӥn��"��媗�kdq 4J5D��(F�Ʒ$�	"¦��1�:Q�6�.D��ኡ+.�5F�!h�&}������6��2�R�Q�ʖ)X.XE{��'h?E�CEׁY/0�`so�WDI"�2D��`�̃	Є�$�M!a�q��9D��� ��"��Ts�
�*�ᓁ�8D�D;U(�
�2�,P`�P���,5D��C�E�1F�����;WYh�k�j D����H�?
<}��iXJ�s)D�`3�/A��Вn���� `'D�8�T�ʤ!��Մ6������7D��Ar$X�,0J%��V�H�Z��#D��jE�L�t��
SF�F�(�"D��+T!�o�B�3�Չ$)�����?D�� �AK!''bt����
��S"O^�Reꐖ��"��ץJ�Nh�T"O\lR���K`|�j���Q�K�[�4D{��iޖx���l��Ӳl��S!�d�I��C�INS�4���9:�!���q��%�nB�4Z0P��V1g�!���zڀxૈ,q�)x��Jw!��N$yb�'�`��ݥ,M!�]9>�<���`�hʬ3#�9qK!�$̂|���@4��
~xaRt���!�$�8��F��
f����F�>O�!�ǕI�z%8�oZ�	�@�Hu#!�!��	 U�!L/x��� C#Y�!�]�"��t9Bݎ3y��F�.�!�$ј.
��S$l�4�Б���&�!��8)�$��e�4_��9�K�4&!�D/?�ȱ ��T{of:zE��"O"}1	.p �"h�=5p�`"O`���M z�r�Q/:MJ�"O�)B!X%��a����;? |ae"O�0�l^�X��͓B )}��XV"O2���k�����~b��[�"O�<;�5�2pa7 ��7R~��"OҜ��M�O��92���$މyT"O���(.3�S6�cs\��a"O&l�%Ș�|c��sg��8s�(��"Ob 8�L"!<�Z��s>=`"Oށ�B�C�b#��;�?>nV��"O2(#TK�6I��RGB�k<=��"O��U��0G��Hɰj�r�pYx�"O�U"S��9��.�bL���c�'�2��@3TNʻ��EZ�F�mlP��9D��;T�#pW&|��� p�����n9D��
��L��4"��.�К�1D��ceV����� +�r�SG0D�������,�Ӥ��3�`\j+D���D�=ah*ґN%INd��'D�� b
RZ!Գ3Y�.�>d��$D����� �R|t�+�nO ����5D�x��G@YH}jA��T��؃O2D�D�b�^��<9���)fWĈ�J5D�`k���,�B̀ѢP0?g�=�q(D���QT�t����0��!|��)�Eh%D��(��U�Z�۷�M0u��J�>D�X�$n�J8 jV8�x���(D������� TpFB�c�(rG(D��nª+V� �TGd�0���w�<A,{�ʜ��ct�����L�<�s��8��A���"��PmG�<Q!+NDJ�8W�-����hBi�<iw�s�.qqd�@�h��#��@�<�a�(J��1�7N�s"��RFF�H�<�c�^�� 8�t�W������D	N�<)S��0g$]����&�j c
L�<�%�2aP�����A+Б�%�F�<!5$ {��A��Ϧ.�!XĤ�B�<g�Ś7ct��f)֟bh8@��r�<aO� Z����E�f��c'�h�<�5�жf���¦���2��P��<��+��s�8y҆"HHb6��lz�	���?�~��]�e��&�L�2 �.D�4! DN��@�&n�1�B,D��Z!�Z�
,*�[.Y�:M�,D�PPB�Y�B+
e���)st��r��=D�� Ľ���
��XY1Έ4�l�pw"O��{��� �x�E`,F� A�&"O4��J�!NDIy��ъ_���X�"O:E f��0����"� T��R"OtP���1rE�5�E�a��y��"O>=��͎4Z�xү��	w�H�"O(Y��7n�z�Ba阊0Yz���"ONXK�!��PJ�G�N�2u��"OZU��N��^H�!'ZW���z7"O����k�y)�E��P�l{$"O^,;�ș)��������< "O����/S��Ha���A�P��ݲ"O�@k��e����_&�H�W"O�hS0 �wG\���G� ,��"O����Hǲ(�4��f��"��!�"O4k!�	k$��ĀW���#�"O������3e�±����3�~ *�"OF
�@ V�P)�$F��ҴRp"O����	ů�>𑣗�d>��B"OyX�@E�C!� 8�Ac7m\��y�-V6�����$Yl�O`�C�I�^`v�p�	�2+���Jůxx�C�I�C;����NV�#�Р{Ѩ�1*֡�D�8e�a�)�*f�Ź��0��'�ў�>uZ�喊Ȥ��C�^m��"�3D�XY�I�`3����J�VY���Qj3D�4�k�Lg�h�d�?}�4�+��>D���o��8 ����)�,�aC(D�pU�%J.P4�c��;���4c:D��q���Z��SA�G�8���P��*D�	���9R� 9Bƅ�[�5���<D�p�b
�\����F.Z�A�O=D�t��eX����*)L�4��$l&D��ئm�0q���%�̴�"�#D�����_�y8�'*�-s�&7D�������pd�.�fu�c��6D���g�@u����/T��q��2ړ�0|�H�g���HUiB�;\�M����X�<�p�N�H.�t�Q"�f�>���eZ�<)1��X85���VY�ꍋ�OWV�<��-'-���b��O��`�
�y�<�4h�~��E1@�V�n�иVH�x�<��K��g�P�FG�=� Aց�u�<��Bj��(!Q��P|�#��l���hO�'r�m�ѡܴ�joP��D��=�l��b��;� ��C��)�@�ȓ6�x����
*|�llٶ@'�2���~H�T�E
�D�*�` �Ī8��̇�W#`�`i��ep����"6��ȓ7�>T�%�غwE��ѰK�k��ȓE>IcІ�:�h���"^�H��Յ�Ie�'�� �%K�z3�Z�o];d:81�'m��P	#8M6�p�Z&_�d��'n�[0���8�4� R���
�'��MB��O!i(��
���H+O��D�W�d��m͢]C��ɥ.�!�� �}ZQ��0��IѦ?j!��[�'^\��v
�e��i���N!�$����e��8�t��Bd3�!�Q+����d��t����W�Z�!��6:�H�iuhC����:�U�2�!�d�K�F ��� .���]$DK!���kB�hs �����x���f!���u�� �{��i
�O!�� 6<����.ޖ���/��n���B"OuIF@%"���zS�5��"O*p�C��v`�`�A�θi'"Ou�q�O?:�&��$�H��(�Y$"O$q��ZR�촐6
��z((b�"O^ � `(۶�H�W3=EbT��"O�	
U�HX6H��0i�E��"O sr���ʲ�b$ՒO(H�9�"O"�q�����4��u�Ľ|#�JB"O��GD !���Y�hN20"ʼ�"O\a�C�O/N���NA�3'Bl"O�9�%ۮ ��9���ND)!"OƐ!bą)L�@�ju�̓;#R��"O ����E �
�aw��~4��"OT5�B'�3%��ᷥE����"O¥�­�5Ɓ1Ö(wV�=	w"OF�!e��r2�#���0VD�r�"O�h[��r�m�4��%nTj�"O�r����,�(c!���6f� �R"O�
C� z/�T�J\aDY"O��@�U�k���0JI�&�(��"O�<�� ���h��	^`�t�p�"O-9��K 8(@=a�(�G�8��"O���SF�1@O�q���<:��"O��(��@�r����$#�5!"Oz����
[|��a5c�'�F(r"O���/	�c(ֈ�SK�;#����"O8�;S�Γ;�^��T�>T����e"O���5���K@�\�˅&4����`"OV�aԺ$͖�kb��;[�����"O�}z���W�:%0C��2�^��4"OfY��۬~,fQ�X� ����"O� T�Dy��i�N�4��"O`��(G7�v���`�<���B"Odɠ�Z�F9��JTa����2"O�`:'@ڕw��%���A�K�:��"O~�"�΅�	#�z��ּ-}�0��"O챋���z(8�V-/�F�f"O����,ۻ1]��్�i��p"Or]܊P�8ҁ�S�TO���"O�bю��L?Ɖ6	E|���"OB�:������2>�I��"O�ܳ���W0�!�41+4X�"O�I�`�f��
Cޚ{x�4h�"O���ժ�)U0�ɲ"�خAP��q�"O�Ds�jB�fL�u�.�1:�$ht"OR��� �\��m��L�CCv��"O�	���^��yi��h��4	�"O(!A��e�H��v��_��p�"On���z=rh͛��z3"O,���W�h}7bA���$Ч"O�8@ ,|lB �*�^�J�"O��m��QF�z��طz}�XQT"O<�v�&`��0Cƕ�b�="O���!�<$8�eR�DZ�v4��"OL�
��"�̅��$�� ��`(""O�lfM�.U�r��Ӄ�#Et��;�"O<I��*کU������eh��b�"O���Ϗ?4MBA5^~�x�"O���*E/#���iЯϥ!o̍[�"O��3��8Ej�r4�7
x4%�!"O`XiG���u�	�X�cQ��t"Or�����$�.@8X7��A�"O�P۠/�@Lx(s5+��	GF�R�"O� :�3q�T2c�X�GL�=R�֌�S"O��l�3w��zV
]�k3�4��"O���FW�I��ke'S��z�� "OFP3�OJ���ҵ&����i�"O؉'�P�]Р�����r�"O�� Ԋ[8@`jTJ������"O����U$���A 	��\�z�"Ot1rJ�*1�����G@�1�6���"O�p %�^�N�C��j�`�o4D������u�v�sA��h���kA+#D��;�]A��v�ĮN_Bu���Oh���OT�D�<�|J�O� q&D�S�\3��:?��("OAQ�8�d���Q:D�z��c"Oą�1fJ�nPQ��(7t4]�"O�����I%k�����\$t<�T"O�qB��'	�P:��K%vr��rB"O�]�󨏮H��<��l)\Q���B"OBY��i�( q����P�Cd�sq�D2LO��#���;f��#���P��G"OrlAwȍ�[���)R%J$:���"O��p#�a��(X֍�ݰ�c�"O@��#R	�f\���-���pW"Obx�f'�2r5��Rv��F�^���"O��fl:}|�`ѳ��R"O>ń����掋$ ���e*O��2l	_l�w�M�2���
�'���G��;��	Z���$Y�q��'��R��ɦw���Y��[�#ZT��'�r\���ɉ8�<���/�;c�<�k�'��{��8/J��Ջ��\ڜ�Q�'c��H�]2q���X�dόSiX��'><C5_�erd��L�B�#�'�ҩC�#��P�*4nW�	�	�'v����/
_xĸd!ޅc�Ը�'0t�ԯZ&r��@�'ɴ'��
�'��0��!�z�#4��&IxB	�'IV�P��<���5�H��ǢRK�<���ǏSn���ջ<Hxh��	p�<��O��g�@��O�0d"��3�̏kh<���ۘ. ��a�ZX�u`&���y�R�N������XByAam��y"(T��Ί�7�Ε"���y����ca����dE*EIؐCC��y��"Pݞ�q�S;#J괺���y��h8����D�)7��0���y� W51H�Aa/'պ8:3'ۈ��'`ў�'�X�Zf�D5o��=2M9o�,��';�p��[�5��XY�J�>j��H�'��XÑ�6KE�԰�O��b�*,��'�8wa�&/�N����"{�&C��.���o�0�6����^��C��B�0H��E	lG�pfG��jfZC�I�դ�����r���!&ER�1��C�1IY��S�j�8�|t c �)!M�C�	�^�lC���y�V�H���#C�h���#���)&d���C�	)_��%�C�.WNP8��4>�B�	�`c>�� �S�Y�&�x�jƃ$�&B�I��R���/�D͘�+C�%J.C�	>e�<����A�%�fUJ5�L 9ʼC䉫N\��(�T���0�(ɴ M�C�	^�*4���XKpaӢ�G6NB�3�T2�"S�t:���˃l�>B�ɬ%
���1=�%a*�6r�pC�)� �!�π$�r��l�6����"ON��R�<X�m"�M�EN�!а"O�PxGR�^�$��TL�dh�L3Q"OL���ß:-�"����ӕw�0��"O�S���*�.��G*�7����"OF�ˡ�άHS��1D�:,�!�d��x�XA ��)�� ��)�����hh{�n��S�B�
R��>C䉠D޲Dɥ�N"f�ʕ�`�A%��B�:��1��$�Q�Ԕ���Q"��B�	94�-�Ư��l�Pc�nO�mvB�	�o82�w��>��d����0`�B�	6H}Q2C/�#t���g�
K�bC�I8���B#	QfސX��J�1�<C��!6'��fO�@O���� �u�dC��_u�,I0��\˶D��È	c� C�ɎLeP�ڶ@���w���z��B�I�T0�惁~��,1�"�
T��C�I4$a�oLF<R���K�|C䉳<��=���"��Hz�Ŏ�czB䉦0���jf�F5G;n�R��
u�C䉱g��P�O�*E8!�S�٪E�C�	�[�����J��"f�g�(B�I:���SضB�� ��LR.
B�	�m�2��_�
UQ�T��j�B�	2n�v�˲�s���BOî=G�B�,K����p`��C�x�hC�IA�NTAg�&;7(AI/�-g_6C�ɝ��g�Is�$������B�!���RE��es�$ZFd_�e�B�ɒzcĘ��k#p�A�E�[�ܣ?i��)�0@��@څ.�Q߀`�Ь�%=!�$�<C�8UZT�P�g�"<��kƣ0,!��~�4J�#�67�x<�K�>!�[�dz�3�o�) ���Y�ʝc!��� T@jc�ޖL'D�x���9�!��b+��ʗ(�2$>�؃%
ϸ1�!�� 7΁��'�|s��T%n�!��Բ�D3��P�}��'(Ćh�!�D�=��cգTb0$�!��.�!��=x<a�����r/��C& �+?�!�$ҋa*��
�ڲ~(�R� �(�!�ĕ�5�fd
���-v�9�O؅~�!򤁵����0���r`��i]�1�!�S�	�5�B�{�����"�.�!�d�X��d[� &�"�*�A�4�!�dV:����gO�5~{��C���r�!�d��=��D+6
�d=��.�<*!�$�HcČ(N�����G�4M!�҃�P���	Dӄ��v�:$Y!�$���Pȃ5̾M��yɲ杕k�!�D]����s�1]a{dh F!�Z#MҘ��	�R[>y�A�
�E!�ą2V�E�F�@6���+��02!�D4� �� č'��� �7c�!�4%+�8�Ce��G]�ha.-4�!򄐚:�֍���hS0�AA�5�!�d�11�m`d��R.a#c�K�S�!򤋇B|�@api��W4H��i_��!��َ`NU��,�Q�$D���j4!�T�Wr� *k�)	`^<3�Ǆ')�!���[Щ3�ʖf5������!�=:֡pDh�	]�zI CX��!�Y���;ģ�m���q����~�!�� n�b�b��S(	��
�tK0���"ON!Y"hň"�N��nϛ{8\a@�"Oi
��A�6r��U�Ȍs�=�Q"Ot<`Џ_�O�n�Ж)Ƹ05"OD]����)�P�q�t���"O$q�̌�@�`�"�'8
�>�`�"O���&J�.��yPdD���<��"O��I�3U��,(G�2�xAt"O��9�Hs�0����)�"O��ࡨN{[|5�"��n�}!�"ORCs的��ja��=6L��"O"�c@�j�]x!-I3#ɰh�"O�	r��(��p�,�+`�Z���"O�Y����\��,s�,|�r��"O��`S, CDQ+W!l�x��"OZ5ZgA�D��h��Í)����"O2x �M,�ڌ@'�* ~�"�"ON�"� �0c �CA�>_��=��"O�PC�\wv ĉv!�;�^�9V*Or-��ܹ?�R|�QH<v�F3�'����#!.M�PK��q���	�'wf|���M�J5\-�%N	�neL���'�`�r��fe�Ha�LҸd1d��'͊��	�=KRU!�TY\D�(�'�Ё��ㄥh?��Cu�V�gljQ�'�@��gܖ
>(���YX��a�
�'K�p�F��x����b]�Sd�L�	�'�B�J��G��T�b�Ç�:��
�'���Rj�8)|�K�恅�b��'d]�w$��b'��*bq��'��A�B�1�4���� %��(�'U�]R�B��P���!A�aJ�'�\1����;�2�6��Q��'�`�C���>>�p`�� ҏ1�t��'�:�k`W. �X�!�t�z���'	0p�D��xް�r�/�7S�m��'X�����J�Ld�R��4���3�'�tH`LH�c��4ƂZ@0��0�'���.ҽooF�����)A�h]r�'�>ٱƎ�U
��@�D;�u��';r���e�
�X�JD��{n99�'��Ȣ$�<Xn�{sƇ�u>�)��'�X豕�Ej�`��*M1m.Ē�'آ�{Cf_�G��9���R�JIA�'B>�R�c@:C�����o�3����',�(�2h[�6����B_�'X$12�'���i&,�'p����!�2#Vrt�'� ��#_ΎXi�̃��Y��'Q|�#�#/9��6B��P1��'�6��@	9��xZ`�Z�sO&��'�J��μo?����ą[ML���'�f��$�,]���E#"Ƭ;�'� �XS
1;ʽ7�>6�-��'z�qɃ@9�q(�j ?/8����'���#�ǀ{�!�d�/.o�)P
�'1�D�bZ�ƶhq"�7�*
�'j���#��Q�f�2q�A:�0My	�'��Kt�L/@Ɋ f��
��HX	�'�t�ŁMO�Z�;�k�	'J��	�')\|Ӈ ݕl�t���*�:6|	�'1`���G� 4l���}���	�'3Z�c ��;S4����O?rM�}��'k�l����m�\p	TW�b�'L��3�%2&�WI��!<����� ���&��F{��ٕ#�o)Fa�S"OЩ!��V����J?5n���"O�@��B�K��Ɂ�,ޖm0���"O��Ж#J�}4d����VlK9q'"O��p�:u����%OSRP�`�$"O:L�&��4%޴�J%�.V��B$"OE�����@`� ���r��S"O�P�ڰ&���0'o�4{�"O6E:�NXkh�Ѩ��&G���Z�"O$\`5�5u����K@��R�"OD<����5-�D����$�R"O�laO��s�N0�b�D
A��`""O��5�=>|�<[�T2w:�01"O��c��[����K:M� � �"O�p�PNx0Nlx��[N�2!�S"OD�8"9
�2x:�+D�PAp"O(��NÍ'�9ɕ�K���٫u"O�H��/ϥ�f�JV���S��mP�"O<00�l�&E؆���7/�����"O�@8��Ԓ�i� ��:D�^�9G"O�
�Ň�,��r�GܤBP(,�!���^��\�z�M�� ��u[!�D�HD���Ə]�Hp��̅$N!���3
�j�z@��MZD���ɠN!�[$�>���(Dd�y�h��e/!�Đ&ka�	±ڼTrcƉ]+$!�*����DZ�'Nxx����u�!��D�j�9��V�%�E��h��ob!�dY�qc *�ݐN�[f�74Z!� <Zx���I�=��в&7'@!�K��`y� ��\�r�6E(]�!�N�s�� �fF�Pvؕ����M{!���a�li��BU.Pn��7�ݢo!�0
}ά�EE�+;}�4�Dݑ9]!�V�.���矵*u��qsa��>!�$�;1���Õb��H`�akS��%V$!��31n��Ǒ;<��-h�.!�AKmrH�v�H9�P�N��!�D�, ��������B���¢�3�!�$H�_��p��KC�:.�[ �Y�V�!���)���`T��F~�J�� -j�!��̜0�vtS&��:Y��t�6���4�!��j����J�7F중�*?q!�, A�s#�W�2���ի9b!��%??a�2aø��a��п�!�$��aP1h�5.�$ ��ӫi�!�HUh�1��D�B���c��%A5!���� Ђ��H�
����T��7!�dR���&�Q�p+.t�s*�~�!��l�[�kQ�*v��B��k�!��]�ډQ�C��Z������$�!�	�4�ذ륢��oK�)�͊�ys!�D_�S�ع���K>U;<�4k��8;!���`b��$$���#H�3< !�$�
A�$l�iV� �ک���n-!�g�B�i��Na@a�Z�!�B�
�ht�͆{Z\pC3�ۑ!!�� �Ĭ��E�><\!�Op�!��o�.ML�.O1�R M�!��3��Dq����FG0Y�5vG!���$G�Ic`%^�%4�X�Ν�F!�$Ѿ5�L�&c�;i/�`kף�$>!�dR*-����q�,*l�K��ٟ	!�D�!`�����(�m@�Z�AÙd�!�� 0֣D�h���OVX���a"O���c�b�D�HgiZ8�n�x�"O
�BM�0D�ى�*E88�؄��"OyJ��P2|k�P뒈D/t�z�	�"O^�x�GH�|(���M�O�vd1"O���v��$��#��Ț0�V�`�"O����R4�>�1��ƛ#�V8zG"Oܨ�s+ܨ�4�� HQ}��	�"O
3 O��8I���(�f���""Oz9�w�	g3x��c(�`|\�`#"O"��8-����HhΘxr"O���.��
�3!�n[���s"O�$���0��4��
�:4:�m""O����,H(Pp�P)X�G,��"O��0� �D��)���#d+�=���i�ў"~n��W��bԇnc�����4��C�,KU��H��š#2����딺n����p?��Lqj)�g%� RP�R�gW8�x$��zU߂)����_;\��)�$D�LЅ�̧e
h�� �����i-ʓ�hO�S�.F�@"ڨz�l�K��F�B��t���E�"BD$��H�{��B��8*@]A#3>@^؀���,WB�	�
���X�*��Q X�ّ�A�p��B�IE���Ғ�"f�l�����? �#?Y��	]�.�p��g%�]R� ��)�!�dB�9���R塎� ���r�@'k��A<�<�%�
u�|�9gh˞B���P�c����'��[qD��2I�2��R͆����M���M���<���'N���JI�'a�&�u!�0���~�I�I�L#wFX ľ!(`�$v����e�����B����c�*;y��+�dz��G{��ɝ:kȪPF@X`Ey�Ϛ<���
O�E��O�Z�$lq��҅wK<ŊRT����	�cn�А�,2���Pg���hB��|S������LXaaźQ�RB�	<o4�;�Ձ9��$3�$:Hh؅ȓ9�L��ą�z���q�
PQ"����>h����M4d4�� ��-�E~�S�?nī�)K�Ș���y��B�ɸJ�F��fO6+�d0��.Z[p���'g�?����^W���5LC/J,�!*5D��ۗ��8<*�������P��q�|F{��i�W(�ȄfM4S��e�F�q�~�Y�hPX9:Jm�f��N��0[fbC��y�%P�l�`Q��JՄD� �J��y"��#L�|�4�\)<��y��
��y���?h�컃d�'CPJ�"@0���p>��gH"jJ��2I�7�|�	��O�<�Cf�2�����U�ZY[V��r��0=AKZO��ʦ�R"uրH��΂k�x���Oc���l�(m��D�$��;:�Π�0��HD{��I%H��A�źga����,\�@!�$
�i�`P��0��E^'S�'F�����0�4)ńǻU�F\�6�ь$��	���|<Q�^3�ؙ�k׶uI,�9���;��9F��o��#|zp�2�PQ2
Ŝ �i���`�<� F�>n0L@�O&��Z`�<16D8rb<i0c��b#��R�%]S�<ɔ$ӘU�tI2C��"v���RFLh�<�"+6lxP�'�W 7%^qJ�MKo�<��G [���LK��P$�C�<�F��"�*p����`}:(r�lKy�<��Ùt�-�aA�@��
2�hO?�)� ���+Yf?d��q(��Ra��X`"Op���W wg�}���]�z�6p��':4���e�Mdm�ƭ�8,78����0D��"�I�A�x���X�`��B�2�I�<Y	ǓP3��V������	�Z���z�pb����^�F�9�@|R�3^��#>��i�/����lR ;N� p	��gQ!��������fT�Sȟ�w�	x���'��d�$E��A�圿R�n%X�fM�T���<IOIZ���O���B@��%����⊍.⊅��[�� �W�O�t|)c�8]�)Ex�O0ꓺyBS"|�����Is�]�A$���'ўb>��%M�0 ��$����|�TDP�jE[h<��J"Bx��î@i�d@�K]�<-P1AU!��Ԏ5���Ӈ-�@$�ȓ1����Fiͨ Ӳ(0�̛Q~Մȓ(O$�A���?4�I����	R�ȓHDd�Q
Y" X��8vO�����ȓ#���	4a��+a�H�j�����ē���S�A&�e�#۬���b��-U�B�I�X� m����o�צ��!��'�a}��@�.1֥!�E��),�AB%葂�ybnHLT�m���X_ڸ��oW7�y��
, D]9���.L��9�c�����7}"�>%>�?t(�EO�m0X�A@�T�lq�O|��dV�6SD���<d�Ҝ�b&�'�~�\���寂��]�<@h�.�1�L���d�!I������N��	��l��'�a|"�ED`0����>����ID�hO:����Df>��ɃC�Rܸt˗.I�|h"%3D�PK�ˋ�gq�õd>l|�6,��HF{��IՄ&mRhwk��y���Ŋ;)�!�d�=��L����a眅��%��dω'�ax����J��J
��9q�LEZ�H �c9D�t�$"����#Jx��t�8D��1��P%��6CH?:��5S�D+D�\��U5]��y2��3Fҍ�fN+D�����؜&�̀�O�"+���&E/D�Y�c��f�D�Bs)Z�˦�t�,D��в����R2�W=h`tl+D�|	 �I-����`�{v2x�T�%�O���z�D*`ʞ=`E*'�C��4B��/@&�̙�m՘2Zq�d�>"?y��;�hKE��ژꢄ4D�����	�h��5��gȫ2m�U�K����C�	7��{#N^8{���P��D�z C�Ii��y��6)t�k^�RB���E
Te^m*
�K�B/e"��Ɠ�R�h��؍>�� ��K*J��E{�O^2���@�dd�}� �J��	��'����T�.�(U�G��2.�T��hO?A��åe�lxd��2z2(��N�_�<!�޹\�tI��lG��Х�T�<�d�Y,B���� /� �I�j�<1rM���Y�F��l�9��)�#�!��׈D���ݮ!z��f�^�6[!�d^'E���Ǡ�ks,��$��Y�!�<�\#���/tnN�qC  )����~oU�S�O�*�+��;1o`,qL�"��U��'e�١7����@�A0��8s�n1D��6�V
PJ��H�ꛭ8�╋D�0�D+�IN�'�j�8��8%��)�n(����
��y�X"Ib`!QҊ�hj$�ž�y��[.�����/��$r#��)�0=!�
� �I��Ar�P�G�VHG6%�"���Px�
2�F�q'�k�2<r �ߝ���~2�|R�@Zܓ�*e�b��m�v���mȬy�ȓDE`�0fݛ=r�l��D�X�|0�ȓF2�R�+�S(h�EÙyO"�ȓ��!�T<Bo T��㘠$��ȓH�������'$�I��i��1�ȓMR�P��a�>�Kn\,p}��<������O����s�w�}�5`�� *�ɰ�'�x���M'K�����KZ�A�<Y�AU�06�8S�ظV�a:r�C�~���O	�$@�èg#�`�f
�QF����'K���&ѯ2f����S�N�T�	�'�֐���	:!��3�`��Bhz|H�'��@A�Z.Ę���f�-4٨t"�'0|I+��C�/HtAH�͚Z8���'#�� K��9�Ĩ��nԘ"����'
�Z���6iyC��;&�:���'v��̣�h������M/8P��'-5����R��;�π�7�����'+M��ϋD �`�)��|��	�'�F���'ʝu�<1D��C`�Q8�'-\A ���4M�|X��'ʀrz����''���dm�7c�%��-���!�'rV���
?s�@V��}i����'~�%ʍ��a�r*��e�<}J�'q\9��Q��(�����K�9z
�'aV}�	�;��A������	�'�$�Y��ݸG��@@f��~�Ur�'ê(�wO(���V���}c�� D���*ұX�]�u�X11G%0b�9D��P�aF�x�<�"���b{6\���5D��� F(j��IAq%� D(�"d� D��R�ܶ]�h(
G�b���=D������ʉZ�M	�C.��Pq�%D��	%̖ @Rq�%	Rz�)qV�7D�$�d�k�`���ˈX��M+�A7D����kQO�%)n��0[T�7� D��)�ȗ(�<�I��T-m���`��>D���æ����,UO��t{!
 D�8y��}���*�C��dk�C8D��pfJU5� hуS5N`�SfH!D��ʀ�YVL�B�Q# �Z��`!D�d�R�
&�L0:��P�~A��<D�𐁮�7C>���s���q� �E(D���숬R=
�@䎒�1ٔ�S��;D�\��C�$�tt�goσ,�%�G=D�+��$\V������.,ۀ*:D�l�ц̒~Z�X�$�/Ee��F$b��W%,�O����I�q�ҹ(t J*k���"Ot�s
��r�0ebe��:3TD %"O��" V��9Y���:Q $���"O��#��В4��jKݏy�Xs"O*�+�dQ�,��F��`x��2�"O���UQ)�$��ˀ�Rp�؃a"O�����\%J�b�Slڥh��a�s"O�D��Fa�h)vLQ��P1F"O�()��ǌ �<�r"Ce��#�"O��c��`�b��#lh�T�%"O� hN��8�`�%��qTH�"OVy���²G�EїE�1R�L� "O.��2iD�Q\��Dd\+�|3T"O�ԣV+�)ʎ�JW���v��x�T"Ox�+��Z���`HC@�� ��"O� v�2(	��I�s���-���"F"ODXsu�މi@���ψ�j���У"O�њ� H�g���ȃ`S3EX8&"Oz!��*��)�^�YQ��~tz�"O��{@!ξhn|A J������"O�2��/c�P}�A%G�z�B7"O|�� �S����'d�-<�(+�"Oȍ���8R^QpAC�M��Ș�"O�\i%)�.e"��SD�)`�:E��"O��KƩ־@*V�rd��).�Z�A7"O�dXB�I:�V�ڇ��h���+P"OF�9@oԤH*X"�+ȖZ0�+�"Ot�Qߝ��B��j��hD"O� ɥ�ʝK�	b�Dڵ�\r�"O��I%G��G7�\�$��6>�LT e"Oꀰc���6"8�c�����"O�ɋ��:JT���\%���"OFȢQdP��!�/�,Q��Q"O4ˇd_(s	H���*���p"O�-����+?�(�2�ֺRټ���"O�q���$cJ5؀΀z��"O�����a�Z41@)�OI�`�S"O�ĳ�h��h�E&�C�j��"Ot�K��T;<q���
f��4A�H8e\��I�Fh�!�b��a d��� �S��􄇱5|�L�����C@,Y괏R
4Z��-D��B��P�@����aoՎ;+h���)�	8!@�����R<�v!����`Ɉd��1��]�ȹ���8D�HCtDݎjBh�g�ј=1�97IX�GCqO�뤬�#!�qO�aj�w���kC�ז?BD�c�b����'w*01�ʕ|�j��R+Kb�M:@'B�S�F�؏{"�H�P�Bb?���>j���E�&�:�2�	��az���pp�O�thw��P��#���?_��*��O@��l߰�0>�a��5w�ҀED�]���X�iC�G�j���h�P�x<̓7����DM/fC�ap�o�b�2@�ȓ[���5o�	;�@z�g�"q���DyBI\X�k�S
��{v��>I��B�!~�B��LLLB�gN�D��H�Y�L�6�C�K���"~n��?3tH:T$�p������54�B�I��<q��;S���O�-�DC�I73�ʱ[��X."f��3��˜L�B�@�d���ɔ>��Xk�ZP��C�ɋ^�*�3�D#,�r�k�?�C�ɨ��H	���yt��!�B\�C���9���<N���,KfC�	���1�s�
-��$�l����>��'����I�($��0��g:RDQ�'%:�aFE�7��:��� �0�{RB��T��SU�>\�`���ufܐ1C!^�	�ZB�I46ā�äɠ��۷N_9y�h3� <�I�tQ>�;����%T�?�P����L�_R�5��8�&�[V�r H�%�&�V���<b� y��ɾ@����˞2Q�,쩇�ݾA���$�5p��c�O��!�Ï�4p�����2l�v4Y�"O50�gX|�R���/F>(B�)�&�d_�"ݚL��'\8�MN8U�X�c����ȓ|���E��K�`D��e����G�+�	��H����yZHI���I�T�`��@5b�B�I*k�0B�V6Q�RAB�l�)��B�	�7�� �
�vȱq�M2!3�B䉷6��hŌ؊L��a�"�ț�F�tD�͉x�ax�b�
�4��&��t,!�F����x�"˞h�eM�4.Z���DT�g�^�p2 ?[�����Q�����	*y?�trDD�%��OD�[��%���K|� �d �OA�.vRu1��/bւغ�"O�Xh`�&K$p��-� �"�B�U�$���R�i~��>�|�G�Z�:E�e��!Sn���e�[�p2�SY��R	�$�Z�!��,\�P�r0W����[B��3�ҕ��)�h]�Xw�[Ag�E�zqk�Ok���(|�@a��A�RbR�J
a|��xSX����K�6aa7E�J`XD��lO3/��X!�钔uV��䦄�O���bM,?�����Oޮ4�t
��O�`|!A$Ծ5R��Ě�E�AY�I�t�f�2��+O�i{�wW~�idh��7������¿kG���e'?w	�zݚpy5���}�ŋj�fx
�@�'N�~hB昿4T���*��Ch]�䫆$Wi���@Ŋk�d|�`6��f�	޺9hw���A`ԡ�� 0Apa`�Z s6t��	#UL �3AW�.Z�lK��vED2�-:h��2%M7g�b5X7�d�9��+�^���ə?�����?��V)�L�԰� (�(�(���F��A�� =	�4�@%B��򨠥M�5���I��<_2H���]� HI���7Lv����OL��v���N@괕'f��k5�7+���%��03�X%(�B�۪	Ը���̅jZ�9��S<gj��b `̹���ˆ��X������!cZ@�gJ�n�����'F
	�2��?�0<QCJ&یuA�\�}�ш�B�3��1�ٶ�����ڌ"�Q1��%܂i#!,\�	~��ؼ�V�Q$fٲ�ol�ؘpka�<	E��w�d�����H��L�HB�SS`�Y��|��ď�6K�4��S�v�h��g`�J��|����<qB�/!轐sÜ��	7�A4�0>�tF	9+	�R"�-p�R]ہ���H8d�뀬�-iH�y�OԴ]�̠��?
�>��6`�u�BEG|Ó0p��2�o�h��$pիݯ�(O���"��p��
���3j��(X�K�-,:*%[�E�=JJ�E��	R�T �T6���$�K��}�/	�u�ZYs���T�Ă����zX9�ĩ�*I��n\(mmX����u�:��O� �"�B_�LMX-BP(�	(^\���'�d��$�D��0�d�-(JL$�S*��LLR���0B2���$ģ:�1�$ђ���"�y'#L}��ŀ&�I��$�@Ϛ��y��:�jP8��.R>L�1`F#}O0ѹ��A�|�J�%�p��O�ўlX�e̍K��Ђ�X�D �wE>�O���w�	�.�.��B�4X��9Cj��f�|$+D��1�0%ڝ1������q�t�Ӥ�Ҷ^\8c�ҵZ��X�K$N��bg�
�h��00��e�t��^U���,�&^��Q�>�yb���_
��S�nUcf�m
�L�'j�.��Š��A�@�i��$C��q�v�s���e�M+��܁�"K�]
�b54D�� �	O+�,��/E�0�7��
r��T�r���YFη��L�xDT�3ړ"+���3�R(:��+�m�fJ���DU|���Ɉoh�Jtt�N�X�.�~'rl@V��Gr�LQw�'����l�G�a�`��8�� �M�NcF&O��Ԡc�k&�$�u���+��l7$�
s#�y�m
@�Q#�������J�MbcH�"o���㒼;��Xa��s�b�)�dʨ4��,� @����D"O��9HQ88O�qc&,�6�́9ǯ	[?q�۳`u�!�%n9���	�{NY��.E�_�(DI�� 9��$��@w�- �ߧ �Z%�"IB�
R8E9Ҭ�43��u
�', q�v�W�$�,M�AO0�Ђ���!_0�໌��!Ջ~ 
Dxc�5s>dPPaaѶ�yR�S,A��\�seO+u��drDO�&�y���"%�ٻ�.��OB�PI�!�y2	D��eJ�B��)�9!pDT��y�<aJx]���(f��x� ��<�yrHG:L����E!��C�P�y��U�}cƘ��c��$}�й�	H*�yR���7J��i,���a��h�y*#�Ll������GƘ�yR���K������ӽ�����.[��y�*��, ����6��ͩ��8�yr(��q\j��a�X�{g�`�e@��y�=~(-��	E(��I	� ��yrfWn"����{g�Q �(��yrg��y��c�'}���B!��yrf$%ǰ���&��Y�<���ѯ�y��*��b�T�c>����y�'_�4�#Iȫ.�8Up2��+�y��2\=D	���I�u���l��y��1[�%ʄhK�!Ĕӡ�ݧ�y
� �mɠm,Un����c1d�<X�G"O�}��P.����D�6��U"ON�rL4�����G;�ᱰ�'��3&F̓� I�Q��P5 S�i$|���" D��Dĕ(+�\�gѝT�^���C??��#9�x�xM>E��"���G/��:$�Su�5�yb�7=�F���,�%m;�I��e�����'�rh��if��ϸ'#:��E%��bon��D��<�����i'6��E�H�^��h�7�Q%�%��#P6}�t�uL/�O�t��+�hT"ɰGH�l b���	3�lr���&��Ok<d��&�:�G޻`���$8D��YW�W�l�!C�Z�$g�<A�Ew8R�3}��	�d�*��L�.��)�ㅻhu!��O�\�H�mW�&��VX��OTY"R��.����qO*�vm�:���B �l�#�' "���Mb<���G��.Dㅃ�0T 0�0@F�H؟x+����ȢG�3x�@��  ��`~lR���c�����ڕ�Z�R�`���L�&���;g"OB��s	È��%R�� )��������[䢛�P>%%�"|���@�;���h�&`5���f�Q�<�E��IG�Q9�K��'{�
4��Q�=y�r�(Or(s`�0餽(��= t� C"O�8b�>WʘId�=w>Yj�"OX�BJ�<c���seX�i5"OF�:wU ���W��c�ND�<��`��:l	�Q��xL����E�<a�B:e����!U�;ƕ��KC�<)�K�)g��) ��ۣ9J�ԋ�[y�<�,T�30�m	��[�ؼ��ƪ�w�<y��:R��1(�NK�g�2H�գZo�<�"�	x��!�儭bk�E�g+�|�<9%(�>�HAz��\� o`y���z�<��E�U���Bc j��Z���L�<A@X)TU� ��`��a8��Hu�<�5$�����D?�8�vO��<�d.Q
>v��90?{��@9 Ep�<y'a�(^.�ze�Tծ�
s��l�<�B�Мk֬��(��G?��
�E�A�<)熍8�
xB�M>s��  ��B�<��.��)ha�^�(��(�GC�<I"��D v��'b&�q��P�<!�m�4N�\��r�(D�p�b���v�<����9Q�>ݢTK'<��<8��p�<�2(�,�()��+M!E��,!�JY�<�'��T��'�ŻuD2�{�ŋo�<��	�*�� ��S�C�ʜ��C�<9E
ܽo<4qK��<zQ3� �`�<	�얫C�
%a��.x7�	3�k]e�<!��T�5��4ȴ�/a��
�J�<9��_Q�� �W<�N�z�HX@�<�#�>j��b	��Y� �1av�<A�	�h���%��p��B�Br�<)�dNƸ;�����M�6��W�<� 
�D��-��mV�~�:&��e�<��ǖ�A,�X kȖc��ԙ��^�<�@!�3Q��q#����BYfZ�Lm�<�f@�+�6�s��i4@H��"Qn�<���%UB*�PD�)D⨛���h�<)ʕDzP���N+so�|�R��k�<��@�,W��K&�V>�8��D
`�<��	���D�Ⱦ\p�����`�<�d$X9v�L��9p��ѹcnT_�<!�`��"��=�P'��r,S�Y�<�$)�;W�LX�E[<-��2!��a�<� ��R��ۖh�h�N؏Y�\�"OR	(�@�,>	p}�$QS�����"O�40��W�Y������l���Y�"O�HuC�m5*�#�&�&T��`[d"O��Je��!�t��@W)<T��V"O�2!a�p��3/�<?R,ѵ"O�<� �
e�1���M�Nx�@[%"O�x�I��X�>E���D�H�5� "O��6O�.��-����r��٪�"O��ͬ=��̀Ɓ��Y�%	D"O2hJ4Z�H[rH!A�C�~,�'"O�h�����c	V���"��r����T"ODmY�-��{vaA2J;��"O`�i�H��^�����#�}k�"O���UQ`|y+���@��`�"O, �$�)3L%���[O� \zV"O&d��@�AA�1i�UB� �"O<E�%Ooϸ�(��5� �� "O�����Ξu%&�2�lŹr"O��(��c�0�jD#_z��|�$"O����!(�n�Ҧ��O�Π�t*O������
6j�B�)ג+�zI��'yh��%�$}oRd���:/�`8��'��0��#>Rl!`g��1%bx�b�'@�0�a�-c�
T���ݫ�'g�ܓ�(�%=P<�ʣ��� �dA1�'�� ��H-T���K�-_�~Ď@��'��yA�M�0i �W:m���'�4��h�-����n�F	�'#���U����U+\6��*	�'���(��m)�P����3!�.���'/lx��k@.m喅[��W�EРy	�'�|I�7�̜Ź���<�FmS�'\�(�s(�.��؃!��kx�2�'$|���'X�|��h���qK����'� � Ax��R�$U�o��-��'h|�qp!^�R�&�ScaK,�^���'AډЅC��f�Yf��"����'(����K���p�x'ݣRԢ�B�'G�����=D�Z��h�;A$���'Ⱦ���,.9�h�DcQ�H�����'P��/F*M'�$��ϠD�^@��'�r���&?�	�Eޫ6F>L��'���Q��~�ͳeCͽ5�E��'��N�9膄J�c!����'֜iA*QOI�y��,�(W�P�
�'�������\plY����( ��	 	�'��$j��Ӯ����$�
K�@Lk	�'�h6��	'�d�sB��E9� �"O��\�o�t��#U�1!�A�"ODe���@�c��m���
+��кw"O�P��-��l��H���Q�u��2"O��à��?C-LeP��ƞ�24�D"O,Y�p����T�E#:T�f�w"O�u�F/]P�UmK41T-#�"O֥RE2jv|HPk�;���"O� DǏ�V��#�Qq�"O�]�%"K��0���#t�R�"OTYٵMJt(��F�X�&!�&"O���w�% �C�c�#9��!p"O<p���EI�xHD�8��xa�"Op5A�Þ
�f���`�,u�i�1"Ot��`D�\��ŋ'�9yJh�"O���T�YU��(�*W�6��h�f"O� .���7vDlx���)�bMS�$	�N�"�!�Y@*}�5�]F���ԋB�#_�=���YB"i���f=���F��8��Q�t��\=via�ے���ςH 0zi��8G.J>
<1��	d�S�xBz��Dd�+ "�,B �N�C��C�1*�,��n�f��	
�ɯlA�˓8�Q��h�'��ӧ�O�A��FN4�B\��N��a��<��Ԥ-��HC k$�O�-C�F(9� {��ӓ|RJ�٠$\2EBhԐ�#���4!��%ŘM�NQ�3����LźOJ�i���&N k;��	��V-)޶5�`$�OhA��٦!�L��G�/-����)��e���,}(����0?\�*�Jޤ����'}��)����<A0�ÒBϴA�1-HG%�O�a�HĬ.~�X�@�&=��q�"���H�Ӛgd�,1&)M�*�$���`��"�Y�O
U2�@> 0i$>c�L�B��&^(X1��Q�w����7"ޕ*��@�B�pD�*'ʛ,z)�m��*�zY����&Zt����䯘10C|Lc6��|e�	�i(�O�AX�ː�k�����B��s��c�I�Ə�;�$��8t7�.Y.B���sB�O*��2^ �@��%�k�0�aT�޻��x*�Gp�{m%�`���yl6��q	J0V��6Ǘq�q�g�B����(��lq�'7:]�!�i�X��x���Z�r��W�e��O�����=�"=�Q��j��%L-?�d瓘@�)AE����l�3�$K5H+rc��+�D�5J(v��$@;ex�Y�cI׻N���H���X�
�&g�=�~��tHۋaL<���*�:gz�N�>sp}�t��2�x
7Hَ1QRC�ɽY�|u�`	�	r9vY�C�k�2ţ�	W&�|����(��F��~}� �'fP�yA@M���R<[<~���Ɉw���.G|*�!��,`s#��/ItXD���)��X� NB�5� ��l��(����t&��1@��gz��Ey�ɚm��8�C@ w*�� �f{��v�(���׳G7T�i7�C�2K@B�I~$��+��qMV\	5o� "�����B�^���S�O���{���<�Ȁe(D9}6\E��'�~�����s��0eƕ�C5N�	�{�
V�%� ��	u �� ЇB
;3J��l�ZC�ɹUؠ�S��@��.�J2�_�C��C�"R��i�"j[�/;\�9a(Z��B�ɼ@Yl$(c.�<B>pɡhZ�J ,B�ɧff^e#�fsPq��V2kl����odvU�80����_/n΢��ȓtC�R6��1�.rc�˭F�%��/�T`	4F��8�2ġ�j[�{��T�ȓ���[��6&V�� ��"n�ȓD��⒂J2hb�CV��;�,��ȓVw��+��Z	D�f�V�n L�ȓB�f@�6�Ƙ@"ѪS�F$�ȓ	��	r���0J5�Y��ƈ<ФU�ȓA.P�a
�h�6���A
X��@-�੄��&"tp���Ð�"gX`�ȓk��Q�e#T O�
��a#�1^��Q��Yo\�!"%ĠB�ԜI������ȓ:�8�R�9Q�-ȑY/\�N��ȓ,�� `0�aBL�H�~nv\�ȓ� ��`l� ZY���G�=J��X�ȓ�(�[t�\CL@(�$�Yè�ȓC�1�*�4"Щ؆dE;gT���+����� �ox\����;?3����$Ϡ��'��.n~ő��ڛ�C�	�g?<I�w��[�.���n�* �\B䉧W�R?�UYq h��L��(GVC�	�hg���BG'C(` GN�m�C�ɒNѶ�˵�܈O� �pL�[ tC��B�Xa���)*���C2�B�	�\�RU�v�ُGG��Ұ)�C9lB�ɣh`���2G��F�n� \Z�OK�<Qc�%�j���t�h*RF�K�<Q��5Dd֘�0� U����D�<��I��
q	��Z���L) �t�<�u�W_NMx��i��x�D~�<� ��ƅĔn��Igω�g:���"O�=[��G���
��� �:q"O����CLek�`פmD��5"On����@�3��5T��"O>����R�xځnֿe�j +�"Oԃe̕�<R:|z��ҬO9Z�"O��j��tœ�3H�����'���5`̓O `�A�K�=�~�Y�!	��}�ȓ�t5���/O���Q�I1>
��'�r���1c}ɧ�L@B��;E>\�� 9�E��"Oz(c��#��A�����1���r�DŻ��[��*���ߑk�F�k��Ԉ"iDK
�#D�bD_�o�D�z�C��E��[�B
�C��ɇE�;L���ɆP��m�G��d�8��S�Њp�أ?��	�;��ڰn/�A�i��	Z��I5,�j����J�|}!�D��Ƚ�M��.�Zat�ƇXj�I�l�E-�S�Oi� �ի�W%��HbO��*|����'��c�l#�L�ʤ�*(�|kt	.}���Q\������{�$Y*1��iP�a�7)�@�K�����?��Y(4bܩ�$8s��������b
��aǟ)K���D�*#_�pBnD�;f�:w��.g�џx�w�8F�8����m�Q�N����I�j�d�p�̝�y�E��.aڐ�o�.nKTM�1��3��D__ٜ��C,��Lㆥ��k*J�b��#:�XC�I�Ql�Y��pI$�e/�`�qO����F�0�0<���.d�:Xz��A�k�*�K&S�<�ɘB��鰃�H�vIt��I�<ٴd��2���ԕz9���(�E�<y�+�#������ ��%���F�<4lL�mg �c��K!i�6����A�<�(T3B@�CK�6W�	���P�<q�
�XQ��R.�$z��^{�<��c2RNXe�T.�#�����w�<���u&(Zd�H�u��	y$HF�<���0vP�X'-�P|���MG�<���Fw�,��GiB�|�&\���<qFω�#�5 �Żb�f��ȋ�<Y�n��-������,8��a�z�<��BZG��`��O��:�ӧ%�r�<�%����t�b�UH�XT�0hl�<�F��@-ȱ)CF�BhЌh�A�k�<�P� �t��2H*zo����h�}�<���?���H���%��
�<�di?cj� I�#uR^}�֪�z�<�$l��0`��jp�w��HY�Ev�<A��ܚ���be�¿���2` f�<ie"��|z�0[�́M��$��ěd�<�pR�����"R
}xD!��g�<��B�ݙ���_��)i���K�<iT,�i�&h�f�$9K�t� NF�<��nt�X,!�k�B�(lsG �K�<�p��bln��W��=���	�K�<����:]Hy˕P;F���ȃL�<��C9j��A�4��u�Π��&�K�<q�OF�Q��@/u� آ�A�<q�l[�+A�h@�.��YҠ��U�<�u��*K3~���E&m��!E�[]H�����_���{�e�.�2bh��
��h���&D� ��`�GVxh��ǀi���k��$S~���?%?ɉ�/^�rx蘛�c@.ð;��#}"ɇ \�O�d��$��8b� cq�%I�\�s��O�]S'8�)ڧ$���S e�T�%*<��H�I�5��O�?�����_98S�&��/���A��?�����>�`ɟ�Sg�O�`񣂦F�"gR��Ǐ5.���/V��򄗟?W��π � wF�e��h1t���`kXP_��z*OP@��@�O��a*B�SiՄA�2�U�V���"E�WPj�S����CR�	�Mҩȥ�T>v*�]u��<A�זS���<��'o�,)������
$`�E>O�͚"Y?�0Q�"~��j����i�h�閅��	�O�4-3��O&l�����<�'i����5�^%��л�!F?* "-��\��Yb]�T	Ia>7�>�' ���Tn�*B��c���?f@���I�N��I�>/�5�����$u,�5L���c�v�XYS��<Ѷ�ϱ����|����lԱfI�i��.3y1�	CW�Ch��͓?�P4�'l�y���OY����8�:�P�� 0V��������d^y
ç%�8i�@�T2���Ҕ���x��0�'h��x��4E��'��!j⪏9;~�]�u�+�`$0�'�剕!Q�b>q��@�f�J�1B��}%� ��,?1s�(�S�O��qqi.����@Ɠ�r�����dUDx��I��#/�`)�d,K�� ��8%���O�'t�q���ԟ�t��,oXÂ�a�fгw��/3V�������,Y�6���z���u�O�r�)%W(X|@H!�ϗ�nx��ɭO@��bJ�~�q�s��"}��� +h
(,��}�R��Bɉr�<Y0��,:�ֵX$�V)s|H3�CCd�<)��d="͑�i�pRH�;6�G[�<���?=�\H!�`B7()�e��QW�<Qb��QN�ӂ!�Ύ)��	�U�<9�� ođ��M!E���HN�<�� Y�!	B�Z�i\I6$A�$F�<�#$�N�ʤA���9���x2 @�<AQ�F�EC.��c�Ųw�fX2iCs�<1�
�,����%D�ؓ���c�<9��"aR�ȩ�h�+�\��V�b�<��O��w5�6��R�^T��bTZ�<��G�$@Fy�f�:Ӥhq�AT�<�-Q�q��Y�g@/@�ئ�v�<�7m���O�Ez�ʢ��q�<�t�@��8�/�  ݾ���C�<9�H�&.�V�T3���RHNW�<Y4��>�hC�З.v���g�k�<�V'Wnz銲@ݐ9�^����@k�<)q����,�p��,-\��0�o�<q䪙� �R��2i]�{�ޱ�E�C�I��qP���Y7�	Y �^Q��B�IJ�R,A�Ԁ~B����,/PC�1M�,�jc�U�OD�e@�d/l�LC�ɶ0(�� `�8,֘B��!]*:C�	;oZ����¡y>�db�m�74C�e6�Y	��tR��!#m�I0C��Ql��ִk��)�N��� C䉽sD���˝E���
�%�5�C��!*�L��Xo.�E�$;�Љ��'� m1�
�>E�Px�eȑa�xŪ�'��d�2-O�C���B���	
�>�Q�'L����˨|VN��L�	�Jd�	�'�=Kj�o�X4�C�	���e�	�'G�� #�>Ci�#fEM_8�Z�'¼�����D�A��Ǐ�0��'7h}���9�]�U�X�w�yI�'�D��-�H��e�U�><vl��'B�ᧉL�cQH�ceL�$� K	�'+X�Ul 'Y��_)t���!
�'�v4�����`��0А��	�'��嫷c�D"��d�]�
i	�'����EB`Y���"���'�lTirHns<Z3DL �hE��'��4���;ҕ����f$رY�'
��Ua���+�fZ�X�zA�'��-Q5�g������]�^1���� �	Srl�u�n{���d�!0�"Ol *��ӯoL�{qM���&�	�"O�Pb���ٹGm�01�j��V"O��f�QW�up�����l�@�"O^=��%!$X�� �M��؁�P"O�E@��7r��PI��,8�N���"O�1`�kZ�X�d�CV�&G����"On��ˏ8�2��dèy[��@�"O�M`��Q�paTC�CRXc�"Ob�P��ҌO��aEC=|ybQ"O�`��u���x"cˬnoN囗"O�<�����
Gz��-��@*
�'���0��U6J<�FRܥ��'���pABC�? �L�[�x��'½K�B�)6�8�2���"����'[P��e۽H�z�z'+�/?��9�'�X�GK�xZ���Cn��	��q:�'�L��.��"(���Ʌ$|9�'��L@�mI�Y�ʨ��@�0�T��'�kU��E�.�r��v<Y�'����A�4|�dy��C$HR�'����	*��X�^5.~ZI�'�Xx��PvN��Bq�qz�b�'�J��dJ�c�nm�gf��;�(�
�'ަ� 5�U�#V �6�Y'-��\�
�'F6q�Dݦ1�J5��a�{h�
�'b6�J'<M�@��"D3oҤ���'�x�C��LI�GW)9҉��'�F���ͫTͺA	�ɟ'"$&l��'2Pz&$��JR����N�XT��'����AU�@�j�����EԐ��'�T�ҁ��EFL��&ϊ/�"O�i � ��gl�q�A� �G����"O�ab&n�Rr��ۃ.�DR����"O�}Y�ݵk,B-_OT�	!"O�� m�-]G�	��L<Q���r"O���&H�&fV̸�-�,iVm��"OFP��lN���2�6(�L�`C"O:�c�A��C�f��1���=�#"O�Q�D��>%�V�霛X��%��"O� �d]*IĠ�@��_�: "O�D�v@Oz׼��h
�?��͸�"O�mA)��#+���2��y
�"O�qh�"�I�M�ࡕ�~�vl`�"Ov�0�Ί�L#�Ḱ���Z�d ��"O�݀Ƥ��ABp9''�"��sS"O��Y�U�y����F�9
�h���"O����=/�� �g��,M���1"OB��vMT�m�b����6^��؛2"O��S̳�J͑S/�a�Z���"OHx�ʊX'9��KEJ
� ��"O�u�@D%x�����*�5
�-ڣ"Ov�96G2�@�2D���|L�"O�y�1ǅx
]�w͉�3�4�a�"O(��"Ç� }R nł�
�C"O�X���+�X B̅/PQР"O��5��9li:u�e�\�	��S�"OTٹ�N�((OFL:F%�/����p"O�P�@;R�19���/֎!�"O*�XXz��6c��i&C2!�DH�Jwx��AC�i!$@�/!��03T$�t�H�(%�#Eޢ]!��}vfQ��!ЊS�2���D,{�!�$�'ʶ-֏� ,����'%�W=!�� .�y��� v|�,єCRD���"O�tx� T���s��C\�Z�"O�����~)�-!�#�YZri��"O�-�ӥ M�¼� �5
f�y�"Oҙ;#/Y�A�A0��T^\J�"Ol��gXY�QƝ%v=4���"Ov4x�/\�vi���М~��W"O�]��iӅO�f�h�*��e�Z"O��@�fޤGC�$3BI\�e�\�"d"O���G�<�6�⥪T�5�%�""O��Q+���,���)ʄ�
�"O�QZ5C��O��R"c�v�"O�=
4�3B��@ -1��X�"O�=#@���3.V�� �3 �e�&"O���%�Õr^@ ŏ	!l��E"Ob1bS��"�����΅Z���yr"O ���D����͓�y��T"O�}��V��
<�DK���"O0	��J�~X���g]��)s�"O���IJ�X�B	���L��,��"O�0���ͦ$ɸ���I��H2b"O�# ���+�dq� �y~��3a"O�:�K]T(�c�{�8Х"O4t¥�ϗ+�zx�lmv4�"O�!�����D�EY��A lU�A��"OV����/ T�rU��<�]�6"O���Gd׼W%��H�h
9�e�b"O��q֊�-�`����#d8�q26"OX����ԥJ�"��'D�(y�"O�봄E%��0v�̙*Zt��	�'x�ᡦ�1b��.Ҹr�l+�'ڦ�pЌ�W��j�KD�qF<�x�'�&�Zd�J�R�,�����n�D���'C�E����;������s�0�'�Ɣ�
S/�(�$G�eV|1��'sL\���FT���Gf���
�'�Y�wNX�7KLpP�I�0q����'����#�8E���6B��*�!c�'�x]��ၨS_&�1�n�X���'y08��R����նeѾ���'YFDhኆ.T��#�ݣ_�ٙ�'��q�WŞ�#2��!���6\´�B�'+�QA�Ǟ&N�5Z!i�M�J���'>X��LUN�D`*��>J_v��'�����%�a\	;!��=Q൱�'�hP��H�:�����@��(��0�'̑�ǥ�Y�ŁE!��Mpr���'Xz�S�B�.p���b�/֝��'��HBc.�.��e��S���y�'�F��r��&���;�FBH��A�'$6���G'�����ʅ�r�~���'h��[�"IȸB�c�t�:�'����'ʙ�P�Nh1¶Y��)9�'�*��c+��������%�y��T�\\�Y�C`�����;�#���y"ܚC� �r�U"f�(k79�y�Ozaejs-\�I�)�(Պ�y�`��P�R���pS���y©Z�qy����s��Mʦ+���y��= ��8�,W�l��p��Z�yR*Z�/�$�f��..�Y����y���)�<P-��*�i�&w��C��.���I4�ߘi>���m��^�C�	�Q��\��,_;]��)�g�M�K��C�)� 2A�G̦HHp'f[�(�"O�qC!J�=
.�A�,Г`W���v"O��.`�z1IR�D"���Y�"Or�h�cWH�ꎛt�1�"O�a���B'@K�ISDhW��zi�t"O�c�`��9�SfZ=o� R�"O"`Q�T9���Qt��=�k""O�`#DeP����R���u�(K�"O��Y	��W @up1�=,p9�"O^ɂ�I\�Y>ҹP���W�}��"O|���cZ����Qp�U 0C8��"Ol�	5f�%fO�xR���hY`��"O�\�.R�;,��ؒE-�ypv"Oā聧^�b�9�2�R�8��"O"���.�y޺ #��vjj��"O��.1S �@*���.C}s2"OR�%�
	n�zV�gT�i�"OBD�a&�/���Z6dEy\���"O�Q�`��{��AӰÌ"nq�e��"O��p�Mի>z��B��PbH!�q"O\h�Ю|��5�F�� �q"O����XPD��M�K2tK@"O��P   �P   �
  '  �  ?!  .)  &2  i8  �>  E  CK  �Q  �W  ^  ad  �j  �p  (w  m}  ބ   `� u�	����Zv)C�'ll\�0"Ez+�D��8��M�P��<iW+	ٟH�hǺ��o� -���
6��x���;d�N�M��P�H�V��	Aa��]>b������Ӑ2J�mJ�A�Qd�jC�I����F `�}y! <vhX[�Z4Q�x��_wX�R��OvR�ľs��+�� g[���֦ԶA,��aL
��䁷�$��3-N�8�lZ�~1H��ǟL�	���ɒ��I�5G��]�6A�-�]=���I�H�ݴ-?Hؒ)O:�D�[�����O��dӗ�>H`u��5&�(j���5x����O����OF��?сbք�Mkt�'���H�����Ձ!�BI�� �I�HF|2�i�D5�b��*Eܩ���y���0aç>i��Ĥ��CBKB$e��S�3\��a<%S����~�l�D�O���ON���O����O�˧�y���^�<�� X�5�앰���?i�i^46mO�ٚش�?᣿i�PFw�@-#f��O��'�_�);�Yb��I�|FU#G�M�'�j蛎��n�÷�s�j�17� /�M`�,X�|[�q9�H؉s\�0�BFz�
<o� �M��'��blT����Q�C�(���Ū�2<��93"��h�����*t
�hQ��g.��r�#N3H�J''��e��6͚�A�۴~�p4p5d�R�4�$�K��j���'Z�P�!rC���y�to��BZV�	/N[����, ��d��)}�%�g/�a*H�z3]�	��`_*?�B�	�4l��(b���ء/a �P��
芸{^w�!%i
�������dD+��i�^x����y֧�h�L���'�Oxň��߱-@�s��080�s�o�O�����ǟ� ah�0�McʟzAŦ��F~Q���T�1> �2�'}�	������|�	ߙi��Ժ�O���͖�b��fn�tW��kf�)@����D�.K�=���/a&��4��O"�yv�ϧ���BR�T=
��H!�'x:����?	�T�@�<4j ��[�E,L��g�OH���O��b>�ϓi�5�To�$>X��#�K�f�����Mk6%�&��y��ȑK)��*> U���ė*C����B;��+gJY4H$b�*�C�'�F@�ȓ-��"�)��?�zPj`g�m����(ܬ�Ru�Ũ֤�@�ݔ:5
l��v� ���c	Mϐ�auO�A�����b� ,���^���:S��B:�ȓ'$���ș� B&Pr[7�p�I6qb"<E�d�&���,G#Q�Yɒ�^�!�D�3JJ��h�c�$-x��^��!�d�kV`�٩w&�P���$.7!���6�ʭ��%N.%~p�@�Ջ!�0HZY9�.C��ZD��(q���6u!�Ȁ&F�'d�Lp�c���#3��c�<9���?q.O��'��$�z��б�0!kX�x`�� ,��w� �K��}�y�xI� IU�`h�C�ޡ>�T��%��7���
w@\� �8��0k�n�ўD��cH<Q�j ��*c�Y��A�X���æ�+��ľ<��O�@u��oyr�*Q-��|�0щ��'�!�dҦp�dL�敉x�B@j���T�BFg���	ͦ��4��I�74���lZܟ(ϓH�xC��:��t�B�N���cy�'Tb>�f�RV�+1����C��)�G�ԁB����}�iE
G�"~ax���'T�0m�C��fV�I��P�ra����N��8{�%9@��KG`�à����UFyB�X%�?Ig�iՒ6-�O8��g
�0����]�bM&i��E�<������(�@b�ė�e0�L"!v�AD�	p�'?~6�-g��qF�i&��$��� �8�n�c��}3�s�D@���
`��% �����^t`�`b[
�yR� 4or���X9X�^q#ӎ�0�yRB����R���d��ɫ1h���y�%��?�� `��F�&<���.�y�͉�q�����8�bP:��yR� �o�M��G<���JQ)pݛ��| ��%��$�'w��'��7)��5�`�M\0��C��SΒ�.�k�ĵ���O�ej`��2o��'�O*t!�#� h=|x�N�6S��*�F
6\򙉥E��w�64SU��?V1�v�Z&g�f}�G6]��q ���va�3���?A�T��˅��O�b>���O��Dι,vr5��gρWn�JcH�Ӏ��d@�q������Utl����	�!z�'�h7���U'��S�?��'t^��`f��FE���mޗ>'���j4
g�7M�O����Ox˓��'VHH�	��N�g�F�r�B3 ��<�8rEEE*mk�=+�E�Y�����Y ��%�P�ƷVR�{���4e�t( �S*(Ъ�"&�	=E���{e���HO҄�'�ȏZ�[b�B�K!�E�6-��'Z��p� ��?���?����?�ΟP��c�5jq�.�t�x`P�"Or��M�=�hY9�K]c�`���|�`Ӹ���<F�!�f�'�S�y'��* 4�37M�D���'�؝��'��:��i��'>1O� ,�@�1L�N<C��Y���ZW�'�R�s��d��p�Š�.�97��zhax��-�?!W�|�%J ���z.�*NL8���y�DB:'��7��8�޵���Xj�R��OD����:W�8�
��ո��დ|�-Q94���?1-�Ȭ�ć�O@�x�ˇ�1�X��Ȅ'8}�$d�O���B!�X�@G�t&���O(ʧ��ɋ1~(�URÇ
"����d���mW�!*2��X-%鉣~j2�xG%:��~zL�AG�:����49�O0\t�'[��k�H�1§RN@[7A�.�$��[Z�}'� ��A����'��yQd�;.D}�"nS0&����զyjٴ��Œh�eM�zf䄂�˅�N�F�iP��'�e�<(�� ��'��'K"=�xx���&��X�%���1�Q���	�U?��I�~XS�[��Dѩj�b�A�U=^yL���&U�u����(:�;��֊W��6�*?iR�����S�'UH-�2�Ŭ �E	e��Ij\�CS�p���+�OT�@��pbA32!S�D��`s_�tp�O���6���ğ�O��4J���c�ԕ��P.�t��#�0#;:6��O����ORʓ��~>)Y�"�6&��a#`eH �T�ؚid(�b�i+8��Af*LO�H7ꕻz��l��KLJ���I��d�R��u�,*�8=��Ï�i���e��(O�%���Gs���nƃL����it҉z�X�lZğ`�'����"hoN�T�?�(�P)��TD{J?!PE*�y+J5&^C�2��4�WGC��n�Jy�O�7��������3�+��]�Zp�`ZƠ]�4����uyR�'�2:��
�"��~�	(	1�r��}���&		$��	(���4�ax�ݽ'&��Y�h:Zq��g�I'S1���.�����gW�7��q�eB�w8�]Ey�cߕ�?�ķi-�7��O�5�u�˗g���a��:]"�(禰<�����(��� D���~�l�Ӕ`M�L\�E(T�I`�'~�7��!
�n[��ֽ!������&W��n�Ny�ҴKM4q�t�'��OI67�m��١�����\p)ݬ`����ӊ0?��_c����Q��b'$'���Ǭ�x8v�@����:�	5�S�OP�ib��?
���Z�)��KY~�M,�?!d�|���	�������`�J��Ä]�)!�چ=���)΍2Ȱt�`2�џD��	
�Qԉi@c�o��8�cԠKq�6#�D�!6���?�'/:dqEN5Q������$�=�y���0=�Fl�>?o� �� �M��F��C�2"���	�U�R��6.24_�sR�ÄVv�-$��SR!�O�c>c����B�<��� @�_>�$�v<D�ܢ�-P>cDɄ�<O��p7ʽ<���)�'��勔��#�v�)�$'�L�W�V��?q��?I����d�|B�O�	�q�0��Y�,TQ�ti�a� �r�z���I?.��4Ju$�/+GT��EͶ=u<�K�'�c3��A"�s,�zҮ�A�`�%��4z�c�N
(o�E2���?���xr�'��|R:�|trУǧv�);�CJ�!$�2"O½�a+�-~p5�$�� �(���|B�q��m�Vy҈��@@��'����=@V�ƪQ���!%.aRP�\�	ğ ̧An^����>	��
��tj�	>l�BeG��/�݈Óq
��B��1�ȡY���?1�fᑂ�6,1��X%��Å��0<a�a�ğX����M���z�8�D���[�j�ґ��x c+O~�D%�)�'L6�p�2�N�PS,�55���'�ўb>I��4 ��0(T��2����A\�P�Bq�i��	  Ū�b�4�?1,O�ʧ�?9D
���e���2��1�Ũ��?1�Ap�P	\e���ٟ�:3.�!�tE��jǭ^��	�RE����i��7��":(�	aWf�u�O���j@��W^,d�@��M��P��O�\�v�'tp7	�-��o�O�^� @@�!a^�SA䇫S�l�M>1���?���ԟ:�f� 'W��;� GB�H����I��M���i�'�^bc�t�J yw�SQ���`��'�>�� �4�Q���`j�RdB��ek�2~�25�Fi2D�4�p#Ţ��J�E*
$J/D����	U�w�.`B���O	� 궈2D��j�Gߧr=�hk)�A�j%�d`&D�TzU�ĘF��r1;#
1d'D�lbe� }��Ƃ\�p�x�'�<�w��t8���1&��w�Pu���2j%
�%D�� $A���U�%�C�A�5sN�jb"Oh%��_�&��H�� �ZB�s�"O�����W8�����
)\@N,�Q"O����C�7 ]�%���հ���'*NK�'9r�[&o�����Ĳ.���'K���#�Qϊ��P�ͪ+�N
�'�N�1�����2�K�'�<lN���'�FDjT�Êb� H��c\�H\E��'���Dʕ��l�'b��Q���	�'̢��^�:�����~�$#��dG�}LQ?��E(͌j,��06G�1�y��:D�`@ ��Bd,�]�Sצ�� 5D�<� *Ѝ=G$䲢��(�Dq �>D�8��C�"ѣ!�hA��3�"D����i��X�mRP#�b�"D����R�a�(D+Ԥ�������O�x���)�'J�8(y��k5�� r���0�����'�J���!O�3��@,�6(���'pj��숇2Hh婳��v�h��'0.�f^:?:`���n�zSv1��'�%;ǅ�a�b��a�y��]��'�YADj�`�)a��p�t��)O�}���'���ȴ�\| ��0�N��9S��J�'�v�3a�ղJ�p���>-�hqp�'�p)�&��2]��Cg�*�̃�'?��@ƋV�2��V�D9�ĵ��'=rQ;vo�\��V�J�7,b���HӜP�LAzY��A�(�Ƶ�lM#*<��jF �AV���K'
nh�ȓ"��9��bx@=Aa耟/����e�j����Ȅ+��x ��RB؅ȓ^�x!�4F��T8��pV��:ͅ��������9�e��s��YE{�j�Ǩ�<�S�
+"�rܒ�4��:�"O`�Z�ߕx�A�Ώ�^S̠�0"O�\Q�k��)zq#d�L�r��f"O^`�qF%jF$Jg͖�c����"OJA�Fk(n$<"����)�"O"噃	g�!p�U�B�v�'�n�����
;����@v�htQ�;I7$��ȓ)�= ���J<la����ą�8kB�Bĉ
\�V8�uO�;|՘@�ȓNؤ�#�M�wK䘺��6
�y�ȓJ��dZ5A��R�#�Sx�|$�8D�$�H���жD�%���i�ƣ<���m8��3�M1n6�B���x
qU�<D��P��C-��t�̡qD�\�p�&D�@&��^y�ajabJ;D�zr�7D�Z�3E���p�ڥw�>�(�)D�PSC��gg,��j�kb�Y��#�O�T�w�OL�K�F�HFl6��
��]��"O��ANEuWll��Ǘ�&�����"O���`����X�F�!RH�B"O�)�p �(?��S����ҩ��"O�a:q䏖;T=�	�5P<耰"OZⱋ� ,��Q�/mE�q��I8ix��~:۫:���VK��]�̝��Q_�<I��t��ʰ��F�Jܑ��\�<�CDɏ,]�d��,�a���B�<�Cc�:3���s&�.
���ONG�<�$
�"-@�n�]�^!� h�<QDg�4v���u� �g�$�F�K����0?�S�O�Uh�/�:�>٣FJ� ]�d�s"O�9b�_:?m~y�W�F�A��u��"O� j����=�� �������a �"O>�â��c	"��[8g�Fѐ7"OʑhwH  =AJ�MW�E�\�"O��� �1����6���W�j�`�Q���q�$�OrH�Bk�0��;�ұkn^�K "O�$*���.aĈ��.c("Ov��%FM�*)1�X�YS~��`"ON-�q�VKZnU��Y�&C��js"O�U ѹ;���xD��eF|�e�'����'T�0�RhB�(a'	�4 >����'�qr �P�4Qj9��.JR���'w�����@6�:H�6K*4��ʓb�P0��9d���"�I� 9�ȓo� 5: Ȁ��v���<(X1�ȓ�t�+1ǝC�8�sD��n�D{�M������h{���gl񈓬S�cU�1`�"O>������K�T�MϣI�&]�"O�ų�̣L�bD���+$-"���"OJ%`#-��u֠3e˔:Mv�җ"O����왏C	<E��M,[%^t��"O,("�C���0A�W�4�:Y ��'��aË���MHxx&�-���I���r�$@��p�z����^������(�<e�x�ȓ(9�b��y��Q�4���&����ȓr�T0KWꊖ[�]{Q	�qUȥ��I ��g��(�$�(�	X�dB����y����t��(>���������'�\����S��ޡ[ ��Bs!���]��s�\Y7+N~�"TΗ�0��ȓ�v�I�+A��*D�R��?_��8�ȓpy�1e��R��WM�:[@
q�ȓ69��;Ce5���'%��m��P��I
9
�	�M$2�����#�R\�Ê��B�ɧO+��V�ڣ��!3BBa��C��;\{l-۶
�#� }r�R�B�	n���C��k���ʲ욐9)B��	*KP��F�Z<Ja�a�hm�C��#h�4�0�d�b
�hk墖�a4��=��T�O5|�VΛ�Qڹ����[�2D"�' ����
�j ]�	M�|u��'��,;�NR%{�@��@I�{�n��'�ƠR����e>.�1�LUH��H��'����W07H��j4oӾ�65Z�'�Cw�m,,�FE�lAF$���H�Fx��	]�(��}xe(n"�5���Z�@�FC�ii	Ћ�<9�B�,g��"O
�2�cO�ָ*�$Hs��!S&"Oȡ(G�5\X�2$� H���P"Onk�M�7��9 ��.SߺZ$"O`|�DKM��-�� �0>t��cT�  @#)�O
��f+E&�:$�����3G4A+s"O�Q颯D�I(��%�?>V�"O4e@�ҧV$�� ,�(? �P��"O*�9M�4d�i4�w{��!9f"O� �a_�ؽBe��RQ�E�P�'��	�'�e�S��<���##(�3+�i��'5F� ���<K�=+B�5]���B�'��[��*&��)s���N��3�'JRh�s��}�F`��$�x0�t3�'HҜQ�"IT��b��:w%̹c�',�,aF��~�ԀQ�cF�z��찋�$�4I�Q?��e�?���i�쇁l{��Qp�,D�P���W�?����d%X��	%D��JQj�U�MY& �.w2�` *"D�� r@ �� Iwp�5$ͶT]�T�#"O*�
�@R#�	e��>oBh]S�"O������k�X���J���B�'&d�K���S�Uu��Cf̀�3R�<� 	#tx���'���Ƙzc�M*��P���ȓF_���@��fV�񡏜�z2 1�ȓ_��1��#_7��5�Qy��(�ȓ0����$�Q-0Qd!)�#	�5��&'��p%B5T�9@�Ҍhtf��'*��2�`�C�g�T�5����|w@�ȓk��]Ѝ�.n@���[�M��ǀei�iQ�v.����E\N���~���nXGhp�i�C�i�A��b��������"����Q�&�e���4Y�z�I|�T��P(N�L��gG×3�C�ɿt�Ђ�T,?{b�Q4B�];�C��	W��@bB��J��a+Go�0}|B��b�iB���q���&�5�C����8�������k%E�C�ɒ	�-C'�x�! �L��Rkx�=FK�}�O���J�H�*����ۅ
���c	�'���8���c�:�� .���F��'\�hC����~H)�`IWH@X�'j�HQ1M��5����F!�=O�L�1�'�vXDlo�a�f$��HS�Q��'H>iS�W6o�� ��ڕ LdK��j!��Dx��Ie�) �+��0D]b&)���*B�K���t�ˇSo�th�����ȓO��yȚ2P�fx�!�d/`��ȓ3�f���HD��p8A)B�p6|Y�ȓyy��K�I@,i��]�1K�9
�=�Ɠqp̌X�-�\�D��B��r�lx�����ɜ��$D�쒯O������ͳw�hxq;#J9=�*��B��O
�H���O����Ox��4�͕#9��:e�F"�zT���Z��uX��Lā ��i��$�"�I ��O"��ed�(��a�[�4.�h����C2�;�&���^�l��yGN�'O�����?y�����18�J� ��	��E�&����D$�ON@RL����"0 ��c͘,�ǝ|"�i>ɘ-O0�[�h�C�>]�֯�"!����X�<Ч�>�M���?�.�z���O��d�5^'���k������UA�#/d ���[�d����MS���A��-iF��'��O	�5�&�Px�8��k�'��؛'"N�Hv!��߆d���h�E�D��;AU��
k ���a8�y"e��X�IY~J~��OZ���#!�@��ϑ8�zm1"ON%����hY�=�GAS J�
�R7�D�O8aEz�OL0��g�_�u���r��V�LE�5�'���'.�b�G�9\b�'r�'�Nם���&(#~|��Pp��S߶0ړiȐX���tT$��g\�\D�g�'����0*��Ab栲�D��Ut(IHS̷>���ۯL��@�B���O%� ��� �/�d,z@h_1H���^2:���O�=I�'y��Bĥַ4�{4�H>R��'��݂��#)���S$��M�Q��7P����ԟД'�\��I��
v��	q��8@�	�(ˇ4K��I�'o���'�2nz�!�����ͧp:(�ũ��i������
�D�aŢ�
l@�Q�5)C�(�a{�腬^���pe�[/�.��ץť-L8�
рN�9@���a�>lO�IG�'&���NY>�Q"o߷Y�̨S��'�ўdG|���?XTH�c��ķFL%@0�N��yҧ�r�L��K�r(x!:7.�/��IѦ��	j��׆ܥ�vT`�큮�Tmb��<y��Ka"OtՋ0m�gH ��a��d�}g"O����^�9�i(��>jx06"O�e9�镑q�Z��I�_����"O¡����_�y� 
�;O�D�R"O��ꠄ�?�65 ���YMԌ2 �DV%.���Ok���`��_��І�D�ƞ�:�'�#v�A<8W��K�����'m�@����?+��UN�A^\){��� ��*�aO�i���ŊQe�(�"O<���_��t�q�<4,$�"O�A2.�!��-Z	T�؝�"���O��}��C���a"��mߢ�Qܸ6����ȓK�v{�
�
�\�(�n�3a��m�ȓ;���#�^'UH�)�E�U�*�����رT��ےv�%�<����$D�\qT�;l\4p���$�w�&D��5'�j�l��S+�29|ҵ��O4ZQ�'���� i� �=��&�:��'ɸL"@KͥI��!���X���'�2Urŭ[9�480"G��M���!�'v��Xq@��U��,A��7�@�'&�sD��"������2l�qk���H=1P�l�F��#P6@9XCM>�&58��pG���'���'Q�c��g|>ЃD��"q
	��?�O�Z���iu:��e׻<�`����y�@%���l�np{G�D+���kgM9K]xP��%ە���ʧ���-m,���d��x�"�'���'j��M Z*2���O�;]��uK���U\"�'��O?����\�w��܂�+�)}�}�!�Q���hOHl��M�2mB8m��\sPj��|�!��:���O(tb��O|���|�����D��J�`� 2�Ƹx���¬�f;n��D$�/[�X򢊇1k$�#W��.F�V��?���u�	F̧��<�n]}��|;�D�@��ɢ�i�ٛ/��֝7�b�'��D�'��ăG�Щ�v`��`�Iӳ�F�E�8]I��eӠ�$J=h����v��H�?7��4|��5��ܘa蒌7��Bs�[fZ��pn�O$��C�;R��ߺ����?y�'�?a�'�A��B	:�Ѻ��V�YH�d��Q��?)�CMd����y�fB������bV?9z��������&dlTKc��O�P(�'�bƆ��~���?q���*��7u�#���;H�xp�t-��|(d4â�'�ι{���?A�B�?)�'�jp��M�;�N��Ql���rS�9ɾI���׈�&:O:H"��'	�`����O��D��C�.HV,Ҽ-�^��6��yI��`T�r�����Of��κ���y2�۠���4K��#m�ˠ��mU ���Ղ;#ӛ�?O��Dr�ul�k.�����:�V���E�/� 5�l�
E��<��i�<���5O�UY��'5��O\">OLEq26�8U&�!�Lp�ƚ�.�0E�Fj~ӨЊP��O�ʓ�?)�S�g}bE�#7d`�b��[O*���-�yr����t�2Ƌ 6U��x��A�M����?9���?���?���?����?a�#T16Ɍ)��B��Z´�҆��R����'�2Z���IS���$"(D5~����G�!8�UQRe����'Q�''Q���IB��E��ºbf�A
`a4D���+�f���roӕ[h�����3D�� �⍸`/��:��D�B-~<��<D��	�@R\ZqSD�n�d,�'�/D���A�'`�إ'P�X ��M"D� a#�\��YK�bM
`r�D� D�l� �](��I�#B�N��� D����I�iI"�豅��l|a�'m>D��G�;3pD�:%H�/��	4 =D��A\U8L!s��۟dZ������6�y��J�&�˓L�![��@���¯�yb�C�\�b��A�3^���EB���'��M�����`)�%&��[�Z�:ïݑQ�18�Ԃiڐ�U#�9A-������Z)z�{SeӇ�r��S��E�@`J�%�9���c�3�8<�d��1���Q�!��?>�K#�R,�����o�/Zh���;.�^�����6�DH�
((V�E�jߞ(|db�40O��#Q$1>3%��43v�5#�'$"B�I�rW����H�,O:�*c�VL�Zѣ��L�*`�ǕxZ�&)[&o��S�'k�H)��iY�|��0dm�F���&��QaH�O.�o�p�Oڛv�m�!J6Mp��;0��'������S����a��k�<���JZ����x}��
*���\44u�)�΂Q�!�!�I�c]���O8���D�1=0 ���$�x�����[!�D��̠eH�|�Vt#`�� �!��]l|@kc���x���*�<�!�ˡl�yq��8L�����
˷ _!�Dֹ2w�|��Y�2}n�IG��<u]!�dZ�[Ɛd���p����ݽO!��W>]r�AfE�+k��	bg,)N!�� ֹ1�  �=�.9���8ZP��q"Ox�:f�9j�R����A�T6Xل"O�8�L�b0�U��.90�Y�A"O��q�Ş<"�Z�-ȇ{+�dS�"O���peQ�q��Qf��(qj��"O�Hk�
C�@b�qH��D'hQ�,*�"O�8����5h1�Ad<Ї"O�q%���$�àO�4N阶"Oʔ��Nm� �� ("��2"O�	r��+&)�)�V����"OB�ʃ�[$`0x@�2kZw����"O�� �-�4"� ���2)�<�#"O�mB�#(1���D�2:� hH"O�S��q�.(�C�7R�`�"O,pTf�p���b Ua�D<j'"O,1Y��'W(�h3O��z�d��0"O�E��C]� 6�Sfϖ�4v��"O��{� ��|9����X�|,ä"OPA�3�� (�`��yxv�YU"O �a�L��eX�0�Sonٱ#"O���+�����%��%e�d�"Ov�S��A;~�X�YG��"O���*P�>�|�A��9�7"O�z�"�k�x ـa��S Z|q"O��$�
Z��<"���fﮬS"O¨Kр��'�Y�RN��[ "O���Q�L0/ ���G�r�fi�"O�4���
~�4�[4[��S$"O����Ӡw���ӭ�7N2�U�"Obm���]�^J�b�L<qD��x�"O�8�`�Z =M9�f�6 1^9�"OLu�s䛆u�Ղ��E �|1�"O��1G�|Ċ�+��*B}r��t"O�Hj2$ܼG�L�녔�b#�"O>U�3�O�>�B"��-$�I�0"O´2g�-u,�8jg�Q�A�HP��"O`�b���4�&��7M�r�
�G"O(!�biN1>j+\�L�*Y�s` �yr���z���#SkɊ@�*�S�hǽ�y�E̯x���J�D	|ax&�-�yR�G�ke|��׈U�P�N��1iң�yDכ1.�3M�D��l�4(��y"O�5~2Zqn8:�����N@�L!�Bk|�}#���QM�m�wg�^�!��n;���3�_�H�j�I߄T�!�2�AB!��'>��a5"ޥZ�!��ϸ �Bت�@R�W�~����e�!�$H�U�8����=�v��"UA!�$J�Ƒ�ԏ�2a�.�ՀP6M!��)�к��ݗ*u�*`!��U�8�dqs� �k�఑�DV��!�� �z�3���7��ਅ%G�M�!��i���[4
T�.�Xlc@Cߵ|�!���&U%�Sl� 6�U:�h��`�!򄁳m �K�:l3�����!��ʃbKn9�A��I=ޜisC �!��U)Լ�ąƒkET�c����!����,0�T�#W?d�� ��%�!�H-d�v�J�O�5*t�"��I)~�!�D��2�QSӄ�|�%���
.�!��
/�vD���V�t
:�Rd�#�!�D�|ư��E*�B'�	#$��"`�!�_��R|B�jM>�ݚ��B�(�!�d�AE�͈VBg�*�ˍ5!�� �A�g,_B�Zd����8�Naz!"O8d�4��
h��yzC�Y'7�क़p"Oޱ	v�N�wc��[f�N���$K5"O��2�#�
G�}�T)�*7�X�Qg"O� �Ţ����H�;s4٨�"Ol�0'��AQ.��"�	,~X��"O2E˓I��3��D�p��$b"Ob	AP/��X��*��o�HЈ�"O�9�p@ �k�(bp���P,�"OB�hCK��tn����N^�N��z5"OX2��P?��e��CǓQ�Za!�"OP)�s �(n��X�b˟S��dhf"O����Nӑ>��y��܄�ީ�"O(`x�	X
��d��b�o��3"OJ�s�'˞V��;F[}nQC"O��X�B�G,�)��&�]RH�P"OUT�/B0�#�J�
#bu��"O�Ep��G�&�	�D'P.%V��B"O�`uӗUQn�#�P$+ �@�"Ox�a� L�<@�*^��5��"OBL��!����Ƈ�%5�v@qV"O�ԩ$F�*-�U����>���q"O�� ��4W��{R��X�"DQ�"ODa+��	p� D��+X�g�0�J�"O<�j���!4�<ڇ
3�Z�3�"O"r���,ed��%�J��e�a"O����-DꞜ�@� �Q`�"OU�
@ojA��bǴC
dІ"O�0��~�|@��C+�]�e"O ����$���C�*+NU�A"O�A�b�%|����� �6���"O,�9T�
4hPT��ʀ1��M��"Ol��fo�>9�4j��׽5m����"O4�j��#*޴�:��F�*v.a#6"O`��B��W옡G�\&t��	�"O��,P�mGĨ��"�8��  "O����#Nn����w���F!P"O0���dا+:�WO�c�b�J@"O�,C�]� ��݉$N Tr��c"O��!�ʗIY��͚]���(a"O�,k�)��)�4����|�\B�"O�Ȁ�dM-J�e�Iܫ~	�X�"O�횥�I<9ź`�Y���aV"O^I�a��Pߊ�S1��#�0�"O"���3' Rtk�Y
���"O������
�x��B�DKr�`�"OX�@D_�J�dxUHS��"`�"O��4�M>�JYCrȕ�Z�Kʍ�yBI�l	���:j�V��C�\�yB�U�:r�Uh��N]0�㗶�y�I�S[6E��Nېy�R�
�yR"�_�4(@`�F̐�㌏�y��ko`��(L,=��U�#/ȱ�y�n[�'O�l�ŭ�3��H�����y2���Y��Ea���,%H����*�yr�B
�$\)���#J��f�(�y�ެMj|
��]D=@��(d�B�	f���V�6��t��ͣM�C�I�.�Ե�g��hЌ�i� ;�C䉨O�<�p"̚?J�:ec���3�lB��6e�b�qtM*�"ɳ&��Z�^B�I!@��)���f�\��7`�0/��C�	+n�n�� Ɯ|����+R"!�ܓ(�N�X�%�4��!B�08f!�� \��A* a?�m�I��N�:c"O<�1��_�`N���) ���5HS"OM�愐�g�h���ْr��u��"O��P��O��2�Nʜ9��"O
�
�*ЬH@ȸ#d�A��8�6"O�8 �/KH��!g��8W`��˧"O�����Y0����ĳ���ɨ$�!��3�l���(g���ЎH'T�!�$�<�l����"%�e���!�$]m�V����Y����d��!x�!�8\���s��Y����
]�P�!�Jc���4,�"�����d�!� ��5%̀	Z���J�y�!�D �~�M�V��(��Q��A�8G!�D�W��`�
�+�OO5%!����)f!"P*i1��!��=���{ad�� ٲ��
,!��4<��+�iT�H.���!�.6�FH�2n����q E�5�!�D�@,z��t��S�4�kG��!�d�*
���
v�K����q+��!�d��vr4�)��(Y
�H
/�!��"�s�}U�	�/� ?�!�ĝf���0U6[��-�2s!��ڮ��ܩuK0�.�#N�7Gd!�DL!~7�]��NQG��9�*ڨT!��(J����V*�)f$����!�To2TZ2`�.&H���� y!򄍽@��<I�feN��1m��!�dEkz��ҽWf9���D/9!��G�v�p,{6�[�g+ֽ��j]6gD!�ǓK`��i��s<���R�>*!���? (��ҎQ�@����4�!�E�j���R�NԲ>�hAZ��ƋR�!�ğ
	x�Pg�N�����l��7�!��\�|Q����_)=�&@v����!��j�F���] y�Q���2�!�D
R�D{Ăוq�F��$��>f,!�D�tC�P��7&�0�E�\*!�� ��Œb�F��D��cY;(!򄋂4I(Y��CD	���6��%�!��W�\@�<y%*[Mp�(����JH!�Z�K_u��m��ub��Ch�#����	�R����'Ӗu��}A3����y�(T�e���Ԯ_�_;��cBl�y§L{B�@� ��R(�YP�H��y�����`h��{,�m(rNF��yB�W$X����B>"�rL;����y� U�n��:�P/[��p���y�9���ҐD�P`�!�g�̀�y�!�2`���3<��K&[�y��[ I���`/<�VTq��R�yr�ʒyeJ��&*�/y,yPdI7�y"���K��dC��H� :Y�u���y���8q�r`xǤ�6�Jl̑��y�E�_� ���gG��o�yb��^=��0Ҧ�4F��T#D!�y��i�jYY��/>)P8�S�ybH̿Lg�%��2��[B�ұ�y�,�bȠ��`DJ��͹�ό��yboU:
�Bpx�JL~�F5��BS��y2�]�%�@�2��uF�E��U��yR�]�e�3X��9�U�L�e,8i��W&�����,�ye�y������"lB@z�I��ɥ�y
� 4B�g�%H���oR�R�ʵ"O�E f����r�L�9�<�1"O��C爓�.�\a��X���!: "O�D�u'�HO��CC�W/g��9�4"O
� c��D�,�RK�/�¤C�"O4Ej�bH]�L�fHV/��3"O,�Ѓ�M	+<���ါ�.hY�"O�X�܊el%X��˗ ?d��"O.�x�M��>Un�Z!�%/.(�'"O^�3�%Z�;3���p"�R"O\䱵i��Dc��bi���S"O|�(j�*;2]{�c�l� 8re"O>�Y���~ڰ��t�
�c"O�I���وL���{i&@z�Q 5"O�Y�k˱%S���ǲSu�J4D�؂���.t��t#ªJ�����0D�����;;b��k7e�%z��,	4�;D�D�Ν8�Lq�h5Y��( o<D�(�"�[�(�����Bа P��$D�����	��C��L�R�5�?D�tN a֖�j� Ȓ7B"�Q�<D�0��C/'hI�+�:cEFt
�l=D�0h"���k$��j��('&&ʑ@!D�tkB蘰^Y^���Ij6 ���:D��3���v�Ҽr�H�*!�P��$8D�`Z6��������<<8�i*D��a�+��T�Q�Tr�<����5D���@�K��$���L%2�i�o1D�\Z4���Pґ��U��4i&�<D��Ƀ�14�B�HC�.��@m:D��hF�/&������=���9D���qL*znڸ���*a��� ",D�L�W�E�
�Ȍh�I��xu���L)D���U�8���ʤڟP� 27�7D���4��v�6��� X6vu�V�6D���f$�@K�h�̂-;j� �5D��ZdEY1������h���G�%D� 83�%r� �Ɓ�gb|i��(?D��V0x ��c2M�v�L��'D��� D8b�T�1#	�2 0�� �'D�����3e6L)���h (�m#D���@C� �y�+M�dZ*��g D�4rt�ۥy"�P
td�2g�.����,D�D)	��/S��ʆB\y.�; %)D���4g�%� h�C��[��I�.(D��Db�,dB��!2�S�3�] 5�7D�h{�-ΟZ�TX䐡�^��5�2D���k��#"^,0(2Q�<����%D����E�'�օ���T�	��!'"B�ɩ;�ذS懆�
�j�l��K�,C��*}�Q23�Z�8�ᄊX�xa�C䉎z�v���Y� �}��n�?-�nB䉏N�nfgZ)	 �\�'"šW:B�ɮ+JF���ň/_fn r��FBB��:(>4�yR@ڳ	2hFC�I�B䉡��=�4*�4M:0u&��A�(C�	�.��T���
9�$�3TDM�bL C��0׾�:d�0�GώNQ��E�1D��`�$N���ZeE5�2DM��yr�� F뎡phɢUb1���=�yRO̩l]��2�,��H���$�S0�y"�ǆ?�f	#GdP~)V��-F�y����%���1��é?+N�$C]�y"��f�x���HB�o��Ÿ ���y
� 2��U5O�`�1�C7*~� "Od�#�ȝ���H�H��b9�U���B��g��)c��QA/יP(��v�������@\Z��1�D(��
�v5PtN�1�>�i�\*nG~Ņ�4*�-��#jx�(I�m�7�4���n5uٟ~ԁ���%`�40�ȓ[�ŻH*W��� �?I� ��iզm#�dؙs�j��o��/��i�ȓRIj�i1��;fN�9J�ǔ4~��I�ȓ.Ȑ����)j	�˔��%b0�ȓ �
�Kҏ\�,̐���eC�R�L��ȓ#VPۇ�G�(18�[Р��Z!He�ȓA��]I���$1��yD��9ⱇ�?L}���ʠu�(e���=T�nц��nxq�$�6\����C��_1BI��a�Ν;ƈ�2
�$hPCE�`�2M�ȓ%���K��\c(�#�����q�ȓ5�b=�	x&��5&��d��i��H���6ꄕL�&-)фhI��b4��˜:5��	5��so�A�ȓg�(Dp�*���,�`e�ȓV0 �؀-	W��TDȊT���e��`@����h�� �~Y���ȓ:S$�!���,���(�Ոr�!��K��a���{��� �BA�'}t��E�,Hh�˄=+(���?~�\�ȓ(�=��A^��,���@54��ȓ>`���F��,�n��ƛ�D�x!��m�b�Hǎ{�d5	R=㾝��xaJ`P�ɓ�eN���5.�79�2M�ȓ�|X���?9(ăE�HD�����J�lA!��t���9�*ӄw���ȓ\�}�(�"]{�ag�D�`h(�ȓ)L�<��:!�������>8��w�p ��0Ղ1�̰{NV,�ȓ^#6�xdl��Qg`I�!ǋ=�����)����3�lt��ˑ@V�Vr1��uz���4m�90�4tK�*��%�ȓZD��!h�z�v�@����4�P��ȓ]5z��t��#A1���GC�*>z=��6!x��/��8;7���3+�<�ȓoq�<�T�֓r��������P�ȓR�ND׌��f|t��3�A:2�M��	�\�egF3�Vq�@���~�����8R�,�Q�(<�d`�%@����m����3O��"ٓ�a�J�b��S��sr��0R�V�P�<?25��HM�� ���jnD��@VN	��$6x�2�`�*X�x����$�bi��^�TZ��#c	�xG�	k8u��|�v}���sgJm��;X����,�f���@��j�3f�8�<��QK(}�ufD\����䉄�dmI��r�����-S7}��� J�}3�(��\�|���2E6�@�ߦU��фȓ	���2��P��L��h�.r*��m�N��'*ĵ]6���l^(j�t���c*j���R�F�� 3�/��I���ȓ{�Ik҈���x�A��?����/��� '�I�)������4x���\4�qJA�8�4I���ˆ!*�Ȅȓ[�҉A�GB�b$���m�n4�ȓJ]r��-<�H��")	=jP�5��S�? ,H�k��CU���.��*Ҟq��"O��
�LͼT"��Sq���𕢶"O������5�<���cךX32ѡ1"O�Y�`�DoF��P�U�f�h���"O Y[Q䒋<�|����T�
(�y"O<p�Y��d��� �T"O���ȨfNd���
5#ǔIj�"O�̓�����j�>s�i����#m�!�T�Y"l�"a��h�+�$I�!��@�:�:�i�]Kb��׈�u=!�S�dgp�Bf�=E� ��%]�w4!�߰4 ��1J��1tM(���g�!��سOdq�`FA�K�P�9��S� !�_53>ʉ���,(%D|��|!��\� �x���_+2� ���M�!��>3��q�@��Ln��*�G�!�� ��$;sA��`O[�×�!�$˵~Qj��W�*@vA3s�W'�!�� B��(��g��#�����^��!���)��-�f�P�#�nQ ��(f�!�� $8��f�z���b��&&!�5�r���ґ+�V�!��/�!��_�f��Ũq�P�0���O��U!�D�	(��(����2��
�G�Ui!�䏆h{P��&I�t+2(�G`AM!�$ޚ��{�����ӳ&cX!�N�v8��ƬN�M�,Hj`#B�!�Ѵ?���2��)mϮ�pϟ�_�!�䜬%���C�[0�{�cޖC�Ɍua������x?`��ǦB�\�hB䉈}����ӏ\�⌐�L�p�C�I���Ģ�j�vm�`���B�S��B�	
S�`�Xiэ!���p1bM[��B��/�а Q� ~��@ˍQ�$B�	-r>l��pD@8j�J���ԁZ�8B�I�d�>]�׭5(BMZB)/B��3_Ҋ���ԍ=��B#bSv�C�	�=� }�o�:A�ys�_�L(�C�	:@mZŊ�l����:������C�	6W|�P��l(�I��*H�7��B�ɦn���@�?x>�]��� \��B�I4�}�X}��
 �Ӿk��B䉌5����9j&>��5	q�zB�ɩ;�6l0g!�{t��B�L�0�JB�ɗpz��'�6&�j�Ʉ+�zC�ɾA�Q�1��nA�q@��/`C�8f�U��¿%� 4M�70�C�85�<� L!8�� �t¥o��S6H杚5�!F���� �!��d�숖�[(��|��S'�!���"s� ! #4�4,�����O;!�DT��A�a�>y��=(�$.W!�<�\X���'*�^A��j�$!��Evx���჈�X�+TD��K!򄈭ft(�Ő�m:d1���^!���	��Xٖc5��y�w��5z!��BVaV�u�	U�<��2�Z�s`!�DҮ����%��y����b��"c!�Dז$_"aX�h\":p�Z�&r!�d��"LsJ��+u���4��X�<I�$-�xB��/���۱Hi�<q�KB�n�&m����)'��K�F[�<�e�S tln|a����;��s�<�[� �[�Ϭ������>0�B�)� �����B��l|��+-C �%�"O0p2�̛~��1�,s�0�"O:�0 kA��#d�+�4$��#�6pQ`ɹ���L(<O �@.�k�"0@C�,��y��"O�+���6M����N�$�*QxF"OLX�����d4�n�%4�<}��"O���2->A|�T,�0^^���R"O�	H�F'/<v@�G+�f��e	 "O�����8P*�՚aJ�=i1�<��"OƤ8�.6Sɦ�q6�JR b��e"O�X�u�ɰj���1�A�{�ѥ"O���$�;_��5y�)�<��C�"Oj�rsM�<�4��IS�U�%"O�#�VN�}��犬JQVM3�"O��Ã��&�nUcA�[�r���"O����O�?0�!���m|Ux@"OЌ SdURk\��!�� ?x��v"OJ��7ܑ�i		%��9d"O��3��ʪB�d�Ȳ���^�K&"O�p�!iI���<�a��&5���c"O���AL?\���G�U�B�p�"O�a�� �S���r����PS�"O�a�#�|{���G���	 "O@��!	�u�tps�B¶�b,�V"O�9�\(+oZ=��@%6��0@�"O���TDŽG�,`*��-�"C�"OV�a�Ê^���U�+~⡸�"OES�D@�9p��*M�xh(H
3"O*QGDX� �F�:`g��3n)��"O0�j'�ַ{^�X�C�x$��"O��R�K٬|���F��y|�]J�"O���!<.������(]��S�"O��2�J1Z|]c�i�*Ӓ%�a"O ���"9\�R��S�*B��"O�H�%��y����&q1�"O>�⠊�pG`���j	(�"O8���ӫK&����L9|�\��"O�����F6�LQ�D[%_��Pu"O���@,��CŌf����"O����Q9M�܊��e��ɨ7"O��7C��;p���b�Q�F쀥��"O���(:_D�+5g'+�u٣"O��9�U�-��qQ B�l�x��"O�P2�Q�� M����DA�̊U"O�E�Uè�����-�,�p�"Ot��UB��|hh �6�u�RX��"OB=�e,\-9lfLIЭ�9�v��$"O�KR�-V�t�pl^=�F��0"O|�@DI]�-IǪS�!E���"OZ|/Y��(�A*�!�X��FU3�y�ʊ)H6�`��dY\K�$�y"�@�@��ԧڋU�҅�GL��y2��<�l=#s�^�?n�x����y�腌0m�ط�"8(8aXwꗞ�y�l/�J��bl\	`atX�V��y�.0_z�kGl�Z��vƐ7�yB�!z_�:�Ώ�Mn��s�L3�y��\"]����k�8բ����"�y��n�NT*`��'-�ت&iK��yR��# u�d��"�NP`� ���y��2!���׼� ���́O?��ȓ4���!c/s�V5)���2:�V9�ȓ��z�D��y�p0 U2&����s
������.1PUZ�#��2� }��S�? �9!BݝFx��g%g��|�"O�h2�O�*G28��@7c��(a�"OPu&O��`�0�2��t9����'x�@`c�ŌU,�A
�j��4ʝr�'JA��	xUF��IH4$W��@	�'�d�;1e��W=�����S��0#�'~(H�����lԺU�L�w6 ��'14Ab�o	�$��@uDSt\p	�'1<��p���}��@N�e�f�(	�'�X���%K�m�L�IQ[LyS�'��y@&؎W�\i���]Le�
�'ݚ�H�A�Gc
ى4�;Y6��'Y�T�W��M�4	D�BXL�	c
�'���0w��'� �@5Wx��a�'�(8#T��5r�؝�#�R�"��'��an؈\V$��%��Wf����'�ڹ�E�B)�Z��F+T`Ņȓ*���2�@�p�h��P'tV5�� � ��OuS�P��b��~��ȓR���0G(���Z�m� �l���Q|����su��b�i�y�dY�ȓ[L�A#`'օ{~耴�ů*����ȓJ��H��j��0� ��bmL�Zi�Їȓ\!I���	?}6�pA�� �zi��e
��h4$]�H��u����6�p`��J��l��� ��X��+%�¼�ȓ#.\|y%b�9�\���԰s�H���u�����n���}�DDD6��؅�#y@y�P��6
#�M��i����4+B�ÔÅR-�Uk����SܴY�ȓC�� ��ݟ.4���KZ�P�ȓs��:�O�֌���>g)T݅ȓ���*��m�|�
�F�7B:P���p5�� �䔪r��]�w-��5��݄ȓ}$l�0V�)p�����̱Q*��ȓ5߀HJDꈊi|�TA���!�ЅȓJ�\�D���@t`��ЈP7�-�ȓ�d�V��g�F�&gow�Նȓz���H�/��[afP{�n��9WX0�ȓpB���@Z�����R����zBV$a�#��5c�*e�i���� �tb��7F�ir%��@$�ȓ+P�lid���cRq�#�����܇ȓ]�>�C�d�n�Qòm��Ӫ���B`�zD��0K�=#"�B�aA�e�ȓn*(�3`��P�Q���P�_h�@��?���3���H�CR$>��_���ǩ�3��� ��'��܆ȓ3��i3Wo��g�N�8��[�t<��ȓ#EF�@�,|���@ �6X����6��1i�H��1u܁0�lGTjp��a~�� ��EC`�9�UQ���ȓB�D1�h�,fE���(e5���ȓR������a�켹��˶h� M�ȓ
���̊8)B.x���E+HJ8��ȓA���x�^U���W=n1���ȓq�Z� adS�9�e�۝\0�ąȓC�qx�Kڗ'Ll�	�K\�J׌!��yU(P��LK�.Z���@�
�'\ў"|��Y���IboK�����B�<)�&��A|q�c��Z�hI��A�<1��rd�^�H�<��"�Yt�<����,@��X�FB�P��%(�s�<���"6��1gn�zQC�m�<� ��qGM�w�HA�O�^���3"O����F�B��r�΍�z�rP�"O �±dߣ5jN$z%�#+�pX��"O��d��"�(��p�P!*�V�["O���.��$i��@OS*��"O֑�G�W�Ų�fA�֤�*u"O��KB���|��E�'3�4�I�"O�1���|��Ey�D��� 1�"Op0�*߭���;� 
��@�B"O��fшX�,�`��6E")*�"OFi�P��٠�:���(�R"OR!��{4hJ����1�d��"OJd��%��H�=Z a� �*e�"O��kUw��(�/k�T=�"O��UD�%X���`ρ1��5s"O��[ta�+����[c�R(��"O�sV��.x�:����-~���"O6���&J�N<!F�JJ��YB"O��@�#;?��a֣�C+� q"Ov�#��q&Լ���Ӆ���"Ot�c\jL�zEaĶ;��8���A��y2�[�:+�Z�F�AV��P!��y"HJ5ehR��#ں%��|U+@s�<ag�**���O͍�F���E
X�<��o�S=�t�0�[�I"��e�x�<q�EٜN} �EQC2nTpE�Ut�<�,��[���y��N$�.��4GL�<ɳ�G�7?���Ǣ�:����Ph�F�<�d����@>h�biᕫ�g�<�#I�?U����G�'�� 9�Ma�<�Ӭ�1f��}X0IA��� �#��H�<I�)U�D�Pزdb��J|�-�Ռ�H�<fDŕ={����,�'�)���}�<�0�#Q�JT�e�;%���8���{�<it��l���T�ضG�,mxQ��z�<1t��^���Q�����e��u�<���,?=����L�&x�l�vALK�<��N�H<�1��@�r�Q��k�<���3u�<��G�[v��Ȋd	�g�<y�m-^~���@1�f}�v��n�<1�eՅ'�i� X�e�B}�eaMb�<�e mfa�fa�%b�`i�7�f�<A���w��a2�g�:
�HT�1 �c�<Q�O�GsZ�Q��93(r���Bu�<�S�_���90/Z8�K�LY�<���ּ<{� ��U�+�0���QI�<�����:bbP��I	�d�_�<�RIԣ�����gR�Y�0�G'WZ�<)�셹 .��a@�,P�1x#��J�<��nԘ8o���Ќ�2-΀�i0�E�<y0�LV_X�z��o����ď%T���%��:�Esv�E{�\�)��(D���v��
D�
��'��.�2���&D��FeK�X�*�Y��E��"�!(D�P1���'�@ᚖ	��2L̴yc'D�����C�଺Q�ߜY����o/D�$�C�8e�%�^%�f`�d�+D�LR�oW�k��	Ѕ�ێr��Y�Rn=D��Y�l��(��w�Z�#��x�!8D��X�ɷ*dj ،�V�S1�5D�ę�l?IL����� ꔬ3D��l�K9Hi��ǯCª$�YaC�I�VDdx1�䑶:f�2�� ��C�ɼH�|�V&Y0 X���F�C�)� ��Q�Q�@4K a��v ��{""Obp��폭P/t�:A�2��g"O�-��%הmz"yieG�д8�"O��-��'� u���:F@k�"O���DQ�T̛�g)=^Ni�"O��v���p��f
	cu�,�"O�)�E:��}[U� �\��3"O����A�}<�y�Gj�gI�es"O�uaT����J�i��6x w"O��T"��[XT�A�H�&NV5z"O�H� ��lz� �⭆�25��3�"O���ã@NH5Q�OW�;2����"O6|��G�^ݜQ&�_s ~��F"O�P�`��#e2%;4�SjJG"O.@�4*_�so�u�&,��"O��"7$�a<���G��t��XIG"O�aC�NT�5�䲴�Ņ�:�"�"Oĩ�G	H�<�ɥ��6g	d�"Ox�;fFN4B���C��1����c"O
��P�^�p��g��9��"Od��F�����^%,x���b"O$�ۅ[�[�]R�i��f�܋�"O`�ڄ�ݭH�Q7�7�x)ç"O���{ b���
�>����E"O�]x�I��Qz��!`.��ʴ�f"O������9��Q��M��.|^�z�"O U�d�� y��+3��8^a
x�s"O�`�TBțtB�8
#�Ag,�)I�"Oti���r�	!��T<H�<Z'"O�a�g�Y)Ԯ�ӊ�(x�J y0"O�T"�%�5isV��婏�)�4�s"O�	S�+D ��a��狽V��Bq"O<��r^$Xm	�f�6~��`"O�A0��%\N5*����K����"O2A3�K�� 0�#�
sT��E"O��!���xQ�S#�?0Q�@�q"O@3�~cl����HT��в"O�%1#� �H�v�:~�d���"O�i3EW
}Q��R�J�%9�"O>0��W~!H�B�g�L�0S"O����Jh����T��7�h�pB"O��� .F/_G��Q�`H�m�e��"OZ�b�SPS�� q��U��e�4"O���rkA/ :!≇9;w�9��"OBU���{q*0�WGG6uh�H�"Oȉ+R�[��D��'g�OOlX+�"O�쐹zp��(��T�<됍P�"O6P�sGD�a���y�nk�@�"O�]4̔�?�}�Q�''��� "O�1q��@�,�rH���ȵpfh���"O����yz�f�ǡc_rp��"O�y��勮y&�$����6GtD�"O��X� ��?��#���.r�<�kG"O�]��b����0����"bB�qW"O���q��4���c(O�T���p"O�0jAKա���qFiA
e�hhI�"OR���	2FG$4���f��Х"Olp��Z>w�b��c
�A��A��"O������&���'�lP�a"Ou3֌Ȼ,�:#G�+<����"ORt�0#��r=���V�X�ror5R�"O���ՁV�ݞ�GNߔ?�$A��"O�PZ��6:�����&)�d"OHm:rʇ~���D�+�D�w"O� @h�W)'5>�=h��ИaFRmI�"O��H�@�P'�4((�m��%!"O`�Y�"P�QB�ѰA��\uLpb�"OV	C��u*�A�`X�i����"O4��d���A��9VN�d2�"OVe:��W"4��͢��1T�,CU"O���3Ȕ���:M�9>MP(�*O*m��DϪ|�	Q�i�!�Le!�'c�Mç�T ^58���A�D���'DL1�`k۽)�,��%���g��{�'�~��	!7��(j��2g�Aq	�'����ɳ0���B��)3���'(��8�a�6WFH$�PE��q`ư��'�[��L q��lR���m����'-"05O*��:�#A5r�>���'sr,k�e2gN����L�3�l���'(�}�f
00Vt���-I|�
�'D�����ۥO)�Ax����_~i
�'s@|���Ζn9|	y���X��h�'����fs~:�:�\�s܆T{�'�A�B�(ԾX2#�&h�,���'f(�yC�ї=T�x�HO]��1��'����a�"qZ�	!�ժV�ڤ�'��|Z1���$�1�U�U�bX�
�'0@L���=D�|�#QxUN�`
�'7���S���c�	�zk2H�	�'�JU�U�vǜ!c3d_�r��M�	�',����c �X6�ݳn���;�'����%��7T��OͯB ���'Np�D��\!C��C���'��k��I�p�H���y/ȅ�'Ɍ)X0���Ѧ9!#G�@�n}��'vB�Cor ��i�/�>�`:�'�4��*Ab���C3�� ����
�'{�����T"$et��)B�~z~yP	�'���:��^�v���j�I�7j�=��'�Zp��oǏX`�@��U4<TyI�'B�-�`Õr4z<! �R*�T���'*ʴhV�˳S�&�I`灧W٬<Z�'An�:F��,�2�����S��E��'v6%rA�q��-{Ǎ�	HP 4��'��uk��X�~8l������]�
�'��E��*
.-(a:V�C�,���'���Cڿj��	&�K�mu��Z�'q~D`	�~HA� *��| ���'T�E҅'Ϋs7����E�'n� 8��'���� �
�m�IRX���Y�'w���aA�x9��P�Դ;��x��'�֕i$��+jh	 ��H]��a�'n���T��{������2:0�	�'L�}"S�5���!R��)%�!)	�'����%H
;S�	��"�Re�'�(�A��֔S����!oC�eHs�'�HĚ��C�D�Mڀ����(�'�ڽI&�%6����$V _2;
�'Q��q�)ܜEJl|H��0X�:)p	�'9�d ��?>��ua�)=B����'��X��:8r��!L�;�@H�'p��j"U�8~nPy��*�����'8�H3�B�!I�v)����V� 4�	�'Վ�1��!e>���SȌ�B2Ԩ	�'z� �b�M�`�0���d��x0ޠ�	�'���[S���w���aa@k�l�'P�us��L���{F,�1vz !��� fM��c݈����FE*qS��2"O��3bɟ��Q)C��X:8�"O��aPᗢ^�&���3l�hU�5"O�H��%�?�����C��4˾�)P"O����t�fH��)́s&y�"O������L#\��(�w%mG�VX���ʐ5&�T+r���x�� �3D�����؈*b�7�\�U[��]J�<9קėZ�͡e��7���r��{�<��j�z�EH����a�jCJB\�<�]�\26T���7af$Ò��r�<�"�Sߢ�ҲDر^; 	S�� C�<Ц�Z;�-�$�ͱ5T�����@�<�JF��*��kƨ1�a���\w�<y���?U�ĩ�V�EԄ���{�<�ˑm(��t@\�P�2���AQw�<pBP\>.��#jђl�*����h�<�1�R�1v���ېnt���e�<��*�;���;,��YcBēe�!��4">6�����w�@;�g�Q�!�\�-�J��Wb�i��;� ��4X!�@<?��p�v��"�8���1U!��˸>Ǭ4�ևN(f���qp�A4,!�D�y)20)�ƩK6��AJC�R�!�]$q�2u��@P���z�kY�!�{֌��$I�+�̀�
ނ0T!�DڅW����F�������#!�d�2r�������7�
�A�؀#�!�dK�A�"i#�N·5�
H��e�@�!�d�5$���f�~��ӀM=�Py�� �D]\�{v�-��D��E��y����H�q��cR�
и�	�Ԕ�y���/�.`a�f����tI�3�yl��*&��F�,t?�L*���y2M�5��1�:h<�8�����yr ٶ;��6��6M�D0k�bO>�y�jڄ!b���$Uƨ�!HȞ�y2��';�<��C�`Xhґ���y�L���b��ǡ��,��]9�'�y2Bvg�Pq�(^�^*%{�!�1�y���Y@��h%�ꤻ����y��ۀLu�lxժ�� A2��y��ϼG
��&���1f�+�y�MR(��c��u^�i`Ņ���y�蚁P�j���%N?�-��;�y�`S;5�Q7H
mR���*Ť�yRnJ>7��p�X�i�����@6�yb$�/�<�����|�B0�C]*�ybd��Q��!�E��
���JB�=�y��V'\�bU�u�,3xzag߂�yR��1�m�'��*�����"�5�y��I�t��sጋ3�]�Í��y+�R}�Tc$
SԞ 9î�y��ּl)��'O&�hs�
��y�NF�s�T(�&ʝk���G�V��yre '��Xb��m�|e��J��y2̊����_~�x�A��yR�W"K��0W��0^���0�O��y��$#<Ty��R�
�$IC���yB�� ����h#L[�@x�+��yR�ȕVц�i�C�w�qz0��
�yҏ�$kX>`�׮�p�:x��yR)R?M���cL�bL~�ꙁ�y�Ɛ�>e��D��)5LAx�E�y
� �=�A�
Q<��;�ᅜz�!P"O��c�����ꜟ���Ґ"O�X�1��O��p��B�	�����"O��Q�E�>Ei�N�3�hU�Q"O�Bu`�|I�J�*�^�ptJD"OH���� � �:���h"O"pKW(I�j՞T!�ӹq1�(C�"Oڐ2ōȺ?h�Ÿ��_�4'�x�P"O��A�hψ+�+�	��Pv�hE"O���� �}���CGB�G�T+C"O��z�˟5�H�8#����J��O��������M���M3�_>�q��T����������
%:�(���I�F�Xq�e� \xԛC%́	qD6�U6U�h賂�N�+��)h�Y��m�9�>��'�"2�xBCn�&�����آ�H�g��7;�����֋Dsԭ�~��$�J����!;鄨B�.��m��U$�d�Ѧ%�,O��ޟ�����bơ�+�/0���?�~B�'�a}2��	3����&��) �<]ⱮG�(O�Im�/�M�J>���u��Ʉ{�}ct�Ǽat��`.�|�d�O��T��:�P���O�$�O�ͬ;�?��>�01���M^HcB�HVZ��`''N�҄��DU���[��:�&9�fJ4���jE?=�H��u��?���q�c�)�F�{�Ț�v��`�0��~�'$���'!V��UOY;�ȅ��V�%��(�O`�y��'_$6�C�'��$w-�lK�#�0�B�s�vL�O>�
��X2p��%n[���@�BǪ-m�Ŧ-��4�?Y��i���O���\>�����0���b�I�pD�}�Vȕzު���̟��	ߟ�ɠn����	ݟt���S�n���ՕZh؁�ƲB��Њ�q�T!Qf��(톸Z��U*7Ñ��:UL�����
 $FH[u�ӈn�1�*˶$Dh=����m��y%a��HO��z�'���c��0����&N�~F�v➾ ;��'������'�p�I~���A*Nx���hh��r֊���yR(�K�>���Fį]�h��Ν�]���$C����4�?�@�irV$ag!t����O���w���r$���J���������F-k@���O��D��\�T���%����Z� �ÝO��@�41t�p���� ��p!���ê|cZ�!��W�#�UYã�wf�ZC��qrZ����0��5�bh!ݾ�Fz��Ը�?)��i*�7��O��'�t({��Ȝvja�M88vv��`�'��OT�}��Т�
5(�6=puCW���g�����٦��޴�M�2D3wk��"�'ͨK�������~?�Ȓ;a>]��?(�N�9s��O�dd����#��)��t�F���jĖ]� ����Ƹ;!�BQ��E�ל9sI��ݟ��'��]c��lXP�E�|"���SR�t�ߴ)n�ૢ
�tDX�@r�O��-�S�@8 ���k��kV��ρzB��P�պe�FM�?��ilF6��O."~n�Dd(�Bh�4ų�G]" M�	ݟ��	{؞$��,�$x���C��Q�q�d�&:ʓ`����y��O����O�HX����3D�̨�D��C>~)�D,�O
���E�xT����Or���O ��Ǻ���M�eŐH_�@��M��o;rp ��d5��(w�Ε~�p�%��H���O^0�Dx���8�(8"���P�ȠdQ�XX�6L�Y#LU��+n}�y��p�ĭ�)=�c��
�N]-��T(!���{"��1Q�>q��Bʟ|ٴR\����'k��h�B�ET�1!��pT�'fay�fȗU�*,�A�L��bB��jx!mڕ�ML>�'��H>�۴-�<� @�?@.���SDӂ.<�%�$��O����O��D�O��<�t�i��%�r�'�*�k�"h����˛��!�v�'��7�-�����$�O\���O���W(S7;�Ftr���(R)P�M�!��7M/?A��D6g���|�;#�B�q�¶��-�1�.�fDϓ�?���?���?1����O�t=(�
�xO�ysg˛	հUP��'�2�'p�6�Ά��i�OX�o�^��&z���6��$D��r�) �C��}&���	��S�6�Ul�p~���0<���Ғ�3C��Y�A�.����3D�|�\������������3A
e����E�ƛ ���ڰc����gy��f�0i1n�O:�d�Oz˧[�ܘ! ��� �cXi���'e���?)����S�$B�bZzIؤƆ!q�X�jp�D�� +����al0"�O��+�?1Df>�D�)ͮ4� vE�ԉ`Dy��d�O����O~���<q��i��m��^)N�lY0 gс~@�@�HF?Hb�'$7�(�������O,9#b��+����G�nx
���O4�D_?Q!V7�/?��
�v����0��۰R
tIZ�"�V��w!R��y�P�\��̟��I˟ ��ܟԔO%U��MT�����sA֔j��t�&=�q�O����OB����D�ܦ�;y[6���ӤD.�+0�� ^t,���ΟD&�b>��!��ܦA�6��5�uo� D�
(B�j�7"<�\�"�M�O"3I>�,ON�$�O��4eR�Aޠ`�GC1�0'�Ol��O~�ĺ<�W�i@^����'�"�'�Ȁ� �?Q	D��-@�S]"̨R��B}��'I2�|��_�"�h�'�6"����\�x`�O�}�GD�(1��6M)��Qa��O Ar4��j~Xhp��Jv�t�a��O��d�O��d�O(�}λ��\R� D�yj@�'ʙ\`���S'��Bڞ(]b�'{�7�4���O�� 1l2��HH��eH�~
���OP�d�O&� �t�n�9��a�)�?��ݴ/�\�����Q��cSIT�Iyy��'���'���'��'^.N]�8{E��;u����l��<]�	.�M�ä��?����?�O~��llP��(��@ 4K�h]>s���yRW���I⟈'�b>	�,?R�����,ՠG�u��C�g=�#�9?��a��*�p�D�3����D\s=���lG�	���d-���˓�?����?ͧ���˦]��A����c@�	
��e�'<��Q���� Yش��'#$��?���?�@�"����,�&?�!A��(�(��ش���mS�)p����O�����I��1C��=�����J��y��'\��'��'���IW�0I����G�(e�e��+�dEp�D�Od��Sͦ��h>�I�M�L>�����zsm�4�@Â�Y����?���|#�K:�M��O�i�b�׊{4� J�F��,<Tk���_tR����1mƓOV�S��<A�o��]�.5+��{���۵B*|MGx��`Ӡ�b1��OL�D�O˧9c�H�"��]�T���,��B���'����?����S���"{��tR�*B�C���Y�N�X�@A���^	�"�	0^��S�zFR&�j��بXq����%sS(�1HBNC���M+�E��w,��JXn����]��lQ��?I�i��OTX�'}R��|�
up.�.|`���W=	���'*�E�i��I�B]���۟��S�? XQ�l[�\bءFNX�Y7�y2O�˓�?���?A���?����	�>�� ��U�L����!C�nxYo�?N����I��P�	~�s�����Cd�Z��u1���94Ռ��(�	�?9���S�'3�xD@ܴ�yb��.m��9�4��g���3�����y�Iq��	?sA�'w�	Py��|p��[2|y "�ɚ�0<��ii��u�'FB�'�������7��&i�t�X��?��'H��?����w&
�ũOn=�R�+�i��9�'�zT��S���4����~��'g��rmVzªu��Q�H�*r�'�"�'B�'@�>���51��Ţ�(|ڼ��F���i�I��MÆ� �?A��Z{���4�0��̊7�@Q2�²G�܌b ?O���O$�ĕ��6�7?����2=����F��#�S���t�'5��I%�ؔ'S��'[��'���'k�B�ʟ"O���q!Ŭdf��6W��޴/�*!k���?A����'�?�1W3����aM�����ff��,���柌�	t�)�Su������4(|p�ʆn��?R��Q"Z����b4���O�a�N>�)OX�״p��eݦX��|�fH�;e�����Ox��O��4�n�*s���"^(b/��fp�. @;P �#��O��Je���8��O��D�<���<v� tH���4** ؁,�(>���rݴ��D�S�T�J�����D��̉0/^H(���� ���T���~����OZ���O,�D�O��d/�/���Z)�9i�o�1 �H�'�� `�>q�W:�n�^Ȧ	$���b˙�@���"�ڞ4Q�����[�����i>�2ͦI�u���Ġ��AL	$[� I��a�l 1�'���%�,�'m��'Z"�'��5qu H�g<n(�U-˧[���1��'.�R���l�+�?y���?Q.��x���9+��s$�0=�$p ј���O����Ob�O��P��Kw�	aSV��橑o�:�u�_?e�@��5?�' ��dJ���Y�(��D�	s�����$�"s��A����?9���?��S�'�����%ۄ�2�099)Ɣ#�ʴZ��[=V5�$�	ӟ���4��'X�ꓺ?�	 �IJ��`7KJ$Y�h<�!n�2�?���8��Ѻߴ��D��6$�Ɋ��N�2C��C.�:�뒆�yT���I��x��ß|�I��O�de��T>tR�AF<f7���s�r�y���O��d�O��?Qi���ӧ�J�Shts��]C�A�ӏQ�?����S�'t�Q�ٴ�yr�(P�� M~�$��C�;�y �����ɀ[;�'��i>��ɂ,���pn�'#�z����cr���Ɵ���ğ��'W^6-
�r�.���OD���zmR�Q���%)A� ;rk� ����x�O���>���4,汁q���u�D��Ɠ�O��G�(��!�� h��2I~�h�O�z��H��@�S�X�V���^�y Aj��?���?���h�L�[?���'#W�;�Nl�p�ȅ0��DH�3T��Hy��|ӈ��3n*� Шƺ"B�ڴ��k4
�	����'�z�#e�i��I�M��U��Ok�_�H��c胸Iz���f�>3��'x�	�8���p��П��(��`��I�'}|$�ň>��Ԗ'Ӭ7���m��ʓ�?�L~���x�B%�"&�b���6$[��RY���	̟(%�b>��W�T 
[�P�T��#cV��;�a׿D$T��EGy���]����uU�'�剩p��I�$oM�)Z��xeQ#l ��ǟ4��ğ��i>Ŕ'^�����"N��7e�q[�: ��F�U�P�� {� 㟤	�O����O���ˌw���"�̐�U�xEI��:��t�C)fӘ�v���"c��\�>q��v�4�;R�D�mR�tc塙�q=2���� �����Iҟ8��K��%�6���<zq*ċ_+VڰAx��?)��a���УK�ɚ�MKN>�g$��k�`�� /+�)Q����?��|�A@Ѱ�M#�O�n����p�RH�j�dᩗ�ݤ(�8H���O �L>i(O:�D�O��D�Ox�y�+E^���`��S�{v��ip��O<���<��i�r�ҥ�'�B�'\�S�W�XQӏ��0�&#� @�`�.�������?�O�a%�$���ga"?[8:�!̅ࠁ����9^�i>��V�'�\$�HR�-M���F�͙:�	yp$�쟘����\��ԟb>�'��7��2N�!M��3;l� ֌�� ��XZ�`�O��K˦��?�AS�4�I��	�bW@~B�
�$��t�	ܟH ��E��}�uGgWAy�$uyb��(4�=��.Y�{��@���
�yRS����ß�������	ҟ��O��A@K̑j'�%����(@*�`E�tӀi�@��O2���O���0��æ�ݙ>�Ԭ8,:p���-���*��ҟ�'�b>��PA�M̓'Ѱ��$Ac6�kQ��5�hEΓJrL�Xv#���%�$����'Y!�q��5Tx��ޗ,�4�x��'YB�'�RX�TP�4.[�8
.O��D�2~"%s�K���Aף�E�`�O��$IY}�'���|b�O/[R�<{R��9��!�"/Ǜ���?sĹಣN�2��������7�.�$W�5���h��	QV@A���Mh��D�O����O���3ڧ�?!ǡ�
^R<�"�V(	����W ؠ�?��ij�e�'�r�`����] s�:�a��]���%*�*t��	��0�'�
���i�I�]��RW�O�:� ƍ*�Ξ;���/ʎG*�PC5���<Y���?!��?���?���< ��V���6��г��Qڦ��3_|y2�'��O�ҩKx���K�+�S��	g�]����?����t��Z$�����	�*�*���9�����b��I�:��z��'9�5&��'[.�÷�.,��٠Ṃ+��̱��'Z2�'������T��r�4~3b����BL/r�k�	�4}�<�0@,�?a��i��O��':�]���L�4D�T4sR���b��$�`���VMt nk~�,0m,��$��Oew�HQ������O�Y����՜�y�'EB�'N"�'���)L�6s9P.C-8IV�˔E-v����?iw�ip��O�҄u�ΓOh��dc��3H�2P# �&��x
3�&�$�OT�4�=[F�~�f�Ӻcf�x�&�
��0Y `ep���x��(���%���O�ʓ�?Q���?��6' �b���瘝��JR�Ա���
ٴ�����r#D�̟��	埔�Oڄ���AA/�2m���a2�O��'���?M����,O�����AҚ!V���J��:�X�q��ۚ(����ԇ���x���|"��37ڨ��vj�U���;5�Q��x�.r� ���˰�N-�f�&���p� �p���d�O np��y��	ΟD�$��yi�U*4m�WI^��Ԁ\̟��	��qnZJ~�f^
m�]����d��3w�x�`��H9v
��#��<)���?����?)��?�,�� YDb�/|j�d��A8xf��0@٦��jMTy��'L�OrFf��.��<��c/�u�n�y$L�#�R���OF�O1�2�!fNb�������1��B��xsk�!P���	��̍qP�'�v='���'���'��#�NA Z�^��G)֬P��I��'��'��X�H2�4,���#���?����Չ�� �2Td@k��Pq��"�>�����'
���.B�Q)��X ��&x�����OPq��^%b�إ��I(�	ߥ�?��i�Ox��C�
�:IJQ�ƴP�\SSi�O`�D�OB���OV�}��Z#"9��ŝ0|�Y�qj�4j2 ����.ȲK7b�'�t6-'�i�(s�@�2�|�zT�Οs�J�� jk����ʟ��I8H|m�`~b眬R�<��S���L����(C�� �/JV��q�|bZ���П��������$(�C^�)tFp��&�8Cx���7��Sy�kӄ5ӡ-�O��D�O�����_�|�ȅ"���q���G�:��'1���I=v��p����Gc }p�M5�1�Չ%=�˓yH��d�O���L>�.O���ƍF�j�J2���i�E�O����O$���O�ɧ<�i�  ���'8�}ap	��qȴ��� a��T��'��6M/�	'���O�ʓ����)
:
����
R��(�"	�Ms�O*H�cD+���.�	��~�p��X7)�&�CC���KVd�h 2O����O����OD�d�O�?a�� Cbt���LΘ?�BA@������˟���4Z,U̧�?1b�i/�'u�%�4�H"m��L�9��\aЗ|�'��OZPXZ#�i��	pg eI���
��sA"O�l� ���D?�Ī<�'�?a���?���N,V/b|!@CM�[�Y�a �?�����$�ͦ)�V����	���O�&�fK�t�4���,эFɪ���O��'���'�ɧ�	�
pcH��w�	$t<���g/��5�A�}�"@�ɺ<�'s��]���]��@)]�n�`XZ�ɂ�Pk>A��{���HNvm�'��O�Fd�`E��X���'F�JgӤ�$�O��N{�ZK`�G�v�����J#k�����O��Cr�k���W���S-�?u�'�� x�b��d��@ 7��t�V횛'.�����	���I��d�Ia�T�V�8G�=�L�'s���P �7I67m�?i~���?H~
�3i��w�hS�)S?����#ʙ'F"E�2�'r�|��"�"<�V=Ord
G��)(�r�Z�D�)�f:Ox��K�,�~��|bS���Ɵ�9��
(t^}��*�8tP��
ܟ�	ӟ��~y�xӠ`b���<ٛwH�|��͍�!t<���/,!	��â>�����'Ƹ��Э�%1T��u�҂�رy�O`��v��,M-&�K��1��\��?a���O�s�ٱ3���:�C%(�0�ӡ�O����O���Oܢ}����(�	��KF��(p�m!p��t��v�П�'A�7�=�i�]2CA�O�ȹ[�*�?>R�c�c����۟���9C��o}~�ϟ�����9&�t	Q���X��padM̬'�'��i>M��ΟL������I;^u�GF>Y_���kX�x0�'�<7m�%}²�d�O��$>�	�O@	cd)�5OvH�r#B�@�Δ8m�v}B�'��O1��\�MS'>̰r��5s !0�݉��UY��<	���4q%��	������U�M�HxR��++�peS^Q>�d�O��d�O�4�"ʓS*��� (��Y�B2�A!��?xx�*R��; 0�E�����Op���Op��	 �ЈY����K�lu���^?>d�$KbӒ�2f�ҁ蟂�>5ӣوd���ID�ˬ9�rY:�[DJ�����NP�|�����Y�P�'ӂp���ŧ̢%��z��Ol�i����6񹳀�q%���(�=I��:iԒ >`������Ny�(�1�d�Y�ؿ!�1ؖǒ���<�3�S�#��-�3��E�ފPYFh���˔C쮭yŊļ(�4i�� <�ʤ�G=U��x�~�� ��B�B�P��\�Q؆�K&n
�ul�%�@3I/�E�E웺j����ug�:t� 9�pi�6�.M��� /�P�D�i#��'�bHO�*_�ꓶ���O��	`F�b�E��Y�4c��!�c� ��G�I����	̟Q�8� +��{9�P���MK�ԤRT_�x�'���|Zc�5�d 2I�`�dJ�O�ֹ/O�0�R�'$�Iߟ���埔�'�����T�KS8-P�`E��]�I�N득��O�O�$�O�T0�a�
SR"��s�G�0�|a"m���O���O���<1��N�A���dx���E�k���A.�8?Ǜ�\����G�͟���9"����I+<o���ADSq~�ؒD��h.Ź�OZ���O\��<)B��hX�ݟ�gOԒ/�YɧÎ�,E��'�
�MS�����?Y�`h<�����I�t
�t���:@3����4<7�O�D�<��:qJ��͟��	�?�H�@�Ot�q^�N�(r�RG�&�����8��m[�����&BZ�e�b���n�fy"K���6��O>�d�OT���V}Zc*l��̰p�*@��ƭn]\b�4�?��RR���2�I�
^��8��f`�q"���F��G�&7m�OJ�d�O��d}R�4�Ci@x9�K'N�(r-ó�M���Z���'�����0���O�*+m�ٰ�3�X|o����I�� �q9��d�<	���~��5'�ba�d�4ˠl4MS���'�&X؄�|"�'��'ל)�Q�I]h��FB�� 3"w�����5P��M�'$�	��<'����B�يv��p!$M/&�`���>�V���?	��?a/O�et�ە`���뵍�5�H��3��k�hP%���	��$����u!ڜ�^A �EʺrZ���!��M������O8���Oxʓ'��@[7�H	� ��L�zYHƋΘ?�A�@V�l�I� $�h����'� 9p�/,�����	�/}Ԝ�3O�>Y��?����$�[��&>U���ӟA���'��X1�)��M������4���d/��hӵF�e��E#ab�z�aΏ�M{�����On�`�ɺ|���?�����A}�"0AVǕ+h�<IxB�����|�'�P����0�G�RS�(1:2��:"�ybF^���ɓ����	����	��\yZw�V������a�10��Y�{��H��4�?9(O<!P�)�Ɍ�9N���M��i��흈z�G��'���'3��Y��'9@��l��<�D��D	ޢ-���Y�^�2��3�S�O�ժu�<wL���в}2�$c�-z�N���O�D��gM��S���>94��	d��|;d�_�%:�jA���቉��O�B�O��c��<	4� �Jf�q`�,��v�'Z@p"\���6⟴q`��KD"I�"�@0�b͝<�ē+��|�<�����d�O��Re���|	�҂�G0�����)V���?����'ZR�O��*����jN3F�N0;$�i���Y�O���O��d�<����M�|j��Lw^A�a*��.j ;��Yd}��'`r�'��I럄�O�BDFA8d*�k�
�����oT�fI��?�����On�iPA�|���!���^��-Yhԫh�J��#�iq�O���<���T�I;z��H 툡jJҐ:5�ùJ��6��O�d�<��!�IY�O"r��5�(�>I��@B��W'&�p�( Gր�����O��d7�9O��P�T�@�&╲bl�p�MCJ��&S��1��M3��?����]�֝G;�A�%Hu?��e[��Z7M�O���x��3��'��Xs�KS���\��3eB��Wa\6M�+Yh�Qo�ß��	؟������Ĥ<Y2��%�E�Z���H��66D0ڴ	�R�̓�?�.O��?���
H��aI�φ�.�&��-˓`ע���4�?���y҇4&<��ey��'_��鎬J�iL,i������G�^֛�R�4	"�c��?�����$Bd�"�棟�8�&�H���#�M������ W��'L�P��i�U��G^�I]ڸP�D�xH��>��-�w~��'G2�'U�W���Á�DdƜ8tmU�T�z,*��B�Ko�S�O���?�/O��D�Ob���t����0�,q�D����:�=Op��?���?�-OJB �|2���7yP��"�B��,��w���5�'uRP�0�I���ɔ���I�o��kP�Q@x�f��.<'9�4�?A���?���$�# !lp�ONRl��bJ���e��<�Q�J��7m�O���?���?��H��<�H�x�D��/wk�b��T�H��H{�����O�˓=�Tb�]?E����L��n��A@�4h�|�4�|��|�O����Oj�ĕl��D�O��$�O8����$��j� ��1��6M�<��K�]͛��'��'��$Ĺ>��wG�l�1�ܭ �LS6�M39;��oҟ��I#D����!��m�v`��I�t�j�� V�^��7m̅&�V=m�������,������<Q�C�0.-(����Y~���U��6-T4=��Ob˓��O�B�C�/NDѳ1+�#y����.D��6��Ov���Of,j��Q}2[�H��B?�A
�(8{�|��J��-��ǀ��'�D�y2�'G��'D�@�+z
����f�3YH�!3tB`�r�Dy�&��'/��� �'.Z� ��(�/C0f��<��g��G��t	2^�|��e�0�	Пp�I⟌�Icy�&�7]I�C!�)dh�4q`	�O�)��>+O\�D�<	���?y���[����h<���Ƽ(p�Ac+��<�.O����O��d�<��e
@��J)#�1��K�N��c�%���T����Wy��'g��'�.y��'H8�c�f7v���d�k�:!�`�r�����O��D�O�ʓ;�t�I����5�C]|�* cu�ƚ
Y��C��M#�����O����O�0OR�'����rM
^�^�!@�i1���4�?����N%m^�@�O}R�'���k��ZJ�J�	�?��m����VNd��?����?��x�T]�4�����ʖO�&YQ��ug܎{;,dn�py���;;:p6��O��d�O��I�N}Zw�P��A��e�*� ��ː��۴�?Y��%���:~�s��}�L91�F�ȡ�ЁS^q��(������M���?����R���'\ʥ���=O|��Xc�c�tA�Ĳ.�PpB)|����ty����O������u�٢D�i���c����)�	����	H*N��O�˓�?)�'�E����EDNH�S�V�ߴ�?�(Oj	j�<O�������@��VI�Xs`�|7M+�!���M��AG�(��_�X�'�R^�\�i�պլ�7^��Ի6Â�`j5�*�>1r
S�<���?����?����@&3Ft8��J��)5�Ľ�P�qDXS}�]���Ity��'$��'tR4h�I��]�*��Ca�0+s�\���.�yR\����џp�	qybg!Q�x��R����N�?��E�'M�89DT6ͣ<i������O����O��b�S��z��L�l����-V��+�DӐ���O6�D�O��ch��f\?�I2�Tm9�-�XWH]�UB�"m?t$r�4�?+O��Ov���;d���b?Òt��X��*F�)Z✢P������	؟��'�����'�~���y�'CJ���7�V�N�'Oߐti�]!F]�`�	����I>l>�G��'��I��F�TY	i�*,�����՛�X��PD��M���?Q���2�U��].?�0��6"ҷ"*�A1�AK4`k>6��OD���v\�-�$%�Ӗa��ѐ�mΐ-��s0��Z6�U�3s(�m� ���<����d�<q-AI�(Y��f�6�<5��BA�b�v�F��y��'2�'����ּHp�p��_]��
ɧ �0Xlٟ��	󟀛E%�����<	����d�1!�neR�LF &�u�Y
�M����� l��?��	�4��1!�p��s�T�f������9%R�rߴ�?�N�d ��ky��'������'2�� R�T��U�c��6Ύ�d).�Γ�?y���?Y���?�)O>���m�5d_.��$�;L2 �1�@�܆P�'��	ٟ@�'��'eB�¡ǅ�PJHI�2�*u�ƴc�F�=�y��'���'urQ>�ɓ'� ��O�j5�B
ѡ X$�DݱZ;�`�ڴ���O���?1���?�i��<	eL�6�
i:%�aE�,3���}A���'���'p�_���#�
��i�Ok��Z|ƙYW#̞/تi�A�T� T�F�'���ϟ �I���X��i��Od�8d�ߞC}"�HF,�=|���i�"�'��ɣ;�D�)����d�ON�钡ek��*Ԋـ*B�YK㩜#���'���'�!���y�\>��z� ���$�J�!A�(�Vـ�kGǦ5�'���ĥf�����OH���H�ԧu'�_���*.��.��F,�M���?Au��<�EP?�IB�'tj8Z� ���j�Ar�Dg�:Imڕy@pj۴�?9��?y�'2n�O8�Խ��դpN�H���H�	�.O�"�|����O`tI�
��2Lk�h�v�j��d	PѦY�	Ɵ\�I#
�.�1J<���?I�'p$���S Hkt�`�O� ּ��4��hvP�S���'���'��"���6��&l�3f�EQF�`�����t@%� �	՟�$�֘�z�j�{��Á6�|��wO�5i��<�� ���d�OF���O��[HP�b/Y�<46-2W�C�]'B=�Fc�T��'���'��'���'Z��4
�z���_}$��Q�I�c��X������`�IcyR�͹��SV��&�[=����mޘ2�z��?������?���^8`�)�[H�s*��r�^MҲ�ӎ	4؜�S����؟P�ILy��9I��윊B�
;9پE�G@�O�8@��˦���s�I̟��	�	���G�̢BB[�#j�TpрB:Qy���'�bT��#0&���'�?9�'��Y�tBЏ���B�]�$�x��1��O�Dд-o�?�$�?� R'~pza�&�֜�,���eӆʓ�pXP��i�X�'�?9�'y�Iq��)j�+B�Z+6�!��C
(�J6M�O~�$�51����}b�)G�C'���E �|���æ=��΄4�M����?����RQ��Gf����ƌ�F��8�WR���o0�j�	Y�w�'�?�D���2L��F֤{�lH �nݦa9�V�'�b�'�Z	ҴC'�I䟨�>��ps3A����ea���"*ݪ!lZ_�I�7!�QCH|"��?���<��X��	P�x�STR�'6F1���iB/S�wr�b�D��X�i�����2X$Ha��
Z�d�� �>�V���<�-O0�d�O��$�<q%K�+�Z�"VM'+��3�[�B+��p��x2�'��|"�'�B��]�j]��N+1��y�(�o;���'3�	��	�Ȕ'd��6�a>��Q�+q(��I�$� ��>���?�I>����?���Ŵ�?q� �t���=n��� ňO]�	BQ�����X�	Py"��2}�& s�n�4Z�`���Q>n�@��d�ئ��IH�	��ɾ5�8�	i�D�f ��6�ێ��F��?1p��'��P���aL���'�?)�'n ��YCJZBͣ!�%�ݑ�xR�'K�@�(i�O&���VY�D��'2h�Z��D�6 ��6�<��f�0x��fͨ~����B ��0�1h_���ٹqy@��Ḡ~6M�OJ�$P>n��D!�/�Ӈ ��Jk�L�y��J�T	N6�I�bh����O��d�O��<�O�Ƙ������B�=N�����>�"H�y���O⬎���(�8PAE�%J�6��O�D�O����B�[�	Ɵ���h?���N"X�	��W�t�v�:��Z؞���ޟ��ɝD���D��H� ᘔ�f�m��4�?�v�S `��On�:���8��L'�N�����#���Hd�Iɟ���ٟ�'(Z�qկ��jh2U�m��h9��,�W�Oh�D�O,�Oj�d�O��Rp��L�����Ị}�,��c�1O���O�˓�?)f"Z��k&#�,u[pd@n��TCc��M���?�������$���B�iu���@/y�\�ѶC��F�
-ڮO�1b'E(!���'�"}�%؋pi@ꐯa~�š��s�<Ʉ��L��� ��o�X!ae�r}b��)=�Dq8ӆ�-n�YB�M��pRP�2��9y��#$�.��S�	��?���c��=�P�r��:O���`�#L���8P��5mP}�7���Ta"t�	�����,cר)�S���!��hi��߽^�6�R��56!`4�N�	J���&��k.N�l�����$�O��d�;u���r�D.�� �MV�?WD�Z���ON�OF�g�'�}��>9�c�9��HB �E*�� �>Tz�;�?O?��F8T�4��%�.Cze�U�mElL��d�O�h��ʌ��'��`K�LUt}��D�v��0��'���8�sUvUjBNˤ\B,Iуĸi�<�Gxu�Xm�S�O0�$��47/��G�1i�H��'6��/s�b����'7"�'�Ga�u��ɟ�C��p�Ħޣ��A�aJ���?9�߅v��{ҊT�+���3ړ_� �W��H��Ò�Z�$f	�F�'�T��W�Ǹ����S��jF{�C�&S"�@7�܄<WW��~b���?q��hO�ʓO�=-$�5���N1����B C<q�m���d�
(/}������c�2(q�i>q��Qyr-��p6�	(�qV�����3K"J���O���O�����O���p>�JAl�D����T���Ӡ=�v-y�邾2�:<*6M`x�l ��O���+��Js: �e,@�^�h��i�d�Ptf�ٟ@R�Y<Q�y��O ��G<���ʰ��T���#���=q���/�5*��zdqC0bJ%|�ax���P�z����1ӼP�e�. +
�I��M����ٱ~8��O�"Y>q����=�L*TĉD��!Ҡ!s��m����	&%u:�Ht�Y����[GP��'_	@�s���9~��l��E���Ey��D�kf� ����Nr��>�H�h�ESL�ѡG��&{M��.*�Z�X���D�JA+�(Qy���rJ�!uy����^�<!��VN깠��T�
��hs'MVC�f��I��ēbH��e�S�Np�P3�%� !����	py��i��'��S+A��)��՟��I
U%l%�U�W(8�u����/���HG�����<��O sA�¿`Azu��eȝX�(��B�'�"<E��I�p��6oH�T)���e�4I���?������O">��ֵ�$s1�ڱW<\t�Ps>��O����K�!j��rb\#,����\*�hp��4���$�x�p�#�AB`&�9���#X���Ox$�A@�#!o,���O����O�=���?y��E�H��Q ^�"����v���2)�!�څ����]�)�֋';���)�b'_���$ix����K�iz�����9��p	��/T���őo�R�'��YPbT=}��d�e�L�/v���'ژ��bֆ@F�T"�=/?hycO2��|rI>�0��3e���د&K@M�EN1:ȝI�O��'���'G�!S��'2�'	P!8���2��5�۪�D�X͜�2#���������*A�az��i���LػK4�y�����9 ×:��qR�O16�lU 0��DyR
O��?��Q�.��f�:vn�`�S�ܱ�b�@��i�^����R�S�m�;��y���[�q� �eK��-��c�O�̝��Ϙ&
�l���iI�Y%^Xә'���ev�*� �])������O"�'6�F��G,�$n��U�č�/�D]��F��?����?�aOS���4�|*��%I�pc��]!�=ô�:�(O�
�O(	&4#}JEb�I��֎�%�X�q�A�'%�����?9��?�)���5-"IC�`���Q�B��b���O>�"~�S�? �!K�ŀ%�mr�(ҋ&�~3C�'n�O@�����f���)��2$�
���{x��0b�%1!���gG��6l���.D��Af���8���� 5~�\�!9D�L;pCќ8F�1Ԉ#m��z��<D�@!R`��]Ϟ��W��A�!�=D����� '���I5"�0(��h�*O>�fKV�8��I�V�"F�@��"O��At�L~퀸{�:A�y�%"O��C�	4D��h?����a"On!B�*�6��r%2_�<��"O^̓�
_7\(+�㖅T� ��"ON\k`� 8~�q��|�n�"�"O��?6I�4���M����E"OΩy�]P�y���j�e+�"O����)��c�:����$�< "OHM3Ň�t`����# ����!"O�M�D,Ǫ68��#䃟u�x��"OD�a�M�K6	�M�(_�T�&"O��H��X�l��9��,޽QC�� �"Oؔ`E	�M���1�!DC*0��C"O��`�V�zeT5D�͆T"9ID"Oάz�N�Wm��XjЫeR`���"O� 3 �ڂp��̂�I=r���"OL{Q
������'�]q�(Cr"O,���F�Q���u��5U6�K3"O*]S�F ��`@0� fmr )�"O����0E���$�ۀM^h���"Ozu��=��$h�3ESZ��"O����ϙk	�S�G�EGF}�"O^1�D�/����׆�#1�՘�"O�RV+]�l�LXb�/i���cs"O�K�K��V|�Qb!�s��<ñ"O^M�Cƅ�=��X��bȳ��`� "O}�#C+4$
��r��K��T"O�h��*�D^}�#�]���Hk�剶ƖH���N��Xq�t�Kb���#�ʑ�6Z!�Dʁ3}b�/(&��}��	��rY�<��c�%b�qO?��=n��̐�BY=%y��0�A!����ӈϞmf��rq�̥R��ĕ�Bt�Ls�@�T��-�u8�eY#K�}�����I�(��y��6O�@��F��b�Ƒ���J/u4�#"O\Dʡ!٬9��) �Q1��2�,KLd�!��"x�p�N�
�x$꓂èk�B�	�r�|h#F(<R5bd�@B�PID�hgʆ4f�r�"~�I��TJ�iy�Dh�@\�W��C�ɠ�3Ў �^cB�J� ۡ>1�OR����7��.%���[�l�)�!�DA�c[L�S�Cz@���~!�JѤ�t�?o_���H�>|!�D�Gp�a�̏<�z5�1��M�!��E-kV�B�ÕG�~CU�S�x�!���bc(���Cf�
��DhG
'�!�W ����Q��l���ǃ�k|!�Q�p���z6O��~X��C��3Ia!�$�(d���v��f�p�e��[!�ͮE�ֹ�^�4P�@c�ɞ T!�d� Ʀ��f�+C�ba�!��mm��
(�P�c��/>�!�T1���ZT�Fu �*5�!�ZP������b�ػ��W��č5�5��ɘWݦ ���V6��9�gZ�A�D��$S�m9�S�'��� ��%�7C�OZJYQ�'	tmc��Y�o��i�uN�/5E2u���$R�=dM#��� |
���kR�4�"m޾'v��"OLh�!G��ִ�a+A�{�0|H�Ą�zı���Oܑ���O1��'����D�
t%�}�U�1����	�'���
E�U���$�*R�z$q "���<7͑�9��`��8����2V���2�W�X��	5e���t�i[n����<I5C	d}PBʔ�d4��p��a�<�&H�+_ҥɃ@�*#�����'�_~����B��is�݉�H�i�OVly�!��G��1�n�8|T��'\p����^6f��4�G��<O*��F�A�E#�'�$����ҁ��Ϙ'��� �:<�n� �/Vp�� �'j� 1dӼPf�A�fK�^�L�+���%y�6��	
i���t.�k�OD���LR�w`���IP�`y f�DV$[n����M5k��%9!�{��k�Y�~��G�T��G	�>�aPNR����2F�&@�{Zw�lJ�>9Fh@�;�2H�`��0��!(�G�c�'e��'�4I���@�2��S:�=��� 5��E	�0W��E����OX x
T+�(^� ,2Z�ֽ��i��h��P�#�,%� U4�BB,��B�N��bTMC$  �b��@���3��B�^�8�2�f/x��i� CXp5����<�~�<O��@�0fC7�FJ1Ob�mM*�f!����
@�A�.V Q[֥ El�L?���|B��6裂hs(��O9h��D�8L��esre�RO2踒�^�_����0�*�kY�]����3G�Z��qᑢt�
�b�5P;Z%��j��Z��Z�(HeA�@�v] ��� g��Y1�LX��N�/(c����.,+��=iN�S��Q��8DG�� ��?) b��zys���J�r��V'�"b���^� ��F4e�l����'�ܙ�SJ.P^�E�;A��� �%�7�2�c��C�,M� ��|!4"�f.�8`������Yd��"P��e��ɢ"�';I�q�@�D?"%��[d>OBx����l��� T� �%&�Ƞ�|R�L�W�&5�e.��$��1�	�(u�U{�fB�_f�K�c��䓟�O�*�٦�-��8gm�9R�&�0��zh��g���� �e�*�hO��Gf�>�2Ұ��m9����+�T����|�#0E"T�±U�h��`�=� )�N^?!�G�)K`���Mͨ'I`��+A�hO�Z��٫���ϒ�ʑ#Fb�ӭ��Z螁�r�(f�,ҕ�{]jy�'`�@0�c��\�X��P�O�� �
�9t��6�D�qA��r��#Ñ�z�t�;O�:� |�����Y1=D�sN?�O�����İ3k�����;Hlna����OO��'o ���IG�Wt�<:5��:E��y���V�p@*�(�L/~my�C�#"��!kw�����Տm/�'�"|r�M-?N�\��<4]��
K(X����`�Z0�G� �.���1Et C�Ȋmɳ��3\	X�b�X�< �R6vLp$bU�B�'Ԫ�KQB�z�q�UF�.(�lQ��I�8�J�"�JO:��Jԝ~A��,b����l�� �T����QX�D~b�ť$#��D�����]�3���K�,�+4A��(O���	�dIB`��J4,Q���`�.�<���\p�T�) Bē6J&��j)#��\�I�L@����d���*w�@�z�N9�	H$rD�vD�-K�r�y�mW��"0�@�OlX �ރ��$W�-�ʧ��d	44���qㅽ���򉕏E��AA��M<7�^�4�',|-�;=�6����1<����؃B��.O�@���
#�
PJ �+�n6�aA@=.��s�K�lI�� ���O,	���3?��}�%����S��p�@���r�� _��Ժ�'�Ӻ�Z`����HA>D�;k��D-�*��%�nvB�06C��<	w�	�.��b/-#��|�|�'_��H��m���{S<��ၩ�:+O�dϻ2��/��X{� �vў��#�HQ�L���I#sgB}�O���dJ�'��9꫟!V�W4��)$?�v(H�qa`,p@,�6:��ф��.��6\Oz5�$�w�b�K�H��'�Y!�m�?\l��hf,��td9[t
�5R[���NL�&F���T>�������~��*Q� hU`�"��"�����(�R�iQ�V�ʰ�`S	4�01;��ŉ�Z��I�6�B� �3*^�ΧIr�<���X?x��!�c�${���1���<�S�2]����';+��5��*(��AE�ގu�"�� �Lx�BZR+����Z'��N����۠LYi����D� ��S�s��	.U	��i��x�2 C6�}�O�<�O�~Љ4'���	���F����A��\��^���2�b%*�-[1��К�C����dK�n��̣�{��~�Ar�����:F7,�����nxa��T+�XKtp���Q$�&!0)N��'"& r�!_���'�"ċ�O�� [h}����!e�<�4�Ս�y��އ(.�V��s���G��u����>3T���ƩS	�}��^�|x���/#�g?)1�K�ZB�%��a��p���v~2CZ�CBp�h[O?�1(�?�@)�ٱnA�P�"1H���O�=��7LO%bgZ�d@�1�b�5�(��F�������~BH��vr\q�=�S}&(4�'����w��y����B�,9>�H�����50s���$ǆqۈt%>� �T�H8]-
5�E��{�\0e��;��}r��$ұK&�	�/<��ff@64s����!�1xb��C�.�eA7��*K���#���^�1���'dԾE��i�>W��9+��<S(��dCl&xP�FFK
g��Z7�ٜY#6��b�%/�O�^��!c`ͼ'�f��;u�"��ɀ6�PW�ڀ�~���I�?L���~�#C#��lc���+�dʓ����k@d���Ar�R@�4��F��7t�)��P�A*l����,@HZG|��t����)X�-�ڝ� Y��y()r*X eg��MI0e!1d�"�P�&��%�iڐC6R��a(��l��6��-��xAI"#"��*�J��f�\�WĐ%0)�]Nl�D|bN�i\����C��~F�
�	ġXf�y���'ɐ��䚇s�	b$��?�~=�Y�Ȯx�ӓ;?�ͻS���qU��M�����1,�p���V�8��� /��5�en�?(8���	��PT"#?!��3c��C�!T��~��a���]�e�h4��P��Q�<@�@ �K=��a����
��1b�'h�	Γ5Ă��Qo�C��|�e��)7���'�����!�n1i��H�>��!��D�(Ѳ��-��"]���g��y��lː�E�n����7볟�=�	.5��E�R�J����m�\EQ�4j�@�p���[���Ę�'$]rNT�j�P0��t5���tJ�7`D�H�>��w�8�3�% �-6lC�����hp�'J8�1U��{L�T���F�UՐ}c����O��a��B%u�z����8k�!)Ŀi6���E�:�
IP�_�:@�	�o
��"R@��0}2�t�-Gh�"���q���03An�$��m��)���*s�E�2F�]��&�Й1*����T"L�
Fj�g�'>�,��4�??)�`ߎ��X�a�{J�KS��H�'Y`]�1��#\a+r)�4F`dQ��\����K
=X t�q�p�*�ʟN(.[�-�>l���:W�<E{RصP]�w���m/��D�a#N�i쨬;
�'x`�WM^.����L�(�J!�-O�!J�q��(�@� ^X�T���ɏ\���X4m���N���#ERt��DS'5�HpY䉁i:~�аl*U[Y
���_��xYG��B��P�큅 �~����uQ�PN��0�t@�@Kxc� 
D�5 �x�R��Ae�����	C�(ja$���TӿD!�Y�<k�t�KWR��Ă��8���˷._a<tt#1�Z�`ي��3?��-M4���8@$R��0�-D�<� ���p�B�M
�)HC6j
<�,C�p���EI��%	U8�0`�B?<sl�`D������:\OP��V=+���*q�|	U`��ܩ��g_t]���1$�闧�6Pdhԛ�j�L��mҴ�:D��r%o����C��/e�2��3�:D�����[.�ve+5EˌA���j=D��A��6V�ȣ��Md�M(SO;D�l�f�Bo�B-#E6 �B�:D������(,I#"��L�p4��8D�8�w�?2��u�J4%�2�&�#D�YGO�z'� m	-`
.�[��%D��i.��M� �D/H'7���0Ċ#D��i�fȿ?z��*b�
4���K#D���Pe�: ��p�TA� U�e��i"D��P��ͨw �� �
C�
��E �?D�xK��I%s��<	`e�+S28)�w�!D��;Т҃�6�aT�1=�f}��3D��sk��km����۲�h$(1D�p�F�¡=.��E�i!B�;�!/D���ď-�	�p5�|�*1e-D��h��W�~X+��,4@H%�)D� rd��=���,�
a�@g'D�D	0��P���I�$�8��`�$D��Z�l��J�^<��F݀@U:�L'D���6�=sJ��v���,�@T`�d"D��@�oGim�3d��{�*i2�2D��g�=g�TP#�Ҩ5�^9I��=D��2��^�3t�4c��B��0�Y��=D�X�a��:���a�D�9�&b?D�(���""�f`{2�� ;t� >D�D�q���n�0���*�~	��/D�� \���b��!:pou�@mɆ"O�ŋB��=Z�̂5��H��"ONݠ�"�1.�ఐ��I�{��a�"O�ɱ�_�@��A8��� e�2"O�T2�W9��:uU�
��"Oĭ�����Ġ\".j%N��yr���a�r1Hp�#ð�8�$5�!�d�-8<��fE��%x��hE�9�!��R�& �Ң�����X�![�A�!��дPX�r
�[NB9��S�$!���x���u2��ӆo��	!�Dο/A`Hr�J�0{\U�#O�� �!�$l 2�C�-*W�rqHC-���!��V&.@J͋������jW!�$��H@ �ړ'<�B�+D!��zް�RSe�B	�<B��	~S!�D�7j�y��)Kdu�բ��.g!��܀h��呱b�2(Yư����;�!��̘["��kE/�*M= �̈́�o�!�$�2T��
��Ϟe;¨�`�ѻQ�!��
b��]�F(�,�[K�V�!򄔻q�R�ɅN�e�(��!�<P�!�d��j�>}��	@�/D^��`��v�!�D� \�YF��[P`]�Go�6�!�䎰�i�H&d������& �!�dA�+f@!-�Wn���֤΀b�!�
�$�f�Z��P���%¢c1V�!�� +r��.M 21���ғ�!�[�,:��%�B-�Ȱ�DKơ0�!򄉢~�\`���}�ɒK�+-!��׆~y�Ua��'p� )��Iж0!�$�+S��e8g�O�+r�%ɂI�"=#!��ٱ����wg�oU�cб:~!��W��A��Ϫh۔�`��ձ,n!�D�0Ġ|(c��#6�������!��O�,���z����$��ň
L!򤑖@%�8�ďԤ͊e���4!�$]"�V%��oͣd0���7(!�8�V���Ƈ�|�Ԉ	�ˀ%!�3;�R4!���x�d���nBx!�O������@���U��˸_!�dǼ6��Y�v�R��,x�#R#�!��9�j�Sq�س1�ĥ���(o !�5y�|����-�2�0���8!��6$�`}�`�B�9�P�홢�!�� 6�*����,PD�Pk��UX!�DI/j�s"�a� b��U=-!���Ĺ3Ig�`��`�ڿ_!�$@,��0JR���HX���ʅA!�DR�ʤ���mJ�]<����V&�!�D@�2���2MX�p'���6#CIx!�M�o�0HS֏�m�\�� �� x!��n�����	&�İP�f[.Ci!�I�Q�b���O��V���͜J]!��Z�|�Bt��XI<TQU�Y9>!�dە����ֈ6�JX�%� &=!�$_"_;\ ����>P��t� �^�	0!�䕶V�rՊ0�J���O4@�!�$
/�� ���u��c"$gU!��[+Uń��'��=V��!1W0)D!��AJ�����'5�����-i9!�dF>3�0��� �P"5UN�y!�dB�%�D�(�J�m{0\�rk�W!��&|�x ��Qs������ !�� �`ĺc�*���,C���X�"Oĸ�'֠Bs�ID�Յ5���1b"Op�0c��{��y��۝��m@p"Ol�Tc�> �j�'h0�8�"O�K�cR2�c"f�{�>���"O�k���9~b�����3"��ȁ�"O��R#חkz��0�.�4`�Ʃ�"O8@���D�a��Pu��� R"O��8T�2� ����	�u�����"OhT�p�	�NCFU25I����u"OF� 6㏺of����J�j"$�s"O�m��E�(��X�1��t�rSsO@�䁇n�P�2�� %X<�{���x6!�_�E�Hȋ��ؐs� wj�b�!�dE SF@�����-�&<�3�>?Z!�d�
;
Xt��G�� ��X����2e!��+p�\2���az��0�\%9�!��I4��c�.��j��3�C�P�!�� [BU�&��L��ɓe��d�!�$�%g��}1�MV�z��h�%+� 	�!���*��C; �t����M�!���U鸄�ņ�F��$Hq@:y�!�$ s?l�9�g��D�L)�B�M$;�!��^�~X&h�J�3lm����A޽O2!�$FHL5���N�4?,��w1!�	��j�҉P�Q~�#!��[O!�U&}pF�S���0r��F>!�Ĉ�|Y�1�����o_;�<X�ȓp�0 �c$N�g�`mPu`�Y�tY�ȓ%D��q"UCx�a�KE
�U�ȓD�E�tI��ڀO6��$��oɐ&ǌp�P"č N@I��x��<���53/r�(Ç���轇�	Q�'y�MP��Li� �0��D�$��'��q˔?��ؚT"M�O��ȓ_f�z6��76�B ���+K��Ņ�\:�r�J�4:�qh#AL--��X��I˟$�dQ,?g���S��]%,��VO�<Ԭ��h�>D`��/���B���G8��FzRAׅX�<C�Q�����y"�ۢ����K��_��8S���y2��3+N���GH(m�@iYb�3�yR��0*R��%�_�s�XL�L���yB`�R,yi��(>��1���<�y2HZ�NB�L�l\�4tn ��L���ykK�A�Ƙ# Β1��0NԐ�y�b��n�Y�ծM"#��i�$��yb	��k>4�H��	�P��3�(��y�h,t�\y�X�zr����#D<�y2߇D����,p�z�1����yL��06q��k�^榸!����y�������S��R�!3b��yb+��x��X�m�D�
��C�B7�y�h�D��h3�G��f����рK�y¨�q����ō�*Y�aSaI���y�ŋ���h�ˊ<A���B���y2`�-,�"�A�8�Pl �&��y"��/wh@�CR!A*m (�Ԩ��yI�aLy���.A���Eܷ�y�
�4'���v&=�"�OV��yB�J�9d�m�D�F}VJ]�#A���y���0Y��q��nڈ	3��=�yb�7i]��[���1l)j���_��y�kC>Mz�X3cTc�xPa�?�y
� �%X�԰j�n�i�A�'����"OĈ�V�K�o���r�ʐZ�j���"O��!����Z"^,�ƥ�;���q�"O���$�[5fE(��&��"�"Oh񠔦҉h��ӰL�q�B���"OZ�"��4����_���V"O�A��1T>�:���jb�ѱ"O��y2@	�C�	r1GO� �,|��"OLd�f�L'$��[c��u�8��A"O�L{6%E�ar��+�)�+ێx�"O -d(�h9�`kŧ�����B"O�<b�
�*Bx�&-ܩN�z�x!"O�{eoC�$#���*ZV�L0�"O��ۅ���T�0�9�,N%W.��"O�1(R��J�)�b)��.h`eq"O"���!F�he���+kv@<��"OR�Q��I�U���=sgv]��"O����ʇ0���R�F]`X,@�"O<���@J��x�ÕVQyP"O"t���~�bЈ%�[9t8�"O8�vϗ5���Ґ�N�]�"O ��$Ǜ&J��ѧ�-6����g"O���m̹��hH�hM!,��"OYK��B���QI��L�%�s"O���N�Hߐ�R(ǽ;���p�'��'d\��eŪ.��X�U�
p�H��'�T�	F�?��,!��#}�t���'h:�K#���p۾�FG�s� [�'S���F����gVe�\�M<�����K-,&ؔڶ&�XN��#MR=P!�@�CP�h9�`�m���`��
4�!�D�����$MR�?����
�o!�$�/>����Ȁ��5�O*3	!��2d�b1�bC;?h(<�5�ʞ(�!�D܀>7<�r&�Yr�q�A�/
�!�$�"@��� ��i`����O�p�!��=>�U��
�!>A0�3�oR9@�!��
16^�`%F�<;l�cP� o���)�O$(
��[:B6����2U(F�c�"O��UR�4y灈&�$9�"OB�����;J�`
c��W!��"Oޱk�H5?l�Ip#�yb�f"Ofy�&J�f���"g!��=�HL	�"O�e{%��%��,*v l�z���"Oq��G�0q�,���1��t�"OB�K����]��(Aǅ#&����"OL�u@�sش��}��2B"O2���D�
��)�v��TxD�q"O������
>��7j`���#"O 钀��}�:�%Cc.�9Q"O��#�b�	����2C^��;c"O�A8�O[92��4�qb�Zd"O�$QF�O�j(�`��\Hy`"O�� ���(>��u��؞FB�"O�D��%�I@��p�� 3�%�B"O~�j�";��$ ��e�*r"Ov�����U�M�c�C�#� �Pg"Orݲ�>V��A�O)�p� �"Ob	�E��=D��۵-�	����F"O��wI�-��#t��+<Dtڣ"O��)c-��}�,A��.^+h�� �"O$U ��[1��KTo�2^8�v"ORP"��P�{2�pv�ճH�0�r�"O��k�$(�)����0X�"O� �q���Ք�D��� .���s�"O>4���Y�h[���D!I��"O8�$2z�`���i�=�C"O���CL�u�
�
.%3"O~��#�˶E�̅��������"OX���`�X9$�ȴ��;Y ��"O���ץ�F.p�d�ȣ���"OL��+V�s �	I��L{n��"O=Q4@��|����k��Ap�t�U"O`|@r
Lޚ�3K ���u B"O|e2���
?��er�����p8�'ŰQ��8<��+(�ȹ`Oh�<�e�}�:1S���j5L��d�<1R����q����>��P�%�F�<ɡ�L	~R�p�N�L����#RE�<q�iJ�-0��V#�<,0J	� �l�<�Q�_�T`�Y�R��h	f)]�<�FP�;�D9��	�pv�qW�<v�ŎH�}���A���K���K�<і� '\��![�O��5[��JI�<!� Ӟ:�Jy�f�	w6P���ZG�<)D�W�E��H�F����ٵjG�<�K\(���K ��=J�,�	��F�<ƋX"{�u;R��8L����X�<cX>@�rYP��kX}z�m�W�<�QL�@���x���p����@�Q�<���H����z�VA�
�ymIQ�<!�M�*�z0��!�F�|�YC	�r�<�u-�9�J�yc�߯WJ;�U�<a�LYYx> ��aO,b0Ĉb�C�j�<a�O�3|T6��FS���u��e�<�g/R�$�S�[S ����[�<��EG� �r���S;��|���[�<���g�vIKeQ!h�P\��o�<���R�/�ژ�F��g�<٢n�i�<y6a�Z백+A�̐i|(�&GM�<�'ǋ�|�����ǎ�����p�<�ҏҜX�LY�F���f`�ƺm�<х�E�H!�Y0c\;>�pH��o�<i�c�A%�sv
Ze�����l�<IA O�Ld<�Q󢒊,�� �Dl�<	V�5a�@�[�'uL`X��\|�<�'�z��40�kT�Z����!�x�<��O6L\̚�ǽ=�H�D/Ku�<Q�`�3lo(Ԩ�����8���p�<��
��9�����6w6Ѱ��h�<��%\�-�z�/0g��G�I�<���@�@3�ҁMȣv���)�k�<E�٬3v��BT� �z]�� �k�<�5��1+Ԫh����d�j@XU.r�<i'�J9p�t=8�OZ�5�`lP��j�<����N@��T}D$�R �d�<9��K�8����]�`��$��]�<�ǌ�Y��T�B
�����V�<yg�U;���ҤN��{�NYq�S�<ٓnӠ6O*�{�C+�ʄ�1AM�<�����P:� H�m�a��DM�<�e���lDY�7$��;8Q�KL�<QU"I}� �%j�-"��I�u�I�<�$cb��L(d$W)Cm����E�<	�jO\�
m��.C&a���4A�<12��S���ĩ��y$����˞|�<��� �r�X��ȿ{��MʒfGz�<�F&�=�&�k0��R����D�u�<� xU{�ß�;��4�&ی{�c�"O.�C��AH��p[$�/]>�Es"O�T��%(�����͍>�f���"O���Fj�������H����"OT})n��
⺁96�m ��2s"O��Z�MEM�]2&�� !��"O���C�S��q������"Or�;�I�_ 
�O�	*�P͸�*O��Ӏ��3�M3��O<q��h�'��i���
H(�x����:]�p�
�'O��xu�N ��9k���a�R���'W��feJ,o0T�@��=/]�q�'�� PL �������䍸�',t�:�(-%�,H�dڽj`6u�'B�hbJ�F���:6�[�8�"�"�'&,�Ƞ��7e����FR�4�b!��'�� ⁦ֆ!�����m^�"�L	�'�~|Q�R���ީarx��'�Nm��� �)��KT�U�(q�
�'���
�H�)"�{�KεR���
�'䄥hQe�=r�.��S�@]�@\J	�'T�{s�X�:�b�@V�G��Z�s	�'v\� ���/��)�el:3V8}��'`�A��S�x�I��z�.t�	�'x�ĸ$�ʭ�����o`����'��:���J��<��#�-mN��'��Q7͏4%8�0���3���'i�X*���!L̤4"pB�.��
�'hLx��Q57@�	,X<�@�2�'�P;0��,6>@������-"F��'�!`�������Ű+��B�'�b]���R8P7T  ��!)����'2R�Y�IR�$�2���N�,b�:
�'V �{� Bb`jɠ3��b����
�'��Y�m��)�
ɢN�4̃
�'�"���ӈWN&P�b'M�5��:�'x�B��S:R����PD�'��@��'1@�'m�#Hv���׮Ӈ"���8�'� ���� �PJ�@0ɚ�P}��'�К�	PvD��N��:A��'�0
��pJ��0�����Z�'P��k���?vi���޼s���'��"6��"z�j�1` ֆi��E��'����o��l�,�k������
�'��̉ӅŦMV&��q�[�g؁s
�'��j��8�t�R�P\\��a�'���H��%9m.��D^�XJ0�y	�'��%ӆ����E�Ύ9S�8j	�'�\���+K8��4���?d�	��'��R�N$z�ec)�2ҡh�'\���NV5U����A�A!1���:�'��ł��0)+��t,��.�,�'�<�!���+t :D&��+�1�'1�:����!p��JR����'� �3DX�Y�9p��]vE1�'AFѰ�C��\JjƥN���'s�@�!���$,�$�O4����'�Z�1��٢m�^Pď�>#x�	�'�^̺�'G=Pe���@�N��Y��'c�%J��	�x�N��F�QԹ�'}
 �Q.�&�h�F#�2�`P		�'->x2sI�(	z��k���(��J�'[��s
Dq���bI�W���'ݬh����ak�1R禘���� J���f	c��$�2�S���A�5"O�����M&ـAa!`�N�A"O�P��C�#eFY8��sx�k�|�)�ӝ[)���φ�D%��9�O�*:��B�ɩKz�	P�ȣ4.��r��^G���ݽ6����g�[
7֬��	D�P!�dA>;P2y�c������;1!��+�Qٱ�ܥb^DRqnݹ)-!�DԢ*TH<�q
�F[�\!BnQz�!�D�D0��aKT�41f��D�<���
�!bR��}8v���I�(�HC�I�0���zէ�LJF��VJ�`ZDC�Ɇ{����sHT|��X4�ˊf�C�I�+���˵	ߚR5��[��ȩl��B�ɔ4��� �O�#U��13��L�lC�	�h0q�'H�4co�0�%Жl��B�	w�%��@�(�����n�Q� G{J?��!5I�bف�oڪl.8!��'D�ԑ1O�*5AP�(�"حo�	2$#&D���Vi.��!Ud�>|eꌑ�A6D�H��ᛏu$�З��� Hw�4D�tqwJ��L����_�Έ�'%D���	9>B`�6DL��|@i�'"D�,�r ǼZ@a�`��B��3��C�	K;�t��c)j��HA�@>*��C�I.&|���B�K��ˁ	��x!x�d0�	u��~B��
�Ҽ'�'�Pź���y҆�+G�|E�g�++s0�ص.��y"ߦx�`����%��TiB�V��y�* �
� Ѐc�V�R|��
«˒�yrn�ze�D�d�6{"�%�"�̠��Or#~z��X!��d�84K�x03M�<qT�%N�t�(�	ȳ6�V���K�]�'ax�P�V.�����6`��܈3f@��y��J�.��Cp-�J$�Ղ���y�!^�\�Vђ X�8K�}ٷ���yB���#8�c�ٜ0Ԡ���(h�y�@Z��5Ar+�!�T�wL��yg�p�,����"N�*��Vf�6�y�V(]_�<�C�H݂1z#�2�?����䓢h����-:ΰ�RΎ�V�4�Q�_!�$��!�T�ʌ/{.|BF̑�y>!�$\+�u����Y������8!�d �,H2u��� �~}��㓀]!�D\Eq$�97�Ap���IS�{b�F:v;D��9Q�9�n��^4��'��O?�q'�
9�p�b�DŅ	^ք�1n�L�<��NC3\���Č���y֪
G�<��FC�.�,�B��/D|X�R IG�<��XJ�X(¡�Q�*�:KA��<y�TޒH2�ԇ$�����y�<�#!A%@�� �"L�\�����Ayx�LGx�del��ąq�4I��.��C�	=pv�\�P�0+d�гAޯTجC�� Z��@r�ԀlhZPj�HȎi�B�	7Qv$}b��C�P����e��lH�B䉁bF�M����9ӥaX��>B䉹cY�a�an�� �k�\�5k$B�I�B��.�:VV�q�c�#!I>C�Ik��B��ܰv�`��C�F=~B�	�s�@S�d�q(�q�$-�+�n�Oh˓�h���I�yIZ|�	ǉh� y��h��,!�dD�]X�pS2͓�e֊�[Em�9-�!�$$&l��c��)3�ܕ���`�!�� ��W	�ID][�ܹ&�bl�w"Oι2�΀eXfdQ�oǕ�hm*�"O[�+J�@��+n2�9���'��{Ѥ�w%ƕI(vH��	
9�D��I�RT�%(�	�	\�"��t��B�	
�����(�e�F ���^T�B䉟j�*��Â?	�8|� ˄@�B�	���,�T�,cr��7ϊ"TB�	���Q� hO���� ���qB�ɣ4�4��3��ʴI���L�Ԣ=!����'7�	E�w�e�d��(n؎<؆%��Be!�@$~KD���×:�XȊf���h2!�$J�9J��`j}��ǂL>z�!�dQ
G����2H�t���Y���p�!���H�Z��"��_ż E۔�!���uDB��������0� I�Q�!�$ǐ�*�u&�Ů:�bջ&\�'ia�$Ο*G,�pN��M�4sG����hOq��y+�'F�3�@�!k,1�aZr"OH��ͩo��jG&$�I�"O���"��?�pň�=�x�"Op1t�W'���������T��"Ob�O�1�bʑ&�p�l8'"OJq�1(K�'�%���["~�k���(ړ���H?Eװyy��F�#2nmӐN�E%��)�k��5c����@�e�3c>
��	�'~ ;��\�$PȤY��)V
�	�'�� n�.%�h���Q�;�|�C�'���8%��T�"CA I
L��?D�H!-��k'
) �( ����;D�@�)^~�K���Mv��5���O�⟘�<��h��_ټ�
1�[�N�\a��|�<Q�a�rJ�fD8 ���@$LQB�<��L7E��="·�\}b� ���c�<� ΋�]�����a욘��^�<�G��g܈�A�i"�(�`�<��FY�X!VI����a��`�q/\�<���9Z�L��fL �l8!�JT�<)q/ƀ����+ƲgW�����O�<	p䎱8��(�1jįh�D�K��I�<�D���SD�Avȅ*r#���"�AP�<�% *�����1q��l�'�A�<��'"L+'kŘB��1ge��<ID�ϯ�̉���/b���A�_|�<�$�+D`s�
����26�C��bI`��VeL�C|8A1���>O<�C�	?��B�NV
��Y�P�H�cM�C�ɞ3�z�S7��|*̵Z�B��C�ɳW���B��/;{�	#T�>YVnC�8;p�}���מ��x���
|hTC��,BD~�y%��3�\�a%
`8|B�	�Y��v"��ps�^�j�a��1D��XG���U��C��:%�AI1D���AK=(������Ԋ#��m;D�9��4`&x���.� ��8D��A�D*m~(��tZ�<7�%+��"D�$��D'k���#C�תҊ�i��?D��2�eQ�BA"�/�4)�D�i#<O�"<1�ЍIx�q鋃��IY��F�<A�(�V���B�2	� �&d��pD{��IV��L�ĭ�1L�0�P𪒩<L�B�	7��i��ז��LB)l�jB�ɡ�0��^�
\@Ң_�O�C�	'!|9�ڙ\��i��I#CRJC�)� �Ka�5q��!k�M�'<��!��'!�I-U*d�0��V�*���4�jB�ɩg�|�Fe�	�� !�e�K�"�Ĺ<�(O��}���(�!/�!Et�!��nY4��ȓ$�]
�NM(��y0"U�=o ���C `�N[��D�#�x;˄���4@���aH[�
<I`�+��LՅȓd!��eF"2��K�[�ȓV�@�A#!Y�}X� {�
�� d��ȓ0Cj�#U�M?�f���V�����?�ӓ��Fl{"I-:@j�j�'�!�D�G��P DQ���,B`����!��Q&N,�A�\9V�*d`�nי$�!�D��δ�u&�#b�r|H��	�`�{r���&r�5���y�(���	�0O$���E
j��#Q�W!`(����|��'���
��ɒ3�U�������K>)���i�=]���It��u�4���S�ht!�DI><v�����U"wBI"<�!��E&!nru���I
#���1��F�N�!�$�":���HFM�b�T��$�,t�!�ԩLF<�`���%�"�2 V��{b�$�&>�L�����V�2H �	��!�$F/�^	j��-D�Z�D!�3�!�$ �{>�$kPm�z��l����d�!򤚖BW�t��l�.6��cE��Ey!��]�ظQ2s J.F�@�����!�<o���f	9$<uѢJ�	v���8O���e�ZH%�P��B]�2s�p��\�E{r�I�b�2���U8����DzC䉓r`�,�|��}��I�P�C�IXH�b#�1�UH�`��>��B�I��F�h�I�|���q�q"O��b%�gբ4���ڊ?�H)�"O�=�T76�p@���J�P���"O�P挅_̈H����]�N�˵�'q�D�3�אt��D8eb߶�B-` -D�X`f���C�>xr]�s��p;*D�T#��;I��	�d�-�X2��4D�$�q*��Ps�M�AhI�P|�S�6D�`(�B�?c��=i.\7:�d�s�3D�ls4�]�	@²n�.�v��t�1D�����׶x��dA�&ĚwB�P�� �O��=E��K� 8X��ܤ"�4:`�%!�Dm�JaBf�ƣ?�<"4�%�!�[���uD�ą[�AX�_b�!�G4�Q�υ$LT�BcӍa�!���5O[�mȒ��I��Ͳ���.�!��Hm;��v� w�.a�A�5y#!�Q'
Q�#��dÔ=K���!�$E n��"Wl�J8�C�B�!�δ��#΃vxB0(P�Y�"�!�$��4��]a�,h�T {�!�SMCz�	�L��.�tʢkz}B��$^Z�5	��@���Jv��4��B�ɠ6�*(�NƖv���Q���j�B�7[� `vApG��)6@��@<C䉡`�`��L�I�{�XC�	G�d@S7̄i@6e�%J+V�B䉾 À �b���ItH	xBTB�I#dސ�hv
]>O�,��Ɔ5ZB�	K�V2Ƌ6L��0�B�ߨB�I> Q��cu�LN:��w#�J�|B�I�S<9(U䂶g}���+9�C�)� p{Rc�*lNL5�d�RT��[�"O�Ѩ��ޭF�6����6>b<Yq"O��p�À<=h�r�-ؕ	.R��7"O�cp��tG&� ��W�k@y$"O��	f@H�SS�H��#�hܨ��1"OrIZ��ƥZF�99���Y�v�2�"O����� ak4��`��Ԫs"O�D�+��� ����!����F�O�@ I򪉩xVJ!�7*�Tkܔ��'�\�I�)���T����J�D�֔3�'���@4 \��d�75��@�'�`��wf�2!c��[���4�����'�MCfO�\W�-�a�[ 3|�D��'�v�1pL�pj��1�n�.����'��|P3=b'�#�9�00��'F�#�� t��(q��8���'�Z9�1�ۀe2�i�`�Y�xW2H�'�t�IU(	�fy�WA��=>��8	�'d��S)��.2�:�D�#.�5	�'�|�QP�/�v܈V��S:4�X�'�f�c���.��0�fE��G�Pd!�'�0�]�p�t���DyH�q�'�D���醲FF1�����Q�'C�l m�J:pYгǏr`@��	�'��S�g.$bm� �+`��TB	�'q�렢Q�O�����!X ̀�'(�mՂW����ζ_��@�'i�9H����q��a���:�t�i�'$n�P�[�QB��*!��?}����
�')ʐq1hޙL�
0� K�L��S
�'� T�*P�O�Ą������<3�'�IR�J��E/��� c7xA�
�'֤t��d�>!5�]�i�,}�t��	�'r�z"\+?LTqI��+t���h	�'�i��G�s#U�w=�V5z�'*$ ��t����ug,*��}�<񀥗tji�PA�v����c�|�<y'�e���@C�>$((iB���5!�$�X
XI� ��O� 	����d!�D�8�t��R� �:�*��v_!�DV�&����n�.�.x:�H�F�!�rJҼ�ŋխb��yQ��u�!��?8�Z\A4�͖W�*�K6Fľ@#!��5~݊$��%����RD$2!�$.-D�E�dQ;�L�11�_;(O!�$Ő'�*��z���1�gٚ35!�D�g&�"w!9O�E ��ڈ+!��Y\.E�e��z=��6�Ռw�!�D�T�.��vO�;8�,��&R�2�!�A`�\�[D�Z���(�f�G!�d%]�,e�TƘ����� �9n!�d�u>�,z���^"�aڂs�!�$Z�J�:�nܪbD(�7+21.!�d;`�)`p%)Y,�1;7��]H!���yfM��iwܤ�p [A�!�D�M�8T�6E�#.(!�e@ڸf�!�fNBn�c�XO��fm!�Qw��J�GOO�03-�%�!�Bu����ġ��2z��J5�!�Ă�:�찕��6vO�!�K\�!�DX$i4�H�#Q�
M�eS�j�!�D�%x��u
!
�T�Z1cI�y�!򤗸Bj�B'��!2�`�rա�%:�!�D�'��u�d&"[�!���70�!�� ġy2�âi	v*��1`� cs�'Jў"~`(��K�V�ɣ-Fp�bB��y��Ļ#� eQ�\-4��ґL;�y�%ıyi���`��M��y"��o`,;��E�	U&1!�	G��y"aVM�$�p��<.��� m���y�˃�y $�ă�%4r�� �� �y2lU'iy]��eK5r�0c�@҇�y"M�=)l�+`���%���yR$�m(�4���	�@Y�����?���0?ŬD"�AY�͐�b��x6�Ux�<�f��0=�*xA ,I�EC����J�<���&$���Z!,�0*l�ѱY`�<�J@#�|<��G��z��"g�<��"Vg���kCd��cJ�ѐ'�J�<��P��l}Y�B�H�0��	A�<1Cљ^�$%��֙v����@��@�<�jH�Y2ڕ����+}�"��#�Ht�<�GС#\*�붬�#e&��1�o�<5G�dd�(�
���@�m�<�`��5��BR�5�7Ɇj�<�b/?�����َ8�X9�3)�K�<Ѷ�Ւ1�:@��3_b\u��$�C�<��V w�ȃ`-�.YLH��C�<QТ�`FDp�E_�?In�SH�i�<�eHޡi�i*e��'<�@��&h�d�<�FE_�tj�O�2rG�\y�<q��$;���,�qc�E�3d�{�<9J�!�|��&o���E
�w�<CL�>{@���F�ޞ��l�vE�v�<�`C�<�Z�B�J�VȜ�0�ȄJ�<qC���R�3��t�`�N�F�<a *��]܅Y'"��H�!;g
B�<AF,��-Nh��b���G�b�<��#�n�c煈�Tb���X�<	.<y�~%#��� Q������y�<�&L�/3RٱP��� �dor�<�3'R�};�e�S*�,�(A�r^m�<������4� `P%eݐ0,�`�<9@�w��������ٖm�`�<��̚k���B|����g&Se�<�E�1)��*�R�2��@R_�<af�I��@�`�*n�|�""�a�<��A.U��Ƨ�(~1BL�ρa��d�|ȉ�ǮG�=�p\b�nZ	!?��ȓe��`2�kܴ(2�kA�Ă?Y61�ȓ4���A�:!z�;��Ά���ȓ)�$�x%`N4I�<���T6pHń�K)�����2`��b D=<�n��ȓ5�����O� �քb�ƞNHZP�ȓ+^
����W
�X�GA���M"f)�v�G�G��������B�GZ�<�wɛW���Pk�6Jp����^�<��R�MF�b�J�0 Q�u�c&C�<�A!�
T�0(T��0ߊ���|�<Q���`}J��F�.t���x�<Q�H�6qX��1�B�9�����Ur�<A��^�i�@qy5�M�6!4D�� Jo�<i&���p%��Pp�H�{��<�.6D�,)�@Q�=�4AC֢�.}�H ��`3D��`4鞐c|�l�2%��q�jg�0D��8��!�4l;7I�:è�Q�/D�ȂU�K�z��HђG7dy�@3��-D����$^� 8�OG%NB¤�!d/D�� �1�atSt�{��5H!�'�H���Ӊ��M�U.���@piq�,D�ɷ�Ï]a�Q�/�.?j���*,D�xҨ��Q7�:RD��45f��J+D��*���kWl�P"'��|<��:#E*D� I�/A�d����è:)��C�&D����Z�1yBQ*�6p�d\���6D��j�6q����o��
<�Z�:ړ�0<��o�|����V��S�6t�S�~�<�E�TV��ꕪK$^1@foE�<��%^7	�*qp�,�G�����S}�<)f�]�@������A�*��as��O�<Y�CB����d@R��B�BHp�<�T�6�Z,!��Y*��WҌ$�����KV��Q�]��\�a��2�R�$��I6"n��36G�9_���U�.eX>C䉘{����t�dH��0�XB�	j��z��ʊ"|�|ӕ�{�BB�	�KN��ȴ�
W,`�9e��Xj.B䉩x��lGM͌�Kq���`B�<v�PR��	'�h��o��P�PB䉊c<VD��.�:t�(u�U�ϢO�F�$,�D(�S�ɐ�4%��)�R]�l��N!�$�+t��ӠoO�!i���A�I�7!�d�
{�@�J�I��AvTi�f�!�Ĝn���I�o��[^�H��KN�!�Dݷʲ-�&�_8OZ] Є-6�!��2m�!�:@KdQ(��B�z!�D�$4�`�p�L�8H��*�◜r$!�D��\�2-����5�:�A�p!�"6�<��ƞq�Xtp�@�)!�$��Ɛ]2��0mtR ʁꀎU�!�d�S�y1��>���;+�!�d<#��і���#B��RW(�: �!�$� J!T���+��?�6y��Qb�!�$�58� �*�/u�B��P�I�#�!���
$�(h0bϢ;�>��%��|!�d���8� �ϺR;V%�C�	x!�$!?��v�^8�E��H�!�$��+&��; �D�7Bµs���qp!�D��)p�,B]L��R�H!�!򄂔8�3��8L�aC'N�	 �!�Dʵ= �y���L�=�,�*�,�qp!�$/:1R˕%�u�jyS����-!�db�d �ԦP���U�TAƳ�!�Ą)�19�(FO_�]�j>�!��W?'B���̐�T5X
�'^��!��{��P8p��AE�گ!�Q� 8�F�B����m�	<�!�d�,M�m� �B�w���׫[�)�!�β2���!y*,L˕		M!��3��ã�'E��(�E n�!�ڢ0��D��(V���YAC���!�� kF܂�/��D6L����!���V���ؗo 6w5F8*�DV�i�!��R��!��KK^ĳ�#��6�!�.h��@�X&�0���#�!�$F��(��UHzw�i��� :!�D�'��MBsN�/]��WB !�$Ekf���֦֘$*��P@
!��	�:P�7��)]",��+W;R!򤇀-Ⱥ�{q�	84�"]y6�=&!��"&�L@�EM�<��a�V�.�!�$�QE��rG8}s&}A�	�4�!�� v�A���mn�0!��"��E�"O�,B2W�&d�H[P	�CK洈�"O����=u7�����J2���C"OR�C,�;�t�!�� /��"OJ��3���OZ���A3?���2"O�hQ&��1gȔ�E�)�%z3"O�)�FH�",�Xcg	�AlI�a"O��y�J�� Ձd,�7�2�@�"O0���O�3�|��$L�!k��0�S"O�0!���T��bD�_��lYV"OL%�FM�𠘡���%d���R"O�H:pl�9���5��1Xc8l�u"O sW�F#R`H�TI��G�I�"O���LG�	!Fi�d��Q�c�"O��á�,O�p��GN���!"OZ��7-#I���j���sgn�ҧ"O�)� ��ME�R�d �T�|1��"ON+6��,>j�RAS��6�"O֝�jՔh@NĀ�b�i�Z�ZC"O�mk��u
4�0���e+,X "Ov������J��(s���"K�x�+V"OL�9�G��>��/��G����"O����&
	E�]�&%D�;��݊Q"O�{&�L�tLDЁ��ˤz��bf"O��7�̈��Iꡦ�=�Мcg"O`�j!M��ciԎU-�­	�"O(�;W�Y�JJ,$�� B����@"Öi��kر�5)מH��5"�"O~�����%�����h� ͪ"O��!�����D+@
�,��`��"ODi��E-cX�ݘ#�C
@��U��"O]@b!L�	g����R������"O��2+Z�p�Y�OM� 8K�"O��B���2sHq:ƎC%w�>�Xp"O2���bɽcH���W2|jbp"O&�B�S�lP�?mBH3 iU� �!�$��]��E{3e�j�`���7j�!�䝜K�,�w([!3�5+ag�w2!�d�2d�"�K��Fe.]K�H�7)!�$@$
��,�d�6|�u��O$p!򄓢p����Ŋ���Г���!�D�G�~���/J��A'͖�e�!��
�&Yn,���E�EՑ#MWY,!�dEr�<�ŧP�yl��˂���!�$V6r�(���P�(_���.2
�!��
z�Đqaʒ�D�4�R_7{q!���R`��#:�w�	P�!��Άg�&A�$F^� ��B�_7_!�dX�/���"��1�**ƨʭ7�!򄊞@���a�*M2t*�(�|�!�ۖF�$��ħH�����!�ğ����6"
@,�I�f����!��3X	����Ǒf!҄�#I�!�!�䏻��8�
 ��B��%i�!�d��X���9�����Z���y��)�o�@�)�NFф,���B���
�'S���0��R(��D��
�R�[	�'Oؼ�ƈr,�bs�Exdu��'u: ï�:xtq*�B
�r���A�'���q�9I��0Ӳ#�T�l�
�'�z��Ъ���Ԡ��J&P�X��'JȹPqi�.�2չ���/�E��'pT4�(�Z�d��C�Sbq"�'0���/P����aE�S	XxPPs��� aH�зB+^��ᩞ�f�RŰ�"O��B�%,|Z���v�ؘ@gڔ*E"OrXi�,�&��Ț'
��*����"O�{�V^��#�x��}��"O�Y �^�~:�R�([>�n�c�"O����4_�����Ҍ@pHDy"O��!�_�&W��1d䉁Zg$9��"Oȡ�i�>@
z�St�[1����"O�I�m�kΤA��:@��ѳ�"Oڝ�V��=JL�Z�̅&� �bt"O��笐٘���4����3"O�d0�m �.�h�*p��_ �2E*OL������9P���  �'Vf�'ڦN�R!�f��~Lt,��'�,��GMC�<��l�e�ʀh����'x!�B�r1H��(��`�	�'V�ذ��	l���$��]�
	�'܊MP��
�X�È_h� �	�'L��	`�)T�����J�:Q��9	�'�4`cB)@�pJ�x $�[�H J<��'˪XXժP+ST|���W"H����'�j��
N�7|0�8nNBjd���'�\`��UO\�d���3j~��'�� �͘ M�t��%�;(���z�'�txEb)�����T�"��!��'O�9�#W�zL!"螹e�6���'bN�Xa�GN"�`�� ߳V�4H����hO?����ޞ5~���e\$E�����Xr�<1Q�J
&���Z��T9Jꚬ3Qa�B�<1�&�&���[���]��$ Q!J@�<��ʙ�`�
��U-
,`�.�`b�M{�<��c��n����,ݹ�Bo�<����6kl!��L�6]�ya�(�l�<q��3
R�WP�"��Ō`�<	�k�	e��$cТ�T�Αa���g�<�w�[T�!h�U=� �7.^e�<���}}���J�((N�Zԣ�_�<�b�B�r�e� 
��u�G��c�<�-��.��9�ȃ f�!�%�b�<aL�
/n�5�`�qC�1HF�]�<��AY�9c�<��d�?v�,���.�A�<��^%>|�#���2�$�3 X�<A���<e#a�</Rm���V\�<���\�pU�Ʒ/�`C���[�<��YA�A��7Az���s�<�s��l�6mblB0�����`�F�<�*��w��-!�Q��HH: l�{h<f���\5Y�[����cF�y�Dw�f���Q� ��e�E똉�yRh�%IrA�u-T.q�T!��h�y���T���(a��]�~�#t��4�y��ǆ��Q�j�Z|��	����y�v,�R�N	�N�R�R��?�y��G! �&2M9�`j��=�y�+�D����P']�Fj���M�-�y�ͽITnP`�C�L ��W�y2��up󴅪1�^"�J�'����C��	�6��QCX!d����'��iRÅ� RHщCoN�bGR)��'�r�����+p�9�0W�|Ԉ�'��+�'P���� �KH�t���'�uCs���� /B#�L�A�'�h��!-�����W���*]H-��'� ;�O�e�qq�gO;o�>���� ~���s&Y� �>m��h�@"O���`�0%����/�����"O ���A��@��#¥L��1�'"OzR�Ƌ3T�љ�eKn�Є�'(��zUɄd�|-����15hdl#�'Y��{4ET
[�*�`���ţPj�<٣`P�`vH}�"K�H m II`�<ai�av�w)�7�N����N[�<'N�:�xX'��j��X�La�<!��/Z} *VOѾ�NhX�TS�<�5D �D��`��6-X�yd`P�<1��X���8���P���;&�M�<�0#�9�LSfX�!\(�%�
p�<� �4e[��͕x`I�T��k�<�e�J�x�f�;(C�ZMR ��Sc�<�t��=V���@���ʔ]�<�*��	�>=ɶ��!l�}��g�Z�<9���Bw�2���)u`�� ��q�<y�	�4k��PbB*�#[#�5���R�<I�#�9L�v�f��p��H�ĀV�<9.AVh�l9�����`e�N�<LK�{����&��=�<<�%j�r�<��l�7$>���*��E�P�r�<I��[�^��襧�6Aݖ@�ơGq�<��� ���Ċ��< pp�)��@F�<��ǈ.,l8��v/�#!�)��+
B�<��
�8@�\L��d�4p��R��L{�<�b&�,�(���jxϜQ���v�<�����q%H�p�SCs�<�5d���@�dL8 �F�Q'��o�<	�CZ"Iщ0��
N�,�#)�o�<9d@�аS &�u�i�<YK�%���Y�iA՘���GJ�<����[�FXJo�����Jk�<a��=h��Z�Ξ
P��QIP�}�<�	�==��YpHR"�v�����p�<��KD���,���
��&A�I
n�<QU�'r�⹁t�س�aF�<�ݏ%BDpلoO�x����Y�<q3��)0�p�C��>���a9T��J��-q��,
1�tN*D���r��0�|2ÉEV��V &D����ѩIk�L2WF�yy���ƨ6D�P�D�j���V��R��2D��rkV�Wut�#t`յ~��(14m1D��V-���������
:q!�d�+X�ԛWK��B�Ƥ3'l�{e!�_3J=d4��,�0��NK�[?!򤎃~FȀ@oA�U`� &�,B!!��F�e#ye�?\Q�5�3cՃ+!�Ą�qs�2��g7�QBX�P�!�8<��Yԭ��d����%t�!�B G��d�f��o	p�h��]$!�dZ�pѶ�T�:��a�f��!��D�U'�I��_d�J%�� x�!�$��E�>�I�n�D)�! pB��Q�!�\�H�5�+lr�RƆ�7lt!�D�G�j�`ҁ�
-�R���"��!���N��a�` ���@aU"\�!�!��(*�V�X���� e�	9!�$�_Z�[�ρ�a���Q6�@�K�!�D	3I���3)Ͻ3�)�f���g�!�A�l�r�XBE�,�+&��E�!�$��N!���
	�iɊ�M�h�!�� ��Z�bPZ�j���)_�fQ;U"O><��F̯~z��XDH]���EC�"O�|��&=x���8s��18�6��q"O��O\���vl�-`��P!"O0�Q�.�$K��XS,�<q�D�"O�ъ ��<��Rk�h<T��"O��  d�5R��x�鑆W�ʙh�"Ov:�TB���ai�x.�`PU"Obx���c������h�
�:A"O
��f���6zaV����"O�EA��PqО�Y�b��H+��t"O�����:젣#���y�Iq'"O�ARR�O�]M գd ޯ!	�}�%"O���$)�}�H�p�K\� ᱷ"O2h�bD��b���:G"O��'';'��Ļ�E� N$�"OB���aUgNTs@�c����"O���Q�L9b^���/M�U��"O6|8`HU�h���Tb=/�y "ODP���՞0�<�3�fËXs�}B�"O��g!��tdU��|\H��4"ODp�/�⭪�d@#*)�"O�(��@_W�x�1B^-8�.���"O(���R�^��f; �^ѣ#"O�0���n�bђ �[�=TTR�"O8���ݪ�ְr��Y�m!.�3�"O�̈��$�����dX+�Ȣ"OlI�v ߥhE�UP6��PzQ�2"O��ca�׋"�nDQTL՝a;���`"O�YZ�hV�.�h�e+֥�Y�F"O�P����܄����d�>�a�"O>��j��,xA`�CԒ����"OD$�߃g/��� ��G��%�"O>iCve˙	�����X�@��6"O�XB�/@//D�x �͆;V���j�"O&i��,�zج�1GBF<�Y$"Or��4e�.>�A����c�8��"OX
��~��0�E�'(6���"O*��%փ2��B��]9kk j"O޽b��&2�R���DB(,MdD*B"O��!��	�`)#퉷"O�qr��	z�����I4���"OL����\�/DUCa �if��"4"O�AXQ�9u��kch��*z��"O��ς=��)G�'��y� "O���MG�O��	h����Rt�!�"O�=�� �4P���:�j��"O:�'�½{�N�y)�����Y""O*��FI�P��P��.l�p�"O�1I��]����c��*���"OTx��至D~0��#IX�Aӌ�г"O��x5JLH!"!��F:VD�H�"Oֈ�ׁ�rǌd�5��^3Rbp"O�3R��Vt���Qg�9p�G"O���A��>��D�W��l!�(B"O"ŲM�At�h����1[\PW"O�uBs�V5)���U�ʵl � �t"O�`BC���Xs W�2�:Tx�"O
�[���)Gh�@� �4I���"Or�@����S�O�_��dK�"O�Ɋ��O�`��������)r3"O��ː��8Y�Љ���Jr��2�*O��g��7>/J0�ը�5!~L��'7�`�&��@>Z8��,:`V}	��� �Q��έ&ؠB���,��Ī"O<���*a������޼��"O
�2��jXۖ��^�(���"Oab�������*zy*<!e"O ����99Pĉ`�f�<v��"O2P	��D1��@�F܁N>�UK"O���v��H	�惡*�<h�"O�Sp�Cqf.�IqhPs"rɐ"O�9c֡�O���F���9d"O0l�d>I%f���@<�q"O3ϘF��{�ǸVF|G"O�2w�.Uش}1��rT84�R"O�I9�B�,�:mx��خ=�����"O:�r�cQ�))��0	�vК�)�"O"��m�0"���)[ݴ�"Oz=yg�7t��@�,�1��"OdX�t�	;���JY~�i��"O0RFD�?i�D�[�ȓ�O(	@�"O���2��"@a���(~�K�"O�`R��ÄK\�g�g����"O�t��8n�h`��%�c�FN�<��Q$ͅ�3�Еb4�?
|h��"��G�7ܶ��#N�<Yn���ȓ#=��`���>���C!�Wu>���XZl���G3�l���NԷG��\��?��=Гb��(��{�G�C~jB�3@��\"��ځvF�]�gf[*1��B�I�'"�����f��#���)��B�I�x6���Ot�q�C��v��B�Ɂ$3.dgj��+r0tW�@�b��B�I�0ᚰ��GBpa��ʶƚB�d��9X�!ԃ.����� (7(B�I�{����ٲ5Bt�а ��0B��b�ʵ�d�J�8��焗2OnC�	�����ؒ5V�	��C	8�B�	:Z�XU�C��s��y˜!\͈B�ɿn�xG�& �����n�)b�B�ɿZA�ɻr<i"4 ��-�^!�B�I�g��T���]I[��� �B�I3��u!�2['  ڱ�(8��B�Im�t�2�s�����V>h�B�/TO�(�
M%E��k5���Si�B䉎=ތP�H�4��%�o9A\�C�	�v����j3(�^A�ә D�B�	qh�As�AW7�0���/n|�B�	�[��=�sϙ��@0a�ՀL��B�I�n�Az�F
�6h���a�C䉽@hy0J	��e+s��m��B�c~�����F/d�_�ٚӨ,D�0#��/���k�bѾw�:�v 5D� �֡Y�YA^���,~8QH0c4D�\Q�Ј �N�Ҋ�
K -
e'1D�$X���J�����Q!b>��Ԧ"D�4�Dn�bh+�Q'I��I*A&!D�h��!��T�`��Pm�+�p�SN>D�HrD�F/e89���WtP�<D��x�)P5T�\㠡C+]��Uڢ�8D����j�v8��N\�1��#�7D��*� �R��K�#{��=���(D�����
�uk:�
g�	���ɀ�%��0|�B�;�bHUCP�n��Dc�l
E�<q�^`5<�A0���H!���<����Y�-҃�U��R[�ē&�'jqOl��,>_ƌ�`�y��ʇ[��
�S�? "M�2
K��l *��ӱG�0�b����>����CNV8�To�w�D�B���KD!���5Ä��j�z��`H`�ɱ\C�d3�S�O���Sf W�C�E��π[dc	�'��YAf��C��0,�/0�y��~�9�.��rd+�0,�����U>�����I�<)s�b����Z�$�E�r�<��]���[���l�:�r���l�'??�+@��4$`�`S�:�`8D�쩱��al�Q@f�H����4D�8���NtH�@�1`��8W�.D�HyE�3����$%��bF�!D����@=���Ɵ��ȴ3U�>D�P�aI�5:��%y�c�GC��ZC�/D�<11��i�X����~�R�I��"LOP��٦��%w��10��#,^4#�. D�S�+N�6`�)`ש"n���c�>D�X:�
ɋؑ:��� ��vn*D����n3�qA�g��p���34��Or�=E�Č��R�
�S0�A�����hC	��}␟h��JO�1�A��Λ!���6�%D�����
�x�r1�ǨM)<))$�>�Ԟ|�U>!G��
 =(B�Ȇg�&u.��5�y�f� ����nB_�@@�M�����p>i��.�z��^.��C7�Kf؟Dh�'������|�}@5ߘ6�F,��'>���C��dD�t�n��B(LË�&�'4�)���)s��S@���'a~�9'؄�X K�
�2Ȩ����yҀƧ[�|P�B����${�⏳�y"
�8i"��X�d�	����bM��'Hўb>�s')��wM�l�/œ\ &l0c�#D�$�#$�-J��,[VM���8!a!D���$c� 0&5�S��r�B�0� D�D�6	΢�Z�iS��)(��k2D��1$�G��X�t��r��!� e2D�tp!�E9 �6a#�P�!e���D+D��[��7>����n�+?���@$*�D=�S�'�􀠡�W/L�������c�����O�$����s��� gɨl��,�?�ӓv�l�Fɝ�q��fX�a�~=�ȓ,����@�kafD��?B�H��d������%q�9����IY�K �8��M"\::��/Ӷ1�R�Gz��'�p9��@Ļn�ư@-��lzm��(�S�$�ןr��\)$�*�X��:f!�dE0}�V�:��H9&���jdO�:`1OZ�d6�IW�S�I��E%��U,�) (���$6?Y� 5�������D��Ў���4�'�ў�>���VY�H䈂�$��o>�Ĉ��6-�hV%�,��=��@�.��O���$� r8X��F�2�ʈi��Af���`fa� V�v�u�6ϝ�Z>��+���(�yC�3t$�l���9N����ς�ē�p>�U�]�N�{�O�~*���K�K�<٦*\�h:2d�MY48��x���K�<їoĀB�|}#��9z��d��AK�<&�C�8�!�γf��CA��<q��Dz�)I�鈡qt���b�5��l��Mv�ó(���UK
-D��2S}�<1a+f�Bm8c��1E���e��@���ē{�$6�$��|�C��$N�	�ɓ%١���h�}�G�^&���S�KE���OBFz��t.�4h��)�t��9(�]4�����O.�~� �(�$=p�ԋ�B�d�F4"R"O�H�B�<!��X&Q-r�0TB�"OF��U`N4
P�Y�KCz�JP�"O��iA̙3H��J�m���#"O򨉲EE&>�z����ϧl��8ȆO\m	b�]�Pss�%��%��
Xc�<a���_#&�SRr��`k��PiX�HFy�
�Z��,��$]J��5�y�a��bA��7!���$S�p=����#�pa����R#���d��!򤎑f�"Q� }pb�фc[�ڱO��%��D���8V��HX2�ٿD�d�V'�W�<�D'E[� $�E.D�I��a��/|�<1�
ĒC�5J���6ly�hʓ(L{�<�L�*0ҡϟp�L���Jx�<ɧ(�p�d�����p���oj�<	�	 p�8m����= U� ��\�<�A���޵KE+�I &)aA�DY�<�BP _�� s��65RT���X�<YQB�X��JE3PD�v�n�<�l�>>+��($N�Ay$Y�!$ZS�<9�G�6����w��0N]��#�R�<QO�9����ߓ}A�Re<��B���O��H#�ϕ�������j���K���'����W�:к���ܾ�ļsÓ�hO\:įX�OU4�A�@�R%� ��.�Ş\e��Z"���1��0(�;��1�'�ў"}�C��0;��y:��~Mje�b�\x�<qƊL=�f�����.b1�HVn�<�e��s���#��j`��h���<�'�ўb?բ��IK�@T�fطFIl�;uc:�OF�Or���N@41!KK�NP  "Ox�*@Ö>�p"W�@���1��=�S����y�@ߪW����B%]�M#N��-�S�O�$��a�֨!��L�H�.kG�d�!�$?�	D�V���`�[�j$x�� �4;0|�'�a~�D܆%G�D�712|P�I��y�8��:� B"bYMZ�b]�y̉�u�l1��W�a(v5	Ŋ��M+���s�j����'OJ8���R� �X-��"O4���C�ztd F	P'd�M��"O��yA!�)6 D�G�	)�*����	m����'$�t�ҩ
������Q)%�$��SF��G�&;h8���	hw�n�~ܓ�~���i���[�n�09rwk\��H��''��&�,�di�֥�P���'aX���B���(��D�*,X����DVs���)�.��t�^QD�փ0=M!���{��O�ca��J��1�`��)�矐����oD�, �,΄@�
#D���`(˜6���en2�ʆ7D�����FL<�(�a��S�9�2�2D���ąB�
!`<����)ͪI*qH1D�P�pL7u��-Yf� �v]R�W0D��/�l��-�:M8�(�&A���B� +@����:tp��V�_�Ma�C�	�Y�2Q�t�
Q�5@6��'B�B�Ia�A�Ő�#���&+�7l�C�I	���i���:R��5��M&�C�I�]Ab��eM\*g��G
��8�ZB��6U��!��:v͉3j�~6B�Ɍ*�A��N$C[Xa��G&!!&B�I1&P y{t,R0q~$+�'�B�I�����#�z!��8ń*~��C�)� ��RŌ�2�"��%gkd��"O�my�c�9���h�C�v[�l"Oh�8ǁƿ�T�P"�_3F`�X�"O�u �Ɖ�p��E�M9@;���"O��ʤ�G�LF�燷q9 9g"O����[J�T�@wEr*�-0e"Of �Ó�M�>��Gگ��Q$"O�Q��D(�����g�K0���f"Ov��Ă�ic�I{a&���B��"O`�ӎ��7�H���j��y��"O�5�Q��-U*^	Y%"O~�h�d��-/X�����1���z�"O���`��5A��:TG�ȼ�K�"O�x����#G� �0@F?v��h
�"O��a+)�U��B$�x�� "O����
5���d.�*�6("�"O�����H�K*�ac�]�9��L��"O���S�Ӗi�h�Ѣ��;�V�"O,��d �Kz!�hR�K:v�9"O�*�*JVq�],u�.�!��
�y"!Ս�JY�A��Z��zCh���y򡆂L���`DMf��QS�׋�y�B�7r����� p�0���yR�VR�n��@�\�^lF�Qd�D�y��	�H0Z'œ�Q���
�,]��y���*���:Ԇ�E�L�#����y�'+x�0ٸ(�B1V�L/�y�*� l��r���w��;%&G��yb��'EB�R&Ej���)���y�,u����5$����EC̜�y2�.XL,e��=W;����C��O,Z���p�h���W�,4�6"O���!�U6}: ��3��0c�"O�}��g�+&�(�	�a�� �<3U"OL���2B�Y*�a�'b���4"O\�T�5+�D� �ڵ4��p"O�T�`ߞW�r)*���(6�<��"O�$�6�!:�`�8 �Q#��x�%"O��2Ǫ"VX��,��k����"O��[�i��;�v�ʃ`��&C����"O�T��〕\;��U��JT�Pd"Ox��J3r! 2���j9��a"O���M	RA(\�e�юlq�]	a"O@���$Y�r��2�U��z�"O(��$�K7�P��Ꞃ(″�"O�@!1?m�E��,Q�I�"Ox5�3�R&�J�h��G>r�>��"O����Χ(�.���j.y�����"On`Z���8i+��J}�Iڀ�yB@�I�Ȧ /ؚ����3�y��לs��J���r�Z�� C��y�b�8L����1kp��Si��y��VZ�X�	(̌�cC�R��y�*]B��c����j���C�l2�y�,[q�؜�f�-6y�a�HJ��y���
9�Iq7���*��0�/�4�yR� �z¬�3�b^5�%�ȁ�y�-*1`�f7�x j�掇�y��I�W�V=�M�
����1����y�.
Dܫ��Uw�T��/_�f�P�!�}�S��y�!	�<I�+s�D�����y"��:qhv%H�kk0x'À��?���~ظ�u
%UM�0��UүAM�ф�	�G�)psa�;�R`T'�M��FH� ^��$I��y��щ��9��LW�C��B�I��'�ؙ)rAJ9C!�F�� �����غt���-�F��xBd"Ot��Q�%-�6��0L̲[����$�ǿ�hp��(3}�� �g}"�P*�"���'Z3�-�5�O��y�/�]��3aᇉ!�z�hɅ�MS���v)4�a�#|O֨���S��i�M�X��	� �'ﶵ�ӫ�6d���I!07[�Љ�����2Ǻ\�ȓ9 ��r%L�L���RN
XB�=�>�ǖ�~� �f�5�'l\���C�M>`T�����F�Amt�ȓ6�ҩ���Y�k*��+r�SO�4�C��]�:h���N�l ��Y�� 4��~�\�S�$2�V���G:D���D� 6hE�ĠU� �C�O�B���LX��D[F�\�'*�
(ɱ.H��a|�̎tCF�h��mX���]9\5(��4/65�ȓz�f��rF�U8h�[Q��?�@��s�"h��:�0��䨏j�,���aj.P��To��	��W���ȓ^�r��Lښp������Rm�Q��!ܑ��*1�<)���_�4B�ȓ7�R%�ŪK&
���I)}�͆�Z
���+�[T���MܨS><���JH���숈p�nQ�o)Gy���ȓق�{"D�b�� ��O�FxΡ��h�@���%n�i����`�6N��X\��"~ΓMP� p�`�)|����L	f���
i\�x�K�
/-NPk���`�1������ؒ�Du��K�H�CD$�ҍO=��룣5lO���'�C1v{~�J�I]d,��"9K�U�4� |&=��e�2(��I4=��xB�^,R벼��P�c�	!��e��sr�i�f�B��]�!'�1�O������iO4�9�Pc�m%�y�f*X����%V�G��kaM��Gi"�bA��8-Y`�k��@��,AH�&S���O�]>dx�"��O!pCH�B�I�=5Jx���wZac  K�={���#�D'k_��(�%�6����k�� ���( �OF!ɢ% =��\:�(ͧnI����'%�����X�>�Z��K�(/�4+��fÚ�&���0N����
C���Kv�Yn��h+���7
!b�ۘL|��P�'��{:���ɳ|�.��!L� hkRɱB�؈�ݮ;#ܜ��#�4���+s�G�QhZB�	�r��l��g�1JS�-Qe#N�ǌ�y|�d�aY�aҡŘq��`���D�d�)AU�P6p}"�RB_'v���x��"��:v��i	��S/E�i�-c�1h�D�`8�^,���356~4Ӗ���h���E��''`����:a�����G�=���{�l����.,=0�I�����!Z��[�T$T��¬^�R�Iae)qE�(����"��e
5\O�P�JsN�q��B�j����Oj�P�2D�&�tcd�d�-F����,�J?T�x��B�P;�T�R&R8�
�Cs╵j�y����%.g&�[	�vN�9���`��EyB�����I�4O�L!V
 �F ���sF���~���=gx��]�e�&91�C�Wr�ڶ`�_���D[�\X&dQ���O�Q�gG��%z�]�щ)J�Ac�a��{y�Ur�G�5����4 �6"�y�7|>Yۑ)�(N�q�z���[T�W=��`���T����u�I�2����7�U�'p.�����䋈�{�Z�f��I��5�ŭ�b����狼`�, �$j�X�0�2��+u��[���HOx}�wF�2q~H����-w��2&���{`*0C'�+��� 'I.c�^����a��O���¯�M�V/ДrÈ\ �`
!O^h��g	�E�K�gN �q�FM��H�&�X��GG�i%@�C�䁮H��!Rm}p�h�6B�EK����iB��Sn-P���.v���O��T��ja��$�Z���(��y21�p����@P�F@�\@NJ�MA%*C��I�JD�u�(�T�7J�Д��GA�	Q&!���ħ�M[m�1:�+��ء����D�B��4Y��2@�[�f(T��_�B�
i���;���AV\��)(�P�c�����9X��.m�̔np�1(;����g F�*��R�"5NAk���.��1�ѫ	*[�$r��4�?�O����U�!2@YC��.��C΋B`�ԱWa�?$z�c`��!m��tƈx������f�(���� T�E�������18^Ya���[t <i�(]�g�.�ɕ�b>�*c	��Y���s��3<g.�$�:|O�9��8B��:C)U9n��'�Õ#7��+^�v��%g��h��b�>7�Ul��N�r���'�T)ps�
�k<�eR&퀕E������ğ=���r��,�'mxj���H��ԛ&��L���W!6qnŇ�	�e�:�r��S[�a��!ׂGnQV��.&��"~�I�y�� Pa	��x^��'�T�o��B�)� � ���f�L${@R�/�T܊"O\��Pj�eq����\9Q�l�c""O���F���*����[}2DA�"OQI!��2A�(�C���`�^�)�"O�yc�	T�1+�y���+,2�C"O��y��p�0��F9p�8A�"O�q*&!A�7n\ij!�>e�tK"O ly#./���H�
H\xu�4"OR���M3�Y����2y@F�xT"O^�r�(Ͳa�tD���
:�4�"O䨩���
_$9�1����~dc�"O����hX'(ې�7h�V�"O�5��)��$ �`�*��@k�"O�h�AI�!f�$�� \�k��a�"O�a J>�.Eh㏜	崵��"O�!�uN�m3�X�U�W!;
���"O6=��@��4��� w�G*k<���"OD�2�7O���6�M��rhw"O�I���E?S�=y��̙O��ժ�"OT�B�']v�(�sr���.��e�'�~�@�K��qє����n�np������t�ȓ"����*�[���Bɖ��2�F|B��0VUar���l��v	�B�������Q�!�V%r����ȡ8ऍJ6)�&u��n��1Нr�Dӧ��Ru���:�|!1��	�N8Y3��#D��ȔƆ�
�)�G�8{������<���'��ͱ�?,Oh���
`���1@�*|Q�'~R�W�^�2���R���dC��IlĠ3 �aH<y��)}�6�a으ZmT��%�Ih�'�T�3����e	�~
w�Sx�*2H�T�9�a�`(<1��+P�j���٭U\����tY ��φ�h���:e�H���	M�O4�HYBoٮZ��(��d\�P<E���'�rźF��.'��'�|�Z�@ۄ]����ȔA���)Or���� VRTQ˓P:FʖÆ,o]�2`������'��a�w(@<kK*�O�ӓ
���2գ�-Wȉ�2)V��8��N�*4���bO�Q@i�="��C&��{I���ʛE��L ���CS��6,*yR �d�i�= ���@e���ukY?g;6IRV�1�O)8 FN�S�|���М2ʞ���Ó��5[�(G��9��9��M�O�t԰�DO�j/>�
�F�^ᓊ���>{���4�T-�ħ]|��DK&2
�V��/5fU��3e��ae�҉.�XA���>�8�'%�(3��\1^D�OQ>�b�-��fʔ!1!@G�:�P�$�y��N�Yo�$�D��3�����(��'"n��F!4>�ϸ'���)�d�T�ip��;���3	�����Q(ڌ6�BY;��rS��J�K]&���@34�O:(!P�s����녱f�J`�B�'����_�\.�'��=���ׂ��Ԩ��~���:�'޾��hʧaAV��ɕh*��M���*+(�qO��ݓ�$E�xg��PLôT�����"O�K$��*�b�����$����"Oj 	�d�k/�����
�f츠"O�@i��(S�f��U-� S�"�"O�|
P癌&2H��������)��"O���f�5x�P����j� |�F"O(@Xb�^~��qs�D>�Fd��"OX���SP��:"eW,Y&�1�r"ON���eӱ}��$_�83*��"ObM��ʂqZZ�I�M��:j� �"O�� �Ө>lU) KO��xh�"O��J$�D�|4��ዃc���"O�F�5�H��AΞ??�* h�"O���a�� r��ք�n��Yr�"Ob!���5�n���I8:��pT"O�:1�H_ HLJ�C�1־��b"O� <�ci�xdj�D�=�0�R�"O,Zvɟ�2�jI�֤^�_ZY��"O�t#�MŊx�1�q�˦k܈"O�@�0�ءPb���F��r ��"O�d`W M�#Z� r��cu@P@W"OT�rʙ����Z���j���X'*O� �D�����+��CE.���'�����K��F�X
�e�1<�T�	�'�er�m%�*�9�j�:
�q	�'���a��$S�����_ &~!�'GzE(����v���"g)Ա頭Q
�'�8�r�
U�P�2��qa���R2
�'��%Q�y{�<cc�X��	�'oʙ�"/$(~�<X��A�#���A	�'1�|	�)ߠ|	�,jܫ%�$�I	�'��4Η�eJ�kq&wL����'���j�)��7�~0(�.b�ޘ��"O�%PΙ��P��A�:s�BD�""O�͙��Eu�������p<��"O�4i#��� "�0eJ�,6�)�"O ��Q�H:*z�Jq��O� �x�"O�Aq/Ӣ9�t�6�K�5��ˡ"O��[� I�&�v��%������P�"O�5[ROIJi������+Є�y.ȏf��\JS�P�c�f08� C;�y"Ș�~�L��f^�:U��Z��y)��6�HDѓ��($b�R��
�yR��i�aa��M�����y��w{�̻2��E�|�6ꓥ�y�H�=6|�p��1h|�ƦZ
�y2��#�La��C+I����*�y� b�Hdi��}�D���yrfìS����M�(��x��O��y"1��\#��&�.@"" ���y���9E��{�fB�nV������y���Z|�u����r��{�-�<�yR,��k�|	B���v���p� �y�+��!Ѫ4B��~�H�Ϛ4�y2mݣ(�$�2"H�j�`w����yb�e�LA��eֻ~F2@��(���y�Ŷ)��}�1�R���}(��� �y2fZ��L{�E����Y3�T0�y�eG�@���bj|��T���L��y�K]�,߄�:B�L�D�<܁$���yM�.m-��CQo�6:}Ĭ�$�؋�y�G�d�<�GK�L7l����y�/~7Du:V+�
��d !�Л�yb��.��(�!Y�y��}��jF�y.����s|�*-)c��+�y����BbQ p��29kā( ���yR�E����1�c3�%PJ�5�yR�*&2��q-�[�<�w��y�)V�RS�+��WXJ',Վ�y�ޠ8�i���p��1�#���y�C�8�`����أ=���b�@�y�狂rF��:6���5���҂P9�y��<m��U�R%���,F�y 9���Ό�%��|Ҁԇ�yr�Y�C��8֨��.�*k��ז�yR�N
2����G��3q��(�.�-�y��[�b�M�1�[�E�d�(��y"�M�7�������<~��MJ,�y���1*�H"�B�)
B}�r��<p�	���H�S��y2D�#V�h�s�!�q�°�y
� ,�{��=���qc\PJE�g�'���#Aڸ6a|��,H�t��T>j�A�-Y��=���ͺ+R�=�w��O���՗}ɦ\�5�Oc? ���"O� +n�5T�00"�!. 쬒���	8��3�lD��h���PI�� �����`�6:����"O�,8�T�VC4qrƀ��O����K�eRPQe3}�E!�g}�%˂r��+�B�`�4:Qb�$�y2�a9�l�-\�H1�[����o�ڄ��E��+�{�g�?#L�q�h]�F@���@��=ن��D.�=��@�O�ȩ�c��H�(�3�ș�'"r�0&"O��r�)G�Pcn`{`��N��Q�d�8Lv<�
A��h�,��抍�!��e�a�
14����"O�
 D�/u5K͞u5�$$���(R*׻��?'�>�C��Rd��?q�(�ZW�R�]
f��f|ƽx�Қ)^!�A��$��P���V�*��"�Ub�P#w/ �M�	���Ϳ�����/�0>��%g7~��;����+���!���$*1�C��=���U?=\4����'
��xS�"O	Q5��x � h��Ow�5X�"O� ��S�[y$��7�ˈv
��Zb"O`�Sf@ªs;.�h@�J��""O�E��C�t�dh����X��"Ob�HT��'�z��f*X�jHa(�"O��ۄcS�LV��㷇K:z<P"O� KViښ7e�Vކ0ؒ�"O l�$a��HeIG�TXReS&"Odl��Y����!��"oN�ܣ�cF:]�}��{��9O6,w�S.:�2l�cL�&�P("O�P�P��4m.�Ց��I�6�ȆM�O���mſ80Z����#%��l�dS�^�V9h��+x1a{��+�,SUoF۟��5i��6#�H{7���l�2�rB&D���*E�<,�r�IQ2�Ѕ�$�ɔN&dIh�oɫ6Z�>��N�D�f��Ab��c�"��6%<D���-�+�H�h�e�9I��0k��?5�z��+L�$Ax���d(:J8Y�OD�_�1���X*�!��k*��ۦBB
%LDX��Ɗx��F�Ŕz�Jx�I����%��u��*À#�L��
3lOVq �ğ��Nu
��r���䂴Q�� ��m�'k�>��ȓy���QN�#(�T)�d�\x���>Ɂ��/��iG�&�'7O�Ub3��}�x}���F�q���ȓ���e@��l������!� ]�Q��(X n �N�F��OTa��MK�TU����:_&�`�
O�����Z��\��]�lgd��Wᑐ�\x�
���Э��>��T�CTR�@��^�_�FD��	6�r��JD�%��
$�O��Χ$J����&�}�0"O�Y����'1�r�ᄶ@)��*F�O>�I��ݡ �b���<�'u�$��6%�Qɰ������t��9��$t�qn�O��dZGD
�}��޷d��԰vFL�����/��5S�FG�5f0c>)S���7d����ɘ�)�!��P׆ܦL�|��s�N,�4�G����RL��6��\�RMI}�P�J�6��Ě(n�\�s���AQp�N?��'P�����J5qJ�	��f>@8Ab�L�O����!A�n耜C�($9�v����uY��*^��I�^�x���ՔMH�1!"�~�#ܔ9��4("�I�'�B%sC�<�b4���
7����ĊԳ4s4i�é��X�Si����IO%��'l������d���5{�-�f�I�L�0�P�K�FX��2q��\Oః��Śec��#�*M+�8�uD�9}�@�6f�>Q�а�'x���'(�X�z��/7�嘖d�-�|ٛѬL�=����
ߓ��ܹ�(Ȩ/;�͠F�R(�����	z����k��=�>�R�骟��s��Z ��1�T�MU�'>�@�3nr�P�r�W��\p�f�.JVt�Q���ʏ9�
�PE���=ح���Y�S�`(T�G�ן
� ���FUv�{FB��||j剐�O�$�2\1"���*`�F��i3SH�W�H� �b�RV�j�x-�a��pD"]>Aʕ��m�9B�O��	�+�6X&D���3bȼ�3����Y��´��>�$d5�����4lZ`M�ClI˟XӠ����U���8����,Ov��IF�Z
t��J���8ţr.N5d��{��=)��HsVƸ[����ý (���,O�u�,tQ��Ȋ;�@�Q�+�'.H��)� ��٬	�e��듇TT0���
g4j$	FBs�O�>XF)�s���S �'�H��'�Xĉ�P�8�8��'�t�8֪Ŝh̓�{���'`�	A�D;N�v��B#�<j��x[�'�XM1V ރo��8Pb`^�|zՉ�'�\���<����A���I+�'b\���ɗq�^U�����'��MҠjC-"?�L�c�S=D�%0�'�����*]V��r/�0�0q��'e��c�T�h��I��d�)P����'�:|[��*������LP�'�d!�BO����Fˊr��)
�'(�����l�$�W(j�&�	�'��ըD
����!K�� c�:`b	�'*�\�!�?'Ǣ1�4^غ�	�'Bڽ:�n4�P	d
Qj�8	�'���
�E�r0$��KIF~��'g*����8N����*�
B�h��'��5 ��m_�,8����i�R��	�'Ƅ�p��J�((�LQ�<��I��'_J���%ͰY.����P�|Yq�'|����/F/D�<)�3䊗I�z,��'�Je����MY�d(D�ۍF�r�'�م
Ns��x�`˴��I��tP�Qx�FW R�H�*w+;SN`ZueI�-��B�I�X!�#�MW5==6 ( fK���">�1��!r�ᢎ�d_�ERVxS��(��ș�� �y��4�x����E(\�t�(��
�?	+W�;JP��o'}��	
v�����+0 "�K���!��C�	,H�b� (��Xd0ʈ^G�˓U�n���`* v|��Ă�+FY�#l
��X�	��ýQ��}�D�T�4��A�C����bI�0r�Lq"݃S��4��KD��E�&Z�R��/�$@.�D{�b�T��Q��)s�'*<�lK%(
�/��I9��n� �b���� $����Iʸk��D���Xt�y"+�X����N��D����V�¡��j��{hr�P�ЛaxNM�T�^�S��|�MWn����"*.����	=��D���@��p����<��#�4kXӇC
����zy_6/Nh���^��?���'G�Y9�Y����&t�QYW`�+N 9�K5YY!�d�!y���CE��U�$���	�^�O�%��	�#��*��O�y�,$��0FIr%(��jbDq�ϖ�8���ӱ L1K `D�5'���E���^��E�H�AS��[�x➤E���צ�8�S��	f���Oյ��O&0�$o��I*�M|z��O�`�x0P2,�)�P�[�^�<��Y�N�ȁgF�Pkb��t��Tyb�ǟ�Z���Sm��S�i�$����V�+ -J�]�\��B�	&��0ӉJ�MA����aZX�pI�D�c�B�'�*�%?�(
�cސd�����ItX�1�M?�O�!"��^)H�Qb��R�%�<��c8COȉ�������?�$ܕput43��7$�	���p�����;��%��y�eRd:��[@)�Q5��� "D�Qb�̜R��;�NA-:��x��%}bF�7Xp\�=�:I�������ٽeE��D_Y�<��dJ�E����G�N�m�*@B�,Lr�<�s-ߊ��eHV�-.R.�����a�<����%<��ЦAT(�R��v�X�<A�! �}[��;#e֨l��SJPX�<�w��n�� *@�Qʃ!c�<��iá�%f^�8|"	ЧD�-&4$B�I�h�tĺu@�< \F��w��K.LB�I�j6ꔊ��B��Qa�aʴ5�B�I�7\\e�󣊒 Ɇݒ��H&$��B�	�Q�:�)xl��4H�5`s�C�I�iM�ȸ�d
 ̤��w��@��B�)� l�#$J5%(Z����>\�9�"O���c���el씁�FI�UЊ,RR"O���SJ�bjp���.�+"O�͘W�$T����^!!'�\�W"O�@Y��8n��eڠJg*��@"OT��F).@�OjŒ�"O���!�9A���J
M%"O����VY�މ8�kӸ*�����"O��c�	c������7��93'"O�DX�	H�y��Y�ȿewr���"Op��c���6Y>���OV8-""O�<h��H�J9�ě���5H�,X�"O�?����bhĮC�� C"OVt�V��r� �@R(�x��	��"OBy��)+���[��dX�e"O�"��n�$�Ó�@���]b�"O4]�3酆h��Da�怜U�D�K%"O��Q��,4�A�B�,����"O��ڐ"�D�TZw��+q�ҭ��"OXM�Uo܏d�F�i�;x*lC�"OzEcG(A jlX�f�9a�Hq"O|)֣RH�&�s$EV&Q�Ip"O�$"���>=���ㅅ�)H��[5"O�q
Ƙ˨�SF@�<��B"O��U�RfT�ņ����f"O� xrʘ	=�"PJ#c���� �&"O�Ǌ#��a�D5�b9�P"O�y��C9}n��Pd�_>~��3�"OԵ+ÉֳeG�%Zơ�*GQ$(
b"O����I�. ����_�F_���"O�԰ +UGh�J�W�Y�U+"O���h�$j���D��G���"O����ܜn�X1�B 7(��qi�"Oʰ�DK�e�.y\ �@���y��q?&ec%�qƢ"�ć+�y�"�������1gpBd��yB�ǉ[R�;��V�P���i��� �yNʇ>�8xPo���ea��͕�y�@H  �(���O��1��`����O�=����t�¥B��q[����"Of���I<Zk||+���)t#HT�p"O����(Ȏ{��)�"%_tj1"O�Ir�����P�fX/>`!"O�qQ�#w�R�����1"O�퀖�����g��K,)$�'J͢��i�kq�
�*��d�C��-|A)�{r��?��O�O�.���5Q{`�2���*�
 ɒ}� Ԧ����* �,�ɘ�Qz�9OR�ğ z� ����$�4 Q� V�왫�`�zL�'r�<�z�@�fŴ'f�H��#�{�05�%��$n�'��e�S�O3t��p�+Q�Q�0���Y�
ѪM<�rA~��E�O�F�q���<0U��k�X�L)��O慈��_z��&�"}�D��I��E�θO �#"�ۤM��l�ܴ"����Oa�� Z�2���F�j�x�#D�u��"�h޾���V�@G��Z�9�Z��@�	`� �z�n�<Ϩ���'ռ��+.'��K|���͙22�d��	7�r�aa�_"UiqOⴸ��*�(O���)|��Aeh�	[4쉀�Ggۖ�ҧ�]�$��M�n>ɫ�*��� ��~��hP!�<j����k��2��6�B�( �~�H?�X �@���f���6�Ƒ�a�	�aͮ���&���a�4#��u���3i �u ����L؇2����'��ч�7e�<褟b?	B���v��kpB��D�X��3b�>�7�ö!bע���zөJ��aH�Y/\��M�7�(59��Z�ǂ���b��M���ӣ��4��@o�����ۚOu�y���F	�l���J�|��	>'6H����)�d)��i(�r �+~Ҋ�ʂ�A���'��Ʌ%�4�ϸ'q�E
�,O���Gks�J�.�yrdI��(��!i�H8�����y
� V�8r�F?Yr�=G�@�5���v"O	�X�!A|�0G¹bv4(�"O�S�P#[2p���_=B`x�Qd"O�;!��i�� �%��"(�0KF"O��kJ�=a� 9��@�v,!�%"ONl����;��)Ⲯ�!`	t�sf"OX���D\F?�US�B��l����"O������D�V���盤�l�x�"O���e�����z� &�(3"O��(0 O��f�) ��V�2��4"O-+
G� (�Aw
Z�]�}�Q"O��h���F��hh_;P�В"Ofi0T��(k�(��T'�uK�A2�"O���!a� |����猁	Z�-A�"O������]����åU9f�{�"OT��BB�F�֡:�F��]�2	�"O|y"T�Y's!���&�L+��4"O�E��nDM=x�abc_��-�"O�0��-]}P1����C��j5"Ol]�u�A�q�X���]�N���k�"OX=�F��C�3w㛿4����"OrL��P2-��D�`�;�,T�a"O��&f� bf��A 8G��k@"O�y�Ղ[/y� Y0D��}�h��B"OT� ��:�"r�C��Ph�"O�3'� c�����ԋ
⪍�"O�D�� Ʊ\>�S`�=پ�"O�D8���$e��7�)&�$�h&"O
���D��������{E�ڇ"OJ�(�a��'	�D�0,ש4$C"O��v���8�c'KZ�3�j��#"O��f؞?K�C��D֚@�A"OB�ȍ2.�tp�
� 2��y�"O�e�kDn�!������(!6"O�u*Fa�/��y��S�a���7"O���`�8@�6�E%����"O�@PB�7;���l؀l��I �"O�!bv��.j�4�2k�"d�c"O�q9�-Fc0I�1/\��9g"O�a�I�[�Ќ+�#I�1� ��"O\)f Ha�];4�ϓ ��m�"Ol|Q�ʉ%���%��Rx�m�"O:���Y�#Z���S�a�!J�"O"�P�k� �&�[�+Y�ZH(E�"O�g� �������2�a "O�9��X�Iô�P����6=v@ȡ"O(=+����Q`D507]�q"OP|��h�PyV�eh͐3�]k�"O����'R�D��d�t���'(�Q�"O�����:V���@#F�7i���#"O(0Ȱhտ/��k�[�l�����"Oܠ��*Q�R^؀�D:A$��#"O�ar��B;{��!�e�<��9�"Ob�1�h';�<Y����C\4ia"ORY��N�\�8��ۙuT��E"O"�B֩������Z���mkF"O���+&����%U�+��]y�"O�	k�3�M#���'j�=q"O��3v���ts4��$qefm�W"OP�h�)�,b"DpE�:VG�y�"O t{-���%�Ҡ�m�
h�u"Oz��V%*z���J�$p�>9j"Oz��쐺A�2���h�5X#N��!"Oba�ƋS"3�b��GH׽r���"O� f1��%(��1��E(� !�"O�䚐�ьr��	gƷO��AQ"O�2 �$
�$�IĈ�,��"O��Ď$F��q֡C�
3�c "O.�tJ�a 0RKP v��Xe"OF]�q*/O�e�@��̉�"O��k����ǆ�9�(ehE"O�$J�`1[�t��g���3�赃T"OX(��h��Z�H\��A�.�*<�"O���p�āشYH�]�J�1R"OƬ	M�!%Tqᑋ��s�"O�"�K�{根���W!\rJ��r"O��#��̶(sj)�%G�mf���"O�����0�pad�ܰXR2���"Oڄ1�`�Qk�tTکZ�8"Ot�h��I�,���x�̉btT��"Or�C��B�g���У�"mI�3"O��%�1�i�P"�zl���"O���WH���yJ�k�[O$H�0"O��S�.ςn��p�!I*���"O��"��E�/��I�q@�8D�`ڴ"OJ��w���u(e@�#M*�Q0"O2{B�G[�"���S��M`�"O�� ���C�\|k�-��9 �"Ob��%+�*i3&�I��D��ڔQ"O��ȅ�*mlq爞�\� ��C"O����. �#J���XA[�"O���*�+��qóe%c*V���"OdU6*׎N��i�6"�c<tm1"O0�ш�hM�8�U�׬'PZ�"O���ŋo!�0pbD����zP"O�C��}����p�߹r׸Y�"O���׌ͰL3�����b��h"Of	�A�W�G�������!]y�|K�"O��Q�΀#oj�Y̜҇�] �zD"O�����5�f��w+�'r�4�iW"O0՛�	G��(\�f� @��8�"ObuSQ��W�Ĩ̀Kb}S�"Or��!�y��	2��(Z�5��"Oµh"}�꠩#c]V�6-��"O�8�厅'A��`�Á���0u"O��ЈI�Qov�҅����S�"O����g9V���4ċ�.2����"OD١e�1l<v9���D%%^�;"O���i�!�*��$̯,3��:"OBգ����8y@$;	v 5SD"O�JG�?%/�B��2N9��J!"O �h�$Xj�� �ee��K��1�0"Oh{Ah�4t�0E��B�vH<��s"O"���5��욳��'�����"O�+��#c(�9�s�̝C�`�B�"On�P�Ϫ����B�k�d)r"OB�3���3���X���&hȠ�"O�Aa�a<Xv�ie��m�]��"Odd �εTM�ठ8B9Ѐ�"Ora��/�й���X)���7"O��ӵ�I�a�X���Ɔ]R�x�"O�̙�d�f62�%D�@z���s"OJ�s�� �Y��aI�֯Ex̵�a"O6D��P�b}�l9�͙wԸX�"OVS�O�!�R�1�f��(��L��"O:i��䙅�4��c�Q�}�VMC�"O�˥L���J�f[;ou64Q�"O�(�p-Β]�<ԅ;t}
<S�"O� �S6gN�Q�^X�e�M�(X�"O��1r�8^���w�n&
���"O�X�$Bd����?wA�d�R"O��ի�Ss��	��E0 O�`��"OX��jG%���\�B��h�"O���4+��d�dQb� ��_tl8�"O>L�$N6cl�Cs��1܈�"O���5L�.@���鲍K ���)�"OH	Z`n�cX.�[�ꀆ`-�B�"O��M�uj�Đ�β1����"O@e�%��j�>4*dF
i\��7"O�B�a��j��t����e�L�Q"O0 FL����+eC_=%k|\��"O��P�lO0"�5 #� �h	 `"O�dA+F�x��4�VT�"O�ycl��C�a ��3�b��"O��ڵ�J�3`�E@��-C���"Of9��G��<����=G"A�G"O�8�Pϝ� ��ipn�F�|�a""O�`�Ua���@C̈́��8��"Ob0�j
(5[F����(s��Z
�'%>�ys�٩j�A�?0��Yx�'���R$^��05�L�YsP���'s�t�G�� N�6�w��XRn�y�'��|c3�4b����0�\�XɸH[�'P�m[D �$T� ���[W�D=��'+��؇'�A�xY�ʜQ���#�'Jmf�[��=R���>��Q�	�'{Z�c^'W���:QǼd
$(X
�'Q,А�ٚ��A�ȡbO�2�'R
C��5W��iK! D`�8��
�'J��@���$Hh����H��P��'&��A�Q7 �pm�s;���
�'Ƽٸd�1}L���(M�`�fY�	�'����� ݜj�R�駍� Y"�Pz�'&4L����/"դ�W�[+X��y��͕9!��h�O\r��Y �D�yR.ّ\�� .Ykh�Hx�Y8�y"k�z��C�Ů`�l��AiĊ�y�[*>L0Ѕb�Y��\S!ė��y/J�1�d�a��~ڐ,�@���yR��vЩ��Yc�(������y2mOOL	{4�9_���PM�y�N�,���3�㚼^x
����yZX��`
�� \
҆l�I��I�'1fy�r�&1[����Nx!Zy�'���5�O���ehr&�e	h���'�x2Ô�/��uoE�nS ��'�|l�!���A,Q���:n��p�'_ذ�c��n�xw� f�l�
�'������,JX��q!�X֮�{	�'O��:�GY�g��*q��b0\ĳ�'آM@�L��Sp��7�V혴+�'}t5���[�ɜLi��m1��'ղ�G�1d�����!gꌱ�'�¸G"��'H:����Y�>�i�'caK��ͧ3/2���+y2X��'��!G.�R����u�΀_���A�'��R��)g<2a�	O܀��'M^]��(� z�zYSw�\=@�0��'�B`���M�"�G�;D��b�'q�%��H�{�IA�b��.�Ȑ��'�p9Y�ê��%� �̉qP��'rհ1g��!q@�7��%]��p��� Ψp�陀�9��LK;�N@��"O�%�S�4Ejm0P�_%Qc�@"�"O�i���B"S�����&>T"D[�"O���5   �P   �
  �  X  �!  �(  1  Y7  �=  �C  1J  sP  �V  	]  Qc  �i  �o  v  ^|  j�   `� u�	����Zv)C�'ll\�0�Ez+�'N�Dl���32O$����' �
�eřq��退툅f�P��r�ޖ)�xR�h��

��@еh*���c�Q*w�W�?%��l��?�C�NǐM��8�M�Du>!Q��]�oy$`��l�=s.�ە���+b�Y�$����u�B�7~v���'@jG
���2 ����33X���X!c�\X1��O̔��lJ>�r���$Z��e����՟\�IݟT�IşxA"K*��8��
V�pՓ�#�џ��I��M#!�����O���e��b�dj����M�3dv�����L�\�5j�O��˴�<y�w�����'jLM���<��'	E<�1���]� �����O�x����/��M�bfˁG����X5�ș`"HP���F�'����\t"��ʟf���(X�1ɲCM>oB!$�'i��''��'�"�'�BQ>�ϻ#����e��IN6l�5J�r��I�M#a�iv7�Z��}�	��M�#HɆ�����b�ˠ42��ciC1o(xYn��E��"=����+�"��#�´o�<-�ح��+��L9�g!�/H�V�o	�MK��i5�4���r�R�\1����D�z���9�/^���)�'PN��M��#(� �5�"B��`�F:zP�e2�h�Vo �M�B�MV����=zF��H�OV���0``nט�n�c�i��7-U��Q��kL�{2�Q�PeG�T�:�s���4�V�	�` #iڌ�E��/R���9�i�' ��2�H��M;`�i��7���yv$�!|̎\�d��F��a�� U,C�-Bt�-�|P����I0B�k�E�\�y�����$��v	dȓѮM�)�L�B5b�i���D6�	ߟH�I��^���4��i"C��1�.��<e�U��O"U���	���ͧ����|�����&�ǟ���Hg��t)]�ZI�T�A�L30�ܼx���ٕM����m�	@��i��̃����v/�2	��xp��$��2U��'@(�g���@�6z��p"o̵o-�@�	�0��K�S�'�yb����N�I��5��T?��'�ў�S��M���ϐ9��ۢ
*7.h隒��6���DR�A��⟴�'��$c I�/N�=�D�p�]�ȓ&hm�N��N�-m�(6�� ��'?����w�~<���0��#�'�t%�#�4s8M� ��y�Ա�'�����i�6Fr�@a�4[����'�"H��FU�#cr��k��L�!
����Gx��I�2��L�c���!7li��P�\C�	($�b��E���f�6 ۺj� C��l��;1�T�v|*���Pz�C�<r�j$�KӳVɢ�����<��C��
;��O�Py�,���C�&tcؘ!�FI��t��n��:���Qo�ky��'j2W�`�O�	&�|q���_/d��+�A	y�<<2Qd(l��Q V�uxaz�� ��X�!M�/sa�p���N��Q��&�>)3���-��@���-�ў�[�̰
Q�B��[.V��D@M�M����F����ī<��Ov#eM�<n$5���~Sd�+3�'��y��A)n�.�;�O��1�eJ�b2�c�V���uߴ���0�o�ן�͓PE��]�t���/��/&���eyR�'��5�^�4�S�	�����4)r(\%KZ��J/2�]��
�7Wax�E��Y���/9N�L��5����īL9p���#լ��|��- ;� GyB�	2�?�ֳiu�7m�O��P�e�I�x�PN��T��Yar�<�����(�̰ؕ�3hm�dx!k�:G8�f���O$�}j��i���y�;����TH�c-���&|Ӛ�Of �q-��Fp�㟸��0,�@��\\p&E��,K
:~b8��"\��1GE0@	�i�� ryd D�<zQJZ�/�`���]�Z0z�a<D��:p��-W�����d\���R�6D����8E�<R�$ͱ57����$4D�`"@D�s� $[�-Μ]_*4�'
���$���a���?��IğD�	Ky"������.�	zU5ZC�B�YwjyQ�IQ�v�B�:0��	vU>�GxRJ��AM�1  $�:�~A ����\I0��U�37 ����T~J��ԭY�gn����l>(\�cC��+̌i���^��^ ��42��-�L��%��OT���OhhP1�[�1H�X�h�-�tmX#.<OJ�?�v(��r��$L4:�B7�ןX����M��i�ɧ��O��	yj�٪5䍉i�|*��= 0X1���-�M��?�����%��J%��E{�ޞ1cƴ�tJY�cN����խ.&mYa@@0y�Z��ܖ'��h�f�Aq L�;i�6��/̖F�sgV0�TlnڮH�2Q��剅��$2���Rr4�a�'�;�� � �OD�ncy��'O��'���'����Wl�};��$r�(�p�Z4b����7�I�<v��
"�Z�g�I	�b�W�~�O��n��'�T}�U�u�`��O��4c#�������S�XBń�O���E���$�O(�Ӳ!�r��-�)� ^@��-�kIR�;&��gdV�:#�'^��j��d�6]�]Q �_�{Wp5;�GG&!8ax�h��?�'�|��5���Ҩs*� F���y�#\*�DȢG��fJ��P����?�v�'��Po��+�p�rE���eL�K>�vj��aM���'TRQ>�c�gߟPX�+$y���':Z��ծ�ޟ��I+[R���m�S�L���@	�9I�:0e�OA�Bu�!K,?Y�L�F�����+�G'���V 3v�ŠԔ�$����O��'�"|r'&�.x�`a��,��"�N�<Q"�B�l�$02���?*V,j�v�'L�}uᛙ/�x�Ӳc�8W
Y�B��M���?�:��9�w%�7�?��?!��y��Y���G��\b}���_��t����?��[�+��q�,�Q��B�*ߓΎ�r���)���C+�3T��H�O��h��cf1�1O(1���y{.��r�΅t.��c�r�p�n�ޟ��c!˟h�T��,O���OC�$��l6.�<���8]h@�$�-V7�㟴��w�'i��O��uKxq8�J���.����?�@[��'k�O2X��Z����(���(=9�\8�#Y�Q����a˟��	͟��	��u�'�R�'��� �!�&!�0!IC�`�Ś�-��%�R�aE��T��tp��'�1)!�Hj�S��]� ���Gc�L�����̔x���	Y���CgACx�'2�㧯��P��|T���Q�:��#	7�?IP�i��b�$��l�'B�XJnßJis�*��-�������?�L~��y�		`���,�?{F�H;�D&��D�O�n�ٟ��'9�%lw���d�O�`���I�D�JD���&yDt��`�O���P�e�F���O����r�ҕXJ�&���"�`�e�p+üQ�f�����0�hA��%-OdK�-��vfH��/�9��m�=�]k���V�{��u]�ƒ(FQ��j� �Oz���ʦ)�	�e<��v�/�فE*oE��?q��O|1O��
Cf��u��MV���$��œ[���	ݟt�?�ON&�$��V`T��6�#Y�U�TO�7o
�Q�X�� Q��M��?9����(���?Y���a�6	�Cl��*��+�Ŷ�?�6�HH����>9t è�b���g���ȉdHS~��?�O>��`�H�B��A2_��H���3?yG$�hH>E�t� ��r�ߖ��yYҷ�yB���*�^�+����B`�"k4��OTD�4-Y�x>� ���Pzi9����WћF�|B)me���'��'U�	�h:r zn�6���,G6"x����l���)��l؂Ŏo���d7x��� �H�GI�P���`Ll}d�$X`9���yR`F�~� �?b]�L�IS�F��d�F��%���$T���gy��w�����8�,}���F��К��'&~p��D���#<Y�-�(�Ÿ�-W��A�ȅ矌��3��į<��������d�$Ѐ[�B��9��yj��N�D$��S#�������P��`yV>��'1�xX���q/l=��/O���Z�(��Ĺ��I�q^v�ytk��x~�a�&%r�0�$���t�摠��Z�r�Q�d�Nj�'�]�t��o0��נW�m�d ��N2�?)��3���'�����?)A�φ1���f�=_��Y�#����D:��ǘ'ba�fK�=��e!%N�!Tb��O>R��!7s��W���d��uG�'���̲p��uRwB�7\�pb�`B;j��Y�D��ßL�ɣ]���/ʍ6Ԓ��CH�<�!۩?��E��:��G��p����f�1*׌�؇�ҥnH͈�0tM�e��I�	����BO#ZbV�F��N �?�v�i{��'Ǣ�
6���Z��D�i]&\�b�'B�'O��'��OV1O�h��*G;>�TЖbPCD�x�5��.��|b��'���C�YV�d�G��*�H�����:qH�l�b���|��4�?����r�pCë�7�(M��oŜ�?���<�@`���c�VX�G��?�����#>��	�G`��K�>s�I� EX�IP>�+��ʚ�(����,+h��x�DEh�U�tg�\~Ү���?�S�i�6M�Oj"|RQ�3Q*� �lG:��
�+J[�I��t��Z����=Z�D�i���f�P�)dl��hO\�d��u��4��UM�|�B��&�F����h3�����WkґY���(O,t��<?�P���e@!�:��&"O���q�\�OV d�w�� �Dk"O,�&Ƽ~��-�7�J�~D h�"On�rM	"ZJ� &!u��	�"OB�	�+w�L�%��v��p��"OX@�1�V�ԁ�S%�Xp�T�Ш�/�O��Y0.�Oa�13��� �uY�"O� $�JD��B|(DT�Ϛy�@"O�ze�^2-�Hh�P"ƺ���G"O�Qc�	ݠ��Kw��b��s"OP�����tɚ���oB�?�J�7�']���'~>XR��Z&U�bM��_�h)q�'k(Ajw+�	�>���%l�аJ�'g8�����( _��2�ß_����'x|�y��U�s4�M1' d��'G�eH�ȟ��軴���p4.Ƞ�'5�X���X�(I���a��1���ą�W�Q?��
4$�h����Br@� 9D�زPk�'F�,�Ҩ��?��q�:D����i��R�����	�!^�9Ԏ7D�\JrG�f ~��0+Ȭ[��3�B8D�Dbf`�8�ґ{w
�$Q"�ل 3D�l*A'I�@U2����!:
<�Dg�Ol���)�$W���">E�,��bk��Qq`-�	�'���B7���b�����JME�	�'Q���f����4D�!�L�	�':^��$�7�U�\U$%x�'of�p�H�"e(smK<O��y��'���X�Aߔc_| ��x�Z�a.Op�
��'*�$���^_�1[��'2�i�'�*h�6��,L/QI���{T��'�b!���,E������/�xi�'`(�j��	A���Q8Bx��	�'��؀U(�"��YA3��6+��Ā
�T`9�3���Ȧ`@���p����3�t����Y�� ɱ
J�Y�(V�r�����ȱ�2&�d�X�EV�ܾ��ȓnR9BĆ44��T�%�3���ȓaڞ��я�2��u�"/�1\��5�ȓw'V� �K�,U��H/&}��G{� 6�����I	��D[��i2eC	�T�1�"O�`��"��-��
�cԹ.��t�"O	�քL�n�u�T��8;���`�"OrT��+� ��]Cb$H(���"O�=�D�X�n�*jVCV�{����"O���L8%�j̹�b��m�<�ȕ�'q6y����#9U��r#X�t�j��
�1��Յ�U����e��;��˶䖅/ez�ȓG��)`@�Z�
�*�� ���Z���5��[�G�d�n� �C��]�l��d4d	A+� �9@���Jv*$�ȓ/P\!�C��j˸i�L�|8(H�'�T�	�k<1E���5o�UQ�l�{��y�ȓm^�LS�n��8���0��}{�ԅ��T�!G�V�3���0b�Z��Ѕ�\庅h��F�PՊu/B�FP"��ȓnVrHR����;��]���raƕ��	��8�	�&	j�cjK(�����Cs�B��) H<�u*��l�΄��F?�rC�	�y[,p�j�N��(Q�Ϡ2�`C�ݤ�+4m^�w����M�+a^C�ɖIIBU dذa�j�G�X30C�I� N�d�9EF����T�=�#�Wy�O�ԉ�/҆nj6t��mZ�Fl�'�����э��Mt.mS�"O�,s�D"$܈aąi���'"OΕ�䬚���bԆ@,Y�޸��"O^!�"ȅ�HYRՂ\3�
�f"Oz�§����<9���m�8s�'���p���e� ��r�N���0��E�a��h�ȓ\�n2���H#�)�ƛ�F����S�? �b�ϯS���3�͘V�Zhpw"O��K��"i�ܓ��P�c�Q"OR��6�\3S��-h���`!c!"Ov�we��9�
�N�2p�t��FZ��ЗC$�O� ��E�SQ���歁�4�Vٕ"OH�0��6w�Yy�
�!>s�Q4"ONY� �����E#X�T<�P`"O�� �Y]�i[�l��6\�"O����OJ�� i�S&�R{^���'���j�'�r�:��T�١��9v.�q�'޵�e�]	͜U�A�Z9R ���'���R��s�L��#Ő(vv<�t"O�q���?	/��a1�3=gb�)#"OHD�4��6p�M�e�@�u2j�"O�q�v�}�Y	Q!�48��0�e�I>
#B�~�n
$H��a[�P �	z��b�<��j��*{�$W�:�^��Tj�<1`M�����"N�X�.�N�<)��m���s1jؖ:P�á@J�<��
C44 ��0i�[aU3�$�D�<���$��"�H�Dbhq��I����b#�S�O��aH���Jl40E�І,C�Y;�"O̘���[�%9�s�L�:4�S2"O�����H�#8̐��ʶ%|��C"O�q�)D>5�H����Cj��i�"O%c� �BN�m	��J#_�l��"Od�����]���Y�$R�x�]���T�"�Otٓ�d���Cc«UОx�4"OD�A��IlӶ(�F����"O�����ͯq��$#�E�(l	ja"O�T*Vi�\��<h₄�H��ܑ�"O���h�`\�X�O(<�&�u�'G��K�'h�U{�K2* �'��M
�j�'Q�C��& ��VDE6dH�'#�l��3/�2��E$�>��i"
�'�Y���O��ܺ�� 87:��
�'��2�Y�yI�W7@u�U�	�'6�yv/�,G����s���7��̠��dY�H�Q?Uh�F�`(\�g�K�~�ۂ�?D�8�`E���)���E�a0B�k+D�`�s���dy��e_�-3��f�.D�3�g�?@�Z���"�<i$�I�	.D��H��X:vQH�&I	���(��,D�<ʗE��s6=���œ8���s �O
���)�'=X�8i�׽�6ds@mN%"��1h�'2$�1cc�3�J��gJ��e֦D8
�'~����LTDF��gM*J���	�'��qx�d�)'|#�I�l�jE2	�'�fԢrK#utV�A#�������'R��*al@*P���hs�6MV|$�/O��Q��'��x#�&ӚNѠ͸��Z+L�Bt��'%X�Ar!љQa4��G�[����'�x�"3�Ȇ	<F��WG�'!��b�'���.P�NY��+���p�����'0`�5`ߩ_2ܩɖ���\Dm��#庐��qx���"Y�L��Y#3���[��$�ȓ'����`ҡX`���Q�ԝ�ȓ4����DD�a�43�U���������9�rYS/Ͽzn��ȓ<������t���Ґ��\P����>�H�iC���ej!����<E{k����@K?p�D]����=���G"O����&<�̤x%���*�ZIa"O�$����@\B�2�V�q^��"O� "����ܵY 2��4@Q�R�za"O���W!R�3,�R��҆NQ���"O 4�îK\�\�c��=���"�'D�:����U�U�R��:[F��	8NɅȓ
�4��ޱzp��JPM�<-1衅ȓ2���թHU6=q�:��M�ȓu��Ɨ�n3�U 'W2jm�Մ�Z�q��lȽOmJt[�
_��@�ȓ0N�6BdG*��X�t���'�n�R�r�¸�v�G�r*|�
RϚy��ȓ:�zA�SdX�nE6ț@�c� M�ȓ,�+��u�젛Cl��	������H܂>4ĥ ۗU�^ć� �^1ya�H7T����ƍC�dJ�����+�x��zʬ!��%LRQ(y�eHM�1�nB�	�{�%P�F3;]V1����oSB�	B���S�~D܈3Ea�;=��C䉷a����1O� �D��v��B�	�-�LY��bUdb���Ť"�xB�^neC�J�!�t��f���P�=���[h�O��H�6�*G~DE�WH�g�=�ʓT���"���MV���h� :�E�ȓ%���2��p��C��Z�y@<��,��Ɓ�b���b�kʁZ<X�ȓv�u��>!P�	 �D�p�-�ȓR�Qԉˏ'���S�G?bZ��ɪ?bF#<E�DŅ�W���& PEpF��1`��I�!�D�/D�2yC1��	u�u�,�d"O���GL@3��h:�h��Z�B�
@"OT��pn,n�>-Kê��%�`��"OT,b�B�,:z����)'޹�TOP�3�#U�șh��b���t��O�1��U���o٦�+4㝽(>�dNϺk��Z�aJ-b�����ʸ6�t��Ù/�?�֦ި�?����?a��G�^6J�Ǝ+������i�.�tr%�; P��.����O�1CG��-b�r�*�%(WcW�~:xX�̈�l@��Y&���1��9�)���(O��ɦ�'r�0bU#N4e,pi�ʹX�Խ�$V� ��ɂm��es���ܹ��g��v�Ol�=�'��8-x��x��)��T�@̘8�@��H�HGN����P���*r��)Mhx��U�U.p@)��n�D�[!Ʉ�g&>�Ƨ�l���ȓ?��m���Q�hDv�%�ӓ-6B�,;P�yc�N�0p���kɃu��B�I1�4pV Jd�=qe�̋ui�B䉴HGN`���M*|<U���L(I��p��	}��~��
�]8�:�H�7M�*�����y��5
hAr�U6K�.sj�'�yg(#c�ey�Dף7����!b�)�Py�\ ~��zG!?'��x+��Ij�<�qL��`I���(n���y�%D�|�Ԃ�;tM�Th'+�7���#q$�OfA� �'M��h�KX^�Mzoū�`��'d�ɚmI�����b�	s� Z�'��0�ve�Su����3T�\B�'���4C^i=�#�˝� ���'ty⠥�8I>V�1�8"�(��ߓgp|�Oh�B�ǟ)c�l�#!�6��p�e"O\e[áI2D����À�A��f"O��k�FB�� ��@�ո���9�"O�Y��Y�X)H� �W��a�"O*1��&t�͓r�i��QҔ"Oz<�r�Y/RT�%c�M�� @�e�$ʻwC��O�6T�Z�~]j�V5{�����'��qq�㖟�b�S(�)b�d�'�H@Y� ϡ�|��'cV�aj�Q��� D��B�ͫ�ț�E�"pȂ��"O����暈Zߘ�d��<�L��"O��@��԰A.�2�c��!S:M@gP��O�}�`��a` j����� þ���`�4Zb��I9`�s�ԙrr�Ԅȓ,O� �f�Ձm�:��c�E�s� p���>Q�P��L2T$J�Ղ�!�V�E�ҵ��bL�H&��&W 	!�d�j	��Tǜ�KӦla��.G�b �p?)3iDm���!�%�,f��yt�c�<	v��a�jwcO+$�(:��y�<�` �(D�hU�v�֎[ڈ�
�v�<QBf�4P�>$���P;����-�g�<1aD<}�����V���:!��b�'�L|�V�~ӄ��O�瓭Bo��L�Z��8p`@�oa��DQ�R���O���K<u��5�i>�d+J�+��%���T>tx%���(�>���D��g���t�ՉH�\��5�K��O�����'>�?��M���%[���yD���R"-D��ha�.<�H��5�N[̔��m5�O2i�'v������zBJ���kPW��,O����OB����Ob�g�Tdx�%FG�Lٳ�R"O�,؆�k�'4ܽq�g��H��@#���6C�����iG�'���|Z�.����/� �F��~~2B����:}*���_�uv��+у׭gz���q�n��uI��7?1��>�5��p��OR⓱��S�F�DH��%[:[��	��>�U�O��}Γ)��Q�҈W�܈��T`I[>�89�K�j��T�Dˢ^��W�Ӌ�P��I>95�p���)*\���(m��z_V�F���]2&������*yMڵ�`��́����ɶ���'�J6�CJM�����0`�IC��A$��	W�<�'�p"���L�b��&�*V�l=�iɶ%��ɖ7n�S��'�@ź�OFA1!��ű���T���rȍ�\\Nȳ+OV�S���ș�O�.�b.
��n!����<S�V�����~�H����?�	.~���"J�l��dB��*�EiU�K ��dF���?Q �=�sw�I�v�Jlbua�K�<��1��d�s*nl��5�NѦ���Z�	�����Ĕ�MCF$�;�h��gA�>	��IS��P}2�|"�~b�E�"0�)e D�dh��FK�<����]�,�C��
g`�*�k�F�<��)�(u\�(dG� f�Y ��z�<ᵣ[T�=-�d��p� FN�<A$.��Yx�ȫ���8���U�<i��Λa/z�wo��v��A��S�<q��un�hFGBsk�iG MN�<Y�D M�Hd�3���z��ჷi�H�<Y��L�����m@	]%RS�_�<��BPk����W��������U"O�E����&��%7��u2�����fI0�B���\�J�H��cȆ f��qQ�.Rl!�ڭ-i$��O��p��c(9�>Y��
GK���&�0a"1Z�,�cE$��tE�#t<0��`�+o��!$LV�|���AE�"���H�L%��Gg%�0B!��y�la�$��.e%�q�I
-Zȡ�"Q#N�!"1'�!z/�����|:�����%HL�3-ExQ$'7�#�;ODz �@�M/Eb��i_=6���y�͐o�^=qu/L������O�L�%�`��k MѦ���|����0�Ë�U5���c�(@��B�x�"/ek\H�R���$��x���� <Z��"'`�DɌ�MM��TسB�R��*���d��9��ΟPE��i�Î���i
�ϯz����'��;T��:�v��#C0yXR��%��|z��ɰJwv��D���a�ݬh�,�I�l��ɹ �Fe�/�.`-�$,�@� C�ɕaa�ؓ2Γ>>6�
$b�0��C�?`�L�B��j81�7�V�NC�I)+�2<�$%�3I"�i���@S�C�I	��Mh�c�(v�T
1�q��B�ɢ�x`�	�+�D�*ݧd�.B�ɗi%�q�����e���Z�P�M�TC�)� r$hoK���W�ÂQ��L
�"O�	���?W���
�䀌za�x�"O��Wf��P�v��ՊVF��xS"O�)G�Ý0���HW�!F�}�"O��õn� �`i��ٷW/�� "O�̲ `5��`1��JOL�{""O�IK@M������LJ�XZ*�i�"O�ĉ���F�P��W���9�\SA"O���#�82�j��g�ߪ).zq�"O:(q"�L�t���4��!$(���"O��1�����p������"O���6�Z"W:��a�Ϊx�LP��"O�lR/I^�t!Y��^�(�@`A"O���d��i֩�W�חop(��V"O���;q��H@T�*Vip��5"O��A�N��$�J4�s���Y�q#�"O����e2��mɖ:�6��f"Ot�����i��A�&@&(�0��"O�d��C�"` �ي[Ϊ�(�"O�
r�J�,Sbi�p �}`j�zp"O����Ю/�~)q�ω+YL��YA"O��ԑx�r�� #�婰"O��а˧:�P����s\J"OJ���Ʃm��m[�햄_�p��#"O��Q�jנ(D�#��O�,f �"O�5�o��hT�w)!
��z�"OȜxӌ��zTt�v�Y%0��!Z�"O��A�kB�oD��q�$B�"2"Ox��bB�w�hU)��^�V��x�%"O`p�`��{��VOA�+�}�`"OruQ6�Z�@�Z��'�O�.=0e"OX�ʰ��K" ����=Y�VD��"O8�˓�V~�4��T�^�@q"O��TH�v�����ǽ��q��"OrX��@\Ȏl����%e��"O�|$k�"kge@b.�wa�Aq"O�-��$j:%��X�J�X�"ObB�.\#�B	�]�"D�Rr"O�u�eE�(@�R]��e�#��x�"O:Y��,��̠�t$P6:���*OH�*���5y^���M�Y����'���(r��.qp"�|8����'�����0(W:���	�2��
�'�`�Gǝ6;p���+[�(,���	�'���*���<3qgɎV�|���'qLS���5sF���K�Y3	�'��h:��Tx�R4��#
0�:�'�r��6�03S8hk�..8v2�'S<�{c�\�Jd��R�H�S���'��u�U�S�4|�Y"ADT=�6��'z��@�B73\�k��^�7�Ҍ�	�'��M��KU*��	��22�U�'� �d�7UY���r΃fϪ�'��\���I7�U	��˽bIxM�'�=h3k�5	�� b�@,ZP��'K^��6h/z�lVGH9?���
�'���#F#@��頰)��*/���'�.�3��?2�<�&�M?q���A�',�](S�Ƥx���� �����'|Vi��/��R�p�e�DLڥS�'�z���֗��KU*Ա��'�,�3R
2���I��
��Z�'%�,9eDD�z���*0|l�=:�'������
��h�5k�m�h@���� X}�f�޾!@PX�c*|��{7"O�!��:T��sQ�:K��u�1"Ot	�����?�聒W�߾J甸ѳ"OR�+v��~Y��� Դ��"O��#\�T���!�ڼ)�#�"O��ѥ�L7k{d����k����"O`�:P�
7L��k!��os�D�"O�����;.��yH6�]`Bܑ#"O\�yQ&�6?؅��BU:�pW"Ot �B�Z7~Ea�����/��)�"On�{��0^�"����R"O����-�1Rt���d�'O䡚�"O�H�2 �v�p$[7|�zm�""Ov�	�O�1O8�{SM;��$(w"O���7"M�yg���P��m�8]"O*ifE�]@pÀ��q�^�(�"O4}��f��E��yY1�˂]���!u"O|0�ׄZ+~�2G�F�ı)�"O��k�V��>�sD�V�xphW"O�!�B���*(����=	@�A�"O��zc���Xɺ$L���q�"O|�꠪�f+@���-
	�ru0�"OT�EA�:\z��v-��3@!S'"O.,JuNؔ�����n՘W<\ ʡ"O�Ku/	�5麸��:6�jF"OJA#��z��N^�u/<�S�"O�YkF�2(���c���i3��3"O��(d/�4���@�^�4!��S�"O�:�׌d'�$"��Ž�@b�"O�Z�l�Rq�Ɖ�;T+IE"O�Q���=d��)���*D�s"O��@o��7��&�ǐ7o
�
#"O�1vN�9��5*�a��`�I+�"O���Ǌtka�@ߧ=�,8�"O�`5�P82F�Xsv,J!-���"O�lقaJ�z9��*O�b��q�4"OzĚq�@-@�2��h̖=���2�"O��(��B�s�~�Z�F�����#"OXA�̔9vS�iH������"O�x��^;:�2�{R�M{Ɏ|��"O���
\�RB�u3B8���``"O�$[��Q�Jظ���)y�"O�e�5�I�u�RI �cY�nq.X��"Ox���n�"wo��Aw�^!oX@$��"O�A��G@�Y5t-�@O�*6��qV"O4%�#��  �e�p΁-�P��"ON%�Dm�8t�16N˗�`�ä"O�YAB6~��j��P2��A�"O�I[�h���.����c��y{�"Od�yШƳj$��`&ӑ�4��"OZ8K L[)p>v,���F �%��"O���GE�M|20��� ����7"On �U��`w8I�rBB�%�p�$"O
9"+��#�.Ik�,��$��"OL�x��×|~�Ӱ��zir��p"OpI�ޯ7*�)��ɓGƌ!u"O`|J@M�X�\:�ʇR�HЫF"O�|3d�G�@��3s隰o`�"O.���~���*GG̃7@ �"O�(�	��1��Hk���3��H�"O�l2 �0v�S֮��o�Y�"OrXy����p��L޳k�*8Re"O���uG9*rul�OO�0q"O�1� mBr��q�ڭX!&H��"O� >�{d��4�@h�ˍ�C�fQ��"O��`lAaЈs��Z'E�QC�"Ot���+3�Isr*ܪp��s�"O&��'�X���i��z�~�'U��A�G�
z�Hp�נ�
a�'c�PKt@����� y�,��'�x�sL \��<Ȳ
t-�0��'���t+J�jj0Ahb��3;��'�(H����k�jt�A	)� ���'p�(�cP]�4 �G� �ʰ��'ZD1r���r(� Q�_9`j� �'GN�qp�'j66���8��q��'�x�(�\�n/49c�^�\eƝ��'�r`���B�}�:pP�� L��C�'��!��v�IJ��'|�z�0�'�Ɖ3��5?��S���m%�"O\`s�6u�V��b\�\���r"O���F�&��F�xP6e�e�u�<Q���t���3G��L�\��,r�<i`�[$2�)�)A��8@��H�<���H ":����;���H��N�<����"m�(�:V�:~��(��IHI�<i��A�m0��=(��[4�F�<��+P40�	�"]3*m3í�J�<Q!e�2G6]���.�8[���J�<��#ҚN͒,�1�؀m-С-	[��dD��c�6��q��29!�d ΢��6��|� ep��ЀR!���N®�(�i��f���2Č0�!�䜗j�XI�eT )�N$0D�X�!��P�؂K�5vQP�K�#�8�!�d27�Zq�ƃʋ8�8K�,,o!��ȓyn�ȹWɉ�,'����b?�!��E���ç^�<;�L���h�!�D�KC�$�aG�1!ҁ�'�)u!�D̂V����# �*]8�m�
q!�d��E�b䰇A�.z�:l��&�<^!�D� ����� � ��\UcÖu!� cIQ1��ԫ;����a�5`b!�ĳ(.h���֍O����jʵNC!�d�rm���$C��!�$��"8!�DS�@(-ؐã0���V�D0!�Ɓ�X	�C.��P��!I/!��L<d����P�2`��c!�G�Y��<��$	,PŴx��%��} !�$��v�P��I$�5��ڽtV!�dǏ|<�[
�Il�`�e�+GL!�k�|(� Ɏ�F�\��ۓf1!�$	1&^�D�b� }��5#R�'D!�D܁J3j�x��O!m^��Ô,�uX!�����s� �MF��T�N>U!�d^�K�i҅�bA�s���	�!�:��x�	�.h>��" �#�!�I&�*���g�,|<�Y�c�Ο�!��=7�Z��`M��v rQ�G�Y�!�$M�=~UcCc��������@D�!���KQ.�(S�X'�6���@0 g!��
&u:�Y�D�D�`	ǪV�!��^�;f�Y��K8�u

��!���Q~��↣C:���S �*Y�!��İK�lA#��F���`ΔV4!�$E
pP0I��EӬ�AsJ
!��*Z�\V+�q�����P0EȬ���� A�� eI�0I����$W������� �\�1pS��!�� r�hP�>�̴�$�4�MА"O��Z��ܶ.�(\�P̈�\֞-r�"O����ͷq�H00u(�-Ͱ�+6"O̝(��L�aD��l�%�A"O��Ig&_�n���r�ՁK����"O.��6� �z�2x�D�@��T��"OL�r#��/ܲ�gE�A`TQ�"OV1G"^��5�<� 4�V"O�t�����d�s̖�SՌ`ِ"O �(�$�66Ӵ�%�a�(M��"O�P3�\8!�l�� )똜�q"OF�3�Ē|��9��JF^�B "Oĭ�vɁ���P0�,�&\��s�"O�ݢ��߂6�:�* �f���"O�`K5��a+>��6�º!�!��"O����9�t��r�õ���V"Ov�R�ɐL_Ԕ@#+'}��|iG"O0�H���"xfBͰQDФx-"��"O�� ˸cu&q���2e	Թ��"O$!�`��\m
쀧�)}|e��"O@D��m��%���IZn���"O.��"I�9�t|Xr��4�zd�"Oj�E��G5�Ȣ$�3
�\h�`"O��)A�<�P��݌)��`��"O����I�C�*�H��C6Ǆ�"OXձ�'�r�Q�u���`%�Q0"O��*�IH�chB�rNZ�7F@�"O�m�e
<����"@�0i�"Ov�2���o��}Rj>{,a8�"O ��U#��?�XјԩɅ#Z``��"O0�8�����������xCN���"O��P`LԴ	��L�F�g�,�x2"O�eZ��K�e�h�CD�:g�=��"OdQ�o�4�&=��
!e�$%�d"O�4y%'�q��A�'# k���"O�S!&
FM�yiql� &��u�s"On��͢X;Q´HR- 5�*d"O���'�sg&<H�M�.0Uz P""OHE{����	q��J-��DKdaPe"O֜ڑbсf��x��,ߘBD���"O:Mb��Ҁ
�`|x���`�J�#"OP�Ô�LBI#��>���J�"O���⥏�,�G��/�$�#"O�|��	ڳOl��Ņ���Rȸ0"O*d8�L\�r�X����I�Jq�"O�qK����T1�MA E�f�6���"O`�����4��d�%#����V"OR}d�� z���C�ĳo�T�6"Oh��I�w
����L���ؚ�"OH��@���=��,(#䈓[���jq"O����ĝ~�����P�1H�q�"O�(����<@����/�����K�"O�,��E&Oɚ�pE�և����"O��Wᘏ"|T:`��E�["O��hf�̞�,��'��.�d�"O���UESA��=CpO|}`pX�"O:!*$�I�>5.�3���?sqʍ� "O��S�E�|Tl*0�ȃ �FYZ�"O��3�㍿(��4����=�x�x�"OV�h�̀+A�p�!�"P� ���["O6�3�j��y""�U�)��r�"ON��cQ��dH�d
)�x��"O�a�d�*jE0䍻B&��v"O:�:󩋽J�9zA�
�\��졀"O� <%s��g\2��Eo�8A�V��S"OB̫�>LD�`�L8;l���"O���A��"�|��EOB�#F,{�"O@���D4���Ȁ+�,�����"O���h��~��L�ҠIS�"O� �5Ot-���R0j>2p "Ob=�o�c�
`1�"�'J�KF"O�e� �3l �J0B�:�XQ"O�Es�`�%���R��P/~΀��"O*`C�%);yp���J^�?z�w"O$�pFA0S���)���3k�aJV"O�9CQi�4n�|�{�K�6cl]��"O*ъ��Mm��B5��$EtJ��"O�iұ)E>~+P��%@�GZH8�"O���ǧeϸ�%"V9d���"Oj��J� д B B�%"O%������q�B
@�0ӂ"O^�� Ս8;��홫zb�8�"O��������.��#��<B�"O �ʷC�U� `�u.�� �#�"O� �G�+��y�DC��6�4�P"O��*5o��n�H�6��u�+T��yR �� x��Ɵ6N˒e��yB�˭/m4D� )u���R�]�6K�B�ɖn ԑ�*��*��BeB�o��B䉞&漃�Ņ�W��YW���Zo�C�I |JB@�����	L�s�2'�C䉡�X;6k-��-�P녣=B�ɴ��Q;��T)o����􆏊�8C䉦1�U�'� -J2(b��x� C��*�h ���\�n���
B�OȪB�cL ��a��N�l��� �jC�	�te(I����*[T��љav:C�I$2��iB��90|MZvbQ�5�BB�	�}�P@������h���2B�	w��yeO߅[D
=��- 0tc�C�I"ɨP���T�ޱ"%[���B�5 ��q�/�~�(�'Ǉ~��B䉯�u)�h�)x����I�ՆB�ɞ5>.!���?������]��B�	�[���	��T=lQ
�B��_gbLC�	���o��w�5�5�[>6�(C䉾�b����O���"/�6��C�	W��=�_���3��5�85��"Oĉ`ᯚ�^�l���`L����s�"O�����+X�򽐐�M!@(��"O*�B��_�X{��
�5v���T"O*���DO� $�2l�P�L@R"O�iRD.x�"�ð�= ��z�"OX��Ռ�/\�P�;�'�m9�X��"Oн2�KF.U궡�P�W#I�!v"O����)M@�����KY����"Ov,��oT�}�
y�#�G}��Q��"Ot<ҡ�R�[��}+ �"fB"�#7"O����VU�VL��̌U����"O��SN�aJ
@�u�?jY�tQg"O�3ta^i:�0�9Tp])�"O�)�ǔL@�ak��7�D�J�"OJ�K��R#XxHQE�#k��Ųp"O� {G�"m�(Y��Id�U"O!ҧJ�:���{�Ǜ?}b�U��"O%c�a�v�@4 ��£ -iW"O���퉾k/�E��e��5hRV"O2\�2�{Z��� &���`"O� 2H�ЇƺI��lڢ���; D\P�"O^��2��<mnq,�Kh~�;�"O�0�bݸk� J\H-H��"O���wf�L�y���9�|�"O@����4%hX�X�%V�'4� ��"O��j��_�N���#d�d"J��w"O(�a���[Fd�Vj�=;�q��"O����?`�=���v*4=�w"O�	3�A_�{���5�N+�8�d"Ox�h��έ 1����<�\
u"O� ��2�T3�cB
��Yc�"Oh@h���b�,�-\YV�bg"ODd��)��7m-St�+�"OB�#� �Ak4�
�E�?NY��y"O"L�աQq�*�˦dQ�MP^ؚr"OXHa![ l��0����sE��"Oz�
@�
l���/͚t�{�"O�l��NJ Ne��DJ"!v.�rq"OL���(9���w�AfF�IV"O��0�ٌ 6�!��ݻ:}�0�"O�D��K1R@Q�Ud��.x؂"OB��N�#d~ a%�v{��`
d"O���M�9N���a'ݮ@���"O�p��@S2U� �O�+��=aT"O�����R�G����C�J�� &"O��hÁ��7��=B�Ȅ
�l�0"O(�s ���48L�s�A�M�TX�"O�!F���@L��S��7j����c"O�M�`C�1Op�y� �YK��z�"O�u��f�%����	�)x� ���"O�̙�#]W8���$he��̰6"O�|Ô��>t56�hE�"qd ��"Ob�����j�l���n�x7j��"O>��b�L��i!B�_3$M�W"O�ۥIܮ`��8B�Ùy$�:E"O��8�G���*
���40eJ�"O��9�G���!�����^J@�ۑ"O؊tc� FĹ�Sf�t��l1""O������A�֗\����"O�h���#Iv�u��*#��� f*O��[�o_�r9b�u/D�~V�Tc�'@X􃛵p����P�*6,��'fv�Qa�̈́:�<�;E�
#���y� _�R�Y�'ˏ+R���ZD�́�y���m��oO�]�@!(���*�yRFC!M�.];�L[�-l�e��O��y�B�4'd�m�%��R�AV�Ɉ�y����颥���߁&O5Q1Ȍ��y�V6z�t �e��\+2�����y�b�]��0�L�c�v���	�yN����Ө|�,�3�"ހfI!��0C�PI��.́�Rhs�4!�!�dV�Y�4a�+��q��P�3�=^5!�G#Y�"t���.Km�ST/H�x!�DƟj/�;�h�'a�4x���}!�d^H����WVj�T��6�ÅKM!�$ۜt���4��4B�
�$�*$!��^+(Q��IFp��paΆ�37!��]��ӓe��:]�.�3!!�d��w;�&�ʍU���Y��!�Dٕy�̕��/��P�0C��W�!�D
�8����M�`���aE#�!�$��
>��:�n��`2 �Z�Qr!��9p��p� �"DN҉�U
K!k!�� H��E�%
QT��Żs<��h�"O�0��3_���2-B4%T���W"O�Cf����L]5VH���WO(DFxPK�hɀ1�TUb��0<O�؉%%WR��H5B�����1"OP	 ��R.c�l�����F�,�"O~q�Ua�L^�V�� q*]��"O��bY+�� k��ܕbl(���"O՘U
C�p6��;��#N���r�"O��`J�H[��b�,J�%��ܸB"Ot���ORiN�A딚{C�=�"O���R�'��x��/]�S;��4"O�l��L� 8,q��c�P��"O�p�E#�%�H�CT���u9p"Ot�� =];J��Q� �j|�U"Ox�E�G�\)E���O�r��� "O�0���^�E��9��O!����e"O��V��_:�h��ԭ>V�yx�"O���eʈ8���d)Y���%x"O~�+�oT�g�R�BӇ� �`LѲ"Ox:A�S���3���N�b�y�"O
]�)A%PG6���KTL���x�"O.]ᗁ�;�|�Jre�(u�f��"O�,��.R�'�V��t�"O�0C���&>�d̂sÃ����"O: ru���hz'b��82VL�C"O�:&��K���	;"O|9E"O�<���A��Lx C�i#�T"Or02�i��ud̓�얓k�.��"O���Dҍ���C+A�2d�\a3"O�h�C�Ԋ]��������/  i2�"O!"��w�blڧ�}l�I�"O�����2q ���P�8 dѢ!"O�\���8�>�{5	U�(hC�"O���b`�F��V���=�Ñ"O���G�*�ΐxt
��uXx��"Oty�gaS�vX	�w�Q�jl�9A"O4hag���f�# L���:#"Oڡ��)0[l��n�/��H�"ON�:��Q�d���;����jɁ"O�`�� �	h8ĩ�I�'QР��E"O�`��u�����.@�qn�u 5"O�qC��P�J<��P�64> w"O. cu�;u��Iӎ�:b0�+a"O�=��)Z��n(@�+�8 �#"O�,c���3�m3t�W����"O���V\X�ԣ1fAl�\Ѣ�"OJ��r.+��L
�K@j
�`�"Oj���a��0�aqh�`��R�"O0Ѫ�F�\`��qU�K�q�6%8"O�͸f-�#k��E;''�' ӄ�H�"O��Xp��!���A��漳G"O��e$Ʈ>c�3�C3s�RPc�"O� Awc�0����e��V)�k�"OȽ{��:/V ��T#�!S�"OV�� #����0 A�%�qx"O2aZ$ �L��q�B#E��S�"O.�&f�8�+`�^�3��I� "O$�Ȝ�gPdp� �l8Ġ�"O�]3���҆�@�� q2���"OZ���I��)�D`3��\�%+�1+Q"O�tJ�͜\����1��?1�yw"OƨÂ��5#��Ӊ�d���"O�NTd�&���q��"OAc�aJ��cdR�R�x��"O� �A9�g��1e�A�%d¸u��df"O�(W�J���Qfa�f1��"O���g�R9���aN��(�
�
"O<���O�`��ْ�������f"O��)E�_�3�ĥ���^�,����'"O�$�d�����;ń�,f�0P"O@x(l�%�\�3�Ƕu�@e@%"O*|2���94�#'�5�b	2�"O�!��R�Լ# _)�j("O6�у"[&%*�9k�O 7.�8YX�"O���ZC�mQ%�ۊ�ʁ��"O.��_�n!jƮ�6]dXP���F��y�C�0D�Np��Y�>�>�:�Ȁ+�y�D�ybxTp238�d�"�Q��yҋ	t�tf�ͪG��%i�ID�yR�Qh�8�y�D�l[���'jܲ�y2���Ӓ|��昹h:�H��ٿ�y"
\7���A d�>["�X:�����y�T��-�0��O�h���#�y�KB�L�)��MܫFK���'���yr�T!k�R	ئ��8�f�1�K"�ybm&'j:`s
A@�������yb`
Qhb�����;�
8B$F\�yr�7Dȶ�h�G^*|�����k��y�G�EIH��l��$p����C?�y��;K����(��-�0�L�%�y"�
"}y�Q�P���P¾Y�PeY��y��h�b���mZ�F����Nż�yRAŮ&���"�>8��Y$�߻�y�瑒+z����Zp�Q�3nK:�yBI��'I�P6*��8�c߭�y�"λ!J�;Q�
-#�N��C�T5�yr��cEhA��m�v% ��(�y�/�\�h���ufv��`�&�y2�|�$+A͊0� �*�yBᑸ4�(k��Xzp��y�!��L1ag�Ԩ\��|���yb
��<�X[���=S5
��C�T��y��v��'�F�O�� yr�ѣ�yҋٟ���2�A7���l���yDR�&Z{@�N�"8�Yq�֮�yR�']3
� ��5��)�y��SZ��o�
��t�d���y���;|wk0f�c�0�j��yR
�+9鉓�Ida�4���Ň�yb[*�8}�bn��eʸ��j���yrƈ;by��j̏a7�Q�@�%�y��|�Nl�!Q�S��=*��y���=���i��T��g�^�y2a�5x�%iq*��p2,�8����y�툴x��K����ĕ����y&L��~���e\�ڀQI����y��v)�2���������y�L�g�\mKC,F�"u��S�y2�
�V���͊�Q�l������yr���t�u����'N?H\kW썐�y���~&�9A'Ȇ�>4���B���yR`��K	 � 6��@X�m���7�y��D��	�n�F�ű�J���D���Oٜ(qQ#O�&_����'�29����')�1��`˧hut�i�k�3[�!�'_Jpq�B[�G����@�4(���b�'
�������4q��92��
�'���g��hfK��dY�H�	��� �5��a
Jc�3vҫ$�HS"O~I;S��vt�*tA 7E���"OR�1�[< ����#@�;w�V٣""O��s%�l#��t�_�^x����"O��k3�94Ҁ(넪P*<qr�!R"O�e����S� 9�ԉYkbp���'k�Y�A	�X�6�K�C�y��9x�'��@�v�ԧUvP�/�u�`h��'����5��M@�:ԏJuv,0
�'<���<<��L�� ID�nɓ�'��\�q'Y�I6^pHZ�f*z���'*��s�Ļs}LdAG�	n�$��'&�����1;!�,RKMU��"�'����c$¡^�Z��Q�I4��M��'�Z͓��O���Hڹ2:؁�'h6� mĤI����T.��xE�`��%� �&P���\�^�ر��j�<�G�ɭG�\�s�
k�9��J�h�<����'-h0�ta�-4x�d��c�<���(�q*���0$cI��ЅȓW�A�2�P��@<�%#�dV���ȓ#*��2n�p1k��Bg�������C�f4:`YL]0�\���n��1��O�3.�x��E��(d��^�
}�N	�ޙPG��|�@t�ȓ}��Q��IC��R# ~}�ņȓ_�@y��g�8]��:�-�\���u��������b��:�٢1�+D�����>�l5��bD�u����l+D������ �X� ����%D���t�S�R�9�3��	a��C��6D�$�&Ꭰ���Sf!�?~�y�"D��BL�$|�Se�wȑ�s�<D��z'���n�\K.F(4&h���-D�����X��<Zp��%6DM9�A>D���-�JA��@33&>�s��;D�t[�F�Rw&��I'?�4�ؤk;D�ɒ�BD����X�F��qCa�&D�Px(S"��䡄�*҈q:Q�7D��c��|6)+�}d��7D�ڲ,�%\�bͩ�nZ$X�J��`4D�l�0�y�X ���+D+$��W'3D�8�#͐[�|�E� E�ȫ��2D��c��%���P�h�0eB�=��g5D��+¦Bk��+%`%zb<K�3D��i��L�S�)�Po��^,S�6D�XS%6t��i#�E��5q��Zu 5D��i���>2N�"�@	�#̍�R�6D����w肄����[��C��3D� ��Ҽ�h0�&� �7Ι%�4D�H���w�d�[���8+�t(�g?D�@��NU��<��F��>r�>�A��?D����,�i�:\�b��Q�N�y 	=D�Ի��E�~r��12FZ!!��R�G%D���Gг'�0����Y�P2ff$D��S#��V)��C��o;��V�6D�����T���B�E��� "�?D��iP<�9�O�M.�p;#d D�d��
"@3�XG-دU����=D�0x �̇YQ�}�͑�܉c�j0D�tH��ǽ�j躳���p��ѣ�c.D��� h��m:�6`�V����6j!D��æ.V�aڂ��2�V}��B�?D�4�W�ˁ�v�6 �<���ď8D�� ��a	ty�q�A�2�B�b�"O���	O*�A���gի�"OH�1��ɑ]���9E)���2"O�}(���P���D0�i�"O�ͱ�ƣ+4pA�)�e�|�"O�a���N�vE���-L߈�J%"Oi�S�[7 |�`FȄȄ�"OX��5��	R�@	c�_�Dx�"O�ę�苮������)J�M�$"O�(@�W�5\l�Y0��'@hd"Oԭ 兂(i[dX����$_Ɛ)8�"OHy
�&�Lg$�C�K��n��4"O���C@��4��e�1DֱqrVHu"O���C%E6*�`�S��ˊyL����"O� :Q�܃~�U��"T��8��"O�]z4o':�Q���֓!���@"O�􁄄���b����$��]q�"O��@�VÚ�� )_*H����"O�Pqʝ�h~QY���e��Ś�"OnJH�^3�h��������"O��C���LI�Ϛ�17,S�"O����e�;�%Bu�-~�	�E"O�[�EO�	�p'K�)=�8���"OV�ٗ�O0
<h�%�� u�~0P"O ��6)ɐA��ء�ОD `��"O��#�P)%Ÿ郥�]�J��G"O�$[q	�>l)hV��1[�i�0"OP�Xe�	Aqƈ���U�=�ެ!�"O�%PW�H�^,�k��϶4��"O���1J��
n`�f�K�����g"O��Bj�v�+b
�%;�����"O���Mɦ��1��[5#�L1K�"OhK�kJ�}�ተO�RĨ�"O��c���
y���J�͗)%� @0"O(�ӣ�&�ly�B�5��ͫ�"OdI��NŬAn��������`0"O�\;sF�#gd&���֪:M�U�C"O>�ö���9ż��‘�n4����"Om�U
�kF<�d�8/ܙ��"OVQ��ăq��H5�3�!��"O$�֤�\��4H�BQ"��͂�*Oj����"+�
Q���J8�t�'��0yW@��O�|�EDNs�$i�'Z����V��0{u��E�T��'�dux$$R>(�tO�6;V�B
�'<c�I�����GJ  ��'�6�S�@D�\�\94�Yza����'�K��ϗ=�d4z3�ԡn��(�'�1)�o�=�!��g�h�>���'�ΨзJ��YP�b�N�4w[�T[�'I��B���*@0�շi0�@�'�����I/ռ�0r�@"U] 0��'����%�mv��ġN� Z�}��'�>Pa�#�WY���T� o۞�y�J�-��&��B�:�')Õ�y2��)�d0@��A�3���d��:�y�F�+��1��1���N��y��VN��!LI8:n5����=�y��,_��22�F ����f$E��y�6>���D�Ћ�t�����yR�	�r�<!XS�[��D�q���7�y���i�:�9n¼Gn9���y�$Tİ@!��"�\�`�#	8�yrH� �P0`��:x]��gC)�y
� �١O׉y4T
�B�k�,��"O��r�_�"���q_�q�dT�!"OΌ�Ui�#u���V S�w#X%j"OF(���Q�K��3�(��2�,� "O|I*�!�We���r������P"O@��P�]Ϯ��%&�
	�a[��	i�O~QpD��Vd�QK��zH|��'p���$&IΝ��H��t���:�'�B�@xA���?
��'�TUb� �+$!`YqP-K���s�'q.�z�+��
�z������n�V��	�'�R��6g��OlaQ`惑#�|{�'�"�2Jڥ�d��W��> ~N�j�'_J�)���  M|�I�Q�_+�t�<�B��2I�5�d��N~��p�<I���;!�=�d�Ɂr��=�lUi�<!�N��y)|isFY�\^� �d�e�<��߸d����A�QA�2�I-S_�<��IP�vdnP�`�Ը+æ��Ǭ�Z�<��c�v���2 ӵH4��R"�j�<�@��^&���aֱVu�����L�<�7J5m*�Z$n��n�0Pˠ%L�<I�H�H~A㲅32�83��H�<U��@F��#׈ψ+j@8P)�L�<�1�R�iqvР2���v2���D�D�<���4-�{U��:�t��,�J�<蚷3�hH� �P8��H`��C�<y�D'K�tAKQ$��0�3�&~�<�B�ְXN�%���+ ����[w�<�U-ַD_��aq!S
'��l�aa�u�<q�n��P_DI����!8
@;bng�<� I�-^�� �� L���`*v��`�<�C��
�l��lI4x��2�F�Y�<�Os㖤�FV��lQ�a��y2�ϊ(Y��K#G�u7��#���yb�A�e�r�2��i�f]��Ѡ�y�E��t��� �(d�@D�aG�>�yBb���1�E`W�\�X	��]��y����d��hb�M�}W ɋP�A��y�l^1t*С!�K�+�La"�bĈ�y��Q-T]t��b�2}xF���c^�y��~G�9���w��B0ő�y(߲`�|[�hwk�=��� �y�k�8�ΝrG^+N�s�"ڀ�y����q6F`@@@�^�閭��yB�PC��m�Rm�(v*�l;����y����;��]�4"gJ. @5�:�y�� ,l��,�✪W��m�i���y���j{V���&��̙��J��yҥ���<dÀ&��1�^4��@��y���GE���ņ�%<8��M\�y�(>T�A ��*�81�W߼�yb�0w�&Y3B�+��m�5����y��Da���X�%V������	ܯ�y"d��[jD�)ѷ����D��y"���/�D�����.���A�ذ�yr�,dx�� !�U8��F�y"c�>���1Bļш	���^�yBӠ�J����f�P7����yR*[O|R��Aŀ~E�R�@��y�hW=2=L�xQ
E:}E��P�y [�0+R��5��#RQi���y!�`�����ąH!����ć��yB%f�&�.��V"��hr`�*�y
� n��� 
�iv��	'���K�l��"O �"�F��)�д`��=��8�"O`��Ñ7��8��B�i�T���"OFd�w�P�b�2=��H��)�Pa�"O\�k�Ā+Q �I�չb�tj�"O iK�\j�1��I�R���B"O�`Q^Xe˄�Try$��dI*|�!���82�
�;@nO�>v�]b���K1!�DD�/"4H�c�=5�&hs����;2!��V3G^V�akS/ߦ�)3,M!!��0$ò��C�B4y$m݄N{!���I�m0��Q�{d�d{��)On!����@a�f<����HU!�DӰ6�������1mJZ��L�wB!�Ğ3���pv`ͣk9�m��쌪1A!�$�4~�̰3Oѱ38���I�	o.!�d�+m�|�D ßW6z��+V2I!�d#"��G�X�tTM�s��5YT!�$��tX^�J'C̡=���a[[!�d׬Z��e�(��8�W(�LF!��F#4��a#�]�3�V�� ��B(!�D�$��lRR�ߕ�0�tB�0m�!�D��Ͳ<�g,ƖpZx��fBM�!��4w����f� OXk��G:r�!�d˔]����Ô`@�H�E�D!!��$�LC�CC1V�"���#!��u��Y���o\�1`Lˎjj!��ԭi�>����!+����E�$g!�U&��z���L
ؕ�a���!�d�#Ĭ�3�m�"���+@EU�A8!�D��^���Q��� h�h�"�-!�$aE����Fw�D�!�%�O,�ȇ�iR�Av+�w�U9�@��Aâ0��t��XNF9H�BX�%Ƃ��`�ȓ3}�=y�؇AE��z��SYp��ȓ+��a��ă5p0BD�D�]�HՅ�D
��u#��(�q�jD8?T@]��@�屃��8#D�(�i�Jb���h�^�/��2�ȋvnV����K�<��(I;b���@����&�X��BN�<y�J\=&�mȴ&��`�]0�#@M�<�%*ЊwHZ�)vnnef}��F�G�<�ӧ\�xҚ�(��Y�D%��kơ]F�<�u]�ތ�%�H6�����)�<)�b3I�vU��9 2 ��AIPx�<��/	��]!#�6Z���wo=T�l+a�$U�|t�0�.6�\���5D��KD��G���Z�G�;:�}�3d5D�,V���C�떢L��B1D�0�uGZ9��`���+�����i0D��C$T�.E�T����:�.D�(*�'[7�~�9�dP^��QqRO-D����OE�FXc%M�0��@2G-D��Ń"M�8�⋮��1Q�f5D�8��@�hF��`�H�}f���W�4D��K��̃p�`a�s�R.+�}�23D�ܩseT'0�q�T�4�	)C�<D�D)�ˌ?.z��/Ґzh� f(D������� v�Y����08�8!S��8D��ˣ��;GR|#L��skR�(��7D����W�3�hyB�)�Q:Rᰱ�'D���b��������,X�<0$0D�����^�Q����[���xT�-D�P:�c�3��7� 	}�|uy�9D�� N0w@�c��� ��<T�"Oؽy�#�7IȬ] sn��$�d5"O�{��O<$�����BR�!�T	r�"O�(Ca��)2^�����#q8��"O����9�Pc5�@0�"O2�3�e�v�@ ���.��V"OluC% �<!ZL�$�8r
��e"O�Z��U9Ga �!�A� [n��"OF٠W�c=0iJ� T0n< ��"O�P�D�)^M`��Eo
l8d���"O�52���#b,ʍR���Z��u��)�O2�sc�X��MìO?�I�i�8�voO
5����f/��Q����cF�R���Y�N�\֦5�%P?j�>!����0�w�_$Dg�P
���]JU�i�PM���Ęj�I𥟯}�ʉC�s��B��~���2��%�-�Q�wӒ1��'�7MC�����s��M�5��"77���v��|�|k�ɔv?����$0,Oΐ2�K Ek)�g 9zĴ$i3�䦑yڴ��+m"�)]w0��c�,ֱ�E��
d�}���<�&a"���'��9#!�F�ȡ[��ɨp\��2h�"�4PQ�Q�w�<�������Ɇ�O�hg���q����U��(��@E�&E3*�
&,QIچ1*�G�!=5�(�O�����.����M
<fb��	��H�Ƞ��HʟD`�4J��gyR�O���9MҘ�	3+T#��a[Fo4�C�ɀx��P ��ɋ'�
����7 d p��il�7�)�d��B�)�<���]	���{���+������b.�y�'Ͼ��<���1�l ���6T'V�A�90+&Q32Ϟ�(u�t!b���D*PD��0#?����'����
�)� ,�e�R|��0AF��g�&�0���L%�5;���D�ҽi2�aЁ[�$��C
M�'u� �d�G���	ey�'*�'�����x�,ĊW2�hЕ�~���"O~0ذ�]�@�$�����P���O��oښ�M-OZy���������I�ӓY-X�4&IS~���7��P��}�v�D��,�� ��N���>���󒂄�D�%���&(�j@鉒'&�YSDD���3C�u�҉Q�O���S�z�p�;��յC9>={����2cӐYo���O�F8V�	�h,��+���84��O�˓����O������gԓr�ˋ\ $0��'����uӜ61'��X�P��/z �:�eY�������o��0����_>˓��8����j�{2ck�(ʱ���2)�#I�Z�:X��C��+ʒ ��i��Ɍ"1��`�0B�$�Nd� ���MK��Ux����#[�x�<q3��E��|�1y�������xa��[֎�
O�D�n�yC��d�Eݴ�?����i&. :s�_�Ah(Yg�՝0���'�Q�h��C�S�4�ѰBq������$���ڀ�E �(ON`l��M��;`���'���N��Ȇ9
@�Sf�S!�|C�gy��Z7K�6-;,OjC�YVh���0`����e	�vE `@�"�R���e^j��5h�|+W'�	Ff�c��R�e�@DBÄ/A8�r��8B���je�J�F�����v�dȭt�R��
ѹo�l9�f	��� W�����O �$���	Ɵx�'J��H��+�D��%~�Xh�>iv�S�3?�����bΨ�2�Ӥu�����i`6-8�4�@��?��jӊɕ�  �    r	  �  r  �   $  b*  �/   Ĵ���	����Zv	L�l�H3R�PΓ���qe"O��r��<���*�a.�s�"O��Ѷ-��cU��`ȋ�}E<x�� �h�(�BVZ���y�E� ��)�&rq�X0͎�imlآ@#
�t�t�x7
Y_���A�^,(~
�D̈�I�x�P�+�'&�ĕ""&�DФh9�Rs�z����[&<VZ���Ϗ�U�u�㑘B�y��e�?7F�e�N֊'D�q���8�:�mC��?)���?�����*D������;<L��1�C�I�� �I���y�&�6,����bܘ ��3�%ҹZ2O��V�J�W$�8�S�P�%�Ԭ�p�T�g�:!q�Fx����5a�\&���r��o$~e� Ī�����<��e�ɟ���w�'���;:Ǌ�;�m	�X��J3��n�!�ű��)1E����A�L�!~S� l��HO��O�ʓlC�#�$K 3��#hH�op�b3��;=\����?���?AT��z��O���U��%����cf����rn����[t��9�`ݤ|�����#Cm�ʣ���j9zQo�#@� r��Q�z%����>&���oZ(-%��)��bѢ��5@gHe�%d�"5���ѐA��e�n��M���D�O��擓\#@����ǯE��Y⒂٧&�((P��D�O���2�i���Wc<n+��4���8%w�V�dҦ��Iry�DQ>U	�6��O\�d�OkLR�Er��r�nͳP/�����g����.]b��'7�[�y��Y�6��W�b�'��� uI��9�J��%��9D�+�ў �O�	 i�����/c��	/I���"0-���+f��/c���ʦ��ٴ�?y�O��8��ƈ!d������'deK�498�����?-O�έ?�K7"j�d�(@�`���|��L�Ă*,b�'�ў�8��$�f����LK	uDb���̏j�`�'�&Hh1�`�����O��d��48�a�Or�D�
@*zu8@��0�\H� ��w�@lګ'nޔ0ii�%+b���O/�S_?���
�m� =X!��T�6e����L�uiޞ,�<�_���|��
�X���Q�	�%�$���@�$i,Q�u��X�z��һ?�r��)����Ƛ�'Iq0���A	Y@�'�<\Pr���D�O��d-�S�>Xyؓ*x�����Nufb� ��"���<I,��8�0�_�+��_�v]d|j��ʦa��џĊV���}��ҟ�I���\w��@ ,r�,p�%��;��P��> >��6 ��ɖZ�]���A��a��A�+;"�Y�E��I�S���d�i�zm*6����R`�Q�Ɋ�0=���6d~�h@�D�$z��P�
o�<�$�=Xy��8�%�? ~�|b��Ԧ�K��4���Op�d�=aϴ}ːN�1Gv�i����.��<��l�O2�D�O�d�Ӻ����?��O+d|{��h����B!V%X�.��fC#�M�&5�O��e�O>ݑ��;F�RA�BF�#KE�����'B����m�P��>�� a1&�,EF>�9V"O ��(U�b���
���}8ำ�"OD� �$_�4D�Ȋfm�C)8K�R�X��4��j�p���i���'J�	Ь���)����%Çl��q�C�<.r�'�2�ƻoU��ԟ�=��S�U�*R�'_ ���ɒJ�`�~�J �v�@��v7hٓ�E�'p�"��5�>�:4�!ɖ}� �5/���3D�H�&�>xS��3���w@v���-�O~�'\���PG�+,nb'b_�3&`��O�X`s�+1�8��3���a�!�	U�F�с���HJ�Y��
�H�B�Is�\���$�h*�l�S
V�p��C�	�U�6�Pv%'^tJ�7+�a�C��%a�
��'n�,e>�a ��V1�C�	Y�IF��'y ̏��rB䉞^g� ѶG�:���*�D�XB��-$r�@�k%*IcUHP*}�C�	;6qf�kcc��B\�Q
�nyC��5C%�|���O9 �&`��I��ͅ�B�0��-7a1��7Xp��>(������}�. ���Ba��ȓa�<�Ã�����b�Q��ȓƬ�"Ȋ�dy�Hn�N�cXXA��`]���6,GI�!"�jm���i~����>_^��A�� Y�����7
01� �̐<��m����>MPɄȓ�,�+�l��X��LI!h�9|Z.݆�cWve�0m!�YBA�23���c���T�Q�B�-`r�Sg<>���S�? �-��E��p b��M�'^���"O,`��g�����'%C�+�"O
��V�A�"\2aP�`ŀ`�"e{B"O��;�	Zl�*�+E��2]��?�yr������EY2A�����/�y뛪H\��Â��@�f��'���yO�K3��Y�	|lK��˭�yR
xi	�#�?0��&F�hk\!�ȓ}m!3#��JӦi-Iђ�$"D�DbɃ�g����D��vE���!D����G
3��lC���F�vٛc&/D�@X#�"�($B��O�;�YqP�-D��ѵLӜSO�A�!jZ\X�젔�)D��R��>�T@���8t`��Q )D�|��.@�����K�w��ZO7D��#�To}0H���:?ޅ:�E4D��r���,Ӯ�	�ٓF���2D�$�ǆV�  7&�[JT��4D�h�e)ӥ]��}�gD�_� 0qql>D����%�Jyf�-i	����yKY�Uq����iǁ}G�M���R��y��*T��&���Z����'�yB��:�Ȕ+��1Hì���yB]1_����@�7�6,�i��y����W~t�����*C�4Є�[��y�/�	�Fԩ��Q�+ �E=�y҄
�3�ʍ�i�%Q̉c��Y��y""ށ]�� ���]&V�llX�� �y-\�t4��D�� �����چ�yB�Q�̱p���R��EK��yR���,���^U{`�ǎ�y��ܣ����(�xA,��#ѫ�yr�L�B,��� ���mº�q�$��y"FL�� 8�� d�tQ������yb�EYҕ��(ר15�]b�,R��yrD�>]��P1� ��([���v���y�H�/?��Xrc�B�(tڱK�+N+�y�B�J ��0�ޣ&���C����yb�)uH�Ha·#����JN	�ye��5N�i �:Uvv��L���y�H����1��@K�B}�����y2b�8\���C�76���IRo�,�y�U�X0���1/�* ׀����̊�yBϡmZ2���ˈ�@PF�B���$�Py��σc��(G��:� ĝt�<����*�!�T�U��L��MKo�!�$��V2�����)!6���e�2uo!�?V�)��7O� �'eσ�!�����c4l6(@�0`劊�_f!�d9=��)�#E�*�Ԡ�	ŽE�!�d���h|�D��3 "�A J	0%!�-�`�Z2FDiyDs׉;6m!�D�3"$�ҭ	2{���!�!�ȕ%�ec�Ɔm���n�9K�!���(����D.&4H��ǟD�!�G�+Z�C���~*��B��J\!�ҞMtm1��'f"�ReS!(�!��B�SԊ�ztk�/�����G�O�!�D�/N�Ԥ��R�\�h����ʵ�!�Dˌ5�z�To��&��e�� f�!�D�a��A�Ǥ��|`R&���!�D�:MƎ%ضKΡ3xDY�bW�`!�d(Jn:�`�+& ؊$C՜|}!�dl�jfn8@7�X�d�ȹC����� ��KÆ�P�ܕPvO6~z(!�"O�$`�G��M�Qd^���bO2D��o4b~|�#��ܖ����?D�H�D&Iֱ��m�"f�h!�O<D��P���7c��!����5�4���;D�4!w�؈Y���{��ՙ2\Ġy��;D�t�'.F[KЂj���K�#D�BS�Ŵ�%1A�T*���6D�Th�	5�6=���o:�<[�/D���D�,측I��گ6褒�/,D��J!F c� ���Ư��d)D�<�D� _)�܉�.X�I.�2�d3D���r�	(dw�] �7�(��Fb?D�$1cc�3"Y'T'�9 �'D��Yq� tJ��"A��5UR��!�'D�|���4p���R�� u��I*D�`��Q�L<<Րe�!(�4�h`	=D�p�Ŋ��3?F4���<j�Q��(D���#��L"^9���B.���(D����=<6��̜0���B��t��Q�k�Mx�hʗ�X�^�d�e[$�n�z��/lO�mi�L����	;=�l�B�ĜP� Pf�*��B�I�4b�Ol�<)�[p�Agk!�"yD�CccQ�W�bD�D�H64Gd��䫆�\�\�2�'ݚ�y�
�vԨ�ʐ �[�8t�1/��kC�Z�L��ɓN��#|�'wx�'��.e|ȩ�Ǎ�&f�1��'�@���G�O�2����8����K�~E��!�:K�:���''PyB"��"^�8��@�>zh}a
�ż�s�Ǒ*d������
H*��t�LL�H��ulB�_w���"O�\8��0�����]4e8e�>Y3c�(Jp�qa��K�� �/�'S�X1�0��P�aA��yl�%�a��NT^����ER�U��nNY�L1�@�e-��4I��3�q��'{f8�Q�..���ׯCyĥQ	�'�f9�U���PJ�0 �6�0E�X�N�	��� C��p�i+��y�e�A�|Ё�ۥMnP���J ��0<I��._.lp��������	Ā#� ��\,�Yc'ĝO�՛���qh<y��БP���r��4��q	V~B�	H� i
w�(l>8bc��̄��NLo<p�"Lx��w"O¥*`�xjʄ�!½�H@s L�BFp����\�l�"�y5��$t�1�"�O��pu��?	���e,f�T�O��rq&�nN�m6���y�dȊE=&�	��,˦ �Hٙ�E������d3-�Q�P�p���t��x��WJ�4A�ƅW�'��h���#� }3��ͺ;wʜq#�$d�ՅȓC�<�9��\�=_Ĵ�5KņwyBQ�O��k�c��Mo�v���u�����I�'R��3Ed�/����nM�$�!�d˭Fۦ	I!r��uƙǶ�h�e��Q� �O��}��&���xs��D-r���^�	(Fd�ȓ���{���E�n�)w.ܰl&�lZ�<�����-}e΄��I�|D6�A(!��U��?l���ĝ ��z�/���?9�$M%�8���L7M>��B�F�<QS�V�O7|m9G;<t��C��B�z�� ��j��*6�|D���_F@8A�* �j52$W�M��y"B6j��yY«�d[���F��h��a��"�w�	��H��ɨ1i�i�P�݈ ]���W)	m5:B�ɢ{�:�h/G4��b���'}bL�	�Vq"!���!KN��� 느o�j2�D2L
�C�Im�� H\#&�j!ڡ���vB�I����a ��BOF�5.\#Wf�C�Ɂ�v�р�G`���f�a�hB�ɔ6
Ta[�aS�8y���� �K%�B�I�7�ޑr��L9V�4��c��=%��C�	�i��9��&Q7Z�*�� ��qϜC�I-�. �p�H�>��� �־"zB�	�{G��Ze��!H��\jd�վ�4B�)� ����.V�<
��8�n� r�29;�"O*\Af�Y\�iC�o-z�A"Ol(vLT4R.d��oߧ+p��"O"�A�Z�V��n�6jE"�[g"Oj��cO��eA��W�Q�dhY3�"Or,QE�&s�8���`X� E��+�"O8uS`� �7H����7\W.��1"OnŒ�e�zo�(��1 �N@�"O>8*tǄ1�ֽ�$�)�L ` "OT�#(̌J_Z$�&+�"��T !"O<�##�+H�HT�)��MS'"O��d��U�0Z�	�6��1)�"O2�)X -GIc��K�o�}�"O,� �NF�q:z@`v�2R��iJ�"Oƨ��L��0D�H�m���Q�"O�Q2�0�*5��|�RH�r"O���r��?�R@����L�n�8�"Ox�1����(F�.d֖ɀ�"OT�/�5;9<y�v�#t�
�9a"O����I� Βq %���X�d"O��!�L�7��C�` S�<�@q"O65����#R��) E�A�<&�8h2"Ol��뙳[j��8�N@1*:��6"O��	��oЧ�b���"O�Y�C鄦H#>0�ǣ�%[}>�1"O"!H� �|x�K��&���"O���߲x�I���/Z�|,��"O��kT"T� O��K4H�
�P5"O��s��[�:��΍��h$"OƘ`܀.�e �9Qxn��s"O ��ׄm.y[ 
R@�<u"O�EP�e�f�1��@F��v �1"O�e#��I�2FD����Y��2��"O����h)�խ��J[�"O����cA�Jw���e��,�:� �"O��"g��*��̐�n���F!�"O
鉥,�/t�aHTmR:֩f"O��&K�/@a���2KU'}>>(*'"O��!�mke,� �=�29�p�<I��p��(�F�E�[I�C���r�<�7�����֋ʔ�r,i�NE�<��!�Wyb�21�.s�eR�J�@�<I�f�T� )���%OD,r�B[�<q���G�fp�s 
�}��)�#��P�<YW��X:�����:gr�H�b�<���R�!2
�i�!�TG�T0�ɉt�<)�n�.L,�7g��al�<���U�px44K�O
\�;�Hr�<9¨�#����-����S�Fx}��.N�h!f�N�RuB`V�Ձ�HO�\�WH6r�y�������f"O�)���Ȣ-R��y��۽}��\y3"O��0Dِ[�*�z�T<y��Y�"O�Л�V��be<`9���"O
A�� ����0$[�#4ژr"O�X�`�^]��H֣N�|�:��2"ON咣N�#���0M�-Sb��#"O�K�	�,F�J�+ÂԝYR�`"O��3�W5q0�2��&k�����"O�ѻ�l[�A� Ȼ H|� x
g"O��B箏�]9�1�&_^�j��"O�dq���g������]�uҶ"O�L�R���,4�X�%C�=r�p��E"O�љ��W=e���)�B*���"O����k�"Ty�+�H;��7"O� �y��B+v����OD6 Ȁ��"Ojȃ�Čl}0����I.v	��"O Q��哳8"�S�$�+�dh+7"OIcW%Y��-�w㓠=|�Jg"OT����k�z��peL�1"O�ŸL"8�"�+��R�Q�"O�Kt�9R�����Л8t���"OĹ��Ɠ�o��*���,��Q"O@-yC,
A�Y��Z ^�lA�"O��[W	�����(V���y� �3"O�i-	�4��b)�~��3�T��yT Q� �����P�^L���
�yBU-�b��@U��:�	���y2��fr�i3�/B=�.4��%��y2&�~궝2%���Hq�:�yb��|*��x�"DqP퇾�y���=H��7�m��ز���y"�ӿ;�8�����"g]l� �����y2�	�_VE9��ƶ^�D	��N��yReȹ���)J ���a޷�yb��w�%��ǉ'��l�D���y���%)J���fW���%@�����yB�{�^=��* �XMd���y��֘�%Q������c��ybn߇&��R6�*~{���,�y2���lA���G`��`U��yҧ��:��`� ��h}~\yDK��y��<=��hPoD�4Rވx�φ=�y�1M����*�3a\� I+�yE8P>p0fR�/;F�	��ǰ�y"c�/N���;"��7+��d��j���y���a���c��6c:�c��ޅ�yrl�	?����J͈3��ז�y��'0�J��D�\�J\`3E��y"Kם1�p1B T��<P����yBi��B�+3�A��J��y"&p���c�	t����ݍ�yON���{���9mu�%�yBL�<�,P6���,P��B�K4�y�D˖6����p�Q$Ehrr�ӏ�yr@^�tw�Ju���
CB��y��E+*yh�kD�9�&��J��y��S�uz���ҡN�p�*��y"lA%��['�K�I|�(@����y"F�f��� �<��,�4+Q�LK��Y�����é�� qSd��Qڒ�!D���!V�nw�ș'�#3�H���bl���B
�Q��d ɿ0�9h�/_�7� 8��	���K� ��&'�0@vt0�"�� #���ȓp��i��j9~�RP4�#K9�	�ȓ>�0�0��v���[д�ȓ[
R����%V,5x��u�D��ȓ+��[�Õcu�h�lX�*�ц�	���키f�̉���-���ȓ@
���w�ٺ�v��m�%>e>)�ȓ7�������,Ё`��z"�ȓǶE)�Y�RĲ�� D)J�pe�ȓ*<.H�1��LɃdL�����#�> (��F
3DIrƇJ�&�ȓ��c��U�]��x�f E��1�ȓUz��be��	"����,�����(:1�޴|��ѳ�V��0��}ʤ�X�����2ˀ�IL����m���F�Z�4h3A�<�����S�? (�B�n�=I��	��ŌicNi��"O����V�_���B-6x��qf"OL�Jd�A�s�:��Ȳkc�y��"Ola�GD�0����Q��"Od�
@m�~Ӕ���9�x  �"O�����.�5#�DAz0<�u"O,X&&@	Mxj9�bIƺm�XBS"O�M�q%d/�] $���+$"O���KM*Z΅�5�٫>�d	��"OYq�kݓHcf�`�㉁�L�X�"O�qAƄ���@u`N�H�v\�"OV�1a�[�8 8�BMJ$n�̜rv"Or	#R,N"��<�ұ"��+�v�<�a!Ӷ��%����-���I��p�<�!'�QՂ��سp������n�<ᇠ��I���1�E���P+�i�<��N�J:I!���-X�6Eq��e�<`�R:5�biQr/�P%��(6L�<��K�4� q�	ĺkw�-C�J�]�<a����,�R��3]�0Ȳ�#R�<I��ĭ<h���1c(T��ÍT�<��԰��i��ݧy�TU��`^N�<�, 6�j��1���E;�t��eGS�<IA�.Zt�)e.W�I����S�RO�<�4�Z�!hYЗ�ȿ4��!	�O�<9a ��(�Ń���e!�Us�<�w	O��L�a��8��@bWJ�<y��bh�`&
Y��m��cD}�<�Pb�_�əŃ0�z4��z�<ѕ� .�����<b�D�(���z�<!�j&:DhY�j �68@#jO�<�F�C�0�����T<��9d&�R�<i�ԑ�\�ۦ"��,.T����x�<�P��18�3����r};�ě[�<�cպ$Kz��f?)�UK�BK|�<95HI3%�J�J2f�9't��#��u�<9'��')��x��CN��7��u�<�p��1@�L�ج�F"�E�<�S��[0 ����N���  �@�<9���U�8(v���3�@M����D�<��U��*�*u��^}�KJF�<�D��	_���m��c�^53rZ�<�C�J�mv��@%�rv{�L@W�<�5�ޠ ��Ȑ��F�A��mǥQ�<��#�`bL�+-[vm/a�PB� KY۱oT9�օ��`� B�ɨ?z� Yfo"�@��X� �4C�ɢ�"��
I2<���*�!U$t�C�I7,�(=h��ޟM��d�l�U�>B�I%�|�[��*�ુ��a�C�I�Kmh)�S(�"�X0�EM���C�	6_�t��ɦ%��� �Ǫh(�B�I2d� �8�Աg���0G�c0C��.dc<�r%ɗ
i2�\J��C
yC䉘����fG���3���B�	�q&<9�2C"V�J憔4I�C�ɊVB@�� ��N
T)q�־9#8C�I�
���@�l{�d)��� C��[|2e�F���g�������Qu4C�	�1���`�N��� ���C䉇'���!��(L��4C�¦
�B��*	+��R��x���c��VvB�ɮ|mL�8Κ�:#�1u�ιS$�C�I0&{Py����6z��f�!X�B�)� �`G��6�l�L�,NDP kq"O�ՓVj*B����L�o�
��u"O~DV�X�]�˱a��9�8,X�"O��r��<�"�2���=ۢ8p"O0��u������NP�(`PR�"O(�s�חe0�<{%�
\��t"On�<O)J��G�
�nK@%�O�:�y�8CVQ;6��;צ��GlY�yrc��&�&�H7��6�\�w䋣�yb�R+I�ZT�� YS��Fό,U�!���m5���ՅB
q�Sn[.o~��dB]�Vp17�2������
�yR!��S��HE��#�x�g�V�yS� �0!�4hό��PBi�,�y�/�JD�c��*q1�6j���y���/�F�"��z��E���y��I�~��Am��nvH6g±�y�nκZ_�p���Z�%��K��yBa߬!G���b��T�Re��MR��y��di�0f$��yr�{  ��y�@JyڝSF���:<���y���!�0�cE�66���Snی�y��H�2n�qs��(�S#kR�yr#X�v�-�vDO�Mni���yr�ێm6����U'DĨ�(�-J��y"lR�	���@��@>�iZ�u�
�'�x�@N r�&�CBş/�R��'��(�d\��>�H!n�7"3��p
�'�`��5	�lD�;��د�h
�'ֈ�b�T#c�ɫ>~�̭�'�H�I%%�$i���%JZ�^�2�K�'�8țB�>1$����BxtQ�'�ة�e!�r��)�A��}��9��'�
��`i�'d�<�Rb�̝p���9�'��*��V���Q
���f�l2�'�HaB`CP�~��4sR\�U��'��M{f@��$�TŨ6+�?�m��'`n\R%e�	��A�D]�LD���'����âW��CPn��Um\���'��zс�h(�yʏSR�#	�'ќوAg�8K�������>B��@�'�~�Qdn�2��-ӦõLB�s�'ܸluh��-�Vm8�lʑSʜK�'�����S��#c�טR�� �'�&Hkj}7>Hp��Y�Hm�Q�ʓw*̭�gИ� ���H,Nb1��M���8�/�m=Xd�7gP�S�d���e��QR�ڔ��A2J������ȓG20`Q�h C!��V�*�H0��F�̈xg�
�n�i�@K� "���M	�oN$-�l��m�$�X��ȓ'B��ZQ&�XJD�{��C5~�u�ȓKi
��P��X��̱&di��Md"� � @�?   {   Ĵ���	��Z�ztI
)ʜ�cd�<��k٥���qe�H�4͒6R64<��c�^F�Vn\�c�5��Aߦ#���y�r�7m
����4Tr�Ī<a�O�6-n��)�䈞$�p!��ʂ�#25a��8�D��ג"�qO��N<q�Ւ\�p��4�p�ض�U�
�ǁJ�d�j6�7?�d�Gk*�8λ<)T�A�9lPJ�"�<��+��D���A���a1�N�$yb�E�9�����O��C�H��U"�ݚ9�Z�I/�8]�ÏJ2���/��!j���휐U0謻L��I�; ��cGmT?�'5iR٣1��vv6-D�����%)��R�� l�$*c~q��׼����3�Љ�"(k�`�:��@�D!	�B7����s��-�qF0L�a2�c+��u6��83Dԣ�yC�"ܙ�<�8����O���������ď6;"D��"��%���,ya�>I�� �)h�(�s'b<��`��&��ry�a��$��Oj�s�A�jdZ&��5�X�ƥ��N��OFpю��߈���I�Wz:$@�E�x����t�ʽnL��~�ܺp����6S�5���;�d�Y6G4DE�9���D���O��j��L�i��fڏ2�@���X�t�x�<9�k'�
g�O~H'�7i�]в�~����i?��2M#�O* �<�1&�$3R5��o�WG�-r,܌�~b�^�~��B���ʼ���N�M��Y0 ,�ta�������q���s�/�4#<��&}b�եRbܱXfK˞mv���!؟��dڲ�O"L���$È1�����T ��R�)�2N!�D�<z �  �x�F�Q�(�����;�B��凐7*���2�3�$��^�A`Ώ�s���,�)�!�$��)^�CS�G�i��Źv��b���S���t�z�b�L�+W8�"b�'u��:d�V(M0�@�5ޜ$�`��{5Bh�Z�Qp�%k@Ӝz\\�t
�O���q�
N�H6���ݶ��xr㄀QPH:!I� 벭�� ������ �ɲ��#�J�:%h�#T�����ǝR<]j*��j�@�t����yJ$N����틁y�(x{�KΥG dA���ȰH[�n%/�rȻ��4�#�D*u�� ��([����j�o+��J
5R�D���<
# ]��� nG4�{3�X��Pȡ4
�%x 	�rL#<O��3�菃J=�Y9P�;ZM+�    �    �  =  �!  �'  )   Ĵ���	����Zv���H3�$C�'ll\�Ǔ&zn�ɵ���,
�a W)�>U���=�Ҝy�瞕y�8�	��(���CI�Ap���A�
5�0i򊎕3��qŅ�k�v�H���<���Y�J�$Æ��eϤ�	ɒ�*H����הq%�&��i�a��V�y�`Ĳ;զ���lap��7<�$��,�?Y�2��r��b�D�٢ �[�[��'Z�3ekX�RlH��S�/x��	�'x���i�
|���k�*�"I	�'�ҐK,@�����B������'��m1�[�,\��Ŝ�)$I	�'���3IA�71x����#�L�	�'��=�3P�-j䆕7"�%K�'��|z��üH]X�Yd.��V�:��	�'U.i����z;h,�(RU�,��	�'cpT��`5ʄ��ȇ%`�A�	�'p������)x�����N���'��C��Z�AT��ǦE?jTLc�'F�I�W��'͚�Q'��g�
7"O�5Ag�A=]��� r�J��9B"O��2d+_x*�\�R��p�Y�A"O���RkٹK�ѱv�	�Sɲ�c�"O��R􂎙LxZ���I�t"O�ՀTg]�.��@2ə)4�}k�"O�������0}b8%�C0C3�8��"O^��$ݫTA��;7o�02�k"O�hjG�_ ItB�{��E.W���"O�M���L�W�bdq�'دx��ٚW"OBP �	k�D���R�6�c�"O�0��BE�+s��W�m��M)"Oj�xDE/*E^rsʄ�5M>�cw"O ]���<s���+��=i��0�"O���em��hWņ�f��(C"O�E�N�[@0���5X�D��"O��@�6O�NH��$�j~��A"O��r3'�7��!��m_h
blhv"O�h(qɎ#Y����2L�`~���"O��bUL �t�Q�\$cL`�4"O�٪1O��,0P��F?&�L,��"O���*Č-��1��� w��3�"O�=X�+ׯ�(���ŞD�\�G"OfT��c�j��=�֦�v���ڵ"O�eS0g�)wl���S,w�X�"O ��)0_c���gF�eX��9g"Ox�22�×p�V��%*��$:�"OĹ�6l�r�J��U�_*H���ZP"O��a#�
;�`��jT4}~��8�"O�8B��n?&�KV�ޮ}�u	�"OL%x���J�Lq��Hڕ�@��"O)S@�x��C�^�tކE@�"O��ؒ��Q4݉�g��N1F"O �V�5��d[QfN�l����"O�dbB�<Q:8|R��V��p)��"O�}��!�#u�����+�d�@��"O��ã��K�|@�S���:*���"O����N����s2�ĝ.��
g"O������Z�4�����2y"Oa@��Y�d����	F�3����"O�h� �/�,d�Q�2~c���C"O���6D�r���ME�H}��1�"O���v��7���Hb�T�"O�,�&bK;)��Ҷ"Q��(�zg"O�T�Q�یqY�q$�P+[�J��r"O�@���0j� "��%���2"O��	�l ]��2U%�:�N�2�"O����?S�Pz��ܸRB"O� �j������S
�B�HE�0"O���0JJ�PAX�r$�T���[�"O��������ԋUd$w�:�pd"O$hKF��� a�����ؽ+����"O���5�"X�0�C+T�y	�09p"Olp���يnIB���'�,O�}qD"OB�C,�7w�.�Y�&L�V��$�"O��@���{�:���n�K�f��!"O.��q!ӶgtXjQ'[	u��@3&"O�|�g�9E��0"'�;g4��"O����L
���tޑ)��9��"O�!�
ڣlŰ��e؆���Yw"O��`-*$�	�䕟z{R �1"O$�g���g����e���gbi�q"O���MX<��T*N�C,�r�"O�Ux�hQ�����B�Dڅ"O�̀eY�:�+C���a�*	rW"OZ��5n�/Q>X�K��4'�t#�"O�M	�&��}��M1GhDV��"O��(֫�(IN}c�] �:�"O�����X�Ȕ�i���0 -��
�"O~��CG9p�J� d!��"Oj���h;9W�,�D��z1�a`"OF}�bC�&�< ElIU����"O�
s��2��)�!�Պ(�@X��"Oi@4Έ(2��8#�1�HQ��"O������+8�VP� ��x3���S"O�p�� N�V�S��ɻ@	�0c�"O:� ����%�&�I$�ΤnjV�"O^��tf�+�u��JgO$ �"O�3��?숰z7e�$y��ܐB"OB�b��&c ��B^W��C*O�S4�Đl�<�!���y����'���4��26����'�U4xR���'�0	iH�$k�$]�`j��j��x��'��sN�;!�l����c�V�
�'���ቅ\�YJ'ᔇH�2�
�'�����	�1O�l̒��u����'��T %�ǚ�ʑPƂ�(�d��'F��2cM��>M@F������`�'L�q�u�����oK+iU����'��T�V�Y�z�:]A� �q8�e��'�>�a&��?<������'\,\%�	�v>�`-OH�SgjG�{/~\�pm�4l���"O`���<]�PL��*B�{�@�1���P�� �E*,�'g��)�D��$e��ʆc��E�`T��u��!˒B��D�h�B׍�4i��$Q3��l�D�I(O�D���3?qBl^�GV*aX��Ь,%@!#�e�Oh<�5��3I��$�'g�	���+��ЂS�<�@�Z=���"��'�a��u���pD�P5`<�R�Tkb��D�*��y����R.�hӔ;�� BHR{zLq"Oysw��=��$)v ک_x$�D�>IV��?�J���/n������!Hx�2�Y�^��ℏپ ��B��(W�Ͳ�l nU��/���Q��7�5��9 �T;ǿ���W�޸����cre��q\��!� �59�����T*��_O:$eHɉ�V�QY�'OX���KB�T���e-u����a�ò�Fi)^�	L��: �2O��
0�X�qBMbd�!h��2��F8bƔ��fJW3<�l�X�C�'�nC�,Y�8���GQ<V�kq�6x���y�D�Z�խWX�\#CN��o:��G3Й�b7><b�P�i��sf�C�?z���QG��Qr���`���K>%@��r��i�.�z��l���n�H����r��m#$6��,��ɒ]�IZ6	�$!� ؇#	��椀�% H`D��~��|:������<I��ϺX$M'�
?eF�@:IYq�'kbx�0A� k|�S�%E(�� 5*���b_:��!�T�UQ��Ei!4��9�/(&�<�SV�W���d�<�GI9X�8]�&j��?�N�� ��
��,�3��gu��
��,9�	�{�<irM_�s��!vdv��PE�fW���4��>"�0bfA�A�Dq�|�<�&�ߪ?��C(O��t���%�v<��c�^��QJ���K���,R�`X��8^u��5a��+����O�/���0E�\P�$��a{��#J����i�R�"���g%1�⩐��YĨvo/D�\z�o��3�Ԡ��`V@��� #9�Ic���Ar��A��#}�1nB�A���(��$�`IWK�<i��A�5�J���a�^� @�̤&X�Z礄����F��(��I��8�������DC3H��9B䉘X��$Q6iX�Vؘ�Ԩ�>@�6mC�dJ&i�S��i�i�U�  h�i] *�B����)\O�lX���(�\�x�U�Z:v�� �+�l�.��s�4`Y���:�Q�g�Ơ���?P�G�0|� c�@���a��B-i�L�@ _g�<a�cU�X�\����'u���Go�<�!H�8�>%�T�H�JSFA���b�<A���p<B0��O��#�|�<y� 1ʠ̈w��BiN��bd��_�찳6зwL( �4M[*;��y�ȓO6��s�KR�3<��E�Ǣ�Zp�ȓ���1q��%Q񔔓��� [����xZ	U'�jG&�pC��\H�ȓ8�h!r��q�b7��Q��I��,�@F�r���a#�-G6ԅ�] ��(���9��)Iue߂,���ȓ<҆D��-W���2��dPR�ȓ+�-z�m9%o��Z`Ƽ��ȓ$�R�M܁3Qq�K�%x����0N��#�9�͘4�ZE�D���'4��qwE�9	d,�mi�
���'~�1A�YGo�]y�cyJ"<1�'(0��a����U�0{ڙ�
�'U�U�UnCHw$�AЀ�p����
�'*z��!�N��}sSC�a�8�1
�'B��pcKːd��tRs�̲h��q�'��ԋ��2D��L**��4��'���,T�k�m�RY�K���'�d�c��c��Z"��=�,�!�'v��I�X����5e��*�L��'�&��sM�q6��鐾u��d��'S��x��ԓײa�D-ڝp���r�' ���vLmr���d�<$�	�'���s���h��h��S	\u
�'��|#�]�%��St���W��͐�'�8d�be��!9Z	��\���'=4���@]���KԺX��'ڒ���G.I`@�#AЫ6�0�K
�'5�5�!��@�����6ϊę
�'M�HZgC��}@#@��5#4���' LA���=1,`	`T�$��LC
�'a��@��.9��0C���aCMW�<2�DVd���`M;O��l���M�<��H�N�jmS�j>��qK�.�d�<���~o�0�B�B�-��	����g�<a d��W�Б�C T�u�܍8eb�<��jp����sSR����R�<A��4��g"V/d�th�nKR�<a�	�T�ze���)==�z�7D�I���v|d9�oP���F�4D�� p'�� �})�%�22��8С&D�\(A�sI�$��l܂,��C$D�� ��R�䟊3N�4	��m���b"O��9�M1j��t�2([�g�x�"Od$3�h�'WbA�P�����C"O�ܡS��AW�Q*�NE��"Ot���+��hB�Ծ1nF��"O�U"�Jݛr�I���$�<hU"O
E���=q�H�#u�F�C| (9�"O֥T�ه	E��W�6l`y�b"O` p�!�-fo���gH�U��ኧ [��c���`X������,��i�k�<a���H�� D���WߔN%��P�ͬe�Tt��2D��I�Hƪ�<�A@N��jލ�6j/D�|�Ӥ�a*><8��D����1D�¢Wx��Q�#*3o����ǧ/D� ��gZ?���M�=2��h�"�.D�`ñlњ� hf!�/`ȈHb`e.D�t�$�V�e�Ja��A��x�l�R�*D���㘉�����J�n4�'�&D�\�@��ޖ貂��7|�S7�?D��aV�ǘH/��`
W��}kdj<D���ƪ���!�I{��J�.9D�@��IB*�9���&+aH%��9D�|9���\֝��G2ژ��.7D��x�`M�LL�J��0j��� 4D�0���$VX��e�K�j�i��3D��#��9{�h� T(�� �|��!3D���
��G+�0�`Fd�vH1W�$D� A�*22�cF1�.�ZE�7D�0R��D0��cb����0W��u�<销��$�*�-���'�o�<�e��f)�|�&�D;	U�Ի�
�c�<i�hʬ�����C�|����/�^�<q&iB}��QɆ��j(kreBs�<�g*��H���;�l;y�:U�T� V�<12��Go�	���'6�X�#��O�<IG�	Z�ZaY��ր8~T9�`�<�P	V!z��0�K>rĢ`;��Z�<	���<s�K��I2/�o�<��b�,��A�u�Vڬ�u�i�<�b@�}�Hdg� ����D�b�<��Փ7C��Js@�R�4�f�\�<���	u94Y
��E�J�УF�w!��I�P��`�j&, � @��i�!��%���౅�^��P{ы��a�!��R1v�-��H{�"�P֌�t�!��m.p���A�3�*�s�Y��!��=�R]���I�	���`0�!��$�i !KU;@ִy�7o�m(!�E3s�tH��$׉5Z�[��V'Z!�D��v���t p	�8Q�H�!򤑻<+m��F�C��`P���!�DՐ*2lE
%%I�uWV=�t�R�f�!�$A�4�U��O V� �@��:3�!�Ė$k��	�7E��чË�-�!�D*�$�J�;L+x��->y!�D�2	M�i((�t�_|!�$�3��)��HD��M��PyRƒY
��@c.C�$��w闹�yB��%h��L��ݥ�&%��!���y�O�|�a�FO�	8Ҹ�l�	�y®\0�rpS1	�(��Y�@պ�yb���l������w De�)ƻ�y2�C�"'R�p$O] q�dTY"�0�y�B�,"�����@[��TX�N�y
� ����5Q1hBFlB�*�<��"O,q���%ݖ�!ª�";
(��"OH܀b''8�9*C��c	@�[F"O2m(���4j���A"��<�Z�"OP٦�
�oH�p����C��"O2�(�	o���8}�^Az�"O*<�����W�0oH�f"O�L�F�t���Å�PE���"On�1@���6�8XjG�N�E�>�W"O�L�T�ՠ�K��ѿj��0�"OB̢@�e��9b0H<-�)��"Ob���ٱ$�R���
�`1P"OR����S�j/jũamęr��D�4"O��z׫\�U��tX��ĽU�`P��"OLI "C,,oR��,�N�l�"O��B1KR32=,�K��9�;r"O�xhDns���mZ�!�b�S�"O�H��F�S2��S��`��Z�"O\�+tCþI_�ț0_�8x@�S"OX��PB��9�F"kb�B�"O�<�`m�6x�����D�<
"O�����4v��mP) ���Z�"O2�ZB R�d�
h���^F�4��"Or�� �-nX���	?�!SB"O�h����XE�f��O��Ї"O�1h��>b�^���Fä^b�q�W"O,���	&��i����FI����"OvI@!B�'2��Ul�66A3�"O��� �:590�!"��7Vl��"Oܩy�j��R�	A�	���H�""O�iq��Rt�M�P(ݭY���s3"O]�SEK�R��Lc7
B�+O$ա5"O�`Kr�=8�d3��ھy:p)� "O���¥�ܶ�[��.�,�p�"Op�KC.t٪5�q��vm�"O���)=mm`�䆚X��q "O\hB��@�pT�"^*rh~ ��"O�E)��D=*�4	A@Ւ`V�5	�'�D�r��X*G"�+g�Tm��ܑ�'�Ds��`SL5Td`�	�'���ǪܲY�HX�R-A�MY��
	�'�0��M40֬�b��L���	�'���5��"/�<�Qf��L�H���'L��T�N�R@�@L-yJ0��'��]��� �t��\!tcX J�'L�qQ4�N5r�푰��9k�ij�':�M��H�0���퍰1G��
�'X6��G�)�i6��**�z��	�'[f��R2wB
]���?40f�x	�'KX0j��l������L</9|��	�'hأ��>p�����,�llb	�'"�BgĚ3��Sa�K-_����'
p��U��	dL��u��:Q+z �'��@��J�!f��!%�=I4r�1�'��%��KI�!�j����0g���'�.J�� <�l����,[���p�'Db�)#�'3n4Щ�JτS�z� �'0�h��	�����D�K��!Z�'���j$��i��,@���8�'Ċ��CcS�R����A$��93�'*���%�`���C�(ɾ��
�'��3h�?(�y{ŀ�'��i
�'��}���I�_�؀Tf'u���
�'��@�͈�6���)�lއr�~��	��� ����˩	�����ã0�\��"O�`�Q�;������;3��h�"OD{���9d�|�3ƭ�0  �L�"O���eE �M4O� n�b"O�}����:P��9��]�A"O:��v�	�u�Bd�פ��7���3"O=� !�K: |�v��&XN 0�"O�=��-�,[��Z
Th�y�"OT��gيr#V<�A�i��-V"O4��7�,Sb��׭�-6�����"OH8G<l���w�Z�zّC"O������( +�|��"Ԕ-�(���"O��� �P�{6�Ł������"O<�6�s��و��1)���"O�X�b�1Q�Y�Re�?WǸ�+g"OL�nȇ^��)�?1��"O%�r�ؐ{��`!
�?F�nt+�"Olܸ��&Y���PUJCjv�E"O*��f6LWmȠ'&Q8�	A"O��*��˽u$�A����)A�}�s"Oΐx��.sk�p���D-�����"O�����)o��x&�(��p"O|}zf*�.�ʝ�vV	L���D"OdM�F���x����VJR��"O�mIDA�|�bY��K���E�E"OT@�1
µQi ��'�u� -r�"Oz�sTۣ@5� ��_�$�p�"O���jI��������|{�1��"O�p��ORC����N�ws��3p"Ol��B���#��l3wO,_sX���"OvܑEI�FX�<YT�ϫAb�X�"OT���2c���d/�L0�b�"O1bo���$rW@͕<E�D+a"OE���.&P���,��x� g"O<U�ԇ�����+ԩ��|��*#"Ox�YtJ^�­Ɲx��$U���+!򤒚(��a��ʛ�u�;֩[:7g!�d���TUBİ+p8|zB�H�"P!�$��,o1�t�|X�����!x�!���.2��e�އLR0�af�/G�!���q���J&���!T�a�D�h\!��G5}��ia�e �d@ץ��>!�$	,�ݘŦ�3nuĒB�!��
"���6B
T��"59�!�$3wҕ�̋!J�p�!*Z�!�dʥb�z#�ף;��aY4FM378!�d_ [N���7�S�Q�X�q�eH�I(!���?f�Ub��12}.9�A1�!��O8�&@�	Ta�uIWk���!�@3"QrH3�.%����(�!���r����G�	�<-����+x�!�dQ9a����ahXT+�T�A�� �!�DJ!�td��-�K,��g
�'�!�d�
NL$3�+�0'v	:�b+,!�$[�lWz����<V��9a��?u!�-��t�
�V�(�K@D!��؍S��(���G���
�'̲�!�DD�C.�P[@,�&@��玬!�D��v4���K�,�V"�M�$!!��D	8�|m����!�U�I�.c�!��E�z�@TX��G�D�h��n�!��q`Z�K�"�{��6H
'B�C�I�-�t���dėr9 1Bs�
�Y�B�I�2c$�tk~�M�Lݲd��C�)� �a�� ϐ62��� g �w�D(�"O9Kq���k�:�(dM�.���"O���2�SE��)sM_��ً"O������#�j��o��4Sz( �"O();�r��m���o3��"Or7j�4R���L� Z'$���"O��qUaؠXU�0��+�<q%n��%"OLD6��i (s��Mw��p&"O�2A^�3d].b^��"O�������}�J��D�]��Cv"O��I���&��p��cX�:4���"OT*�
V�w�Ԩ���.�
�"O��yD� 
�tUrp���)�L��"O��;d�  �P   �
  �  !  �!  n)  �2  �8  ?  `E  �K  ^S  �Y  `  `f  �l  �r  'y  i  �   `� u�	����Zv)C�'ll\�0�Ez+�D:�DlӞtB�8O$����' �
�e�� M�A��A�EN)�%@�V�Ag���HY�푸T��@�a�9	֎�?��o��?��[�_�8l{���)�n��ç[#Y���� ."}�f�4(���@Ғ4�뎛�.t����O��2�J��NDcD�ԁ:f�mʃ��4}Ѕ*b��ȟ�S�	 C'�p�$��M�6g��?	���?����?�%��"�`����'\*F�BP���?y� �ք���iL��`�����?=�	���S���_4ȹA���'=�J�$�O��o���'��zd�''�A"b#��K�#U��rI���4f)��4G|��i�F������j�t�u����$h��>��'}�'�$�-x���ɟbaz��#C�x<�gg�i6Ό���'�R�'jr�'���'��U>��;:��S�bHyp�Z�8���*�M��i�P6��ᦽ��ΟQց�M��'�?y�1��X͏�_�ʀ��!#�����(�X�O���L
���[���1�rm9�N
?��K���!��)�S��/�ƥg���l��?���15��E%^�X�zU����4��p�����Q\h�ݴB����CA�"���2�@�!�Z����@މ�ѿi.6MK�rD@��,�R�MsV0�a�v����$u��8�4��f�f��vi�yo����ݓ
���� ��Z���;�/��j2�9#^G?>������q�&���9ش��"~z	��E�(�l	����,w��ř�IΈe�d	�Ҧ�68���D�}�愐�왹)P�P'W���#��O^㟀��`E!�%��,��1L�����ğ�?����?�6�H�zk��?	�Bdt� $;�B�H!L�O��?������H+O�(ĉG�`V�����M4�Y��X"N	b�  �M]�p	Óe���2sMB�s l�S L�M#U�PcTtPУQ�xAF����[<
�џ@�Q �O��dFny���;m!�q25	��sT��U���?����?�����0O �+a	�$8f"��,A�89���$!��|��i�ށ���O$��r̂�9;dM�! }�����%HS���jb'��!hޘ�qf\b�օ�Q��"�yr�ݬP������_x�bfE[��y��Q5�
hP�TfΕ�R���y�nZ�x��<�"˾#q������y��=z(Z�B� K,nGn�!Qn
�y���/i��i!�	̀i���[W�V��?iAAAi������PPN�W$�YQAM�)#IBB�	'îЋTJZ]��Y6�7��B�<���l��.�~�U@ԇ��B�ɀW�uC�O���AkI�O�&@p�'NR�4fN�R-�P��2�lЂ�'L2����O-oc�͉���@�!Yv*Q��	�4��Yy�V>�Χ Ůe��#Wb����T9t�rEB���yE���r��G�	��	-;��KF)6�b�Z$��ut�5K��0<Ў$K-�v����)$1��F{2j45(D�1UB�)�0m����I���!��0���0?��EC4��YW )�4m!��򟈅�IH̓�ָ�����ߞ�{ ��/L{h����Mӝ'�VrӒ˧:H�|�v�'S�$ñ9Y@|9�ȵ=q~qI�J.��T���	ϟ�ϧ97��q/G�e(
d��f��`ɵ���	~� (��{�l ��z�1���s!X�S@��#L8e�0C�=l@� +1�
c��H�s�L��lʕ�A�%�Q��RB��OfAlډ�MS����svf�Y�&8huK؋;_��)O0�0�)ʧ�,��K�^/@$�QN�8���?y��h���l�I�N�s@�>̼�� (���4��9Pb*��6��'���/�=LJ�W�G0{ ��K��	/!�3/�h3��:��)��ˬ�!�$�=c�� ��gC	����D�!�DO8WBZ(�hʎI,���nV2m�!��8ʨ�"��&GdMk&*P�)�!򤄻4q(�`e�w�V�"P�Z:]�Z6�.���29��?�'���b�'D,`m��:�e�:7<5���1B#5 ��G` 	"2d_
��)���=pO<�̄+\X���!C�0֪&q��,��#�'*'0@YSh 1o���|ZN�(Y���;�~�[w�Q�	,$]�vA�L��d|yBۅ�?)�����?���PN�a�M�9����o��Yϓ��O���"�� r�*��aK7i�"y��X��P�4UV�f�|�O��]��H���y���`g��
!VX��5�و��ߴ�?Y���?�)Ol��D8Y0�\�pF�9���Qw�
a�H�PU�𡈔G�~�X��"LO���3����M TIȭ����<V��(�ږR�x50�������l^�'WQ�rrE�H�e�ȫZ��C&߻9Z�D��A�'���'���'�ҟ?1:��V�c���Tˏ!b���h!|O�b��`���0L8N������F�<�?�D��}��Zy��E�&�&6��O����5��(8�n~��)��.�a��O��d�)���D�O�dKe�~���P���Ё�&~�� v�0k�<�BEH�0;�ҡ:��'nx1ǚ�r�`Y����޾6��x'���8b���^�um���_��(O�A���'���r���D�'NB=� U
E��42�i��6��ʓ�?���OG1O���-�6�q�&�����Q�U����̟��?�O�l����l= D3�@4D��p�٪R-T�,�B�7�M;��?i����ׄK)�?��A�A32��Y��`�U-_�?��U�N%J�ܘ��>����3's`x�ƺ C�/�Y�.�O�z	Ex��)7pΈu�F?\"�R +�6^a���|�H��D�)§}j�h���V��-��c&~��ȓ>�,��I�(�L�:$�H�4�GB0ڧ�$1�����d��Rq�$M��Xٴ�?���?����&m޺H���?!���?џw���r荳r���j
\f:4`QD���?!�P�xذ�`����Ʉ�V�	�G^��:���e�3ݶ�ɠ������ZHx���dԇ54Z\��G�-��Is��<F�D7��ͦ���(eӜ��	�Q������0���F�,�#J^ǆ@����OԠ�#�3���?iFx�e�"�`8�� ̯n��L�f���?������OyR�'����'��	 j��pYB�H;�SC�*L:B�%� p����\����PQ^w���'7�	��0��󑢗13����v��
Cf�O4��$��
��,'C���ȴ+�1�!�Ė�����I:��̠юN�_���B�'����$>y�DpX� ړ�6�����!~�!�ކ#B�ȴ��O���$
"{l�'j7m4���G�*�n����I�'b�-�֏�,�8)�qFW�����Ɵ������������$(DI��)J���Q��n�B�ͻ�@���.��a������	 a�ه�I@��܂���!H悀��	BGbH*r�Ȳn+|�������S�˂�vF���ɮ_Y`���ަ]K(O�X����P��T��NQ�%���]����|��D9��[�)�T�Ї�!~ݸ�f�[ٟ���Zy��i>i���I�~�2�cڞllBƅ	�hHP �IKy�ݬ+d�7M�O@���O
�	H�_(����镊V�)d���+F{���OH�⁠�O`b��g�$��$-BEE�`�Z�2 ��8w��I*�B#<E�D��`u�-`����H�!�`#�����Q��+&���%~-�X�%,
�`�-���B�82� A�H�	q��b+ի�4�?�w�
L�6P2�=Tl���P�gO�lZğ�	ş0" ��+To�A��ԟ(�	�8�;#[�8�ߊ&���u�N�!�<!�n\���0Kރ~O^I����i��J$M/�	�^�����ӑi�ܸ�"�1,Y�t�R(Fk2�O"I�$�'s1�1O�ܡ��E����AP�Tp��"O���RgZOfV��+c2��[�d���4�ܒO�����)6X����N�ny8�ӥ��*Ud�ݪ��O��d�Oh��������O���T�o�!##E��>O��Cc+�� ��<X���  Dy�B�#4�l��D&�j!d �<ĩ@@'C"�T['�ڱra��)3O�3��3��,L�������K2��UkF�O�\�R��9A4���'��.�d�OX�d+�$}>�Q1�	vS0<�q�]�u��a+"�3|O�c�@��Z1viZe�D�P�spYI"�,�$�ۦ�ڴ���K����?q�P]�,Bq��:4j(`A`!���?��X�Z�#���?Q�P����˺��di���M	+e6�{�L�P(�c�1O����Qg��R�Ԃ#�JQn:>,� ����5M��Q�8x���$��>��'p�7�O�0x��0G��l��O"mP~!ӥ�<�����(�p����G7�Ѣ�A��z��U�XF{��d�s���`� �Bj>��j�>B�v�q���ͦ�'��0&�o���D�<�)���dQ0U�R\V��'�b�����9���OJ�y���>M���W�a�\��$�S�.��YXB�@Nd����)�`��M�'�8�r�_�'����ե��?'�P �)J�\�(���Cm+$�gC /_��	�*�J������4�?q��� /L}�A펪P�����(��'��'�ў�Ӝ!�d�"pG
� ����g?ܣ=���&��&�vӪ�OX�§�}���a���-���7i�OV,+�g#�i>�<	���w���9 kM]�
X�AC�c�<9 j�9��Dj�MM�*B�Ed�G�<i�'�U���e��E�v�����i�<!��G|� ����]�����b�<��,N�X�^�i�)��A8�,�F�<Y��)&,J�(]�w��u��@yB���p>9 ��,s��SFeA>gdp�d���<�  ���φ�k�ʙȢd h�z�R�"O������H�3jԀ$�Rm`"O�0�ȍ����s�bW@�����"O���Bl�xY�K�2g���"��'sjA��'�0!a&G�
�d����_3z�J
�'�zՉ��)$�0�O(ܒ�	�'A�� Q���z��`�!��+�µ��'�,�d��.J�����P:�)�'r��Vh��s-�Q�0K���`��'�T�т)'c�
�� %�
q<x���*�Q?���4)�$�S�'�+s2�*5G<D�dH��j_�Qڐ'\:��)��:D��)G%�� �-�#h��|Ƣ�I��9D���'LӃjxb%�4Z:���`�h2D����˦-��y���S�}�.H�ah#D����W�3��<ItnS�?��k�@�O����)�'_sl j%d�3t�\j$�G�h���'�B��R+�{���C�V�Kդ���'ЄHB��3��8-�H%�5��'������� �<T��Ŕs
\��'�hI�e�S� ��r�-��P��'*����.�N��ӌ]K!0��.OD���'1����eZ)b�U�c���t���'�.���VS��D]�e�*]��'���(���+b2�ԙ��ԡ`��AA
�'W���\0�@��qŋY��Y	�'FDJ`*
�$���Kp�R;P�*��/���#�ZUXP
�\HXSq��
&!��?�^dydb��� �bvL��W�`Q��Tc���&��(�.�r�h�5:�xP��[Epjw��l�Q���-mL�D����Ra�T9H5�[P˒@�Ї�a� �y�*��U=�f�Q��~UG{������*ī��.$2U��F�	��rg"O���0n�4Fd�P;�7�b�#�"O���U*K�8�N��U�ɷh3�H!2"O:eZ�(ց'n��0���M�dL��"O�����Ї{��$��DZ�O�4`�"O(�
q��64����b	�d�����'���������>x:��sM�����4�΄��$�䙢���ZN�i�C� :	.̄ȓU�쉛�E�]ր$�W�٩.mD�ȓ?� �*�~�sբ�,V��D�� 8U�դ��>3��#c˰�2	��V�̢'�H�v.��$�I8��\�'j$D��1B�I�!)�=�B���C��9��8���vA�6M��-C�
��mM!�ȓ0]�a�;��p`WL�#�04�ȓ]�flQ#��r�yq��D�<ufl�ȓU�A��H���� P(Ֆ4�Ҝ��	)Kb,��d
UQ�)�>ԅ��GrؚC��E��@��P5d�mP�7��B�I�4���\��p�C�͖`��C�ɮJ�ҍ�s���@�Z��w P�G�C�I[�$�b'�E(!sVĂw��<C�I*s�2���O�2�*�,M5o4�=)c%�\�O{�jC�%�n�S�΁'�f�X�'�|Kf��[���!G�o�8 ��'�q�ΐS\�h96�A 8t��'��=���Ȁ]4��q6H����{
�'D��C�ږ9���pƔ�f��	�'�xi�c�^����NP�$lc�D�8Gx����BP�"3�8i�.x�%NpF2B䉿g`n!K�A ~� $�5iL+
 B�)� �e(4�%7��˷��\D���E"Ol�Խ?2����V2���a�"O��c��{m����3�ش"O���`�фai�`�fD�^��	�Y�X��o6�O�P�!M�>�(M�P��(�Z���"O���ELJ;�6���8c�-i�"O�T�ѫc���!��\7��(5"O:��򃇯����,�V�.\+4"O�I*����EGD���[::  ���'���Y�'����$H�rFd����C�fX�	�'oh�*D잏%"X����	P���	�'&�x���,��)�DЊ��	�'ƹ�� �u�R�rȗ>�Q��'��0�nR�J�&�pf�N/0t��'L�T���/E�V�����8I�!E|�fV#���<���M�5�|xp��
�^n���B"Oj)1e�K�0g�<p���N�$m��"O�5c��?����<?x�Ma�"O��A��ظdfD�5��l\H1Q"O�A�n�,�,)���U
�Ja"O�	s�5e5�����P�!�V!���'>򬨉��S�OL�%'�O��h� �Jd|��E�����%oޢ*фηh1��ȓ>�(4P5�0�����1"����dTz�sF�$܅V���0���ȓo�<��Ō�P$�Ʈ�H�J}��m!���A$T#)l���չj\�,�'r�YK�:���ju�&�rUڴ�U���P��D{�����7��j��B,-�B剅�����L[��ɯxṯa�"O&=h��B?I���R*M�Q[9��"O�1����7/�.�	R��!X��Ks�'�N\��'7�9I7��&|Q���t�tp��'q��6l�;HK����GZ�sj�՘�'�Ω�W��=wC��3��lY,{	�'��Ҋ��{Xvأ�MFO#|��'��p��nL	p��%3&�7���'��-��.Z+z}�.+l�)[���N�Q?5r��šH�$q�$m߰H�vӷ�"D�(@���"��|Y'cI�>�M�`�5D�����@�I`]��d��S��K��4D��S Zm��ӂ
� &84t��<D��Cbב|�r���I�OV��I�=D�t{ �u+����͇2n���7O�O2ͪ@�)�'3A�ф-K�\�� �M��h��D��' �AG��w)&�� !�W<H����!��=e|�Pe��ta�F�\�<�����N+�!P垀O�f,H�ENW�<�7�ũ&r�$c� �=H���.�k�<!���'_�{�2�Deh�_y���p>�#%�c�!����l��|����v�<QrG�:�@�VcV#x��ySV&�u�<����<��y&"B��T�Dy�<Q�a͗F�����QE��R0 �K�<�ԩ�62�1�A�g`<�qV�Dx�0��쪟�`���#���5�_�M��l`��"D�̀W� �X���I߈*h ���!D�@��U�xC 8ː�(8�D��"D��P�"Td�P���lu%t��F�y�n͐9��a�צx|2M�!��'�y�L�8y/. ����vf�z�c�9�hO�(��S9�����c�.<�
-!����3zB�		 }���ԞX"��rf�5cu:B�I�	e0�{�iˍR�੅ѥf:8B�)� �8��6ZUDD�A�O_�X�$"O�d��I��rW���!#G"u����C"O��"�-ȏFR�@��͌.�t����'$|�����6l�.���%���J���IX�ȓ("TD�E�7^w���/�'c�I���z,�"��(I�8�*���	<*�ȓ5&�lB4��-}�A¢$
G�͇�yE��C�f��Q�&qqA�Z�k\�5�ȓ�<�@ï׫l��8�J�|�'P�M��tk�����v��Y�튇iV�܇�`֠�h��/U0���Y�-�
���/ɀ@�aʱE>y	v��Q����ȓd"�uHܚtfb0�W%�(�.���.S6��5W�N���l^4i�$Q����Z��ɄAȴ�b�̙J�H�B���3��B�/Y�p�r���"Di&�c��A�B�I"S���
�k��8cP��!X�B�}�,ܘ�G>*���9w똠n�!�DR����D�0R��GJ��8w!�DD5n;�,"� /�.��b�� +Dў��b$�'��l����2asp	Ƽ7�B�	:�L��U�A�4���X�1_TB�I0��s�ȓ`���/ȮTB��<ސ���fz�`%�F3[i�C�	5Ąh��0|F��X_I�lZ�'��4LL
M]F�Z���'�����?<:YGx��	�%zݩ��1S?�ZI�S"O��Z���4^��YU� �tg*C"O��ۅJlpMr����F�"�"O� �7��\	�5I���H|%'"O�h� c5M{�䜻�d�����C�Iji���I"-[�`z�&�4W7�Aqi�O}�̫J&�$�56C�4���і-��Dm�����	��K䉘���͋2$Ӡ�$��	*@f�	������� ��c���=�]a"-<���ͧ?�r��-8[�Μ{���<S1:F|�bݒ%�n�ymQG]�� u�K\
��Y�17n�#M�tB*1I�a�u�'�r0��8��v-=��֋Rq��i���/0R7.� ��I�x��$@g U��**k�9�c�� k�Oޣ=�'��ɮ$�.U����<-e��J ]�`^�ʓe ���i���'��S$Sq ��I�ӄ)Ǿ�X�b.�3&�V١os��S�N.�B�R���$�v��G��z���	�!jh܈2q �B�l� @�@�#y�G0*h� �!-��9�"�:ܨ�:�dŋ�F֬Y"��{�v�P57O�$h$�'R�7��nyJ~���y���jaD�!a%$ZX��C��y�jڊFK��Ё� Xڛ�.��`ў|���	w�-���Aj�\t#��D�QK��d'����OVCC�h���I�O��d�O�U�;�?�b�F�-5�	ۇ@�)Ukl��uχk��<���'[2Q+v@�l�<,�͟���Mh��6�Z�J��/2c<l��B�$$�2��2�l]�O�~��E�}��@?�l��DM�1u�\�#͈� ��I�b�j���O���8���|�I��^�R��_,*�n`�� Ph<�#E�-,F�AH]X;��S�G�1�?!5�ɖ�M����'_ -���A܆�ke�X6$�{�?d���	�b�x,,����IҨU<ܓ��#D� QcmK(<�X��0b#$�:!C>D�$���F�fV�*ffOc>�6�0D��Y���^W�9F捐`�`�$D�4���s�j��!-��Н��"|O<}�V�>���O�:ˬ�h�Id�=�b�V�<)֠�3����#<`|m�r%�J�<�%%�Y������C Q�,���G�<a����%���R��{ef�n�<�兓b����T�sb�,��i�<y��O^��!2"э(����e��M�'D�DxJ?IX�`ԓL��FG F�fQ���:D�8�&�0�5����B�!���9D�,�ƟY�i�^�j���Y��9D�� ND��oօk���Rh�g�MY6"O���f1*�V��%�"d�D"O����H���� ���1�iȚB�"<����O�ܢ �)Q9�s@D���@G"O�i)6�H0��aF��`l����"O��I�fFN�pi&;�<��&"O�|ӍIlnd�0#٤9d�yHA"O�)!�3� ��b��FM���`�'�L@� ��N�|A�H^5y�r�Yf�חf��(� �+�"�'&"�i��I���'v<~����cHX�R��#���fV,cS����l���'��d! Y�r^��5c�qB���V*�*��r�c�2mV�AQDB&,OZ$k��'��KĎ� 6E��J +��`v~ � �'��1�'D�h��&�3q���d�0��tB�'���P�P�]S���r���g���+O��n�ןX�'��E���'Z��'1���ST���h�>���
��^:V�2`�8���'�b̉*h��0�")�.�r��'��I�  ����Ȯ(T+L$O��	צ�\z�gԎ�jI����rrT���N�v�8���$;�j`�kIywQ���w��OR��0��&
Z��a�֫neHxP���a"�D�ON�O��je#���bl8Ċ̚�&���	���hO�I����4 ��,K5�6ݢ��Q���tI�:,O��d�O���O|�'�?A/OR�YeD���k��7x�c�d8O�=�U�K�=|"���.n�J��l���M�K<YgM$�iB�.���+/B�,��bl�$:Hn�ǟL�e�<�tA���L���?	���<��Q�q�.es�kɈ#k���H��H`�L��4�?s$M��?��'�J]2��M�;A�s���%�YFh�i�0*�C愺n��[@��'�2�#4O*���	�?�	�<��X�Li�����f֌�B�T=3y���	�410FN��ϓMo�	��ם(���zW��A�	�V�"��u[!ga2E�?a�]W�%��?�I���S�Ի���k-r����I/<�t-�ф��?�VWП���ERH���<���Pnz�"Xw���H�ȕ&=g �ҮT$c��	޴�y���?���=���O��':�$#�Y��H#��ϗ;�z����A!�,��>O�P���'�2�rݍ���<���jnZ8?�^`Se-M�Ixi �*_{�d��Ʌ6�MC�'&H�{��i�~6�mN�s�6M��2�zj�6+�1�`�T~@���VP䦅13X�<� /���4�	�?���<�G�J�|"s*CNP�	0GH
QI�.���MK7(ȯ�?A)O���O1��	R�!j�!'I�zP�f��e��B��K�� fBܜr� e�$�@���7M�ON���O���O(��O*��O��d5��XB!�[��:d�E�C�v�֝oݟ4�IDy��'T�O���EĲ��S�7gL���n��X7�c��'��Ey��Þ'x�C�g����DB���y2��es�좵�He�x���
��yB�ր��ED���(����y���/�x�D���6Y��ߑ�y"Ip��Q�Zj:D��,E�y�M� s��ih�l�L� }#���2�yBn��~+��s7e�s�PCL��y��A6�!�Fe��,��hA��y2Ԭ#�V�#�
Bd�>Ԙ��O0�yR%D�_d�9r瘢�`��B�)��'���f��V�OcB,�&��_��{a�P�t���'M��6�ڏo΂���$D�\ {�}�.ѢĔ-	'�[2n3�s���v�:}ʁ�ڕ~��m+% �$kHQ4ȅ!��PV&ڽ$E*��r�K�tHQ��WJ�#����ϊ?&���� ק-��X�R>�M3s$аÀIYWG
�C���A,ݳ>W"Q��BFȡ�ަ"���
�]j�ɴ]���3����d�6�@�&B�I%f�8���]"B3�4���[O.�C�Ɍ��-V6�a�CI(kP9�"O�	hG'�F+8�7b�!�0q��"O�L���#��|�d ѩ	����4"O6ā��	~�6Y�a� 
�b��"O�4�ң�5�*�+��R�t\@A"O���m��_vt8&1ܪ��"O��S醲��I��~�Y�7"O���f�FU=�@v��,w�8u��"O�z����V
�H�fg&%��a
"O*\
wI�O�����"}��;`"Om���u� T��JR7d�l�"O� R���\� 7�ЧcB�Z*|���"O�T3Ϙ+����i�/'lp��"Ohh�p�͕?����D�G�l�`"OƬ��-����Q� Y�X��Ԩp"O}YT)H�|�M[��I�����"O5�Q��U"(��7��eݦ�
�"O�4��$AY��+� }�bP#"O�0p���s�VN)e-�P@�"O@���*n/��c�,8%@0��"O��Çi�&�dpp�K�/vгs"O�y�aMԭq��ѕ�,`>�h"O�H�GJ,H@EFk[�;��0 R"O����N�/���錶z�*E*"O����,h�{ah,����F"O�U���(t����L��3c
��"Oɩ���8��z�K�&3F���"O��HW	�Q�|� ��4&}��"OFUj��Ɔ���(�!���2"O �(f��,�H�pՉ�1ע,��"Obh"%���|��ibӟ �R��"O<q2ph�.n�2�Ǯ�N 8'"O@�cDb���f��K�<=����"O�Pˈn�Ј"��$�� "O���Tf@�fO�)8���iuf@Z�"O"���`�L(.� �bĴk]�8"O:@�F* u���ҧ؍WJjC"OV�8��ܴ=X�����]�D֬�v"ORw�A�.�b$#�)r1 \��"O�T���3#���`1k@�(�0���"ONT�Aɮ_o��ȲI�'��#�"O�<�%���
ᠼ��*ޮH��9�4"O������?5��p@��T���H7"O�숳�S�+v8t��N_�r�2�"O�ICE���T4�p��Ȑu�6"O�@(�)XX`�&.� 7r��"O�9`L�f�<@Ǧ\�,H�"O.;��"��� �l�{ڨaQ�"O(y˄H�Y4̘��CK�P[�"O(��lȟ9��|#��8��4Ӥ"Ob�Q� �1��qJ3��'Ͷ "O�\� ��nL�u���~��� Q"O��d��*3��sh���"O��p��i�F,��h�a�l�a"O|h*�мI��V�mUd��"OԬ襏��w�d$AAU'd8�)B"O�`��m��3:��1���l$�͉�"OxY1�k��xZ4x0��_�E�\)�u"OHDۡ��9j����*]�yE��Yd"O,��&�ɵ.�~iW���p[��'"O�ʆ�˴���Q=fo�M��"Ol�q"R�oD�݀���?��I�"O��C�;��@K� ���t"O
p P��T���ؔF��Q��0�"OP!I�Ɓ&v�`����Z�t�}x�"O�A�+��=� 80 iõ?[:��"O��ࠢP/g;<Mx h_F>��p�"Or�[�aT�~��!�1&�6 Y���"O�*bI�lP� :�BY�O"}��"O��p3
�K"E�!��x�4��"O^�j��+,��e��aH'�t�"O�ѰW$�j�N��o�>�F�5"O����B�dan�k�H�{�c�"O6���n+k�����N� 4���"O��c�
)O�p`Co���Q�"O� L9y3�J�jc�h�4aЄ)E�e�s"O�T�ga��+��[3�UU@�\�"O�)�SI�ȓc摲t3^l��"O�K�ã8�ĩ:f�L8)�<�F"O�hJ��L�y�@��P#��d2��Q"O :���=(:4#�Qr� ̚u"ORDQ�a�
l�a�P$��u�JX"""O@�␁݈:��f��	t��� "O��VN�2*��d4HTDo栒�"Or�����x�6���O�����"O��� �ݖDDt����D���CS"O�ؓnK�6x(I�iA��L̑�"O���"]1.� � �jU"/ά0�"O� �+�;`x�*RɁ�P"�-��"O"y:��Ι��L*�M�$��"O�ԁ��B������ݪv��h��"O�YX��T85)�$0�� 
�D��f"Opq�5g�<���`N�}��i��"Op�>���;Ql�?�<�Y�"O���a�W�	��l9��_H�\�@"O�ɩсɉh,����cf����R"O�h�E _�U�P�"��(�n��"OI�ǟ���ds0 �)4� 8�"O(
"f�e&�� ��[z0P�"OpY����B�)KS,��<�R@�"On�#��&	�^�)ӫ�:oi~���"O8�`�� �m�ri�r�
�,��	�"O�Df+��G���jv�Ρ�Tk�"OX�ے*��
p���&��.|�"Oƕ��/�6���E�Y�!	n�h!"O,� B���x���
�sp���"O8�ʧ��J��PP@_3\�B��d"O��"Dō$u���2C�-��t��"O&U�f�C��L E��:��l�w"Ol�" M
	G�vx����q��p2"O�胒�3^��rǧހk�6���"ODY��"�~�J��Z�|i1�"O�Q����g*�c�̋v5���P"O��ꆃ�
wk��!�ެ���s�"O���cEǆ�d�	��Ư%C���7"On)�ӏ>]H��v"Y�*��(��"O�^\2�+S�>� ]�Ď'1�v}��bZ�<����,8����F?k 9�ȓD֬���#����gf�]\F�ȓpZ�|9�ʁyL�ak�
����'�\h��V!s2*��f��|\�C�'�z�&#˝vY�c��S�rˌ���'�h-C��I拉I#�q*(�9�'��*O��f�Z�$�1e7����'R(��� �!eb�b��\�$���'��x	��P1� %���)��'����98�����.��4��'_ĵ U��]1����.�=�|�B�'h(��.I�>�=It�E 0~M �'0\���F�H���``���`���'��%XRAÎy�n]��� 
�x�i�'�!�uH��C><C6�Z)����'))���E� �e���{|ڝ�
�'� ��U#@�D���b�͡m5�M
�'��!8��7��`j�2X����'V� ��&�����[T��<Z�'���;%g_����C8`�{�'��m���%!�����,S�90�B�'��ey�%_�w����uB׃)KD����� ��7�T�tr̔`k>*�"O�#��b����蛮��2�"O�dK5���Ҹ��f��F�2u2�"Ol��7��<�]��ӱ�* ��"O� �vD��0Li�b�'8W ��"OȠ)���`z���KA'<��"O.�������"-�K�&"29�"O�Hf�
xȸ(�����&��H�"O�
'j�*/
u �+L����"O�u �'� B��i0�ԮY=v�d"O Ak��*�L��N�^,$,q"O���	c|�qK�?��YV"OȬ���S�!��UR��"6���"O���ԍ��4㢠s\)xD����^p����O'�%�oژ�ȓ^.��@��1�D����}�a��/O$A�kN&��ScO���Cq`�S7�ƨN�F��뙜{��|��c�.�X�B�7Z"<����EI� ���|s'�8��DC��� ���ȓw+�\��l_�n�<�C���	c�̅�%��\h�L8Y�F�r7��k'��ȓ ?T�s�&ߡ*7||�C�:M�@хȓW�ݫ�C�:FvP�����'��!��<ښ,[�hE>V*�� �('��h�ȓJ��� L
3�
����1b�]��&��m��.ݐXM� �wD#:��I��W��e tɁ�(L�,!�+҃N��̅ȓ��Lf�J�1S�� f�F�����B��LU+��#uR	�d�ʥdX�m�ȓ~��(�& j���+->�ȓ-e�u�7Q �Z� �68<vY�ȓng�y�qȅ�/�8X��	�;E��ȓ�8�C$N9wL��aA`�7K�$}�ȓBu��H��@ �|�'��z��r����낟>%� S���N� �ȓ�T���,B�U䢠 4�ۄz��u�ȓ2ބ�0̊�$��E��+T$��G��X���$&�ْ	�p&����O%�@WkҵH��=�"L�@���O�����,F���C�	0	
���}w��[�ȁXa�d{6��5��	��7i���/�<���H4"�$@��C�>ip�e��̕+x�H�Z�n5*�2C�$:��@2.��|�T���K�\pC�I�4ިK��o`)T�O�cl�B䉽O�ZH��ʵ���%�L�% �C�I�VT�	`6,C�)��Q wk�S�C�I�/�vr�p���0���ddC��"���A�����X#���ϊB��#|{O6NZ�T	�㈯h)�C�%IR�81�I�����䃆6q�C�I�&i���1���^@�U�]1�C�ɜ	�p�	d�B;'�H��Q�+�B�	�F\��dރxy.|�$�B=V�B�I�@z�x���O	-^ ���(4�C䉘Ɯp��o��>�������5�����ڟ:�D1䀃�]SD����7�$G(7z*-)g�t�b�뗫!,�!��v1��.�:`�@@�!�d���y��ˍ7E8�����F�!�d�i��إ�d��T�JH�!�� x�,d� �|���a�ׂw�!��J�=�����4C��IQ��F!��Gb~x� &.K�%ac��rl!�� �X���]&�Ѳ�5,�Cq"O$�*�D�Xs�D�l�
�'�j�3'�6#)t�`�V>ou �
�'-.�R�Ƃ)t���CCd�n�:`k
�'˜!�f�+�h�iGO,p{���'��@�"�<�
w�@8ˌT��'��s��FL��`����9%>(#�'�T�jtGQ�M�j�+90���	�'�	 i�c�&��ѧ��~8�'���"�+Em��0A���,8�',Й�p`����<��W|�1i�'� sa���TȺ����W�9,���'�8((��	
K�^Y�'g��+��Y�
�'1�]H7D�_7�@ڒف ��B
�'x@Q �!E*o�����]7V�f���'�fԣV��78��āɟ�cSx��'�8�� )�l��� ɗ�H��`8�'i��0�
8E(r,Q��H�����'����ȅ�n��d�ܤ}:�
�'��| v��/�\14���v��I(�'%X<P�g!:.�K7��i6
Y��'����3��Y �X��4�P��y�ɾ{*8xC�9�`��d��y�G۴A�ʠ���+��H��ǫ�y")Yc��wDǺ"�Q�f�R��yrm39ŭ@7�hQz��D��yb��4�N��[);��� U�-�yś���,z�.5/�\t"d���y���x{v���oa@,���3�yB��BMС@��0eܡcRf
��yRO�xn�kg�SHLa�́$�y��N�����
H��,;QE��yr�=NIJ�Ú|�����E��y"�L#4����Ўs󆅳ćA�y2��0B�����[�c#P)�d����y̙	�|d��/W�*�a���8�y���q�������Z������y"�� �8	�E��'r�T��#��y����|�p�K�S�b���&.�y"��33�~�22�K����!B��y�d��7�\�W���{����%�1�yRC�`�a��I5���f/E�y��	�J٩!쀴���� ��y���Hc�YG�B���h1�⛉�y�$��Y$J�[���
��5K�)�y��K�Q  &�-VhrA��A;�y���"�T�2@��4Tr�5XCș�y��Q�E
L`�"흾D��#b��yR�U	b�M��J��'�Mc���yr/U�i|a����-�l�Ej���y�E@�#|��P�Mi����K0�|�ȓ��ԃ��+n���F��!D��ȓ)�H	P���4Y�(�k��,�ց�ȓ+B�X���0J�x'�I|�N<��4*R-v��G�n���OT��ȓQh���c��a�¬�Tj/YH8���|�6e��6]��"�!?�%��#��u�E�8	��J�(˄C�.����t�i���c�$(���E���ȓ�a���!<���OڪȈ�C(D� ����vDb�+�.Wg2�ѕc:D�4���67*��AJ��efN}c3�#D�쉄F3$��"%�����&D�<b��΋}~�@��w!�yѡc&D�� ��a��3��"��D� uP$"O��glD�e,��F�&�!��"OBa{�)�tAa�)L<��`*O��Ph�p���0!�SJ,��'Z�a�Æ�
E)pH��3T�
�'s�a�v P4�T��q��u�R���'�jؚ�ǡlĂqM�T(��'!�`��E�Za�`W�Ŋ{�'�ȸ��bΐu H,�P)H�`o�:�'�J�K@�~5C  ��d�%��'Xв0�*�4��Sƍq2
�'����&�.v��ejRb�u�B=h�'�<�@���2��%��apҝ��'E�lɱAÃNY�����Uo�����'�ޥ��Ȑ"=8,�1`d��f�X���'�Y0R�� !�A�h�1
z(Y	�'�rY!�듫G��,1g�
�� ���'���`��A�'�~̛c��*;���
�',��A�߱bf\3"�ߣ/����	�'c%Z��ߞܠA��#�#w���'�f�jY!�D؃LÇR�C�''�Ժ��Q (�f�Pv)�.3��
�'��q3��)lZ(�FS�'�X%J	�'����j�%�����._Iy��'E�yb�	�mQr4+�Ǭ
#�8�'fИG���,Hi�^ �p�k	�'��lr�[��*���A�D�Z�'l>Ѱ���8�b@��#@�V��'!�%�U�t�М�4��E�r�'���6�Z�JZ�� �!B���'��A�Da��ZD��B�o�X}9�'D�H��D��k��=��(�
xM̔�L>�� �*�0=I%���xn�@/�( �R���Ö}���a'�,>���0�#��m�<����4M�MǮ�oH<�$e�"�e�A�(YZ�!��Yz�'i*Hۆ�X�<t��%���<�bT0��~��(0 1�!��r�ʜ`�l�+!����b�D�K�V�D�S���p!�K�Z�,�S��MkbEr�<�r������P��r�<�̄SI�09�Ǉ0%;ȬS�$��.;����|	Q�����g�''$�D�*��2�K����	��v����S��s�32�F����� B�0�f G\ 0!��'�h9#S#X9,��أ��1r\���D�v���pB�V�2؂8�C-7���'dX^�kb�I Iݘpa0�D�8�B�ɣ&��9�qňA�X��)C5o�<h��3X�P�p��82U�B�1�g?�%c��74sW&�Ehz�C��|�<��dBn5Z�<[Y� �	�z�6� ��@�U�����1AҞ��h�'J�c�O��yw&Q�ņ�b"t�ۓc���RSR�N�)8��9�ԅ�K�BlHb #O�S쌰�7EM�0�a~�� '|��%Aާ,�z��#㗗��'h����m_�3��F�$9����t���ڱ,9�x9�"	�qW*��F���y��\�S�y;&���d?V���#�"����4폗#rX�H�k�	8�6��,�y�c_�Hj6��Ŏ�F�֐xf�R)�yb��U��S�O��S
��⚫Vƞ6mP71J�huBQ7a?@]qѲ�x�D|��\�Q!P��G����M���=�g阺c�޹���r��iӎO "�Qv�Q lT�q��qm�u��M��*W!�8+���2%��X/��?!�U#Q��%9Q�R*1��P;aB]�)�=vڔ��)�x��L�A�I;B�!��["%J���Z�b� Q�� k���U*� �Z��Y���O}��KP2|f����/�>v��	$"O�ܳ����h�l�A�h�=b@�I���]yBكw� ;7,�v��d\8 �MRU�{~�;�هCu�~��@�1ad�5Cƨ����\1 �l�b.H��d����3.�Z7��@1�x�1MW4t�G|r��;kF�� �4��O5Lz� c6J��c�ƙ�5�)=D�� z�ɖ��S�Qˆh&l�q��O�i�ƇJ�p1'��}��0:��
G��'=����'�Yg�<�a!����ԆI�ȡ���`~��L� �A��'l؍C��s`��x@@hiDu�
��.�ر�b�7X3b�!����܈�w��3e�!�Ē�<��*Q鑙q��	��!�!���(NE��:Bk�;F���3A�	!��M�cJ�р�}�������C�!�dŘX-����m�,a���)<!�B37p1j� F�wn��p�C�+!!�d�0���� ?I�ȥy�#�;*�!�ʣ<�0���43zz��D��!�$U-�<ܒ5�۞X���??�!��� >	2�#� m��)vF@U�!򄙛q,�(c"$�G�ɋ�/֎^�!��^[N��7G��@$�u���,R�!�$��4�Y2Kݩ &JHR�$_�e!��P�b�RX� T% NE�����VK!�D�o�RL�� ��5.;E!�DH�X�Z�pr�ӫ(Ȭö�2�!�d�����;T-!5�a'�K�!�U97�(��"�
DG�I$
�!���a����A8Y�rp��7y�!�d"E��a�O
�0��{SgһR�!�D�
3����AOaM6���V6+	!�dO�yHе��G܍>���'lÂz!��No`eг*�0@�v8bgAT��!��H��1�O�;x�Id%S�e�!�D
�<�����gè�xA�S<U"!�d	�����1S���ku��	�'Ab�Jf$�=EcpL�"ƁV�ZY��'�����</�i(����"�,�A�'���Ƭ˲J>��Y�[�����'Nd��=:4"�C6Q_P���'�XL�˛���,�4>�RK
�'�`p��z�iBV���
�lP��'�Ppa��,o�6,b�Y���$��E�,qI��5�Za��!�m�
m��-���↘�
wJ���)�� ���.�ڱ�͘���딊�M箌��o�
��`�D�94d��)�
��ȓ���w��$8k�L۲���`��D���X���["�!�i @�D�ȓ[��eYE��*C
4��e˻f}�P��eF,`���,�h����d�t���OH�A��y�h��)3@ͅȓcsi�)Pm���ʯl%$,��]ilQ�%�4[�����E�vF����q�1�aN��C�X	4fٹn�l��#����,���!`�1[	���ȓe�V���b�,lPK���(n�6��{���� �$h� � #JM:��ȓT�V��1�Xo�N� �jY�	�a�ȓZVH(����8iT�F'��tޠ-�ȓye.ț��M�UNjѰ���.�V̅ȓ ���G 
��}pdd.?Ϡ��ȓ���H�.YXX��_%WB��ȓ}|t�"�zR'�F�p�6%�ȓk�,*�%�$Kb6 :���	\H������@%��SO�M	���<^?0%��b���ҁ�%�TyT�\�v<��=)Q*V+>����H��.�`)ã�s�g �k�ㄹ]��!���,V�bB�	9X�ꥂR�� c��_��~C��$��&J���8���1Qܢ��"O� "�	�HK�YȈW� &S�荁"O�qhW) .(D@(��ߝm�N@��"O��)�˩md�P�e�5a����V"O0�h$�ծuB�Xk����J�:ek2"O�`��F�P���1F�@. 0r=""O(u�P�
$2�HO�ؙk�"O���&� "���W˅[r���"OH �1g��1���sf�62���;u"Oʁ��+>V<��"��"`���hS"OH�y�M6A���DH�~�ġR"O�Уe@	h�ah��J�:�� "O�aHDiªf�0,�$@�$���S�"O�@��M�4��3��NB��e�a"O`LSÉW?Q�ġ�!�G�\�b���"O0\�W�P#O��(Ԩ�F�����"O2�Z�zOb�p���~$�T�d"O�͛R耄(:8K0�;�e2�"On�����R��L��,H �V"O��b�լ]*q��MJ�|-!�"O�u`�ĭ��m�f�&k�^�h�"O����<�^��chÛy�l��"O�I�uK9@�@�����\nL�i2"O(h�f㟱/���9P/��	?�Y@�"O�x LBF�~�s���	��,"1"O�%"�(�ea�.:{���"O��L )�`ԃ¢lJ�1�"O�1�F�A���yp"��!YXx��"O�e���\Z�y#_�n��"O�(q7j�1O����R1��%�p"Or-�Q@��4��8kd�^�����"O�%��ER��4%H7*@�<�&l "O8\��.�8lѤ�J�)����1Q�"OX�P���I7���(ԦU�t+�"O����F�)�U����U~�5IB"OH$'Ȁ�C�0�Y#ºUw��"O^�x��7#L|k6p��2"O(l��L��D�0H�R+�5@2H���"OX����Xo�zq��
 ��p�a"O`-����'q��X��	N�F:�"O��#T�t�yJ�k�9�<��
�'���I��2��LH��Y�+�����'���X���z���W.m�'�ܑ��+�;	q��;�AɊG�ؔp�'�(�g�F�%5r����F�L���'����UŖ~Ű�X�C��Eqz�Q�' (�c�/�|��ìF�3��Ek	�'������50�l��X�B��x#	�'�j��'S�,hB}�( <4
��r�'Z(e��GwU� F����s !D����<6֘H����iw�	�C�	��L��fI�2�2�;�מ=��B�I+g ؜xQI�(���Tہ3�B��*>bx @͆&M�� �	�7�JC�"
��(@HG$e㞡��@o".C�ɍ�T�H��n��8h J�)��B�	/��S��2>p��"0"ٿ�C�I-�>�jS&��I^�P����ҬC�7f�RY��ͱ
�:�B�m�(2�C�	/̥Z��
#0���B�(ŒC��9 :v���,ы��`�c�f�^C�I&qR��0R��&D�@aq ���8C�ɧB��E0s��/!	[�k�|��C�I�"i`tς�r�e�+AD�C�ɑn�>Z�"�>zu��(A�\ΞC�)� `�1T@�`qFM� P���V"O^��7���x>�\�7n"�(""O0,�����A��)B,�5i��qv"Ot��ԙwb tX�LJ�E�|��"ObH����"H�l4�P� z�.aB�"O�(�� �ҵ��k�u��`۔"O�vJDAZd��3b�M�"O������_�À)R�6�x��"ODx��mG�BY$������"O&�2��k���	�>��Z`�Ro�<i���#������'K���C&�l�<1��35�l��G
b��(��l�<�mŁ�@i����ISԸ�Ѣ[|�<!Q�5��)���U|M �P�<�4�O�{cP	�I��u�ԐP��K�<�P���O?��(�/S{Р��g�I�<1�"�>ʾ4i��ݪI���UGE�<Qרx�f܈W�W�
QH�fL�<���� �(8gŅ~���F�<�Ō��&��i��왩K�P=��#��<���F�M!d(��/=(|�1Cz�<��`!�&�W
�"i"�� �S|�<��ʈ�x�����]��Aӥ�Mx�<17�Q�vk��)�dө�>����t�<Y2*;
���(@�v��0�b��E�<����VT��kZ"�9k㮟�z	�'���ӧ�3��뎪wɮp(�'��<�V�7`����l����'�T���e�4_�@�ۙb9�8�
�'h���,����5ѳ�M�&�z�q
�'�ܑ���%;
|�+���.-Y�%y�'���y�K?S�X\QB�ƕ(�R���'1��ucR	�XQ�f��%���p�'��EA1�
�,��& �-ıK�'���c���y1��B����M�
�'��Q#�58���#TTp�X�z�'W��3�ػ[����$��
|�x�'0���tA��� M�E)�$�;�'\���K���Ʉ�$90�'h�B�hFD�h�	t ն5^�	�'w"89#�5*�"3н���'��t�׆��4fE
�`
p.(��'DЋ��q�Q�����~X��'���R�)�	(P@�A��^�TMq�'��� $ML�'����t��!��AB	�'��4�F�n�T��>E�<r���yb���H2�Q
m������#�y�,�tI� Gl�u��{f�0�y���+>��i(v���b�����y���q*�T�uCP����g�_��yRN��,A<�� Y�s�.%�Vdݱ�yB��5�J؈%FK}�f��(�y��`] ]��l�t��)uB��y���[ʸ
(��l�@��ɖ>�y��Q�jL���X���AE����	a���O#6H���I�a���2E,�2FE���
�'��1��n� T��=rQ
�'fdix��]$7���T
�*q2J�r
�'�6�w��n $����; EʅB	�'����'��6d��xia����n9h�'x��k��Zza�� ��J
0D@��'�\e���N � �u��D��'�:İ�V(�&��lB*EpȡR�'Y�$�gE^[����4J�:T~�I��� ��K�&�8(6N-���3�A�#"OIy��3 @[1*d\��"Ov�&JL'G�Q׃���>�؂"O�!���T�z��"�^���"O�sT�v��}1f"O	3/(��"O�ur�[vh�ѱ��^@ !�"O�l�G��%(����� F���"O4ls�al��ɩ�m�{���+D�P�� ��<Y
�3�)ۛ$�	:G�5D�Ȱs����)Q����S|��i3D��j��Z�J�,�@vf�Ph�"��=D���@�Q����������<D����K	mђ�P��,T �G�8D���lF3@ ǐ�A^$��!D���sᏒ[F�t�#ɍ�ܡ���>D�0�fS����Z�G�f�1�u�;D�T��ϵ��G����2h�'�4D����� 
];t�N�eD��x0�0D��dk�2;���X��C�l0 #0D�Rw��#/TeI�!�)�p+�)D�b"͵��!Q�	#8V�	v�"D�ȫ e��BC�i��*f��X�2�,D��P$Μ-���UY憍�~��B�/H^Y�6��;v���@%a��REB�I�C���f�C�3^���	��`�C�I?޼�zc"Ӭ��,��l�s�C��)��y(�	�taS'�<��C�I=��Q��"��B��I���I|�B�ɣ.fDj�h[h��5�Ï��ys�C��0ZV�kQ�*F�=�P��)L*B�I��t]�P��A�R�H#��4;>B�	7:�L��'M=KdՓ�O���C�I�}#J9�Bh�����N�K�B��W)d���n�a��-st"Q�;�HB��-6r�m±� �H�3-A3��B䉾$�,��D��+��#�����B䉼:�P�CG�.
ʽyeH��B�(@�}S�L�(N���m�?TC䉄:��`e��+i�]�aVSMBC�I�c�Iz AQ1����&�7y�.C䉂\*��h�KQ?wB�'N'uC�7sT5�زi�vh�0��!{�C䉭~X�H�Rk=>�pXSC��=[�B�	�Ah�e �@�Y���I#4	�C��,�q
D�j�=xE+rC��4?���FF
$9���ˉ{vC䉜P�$� ��ΓCs��J�K�.*>B�	�m;ܙJ���*EӾ��!<�C�I$)�6`�2��pF � aZ��C�ɫs�E8W��d�<��GD���C䉼V�Tir슴{�:5�����C�ɛ�@2�Á=&Gڡ�0���VK�C�ɂ{�"��W�uM�iLK��C�	(�H����L?�V�z�a�"O�C�	/{5��k�jD2f]Ka�"v>|C�Ɋ?d�1S�lL�!��!3,Ԕ3�
B��F|`C�gC�N�9A�?=�B�I1�ܬ�G��	\3BH� �4m�B�	e(1�#Q5���!ؓ$(PB�I4P%�K)�2v�n�AīT�@B�	;6�	Ж���NT$�ckw7zC�I�V7�ũQ��K+�p)�(P	"GB�� .b��!bFŬp�%��(L�DC�I����\��R��dC�)� $djR��z�ӏ�-��b"O.;cɆC�He��(�:���`"O�`��-ʘ$�|�P�GS�$��耆"O��"��M6y!60��G
=3��;�"O~�S�㓤6��m%�� q
�x�"OZP	��38� �"��p&MX�"O�9V��$Cހ�àS�k��0"Ov����ʢ�Tk`�<e�3�"O��������Z�.'r�Nxr�"O�����59 *� �dB/R�NH��"O��%>r���[gP~E�""O"Q�a��2=�9�@& �#_�0�"Op���0of���Ë��J�8�"O���0H�*�|�U$p�TEB�"Oh���kR1�Α�3b�!����G"O�����%;KF��U���{qr ��"O�)G
�q�X�+�/�5\Y̍��"O>03V*�s0���ͪ=`�R"OJ�J� O0�h�J &_#.��"O*|ä1�>Ts�P�,�U"O\yIU��?���Y�nN!�&i E"Ob!#��	��țTn��\���u"O�ɂ�m�nF9c��֢_rQ@e"O��a�jɀ?J��1�;x5�7"Ou f�C+�a�e�һ7���Z#"Oe:�cB1��]�Ɲ���Pxa"OƸ��
��\IL���ŏ��qB�"Od��� �+�Ny������"O�DPCG��J��U&%��r�"O���$+��h�PwNS���ha"O0�U	��Mc��� ��2�PH��"O��8��/����,�����y�CПaؾU�&N��p�S䄓�yR��,]��D80+�ƙ�y���_C:�s��U�йCƝf�<I�V�;�2! �V?J&f�i�j�<Y��ã!Y���'ҁ.f�9 (�n�<)�@��&qx9cqʼyބ�Z ��m�<�D&ѥP��Ɇ��:O�2�:�q�<!��bf��AwB[5 &z��c��w�<�3#9�K���[~��b,�N�<���4������ن�0cd�TL�<qfh��T�.(��ɜ<c(�l�lEL�<���	pq�vN$�$���gL�<���^�I\ܬ�c���1�Z-Gl�<I �ҍ!G�aY��  L�%HÆ)T�ty����}d���7*��������3D��֥۵+R,k�l@8�) �4D����K��.J��ԁ��?ݐ!�"+3D��1Rf��|#��ܗ#pyr0)3D�|3!���F���(Aꙡ�4	��`0D��Ѡ�ݣ�`�@d	S�bAT��qL-D��B ��9
 X��Ԡ&�n���5D�I����Gf:��͏����!n4D� �ֈё��<K%o�>�
9X�.D�`j�ʘ.B�61�!����.D�a�a˾'L�2׎K�+��k�	2D�$��nJ]�B��8�ش���,D���#eH�h�T�i�VL��d\�y2���x���Y�����M�ye_����DJ�)nxqӃB��y"��i�z�r4�N�'�}[�"��y2��.�Tٱ��E�Q0�eݲ�yB̍%%B�Xk�a�(�f5j�+�y
� �ر��&$�0�墖�$ԩإ"Oh�YC�k(H1�塏2u���#"OL�"眾'8 Q��]�.I� "O����K�k��-�Ï���xM��"O�"J
^:�:�h�� � �t"O���'K�aA�!�g�|���"O�r.� Z�'%L��0"O����f���f�!aD\�B� �"O�@� =�.L1� �&��H��"O����	��L�O�51�F��A"O*�s&h�9���	�`?�!�P"Oz%
7#�[����fE{9,۔"O��1pl�1l�b��eG�1& B�"O\�a���p���e��(m�f{s"O\�끤^'(��l0�ɛ{���C"OxX��kے-��{�DЧm�dsB"O*tA��ӼM���0�̘�%�Z-��"O2��J_�AN���A�(3�`�:a"O�`*%)�3��E�jЏ˔=*�"O���%����� ��	P2b��8)"O� c"�W"�v0bS(όm��])�"O@�� /ŵb��)p'��9���zT"O�d�Sl�6a"���F���Q�"O����!x��Y�!�`��k�"Ot�Xb�X	J.�bA��D�R��5"O0��&B�$=��o�>MN�X�"O�H'��,;ν�� �g.�MZ�"O�)@$	B5:	�,h�!� �x��s"O�\� �-lx�(1��Q�eLHd�4"O�5� O�.z�� ���N;Đ�"O60�O�R	��"�k�Aª�	s"Oh��V� �'�	�A��$�(���"OR0��>t
d�F�-�VP2B"Oά+J��\��m�u� e��TrU"OX�m��tI�pC�O�J����"O>��hٛ�C���,E?�R�"O*�����a�����ȍ�\�
�kf"O�eeݯAƤ��sF��5��"O,u��9w����F�<3 ��@"O�A{�/�=�բSf�<��y��"O����>�p �J�V:�1�"O��el�23��m�G��:|�����"O� 
tX'��@�f��}����R"O�(qC��l��uI�I��D�t"Ov��-�5:t�Pb�C�8�b��"O>�3�P�0��t�}*�xpq"O�LH%��6�%�DaC�|!��*�"O�(��!<��T0�
z���w"O\(aw ��2/Z��/L�2�B�@�"Oz��֫�]�^�OE</���st"Of� a�>�p%�5P"O�H�%I�z7�)���i��qw"OF�   '"����a�y��9a�"O�zǫ^�fZ��W�ܺ!�`�z"OBL4GF�Pq��!���8)0�"O�3��� !�b'`�,F�<}1"O:���l�fl�aR�ۮ:�B��"O��5�ѹUneP��ʞK"�̱�"O>Y룣N?[���P�_2p�D�Rp"O*���)U�4�2�#װ
��a�"O��@Dff�ز�S$��� �"O�c��*�
�`Z� v$P��"O�`A�叅N~�!1����/bV�"O
�Dj��$#�1CB��;aL&��'"O� Ĩ	c����U�ߍvH�9Q"O�e	ԇ�v���:�ʈ�E/�xW"O��˜Lu�X{g�_�KxʘQ�"O��rv+U�q	�j<	q�(ȣ"O��u���F��� �	ޫ(���"O�� A�O�X5B�
Bz��"O�i��O?{�lu8�ϐ�mi�I�"O�!����R�tȳ(� �x ��"O���S�HQ���D�D�(�"O�P���L�l�HR_�U��!"O\�2��ȫ}�.����ؖfN�`��"O&L�H�B�m)&N�$wMT89F"O���e&
Ki��!���>1-��"O`AB#j��b��q�� E(bZqC�"O�}��)\�����"v���*"O�a�$�V������6�bh#�"O� �ŗ�4�8��=tĩ��"O�iv�?c
p�Ce� �Ĕ"&"O��җ.K#Hx�1��"�4W�V��"O�����A�V��J�6`6�2�"O��8ÇȂn�������D��!��"O|h9 �Q<2d6y�­�y�P��C"Ov9����-�����H�R5��G"OR�RT�O	S�����1T�I�V"O�A��OCUz2`�cd�I2�"O֘��HS<E5t�����"�8�"O�@�N�?��ۧF�Lf�R%"O�E�@���drb&G1W*Q��"O�E����:w.H����Ka�r=�"O)ɔL0L���A惫h�~eK�"O֕ȗ�	12T�Y� �U4'�d�#�"OΜ�7-��}�J,��ʁ�}�yц"O(�`FS�X�R��V�E{y���"O6���L�w0�$�3���~�d1S�"OB���f�07-�)��׫x���y�"O�4 �R|�\*�+�le\��"O��X�H(:���A���F��"OlD��H4k�8a���nd\Y�"OX������.}˶��7��j�"Oj��F�^9`�`�A`���,)�W"OfU�#�ƹs5J��P(�)��0$"O��sq�� X���)�	q���d"O,�S�D��6U�qe�T�O���A�"Ot�'+S0�J��� �^ ��"O����)&d��_+��P`D"O�QBPIN�`$���L;�z�(�"O��	�g�$CQ�!����_��,:�"ON�:�k" *Us��I��|=��"O�����8<���aO�7E�*� "O^��'Β�'�,���Ȏxj�"OtS��
?S�XaQN��&��"OҠ��f�n����H�2�b<�b"O�4�lQ��HY�5 ���rĈ�"O��a�W3�X�!�(Up ��""O���U�U�*�f�%�ܑm2Ÿ""OЅX'�>e��4H��iQ�`�"OnX�7�A�z�*]Y�盍xE�""O.蠃��Dpt�C���E�	��"O����C�&8�H�Pȁ�	�1�1"O(��.C���0�K1����1"Ol`��"
(3�8Ɖ���h �'!l�Q��W"ȵ	e��&aQ�\*�'��<�����;�r8hOPc�	�'��8tjhs��S�ڳb��U�D"O� t���NP\�M+Tg�8��"O�U�`	~W���+:z�.L:r"Oh�ʄ���R2j5d�l@S"O�x8&�΍c#��1��s"Q2�"OM*��S�i:�qHjlѵ�	�����Wۛ����%Y,��SfM��:i4�3��C�A$qO��4&*�c ��/Q6�UYQǐ�]h0�S�O}ƍ���LTz���&�/dklt��D���L�������Ph�YT��o�8HE�L�@n���W�%9(#=�QiBޟ81ڴd�V�'L��&�٪��t�2+e���J߬h����<E���7~�Yq���i�Z��:Y�����ɦe�ڴ�M��gt�*9�C�J=��
�b?9�DۚFT�����4�`lO�	""T��!�H�t"p��A9Y���)G�5)�@dS���/v�H����M��>����Ԧ�BB ����i���f�i� 3P��t%�CUA+�F�	q�>�*J�T ��V�zY!+�h_�c�6݀
fB�'J$7��O$���yB�d�3�H���k�#He��Jq������hX��a���o�,JG
�>v�Vqs"<ʓN��lӸ�O���}�2$�����KF��
̓�/� ��$�?&�H�n�EX��ht� 7��l9�&j|�|�aЖt���1P���x�aB�`t�`��7�6"<ɱ)�"A�.�P/
���U���!s'M�d�I3c#��p@���O@Q��X�*ٔm�0%:�W�VG��@�	�?�v(S��?a��/��gy��'K��i�"H8Fg�J�윸u��z�@��#$�L��C
!���#*R�xv��b�KŴIś�gz��O
�i��˓>��$CJ�]v��s͖I�HD�	��fR0��ϓ�?�%-��\>�T�R��5BJ�gà]���v�[�*��s���ܓ&�#�`���p�$�.��8�F`��3�!b�&�$�:�J��+L|�	K�&P�Q��,���O�t�㇚�cg�=k7�ݛsi����lU�~H�m���ԗ'��Q���~b�/�U�p0�"�/t�$	q�<��,Bp�|����qi�S�&�l?��i�7-�<�dG�QI�V�'`�O���q)�NΑ;AG[E��h�{��'x�[�	�r���R"ȑ�&�S���|�&��n.�maF-��>9*��A�'�����m�,�X�2Շ�g��aR��?Mɀ*��8a����	C�h� �xP(?�B��`��,�MCU�i�2P?	�UdP�2H��`b7:Z��Y#ϝ��?	�����'r�ɬr��tA&��	#7�	�Q� K����D�Yy޴�Mo����CجKyd�P�0r7m���(oߟ ��ȟ<�!D.���֟�mG�I�f�oJ���cW�W�HA��.T	3 ��<q���ɦ|�'� 4zb�ʍf��L,q����_��m3Q�\��@A1�̸a&�0m�?�`��ID������!<QE�emI(q0�����h���On�DϦ���F��Mc��j܆d�f�7�hFd�?A���?�"�$�T��5�r��/|�Uh�4E�Q�@��4��V�'�~6�O���kݩ � '$�J�srn]��!�����İ=qĬ�   �   �   Ĵ���	��Z�Zv�
�)ʜ�cd�<������qe�H�4͒6R64<�bʄLL�V.��Qtx���T�&��8ɳeK�~�7�Ȧ�����y_�|�'i��7O�8ɵ��==@�zamZ�B�U� �d � ��aԯ��'� ,%�`FL%d���o�)e~�܁@EP�53��A���+,��G���c��V3�>�*D`#�I�9"f˓t-CE@�>�H�{�lӶ5�N]r!׮6��<��>$��$Sb��*�q�����+�~h��XS�+�����J�n��5��.Y�+�����'r@����ܶ^��ԟ�!�G̛=rL���c������4� �0#�8������s���h#��0�ª�O>$�į�=���#]��kQ�N[�ܔ�WL>~.���ҋ�^}L0@�Ǎ�z�qO�!9��$ۼ9���#ؘ ��)��ƒ�!��Ex��V�'�x%�'DP?�FԨ$BF�'F:ysO�p���n�qO�A��B9@Jh-���ע73���V�i��Gx���m�'.x�������|I����SV������'���Dx©_J~��	Q�YAC uQ��x5(D�����Oz�y�B̚����a�j뚠P�D�8;�5Gx2lGJ�'��	���4�A�1N̨�B��-$�b�0�V�	6f*�'l�5z��׼
�i��Ǔ�Q��Ÿ�'C�GxRdC�	�~©��3��(2h�W��!�'�2d�m�5OX1����q�4[�c^i}�����x� Y�?ɷ���T/�����#P�	b	�K�y�#<�%�*񤆽f�7-)�M;p�J��O�������OV�Hb��){�Hձ�hי1b���"O�Ⴖ�  ���If"O�L�� ҥkf��#�٫D��:�"O�%!�$�>8;�Ё�Ɗ�gxa�"Ot@i�a؇2�b쐠��P�.a
4"O&y���86eL�� M��Q1"OZIq�C6���1�`k<�Z�"OV��sa�1 i�XS���-i:���"O��c���/Xk:�q�nF�+��"O�E!f�<i|��"vM�e24i�"O
�KN��B��J��8H�"OH�������#�_ 9�dI�"Ot9�������B�ׇ]Z��E"O���H_�X�E�@�S�W�DXa"O��B��]�$- )r����^�<ໆ"O$�x�D/m<�AfB��k���"Oi �8F
�"�O�o�2��`"O�iP3���P�c���T   �
    �  /!  �(  3  ";  fA  �G  N  IT  -\  �b  �h  o  Su  �{  �  6�  �   `� u�	����Zv)C�'ll\�0�Ez+�D����M{�	�<�4B^��H�P*@���Z��"F��B&�0Z��!���L,;�4`��>LJ9#&�Z7�u�
�@��t,����I	*~�<:e&bp���e��/@���\������9L����N��c�:�]�J=���SП��b�D#qp�h�#/Q�N3���K�l��| ���?�L^�d~F�;�F��֪�E.��'j��'��ʝ9�T��䙨_S��D �i�B�'
ft�}���?��c�/�:���?�e��0'�����א<�2US��3�?��w���'g�	��T���������`��6k�n�B�c�*tr����O�'���l�l6j�	� %�Phi��z�&r�O#<�'"�x��#c����(�]�ˆ��?Q��?1���?����?i�����e�)A�g���i��#Ҡ��}���O�pl���M@�i��6�O���%Y<>�n��Z�@u�I�XYn}��_��Ī���ZV�DD{[�>���,j��T'R�Q}B���͘I�d��Z2Mt2�R�G���mZ��MC��i��$�Of�u�P5���a��(O���!!�l?���Eh�b!��34�<���	~���!�,�P>�YSC¦����mZ�I�إRL<u���ԧ�.֑Za�]2"�x�"���M3��i<R6-ֻa,<��Ĕ<��[��P�q�R�c&NU�h��!�*�k���ơ�c�M���T<'�Rum��M+@�i�d�wV]x�PC��4)�)���"�F��/�cr�Y5M�:<7��:�)f�ȶ9��їG϶MD�d=���2O�)��*��p�e�~����B���?Q��q��L�a�i	��* ��,S�LY�ph���,4�p��<����?ɚO�,HE�1**�q��-���?s%ƞV�� ����s ��c	���0<	� G�q�l�0OR[�V��4a��h�P�^U��cc�L�����D�I6A�����O`��'����#��.RC���<*����?�������Ot�D�FdZ$�7��E������C�|A�OR�=�'_3�FB���(�&�0)���R6��
��7m2�I�c ��?��'Q�E #�Vt[jA�&��o;|�
�'�8�1�^� f�XE���g�
�[�'� ]b'CHQE�K�U�8��'��H3�b���,hc�(�}�<��'Q�(���UP:^d��a�BMTD��'aV8�q"P&8����N�2�H�h��e���Ex����)TJ����]�!�<����<gxB��4y�R��f��(��8�V���RB�V��+#E,d�P�JP�I�B�Id���s&a�D9q3�� <'�xB�	�hh���A ��V1�B�	8s^B㉤DC��c̎�J����C��C�H�R�ry��'�2P�̗O��)�����d�;AEEZ *
TԪ�2���Y �;G��2�az��7"���LN�Z�H���#�rԚV��k�.ĨIHM��Q��6X�ў��4e��.=�`s�N3a� �ҥA;<�&����I���<��O�QRΜ�d_�[ׯ�-Zb�!�'��y���ϲ2��[B*�]��f,�"hG�*j�@�	Ԧ���4����0��Em�ϟ8�S�f��"�eʈ�"b�I� ���Nyr�'��9�(�D:CVFXy�o���"�%(���m�X.6]���W8]�ax��R ��E���?y��"�!�a�H���J��^��h3�CB��S�H�)��TDyB�M�?A��i�
7M�O�lɥ߉W�zIƀ�.�X	R��<������(��\0 ��%��yD
�/mV�5�A���O�}zT�i����I�FV�0��]� U��1�x��O��b�����`�ӟT8�R�]kXi�e�Fa�Q��6�dI�%�';C4̰�+[�t��}��GwƼ#ȼj���pl�%rV>D�ȓ���K�%]S�a�"c�#V�`�ȓy����WG�R|����=�E��p���&[g�t��Rˑ�}���@ߴ��7�
X3��L�hw%]�3�ȈIco���D�l�6H:-9c	 ��P�P	M9,�ʧ�ұ/�DN;�x��U��9$,Xm�'�^������nB�	B���}� t���]M����'��㪄�p�:d0Ԥ�E����o�剓/o��:��O�D�O��x��^98���5��sg�ɱg�9<O4��?)�&��X����+�c�8h;�vy��{� $o�w�i>��xy��U�#|N����E8�"��L��0K��d���OT��<)H~�����p�f#ȐM�I���TI/ ��
�
^�"��0=��f�60����媀�X�T�2@ڡV�T�뜲M��,�F�H6!w���Zy�UFyB Z�SU��(ġN&����TC+=7�������P�d���������|��_�t���u�G5}Y.���͎�/�^���7�	1;����2�E$B(0�W��h�Oαl�ߟP�'Z���g�����O���!���q���9儛�so�9h�`�Oh��K>(N���O6�S*F�p��:�)� 43�
D�t�w�l΂Aj��'뎐��DB�{rơ ҏ×m� �H���&axB���?I2�|b���])�l8���Tx�c@�7�y���_28�.v_�4⑪�,L������3�?�e/�u�(�9�ƀ!�.���`AO�	Or��ݴ�?a����	ҏ|l���~��� t������T
sbD�D�O�9���F�T>�'>t��Hok9�rb�+Pe�� �OX�g�)§U��];d���
���V�,�X�`/?�Uh�ҟx�I>E���^33׊��AI�$>��*����yB뒆^.���Nτ`8�C�ó��O�DG���K�}�E!�蔢Ee(�.]ۛ��'^R�'H����I���'���'��.�qTQ*PO�|k
�d��\�1O���D�'���.\�z�hL�b���4��eۍyl͠�0=��h�M�\	��{ܤ��'�܆��xؤ��Il�g̓�ba�!�p��MJ;vK IQW�'D����M�0i�DzoĲ�0�ū�<i��i>�$�d �hҊ_��LJrG���#���������?Y��?Q����.�O���l>Q��Ȯt���Wǅ0KZ���	�2tB�	?C��Bejβ;J���B�#�Vh��<��be��;�d�q��:|����5��7G΀�$�B���2�F3H�$���mT�28���b#D� ؑA��j��F�L�L��� �D��$��R����MS��?���A�yEB���K5p�X/�d�O�����O�d�O�]@&$��O ��HL,5c*�]'d�Z�pr�Q�j��0E�+"����O��z��� �2=�,X2I�{-e�u�ظ���iEǇ�&���� %՜j���(Ol*R�'�z6��eyrE�h���r`�'H�BM����O��DSHF����ˍ]N-bC������$�OJʓ�hO���Ƞ$��Kb\���V��,Q �O,�_��qj��i���'2B�O)�����'��H� �.Iu>���c�4������'kR�yZ��T>�'�Z ���9�jx����
��	b~�K���O>	#b�q�TU:J����S7�-?�4(�şT�O>E�$���S�$�s�o��:A��*��y"������ K/yc���e5��OЭG�ĦZ7�X9PL=s����s�/om�F�'���'y��;����e�'���'��ʷ-�8ӓ� �,A���N�p�1O�����'��DN.SW�!�� l�3�y�f�0=� K;&B�Y�*L58"�(U ����;"���t�g̓l�	���.��uH�gΈ;�!�ȓZ��%���#84���;*v ���Dz�O�'��)���
nC�p��L�OH� �E� Q�D��'�r�'�OG��'R�O�j�Y 	�&)�����}�~$�� �<5N�I�ֺG7az�N��9"Dړ��!*2Qqτ�*(��å-+�pHa��)TL��N�q��Gy�O9��b��Ǎ�� �C�"Ha^̱��?i�xr�'ҕ|R5���9J^���ɢ�GD��Qg�'O1O�i�n�c�iP@�X��Cђ|r�s��)lZ[yB��?��͟\#�,��r$t���Y�6RC�������{�-�����ɍPE�U���Ry;���kQ���`��#�w�
�zt�'1.	U%� )_�p����d>7�����ȍA���jR;ax�-?�?������'
v�z�m7L; E��B/w�P�fU���IO�S�O~f�+��_�?���a�!F�<}�h/O��=�|���i������{�"��B��gu XH �m�>˓mk\|��iC�^���OL�Y�I�h���-��h6��e���'�ڍ��"~"��C��~���)^�'m6Y2ҍ����Y�DNJ�$T�G�]�7�Xu ��À<}*����D���m�j����ă{t0�m�@��	���d����Kܴ�?)��	��a����ܩ��㋅q�'�R�'wў����v��GИagfq�t�B~pƢ=��bg�&�l�`�OJd��'U%ዦ�G}Z��Q��O�����?�i>�<�a�Vn�L�4�Yp�
����T�<����h��ir�C�����\�<!�hhX� KƑ	���a��Gq�<��٧@�f��U)E�b<�aq��E�<�eK�!�:�P��ЀP(m(�,]J�<��()l�D�!�N',���0�F�aybi_��p>Av�	A���@��_#L����_�<� l�Z1��a����'Q�����"O6�z"׆2�"�It��oz�4��"O4����1&� �Ǎzx�А "OrD��L��^̢g�_�m��ͳv�'7>0H�'C&�"�D9$�m�u-G�k�fE�
�';Ĺ��I�K2�k�$@7j��1�
�'t`��W�W5 ᫔֨�2�!
�'�>�F[`Z]h�Nת��	�'�9�؎���ˊ
����	�'��<H�g::�곆�m��*��DW�C�Q?�Z�c�,b�tre#N%$eC1�)D��9U�Gm�D�q�Y��p!�@-D��IR��d,0*FC#~��h� +D�,�����dq��GҞ�Q��&D��1s(��hj�	ΕF��:��0D� ����Z@��G��,E��	���O`a�'�)�'s�%j ��^l�zroP�a�,�	
�'7x��UU-r7�b�P�1��'�R)�A"fh��B�ʹA��d+	�'{�,��(�Yð���'��-K��b�'n5+�-
*t<��E#�����'�&�����vb]"� O0H��AS/O$�s��' le�U*���q�"�Tʨb�'ʼ`֭�	K��a�rNڎ|�\���'?VD�f�@�g��I�Ȏ�7iq�''BixR��}��)
 H(l6jp�	�'�Np�z�"�r��;ul�		�D��i��|�n��F��L��gDÜ�8�ȓ}��&�ž]�*���MȚo��P��

���H�-bq������^U�˗'�,wP� ��ٓ�<��ȓ��qG�_^�����uڨ��ȓsdTB�@��)1A��2a.	D{��樟��{�#�{T5 S��t�Fa"O ��	�R����o�j��Z�"ON�@�lY�T����a�V�@"Oh�H���
��!b�B�/4�~�P"O]At�
�#Hj� �3���b"O��"�*=lh��D�An����&�'M�])���e+����$�x�&�ŊH3ڦ��ȓ}��+����w�����҈`�
�ȓZ��|��)H���#₪V�p�ȓk�Όb��^=R�*E���P�V�$��ȓ[nP�\Z4)�%��AQ�`m:D�A�T�K��+�����Ղ�<�$@�u8���S�Ћ��l�$�$p��\�F�"D�|�R)d���B��*W��m1��=D����E7%�((�EE�w�D�>D�d1受	}rث �B�Pb��	:D�@ҁ�R'��̀c"*�+�g:�O�I�"�O�ac�L:�HU��7n��W"O0����/.$�XA�HDR� � R"O�m���J�+D���f���,kG"Om�� 'S����ek��^n�d8!"O��6�
�
^r 8f$�M_Xp�"O��r�#W{ޭA	X�r@Pg�I�S"�~���ڹo��2$�t�H���JSL�<�6I��fgZ�03&��	;n��_s�<1B��!s�"e!����'k����"O�����&,� �Zq�ٍ��8�F"O�$�BePͱ�I�p����"O��p�B�L��t�$�� r����'�ڝ0���
�>�QGKI�$ �����.���ug�1�._3�j�G!h����S�? �\22�R +6�4�1n,�a��"O�Ep��ü��Iis
�bL�"O~ ��Ë6o�.y�fFѡZ�2�"O*E3(̍6��P$��Y8�Q[�$�C(<�O�����5Ѷi!�)via3"O�[#��<!�]�s&�0# B��b"O��[ /�r˴x��Ix����4"Oʝ�diϥ9����d$�&3�`jW"O�e�feM+K��!�lA�۪�c�'$T��'#"���@@O���6�B ^<Bu�	�'�n�rGؗ%��Yzf�Q�8���'�l��h�>p�4z�.�.8l
%X�'bl���4Z]�UK�DM�"��-��'���'K�)�,�[��	�-Gl�b�'����Pe�ѱ�����,��䟂I}Q?��v�[�)�Z%�d��4�Dl���>D�Lx�[�q���a�4�6<S �'D�4����8��@{�i4'%D����"����#�ug/D�Hy��!���*'�K%lX��)-D���&��P�I�k����4��Ot��e�)�b�N���1Z�%��G2j�X���'Kl!���{� @�Z]'��'�	�ӱ�����E6&��<{�'V�Pj�'�� yЮ��*��X�'�&�{ҫF4��R�B�ţ`�<��I�2�|�{��]�o�d��Ԃ�ayR��p>9�+H	hM���0-�4�J��_�<!�#QQ:茹&��)�R�zF�W�<9�k�b~�)��-�|�,�R���P�<�j��5��ٴc��p���떃Tr�<i �Ňn�I��g/H�FH�Q��Rx�����p��KW+e0m����T}I�"D�X�e�MM�͹!I�u�V����5D�AWH�%)���S�PHd��4D��DE_5X0��E��#��ț(0D����KD�?3D�I����.���:pe-D��c��a[v(0�A$=�Ѳ@�,ړMf=D��##9p�L����+�^p��Ō�y2��fF�hEg݊KD��j���yr`n�ё��Ю@N�	�p�Q�yB,�A6��ˢB֋@��a#�ƀ�y��ԏ�N��P!R8	�x���?�y��X	]s8���L��8��*/�(�?)�h�w����tف@�r���&�$�.�H�#D�|[��
ު��`��1�A!��"D�{gBQ9rB��j�k��X�2�"D�8��"�4+K�d���5�t�j�k=D�@P%,�()�d����'AyE1D�t:�CD�&=�aӓ@���Р�<�ÏXb8��	�
D��qfR�@G�܈56D�l����i^�d��I��=�
4D�Lp�g��7*굑W���_��%*�(1D�k��9@�M{#J�LH���3d$D� ��E�u���,D�� u!b'�Oވ���O����E�
C����3 �?zꉣe"O�X0���|��Pr��G_�-;B"O�p��*S��AĒ�k�ԙ�"OHp���]�y�>l����1�P��"OZ9�%/(|1�W(��D�q���y�.��c��`:HZ�����V5�hOI����9��1 �L��"����&*���(C�	4��G����\J�%	)�B�	K���᳭�"Hah�G I�f�B�)� t�:q�Чj����@�B=�6�p�"O���#��@����F/� �����"OA��k	X�ɐ��)�2�0�'A�,k���/5��cC��:Y|�� ��&�v8���DA�CJH���� c�\yz
���.0�$�a��(� qh�K�����ȓ%�	i��kr�0�P1D�ܘ�ȓ�ҸC@KX���� 
�"�Ą�s
�`�`�G�mD��P�)���'��I�
��E��i_����4!ŚEӌ,��W�����D��M3� �"�ش��$B�܋$�W'{�)B�I�q��S���(j��ٖ�ޛj!���O��\ V�?[60�9�,I`%������.N�Q%�ʿ�Ry�4ʉ8��B���,�!��35�f�CS��DB�3p����D�8�[�KsFB�I�wZ�q�f LO$��R$T4�6B�	t���RA��W���Gϐ�5aB䉀�:���)9���	��C4�=)ӏ[�Og"�1�/4P@La���Z.��D �'i�M��%��b�	P���~��'���h6/���F�����u<�t�	�'z�(�C%P7��ᪧ�ƚpl��y	�'k% �K�����Pp�@U�L�'X��hK�V��yB �@#8"h��YN� Fx���	�I����΍�W���{䢟���B�	�Q�͓����x���K�,ƾB�ɷ�����G��h����P);˺B�	w	��R��4i� � 
���B�
��,�����bԺ&"Kl>C�ɒU��$ȃ�ςe�a`b��<v���}�$	z~R��<<6���{��?��	�&7_����-�?�4=y�����?qa���?Y���?�l� :�x��+.1���������F�5��hT�-�TI������Od� �%�1���#��3Y	�q��O%"l��Ɍ�t������T� �D	y��D��2��pӎ�'?�pw$��4��q�#�<7@jh�#�<����0>!!���:(���NE'I�"s��p�	k����g�<��n�&9�بpI��&�P%��QyR�ɖ#��6��Q�
���|�VE
�����}%���!U:3X�꓁�3ʹh��J����ȣ	����-DB4j)��b>I��e���v�� �Y���Yf�d�D���
�:PV	�m�W����w�ӖV �qCW��7/*$�$$^�l��ɶu�x��⦅!*O�O��4?OTQ�s ܆#jp�Ȃ!ԸR�)�"O΅�$�  X�
UN��J���s��	�h��7m�oS���J^	O��X���-��< �*�OD�䄃bYY����:�D�On�d����M��`���S���A�V�lP�"�a� ҃]�������.M�\A㈒58e�Q��<�t�HΦ�[g��z9 ңN�ThB�u��ԥO*i(r�A�:B�l¿A��r2��$���OJ�$�Of㟜�'@�TX�1�W�o4���fMO�6FlԆƓs8>0�c�fPYhV��K�,)��B����)�4�?��y�M�1Iö�� Y��iaS���?iÃTo��4)6�Nr�m�A�>���fn+D��	!-K�?�e����+e6�q*O�=����<*6�J�〉��"O�qI'�S�\H�*&�H!H!�Q�0"O|���.�;0���S���&�|�6�'J��M��kӥ9q���A��>�J�!�	3D�`��H� ^��i!�~43�2D� Q2�9N ����܀}>2��2D� �S�<P��;�Œ!u��,D�<�P��K^xA�C�zC��:w�+D��K�.�,b�^|��& �*v銕�)�	�"N�#<����c�h�F�<�r��@���:�"O�h���ȇd�X9����\��"O��V�G������F�K�U��"O� �$��+̊���Z�Nq�$"O႗��f#�!�5���w�~�"OnPi�Dշ|M� 1UC'D�(8���*�O�}�:.�A��
$�zT���c`��ȓ,`x����Ȱh�^!GI1I ȓ`��`wiW�n$d��mI�qɤ5��f�P�"D`���j���>_nL9�ȓxHX��å�����
�854e���;���2�Q'6�\&J�"(�\C�A%'����A��p���P;ZwcR�'��i�$�VP@ՀF,'֢�c5IO�#���%VFΤD: �V%l�8p��8?�B��w���Mw-ʱ�4������'K��q����+����
˓L�p�	!&��hS�5 f��af_"sRE�	ӟ��?Ɋ�)�2�����,�-��� �C�/;(C��/*��R��ψ]ي�H�"�p�R�@ܛF�'p�KBꮟz�$b>}��
O�CB�(����.�3&�Op0�#$�O��O�1���
�	b.���l\�6�8R�	>�H j{&]:�qJ$dR7>�K����k�x'�8bpHM|�~�Sbb���__T�+�/N�}5`�ێ�D�11}r``���'?�㝯r�d�e�@Y��ճ��<!���0>���K�:HYgE�%q�)�*]�i���TC�<�`�02��e�1a�89�����l�Ny��'��6��O����|:���d�(�L0��%?�1�G��+���D"�P#���c�� ]J�(�U�?$֐�?��4�ē^��b�)$�ͰPRN�v
c�xL��l�Ԧ��I	Z�nE�R����؟���ԟ�̓+�@F���8��pG�M6ʴ;@�/�M;�"�����yB�V��������?��]��%:�n
�NDP��d4-N���'�b��!I�$u��I����ҟ��y�����H�~�!�@�Ns��8[����I�������<���Bnz�U+��;�e��i��x ��T�^$���X���ޟ�J�k�����On�d�����	JB�@���Pʖ`AdiT2s� �	
p�����Oĵa���O@�I2T�h�s���麛G�%p0���2b���g&����c{�h�������7*��?��Vp�<��҆^������2j�0�H8�y��@��?I��3���Ox�	[��s��!��`]�y��:Cn]�#h�f��N��l��<9���Mӧ�i�f��ϟ�����T�xR��x��s��(Tb����Ц��7AO�<!��̟$���?��I�<�_�|����p���R*�4F������Ы�MKE���?�.O���O1��ɧ%N�	G�U&�j �&sxC�"kT�����Ȗ(��1�̙~#n7��Op���O����O����O��$�OR���7F�\ѓ����cC~+���BG��n��X��Ly��'��O���#������C{j�h�$�<c�&��Ey���"<�D���[�#�<��O�y¦���,b�D�����Cɻ�y�L�Ȇ��v�S�^n,Z�b_�y"G
Up��K��ձ\� Ya����y�M9%����DY��"�IL��y⃉7J|@��\�O�~�Z���y�(.3��Z�_"GWh\Q�`�ybi���
-x1�Z�@��q��yb��E�xQ�"�ɒl2�5�`+�yR�O"�HbG�W�k~
�Q���'q,��0�E�����8[��ڋa�!B�kW�d��)#s*O���R��Ki�q0�ܘf�r�c�}B��!��DK�#�w6����B�yw�Mrq�J�:*�\�Aj�' �h��FaE�c���i&̾
�N,�2	U�c ~d��Q�p*<
�l�=�u��fJ�_�8�� ��>؞4��F��=Kr���B��#FH�{{,�x���b���@*jfL�`L+/��ٗʑ9{��Q�ؔ�M�ӂZ�}p�0��PVbq�R�> ��'�Tݙ����1� �'z2]>��O� �(��B8�(%�Г��w�O��C�d�4�F��U�O����,BӲ}S�R;{��92H<��x{ܴ���'��'��D&Ă.h����)_6ֱ���X�#�'8������I7z����?��W(xl�CȎSG��!uU"ABvL���4���'����	QG&�LA�d!f%�*y�������f���'��'�����ע���?���?�_cM|�0�k�� ���%I��������3�(�
Ҭ�O �pcF��o�$�DI���$��.�.��U0�K^�p@��iI ��M�b�i& p��O'� #�|�i�e(�3�J�:�kZ��(�A.�&�?g�iE�eI��,O@7-\5v���+C�"�:���*��G{��I�ͻ�"��s���ƫ؈^�<m!���<�?i�C�Iay�\>��I~}�Z�	P�D�W�N��hS��:,X��& �����O��$�O�H���?����?Y�EP�>̬�)&�u�֍x��ʰ*����� Y�]($l�0=y�� �f�9Qfl��?#dP�0��`5��f�?ڮ��0�
�y��E%0ʓXW������.�����H�)k"yH���L�ڴ#�O&��+���i�8K��̰\J,(�"�ֆf�������?�|H<��g��wv��AѢF�d ��z��׭j{�	˟|+�4�?i/ON@p'mɦ���ͦ����ʷuhܜ��$�k��jր9�?��(�������?�O/,���ēu6����I)��:\Ht��ɳ`W�b�p����Y2�@9N�'��i4C&,Oj�"�'���'y��rQl�8xdl]Qq�ˬr�̳�'���B����� �V�uyL�
�'$� ���Ō;��H�@@�*{� ���{I�'5���5���7�'v�T>��w�ЦC��^�o��f雵m f�{�&�0�?���i�`���瘧�Y��k�䘘B�����WXnAӲ�=��A���b?Qb��V��Ҽ3S	�>y^HOd1���'Kj�O��0}{'�b�(�*��^�v��� �"O�9�"I�Hk�(�OD�S��ȣ�'�ޢ<��I�C�A(x��-J�rH�7m�O����O^	��q4��OB���OiѲ�@�S�u��]!�߼[��b�@a�)3,O@Yr��:*��(a��`��[���Й�ayR�@�3=l��*J�.���  �)kei'��  ,�Oq��'|B
�!�U�"*�LX�wv�b�'�(-���@CS ܃����%���L��C��4�OL�!'�ϲ<l�1#�u;�}���Dx�<�Ăڟ8�	�����3�ug�'�9��l��H�/�dI����>Zu��.�����ӊ�|Txy`��Y��p<iU�^ ���}��Ƃ�V'¹A ��-l�`��]l�`��1O��1���P`8�ѢԁT{��r��6sJ�)f�V�nZ_��^�q���d��.d:�Ӕ`�;FJ�z�"O\H�Q�}-`E��dC>o9�9�� ̦=�Iby"��@�'�MQ���$�R�A!�,pP��"�A!2�'�8 ��'�4��H��	`2h��`�����}����6��%���6!݀�p<�tL':�HB�)��Mf�i���%e��*ԫ�!E�P��������D��9B�w�@x��:�$iA쀏;#�4�7�9l��`�=��˰<	��sB�a��C�0��w�V�'�ў�9q��^�>:p�&�(�r�@����<��>)�n�"��}:c��v'D�;�Ȗf�<ɥ�](<P�ө��<+edYe�<`m�1Q�Hh��~%���,�d�<��4O�xBco�x@&��u@�b�<ѱƟ?��$��O 2 �QɅE�h�<�1��11��-���=t��$��z�<�g[?+�d�Pz��dᓅu�<��kП`TJpFZ#F�L�B�z�<��cP��(͖�i�R�ʵLn�<9�cS�Ra ¤��7x�i�<���X��D�&�Y�h�ݨ��\�<a�b+F(@�C&p���#�d�<鄦��M� 0@bLZI���a�<тi�#g`,h��낆&J�V.SS�<�� 7=����#��m�t�CF�R�<qp�Hc �k�J=K��ɱ�]L�<a�
F{'ڱ;ciܷ5�L���SG�<2"V�<�j�U/ϲ,	�0��LB�<a��ۦ\ƎU�%XQ�fu��EWI�<Q&�2"Ѩpe�
XP��� E�<�t�\!�:�pl����Oٗ{	!򄊤|����Cg��3�v�	6d��z!!�ȴR�h�h�^F���@>!��ËGLp�c�&
�?l2*�4o!�����{!�&1`t�b�1.i!�$^<L�m��O+�Sq(ń!�dW	l�
��FiJ5I8\X%�C�
�!�d�174��ۃ"G9$�(Y���x�!�$�0b�ē�ۏ������#:�!���H@�xp@�8lj��̇�D�!�d[�r60���A7��x��ܐ4H!�� �u�`̊��������5�!�"O"5�w�&2���Ań�)p��S"O(�A��MA\y2N!�`I��"O,XHע��i�j��v�P�#_]H&"O�UsD��;;Ԁ�Zs�#*@��"OҸ�p�M�q���G�:|3X�+a"Op��I c�������D�h�"O��h!A	1"��çE�DF�"O����� �)!�����k"OT�*Ӥ�.���)����,�p�"O�T�1��<�X����8X��"O��vH�	���k���u�Ҍ#�"O�Y3�h�h;�uR�G��%���"O`|R�튤$��i@�$�Ɣ!D"O��)q�ZB~��@I�:0�Q"O���ߙtx�9���qD@`�"OX`+(o� 0�O<<=(4k�"O&�� B�XnJr��	�)�"O���VK�$�>��ǻ�4�a�"O�tXը�>Nj���-C�K���`"O���"r���+��xjF"Ona� ʘAܨ��� �&Ϡ	�"O�=s�-\�G7�I���!k��Q�"Oh�ˡ
�U��˄-F(����"O~�Ȱ�ІU�,(�,�(�t�Q�"O�D�BZ�q6 ���G <�R���"O\���@�0orm�gk���%�"O�\P��ϝ8�AZ��e�"q�f"O�X(	W���'�g�H�9�"O�����n
J�E�3\(��"O��JcL�C���Ы}�3w"O��8CB {b$�zc`ӛE�2�:0"O��_^�@���@�N�B(�C"O9�w@����0QFؓN� A@"O��Ŧ��^=�D���"��P�6"OB՚�δ~���0�:$��T��"O���\D�'$ʬZ���y�"O��9���3Q�>����ѧ �Qr�"O����H�����#6igh!1�"O$8���$
�c�L#~�B��"O<�@����D�pS.��mC��#�"O9�C9~n�a��˼@1��"O8�Hć\ ;�@�ׯ1'�t��"O(���˻PDT(�"�-3ڴk�"Ol ���D�5�*�	s�M6�`T"OhQ(à0w��� yQ�"O,�r�K��h�"#� �	�,Z"O�d0�䘔~m�)"�o\U�i"O��Z�,ل"�9�4 5"O�E�%�ҵH���C�A�#�d�x�"O}�h�)�8�S�o[/F���2"O~M��(ŀb4�<pA�9N�&�6"O�K(�c�!I�wlMs "O^�u萡�ڝ�g�g]�,s""O�}�$vj��##%��>Q�L(2"O���BgݫvȆ���#ǲA����"O6@�L�N�{�BJ�e�4zf"O���D�*����A �PS�"Ob�+�b�&�B���&0��0�p"O&m#��ϱuU�8�f���@)��"OdժģVl��I��� ��0e��"O4�" OC�	�z�k���h�4,�"O������}&�!+��ɳ��H�3"OJ����1b�z����$��"O� �@+'�O�(|hU��7��u�!"O�a�0EӶb��R��18cXE�U"O�I����4f���e��&OL�i"OT�tcQ3{��]�w�¾�L�W"O��� G��Dكl�8��"O�sT���:�f��q������"OFI��M�4�r��a ��~0�e"O����Ȇ.�2 ��.V�Eҵ"Or@G�6E�@��kS=��	f"O�̱��V�^�k��?j� ��3"O�;����8�,���J*v����B"OŢA'�s*��)PMсʸ)8�"Ol0�b%�����l�w�v��"O�� 0=�49k��ֵIG�6�-D��#�-(6�)!��C��X¥�-D�p�G����D�GA\�DĆ!�3�,D���t"V�+R�j�D�q�j���=D�0s�	�n1�M;KX��l6D��Rf��#r-�Г��͉M�J���H7D��	 ��O�jm��l߻0X& t&+D�t�f�7�X�sa�:?H\� %+D���G�i�$�`���`j��{A"(D�T
b�Ә}�b��A�L�2���L3D�,H�nLrX��Q��>%���9t�#D�#��!�I�F�W�`��T,#D��kvhO$6��	1��|膰�E.,D��{©I�&
h���A�cD�cf�-D�k���`` ���_�VX8��l/D�8P�a��k��%Jf��-y�U�+D�$K��&*�Ȝ��32��Ӥ*D�x���U�]�D�ӡN��iHT����%D����Q3����B<��TYBM"D�P3Wg�?F.Lq��-�)C]�)�"D����E?m�l	�H[#RԮ�`�2D�<�͔xT\hzs	�$<�ȳ�1D�d��ꕌU�D���
\r�Z��*D���
B�mA��u��0�.P��#D� Q�Ԧy	�%���n��2/D�裔���HTѡşw�N-�?D�ڢ��8����2]l���k=D��"�l�� �V��@!��aɱo<D�1S
�&'NЀѣ��XR�M&D��D�K	j�̀(µ_�>Mr0K%D��EBI�S�:�H�G�%mR�QZ��"D�2���^��W�\0�����!D���Hӄ~V��+s@E�X����2D���a]���l"@g®;��@1�.D��Y�n̐\`%A@�=)��H1�?D�T��+��:�I�ˀko�}[�>D��E��9e6�"�r Pu�`�<D�laL��7|�-���/LX��hǋ8D� ���ӭm���H��X�1�d�1D�8�u
�1�F�)v(��q�x�6C1D����	+VR6�p�ES�+w��J-D���0��Q��TKDc^���r�,D�xREh��L��	r���P�b��(D�<b�IкB�H̊�E�<v�`ȡ%K$D�03G.�8ejH|3���!}�8,�Gc<D�`�f�X�ln$@�kKo+�mX�<D�8s�j_�}˼�psd<G2��/.D����%�\H�0*�v�\�"/D��#�jQ�+�&��@�N����&,D��a��ɢ-�L�H� C+�"Dc�)D��!���"l��Dߥk�����':D�� ����^d|��#�Mr�v�)�"O�t*WES�3�꡺&�2m�p( "O8љv�'/5.8:s�"jP�@J�"O�q�åH16"F8#�KH�P��"O���(�#CR����2,6Y��"O����
*U�����h �f��S�"O|̐5 B�w Jt��FW�=� 6"O(��瓴8�N��V%�*`�|k�"Oj��A<48��qEE9m�h�;$"O]A����p�%� �L  �"O���o� <��\���E���"O4�K��oDF�����65��bc"O�����5B�m���L;^Ѫ�JE"O����8�r��T�u���{d"O4�A���Pcd!��e��d{�"O� uS�VYn*���A�����"ObH鶠D�kd��&ъw}��"Obd�m�1����fM�dΕP�"Ov�!o�,K���$�{����"O:��An���b��IP섂�"OX��b+-7����%C�6�Er�"O: ���P a"��v�M��B"O:|9�F�NڰeA�F(xu2M1�"O`������������bm���"Oy��F��I�L��E�l���w"O�C&��;�����Έ2���8"OvU�򮌳l�d���A$T?��)"Or�P�FL;����F0-;��@G"O��`'��5P�C�푫[C�Pc"O!1@G�$�(�f�+|�
�2�"Ob�PV.ʼy����#l�z�"O>�9V/ֺA�.����=S�l|[�"On���������;aA�Q��"O�� Q0��`�A 95l�%"O*�[��|�����O��21|�cs"O� �D@�;D��b�ַC��	�"Odx�EE�,?�6H� C&[�.H+"OMӆ+D!R6p[ �ʧ-�Qf"O�� ��I�����[�e�&	*f�$�"Jӄ���F�uI�k�D��'�(��Q�����<8$C�o'f���'L��Gj�C1�tK�H8l���'\��p���M.�	D�Cld��'LX�)4����@�P�Q	�'i��en̵9c�e��Y�&�K�'6�x�s/O��<�b��7(�)�'��	#`�K�����
[  I�(�'O0H��Hѝ9蠝;!FңPV\a�
�'�
� ��4L�4H���@+����'f�|j!\�X��ڮ~����'�ּ��GƆ,5j���(�5{Pʬ2�'�L����ۢ�|1�1��s�d��'�2�b�FU'TqB�!����o4���'��I���O������d~f�0	�'�>H�e�!��X0��&��TA�'4�\�ī�	"N@y�"�
����'��L��)Wvr��ɓ�p�� ��'F�ۄc0T�h�!`��g;��y	�'%B��6� � �ج<Rh��'|&Y��H݌C] �Ȳ��3c>�'��p*W�XOQ@�8��Q�0đ��'�����i�@���c�8�B��'l���b-�:AV8�Po�8�����'�t�tϱ[Ed�(�X� ��t��'��Hr'���y�Xچ�0p#��J��� 8��`a�Ѥ���ʝz�-Z�"O�h�ŝ*�rhe(ɕ5>�Ic"Ob}; ���O�f]p��[�:�8���"O�)����R`�r���F��q�&"O�X�L,∔�pk]&��P�"Ox��kŦ>���� �(&�fQ"O` ���Gp�.�+@��%�Ȭ*�"O�+%)�2J@��VA�N���"O�2qI��B�5(Rw9�,0�"O�"���<Q^�kw�2$���"O��"v��=?�AF�"V��"OnI���]�{TP4K����"�9��"O�K`�=(䖡kW�ْZh�t"OP�t��#-Hp)�|�qyC"O�,"We�:J��QV'��j�҂"O.���`�`Nh�/њ#�<�d"O��+r�O;�6���+B ��"O���4�݂{+2��s�ڐVg
|�"O>H�82<�t#�;�l�"O������9k�e�w��^Mm9�"O \h�C��Gl����ӿUp5�s"O��ԧ�� :.i����.'�"Q��"O|L 5�H:�E�ƍڧ�bh;6"O�m�p%��8^츙�+T�{^�C�"O�-��I�\.��τ .jY*P"O�0Pg�7r����n{�#R"O���7�� �:���c,�7"O�\P�G�i����p�ŮYa
y�`"O
�( ��
XN�*�Hܤ#�" a�"O���v��\L���,?����d"O4��5 �u���f���1�z���"OvU�Q		|m��E��+g"O����)H����DM ���!"O�� VJG�oڬ0!A�[�jpD��"O�`�p�@�]�Y-ye��cC��y��a�ڈ�4�҄hOz��&�yr�8e����-]����{����y�L$7K��B�^�l0Q��� ��y�E5v���PS#����s��yB"�qI���GU�{�1j�D
��yrX�g��$[1��+��x'�y�.��V6mY���Bi˝bid-��'��Y�T�:�y��l�����;�'��=H#FX�e�b�s�O<
�~<��'��[�L�yL��Rƾ7���'�x�H�߲j�b8�F�g���#�'(��wdYVz]ఌ �Q
B���'�fm��c�(_��Y��C�,I��'?�\�G�ԛd��  W愼x��;�'0��Q�]�iX����(k�e@
�'Zn��P"��!_$Ջ��K(h�a��'@ʅ)C���N�3��IXR����'<����C�,L$D�+N�J&�i�
�'����,�(�@�����E˔���'~����΁9o��I��D��X	�'u��BB��~_")	�BP	K`b���'$^ RuB�(\���i��C�F��	�'����g�+"ߊ��q�T��m�	�'��(b֢ˉ/=�82)�+F�f�'�j� @ͼ:)���w�H�'Q|-���[[jdH���E��|��'ӄ���&�����B��|�����'|����G�:���/X�u��'���x��π�U�F�`H������ �Qs��v2��b!ʎ�͌m�e"ON����lЦU
!�W<O(�P9"OD��Ǒ� 6Ԩ���'P,Q�'Br$�AZ�	+��<�!�'�\Ш�JɵMؖH�#���E|H���'~�`��t 4\j�M}kz�(�'��X�q'�.��x�ąP0KgP̉�'6́4�VUxL�gc��J4�Q�
�'��Ə�C�����AH9L]��
�'�<�e�T%D�jXZS�D3A�|y��'�FE��� E���qR�)��
	�'�0�r�� -��&�A,ʼ�	�'��+�kF�Eh��S��<"�'�Q��
�Bfv���Cu���K>���0=I���ߘ�d�	,�^�J�h
p��$�$*�b��d�ߠ=f�ys�ŉg�4 �,�JH<����D�:���V1'|�rg��L�'��/��N9*p�Q�	M7l�襓�CQ4�x�-nP!�dO�p���sg�$%��Se��;q����<��-���?7*l�S��M{����,ł��!��7Z�EZ��V�<q�j����9FɷN���c]3g*�'
�#Ԑ}�@��(q��4�g�'e:��
��'W(���F�H�ʥ���jDS&�r�N�KR"I�t_z�0�!��m�riL�d���J��'��F�H�Q (�y�[�$pʌ���xa��j�
� E�ޣ]
�OH(MQ�G�e��}:@ I�L-Q�'��Y0���D|�3F��\+�X�E#j�+�Hԧ����)ؕ�h���()�Q��0x��	�鉶�!�dȓu������J% ��4x�\n��=[�.<	o�U T�Y�w/ȴ�"�Oh��:�눨��Mh���&�9�tD0lO�P��h�g�	8q��1)K��@��:^�^����>'�,��L)t^����I�Y�)��"��`��t:6+^c �b�̈S�(j�
e[���,
�L`��h��+�0���g߉8�Q #�$+-�B��<2������
�f����ùH��!G��,���h�fϽqp8�9�t�OȖ�	������Q�K=�"u� C�C�I�fPd���F^`�X#a�\-�Diڴl�v�`��,_�$�ᖣ�v�ɒ5��Y��Ў1�$�c��E�|��d��$��õ ��e�*xI��݀TH��`�e<p���
L�$��J�,H���bG	�	Jb�Ac�ț
�ܠ��"�ɣ[PP:�"�24���
���w��O�.�d�2j�	r+�=0�
�'����@�E"iX%F6�+�OH,E@�
qb�����Ha��~RƲ��]�ㄗT�bT��Lح�yBD�u_
��Ӌ�&e�9(�0���J8�c�T�8�����'�Ę�3$�����- $H�q�R��9� ��%�܌���S�[U�Sh:�xZ6��8QaB/*�����;&h1;�&PȈO��C�h��v���p#�	�¼\��N�owɫ�\�?�!�N�WOt�Qs��;r�4wG�a�L;u�$/Y1w�)�'��9�)Z�- �4��-˒B�k�'(�q�0�n�`q���!�����O�(��*���v���9��1��ڎH�����)j���D�u�rq1��\$�TD ���p�@�Z�<ѵ*����:"���B�� �h�ȓ�Dd�Ti�n�t��B�Yz�<Ō jTJ`�cbY�}�����m�<1�A�#�����D�j��lħg�<�R��1c��ci
S5x�Ť�N�<A�M�
�4x1gʖ�
!�|X7.�f�<1���9:� ��˖V1"�z�J�{�<A(�<��(��chͺ��y�<��!%��K���!]պ�r��n�<1��5h��IB�M%I[��1 �	i�<)��D�F�h�ᦄ;f��p����c�<!G���(�yySd��%@YI!��}�<� b-EN�[uGF*
�(�҅�Jr�<� �L�
xE���AL\��"O�L��AS);��I��^�'& !8f"OdUELS�0�ġE�ܻ4
� U"O�	�g�`�!��iU2��XK�"O�� /�:�(FR�;w��g"O
�r%by-&�GB*.]�y��"O���'h��m]��jW�X�CBj���"O��f�5�r�`q$H�^���K�"O*q ��6����%�i�gjO�<ѐ \I�m3&�J*�<RפN�<	�d�x�"$��ĝ_����Ī�L�<�di�5A�p��g��G�PA��V~�<�#���4��%	�p3}��l�w�<!�YZ�"�	b!@?7�� �$�u�<G��TF~�x0,�LW�ň�{�<A�ܭ>�H�9@��jF���,O�<�F+� [���z��I2�T�H�#t�<1��N�*�:�@0E]*���A�p�<	AP@����J
�!A�Sg�<	�A	�1�R�q���/�H�E �d�<i ��\��0�� $��B�	u�<�%bɬ��<	S��|d�ѡ\O�<�7�4\]��cF�%�99g��A�<	��� 0Y��.�ypP`k�.�\�<A�ܫx���u�EJ�������q�<��#Z�!����2i�9>"��j��J�<A�'
#�`]PU�2H����,�`�<Q"o��9v!�f��:�,���^|�<�Ī��v��GaH.x�8yH�%Zv�<�aJ�);~�Ę���L���D�}�<ypn�(ق#���yt��fFZe�<Qu"P 4KQ��J�2���堖Z�<Iϋ�V��}QQ��.Um&��!�X�<����襑�Ń*% �t)�W�<�&"ܸ/�})'L��e��Z�*�x�<I�̊!"��H�ښd�~��Ҋ�z�<���(r�D���LzƖ�1�Oz�<�4��0�Pp�*e�p���]�<!֌��j>��nϠp&ؤ G�X�<ᒊΒv��4{��=5�����ȋn�<iI֧T5f��gL7o9N��W��t�<���B# M�	Ƭԫ\��Q��'
h�<0���t��iv��o�@�1�k�`ܓ`�n�7b�y,��5�G�{Ͱ}&��Î��l����T�8�7D��;��V�.�N}⃡ȜsV �#)D�a�L� b��zB��"�z+'D�|q�$�!"N�� �?�����?D��X�AC�b�&�r���%���0�?D�ȩ5�ĴdI��y���h�z�J�(;D��Y��w��I�A^�76�]h�<��O�k �2T��*|۲z�<��b�"Ҏ��'!��zk �Zr)w�<Y��R�  M��g�_�d�0�g�<'��XnFP�� M2i����Y�<��G���H2�F��P��U�J{�<! �ȋT�����G����ٕ�z�<��J4"+��!�iD#>},��5ĕx�<y5̗�a�|)��i�)iQ�`QR�q�<��/�,��f�d�h�$MWG�<a��J;a*d`dZ69t�Q�iC�<��/�G3��N[/`R���g]h�<�d�_52>��gc�|�  Z�<�����vf��"Q
ڑ{gp@I�N�a�<�2��3�x�-��Ȱ�G�V�<� � :0�S�r_�E��x���"O���	M=	l��`'���s	���d"OnB���.f  Em��,�
,�"O(XSMC7%5 �`!��$� (�A"O���E���^0�hwD;/����"O~�(�[<!&��$L[.)s��a"O�#F�B�AQ�<҇d�fϊ�w"O<�q�$@�C��-����[4��$"O�]�&��7�@L���;.��"O4�G�°k*)�K�q�ձ4"O��:Ǯ �2lq-�A%���f"OB-zq��<�$��)L2f`��"O�M�VH��e�3��4�G�.g!�DF�^W�E�DD�3!1�P�7�@�J�!�Dե	��3����x#'�9D�!�I	)D�D#�'P�O��˴*E�!�ܲ\f��3j��.j�T1u�B�.E!�$�&EBI���Wq���.R2�!�[�c	�\�蛦N�J#�4)�!�Y�e�J𫲨
!i4��爌\�!�d�T����A�|�kp��N�!�D˳"<hXgE�����Ғ58!�$حg�T�phG�>H����!��Q>���Hgg�{��h��ۉx !���`� ۨ+��\��kG��!�D�r�h��!�j��i��48^!�D:��!T�Ú�`�3 N!�d�W7���w�j�Yk�!�(�!�$�Y��� ��{J*I�V�5#u!��zI�LâoH��]�4��%"�!���z�� ��-�%��"�!�$ZJ*�*�Uu��]R�#P��!�$^���Q5+�f����7B!�$ً<�b);��]L[r0�''�,-!�dߝ?�p:��6ܤ-#Fa%!�d�s�¡g������3�f��j!�d�����]�9��$���!�D]\���3q���)x.�'d܀#_!�dP41���jE<(Eta0�u{!򄋱�E�� 97��p��6Lk!�P5@4j$x!�:F>���U�}}!�DMb���@�;G6�ݹC�ңU�!���SP(lA4�^";�,�5/�!��K��M�4�k��a�H���!��>V��cӫ:YB M��Iæn�!�$+�Չ��W9)Ԫ9���Kw�!�$R�:��DjE��p`4u)�g�o!�䚹,b�A�
+Ly(� �g�\!��D'���Ke�V3f�D�qdˉO!�Č�r�����j�[y3�����!���NP��El�&NV�2� ��r9!�$�(*ʬ�2�־B��J��V-l,!�d�
P�BU��c�\KJ�S���>ft!�$�9f؋��?f,����� �`r!�AA��1X%�]�^2}w�R�s`!�Ԣz2����F�d!�E,ٳ R!�$��%���A'�Z�\���Z0�ʁ�!���(�2��-p�쫲��+iz!�L:%K�uI�F�z	�M"0(T��!�D�T�&�+�BG�w�j�+��#[�!�] X�6�HEǙp�A�A�O�!�$�&(0u�F�.=������&=�!�;N~6@��aV�X,��oQ�o�!�d�u���	��&_I���� ڡ"�!�� �x(P͐%beyC�N,F��U"O���1a��S�@a˦!4x-S"O�T��\��8"��q1��"O�Xȥˆ�hШ|B ��1x�$)�"Om@�E���!`L��0��Q"O@��NC�dP���)�X`�A"Oh�B��a�F���G����B;D��
�eC* ��B�Fr�H�`�p�<�c�
?K�D� s@U�B�Nextl�j�<�R�Q;D���B.Z���E�j�<��H�pFQ��F��\<��DI@�<�s×�TJy`�"Ƙ6ǆYa�i�x�<i��!p^-�0�K{-��Z�-�H�<���	2����Q�W���A�<a�]� V�ĉ��ҎI�d�)��~�<�Î�?�����E�m���a�|�<i@�s~ ��Nԉ`��mb��`�<W.�B8d�q�:f9	
�v�<�Ĉ�f�R�	��V�(�S(k�<a̔*���8���9H	�,�Lm�<�WO�@߀���B�X6�D��G�T�<1�)@�n����G��I+�<���
E�<�F�8L�B�@�G2w`�⋟}�<A���:�z�ׁD��4��,
z�<I�b�ر��&Օ*t�ɀ%��t�<1�U�sɆ�HB��h�}�U�q�<)��(&��$�Րs�xH��l�<�1*8E�����Q
ؐXsOQd�<���*%��ҝY�n�3��[�<���$�B9�Lʨ]ȱAW�<��bD�@(��[W���b�g�<�R�'F�Z�#�`�bQk��h�<�f�ͮ{y ��r���aAN��6�He(<��4:����& �Z�pI��D�-<��ȓO�m+c��;��@v/� G��d��=Y��C!N�Wp�\0#�B( �ȓ&��4ۃ+��6�D50� 2�zh�ȓ@�F�f��L��a��R�L��W��uˣo�B���RlE 6���ȓ~�ܘ�%
��#����̣��$�ʓyz(�G#��A׺8���-["�B�	?	3b}p���MNڸ��		�H��B�I�-�F�)���.\7 �x�+H�kS�C�I)#!���\�@ �i�Z�V�C�ɠX��˷��P��%�0O�8�C��*k5�!�(L�I-�y�2�Ռ/pC�	
i�t�ԎǊ|���� ��=>�B�	���m�ײ��`��(�I��	�'�p�S�ӹ,�j%��&C�<�+�'��l���m�����:lk$<�'���Hb�%>HM �$�{����'R��{�eF��^�B���E�Z�S�'�|��rM���6�`C�?m�\h�'�z�h���*I�$��'']��td��'r�c��V)�%crDCr:f�H
�'ێ�B,�"��"b Sl���	�'�8s �s�,BJI�jo�{	�'���Do��,E�l��C�<ѥ��"y`�I&7� ���}�<��b�!��U��cH�L���L�a�<Q�n��qPc��Un����[F�<��䟽0�҄9`�ŗKI����X�<��d��z\�gΑ��4�0h�]�<�w�W$��PlZ�'t܈I�g�W�<� ڰ���&:����<@��k�"O�'�aD�I;�%�	��Y�"O�K��Y�N.h�����2X�"O���1�_' ���$�ל���"O�)��kT41q�ÐwB4�p"O�4��OP WX}�bi+b�2�"O�8�W#?"���/@<A$݀�"OV�q��Put�� 3o���f"O`�S�G�U"LБ�-x�u$"OЭ�B�Ħ ﶑�VG�r��h�"O���fkef�čQ���r"O8(���)��aQ�M
&_��I�G"O`-�p'�8Br�Uj�
�lW8=��"Ou����[�1�tO�-
�h0"O�{@KA��ҍ@ 00"O� �Ì��s�쑕���z�b�"O�eiTM�	�>L�l�#'��$"O�� ��Z���C��'�"�"O>L9�eâ1y���gۙ�\��"O�ݑj��M��J7&X(A�v���"O��0؄Eդ!�b�$��ѥ"OX��r�� c�x���'ǽ�&�� "O�X�����H�d�AQ��<Lm�]��"O�СP��%X��!�R"$W�a�"O��*�чc��p8A%hL\�7"O	0� A�bmR���Ĕ/k.�|�'"O^��@ _�E�������9�4Y�"O� @�]f���iFb]����"O��*7/��D,��7��7��)�"OAZ�E1;eTH!#i�`�^]��"O	� h�I/�H��HM�@�L�yq"ObУ���xV�i����:�r0)q"Obl�U)�X|D�$�D%���Pc"O�u#��%9�Mɓ�O�/]$h��"O��r�����@�g�?�\�T"O�g�I�;���[eMU�D��LKa"O8�Ƀ扚�<�2��4:m�X"O�)�g {j��Pr&�\���ذ"O��I���օx&�7?�(�8p"Ol�: �	%�&����)ce��P"O���U�ة2��{aBxd"Ob�!��0�4B�-�qc���"O �R� R�g�
�����~OҜ�s"O<��� +��I��[�$h�!��"OL\��A[�e��L;���&1º	��"O�-��
�	x���#�	�,�"O�(
p��(i�8�!X&=� x2�"O��@B�*&\��ʵ�r��2�"Of=�3D۹/T�p��m��mA�"OvI�^�i�@+,X�\���"O���p�Ih��P���;9��L��"OJ�8��1}:ՙ�`����m�"O��!����l�q!����@}�e"O�RHI9�@�&��ꩀ"O��GX�S0𴃑�O�eN��!&"O�a3o�vy6���ЈR<�8�"O��	t�V26l��a3,������"O�U2���R����SM�-uz�:r"O�[͎"H��h�sF"k��a"O�6i�~������a����"O}iQ�a:p��GA�Aef@�"O>��r��^pp��%Y�	K�U[&"Oy�~<��E  ¥:B"O�Չ���6���r��q���g"O� ����_'� eP�HT, �ݐ�"OA`J�H�( ��בy�z��s"O�ᨓoUuq��@	L����f"O��PR�[�X�`�H"i�,���"O�m�sG�z�Ű�@�"�0�˅"O �`GL�$8��CZ=6����"O¥�7��L���	�(R�r�؅"O�Q�6#��g;�$I ���T5���"O�� �K$9`@P;{=d�"f"O�|! E:
.($�手&}���"O.]H�퍍.�"�CQ�.���U"Oqs۵q^��@ [�~�qp"OV<�fM9"W��׮ے��Q��"Oh����&��C$�2/&��%"O*X"6KÃQ>�ِ$�(r���"O.}:@C_�={P�$Şm��@�"Ot���!�#��@qcCA/\݄�3�"O����];.ٹ�,
�6�
�۲"O�p���B�.B�5�ܼr���"O�yr$��	���΀k�j!*�"O�ԂvFK0�����l��<q@"O#gI��-��̐P� �rղ�"O�t��l�+Qʚ<q�͐�~��K0"O�1���	a���hV/��:m@���"O�i:D��$�V�(�oY`�j�Rs"O�¦L�~6PC�'4�|<��"O��:6�ڊцX4��&13��P�"O���A�I� ����|��c�"ODE��	�/A��[ 牟+�����"O,�9(�Fm:���J��8S�"O����}�`�^0~&1YS"Op�p�\�����t$W�͓�"O�,KA ҭO���b$�Ѓu�G"O�`2���t)��˹1
r��b"O�̘���N�8�{ �_�<����3"O�P�@�H�,(0
�/2�v���"O����L�1���bp��#m` ib"O�D+ ��2sF\��!�٤@S:�hd"O��k���R��9Z�GЉu��q�"O,�hWQ7c*٩a�K��!�"O��36N9!�����׽]��[�"OR@	օA4�PsƇ�
yڸ)j"O�I2�ˎ!j �87揎\�Ή��"O��#ϕ
�@k�D��&��Y`"O<�x��U�lء�#�m����"O,�#3��O `���/}����"O���kT1p031!W 0n�U��"O�x�Ae��B��W�Y3]�d�$"O��sE��7ozU��咮O邴:�"OE�4kN'rݾ	(δg�lx�"Oՠ���7�R��S��S�4}��"O��r� ')X؈v'%�Pl�&"O�A8dl��Cwh]�0�ȶU�^a"ON�k���[��͈�yVɑg"O��!�ώ*�00�ڮW<���"O���@
�i�X�{�*ҧX~Ic"O��[��l�au�U�	]攁#"O���e���U~m2�IC�wE��b"O�˖�F�
f��"2�̢V"O���wc��-y��Dl��E "O����g�d`�%]�,��PJ%"ON9R�`��C�.�q�<N���R"Ot3ӌ�N�8B���!f���"Oҝ8 I6+�Ę$�H	Y�bg"O� D�v)�.LhA���L�TR~��"O�:�KT�U�|���(1:Ѕ�F"OЄ��Ο	�ҽ�uH՞�"O����*Fj%h-�ӤW_�D��"Oʗ*V�%��␰&��+� C��y�X0J)��(�-�(͘����y�j��6��Rl�4%�t�ՍY=�y�\�tU5.w����P	�yb����6�*C�ٻS��)���"�yb$��R���L�(H@�r�^,�y���}��pTl5������[;�y�$�/���1";2HL��bi���y"�Ԟ`���Ɠ6+r�IJ5�y���DX�쐖��5EHH<J�$��y��=���sJ%h��Rm���y¯�0Vk6�@��p<�)	2���y�	�*#h4#d�ݳfnP�2F���yB�M�!���7�Pt��c��	��y�''^$�8ql��n� �ꗨ\�yb��^>1E*�l$�[����yBK_#\P�!�_�Np�N#�yҤݳ%,����B�ЀY��dY��yb� �C��p�0*ڐJ��Q0g���y�͓�L=
=��L�^q	���;�y��		������F�wJ����!�y�^�'u��� ��!E�ԍ��C�4�y�
�(b<��Q��7�4U�[��y��K�J�,�����4cֵON��y�)��}*tcF1����G�y����4rܽ�����\{t�9�y��_$�BГb݄f��q	$薘�y#
�ꀌ�Q��Z��[���;��<��7�N����-}���;�(�>kY!�$G_����kP�'��݉4B_6C��C6���?/��0��c��,�7ツ|��B䉊qj�l+aH��qQ���F�O�,��b����ha:v
�m�
 v%ܱD��]�ēZ�$�3��	�1�e��3=��Yp@"O�� ���"'���X�� +��'�j�<!pkI)m���p�^�HKZ8R��U�<q!�ݰuO8���.q��� �{�<Q�b�����8 	�.�����Vv�<�� m�L�3��/���r�/h�<���41���� ���(R*xJ�" P�<Y��ٔM{�	�`"S�<�(z�
s�<�w�[4Sq�t@�� (u�	Vd�p�<IsDS�&4<��MM#	p��˳ �k�<�!B��R�ťX��bo�B�<)�;-����a�n,XI��(�{�<a�ͯz#���c�6�J�`� ]u�<1wC7[��}�� \$JS�dꖎ�U�<�U� �Pj�y���F��R�<��	�2 W�X��A�8�Pt+���D�<���K�s���2AF��Eߌ|c#@��<)�>4dիG�S�$AȽ:��}�<QT-װwV�����Q�1LH
�%z�<���O�fz�U���<c�!B1�@�<��m .NU�1)w���;�J��2,WC�<9FoV�r���'I�r��`#wd�{�<1UmؗF�����N
�x�`[p`x�<I���"E�QX����n���jr�<���ߟ|ƪ��L�6|�9H�Rp�<���@$bRp�D/�Z諧o�n�<yƍ�d6�Mq�!Ɩe�Lu3fdY`�<� ��2�.�7n���`�ˍWm6�[F"O���4�L�S�Kc��d���V"O*�U��&(�q#�
H�h��"Od g�'��ak��h�ļ�&"O`;�.��\/��C���]�pI�"O4�P��$j7��QAϡ	��t�u"OTY8ň��+��*t�E37wx�0F"Ob���
�N�����χ6nԱ �"O���f@~�1�J�sT�Y$"O�	q�f�:�|3���%�H)�"O�\�V�ۓg�|��$�@�? ���Q"O6�G�
2hۇ�I�Q�E�w"O����Ȍ''t�q���8݊���"Ot���OI,F\L���nE=��UJ�"O��:D�R�bZ�%@d :Q���{"O l��E�r 6%�!n["Y�`T�!"OFy��*L
j�bi�@^�$
X̺B"OxtRP�A+�,i�����.����"O�E�bу�z�d`Z�"��q�q"O���Z�d�H�.�$��q B*O �+��7-`��U�R]�D@�'�
]{�dI�"&~vE
[���:�'��A�$ �>�QA�D�Q8N�S�'�T��Lӟjt���;Ҍ}��'n��c�O�>�8���W�4�>
�'�V��c�
&��,�aS�2�%i�'�B�ۢeR{��sQjʖ"����'2F��P6\+g�6
$j��e"D� *�B #�x��!�N�P.L(�B.D�k�)".�8Q��9�&X��� D��y��4��(�&�y��أ.�g�<��N���R��fKРs$b�<���T5 XDz��tE#kXd�<� L
\y��aD�WR���!l�u�<����=`�i�ȁ�k����$͋y�<��$_�+����ɇB0d���#�j�<�S�F8T�d���I���h�T��N�<YG!��u��@	�-����G�<�Q*+l�b� q�8�a���@�<��l#r�L��VR�,ʒ�
�<�!k�j�D���[�4rm�}�<��I����i���v��X�W@b�<!���eTL�J��Ā6�`L�ł�_�<��>��{-�8e����R'X^�<acH�W8��B�U2:�5�BG(T�@���c�
�p��דO4�DSP�0D��cC@52�B�al�(٠P�3D�����|���B��h�EM%D��;q$'16Ȓ0hEib�l(�!D��Qj��#bސ{1����1E�$D�V�;V����gJx�`Q�c!�<�O ��["VHq��4��O� ����\:~�@���E�4T�m*�{2�'��5�%���:!�WL�'E�$ ���|�'�V::�T�S�D2M�,�� �f�'�Q2ViՆQBQ�U���"�� sӟ\���j�.#�T�7lW&q=$F�ɰB�����צ-��4�?q��������m��KP�\<�0���d�'��)��hqĭG�c��_��`� ��o�a}2�i
�7�pӮ�c���>��rnP�7�R����O��92�\�j���$�<�'t]�Ɲx��И�Q��� K+�Ձ��f����fh���؇BJ�qiŋ���O���;j��O;E��ea(\��J�o�*M�&i�N�XDL"�Z�B��$������C�{���iqmț)xR#�ii ]C���?D�i�R�?5$?7팖86:�"�m��!�M�{���O����~�ր�"8*m���z[Q�0�4p6�f�|�O��"G�Rx���\=28���^08�'���v�<��DQ2N���bJ*ES���"`]�b2���'�C6x�{w�w�{uD�?���)� .8uAC�Jǈ��rg��T��8C₪AT� eʆ ����	F��p�'�D�ɖ�Z0C@~��� �I��Щ�)�O�;$�O��$����Y���I��Dl�!R�,غ�i2����Λj�NJ�'���!��>]�Q�ÎU�9fz������1��4���������}��!�A���I9��L��"�@QiSf¥t��d�OBY`��>0T�ɲ����cpm���2!�� 3�T�R��E�[�m���b���΃W��0�Յ��hib�Ivd˪z�:�1��� ��䣕�VGj(MNC�'f� ���J�6�
�F�2.z`���A�g���%�[�XT�f�'!�	�4�'4�� ��F	g�ڠQf�
�J��1�"O1�J׼9�����d�Iq��Od1n���M�.OV�K7l���IU�7pQX��D��$m�ɲ��U�;�������d�~e�1�<
F��jS�؄{�x(9�Ȝz@H�)�}S�L� �>�(V鉡C��YG/�Z9IW��Xv���O����!K�H}���[^,؉�D��O���r��mZ���Oh�Y0AS�T��PעF����f�O|�b>��IZ}��ͨP�LHi�U�(��h��@F7�p>�2�i�7�m�T	7�T�8��:��X�K��M˒FG�z����'@b�'��D�%L�"�'ԛ��v�*�c�5*�H����~��e�'b~!��W��yB�'���[�,Oy�'�%oj�mp&�I1`�>�ң�iY$��냡�<�8NW�G	��1�&K�0X��k1��:�J�-�,��q,W3%�~�*e�iH�ݑ��?��i���sӾyppAQ��#�-`G�t��$�O��(�	f�5��9s�G&Z�$\�@�)0�yFybOz��o�ɟش�?1�'�u����ݎty2I�-^�(*W1EY�Of��$�?j 8  �   f   Ĵ���	��Z�Zv���/ʜ�cd�<������qe�H�4͒6R64<�b����%�0��-�VEC�A3�0�qC�MӐ�iU��q�ؔ'��	㦱�1��9�bY�Qc.��5�L�}�F���K�L�
Tg0�o��'d��q��˕L"�F&K&�ʘC� 9 ��d�6�����U�B'�����	R}vp��3���=V|U����b�T�Q̖�x��dW(��M�#�d��TĢ�OV��'�N��4"�6Ʉ�v$Z9�:]9��َ=����"�+;�`���]?��	;\̞l�7C�?eNѹK�mMV�y�T��g���?!Q�(�赁GJ�O���	�@���Dj��}�Tʓ= �Įj�i���65��)�B�$M*m�F?�I	j��)S�I�r�H��j�H���9P�T�O��������dQ����˰H~��[7,6'��#<��-�	K_y�fm�@�� #��Z#J6ԡ�OҀ��X�/x�pp�_4�zh#&�#�����$W��Op�2�Op���X3T�����d������_��ȣ�ɕ��O���d�;M�n��w*ۍ5�:�!Α�O:8*���[��?i�g<1����Y������[̓m�d#<��-"�$�,F6�E	[>G���	��hi��U(�OJ��J<Y��O^PJ����}���QN	�H� H��'7V�'���Z�I]?��O����t"RX�$yӶ��?0a��s�{"��g�'$$�O��5����4oK�2�N��]� � ��d���9�.�,������8��a���5D�� H   ��ł%}r���&"O~jai�3�HI��٤uU�i�1"O>!Ȓ ]#0s�h���2Sp �g"O�|@�� \lH1�t$�e��F"O�P��(׮cYZ���,��_��"O>�Ke���@�٥�	2eH8��T"O���A�xz��q��D�G���"O��3��Q/6��!sƭ��=���v"O���ťl`�t����A��Y�@"O�p�Hϋ%"���vH��"O�$o�ٶ��¤K�}� ��"O إ!G��Eq�C� ��h�"O��*p틎+�ԱH׃	�F�,�b"O�ER�n�R�S�?Zӄa�"O�s���>殡#Ǉ���Mjr"Oԥ�$��)jƃU==x�"O�Ő�E5j�R͓�䗜/�ȸd"O�hA�bv��UP   #
  �  @  �  b&  �.  �4  ;  wA  �G  �M  VT  �Z  �`  "g  cm  �s  �y  ـ   `� u�	����Zv)C�'ll\�0"Ez+�D:�Dlӆ�>O��JB�'� �a�0�R���%S�A��$j�醊~�Lhj�E��]��$K�W����aݩrGH	�?M2��?�Rc��Q��M��j�0KƮq�d�5@�ԉ��7@�D�՞U�R��7�	��uGiГa����'�������o��+⭒�Z-8�5�̦C�"Qi���O��Q"m�&�2��S�Mզ庠+Dȟ�����������P��	+/��jC�X
����
���'��O���Ҧ�����OL��Mn�4���(5�pȡ��)DL��%���O�1��@|���'�D���Ђ��M.I���S��7<_n��	-ғȈO�6M�&���r�G�v�X�7I�_��m�'6���H�5�w�0* ��\<�UN�tb�[���ϟP��ٟ�I��0�����	\��3���"�Y2_.@qb���H����'M�7���Yشx����'��$'H6휓:8��d�'�$H��`D�a�(�>�`B䉁Q�>}r�T�dP���`�����c���Ϛ�0��#*���o�,�M�r�i����Ofܭ�'ID瞅�B@L5�l�F��5  ��:��y�X9�&��*�HB +.g���b��O�⟠jr��?=��T`N��$�`@
ڟ���D��xX�j�v��$�g�@��p"7�*���?�����O����wO��L����A�1��!�,O�=E����2&�pX��M�m(���SE�7A�r���������M�ʟ��+X�Oɼ����¦�L}�0�'��şx���|��E])E$�9�O��$��}u@ x'���%� �r͗�m���d�#iU����XR�\�b���OdH�6Nߡ?":����5��]R��'�
����?9�_�4�� ̬W�2��0L�z�y ��O��D�O��b>1̓ �e3䧁5���8�^�`��ć���M�� �5$|t�
2��):\��C���t����=/(�⟠�Ӓ44�!��"�6Tȹ��@��d�d}�ȓo��<TaV�(��e�[=^o4%�ȓ�C3�dc,�R`�պ+E�u��0Z���u�ʅ=@�@���}��@�ȓY�^�&A�.�@ b䡄n���ȓS����VT#�L0�C��E�	1>�"<E�tj�o��4a$�:�1�	R�8�!�$�ʲ���w$��+'�)-���ȓ*qh�3��͎��UZU��$KђI�ȓ`V�MA���@2�e�s*D(�������	XbN��>��PS&��썅Ɠg&�CS�¯Y�(QA���u�� ��R6��$�O���<�-��瓯|��Y�D�N�^�B�╣�A1�1���ɬp�.4��	=G���KC��J�eBA*�r|�Х��.]�x��C�='�֙b�G��m�hxG{�mE5?<���z�V1ܴxun\��d�Ӧ푉�$�<��O����*9���eV�<ծ�17�'�!��JF�$uy0�O�"TF��фF�!8�Gs���ͦ��ٴ��	ǃcJ��l��̓%��uS�K7~�н�0i�'JȜ��	sy"�'��1�f��
Q"U؜�����Pl��9kdڠ��ISz�1��1ax��Ț'F8��E��F��sd,"�TyQ@h*(���;���#�lٍ3�ʽEy�ܛ�?饷ij7��O��c�uB�Tۣ��V��仆��<	����(��uY���[�@<;T,�LTE�	@�'��7͌)N�y�QG˩L�|�$��3��n�Y�'-U�2�]z��JG��;h=ɘW/Y�R����6�y� ��;�����t�^��C�:�yB*A�E�Go�s.�=�ҨF'�yRl�q���hfˍdw��R��yR�A:�M�r-�\W����#�yR��6^�5!���5U6���3�(y����|��T���'��'A�	/%B�L`t��W���ڀ+g�f�[ ����(%� �ѥ�Jt��ɍ2�"q"��X�J�@�mմϨ]�p�^� ���	ؗ�F5�J6��M���کO��!�x$�dH7$�I�"!16�'��yd$Q��R��p�I՟0��G�@1�a����
X���bVQx�`���J- �2�{%&��$M��@����Jߦ�ڴ���|B�'��D	
)q���DHk�p0q��(�*q0����u�IΟ@�	ay��D�9���g
�U�Z��t�ј->������I��qF*Hz0az�ė<<��\+�K�-�l�ؓ��,)A�	Ȗj�!�L{����ɺF�_��"=9���Yvt�f�+�0���#al�	��M�-O*�$�O����O�D&
CCPS�L�f+By  G�g�<�Қ8�. ���T4_�*��-�M��M���G��L m�B���s�d��FO1��4rm��F`��Gx
� �iE�@��U0A\6č5�'A|0���T�<����� �ݓ���-?:ax2O��?Ad�|�+�-ݜ\ig�Z-w�W���y�d�>I��[�p�v}��M���?q�'A�s�:\�������3I>aD������O~��je�+C��!��^_�R�
�O��� �)�'M#�4Sˋ�<@�I3#��.!���'>^�����\�y�BT˛֢��x��'&<,��O3ɧ�بՄ�CJ�aB�L4[�(9V"O*}X�4<G��!�3k�0���/�h��DR/݋h}�8�sAқ+Ű�a6 k���O��kt� �3}mZ/s��
��4
(*U*ԭ�+�'o���|�(�.3^)0�![	P�l<�<	0�VP������X@֘��
;@Jf����[��:BJl��5�3�,_�����@�>�A"�EŪ�0C�*��РcJ;A���ʃT���Vґ�"|B�-T�\��ŗl1h�Ye#�%+��ոi)a|�
;b���҃ͬ#�Q[� =���R	�'�$󐠞4x�a��陇���q��P"�x� �4N�]�L�yK}2�Lі;�T�b��UO�"FZ�M\
�P���bt�3mD��ybJV�&�֭qaaǧK;��"T���4ıO�f��u�'�PIrj��J9��x�L.N�D�K���D�O:��O��SA>�$�O�4���oi�Dc��"��T�[�\Aax���#����;y��A{��'@��N�=(�B���L�I{v�(�r��y����M�X��aIK�o6b�E�^+�
�a�O�<����=��T�t��ܓ�̒iu���f��"�?����D0��|�d�'X��B��j���L�a��R���ē�E�9lZȟd�'��OYL�H���7`O:p�&V9)U�p��h�Ǭ!�S�O��qK��g���];�+j ?��N�i���:X�"BL N�AB���'�Ĉ���������O&�%�"|*%ܢq=�8����p��R@�Bs�<	��M<@G�d��
�,OJ�z���d�'��}� �H0p̤۰�C��f�B'��"�M3K>լ������I4H:�iS��0#�iYs�.s��c�t ��=LO����u�(�m�"0��ʈ.|az���#P��\���c@0Ⴏ[�:��'H0�����Ϙ'(�Ei%��a~,5���;*�4�
�'��d(���,�(}⍄r? �)O�!Ez���N>(��q'�8z�Q�d���� C�O����O��<�+����
S�a��h���E�g �T���� �y��~"N�%]t����Jl���:f��M�PaBY��}�db�E��P�#܁�^���ˌ�\!��۲ b��$�OX�$�(����$� ͧ(Ϣ�І+��{�|x��(��?D�dAm�T��a�IߗȢLZ�;��覥�ܴ���5A�p��O��	�Z�x�����F�,��Q턇2K����<���?q�Oᠤ��?}��'��z�iXu��%ٔZb4\A�3�'��4�Gh�.;�ت�,W�fn�7�&X��k�F�`�
T`G�ܻ�ax�h_��?��j���'��`�KFV�0!��bZ*n(��V����O�S�O�,��O�T�Z h�g"���*OX�=�|bղi.�a�1�H,h��2�t�oZ|y��om66�O ˓����O�(�d�� 5���LU^����O���N��Z�`A�ZR}2�'u��U1�,2��E��$�j�4���/ ?��.E�2�0�c�eR�JP1��T\���⎄j�vq���>�6������$�Mӱi[r�ӆX|�9�Z�3;JIS�o� &+L�OR�d�O@�=��Si�=[�U�����0u\ mD�c�|�nq�I�?Qd%زK�D���:��U�%�U��=R�N	�?�g�'�F�"L1��X�/'�f��'��X2�D/]T�
�S�^���'w&�3��@�p���B�Eo�A�'Rr1�扅"Z����%O֪O�J��'��{5���m��	u*%r����'����e�:��\a�l=B�Dؒ-O�y��'Լ���A�+wb���?�ā��� ��S�Hׁl$�+�"��d�v"OT�CAR�\�@�[�S)k�8�&"O��Z�(��Do��cЦ�  �@q"O�����o��Mq�D8i����s�'f^=h�'̂D@4�#f����B $a6�k�'�"��O�]N�i�G��u�M��'��rfB�^h�HBh��?�p��'����7o\�-:�$�f0��r�'Ty���T+R+�hd���!}8���'Blj���hc�1D�Œ'�@���Z�$Q?�AV�P6n�l G��N�\��O"D�Ԣ!�1�E� R��h1SJ-D���c�*#��0��D�\J朢5�-D�� +�u@�p�N·j^�<�u�6D�D��/ԠGo���H@��a#�4D�� 7�Z���P�B�`1Z�2fG�OP�Z�)�k�<�h��S8_R�*�N�Mn����'��}iȈn�te��,��Q���' N�Y���:o�h��J+K�����'o�����si��P7��D���
�'kB%(��߼A�A���Jz�J
�' L�b1���kD h�.�F^��A+OP��W�'	����/>-�={�FV�:�B���'�X���G��f��pU��-����'W�T�Nʐu%�x9�H@ #6t	�'�T��#h�8`t�4(U�W�J�ш�'�I�ӈJ�H�4Mʄk�n��@����%6��,����Ju*�h����NlpH��K�|=��Z�B��=D���T��KrlY/�P�ʴ�h)���F�v(���߈E�l�:
u�>u��vy✻ƎY�8W���E��3����ȓo/�����ƣD��m����B0F�E{4ݨ�������Zc��)���	�t`�U"OFy�#��*�b5:f̅=i��G"O2%��hZ�7Qx� F��<�L{"O�uZ���GPX-y����Q⒑3c"O��1%!��0�R�Šѹ&��T��"O�<j���;=\����.��U.����'u�A(���5���C��V$=R�s���(���ȓv��\B��U'm�Ƞ$��R��ȓV�����H;�м�� ޞ6�$�ȓ4����D�H$4�p��
��4��o��$
���F��WM�f�指ȓ+<��%BH�۠�kR%D�
��'�x�o�^9����G��BL	S#T��Z~��q�jH�D� ���S>=�x�������X��9�Ro���ȓ1$�����+e�`��A����� E�<�WL�e�i���;�T���De����=�j�I�.ʬF��:1)ՕZ�B�	)_�ܹ�)�5���׀��=B��!�XZrL��@���#pb�nB���nɱ�Jܒa��aE�ҜjFB䉛��;� Sl�|b�*s�NB�ɲY��Y���D�!s�1js�=�G�IW�Oh�اgŀ%'�\:U�>��)�'�0mi��4ntb�`eT�bm"̀�'���)u"�"*�pA&K*iD�A�'*��@TgS<��� "��n��0�'��}�c�R^rl1W��kn����'Q�=�����a"�U[� �d�}����Dx���!�P8��m5�v����W��B䉻%����f�rv�@��㔺��B�)� �ʲ$��-7�|���2�6ݪ�"O��*ҪU`�L�VcB�IRJ�	s"O��3�O�%
O|�`��I?<�DP�"OXX�D�
MP���G��,W9���sY��b !�O�����i�@$(�DX�1Kи��"Od�*eL�K��@��#�.oܼص"O��*� ]�"�*�x��A><��Aa�"OZ,�%�Ϙ�n�2#�ǸXVB�!�"O�E�B��J,T�RK�]�`qhs�'c����'ˌ�t�@ n�h��L�}�h��'�4�@�7&� �+
KFN%��'�\T"X�;���'������'2��vIM&a!ށ�u�X��l)�'K�.9(�4x�a�(P\=��Hh�<�D7x4JUR&i̥T�����b�'u�����)�
D**E{'B�n�R�������!��A�������Dq,���bH�@�!��֟nyB,{��J;�8�8ϑ#j{!�D��q:d 1�B�v�����^��!�DO�c��[�Ϫ���g�<�!�d\�6�ԠBS X�R�V�RT	!R�r�ҕ�O?a�3��2��hp�kùl��9׉�Y�<�B߈�`
���;{�0�V�q�<	��=/N���'B8!�؉Z�-Mm�<)� �W���2�NY�#�h�<i�ӻ@�n$��	�ܢ�
�~�<AUi˓ Z�}zR�N0g`=�G�|y���p>��� ="��@#a݅6�%�d#|�<q��/���QR�@�����!�L�<�c�I�<n�;Q���2�D��`c�`�<9S,�+n�f���՘i��y��Y�<Iшڒ7�ޑ!��֔ i������Vx�dbgc�����A"s� ��)���iQ! 7D����hY:7�
�T�Y�G_�%��h'D�|R��K�b�q $�7I8^�Q®1D� �W�	(�0"�˖,?�^m�s�3D�S *����X+�j�1G�E�@,D�h"�ً�\L�K�3�D\p�,�L�d�E�T�E�0.������bSb��y���j)f�b�Z��Хz�-[-�y�L��m�>���;_h�3�O�y��#!p9R1��7o����yAJ�ĭyR���5Hx� �_��y2B�&*�5�i�-��ࡌ��?�U-�\�����x�  1l*�'�NH,8Yǧ+D���)P=]���#�
ȓw�;D�L���3�b�r���/M��0�'D�x�t�
:M�EQ��-���6�7D��K��	G�a
�c�rX��V	4D������?Kw6�2JJ�s�l��c%�<!��W8�����ǓA��X�Ӭ�5R4$��2D�TB� �~Μs�N��S�,0g/D�XK )L�I�+�ޥ;vN�	 ��#�y"��b�1��H�4�5E����'���-�5G�6�Ar"�&3h���Y̖`��q; ya�	�K���'k�7*5.h��D�<S#�V�+:��qbj�$W,����(��CP�6�Ja�g�U��x��ȓ+��ж��lD�.��T���^�Z����wl~Db珓��d�ȓ�D)��:"'ܠ�Bfw�=F{ߎ���BT��M��0�p�a����?�  ��"OD����25�U���u�J��"O*�ŏ�90ZF��$дq�"O� �`����V$pQwB)un�)�"O����_�3Ѵa�1���M�L�"O�@I�@�oҤ��u����VQ�V�'�� ���nR(iQ���4�xǈζrunфȓIc��1��TB�Ѐ+�lٮ*nX�ȓ:��*��Oc�u#QK#?�y:�hd��TmMc�Q�h�p�ȓ5c��W�E�d���zT
�&��ȓWX��Ѱ͈$ZN��r(�;	4��'m����1�d�Q�c�¤��=���(�9�dMQ�0��kĮ�8�ȓ+�Zmӡ�Y�&$�Yڱ���Tq�L�ȓB���CB
LI����'Y$����E��i�����nd���$蕸`�~0��IC��ɺ1`���h&ec$�;�O8$C�I�zd�����,��|�P���aQ&C�	(`��[�Tl�m��!O@C�	�-`h�;ƩKK��h��n�bC�I�^p�$��-�
�j�h	/
�XC䉔v��BB+pN�UxC�ţy�$�=i�J^b�O�~DxTHR;<N�B@&�1� ��'�x�R��6e jL��ɏ
n�Y��'!|����[�_���O �-��1��'P���4�1jAR�C��Ѯ"ef(��'�0Ad���=�mH+c�q��'�<������7����H�i��'��H����S� ��C��mp�c��2Ķ���X߬�����<��aDP�>*���g��IRg�7~,��s�KM&#����N Խ�� �҂ə��Q:$R]��Ғ�#��<^�������6b�]��@�A��<6��h��Ʋ*h,!!���	2����q}��%��m�d�c҆ϋ>�!BG,=�|B�I/�tL��k��|��̚��C)bB�;7� C�L60Yƕ�WH�^�C����y�C(!w��	�
$j�&C�	�?�`mj��D=t�-JѢ�u�RC�ɉu��X���5�Ƀ=Z*㟄K�4�S�)��E7^8�K�3]����j�55�!�DY����׋�<S���ҭv!򤏭w2���h�v4���
�'c!�>xٸ5['HЙ4��8�@Ћ�!�S(i@���O��7�H�k�!�#�<�H�KO��Ua�성�^�I���"�g?�a ��B䈘��G�� �-���V�<Q��@q��`qdH�tt�kw\]�<1R`W)U�������+ U�#��W�<�P�\�EM����Uz)�em)D�<@A�I�"<�p�EH	/ъ���*+D�ȋ��
+�6�	�'D�!y~��Q��O�]KE�'��IIM�\��P��cЈ(jX�
�'�\�aH#�t�A 若/r��c�'.ĝ	�;l��q㋨%�h J�'84���"�N0P�Ol|�'p�Iم�%2�V	"���<�� 1ߓO��O�� 'dK�����ǃ�"(nؚD"OH��7�m�]1&�\�|�z�Y�"O�؁��>d�09��C��bl��'q�(�����p�~��'�A�e�8�Q�'�j0"h��r ��)�P$�'�r`a��K@���8gMʬ����,�#�O�'f= 0`q$��<5�ja��ņ�`+���a�ٓpG(���8+����^Nɸ� �7RH(<�� ��1��S�? � �b��@�)7h\�V��"O �xcCX?W�N���TgB^ �"O��sAǤ`6��`Z7E$d�2j��O��}��XB�(Jwdֲ(=BA�%\�2�8�ȓ\�:��o�z���ˡ
��f���ȓz?
���E*<1�S�IԨ�l5��=q����g!s�d���f�xRbP�ȓoņ���T'��r�J�, ����M��� �@Z���!�.A�h������~�����Ff߈����-.��P�k^�\�!�d
+d��8��n�:f)���
VVL!�����p�$�ɵW.�JQ�b!�d�2&>(e�6E
�g�.����ho!�䀚��d��L�{����n�ł"O:)Qrɍ�,�(�v�ŅPъ��f"O��[bZ.G��ق�[&a���X�"O���V��H��g�<�LՉ�"Oz)�T��Y���� ��W����"O,��/Y��(�%�N���c`"O`s�m�1b��j�
��|�����P�(���ؖ'��j̧�M�w(�2w&<�E�V'`:xp���$�0p�N�K{f�W�Y���Q�?��@�	B̧/5�����Q��L�d�B*O}*��C�i�j�	��P���'���'���hR��%�24J��P��
��,���c�.�d��z��y�P���?7��R ��5f �L�­����I�����H\2@����� �Tʅ�<aXwVr�'I���'���6�D��6�,4̼l��ɦKu�mi��'^�ȋ'UB7O@���ޟ�^w�P�'g0.�{V��T#܍C���	 ����>d�����O�8��O���'���O�b���A��3Ī�QJ�|j�d�
�H�䞳CSr�'��g�'���Q����u7�m�Ѻ�Nl���PD]&w� SeGeӠ�	�k��D�O����?1������4;:��a�
�@b�][���XLfy����<a�Fʟ��'�u�'�����is�,�Q�(m�T���W��M���!1|7�m������O��ď"nv�S��G�ޝ�C�R�2M�u���C3^�`�ߴ2w4�!�'�xx���?!�'�?�'%��ɜOu���!��nX����Rz�(��i� ��'�������)�>I���8-=2��1i���X�o>B�I-A���N��Q��B� ^�26m�O��$�O��d�O��D�O���OZ�D� �αp��
�-�r���V|��m����IMy��'��O���;}�
��B�N����$o�,^��b��'��Gy2C:]�2AC��Nm�#R���y�iE!�89䆆�sgP�S!��yR&��L�hc]�8�t-p@���y� ��y� �� *[��w�G)�y2*��V�#7�ۅ��jF���yR"�oR�Ha��u�%���y��A�P�ber�rL��H���y�h�<�������J@Z�[8�yBa�,��9�Q��aV�1�i���v}��Ò�o�h���E̝Nхȓh�z��o�F�V��%NN�=O�$�ȓ��d��khIá��fA�d�?9�L.#$�#�4%
Ȑ���A�	۬��B7�h�"��8Ir�ٰCH��3�.X*P�s�F�/�$�bN���cf��"}<q3DG �l�Z�
�4l}�Y�ņ21���xR�R|((����SxQ���-!���dd�u#٘����XQ1�|��� x"�
��|T	�v��y��+B9l��mt�l<����y�OS�'T�\ٳ!��gFp5ap�Y��yb#N��čS�a���*��5�yr'��[�����^�'��`���R��yR'�0tc�DK�
��%.dy���yb	�}����J�|x#�ފ�y��Q�K^tܹ�H�DU9��K.�yR�� 
0�\s�����uH�cͩ�y҂]k��0��O�>0�WX��y�EZ1{���c���M)���B+Q�y��$'̬��Q�R���Q�E��3�y�۪_�8��v�ȕ=���v�6�y
� �J@E��RS���4���|��Y��"O�ؙ��I�e��i����znX�Hu"O�|ja��/B�����Zk���"ON!�Se�Uj���-R (Z�"O�2��S�\�ӠBT�:�B1U"O�43��O2?�azq�R\@|U�P"O��7ODZ���8KV�P��I �"O2��T�.�ȟ�Zj�!"O�I26�?L���Y�&�xM68)�"O�tp`R70.>P��E���٩�"O����*
�5$��Q$�s���&"O�(IakZ+�2-a�����HG"O�5c
A3�	q�B�-Q� I��"O��(�*J&D�Ef��h��(�"O4���C�L$!1t⎚¸]�"O�ͫ3��4c���s˅,>��3<!�D���RϚ*h���1d
�CU!�dD�hOx�J�(͜U�&	)ͫ\�!�D��J����b�Ѻ$��!)�hͩ>!�dI�Im@� ��CflNt�@HԤ�!��Q�Dm&X�fL�X��æ��'�!�d5@�HQ7ꏒW>�(��%j�!�$BQ�4@���k�|��$AW23g!��& H�����ޮgն	��N�-H!�� ~��-Ps%�}�:�Q�-
11!����x�TKK�����Ǣ9�!��,\3r����I�4�!aƫ!�$�5=.��Q��P,?�~E���G�!���"i���W�&f�=�IEk�!�D��k^�&�Q�@I�e��,R�!�$
tO��QbȎ�j� Q�TH��}Y!��Q��f�#�I�>D�6\	���^s!��>�d�R�ֱP>4%�����k!��q���5m3ve��DK�m!�$�'Z�}(梐u�����/g!��l� ��'n��K���� �
5+!�$�7:�\"f��!��lX�Ȍ�mo!��,290��A�]�>��fJ��n�!�d�΢�����$��8��HE�H�!�)|�9V4��tYg��#.�!�$յ:W��
�(W2Ր��9sl!��ݐ���aǗj9�T[��� 6!�D�3<D�#F�W4B	��CS�	?�!��wj��Z�޾�������!�$UP�|��Πp9 D0%�ĿO>!�D�>M�@�u�Qb��.!��Z�S@� ���u�!����T�!�d̰|���3ժTJ�`i�%]��Py2퍒Lp}�]S�-�PaP.�yQ�U�pd���"J�X�G�ۑ�y�n�8�&x�S	��:�N���d�6�yB�-��)�ր� 7f��E�Ó�yr4�I��E͡2��#P�Ý�y�3�r Zׁ[�8z,X�.P�y��⽀�E�=5�\��F��yb��5��e+��Ћ]�ȓ�� �yBȋ9o1r�K�kT�(8���aZ��y�e�9TĘ�0�E''F�D�&�C��y�π���`�E��4�x#�͙�y�Z�zx�2c��$��2-��y� �:e]��Rb�x���r"��y�K�a�����A�o�zX�@�6�yɉ9X��B*
<{�AP����yl�(�u����&9�$�ѣ���y
� �X�e�2+�u�%�_�U[��	b"OF��R�mS6�XrjF<�D�;A"O:%��q���y�
��v�� "O���t@��J��K
����Ʉ"O�y8�$Ƌ+R��Jt(�]��}��"O �`�����xC ��/W2���"O"���]
���Cń�=m�H"O�-� ��h:%���;wr�ó"O�h���ѹD�لb�_��E�"O(1j�'O�z�v�rt"_//�bԒ0"O�Qi2�x��@IS�b~Z)�
�'��9Q!GT*+�Mۀ��0�y��'(v8�B�ȼ6��9 ���#-�d[�'*�p����Sl� e.ʑ�H�#�'��ct�ݵt�9�'�Bw��)
�'��=(Ba�Pft�yvj�g:�=��'^����) �z=J�#I^U�'�D}!�]8��I�4��-�te��'�,]*�c��������0��|�'�ƍ�`ưYF�x�TFG�����'�^��G(gk��#!B����'��Պu�&�Q��-3,�C	�' ��l��3<�EJ��&|�L�Z	�'��g��RA��c���B����'�NܙF�53,�Z�ͅ*d�����'���0�ג@�(�����^�4\��'�Cc>T�l�Y��4�D�{�'
@�!� S%:eaၬ4� ��'B͋dF�
K�4�x�Hă<�ʸ�
�'�z�2Ύ7Q�$�3ć=6(�"
�'Cz��KU8��Sd��
Z6t�	�'|�L����h��L	�|�2��E�<Ypl
?�v 0ƐSl����~�<�Q�%E,�:�&�U�2�t�b�<)D*Z�RR��@&#P�M���@�.�X�<y֬�25/�I����+UѼ1�+Q�<��P�b������*��=�roXG�<�-̙F�^��#�&.����RF�<Y��~fT���R�8��e��D�<���Ђ�����D�>T3��D�<�s�޵+o"�j҃_	6�R|R��D�<	��T�#�bD�燈q�� kU�@�<��ŝ�Z*��N=H�`�W/�<�p��u��� b�Ճ~>y�Fw�<!u̞"!���-��sw"��F+�{�<A&I��{ڜ��(�<e�N��(W`�<iGcҷ<�$�`�D�)�-P�G�X�<���5I0��z�AKk�fyB��J�<�U� Xh��ƟK䈈��)X]�<�bjpL�#�FJ�z%%LW�<�ǅ�h�@aPb�v���S��T�<��W�\���cU�!r�`�	B.�R�<y�5-"�яßC�ĵ�s��W�<C��h� ��o�_�LQW��X�<1s�˒/�Hid%A�0����s��P�<9bfJ}�t��xlv��g�L�<QƭO�*�4�q&��iP>HpVJ�<i�I�:6qa�*[J}�t@�br�<F	��Y�F4s�(I#�L�x��s�<1p	Ė)(���t߻m^JM�e�q�<A�C<9zbY�#NY��8�'�Bm�<It�f�T8�g�<n�5�u�o�<I֭ g$���@�d��Q(���B�<�t�Y2C�~����Tz�A@ge�|�<� �5y�+��4��U��s.$�"OH5��� IC>��A,��^�	r"OXU��k_�8��h�'��{r"OxlKrh�1ur)�-�#x~�g"OLxل��z\�0��O|�RQ�1"OlU�	Y�:�^�1�}Ӱm�%"O�I��
20lِ�N�]��4�3"O�`@��O��Q��6 �q �"O�I�t�G�}�9'�>�!F"O|A�����z��e��&�$f��+�"O�j �1y5���F�>lS�{"OP1
\_1�j���7f��"O�5#��ɩ^�I�`���R�J�"O��K��(� ib��`�D��"OR�2蔫4"!�D΍x��H�"OD [���:xT%���N��S"O��(`�~1ذ����6,B�9A�"O�$���<��`�޲8B\��"OV]��0�����&�,\zԐ�"O�}����p��E`vD\W�	��"On�0F�ݢi8X��bO�G��d�0"O��Q�"��2���G�������"OB�Y�+�??N&�J"C �B "O�1c�
��W��S����(#"O�ѓM^�]�hP@�ѭ	��*P"OxȘr�X9}R�$��O��	��"O.���F��o]~U����V���"O��t��"5�� �5#��Fb�X�V"OB%�a��(Z�B=�왱?^F�S"O���sĀ�8�Tpr��ɤdC�h�t"O,�:&�ڳd��U�e2�D"O�D0����b�u)��X�~��M��"O�;`�I[�*yc��
~��"Oʨ�F�J�E�(!�� D��a"Od pǪ�4���ņJ�x�V���"O��#`U	w���Af7vp��"ON�Z�>j�0�9d�P?X��"O���������������"O
��eY���MAV��4"O�YHf��`Q�-���A�EѨqy"O����N��GѲPx�͟���H"O|	huj9S��Q���o��L�P"O��c�T�'w����i��S�xQV"O6�2%���(̻d��8Y��P�"OD=�&KH  �2W�P�8�jH	�"O��L?*�X×f
Oۂ!Y�"O���w�H1D+<􉤅I=��YS�"OT�cC	�6v�fQ	��þR�� �"O�U��lU�&���#B�
m���"O*�Ҷ��&Q8d�S��̭�DQ��"Ol��C�ī8�TY��DY�7�z]	�"OL��Wf���d����-Ԯԙ�"O�y����04�H)ySCv��(q�"O�}��g���� HB�>Β!("O�1SíC�6h0�Г1��"�"O�ya��<t�e���� Lҥ5"O�)����/]ƴ�ccZ}G�D���$�����TKY6n��3�a�8��'���"Ad:e���"gS�n>��'+n<��݉,��UC�d��)Y�'/�];�Z9��X�W�V�nB �x�'�ּ�@Q?ln�|iPO��g<�)�'5^w/͔��`�E�cg��;�'��`�E��vzV ��j��P�x
�'���d��6?�%�����[r@U���� P��LÊ*��[AP�҂"Ox�c)�O�"Հ@����t"OjU	�@-P8�`*sg�8���9�"O�a&)
�1`
���Z�p$�"O�$V�@5�~ #��H5T��h�"OtP"M�b<A����i�|�i0"O��)�'�N�*8�äM8/&�0r�"O��Kv)�;b<)fD��S*���r"O��g`�(����*�;G+D�c�"O��bg��z��
d*�,Y ���"OT�{ h˥��q�j�"�dЃ"O:!��-�Pې���ʹ#�NT��"O�c�a�-&�A{�N�6*��rp"Oj��g�>g�tRƮJ9���i"O1�.ק&�<$��v�؍@5"O�d{�)�3��=�&��\UpLrr"Om��]���}*`���obB�	F"O�<��-&b�����9�"1P"Ov(vgJېౕ��+V���V"O~,��WfS���ρ�{�d��w"O���tȟ���)�ωt�2�8�"O�jK���胷o��D���V"OTey��Y
�t9�HQK� �D"OB�������,���ʀ3X���*O��[�-�H��܉�ܾ[����'� ��ܥS�[��C�J Y�'����!�z_����F&��
�'O�� q/� 3�u'��wxn��
�'^�,���QyZ|9��y�X���'P�0*�S�jNb�ڤ
��C�Ph(�'����#�;[~�U�!/[�Ag܀��'��!�3!��W�H�"�AFq���'<���t�F��|��ʕ:D>���']�!O��F�z�E\:hڎ���'N�Uk�Ο�Fd[�J>f*�1����O4?�iab��nv�	g&�b�<��9u��h���h���®D�<1�]ʸۀ�з3�͢�_A�<�!/JY��J���^(�\�<'�.q��a�f�)��Y(�+d�<!%��	�H�P�@@މᓫ�c�<	#� =Hٛ�L��[��E���t�<� ��}�r\�vѦ�!�u��i�<�2l�s�r�"@��9���2d��@�<�W�\4g���)Am��Eu���h�t�<��̋h.��tǊ+^�896I�r�<Y�IԈA��\�sjƒ�"lpI�e�<���X�<�pZ��Ն�DI Bl`�<��̗oD��b� .�`���<��Fər�`�b��B�h�*��E�<y��جq"n�c��fk
��QF�X�<!S��.�!GD�.�\�x�\�<�gI�)G%̻�Þ.D�<����UW�<Q�N�)X��-9�,�:��SE%@W�<	�ծ
�|�!�eĿu�XU���\Q�<���|���C��ih����EU�<i���[��A�M�=���1�e�o�<����.]��(���Ё	U$k�<�ģO=N&z�` ��z]���b�Fc�<Q���$B�ʀ�hñ<bly�n�h�<��ԍk:p���ی,�nQ���X�<�򯖣n���c�N� 8�qa��Q�<����2wph1f��'��2Ǆ�h�<�`Q
P�|:f�$��ӂ�`�<� P�r��_�V�P�d���"O���G�����:p��">D��� �&����e	�By�p��G=D���`hȵZ�bցV "�����9D�t)�֙B�0��!�("��6�*D�P�,��V;��s�׾b�	�@�(D���m �\�1�҇}w��6D�@��C�,�Z�j��%6�(q�q�5D���0IL������O)K�zT�)D����_0<�TLH��;>|2쓅�(D�8EB�#�b�TA����4D��)T��*'U]AG�Q8��ѡ&3D�����&B�TZ"
u��qj6�?D���$G#���� ��!@���?D� ��	�ɂ HЧ�}��I��<D�<	�R�*�Kq�T�dN�`�D/D���5�D-Z��q���Q�6P@`#�9D���Q���(찰z�͒�UX�́�"2D� �� ���S%�ђ2?leP��0D��P3� :^X�{@�P��F�Y4f?D�y�e�N���g� |��C�)D�`ɒkH�}@�-��jɑ}&�"7D��yP�"D�$�BV�ö2=�Fl5D��c"i�;`2��F���4�����'D�0ӱHЖT�f�q0��=�@�:D����'�D�n�!����8���x��-D����ۨyl]Z��7-_�@ش�-D����г/�<�ZVB�����(��6D��B������1z��6u�beH�i?D�d��D�9Q~P�+c-|��q)[�!��R~���h�$.=�E�ֈ8�!�$ӯ������	"��SGo�!�P �u�䢚���Q�1�{}!�K�(�VA�7O�A��̋�@i!��u��y�M��-�nMY��K�M!�H�t� tX�H;
�<r@�+0�!�dM>ReJ�b2�0.��:v�!�D�M�~Q
�U*��A����s�!�d�;1����oM�x4b�&�;�!�d[()��=S��re�S��;�!�%n7r��Ü/w(@y�I�"4!��@�x�lx��N�Q�l��"�؎#$!�$�,r젲"I�D�2a��@�!��V��tbS"�j��4��(O�)�!�	�m�)�����~�sD-  �!�ɾ.�T��R�I�\�(��,��(6!���`�c�̰;0�<�3���C�	;�R�)t)@�Y^���E�-�B�ɋe~��J�ϊ F�����,�B�,̋�C�	�^�B��4*c�B�"t�.uyp��'�>t�Z+4DC䉕m�X�HNJ0�nE:d28�C�	e~���2F0�)Խ�B��2j:��+` _)L�Dief�~�B�	�-��m�El]��qU��HCRC�	�SLD�й0A�f�0TΎ�A�1D�X�@cЩØ�0�#uHL�tB"D����lT�R��\���SifqIT�<D� 2�-��<b\HD��&I��a���&D����>n��aW;?�d��!� D��P�M�
�({�e�����h7�0D��Ӥ��E�����S�]2*̪&0D�P� V3/ �e��S�"$�9�`�8D�� LכE� -�`o��B�<k��$D�� v�E�h�E�W�NM�Ѓ�"O&���DF����ΰIe8��T"O|�0�/�f����<�B��2"OZe�S��۬��&��/:2"Oh����N	(��3��(��:�"O���GJ�$��պa
ǝu:�*V"Oڤ��#I(s��k6i�3C�-;�"O�p��C9�j 3�ńv{"�"O�����"M�0�c���\`d �"OH�a�K�5<~�Y0.X�3����"OX���f�\MB���&
K>|��"OT��`L�A0���W�����"OLI8�څ:�戹�d��B?,��"O:��cD
, ����
V/{B0��"O 0�2��/S���p��M&1u>���"O�I!��9��Ͳ��$.�$���"O��#ׯ@����Ri�x�&�"Od��`�4.ZT�s��0J:RDq�"O�L�U�ҽ3R���%fť'>|x�"O �⠀�_12%g����H#P"O�0C@*
X-�YCe��tS�9��"O��CBg�s�Ґ�0e�_����c"Of3�|��
�$�$Ԭ�c�"O���Gдfi����DB�\<���"O� R��4Oyv\y3j�wx�q�W"OLlxd/I(Z<"���J TY���%"O�R���D\FM��ID<YF���"O�M���ß0� �(�ț�b��`�"O�͘��A:b����o��g"d��"OŐq/�r�N`'D��rH1(�"O ��v#�5&l0�B���W"OT�s���gyxh�n�-2��
�"O��І'� ��#-�?�@�e"O���rkV$(��K�U�`�"OX���Ν3_k�كsm�{&48�1"O�=���Цhj���*�����"O����N߰%��`�eMά��`I�"O�i�+��tZ<�[�#H<D��3#"O���r�B�]Ƕ�"%6T�ё""O@xK��ϡu��`�bLKT.���"O�e��*�%zzj�8��\�X����"O�[�E@�um��C	�
C�Yx�"Omd�	%$�x�A-(B��;�"O�Q��+̊[�u���֛��ɥ"Oj�vN�(o,6���L� ��x�Q"O$�ä��D2��j�㈛ �tzE"O.x�����K�]J�"�k�V8�"O��:rO��z`�$a�ƒ��2"O�p�U�sXJ�:Dg�j�Fx�d"O�;PE.b�2S�ܢE�ؚv"O���.�Hp��J��5B�"O^I�:O)���C�{�{s"O$��,�:eMd��A�S8d��"Ob}��&R?�����4g6�3�"Oܵ"��(1(��9��G`'\,�b"Ob�!��L��c�Hx�Q"O�Q�3��!u~Xx(�� �ج�c"OX��C��.e��mi铯F_Vt�0"O�e��O
�	�H�u8�H�"OV�H%@�f����Ϟ>;4bi �"Ov}��(�.Y5�h	BoJ4�P�$
-Z�( ���f��ɫ#CC Z�'���QSo�z:ư�R�P�U�l1�'�܁��S�Rs��x�,F8Q$��'ń]��n:wl���q�BV����� ��'N�)�� '���0L2�I4"O���"���g�6库�38����"OP̐��Ax��� 7#����"O���@$��0 ���_2v�lk@"O�<z��=h��x�a�N0|��'�X�[���8�pX���n��'�l-2@��HW�)b)�PT&�b�'F%a���O*,��w�.Lx6���'88����<,�WkVG�6x�'�I�p�*Q��S��˛D��[�'� ��%J����i	S��A�Qh�'f��7�J�%`�<("d�4b���
�':�+��1atj��q��Z�V��	�'��,Q�m��t�m+k�&&ư��'�D����
W
��c���<���'�"���N%%����臻_]��'޶� �	�!Dt8C�]Tʠ��'�ȭ��Ce�<k� �����'��XB��-v��9G�Ο�@=;�'��!��Bĭ!/���v���x7p�x
�'t����΁�K0Y1��7{5hT��'@�,KV�W���(!bB�;b�:`��'I$�8QC�7>��dj$K��
�'�~ɓ�˟']���3tNԺ ��3
�'x���P+��4<�YV��y� A	�'z<�؇����r֧HZ�����',"�eǇ.aw�I�vL�Llxj�'�va�C���^�t��	\6V9�K�'T��FbĠ�6���@Î5Y	�'_.����9Zޘ;T�_�bx����'P M*E%Q�zf�}h3d��C���'M6���b����KH��A�Zu�'�ZͺW��+���ɑ�7�^�h�'���ڰ"��A�IcPe��&��'q6��7��A���(@_N�0r�'����Я�Ql`S�H'�
(��'m|�q��׊~�ޥ�v	�Y&P��'Դ������_g�l+��A���'��3TD֪h�LH�`�[#c�Q�
�'��'h��@�lT�p��1��Q�
�'��Y�aɍ*v��g/�0�F�
�'`�w�[a:� g��W�T)��';�,��V�\�v�ӧT�fD�<i���l9�4���P
�,x�%#K@�<�Tć���	��W� ���#q�C{�<b.��V��m�o��+vg�B�<��nT;2���6�G�V�K2�W�<�qjI�MJX� k���B�ccBS�<��J\�D5\�j��n�Hp���R�<1f�l	0���he<��v�<y�`�
)[����3K��I�{�<�r,����AZC���x(�t.u�<�"C�-5�D��$�f�1�AmI�<y@�C�U���(�oQ|Q8%� �Q�<�D�H�/��|�j��Fl��� �P�<A�`ت>��`�O�<~|�cF�Nt�<�� ���X�đ�|�[�*l�<Y�)MC��#dض|L.�@v�j�<�%A� ���,�H��Hp�bP�<��%o�2�3Ǐ�S���"/�O�<�W`T,B�BE	ۊL�R$C��
C�<��e@�rN�@�Q@݅%]�+W��B�<17�N7R	Z��^�-���:P
_~�<y����UJ:���E��0�f9aT�s�<� &���0s�����	�)�n���"O���� <]pt�A���1U�Hȣ"O�9�6
�R�-SJ�.���Q�"O�bP�ߊI�����_�5"Ox;��l�Zԩ�$�@�"O�2�I�a8؜�b�4SI�@�6"OP�yרN�w$���PJ=:?�$!b"O�d �K���H����/y��9��"O }�$@1�j����8q*�yR"O�9Y�E����I�ɚ&� ��"OR�y��ňl����I�xT��"OPM��aܘ]	�t��ھv��$ �"O�a�+�/wW���g�0u�]�C"O���LB�.�εX���{hfypr"O0H�ϭ����$D%i[f(I2"O
%��˛�~ڸ��pZ�x�"O~��*� �D�J��N�LX��p�"O����|��@ϧC!2�	�"Ol@`#OQ�{�D:7D�v��l��"O~� uE:��]+�mV�S�����"O�H�fě#�&�a#͆ [~^a:�"O�pb6��?v$]J6�,uW(x�E"OБr�'�>
W�t��&D�ZV�%��"O@$pg*U�<\<xf�S�\ݪ�
�"Om�($'��!�fI^�T��V"OjAa��(��`��`��!ЬE!�O�p����:J]�E#RA�v�!�D^a)�Y(!�1aX�-�I��!��/&`)���y0lX��DһW�!�䍕|�m�ӡ|.��"�05�!�B<���MûLoș˖�^�o&!�@�2�RM�6�e=�0G�S�!��?�H�*�D�"�#���!�A+w5~%�u�I6i4i�[��!�[�ޜڑ�WJ[Ry�h�"R!�̬H!��J�̙�"at1i�I\�X&!�G�S@��u���U���qG���c�!���$��1��R�K�h�H`���"!�d��|M�惨[ܘ�ӇE��!�� d{�U� ���>�֜2���Py�j�s�:��DsF����yB�=F.���cV� L�B���ynN�B =�s�B�i�6�3��B��yJ�\��$C�-�2��QH�yR� B���(5�Ob�H��́�yb���<�˒������F\��y�O@�{C�(�K��h��_��yb�_�{��S�P�}���vo��yr�Մm���!����w�DI�.Z�yh����e��"�z��=2�\��yB/͞�]��R�j��ls��X��y���	G�qQF!)UR*���\��y2�7r%�(��MD\��EDH��0<!���Ըh�PPȥ�σ_I��L�y
!��O�H��UcS�;Mvus�
L$w�!��_"!+�����J*l �j%
͕FS!�d�߬��f .3����� �j�!�d� �Ƞ�fň	�ڹˠS�?�!���ox�\�p�T��h�C�{!�C@� ؂��ɏ-z�Ę���O!��]Gp��!Uf�+5��>?!�)j����)~S�ܱdA�4!��~1\�R4.@�S��-#� �'}!�D ��]����yx� �$ty!�� ؁:�:�n������ �
�C$"O윸u���U�ȧ*����"O~Q�ۛF��:"Ϝ�x�N��"O�L⑍�+���B�L<�Jt+B"O¬zF�p�@��f㞟~C�mX�"O���wO�3A6(�#cƂm7x�3"O*d#U�Ĝ�5���:$.̓�"O2�s�J$A����!W�U@@Q�"OT@�P̝'H��#R+��^�D̉"O6�sC��@D�@��O9~��qv"O��CP��g+N�Wm���`�P"O�a�Bo��/���+��Ҹ�&"O C犋)T\:lH�J§_r�)�"O29�G�Ƕr�L�*�J�6d�i��"OlY8��� ((�bv�Յ-}~-K�"O
Xc���!���GbB�8u`�s"O��C�6��
���n\�Kg"O���ǫ��L���R�@�I]�,p�"O�@�f�,�����0?X`yt"O�يe@^;�ؼ�非!;�3�"On-��Ύr�H	Q�.BF}��ۇ"O�\�i�&DJB0࠭�9P���
�"O�I�"�Qm�l����1f��p��"O.HP�.�/����#�JǰA��"O�T���6���0�9p����"O�]�F���S��Y9�F�*`����&"O��BoT+-�r���F�
�^`�"OVe���,=���`��:M�!�P"O�T@Tb�+-�qP"eS�E=v �"O�lq��1��8�U��,3�A�r"O��`%���MVf�����!.%�@��"O�=P��"Q�p�RaQ�8k֭ "O�#1���G~�����<[c��AS"Oz�{�$N=�NL�#k��TL�8�"Oj�ʇ���U��yf��`��2�"O �r#J0(R�,�P*[�}Ҥ"O���rML�9_��c+M�CF��bP"Oj��CA���$ 0��'D�t�"OH�"A��R�艢�n�w1�ڂ"O�ѣ�#M�X#\�qD�®
���"O��c������>NEc"O>��%�|M���]�D����!"O�=��`��L��\9� ��"OJKtc�"�n�P��0g�
U��"O��EY	h�`Z�M�a̖��s"O��� 퇸l�`qc�*Wcظk�"O��P�Ձ�,!3�P�:(d= U"O�H���(D��\�fX�y`��`"OL4���+g�ɓkP�3+ L�R"O�ea��20FEE�I�pz<��"O�Xu+J�.g�ə�E&Krƭz�"O:���O����
�ReV�q6"O���"�T�)�Z	iSc\2o]��$"O�D�r
� [���S���l9�3"O�9@4�8iZ�|i2�9NS �%"O@e@�D2YT�Qo�=}D��"O��c���8��7�.��,��"OI�JE�/E�l�E$�"OF�hF�Q�6Z�����p�r@:T"O~��
,�����"T��E�"O�(@/�:)`$KE�9>�3�"Ol�)��&B5+�ݜr���"O\x��T�~wZ��D��:.��UA�"Op�b�KM�3E�E���K� ) 5"O� �8�ҹ,��y��BC�3�r1��"O�x�dJ1Pڔt�&BA*�N%X0"O蔨R��,:Kj����)�~$@"On}ȶ��e����2Ǩ�*h�"O:�iFC�w2��2�Ƶ��-�w"O���v	Y�t���KB1\����"Ona���� ����YNh��"O�9gG�HJ5�3GӶF�$@H�"O@9��%Q����g̓<o����""O�A�DD9S@dё���6��u+f"O��!ߟ}U�Iqg˦vin�"O��8$�tC���F�,g�qC"O��3Q�[�p#BUɖ䟪+G�Qj�"On�HD&-jB��c)>_^��"O\��P���l��1Q
O>%Ƭ��"O�D�l 6
:2��K�Z��V"O`�0�Fw-�a��<Դxc�"O��XVi,Ф�ڶ`ѳd�d�!g"O��[��ˀG��e�7U�g�����"OΘ���ɳ�
���
�Z���I"O�uHB'nYu��Ф=���V"O.�s�j�41 ���)�P"ON\�V��%'���ݨ�B4H�H%D��� +���ݲ��%�x H�a?D�i�V���TVm���v���9D�@���Bov���B+�3�0mya,D�\���
K )���HF�|��(D�@�V�M�g�Le�Ug\�i��D{��0D�D����TOXI��W=�@�+D�\Z��0	��8b�3�آ�*D����n�MD�ɵH�p�����%D��s!!��TV a�B�)Ĝ32
$D�X���-c h��2K��o�Lݛ�@$D��"{��sr�((��pA(#D�l#�ů3���8�'Z�H>ƨ��� D�pQW�Z�e���d��08e�#D����e�9S/,D�tU6iF�=�2! D���� 1,��=C�CT�%�$D�����"̲�2F��"U���j D�h���@�R	�(#6Oۄc&f"A�1D� [�C��Fa���"O�5�JQ��m0D����,͘��ԾkB�Ų7� D��"&��>7>t{㉑�(��% dd*D�� so�-)=�l+�+Ϸ�n��*D��whD1L*���GI�$� ��%D�� �Ǒ�63x������Q+�>D���$�`�!�F��E��:D�h�%(<4py`%�-D��UȆ�#D�h۱dX$$~VdY7h.FuV�!v=D���/َ`�ع��a�~!|�2#�'D��AEL	6���g�?a���*�$D���֨.��\�'�ݜ&Kvm��F"D��rա�1)�b�xׯ!�����!D�8�W4��TϘ-Aͺ鈗�#D��3e�[
�� Y�%V&u���G.D��9.ׂ �a	B̉13�ޙkT�(D�(��!Q޺��䦛>9� �#�(D��R� �cR�a��N�x�2t'2Ox%;�F=Zb�y���; � 	�'�,����/pJ�� Ǣ�[��Xj�'@x�htA�mƪd�.��L,��C�'���:��"s����ˇ�{��p
�'���c��T%k]�h""��ct�1r
�'��}+ת �0��z"!ڶSL�]���� ���l���r���׾���#�"OR�M��<��! U��c�^ [�"O|�� ڭtt�U���P�I�"OI��"�+�fe�IOk���T"O\����/�:�[�K�0���;�"O��b�Z�r/�aQR���v�:�"O�����o`iJ��{���"O�%�/��o�fySA�`�H�C�"O�;łЗ�D�K���m�4=q�"Ov��qΏ�A�v�9�χ��l��w"O2Q�v/CX�deY��/�tE+�"O�)ɠ�[�C��M�����K�N��"Om��]��qI�JW�q��M�W"O�}8�m��?0 ,z���&a�S�'��Ðj��m�\À�1)Tڱ��'��䡒Ν�UΠB�N:%Ӫ���'��ЅR@����h��*�'�l˵Bι0��i��A����'��Xc��̏9j�Z�JU�
�Ё�'�d�dDX@x��w��q�F.D���)�9@�S�I0���b�(D������W�@�Ӷ���0bX����$D�`��@:�r���/E��ذ��%D��h��Ѷ?5>�(D'��3��X��� D��ъ�;m�tr#� x����2D�����M�"�J��^�r�����:D�t�Ed�mI`���P)M����!�4D��㤆�D.()��M*��03b�.D�T�.��/Gr�Y`� B��4R2")D����B��b�ʣ4v-�Bk&D�\��H*f4N�9!ɆZ�T�u�"D���-��e*L谢l0c���@h#D� �g�ئ@��*�A���3�&D�Ը1�$@Ĺ��Q����$D�칶dʴ`Ԏ�p�C�5!w�K�b"D���f��`����N�Lĺ����+D� �d�_?,l�d(	&n0�&�%D���U	��x��(H6D]�B�2���#D��H�!��n0DA5(�$j2���,D��iS#SƠ	��O�������>D���P�څ��	�b�ƷG��8�%.1D���ǭ̋@L�̀pj �0D�t�qn��f ����U����.D����عA�����S6Ps`�/D��	7j�����c�@�P>M��*D�Ȱ��gg�(�ġЏ7J�`e�4D�d�@�X:j���в��<2N��r�3D�|�A�����	�*�1V�b�h�C2D�,�f�F6'
H�t@C�Gk"D�H��G�:�^-*VG�,#���!D�\�0��~Wf�ȥŨs�m`�� D����Ạ,)����^�PMr����#D��� �# ��PQhܭm�00E�>D���'F��Y�N��N�%Uu�@A��?D�u$�v���xÆ1������>D�H���un��S(�) \D(�'D��� ɴVU�eá���3iZ��)'D��i1�N�<	��*���QT����#D�(���F���3��ҡ���h!D�H� ��\��X��Υm$���:D���r��o`�`�̩>�&X{u*O�dS�
-1)91�ȟPV� 2"OR���'�7 ��1f�=��܀�"O��3#�1�4�h�O�{��{�"O� �1w�\�"K���-V�~�T��"On�����	MG,X�C�/W4�ҁ"O@|���SEXd�E�!rN�q��"O>\:U P�Y��H2����S��2�"OFX:��3�F�7.�lh��"O��S�/ޑa\Č��#��'�����"O��ċ
8[��yAbZ.|�h3�"O��XT���8ՋU
����H�"ONЧD�'r�f�U�r�K�"Ou���
�T1p�D�����"Ob���.��T�ht�U�6��\�"OlL�U.K}�ԙ;�JI�)��=��"O<l@�A� 7;f�(�T�N���"OfQy��:?�0)as��+"��a��"O:�@/�o�@̚-F�X����"OlkT�V�~Y9��4>s�<"G"O��:�G �W�BԠ5�˱`^4��"Oi���=QmX��_3Pް�"OfܺSJHd~��h@�7M�U�0"O�)ZQI&\ή���>xޖA��"O��'���W\�RoӼ�J�s�"OR�AF G� �����lŘE��ܚ�"O0�<"X�v��9[��9��"O!8E�2-r�4 �H!���	�"OL�$ZM� ��/F����X�"ODMZ4���"(���N�e��	��"O:U)�"B�b�� n׋����"OM"��-si����v�"O*4����a.�(��� �T"O��Zv��'oǸ� ��4+�F�2�"O�S� �%�L:Eg�"Cx�eɔ"O|[�T!q<dI@CM;aqi�c"O.�U��3��t8G�K+M z@XA"Ox}� ˏ7k��]�2ʬ���""O> R�fp�����G�b��T"O>p�F��)�L��E�
=�pg"OT��ba�r�l��ƺn+vH0�"Om��D>B ���dԪ^RѣD"O�<�,ވ.c��9�Y�i����"O؅q��¸y��� BN�D���"O:����"�\4p�I�i��t�*O*L9d#V�Z��pd�E�K�J�'��i$�� r�@S�ϋ:��(	�'o�@����<z�
�}֎�(�'/.@�a#�<{ia�N�$'.r	�'<.�
�	9��4ң��)~�bm�ȓ<���S�ѓB���cqEW%k&ԅȓn�^���JB�0o&P�L6o�����
M�dY@ďwZ�k���;?�͇�n�ᲁ�R2��f�8xY��U0�j�.��R�,$kP��2B@Z��ȓ��0�#Zn8�����ؖ?NҴ��L�8�k&���$���Y:�Z���t���B]���+D�N�R<��"���3�	9N ��
c�R�rԄȓ[Τ�W��XN���'�:����_LPz���!D�� jWh
&|̆����0h��%m*%�1�]���ȓ%�������11�  R ANli��ń�V�:��{�T�8��<��r�l�����k�y�P'�*���oO�0ڥ)|j��*G�_=(؅�bФ�r�E3t�`d`�eBD�����d%�sh\��aP��K�?m���S�? Z�ȑ釛8J8xD���^��4K�"O
 QU9/�D��b��2[��%��"O�m��,�DhB��  �Z8:c"OR�9�a5.T�s����8�{�"O�ȩ%d�6U�pܱ
�������	ߟ��GJZ�j����'��T_?���A�)Vȉ��P t*)��M
,���?����4$��G�?7�V�{94���|b��M���@Ji|���l�'����!?gr	R��w>e�G�X-fTL+�D�w�����L/b��u(�&/ғ6{���I�M�7��4�i�pǙ�iS2@�Ca�?m=*m�p!;!w��֝P��?�ײ��#R�k�P�+-��ݙ�2�OJmn�$�MKٴR/@p��lbA�脠X�4�rs
Z?q5�˄M/�6�'��V>Us�'��T��Ӧ��u��0b��K�AC1?U�C��IR�J��HK�}����_'f%^D`�I�?!�O��T���|	B�_2"�(u�"~�0��i�M���g�@�CWn�H���^$U!�k��t�dH'肕&\�]禓'���N��?��iS��S�c�ܴW�T(���	.*��4a��[uW���Of���S�,O\��m�5K�.��C����IŦ=��4�?ٲ�i_�غ3��Yd������?,�`���1s��'�P4	0f8J�2�'���'#���xmZ;^b�a1��8#:����̙4A�]� �"~��ㅳM4H�bU��ja7`�̚m���*1�E�K�I�
�r���0^�� ��dg�����e��CG�Fb�t`rd6%����T�:����/�>9L^�����:���?1����D1�mi�/�b�HCq���3��$�O���$C+i�u��Ǥ2*uA��F�2,(ڴB4���'�6-�O���T�'O�\��%�#TV�C��"T�̸�↕PdJ�A��?Y��?	צ��?)��?CM>	��4K������r�Wb�^d�ղ���)z�1b�*�3t�uZ���Xx 
��� f�Y{`�7	�v�r���`��p@�)0Q�����	�v�(�ă0c\���գ�
�A 7a޸f>8Y�¥�����qy��'��O$�'jU���Р�}� ��5BM\����u��!�7�Y?5���H��Q�V����1݂��S�i��	6�豩^wr�'���i�:ɢb��!G�z�#&���ed(�D��,�?���?�&DK	pЊ��A�H1v�z
��1Y~���M:b0�߂M�z� �&ߥl1<"=ɳ�N�!��C��Ϯ}\�Pa	\6/p(гR�E�J��ACC1�1��ΗS�������O4n�>�MC����Ʌf��y0�#�\�uh�I٤ �\t�Iʟ%�"~�	<2%�ӆ�=q*�
t�R�4nz��dʦ�h۴�M��	�s��*."	��m?A.(�qY���?�.����E�O*���Z<��aB�5t�D3�N�<|��� ��'Ap��Zs�A�1��i�� 8����uן�˧��\c�>a5䂤M�Ĵ���^�!x�ܴ�Z��E���nJpQ�#Δ6��}`!lﱟk��(G��dG�/�h�o��V����?!��i��S�SM�ܴK�ܠ��cB8����Ն�T\�=�����D�M�Y]�D�7�[~��Y����(Odm���M���Զ�,�ԃT:]��x�*MnYhBg��T؞�S�   �   d   Ĵ���	��Z�ZvIJ(ʜ�cd�<������qe�H�4͒6R64<�b����!$My�+�D��`����M�'�i[B�p�\�'x���͓_�������<.p����_�/Բ|ǭR�K��у%�	�.�' %�F�ҞK�������,���#�� ��B)\5���I�X*��+�>��Uh� YO^˓y�� ��5ܤ1��l;Fr�Jj�s��lڲJ��`�}�V�{�.�>�?�fE����GX��҇C?qix��㆔�,�~��'����	(�X�a��b�t�'y��c��3��4�׫eÞb�I�,<B� ��Vt~r���>���C�
�?���'0�����
,?R� *Ot�9ӂV�"��\Sc�X�W}*�r E���'�|EEx"H�&��°�K4CR|���� ��#<�G+�u���a�B���< p8�O�""B��O�ሏ��_��'ق,�J&N� �P*_h*R9�4zU�"<�EO5���*S���a;
2�aԴr:���u�q�"<�'n"?�G�2K��=�e�+n���q��my�WR�' `�?�D�"C�	26%G�"Y&+J�#<�"�6�wS���U	,B W(�#@��3Ζ+�1OR��DO*��,}�����A=��i����m�	�8#<y'!!���F?adn�3<� A�DX�'�0������8L�@��9�'���?��6�"c ��c��T�W�^�r�;�	dP�(�r�>Y!�	,��Ek���C�B�ԉG[}�!�D�'_6�Dx� U�"�!v���S2XS�Q��y�� d  �Q�<�LT�P,h�!bU�P�:�[��q�<	�	.XP�S��ňb�y�"��q�<a��ݒr�&)X��
�d��f�[l�<�I�7 :fa�k�8���ʑA�<���6N��Q�g��V}�`�+�{}�Rx��	���)a��FF�_�����%8�O������<�N�LѤ0�&mj+1�o�<qS�D�;	�-�DI�D@h(0�KZC�'�rHi�0�k�uc2�1*=
��� �2���O�����G��d$}�ek�.����N�i��O?�ɝDB%�� I(�:X�R�2"�JC�r�($K����
�2#/�0J�$��I�D;�@��$��#��lx��b�ߣRt�Ň�&v<�p���A	��$�\4 ���O���b�(@)*�!�92A�Ѹ'�J�D>�Hr�'IH�    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �   ~   Ĵ���	��Z�tIJ(ʜ�cd�<��k٥���qe�H�4͒6R64<y�b�l`�V. 'Oo�tۖ�h�B�h�#Ԙ26-�Ԧݘ�4B,�D�<�O\6-c�bb��&��RA��M:d�R�A�F�B�҇��)�qO��H<��"��"�v�2�4x j���><v�Z�+��[i���'���(���'�ȡ``J��]\0��'�����A�9��;W-�1r0�ӒI��_��
�4y��5s�'�4�v.\�<���|"�MZ������z�b�Y.8$4]�P�άyq��-w�x�i	�L���:^�DH���;��q�af�!9�V
%aְ���#ď%&��ImE�1	��l,҃�O�ye���[׶�q�S����,�(zb�K�(W�G1��Q�BXp�/��R�qOҹ*���[�@�|���A?X�^�"���+�,Dx��Bf�'�P��'�D�e�ȉ*yZ5��%;�
q�N�Hi��!)�qO`��
�
o��y f��6�q�2�i-^=Fxr�T�'��I���ط5��a���hk��_�'��c�����$ ��?!��p��	Ŭ.F�q_�,�`˓k�D#<!s�)�	���4�A�V"P<�kV 8"F-Iq�	�%��t�B�'[�-�u��(i�4i��l�J��yR�Rb�'j�%�,��kP$��Ġs�Z4[n����@��s��i+q�'����7O�"	��I0�d��wf�>DJ0��MyR"^�[��%� �|r�@?�-A�O׾�a�#Z�`E,%K�Z[�O�|���%�(Or\�N�(�.�K�Tܓ��!O+.��d�>��!�4�#<��
�T��qC�Ap8��c_|�<qR�� 2  ��D�U�s���P9�9{�k�v�<A�I��8hZh�$��X̮���)WX�<1RK��l���Z2�K�̈���Q�<�⋕{����U��c�:9���U�<y҄�=th�!j�fW��F�`4D�O�<�W�P$b$ք^����aV�^I�<�7�G�*�<0a)�)pnY�BO�D�<��I�6j8t��3J�2�����@�<�3�Bj�zͲ����*M��Dh�~�<)6�" �V��"-ON�!�À|�<YSN�>�V��	ؐ`5>�q�kSz�<��(X�Kyl��ve�"�F�+��vx���'LD+1B���a2U��i��d%O���u�~R�"�ܞ����"O ���A[>��X`�DK�{�La��"O�A7C��}�D���D	U�� ��"Ol��� o|����B�R�|T@�"OВ���3ZJ�h���7x�x��"O&��m��c&Nb�� �"O� 8��� (j�|Ç䒽pC�d(�"O�P)�l\��J��7ߠf���8S"O�,���!���a��3 �LI�"O� ��*w`з,�Ā:�D}�
���"O����Nɼl�������E��S0"O��b OԿ4���a��܆&��9��"O��p� �w[�`��fҼS��=��"O����I��$	h%�랖D~���%"O|�X� ΰZ�� �C
jN؂7"O�9�
S=k����d*�Ch�|P�"On�y���3B�P�Hu��}(��"O~���)œx�.q[�	E�m�"OY8��	,J��PfߋX�e��"O�u��H�(��a�ܳ��("O(�!�&�6�3$�0i�؀��"O����$\���t���;�"O8�ã�+|�L�*���g�2�
�"O@a�vHc|�dC3��|�h�S "O���6![�g삡�$�&���"O���'D_� �WD0A!��z�"OD8�1�Q�!,�TB�$<�L��"O,��^�K��L8�&O�B�09"O~i0D�"�ZX�ͬ%��$�w"Oj�R�k_�
]y��X�U��0�"O��R��9x�t���mI!I���U"ONA[%iEo��t����F�0e�t"O��4��uD��	8*�Ќ+�"O8xp�G�^��uږ�\#�*�J�"O�<kQ�ǒ&����A.^����"O��@4�Z41F��p@R P ]� "O�0J�$��f*T�ϓ.Cab�S"Oz�P��� wΪ��mΝ����"O����ʰ;2�ē��I�߼�1�"O
0��D�5��������c0`��"O���g�dNԴ	0��F'D|�"O��C'��su"�B�Ȑ>E�}���D(LO�YQ#@�	R`���OL�~��pI2"O����\3$I�yXh�f"O>�86��L��xKfΔ�_Z ��"O��p��||<���9iC~�S�"O4��I��"$��l�>O*��� "O21�P(8�rt�LҰ5z�A"O��A"�Y�T��@ ��-qX@Qw"O����홻%�Α)�(�̄$#"O�	� � �BZ�g��d%
�"O�Y�
�8b`XR�o����!��"Oꉺ���BC:IN���uH��|�!�$���`u����={B�h:���!��ğ��q�.T".�=��'_vz�y��'�1O��p�� /�U�5�?pQ���"O,�**��l# �85�I�(J�k'"O�d�D�m7p�����O=D�)g"ODLi��ЗA��UJ�8_�ԡ �"O􈈆!�@�V�����y��"O�LS��J]b���f�lp��I�"O�Jq	�.i�r�`��n=�I矰�	çrwR�Z�!�i[���G"Ht�ȓ]T���\�"�T%#�E]�^h��*�~%��H1DD�q�Ӌ���ȓ?���TJ(
�.�Ag��+�ʐ�ȓI&���C+|���x�$ɉ�p��ȓC@`R��}�"�
 �̯J`��ȓIW��7�LY-��{SL�@�0��NNl�j��2G��	q!I �t��Wԍ���?ٴ4`�%��!��ȓt��k�cUv���OU0�z���}oj�"�拍��S��Lc/Ć�S�? l��5�\?�!J`HYgܽ�"O>% �b|���  IN��"O.���п7҄�SL[8 />�q&"Ox%A�#κ'e�]��N.X&�m�"O0GD�.�t}hւ,X�+�"O< �s�W)�جw��k`b��'"Ou2�o[�\�D)�gU
\U�� "O�Hx�ϋ!V�N�B2G^�{��v"O� R�c��{��P��&U4��"OƝ٠"U,I@ �PB1n+���s"O�����	/6�;�B	_"|��"O��U��,�	إ��9�T�0"O`�S �Bs8���DJA(�"O�e���B�m��|��@�y�n��w"O:�����
.����!J�ē5"O�TA���$�|�*BׄAН�"O��ub�R0�};�@C'�b��"Ov`"�,C�h���@���Je��T"O�<If���%0$X,W�`�)�"O�y{�/�Nr��A<y��t��"OTH���=�l�ʦ8���z`"O�����%�Z� >9ҒU�g"O>�Z�Ǝ�W��@���:�B�2B"O�q�5�[
~�l�o��a�i�"O�P�ii�J��-�t��I��"O2�b��]t��X���M�W"O�6�P�k���z� � h�~���"O�d(	??aDٳ�P>Y�>a��"O��X���(�lh��،s����"O&�vI`; ���"ĥy>�m�"O\����[��<��!ޮN/0��%"Ot�4�/}t�z�� W�HI�4"Ota�s@͔=R�	Ǭ˨#�$�j�"O:�q�횋P�E�ԋO�S5V���"O�t�����Q8�%`*O b���"O��kM��0���2S��0la�|��"O�9J	޷T�
���ac�i��"O
��e��G�ةq���2va\T�"O�Lx�N%t�D0#�֚"�(�"O�,�C�0����b�,I���"O<�āU�A'0�:Adçy�`��p"O2�aɂ�^��[f۷NYf�i�"OȰ��$O�<ĔAS���-��u�g"O�,�B�)�2R#�.��hiw"O�������)�7�U5-��Å\�T�IK�S�O��\@� dB��qgX@+.%`�'���`��оRi�8Х,�=�2uK�'6�=b Nؒh�E��O@��;�'C��bBN�T����\i�'����,�Z����#M��6ܢ�'5����A�.7ɰycE h�|8�'�RAGӏނ	�2�ŚtQ��Z/O@��)�)ʧ�B���ΧYT�\���]1�\��`�L�¢
*(�)��#!�\����Ar&K>C�f0Ɂ��8a��ȓ2�(9w�D3mvI�]�UxL��ȓ7��X�e�.����3O�J�d��ȓ 醨��))}�� b�#4�ȓ|d
2�ġ:L\d�t#�$t��a�����1Vz�@ �I�g;�|�� ���j����Z�.�#���)���0��I�5C�T�S���i�l���.�X@�򇉅n�N��e��%je"T��\����:�� ��"byj%��S�? �y0��]�N���Y��3jq����"O��p��p��pJTA)k@����"Oa�	[�L����t�� \949`'"O%�C21Ը�Ue�8s���"O昀� �i�`h���!H
�"O��i6!)ekL�F�Ն)��
�"O$}�512��C�X�x�"O0	g�<~n���`������'o^��Rl	�<�݈��Z�ER$�'Ђ�Z2�� %��T���U';Ҭ|�
�'�t�ä���P@^�9�
��g�2�:�'�6�P��W������oM�S���'5j\: '�6[\��q@�$��Q
�'8��*EC�#��ps�,��t�U0
�'d�esv#�R*
�1/��a����	�'� 0�	�<Q��a�0h:	{
�'Gb��U����|%i�	ۦg�e�	�'X��+X�jy)��C�k���G��`�<�q&��|�d��̄/ar��w�`�<��0��@��,EK�q��I�Y�<&B��6EtM:3��#u�X}�֭�O�<ɗ��8V��BL��}*ZQ �g�<I4˕�>�`� V�V9�eA�^�<�e-td�(�7��^R~$��+b�<!�9�J���R/k����/�u�<q�gȣg��Z��7��{�TG�<!$M� )J��7�LZ8�q�Jh�<Y��m���郞��u��m�< dY
.���՛v��"���`�<���T�k��xVd�C=h�z���[�<Q5�
6-~B�&����dB5�DP�<	�L���p���_@��r'&
u�<Y"O��'�p��ǖ@�䙥��i�<q���VQ��C!7�v�Y�UJ�<��U�j��J���b�(؋#@I�<���P]�ڔ*��ܲEQh\e�Nx��'?,�(A0�P����L�t��	�'�:(!�*1�^]���L�3 ^H*�'d��j�%�	-�d��p �~���'� ����\�ntc��_6�L�
�'�@�!�d��	�4�i'�F8.�F���'t��%�A!~�J�f*�= >��	�'{���,Y�?�P��2m����t�	���'q�}��-U�{�Z� �jQ��:	�'e<	����%>��������'���R�ѺH�r٣R���߂���'$�+���"K���pO�#un`��'��쁣��
K�2Q����!V����'p�y��B�3d�-��%�* "�xi�'�%Y'h�(@���kR����бr����F&L���qf˚M@l�b	�I�!�d�>w/.�㔦J�tD6�"�d�L�!�@e�Y���8�1��
�g�!�d�Q �%������g�&_[!�$[�9t���_8i�V	��b� 1!�qt�4:TW�U}^�
�AG,# !�<, Q%@�@l�����F�]k!�A!��	�a��wX�m$ �`!�d�SH��3�o�)BFpcc�݌Q!�d0g�QX��@�E�Y��o�?H�!�$�#"�2�ISbB�u�,8�h�%T�!�W�A/�=��مg�j��:&�!�i�jYZ�D�� ����B5�!��Օwa6��2�C�V�z䇔�5�!�� �᳗b��5ߒ0!��	�HQb�"O�-�C��;J^Y��	�6uԴ��|��'`az2݋v,�(j`L#S)p��"`��yr�Q�:���H���`�1�F���ybg�L��Q`��]��0�@�yB�."q�[��A-���k�i��y�ᗃz�%D��y��Q�:�y�ʂ8621��J�=qo�)������OT"~b2���K���"e�,v7LP8RC�K���0=�di�:Pڈ	�"פO�HX�g�G�<q���^4�� ��"���P�B�<�!I�P�8���5x����z�<����r�`�u�H�H�@Tq�<�M˕R1�9C�냒QK��v�R�<q�,:(l�h� �3��0p��IJ��?�	�'6��ɰ��B 56\�^�VA�u�ȓ��h)�EX�k���k��H:l����Q��ab&g�HR<�9@@�l{PU��z�P��J�W�8��c�<@�z���J%`������(����|���ȓA2ĉQ�>&�pR��2�:9��a̓2�B��n��^`�Y�Bl��s���G"�S

��4�֛�Nu��!0ԨC��4A��bG<k?}S��Ò;��C�Ʉ����hU�`�1�6�O��JB��<U���Zf#��)JDK E��
�FB�I�zx�} ��(5v�hn	�c�0B�ɸP�$i���@4A@�j3�\W�ȣ?q��)Zݶ5`��� xr��v&�"�ў\��	�h��@��"��e��Y��H�C�I �ιc�E�K&�� �K7 TLC�I/�␙EH 7L��U�E,N91 C�I8g�ʀ�+n8�%JᏜ�C��2A����w+��G<��iwꎲL$C�I <>�� ��ɿ]R��gE�����d*�)wHh #(��#�8}�"���4B��H !&�����4#�@'��F{���G��U�
e�DBG�������yr��L%��j�W�y�t`���ybAA�.���9C,6�x���OX7�y"�@0\$4������&FB�Q��y�&@j������JG�$B��S��yRf]�l��j��F�@# 9䎏��y�)F-(E�Wh�9d�RC˝0�y2��m`�i��s��1�@ŜpI!����Х2��P�V�����I1!�Ğ0L���A��޼>��qR��#00!��&:b�Kdș�l�8,r�&ײ*!���]U�u���� 
u2L���; q!򤟦j�F)�4k	�+c��g#I�:�!��P�pi�a!�*U^�ab�*�!�DǑP��(qb��o:������~x!�$ԭA�R�z���@1��ի�rh!�D
�\�D�!��*�Ä�
]!�d��aͨ9�����F�I�Ĥ�(p!�d�=�vթ��d' ���eD!�D��=���#���rg�}�g�!�$�'s�ࠃ-H8v�%���!�
*&�4��k��a�@�;!�$#p��0hС,w\���b�5�!�$؈��D[R)��|S��^!�D�^FҥJ�Ê*"T��.� .�!�$X�t�L���iǷR"dU��ݖ{!��DRm �h��jb�\R�� t�!�� F��eG�]��+r�P�BߺQ1�|r�)��;9C|eb����}Ė1B�N�=Pq�B䉡;L~�Kw�Ʌ$����&U�b�rC䉍>�4ɑ�b�h�A�D�h8>C�.6ta@�8W(��2.TD�JB䉳OW0a��O۩b�I��b��H}�C䉬,�%���_ݞ��Ev�C�	�
�n��%#%W��sD����B�	�>�~ɓT���,����H*B�	;��4��1QɢȰaKD�2�bC�	�@|d8b���M�dI� ��B�I���Ű��@�i�((�%!��_HC��> ��`c`�v�(|��e�?@�dC�Ɉ>2|�A���-W�8S��G,Z C�	�1W�0$퍫]]D�d�<;hC�I�_��8UK'Z9\!�w쑝Q��B䉒,M:����O�Y-D�d�B��� ɝ���E(�p�!�"O ܓ2��,Nɮ�	�f���Ca"O������6�L�#��o�ʵ�T"O�:� L�s���9Ab��v�"O`���e(Ǣ ���Y�#%���"O*�����p<x Y���!��`"O��CM�R�.mbBBW~826"O�Up�(��
1 ų�(zYj�٧"O��!��q������qQ��'"O�#��J(lb�j�)?=x@"Oj��GhO����J�wN�Y�"O�d ���+��ݪ���vM��h3"O�%hf���5�6D��M_�>���Kf"O�YKV�-4�Z|a@ύ(%���`#"O�Z�Æ5�pq �����L��y�N�&n��hs�Y�5@00���!�yR%o�U����.��h�Ȕ��yb F���P�X/Q�*�RC���yR�O�ѣߵ7m���n	�?��ȓj�l�۶�?z��}k&ÒGP��ȓ�|��$��5V�I��N�P-�܅ȓ7�*��(�i��튑˓3+¸��ȓsن8��׆G����E΃-�<5�ȓ�|�)�#�R�"!д�]�f�4��ȓ4��3�-�B�}1�ȜHVDH���t���A],�$=c�ѠS�Ņȓ#��Y���I�NRTc����fQN-�ȓ^�b�	�lQ%<�"��p��E�d�ȓE ��
��XP'V�q2� 9x5�����l_&=a�t�ӱn�0ͅȓn{����C��$C�
!���ȓ�T{�瑒2�l��.60\�ȓjt|�gP5
�����pS�p�ȓ)��P����]3�@nRY�ȓ��@���;J�0;#��/hB��ȓ4ƜeK����/�4��Ƣڭf}!�d�20:�k�F�[����E��/!�B�kq"5*����(�@yZ�KM�!򄈱�$�JP�ݯhu�al�	!�d�9mԖ;oO��eHG*	16�!���.-�m�L�$& ��)_�*�!���=,qn�����{|��G�ڟi!�$ܫ,u8�:b�Ѿ���P"�,-!�ǌ�
I�7��<|�4��Вtm!�,:�*qm٧/�|��ʞc!�ɇ;�ҕ+"� B�8Hҩ�<a!��(V�BŨS��X��C��!�� �Ũ�kɚ+b���6�Ӡ8M<MYW"O@-�Eh��GKv9�rG�2נ���"O��i�A�~H�po�����U"O�	���U�� [�+��<��#"OJ���B�x���j�
v�,a3"O�@�D@؎h��p��RchP�@�"O��w�Eb�xDk�K��;^raH�"O9�S��TՖus�HB�~'�u;s"O��kpH�(<8�ၰ�]�I!�I�&"O8-�嬅d_&I"�e��8���Q"O�,[%	� �!�V���H�x�"ON�c�	�vt�aI�0F�p�4"Or�#v�ӸVa�h��4-��P"O��ÀFO7j�qJa��C"`��6"O�\��I�5�~�� H#C�d �"OD5)�(C#a�J�Z�'��{IV1a"O(Y�Ƣ�5b"�e(� `���"OZ�SKX�Z�L�a��Wۖ"O��Վ��!.�"v��=~��Y#"O���G���X*w�3n7\��T"O��B���72h�]��)��J��k"O��ӲSt�&	��(
�cb"O �Y����L�"I�3�^�S�d�QQ"OBM�Ph���)r�ֳ%-|�P$"O���Q��r0Ec��� �|@"O��p�o�!F��Q��["d��"O��sda��%5~�`U,iV��z�"O:	�Ɗ�8�dI�#f����("O
�	���PW
�2a�2��$"OH�J��
3����hI7O����"O�m��LtP�Q�Ι�Ol,�&"O*@� *��@��y��5�"O&�#���u��Y��?�:��"OސZ�I�8=�ԐR1S�c��I�"OJ-r�䇓HV��S�(����[�"OL9�J	�<���sG�$�0x�"OV�@�d��4p�#���hն��D"OPq֬B�G
��T��I-�	Y�"OF�"� �5r�b���fܬӷ"OĴ+$F�f�*B�T�M��z�"OzyX�遛b��+u�����"O�T{�O� ����G1Wt0�"OzH(`�'xl)��_�n>��#"Od��!�3�0�� g��u*��[S"OhI"� #D�p91���h�1ZW"On���V�r�d��hȝ(�vT�"O�]�4��X�,���fٝ~�Dܘ�"O��y��ٿ#.t|ʧˊ;*T:�:"OL�C��,�LT�mְgO��"O��4d���M��,Ǻ2O\Y��"O����W ,D��
C�s���+�"O� ��,DE\d���JT����"O���dE� p ��V��3r5��'U����H�\"8�W焊G.�"�'��;զ� qu.��Z�j�6a��']�E�#�I�h�<qc�� ?\M��'�v�wr��[�a�-B��e��'�V�)�咇�L�iT8<*�Ը�'$f�A򨃤y׬EA��1-��L��'H*�k�j�2Cl8�ʐl��+����'����P N!�00�*Y�[	�'!��8��
/`��2�� :M���'匕�. ����-"R.��"O¨r�'8b@�y��Ǒ
o)�e"O�  �8���a��m�fm��&Er���"O����e�z���8>jZR"O�P��k��t��cf׉G�x��"O$ �g,E5/N���E� ax�"O�Ay"�B�gߞ�sd��RE�@A"O����J��<�h�JtC0JC�Hk "O�T�`E�S�4�b��S>H3a"O�}�� T�D��騐����M���"D��C�`2K������`���3D��ƏZ��H���G�����*3D��4AŏJ�"P�H��K
�Qx4�2D�����/�
Q������B��/D�|����P��e�Z-@g��h �/D��e.ڵh��LcF�� G�4i�f�-D�(y�OZ8<�zq�U#�$��1D���� 12�\�k�`Q(���e,D�$���8z���a�S
����(D���l�|3fK��l[�Hj��!D�����R^¶���%> �����#D���qkA�ل�C�(M1�$����7D�@�#�8q��,
7��:M�����/9D� �5���]���pǆah��9�j7D������%"�̹7�Q]xHqAIb�<�C��4KO����	ژh��嘥�IX�<�dK��d,��tǜQT�MТ�K�<��"Q�l��8fbN�{ɂ��cŖI�<Ag��������ܾ!O�aA1dC�<��fJ9����*��I� !@�A�<���3�xx���]��]� ��t�<��KM�=n	(��X4�셁D��m�<���A?p���8�������`�FA�<��)N�V�nY( ��;H�`Q	�A|�<��סFDv��@!�Y�||q�)t�<���#$WH�PԎZ7w"�9�t��m�<�1d��[z��33��3 ��1��Z_�<i"�Ȗx�bݢ�hX�'>� ��^�<	4N�n.���[�0�3��Z�<y�[58�p0��_�:��SG�Z�<釉*k��ɓH��8\AYcG�X�<1�@~,ze{�Q�Dw �j5�X�<���ԪNS�0� ��&,��i*p�RQ�<���9Ąl��`	";2���b�<���-�*ɂ��8�(��Da�<���V:v�N"���\���`�r�<Q��U�=@!�R/�G1T<��cIo�<�SfX1_�t��$�!��aE-Hl�<yA��2"�h]�Sh���ܙз�A�<A($E�JT�6���9>�Ҩ�t�<9�!�0Ĭ���}%�蔌Ae�<p$�(taPo�WR�YHԯ�c�<q�j��?]d�!@��8�#��Ut�<QuCM/xn�:����B׸ZrBنȓ4A�¯T�$E��Gɝ���ц�=�����m����F�%*��݇�i��A��HE����b�j}��S�������HT�֖�<�ȓ�X}ÄK�.��V�ۑ ����ȓa�B���i	�z��ro��\&���ȓ��\@�ΐK��岷�P����ȓ@�~-��%P��Ja�R%�"���J+ � �\�6��cI 3x ń�L����L�#�&� ֹb�&�ȓm���Q(�7y��<�Ңa!2kKG�<!���ް���ܸa�rQ
��<� L�3��\�N�6�0���
@�*���"O�\	��T!'wv=�6�S�-甬��"O���T<B���$I;ֲ��"O�qQ����.�4 �Ï�K�=C"O��S a]�`}�QJ������"O�}�qg��H��t�#m^5k�F�Q"Oh�86C+%B��*BϳYE<0��"O`hHa�F+M��G��� >rX"O��y�,rI�.�'6,�B�"OPu��G&��{�C����"O�8R��< ���C /��&�T�`""O��JtL�QJ���sC�i�B��"O���F!DV��1)�!A3i��
�"O\�`5䔉S��d�b��A�t�Z"O`D�s�  �<�#Qg*��"O�}���C�OϞ���AF
\T�aP�"O�:iƲi��˳.[�L��\Z�"O,����
U_�di D,�άZ0"O41{7��=h��\�v��+M�����"O����'ބX*:l�R@7nLMB�"O���P�#"�pCD.O�@�az�"Ok�*�T ���,�(`� �"O�0S�쀑*���l�)!��3F"O@}:�����(�j�"�X��"OZ�{n
'?�D��3�:���z"On��T�X�M��<�2�H*�ZA� "O\T(&��OA��îP�sr��8""O��	P�Ln"J\���> ~�L�!"O��j�WfT4 �/�Cw���"O��	h�d�d��\q@��"Ov�{�l��б��o´e"O���)X�G,d��&�ΟCC�i	�"O� :RO�@_,q�Ǌ)d#*�Ї"Ojh��Ę��M�G�;��ӕ"O��r��l6��@O,�� �"O
LP��e�<D@��O�I:6�"O45Ѕ,g�	�1@\! ��� "O�@yU&
=�H�6	C%-�ŉ�"O�P�M�8 (�k��L�G����yB 	�{��k&n�>i�ⳇ���yL:Q�V�X�M)`�@����8�y��\+%�\���]A�q9Gj΍�y�/���>4`#.�V�����n�'�y�aĘx�����B�K^b}���y�MG<l��ٺ����7 ���ì�yB.S�"`~m�2�A�'^h(B��y�c�Jp �V�ܣ@�)�w`Q�y�˓X�|�`*i囶D\�y2+����`kC�HfB(�	?�y�cͷSF���$B�\�������y"hZs��86G�4Qh�$(6��y���2%1ܵYV��Q��p���y�D�PY��1q�F:r0���ǋ ��yr��pv�`�G�ΘcH�j���y�n�+����_�	�V�CF�Ȱ�y��4y\!��/�t 􀸶�ِ�y��V!+,���M(�j�UHO��yR�2�ޙ����M��0(O��yr�ɥn0�2 �ģ%6 �CJ�y�I��P�yO��V�@�P��y�ؖ6�je����V�V�IQ��?�yr�S%{�x���Fz̈��C��8�y"F'F<�d��	ۛx��+�Ɛ��yBoW��ָj ��s��Њ��[��y
� �9A���lm(�"R�75�V"O���b�
\�e!���/2���"O P�2��3������y0 ��D"O�J��U>/N���2,T��c"OB0"|P�8�I�$�����"O.�#%L9y쑢�a�x�� p�"O"u�"	�W��qb�5f���""O �Y)P</�\���}`U�B"OT�p$Ӯ$T���Hp]�I�7"OB�2U(�/3	t�1g(��L�j"OĄp�GN%���7�˟i�(�"O�dQ�\�D�P$8���&DX�0"ON`���ȈR�l%���q��� "Oੁ���%'���jg-��z~�s"O�{Ť�.+bR���KN	�\�
�"O���`�ܠ���{Ɗ��z�|�;g"O��C��;a���ĩT��8�"O��ZNV�IE�u�%�{{4�@"O����!��K���7@Y�0��"Ot��gM���9cK�J����"Or�#��V$��8;q�V�}��0�"O��&�Ӫ}5��@C����"O�qɢ+��f��t��*x�Q�"O:ɚ��W*o&�!8!�Nr^� "O&��1���&�����4�>��"Ot�A���BA"�3�6A�P�"O�嫓A�[�������s�T�a!"O�$v`P�Fm�`.������"ONi��j˧y�Vŉ0(�Q��p�"OҔ�1?hd��'H�&v�>��"Oր�F��Z�z�S�蝰0���C�"O�)���eu��*��|�bT"O^��1�[>Z�X���*P���Ec`"O�`���JL�� 8n��L a"O�<�F���F���j�3�(�!"O���AG^�Wc�ˡIǊ6�h	�2"O&AP��
.mP�9 k^�t�5��"O�%�����[;~490����z-�g"O��cqA�p$�8'`�=,����P"O��`�T�=~~�#�nWC�DP�"Ox"�Ƴ&�RkI� ��U�7"O|H��	�	:�t�8SJ<~|yb�"O�p��4,Y(,@�	���is�"O^��6�I-�b��k�}��	� "ObyQ-S2�$M�$
S,���0"OD����u�Р 	� Y����"O�@Q�NݮQ�ҡ��D�B��<�"O$��ڸ|}�Y	Ą�	c�p
�"Ovc�Z�l~�	w�E�Z��"O��fa׺n\��P� 
4O�a��"Ob!K�����\4�y$y��"O>��W�(6P-0�ȊA#x�f"O��z5O��[�����Q�D+S"O��b��w�y1�/� �@���"OH� э~��Y�Go�?^@���"O�!Aō�O↼��]�r��"O"{��&�`���];(7�՘�"O�A�@��s�j� �_A�yj�"O���򥗦#��Q�DH�[2�]+�"OΨ`A��!%��1BÒ�*x��5"O�!���#J�	�C�
����"OV)FL�0��8CU���V^�:�"O8�Yp-߰� ���r��P�"O�-�T�:���m��b����5"O� �HqQ(�9k0�qZ��	:�i�"O0���MW�t>�JCM�c��MXV"O�T�b��(7>�k1�,	�h���"Oҵ��ӅFO�(
�㕋\�} "OjD�r���h7��եL�"�@u�a"O"i�'(�6ڪ��n[3qў���"OV}sv��;Nn�ڱ��:�0�{ "O�,�iب%\�x �g�?,���"OD��iG�$`kw��W�PH�E"O�9�B�^�&!A�A�n�Ka"O�� �@C�$���o�RO��"O�i����0Ce����hs�h�+2"O2��(R�~�Aᐭ�7ۜ`h�"O�A�� �Q��{b���(��"OT:�ё'���b�k�;y�0��"OP	D�Gˎ�h7J��pLu��"Oz��fI�B�L����Q �}��"O�I���c�� �bIV�:�Y�"O>\[Q��`�~1�*G�V��tڤ"O���҉DN��3�*K`aZ	��"O4ub��ǡH&�E�C�ܿ(�
y�"O.��5/ ,:��S�³T�|�zU"O�ɲ �T�]��K3Q��"O,� ���BG�:UdM��㛝M�!��Q�e�)��2<r����!����,bqgI�V"�9�UA@�)�!�@�z�����."�<�QV�\�fF!�"sr0	WE�e��A���&,!򤜎T�,$k��#LlZM�$D�h!�DTi�ɻҨ-u0t@�c	�o!�d���F%�G�!~�(p-�u�!�:��I㋚�$��ݘ
�!��A6x4,�td��tm����2U�!�DK(\1���1�����	J�!�ė*U 	��ᕗ^Ķ8���e�!�D�&�2- '�C�0f%��i��=�!�$��UL!Pc�{�|��)���PyR(�2hX�Ls���oVZt[b��y�K�-Ҥ8���� ^����� ��yҌ�/KW��Ӂ�#Y1Q�R���yBۭ�jԙ1#���^yyb����y�o�(x�F�TjW0��bsB�y	�=P���&��7b�R�U>�y�BϏ3�>Գ��.�@�����3�y��G�^�����J�z1�ᐅ�y�N0
0ir�Q�t�0�
�����y¥A-G_�e�Ǔ�@jU"����yR���Mn]�蕊����m�y�	�n�nDj��T�xϪt�&����y�D,K n0��_��iㅅ���C�ɳ;6+o]J"����=М��'����,��;Q(pk0���a<�-��'~�y���[= ( R�l�V9�
�'V�=J�a���5c�
QǬ8��'��i���0�����J�n{�'�:��@4I�5�ț1�3
�'�̜ia ʔa�j�3%A>�L83	�'�� �/3����`K?Nꈫ�'�j�b�ǚ�a"� ���=X���
�'X��j�>��P)�$��|h����'� �çh(}�|���ʿ��9�'��X�Gc�"<� �@Ջ,%@��6�\,0��
v{R�{WFMx�t���A�S.Ze������
9Tԅ�S�? ��� P03�V�Y�ʥ~ȢD"O�]Y�>Cf�="ֆ�,��9q"O�U�d�'4Z����W��aI�"O~�fiH�A�����?4V$�aG"O|qiT��~l�Y�D��)@v�&"O�(�F�2*��lY���
GL
��*O�Е��h�\�2!�����
�' t�Ϙ�Bb�R�G���{�'�F5���TG+���Wn�D��EH�'@h�ȝ2�}�PKM�oԎu��'�㍐�j���V���a�L@�'t��S���0�^/X�ੇ�=�z܉A��_�� 9�)̓\8���ȓe�ĳ��ݑl�<J7�&k}� ��H��} Ǭ�?+�.4HS��1$���JO�(ɥE�a���a! �B�)��{�kƎ��@��F(��v� �ȓ:7I�D)?Ρ�lV�3���N���9�+� +�6\ G�
ݜ���7}���O	�AA,�Ud!��@$��H��|�ׯ�*���`�ް�B�É�h-@�={��ȓz�� ��2N��ȓ4�K�7,�i�ȓ'>�X��&�.��P�7�(I�ȓ/�,�:6ףg���#w,ӈD��H��#;�8�V�ɲA�sá�WFE�ȓ$���FB��>~l�ȓ%�RE�wk��t����@&ي4 F�ȓ#\ �#/T�� ��ʚ�=�޸��M��Sv�- #���Eك&�0��ȓ2�b����]�Hf@�k�ޣ:'t-��TT��2���@�"mN�ϪلȓdN��'e�6)D��B`��n�<�ȓV�Py2�@%њ��Z�&X�ȓV���H䀅'��⡦Bv�&��ȓ@&��e�
�E��D�ԅ�i�b̈́ȓ���[��U�vפy+D��a��M��wܱ����	x�����	�lhD-�ȓ6��zRh�i&P�
)���ȓ����ȉ�>�d�'AZ�!��l�ȓq������7�PAx�aF �q�ȓo���qM�4i`�mȥU�VT�ȓs�FH�ŬC�[��҃�|�p��PU�U����%�ԉ�K�(�ȓ{EN��Bo�%����b�ԅ<�@�ȓ?��p��/�aB
09!� �:����z^e���pNl�(G�P�V��ȓq�0 #Տע4�����]�@���$����
�$�3�mQ�6�����7,.�P gC�:� � �f	�Wo���:Z�x;�� "
�@1@��ދJ��I��t��a%�{�8 `�/e���ȓK��1����>�\ccL�S����,�Ry����9j\�����[X�L��x����#��<1ؔ�#B�ftZy��g6��glD�&�����iiL��ȓL��-��I$;�2��ӧ�1H�8<�ȓ8��,�&m]9Y��{7鋖Tr�<�ȓ�|#��=R~�!��̝'��)��&x��&kϛ�n	i���7��ņ�jb(W�q��_`���ȓD�\�����	KO��	�J��XXY�ȓ|A�X�&
(	r�
DK�+TH��g���c��d���"�)NC�)� H�Cdin���ʇ@ƚa"���"OxM�E&Z���ŠL y�]�"O�|�7��.z�`�`�C���"O�4� \�s��Rn���"O�M���źdp*����>/YĒ"O(L@�o%r*TYc��.K��j"O���w)w� �	��ݕvWʬS�"O��	��6z�Ljn,(3Rp��"O��4�_0}yJ�X�M�]�"Op��ԨV�7�6 ��
���K�"Oxx���ʤ��"C�<d��d�v"O�XS� /;r��t�RHan�b�"O��0�zD@����8b�����"Oha�7ʀr��Q��c�5�Ї"O��3p)�	>��V��	v6�2A"O�y豍ƓEk"���HT�kKr<k"O
��玨~Z2&� K,�%�"O:\ZB��	={$��"&�D� "O̫�Gk1P���n�"1l��'"Ov� Í�}2���  y�^��"O
E�I\�p�|�R�"�2p��"O�0�@D���u�P�z|B�"Od�����#���`�\�
���1"O������%ML���-�f�D�0"O�����\�f`C�e
�Ph}3v"O��a�!�5[�$5�%���d�K"O���E�B�\8:�8�ҮO�!��� �zQT�V�mN�ř��%$�!��6i�5`%ɔ*Lڑ�"��M!�dC-!6h`�2�*���nĊP�!�$Y�5�x���VϜ|㴇��^$!���(<"���`�8
�E��G�T!�H*o�j� Ì^�;��<��Ǖ�b!�7O�h��bV��zi�A�p"!�D��]�p!�H����$�s!�d�#=��;EF��U�8�p��K8	!��?%J�ɷ&��tg���虄n�!򤁯7-��!c�X���>�!�D�hC��#���4 �y/Z�(�!�$�	��k���s�t�I�!򄍧.0�Ei�A�cj�� ��^�!�$�2]��C�MV2HR��s�σ1�!�� �aN"��$GW?�퓐CE��!�dI�H��!��ܣqB�I�#�g�!򤅧\��тӮ0W��%¡��+8�!�dMH&�2'�
�Z2U� L�n~!��֋	xt�b�C�ww��(p�$2w!�dC����PWIi�X� �H�,w!�$I�"�z�x�	 R�X-�al!���Ȥl��#����'[H!�䝬=��q�m72�P�0�O��x-!�$��j3���B�� B��j�<��N��k�ŉ�f�:��.���ȓu�������r1��+~�*�ȓ%[.C��(�D�"� *-�`���th8�J�˘�f:�*��@?9C���A��=+�F�9ڎ���7T�B5��@�R�����Vd$�+pV����dUf0���9�0L����N�ܥ��-�d�t�ӇWv��ۤ@X��2-�� �@@�gI�L�J�I*�LV��ȓ ~J��R7U^�9䞼����a�L1�`�-���r�ݠe�\��
��j �øG���j�"^��Ȇ�S�? �=���� w��\��:��(�"Ol� ��;gj��#Oэ�&�P�"O�"UA���r�C��|���"OPD���� 6)2���U�4�A2�"OD��@/]"<�"��6�ˏ1 �ʴ"OH�yA�L�$��f#��B2 !�"Ol96(}�2���#M�� 
�"OZqɠeF�9��[�,ܪ#�jK�"O��d����h7&^9!U�
�"O��"���ifB������K`�rS"O2�$K^'1����}B^��"O���G&@=����±)b !�"Oz�
r��x<��q��f	l`��"O�bk@�^�na����,*��9�#"O��ؑ��d)�B����t��f"Of��5�Y��`���#*yXa���?D�h�@A�$*�h�3i�.-� K*D�\���5�p'ҝ)�6��'�&D��R��EN=���c�ì�(��!D� �Ѕ�g���BGhB5����!�>D��:gA�OLT�DdV�U���
P�;D� ��	�&gP�C�O<B�\M���9D��Z�/�ѸT;� �<�~�h@�8D�:��ߣP�^�q"��*v�p��G<D� ��IC�s��$("����<���$D��+�AE� t��(ǥh��z�f8D��s���S���s�:Fx�p�#<D����L�S5AH�o��&����9D�<2'$�D��D�����b%D��i2�H^%���G� �ɤ���7D�H3R����V ��L� px]�0�4D�ء�ر�6m�#I�>f9�w�0D�P��G k 0�	F������;D�����y]�ah�1V���$.D���Ȃ�Nd:|��aA>�d[!� D���C�� k�@q�dA�ckhQ$T��r@�Ymmh�9�-Q��8�a�"O�]��m�C�*�@&�E<�0���"O�<�o�&L�B�KS%˹8c,��'�(]"�b�-V��a#�P'iL �����!����-�4>htER�H !�!�D�3/�DC��|G0A26#�1�!��V�^&Д[�͟mMLu �i�){!�G�����z$vx�&�H�!�1 ɡbә�4��!�DK0~9N��A�ث6-��A����!�D��
,+wl�,SPa����9�!���k�"urF�	�L	�d��6*!��XlN�SQ!c�h(i��W!��6庵�d!F�p�^�z��Y,d�!�dS
��[rW<���H�H�+�!�䚥N�z�'$?G|$�A�Q�!�D�?C��C�,Ɲ!�����a��!�d�-#:����-(ʮd��C�:+�!��$An�ȃ [1{�����Q/Za!��W�/B00n m����!nİv�!����=D*�"��7(�����!���z��9yu���������5�!�$FzN�M2q�I.W4%y�ϑ�
L!�ė-'�.)����AD!��	�'�����ԬM"�p�"a��R �3�'�����"v��e�"k�U5����'pԁG:=���AG�ZM$�ϓ<��ag�V��D&y���$	�e'��Q
�qs!�d�?0�����=s�ء�j_�1��'x�\���?	`��� ¤��.�b��tp�f�{�2�Yr"Oڸ�j�((4�
��t��SPbͺ)�B�,�(�9�`$�3��ۗ{2QU�?MH��A��T�E�!���y��2�PR�x�yeÉ�A|Z�:˚� �5�XX��(")�4�HX��G!F��ط�(�l�ttᥓ�A]�)��jb7Ÿ;��@�0�2. }x�!p�<9Dh4`h`����`�sy�ᙇwPh�#'���i\
���(���sM�x��9�!��8yg�`X�kA801�EC��(u� ���
���3#޵Wq
�:�Y>�<�Q���ű@��+��Lkc�UHX����F�0F�ɓ	�6�]%
֣�x�Z�I[���0[@y9E�Vc8�:F��� �n{��!��Q�$�q`P�3|4��Q`D*it�=�Q ����ƅ�m�}��K�+�aҴ�y�X��z5:Ƨ�
���!3���I�"`{T�	1	Q=Lxu r�l��ygA�h�(y��צ�~Ma�.�yb�Fo���*�e�}����BX+�|���kX*AP��W��2$��Z��o���Fy�D_P��\k K�pǾM9ҀS���=GL�'.�7$��U�:A����v2Z��Р�bt���]ݮMr ��a8�	�g��ed���tn�uK�����;�I�Rq�U{�F�����3	�j��0;5G�?�°"�m�:I��ƑP�qҮ<D�4J ��p���I�MK!>�ٳAi\����bg�C֪(��iѾ��-j ������@ߙHY䵰"�=4$Q�4�w�<!�.Ҫ�q�#j׉(���g�֮$�6����P>�h�����-{�r�"�Nҫ|��<YքR-xh y&��z�Z�*���i��L�QC�������M�P|+��c@��'�Q�]�p���4U�"\s���:�p>��	7�8�RM��-:2�ã�b�ũaϐ�H��6	U�o�"X�a��I�qQV0I���6y�W���!�$�1\���C�e�,�p�E�H��<�%�^�SU|��2�M�qU�U��0��O�*��;�Z�����8����ɞ:
8D�ȓ|���Y��Cf�\�RaB:q�,1�7)I��* �)�.0�K��ӡ|���aP�"ʓj� qK��ͥYIH�yb��9b+�!���j�|��.��c���JTMA0m~�����<C�(h��
f� �vN�-ւ!��"\X���6nA:�I����	�=�h��K�<�r�F�v�m3� N���謟FAY�R$���@g�6#���D"Opzt�})�!�0+O8�a��v�|  �'��)��D�0@�P�J'§�V��MXa�c�#d�n�(p���6L^C��-�h=�#$��$�nM��4��l�R��=E�s�5-�֘`n�ٺ���N�.:V����#'	P��ӟ��{� ��wj2�9�M�,9��D.� !=�A��@��.A��c��,A�	
�� l ���(��Aѩǒ8Kh	Ex2�-#�hɑ"����Xgh�����ah��oOЄ�B"OH��&j�>���Q��V�{OF�T��)m�2��͍���S��?tR�5�Y[G�\�VM���Kv�<�R��98�N� �EXr��f�p�<9�*ÈJ��X��A��\1AM�q�<3�ސ[�����QQ�t�E�n�<��k=\��)�i�?�`��RC�o�<IM]���yqh���e�A%�d�<��+7~��W&�*8���Dz�<y�	;m��*%a��e�E��`�v�<i����j��+V�!xvB�P��]l�<��Y$n�: a2M�"X��U�� �D�<1ǌ�'ǘ��T	�=��9�	_A�<A�L��:�F�R��W��ܼ�F�B�<S�ױt!��0r ��4�L��M�{�<�Ģ��d�!�Αei>�C7/JL�<�CG�*F1��޽r�4"� O�<q���6eFua����%˕@�l�<��\5?���WI���T[���T�<9�+��d�0�`ې'��H����<9@�ǈg�(�b�ě�88E  ��m�<ѵ$��t�)�:F��DX#��j�<	3���Nu���7�B0MZ ��De�<	�f��$���� �,.�n��i�D�<� �LsE��L����_$~E�T�"O�(Bp�ߡ}��;uF�"x>��HT"O�,)����r�`[�f;7��@��"OS�%�7임 �ޯ*����"O�ڲ�!H�<٧ٕ(�� !�"O.�f�A`�
A��#�R��Pq"Ol�b��9:�c����SV��"OB���N�3�hX�!\�.F����"O�Yє�P�_r�Y:�[�i� �"O�EZeH�3~� U²�4@G��92"O�@��·W���B��A����"Op�ۢ͑(`�,U��ѓ\���"O4|�r��$?,�1׫�3d����"Od�I2j��c�RA�F�D���U�G"OT$��
k皔 @�PZ�0Y��"OLU��ɉ1�$�YBW.(`ڒ"O2�[G�܁`�H�(�s���e"Onњ���b�CF�ߠ��D�U"O�U�����ؚE�<1����"O�$3�ț����yb�5�mk@"O�P�ԯ�'���!�G��d4�@� "O2,���8�}k�� �"��"O�Rab�,C"���1�
��F"OX��Ī$:>D��d�=gPI��"O|l�w���Lu�����ˉqH��;�"O���M�:5�Z�{� Y8O�ܰR"O������>Yu����τ�s4d��"O��yc�A�[(1*M��f?��T"OԠ��9K����퐮z� "O�<��"]3\�j�P5LK.�IY�"ORLr�Z��Y��k�#1^`���"Oh���"3hȹ�)!p>zź "O,Mkp��.%�V��F9Ctp��"OJ�R� �v�����G�ok��3"Oƅ�.7DQ���Z=�0xg"O ����?10�V�J�L"�["O�t ���[�$���&חV���"O�TYюW2*h6YJL[��"O~���Ht����#*�=	�:��F��'w٪�ڍ�	�Kd�)c	;D��1�HٲJ!�d�=j�����˵ l*p��ԁ24@ѻ��I?��gl�|�'�$!Ă�V�`˅EA]3���'@tB�eV�X_��4�I:W���b2j�E\n5��刡LA����	�`���!�9yYDT�%�խZ���d�*r񺜀D� *Y��ۖ L�.�![��P�4���0�l��*���!��ېI$
���F��f�'�$�G��	<"ђG��3t4�F��)Pu��h�+��nO<�Ò��1�yBh�X�vq�F*��t��1�&�U�x��8�厗�n�t�CG���i6P����L>��n�Mc��i�%�v5D"�(<i��n�|P��B�p�9g���Sa���&��pҘ�`T·�q%���G1�������!,�!��Φ/�axR�ߦ<� �(�mX�z~$])��a� �`�T��h���� �̵!�Orh6Ι	\͜-JT眄wU¬�Ɲ�<C�N8澨9��H��!���s���xAAaKG�]0��IH�~x`݆ȓu�HCu@Ŋ-�b�&�Qq�A:7K�7R@�ಯ֟[k��(�G�f�'��.Gf���EW$B\F5y���KV��.Dn���*݌?�n1�`�S�6���X�����C� =(5QC	��<���(D�`��ƥC�u`tp�Bs�$�F�6*��kC#��w*��ʳ'��w�u�%�]�
�ڡ��-��\�Ɠi�0�#f�\��%���R4cS���'���cDMZ�m;D!�m^]dΜ ���L�`��� ������	4�!�$�T���x��`�
t��(q�dG�Q��!��0LƠXLC1�ĒO�`��iP�l(��u�$=�0
O4]�$"��v��9�J'�%��^�8
�c�N���0=� �PB0��=`��ls ��6��@���'���
�A9��T�sF-����4�Aa!�;{V\[�H�I�<��g��&�h�Rp�7
-$��M�ɃoR\v%[�}����$^m�Ojd�d攈c���6L:f�����'�(9�Ĩ	��`��Mv�6*ҒEJ�b������ � ���ē� ��슰(�@�"^sBh�Ɠ�*y��	��.u���ՐEi�y���R�yԒ0
щ��
�Z��䒠pL��/�I%z3v�zr�z�#�	�Y����<�g+R�X��<AR� ~HiR!��Z�<� 
:>��T ���,��g@J��@�c!�v��d�!(�B\8��^�y��.�>�I�)Cy�~5`��ѻ_y���ȓw�@��"{���×0*k\ ��_��c�"�$h�"��%l��<�ȓR5B�+�)n�+-"n�`�Q�"O��rA�I&��óLs˜u:&"O�ѡ��՗r�`Q豮[�w����"O����D�?C�Z�;6�]<��m�T"O(��q�Uk8�R%�
2����"O�)�'f��lF��&*B�*�,1�d"O2p� �(�X��P���w�1�P"O��%�47�`1C�,B
M
2,��"O�tt�2T����A��q�	
v"O �Y&k�<������&h�Q"O�)3a�)Q6`	aC/�zeb=��"O4%����302�{�,�#zEΉ�q"OdS�l�s$r)c녂G���kG"O�p�����*zpu�j�8st��[ "O�}Y7Q��R��d�Ot֥�W"O�̓���o0~e�`�!P�D���"Or�C�ʁ)M��l�� ��p�Cp"O�q1�
�z᎜c�H� dy�xr"O��8hB�о����/fb��"O�a��SC�F�pǫۏXfN<��"Oΰ��a�;%���bQD���� ��"O����C�h�:T+vĞ�[�z%�V"O��r�N�0��X�	Q�a��8�F"O,��r`�#k����ȗ~���f"O�u�VC�;pF���7a^}��"O 9���t�Q��V	)g�ċ�"O2|�2%�Z�8k�)��at����"O�EPT�D�MZ�И�'6P�{�"O*�s#�V�O�u��ѯd����"O�,Z�M�:\�,p�Z8iT^Lq "Oԉ�c�����r�.��N_Z4��"OvuZq� wƴ�'��%ʐF"O��!ਛ/n6\X��ſP �q�"O�]�Q �4	N�� �M�[���4"O|�
GEU�lf�8�ϳy |T"O���I�W���J�&ů\QFy
A"Oh���zҥ�g�[=*�b�"OP)CD�B�iu�\�a/y*�$��"O�cg���>���J�oT
P��"O���P�Φ0��уM�7
�4��"O JN҉�6�Q��D��.�"O^�8�V�Z( @8t��ag���g"Of�7`�*�`�)���W���4*O6����ܱv���
�V�s��1�'e���C�	���cϝ	�f�S�'E��1A`ʐy;Z��1fye����'�Lِ�cwJ��PPѱ$���z�'�81j��p��m G�A;���'��cƊ	#JR�0:'@";�$�H�'|~�DI*%R2��fG?�h4I	��� R�Jt*R�|.DT0&�,)c!y7"O�)�k��v=5��C�?ri�t��'<=��׿��	%I�.IC1�O	6xձ��� C�I=7 ��R_"�8M42[�O@�ib��jg�t��Ef*�0�g��p�y�o��g?�B䉺�Tͩ�)�?H<|9� iU�(}��Cq.U\~�a�+W�T�}&��W(��'���"�1g�h`��+����Ø+}N�H4�>H�Z��a&y�h����GE���K��Eʂ]$t�վ��b�&�w�@Ah"�Ō��]�J�q
g��V���o�J�E���W�<Av��8sD�!�w��*��d�Jgy����dL���"�>,�����	�;|:%q�Ƃ+H4�`�C�f�!�����[d���o=�с��D�I�t=apAڸD��p����{�Z��]>�<aa-��u��Y��)V�8;�Xh�KsX�H��D�5d(�y���G@�F!�g̍.k��s#,-X�`xxU�|��`��	� F���+�e���p�.֊YJ�<١%T�&J�ۥ�c���(T�����O��	�@�&�����6VX���'���w��9\���-�8ĩ(��x�ց[���1%vd�q�I��E��w�rd[G�hW����Z[(�B�'��lĄP��* ��/��u�h�BI��A �#I��R˟4���o�'�Fi��#Z@���j\�t_TX��n��Y
W%D�n�PE�+�!l����@a��q��i��d��%j��^�I���P����&�]�Ipu�fb�f���D�l3�v�c���8^�:܂��51�l�SSY�@�C�^�(�V�%\}�PC�I$	��`��b�K�耺t�F !<U�`om�"A�F&S{^a¢���.Y���4�sޅb0�U�Z�b����u�j�#'=D��hB�+�G�4���$LV�a[^�8ⴍ�t#�/�J�z�cF&G���0��J8 �Kt�X%�@����5���d�9,Wfܢ���6 H6��t���c��y��̒�{�Թ�L7nH��Cv��5Y�$!��I"c�(��F�Q��q�%W�DB㞰����'�-���j?L�j�L�)���0�O*��R�Y�8Ć��k�?T��yC�'�8�"4��mA�XId�<P�zlƩҪDL ��$�B��kE���a�0��~��x���T��sƞ��vg��F�D�b �,D���-̸v�]����(0��A%i�t���;'�i��\Ӳ��Q�����9r�Q���'�~<�
f�XC��b�7\O�	A�%r�����D�thVH� g�iؤ�8��^)d�,�AFĦy��-�K8���q�_�jQr!���U�Sjmke�#�	(����`�f��}�����dȨ�k�t�]�E����ȋ���@a�
�yҬǙZ��BF��Fw.`['*5p�t���.��`͸5P'��v�:M;���k���-�!��
$qiJ��nD�M�!��G�E-D��3�%Ji�A#A+E�3�v�S���<�@L����5�Z����D|�EA�JZ�#%AC�Q���rPEX���=	U͟/S�����AKx�Y�͔.J�x�t���WZ���	�N��	a@v@;��Qfѣ�I�+id�#<i�;.ƈ��F�Sy�O��Q��{�>4��f�!FX�];�'��!q҄٩dH"���Y'7�F��qO]&O��Z�Rz�)�矼
��%�����_�q��\��$D��+��<,��9GK�h�
ݛQ�"D�P!���s�v��@�eF�89�� D����&Ǽ_v@��n"tMR)� ?D�\#�FݏB,�u�p�q$}�cd?D���E��:�\-�fC�S���ڷI1D�xB�ٰJ�=�[��40��L�!�$�PMz�Q�Lϔg�MjA����!�dJ�Oc�)(e�ǝ	�����x�!�dӪ}G
8�D�=*Y>ݐ���*De!򄏛[ǆ�p����x@���&�#?a!�$2�	����7DT��(�84U!򄜫YP�@! 6�������:G!�ĝ3��Q�m��<����-�I!�$<vpƱ�5J�7)R}�흽P�!�YGB�뵁9?�@�\%�!�H�Bx�A��� f���oB��!�^X�u
�@�N�>՛�?V�!�� H�8#�Ϩ.�������H��"O<�YS���@6`�2��<���"OHU�A��_`��,*	�}S!"O��#L*RL����!��n���[u"O�YA.��U���ˁ,전�"Ovyc��ppSS�I49��"O�x�/�t:�h��%/�Y��"O�AbU��eD��
Ts��,e"O�)�V��/)�(b�j�3��J'"O�aCP�2�2H1		��!S"O��0�ǻ�P(r�h3�a�R"O�3 (D�/,
9�ѧ�M��@JB"Ore���L�D0 -8�������"O0DR�����|�*�G��w����"O�����$��xYW&A�T����"O&)�e��x���%�����"O���ូ�Q�O��g�d�q"O�<�P.�DX��J!a����"O4��B��}*8y-ȈD�����"O��FYp���B�M�)
@}Y�"O�i3��$+,PP�6&�p�\}��"O�u�b�ށBl��)��J�
��!�"Oz(c�_�}P�Z�gU�_StJ�"OĘ8@��T$��D��@���*W"O>�s�cI�1R��PD�rQ�X�"O��P*8&�,��Gʞ		@�qA4"O����ZTX��2G*���"O�T8ң��/�QF���]�D"O�,)��		~Z�$SV�F��rA��"Oĉ�J��^��c��X�A�p�&"OR��R�!Z���Ыk� �I�"O��"�ŽT�^�:dM�/r�6(ʒ"O�	bu�R��J�.N_UR�h5"O���Vc#����l��s312"O\m#�L�6m|<(ؔs#f r��>D���,�w�	j�&Gu� ��"�:D�X �/���Ƭ8��?
y��ɶ�?D�8� ��#~[1�2>K���(D�䛃�[�^(��y�R�F�����) D�9d*��/,���BM/~HD��s�;D� �a�Z�H��5���)L�f�2�9D�xa`��b��[@\5B|<i��:D��ۖ�nz�8	d�� i.H؋b?D��I�eĜi� [��W!FdLB�N/D��b�ؽL�V��'l�lE*D����.F��Za!�d��F�z��&D�hI� I�6�J�k�*L�
�����$D�x�����T���3rf̂,D��3EߏN����K�B���� D�$�A��2-��zW���8��<D�xs1 鶴�5&ݝD�
����6D�4ĂT�-�-�]��0��8B�	�z��L�k:@�J e۶)FB�I���p�W�eB� x�W�$:B�s��$q&���8�p@��9SB�	�H�vE�C �Q`�����Q&C�I�� I�bذ�d�b`f��C�	1ne�zs�é�����`�=�B�I�q�D�1l�96eHAk��A�O܀C䉩��L3S͜L�N5�C��m�~C��f��LD��~���&�6QMjC�zZT
�3M%���o��bgvC䉟s��3�-^3k�U�@�	/~W�C�/?L�H�c:&�X�с�8�<C�)� ���T´C�uC�m̊��l�C"Op��3�;v�;Cl�{��љ�"O��Bu�ҏ_o� �,�p���S�"O�]��MތH/tS�!n�x"O�����,
�Y;7l�a/�ę1"O��hW��(F��Cu���[!"O\���C.v�I�'*<���"O��#�P����"�$6.�2�"OI'$D�z�x�x5!D�h����"O8k�@<DZ�$����<k�"Oz�J��;|C��r��{G�!"O~)	��F9k��|���SJՋ�"O<)��G���6a����aZJ	Y�"O��B2�;1�A�a��"���
�"O��{`@�)�\��/iwԜ��"OVؚ�+�b# %P� ���2"O :D�4K�tض���9kBi��"O��jo�������4m\2�ڇ"O,ܰ`Ʌ��89�����9ؔ�"O!���?^�ҁr�(�Z��<3"O`@�C��6}�l��B"5���@"OF���2 ���K"�A�!���j�"O��ѱ*�+g(8��oB��� �P"O�}��͈���bcy�"O�0ʷ�3�:�b,	#(_\�HA"O@-y!O	a�)4="D�[�"O4X���}�RHt��'�]ʢ"O������Lɘ��ۋ�I��"O��Y�A�|�*�8D�� #��Mb�"O�\:U��+��m��'�(�� 4"O�]����`�ҥt�ɉ�X��4"O^�Kd`�,��m!0e�F�V���"O��"񥆉|��,P��FPt�xA"O��' �:�Zm��E%29���"O��A!IQ�����4]-r90"O��V��'�\����w0�{"OVɋb�-���c*�j�$*�"Oh9�Ř>*�����
�z�����"O�ZÐS����rE~�\��"OL�y��Q
��ue ]�`�D"O��4͵EO��aD
 0��k�"O&�$R1=t.��֗S5��� "O$Y�a��6xA���1<�
�"O�E9���$(�9�nO$_>.<h�"O��8g���M����a*ļGJ���"O�E���Lrb�8��U;D� Y��"O�x6�ҜX��a㗢��� �2O2���ٵy&$��1���$�1 ��ɫ*ϒ����,@�X�$�V�f0B�I�.�BMjs�_&?�����('3ZB�o�n�x��=*}�����L�h�C�	��� o\��Z-)��Ȗ����(?q��U�~}�5��M��`�<1ԌˊX��-q��UQ�H�1U�
w�<�a�¢��@` "�k���S&)�l�<�*j.g�=�.Ԫ��_e�<ɶ疼KpxH2'UM�ܐ��J\�<�rُNHcƝ=S$pZ�bRX�<�g,֢?%v���G WE�	��nJj�<���7h�� ��DP��	d��b�<rDث��E�2�r�,^j���E{�G(�����"	�2��x����u��<q�����'v���yU�C�2LP<����&WQ��9�V�4I��ا(��$A�أx�}z��Z��76O�9�'
1��?y�>0nԐK: ���E��E�f^��D	�����?� ���Ԉ;?.�Ivcէm���Z���H�'
v��i�'`��p�A�&��Ua�.��Oڹ��i>��\�`y��S�/ت�����!pz��%�P{7��o�S�.PX�g�ݺ>��S���'�%�'���a���ӟcԘ����! �x|S`�ٿZ�>����(O?1�WDϺd�	�	��ł�"ac�<��?3mZ��kMe�2]
4*^�<Ys�  ���'eV
K��,jEq�<�%[�M̆���d��#u�� ��v�<Q�O q���A(��(�6��G�u�<��d��*��=�t�zA�^p�<U�K�N�0��q�5JӁ�v�<���%(�p�ڇ�w�p�³#�r�<A�čA�Mh/	s$��+��s�<�0�\�P�2��@�߂��!BIW�<�� Й-�0�c��,+5�CQ�<�AI b��e�,j�x��&h�<�r�S��Hf
�*�T�#ĬNb�<�p�O��t���n�"t�ƽ����C�<!4�TPj�!]:�����=T��J�M׊GP�[��(1`��,D�$��h�4���CF�0_?��;�+D����n�?U��P�a��t)�	��(D�v�i�ê���j,�+^Rܘ��'c�0�����8�ʹ匊+j��x��'�\	/Cd'���Tˉ8_(rt��'[D��@�1~t��3����2��'��Ĳ7�ù^�003��%Py�i��'z`a�� ����oV�xXҁ"O�Q��R��m2���e{�"O~���
Ւg|��f�OV�8m��"O��{�jP%H���S�|x�0`b"O��"��t[r:�o#O�\"OT��c�޼G�D����G��};"O<� "Q�Ԁb�G�K��9��"OF,KՇU>�\tq��2\{�"O�Dį��@�y�i�6)�NܢT"O�3�Z�i�D�V��D�aW"Oz��S�L� �q�����p<�"O*Ⱥg�?}�x�Zu%VT�\y�"Ox�Z �I3"\���� ,:̪w"O�$U*.�:�c�@�#m���@Ot�<���4\ܦ�S��R �e �iF�<�0�<QLxPc��X���t�C�<i���q4�rD�O�S$BY��|�<���W|�qhEF�	(�\��NJp�<��-�8vA\�����f3�4��YV�<IuaN��{&b�*�n!s��\h�<���:H
fLЙ�4���Ίm�<��@'NO�E�D
H<�!�:�	���S?�b��v�C�!�d�;�Ԑ˄HG�a�Tat(��=�!�d�)U:,hF���p����>�!���f�p}�$+̀{�d�<D�!��;�p��C�� n��i�cܓn!�1y�J�" ��J�����4x!���+�ΐˑiBS����T�'
!�B�=^�yжK��+�>i	��I�X!���(}���#T�2]*6�1a͌!�σ.2 ��ߒy���cj<'!���x5f�s�)^�+׊ZD�C�{�!�$�|O
͡P#�M�E���	>�!���
�3qO��e���1%�ՐF�!�� �,��l�0���!"�M�!�� �4�se˥H�N�s�)��aQ*��"O�ɘg�ωS��E�O�{1Δ�@"O<4BfIE!g��0���DЀ#�"ObT8��Mӄ�x��>�@��"O~��@��Jy����(��+�"O�ܱP�GC�0��0[ɪ1�"O.��"i�&E��ð�>�.�k�"O@з��&/6��j��LĲ�"OX�C�jB
8��i�>��9;@"O�ҥ�%HcV�۰g��i�DQ "O��`Q��6Yd��(��[�B�Q�"O�lySǅ\��j����\���p7"O&��`�M:����83��ɉr"O¬�0�)[�X��W �F"F1��"O̙��A�"_ܲ��ɪ��/E�yrN)
Ll�����	�~�� ��yG�L<b��d�BVI�`������y�
ڀe�$Qum+c�<ēE%Ԍ�y�X"�YG�C-^Ȇ�B%O*�y«��l���b%l�;f���8 +@�ybM�2<�LAbq�-
^�,��
�y�i�d���r�9|�´3G`�?�yr�7|���8�h�KB�K:�4�ȓ_nq�1�ѷ	N$萦�+O���ȓh0�"�����['Z�9[�̈́�~s��b��!�r,a$EB�2�:Ʉ�,,x2V
����i����%�0نȓ �%8�mX*���V�R�5����!!g	7~u�����ޒ
��-��{��T�&̂��ʔ�We�)-�l���$�.y�p�֨Czm�f)�r�L��t�RI !��+;�4�F��ni�݆�7V�m�"��Q�F��e�%���|g�� 瞹+�A�SI��j �i�ȓ?�*	A%r�lx�Ğ�_v�����s�K�����E���i�`���-��1 !��R��72)h͇ȓP�Ј��ŕpf�u�i�	hE���(yy�B��WQ�|�'���8�ȓj�"�Y��XZ�P�(�*n깄�~�*����	�y���TBD<XSd�ȓ*q^��m��h!<0�&��k���ȓ���1���{��)��ί>M(X�ȓf��" Z�h�b�[�wX���G����׋E�7���$Ҽ~�怇ȓx\t�h`-��7P$�s6"\"h��@�.��b��	=�|�U&�5��}�ȓ7b� �I��T}��	WKP�r�J�����QCːx8�6�3A��9��b�� ϞY�at���捅ȓyŎX�s�R�q�X�x��A�5����^�bd�d�@ ��bBi��<�F���elv��S,�gꌨ*��� �Ą�a7�$
���T�,l�րB�4���qr|˂̀[w��!����y�ȓ	>ژ:�I�es���.�(Y���ȓ_nD���M�8�%�P�ը�2�����cGGD�J�, �Rl�ka*M�ȓNX�z��߁	_$��jӔR�\���0���g�TE�4��c%��sC��ȓ_=4�RDwfe��KW+E���ȓVs�T[��?/����R/T��0��G�r�J�
aĐe��@�7rp��;��Y!	�01�A���S4de��S�? ���O�>+�TMc��	3LY"O~��#cP�Qy�tP�h�
N4Y2�"OJY���N� ��8�i@�dhm�"O�e#�AYN	��&ޮh슑�#"O0�a�k4m�~�c(ҳ
s�}��"O,2��D1,a3L�:;�Q� "O�u�L�� D��e�"Qƭ��"Oޭ[��/�>�D��RW
̊A"OX| f��&q�8r�M|<\�P�"Ol%�r�-%�uʢ�!4-"�z"O��pʍ1m��M�D�A � C"Oބ�IJ�,a��Cm޲|z��"O>�+�(Ē_d���'LJFRF49g"O�8�FJ�{A���*�<1�=�u*O<e�#���KO�M���f���
�'=�Q��#�o���D�r�ؕK�'*|H���M�5vјU!�>�&P��'��%� �!z$t�����G��k�'��G��%�����a��P_�eq�'�����	Ю6u�� ���I�H�0�'���Bl�=���1� ҕx^��z�'njQ�#�!=�TE�F(H�;�xd�	�'�0�ڲ R�,\�+#��?3���A�'��[�l�;ޔt钣%1�XZ�'}d=q�OT(+l.������(Bd���'H60���̅
�;�!V7%:&���'�jh�C���&<0Hpd��(��k�'&F�;�Ζ�5������$���#�'8
0��j�c�m��5p����'�,	#���d
d}8��ye�a��'�ӄA �"G>���mϚ{��IB�' �����C��V8��d	@�G[@�<�&�t����7P��A��x�<�b������(�i��8��ae/F~�<a�fG�`Ɇʧ��
7�N��ZA�<ԅ:S�6}��A�npj���g�s�<A�o1p�u�0
8�l$au�Pl�<��N1Rm켁`!�%V�p��	B�<Yq�D�06U�a)N�q�v�#*ST�<�E
�
A�]hP�L+"pP���P�<��ŋW���	��I�x���+�g�q�<7b�'Z���he H��b��Øm�<9ԅ��K�\T�F�ucd�`��!�yI.~�8�I�G_
���
��y"�,7Cz���^?B� tH�hܒ�y��7C�\����F�"ȑ�V��y�%SA.���J2Bi� � �D��y��b�)��CR�:����ǆ2�y��D+v�^���AL;�ptYrb��y���	�@ب��S�d��ac�B�y"	��j�Bd�T�^�`J�J񫑈�yRf�.j�1F�G�j2 ��֪�y"Ɏ�=�e���K%��M�u���y�fD=���S�H*O˒���I��y��$����hKS��� �0�y���[����$Ets�ّ����yR/�=��Ҥ�O.W2�4�_��yRf�D�n}��K�op �	��y�j�)5�n��FJa8��K�AR��y�Ȁ/I<�0eŔ�{�`��P�y����f1� ��M�k�hI��ˋ�y�oA'!>������dq��T�
��yR��zGJ�B��n��1����yb�?%�R �7.������y
� ���ЂE�'�X�+�.;��2"O0z'�T�[��U�K���6�"�"O�dxV��	�^A��*ɡe��I�"O�A�VgV�m��u��	�$DB$� "O�=��E�#���
--�\ �T"O���biQ4j��-�t� V�z�1�"Oaa�bU*�RP;6�� ��٦"O��X��ǆe=@
�k�=� P��"O�I��6l� A�0�
, �JQ�"O
a�� �Z����g�'g� AI�"OĀ�f:M�T-3�
�[�\�"O�����Ǫ?��^�D���4"O��x�
   ��   �  z  �    �*  h6  B  �M  fY  �d  o  8w  T�  ��  �  R�  ��  �  )�  j�  ��  �  e�  ��  �  r�  ��  ?�  ��  ��  v�    � t P  �* �5 �C `N �V �\ c �f  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����O��=���Y�+�F���eIq���JK\�<1!( )�%p@�ř'#�ܙ�TW�'w|��I�E�J�����{�)"�/�F��B�IX��-Iӯ�7�ة5�Jba�u�	�'XJXw�
P��-��I[� �l��
��� ��{�*\">d 0� o9f�:�"O8����e����!(�"R �R"O
=�kZ�t�:f�C(kA@B2"O���1aT�l��yj'&�8l��u��"O�"3�	K�,@A�˽\u���%�'�剁IQ,h�A� 
��T@* �L���'!`5MV�+�z�i�ݕ.G�P"��HO���Q��cD������z-�"O�܂���u�0"
]�8�Z���	��0<��	XX���0��r;�}k�c�F�<	E/�����b��B���t��E�<��NʭZ� �被�������j�<�R�)����ɀr����F�e�<IcY�n��,��%�T$IUF�M�<QCK�@�������Ip��EB�<�e'��%�!A�*Q�)�THX�@�<Y�!]2yΈ��� �I/�P����p�<٤H�<��y��фk���Bn�<�1�D|L��a��=�m0�yB�E�`+X����I��A��y���':�kQ��h����y�+�F,|��Z�0�i���Z��yRE�!���h2ԋ+
����y"��;(?�h��c�!T��	i���yB�N4�M(���M��9�����M��'7��b)Ÿ4w\��!��=L`����'@9{�`4Lb�,`�թQ���'���(6�Ӿ�x�J!��:����'*=�� �g�H0�- <PMz�'y�0�q��.)(�� ,׃
��"�'n�؋��O�7G��\�*T����'>ys����?ڔp��o֜��C�)��<Y퉟:��|�go�)r)l����b�<!cn�/@���bd��u�*E`B��x�<!2悑D�\)��D�2�svMIu���p�{�cY>/QB��e��0"U𥣗�y򥟏=Ҧ` ��Ns�X���=��'+ўb>i��C��0���2���?� 	 �M7D����ǔ` <2A��c�� �V����xB�Zv�L$��,Ωw��TI2KK��y���c�:|�!K�>̨)�d0-M�=�'9P�	Ǆؑ0��H�Pm�;R��

ד��'��a)�A	>#�����9!�>D�
�'�����I�O��� 䌑�q ��'p��˲d̩��,�@f�Յ�;�yRK��|��� ��wI���V���y2���q�h���F�.#Z|XƬȻ�y���L�\�c.M�%�������yRdհg_�Tٗ"�>�IEfނ�y2��^r�9�%�/�0�0e`Å�ybOڪQ�n��T��"��Q�տ�y�gS�+�T�sdo�3_04Aլ��y� �?/l��nK� Jǝ2�ў"~Γ�j��q��	���[�
�)|R��ȓEA�y�h5T����Mȇd������?9g/�r_8��֎ط1�@PgDx�<�U�ъl��fS4+�8 d�r�<!�B>p� K�V� �z`��$F{���Ŕ<M\�0�	��j�d%��7�6C�	����b�)u-&�:��]5C��/}����LϪm'��9�Fߟ6 D����<Q��-se��#�_>v���z�<�N�	s��L8'U��hS��t�'#�?�hd/� d,��7\�xiSp�7D�� >}6�ͫP�D��#�շc�`��e=O��Dz��IG	�������������D�Q�!�$�]�X�k$">n�R(@'.�&F�Ї牑I�I�@̙ �`쏨V�C䉪&D$![a�!��E�	��B�	�N�@�0s�E�$$K�	��(�pB��Z�Vi*R���N���F��C�I�q[�0�*��Y�0�I=��B�ɷ)�b}�r*K��
�ę3�ZB��8Z���B���Y�&�Q2,6�_8��?a�@ăD�X�@'�!&^�vc�}؞� �Z��j�41��p���-VH=��<���ȓTZBmqB��*J�����i�&�m�/1�	[�Ok�̸��&Ze�πri�	�'~l���G�E]y`D�B'T�
�'R�}Q��8k1�X#��)3���	�'3ġaǦR��jY�ťܱ|���	�'2\q�Y�&S�$T�BvRt1	ϓ�O���#f;�6���F	{eܩ9�"O��x��Ž��,Jc�ךw}�!㗟|"�i�2��>}ȱ�U?Eɴ���Δ��@�1�Cz�<�gC� 8�`�_'/��I��u��u�p�$�>��O�X��̙ƌ�(1�q��2F�zC�^�C��R�z���!@ǐdJ˓�y��S�\T�d�����C�G�q�:C䉸:��br�ʄ0�l��G��dC�əZ�*!h����`�H7cǚd��B�	�>x֤b����R6� Aj��(��B�	!g��F�P�(��q�M�(��B�<6e��b�D<h�p,�y�B�	e�̉����<>�Xt���J�CƲB�I�Y�X�;��ݡc� �;e<]�B�ɈZ<��4�T�����$�B�	�Qiڹ�R�D6U8���_�K�ZC�ɐ_�Ȭ�JK�QT��wR -�"C�ɷ8e��X��F��Ԫ��"6C�Ie9he��Ԍ��ȉ���3lg2C�I�6��$��CT�P���:�%�7^`�B�ɶId�h� z��L�< ��B�I
T-� 
���d(fp(@��F��C�����
�/"�bV!.��C�	�	i����S���t��&��nz�C�	)��4��J� `��f��6B��.�����A*b���ʒ�n4�C�lR9
$�I�T�شk��B�	�+� � �BO25h�!�5N��Fk�B�I�jhy����8 �!�*Ћ�C�9S4�@��4&��p@�*W��B�ɑ�H�CA�u���+�d9�6B�ɹ!hآ�R�tȐ`��=s_>C�	�~���'*�=;*�P�`*T�-QJB䉠6]D�jt�9:,�T�k�?t�(B�	8Y=��Q�N}�,��lN_#�C��"�*Hs@�C�l#����L�4/�C�� X�@Y�cƇH��<�Gi-�C�I�<�Mp4!��F/�dA�f?\e!��� s.�IeD$-,��GŚ�@/!�ă�C�5@3l�})r�⣍:i'!��%	�4Xg@\*&$X�c\��!�DΛcT	�m��.���!@\�!��]e���ZP���J}rS���0z!��P��[���;w��P�Cτ:f`!��6�$)B��.�:�P��<w!�d7%6���bސ����v�Mb!�� BQ2Vk��48u#��5[����"O����(ð��4���Gߴ @"O�X��/ݷ���ÖHڤ6����"OAQ͆�a)��PDʜ�_Q.eS"O�Ժ�坎z	��;��k ���'r�'���'�b�'��'a2�' ,x��u \aZ��S�+GT8h��'q��'C2�'B�'b"�'���'�T��!�	�ȼRm	%xmF����'��'�r�'���'�2�'g�'�&�Z���=7Й��)�
	���/�?���?���?����?	��?a���?��E�)���Eo͕v.�����?	��?���?��?����?Y���?aAO�+P`�|8�LN�n��p�KR:�?I��?	���?a��?!���?���?y�$�3X��[��[dd�Q)`D�/�?A��?)���?���?Q���?���?�� ȣn�$s�[�S�t0��Y3�?���?	��?Y��?���?a��?��׏������[Z�*��D�L$�?����?���?9���?���?����?���C.8b��"t���b�S��?���?����?��?q��?���?Y�f�L�� ���)O�z��TL�3�?9���?)��?i��?���?���?I�e�N����ݰ\��	��%L)�?���?���?����?����?���?ač��d�4�j��@�^��,r!�E��?���?1���?����?������'�B�Q;`@ah� ��0�%�m��B�˓�?�.O1��	(�MӒ��5m-��*�.I�$-gAOuL�X�'��7M<�i>��@����/�v��,� V4ȡ1�����I״�o�b~R:���SD�)��[���f�G�E�TC���]�1O��ĸ<ɏ�)�$Eڐ!��J�
)��͈î:�%n�N?^c���Jt��yg ׂg�H�Ok��ږ��cF"�'���>�|�D�@%�M��'��ف4i&�bT[�&@G-��'�����Pa�i>�	/��l��冲s���ȕ*_�O�0�vy��|B�a�����_�>��#�㐈Tt��M�t~���Y�O���O^�Iz}bO}x�� �Ds�q�U�Q����O�A��*�#4l1��E���4l��d�i<�#W���h����fZ;���D�O?�I�(�&Q��!̫e�8�ףހ8���Ɏ�M��MXg~��o�t��%�Lx�Uɀ=%$�iRb�%u(Z����I؟̘�!�����'m�)]�?-31�<6K�D	W�2@%aH;a�ў�Ry2����X�*�������4������Ȧ](S�2�I~��f���$�H�sn��;& ���
�R����០���'�?i�^i.=+��F�( �AЗ.C�,!8�rnߧ-�j�'�U	��Is�B#T������	0%�9т�P�H�"�9%v.�d�<I)O,�O�lZ�f�͓U�iˤ"4��ʳ�C�2y�X͓J�V�4��$�OJ���O���Y;�
�#	 �(�3GB�J 6�f�ts�ğ!6�O����8(��H��s⍍EB�Y�#f?��)��<q���d�<E�4j�6g�����'�6g6Q���\��'H 7�~��	�MKJ>�0 \�<��1���.��j3�� �yB_���	̟���3��m��<i���?��Ѱ.�J\�`AV�Wnn��2�o�����hO�ɵ<��hD8Z��	̽k!b�
"j�����5q�&
���'E哜T�l�N�5e&ֽ#sM��2��m�������	�<9O|z�A��x�t��X\}ٱ�$G�.����#!Ƭ���s~2�'B@����g:�'M�<��ؼ-r�r�%�X5&4�5�'���']��Oe���M��$�2� !=��\ʁ��2$�=�(O��nN�9��I��M#ɝ*����)�� �Q����mZɟd��#�a��?a0O\�G��1�1(b~Ϙ!Qhlp�V�%%��Ώ�yBU�����$��ڟx�Iϟ@�O6�����]�Jl�a�(U*,� `���ʦk�O��D�O>����DΦ��3���ӂ�A�<|;`�Ө;`
��4h_��0O�Ş5���ٴ�y"0a��Y{�H!n���Zc虅�y�/��E� P���ݠ5��'��i>����F �$%�%x�bI)�V�DS�I�	�����ğH�'.7�F�|� ��O��$Ux�(4#���1��yH�i�$#P���O()o��M�'�ɝ��J�
�"t��)9e�G�3�
�����B'b�P�$@:«"?1��8�٩\w����v��	X�K��~�*rf��Y
���O����O���|*1@�N���'��EL�Zy��e��&)�hX �'�"6-�T�(�
z���4�������ej@r2��FX���?OXHl��M��'P�-�ߴ�yR�'f�<A� Ly(�I����Jq�9ᤍD��De�a�pN�'��i>��	����	��4�	��lpbQ�s����߼X]�'��7M[�q���D�O��<�9OVj�x�D�(v��!�v��>j�NU�'�R7-MЦ���ħ����$#hX��(a�J����߮�
$;s�9qQ���'dEj��'A��n�p��Vy2C]T~0�$O�@���D�@
��'r��'��O1�I��MkA��?9��������8��2��33�����&�'Q�'���?��4�?!FA
4r�^<�E�6�2X�IS4��۴�y2�TK�29H���Z�:���_wo�]�q�? D�S��@+b��r�M��g0j�;b3O��O��$�O8�D�O��?����K�̄iA��-PRP�92L̟\�Iڟt��4q�m�)O�lf�	�������U�u`�!N������mٴ�?9�gE	�MC�'$FY��ě-�=j���t�"���ϙx$x�G!ۧ4.|aJg�xR/�<�'�?1��?�ģM,R~��c@Y7U��!i�4�?����A⦱S ��8��蟀�O7���c
���t�u���m�n؀�O\��'3~6�����̓��'�*�ʋ)���z�N�tq��K�j���82��q�t��'���'�h���Tz�K>���G�\8U=&eX�j
{=����ܟ���ǟ��)�SWy qӨ��n��DWD�J�]3#��Rt�C�|���t���\s}s�,yID�ӭ�Ha���&=`��4$�զ���1�|lZ�<���J�}�3��H�(��'-�)X!i$q�h��J�)WI��'��	럠�I؟����L��F��Q�&��mٖĆ>a����6)�,7MX0:ږ�D�O���;�9Oȩoz�M���5�p�@d�5�V�ː ɬ�M���i��>ͧ���XL����4�y�
�*��5�` 
�R�= Y�<��e�2`�!�U�+�N�M>�)O�I�O�E3�Kb�89S׈��a�����O��d�O`�d�<Q"�i��c$�'4��'��d���œsvJ����g=�Uɴ�$Fy��'#��2O��
]�	�M.v{^#`N�ϥ%w�x�	�=����q`��V$R���d�­�u���O�պ��˼$=
�Ci�訃'�O&���O����O*�}��
ܜ*�%N�s�-e$ѫ{D����fD�v)�)e��	��M[��w@�)&�>N���UH�;MnԘ��'�X7�������Gq@nZ�<���FJ�x���V��Sq%�C�6��C&75�m�#D��䓷�4�����Oz���O��ēz`���B�!:c����52Д�z����7(��	ϟ@�3��$K�dɥ��j&�]"` �7��I&�M�'�i���3ҧQcF� �G��tG2��`�4�a*A�E7z���'8hH�t��ʟ���|bP� �R%�1Frh�(E�b"F=;�+Xğ���ş������]y��{Ӕy�l�OX�Ǆ��!�|`$ӕg�f�ْ�OB7'�	���O�6m�O������Q:$���E�.Վh���\��7M5?y�M'?h,�	0���56�۫w_��U��&
`ޡ�D�֊�y��'j��'��'��	κ��e����<#�HZ`��/2"��D�Ov��E⦗�#�	|�po�J�I=4� I3�
M�#�CV��$�ϓ����٦���|"4�8�M��O����E+�\���x��"@*M������x�O��|���?���i���pd�K�h����
�F�����?�.OF�o�/0�Zd�I��`��b�d�'\�A#	B34k���2�����O}2�r��o��<��d#A `�9�L�
~�"��d>r!d
\:/?�]+�O�)P8�?�WH!�dB9`Y*is �ya��s�4r�����O����O���ɶ<��i��5��ゾcG���ra� yD�8E��i=�	٦��?ٰT��ߴ^�"�J3�]<ob��5�
D,����i)�'�y��8O����(����'?���C�B�c6�R�.�\a�f ^�"��zy��'�"�'���'�i>Ї��4�(����^����D�T��M{�ɋ��?y���?)H~j�'���wG|yK�ʎ���A��� Ö4*t�w��m�<)�O1�b,� g�*�Ʌ@�D�C�M�B�(� G@4��I>��|!��''4D'�x�����'L\��
X6\��FR�
��iR��'�r�'
"_�$�޴cV�|K��?���r���kA�E#�9v�݂P��!9��J�>鰻iKB6x�@�'4�Z��2C�aB���"A�����O�4Ò�M�:������	9�?���O�$CD��pT���p�� ��#��O8���Of���Of�}���#��Z�5:�xH���w��4Y��F�܆j�����?�;i���~^�AP��V!VXHΓ?���Kk�Z�Ā��Z6M2?)���GV��� '�b��]C��G�X805^l{J>/O�I�O���Od���O�	�aTuT�t��@�i���`ζ<�b�i2�pZ�V���	]�'=uT�q£Ĥ:�jt��e��+�����U����4}\�5O�"}�F���D��U�>���D⚯b���ñ-�}~�ą_��=���{��'��	�>i��8R�N2D|x���/S���Q�	ɟt�����i>ŕ'��6��h�6�$ �(o�i� ���p��6$���f�⟄�(O��{�[o��L$���+ ��)*��A&
Hhź�1(��H�Z%����>1Yc�>�{�g����dׁ���!�'~��'Q��'���'��H3D8���ذdC{��s�g�OD���Or8m��lm�d�'�V�|���( 	�u�[��f���I�'����c�4�?��l��M��'�r�7(9���4�:pD�D�0x� ß�Q�|�P��ş���֟P����X�*L���	<fw4�V�͟\�	]y2By��x��O����O�')��Yp.G�s�0����y����'�*��?ܴ�yb����Oަ5��� 0=�!�ei�B�T#E��ԉR1�؁�O��i��?A$�2�dƀ>NT�u�C�\g�c��;I���d�O��d�O���<週i�$GH��7�̰�A���<�*����*p��������^�	:��D�֦}P@Mڱa5���C�X��(��(�M���{C`���4�y��'Ɇ�{�(��?�c�O� ީB�G�66��:A`ċQ|���66O<��?���?Q���?����i�+Ό#5*�5z��`؛*R*lڍ~�D��	�0���?���~��y�չsۼ���c�;")��Q-0�X7m�֦�̓��4���)�O��h��i�T� �N98��3���d�C��8O�rퟌ�?���)�Ŀ<ͧ�?��L.#� ��ş�V2��@�R��?i���?���d��XkLПL�I矴����~�^��� ȴ[����A$j��z����MK�i��d�>!"�Kb8$b�)�i7�!�aÊH~B�S���5C2�F٘O��)��YE�%*#���r�R`NL!#(�QB�'���'���ן0X ��@��ȋ��?*x�p�`E�����4)�*���OH6M/�i���f�-��ղ��a�j,��`�Бش:����'��Ң��=��d�04��q��jD��:���,a����Gi+�37�:�$�<ͧ�?����?����?� ��7�~�;��
!��(�FNO��$�П0˰��<����O�`�L;s�.m�2)!����>�A�iS7��q�i>���?�
W�L�b���(Do�
_zPE)H+�k��$gb�IU��<
Q�'���$�8�'��s&oڋ$nIЀc�/n�"`� �'���'m2���DZ��ݴ]�Y ���Hu�P�P���Z���3��)��M[�R�<����Mk��R��*tʝ*�f��U����D��M��OF���.A������`����K:M��H�8���,A��$�O��d�O��D�O��;�S<C7z��A@�0E�\"E`�*��ɗ'7"�w�v�*�>�d��Ӧ�&��8D��Ti(ŀ�ʎ%��l�F���<Y�Ov%mڦ�M�'`��,B�4����!2�(ɺ�+�Op��(ãК&PH�Ycf��n/8��'��i>A�	����I C���Z�-��-=�e02�Z%~������h�'��7-ߦg��˓�?�,�B��A�`���QoٶAt�=�Ӕ��OB0l�MS�'ñ��5p@�q�ij @��_Z���e�[f��P������i>�I�'$�'��{�k�ab��i4��'~��������Iȟ��I�b>i�'��6�=kƆȡ�⏋Bx�@C�F�~��Ku,(?��4��'U�����Q�ExJe �<-Av�b��8M7��Ϧu����A��?Y�ժd��	���D�m����G��^Y,xBp��N��d�<���?y���?����?�-�T��p�§�F�!�C�`B�dQ"�@ݦ!��韸�	ޟ�$?��	�M�;+�$k��4�,Ԑ�)�#0�Ʋi�:6--�4�����O��F�u�|�	([�N$)��9)������{ْ�ɐ"Z�Q�"�'Y�t&�@���D�'t>q��C�h5�Qb�;=���ҁ�'l��'��]��ڴ<��	����?!�� �p8��˙o(9�!��b�l-A���>�@�i6f���' ܙ �J��lա�� 9H�yÞ'�b�V�:c|�H�n�=��������oHB�$F�3�$�!��_]ȈWD�:W��$�O ���O��D!�缛��]�6d��[��'`X��"ʸ�?	�is$��$��m�P�ӼS ��"	{�E�'�:)6�T��<��i�.7�O�����u�6���papE�))��tc�j��"��/hq���U�_��'�`���$�';��'f��'Ӭԁ�'Oa��H5���K�l �^�Ęߴy��Y:��?�����<���h���%U�~xΙ��e��\��	��M�Էi��:�)��N��N�qKr	�򁕓u�d��;%X���e샠?����w����'W�&� �'�p�ڒd(eܤ(�g`��N	��J��'*r�'^"��DQ��A�41��!���KJ��SS�� ]M���+��&N q��M��b��>�W�i-�6-�O��[R��x�� 1D�t$��'�\�	��i_��O�A@�$W��r���ӣ�5��Ө>��	Vi;c�$�I
/�y��'�2�'���'�R�Ɍ��|�Eg̢i�h)�aJ�`!�ʓ�?��ihP�ɟސn�f�I�B)I��:�L<���WN�r}����O07=�j��dh�l�H��)Z���΂{!:]n�2�fB�]k��$�1����4�����O��$W�TkT�Q GD�i�Ɖ��;d���D�O�ʓp����95�2�'�r\>�8ï�2	rh;qW�
�1��*1?��P����4Dn���|ʟ��@B�K��y��C�@ΩP�A���~H#���s��i>%���'�T-&�8��Vx�n����8^�ppH&���	����՟b>ɖ'��6M� xW&l!u��h�v�����?�$��e�Ol�֦��?�QW�ȱߴUꂹ�fCA!-F.y��EK	
{5Z��i���ΰH�V��h���P�"����~:ƀ,B�:I"���8U�hH8�AN�<),OV���O����O��$�O@˧=���ƄZBB [�(���L���i�hm"rS� �	_�S�<I���#c�^) �ޭy�R�
A�$jC(%�$|��Ij}���bI2-l�3O�H���$|��UB�@�;��m�7>O�I���?��N>�Ļ<�'�?��K��>�A�D� .�~d��L��?q��?y��� ¦ik3' ß ���g �6np��v
]�Y��J�d�^�[���>�M�d�ir�>�,���Ȣ�!Q�uP%z�.Ec~�!CB�hq�5@����O�jm�I��C�1-�|؃EV:JG$T*5��4Sab�'��'���s�-�����r	�%j+`t CH���"��Z����':�f�4�\�a�iA* j$x�=p���9W��d�ꦝ0۴p�mӏZ���0O���3�X��'	�� �BQ͎l��hZ�e��r���+&�D�<����?����?����?��E<g�.�S��s��B$,����9�pc�������%?�I	q�����+�7PVA���2;B�h.O��DkӞ��s�O��Ȑ��N�zI1�҆H�ظi�%ղ{_�<h�O��q�&*�?a��=��<i!+(?9���1-B@6L��?����?y���?�'��$�ͦM�Q��˟�0�oJ<�(� �B�6-8�c壟\m�J��4x�ן�m�ȟ�1��͑x��a��S'WV�A��UU�
�n�^~���W]J=��k�'=�k,JKPB�� l
��}{�O�
���O���O@���O��� �S�he�`�AL'u#�A�ӂS����	ןD�ɮ�M�"�Ԛ���x�|�OL�
�$�#s� �pq��h���t�0�'�6�Ȧ���N�~�l��<��W�-y�\Tܹ�ȏo��e���
��'��$�t�����'q��'�x���E1f5���2�$��-"�'2V����40D��i���?y�����\�(by�FB�_�Xbe@ J��	������4�y�iFU� �B�"����ĝ��vdAFŗa$b(:Q���ӧ1�B�Q�ZAȬ�r��!
(JԹGK�����P������)�SIy�u�ذ�������1C�ln� N������O8�m�W�E�	%�M��ٶ
��)��$(��3ŧS!"��'1�Ұ�i`��O<��AD����x���J3n�##�ȿ&?�y.i�0�'���'�'�"�'
��1I��A"7�E�]ghY�N�mJ�K�4@x�����?���g?�����2#Աux�!��@c�<�4�
/7·i�d�<%?�84��'iT�ɼ(a"�G�K<�ڝ�f�=R��Iz��|���'J&�%�x�����'^$!e�*gRHQwD�0x����'�2�'�U���ߴy�:�k���?1�;qB 
�.P6��E`�
�N����>	��i46Mv���'[���酮0��8#ӯ�y�ƨj�O6�qP �G�
�I��ID�?Q�K�Oh=�3�R<J¥��H7���rw��O���O"���O£}��o���� �O�?V�����VX����v(���:O7'�iށ���ݐ!��1W��d�(q�Jh���4����'��S��B'��dT2�4s�'_�x9���WU�]+��ӰKŚa�7��<ͧ�?����?���?i��ū[f����QuO.=�C-&��D���	���Qܟl����$?e��<0��$�Ѳu�0	7h�_b8Y��O�oz�޴�yR�S23K�T�AŢ$rz��h>��(f�T�o9t�*���@,�O4�RL>�(O��Q�;t����7jZ4�Zщ�O �D�OF�d�O�<i@�i�F!�4�'
����E_�c�.���2W�'՛���~}`nӬ�oß�����	A�����,A��Kݕy3@�o��<!��]��i���'?���r�z�Ε)�Q@�)�F6�B�J}����֟l����4�	۟|�
��V��
��#�x�Z�� ���O�oڮh����<��4��'��L��a@�d� !1d���&�F�A�'��	�Mkg����@��-1�����uJ���թ$��#Q�jؚs��\���#a�'�<&�������'y��'�X�j�$�B��ؠQ�H�U*\�(��'�\���4sU�"��?����	�"	,:���L
O)�@a�HZ)9��I��D�馡@�4�yB�)^��qJ��.��Y�v'��U�G_�t��q���6*��w�	�Zb�*�2HN�t[�&BD����|�	��)�Scy�cg�� w��+[^E[�'՜g������V�j��MˏRj�>�ŷiT!p�h�0	jd���(Dj���@Cq��䟇1�7#?�E��$1j�)0����Rgf\Y��Y�Z�Ԋc,U�ybV�`���h��̟X�	ӟ��OT<p1�*�Є��&�:0��+�b��q:���O����O����t����AWXp��OtP�r���0H5o��MÛ'��)��3�:m��<����9��Y"��َv�.�2�O�<�3I�%3X�����䓳�4�����m���`M	�3B�`;d���<j���O���O<ʓ}��6�	�!3��'9RJ�p��q&�Ӭd���fζg�R�|҆�>)��i�>7q�x�'A���ub	� q�x��-b �3�'w2%�8W�ꡊ�
�6��d럪�{�|���$�7B���7x����rbF_�B���O����O��:�'�?���پ2�� ���$�z!8�F9�?a�iZ �2��'���xӖ��ݴZ2H���DG@sTQZ燑� ���ɘ�Mk0�i����7wn�F��lZ�Q8!���į�>�Q_ux��R��'f����|B]��ϟt��柸�	����k�`�޼����S$��ᰍ�ey�y�xxY��O"�d�O����|Γm]Bz"ߋs-Z��ϝ�?"�&W�p�4�0O��:���O�rЎ�@��T�'&c��q�T�����l8Ƃ��BQh�Iiy���*m���|��ٲw�H�M2�'	��'��Of� �M��ˆ��?Q�	�<�V5��;� bC��W?Y�4��'u��5����n��\�U�V�@p(�0h�ޔ�G�],rj�4#G�r�.�	П��Eb�0����0?��p+k�X3��=hU(�h��''�,f\���O���O��$�O��=���s'�H@��2^uR`ƀ��H�`��˟�I��MdZ��dr�P�OF|���-�`���H�*�ͱ5�d�0�'������Bp�������g1� �py�O�-��f/"�{B�O�?�C@,���<ͧ�?9���?)KE≮Dc� v�M��͒)�?����?9�8�d����?Y���?1���4A�2�h�W`�>c->�C������$iy��'���On���JQ\Tx�$��)7���'�OϨ� %��D3��O���R
�?�2�&�C$V�J7�D��|0B��X5�����O��d�O��<���i� �����t�n(��Zi�&�0]�*��I��)�?�g]�P�4RX��Ʀ�$.��U*yP�a#��i�R!��G����pcSeR����~jÀB8CO�5�F�2���� �b�4j�%[`h�QC@�<"�Ȱa�I�hgʕ���8��`c�	J���a�X��py��nG����K��+�VE�Ў�e�ND�`kJ��h��S�� �h'M@���d1h�1<���o�`�g��<�BgO�5���`�6eQ��L�!b��A�b��t5N�Se��LH��L�!��a!e�'?�@*�/�"�� $0 >�xв�	�<��!���B;n�У�`�3��j-�>�r�s�'
:4��X�HS�q�	�FƜq��@�a]�)HD�NЦI��؟��	�?yJ<�'XuN�� 
�*�����Q�|�F���`��'��G�s�T��Q�E��AҰj��,�����V� �޴�?��?q%�_�I������'���͗s�zl��i!SV,ŉW*3O��IWy�����'���'�b���X�0��
!z�rjeE�.�7��O^�pWo�N�i>��I��\�'�X�02��`�VR�lÉP��@�x�b�D˶<�1O0��O���<"b��Q���%��,�t�ӱ�84]r�XR�x��')��'���ϟ��ɾ:qFX�#M��@��@�ֈƷ,&�eC"�&�I��,�	�'�L0aci>�9�G�Į�(����")�`�&�>1���?QI>9.Ob�afX���2�� ;
L	d�B�@�Rq٣c�>���?q����d���<P$>�b�ˉ��dR�KV� ���Єk[��M����?�,O�D�Of����	�7+�4r�I�dϐ�+��Z#9�lZȟ��Iry�������k�ּ[�(����T��!�G�%k�'��ɧ1�,#|��O�fbѫ#�4Q[F�3@�^(�۴���-�,n����i�O|��`~���3o.&��f��.b�ԡ
��A��Ms��?�A&
���4�@����'͎��:H>�����W�'�F���4U��s2�i��'e��O� O�I�j����"J�$�`��#�4ja��mZ�Q�����D;�9O��<;~6h����<O"�b�v��%Lh�N���O ��P0M�T%��S��2;���"�K�iµJ�=�6Q�']�I�T�c���I�L�	�4�>��4
Y1"{*�8�`N�C�����4�?��#�dd���D�'��P���+�	��*��T�"iڂ���M��Z����<���?��� ���X�	�7f/�� ������S�j�N�	����Id�'���'��!s��
]��1pP�C�1Rx�&>��'!��'��Y��Bg"��T�>�$8�����0k��ݲ��?i��䓦�Վ	�ɷ4{:����-o(v���t&���?���?9)OXE��N��of �NM�&�1aI���ٴ�?y������O���RvP��^��H�M�&AC���7H)D�9b�iG��'I�	�EDjL|����1C�`�8&'M�c��<�wʇe$�%���'�ȵ���)�?�J�ؠbf�Q"���S��I�Q j�`ʓlȘ"A�iQ��'�?I�'f��I�8df����ɑo��h����1�d6��<����L~ʟғ���m�	:�v�4�03�q��̝��M�`�����']B�'M�4M3�4��avFI�W����O�	_�U�����C��5?y/O������O�P�n�x�8D�!���<dT��N���}�Işp����-���D�'k��O�PYC)I�`YuӥƓ�2jp � D�j�6�,hכ�D�'0��ORM�M�L�gü>!��	`�i��M݀\��	�I���=Aƍ��Z�xG͛�/�z ���}bmT9o!
�O���Onʓ�?!����AH�8�A(ɺT��$`JJ��ݑ,O@�d�O��D0�	���a��~j��a���1.g�5�Eї*���P�5?���?i)O�����Q������$m��d��|ʒ�c��_ ;�6��O��d�O4⟨��=$�4@(� `�T��Fm��>���;�d�C?�As�R�H�Iӟ`�'��c��z���T�6퉰1F<a��+���typV���M���'��a̎��A)J<�i�Uq��(X�%���	���Ijy"�'F�t��Z>!�I՟�Ӯ	�b𪇂Ίqe�Aa��(2�"%�	�<������b��' p�1���c\8�3��X� ��'5�#�5�"�'��'P�$^�֝�~\>��F)QS��҄�|M�{�O*˓kl)GxJ|�����U�b�rAP�%Eb�P����!7͝ß��	�����?}���d�'#�s�	@"����JV�B�F�Y"w�"�x��]
I�1O>��	4 ��4�S�-��Hr%j׏3J��`ݴ�?����?���	��4�&���O\���s=��!�$I�&�2]�lu��y��Cd��f���O���5��0;ƬݠQ�θ`��� vTx�R�
��,O����O��D1�uR�����h�:�a����szJ�#�JM�!F�\~��'r�Q����f%VH� �D�F�t(;CC��3�E�py2�'e2�'��O�d
=V�!�����!J"�E.����Z�6����8�	yy��'�mi�ܟ� �ܢ�!��fKb�G��Йٵ�i���'�"���O���FH�6�Y��e^1_ںe���\�����O��d�<��qN�#.����N�(��[)�JL|��E� t&�n����?��*�<�F�h�I!�������5x^�sfF��27��O4˓�?q�D���)�O������9�-�jcBy��٢[#�A ��m��?Ydk�-?+Tp�<�Ouԙ����~J��"��)Lh�O*������O����O��	�<��L��Ҁ@�m��:GLk|���'���0o�ƥ�y���J���R�*ч�<�^�	Q듓�M���*�?I���?1��J,O���O>�X�l�<3kr�2�EZ�L��9�3B��r'�Jc�"|j���~)j�b�:q�
Di�bW>E�N��лi���'���U�i>1���\�g8� @��HD(2���(r܀Ȋq�D�>y�~5%>1�	՟��E����&Q��iU�_�B)��l�����sy��'���'�qO���uI�:R���@�ԭ`�W���&OU�%Z���?������O0�d�B��j����Zs'�.H<˓�?���?q��'�4�牖�7���R���W���	ʵNa����O,���ON��?��ž���ɂ
 ��ᇁ^���S+�;�M���?����'B�M^*ٹݴ`+�P`��2[��@���&@+ND�'9��'��ٟܰ��]���'`(��!�b����G��-�m�!�h���:��ߟ�bm�&WHOVM�1�R��Y�́�LRH�h1�iU�`��#T&��O��'b��b�zf,�h���T���G(�8�c���IJ�eJL:�~
 ���C�`��į�1$�F�b4�Ds}�'�v<��'uB�'���O��i݉z��b�����!�|u�d�>���#K�A�DTw�S�n�*d!�I
,�Q�T!E��mچR�0�����D�Iܟl�Ky�Oy�#K �N!�"�؋D�A�R�S�|6m��N"��f��S��:ՎX1WRx��h�R���v�׭�M����?���!��2-O��O��Ķ�0�f��f����=:����CҌ��'��q���-���O�$���D��'�:�A��"o2���lӺ���<8�ʓ�?����?��{�$ �M*x��eL�Y(�Q0�f�����S�"5������I�|�IEy�I6��ġe�ݴn��y����z$iC�-�d�O���*�D�O����W�H�YդƸq[`�R Fo*
��N�O��D�O��D�O��D�O6�D�S+�	nڭ9���y�DL*��ؒ��06�\�N<�����?�2B �=/|�JB��I�9#1�Q7Hƴu�i���'1R�'�剞_��1��P���.�6�i��0L2`�E��o�ޟ��'�R�'{�A�	�yr�'��$O>��yS��!d��I$�������'p�\�������)�O��� �PB��:��9��LJ n�T��jZg}��'S��'S:P��'��	5k��@���E��M[
��U�`�ۊLz�\n�cyMF�;(P6��O�d�Or�	�J}Zw[�$9Ue�~	��H��4�?���r�Z���?Q*O��>��@b��(q��WƐ��HE�u�i�*УE�ܦ�������I�?遫O����)�G��e������!��0;�i�b�`�'�"T�����p4�@"�$��ch�����7��ղiE��'r��[\6��Or�D�O��d�O��B�)�*9P�G�
kh�k��^�X*�F�'��	�29��)z��?��)ߚ�o�/x���QM�ĳi�r�/�6M�O��$�O����V�T�OH�'	?u��9�Q�Ǚ":(��[�P;�$j� �'���'.T���J�s��X�pa��]�Z�q�cʏ
��*�O���?a-O��$�O���Z)7�C��;T��M�w��5v`�5X�1O���O�����O����<������I;E��Tb�f��6z��$R�R�&X�0��by2�'���'\��!�'��ј���l��8�5*�-%���?8�I�_����IΟ��'l��+�D�~��D�T�Ϥ[z���	�-5t��E�iBZ���	� �I.b���̟����m��ar�*8z5>`<��n�����	Ey"�T;0�'�?I���)N  ?���R,[o�0M9���8���֟|����`���h�p%����
���*L!~�`V��V�f�nayR�%2��7M�O��OZ��x}Zw�t�%%Տf���a�Z�g�x%��4�?��l !� ��S0Oz��}�����0sT�BkN7��Q*�C����*rCN��M����?���g[���'�D���˰y�m�Ձ��B"s��D�ہ1O2�O��?u�� ,�֍Z�lX�WV���lȍpA���4�?����?�q��b��I\y��'��$@0�:�js�ȬoD����M�."��f�'l�	�r� �)2��?���0��$`��	i�����,͈�ã�i����Qش���d�O�˓�?�1=s!�o�=0��`��0�Ҵ�'K\$;�'���'���'@�Z�$zu�[�$�"qC�X�R�������S�O�ʓ�?�.O����O�����<���TJ)6Ͳ�"�ѵ;�}�s2O��d�Oh�D�O$�D�<)k����
q��2���:��"!CB(5��^�P��My��'gR�'��C���WȘ6d�N��w�(J�h4�i��'�"�'��i��с@^?���B�����I6n��E�����n��dZܴ�?Y.O���O�������O4�$��~�3wlT��`X�&�S��<x���O��$�<a�
�T���Οt�	�?E1� Z�h'��.���qE	V�&�-��T�������I,_����?%Ac`��uc�X�&��T�>�c��s��gġJñi���'b"�O�>�Ӻ�r���U��J�m��\�G!�������h{�(`�43���=�ӁCM����LW�k͚�k�J@���7�ϭx*�n埘���P�S;��ĵ<���)�n��V�U�����Ձ�O��?��I�{���۪n��Y�*�lq��ܴ�?���?��D#���jy2�'��E1A&�h��ȣJ�h��fA���V�'�剧L�)���?	��1A��!OE�6�c�'G�8���Ÿi0�G�/`4�Oj���OJ�Ok,����ː�T�e\� i�	���"�L���EyB�'���$�Ag �8�f�J�Vys�,R3p�*��i0��O��1�$�O���90j�:$�C
^"�ز�*$#�Bh+��6���O*���O<ʓx^&�K�=���qV�����.5��)�N�H}��'�_������ �	�"��r4��фdN�6��YB@�Γ\�
��'v��'nBX���܆�ħ/hH0��@#`�h	��R�3��a׶iq�|��'pbB�yr�>1f`C���K��H�̌�`ud�ئ�I��'�XM:0O<���O��iA8WM<�9$�O�T"�&D�0�:}%���	ȟ�X! ���%�p�'j��CmH0 T��f�=F=F�n�Py�0��7�Gl�t�'O�$�>?)�N�*xdT9ʴ�E9tv~�{gdTЦm��꟠�̇ϟ�&���}�g�8_r�Z� �2�r%H�C���W�K��MS��?1��*�x2�'�`���h�7_Flx�*
h����r�α �7O\�O�?����q@e[�oϲ�B��ڨ�F��۴�?I���?��N���O����|0�b\�\�%I�!P1(� dz�Z�O !�E�t�SƟ��I֟�w�G(R{�Ih��B4�ڵ3%γ�M�EJd]h��d�O8�Ok�W�C�h�ô�ث0gܠ���ܓHH�ɐ%�p�IDy�'wB�'�ɟr�ق�݆Y����<a�@�1g���ē�?�������O����OF�J�ə!9;8%�穁�4��2�&�l��<����?L~j�	˛(C�I�� �~�P'��?eF>�����-%�������Py�'���'��й��'BR���F�9�2�+���`Ѧ�qK�>����?�����/5d�%>	�QM_��.]�5KG�'�`���+�M#�����?)�^.�� �����~���͕!��x!ĕr2���iH��'��I�!b@�N|���B��Ϻhx�hAƁ�L�n��P�H�W�'���'<��K4�'�ɧ�)�7/��[�H	�|mlY�/�=SO��V����҇�M��T?=���?���ONh@Jɡv�v�`�K�H�u���i)��'�Jp��'�'�q��ِ�K~�U��n��� !����/W��7m�O��D�Oj��Iq��˟P���H4B�@ Q�S�B��˕�^��MS�l���'����R.V�;�%}�tRT�FHG
�m�ៀ��ß���H���?a��~rK #����܉t`$���#���MSL>A(��K��O��'�҈��L��8yTGA��M�c.).�7��O:���B�r�i>qGy��3���q����Tnl��sT����Y',�t�D�<a���?A����DZ-��e
�˙#_DJe�v��E�< ��f�IןE{r�O�A��I��J��k'�P-sBց)��i��'�r�'cB�'j員k��	NȌ�񶅏5��b� �f��M�޴����O�O����O�)�!�]����
@ �T��,�y����%��&��D�O��$�O4˓zv>����4��$x�M��Pf��� 2��)�7��O>�d4�ɠ~6�c?m�g�Ƅ[Y�4;1��'�hȚ7�p�<��O��d�O�@hA��O����O���L�`���Q����G@&���B`��П��������&�~�iaҕ(���Q���0�j�mZR~b&�^��v��~����"2��@���§�irA|q`��i�����O�i%�)���b:���+K�D~�B��ǯn�`���	z�6��O���O4�IPV����7G�4Q�\B�mD�C!����̘�M�q��_���F��Se��Qd-Y
J� �S.�l�� ����@H���<�ē�?����~���x레zf�	��T�h)ބ��'�j�+�y��'��'��y �G�.>�:C�":\���.q���ā uf�&����۟0'��� �R԰B&!p2�`�n�`��H�ܜ�<9��?�������n�٨5,�<D����J%�A�v�;���O���<���O���E����a�9r	,�K2F]�=J���D�O���Ob�(4�O���c�Mx��� �5�D��O����O �O����OT �U���r�F�Z����,ϕRC��SD�>����?!+O����6YQ��ӟ���j	��޸q%k�_�n���9�M������M��	��xL�~;����`�SM`�`�쑿�M����?	(OF�����ϟL��~춬�gl�9D���Z��U��� pL<�-O�����B���N�Aq ,ҐlX>+jpEc/H��ݕ'�x![�Az���O��O��8M\訧��3y��Cq�,uܐo�Kyrh��O���abУЕ'�bJ2B��2\��rP�iR�l�R�|����O�D��'�<����� .p���]3�%�f �gl^��ijBx����۟����Y*��z��% �1#$J��Mc��?��^�x,qלxR�'���O�)�i�p�\�#  �
�����$TK1O��D�O8��צ ���bl_{��H�f���"��n�ן,�������?Y����r��oQ����D	=>Զ��j�^}r���'r�'�]�Q��.=�qBd��n��y�)B4R��K<����?�J>�L� �a��X5�`@�=iIŬ+��ɟ����8�'y�iCE�k>��,�Z�
`ـ�'}�B��N�>A��?iO>I.OH0��R���W
߽5�p�2Q���5`�ɓg�>��?����S�'��&>���m�<z��r@�ހT\������M����䓾p<��)59>4�$��!2�n@J�`��]�Iӟ��'5���g&��O��)�A��d��:��Q�����'����IƺA�a�������1j7�<����64�&��~����Ԑ�̙��R�
��1�Î�s� ����`��B�	;:R��TO�x-�V���_�7��"M��Do�ʟ��I�����+���?���@<�z6�ך~���J2#_�_�a�'�x��!.��)�$���	l�8�p�l�$�Oz���N�&���	ߟd��)���ucR�d�Z�I!�V6H�Bh��؟T��۟0�1	���t�f˷>��3�gB�M���Thi��?�CT?��w�I��X\��F�D�`� �۽:)���O"��][g.�@"N�W�l�OBL�a��Tq�y�ᅩ	?l��'�~0jk67�28�'@���[��dI�g�uC�(�1{	��J!`ٵ<�Vd�6�ֱ\3l�jU��l}6m0p�T>� �kt@��@���h��p+[dUA��ݧpkܘ����X��q��[��-���Yc��q k_��Ja1"��,���WJ��d�ҽB�/�->��`��
�C���n�)Â� р��,����Dr3�̈�̈����ipoڞ
8="'�'���'�Qcf^8bLL���%?�|���WE���׋*C"�� ҿ%���T�A�'d�Y"�%b%�Ӧ��d�	P�B��-��Po��l��1R��; c��P'm�E�'�p]����?���d��>	�B��׉f���q&/���y��'��"�,�l�S��B�gD�;� �'� t#"l�0Ft���c�7����'�Xȑ3D�>�����\�D�P���O��$�0p���HƢ�,uwc��"NRIz�H�n���qn�G^� ��|����O�����b�nE�����m��T�D&A� �5"�>h �Y�𧈟�	 zl��1 �+������ ����'3"����F�O���Q!&u٪l��aѠ5�l�XR"O��Y�$�2Z��Y��Vp�i��I��HO�>y��c��q��%����8���I�����@ ���	۟���͟0�]w���'n��r����D�ѻ�B�MM����Oxu뇨��{��t���U'�������h=��E��'�R")׺H��4�I>o��� 1��8�������$UgP�%8a�X7E�v\PV�M�%���	C���'[ўt�'~ 
d��Z��#�߹���`�?D��b�⊽Gi
$�����(��]*����HO�DyB��~�X7M�6}b,�qK��k�F�C�O��D�OZ�d�Op�Hm�OT��y>�cW,Z����Pӻ:��be�� ��d"�LB�6��9� / xx�$[�k���$�ˁ��O2E0t���|\T�ck��X��M���]x�H�ck�O��$ƟzK<�&�#F|��4%�,{ �=��D�m� E0�	�c�\����@� �!��< ����+Ȍc��S�#��'��d�d}_���5Nɬ����Ot˧u1�p��<�>	�ucO�w�&}Y�#��?	���?��^bT���r��-4�􁡵�b��S�C���s#��5�Bp��T�+簢<!@H��u�dB a�/8���$�~���CPc8�Phɛ$z���UH�'�V���Fb���0���9@�O�#p����q`S'w��	Ɵ������qxPc�#tm␰�f�	AC���d[J�I|*��P�
R8 ߪ�P��`����1M�|��ڴ�?����)�1U���O��d!0�D%"���?reQe�D��1���;+
}c�9?�O�1�2�γfh݂�%R'�,�k� ױo�z�u&Z�;(b}뢙�"~�	�>�H�P��4N�*��(Xv���'���H۴}䛖�'�?�D�.*"�Q 6���NnB�����;���O���W1;؍�qM+)VljT�T�rn�l��V8cnr�$-x����HK�^��8Qr�Z=I��d�O�qqSY�����O(��O�<�O���X a��EJQ�,YNv@3&���d��#�z�+"I4��!���n�ذ��+,h�l�sd4.n���C�)��]�G+�
 #��r�?�=�tX&KS��y�Nگ>���Z��J��?�$�	��?!�iUV6ݟ�̟��'�2x���*B�����$��YX
�'��`xR$)����LL�	-|Lj�D3ғVe�IlyR����=� l`� ����iRƊ�8�@y��O����O����{�b���O��S�aF��Oz�r5ކ}T:��G*Ck���;5�'n�k)O�́�b�3AV)	)9f{��"T�'����?���@��kFǘ5N�	#�a����?1�������8ax�x�v��	GΘy)C�=(!�$Sw�"hp��E��07gNd���]y}2[�|ʰ/9��D�O�ʧ@A�4��,�18�;bHC?+d����U��?i���?���[=O����/Y8 Ro�#��0uD�Yv�ڕ,�>-�qM�zQ�����!�8e�ԏ,����B�?	ҡBO�7N� ;t(�DN�M1� ʓ0� h�I�M#��	�����K !ն*�^���KZ�$�OZ��$H� �� ����*��Ȃѫ�G�a|"�)�D݁N�x��M�z���L�'	��'��Q�'��\>	���Tݟ���,��nD2�0�A �1
(�W�ՆY���!2�5k��"�D�	�?�O81�2��, 4�e��i-
��+��LCq{���	�F|�1ǉ.E!����O�99����E�C +Ɏ4�aYr���$���,O�O ��U�� �%��/�z���Jns#�/D���b��^�)��ο{`~�s�g(�I��X���$������%t,TX ch��2F�4��.#Vm^,��˟��s�K�r �I�����ɟ�������A�\h�&@�~F�l:�!IL,�d
f�<��Iui4 S<�8�sK��E]L�	r�&Lq
�7VΘ�LX�6aҪK�!�
�z�S������?��S�'x�V��p�f��I�9�A�T;�Ҝ��g D��[�F�5x�(c��%'���3�B�HO��n~��}��f�ͫO�N����lw�!�A�S��'�r�'��U2��'��<�6���'�)H�r�:xPqk�wH�1cV��5�p>15
Thy��
J3����G18_t��+�#�p>)�����3�xU�`�Ȅ̰���[��C�0{�$ep ֔=���Y����4�pC�I./�F�PKA�,��h"ą�(\#��I���'φ57�f���D�O�˧tQ*��ddN�zY)� ��(x(�HM�
�?����?	�c�V�,�b
�8ոٱ2Ƃ��(th��a a߿swT��D�*0�<�R��1t�pP#Ö�D��׫����T$8h���)�F-0Z̄Ey�AL��?Y����ڨ0s��izh%��@�a&!�à6����ѵDwt����A6p�a|R:�dI�t��D��6\�\ ��۰T�1O���K�%��BT(��^T"s���>Q�!�䃃y������J�\��`�	��!�D�D���ؐ��$M�zP�Ԉ� o!���9����Ee�Tֈ��(��B!���:��pP�F��*���S!G!����0<�IU�ړ8�$[��6]!��0V��B���6�dE B��!�D�6 㺀qSʙ0/�ơ��G�!�Ą�4K��ӂMGu
�K$A_�2�!�dI�~h�J�ǝ� �r\1q�ݯL�!�D�W4:��`!�)(ơ���!��P2}fq�"�vhq��!�d��~Qб8�L�$�5�'M�T�!�H�N]�D��2�5��'5!�G��pqS�m5 ׎HB�	x!�dƊ7�����
Ia@�Y��li!�9r{ YB���(Q8��%D�Q�!���g���K/U�����K!�DԟwM�H�&�ՄIM�eBd���&�!�d�V���1@�Rx�bcX�{�!��^b �`��B�lXc��)Is!��QwDm`��&����"k� qb!�D's��ai�k؇P�F�yf�`!��{� b/E%{E�H;#h¥8q!�$�H�hYj��)�~q���me!�(p���f�ػ��`PAfB^U!�*D�pz!�>1L|�s�J<X^!���7���!F���r՘'/�[U!��OJ���kƄt�8�"��	Q<!�� ���DA�A���h���Ls"O�6�G�6bf�OF/5fx�'"O���C*#|ެ����U)@�I�"O�e�tWt*)�����lHsQ"O �ɴ
ӎjByX�n�!?�9�"O��b��3m�@�wn�"k�<#E�'�̵	ϙ-
���'R�Q�R	s����� \�l)h��
�'X���넏DĄږM�Y�d��O���%�^3|��0��Fś��X�N�H7�إIYv�ȓ�>ԓ�*�"]�i&E<uX0y��S������rZ�Q�'Ҵ�Q��c�
��\���d�>w�FII��X<a����N]�4 ��(a�̏}ˎ���o3�����
�?ٱ� �A ^|�0���4�
%)�4<�F�;J�n�J4�:O(H���P~_�PPq��<Ʌ�ޝ`�$*�_;zk�A7攜<Hh�
�HY�r�~���
!��<i��V&]q=��
�03���GW~��
O�v�Y`͟0n�Ɏ6h��ڷf�%_�85�r'�<&g�=�v`�&p[%$zӾ̄ƓeB���Q�׉dhjTP��"l���DL�qm�5�k��I����s��OD��
E!?y��@ܘ���
0�(����-v!���S�бC$.��f�\�Rv�����h�+d�BYk��]�\�DϺ&8���&��&l\�g~�Q��&)���د{2�H��N �0<i2A�fG~ܑEL�6r �B� ӧx�,��vK�AS��8P�_�C��Ê�PX2)Q�cu~4;
�[��!(�Wb-
��,B�"��'���X�LDzccD�R�R�%i�����L�v�P@�^�: 8��X#CD <�LݽfH��f��A��jA k��h�@ �PI0c���j/���)D�1
��	#Iz@��f�i�D ���nN�Y�rd� ����֧Ջm�!�d^�`���$1p��=�S<qDN���eԾQr�O�3p�<�A�ܼ^����,0=�< �#�d��I�mK�j�)}&� ��
�X�ax�eK�S�M�7�}��İ0�и`��E��*ܤ���׷p�"�U"�;L���'�T9O�|��'֒�e��%��x�G��3� Ȁ�Ov��2�>� ��J�4|�7l�<+���,h�H�
c}���G���j�;���*��䂅Y�>8��b��6@�e�D�Y�>Y��ⓓz��+wU�U���sӾ�d�@�a�U��Լ6T�C���dLY	�Y�F��Im�0��
�s��+ ��z~��S�q�┡UJ�S?�O�5�׎G]�a����A��=�B��,g� 7��x�Pt��D��{I�}����c`ax���d��	F��~$�]�=6^�+ ��X��tzF!V$u�x���딚F�j!��Y�'�bDPc�'�^�)$�7�i>9[�3��[�aZ�_c̔{4N+?��Ӕv7ֹk�`�6'k�U�fk��?� m����Ė$b���C�3B� 8p'@��zFl�Ȣ8,��>E�����E���C��J2�,�slT0YY@@�4^�����O��-�wdD+�y�eR+&�|��1�Cq�����8��d�?���ɷ	-�M��D�r�V�P���"�&���c'�+=�m�kJ�d�t���
�"/���ݤZ���oZ�Wv�(äL�&V�Q�vK�	����UX�0@��9�$��=v���i�i�COP�*��?R%Y����V�I3�ՎB��!8��'�+ea=�i>U��L�^��=��I�{m�4a��9�j���b1�u���f�8���M(.[��(���2C��V�հg���/p�є-N�>�j4 T@W)y ��;Y���w�V#�t䓖�o�p�)§"��D�� \�{�\�A��-+��	��CL�ÑM�?=.~�+%F
����'�\�jSB�4N��y�Hχ7�AsW��3����c��1��>�g��Y�}z�뛮=��� �!K�1
�T8�-<�yBi��f>�hR5ɍ�(����q� �HO h�0�F_�4�|�[9�����)ђI�1F�Dn�<!�͗US$8����?��T�����b�$W�%�"~n�Y��`��_��*RMU��B�I	A�LM�-Q''��T��JR���(	:8K�����p=1pk��^V^�{E]/<������xX���-S1�n6M��	�Lq�
�	����C���!��%<�P$~���8C#
(]đ�� ��I�>}��,D�x!�v�J�8�c�6D��!��3!:,xX"(N�	��TA���O�1��2�O���5	
xyb�
`9�X�6�c�̫ dJ+-�!�̈0Gh�	��noJ��$J!`y�I �~B[�h���O~qyW����I�C���;��4m�p�dΘ�0?1cD��?�'�	_�`a0�Y|( �#�	��r��'�8��G	�<A���O[h�#��v�X�b�af~	��i�h�+7�	�y
� (Y�@'��H{b���"/-d��ض���L�"����'�桳�g1F�X0q0��{�Xb�'�Va��x��4��Ƅ�R��q�韾*������;�8H�v��]��c�܍l�r��	�'E�ّ�d�lV8��˄gr�9�4{Ґ-a��i��r%͈�=e^5��G�a�y��gO���N`��g�s�(�iP�]$L9C�'���#t�'(@q���S4#y�lp쉟r]���od,eqo�EO��kS�.��)��|�6:�x���L���AeA!�^��Ҫ���OR�;�A!}R&[�V^�6��@c�탶d�8^�m�5J[;���J���<lC!�c��^���A�'�m*@A�*0BB��Z�d�ѝ'�ā �>٧��%��J�N��ū;sda�6�DA�Fe�T����}�&�W�VH<9@hN���1���#>�n�j�]����j���M�p���_��X���=J�r���J���5Y�\b�;E������`E��0?!S����?�'�D�B��X�#��	C��{:^h�� �!�Ψs�� GP@�O`-	�F�1��<�b@(g�Z�%,*��X�&f��D|�ON,He�"���i�0�Q� �#�x��blIe=>M"A� |p"�F*Ά�V�Ҷ��<i�J�l�bW�,�qqao�A��$˖�e�>0�M
ț���; H�b��,�v���%�b)�Э�Uh|�蜨L�B�
�'2��J���b��Fa\k"Ԕk�4鴰b��ic�pZ�
1�J�&+�4�"���Ne��Ƥ ���l_�t!���+�8,���'����$}˞�i4�X3�,d����G�1A0�؞Bۜ!%�S���a:D@ K��SV*,e���;�D�3TG���A�ԫ	��S��S�JL��s�☓9���x��'J�qR�y�@<!Sm�~V�25�8�����̍6�F��a�-W����Q�X�[�ay��U?l�&x��bA0B�n�I�mВ�?�bc���!����,���EߟX�Db@2F�~�	mѐn�HՃ6!N����!��=�D��E���B�9P�)�aE��|}����?a�7%��DÂk^L�t/]9w� `ÛGq$�f�I�����^HC�"�0#Q�ِ6��f�|d���'M&��&��+)X��T� >\@��/Ոv4te�T�	��-�CŻ
sB�*�KV�J}z��P�O�@��'Ũ��X\�B��
�Y�
}�1,ՎW�d,Ez"k"l.F��GЌ �b׋�ybbU�ܥ��U9k0�7	A0q�\�e�J��1�ۄ	�bX��P�*�*ᚑ�J6?�xM�O�pKĩ�Y)��c��'PT�R��'�:���K27�98�M��"Q.� ���`�ɞ&��h�	"��xO �S�LF�,^�z&�!�M��� =
����Z�TG4b 	�:&
,�'h��|
�D�#��1)�x`hfl�0(���P��"b��?����Q@^�/Z�����O9��9'��Fa*����^W<�Y���,iD�����_X��1E��S�	�@��Y9"j��6��� �@�#<!`�Jl�vL�2K�<"��h}�b
�>lԋW�"�ޥ�2�9+�!���G�|�pAj�\((���	˓��M�pM� �SF���Q]��XD'�NW$	R�O�%��(�m_n}�I��{��	c�N��*sb��m��kQ�4��$���ֹ;1_� <����HLC�h��l����=���e�b�`�E�;kI@��u`�">\�A�'��y�*�G3У��29P��&���`(�i��㊣>8``�K8/4����=�O�x�%'�Xg�Y��-�A`����  y��mrF_�%���X���L��!�3��G���[.O"=�@�3���nX�44�� �8**:0;�k��M&��U.�g�':�D��	�4�DU"��kM��'��7�|�d�BpI�+T��U�1+����|�+O@�R�ƮV
 �r	:]� |Rf�Ĕ7�>�I��R�&E� K�L}L�s��R� W�i1aC�I2����?O>���I��mХ��:���	W��%7De����/NP9C�G\�-�\�CU�Nbآ4 4lO���EH=/.`� S�fl�j&(��IQ��mڧ�~b�V�"
��,5��X:ua;Gb-��5v��[}J�i��P�6��IǶ�8��Dm�kJ�8����C<BK�A��F�u�ʨ#ԁ��@���a0��$�~�S����(O��iM�rjT" "� 1x,��߅���;`吒G�$���s�'��x�D̝O�$�1���e$��sӀ�m��%����Ê�F������O(X�~�YVQ��B�4;�pM��fX�9$v��0��*qU���W�gW��ҠL�]fX�S�;�xzrm�MJ�m�a�u���9��|�&K�0-d�!%J]�?ƈh!QJI�	I�U�r�L$����匉�����^-O���d�H�=zbd�7� ]�w�]�*)�Ȃ0���<1��~��E�j�L�:�d�S?0|��䬟��LՈ�bz(��"�L�;*`a1�'�j�S5�a�2T!���'�^��@�Z����o��d�� 9��J��d	`��	!~�KR��c0N��S�D���Pbg�� �!{6��i�$@�l����ח�OT���k�]���6
Y0f &���<��HM	EHP�+�ϹfW���g,�(}�ԕR������)�	�8N"��GI\+�@�i���[�X��\��BЯ(&�͋ �ψ����%��K���fjΜH0��*��'��,3�O�RQ��ʐ:\�<��J���`��O��Q�揍?C��
0S��M��V����G� ���#g�>w��)r��v�b?Ak��W�`��3��R�����*D��%@M�/��q١���HI��X��U�����?�$杴d���T��M>�w�@�� }��E�����#�\��$�+>�
�b��D��Q4��ai����`V�C�f��
�����<� TX)R�	�N=B!v�B#6>���I�g�:�
�l�K�I�T�^<U֊�7��N߈�B��V{d����f!�M�YD�A-6C�u���U!4�!�$Y�6��vnƅ+(t(`l4`w!�d̑�j�I�k�;%����&|!�$��Wa�A�VO�|Pa �Vq!�䊭a�U��(�-2h �V�P�bY!�$��� ���NT2���i[Fo!�D]'F��Q�YG��1؄8W!�$Iڬh�D��;T�xd��� %2�!�T�e��:�NL�@�L�A�R109!�$M�H�tMr�iÿF0�ѣ�տY8!�DćPOf�R,R�b|���.��$X!�@�it����4�^�Qg.k�!�d��de��Z�l�{��i:��:�!�HW�}b�-�T�����o�_�!�AJ�q����6i5+G��?W!��� �ni��/�,6���nK!��#+� 8�D�;l*tL�+ԣY.!�X�z%�I��/�@�|SD�T*�!�V�v��]�&m�"���|�!��8���@�${�(;�KQ�T�!�D_�7�4 #�a.Ĺ��.&�!��N�,�j0��ͩU�N�y`A͍^�!��ȱQj�"��"?,��k�x�!���B@�U/h�QB�GW"!�$B�}�TLB�eS�Y�BA�]�E�!�D��B:h�2���zH��mD	!�d@"Z|�9�2��|���,��!�P6~MV��(��/r�(sbl�s�!�J�vQ��ҀŁ�<YdMZ�@J"8!��H���)��'�� O� ��!�䇡O�	�`P�h/�)NQ$u�!���&N�8!�f�W�*'���4b�{�!�ͿIʜ<�� g	 ���U�" +�''<���A[���P���<��'�<,zd��[TT�;��Z�{�4u0�'�H�20�βZ��$sw�$!��Q��'h���cG ]��A`��b ̰��'��i�d��r�Y��Ȇ�,�x���'���"W��W�%qgǗ� |	��'��@�!�?��K�H�D`�4!
�'�X�����>�L�h7j^$R���	�'!*Il.jXV���,�mu��		�'��x#tIM�1+?8>�;�'�d��/�l���;�K@�1,p��'cx�!BE����Y��TX���'�~��f�*-�H�$��4Q8�I��'�~�Wᑈ~�ؽ�F�6L�K�'"ZŢ ��wFik�
�>�$�����!K��	f�+�@0Q7���<Y�O̭:W�u�L�EW� ��g�<��A�I���H���7rx��3iz�<i��N�$\|ŀ��R�Y��!���x�<���7x��ido�t�l��'�n�<�'���!���#�F���gMi�<�7*��@Ȃ�"]=�l�E�l�<AD�\�D�j�����6;��c�F�e�<I5�Ft���W�U|����K�<����B���
#��3�]'�o�<�P�"U-�s���)(8�����j�<ѱ'Q�tn&�aA�>sf�P"G�e�<	r�Xx�L|X�(��_��E�b��_�<١���v�5X�U�k�^�<� J\هDw ��#b��)���X�"O(��K=si�D�t,�^�T���"O�����J!c��g���ZE"Oح�g�/=@ �A�U�D|����"O�ب�R%f�2�gJ��r� �"OY�$�͝n�0�Ce��b��T)r"O@|Aa�/(J��H�-��0�(���"OV���Z�M_|��R+�g�>���"O.����ȕX���k�	J��<E{�"O��A�G���M��(��=��ړ"O��(�냄:�ЈHP��ʼ-�G"O�H�/���J�x�Oڈɲ�z�"O�� �AG�����2D�a��"O4��ᜧ@���f�;���"ON�0d�]|a��lB
	���"O���RNO2�2u�F���业"O��y4gȾB�Rd��}�A8�"Oʐs�M�a�6�"�Ci��� "O��Wɛ�M���CCX�`���"Ol�W-�"Y18(�@A+-��R�"ONMc���4"�,jc��cĨ���"O�*a���$����C��[↩;$"O|����a�@\94I?W~��S"O�\��F��2i��:#�fc"ea�"O�U�6AH*11e13�޵FX�,�C"O��e�"uߢ(���2r>^X�$"OH��GA�_�`��aW��n(� "OrM��.kk ڕ�Fb�|�j�"Ol<� g��i�H��@�U�Xta"O�eؗKX,��񐁁�N"�&�X����¯��ª�ha��QbB�Z�N�y�/��fB��{�G[�Y1�تe�@�y���vŚ� �.&Z�u"B ��>Y���y�ٌ_.����$m(�R� ��y2f��Q����!`
>$S�텨���hO����{%�5�@0W U�}~м��"O&(H�ㅑg�p���ȸ_j֬2�iR�"=E��4��uɅ�)T���	(ڐ�ȓ[V����1�t����Y�H�ȓJ�,L�t�]>�:Y	s�\&E_�y�ȓ[uz�rj$j�ɡ%`Z�(��A�ȓnӼ}R�˅�Ff�Ճ�{��|��f��ĺs�R�"`0S��-n� (���T�"��1H> ��V'm����	J<1���5QJ PR�J��,=��/�I�<d�K���	��TmZ�)Q�_�<�F�kאհ0mOd|ht�ǬE�<1p��#Iܡ c��V�"�� F�J�<9�K�M2�� ͘3
p��O�<y���$�c!��@؂�0GN�<ac�X6F��i�hQ�W���h��Q�<�QBԉc'�A�N�>�x����EN�<a�b�2�T�   D M�*�K�<�4GӒ@�"��<�2����JD�<i��`E�TrS(6Y�9�&Ɠ�dD{����2�H�P��E%X	�}Fl�<i,bB�E�^����4w�L3W�4T@B䉚3�&|SK��a.�)l�$gf��d;�2}=
9��dV�/��zŵ9wrC䉣��qv��9?|\��T#ˁUg�B�I�DV�sp	Q�g��{�C\h�B�	(`tN���偽Z9>�Ae�,GfB�	�	C�9*��	�?l��.S�@uBB�	(�z=2�-��y�ޤ�#�15�B�)� X�VL�$`hb�m�x�ɇ"O�q����fH�x�߾
�>)!�"O y�'�ؠv���b�۪J��L��"OT1��t&�P� ��O�HD�"O�!(w��*�M��ΪOj�L�"O,�#�L���ҨًlNv�0�"O�5K� ��-8���^� %"O��R��1Q�ps!/F�8`�8��"O�@S`�
� ����G��-I�m��"OX�xvD�Xf 0���V�0�ح	T"ON�K�fU�U$ht�*H�5�	"��'��$I54��7ɼ#�`aRc'ʯ_t!��P�N.�ء���x�^�0l��yX!򤖻�0��3\^6�`21�!x�!�d]��\ ��͛�_�|�ðI
v�!��
j(�K���aCG���P!����֡(�JD#�Vl��g�y�!��Z1��*���N�p9��%�� [!򤜬6:�Xr��Ž(�~�B���
q=!��WL���%&ڧ:��a"��V��Py��CP�`����Õhq��`��Y=�yrJR:*F��pAL�V�jprS���y��%$�A��k
�<�\ѓ�� �yB�\�9"E��%؛��P���y��ъ=h�����"���7�0�yB	�{�DX��+	u�RG��yҫ�	
��S��w���aq���y���t�"�@F��A-jY1F
�y q ��ECE�b��� ��M���	V���O^�|Cv�>3�:����ߺkL.�i�'z��֣��'�Υ���7_�0�
�'��!���&	�ԡ�@�Y>����'���d��l��j�L�<M�����'������F�y���<G����'���yW���/��"B��̸ ��'AY���-t(����V��$R�'3�ej���_�:��ČD�U:�K�'B I١�O�cJ���ҡ�W�`�"���8����NZ�>�6\``D̤��h1"O~]����w�˅��w��PQ�"O0�"�IÒ���:%��/��``"O$�*3��m�P����ȓj��u"O�Tp�Q�&l����,U�;���v"O�8�­�/c�X���AO�w��9�2"Of ��B��C�n��ӆ6�h��7"O$���f�ԤHunT+g�L�["OUTl�j���� M�q�v!�"Ohש�!F�� 6 ڑx�"O���sG��Y�`��D.v��#�"O���最$�|�ȦG�t����"OXf��0{o��1T��:�k�"O�a�g��%�6�pF�(Q8��"O^y�"C�&kC�\b4�ć��"W"Op����<!�"�u��M�@"OB�zuÑ3�8��゗	����"OL���@H-C�Zd�V^"�K#"O�)"Bf�>�(-��BP�*�a2�"O X����82��!��kg"O�X��@o/`yJ��5|g��A"Or�k�M��8�0�J$�q*�"Oh"��P�_Gd�AAK<]��1:3��8��	�es�U���7Ga@��*N?1�NB䉯ApU�v��e�z�ڣoN�7"0B�I�-���B�	)QlԺb��$nC�)� �\u /��}D��??��q;�"Otɤ��)S-
p��ѵ��Di�"OʔH㤛�U���!1�2���*OD=
c'YP��j�ʷ_q
�'z�a ۙv�I�c��[	��@	�'�y�ӪV��3�ν&�P�X�'��[��I<y8�j�hA=���'<t|��FN��$Er��)"��� �'��c��'�~����IC��T�<Y)�J�������4_�Tu����b�<)��Y%!FRp��ʔ�6���ɏf�<)�Є ~ ���(�ԁY�<ɕ� (X^v|R�'��[�8�!� ~�<!��.�XكO�v�6���x�<�0�
6��	���J�4�CAQp�<���� *�@ �1OK9i/�貧�v�<a#G�56�x�ȍ25�v�
�B�n�<FK�8.��)ub�3�����
LP�<�e������V/%'����j�b�<)���h�fWJS/�x�D
�]�<�T�U9A�
���M�N���+���b�<JK�#�ԙx�΄����8��UV�<�ʋ6����T�((�x��2@h�<!���mMp�J!�C�3� �$�l�<!b�ک7W�t���%"`T�5 �a�<A3�%g ٠1�
���R��a�<� ��,ۼ�1�K�!-��i���[�<YcS�=T�a	�-��Y��	p�<�4�E�;Y�Q� ���R���Aէ�u�<�`GZ�T�L4�R�4=�
�ea�s�<���	��ֽ�'���U\A�Yn�<��h�,��i��2m���l�<Q.�$<�y:AmD>��-ZP��e�<�I>N�NxC0+�(M�	z��y�<	�c٭�T4�qf�Y��L�ԣ@\�<���!x�� �GjXFEre@XY�<�DK�6��UB�ԓq���HY�<q���J|��%�H�4��Ĺ5��S�<y�%!M�y��Nӄ:�0d�C�Y�<qq�Ԕ(������?�xIQ�MW�<1SoP7-FV��aM?}����AG{�<Y��9$*R���=-����b@{�<��H���9 T���*�k�<	� j�M �O�o�=����_�<�e�R�D傸XЃ
ABb�K�"�T�<��F��C(Q���
=na�$K1.�R�<���=Xr�H�4}6`}�q�H�<�P�U��(ATL�0u�0#�Y�<Q2-U�cJ����-�.~)s4��Q�<��$'h��s%�<Ğ�Z5�^f�<q1fF�~E����Ś�J����GH]h�<T��!1�D�b��K�N���4��n�<	G ��>$gN��.�j׉�m�<1c��$e@�9Q'�	� ��s�<A'-�/�Z�#�_ƸZ҈�r�<����&U�1��E�>i�PHQI�<9��~v9c'�[78P�<��fLp�<�̚,�r��/ݵr��Y壃p�<av�Q�
����CK�W�R<J5��m�<Y �[�o����A)2�d�1ħ�f�<ᠤP��0��IȤ~�����e�a�<Y��\�J�"�� �*L٨�����[�<i`χ�O���sW�$\����1�CZ�<I"źi�ZԐ�gG�r�H�J�<� D����"�.�)R!	#B�`1P�"O̸����3���`���-eɚ�7"O0�
5"��00�⃩[�8�;E"O�5C�Ő�"�A�g:qW!3F"O(�2�c	>���`ԼL��h&"O"�
+�=!U�E�@"S� 2�D2"O�R`�V07
��ȅk (o"�x�"O>�в(��G�}0"離- R`0"O~l)"��e���8�WOZ䊑"ODU��e؟���"��NKJ�C"O^9ȰoD2W�f0;�BX�A]�9�7"O�f�Z�;ش���Х&Gܕh�"Ohd!)�=6�	��nqV�y��"O4(B�!�<^M���@S�"U�4K�"Ox���B�u���2�, �xP �r�"O�ks<��5H�F�P�5Y�"Op;VD�<:�8�`׀'A���"O����R�e	�<S�6J�}i�"Of�b�K�0h�ޙ�U�͙zG@L;""O:����J <���G6nG�2�"O8r�e�)	�8��CV:=Lqr7"O�,�SK�4Q�!�LR'W$�i��"O�4�ߟ?��@3@�[~\�"O�8x����Qi��I�	dظ��"O�e��_?&�B��!�J�V0�f"O���%2�2=( �� �
�d"O*1Y�S�}�h��aJ��(I�"O�X��NHT"X�F�$h���"O6��D��{О�)e�i.>Ԫ"Ol�S���]օʷC��u�H�4"O���#�H
j[�i�rȆ�Z�C"OH�s坵+c��EgM�	B�8�"O���,�@�>��Q�@9m<LH�3"OR�s��u��Jd�?��"E"OnDcs䝱{1�upG�+3h�K "Ol�jpn޲��@#�K�[>AZ2"O	��W�;�D)���R��QY""O�u�!fK�X{�(��@
�Q����q"Orؘ��X(3 �C����"O(�3���?T-��RIZ!w*Z�"O((oL;��0R�HH����QS"O ��D�@</H�Cg��`��}�"O��CEҜWj�)r��Y��d[%"O�ܨ1

#^\5����Wed{D"OZL��	Tn@�yWJF1J~q�U"OJ}�@ o�,;�)9q+<Dq�"O2�kYm�VA�.E�ܫG��d�!��D7 � i�#/���͉�-B!򄏡�l<�e^�n�� ̖	=!�%^*���%!�o�}Ѓ�ǀ�!���`<�p�ƪ��}�p��	�?7i!�D[9j�Lq��
3 ��1-�!�D���#t�3l�>Y)"��.<z!�źX����,�z�t؀ǟ�i !�J�g���Ü6ܢ����\��!�D���a\�1:ȁ�U��.�!�D�DZ�N/4#�<���҂/�!���+�>	�B&"g���rڮd�!�Ĝ%U���qr��>�I���δ^!�Ē�`��9���H�"�� �79!��BN��$�Ō�
s�괹��!��F)k�yA��-'
�8�'	�y�!�D� D(�UJ-;�r�Jd(�4-�!�՜I�0���P"씱8�˄|�!�� ��iA�ٙNCVp�FP5_|l�8�"O
��W��H����4#@�`�3"O�� ��� .ɾ�0��+]'Ya�"O��;ס���D\�n�m{V�a�"OR��U���
�:m�-C
	��"O�� �C7-���G��{�6���"O�h@$�Zy��1�l�&�fq� "Ox�r�+YjB� �H�d��|""O Q+"V2f$a��@-a����"O&�5��sL��,]!p� �R"Ox�XDIV^U�E%�n �"O���(O�#����}���J"O���QB�7��lz��
%����D"O šq��(����AX6Iy����"O��'�J��a�� ^v�<�3�"O0jr��
������#�R���"ODPF��>O���o�&5zDܺ"O� `�K�&<ȡ�s�G��:�HW"O�A�b�=q�\D�Ň8��0��"OZ,ɑNޏu=�<�瑳"o�`�"Od�[T��8Q���r�e[B�)""O`t�����0�K�kSPL��"O���숧F��pz$k !S�N�С"O��:A�[�i"�A��@\m1��0*On�r�ME킽 p��4�$�	�'�P	�nDU�<��6L�a��	�'.& ��Q A�ɋ
4V@`�'&}�fK��՜a�6\�����'�z��㑶~[�(Zs�0�K�'����⭉/R��[�`вd�X<��'��ª��R�岴��&WT���':0����?��ꖯ.P℈�'f�q�7"lX;V��7�l��'IFPq& F���<8a�+�, *�'kЈ5Y)��P��r�����'$��(�/I�a"���ƫ,_�`	�'�`��b��]�����
!A�T��'��QD�.Gg�)���� MV���'�X�T���I���# �xɒA��o�<�>)G䰻�J�R��"� �j�<9&���,�l��d�MF��Q�oE{�<QPpf�9 ��Bi�a�<ф��� @�����>�j@�v˞s�<�J
w  \x��b����v%q�<�b��  �3CJ��BDol�<y�f���4�S�HRT����m�j�<	�瞲!Ҫ�*LR�T���f�i�<����-z��ɒ$�G!X�.u�4cPd�<��_��L�KR��(�8���^�<)��%	� ����p��`r�M�]�<I"��#�y4@�>s
�m�� o�<Q��J��4IҺ/4Й(c-Vt�<	��71�ؐ$��h��i�S�\q�<��Q �$�Rp[�Fv1 �c�i�<��k�j�h��c� E:Reg�<A%�Y�pi"(��fQ�PP E�K�<�0*2T���d�v�D��@
�b�<����FFK�U�;!l�
���^�<QU�K?S}F��%T��Q)&D�<���&z���V	�1�����h�<��e ^�ܜ���ѡfY���7"O̓��+�5�rS�N��z�"O4�����	n�x�D�B (B�t8�"ON��㎶��ɹ0!R�656�H�"O� �sf$#���Au�ҁ'p��D"O�){�G�.��{��;!�!�0"O��aP��T���0aE�<r"��"O*=����Kj�Z�C�P����"Ob�@�%PN�`�`��NW���"O:<;�� &[�pT��A*H2��e"O��p�.ΰ~Jp��G�[+бiP"O���mK�?F|�k��ԇ{�HA"O.8#� ��bQ��B�K	cX<�"O�yY1��;_�H4�#J�+|��p�"O��X�.O�AK�m!��0E����'G&@{.��X�`���4�l���'g"�I¤Sj��|ˢ�і+���ʓ<Yp�S��2�f�1r蝚T�Ru��652@�a��byވq�ܘoΜ��ȓ�p��7^m�ޡ�A��(�*�"O�8�G��*:��0��:B` "OD`J�,����2�`Q#N4r"OH`:�O���,�h�iބc��"O���cPjptHΡh��m�p"O	�Ӫ�eOL9�b��- ��X��"ONm(0EP�jj���e�0���;p"O�=��� Q @I��M�6K%"O�2G��(h��A�7/}DT)�"O�-�A'@P �S�Ϛdy��9�"O:)���G��q2�2�@�`�'4��" o@�@|D��e
m�
�'l�P'�	"!�F���V��	�'<���"*E'[�hp��ゾTxVA��'K汢ק	�9vx���� N�H��	�'Ӵ<�G�	w�ЈS�I�t�B�'"4��iٿ}�HIq!o�Q��%��'�:A;QeW<Zi\�I ؝N����'и3"+�(�I!�*�)����'(�Bfʄ�*6�@ke����'�f�!a�ö&lA�fއ~vT\k�'�6�*&ڔwI,���ĺ���'S��;��нb�js.J�7�!��'T �0��P> zjX�ۭ|
���'$�б��	~�@�:��ǭr;�8��'y�����J�b9�G\�`���'Z�����B?L�☚�*��N�,m��'�H�*AA.o��A��j�M��1�'2���f��4,�:3�;J(�+�',�YAp`�;%g��Rr��B�� `�'��\��K�Z5<����6r�Q�'���̈́�l�x��V�X���K�';��Hr�_"S6��pӂծ^C�z�'����E��>#�0�q�.��q�'�Q�CCݰ(b^�
R��-*�H2�'����@(	���C6��S�5��'�MCn[�Y?(���kǘ��
�'2�ö&?@��$i�(Zi�ъ
�'�n؛Sb�����G�73�F�	�'�tc�]�ot)�7�]��-��'1��ӓ���i��胆�қ_C~xY�'�nѪ�"��h����E�C;0�
�'���
!S�����V/=7����'�D��7�~�ҕ�'�#2�4�p�'Lt�s�&��Cd`���'Wh�q�'�l�;��#5Ǌ�1!��T����'���C��4_�,��DµJ'f5��'	<A.�$mG_�x�DX�'j�i�d�_K�����ާ��	���� ��r``�$K�ؘS��I���@$"O0���@�� �ds�c�7��p�"O4
���=R��'A?u����"O��R���<R(Հذ+���h%"Ol|�-;.���O�2�����"OLX�Q	�S��C<p"��t"O,9�,C5I��@a�+�ZL��"O��
1fM7R�dS#,_�P���"O^l���K0A�PjD+T�?Ҥe��^�xE{��I^%�:-�#�\?C�^����ƻ7!�$��N�0����C��U( ��"m�!�dF�a�,Z��D<1)^��-�!�$
�.n���T�h��sjʽ'!��"2K��b�Իwt�U�E*ɫ*!�DX������4`V~x�%����'�����Ɛ8�\ S��H6�|RH>y���)�	�t��]Z��G ?9���D�;L�LB�I,{"�D����Gаq�0�R-j%�B�I�Z�Blk���%@�@]X ���i��B䉧|���qƀ�a|�QWC΋_[�B䉴"W����#�L9AS��ǐB���ީ!�.R�,A,��/��w*R�`F{J?�Q�N-��(s��]�#�^Yx���<���?q���?����l�����V PJ�B�H%;�!�'A�Αs�F�S=����^�5t!��l� ���5{�`x��(Ğ�!��'y
, �D��=��E@
n!��ӑx�~i�fK�2M�09��EM35!�^h�T��Gy�	s��!�d+�:Y#S��?s���
�@��!��9�>�2C�A�sPԫ��J"�!�$�!��؂�C7 =��SՌY�B�!�Ğ�F�`:��  �m�gč<�!��E�=0��Z��ԍ��wkQ��!򤗕f���h��znX�۲J�	O!�Q?J�,ذ��(_aH��R)G41!�$��b%�}i�D�z�i�-�?:R!�$�5
ūj�&�=S��5_���ȓ����o�b�f3`��\0���l���ʻcP4��rI{��$��n5|�vj�00�8����9H����(�(ā2ČX@\�0��x݅ȓJp�Q�F�&�tL1P�V/�t�� ���j!�@<f<�KnFuEb�S�B�bz�P<����B�"GnC�ɉkF$���A��B���Å�VC�	6B�� Svk#]�ٻ$��C�f@,�Rb��"m��Mj�%]6wVC�>1T���$�:E�бi M�%" :B�	�l��q�1Qw�=˄ǎ4:c�B�I+e�z{#ɓ�Q���2�f��'���?��hOzZ��t���W.\2*�X���)D�@�	�|ވщ��UB�ɧg)D�J�'�=���A�A	"���-'D�| �ܛF(��|�[��L
�LB�I�xI�0ДoZ}�z�xÄ�T�!��U�H�jN�=K�l�I%�$N!�$�@��(�G��%�=�g��
 4��)�U��us�"�2�4�Ї�Β鎰�'��4����-f �`CG�@�m��'n�҅X�R� �J�M�����'�5;�g�6�4����܆PN�'��y�'ID�(�;�M�#^��
�'���`�!F�]:rJ�<=���
��� ��Sd�X(2R��%NO� c�բ��$�O��}��"##2��;,W��P�u���ȓe|�ꊱ4  �7�N�f����ȓp5��3�,��>��&�5$p��ȓ�h����w~q�`O�.P�����0T�DJ�G5>���@H�7����_~�p�6�K?��88EM�(q[z��ȓ?���Rc�+Ym����!D�v���Iu�''f��c��'9d��F�/	�f��'������	o
 ���M�yD8Y{�'�@q'�H)ڊ8Z�Ț�p��!��'.��i�Jގ	���jѿa��M��'��q2D��Sy�Ѐ$茒1�d	��'���)��/*�x�R-I�V2vi��'��il M� �("��<Q��	�'Y�݊Ġ�:(pbJ �]&̻�'�p��D�Ua2XK�	��g$B��	�'�0ԋ���.-�|����S�rh	�'0�3`��#Q���j�H:���'[D]h�jY
���'<_�4x�'�x��O?�$�"�%N��'�n�ʂ�L�4n�k�������$�'~F��#i�}gl��',#y��ȓU�~CQd��b�A+Yt��ȓZ�2 QwbQ�q��#����ȕ�ȓy�(Lz�`�<T�fe���=E����L��K��J�]��s���8'��!�ȓxm���6�07(��� `X��ȓe��\�����P���	&Qq�X�ȓ5X���):��X$͝i�:���9�@d)D�����X�g�>ö!��P��D�)4�V�y��= ���u
l�iKC�ʁI��ـ:�zi�ȓ!�N�j"�A�>��f B:h�>���i�B�9�a�zYT���Ǎ�W����ȓQ�B����0Zn��sa_�_b��ȓ1��Q�!A�Y��bI��{Ⱥ��ȓ^�-��M�s�DyQ!��x��y���.�9��#�xQ��� �a�ȓ[ά���ȿ+CLM����;ô���()hJ5`ΌL�(�����Ar�̅�Z
@�XP�#E#0�y��EVD�ȓ6%򠢁Ł9Z(�pbN9����:3���m���F�������t�$��J�;t� �"�G��N���_� D�6�9n��*7.�48�ȓW��XK��l���8��_�t?X�ȓcA���Q^
�@�Q�*�zمȓu��1:�	�b�"d[�٥a��U�ȓr�$C7+���VpZ!�S�?B���u�nu风К��,
5hA��e��fS��Є�ݝ?/��r��M)D��ȓY<�0K�RU���؟��Іȓ[�|� ��H�*��T�K�N���@���0A &��Ю8`ڜ��E���Ԃ�g�J�JT��)y����q�Z��AF"+����٣|��D�ȓ7�WcQ�W��0#N*\7\��ȓ|�����1w���'�l��i�ȓS�$`��v1��k��P�i�x���cs*u��&��i�b�{�(�%`�L�ȓgO��%j�1a�mӄ ߚ]����ȓg��)~}���`W<!�ԙ��i�VyX�E6�DLռ�f���S�? �z�FވP��ĉvC�Q�v\ʱ"O`Hue�+����S�b�t)2"Of�Q�Hˉqq�G�{fz@!"O��i����P���3B�_C�`�"OVm3�Fd�>�p�A��+=0�"O�ɺ�@L����C�ʜ�]/V}�C"O����M�_L. :��+Or��"OxE:��_�+G>ڕ��9M�M "OXXcu��Y�x0#	`��D�"O��#g�M��ݒ7K�29���k�"O.��vn�!OG��1
��f�0�1"O��$B�4�*=����'b��"O��oK�r��u����΂��4xJ!�䃍Rx�
6����| Ӆ"hC!���'2���`�)$׀T�P���	3!�D d�TH�Wg�N��鍪$!�D�.4�h���@]�x����2I��!�� .�K��Q��EhO�>��9�'�X�񂀬�ҡadJ�7�:���'%"���G8Bv����3z�4��'�N��4�P<jϠQi�`�w�J���'Z��S͞�TW�i�0&�j6�	�'88 f)��b�x�)#j���B�'�,80�"��c�X=ۇgC+b�$��'����A�4G���[�!��o��p�'t��KcG�(�"(�F��<�̙�'`za���54#hl��M�/x�	��'ۨ9�!��-!x���䃤+�����'��DZ� �-��0��]����C�'��l0�"�w4��װ�!��'Ϛ�+�
8/�!�hU~�ze��'N�Kvi��X�v�i�+�,z�(S�'.�!A�F��ū�D��RL��'�).��}�n-�Cȹ
�����'v`� A�Z~� c#�
^\���xR�V�?���ד,��=Zज़��y���`)i��+�A�����y*:�pX��!)0֙��N��y,��6T�1`mϔVlB��pd��y��csJh��/?5:ѩ �]��yb\�J�f��d�	:�������y���$H��������s��C�I�e�qɒl;F�H�!�U"oc�B�I�X�Ҭ˳�1=T� ����vh�B��(܈��F6*�̙���QG�B�I�M�A�0'  �Y�'�ilB�I�K��T�ϵZ�-�2B�I�l�!)�4��EH˔e�
B�ɵY���P��
�U2��Y�`�6q�C��%c��ա���K�e&cEI@�C�I	��ж���>�bģ�ÂZ�C�	�V���J���D�cn<r܎C�ɣBIܭ2�(^�.�L��7aPC�	�op�5�����dl����dǷp4lC�?HȦ#��W�+L�����I�4ZC�ɏ4}49��R�����\�c�bB�Iu�<� �e�H8�&��&8B�ɾ @���(h�4xpg�!
UB�	:#�ԋeڰy��`�͈�q�C�<P���Q�~���J#I��B�Ix��`sjѲ6	|��&*H$3XlB�	1%9���vF��e�!�i�SU`���Ob�Or�}�0�-b�	�,s���&��Y��Ԇ�m�@=#���!��P�"�6�`��S�? �� ���:����N~jh P"OH�{J۩j~l!�ʳo���8V"O@���'_3V�n��"O 8����2"OX uBh`��N6�*���"O��)�C5t��@{�ᅮ4���Q'V�h�'�ў�O�$���H�YlH�K�x^(�[�'��a�Ga�6��C�	Ԥl5��K�'��r���wb}���^^@�Y�'�V1��/2�Z��m�Sshp�	�'O����eN��0��R@���{	�'���RJ&IG
�s�'L|�	�'V�D�K�m��̣S�H*���	�'��Q��\�h����&�C�Vps/O�=�����x�\;
�^�x�cPK�98TJ�y�G>D�D�!��|"|����;���J�!D�D1�G�_���r&F��`���@2?D�<a���!6�M�7��*�j��)D�lr��p�<pG�$hl2,�r�$D�LC��P�x&Q���CGc �+.D�0[�̡�N� �&��kb/'�����虛-�%��0妄� �~��"O��`�b�[Y��Z� cg~�R"O^�#Yq"$���Tk�z��{�<�nݒ#�=AW�,F�@6�[P�<�  J�o��AJ�+��`��x�<I��B�n�����5̒@l�p�<�t���̙�Bj�
��p�R*g�<!a��q���t��	d|����c�<��458�aE��^�.#6G@b�<) N@
#�0x+�,�|�d$�w�<)BD������bJ�t,�x�M~�<��PjМQ󂀁�.<�zT�ph<��dF��`K�O4H����Ƨ̙��On"~[� �N�2M�eS�B�d2�1��y�@���o��EZ��S&=��ȓ0t���	QW���`�%x�|m�ȓW�7n�EF�!Fl�$l6@���*��'i�8 aaP�d����yy ��:1Nm�V�C�/0���ȓ�|5X1�K�HȢ �6�ت"=>���Q�|-`4���B�u*��˭.��ȓp����/��%¬��CX3��ȓXLlp��ӡX	ʡy!֭K�lU��=0>͚����zfi���i�n4�ȓz�A���9˰$�R ��0[�%�ȓ2pF#��@W'j���(�+CLH��N���1g��(i��1�b�}�f��ȓW#�i�F�Z�{��S��/F�0���ė'��d��Dx̬za'F�?�����D�&�!��7R�6yړ$��:�0}r�,�}�!�dB.<�̑����T�ȁ�7	-�!��G�ڀ�v� )�[�M��!�	< ��m����(�>�s��	�!��/'��ڱ��2g�@�� �Ȟ>!�D��nU�qC�1dwb���G�|e�y��	6Iq�A�[:8����E�ͼB�	�,l������;�:6J@�a��B�	��$*��m�H\�� "�B�	�^��� ��E<��1oF�B�I�D�:��dP[�H�!�#7-hC�I�r,�����A�!LD���J�nɘ�Gr�q;��An�YzΉ�a���R�C�<5®��EM0w%�@����C䉜
��sD.��g�x����7��B�)� x�Z���"��]��!Ex�U"�"O&y@/��!�p`���݉2�N@"O�Yx�OA�$!����%pj.P�`"O,�PB�AAڇ��Ҩ�"O81#"B�GX��!$��%P��#�"O��Ԇ�(&����ҖX����"O`U ��X�"9�a�J�<T���"O�z��;v{0���ƼQ<�L*�"O T&▍C��2�mX��A`a"O�M2��R)�f�b���`e"O�T�c$��4�j�r�k���RV"ODڧ$ۼ4A����ʚ� �:���"O�����:fu�(��	o��m�"OVxbE҂tE�适ʗ\���BE"Ol�sU�� (����+[�(����"O�푣��/���CL)�Q	�"O�ͨdlx��r��ZR�I"O��D�Q���ȶf[|��-J�"O: � Qń�Ƅ�E��aӶ"OXEr"�3i$�i�Af�6s��pk�"O��BnK[�^�u�I9�l��"O��Qr��9��m�fDL�y�&,i"Oz����ר>T�Ӧ$z��I�"O��Ѩ��x�Y7#��T0F�S�"O8���'�{���S��Î^+�	��"O�h�`�LL�1� �)�@<IP"O�Q���,9����ےWZ�(D"Ot�F�.?J�4sq��u��D"O��ǣ��y�0�9�B��iRF �&"O���!�%M�0����!)M@�Yb"O,��6m���5�ۼdAv���"OR�� �\�D��B��F�]1\Q�"O��FIZ:�d��/@�)�� �"OBGj����tNӭw�~$W"O����I�Ti���M
&�h�y6"OĈrD�
�Vi�G-�l|�5 D"OF8{u/��0�5)v�N�GSp��"O�%���LX��k6�]�"O���	!;˶�*�%�A-���t"O6x���I����`2��A�u"OX��RnΗd�����S"ODD	�n��,G��!�`݌S�Z}P�"O����^d��Cb
�N�R��v"O��K���#T�zeaQ�T��D�d"O4���H�1C�Y��iX"d���f"OBP��OK�:)�Aà�����,�J�<�u��2I��0	��hy��b`�Hy��)�'|�� jt� ��0��ȝ^���{�&ݛ# S�V"@-�ǂU�(J���q�D���MI3����bpC^��ȓ-(��!PB^J2��y$`ԕ+ڈ��{�Ycn�Y9ʬ��NP�7�]��,�P=���)}`���~� Іȓ)µ�wa_J%x���I�H��ȓP���α1�
1B���3�t��BY񑔡
x%�R��_"��E��wB6���W�h�r��V�%�~ ��@l�J�Kι ��r���'D�p��fe<�1��Q�k��%���ĜF� ܇ȓ@;�x��D=ypν��eƀ,̰�ȓP�,4cF�r�|�1׆�uiP���sy2�'��	ly2��˕�L�Mb& ?o 虲�f�4\�!��0'��Db(�XK�H��� !�$Ϊfͱ�̅�|�䈀�P`�!�� r  F�Жt	���w�X�2"O��R�Ȍ4@Uh�3k��й4"O�᩠,B�G.��pa	�]��Y��'�ў"~R��/P8�L�/u<D��b�,���0>�լ��1��rЭ�:"�� �Ly�<���ЄAO��Z���&���d��I�<�s��l?z4�eȞ�dV�iA��B�<٣B�D�D��BN�&4\iG�A�<��k�넕"�,T�BäX��.N@�<�P��~d���~��ܸ��Zw�<� j�Q3T�bc+_� I��P��Ο��ʟ`$�"~2�^�c0\  B*��9��戰�y�N*N68S�i #��g���yBM�*�r�Z��Z(�*��$��7�y���sR$	(0nBAL�RĊ���y���3l��L�f�\�,�,L
�M��yB�D�kY�9��Q�$^\�r�Ʊ�yB��f�����l&l��ř9�hO���I�X��Q	���-/�-���X,d!��(��|{��{�8�W�,�!�@]=2�XB/8D_�USBK��.�!����(�8��.�`Xl`�!K��`�!��	��BE>|���`�O
H�!� D�@��@M��4s��v�'�2�)���S�D�I�R�*��i��*����O���$�'
�D�ӗM�00�єҁ>�!��>vO�����Vz�AjV��8!�D�\��#�ݾcl��Ȅ�҈N�!�$�3F:����܂i����	�Rt!�$�?I��ٱ�ڏ_Y��ʶJ��=r!�$�Q�����5YYA����#�!�dͪ=Zx��!A8?(l��a@?a!��E� �qF��N!b�q�K�,K!�d� 9���9��>r�P�[�l�!K2!�ա/�f����:U�5�TKG!�d]ff�H���~ƾ�SViю5!�Ě�W	��AFi�S�-�
b���ȓC+��p�n��+*lC���*�~��ȓIBT���Ǿix�M�d͠cVP1F{R�'�&(��$%��
�cY�M�����' X\�F/�ER�U��(Tn��'�l��Bჵ5ܒH����YN]�
�'�}h���;����UL� (J�ā	�'�8س�.4R�e1`��-�� ��'L��c��&;[�p�D�\������'���j�@Q�]�XPt��@�ZH>(O ��I�,s��'�� P���Z�*!�$X�=��c �n��S��0h!�d�_ Rq��g��v6U�E�ƤpX!�Ğ\��0���A=T�����\}P!�d�����6�ꘪ�f�n�!���-)����ΊTڸLBe��U�!�D�h�FHR�JZ�9�8�i�BG�L �'3r��7�Ʌhf��F�	�T!�K9'B�	�jk���E��F�r {��'��C䉁3`m��Q=���t�N�y�xB�IҤ+1��+#dڱ�勽sAC�^9 ���nΨ;������T C�ɺ_o⹊�؅X'bB��"��B�ɟO��4��b���t�0���}�BY��@y�'�ў�O�0��Jh1��ksƈ�R�R�'7�A*GE�I�����47Ʊ
�'e�\"�¯O���h��34pI�'i�z���L�L�сǬ#������ �C�e�)�� !�oP�v@�tp�"O� �'O3l���^2n�Р""O�AH���7�PQ'HJYh�6�|Q�@��ӧj��0��#,$m�S�K* o�B䉰c���H.P���sԪ�}��B�	� cB����D�#���ȀbO�z��C��&�^H`v��	lV��o�	�C�ɩ@�"��ՠ� �z��F��#+D�B�	:L�v�	S�w)��(P;R�B��2 �{UO��	�^Y�`M�V�B�	#|1�,;�E�>>,���/aшB��3\ܩ`l�`�(pa�%+�C��eQ�]�s�Y X� U���P�\\C�	��$K�C�U� ł�f��^�C�I�"�ͣ 
�Z��iy��F:ve�C�	�x���wa�UX�Z 	�2��C�I�5dvU�I�(Qi��6�O�T$���D����� |��j������;�""D��	�b��W�H�ďͪ=��4S�>D�Jg�:Ot9�����-����@�)D�� `�݃:�L@􏙆^�b�pC�%D����$�����
]3��ԠF!�B&��\��$*��)gbX�!�Ac.
����k�*%� o͔?pў���K
ņ	mE:�D�*'��B䉱V�a8�E�9Nֈ!��*��B�I<�RpuI�����H;��B䉼/^�e�Ԅ��`�l0�u	�'dj�s�@�5Kȕ`�DG' (�
�'�)"'�j
�1Z�K��U�3
�'�ŚgiF+�*��G�|���'�(��C�8���!/M�V�Zz�'(��x�dʴFߺ�+�M�2a�'Hd���k��|���B��܋N��h�'�`����?R�V83�t��'d
T��$@�2�JQ��H�'Y�)
eN޽	(���?��XK�'	��+�O�e�����˳u̘d�'���sFI�0?����uL�r�'�:����O��&dShNt	�'*lT��-]>A���"��>Ø)�'����3N�W��x�#/� Z}��'���35e�Cc~`24��%C ���'/<�����+w0���g��x�� �'DLq⑪�IaH��rcD�q��<��'�Pb�"�.���+�ۚ|c�x1�'��i�Bf��c����F�yJ%[�'�NU�B*L&��T�V�r^� ��'�"X"��~�42�����
�'�];P��5<�0z`ƥf/L݃�'���1V�M�x5:P�8X�P���'�c�gE(���G���d�q	�'h�q�bB�b��7�a�k�'���뷃șcݒd���O4JN,x
�'�fSa��T�9Ч�>NL:�	
�'�&4x��B�t�XtϏ�G����'ڦQcD΂#�M��Hŋ7V���"Oؠ:�V ����h��1�p��2"O�F,F�!*�颷�ڜ��7"O�5���W�����O4VP&e�5"O �p��ִx�@����{瘨h6"O��1G��~ʦu��-���"O�PA@����
Ԏ߾N��H��"Oș�d
�] ���$��n���S"O� P�c�4'Ȏ� b�
�B=K�"O�"�k�)�쨠b�Y�!6�Q"O�`�c��<E�qQ���
b>y
�"O�q����*a,�����Y�?�u"�"O\��4OҾ�\h1O��_'I�5"O��
ư}[~�u�T�j&^��3"O4��C$�u!b$ݞ	����"OD%Z��.�6L8�r��Ѱ7"O��P/J)^�ڴBI-��e�"O���2���2��ź�@ڿp���"OA���!>=����׌Y�&��b"O&@��Ǒ h�̌�$��n����c"O����0���C�S;8�j���"O��̹B�<{wBٯ_f��0"O���"a�g@�~^��"O(�@`[�E��(2�	+kh�E��"O
�J���_�F��4��"_P��Q�"O4Q���\8&(T9N���R"O���P�Y�&,�����'G~��"OjP�FΧ���Ƈ<l|�6"O���*�z�Z����0��0�"O���ŮwjԸxe�F^gҴ��"O��sR�/b�r%�ʣ'`��s�"O�-����4�����
�+QlH�"O �'*+�Tv�G+�6���"O*DK�C&}p�X7�H�*��"O�؊�CG}�2hR*�$*e`"O�D���
��U�刏�f�=AB"O �bvb�R�JӍȳG�h��"Oi�Q�(�6��$gӚs�T�*g"O���PT%]�\�qc�j��5�"O\�q��fF� 	.@hU%T��y��e���W��l)(���NW�yb�)4Fa�'�<W�mSW�Y��y�����U]4;�<dw(_��y�["XȦ�bUK��7ߺ�ba�C��y,�n����E.ؒG�Y�𥑄�y�3�D�S"ͣD!�us��X��y���0x|ZQZ�+��Bp���Q�׷�yb��(|D��"�]/V-�JG��y�+��j>`������$��<s��I��y�6'0T��ϗ�#9R�aЊ2�y��yT����n�/�����^�yr)D������)��(ͨ�(��ߎ�y�,V 4p���%�)3�
V�ybE =O��|�S��P�%k��R��y"f%F(�b�0�iʇ%�:�y�h\(���t�08�N�*�!��y���`t��!����3I�E�Ō���yBl�/p� R�
��x~��"�j��y"@�Z�h		R��4Z���R#���y�DD���Hk�U @����c�^��y����[����#��
<��\k�'�9�y��O�Ԅ��e�F���0�jA�yb��ri�=DER������y2h��>��;��W�<^l�P)���yb�?AY�QRNߘ-(�5B��X�y��Y'1��p�7V8n���N��y�]�`�:Q��|ڎIc�OP8�y�J�N��I�d�.tP�����	�yb��y�v�R�oY�sx����Y<�yß :�|��$f�o��M �S�y�kа ��ɹ�>R5*���yr��:�}rMK��|��b7�y
� R�����~���#���MG�y)C"O���[�&|�C=!��I�"OB�{D��Q�`��e֡x���"O��"�L�ef��4�8�:y�"O��*Z[���q�^�0޴�G"O��`��M#��)ŭɟ����u"O�(B@�O+t��@���<<����0"O���OYN�:t�w X��%cZ��y�iQ3��)�bKL7h�&��ΐ�y�cL~%c��8KЎ��'�ý�yR��Z]��i!4Q)	��Y�',4  g���� J�Hz�:Y��'���q�#ӆ8��[��2L��	�'�B�����7"a�d��m�0Q�
�'��	�0OX!'��-�R�$O�X�	�'ќ9bs �t�A@b�0A,$��'~��q�J�L��ZfO�<�����'������*�qau�̞4o�5��'��ұ��3+�N��D�3-r�Aj�'U(E�FT��~]�р�%x8J�'gp+0��� iE�t��`
�'P�uS��-uZV�y��G�p�j��	�'�Rq���8X6(����rO>�K	�'L��"2nP?ݰQ �gvv�2�'(H���B q����L�&o�~M��'U$h#�
�S������a!�	�'g�1+G�
'���BAO�ia#�'ŀT�f
'+ :ABUIJ���E �'�T0sU�4v�|�!eBү#d�1�'�pi� ��j30lID�Źq7"���'��-��c�,Q��{�$P���Q�'l�'$2Ѥ˦,�&� ���'.Z�С̅J��9�V��8�
�'|�,KsT�5��3.�D�gϛS�<�ą�8f��d�Ô^2�`��R�<����]OR�h���Vi%h���d�<Y�Ր_v�pp�Cх7T��)	`�<�!. :�t����<HxZ��4Ϟ[�<)���8���(�*
�T ��p [[�<��ƌ����=�|x�TŋT�<��Q��Kg�W���z��]k�<���O���q�ܖ5�z=���N�<I"�UY��ag!�"��4Z�	�s�<q�e,U�D�bDf� WYfuh�S�<�B-P(@C5b�H Lg����M�<�+S��>�;���"<�p@($C^�<u+� bv�q�t�)GQr���c�<�V�^>;�,�������p��� \�<a��[�c4��Hbڭ:�\��*r�<�m�[����(I�]�P��Do�B�<�G#N)Q�����mm�JF�<Q��˭	%b���O�>|.���$�<q˂�k��)&lQ>WJ��Z#��}�<�E)Z�C�����h�f�����U�<y��lg��F �,8�	�J�P�<���3vL����Ȓ& ��2�LGI�<� �')�b�ʄ�]b,q
�j�B�<� &]�u��̂SF���1�T��A�<��.?G@�5���DqY�I!@z�<e
�d\Dn��@�a�2�yr(ښ3�<91��.=n0����y���x�3�]�7��,��IS'�y��ܭ>	�	C��YfA�fX�y��������@��V�T�3�݈�y
� $u�E�=A��<@�#YTmHP"O��5N��>|u!���V�tP��"O,�a��]�_~@E���E.�Y1�"Obl���ʡw��ZqnM7���A"OVk�K3P�tM��#~<zS"O$��69S�9��?2G"O���*i��"�t�s`"���x�<��˅k|ne�G��~��}�x�<QҊ�:��\ٱ�ދ>�v\���H�<)���.�f��� ��H�D�G�<����*u��Ը5,�1�� ��Ai�<Q%��
)謴�R j���
b��h�<)V��5	�|г�53�VX*���o�<AɺNK�@$Iǧ|�Iz��l�<��-%��)��)�#C�8-*gE�p�<��+�F 4R� �^����3G\p�<A���7'�QSCF�8���W�<���Ҋzt�����]�
�P͊A�RG�<qW�J,Q|��$��p��գ�<�d�ӕG"�ש� a�E�"cV�<�C�ݯ��Jf��m=����GZ�<�&ǟY�}��D��*�4 �P��<�ݞG������l� ɱ�DD�<)
ɷ? ��u �x��p 	k�<�F�AB�p�/��#tf��B��j�<��H�3F&��vX�ln����@�<t�V
�����Vr���B�<i�H�BS�$�fn�>bC Y1@�Z�<��Z�F�-y(��u�YY��M�<Ac�9�0�%��+R%&�8f(LJ؞�=�a}���J�E^�B*dH���E�<A�փSI"qٕ��.+�r���NJ�<If�'հ�iiԳ7�F�I�n�P�<��A�nf��e�ƭ��}��N̓�~R�~���Ĝ1hf����F���k���K�<1J�,*���`l��h!��ǬGJ�<���[�t���K��	�l�yp�SC�<�����c�΁���X���H�<)�AL
TP�N�fĄ�E�'�ў|�' I tTq��B��U*M��'�:p3d�D�g�(�j �ԍt���	�'�"�:��)��(��v����'g04�s���Ȱ5ywA�g���p�')��`���� ��� ga2_Ɯ"
�'GtⅯ@�Z��J�[�7-JUI �&D���挙pXIJb��A܈t#��#D�0��l��=�R�,�/c�| �D�"D�0с͋��x���o/^h������'O��Y���$J�4��xi0��'J�B|� qӒC�I~4dYBW����!̃�}��D�B��<��O4�@Q3lgd���K_�jx\Z��'��'*P��kv�Y����&=�<��y��'B��	,�'^��QT�\y�[W�޶Ʊ��	2!��O������ `��O(Ԧ8��'�ў"~��O�s�ję��t_Z�Z��'5Z0��M۟'��)�i�/K"� �tL��l�r�m	���c8��o��F�����Ԑ��F\9Uh�}�'�ĉ�a� ��~��~⨚�g��P .�e�ȁR��-��>��O�����D�f`H��ŀV��ը�U����ɿRd\ �S�D�F1z�J� %O�~����?�"��9]Y�� ��i�d�T�<�f@Ihdś��T�_�ty��Oh�<ѕdȱD8�u��C�PX(U��H�<q�^+�0�� K�1�ِ&Mߺ1`��m�L��t�S�? "��b��o
�9��
-���ku"O,詡��_�`�3����U����C�'��OpE� �*qu
v֨;�~L0�O���ъ}�̊5B�* f�h�^�!�$�"骍�&&�8N��U��O�!�(qy8�@-"��䐗f�	E�!�d�5Kd�Q���X�ct��^�!�dܖ?�Հh�iڒ�!���={ar�ON�`j���T\�C�=��{R�	�<���	J?a>d���� w�:9P�)ךz�!��?���u�H�x��Hպ-�!�#x�z�L�6kA,��g�^�!�䓊;%�S4�Ɠ.h��g�/w7�'y�|�e��%�l�K&EK�?J�����y����2 �Ā�����Ԃ�<�yb���I��:.
�ܻ�
	���M+����Y�>�H�ǃI��dM!��"R
�i#�P��r����&!�d�i0]9�BX�w:8�!��U��	�'����I^?+O��a�D"L� �� �E��)�l54���7��@8@�{0a_`jF͛�A6D��hA,�rn�{���G�%�&�7D��Q�Ex��
�%�v��P��6D�|[SD�),X[BHDb�t7")D�4
A�3R�"�����H"�Q�s�,D�����/,��s　�q�`�2�&D� � �1��a�iD�N�j�Cw�"D�@���"QzR4S��5kAXeBRm"D������p4���+@CF�xSsI"D�t�C��y�⠚%�ߞ�@!�S�*�d-�OPa�`^1;��K�.�*���T"O�HY҅�#]1�\w���t^�m��"O~�0A�]+?��9	��S�R4��X�G{��閅=���B"`�5vLM�c�֩bs�<�ߓd��xgCWm���w��.? ���IJ�+�91O� ���ᕿ� ��k54�%��2��BwL�w�i�'V��?i����@	�(Kq�z�H�H�ġʲ"O,8�7i��q/2�F׫n�c3"OF(���,o� k4��V��y�"O����߯;
t:���O]�����$4\O� (t�T(D���B��BURUhg"O�P! (R�Z��b��HT
�"O�x��F�l	�	h��y�"O�r��L&'�|u)�A� Q���`"O�Z5��v.B�W@�LGt�A"O~E9��N�!�����(� -�t��	h���	D+*k�p�酁Yk���N�"e!��m�Q ��)��Y�'(V�G�!�K��m&�� B���3%�$<�a}��>�B*�6`04��"�����A�<����'5���B�cneF�^����?1�fWg�h	��b^NT����,Xz�<Y�l�x�&*���.m���r1��Z�'	���O���1�E�l1���Ύ�]O(��'��.�0��I�Jn��A�6�y�C�΂X����(O@��DL��yRo^
/~��1�S�n�I�ui��n���$L�$bn�[UIЗZ�P��%���!��.za$Jr�،���W	�!�V�8��8�A1��� � �#�����?�H?	`�dN��x� P>n�񘶤0D�p�#�	!��`�cBZ%}8>e� �,D��"0�B�y0��p�3r]M1d�.D�� ��)Ѩ�v�љ��S~8�C#��0�S�S�y�h�vܲj�X@��@7ekbC�g[h�ZU�]�.�
Q^�E��xx�'űO?�n�H��a�'>����n�.i��O�':�O��	�1�KQ�^��`#*�� 6"OH5BPk�!����#�5Zٚh���|��`~B9OL�� -ǯ^�TI�1!>t�kB�'"�'6<���)�_;h0�����@��d%��HejS���RSn�Kv.N:�B�ȓo��T�N�>:,^H���[Æ%�'��'��)�Y�:&�'aP����33����1�O�d/��>hJ�H���&�Y�@ٺ�E�'�,���p=ɀ��*E��m���Bh��cFf؞��=с���S���BU��}��T@8T�d�D&\���ز�+�l��U�r�,�È�$q>��nڸlPV���Ο��Ԡ�iU6\C���FX�6�8g��U�#k ��������Y����G:+���s�Pr�'鑞�ce��B������%m�*���9?qF%!�O�ɐ�X0���Ha�՟| "s �>���)�S͒0�A�
鲉�ta���ʙE"O�1U���m��`���vd��X�ϓ"qO�#<�Lޟ+9��y��%WR�P�*�Y<Q�֟�f�����V� %�hX�~r�E�ȓ��9LZR��d:1)�>L,D���o���B'D�,2>tݣ���;0�ְ�ȓ0�@-�qOZ�,��5��a[ 8Ol���{1��a��G� ��a���R ���ȓ&��Ljf'��9�U`kZj��`�ȓ<?��MT(�l����&&�2��ȓa�fHq�e�X����7Ț��ȓ;���3N�56�=CV�1�XĆȓ�P���	n��S�(_�fE��l������;�]81��*E
nH���<��`I\��pb5��9����ȓ2�f��%�|���+Tfƥ�ȓ��b2 �M.�:�#�	pپ0��+}��E�д\cu2�,�t���ȓl���@�\-�`� G��!8�4��ȓ�,{��?<����M��Ņȓ]8����J�X\x�d��K՚؇�Bh<y�0d߷n��5�P��9,6���R��E{CQ-v��!G�,�xT�ȓ��k�, �*8�D��s�Շ�:�}�0Iy�̄*�EJ)L�fi�ȓf����ǂ�\` ,���ʝ,�\І�&:rY�S#�7"�ԩ��^�~'PɆȓt��|i0ڶ,ji�a��?"�\��_hN�!Ƨ�
oij���^�+�̴���<8"'[�9�ڸ�(�5J�!��%Լ���B�&�8��y�HC�I����aޢ4q$�xb�O6*��C��WR̄
7�:(���F���Z��C�I�b˼�)'�˓.mF��t��"��C�I/6���e��X���HʷTp�C�n�!�ѷ]\
X`Q,�k�jC�ɅC*��q�E\)�1C�V�@C�ɪ7%8Ey��8#K�.�s3D=D������eJZ�#��3�6%���0D��"U�H�y	x��N���Kcl-D�0�O�$e�v�q&*�6�ؔ�E�+D�� +�1�8�a���S��cc)D��㓦UL�N���e>5����V�g�H���]Ux�+���/n
f��cF4�d�Y	w!,np-�a	l��m��S�? 8k��'8x�A�eʫ":~�ɴ"OL$�r����Ph�Uf�c�A0�"O�I�@L �F��d��K|�D�G"O�ik��?~ո�S�Ǝ�O~8��"O���f���:��sD�0�x��v"Of��W�~����<_�v(�g"O�uB�Ƅ�2�UY�fɎ��%��"O�8�F����Q�.��s�"O�!��C�+N �H΃�ԭ!�"O��a��A�:��2��F�8��V"OZPs��ԃQ*���bݭ&TD�p"O�x`�%��r�X%�[�94H���"O��(�ߜ��XX�o'D�4���"O��#�=Ԯm���Y�b�ԁ26"O�PqV�K�Ah���a��]��ce"O��$����A��.h��(c"OLIS�I�qĤ�QH�qh$yP"O�Q
�-�|i���r�V�O`�#�"On�K�Ƃ���lO '}�M�1"Oƽ����1/��I�.˂����'��Y���{��=w��y"tm1L�I��c��C�ɖ+Al�i��߯HJ�L뇏W�V��'��Ё�o�/�6��Ӥm��ͣ��ǇK���%7�pB䉢m�-��]��+�P{��=�F���<��кS ��'+�"��Y��3���3fn�+!8����V�2���!3�mx��1�ŭb垨�W��=	�	4�'F��\1e�G�~AP�����Ab�ɱ��	YO�zE�4��'��g��H�#/�W�|�T8�2���Cb��X^��їEN* j�]�O%܀�ƈ���X��w�� [s��E�͘o�"��!��6�{���0�+�wr�\�宆�8�uy*��j��]8��M�Y�z�C��|�&Kut�@��9�ט�X�v؀��O+e��=r�w�B�I�KxP�2%,��"ޒ����9[ �=�Ǖ�S�Z@bm�@���E�Z#H~X�2<O��A`��^,�睑;H�A�weC�m�"ʖm�*��D�S�:HS��I� ̢Dz6n]<<��*��ǲ^�f���c�%d��ͻ�ˈ �?�E�95�p��>8�� :�{��I�����+,��pz5���O��� CD4I�L1m\PU��\�nt��B�&H���3fS�&YLP�� �<t!�x�`K�;i �02��	4ȇ�	�h��1 f��w�|Ĺ�IڙBY~	��i,�7��}���yWi��=�t�1O��B0���YB�LH�.���4 3D��`ToҲ%�Q2MBŸXR5GЈB�*1["K�"�4�@�$Vp�0ԏr�f=J��/�Y��O��IR�L�)iF�l �#UM�di�ff��� ��v�'���겍�9&�-p��L	m�hP1S�W�~�~�:��c(������2�r�ҷW(0���a6��h�zD	#ϗ�}�t�
�O��	pG�Ҽ��b-4K���B�5~TdY�����!�Y�5�[�k8�P�we�:	�K��&v����ϖ�L�)��OU37��@:��_~�j�ɔ.�n�P1�'0�Ջņ;bK�/o� cs�
5i�`��"��/�\��6��12�J� &�h/L��b���m�$3Ӭ�1`�L�F�U�*��mB�^"ⵥZ��ֹ�/]���}"���!_Z��|�H�0��@�3�I!-�� #�H�8*���g%�
� ���M30�ν�B������$�B�̳1�ڝ����z^\�����!/�֘{���O�H$c��WZ\`����c\��
�2��OrTq1!�E�XťQ�׾őwJ	Q���ȗ���?T ����Z�|���X�{������
а�ɷ��	Q��Ĉg���`q���!C�^����*��.ؽZ%�"=!���Y*J�gN��b�'L��Y-�%��Jp�h���}��H��19Kd8�T�V�0����h�`�  �ㄆ�Oh�CN
x��`�JC0;Hb4�d`s�4��É���n��V	['�5!�Γ=?��XV�x��4
$�-qW.��:��cЈh����𢚒p�u����Ib�*T'�~�����[�
lH��ԁ�.Cvh@�A�ٻ(�m�&T�(Oh};�˅:�H=��S�\,���ip�����漴�`ʚ"\b����W
.���nJ���Nɔ��=��iF:�<%0�c�+�D��LJY�|�ɓ�R�@:`qD}�l@(˴@���ƞ8rr8Dk�D�&t���C&(�h����D�ơid��z\:l��v���`b�3�jm�"��Ǧ��UoWJ=1,�2Dpd�g@jX�D"8K�B;�"��c�6ĈT���M�QɓcE\<+!�� P�`�RXj#��V�+bghU��5,8�m�"	jd��R�F�S�D��X�n+����Z)fn%8m@�=���d	#
^�T{WC4T�  !Q�;;M��`�4v7��:On Aw��C�ؑ�n�k��!@�"ь�� *�↦H�8���f��n.��Q��e'xD�MC)Og਱F����,Jf�ǤL�2��DF��~B��}M���$�ֈka2`�2V��o� �aMOT�ѓ"�
4��Q�邬��d����;+��H�o��BOJȹ�$��x���@�%��g�~d{d���L^y��,�fX�R�o��FG�i�%�U�{6�j��ԸJ����KOV�41��	t�N��d�]=Z��p9u�h�� 
1�Q*w�.����,� qB���
�)�@���hc�K�Z�
q"�R;C��1��J7�ʓH�3 �Ѭ,:�4���"��Ď1�5����.$&!��X�j�����eS0���bS���-�'l��BDdP6��b�R����Ǎ�?&X�eB�-!I#�e�2AR19 +�B,4#D�4Yh��d����"�O뮄�[�2a�d , t�p���B�\X� ��3��@��d��Go����$ؼ2�(H�K����ef��ZD��s3쁀�p(ۑ+ۄEh������I���Z�9 �b�P�S-bAI��r����# �,��ju�֕9 U�f�۹38����R/x})���i����4��m���`莟*���1N��MY(�f������ ͙�%�?��ċ>B:`�;D�r�a��Y�	0-
x��x�&$�1�s1���ޔ����5iJ�=3A�N8\�=X�m���X���ܲ�@.��&��2��U�,*u%N+��+R� ����W�}�����'
��G�Ǻ����,*�^l� E�H���3�HI{�т�ŷYx���o>!����a�/-�@@�P�֛K���k��	ڼ�ˌ2�(��e�ؾ�#�ȟ,c ��
_�|HQ��OH��&X��I�6m��,��,5���ʕ�� Nx�\�V��{�.���⏬Z9�tGʦlLi�7M�;"����!��L}�L�v�Еy� �s�*�IƲ,�V`�	�#���'k�Ob0��*�P!���!b���zP�1�M�@�D�4B ��/փR 6�h��O!z�5[N
�<�DКR'�;a���H2g��6�l��pGM�e���P"�I�V���S�넑qutCA�V�0�B r�JL�A�\<y��V3ql9�L� W���k�KD�ptt	k!V�2�HR���>�U�C�F�|1���V�aF��@�\�;�f�1˓U�"���u6l�J5��mR�0cN΂R��x'c��VԸ��2��8ݴ�h� ��Z7�y�F� �2��w�hX��d�� ��!�U+ש�`��]�ĺ#3� ��v
@<@QphIpg֪*����-A�k�
�#d��uz��r�^�������BW~tq g��/����Aٟ|I�ە����Xb�I�-:�9Ӥma��ۗ���䖍[j�iۓ[A#����B%]�Y�Q�վ��g��t$0I�OZ�`��/s�D��`g"� 0B�`0#}#V�2�N�eF^�ml�`0/E�V��A+1̉)5
t��q���R� 5nv
 c�W䘅h@@K
"TRvFI:A�2`iu����G�D�P%I��&x�\ʶ��Ph�D���M�7	�n�!I�U>)��IߧR��A{�d��x�2'�U����GυS��	"�D3�OXa;4F�j\�P��,ç.j@�0`O-���A5�^�o�,H�f��l�*ۙQ����&�"�W�uz@"ϛW��X�$љ`Q>t�%��iUo�<��e� o���#fT�:�� )���	WH9�f�O0]�2eAR�Q	P��+4���� ������M#1@�{�����l2x@h@�)bM�,X�Ǒr雦-F��S�lțD�B�\
!�p��`��W���Q�DO#0�ԝ`�F,����._�%lv����[��MH	ߓY�E��n�(��`��QTL�T@�%0T(M�B ZbfH��M6Pb�e��(	��HЦ��SZT��`�5X>e��@ۏ�5�D[�В��6��+z\�a��_��O���k	7-�=	�9�?���>C��@��� '�*`*�'П=��vlé[\��C%Etɡ�n�c�:�.,����9���aw�U1��䊌|��iȢ�s�:���+�`���W���(�< ,g�B��1Tl�#��O�y�T�_�H�R��r��!X�j�s*�$5l$���ݏ
)xݪU�V�:��]b�F��U@��,P~Ն�I�aND�� �b �S3�ĀL���ɗh4-k�$ bL|Cb�k>9C��Y�&bAf%;�b߈T,ܴh��!}9�<�q��|��h��-,Op<Qr��.��cA�DBS�ĩ�,�%|/�t�'�4M��)T�
(�
P��K�/tHY�4a�DZ���r�'~)�d�ڴk�,��J;�D]r�¨u*� �끼1A���?��;x|b��4jO�U�Xb�O@�髓+�5�.5�ѥS�I�.��Ҩ�='��S�)R"U*����C8-� �c�4�(9��œ<H�(���X?�	*4��@bΏa�f�`��S�C<Э
0#,��x&o�O8�*�]�4��P0"��`�b�hЄӪB=��݂/w����#�;�b��&ϵ#J%�ɉJ8��cP�W�'a�|���B�'�������O��Ar���-G����K����d@�":�����ШA��y��H*H���E���`Y�US}�� 2ÿU/BT�IADcayRL�|�L���� *�����N�W-�I0�-<�fى��/��PQ�b1��DV*̀����P!�y �	�%=R,���ٽSȵ�"���+�qOX|��̕�Q�>��0B�/��� N��J�^M9%�r��b�k�����C�c���J䡔� �pM��̭:H.�Fn��"~Γ3�8���_�?W8��V�5�h�.�8I��5��eS�l��M�7�4��ԙ��`��y�����jD�QY��P�FcU��~rC�9���0��6�uF�B#H�]y�fX��9��\s�8P@r��m��(1a2J��A	��!M�AA���
�MKf)}ݝ�$!т#�-c�����^�~�����:<��Ҋ�D�6xg���cy1j���_Y���$��`�9 ��7���$H�*{B���@H���rQy��@���.0��� (��T?1��>N�C#DN1XB���G1�d�`�����b�B3�#�I7co��q�뉛y)�4J�C�T���B^���%ɥ(�m���I< ,�S��ے]��S�O�ҵ�qI�YP"H8rc�g��Ę�g������e�B�"4,1�zzʝ�����٦=7��ͻ(�H����w�RId �O��O�
��@���<1%�,mԨ�k �E��E��FW�cRB�i��!�Y��$�z�K�3,�jI��m�/$�M�=���:`�t;�ㄸp4�3�b
[X���&��t�r0�NĖ5���p�*b	Z�KdD�t8������Rr�j6��9AL��z��_Z���h�U2Dؐ�އ<�p`��B>�d=~�ɘEĿw�*��
���@GY�)WN�;�gѨ|����ЄT�1�G�R��ȓ7�¹�HV�gle�ĉb���(#�]�i�t=�A��0R�Z�`6���1�ҥ�6�|*A�3u?�N�7jc��ːa9��X�R3B!�Z�zlB �w*F?ȎIɠꇂ,5��GfE3y�f��3Lؕ�z$�"c��xiL ��jǛ;���������Uh�(��0��!e�&<O�YH�ȋ�4��l��+��@7`��Z�];���8t.<�Q�
w�P�ժP7'�f�[��'@ԁ`�,�ki�8��CC�q�ഒJ>��#C2s�b��G��5���O�6 K���+DЅ`ĥ@%P�x�*2�+!*�q������y
� t����N� 1�j�E��"�>��T��I���0�)&^�)�ҫOxd�����}�D$�S��杭6�*��a+�-48cL��TΒO6<s5���O�x� �P/fN���@|��z2�N6#r��q�(]	&6-�=PL���6�Π]?"�KA�8���η w ��`�&	CR�B���/!�x�yB/.2e���dU(&���R��$����'��a��M�Ca��q��A�A�h���\*��Df��5/�4�'��y�Ow�q)O�)�L�fEB���>Y ����Q��I�x�\�a�*���H���-J�X����%[�Y�RJ�˟�	ׅ�?�|M�&�ƛ_/��(���p]����mW�l�b�ѵ�
�~���74T:}:���(l�\�PV��_�&A�ҥ�����D�`������50\*]�B(�u�"�,�l)Üw�*I�U��;	۞�*P.	9m�Kd@��䗀vA8�)3DXc��{r�҅^�nt*R�P5xU'Q)�r��#
G$ 1qQ�Gе0r���o�;�zXB�c�0pA#c�-�l����'!\�xz�$\�Ϭ��woM ��`sS%M&5L�Fy�\!Ǹ�؇�L#��tC�̤0ڐ�ї�?�(u��l�>
��bmH�y�����S�k��A��+-ӊ�ѷ >�,e�,�;���D��@�w��0^gZQ�o�g����'�Ƞ��o�	� 	�Ԛk��pK�)/��M�P�S�V��F%M>w2`B�G�"����&F�;S��[G�V"j A��A�kd\�E�~��~B��:/R0l���&u��

�N���Ń'y�X�a�5k�x��+T�)^$L�W�	 a#0����y� 5[���!E���8�۷�ȧ
4Y��	��Qlh8�A�:{ǚ\b�g�'6A��)K4�2v)� '�BDq�@��� @�Ꭱa��<p2�q�+�)
 1�,r���%�\tY�l ���4xCE�{�X1��mT##�|��f��9_Ѐ�w�s�'��A�F��h.EC�gY�+aT�C��<e��CfAF�9x�����j��֠Y?a|X���-���q]<g ��sv�F$>r�����?���D{���1�gD&r�N�il+}rF�N��"�蘗p�h����57l����+5��Ea��'u��Џ��� ��ʮ�xg���s����g�������%w�?U�# �w�
��t���W�����a��y5(� qnN�8�nR���+0��#������!����;ZV�����rU�H!���F=$�i��;{ɬdA�e���;DCٺK���ݩH���j6`�$I	�Ѱ$�� &K҄�d(J�d�\����I�X҄M�I���r M��uW�a� 	�*"/J�!���	 żT�X9S���5$�-<ڕD~�
�y�ȝn�Q@�)���J�cJ�!{�� }��-�sd0� ��ٲe���k_�>CQIc!dC�vG]�}��!�cT>�QaG�K|n��eb�a;d9�*��ŎW	R����P�e�F\�Q��r̩a@�� @j�a��eQ?i�m���n8�&j]��Y��+!�&tlX�ૐ	��� v�8}R��!���	�z�&����c�p�c�oGUٓ&O-Ĉ5m��(�Q�b�#ը�!��1��OL�);�&%`$��'W`\��'�JpRUE:"GX"�!@�_�(�����A*��"eSd�O�([�k��Dx�h��!g�����I�^�ڠy欟:e������$D:#Ni��i�uB�7@ڃ�y2��%#~Xq�Y	{�~�[�\+��Qb �����O�"~�	�7�x��{��dA�Z��|C�I�z*�h"�M�
��H%C�5&2˓I,`c5lO\u��IH�h%jSǁ�AM>{u"O�@	�B �BF1c��##�87"O�@�%��/��Ӏ�(CR"O��CC��G�d�@���V=���"OD��*�,@A��UO	�+^DA��"O|� �!W��`	�ΞpC�B�"O& �s��'C���3pÍ� ��I�"O���p΍8kI��y�%M�J��I�"O�i��Uy�!�vi;�0�B�"O���Ǩ� ��iR�)�[U�Yr�"O��� %��Ra
#fʒC�hi��"O��¢nUH��Z�%	_�R ڦ"O4<��KI�]�N���ܛta����"O�hP�c��<��c]�_�%#�"O�e"e�6.�U��9/<��q"O&�
�h��2@8\'>�B%"OZ(K��ħY@���d S�.'�a)�"O:P��"�,f#и����(���"O, ��Ȇ<G��`��/T����D"OT�A��r`kql��O�2 �"OLD���%I�H1��aƧZ�����"O�����O@�m Ǡ��AS$�+V"O��`6���� ����&@8��a"O.�3p���$g���CY�ycP-�"O`䩀�H�Kj���኶z��'"O��U�ܒKf���K[���CV"O܀�`T0�|x)�W�
�"O� x{�"̈�H�c��Y�"�13"O�H�-!��!�m4�f!�!"O�|ի��`���XĖHٚe��"OX��p'E�;�@�Q2@�.?��l�!"O�-�Ixi��:0ԃ
�nD�"O��+Qm�&w�p��_���� "O�ђ�f�7�F�
%�{�pJ�"O<�($�F�-n!��cL|TJ��"O�q�tE½0�p�z �/G�5"�"Ov�C ���
$�]r���F,Hap�"O��km�FWBD� ,�34��#"O&1`�kH?��]��J(9��)7"O$�F Y�O�n-◀��u�,�8�"ON�ʂ'D(	���U�F�t�1��"O�Iz��?���i�Bi�N�@�"O��䮕��M0�R�e��,�7�7D�DC� �4���3��)<�1���4D�(�u�O�I|ѐÄvz�	D%1D���G���d��NT�HT!W�,D��yAՎl�A'��}0�@�'D���/���@�
,Ej Z�H"D�L�������WŃ�Q>a�Ӏ D�RE@\�q�(��LL���	#=D�L�lF�j�&t�K�<D�U���8<O$p	$�4�����Y��e�`LX�R1L9LH��S�B�V�G%2I���3?�4��O2l��߫f}a�'k���b'˭J]M򃠕�uN2��
ڵDQ�_ed��μ`=
�;��  �yB��&n��+�Cо
�>�G��y��ъ]ʨ��F�H&�h�Fh<��>�f(˼s���` 3d��1��-Մq���Y�D�j cFL�:�P˓9®1 ���1|H�"<��k=2�xɪ5M67R��R,�s�'��u�e-^�d�j�ڦ��*_|I9���k���
|����լ'�z�MN;gx�}��G~RZ��d�Ǡ���I�/P�9i�lC�j�p�0葮mC����e��>��O����ĉ,W�-I�,C���͖:

x�����Z�҄[��v�<"F�b�Z�q�F�Rt���+4%;p���>�|�p�Ǎ,�JMCR�F/c�\�I�V|�Բ�����&=_�h�Ŏzt|5�'dE�Գ�<%�<dÐKʂ7�^C��(.�V����ЩZ��%@�	1�z��"�'8��U� 1�D4 ��|�{�F�++D��UW��~4��A��O8dʔm̠RN��C+C-.�(FC&O�� j�`��V���Sn��R�HMscA��}Q���޿:��mkU.��p=1$&��F��t3@��4 �=�E
Ba�D+�i	�Ze�����[P�|f	5G��x0�5�5D2v���H�n���:D:�Y�ȓ/������:L� ӈ ���"�p��lI�Jᶐ���ӈ���ܦ)i���P:PJ�`�����E�uw`�CK�;Moԅb��B]`8Jg'&,Oڤ#�H��8���(4�#i�!�D��"q��KF�F3	pt���Iv�-rA��;g`(Ӡ'��&c��4'آw��c&����T����5�B}1
�qa^����S��*I��=9N�.�r4(c�v���ԯ�&��&�@�N���ʁ�z���YAӸm.~}XĪ�^���ʘYy�!ѫ�p����%���^�"@�H�FbI> �mQf&؂i���`��
�l,��;q��ge�1��ߌ'J�h��B�<
�Mi6��k��\��b�*F���ፆ\j�)慉�+,r�m2��2ˏ���g��Fѡt`ӌ+���@�>l��ԝH ���Z=���3v�`���K4՘�A�?	,p�۱cƋ�Jͩe�D!�X�袂ٿ��{��ی^\4QrN�/(џ�2l��l4te@�D�Y�LL�anۯY4�� e	�@���%i%����cȍU�ĠX�遈X�BP��X4��p��
D���U�ǆEَ}��&N.3���a��#k��I��#n�4PY#g\�h��$��03,��A؂6W
�X�'P[��aaG��"�HE��6|&�PU��y,�"a� 5R �p��ҌQ_��I1�-#�PsJR�ف%�̆+�::��eͩC��ܪ!���r�oZ�Ү�q�(О^9�L���up��!͊�QF�����S�C�8�B�ꉍ7V��H���	h4�dӮ���(Ӆ�
BA����&]�'\fH�h�g�q(e�[ "�:��4 *}+1��!�HtTĒ&yb��*�bQ��X��
�4�uǉޘ,����٬c>f��@��ms����֑���ZFc�w��>�'��x�|5�q��F'���.����a�.�%q�n��<�0���W.(��rL�A%����0
��qղiS�z�HD�>LH8�0��T<�<+Ç�+9�0ř��D�&:�� ���hTQf�o����t���<X�eC$
��0T��9x�,Qc�_6>q�*��@��$��'��$1*|�գR%��4(+��<s� �c�Z<*y�@C��3!ˇJ �@��P:Б���7�\�T����y̓<P��&�� ��V��*� \x��F�-[�	���Ԗ!�����%�t�2�>�Xy)��^(z�<�b��(P�%�S��IpO�=]�����`��v(�CSX���_%�$�d����I`H�+p%H̓t`߄I"T� '����R8��azூ���<1e-D�g���*�	��d�����I
V�R�9�H�,S��k�*);��q坟�2�u�'�%��� �]9V�Q_D�p'��p���+#���aT��Dۃs��n:xb2�Ӣ,�"��\c0�5@�4�Ç&9*Ǡ�WG�	*���
7Uj��袩�xrH��R�iy��˧I���y�b˯{��[E0��`�$��F��Eb��gf�sr U�[p��(@hE�Y/��!�f\1$N����P��U"�dc�!� ՜]��x�(�_"� ���4N�2) gGƿ�J�H��Y"9İT��i ut�a��ȟ�]�/�2A�����N
A��c��(�B\�UՊ����$o��{A����	Cu�
)�L@�F�:ӓ#;t�D}s"�%�|��g�><*�K�4^��CQ
F�)t��ІC�8F���S3�]���4(l��@�_+P��h��Z�=ohl����
����¥"�&�*�k�?�6�"(��[%bPlӭt��̡S�/%�&Dڵ �<�B/O�$�P�W�G�֝�?`q2q˷*��d�s�@�a��l������L�M9�XV���;j}*!�˵/��P���A�d��X�qC���^$*�Z�g�|}����\��-���Ġf'�Yh�O^qC�#]C�DT���OU�4�5P8�8�MDLM|��5���C�\U#��B�L ɔDV/Z]�bT(ԶU2�0��D�KFv��w�bE��폩`l��;�具G$�� ��)����Fظ"Z\ҧ������"Y'^�� ���X�����������X�AQkT�=�T�A�+�)�P���R��#�����2�Y�M3��� ���EXG��M!���s�˰�jm�bF�&d��Uha��{6�����(g�pZ6�ۆ��)�M��x̙'�]+(�ؔ�UJL$$�D�Hz�ȑ���^��,ir�,ғpu"Q��*�%��h�E9L��Ig��=��,9��+_��$�X$qv*E���ȑ&��t��P8N��]"''S���2��]�,��̓��9`Gq��((G�5�2�'w�X��n�,$�w'X#o�%@$ggjT����"~u�	�&�i����lM���DO3@�*c�8�r��@���-��^�%@��'�|�C� ��4�3���C`|ق�$Z�]u.�`D���9���D&�,JO����G@�u�CiL�@epź��ZY:�(�@ڇ�?�G'Y8}�n]����(�pvG�|�'v ���9y�~}�F�ß�8�0�G�>��kdf���4�Q�f�0��Al��韰aA���;�f�Z�'D�:�bT72�d��#�)�~	j�4^�P�҆bG�)�jlbeB٭E"����+h-r4�r/�$����/b�9���5��ʰ*T$���k4�P#)�:ą�I��z��$��[D@�P�h��&ڀ�p��4@p�5��e�^�)Bm�|��`�%�BAǈu?a���]0����bN����S@X�n�8UZp�V�}s�ٙ��������lզ�|d�ׇ^@~e!0	�-�LY�щF�~x��E}-��Ph�ǃ�yA ���k��y��_!q>���'6�U�"jx����3�_Ert�r���6)�T�	�,(�.X��
�� 1.u� �[t�>$���iWZ	7 �e��T��*�8�!@��Z��L���e�Z��gG � �h+�CV��ƀ���Ԋ|{ `0��4%7|E�`o�2X���*[2\9�+��G[���u��^��{���]�fxȕ��}ڴ���ƈ���Xs��%q�b<�'��,f�P���5fVnlZ����}߾���FH���|#%�'t�z����PQ���:M�ӌ����\B�ɘJˊ�ҎU&>x��' ���,Y�&�By��سv�ֹ@���D|��	g�Y.%�	7�܈r�$k�G[rr�]�rB��r�g��1G{��� i�
�<8��2Ԩ�$��+a��g����(A���1�,uP�'�\9RԎW��#�J��D�[�\��|K�F+�>�X+�O����]~�� #���RT �Óp^�����;!���Pg�+���d��	x�͇=�\-x��,[N\HfN�Z�`��q���BEŇdclU	��Om�0�R��``v�UX�HyPe 7�8)�`�/Ҧ��te�7���8V,OO���1��+HR�Ma#܌a���!�d�?޴���%��3����i%�����UX�T`�{ �Cq��)ΰ@�ł��0�Jf	 G�&T�ҟ̸P��1Lo>!�>))Q0A�5.�\���� ���r��E���'l89"�P�(*] a��~�e���q"�.��i��GU
(YX,JF�޲+X�2���NxR����Ţe��	�Qb�.��a��g�
)[Z �;���3�L=D�ht�Љm�t���0�ȑ���%Fz���M���O�-W�;��:@+V*f���$��qt��˱�Z,�x�2��?M��t�[�
��W�a�ԋ�o��u}&��`��ʝ����9S�P�nӬ�
��dU-q��)�T��\�����L<d 9ĕ�S�Ö��>z,��ّ�F�!CX����m���g"3|)b�5���ɒt�vN����8xu����
=8�(��7צg��S��?S��Ջ�̓�������B(mc�c
��b��3�0H~�S4s4�pR�����?E��'P!4��"EJ3d�\
.�&YB^>��SO� ��2�Ŗz�:#�b 8��O�"Ub�wST��P_(������B�1�'���r1�%a���hUJi�'��#���'g(�q�HM����;u��Er�B&S�����	�M���h[�d/�i:�47�>�'B�[D�ӎH�yö��=�p&�t�>倌�D�ET�st�����c҄�u��*CdI2U����Hg�O%�ܑjTa�&P�8(���*ڃ�ɡu�YȵY��(c����(� `U hҰ	� �.�&����ӯ7	>u��e͗X�TL
H,�R��s١F�}����Dǟ�8���1S�d�	�xBr�aa�#	��S�O!hd �J�0*(�C��3��ZT��V���K�"18wD���/FpL@�����i�!�1�;/�����)~X@1�d�t�v��O���B@���<Q������d��pWP`�$˽D��uY1�	)H<rUY�M���m���´�����'�RP9�	T�j1��f�,f�!���j�"�匫^3��J�TX!B���8�_�m�C�a�^�1Ė	���P�Q�>�"��D�m�(�±�F�MQ ��4�F^�'��TXs)��4��#m^$_:p�p7iˆ0�<��A«<���y1��5I��P��*/]H�s D�`���  �ݚ��S�4� ᧮_�CV6C���,hy:�s�*@�{��=0$��2�өE􉣟w{�uk��ք*'��r�ɪr�V���'�^<�ul�6G� ������$����!�Z�|es�����Y�+]-(�-�l�4B����� 8��t.R�>��m��,	
n��It�'��}�,j���y4샨N�lux�غ0!�+���Y��kֆ���k��ѹ����ד6�fLa�Yk��E�r��|$����M�q��`X��7�A���uU��`�H��4�dL1��F�aÆ(�dkت@V� 瀝t�<A�C��KN����"�ܥ�v���&=N,���;H*(z�)+h���JL�ӻU����w�h��VEP�R����sě;XQ�X O>�c�;�E�I�=����c�%1�u�ƦS<?��mY��ߛ=6b�IrcǦ}�ק:,/��C�'ƭ?Mh��`���di�nߚ?2�%C6 ����uV�Q���2e�Q� � �8;YЁ	 ���d��={v.�/O�  ��
%`<��0��E�����T�K�0��D*�cʌkX��N.�����R�i>Ia��D�F>�a����|��3?9����)��/Y�*��h�� �4�!��^�l�i��x�敩�Q�=��96`�$�~���l�{���#kߑ`�@r �O?���^�6X��Q�(k)�p¦(św"�Q(s �����&�O'k�J�Y�_�2T��q���	ڠd�[ 	�!��a۷I�J�ǧV�o��ضU�Ԃ�?:�|lX+�qO�	�p.�Qk\�d�M�"����G��my�F��H�,T��I�`l��� �TfF����C�O�,��!F���Q��0;F�jB�W%<� R�DY�o"02���)�(OJ�J2��':�2dD�0i2bS�J'Q6r����G/:��Ȼ�C?*�XB�#�(j��S�ȾO<���Ү$P6v�����/8������˿��d���=cD=Rd��D�Z���c����;7���2s!��?��h��g*B��#(��2nX���5_|���M0 �	1,�J�li���ؐ2���cS�d�jV�z��	���O�Z�eK�xa�h� �H0b5���P�O�@P��g&�<k��M	��<"D�ʝ|f�d� ���`3����:�<M�f8xs�4#f��13�H�o�_jp��G�N1flPa㣛�P�����S�\o���_D�^�@��,dEb=(��Y���y`Tn�2]*�
��� 7Ê���ބ@�P�`��R�"S�d�^��� Ș\=�q	`ɚ�%�����)3���#�W�'�����FLx`&!�B��Њ]�M�^1r�m�
$�y�q �.��A���T!R��ұ0�! �,��m�t"T��8�!��ӻ[��5�^�v2���cmS_���'�`���'-��YG�;%6��un�_~�M�Bks����Q��7H����YZH\�����(�(S��ӄa�%ĄY�*�q�#��E?i@���?G�TbFg�	T�Q��:a���SdH$esF���%��'*ީ+����;@�Dzf7��I�"]��[��_p�^���f^�khѤE�<G��	)7�.a�����AHS�կ���O�$"F�ч�4u��6D�N�P*��b�iX��S&M��pc�D1�,2v��0}�\w��Sᬃ� ���*�HSg𨅀��Ղ�T��0
S�~�$�XF�H�'��(�J�Ħ��W��gh�ab��\�K�2� �������_'��ٛ���0E�������^g�E`���M�6�`dX�~�响#�ⅈ'͆�ܠ8`t��M9v�?�7b^�} |� Q�{0��U�+xڐh��F.u�P�/D�
Wȹ��I7L�t�����&�H4�P��;�H���iHTHx��W3qb�B��Ë>J�'g�̈��ǟ�Z M	�	��>Mr�*�z�)��J��������Y���.3�`@�0�_8|������DӟH�R�AV+U� K��cS�L�	�d�V����Tz�MG�;�1����	v�ݨ�'Ѳ�pS	�'^���#��OB:��B+��q��^7
�`k玪M��p�~�R���2R�S7z�t�
��Tx�<bA�]�ֽB��.Y�^|��ʴ! ��e�Uʼ�O?��ń&��p���ܠ�Z�+�!�dJH�&��r�\(�nU!
�4l��5r[�ĲE�':QJ��5�a��
Ue�L�	�' 8;�i�7m��q�Ռ�-D���:�'�bm1�%^�Z��;�C��U��P�'���ZGg�0�dBX4F���'��`��8d.X�Kƾ_*�;�'a:�zvJ�@ʎy[E�E�Q�Pi�	�'�$-��nȷ�q����Nբ��	�'c���'�ޛS4�]�F���8��[	�'�j�0��	e*�eAvmV
DĜM��' �A�5n�9J�D�ҀY)U��5��'%Y;R*@5p��V�K���'5*q�Ɓ��x���.N��{�'ru����>93�+��,+ T0�'Q���dW�~V��S��$��,H�'�<D��E��1��YӢ�\�w3��[�'��X��k�L�1ė�cn�� �'w�)�.<a�Ը�VꉿQ��;�'e���@�X�%֤HUŔ:Rܨ��	�'�u�M�4<��`��ױJ�P�	�'���?rƜJR&�)Eܜ�	�'Y$�[1��$;��a�Q�X�?�xH�'� �'%�$|�q��Հ&����'���{C�:7L*�*E?�^�
��� �=sd�7]!C�C��L�e"O��K�˙�d!���UJ�
'L*��""O�1R��ث�vY��AL#0��"O.-�E�޹x.����̚='�i��"OJL��A*_9f�!�sL��W"O<	c�D"�d�kݬR�.ub"O�չt䐼X�Q��:0�iٵ9O��@a����{�[Z������8W<6�p�͏�6Ÿ�D��]"�{�CC�w��l�<%>i�a!� ]�6@�'C��% w�Z����� �J4̙;4)��M���=��(G�ƹ�0|Z�ܙ¤%: H��t��SK��M3#c�4Dm��s{h���_y�O������X���3�J�|���	���L[r���Ό�3�V���Ȏ�0|b�ӿ�bDɳ۱M�82#��F�2�c�<ڲ��ȣ!2�ͅᓤ |RXs`�¥r�MZD�����L�ŵG(X"'Θ$E�ʜ�k-����Ռ�9f��m�7=�����\�J�K�A��x�C�Y>*�a����	{�i��S��(Y7LRT�2���߆H�:���O��ᓙF�|�+��&An�@���a���=Y�0�?牠^�@5�׭d��Pg�ٶ`�jO�ñ�H�<�b���D�F�d��-P�lUBeI҉()5�Ec�(WX�
�4J�.M2�'5du���(�'����=��(����l�,Ĺ�D^,�?Ѳ�����f�[I��R
�',�jpR!�R>�d��hM�pF�����O(�[!lV�Z���	M�'���>S�ͻ��֦^\@�Z0�<,�R6 9y�T�ҬO^�ˢ*%�'�N�]Jt�͉ra�u�Д��>gx!�Tg�>y��� 0���0��OX29�B�F3O�����V|�O��s�$�0O�����h�OY07�@<�����u��	�<E�@�K�<>�P���p���)�'W��c�f�� �7lO�Tl*��geɻa14U`��M��҆�I>�M�_�E��X5Barh�d%B!p�0���?)�JW ��)�5 ���8�̀	THBEI&�.� \P�Ο�H�d#��"�O#�DcddU�+��[$mQ#[D��#B���n��s�MS��Vy ��j����f*�9p����J�i'�-��'�����^ ,N��fB�r�ϥOu*jE��JJoB�d 7�Q
	mV��'`�1���8F(&�Q��9OY����	����Z�3|��	�"O�i��O	�d̜���0T�<�"O&��7�N{9J1��m�gm.�"Oz��F+���j��*d�0Ӈ"O�@3�	uQ���;0ǂ�8P"Of�
��@OZ�T��J�´"O`���@�M��BR�+�Y��"OĈ�%h�xpi���Ă�d�"O�-�`D-��|Qf@J�^�x"O2*2��#A�̼z�	�u(i��"O�(��KƉ>RxEP�ko�a�Q"O H��N8�Ȅ�u)WsQp�Q&"O(�K��D�.���H�t�4��"O}I�o�?i/�Y˒���j�A�"OF����
Z:x��q�M�p���6"On<�u�JJ�`��R�H��$�� "O���@��Li���O]$(.t�&"O@D��l�-d��ٸ�`��?/�+�"O6�`��c2��r2��7(t��%"O��w.̉]����n��U�J�"O��9���5s����4-��f8�I
s"O,D�Մ��Qj�q�,WI�*���"OMj� *3?�㦡�M�̠{�"O�i�g�{@�%kg D�HP�"O��pAcؖ*Ұ�xRO8�&2G"O�P���
?�:��1X&f!��"O����#ަ81VA3E��0�&�
�"O���� ��8
���0�M���2%"O�c�P;>�6,����~��Y)�"O��Sff�=_�FK���@�V�2""OZP�di��
:x�8��-^N|��"O�9sfLU�l982DÃ4H���"O:�k��֕<jĔb��ǄJ߸��u"O恁���$K>�=[功�~���c"O� T�Ұ�K2C(�Q�	�e���(`"O��"�lC3	�A ��Jg.4��"Ox��&��N���@���^t5Q"O&��T�-�h|��AĝK"Vٴ"O���b�U��pӳ�ʳ	�I�"O8A2�Z<-1� ��`�5�U"O4��!�X8>��Y%ݛ%1��8�"O�M���	�� x�U;m�a"Oƅ�BџX~+
� 4	~��3"O�!��B	m��B��z�t�s"O��y�lŗ'6ت3oʄJ`F�0!"O&�����6Q�`�^XWT��"O.�+@a� 4�]�SM�:H0-�U"O��"%��6`�e���(K���"O���*�O����r��{��L��"O>�B뚹�q�q�K
j�졩c"O�RB��3����֫Fs���"O&� �Y�b����t'ىP��ə�"O����D���<��f^u{�(RE"O��	sP�/��ePr�����D"O&���*��j��l��$i��IھAc!�$��\��Eb ������m!��J:
X�<��	����b��ȯQ!�8S@��J6(ɐ@h@ �'�Ac6!�D֙lb�1�"͘�	�ry:���("!�Ď"r����f�r��i!�䊘�\9�W!:�R|��!�$l�!��Q�nYn�:�)�z���z� E�!���Jr�1�k�W�f|b��۝v�!������!�銀j���:Vn'�!�È�ʬ��X69*"N�
!��+�"�*7���<����O�2b!�dͣ_d81���V�0i:�oT�/!�D�A�@iyeKȨ1���)þ>!�d�n �NЛ 'b��d��{�!�$�='��Zg�]<�pt: 	�2�!���|�&�#�D�Zn�c�O"V�!�B�0e4��(�^Z��#���' �!�˰K��]�?X�Xf`Ǭy	!�NQ��,�)�nqR�«+�!�E�3C�H	�͌��h�ĥX�f&!򄄟c�aѠH�=.��ADT!򤋓}�
�b�E�����d��!-!�
8d۔=���#��c��S>`!��Q.���C�S�	ᜉ�$f�!�J��;��S�����`"�z"!�Q�aԄ)RC�@#�`U�W,O��!�d�<v�4]a�@�[<��p��� w�!�8$|(��
�d9б�@~!�� ¾`k� �6Z�
=#ȹ�!���!A��oL��+�/K����'�4ŋ�Ė8����f.ȭ�i�'������Y��
	F9� ��'���Y�(֕�(@��� �>!�9	�'g:���B�9�bQ�Dk5
��lx�'0`�I�-W9S�Xq���D\5��'�:�c�Q'!���� �ؔL��%p	�'Q��2��#A�(�F�ːW���r�'� "�)�T��4�T��M���	�'�v��!C��6-��b�"R�K���
�'hx|�T�jġ� �·U��A	�'�lzV���viF%����r�	�'W,�����!d[G�
pf�y�'`BP��\�W��f!�ؙJ��� ؃�"^�����K�*zjܰ"O6�{���vL�ö��
R0!�"Oԭ�) ]<Pi�f�hj���"O�C��A&i&�҅�S��ɓ�"O$�h�-�Te�ҥϢa�M��"ON�`D��=�&��t1,���"OP�g��6~.�}�b��5NJ���"O|h��l�^D 5�G�����S�"O�y�����m� �I����"O|�a5����6�s]H�"On��֤y���vf�,m���%"O
5I��]2E |B�ޔ+Vnl�W"O�,p����S� ��a۞_>��@�"O�U�N����Q�A+d0�e�3"O�斑q7jxtA�~wH{�"O�u9u��3���A�@I��c"O�1H&��c& ����97�2��"Oڸ!��X���!��+u�!��"Oʵ�t�ەN�=B��P:>�R"O A����42�u2��Q-$10��"O��@�	�vY�P ��R6|�a@�"O^���T-M~����,ͮ8�v�C"O�5�`dGN8t �޷TC����"OBlB��� �\H�a�ɡ+MvԳ"O ����8+�H��bgǁ疴I�"O���˴f��Բ��	�.��"O���gX%7�"|����>��ՉW"Or1���M�ԜxF O"&{���%"O��C���Yd������$�$�g"Oy1 %w���Q�-�"WR�Ra"OBa��;h��ip'׏pLx`�"O0U��&˩;Fܲ#�B�>/��D"OB��L�z�8pe-P�}z���"O$hҗ�	���uaDQ�z��!�d"O4�Q�-��Q�X}h��ԉ*^ܨ��"O@���ҫn���eޒ%�|�Y%"O��;��N�r�Nɨ ��t��ɲ""O�PB����M*���%�"%�G�,D����^�5���C��?�(����)D�pJ3�ՒX�xH�Ȑ4��}ï)D��"���=d(P]���Y/V��U�&D�X!牨O*$�j��D�*ef�!��"���%l�$Ŷ}S�Ա!�Ĝ�sx ��5�xE�7� 6�!��7$������>{(�PX�!��Ћj���Ì�9,q�h��L��!��,���� ��	�2�z��J�K�!�dE?8�r-�Ť�6e��a#P!̀8�!��/	��`��P �m�3aD
"�!�Q8Ȟ��^>�j�O?Ne!���N����c���p𰤘
(�!�d�>t�`jg�739�y�lF�|�!�$�S��@��!N
G�y3P��0e�!�X><8�YL�9)2�C�)N6D�!�D\6�Z�
��N�c������$f�!��z( IQ,�b�5�/�Xo!���� 	� Ǉ�b�8�Q�d�!�Dͳ���+����DN*c�!�Éy�~��oX%:��Q�N# �!�Dŕ^~T��blV�;����� ւ0!򤐒A����FZ�i�R���`�7 !�>v��d�/�~L{���-O�!�D�6��Z�GPU��+�م^�!�$ۗ(в����H�ShD���>!�� � `�
VT��Ա��RZ�έҷ"O1!�4�dL)��I���DB"OF0h���9Ѻ��q���,�r9˖"O��HWA��~�ܸc 92�(�"O
�:��*<,AS*�7����w"O �j"`W[�Kթ�AP5y�"O`�ڳ���R��]
��� X�֔�'"O���e�o��)�RƞS{PA"O�,xQ	K|���AO�:gvtp�"O�y*���9�|5��"dm���1"OV�I��� k�X���P�R^�A`"O�T"�cе4��#��� /N���$"O��iٗ"����"�ɓG.�M�w"O��f��^Jx���@�&����"O.�����>0�92������"O@90v�֑[p��,|�\A�"O�8dD[�T�p7Q�)#P�3W�2D�Pq�@�I�V�B�l
�-jz �o2D�8ʤ��c�T��aL?F�@Dc�'$D���k�N��� %j�  ���/D���bف$�
�K	"D�hZ�.D�`E	K�c@v�����V�bp�*D�p�r���W�hu8���nQ��/)D�0ku�W��e��iQ�?�VM�S�:D��d��"�9����B�@E� �5D���%�5r�� �.4)�q���2D�8�2�+)l�l�����Pݰ�d3D������$sC������'s���0D�Цg�Yp�!�R�;�dP`�G4D� j��m�H��AK���|���3D���F�0�Z*��9�b�L3D��I��N�G(Q�蜾���E�1D�l�G�l@б�aY�I�qǇ+D��� ��WD^�wGٕ){�T!�i+D�T��
¿9� U0�F� ���)D��rs$˩b�2��R���E/(D��Z�   ��   �  ?  �  k  �)  �4  @  �J  V  �a  �l  �w  ��  #�  Y�  ��   �  O�  ��  �  %�  {�  ��  ;�  ��  �  ��  ��  ^�  ��  ��  ?�  � � > � �% =- k4 U> cF �L -S pY p[  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+��6-\�c
�<4�d5h��'�B�'���'	�'/�'�B�'���k'�M�=��Y�A�D�S��܃��'���'�b�'���'�"�'�b�'�t�"���#H( �TQ)G��ڟ���ğl�Iԟ��I˟d���x�	؟�QH��&
ga%@B�Z��[�$���<�I�	ӟD���������5i /;N`��M`�
$��J��	���	�������ß���4��$04��)�¢�6���N��|��埬��������p��ٟ�����D{ ��n��0��/�'j��: *]�l�I̟����8��ן��I꟔����T9���Y�`��DI ªK���韴��ퟨ����	ڟ���ٟ$�I럌aF��sk��C�cV��p��ɟ��I����I����I��(�����I˟�������H���-�^�rA��Ɵ���ɟ����p�Iٟ��I蟀�Iğ�yD� XCbE#!�0�� �����Iϟ��	͟�	�������������Ɍ|��Q�C�%����A��)n ���	؟�Iʟ��	�����㟐�	������Pӧᑘ �􁣃�ȴ1������|���X�	����	��|�۴�?���4_J�2���7[��R�Z"Y�VH��U�h�	Qy���O�$n�18�srʙ�2�<I: *�E�+n���D�O�H�'Zb'O�I$�	�5Kւ=U�`�aC>6�'�$�b��i��I�|���O(�j߸��t�ޫc��A��D����<I�����3�'^x��k��=�X5`\ u���aD�i�ҽz�y��I�O��L��y�bnV�(�BY��/��y����OL�	E}���b��^A��1OT0:��"*�x�ѡ�Ɂu�6�k�5Ox牘�?Q�N#��|Z��j�NlI��y�,�F�.c6BH����;�Ϧ-�a@1�	�q���й8)4�k4*��,~�U�?�*O���O���V}R�������wI��'~����
-��d�O��Q	ߕZ�1����Z�h��Ǧ殜pn� 6�@�%I�:�|����O?�I$4�wkO�k���׆G�O�d���
!?�������.��EC
|�	�
^dа%I��y2�'Q��'�����i����|RB�O;Q�'g��w�`	����~�2x�6�Te�I]y�O:B�'i��'�r�h�6*�E�k�4��Dc��I�M[ա����$�O��?a��B\AT�����	z�H�ʳ�VyR�'��O1�|�je�."�^q��4�=K^���
��<��~?>��:����U*b	8Q�w��	_�Tb�Fw^����O(��O��4�������̚/��N�C���X�ʁ�{�F�£f@��y��'��O��?Q��?	�B���Ą�$�sB��G��"�
�4���$Dܡ��'��O��ߡ[�lpr��<g�RxY3)��y2�'	�'���'���iW+pn����!��fȓ�0|˓�?���i���ȟ��$:�d�d4@�;�[�L���;V[�/�O
��O�	O�{�07�0?Q #�&�> ��"� p�R@�0��Rl��4$�d�'"��5�4�?�E�)�N%��Ȱ��`ם�?!���d�ɦճ㢇џX���O]L��3��:A54,���,����O���?�����S��J��(yQb�f0Is����D��A�=c�X�O�I���?Y�j#�dȺ@�x�	 �ƞm�|t2�a��1��d�OT���O��i�<�s�i����%�?4���-�N��ra���YV�Ɵ0�?�.O,�d��t�eZ1ZTV�tm26#�˓&&
�a�4���J�`Q����Bצ˓	��u�4G�	f4Q��Ki�6����d�O��D�Ot�D�O��d�|BD� p����&K�}+�
��\(��@3V���'-"���'��wq,�E��:Ok�%��V����'�2�|����
�_3Ob���! \��)!/�i��9��3O� b�؂�?���;��<ͧ�?�A&M�&ŀ!�θ\iJad���?���?�����Ĝ��*2O���$����XR5%A�tG�@����9~f�ǈe���$�O`��=�dƫv}���R*$�<D���[�I�0`H���O��k%xb>�÷�'/x��I�;�ص(�뜽���z&��L
���؟8����\��\�O<��U3x�r �@��6V�;���sr�bӒ�i�&�O����O����!�m�tD��)k�|����$qr��Οl�I�0+ ʃ殮�'�0�8u�C]z�.ڲx�$8�	�T" ��g#������O:��O�d�O�dV?s�*)�pEX�<7*�	ÆBuR<�ye�V�T�6��'������',z��)]4�����&���^�P�I�L$�b>I�g�Ǉ9�X�٢��$Vļ#�F�5F P�ú�˓vd����OL-�K>.O Q�I�<	T%Z4�P�~�ŀ�!�O��$�O*��O�<)U�i�eڀ�'K:�ɣ�_�ex����U;}�v!��'q��$�<����?��LI��F��&�*����K�P�wk�8�M��O,�2���(�4�� ���O��C����Q �"�;�0O����Of���O����O��?�xӡI�9�|�$���^�����ϟ��	՟x��4p\��'�?����->�)5BH!'qƥ 0����P)�<!������&P�6�)?��"EK��t;p&�	6����o��Qפ���O�O��(I>�,OH���O���OȽ��*�PT��A�͹y�ِ���OD�$�<���i�0i[�'dB�'���W���%�N��(�1�����O��d=��?��0�G�n�8|�Si��-`t�9����z�k%mA?���|
���O*1zH>�C�EI�c�M�aHN��� Է�?!��?��?�|�.O��nڝ���2b�*y��� P���bj��\�I��?i*O.�D�F���� $0����B	y��G�\���4����6�Ը!����ʓ7�@�����PB0a	������d�O��D�O���O��$�|�񭜸�8�x������dΚ����S��B�'�"��T�'W�w�Ll��]�'rp�+��V�zzDL��'���|����A�d*��5O�}�$!ڐy�� 5��f�t�@2O�9����?1�+�d�<�'�?�v��)�� ��JO�$���zD�?����?����d��%���DٟL�I��z���P�b��F��7rNi�K�m����ON��;�dY)Xpk�d+c�,)�u+ϐuh��&V���ʦ=L~�ui��(�I����K]�E��u�`�>h"��I���I����IM�O)�ձ$�ش���]�p=Iu�݇q`�h��@ٷk�O����O����5��8�N��p�`�2N7T�����x�	̟�3$�̦M�'1�\�4-�?���ܨP٘�2gC�}�Ri��b
��'��i>��	П���ǟ�I46oP�u"�sJ
&KM1�ʉ�'[�7��Kk��d�O��D-��#�� `��>/��YU��*���':��'ɧ�Ov�A�RFD:`������Q�����蟀e6D�;^�tZ�M�~��Tj�Igy2��8мqpDҋO&��p� �u"�'�'U�O�I�M�d��:�?�����(g�a16cN�]�4*��R��?�����']��Ɵ��Iܟ$�Si��Ay��WQ�f��TB�� r�xl�@~B	Y�.��D��\ܧ��!��C@�� ���5ks@`���<1���?����?����?9��dI��cP\KD
�_0���èɜ
�"�'�" {� D�B1�&���O �OT0��D X#����Udx`S�%���Ox�4�,��$z�X�ӺÅa�.I�ڈ9$)�Ja6]R�eJ |XF���F���ONʓ�?1��?��(��mH�$^7+��)�t(ȪF�����?�+Oz�n�'�4@��ܟL�Ia�$�	Ġy��� ��\
u#/��d�<���?YH>�O�����H�8A�bR�`FI��!�9py\�QwJ
�g�i>�a��'N�$��#�H(8�Fɓ�a��>!<C`�ݟ��I�����b>��'u�6m)�"۰G>!�|���.�RH�ல<�����'����@��HP���xq��@^��"gdy�\4y����� EH�b���Oyr�߂�Ă$G�,sQ
McreE�yBZ�@�	ПX���L��џؕO'≰ �4p����� u�6tr�{��5����O��$�OD���D�O�n
(�`�����=��M�2+&�6�)��8��	n�<a�A��t�,-�n�;��\�g��<A'�"'��d�5����$�O���)qN�"�%�c�:,�զ{���D�O���OV�E��&���B��'r��)/Ð��Z9i�b�xK۝N��O�ʓ�?���� �L�Z#�ǧU�@�h�Ă�'�4h�V�B�(��-)����ϟ)�'��X8���)KwY�%�Ӏ#�z$���'���'��'��>��ɖ>A�P�BD�8
x�gM��L��\�I��M����d�OH��] "��DB5E̩L��	q�C$d@�I���I۟0z�
�֦��'oB��P(Y�?j2��༒Y�@)0@)�^��$I>)(O�	�O����O*�d�Op����	+h�< f�C`����<q��iC.ة@�'�R�'��O����&B6�����<g��D��.	Dx�I����?�|����hsX��3��?x	H�G/�����Q4'���$�'"R��V�OZ�-�f{����&��� -�$���Lҟ��	ޟ���՟�Wy��n�\�P��OܱY6�1R)�⧢1	
^m;���O��-�	dyR�'o��'@��1g�5F�*6��hP��S*܇/����Hc�Db�čc�S��IsG��ఽ�an�-F	�0�l�������ٟ��Iӟh���D��U�r����C�%;r�Z��V��?I��?�s�iÜ���W�`��^�	.U.\! /�!��)1�E�v�&�(�I���Ӻ~�&lo�j~�KU������&!��M���]0�*���Ο@r�|�^����,�I���S�ȇdJ��G�؅�ZM�蟔�IZy2Bb��tj���O��d�O*ʧ U��"���1\����
X$28H`�'x�	���	k�)�0BR�^LKת��oj�
�N�
#LE@Z�[��������K�|B�$ iC���9�J)h�r�'�B�'����Z��b�4^Ƽ�p2��;ua �����^��<��⚎���Ov�T�'P2�O����3�=]`���fW�iC�' �8���i[�	�.����r�� ��a�E��-x(@�l+h,�M�<O���?q���?���?����iS'_��A�Κ�3þ�	kU��V�n�;��Q�'�2�i�O���(|N��I�O0�0��@L+W�|�$�O�O1�f��A`���I"J�.,�I� [����F�e3F�I�*��H�u�'e�%�X����'n0! � �:��Ip�ozZX��'"�'��S�����6ޘ��ϟ\�	.w�X�u��,������;"�H��?q)O,�D�O�O�p�A�S,w���r��/���:c��l#@�J;����&RH�<r&ڟ��槗��29�h��'�Q���ݟ��Iן��	ҟ�E���'��P����Դ��]��v�'z67-��x�^˓�?ɋ�w�a0�N�[����5EL3]:8�'B�'W�+ne����T�I�Ą�/��+ ��L4��vH��e���&�Ԕ��4�'���'�b�'-2����I��P\P��
�C�)��P��#شT�^J��?9���䧄?c�����2��IrO���&�@�����O��:���7AЈ="�`�>�M�"@�'~PV�`��t�Ԍ�'<��r?QI>�)O:�KՆ�B��7�F�M5NP�4��O�d�ON���O�)�<��i|~u���'5��Eኩ%�~��`lF�j'��
F�'����<1���?��+�Y����1W���$�3���j�'	�M�O�0�+ˆ�(����Y!ZI�قF�@�v�$��a�/6����O"�D�O����O���'���l�Z��_�L���i6��q1f��I� �ɒ�MC��|"���?J>�"iæ�VT&혟 �����EB���?���|
b��#�M��O�.Ȧ^�(SI\58iX�!�,	>N�vEAE�O�U�I>I-Op���O���O��*�U06�I�EG"�
W�O@���<	�i��	%�'�B�'���M~�e�F5n�*��N�!#����O��D ��?5{r��k�ԉ�G�Sf�&���,ڳ'W%F�y����|�$��O��cI>�C��2�
$9SA�.\ؘ%�B�_��?q��?��?�|z/O�`nڻf��e�P�H�	l���9%�L�$h_Gy��'��O˓�?AQ؛R�^��N���k��#���Q��6�4?!5(<u�~������J�V��t#Î��y#�ꛩ"�$�<Q���?Y���?���?�/������.� �Q�ԃ}|�8����u8C%����՟@'?�I��h�jw��H�F�Vn�_�����l%�b>���ڦ��H�D	�e���Pdr��M�͓]F�)�h��@$�������'�T)�F��2�Z�C�v��A�'���'��T��޴-E��P,O>�D%o&�SS�O
#$�Pʲ�
�a"�T�'���L"�:��	^,���i�	тXw�I�X:��h�]�� �$?�x��'� ��ɫp��D���
jJ�E{p��D=���I���I䟴��{�O���T5R�%9��Q(.	��P�͚%��&}Ӵ�A�E�O��$�O���]4$�ar��F��@t��}���	���IşLb5��'��0f�aZ4+�$x��=o˅�"�I��)����4�B���O����O����%���!�Z�k�����/ȷ��˓r՛�@�E�'�B��4�'�x�@��IO�pWl��Ȍ�]�<�IQ�ŞV(b�`�*�/^h}QFlG;lP�w���3�� �(O�@�_�?	��+�d�<�tj�/�t�X�'��@qҘ��i��?����?���?ͧ���Tצy �@�(A���bh�ҕ��	g��37�ҟ���n����O��4��Tc�1��i�@-b�%aD�� ^�7�2?����
8"�SQ���E۷�K�YnB�M�+��(�hx�P�	����	��4��ҟ����פS�H2�lX0N�9A���?��?9��iH�W���	k�d�����'�!�̳�m�6�\�%�������Ӥm��m�A~�&�9b:n�+5r�� t?}L8�����8Q3�|�R���؟���Ο����G>` ʤ`�nB�= EH�ş��Ily�qӾi���On���Oʧ6�A	Sǈ<zф��S�Z�hh�'4�	��T�IZ�)*&�MW�����ԸY����
b"���T I�Z���� 埜"$�| @�[:�5�C��2��eb�K-|��'.�'���tZ��h�4J썊C�JOJ�٨�܃:�
Q�E����?���?��Y�h��6g֊GkK�%9ǎb0(ɖ'�0 f�i���j�x|���O�(��'�l�q�Œ_�BL��(W�vND]�'��I�����������C��C�%|�@�a��P
�Y�f�O�	�6��9�(��O���&�i�O�4� m��Kӣ(����i�x�y���O���*���B��7k��3/p�� ��>��!�a	S��y�m�b*���������O~�ƢPlad�Ѯ^v%W�!M���$�O��$�O�ʓ<w�&�ޓ/���'zr��W7b�ـc��X��q�^<]��O˓�?��T��(�D J�L�5��Ξ���� �c��P�&�c�0���X��a���DY
=���'�Я�ة��2�6���O����O��d?�'�?�G�J�)��X�s�#}�d�y�'ڜ�?	S�ix�y�_����X�Ӽ;�%Ϡ;�Z�a���eS�u�PB�<���?�o����4��Dؔc]0���π ���qI_�66�� � Z9@k��;�ı<ͧ�?����?���?�u�ͽXrj�����0n��g����d�Ħ�J" ��(�I��%?��5=h�G,ش_>���ß�I�ܖ'R�'�ɧ�OŖ;$��K�t�k%�۾cT��ɷ[�>�X��O�	�oA6�?�O<��<1v)��%��va�'g�,��!�ǘ�?���?����?�'��$�J�A��\jU�yG�e8�iޡ3N�0�n��?a����'����t�	埬3Վ&%R�c

:B�t��/	�C�2�m�S~���$�H��Ӌ��O�7B�= ;�2�L[�w����2*ؖ�y��'�2�'���'}2�������8�K�H��� ��>#<r���O���Ʀ)��g>Q���8'�ؕJ	u���+�e��N_R�R��$����'v8��i��ɀ]�4i�J�+ M~-�န�)&9�FeP�g���P�IRy2�'2�'|r��6:{*���l��Hׄ|�f�S k:��'��	�Ms@�_�?���?�(���3�T�A��ԧG�в�ᜟ �'y��'�ɧ�	��{�JTjAGʀ �|�Al�$xje�EOGHX�'�<�'s2�$���&Kĕ��iܗV�t�r�B�3��;���?���?��S�'���٦�针߱r��1;I֎e\D�Y����[���I���	Z���D�O��ZG V����7d��.��-A�F�O��ğ�7m<?��EЪj1��>9��⁘e�j|��$�%9c���d�p���'���'��'���'f�<L���C�M@��K,>�s�4g�>�Q��?�����'�?��Ӽ�r� ^���Y[c8]A����?����Ş=�t�ٴ�y�ń�Fm�!���*����$�y�A
rwz��I8�'u�IΟ4�I�?P���_�8k�E���|$�����IП �'��6m�&1����O���4:u�xMڝW��0Z6M�n�"⟠�'("�'M�'j�ACH�"� ����b�|[�O�APs!R*n66�%��&T��d�O:Eqw�����ks�D�{��ڔ��O���O,�d�O^�}��� -Ӄ��^g��� �_NX��#�V%B�Q�I��(�?ͻT
�KLЛuD��Xe#7gA�@Γ�?Y���?�����M�OD�(�-��zsL#]���܅�v�˰�f�F�O|��|���?���?Q��M�9���B�I^��Ef�E/Xj*O2�m	�: ��ӟ|��J�s��)[�J���+ �!�L�р��py��'tb�|��4�@TWT@�@�͞>�pEd]�z�\���B�����Ⱥl�$��hJ�O.����� H
3���*W��~��T���?���?9��|�*O<�oڕV�����w�0�:dBT3.��$Ț
,ȉ��ݟ�?�-Or�d�OT�d=D�:��� ^17NDG ؓ>�xM��.|���`O� #Q����>��ݣ>|�ڶIE<v�@��J��*zb��쟰�����	䟸��{��M�h�w�S�C
��i���#CT�
���?Y��z$�&c��S��џ�'�4�5f�$T\���g�V�{��	U�Rr�IԟL�i>��Cf�I�'�r͘vC�2e��=H�!�H��x�.W�0'<�I�D�'#�i>��������_p�l $/[0R*�1g��B^\�	ןԗ'R7mD*\����O�$�|B� ��+m=�G	T�ْVb�C~V�H�	T%��'R��Ѫ֭X*��;UCuU����T0H����AŨ����|����O2M>���E�v�P"��ȥZ��X�L8�?���?9���?�|�/O��m�M	�Ȳ��ϔ)o"=�B�36S� 	�B�my"�'��O���?�2C�?"�3�!2v�A��T�?�N�\�ش����%���A�)O�P��dB_�T{��P�v��0�?O,��?��?��?�����i� nl� �iL���T�J�D���nژ_�2,��ן`�IP�ןP�i�혵��2,�e�ŗR�j��s��ޟ,��r�)��Y�(�m��<�b��$s���PJ�C>��f�H�<9W��S ���B*����4�����_(�4͐3!6� ��b�.u �d�OR���O�˓�֮ĒGB�'�BcA��쳥,Ы&��-X�C	0�O�˓�?Q���M����	�>,�P��䣞�ג��'Y�`Ռ/��6��X��~��'����5��2ޜu	�� ���i�'��'1��'��>�������j��ۊU13SL����I��M֍V���D�O&��|PX�!�Ҝ8P2<���Fe����L���H"���릡�'�����d��?iy��΢!���1AQ}�t�裀�5}��'��i>���ן���џD�I�
�|�y6� ��m���A���'/�6m�(���O��#�9O$̒6@ X��Ҥ�)T����K�<����?�J>�|t��# �y�ף��.�)I3��`_�@![n~�f·#мL���\��'��� 	�`1�����Am��*w��J��8�	ğl�I����i>�'��7m�MO����B�dI���=5��x�t�6H\�$�O���'���ygϙ�~�堅���mD\��P�C��0�B��i��ɕ_~�c�O3h�$?���"E�0�ҹQ�|��&o��n��I��	� �I�����~�'4�VؙF�֡ ��50�EZ>N,��R���?i�8r�F`��^h�I���%��z�o�<d~H���21b������o�	�$�i>��r�ڛ����z�j4� �H���l�$�
�)�2�:E�R)˔�?��m"��<ͧ�?	��?�0X\�4��#�M�>�e��?Q���ܦ�Y������L�O嘑�`Y�z:�P�j�r�����O�˓�?)���S����[3~L���R�w;)����,�E���b	.�C�O�Z��?i�H'�� 1-=Fe�N՜Fl̨*@�	R�����O���O���i�<���i(fQ��!��x��3�n��%������'���'��O���?ч*�5|��\R�N��":L+7f
�?��pr�P�4����r\���Xk-OL��p _���yk��q�F�Ŀ<���?9��?���?I.����,�ը3�M9wG�
��������ß<$?�����ݤ�D���3}��<��nx	lM��ڟ8'�b>a�0��Eϓ-n* A�AB�7� �B��Y�O��Γt�t�s���X'��'��'	V(X�'L<ZD�t��!PT2���'C2�'LP��iڴ`2UB���?���y�lb���Up�q4�"Ƽ����_�0��R��X�1Z���-|����'�$U����'�L9s�m@�E#4��2��t- ⟀���'J�
e�54&����0)�,�J��'l�'���'$�>y̓]m�,J!��;h�t9zUȋ(a�u�	��M{�`�.���Ov��]=@�3R"_�$f�= $.�"0��џD�Ißxa�����u�+�'1���T�S<f�pR����D�~�<1&���'�B�'�'���'  ���E�:�y e	�tU�P�cR����4e׆�����?����䧐?�g �w�0�#��,z����D�O���9���(D�03�(fȼ�!�bj�R��}��%�'nhRsi�S?J>�,O]�D`S:.��d����6S�4�T��O��$�O����O�<�ǽi�.ܢa�'�h�bd䈼�ʱpDA� 2�؂ �'�"�d�<���?ͻ\�Uڥ���M�3 �H*`�Ī�Mk�OJ yB�U:���D*��wޡ�$�P�;��C@F�q�B��<1��?y��?����?!��TA
1E��)C�ʌ0{z1��c֒s�'��$rӦsf>�@��O��OZ�C�}(���ԇ��
�~���Hܚ�䓺?���|����"�M��OX9)U�.}N���ƊB�j��Fں������uj��O���|2��?����.p�P�?��u3� \耄Z���?a*Ooڽ$ ���ӟ4��n�$�Z29DT���:mM�X�⧈,���<���?aJ>�O���Iga�="��A0̅*3��!����t.(���io�i>��$�O��OrYТ(��g� LO������On�$�O����O1��ʓD:��@	�g,$0��7)�$S2�;d��`�PV���It�����O�0 �(%oεp�G�q��@C�M�O��䁈#!b7m>?�B��y,��)=�'�y��Z��"5�>��I��yB[��I����柈���P�O��Y����B��r��5G�(I(��t�r4x�A�O@�d�O���F���O��ݿ*0E8�cϭCG��֧]	)��d�O�O1���Q�o��牝l��Xy��uX`恘� ���ɕW�ڝ��O��O���?�8]q��_�U����	0Z�V0)��?����?,O��n�b����៸��2�L����:%�0z����-�?�.O&�d-�ɽNMı��B�=�
�+1��f�{�0Α�#tQ�M~R!n�O~Q���<_F��R�5gk��;hF$`��̅�%Br8��π	@�*��oR��91��qԛi��|�b�'��4�}06CZu�H�C���8Mp�I�4O$���O��dR>6�*?aC"Fh��?�ܪ�aո'��E�v��=9� �&�T�'�џ��V�߈&������5/�:Z��!?9$�i/�� X���Io�'^F�!�dVB�ɳ�Ԃh��t�+O����O��O1�� �gG�I�`dc��S;h�Α+Ѯ�7�P�˴
�<)G�O�r�B�dҪ����ď�b��R���z�����a|҈bӬ�b M�Ozt	��-	h��k٧8��!q�;OP��7�	zy��'���'�tL����Q7�ā5\( ���*ՈYw̛V���+��>���@�_���ъ�nߝ#X>M"����7�L`�C�o�؅�	�D|2�����8f�n���MU#"̤��ϟ��ɧ�M���Y�4�'��'d�����܂{�d�e
�?�:)�b�|b�'��O���i��Ij�+�!��c�];�.l�s&�����'��'��i�)h�R͖�FXj,J�g�TM�Gx�)lӄ b���O���OV˧Ww ����X(QPF	U0jf�'q�	ȟ���z�):sK���Vݚ���&M�.�!�3�$8s���M�']�擟��d3��D$����G�>�4�BӣD�]!�B������!)��u�1(�y�x8��! ��'���D�<!���*�Ӗ��b�(դ܈������?�dh�M#�O��`���݈��D��M��R��!�ǔXizE0Oʓ�?����?Y���?����iL?x\I"AFn�*�*E��l&ؔ'���I�O���9u�f�I��i�IY1D�*R���d"�)擽!��nZ�<� Zq���U?H4��p����Ua6O\A�dB��?��i1��<Q��?ip(08z��R�,۶~x��W)Ք�?���?�����d�զq3I�����	ş��o޸:�80;����tT�W��|����d�O�⟄j���5��%�$ �	W��͓��6?A@�A��9S#�ٴ��E���D�4�?��]O,��Ǆ�2P�	;S�-�?i��?���?!����O��SJ�; t�壓0P��j�Oo�[�~d�	ß���B�Ӽ���4/��3��
D�0�q#`[�<A������v��6m!?I�˕2 ��)�	B�L��z�-�Bͳd �,�cI+�$�<����?9��?���?�I��eѪ���̄d�XRDM���U��5�GƐ��	�h&?�	 �H�V��9*�Ѐ	�+�T�zЗ'&��ɁdY�-:�@{��� �9+n��p���"Q���D����6c�ONe
H>�.O2͐1#�z�(�b(�*R؉r@�O:�$�O��$�O�ɡ<'�ii�)��'�*1RW,�2�#؂�X�1�'��Ĺ<����D�6�fP9u�,�ZaBg���5�S� �^7(?y�'��6�I�	�䧉���,4���<>^�I���<���?���?���?���T�� *�QxS�ӣ �L�q��E�4���'�Jq��(Ȇ��<)���qD��K��2�M��mɧ|9H>����?�'6�����4��$@)Q,�sw&� $��X�64�yH�g��?� "�D�<�'�?����?1U�I�9j��f�
]a0C�o]�?1����[��9�'�ɟ���ퟨ�O�
D�A� �\���f$d���p�O�ʓ�?����S��J ���Ự��x����C�8���a!� %~i��O�i ��?� %/�$�J�
ar���H�b造���	�����O����O���<	��i����	S-� �)dLA�_ϬL)s�:��,�?Q.O�DY��0F�W�'��ke��xYt���O���q�b���/%,�AE@�N�O�~���ք��a�[�Xi^ [�'�	����I�<�	���IU�$您i�p�ڐ�R&6B����
Rv6�3T��?q����y�(_;jìl����0o�{�Ʌ�2�''ɧ�Oa�Y���iw�I5�RA�a��W6`%q��[�r�'� !0�&��Z�|�V���ǟ0�TOG��:�Zs-�h�:�(���|��柀�I@y��c�tq�a�O���O�Ÿ�Z&N�:�Ǭ* �ළ?�	Py�'Gb�|r �)���FQ�t�M�����$��(�qe�ߍ"E1�u8��'E����/ $��d"����$�G��_=l���O��D�O��$;�'�?	A�]�(َu��f�'jX�C�e،�?!S�i�4��ݟ��I����?�;M`mXb���2*�r�f�-�l�̓�?)��?�M	�M��O����
/�ҵ�]
�!�)ՉHiР1!��qړO���|����?����?��z��q3+�;����%NJ/�*O<|nښb@D��П��IK�П��بb�tɪC$ĜD�t]�A�Ky"�'3R�|��t�٠e�1A2�{b\� ��
A�&��U�i/�ʓ07��'I���$��'>�Z�(Դ;�,	u蟒8�ũU�'�r�'�����dY����4	g$����x��p;v�9Sj����?)�b]���	�8�I�B��9 �g��Ƕ�3�߈[�T��m��Q�'"nRՏ�o�M~z�;K
�0U��I�t37��:�*IΓ�?����?����?�����Oe�IZ$��v.,�3�!!0e1�'�"�''z6-� ��i�O���%��D� ,@�#N;�Zd��,!RhH�O��$�O�
�fn�7�6?9�)-�d��� ��V!3tF�5�]AR ��H%�8�'SB�'/��'v�	�D��R����>�z��!�'��Z�\��4l�i��?�����_gP�R�F֒rWzq�.�7N�D�Oʓ�?����S����}z�d�փ3]b����Z=�����E�G���-�<�''#,�	F�I2!ښmrֈ�d���kZEk���������؟�)�Iy��m�����Ojg� Qr/D�P�P�W-C�}�����O8��-���OZʓ�?����a֔ڕ�ς$*�m3�M��?Q��%��q�4��dE��^a��O��	;��z��Ɨ�E	Z�<�١:Or˓�?Q��?����?���򉆦���C�����0(ÔG�n�;k���I��T�	N�ß��iށpd�ͅ/:�	Q�*@�xۗ�
؟\�	p�)�ӈ�0�m��<!F(ۢ/g�R��92��s �<�rfH(���IL�	Uy�'����
)��1�wo�U�,	���)}��'���']�	<�MS���?���?�a�:r�(�n�<�(��ƨ҂�䓍?q+O����O2�O�!ІjM a�I��#�.0�|hJ���<����-H��]�4�d��)I���C��T�lW�-a��!eB��:6�@����П��	�@G��w����פ�!}"�|� O
��Y�'{b6M�}���Oz��/���O�����&�C"&�,tB�����O����O��a&�{�r�Ӻ�BT��J�-E�^��V&F�M��%�P����O�˓�?i���?���?��/�X��t@Rf�t��A��Z�fI�(O�oZ�A1����ƟH�	p�ğ��Td��h&��G�Q+<X���u"Wuy�'��|����A��� ������0̔H)&��f�~H�Щx�5�'�04J�b�D?!J>Y)O���G^Oz���IǾ=\�i1b�O��d�O2��O��<Iq�i��9��'�P�x�k�.�������� f�' �|��'����h�i��ON�b���*��q�tp���I�{� �mZj~���>'�l�������3����caD�{�.]�#$����@�<1���?	��?��?I��D"
6d��p�ņ� y�@޸ 2�'2"�u��8�2�R���O�Oĩ�%�Gz�
9� �n�LYҗ <��O��4��qe���Ӻ'���D���c��s�ܜ��˃�)NAr�c��OB��?)���?Q��n�J��Tв$#��:g�A�v�0(P��?�(O�An�2FbT�'�r^>�IdnQ�LH�5Α1�9{#.!?	)O\�D�O��O�Ӊd=-���MsLic�?6֙H���
"���nڛ��4�r��'R�'-���	��e�: ���pX@���'�b�'��OH�I�M�F/�����bI�>;��X�dݛZhT(���?�����':�I���)�dG�+"����"0#T�QlL̟��	�L��l�Z~�(��������
(ζ)"b�&+�´�c�λor�<��?!���?���?q)��( b��n�T��D������"�ʦ�(�+����I֟�%?��I��1JL�!�]�e�*�'�+����ԟ|&�b>����Ǧ�Γ&kD�:���&u��@��Bӟqy���Yxm����&���'�"�'f�����t��A���҇A\f}{��'g��'�"P�\Aݴl~f����?��,�
HٶgI�d�맊cdL��bP�l��ݟ�'�H�S�7[� -iPi��ZGt`d(?QҠڪ~�I�4��O�����?	�� 0w"P	�E�	�x00�7��?����?���?���	�O"�;���9�=� �F T�*��6��OR1l#*rB����D��k�Ӽ�@� w|.��!��\�$�2(A�<q���?��:�U+ݴ��D��	�j�O� ��*�<2�g��}� H��|�W�x�I���͟��I��4�ԃЄY���q�+�ӲE��dy�Dp��ex�m�O,���O�����ɾl��R�Q�305��!�/B�˓�?����S�'Q�aA��ǡ~\����n�py@�%���n��'�ԡ��G͟� ǟ|�W�� ��8� �F�¹17^ɟ ���D��̟�SDyt�V���O�4z�h������fފ1�4O���/��ey�'E�'��[��C�2�6I*b9�q[�H,Y�������hE�|��4�)��\������?e
@z6�C�H����$K?3��S'�q�T�+�H�r�$����1c]z����F�\����`&@)TF�²*��d�����\�q���."�Z(�&�"�0�T#��c30t
3�
��'2|s铮w��kȐKB�y�b����G�X�L�Tyе��=>���㖤c�����˗W'A9S`��V��[ōx�*�JbcM4 I"�%��-���a�/��.��cѧĳB�R�0�l�Zl��`J:arLˤ������T*� �٘�*�:\�PQ�L�0Iԛ��'7��'j���>�)O��$��P�B��=B1f�Y�(�$�CТw�N�O��z��Do�S�����ğ�itɃ%�t�k���*J$j�����M���O�N�sY���'�|Zcbz#�JP:��d��J�!�O�����O�ʓ�?���?�+OBЫ����8�R-���	8\8Rc(H�	(�'I�	��$���I�
a�Y�d�wl�e�� ^�T*�b���	͟��	vy��̀x�T��N�$���7qG��rT�AM7m�<1����?9��cJ��@�'�n����
Ap����&���N0�O6��O����<Y&ɏm��Sҟ���P�v���t�G?Sր�r�,�MC����?I��)�}����I�i�>��pgA�n^*�"�T��6��O���<q��4��֟���S��IM� 6J����!(�,9pa/�`�	�\���M"Z��?��O�Ԍ���X�B�얰Vծ�H�4��
`��n�ǟ��IʟԔ�yZcD0H��'"f*a��S�BzƵ ޴�?���f�83��	�j���c2��"��%�!�e�F א}��7M�ON�D�O��I�|}"R��C�̎$g�-��^(Wec0�Յ�M���(��'��N�D�3x_�}2h�Y�qZ��4���o���I� �b�ҏ��D�<I��~B+ :n����ӧܴEb`�ف�MsH>y���%�O�R�'@��N9^�H�1@�Z�U�Fh
�Ƈ
ux7��OH��J	H}�Q���IZ�i�au��"���CB�G7v�V�؀d�>9wI���䓂?q���?�,O~�J!_[ ��1��̂'ʄ�X��W"h%� ��՟H$���uW��O��.bF��5�&�M+���D�O�d�O��l1���3�D��� u��!&+]�M�|e�2\���	�`&�����T�'؈:୉+,X�R�����E,�>1���?	�����G�(T�Y&>}k�(��b�� �=5V�q�O���M���䓥�4����(��"Z(��KuF�1��؉��A��M���?�*O��r��T�ݟL�s��Wș�p� aP�'-O�:����&�d�<����?�N~�Ӻk2V@��j��&Xm*=�FgR}��'�>�bC�'[��'���O��i�y"�*m|DL��C	9�mg�Z���<q'��ħS�X}K�E�*R'$���+�#^�om�����ȟL�	៰�nyʟZ}� ީ�5��iì�)���`Y0��7[����"3�Ş�?97 ��dtP��"�XS�MF�4����'}R�'���H6�4���D���Xgi]6&L��t�}���:׋r�z��$�$e��O��d��lB��ۗ+�浊pJ^=r�aQ�>�`��D�<����[�b̌!b(�m]Dd�dMŎd��ODu3㖟��	�\��uy��\:�Lu��B�=Mt���i�'�L����4��O��D'�$�<��,gp=2�`���8�iBހq���o�`�'���'��U�(D�� ��TJ�>,S�0��d[$4�ށR�b�����O��d4��<�'�?���D�xm�x*3�0�9bĤ��!��ٟ�����']��둈/�i^i���
��\���h��&�lZ��$�����'��v8���@�ңE5\��j�PN�oן\��Kyb�����b����kO���r6Ɏ2~��!Q �5�'���ǟ��x�s���8pr/Ӆ�0��v��68��6-�<��a��T�����~���
B���j���4)�� �Ō/l�b�m�2��?���h�O\��M�&&V�P�@IєO�x��Sߦ�q��؟0��ɟ<�I�?����	V�-x$�s�lC�&��2LT6l��)�'��z���}nf@����| �(Q�F�1U� d��4�?����?y�J\ ��?9�Op�A���tj�Ѥ�3��t ��b�';��6���O��$�#\,�u�P�n�D���NA/yop�o�˟�S������|�����Ӻ+�k�!�,q��}7�4#�Nv�ȟ@%����]y�'��03�A1JF�0�J�0���A��L�3�����	[��?i�'�h�c�&'_��Af�V*\}z�4]���'U��'l�Y��y�����D�e��He�M&S?d![U�A�����O��d9���<ͧ�?9�l�y�
k$�ƤC��AS�)��XP���(�	ϟ��'��ɐ��6�)�n���Lʄs��x�L�	)(MmZПD%�T�����'��'`$���+F�ߺ	JG�.���l�����	wy�ֱzL�*�D�kL��(��M���"���@	< ?�'D��П��IE�s��ݤl0+VA�;���* 0vܐ��?Y�� �?��?�����,O��[ l�jR�nS8NvJ%�a/ױ?ԛ��'��I�Fp"<%>�Q`� 
�Rk��Q�B� ,�x��H�CA��!��������?IJ�O�� ����	,d)!DFн' �%g�i-���'��T������=�d$�a�5/��L2e��2�VH*'�ib�'��ē5I�����O�I5b]1�vk�zdBA0�Փ0�R���H?(z�i>u�I����	Cl`ٙ� C�\��Gojt�ٴ�?�C/��w��Iey��'��	�֘$6.� (Z"���#��(J��BXb�͓����O��D0��OJ� )�&�ɩw}& �Ca��C�N�H
OB}�Q���Zy��'�r�'��$)�Kۖ�| ǧG�Dk`�p����y��'}�'�"�'��Ɇ74� )�O�fa�E"�a�h���UR��޴���O���?i���?����<�R+54,�t���H%`'���.��I˟��	��̔'g�0����~���4,n���aGdx�T;�J�������i��]�������	��c>7��7�^�S@ɝ�n�L(b�ۘ����'6�]���H�!����O�����4��g�������{��:�%�[}R�'��'����'b�]���'��Ě���,��Q�Й/�zXmZVy��S�JZ�6��O����O��I�Y}ZwĜ�`T�D���q��c���dGi�z���Ot�ѕ4O�(��yr��L�3	���'��8X�>�z��ЛAI��9^/�6M�OH�D�Oz��T}�Z�pI� B��Mi�6��$J ��M��� �<9H>Y����'t�����9���0�����i�`����O����N���'��џ��QZޕش��
z�t���ǡt3 �'��.x���|����?q�w%6ă��֥7������
Y
(U���iqrd���ҨO���?�,O�������k�Bi�m�@�T�(�PM3D^���x�H�	�0�	韸��Ty҃�n���WC�2k}�pq�BR�U�U�`i�>�+Oh���<���?���a��dh�OT����Z���+Fw�pp�P�<q���?���?�����X�G"̑ϧ&s�
�
-$���4H��oUy"�'�I՟\����D:���X�
3�X����_	�� .��Mk���?I���?I-O�5�o���5�S7k2�Sób���(C��M������OJ���O���1Or���&�pbܥ�D�K��V%�׊oӠ���O�ʓs�fAӰ^?y������8tޔY	3��l@*��Pz
ݓ�O��$�O��ͧX��$�|�����>!��
$��1.�R6�M�/OE���ঽ��������?��O�Y���lЖe.4F��i0ݹ2X���'������ħ<Y��T�,|�$�ȦJ��OY
l��=�M��$yڛ�'�b�'��� �>�.O�tJ�SV�Rb�� Ht�1@UȦ�iS�"?�)Or�?A��@� ��f�d��Ks(VB�P@۴�?Y���?I�EZ�k�	Py��'��$(_�ȢE�=��]@d���}1�F�|����yʟR�$�O��$�Y�.�{�"�w�X9En�ƀl�ş�C1�V���d�<A���Dȼ� �!A1#�p?f���Y�m^�[6�ipB����y2�'��'xB�'��	� ����	�)k҄�WC �8v�� � L%��$�<�����OJ���O�|(�7KGZ�`rbJF��02h�'d�d�O����O��D�OT˓#Dv��0��+A�Z�O��!K�
;8�(ubd�i-�	����',��'�����y�@	w�N���8O�
L9���Q��6��O����O�D�<��fާ�O�N+�A�]�G���{��т!a�x�� �$�Oz�d����7}R��$�m;�+S-'�P���_��M����?�-O�u�s��R�۟ ��$��4���%b� SмQ��S����?q�R�x`��������+8^���&G���B��5(U��Ms-O���	Z��|���j��'�d�Eđ�x���(M�` Fq�4�?9��
�����䓠�O��<x��)�����  m� ߢ �4�?i���?�����O�<�W�ٌYh��5�� Mɜ8���ͦM���l� $�4����F3hx�#�թw�8���G��*P�Ѹi)��'��fȄJ�c�0��v?�&�C)���}2�|:"�Gަi$�h+ �b���?Y���?�P��Hh�=2�n�;������?3D��'�F�y'�4���L'���o� C�")��{�A�xoP�I�� �<���?1��򤛳\�R��գK&$�.Փ=�mH�)_�	���	p�I���I'4h������q��˴��8�Z���-��������'��lc�>� !ٛ7�zx0�R8��1�bͰ>y��?AM>q���?ٔ�O�<��,ʲ)}.ػP��
M�(=;eO���ğ(����t�'O�P!�;�IJ�M"�e���4��;�D�u�X5m�⟸&�����䫗�ޟp�O�u���0��{Ӫ�^��5A�i���'n前/��iI|���2�BG!z�����ֲK���Ժ>T�'4R�'�i�'�'|�I�0�P��5��[$���Pq�V�ԩ�i�M�W?��I�?�
�O���DY<#MD�q�K�J�)¶iCr�'���w�'D�'"q�$)�.ʅgjtL"0�B�#>)��i#�`�!mӨ���O|�d�ҩ�>т��$&����A,ï 3̈3h�����,ʧ�y�|����O�R`=m�b0	�^e�"�B%����	̟��I�:��M<���?��'�&%2��4f�P��.�]�t`޴��M���&��4�'���'�̀��.��c�^�r�̴:�Z�q�t���$J\A>��>�����{��)��z��I�W�U�G��^}����y^�x�	��x�OT�	\�P-�� ��u�� ���E��|���'B_��Ik�ҟ��imt$B��K:(�)�Ѣ?ތnZ1;���?	��?�*O����͕�|�mT1m��1�OL�`\�)��aY^}�'��'��O�!x�R?��RiJ"k�T,q��˔L/����>���?����?���E�x9�,�����:�ܘ���ߙ���§�ݸS\�l�ß�'����Cy"ˁ�ē�T x��%/� �xqOO�ym�An�ßT�Idy�#R�c����$��t `!�\<9m<�˴Ê�_Uv%ۖÞT��՟���
`R�#<��O��)r�!ތD�n�`Üs��	Bݴ��X��`�o$��I�O�	�y~"A�1<� ��ƻ0N`���?�M3���?ɤ�BE�'�q��]���(%�|XP�۬20��u�i֞�E�q� ���OB����4&����'	l��L�5mlP@�,����qݴJ| Ex��	�O��"�e���i�լ�P�ơ�Ai���	��0�Ɋ*�Y�}��'x�D�?5�p9b�柒:p����i�j�OF��A��O���O�P*�䟣?��9G�D�P@F����� 4�J�kN<����?1O>�1-nX-+p�إUD0�Z�bͽ`N@a�'�2lj�y��'���'j�	e��k6)ՠSFyK��WzQ.��&M��ē�?I�����?A�	��b'>9؊�1+D�HKrD(�G�J��?���?����?	v�Y���ԤL 	ʹ(��MN�8�F���ҿ�M+��?��䓤?	-O  ���ix.�:���) ��B��BuګOV���O���<!�
@$%Z�O���9¬� I�����7rN -�g�r�X�D�O⟤�J%�/j�a��P2�h���$F@�7��O��d�O�$ʇ%:�'��$��7��+mb���O�AF��1R��t�	ߟX�'{�������1Ea
�[�ҥ�c��	4�vԂ�i��	�S1Lh#�4 ���P�������#^�L2waQ3~�(�g�L�v�'�2g2�O��>a�/QB����uᒻM)�Qoa�  �P�Ҧ��	ʟ��	�?�[�}�+Ѭz:� ��L�v3:��	�y��7M�&�������0S�<��cC�f�|0$��-(���[W�i��'��	�u�O�$�O�	('E���ǉR�1��dk@-��od�c��*�5�	����ɟ1�CN�hl��r��'m��#6���M{��B�h��?1�\?��Ig�	�hf��@�p���
b����iM<9�+�u~��'xB�'��30qB�
4s
8eH8I-�U�C@����?����?��B��a��e�cN�uL�I�ků5I����y��'U��'�B�'�!Y�ԟ�Y���D,E@=F
�.Y��Z%�iv��'�"�|��'��	�<�7� ��'
�g���VI&2�$Q1�\�4�	����'��%�/X�R�'��OԊT[���r�	^�ʤ�G)	/L$^7M�OΒOJ�d�<1�ɂB�I	a�ڤ�`�V�:a`����;`�7�O���<��.��n�O\"�O���pC��.�m)��G�^p�./։'��'+k"���� ʧ.��3r͐$>h%Ȫ�M�,O���!�覱۬������R��'�ހ���\�T�K���OaD�[ݴ�?)��MR�FxR�i� o����6�6�3��!%�6c�RH��'#���?i��Ο��'bެ� J_[��%��ذ�>cOOx���O��I߂_�AE�=A�9��R#{��7�O��D�O��t��t�i>��Iӟ$4K<d6a�!"����2#����'�D��y��'�2�'���Q�ȜD�X�9���PbR��vJ�>�L�9�?������O��OH)d�Ӥ?�jH��`�?s�؅*Ak]P�	� ���?���?i/OhH���Z :�ʩ�������ȠA�>M\�>������?���g�  �f#<f�:��i���$C�t��?)���?�/O�HJ2/M�|z�*�8_�n� 'C��`0�SoH}R�'��|B�'������䈠H�B�')U3g�Y��Q�=����0�	��`�	䟼�㥙A���O��B�ɍX��	5�Ҁw���[t�i��|��'��Vh�O�s�8.�Jb#��x�qu�i'r�'H剖)m�ꯟ��d�O$�ɉ�/��鳯
ox��S ȵr�v�o�A��>�S��$��b/��}��M���\o�ܟ�	�yA����ğ��IП���L�i��@�Z�O�����@%]Ä�B�wӸ�ĩ<����o���'F�P����S�����a,Lb�0�Ir"�5�f,�G�|��!>;��98�� ~Q&q�B�1D��AK�q�B����h�8񸖉��t嘴���G�+�(Y�
�q����N�e��#��t�H����`��P���w�4�	�/r�����e 4%��7�@+�X�B��� ln0����c�dd
�!n��!�g ��`�ūZ�V�c��@�+��\�F*�wF@`�����	�������ug�'0>��`��ϝ�e�j��6㚂t�� aw��R��YWl
KRr�IGOEL�!D~m§y��(Z[x5P�S�ja�L��N��z��"p	�E���E��-J����T�!�aT�Sd��<YW��C1x-b���ʂ�� �Ic�'��O�U�C쒷u	J5��5�t�)�"O�$�@�]�'4�h$�K�;d���c��ܦ���^y�:]���'�?�Th��V����H/bKt�Y����?���1�`�����?�O��=S �[�]-4��ݫf�֨`�W�q�~��Ť�UWx �o8�؃bLڈik��0a�L8"��e�U�̡30A��@
40ݑ�/G�!��xr���?Q������+�Ve{�|�@ysn�"�1O���D�XǮ (�Ŏ.�ԋ�VD^�F{�O�7��%b��$(���}�l�P�T8��$�<��^�/ț�OQR_>���՟�'��
f(H�b
�1W���p��������x�
�n�$Q��"6�?�O=�S��R4��Y(BV������f�8�'�r�* ��f�2Q�G�1�B�Ǩ�RH�O�Ip�eA>9�� G�	a �!K�tyA�Ob��$ڧ�?)�J��_��%����-�p�F~�<)�.��^<IP#�ŏP�ZL;�g��hO�I�p�'�����*�P�zq�Pd���TIhӢ���O\�����ʧJ ���O����O�nJdT��B	$W,h����S7sN�	��bI���$��d!r��|���+�p���	�>Nx����'��<Z��J@}�ƈ�!����}&�S����`D���t�yk��C����'� 9���|r���М6����O#dY�]�B@"b�!��q�2����ʧ_;Ș��#�0@��	*�HO��O0˓�ta�~T~�0D���t)���Ё|{�L����?���?	�����$�O,�S�tk�P�!�&z�0��!l�1`��!UzB%M=�O�,�� ��E' 92'g�G��ʇ���n���`��Z����ɝ}����>w���S�"h��B���O���������G��v�
1U�)Ta|b�|B!�{�+�`�6$d+CN���'��7&���Owұ�OD�C 0�%��3� �sd
Àe�'v2�'�R0�����:#��U;V̏� k�6��?�����j��pNB�Qw�Q�`�x".C7j"�q�A�3qKH��7�i�j%acT�B����=Ib�8�R
}�	㟴�'=��M�Cclz�̈́�=:Y��y��'.�y(�=�^�j�m��N�Ҕ��x��}Ӝ}��,�7Sٞ`b4�Ǩ�J�����O
�C�U:5�i���'t�S'P�~�I�i'N s� Z�w�̺Q�%&#J}�	�4C��ǵ�c�P'�|�S�TY>��b�L>+P���'�)�Ib�#>}��C=HS�䊇oʧo{4�
/:�4��d"�h��
�/N�WL��HU>�	� ���I]���� �)�Sת=�æ�1\�� R�M1zB�)� �20l.d�&m���_�fHr�;��|"p鉗k�:$���H>3�)����)2�p�ڴ�?Y���?Q�L�3�q���?Q��?ͻ�^<)$�5's��B��)=����y�2��<��gP�Q	V5���*�n�@CC�T�qش0��	�*��Yh�HI5#� H�F�e�.��<q�F�ʟ�>�O�Q���7l��.��\���Q�>�!��}�J�ڔS����z�-����HO�8�d\�_�(��GK=8R�F��FΖ�0��۫����O��d�O
,�O��9�����&4yu�E1��r\
Z`����B,H��Pq6b�K���+w�"}=h  �#�O:TqbJBj�h��ܛd8Ή G��bb��' ��'�	ꟴ�?�vK;?��Ědg��>A�j�<iv E-�h	�`Ä�&� �'-�j̓f���nyٔh��6M�O�$P�*d�����,(ˣB��z�D�O>=��J�ON���Of�Ҁm�(~�Ƽ&� d�?� �+ɛER�Hw�/O�y�`��EĖ/��`@�B0o6�d��*�)��)��[{�\���+H���d�O:�m�� ���5f&`@8աŠ#��f�Ryr�'��O>]��M�"L�э�23�4X
�C"�O*�E֦1�w��YrD����E����膢��M���'�c�����S���e�gOE6pn���/&�����5�p�"A��iX���H���d���q.����Ղ,T���ȓUiT�� �P1Y4ɻ�G��s����ȓ|X0%���Bȕ�"h93�͇�78��eAU�A� �R�B]L�ȓ~RaA�.�p"�BFL��`Ї�5���(H`���a Z'%L�ȓ�h�s�h���D�a�KG��Vu��~�b��Q�߁J:� @�K�5nu�ȓ'�j���� �J^��M�)f���ȓd,<�{b�$l�����~Ϯ���F�!#,�j�T�
���3�蔆�Y�b���fðT1�A��
;	�Ԅ�|W��sbH�E�`(�`��g�H���L^-+���JD1نn��F���x�Y�q��?gT~��`��DHvI�ȓB �d�P+Lc~����[
>e^��6�(�q���+}d:R�O�=��%��_���k�VY#���c�)�d=��S���T�6n`cdF_�
I�ȓ@2\�2��ӋC��1NH����ȓ{�����G�g�|�1L�K�(݆�d�8�Z�L%]�5��	�sF�9��a��q�w�-gM���!�͜&���ȓy�XTv�W��q�"�H��5��(R� D���_�)����>7���ȓcYYIC@�;�X!'�^B��q�ȓ!����3�śqW��X��A�/���Y��9�4�B�RtA�ņ-f2L���IPQ|�"��9�?S՜!X��j�-ڕu|EJ��A�<)���.m�8k�k�I�$�I���C��:A�;�
D�Y��#}:JW+;v��ԅ�h,Ҝ)�
C�<0kГ(� C�E[�9ɷ·�Y 0 T��h��$�st�ũ���Q;����.�D�!�d�0_�(ppS��7m<��sk��N�B�3*Y���X؞��@ND o��r@H��QZ]a�� |O8x���B����4R��ƪ���Z}��.�'h��
����p�U�ڎ���Yz���?��/\�5dѻ��#�'*�$Ce��w&�����
I�)�ȓ,F,ó�i��1��QD�%�'�#=E��G�U
�a���̙C�.y� Nň�y"K�'X�`2�&9�% �n�'�y�kő!S:�h�iC�V@�;$���y���T����b �o�xb �]��y
� BT� M�()1[�ʩJ
D�!"OQq*��B����c��mXS3"Oʉ�Q.�(%�L
���
6�	"O�0�B��6s�P�3�B8�H��w"O4Y9�@�$[r���Ӝ�+F"O�y��U�Y��!����M�a"O�cu��	e>J0��
1'���'"O<�I8U�꽨%Ԭ �p|�D"Ot�R#�L"�^��S 5��q�G"O�+s�i�]������� "O���#-B� ��L
�-?y����"O�9VEЧ'�pY�g��\j"O̔�F@O#\���FJ�^���"O`A1����5Ԯ����}pX!c�"O�q;�ǰ<�}J^T����"O>�ȕ��.n�&\I�/�P
�x&"O�M3T��7u���%H�8��"OZ �Ae՝O�DU��� �{ˬ���"O��q5Lк6���C�ő��*���"O�p�FJEH1|���C��mx��"O*�(���U�~)�f�¯�>�a'"O�)p���&n�8���_�ȕQt"O�9zp�"ÖPSs	<��@�"O�@Q�HMi;,	(�Bލk�P��"OhM��ˌ�M-���a�8M�ER�"O��2�@&�X*#@�Je�ɳ�"O�u"!.��Jm�hn�6�z�X�"O�<s3n+��-�QL�<����"O��w��2D���f7����S�'���a��$�;{\�$a��VY�P���!�DI BmB���1V��fR�o��'k�X����ٝ3R.��ǧ˖\�(��]�@!���GG
��w�/ܾp��#zn�sp���>���P��� d��r���|B�˻�0P�b��S�����xB�ۉk�TP�+�r�Ѹ�P�2'�ƾ�=S�'�.G�y��	3bx̛�@�1Qp1O�S�{�:('$��X�׆X�(ۄ���X	Eٶa�ÎG�R�d�"��4�d)�@�6A������-:�X��-!�D�z�Iv��?�0$����9����FJ~"j��W���0�Ŝ�p���2(ҡ ��c?Y�5�ֹ%ܸ�J�s��ݒaG���cƜ=T�x��퉾$f�A�I�Y�¸r�j���z��j4��q#�;'hvy{�?�)�c`fY;g����M[�mC<��T��K454��%L���c�m1��(Ί�X�cSč�'
���Y�.Kb�{���v���8u�������2$�z�a��!�)a�ٶR��m�T�æÈO"� &(��B�,9�P�̀	W:T�p B�\$�Ĭ��Y��/ģ2������U�H���j!�g�IR��?�fF tV�EZ�B+� �3&��<AcmE�	�E�4�����bV�����$)�S
qm&���k�~��x�� >GH��Z���K�`�Q؞��gթ&�\�у���/��q#�@- �V�h��<=�����r!��O��SM>A �>����4l=&��c	U؟ ��j.<	�M%z�`b�� D|�)C��[��P�c��a��B��'�����ԥ�n�ۀ���x�t�����W��#b�F����U�W#��I��R�,�:���������� D�p0W���t�ւ{#��It�>?锥fvF5�� Nf�ԁЉ�v�O}��WԗyY0y#�-+���'s���CO>7�]�剆-h�R�17�^(^���qF�Ohـ�!<����i&8#���8:[< ���&�z�ē@NrQДϊ*1މ!�EC&]G��@�$%y����8r�4e��E��| DG�bA~�)�D�� V�����`?�A&�Y0k��$��U8��[GFҳ8�^�u���h6!�K-V'����M3W%����/��O��	�N�'n5Q?���M�LE�A�B�h[�lڽ��d���zf^4can���;��Ԩwh%�����{$�x"��66��vm�$�����E��y�Θ}9��E!�p��HZ���%�`��H;�)��������&*�H3TG�t�fB�)� ���To�x��B�*�u2 jܓJ�*9@��L��&J�9^��5�2��'D�T{��.sp R���
j�4-;@k������2)��xa��l�5�A�ϟ|�C�I�P`�@�AO�e�|�� �K op�B�I�dk&l&�
8� ą%i��B�ɫ>���e������	V̈́B䉋���j2N�!Z�d��(�,A	C�	ML��0O�x�t��hϘ%M�@��P��c��R��MRD*���aI+q��E�����������p?�Ǣ\�!��� eI��S����e[�
��^T^��4�'���7�0#^�	rf@ث�\���Dޚxk!s⅟"c�����ɱ���~�BaRP똚Ȗ��u"O.e��X�J��)����.R�P�p��O�u�4O��:Ff��⇱�0|��,R;UBY*p��w�&�20ʞ|�<1$b?S����a�1!���"G*�˓?@p�AF�Ĝn����'��3�A�@'�L��F�9N�S�'�,���O�s~�����V?�pY����[�d���I5@�����犚f�p�+��Ι[�V��$,p����')�Y��05�bL��@T҉��'���,7V�0h`�׭I�,�Q�'�f�Gb��=�N���E�1�@��'@f�)��+� ]���.z`i�'��TQ�f؜s��(��ι���R�'���s����iq#���:�,k�'At:Ë�v=`��I�nq�P��'�ڨ�G�T:J}`��3i�eT@�y�'���� �ڣ���:4��5A��z�'>����Xp�Г�G�)I���	�'Q||y �@�h�8�[�L�2i�
�'�lɦ(\�}��;i��d+	�'�r=����:�:0��8lx8�	�'R8� W�A��U;4-�5t��E��'�V銅˜�c��i��dތ���'J��`�Ⓦ !�8Z3�2�vl��'����%;���q�勨+Nh�
�'�0���)�sܢ����M���	�'��K��9����P�ʡm�>���'$�h3
�+�<B0m��p����'*D�9E���4@�U��˺�� "O�\Jp�7��ٛ�k���^�J0"O��2SB�	5C�(qs
:$��0� "O�C�$k]P�*Ɖ�$d���"O�쑦���=���I��C)%]�!��'j��#6&ܤ
��Ta䆅�:s�I�&�4�J�2��ŠD�����>��x��؋<�`h�g���,��@6��I�;Ny�	�hҌ9;�I��T�~"B�@*{5���!�;2�h����s�<Q�'�R��a�Ǆ؜4>n����,!p��a�N4|D��	��G�_I>��}�I<����B�~`�ҧ��>a֔��Ni(<�b�ʢ}�����d��N������I#�p�w�Ϯ9G������K�tp
˓6�ؔ�"j�<x�l��g�R��}��Ɍ}���D��"����Tf�V�t-RB&a&e(�HJ�~$Ƞ�L6$��QQd��,tj�n�: N�� �.�>}D4�@k#�
c?�`�a�>,G��T��>s�i�h-D��r1��&'w�Tp���N��a��O�O�L2�'Ic�Z�L�"~b�@/fN�<��[I	̙w�B��yr��d���E?���GDL����B
���o��<Q��%6�x��.���x+1�\���X�g��l����u*~-:�	��+�)ѹ��x���D�����ޝrL��ن,�:�yBƒ! R.�Z D�L�C,ޫ�y2Ŏ�1��k��T�` ��3E�P��yri��5��3��4$��H�����y��Dp�Z=�r� "���IP;�y
� �@i%-@�X�,D���&O�0d�"O���u������ H^�Md²"O�<QgK�86	|�J�F�#D(q�"O:xAФ[O {�Œ/��3"O��rd�ԟ=��K.�<�"Ov�+�d��9��u��jT7"��=0"Oޤ�	X�N7��b�'W�3�.<��"O`�b�o����(Z'g�r��h��"O̐3$��)c#�T�0�Oٸ�!&"O� A#/���ʣC��"1�S"Oz���R�]�l����D� ���'I0*0���N�2E�(�ƴ��'o�(2��^|���g���qWJ�;�'�>8����l(��#��eI�=:�'��u�`/�0x?ޔ�,ˈ2�Q��'Ж`R i�s��T��o��-d�8�'�$	��ׯT��	覀ڸ*z<�x�'��D��Mدt&鱧�P����'	�MCU������6�_y��]��'�t32�UI<Q���Q	j�� �'s��F&�#\�:��[� ��	�'�-آ��I�lEk�O�R�FL��')��i􂋩d�ʘ�K�6I(��S	�'9���EKV�`{���A��H�ps�'�D�ȷfM�R�H�L���A�N�<�ӍУs�|p���MY�dR�q�<�q��8舩�5��A��Xo�<�k��E'��*�O3w��ĉp�i�<��D�ҴBG&D6f�(�ڶ��<Q���2!��i�àʍp��bpk�}�<!��1V-��⇌B�*�*�Dz�<���2&�8PƊ�}��8�djM\�<)FOُ:��E	�+�P;�@���Zb�<�����RUOS��)`PjĸY"�B䉮Fgb)W�˶�l�6�"O�B��.���B*<8�:Q��J��z��B��/dÒ��VCLlZUᦫ��[i:B䉢
�qe���<#yh�A��+�B�
0yV�V.
��:Ъ_9Kj4C�	2g�<��N�R������&P�dB�I�$m�!k0.�4̩7��l@B�	�9 �((����l���Ǉ�-x��B��mV&����A�!��[se
7K��B�.c�X�ٟU�����UՈB�I>�,Xa��	F�����,"�B�1xL)$	Ƃ�������hB�I�5��E�l��t�S�ۮ�8B�ɩ�N�eW=��`���؛snB�	;x(Lc�E6,�C��zw>B�0l�$k&/Ћ���J�@֯;�@C�=)�����^XM�����ҵ%�B䉧 �"�W�Y�GkF܊B�I^��
�F�|��EZ ��N~B�	8k-���̆��֮_2f�DB�RGX5��� U��ѳ"-��2QB�a@�l��@�6��r���8s�C䉣�B�����=Õ��n7�C䉭YJ���(ʊB�8u��P�3�B�I�t���K�,s�8EK%��N�B�	�q�X���9�N$A�YӲB�"F��(�EA)K5��GG�#J^B��$0&8a��Z�T��@��C��M�2B�	�5�"����u��H�@���Y��C��27�YÂ�߬Q^$�Z�7IK�C�)� P�h��=u����UǊ� �-�"O8`��%H).4 �悚KZA�r"O�]�#+��C�����*V�W��lb�"O|��U�5{
���J�d=	"O֠�狂H�:\�$ǝ,]u�"O����\:49!5 [w�0��"O.��	9{s�����f(a`"O��T��}��j E��dS��R"ORЈ@J+腣���43Ih<*"O8}�'o�5]���#��wb@鸇"O�eK�(�;r�ڔ����hC�P�"OdM8�ʳFa�X�f.܁�"O�p���1y��|0��tZ5:�"Ov!��L��Y2w�B	����"O�0U*L�s{��#��ӘN)�XQ�"OJHB"@E)9��Y�e�W~�%*"ON���S�4P0�9 -x�"O��� ]?>&A%�A��19bj7D�((T�׆Kx@�a �
29�z�c
8D�\��-L>���Q�d Q��6D���W�K
)�x@�vaЭ��Lf�"D�03�F�7DFU���ͨ;��0� 5D��*%DH'O�p�K5��<r�0y�-D���t&K�I�Z���o��L�`�+D���vl�S�H�2ĉW�t�� ��F(D�HsҤ�/G�`�+���$��� �.9D����<7��XT�Tp�����6D�����9H��ٸ��?T�f�c��2D��+VMJ;/=di���Z7Z��B�1D���d�[t�L�ң*�.�Y��3D�L���Cv�H�0��0EN���!�1�O~�Ob�v$�R����(�/QX�Hi�"O�|�wc[y� �Ibm`*
�Q'"O�[��Fpb��F�ÜuhU�S"ON�G�UN,����I��1"O��#3̒\v��a��Z�yj<Q&"O�-�T_�s9����L��aq$�'�l�̒/�bI a��<!�LX�'�1&��R�v�( ���{�h��'�|E��Ǝ����@�(�D��'& )5jO��F���� .ZƩ)�'�؜J�$	*p� i��qߠ`�
�'e�`!�@.����Gkި2p,%+
�'ef��6�^� ?v��U燂���	�'#\�s�iX5!�#�E��U�	�'���C����I��?����'��� '�K�u@~y4�E�}V@9H�'46Ĩ�F,Km������=xj�,��'(
�(`�؟<�\���0�ԥS�'0ҽ���Hzd+�J�wAx�'u*�h�쎇.�СY�m�:s����'I�t�����J�0�+G=�J�s�'�����!�ZQC�.��:�@A�'���GN�!��$�w�4�����'�$M�.�'F������T�4=�8 �'΀\�'�[R0lCV��0�V�Î{B�'�JX��ꗫS/��CdLĉ?��ɠ�'f��3��M�#8z���R4=�Qzߴ�Px���4G���f�@�-=�q��!C�y"g�)��\��b��*�}8�D��yRč��@y�m�'$�ѫwk���y�ӺW��x[���r!��a)%�y���-t]���C��{�����*%��xB�L<3�"ei���T����Ƀn=:����� 2�iu̠�~�9��A�?.���'��O(]�X���h�B���#"O�YID+�:tA��ɲ�ٳa��qs$��6�S�ӓ[�p�- �F*(�1CȈ/�B�\ ع���1tFډ°	"~�B䉀=��tg�L�V��������*ٔB�ɀdh����
f�q��#A=�8C�I8#0� A"�,U����5_=6�B�	��z��N�y����B¡R�B�IJ���!L������A��B�	\�,�WI�������H3t�C�I}L\ˣ�t$&ͣ��� ��C䉿N�T���
��Ea&U�$"�<FL�C�I�ڈ� v�w�8iq��f��C�	 <ƌ�0�W
��a��7g�B�I�4���`F�ԤTl� �v�B��]k<
��?g~� ���9K�B�	�mp�����	JvxP{%�ʮx@�B�I�;gKp&P�m�v@n�H�B�I7��"Tgρ'�Z8 �M'!d>C��u����ҭ'FT�Q�DJ�a'dC䉫6�P���Vt��y�4�F_2�B�	.?��e�`�R���$�P�B�Ƀ*
:|��ġ@F�N�����"O��(�G+I��T�ÀI��u�U"O��ۡB!P'V���IO�&����&"O�e���A�$�2��F�1e����"Of,�K�VĪ��K��FH����"O����	J�ty&h� ���Q�"O8�
EL�,D	$T��F�.~�n8KC"O���Ch��X�h����\����"On��dلf&�qAN6S�Ѐ8T"O��P�O͜^p��b_�c��'"Ov=Z%EĎI?�$y�U�\L�5;�"Oꐀs`- �84�D��8|H ��"O����+�N���K�, x�� "Ot ��U5��5�"���d�8�"O� a���`, �{/��2�-��"O�)�l>2C<�i�	qd��"Ov�8���NL�0;�a�Sh�(��"O�i�)�c?���V�@6nO^D�"Ov� ���k}����ş�?K��h2"O��Z��̀1�	��W��ax�"O�h�g!^�����%Ջ,��e�`"OZe9�]1?h8x�`��%P�)��"ON�pU��59�y��I�3���"Or����N�k�<�GƈZ��4"O�EqE� /���Yc���p��"O�)Pe%�$}*ܤ`P��5JĨ���"O~ ��)w� 5�'��,����"O�!-Q�r��k�@(|�ֽ�"Oڈi��t��k�U�Tn*Q�"O �Ƒ�v���$�ui,�1�"O4�(SFū4_:5x�eL�BRd�"Ot���J�ga�d���&ot��"OT����>Rd�itၺW�`��"O�H�'C���riуO�2&v*�%�Ii>�v�1v��B5�]?
��0�n7D���dʇnL>�@0"��h��QS�@;?�
�^��0ŕ�CFNA�dV�8a���ȓK��`r3�9���+	5\�,�ȓt���v�V'X���bS���9!`y��?`!����	vO��p���/.08��{�T�2�	FZ1Ǉy r���S�? p1�,�]�ȝ�d�<:�z5"O(�� @ݹHl���Q�B�OHH�"OB!1ƃQFs�1�#��,Y�P4�D"O�P�o�s���{@��.�HM�"Oxi࢈�l�Z�A��Zpx��"O��Iv�P�x���q"�]h�(7"OT��O�m�ƬJ��3%�Tc"O�#T�(.Na�g��r�:�c�"O�MkA�b��w���T�u0`"Oh��d\��w�O�+F�a"O���5��y����3L+�ȸ�"O� �,C�(�(��~nv\��"O��Z�@"��L25�:��6"O8���ǏQ�`d��4bFIy�"O���Kɱ:w��b�����d���"Oj�Aő��>�zF@��=���"O���?��-�$��O�"��"O�(K��J�p�v����A/�α�%"Od�A�P�MQ��u'J nu��zu"O���U�^�jtӂcވDo2�)�"O���+ģ1���A�)V2U#"OȀ�Ѡ��~d��h�MT�oF�a"O2sl�0�8���aծ![��"O���'����Ph��O�App�r�"O���%�Ĭ�Ѐ��%]8�)�$"O��K (\�nh"3�$ϖ:0�q��"O�)��-b�^�6É<>�p��"O�<a���:h�(H\=rM�8
�"O|L�dI�U�vLU�ؐw$��Ӓ"O��S3�JpdhL��D�,~<�t"O�-�:Jtx���r	����y"�1�E���B�+uԽ�����yR��4���bP�J^H1�E���ybG�E6��3S!�eR@4�7�V!�y�]>}�� ۑ�ن[ئd��ɑ�y��=M$�����̼^D$�E���y�l3MT��p�IǅJ����1�N��y��O@���ֈ�2@*&�jN	��yrCǱcB.0`�LV,l�YѠ�
�y��$wS< 	u�	O#�IU��y"����K5�Ύ-���eʗVG!�$C�T��EB��ZaH����)=!�ې"�<�*��9]R�@��;K!�P=J�A�a#+yG	#�共>�!��ʞ[M<l�h��0������!���2H���"į%<���_�>�!�dF!vzE�����j��#��T�!��4<��=�`A_k�
)yG/P�{y!�d�77c0!�M�Z]��7���;�!�Z�@.nHxe �
s� -x4!@9A�!�䎲|*��H��J�`�H�ڈ5�!��*ِ����=.2�ITn�j�!��a�N,�Fb� �Z�;�N	&%!���'�������s�){2�4�!�$����j��#% ��$O�4�!���͚��cΟ	���nE�!�Dه9��H�A��u�p��-
�Z�!��D:��C�f�}����6ʑ�w�!��4^�e�Q&��B�(�)��ԡ�!��Wzj�2��V�2�o�%w!��R�E���b0H)�,,��͑;\!��H�IVh)�,��`�4��r*�m�!�$��$^�b��P�Nui���y�!���2i�B3��ݮx`,@�
���!�� �闥�9p��D�慒)2�N�"Oa�
�9;� [�I*2��L("O(Q�u$�0���c׾<o\Q؀"O(\�U�Q�p�pA Ҭ��GO��Q�"Ot̀���+��`ô-�>Q�hZ�"O�8���C���	%�V�W(Np�"OCAE�H�c���t�!""O�<a�a>
�
�Cs��d{�$��"OTi)�ٗ0,�R`&_�Cf����"O�j��
1|�ղp$�	t���"O���D*eX1C#�Oat]Y�"O�@��$F-w�|�A%���o�:�ʧ"Ob�K��q����?2�FP�g"O���"Gο4gX����$S�Z`Zs"O�X�坳:9�dc[68vIjd"O�������$�bͪn�@a�"O�|·�N�"ʙ�P*71?��"O49����h��Z6+0�ݘ "OFDQ#B�9�z0����J���"O4�K��)$���`�Qs
��"O���ԭ���I���ab(�!""O�8�©F�NpZ���=\`��D"O���u���*Q�T{`��DUF��"O��)Q���ht��)"*�"M/�xS�"O �p�!Wj�v()2)��L�-z"O.l�cD�Q&����GP=,�a�"O�D��N�V[� *% 3��22"OP*2�(�61q��C�F�)�"O<A�d@�\8|�)��ǗF��u"O��B�#G�!��t���*���1"OL���
�?��|�C��r�r��"O.�@����H�V�" ��� "O$0�f���}���i%eC�(j����"O�Q�$Q2Ril#7*�ڕ�F"Ojɓ�ƅ�@�d�X�ɉ(1�R"O��y�`"`<^���I
L05#A"Ol�r�j
(I����DO	�Uc#�"O>��W�^��B9s)�0Y$�<��'�x$����9�(Hs��P1���'{� ��_9E"�eX-�:q-��'����.WQl��E��v�5��'�r���"Q��s��i�b��'^|��7$R�Z.�	Y�ːK���'F�Ԓ�����I�ˀJ."��'�h!�&'@�gr����5G�����'�z8�$`_�U���"�c�<C�N�K�'b����8\�maa�#7����'�Z�e�,Q����n�.A�ȓnM��jǅ
P=PP�n��a:�)��#�@9���ƆP��˅�+ؖ\�ȓyߪE�gW��!�R�J���ȓ.4:P�5nHc� ǦF�bt�ȓ5�n803�U�!o^���]������P�@��N24�3�^'{�橆ȓE���b
A�\ˇ\"��Y��"�R����>L����"�����SZh=q���H��W|6���S���ܻu�&�"�K�0[���ȓQ�� �dn�2E�:�7dO�6Y�!�ȓpE��j��/R���7�U[������)���PQ\��`�Xe�$�ȓ4��=�Ti����xz6��� ����ȓE�D�і��S�T��fN��|@��r�� b�M���aF P�U��S�? ^I�EG#f���B��8���(�"OFr��:�hhГ�HWvN��B"O�e�͎X�buQ� NjT<Y4"O4���D*OK�HPh�S�x3"O�2w�U�'�&Y#�ֳN�+"O�����'H"r�٣�I:m�Չ�"O�9j $�P��:�Z1m.M��"O�9��ԧ/�l���|_F�9�"O��#D/�14�D�"�ꀴ��8 u"O>����᮸��cL*[�<*f"OX=AiΊ	�P��a�D��4"O0Mʃ��1h����Hbu�1��"O���Ǌ�E��3��HffF���"On(@�� &E�`���W�c~$�R�"O�8�N7���F�R��x�w"O��)��
�Bfyʡ��S���"Oz��k��I��� Q�Z��U��"O(�Y�fU3l����@�Ėպ�"O"!b^|�&k":�0ځ���x!��N2E*�(b�O�$nҴrP,�L�!���^f�g�$P9�\�V)L�&=�'ca|��K�|��1
aC��'���P�ly�ȓ36��s)��h'A�Iś;ڥ��=�>�A�fV"n��)��iA�@Ȁ)���8�:'��Cc��!���-�Z���xҌhJ��A��U`�A��ͅ�=� � ƥhAN�d�
�Q�������� �O�!�rz���
wn�?��y���P6���'L�����K�*��ȓ&��b5��40 ����l�Jf8��ȓGOt�k�EΨT�X�%._$(rLŅ�P�J�H��  ��q�RI�!��0��D�ĐE�����6J����\�ȓ	F��!��:t�����4�`!��u�$�1����jiXe�L7N��'a~BmːSPې̈́ӌ-��i��y� ��)Ba�ZU.�����?�y��N5\�5�� J�X�c���yR��>S?Vk����E�(����Y8�y2%�|ՒQ��fK���y2�պ>$ij3�8xsD���(
��y��}@=`4`�Y��Yq W��y��?�}��I���P`ĝ�y)ςl��$K �*���`��y��̟?��е�C�y�j�P���y�I�An�4�M*'�L@ǈ��y�@B�Rb�)<�*��m.��. ��PA =B}0#%�2E��Ij�'��-���2܂)1�#��Y�� /Ov��D��S���7g]2\C���f� X"!��0S��IDœ�9�ڥ4J�|!�DG�Ki0��R,��"�Y4!���T����  �.�`��7!�D�[b4����;	 x��H�!�dN.&�@�� �t�pfe�]�!�đ�Q�EB!��`�aā'�!�$R�[wؐP��.ː�;GDߋm�!��A�DD�� ֳa��p�B�k�!�	[]d��k߼F���PQ��;4�!��ޘbVB�s�#&�P�JA�u|!�$\�e�!��n�o{4�8�lQ�g_!�d�7���ui�6Q�"QzU�Q��"�)�d2���XC�X�l8zh+��=D��J�@�B�.�7"��,�ĩ%�0D�� r� ���#u����s�P `2a��"OF$�al�8�8
6�K�A!��"O�˅)V2*!�̰�
�`�މkP"O����� Mx|1�J˺f�3�"O,\�b�L8vK|�f�x��5�'Rў"~2g��]2�}ZDd�V<(�a�yEB�	�rج ��gȽ�ڼ�%P5Z$B�ɨɶ+��ΧKЈ�ţ�}�B�ɼ\��⅄�;frƜ�p�֘O��C�	"h�N� 4L�5Pm1��0��C䉻d��=x�Ho/"5B��SbB�I1S`�<�6M�q� 9E㐈$�B�	� V*Q	7��Yvt���'l~�B�I%O �g�dB��P�Y�77 B�ɩ?�t<"�H�&h�b$����.��C��L� 3��=%`d1��Ծz�B�	"jI��`r�/[���Q���!]��C�	  �pHJ���=-h��� !��f��C䉴^���S���] ��ⲥ��=	Ó
���A�#��	mI#Q���Ͷ��V�"p���xqn�\
L����l9wC37��*J쬡��<���S�Q>trE{�`Y�!"��1��t�׳�]Ђ��M�om!��-l��Y��ߎ�t�K�Z!��UR��T��J�	X�&��S���QU!�D�1<t��r�HUu�����/�3N!�!dyY�a�Oݸ�1��9^E!�D�Z^�z��;k��y�C��T�!�dī&=�4�p�ɴ�
�VDǇUW!�Zy7f�ST�7��UZ� +�"O
%�&�S�Tt�H�
 �tݡ񄍌Kk���`
!My��0��F����hOQ>ixsQ�e��x�4�*L ����d+D��9� �!;4T�C&jЎ�ҽ��-D�p�&�Dw����Ǝ#�ڌi&�+D���Ո��F�5(0��>s�tPh��*D���$�:���Y�ʋ	mx�$)D�L�u�Τ*�$��bϊ� � 8��9D���׭ }�t
0�	&W7&��t�7�O��	�.��0slR
.��@ ��� �tC�ɘ�ݚ2��)�|"'�/]uBC��>Yd.��Ť��[\�l�BE��!��D��tEЬ*A6ɰ��_\>!��Y�>ΒA���hDl(s���d�!�D�����[ ]3rb���IM)!�ĕ�B`|��JܿW��L�6!�d�+sw>���#��«���!�DB��J��3�+�F���IW*UE!�D�*z*,*��� &�h嫅+O�G)!�$�>�Z�S�ˏ1o�,��
��!�ܠw������^R�H��5C�@�!򤅦6�B���u��q��E�!�$�VBR]�fK�2e�耂d��Z���)�'!%��yDB�"� ��(���/O���$��#�P0aF�ù��0C��gy!�D�q>}#b�3c��m�=?g!���9�t�ʢ&�&/XJ ��چ}�!�?t|���#�IH�a�ń+�!�ľ����Gƕ8�6���4;!�d�?:Ph����k���'.9L�!��L�8<b��"'��o��i�Ο�n�!�Dͤ^��]S�M�-��p)�|!�D[�m�urSB[	0�, -xf!�� `��䠁�x�E�a�8BP���f"OhCQbjV�A1F���GiT"O@[Q�5�X-��n�&�xDJ�O~��D��,\�%���]�)�*�"+>D���S��S<��ҍ�'T$`It�:D���A��b'�$�3�^�iu�����,D�d�B�� F�J"��>E�5�$�,D��k#�3B}\����;*F:X�V�)D��Tb��L�ڱB�l���A�"Գ�yB�cLȀR�F9Ō���lف��O�#~2�f��v��B��,��ƀr���0=	�	
_��G#� U�0�S)�r�<!��̧`@�Pj��T�IX��Q�	q�<�a�)w���c��E�x��z�Yo�<�b�V�4���#�`�n̺��q�<qv��#�h���[X�	a�c�<�sj;?��9���#L]�$���[x�$Ex�#�$�����W~d�Q�F�y����f6��񃀖?q
d�ʒ�yBk�9�١����J~L�����y"`W7<u�0�6� <�j�ӀG��y�7.N���R��2Bb��@S���y�蕣JZQD��Gֶ���G�y�S� �����GէR��X�� ք��O�"~�`*T@u�q�ܣTz&�Z�����%��G{J?̓1aVE�qb�70�^m�:D���1�B7��@(��7 Za�Uh8D� �R�[�POx3)��!6i���6D���N�#P��@BAJ�d�r�4D�*S˧KZ��PCA��`T���$D�h�0�E��� � <�`��2� 4��U5i���2Nil�c��U�<�Q�ر#m�92���h�z���M�<�pj�,�vm��Ǟ�R��(VI�<��-[0 )DC�|(�Y�C^�<�Pj
�<����D0nBE`�<Qҩ(ZT�*�LO�}x��7jR�<�(ڳ�j�S�O"O�t��,XG�<QFLY�wZz ��+�mn�)�KFy�'�ax��vD�W�]�9�¦X��y�(��pQ�s�C F�b1���y+D�w���:!-�@������y2��!;pT$����%����-ʸ�y����̸�$!�A���7�yb�L
"���s���א��-W��y�΂�CL���m�	2n�PF�ϭ�?�,O"�O?��Q4hx
qS��8=�F�OS�<���
�T�����>/����WH�<	'�,(0��� F�3�6���NH�<I���2�r\aRn88x�I��
G�<1$DJ&I��kd
���l��c�w�<I �W�%�I;`$�&P*�	�e�z�<A�jQ�3�и�#iK���HJt������"�V��C�	�?#�es�B �\d}�ȓzD$C�*����Rbg��tM��R��͸�F�9RTyC��d��̇ȓ�0U��N�@14��Un�i���ↈ�VSS����K y�ȓ>��r3�]�Q�l��"ư��m�ȓT�>8sp�
�G#.��4��)؇ȓ�͛�B?IB��@�	 C@x����x2(߀q0�4 `j�)�T��"jĵ�y�V�.�JI��ӳyG��2�V�yR�V�G�M�$-v��XJ���!�y
� >	;҄�����P��}Yu"O�D���t�XJ!�ȗ'n��d"O�Ha�d04S�ٳ�K�W�n��'iP) ��#+jPX��l��aG>���'F�Hw�\���;.�[v$�A	�'[Й��eY8a��=��g��T�̽҈�d&��ai�ȕ|�
�;�ݿ\/�� �"O`���V0�6���Q"n�\��"O0ț�L��U�Z �-�0����"O���1�9,s��q*J��P�t"Or�qu%D�W����aCK2�޴q�"O4��+F��D��b۞X�&D+g"O��A��G�ZC~"� ;�Z��b"O�0ʆ��LU9a�.���*"O���Qm�%��HVd�y�D
�"O*�c iF+ �9§m��RtRe��"OZ����[�gU 1�t)BI�R�[��|��'�L�c���X���)��W��%p�'��xV��8RY���6O&�Q�'b,�p��n���EB�]����'����G�5T�PӁ*��.��'~B���Sݜ���,�+X���"�'��KFԱ���s�S�KÔ��
�'��PfeԃGXН���K�J\x��	�'\����!���74?a8���'�z�*�o��ީ3���o�q�'��
nB!'�}:�EE4Q�����'I�$�mݛe8nY�ad��L�}2�'_�pS��%�,ȠɁ�V1|���'�0�Q�g��HC��t���zr�$6D��Q��.>p]�q�����E�'D���7����)
��܉Q�|�8pE'D�ȉ �"�Ztxe��}�D�v&D�x�T�C&U8"�8��ÂT�R�7�"D�ذ��TA�� ͲR�9���?D���>wB|[Ҩ��z, T �/�y¦ߐ"����GFH��L]��>�O�a4�C��@H��)-�fhzdU���'�ɧ(�+�U�V�ࠩ�K�;t��He"O����
0�歹Oά)i(���"Ob)�Ǖ�/���z�I�iL ��O\Z7�OO�Ɲ���	^�bA�5D�c6/ҡ;�4`�0�?^�6txj2D�(�@��c��a;�狙0�hwa#|O�b���"��'�0�Ӵi0[p�����=D����R�V���o�%5<�)9�o/D���� K�*�U�B�K���#)D�4C���^qp����B�ַ8�\���<��O0)��j�{�@�J_8B��K�"O����DO"*�i��*��LqKd"Ol�8O?	���y�j�j�"p��"OH1�H�>*qt�k&�R�!�B�;�"O�SpJX-z�l���ʈ����5"O�̃fZ�z���H�G�����"O橢�������*c���k��I[�O.���'O�.���k�*��4u��j�"O2���j]B��b�ױ7l�\�3"O�D1��Ab� �����\�02�"O�E�l�`v�N2`�22��#r�!�d�'�r���F�x�D��0.V&�!�ے��tٰ��J�f�%&�!�D�T��-9Ћ�?S�������f�џ�F����2h;���Ci��%.6�A��V��y"	k0F(�e��#]Б�4�C��y
� H���/O5'd}��c��-�����'n1O�P���4<��`���{Ex!�V�'P�I�pW�aC\*"m��;6k�Uv�C�5tL�C�!�#|s��#��|�C�;n���;bjs߮Yk��h��C��>/���&���F�Y7���Ms�C䉡ou2,��HO�7H;�BP�z!�C��=�� W.�V���F�f\,�ȓe목b"V�=n2�)��K�^��'ja~�.S4�!��̩0��a�dP��yRhʌW~TKv��T�a���yȊ�53>����N�t�34�;�y ��^ɰ�%M4��yæ
��y�
Ր3K���A�
�p�P�"ڬ�yB�����hC'e�rѲ���<���dO�V�*� �*�4g��i!r�A�{2��f�Z]��3���m�o�!��O�L���,����0l�59���^!RZY�R���(��!�I�j/6B�,#3ZP��.˰7�E+��J#X�B�ɉ*I�ڗ W�p}QA��r�:B�I0U����	�u6~�A�G"t����%�qz<��uc�w���b*ĘM��C�	�z�5#�n�:2Q��{�E�dzxC䉟69��DS�2r8�B1��
Et���;�	�yԄ�:E�'k�nE:����HC�ɨa(p��7��
������nbB�ɇy�v��"�Z�Z�d5Z��Fd�B�ɴur1K�瞹 �����B�I�2�1��gձ+:�#���6Oz�B�	�s����M�`��dKBZ�B�ɂPܾ�p��I&%���`�E���Du��1vC�3�
i�gǈB
a� %�D �O�颁B���f�TAے�~� "OJ	��#�JvZ�F�_
��(�P"O�yH"O]��P`��L�a�,I7�'��	�h���� ɻX��Z���<6�B䉿<I,D���N0����V�L9D�^B䉱i#�a� �U0��q�o�Q�JB䉩f$���	��3���XG�V�	�B��HLH��qN�+�d���%bB�I2���w�j�J(�6��01|�C�I�C��)`����4���pU怱1"���$!�Sx*�ʘ-H��f��:	�����Y���pW�&�$��U��:0j~l���B��PN�&*�:w#_�o�vM�ȓ;aFd���!�Y��HS�%4܆����إ
�;�����'^ڄ�ȓ�Ld[W�U��j}KA-D&9��t�^��e�WD�����<'<Ņ�|F\�f��.С�b@���ņ�}B��+��X=!�쥩���x� ��ȓE'̈H�fA�@��`��v�Q�Ɠ
GR-p%��Z���qrC�20]K�'�i(�%���S���%�r���R�JUCS*S*��gT������/܊� ��c���񑀜# d&���8�řD�~�b�9t�G*Fh ��'3ў"|�R햪yj��&&�=#�@�I'�7�y�'ʝm�p4s�J�e��+�H2�yr��:(��X�wHR�����֋B���'�az��h.��p&N-���	Ё�&�y�d��wnhT�$X��3#V��y�愎o��}�"떡 �H�h"�M���O.#~� \E��T+�FQ$�D�DS��'����0j�� ��^
^{�Z�D�(��C�	5W��]p���52P��2�����C�	�8	> Ů�4]2l�UO�""�D�=��?Ɏ�J�<Ҩz��K"E̉(V���
!��35Lk'�H�w-i#�^�%�!�$ b^@P��I�~_���gB̙9�!���Q�
�cez�i��ܥQ!�ǔ\�(�bO�_�r8��'P�9!�d=cv(;uD�W��Q9㨑�A2!���	ܐ y����g������g�!���ZvJ�����khj��H93�!�gb☪g��"|�d�Q �!���5��@@@�2/`����O�`�!�$��mZj1�3~��@@�\?�{��d�
	�ڝ�T��wa�9`�n�Q)!�$�'�mi���3#�8H����H!���ƁZ!ȑ� �/P���]�i�o�6�01��+�z�V��ȓkl�蛀�O��:�2凃p� 1�ȓv��y���sn�:��͢6D���R,�ekF��ON�1Xb9D���f��-v�� ���
���`��<���S+Ml�3F-�$$tu�4	b�C�I�FKV$�b&�72�T+ )�c���=ç����H J��h�e"JS��=��#o�}��E�"x^���vȅ�i9|نȓ4�g��C2���^Y�ޭF{��'!?I:�߸F(.u"1���c5D� � c�6�~%�7@D,V��S
/D��hW������1�&�u�PF�1D��6Lݲ��p�b�6
��@D�/��$�S�'�bP���D9���Cwش�ȓj喐�e�d����[�A��	�РC�Z�H;09a"�SN�ȓt���S䂋13��8�O�n��X�'ў�|��"IC/�q�����zx�,Gxb
�'h�z�	�_=�XP*�����0>����!�ڄ���.^�HaX�e�p�Ib�	`�'��E�D�f/�<h ��P�h�3"OR8���X���yІ3\֒�U"OP�8��"#!TiFkE:nǪ�("O�� �D�0j��I��k�*aa�"O�|��ܘ3M.��(O�0�� �F"O� �휤!k�2����0i��"O.�Q�ٸtE���tn�Z����"O��CQ"ֈǮ4�-ݥx��=P"O�0&��/&b��@�ŁCJ^i�"O��+E�,84�7��`9E�"O�:�ˉPĔ�0tA�PX���"O�� lB6m�B|1�o�;P7�҄"Oj�Y��	J@ʃE[D�|�4�'C�I%[@���Fѣw @"p�G�rxC�I���E�T�Աc���Ƒ�//bC䉪����E����Yz�hˏl]ZC�ɫ-$e�	�h�ҥ�T?j|C䉖-9�&��&r����"�����O@㟤�I�&��"hV1�!!V��-0")5�A�<!��˹c^�U���^����!Ue�<iU��?p��N���@�B^�<i����I�Nr��_N!��P�<���.$ b&� >���	�O�<1v̘�<�;7E
�0~��rD	Id�<�� B�/�H	j��NhL��)�M�^�R�Zyb�� �4Hakǲ$���-f�Ͱ�"O��[C��C��e��E	!}+����"O��q�폥�Ι3��>����b�'��h⅄�[�}���%^���D0D�lH�lݔz�^�H�`�R!�cK/D��Q�b��qRI���W
	�U�0D�8(�
 -M����a�A"@I�.���?���O]&�x�) X-�#*\��V$`�'S�A(�,�h���)��I}�1�'��15O��8UI3nP<5T���2�)�$iS�xg�B��05�)hɍ�yBܻH�*��P炲 p�m(��ҿ�y!�:o�qz�̐.!�6 �B듚�y2�A�jT��IЭ#z�s�C�y2L@5e�BƄ�o~�i�a���?�	�'Sdq¤��vf�1�0c�2��0�'��1��F������k�l9�'b�E����WY��C���
��'�V8�\7n��y�7Ё��'�f�k!���0{�a�"Q�w'xQ��'qpD���ܧ��A�e�X�r딬Z�'�0�Õ�øX���#��C`!���'�Z�Z���K5, @6ǔ>W6Z��'����Ɨ5�DI��I5d�v��'{p���FL�Rg�|���Gd��My�'uF��J�,ĖA���ǈ2���'/^嚠�D=X �kV�� _��B
�'6�0kG.����W���J�����yүЦ-O��D@ĽI��0Ѥo��y����h�h�N<B�F�3DԼ�yb+F
Yl�����6?�ћrjG�yRڱ'|E�E�_%\.�ڶ�E��yr�ͽ<B.a��̞�V�:tK�E��y�ǈ>M`�3��U�f��Ǫ�y��&zE����c.f�Qnʧ�y�&��y���.b�*����N����hOq� ��7ǃO���Bf_��|��"OhX�U� �Lܻa㍠��q����L��� n� [��:���
ҴI��'D�`*r��#;�D��9��I���%D�H�C畖t��(R�5-L�0قf7D� )�jN� �x�8SD�j=����3D��KR� ��������j��Oh����
rX�4i��V�k�倁�ҷH{!�ͱۮ� ��T%~a�]��"Wd`!�$Ӄ���vaU$tC��D�Bf!򤁧0�J#I/j��iZ��	S!�ĕ�_������MQ�0�Vf�#&!�݀PA �Ո٦O��-[�8(�C�I�a�80�V��/vy�9�)��ZzB�ɋ(����RJ�#a���R-Md�C䉥k�x��'���!:���D6C�p-@q���Hy����6`^�1��B�I�'�P�Jc�2��d�D ^*BzB��=%�ْ��K�!����U@�~GB�I4v�~����"S�ƹ#��Z�]��C�I���,��$0"���ì�o�C�7���H��t����wʇ*R���hOQ>���#Ķ`�����Z2l�\���>T�L۳�Ӊ)��B�l�G��7"O=⃯X *f��� ��N���!"O��p4GF�A��]1w�I3�	��"O���*��HZZ��,�"y���"O���!ћ5����X�@����"O� ����.��a�ȭ�a*ɦ?9ܵb�"O2�Z�E�ߔYR�H��~��"OT��&eǉF������ ᘩ��"O�4���|��]��.hf�0Rt"OF Ѩ��L�8�.X*j���"Of�!��@�����9y��s�"O|�-!1�U�D��^�XM�|��)�S@8tm9�Ǆ<Q]�"��Cl���6�,�@|����	2̨�*�);D��	T�\�Y�P�[����2Y��k� ;D��#��e�Z�s$.� h=X2�8D�8`uJ&7�>q��B¥C��Ԡ1�4D����Z�Y HĄ�=��|��A.D�<�t,�/,�Ӄܤ6�pQ��.9D���mP�}��c��L`�Ͱ�a1D�P�[f�.���W�uG��3Ui/D���a͔
^r%X���38��3s�2D���Ԥ\�K��X� #п:���Ӈ#D��cD�l�,�sd��3` h��v-D���I�\�V!D�`*HQ
7D�����˺Q3�K�c;G�h���@ D��X%�
S}$�u#L�E8U	CĠ<����hOq��| �NT�C�P��@�E�t%���'����=�r�����-�\���
O'�`�ȓVAx��f)�)�T������u���D=9�-Jl���&G��ȓU����nN�}�Z���J��x?v��g6��FX:>�y��΍7zL��s����v��{�)!�h)/��ȓzc(ĸ5�m�� �%�բ��ȓk�ܽZŔ-*�
$�p,�_$���^�j�#��GbQ	��X�g�P�ȓt��5�BO�($T%�2<�<�ȓDEl�E�H#(��;dF-�ȓ!���@��	A]�Q.�4b���k~2�O�E���2��Z�Lmp�^-�y��Ph܅ˁ��7Y�r0��#�y�ǻ
�.TQc�[$MX�YPWđ+�yB�������D@8I�&B�yrcH�,<ɖ@�;>\�0���U��yr��>J����>�ڰ"��?�y���:2Ӕ�UD=�Ы����y"H��~�z�8��R��C� �?��'�azrb��9�f�	�ET����-�y�j�d68�H�-
	`U� su Љ�y�h^U|,U�U[��D!Uɝ<�y��55�:$Q"FnE���y�LU�S�h�i7"�-hwR�[UL�ym�;D��1�N�]x�'商��xB�� 7�4�Q&��n���r��P�!�D�;p-�	;�i�*e:�٪��L��ўX��'+�hHEn�.�8ـ`	�{.B�2H��co	` �q!F�H.	
�C�ɎJ��X�Ȅ���Bk��
��C�	'f7�1EcN�e�VLKǍE�B�	%Y��S�G�BN0x3��qxC��F�!�\,1U��H�@��%bC���*�q��'"��hh���"fC�I�"��c& F�q����J�l��B�	�xXAm�n��qBV�n��C�	�?�pǃ�-�,�A畗i�C䉆-�Z�)��[.�<(�Tf�B���~;gWO, �e���8C�I�w����e��1�.a ����/�xC�)� �����oM�	�(�3y�L:��$�Ov����4��M0�$X;Tܐ� �m!�V�7#��1�h�_@|����a�!�������n$r�R�-�9r�!��/|��4�3d��#4 ���Ky�	�'�P��Q�ɎfX��dG+t���'.n5j"N
�'���'ދ9�����'9X��H�wad=b"̖�{��=	M>i���'�	�R+�$C��Z.j�7�܏"^C䉟= ��RC-Kp5<H�S!�0,��B�I�1�:MYv �#z����Y#��B�I	<,��hd�2^�E"�Wi�B�	�
[�٘4�P!*��5�TB��DאB�ɨJ�.�;��,���Ē3;Q�B�	/��X��l�(K�$��(Hq4�4��0�%ȇ@X��j�x���T%C�ɏ��H�e�6�4(#�dY�+��B�ɼ��D�@b�tbpL�7�C䉺WU���EB�{�j�)0zC䉲,>� ���C�:�Y�U0xNbC䉊0<�9�ʀ5k!���R"!��B��*u��F�-X��Jr�\�B�	8f�f��*�#M����.�jB�I !ƀ��OI�%���R����;��B�(��A����G���[�!��5� C�II`��c�+0�`�`�Z�C�	��� 2���:��� V�WtB�V��q`�/��7����
�Gf.C�ɚF�X��(�����K�M�㟔���5\�^H�Ə�~d����p��B�ISH���98��8g��}�B�	���i��ܪU���1.PF�ZC�I8���s���&֞i�)͛P�lB�	�xH\�0�.��Vˀ�	hM��
B�I%W���V���	j��#�B�ɱv�d<�0N]-G�]re*�)q>B�9@ �A���&7ܴ��	�
E& B�	�Y��wM[8]o�`B�O�>'@C�ɮs�=;e΍�{���@'c�� C䉳h��!b
Vy���y�MBK�:C�I+8U��(�`��?q���̞3����Ĺ<ir�Ͳ8�@��)S� �WHΩ�ybFO������ O�x���K!��'�az�@ɳ?���"@�-|0�X*1���yB
(�f����V�-�0�Õ�yr���E0r���G]E�\��n���y�l�2a��Li`�I�A�����ϐ�y¬ܿ[��1�c�B�хI��yb��,T��M�BN�)�4�k���9�yB��-=�Z�k� 	 ��E��g�8�y��&_ $9A#�h;�R��y�n�
`ٰ��B� ��0!�Ǻ�y��vZ��#��!.���b��"�y��F�"�I�'>�Yxΐ��yboLE$�T2�+�� �
	A�F�	�y.ԝ p�z�.���(���y�A���dE����/*�s�b��yҀ�8'��x	�+��Qإ�@��y�T�qh��A��ۍ>J��'��yR��+z`�$�ϒz{��A����y��L�e	�Hw	O�yR�8����y��,^�j�Q�LS>}ͨ�sC)���y��F+"TJ�
������P!򤊜�a�@-C=p�����o׬V!�� F��Ў� ���"�j��$ѵ"O�D�F�»y��R���`��"O�볇���� ËK��
e"O�EBf΃KqҰ23��5̠��s"OXq��g�� Y(́`��0�2"O��hs�	�����E�K���C�"O�]X�iP�(\8a"ʗ�q��8IA"OPMrҏO�;�=�C)�&���"O0�I4�
�@P��5����"Ob�X�	[�� K�ނT�lp
%"O�t:��y{�<KЈ�P�b�"�"Oz��.Z�UH^�@@H�#*��Y�c"O��c�e�#V�)�%�>t���2v"ORA{A�b�b�*�.@*^ű��Z�<�c�OS@Ma�C«�Ȩ`�Y�<ْ��hټ4�P�'�hӁl�~�<a�m��c"��j@,�09�f~�<�ffN	�V<�CoB(�<(��c e�<�iA��j6��	:�\��Ru�<���s�~��f��i����5�\�<!���#����E�H-���B��}�<�F�ݨyNx����Z��,{#Jv�<�'���UTD�g�@�o�: K��j�<ɷ	� ��5kw��v&Z 	�� \�<�B�'W��Ysh�h��m;"A�m�<�����83wK̬L�r�B��t�<Y�e�q�B��ԃ���ʐ"�G�<q7�V�h�6BQ�v�F�"#��n�<����,v-n���d�p��"Q�Na�<A�Qiv�1����Г�Y_�<�4CL@����ԨW�N:B���D�<�uk̾e�u�Q(�#(֌`�iW}�<1p#�X����T�'�%�,P�<1��bx5��K@�7�L)��%�B�<�Biɭ<|�y�O*�:����N{�<��m5��DI���F�Z#�M�<�Ά���˦"U�Z� ���-�_�<�F�n��s��xJh��#X�<qt`�2(C$X�F(��:3R����~�<)�Y����-ݖx�Z����|�<��D.D�i�(�.?��rev�<a��:�8� 񮅭��i7nr�<���P#$�\1�ʙ���)�m�<�!�.e��굈ءv��ҳ�Ep�<���08޼��N�\�p�spI�F�<���ړo���%O�4_��UM@�<aW��h�l8ģS:<�P���T�<ѦF�3c����ӡdq�0�Z{�<��$7��R�cZQ` �w�w�<QEa
�jf�s`b���Z��E��I�<i�@�l]�
g�O���8[���G�<I��=e�B��Ȓ�B�p����F�<�g �����s��L#(-*���@�<�H��& ��kײ*�z���G�H�<��4qv�ɠ����oC|�<Q��1_P��S#�.4;^K�Bu�<Q���2uGE����$�W&�t�<�r/D"2�A��Ǥ�¥2a�U�<q׋@� �h�%����kתIw�<q�E��:Th!��'l!elѼPy��aM�)'��$N�p���7�4���j��-����A��]S�f�2�^,�ȓl�D���e�e�(�u'�#�̆ȓlNTRF&�H BLR7.W��S�? ��KfO�,ʎ���腯-#*8��"O���]�n�dHQCg+n��dZ�"OzT��;K��T����`��d "O*%��k�n1�A�F�
p j��v"O��)A�5�A���E�h�=��"O�q�D��P�Н4#.xu0U "O~I�PjV�M̞�C˾p�]Æ"Ot�(U�M�~Ͼs���(fq����"O\��+F�}� �Iq��BbH�3�"OҹB�lI71�8ꐁWSzD1U"O���߃3�0���EW�H��ac�"O��+tcǝ�lݘ���u�ޅ*�"O��G<��`"g�̜XtxX�"O���U���0ej�Һxiʴ�a"O���5bX�UP�$�w\$k�"O<mJ�C͕M,����X ��"O%�΅*~Y�=���ԧ V�`"O�싱�\0o�&��?/S	�E"O������Zh�2bB1f@���R"O��#C�Q��#T�V(C"�9a�"O}c"�A6	��ɪD�_��p�2"O@i �����h�T�֠~�3�"Of"7�g��G@}�k"O���!%��b�@X���ߑ" ���"O��i^���c�m��d:qNV$!��>S�m�b�$4th�{c`93!��6�,B�+NqBQ� ��F*!�$E�:�e �D�+$[#d��J !���>D���e��+�&Q��K��l�!򤍇cnĲRN�@6�%�G	��b�!�D�*����EX�* ���I6=m!�d��V��Z�� ��EE��$[!��fw��p7x8��9��W�2!�䌤�v���-K�j��q�$�)x!��FH��EJI�\dq�غK!�	|n0Y�A��&� Q���"-^!�$ڵH�9�&-$�ЄY)RE!��='�%�t"�p�#�_+!9!򄊩8F��FɌ��
�PKZ�2!�ؕ(���7�MP�ܐ���ӲB�!�Գ'>8�4+�)�t�3늜5!��	�L�p�]��`�c�� �!�$ɷp!� G_<�̙*V���R�!�[�r/�C�@�|ͲT��G95�!�܇"��z挔�~�N��f� ��!��F�ɒp��<��F�`�!�Đ�}�i�� Ob�����¹C�!�Dð)W~�%�"��AN��;!��c2�yCl�=�d��KB!�Ď�i���a7l���e��&^�!���5Mf&�s ���\{&�(���'�!��/86qUH�Q`Lp���ͮSv!��~Z�)�2��	e��*F�Ѿ\�!�䘼1�&��*�2����[�8�!�đ�C|pq ��Htt႓͈+E<!��\aT����+/R�/��|����ᆩ;st�� �X45��`�ȓC�8�#���!B#i�c��,Li�y�ȓ��k楐@Z�]0���&{�����@~���g��*��@�K�y�\��L��y��/�G浻vA��i\�e�ȓB|ĳq)��e����E�!֬���V<��c��9Vj\"7�BZ�p��' *����Y"�1"!+M J����S�?  �g۲x_N�kthC=Zc�t��"O,hb��*6�=�t�R60���Q�"O��ᦕ�'��-�nR��zU;�"O�}:W��x=�Q��� �����"O��ţY�%_r`z_'c�`ѡ�"O�5���)H.�W'��-cb"O�dA�%�	-��h�c�p��Y�f"O��1���XF)a��� �Y�w"O���D�  H)�Qm[!>�����'BF�'�6���I-gd�XW&��[,���'\T�g�ޠ@�>�:�a��H����D���G��g�iߘ�h%F��o���� �yr�+NP	�5dQ�`\8Q����M�ĉ$�S��M��m2Bܶ	����}b�܋/Or�<a�E"e�D=B�6d��Q�<��'&�|�Ē�g���[�f��
G������y�O�$��I��@4wJ�f�.�y��T�61I�-Wt�hU0Wȋ��O�#r�AU�B���T퉱8eՐ%O�C�<�E�h���!W�	1���*f�{�<���?Rd�,SQ���$���ǫWy�<��(��_�r��gͅ&X���.�`�<�@��+|�,��o�;_̰42��g�<�(��p*4�@�I��V�l}s�]a�<��� ��|�J��7i@�2�@f�<��]�3���0)�x�:���W�<��n@<M@�I,TB��b^Q�<!���I4�yp�kU+֐��f:T��P�������{�$��c\N`B�
)D���	��X��6:�L�!�&D��Q�F_�uVjDj�*5T*nd�*O"���͆@O�SWhGR�6�b4U��D{�򩙣 �B$�u��j�ukS�_*!�D2J��hW�,A����l˲0�!�$ڟV���A���|O���S����!��9oP�(�g�Q�5 �H��z�!���*U�$j��X�9p�sd��)~�!��8�m�ч q�V��ɭY�!�D�$�8@`��A�qɆ<!5� c�1O��=�|�ᄓ�C6Z�K%/�# ��P��j�<��@�ඥ�T��!6ehAS�P�<I'n�Ųq�(�<�b��&i�K�<a�DB�$�\�bʰK���Je��G�<a�����,%%��0Z��B�<�t��nl��Q+�����Z娏H�<qq�W�
$�<�E�O�q3�����]�<�5䝜-iH1�M��IcZ2Q�\�<���'7M4��q煦�
`Zs��^쓸p=Q'\�$�0p�f])x6Ƶ:�f�S�<a��\#bZ�-��Ť��╧�N�<�6��UQ��h%
\�^��庂iNA�<�dk�A:`� �"@� ��Nz�<�b�ՓgkB9� Ǟi ���@���/�S��(��\���M2K�j�Q�$�ȓ#I�`���{��r�o!�X�ȓ ��`OĨ!_��k�S�`�Rm�ȓ4H���,7�p���,ו}2"���	I�6��΋�,i,�y�=m�ꑆ�9��  +K?W���,���fDFzb�Ts�O��운H['3�<@��.Y2����d(�S�Dn�\��aV^�1y �����D)�S�Oɂ5�ˀ�e.=��Ǥ*L.����/Orxye�M3�(L���>:.e�\�\E�'�]�ԅX��%j�1D-�����+��~
� ��y�(\�9���0ep�h�"OR=J��	�T�|�"�
ӛ5�Ri���Iv���i:"Fj�LP?}��K�iZ�1O��=%>]1M��W␍�6`�=�
4r��_:�y	cdt�7ƌ�B
B�8 E��OP"<	K<YQC�b�h�Z�O�5���Z�<�'�֍RY@Y��k���"�$S�'ay�n�*�~�A��l����1�y�g�p2n��v��/�hH
$̛��'��$ ��q�	0Y������ތV[ ���h�?arX#?���S/� �I���
iӺ��p΄. y ���O��(R
�5m�r�CA��/���\���'p1O ���}���s��x��m�^�������y� [�yqgԒQ"H �'L���v"��=%?a�U�Ƽ;�e2W��1с� � `��U�]�jpq�!�xLad��K)�<Q�I6�x�Ș�������M��	����&}�d$q4Tk#A��:��x�HC�hO2��d�;L#�� ��4��E8V��#�qO�6m��ا�+��I�Q3rH�83�]&~���S�"O��A� W���s��/qа�1E���HO��D}���5�h���J���c5�ǫ��O��lc?q#W"g����֎V�V0��:#�<D�tI�	�j�b���B�=OK��Bdkx�4�'D�O�>y�3I�"Ĵ���)��p 0+G?�hOL���ڒK|lQ¨�	Y�Q۷��8u�ay2��3A�ȍ�CL�'����ۼ/C�I=.򼂱F�_"��)�\/�B�	�J�ZS�PR�n)� ,��z?�B�	�#~��)�;m����`N��B�	U��p�1�µ7��)	E���v�'ў�?]:@$�C��]�'�G�h�aX�n%D�l��$�'! �k�fкs�Rk≥���a�'rG�"z�LYa�(��A`~�ؔ`�(?w
C�I+s`C�o��Wڼ
5���	�B�	�$����4'�`�h��L8���c���'�T���J��D ���"[}��x��'Lɫ�픴j',#�(J�b�!��']40Pgʘ�X�цe�k��L<�A�����+�@ s��p�2TE{��'.�iӹ_l飒�lҐE��'sX�� �\$��	�X�a��݀�'��]cpƘ����Y��%Yg����'hz1�7k�-?�2����?Rh�	�'*(|ⷊʆr��ȫR-M=H��x�'�t��"ѝ$�P�A���>��'�V����>f��(2P��
ϸ([�'��PHb@ |�0�@�-u����'<����Z"V^�����U슰q�{�;O���Q���sG��J���b�;sa2�i'�V� 5>F ��J^!ԕ�gK-�y�H�Sd�ś��
Wu@�j�����O�~jQ��(T��P0Kݑ)���	��쟬��� �q����֚i����K�RL��x�pd�0�ܳ �b���&܅�K���"`锗"�\�F��O�b�mZB������AB	z����U��&J�M�mL8�y����{B�ñOy���a�4�yҩ
�d�EڗJ2�x!�P��y�	M�Q,�ڷ(��R�r�C����Mk�'�F�*R�P.@��� j�l�a��Y�D�'�q���K�-�-z�ys�o��d&��u"O�%#ӫ[ ��t�� 3���A�x��Hk���O�XI��I'����t;��+��� .�`ťOl� �C�,.����"O���vb�6S��`��)�*$��[�"O��K�LF�\�Re��hҴf(���Ox˓۰=�΋;i�*mS���\"	��}X���R����Op@I5��Z$�1�皔M�mh�"O�(	ňȩ;2l,$jLдdV1�Ox-����d$]�E��ű�HћybZիܾ�y"#Ϡ^���S�*�o"���ŕ��y�!�@\܁p�C�^�$m(Rk� �y��[�*�ӡkK�Z�Њd���'`a{�$t��p&I�]&8h����y] Aa����E5Om� ��̟�y�-��p�I'C^�R����R8�y�)�'��a���P��.Q��-�t� �ȓ~eиʢd�D�r�p���$��<����=3��L[84X�K�u�Ʌ�Bm�����S)�
u��K��`���>@���AW�T�Ѓ��;+������V�f��Ӈ�4RΘ��V�d%:���B�d�ö×*�ʕ�ȓqr��A�_�f{���^�4���ȓdH��ʣύ/x����M<<i`a��$��m��yax(��Ӯ|�I�ȓ �x����po�dRP�Ģf��]�ȓ
�X\�D�_�� ��,��sn���ȓ5�Q��*V 4I�|���z�
��ȓz� �zphǜ%�����^�\��L��r@���O��{L��t�.,���ȓh��0��(/�r})bC/`Y>؇���9Y���j��I�%ʰ5�:Q�ȓIN��p@�G�hG��tj��8���P����t��z3@�A����
}���j�8v�U=1G�q�*�e6����AԜ�PP��7e�M����&-,��ȓ��� lݟTP��hQ葦h���ȓ/b:�8�e�2i_*�Bl�!@��� !�݈jM�=��1@#M�vOHx��F,F��R �I1������2B��ȓ'��C��#M$$jǋC�Z����#h��"��6,p�lA4)S3gt������G期��,Y�ڀ/����x��8*ƽ�ҋ/Z�@'Q��y��[i�8m��E���1F�J#�y2��t��s���85 ����y�kR�u,�0��Ĭ$����ٰ�yb��1^=������]Ƞ뇍�y­��%A��c!�T M[�\��* #�'T�`����d�4�#⤚�}T9��yǕjYƘp1���u���#�y�E}��5�! �Q�Ȥx"	��yr��2\�T�۶dR�u�D��
�y���#��:2E��Hg$�y��
?``eBŖs341*��@��y2ETJ����T��n����y�f?%	ޥȄ�_�u��`��&���y���|p��D�H�b; ٢�)���y.� ���6i�� �P`1H]�y⢀:�F�:��՛���+E�y�d���Z�ѣ�Fx+Ƒ"�f���yb���*]���킟DӬ�RC���y2���yda������E��?�y"AU ;MR0+�%�^n���@����yB̟��B�ե^#��"�.�yn�"%� R�AD�U���@�_2�yb�[��X\PAGA�Q��X@�G��y
� >�p��8�����/�J�5:�"O (cP��'La�E��R�lʌ�"OΌ�b�Y A��!,γB� B�"O0 #�Q���p��H�-�sC"O�t�L�"�L�t�^&{��(�'���� L�H�a|��`@j\�&P�9����6㕀ΰ=��ӗ�l�2�	�O�<K&�à)z��%ɝw����@"O�y`bJ�17Z��uʑ�O�6����dC'L�l}K�/��Q8�#}a�ڀ$�(p�P�B >��$�Q-�P�<qQ!܊S`i���fǲy�B�$օؑ7I��
C�Q>�Y˂���-�>b=lD��FMAjɅȓR Q��%��X�xĪ���9D�j�)%�ДV�X�φ-H�a{�ϛ&0<���nV^<1ga�?�p=Ia@�e�U�?�Mr̿jL���\�4��}���
u�<9%&jV�D��$'���J�"Gyܓbsz	Q#�*7�nD���i_/10
��RbN��Д0u�TO!�d�'j�� �$����!hY!&�P�a�(6��'�D�D�,O�a`��X�D_H���G)s��c�"O�Q��I�g��ȧ�4BA�-�cj_5)U�(A��J�o�I��	�B�
�V�Au���%��l=b���T����-ǌ�?q��R)8���� ����g	N�<Ⴆ�5=��8YeJ��r^�up�e�J����@�E�;눟�LHu=�@)�7`Ȃ����"O��0�IF�iN�9�G�N�|Ј�"O��u�Iડ��e�b� ��"O@�Ҧ�*G-V�y0dІO���Q�"O�!tm�+C ���ٵWu�c�"O��f���h�"LK� v�l!b"O,�pţ�Q�X% K��j`��q"O�Y!E��4�4)��T��s"O��y7�U��Ș&H�#�@I��"O�l F//lk>m�&ǜ.w����p"O�)�4 �7Hp%0iJ�-�ʬЂ*OD�pG�G~P�#�f�W��-J�'�ּ@R�Q�?~��RCE^(E��x�'��L10ƕ	/�+b��PU��
�'`��1d+N;KL��A�=��B
�'5~��r.<HpP<���ͭ4qH)	�'���QdnO�Kg<ɠ��ݜsfT�R	�'v��p���j_n���J��a��H	�'�-�1�Q.l��Q��!\\jŐ�'A�)�D�y���®P�!SU��' wdJp�V��G؊�����)T��S�'(执I `Jdn��H>j�"���cvC�	Xlz�{�*��Fx ��¥5�H�D�n����
��ҧ(�F|cTe� ]H8��%	r=ӕ"O��Ҧ r���S�^7򪤱Ħ��m���2>���������3�	�L���҆+��M��TI˘u(���DL�bPq��U
3�Ё��鋃 TlP��~cR�c�ݨ����d��<�"�	-N4T̅���)~��(`ק�<'�ٱ�@ʸ�v�O]>aJ��%,h��RC�##e4���'�6#L�5�"A����."� �1�bL����,���B���s�4�~3ąt���S���(3�4�qʂ�y���묍14�MRБ��dd�[����򲬍%!�`1�*p��'����������@:r�@���o<v� �S��;�a}��	�u
�9 �_3/Z�|���b�\�3��//����%)�P}9��'!�z���0(T�X�O�O{Δ���͂�qa ��"����W�?b��
��`M�x�EO|��\>4�C��+#*(��;����?Ա�)OJ��Y�pS��͋i�v��MC�
<�Q*g�>�Yam�,=w�]x���U=D����#���p��-�Ԙ���%P��6g�
Ux1�bo��@"��'�\X��$Řh#v��1EЭy|����D�;OT��v�.Y�aF���Il�x��1�Эzx����9���XCOؕr�nt�q��$c�1�I�F=�^�f$��bJ�#����Ǹ1�� C�Ӫ/��*Q�Ƚ |�#�H�6�&����̠��$\\O��''pƜPN]v��H���(غ�Fz�E��:e^�P� 8f� ����m\f7͌H�? ��"�˷^1X0% �2���Gj�$#�L����"S �_�Q�H�~�'��Z����rRdrP$J�t��Y�4B�,�%n�I�ty�O?5N��9�AX�:�����\coH����υlDt��� ֈ]���Ļ��t���֜y�~P�Z�,��7˖:' ��@R�`.&���m�)z�d�{��.Z<}q&"{��K�0l餅�K�|q���K�hh{0癘z���d�1��}�$A1�2��D	f�r�j��a��=���ͨb|&8ʀ�,E���3v�nƄ*�'��
~�z�Z�t�p�0���DW�y�F� gf��o.@T�mS���O��*r�T���䒕m�(��e�C��-'�dP8�����)����K�H�8�AG;��JR��	���L��91�,D
/*A�ER.k��ϓS�D���⁐7\(�)�L��%-4Z��҂�Q�'2�8���8H�@A!ơ&�0,��=l�Y:tꊰ�2���Ĵ\Y��0BҢBut� 3�;>�LDÅ%�>%4r�'�2$ڨ�c�~RD�N.aH�y�g\Ⱥ�2���(���wą.>Zx�X����?��M$	�,#�P.�U���Ə�p�m�0p��хzb�pѩW�I�(�������5jȉ�/ˈu#���U�J��p<�1>,"��"���k$��J���FI�{N�Y��,أ)%���'�\8{�"��X�m�q��T��ڍ�đ�](f�*��D��A��P"�"��K���4�	�y��17��µkM�bŨ$���y���!wڰ���#(J�$C�yb$�9r� k�+��Q��%�y��R!Q����u�1 j�R�iZ�y��E�U���i���0�4�� 	��y��£P�F�,�-�� �E���yү�l�&�*w���dIB��y��Q;P��`�	�B��Q"��y�Ax6e�P�P1I�w����yBei�p���+�6�!D.\�y��F.B��e� ˮ���X�?i�bԋ^�	xI>E��虆����0�ٕH�6	��>{q!���H��%�ҤR���'���`��I/0�,�r`l�>(��y2��)��lH'&�,j:2���e���p>� /�&�К������'ɝ�t}�Tj^�2��ka
�{��~�EW(�z �V�8Y���(O��-�ֽJ@���T�0Q�̟�`K�þ'� �:u)C�)� �� �'�<�k�K�k�S�O�l��dc�B	K�(mn��aŖOA�PV����p�����Tn#~�ɑ���@�K�����.opb�"��L�5F�-�p=�ƅ_ �X�RӇ��k�F6�[�ڨ�+`�Q�Z`�l��M]
[f�ݻ���d݊Y`���a-�? ~�0E��.�N���AN�,�x�	�8��T�"A��Y�HZ1!�q��U�Ru���ФID�Jg��U~���N+*b�N�y�T>5	2jA6� lao�#���L4�=�HY�*�4�,p@���&�ѕO����4e�ސ)1L5F�X��$�ݎMY�q�A�ɐ��)��XBC��3J��z�aŝp�<]�剕�4�dY,@@!��κB�6�ʔ�2���r1�\C7r������Y:������#�'c $h(��'+Ё
�l[3v����T�>�DiR��2ʶ1c!�ػ#OF}�#i$���O�4���&S�؅xWj�8
5�M�p�U�5ɀExR/jq���'PjI������K�b�'F��X�F+�Z� ��+�eJ�o���� N�1Ĕ���S���ɜe�s�"K
KxUp����B�{�G'd��y�����H�k�O`XpB�MNg��F	G�K�
m��.�v֠�t�b�z,�L��Q�)L��q���	7~ˌ鑕��2O���E�'���FA}B��h�QZ��u�$�+x�^��g^�9�,��K����>�`ةD)4\O�H�uI	�D��i�V�G��L��>�$M��i��g$��")��� 3�iM���e��rMb�P1Jb<�[�'� ����AȀ�B�hH�pA3��>"6����|�C��%iA�J.��c�KD�����̊��U==�����(v<�:�D[�N6@��! �Op�{񂄺8+�;��׏��`���'��0��4[9��'�� 	��z`%!�#ӪJ�q��'O�@KgÜ�j2�3���E�h�8L�,R7�K�	��Ũa�'�h�Cv�b�%v�p`�hX�!�)��-�Zхȓ$���QE(F���"$�<��i�J�O`<����.@򵡑�X�'��	1W�J����P�����δt�B�		T�� ��=V��a#��Z>�Sň��M!�aS	1���S|���U��
��Ȑ�B�yM��X �+�O�ɢ/փ1P� 2�O���
Jp����U
!3rH���Q(����� ���6ŉ�-n�i����Ĝ+����mT��H��Ty|�Z!�8@*���6��J:��R3���k~�qr��]!�6(L���K'n.��ċN,��d��DT"M��	ߦ\vhѸ��ƚ��tx���Mݴ����&5i�)Q遇�!��+Xj��aD���8��)Cv�H�����-L�|-[gt�4a���S��1O�!��\ a���We<���'6��Y�ف��Q[d��y� A�0b!8�2$��h�4G1zA�G��$���+�=��Ȕ�d��D�Q0�<E@+ ��bHU�j�Ц�W	(�*���S,��`nS�8��!;�CO 4`�B�	� öe�����u�/���r̛�S0��ѫ�Z���QL�&Ϯ%*5�#�s��j�	��@��% �In5� D���@�
c&�H+�-[H�$�#@ P�l<�H�BO7BںUД�>����a �T��;�ɚ��0Cv�Z�BO&�s��<C����$B<$W��c��]|����cŤY��M�N��C�h�9�ZD���O:�Z����;LO@x�f,�a�+�l�1MϪę���;����-=#� (♤b��A�ca	nь1��c�Fs<`k���2=��s*7D�<ȰlZ�?)�h:wQ-e����"�����3Bȧr��Bvn�/,�4ؐ,�,��O[�. �?����N�����3���=�!� �%8x�7��J����ۀ�r"Cx_40AQ�l؞��w@�@.��	��F�m��� �,|Ol���@-����ߴQ;��K�&Z1��@rTVh��"��f��f��	s4�^�"��?a ��C,��>�'5E(�!c՘[)v��eY�rYf���XV(౬E�E�lᐡC	.o�쵈E���R�QL>E��'%�a�A9&w�2dS %��H@�'x���FK��i7(�u9��@�'7P� {��c卞�inXq��V�N��ѱ��6D�P�7��l��C�ѥf%���s.!D�D2%B�h�P� �*:%Q �>D�܃@^�0�A9
�� � D�tHtX�=O<�vJ�:h��Ds��;D�t8�I��E�¤����wBt �U�9D��`����f�v�%��Yxۣ�4D�\#���[1�|@Iəy�2�KR5D��)AM��/Ѡ�@�=UL�Hը9D��j�$��Iq: �b]& ��FA7D�(�`
�����wk^�	�ܺR�7D�<�&H�uàe�tA�6�6D��/0D���ׄ��]���f�
�r���)E1D��K5Cև���J��W�-@b\�U$(D�4C�o_�m` 	�!�W�O����H(D�dB0��:h��Ď�gJ��1ԉ<D�X�bʑ]\9��=x^x%�r�=D�x*��A(9gu1�(�%yTF�2tK;D�����D'��M��g^nP�ңD,D������>N�]Q�ú*6���%.D���E!J�A�|�VGA�>4Bu�ri1D���W�3�<4��-��Q{T��&f1D�����5284�1�v�hdk�%D�H!�/�lXk�/�\����<D�Hp��9��e`K!"Q&�#$�<D�� ��˔Tj0Yx��6�$�� 9D�\�@��k��!gU�$��5D���1!H�e�HX�/^���)5D?D��C�jܡ!	.e�����)VtXŮ)D��ۂ�̠��l臆�&M@,H%�;D��@�HѸ4l��3�
 ,24Pq%,D��&�؂L�&�Sv(�+��!i�++D����Ǩg�~��g�
95��e2D��rQ+!�R4��m�>z�<�F(7D���b�s��)�柦���Ǝ)D��Jӭ���Ͱ�I�?i�K�95!�D��nMLRF��<���@�p4!�T�K�*�G�37���6�H�o!�� h��R�ظ�(K�1��p8�"OB�z��1NT�J�(ԍq���"O,IA�8&�
��(
�DR"O�5Ir	4s�4�+�D�8����c"O�]S2�4�<05�H&A0��+�"O�Q���
4��T��Mɢ&�YqF"O�݈��O�!�d�b�[,����"OLi��`E�h�h���+Y�]|���"O��0��ܼf��}3�)N�_��s�'���{�Y7r�a|B��!+���#l?�X��`��=i�mG�I2�@��O��\�I(PɳǗ�/����"On<�"f�>IP��@�Ћ6�d�  K�Y#I�3A�"}�A��$��g�שG;`���.T���wL�k������L�vZ{v	�:|ͰI�fH����$�(�剴LMbM��ɛ�$1�Q�V"J:N��B�ɟ2������&i?zM"ƭH*GS4�9cK_
;B�\�VC�%�='.�;�p�!�Vmq"e�篈E�����ZO��{�����׀�I�>��`剭S=,H&�!D�����(�\i�*G��<����3�ɉ�t����7m!��D���y���,�1
%Kd%�yra��Lc-aw��60����4@�;2P����u���1�|�'��+��܌&!\q��M�sxP���'�@�r��K.4��)�j�h���.ԩ5ʰ�z��>�D��D�}y�m�d�O�1c(�C���X�a{"&z-�ͰA��ΟSpB��m}Z�jW(�IPx��)4D�Ԑt$W�V�fE� �)4n$2D,2�ɄA��M��n�O�8(s'NƝB�`t��B�$|���c�'�&�J�Ϋ�
�P�?$�܈�'���ĭT#j�� �ɽ'��m3�'�4�8�#T|�l�s"�</VLT�'F|�7RK1�� ����5b����'}�D2c�ۀEUT���^�U,��'�@��2��A@-��j ����'�B����
@�м�`ܱ \T��'�p�ҧ�C]{�k��}Kx�#�'ɠe��H�L�Px� 8�2���'=ʝ�c(��!ލ��C�
#�A��'�DR�D�L����o�Jº�3�'����I�,R�L�v��F`���'Xh5z��ӭ7�l�K�$ՋKAh�	�'��E�`��
�5BУ�.�>��'n�@�$R�֔3�H��{���8�''nб�n�$.Z9�R�C���	�'VZ|���=�r��c�ˬDed�`�'65h�D��]�r����� l��'�$, ��$�Y�j�3�ZtX
�'�$��N�4ꔐZ�mP��,��	�'_R�AV�Ոy:@a�`S�{-Np		�'���;AM�yQV��%\=f�L�	�'� ِ��1�e1V&.(
 �s
�'�⽠��'�`�
TĂ�-�v� �'�Z�:��ܿ<a	tC�7�����'5�Q��&�'|�Ȉ����6�,Q�'b@4����.).��� ��Z���I�'R4=b��g�jU���8[^�e��'��TI���	2X�	��E�S�zT��'|J47�A���z@n��C�����'�N�#s�q��t��d�#�N��ߓ|O�1�Ю��y��տX�>T��(ѭN�V� 	��y"@�#��}b�C��L\<����(��'q"-)d�ցo8�dF��よM��c�L�G(��c��̩�y�N� b���#BW�G�ĵ@cd�.|�Zf��/< v����|�'
H�"_� ��(�FΗ�.V�i�N��A��/<\qO�vx!�&��<��t��� W��=q�lPm�њs�ɥK�4��)� l����	j��*B�!����&�&�#�����~ڗ땆'K���C�Ԍ`��0�摸1�ҙ����7.�����/&�O`��q�4!��H,���)rI4#G��3�~r�ְf�X�3b�:_���p�O�!�e��~J�*_�� ��oW�%L�p27�I�'x�#䓼Y��8͓K&Z��  �O�~�ab@,ʐt�bj^cOؐ�m�#L�R��O�CB@�g�gy�� T3���) �B�*��e�_���%*��0� �?�$�U�#�p]" �0�.H��1��'7Ib��SǇK�`��)>v�Y���O�vy\���߇�a�@�F�j6�ܻ�	X���u����x\��Ê���嫇�~�p-�{:*����=>�A�ϋ1�:��ƅ\8��p�6�Oh�yeO
30����$@�9�s2��NU�c����?�@�Q8!n�T�20����t �>y�(�&(���ܛZ%Rػ����B�*DF�:�џ�h�?jB+��'�R�c7FW
>`ʱ��)�F���G�a�6!�S恠�n���Dmy��Ι���$^INQ���x�y�j����I<@P�&]�8���VX��`Dḑn�X躃�==�-B��F<�A��4���ѱ���u
���$ˍYk:��ծ(��d'�ρ"����0*�L�ڢM�q5���	�s5� �KYk�-���$K<l�K��v�a90
OXZ�Npur���7X"l)P7EA������~Ң[-����`��?UP��D~>eF��x,pl R�Oq��+D+=�Oj��@,D^��(��bP4	� ��@���z0n-���-�8:g��"��:2F^�<K��Z�G0��Dl�h�(�Ӹ}�ԅ�0��D3��CfT�5UC�ɓ���(Z'1˂�+�AR#/�B�I,IV�$PW�R!G\���Giŕn��B�I�����V���nZD�Ҁo�@2�B�	�zߤD�2�	��HhAw⁚�lB�I+;�Db��^?RbR����"�|B�	�?\t�a'� h�<�႕~!|B�I1
����)��m�@�k�~B��	���� ��X�!���IRB��BpR�j厯tT�M�RA�7�B䉺}�fH��N68��0RcA�,U�.B�I�~H�ͳ��B�5Ơ,2֧7,'*�d\<
�.�KC,*��b�x��v��qpfЬB%5��C����#=G�,)1���� ��'��)j7�ɐgaXA���F8PV̂+P�R0���ٝ*������eq� S�aрL��|���ΜXfr`� M�7Q
��Q�nN7N?�ȅ��%#cJucp��-j ��p��6j�~�<��(�'&i^]3�h�/o*��P� �!;\�8��5jX�"ۖ��Ýş��5�ӫX�qO?�����3a��0�LŽ���3LK�4\iӦ�
u�@�P���.)����'�l��F��9o�FYjt��pJìO�q�gj�i�|���I�\���8b�HJn�)۳J�Y^�d���!���$ƞ�8���E՟�ɱ9���5E	�]�BQ�d�ˢx��ܘb�2��5C��'�Z����VX"E��h�-[�Ꜫ��X�jE�A�F�T[����O�����X�3�u�%˞���|��Ϝ�>��s1I��W�=j)T�'��Y�u��;��K��N�]�)z*��$ �=��d����4^��&_�B�-�㩍lM�S��?!0
; ��R��p,�։>�4�����)*��0�A�j�ˍA��?��m
yۜm[6 �~�4S�bX{?ɶ�[����;�)8LO�- ��ўQ��<'$�S���IPH� 1?�UꉢsF� �JL�����!��+5|�� L��tR� @�`q 6n��0����8�K˧G'�bbJ�&I��H�ы��
��r4��%�e��'�D �@���L15h3}b
/E!��P)��Z^`����>{Aa�hx�p�cH�:�J���N�.ED��'�J�y�J9)���X��\���9z���'�������H�矜@T�X�R� �*H,��X���9�	,��P��_�Ȋ�*�3RKr1p�?͋$G�FSQs!AՓDpA��>��ڊ���(
דz�t�R�� >` �s���9ٖ�O�TG� Ly�9#��T)ζd��o�
c`��U�F�����w�R��B�	N�t�JvBƏex�I�_ V�ؙل
7}��Ծ����}&� �a��3)U�Qhמt�p�Ba(���$����A*�l5�)2�%bK(pr���8�a~r��;ô��SaS�8N�bt�B��p<���O�H��0U�1?�J��mL}�%�ķC���Q��E�<��d�Dy6hZG��)3߸"��D��J;Q`�mR�^�?��hOL�b?E�� �=8��
��SZ��Ր�l=D�`;�-�oO���T�SG`j�۠��"���N�Hp4ea�=?�b?��O� �QP���',���#���n�&tÔO2U�����2c`����ՊG�U��#�O�T�� ��4"R����3SD�|r@�.}�a1�ĭb�~R+�8�X9I���AeZt(���JeRC
�pz�)D�Ň[<�1p�'��zO�-&�B�Q�L",���,���.��)���{��a-�a�qB��쭡ҡ�
N|�������г��"�Ĵ�v���"@j���|18�&�7@�)2KFZ_@��g�!�'?<I�!u���Bhe�;����y"��%��h0%Ɣ&��`� ύzV`���	�[jHA��(���O?Ͱ��$�>�0j��_0E\�p��y�~b垇e��x $��>@D#��_��t�	F.���p�31xP��N�w��|(r�F0Y讵(�k�hrr�Ҷ� ʓmy
t8""�2_綉H���kxj��FgA!"h�SgY�MN <��!bR"(��C�I#S:�XR��ċ#��񌗗/*0"�Τ�F�����vm��@ U6�pj��$�s�}�0�	�
;`+ּ.<�m���?D��ԭ]�d}���
J)>�t�	��Z�I�̥0G��(�������נ���f{����*��>v� ��m4 �P��SiՃPZ��DE�>�B؀eU�u�H����a�"�'�C�'[�w�L����1���<s6�Q�?LO�P[�BƗAb$$HpeԘh%��Z�n����&�-��\`Р�,�%�f��kj\�(C�
�Mٌ��t�	>�d����'D�����7p�I��-��fGR&�)I2��G�5{�vPzV�0a`����ᒚ��O��ΝO:Г�
L)52��ˡiM�4!�$,D�� N|9�݀�HV(��Ԝ
��P��c^M؞�p��X�th�Ë�U�Ҥ�ť!|O!hUl̈YT�`ڴi����֏Q�Lbؙ3�k�9fĐ�� �䀚��&^F���Ϸ^�B,�?��+�	G,�)�;�'S����D�_�M��E.,���ȓgV���o��a�1"�!A�pv�E R(���N>E��'����)B�B0M�|u�'^�}91�:T�:%����,@z
���'�ԩ�i�d�(�(N�;jb�ɡB�{>�p#5D��y�]D���nкV����.1D��c�!�.�B7B�,Y��	��,D�t��C�J'0R'�΂O^t�8� +D�pp�d�:�FL=9'�s��*D��g�Q�>�iɗ�̍65���`&D��XR��m�LQ� 4F�tɡ-$D�h:��C��.d��b�P�Ȣ��%D�p����fȲ=��%�A�88�@H.D�c0n;Ps>pi�e��wj���R ,D�܋p�ї7� ]D��${F�-D����/Ƨƨ=���3o�<�ӡ,D�����z�F���n�X��H�&� D�����cǬ}(!��8N(q$!D��*b�/�rI��d��(��� D���%�ͨ(�����A+��㧤0D�,P�/�Qy� �7[I_�$���=D��z��W.'��d����!b)��4D�d��*�����`�f�8��d2�1D�����y\��f_��P���+D��)WL�9�\�@���,���(D�4��]�6�`@��MU8@��� �)D�T�0�M\��$:GF!�N+D��s�"�\��Y��������)D��x�bB�
�Ҕ)�吳����&:�I0���Q�[	 !8��`όeSc��a�� l�T��f�I�,�\Q�(=D�,QC挈IC4d�8m:	��=D�p34��:"�,59qɉ } Mq�,:D���"�JYc�I0bZ���8D��R�$X�?��œ�+φ�y� *D��S�n�g��]�W@E"fN�k�b5D��sUg���*ac�6�.,�D9D� ��["g|p�va�'65��!)��&�O0��;�$��%��@�J;3L�}��q���w�<��'��)t����}��3� �	Cs ]�D3�SA�=C���2�9O�!B$C���|�;dh�<E�d/�
*x��a�E0VPC`�B�G������ٟF�uXS����E�<���a'�mf�D�M6q^�Ã.�w��l1��g�T>�	�kƒJ�䅠� A��Ҡ@
 ��'��ڰ`*�s��s�H��c ��j��9�&�V�!�|Y@4"O��k1g<(^�b�M��-��t��"Oj)��ˁf�d���>^"��w"O�QS�&C�ڄa&���7����"OTٳQAS#>�`�MҾ|H��"OF5�TC�L;XJ0,�Y�B���"OLj���12i��(A1��`�"OP�: �}�4�0�ـ��3"O�tH��-5�EZ�&�)k����"ONeH��ý�Bẖb�RN
@�G"O��xՆD�G�p�i��Id���"Olt�$B����!+a���t"OB�4I�jYbU2&���V"Ov��3�;5R�A
�KȮe�LW"OX�R@��^֌��e
$q���"O�Z��#��Xȵ���c���"O"l�@�_��Nu��"�/��\��"OP��"���C2�c��q�A"O�=a\W ��N�<?d��`"Oz�R͈֮3e�Q�3ΐ
2ZPPd"O*XZG�W�'��1��F(FUd�JW"OR�ە!֙}�FUQ0���$Kր*�"O��B�m��A�ȸbdZ3nq
�"O��I��8��ZGJ	�c  {�"O6|�&ǅ�K� �=\��E"Ot�g�
h�`�r�C)S����"O����	�g��{�K�@�8��"O�Mֶ$� �n\�Di~6���b6!�D�NC�(Q�o�T}�m��(�5!��ϛ&Ҕ�!	��^�C�Ǐ��!�� �׺�k�UyTx��؄w�!�d�>=�eB���<r�Y�vL�7!�D�y�<����RZ�lq7I\M�!�$�765���·F�R���(A��!�TY�aR6|��Q��nɷ�!�dE6v'hԂ��E�ZT��F�o�!�$
�,��кd��kXɲ]�!��/FqR4��](o����RM
�!��R	<�2#�Z�(tn�a#��6`�!�dI6CA�zQ�T�XY���t-��'�!�䏘�h=c��H�u(�	��fOH�!򤎸����a��,m\DK&���!��>��ᙣh�1-�Ңō�w�!��X�(�2u�!nH�$�YE[�!��3H�haz�#��n����w�ã6�!��.Fր���%'7x4Bc���]�!�ކ+�(M:'
�}ÈԫH�Q~!�L*�����VX���Cο{r!�'y3�-*׫ƵM�(�1��d!��PiW�Ms4��6;6�qr'̾\!��4�ݡb�
�].Td��
6U!�$��s�-�5Aȕ]|R���c�kE!�Dȩq��T�P@�)}and ��"/U!�L�^�>qh���q��4�6�[�!���(E�2�S"lG+2�h���ķJ�!��G#d|$�:��${ �!����,�!�P2G��,��i_*Q��ш�A?!�ݪs��cچkV��3�̏�a!�z�XqfR�	�X��끊m�!�$I�2���E�@+N�5P�*J";�!�� b��@��m�$��f��q�"O䈀b�Y,1OTt��!)�t	�p"O0��d!���E�|4�+�"O�,K�1.2�L�`e�xcB�5"O ��@�O->��������RD0�� "O�����[%N��2$D�'�x��"O|Iru�P�'M49y��И:�N!J�"O� (�"^,�1%"î[�j�ô"O�ь�9%��x�� �h?@D��"O0܈�'�ʾq�3��3X��R"O�}�ģ�2t�d 3CęX�:0�2"OJ8:e�P�	2ף�%в���"O����
�:D���Y��q�&"O��h��<6�\�1��i��E�d"O��k7k/�i��N�,y�쭚U"O,P��␲U��Y�U�Q�)�ԁ�"O�=����v $�s�[&@�h�r"O�@�O�8XD<�Fi�7t����U"O�y�fdJ`�  �(ܘ�~�ѧ"O<��2	ޙD]s��Ϸ�bY�"OF̛��(Nb�R%.I�TEKs"O>i���8��A%	�\l:��"OL	�voU4m|2����k]"�"u"O\��v�G�b��)���:TL��"Ob��U�\�,~�jb"Z"k(|�)�"O~,rR�A�YHTu`�`J3~C���"O"	�a^99_��x�Aɭ���9#"Or��	�� C؅X��Ŧ��`v"O���GӁ
u��0���
,�p�RQ"O�y���.(���J'dї ���"OZ$�VXW�R�9d$A��hpB"O�K�.|� -����R] b"O�iE�ă0ۢt���� dR���"OL��ԬQ$(���cRb�=N�<``"O^�Z5G�fX�[��	"���"O��q�
7��];d ڴSX@ a"O^�A1����4��Մ�9� )r"O�,�!�&xA��a�m�����"O ���X+G�X̃s��&'%�Y��"O"�3��l ��QG�43�e�C"O6Y(��=�B`�!�C�\H�Ц"O����H�[��]�l�=�h�J�"O="
�2_����[ǘ���"O��8����c<��d�<w�ޤS�"O���"cۻl����ەn����"O�Lq+� ?8� x�� ����$"O������j����̼@$"O�5��`�*6:QB^�t�1��"O��pu�E;x��0�S��:����"O,iDA04^� �#��(� �"O&�#��W�_��0�Q�ߘ
��X�"O�4��g8N%���!�($�!4"OR��m�5����� K�8�0Y#�"O<�	FM�2&2�S��Z�2n�"O��Cj����W|Ö��1NN��y������yQ��m�Da� 익�yb��"�1����!S�<�yR��!���∘�`����A��yr��(cW匫,�D�S�*�.�yRN֜<�h4��g�:&2���u�C��y䂦6��T;F�ӠI�L[����y�m��Sq@y�l�+sz�g�̀�yR�Z�7��Փq�5x~���֎	�yR A�r��"��ڍG��$� 8�y
� �л��G�~b��������l�g"O&�!e�I����/1��F4D���O�&L\�͑2hg��0S�2D���S�,?Xh:�)ٜ3��*�@0D����@5~<P i3)\HZ�8Ì,D�4Qu��N!����# -c��.D�����պV���l����@�)D��+��4iA0�Z��&C̬�`�+D��`�$,�\�a ��{�  e)D�hh�XBT�DE_�hA��rto1D�da!_�"б�2& :j�e�֢3D�|�3�Ӻ%��.�;j3���b1D�|���M�2���IP�#�-� �0D�����]��p(a�\6?e>� T�,D����Ʌ�j��׀#-g�|�w�5D�D��I�1�n�B��!��4D��rG%ǪRP8j�mޱ]bNpÐ 1D��Y�3��!3���"z�k�!9D����51�I��&Z�T0D�<D��:W�R�j���������#6D���$�B<�oF~+�Y��o3D��s D�l��,ѱ3嬕j�
-D��H@�
�n��3#��Q+�m>D�8�U#��5ξ�x�B��k�#7D�����E.�dK"dĩc��:�4D�|�3��Kk�5@�Ă!&Zʤ�3D�0����0b�#˅�	ܒ�K6�/D�d��!F5�Ue��!dq{�;D�8Q�IML�i� �e32B=D�T[�@�<ls��������5D������"/TSqh��^<���Ub6D�XPT˜�dZܺ�9u:P����5D�<���0N8�@��#�<�h%8D�4����u.���T��x�C5D���' S���8C���4��q��*8D�� �/S�T�r��W5��(�!+D���~<��I�ː�r&�`�4D����gVc
xc&Y�����-?D� �wiV�d<��FE��v����D=D� ���Z 7v���f�"�!x <D�Ⱥf�rj4��԰$�Y�5D�������^�"Ep�+���p5D�0����Kʄ�X�%&3�Б��b4D�c�	�{��m���Ok���Al-D�L�k�>:��LZ���3Ȭ��-'D�h�dդ%TLsE�نw � *�"$D�X�ы9���+l�)5�z�.!D�$��)��~̾P�b"/�}��F)D�̚a�R�(*`�`�V���e:�$D�\ ��*�C�!�]��X@�#D�����	)�x�rc��z���>D��pb%f�f�b!iщ4�Z��� D��zd-9hTp�1"0!9$+3D�d�̈7s\��D:��!O/D�Sr��
i��H�5@�5M���T�?D��9R���jt���M�Q��)xW(3D�HA�@�:dpę
���M�ص��K0D��f%�$2֠�kQEK�n����,<D����/���B
<1G����B8D�l� �Z2���w��8@)s��6D��&)�,@bLaX���,�PF!D�P�D��� pf���'[&C�I����q�dS�j�A��ϛ�9!C�ɧ=E��D��'�(s��XvDB�)� ,$yë�\�1cb�ъQ�&�9s"O�!օ�6"�8+���L\�+�"O�{d�� w�>-*��1?1�ԛ�"O���%��<�f��ǅ$xy�E"O��+4O5=l�IÖ� N��C"O����9/��y����I�`Б"O�E��!eS��
�$�!�Ѹ*O(���{�*�8QkY)c�0���'�t]�h�y��40Q���[��)#�'°8#�ٖ#�������q�'���I���$��"b�Ž��P�'�Z��&� �x���QCL�5�f)b�'���FP=\�dy@�86�|m��'"����=z��ҷMQ0y��
�'�T�,YM[(uS���.搹�'-�10��
p2�!6�L#+�И�'%� �7��nݞt-�.�� �'
�L�Ib3���P� ��	z�'B0Q��$=\��'�X�=��"�'��<��WEDL�q���sPL��'���J  ����?���?�H~��tݠ���f�;<�\�"�P&h}�}`]��"شL��/��i BT�)�BL�B�d]9��B5d�>����̟'��	�jSdR�'E��%��'3���ui�]�Z(�H�NV�3�'�R�'����Z��ݴ<\��n��c�#ѐ�s-#M̡Q�@4���O}"�'��	�ҎD@��5�xhJ�ƌJ\�(�u�צ�ϓ�?CIMM)������D�*�.�[�|�m1Y�t�3H�1):��O��d�O����O���4��]�"����;!��XB@�M�2�|��I؟���4�M�#���|�I���|�'�!���̚!���&��'e^�-�$�md~�',��dh�)�`�Ѵ�ئV�P�)�៌rq�|�Y����ҟD�I럌�eIT�������9u0։��� ��oy�l~ӎ0q7��Ot���O˧#�:`'",�ՁF*	�,���'�.��?9�ʟ��Yc�ɬ�@��'
�g9.4��
J�.&�U#�靻}q���|�v-�O��	M>vF�3�$���I@7��y`��F��?a���?����?�'�?�����զ���Q�*��( ��гl�Dq��'��U�I���柬�'B\����2�Ԑ���J׬��pi\�u}`<������E� ����?�!)׫��Ya�AҸ�򄑙O��̠V���'"��T�
5�<)���?���?����?�)��ȃ�t[�ق��S6?�����n�ǦQ�ga���h�	՟($?m��-�Mϻ@u�e�5#R�8ݦ���� %�b�
w�i�b6-�w�i>��S�?9r��Ʀ�͓^��,���Q�L�ܝ�"N2C��,~(� �,�O�${I>,O�I�OD!!��<s�U*`Y�Ǿu��O���O����<)t�i(��G^���Ii-av��"+z����b� *�Zp�?Q�U�8�	զ��O<!�㟂(����ҽX��%`4Ir~R���{A�<��m���O]� ���e��A���bO��E��X1�òO��'���'����Ɵ���%_�f\�ۢ�ӵ�V��¢��,�ߴ0��x���?�2�i��O�nv�`���#��I�y����x���O�u�ġݴ���S�С��t��:���Q>]�DHS�]����(�$�<)���?!���?���?����f�(��d,�� f̣a���'+�7MQ�b���O��d,�ӎX�Yp�FB�Y0h9&��a��LӭOB�D�O�	'�b>�pх�&)v�쩇��s�%K�oQ�o��8���0?Q���"3�����!�䓲���Lx0te�4/@4�f�*j�$�Op���O��4�Hʓ5��G��d�6n��Qy��V����[<!�%��D�y}�Ik�d�l��M�Cg_�9+�]����TA�-s	�L���3�4��d�%1�����'��OpGC��K�0�0th̯e�U��U��y��'���'��'���IR9I2�ɡ��.'���:YF"���O�d�����dy҆dӈ�O�B��>�����(�P��ԩ�a�	�� �i>iBD�Ǧ��'~�q"̈́�"
�1�&�I�)r�eH�X�H�ɐh��'��i>���럌�Ʉ|Lx���0j��`��h��͟8�'H6M�5:?d�D�O����|��A�7���@�w���2i�E~�O�>���������l|�����Z\T���ѭ'(mpǧ�
;�"���H�<ͧ})���֣��tϰū��	�HȧeZ�B��	b��?9���?1�S�'������/�-"?�y
��Z����\��	џ<0ٴ��'�Z�;���
]�>�*,���A.q~v�ڐ�̊3��7-�Ŧ��e��ɦ!�'�.@�F���?����PC�m��Y� ��Q��`ܖ��b6Oʓ�?Y��?1��?�����t=ڄ���X1�d���H�9���lZ+Hr ��͟<�	G�͟������F��������m��0�y���B��?����D�O�f>O�����\+�`)(b���|/
��5Oȵ�`�?���)�D�<i���?@�ΑfF���4/�w89c���?����?������ݦe��Í̟���ӟ4��#�7w1��{G�M�L�����Q����ן��I��ēNx�p`N��*�0Ma�a��|�%�'VH!�r�_��!Ҋ��̟4҂�'��,�W4F����d̔.bY��r�'��'�2�'��>��I *��Z��P�f�j,rW�Ä[�2(�I��MK���$�צ��?�;89ƹj�d �4q�� �\��ϓ�?q�����=U+�֗�PX ƍ/w�d�5� �\cd�foH�ó���b�<�B7�/��<ͧ�?���?����?��-�`'���L�D�hYB2!�6��Dۦ���ҟ�����$?��əBz���ɝ!N��Erf+N..�D=r�OL�$�Oby%�b>��`l��?
�}9��>k���bJ�&&���'?���pO�D����dLq�� � �an\�f߻I�����O~�$�O��4��ʓ*���úDg" �/O��]z��3'�p�h��<kb~Ӳ�xگOl��<� ��(����`�Y2�� �
�;2`�i�4���P+g�2�I��9y��� �.�(��K�Ď�@���T�!����O|���O��D�O<��&�S(d�x������(h��S�I�Vz��I��(��+�M�bd���ą֦�&��Hg��8��X JׂZДɲ�A�ē�?���|J���MK�Ol��ߴ����((]t�+hV)�$�{�'f�&������'C��'�l��lё,�p�`u+��O+V�˦�'�2X����4�١��?����iN��L�f+� `�֌O��Ɏ����O��$MD�i>���4��� L�D�yۖ�H�u^�1@�ds|�J��#?���5�������-^��K�C,�EoC���9���?���?��S�'��KǦ}Y ���q�V�9po)i
 ��e�ܥ:���'@�7�-�	*����OR���� w�F�AR�D�~�k%+�O~	l�)t�x�n�r~�K �h��<��|���{1.�2JK.ӬīdE���<����?1���?���?I+��t�$B�M_�m"�I� +���DjE˦�js�K��`��ܟ�%?�ɥ�Mϻ5ܘ�1 ���"��W
S,��9Z���?Y@�x����6`���5O&l!�D�6���(_(G͔Y�8OF��cC�*�?	�l9�Ľ<�'�?�G�	�̢ hUqk�M��ㆰ�?a���?��������2R%���������3eZ�E
�c�M�&\��D��o�C��I��M��io�O��Po�@Z+����R`�5���*�C�.�4-�r8�/��⟬�pM�	���V�K�,��{pf�ʟ��ϟ0����D���'����bÒ9��R��ܣ<�xPF�'kV6-�j�˓}���4�z}z󅊬
��3�/9s|� )F<O(���OҘo1`yoc~�Ɯ->m� ���/-Htq��#Z�Fd:G��I��QŒ|bS��ןX��ݟ`�I۟��#&��{F�ȡ��2[���e��Zy&a�hkħ�O����OT���p��RNh�D2�͓X��'��'�O�I�O��)��Rv���#�K���c[�#ݐ@��9;��	�b�y1v�'s�&�p�'�@�C��/T���c�V�zP�'+r�'�����W���4@�9H��f!���T*���Ӧ��g<p̓o䛦���{}�'"�}ӂ8H@�Db�`�쁊-�0{fFʦHŀ6-g�p�	f��Ta��O�����P`�`F*�/�Tl6�ٖ--�y͓�?���?���?���Oq��B`�16nD�W��)�H�x"�'��'Q�6��-N��o<���|¦X	}�`Ȳ�Z�A�^Y���D/ld�O6��O��]�6*?yS���+W�2�AV̖0B��r�>R%�O$iM>*O�I�OB�$�OR,ZebƼn��i�2%ƬQ*Ha9Ҍ�O��ķ<A��i\�;��'���'�哌��	��*M?9r��#@73UH�
y�Iן���"���|B�9���[���]�a0U���8�v@B�@�!��e�f!�r~��OUL��	�e��'x�p#Pʎ������4}b���'���'[b�O�	�M����U�~��2���b�x�D�B�blB-Oإm�w�b�Iٟ0��-P&[_ʀ��T�y��F��D�ݴ
ˮ�
�4��D�e�I������kM�ճ�IU	j5[`��'Tl�}y��'yr�'���'�RV>ysaI���xrr�է3�\��F�$�MSGEH��?���?�N~����w��@�gLG�R�Ԕ��h!V�a���'�o-��I��
��6�h�8ص`C�Yh>�+^3U�u�bq���%�����G��dy�ON�D��Q��`��g׀ �F�B�)NR�'-�'t�I&�M�B�	��?���?�3
�,v��l�94ZL��m ��'4�˓�?I�45�'���2t']�>��"��ɯzh���O1�F�'o�T�'�)��?�'�OP�m�`K
�;���fϜ�2 ��O��D�O��$�O6�}r����tLH8X���c-�V�4Xy��o���G)v��	��Mˎ�w6��5o͝z�Hr7IY"=c�M{�'3��'��7m4wH�6M,?��,��;ˬ��H�$4h"��</,�`��L�|#�AJ>q+O��O����O��$�OfU��������ㄒ
��%D�<9Դi�L�ɤ�'�b�'��O�B[ˆ\�%/�5�04P��@*P,���?������O�R�(�Xh�l�qh�pf@�T�O�a�O�� ��(�?�0�>���<a���/�j`�2��`���
��?���?9���?�'��d����V��㟴A��	+VJ�rF�5s��d�a�۟@��4��'x��{盖�f��$o�=�� *�A͎d֝��ѡYN�,�%�B����'�fQx3��?M�}���E�e�gC�Rb��s����?a��?9���?�����OhEy�B�(Y��O83��a ��'+r�'Þ6�F�:e�I�O�np�I��%�@̓�-�Z�qhsʸ��I>y���M�'T	�4��DD�+�� ���!Z"Ҡ2cfn�@�B�?�%-�D�<ͧ�?A���?�ŇR��4,�&�E}��)��'�?����$QQ��ǟ|�I���O�x=r�.�$ݬ�`�J�:�@C�Ojt�'�B��?1I�)��l��䲧ㆂe�����T��2��5��{?�	���dN��� ��|�L�8�IRE��oAf�Sb!��'��'��$U����4jD�Iȥ��j�L<��ƀ�� u! Kք�?���ig���d[}B�'���ZF^N�|�����ȰIC3V�4F�UĦ��'`�=�t���?i�X���c�-���U�fI��Sb`�ܖ'���'lr�'B�'*�-�Ah��ؠ#p8�D������4rH��?����䧰?�T��yg�K�rvW��(apA�O��X�����I<�|�C���M�'��=�@iL�g�i�WL���
�'��Ly�P���0�|�_���,��;�n�v�,��%�������	��	xy2Kg�X��D��O��$�OB̋�Cۿ�������i�B�cf�$�I��D�O�� yg��JI�rAJ5*v�,҇�5?��%�G9ɠ����@;����?�����>���0k��N ��`��M��?!���?1�����ݟ���V�%ҨA	F4{��Q��ɟ���4	��Ũ��?!��i��O󎖡�ڽ�e[!$.6u𧗲O���O��Y&�iٴ��DS�n!��'�@�,.�tqI�9��ш���Li�'��	ڟ����(�I�\�I�K�����ܳy�"�yS�_�bՖ'��7�\�v���O��D9���OH\�@�ήɨ�h���5��UP��W}BOg�,�n?��Şi�"5)�� +9jiʗ!¡i�.m3R��H���'�h5�v��3�|"U��ڤD��v(�{�lY��8���B�'���'��O�	�MkP.��?����Z~\��e�4���G��<��i��Obh�'��W��x�N�>@j�`a��zɮ|K񈍡Yy@9n�T~�-E.6-���ӛ@{�O%�揻�,���O�~��ث�M��y�'�R�'���'�"��s\Fh!D���!ش���N����O��Ҧ���YyR�g�,�O�0�LQ\��(Ӓk���a�#��c��⟬�i>�����Ħ��'v�zVϸ!��ʮSî�U�TR%T��I#yq�'!�i>U�	����	���1pe�<M������/�6��I˟��'P�6-�>�\���OV�Ģ|z&`�	\����a���0��aҴLW~B��>ѐ�iO 6Vo�)
�����`����"a��Ć8r�zQX�;:��d��G�埐�&�|BE]w��`�(�-6��c���pz��'���'����Z�`��4C�X㜫Pr%(bB�F�`S�#�5��$�ʦ��?IR��l����A��*������O�K\��rش �f@�YU����� ��+��T�~c�D�O3\ "��t����<�,Od�$�O����O����O�ʧsAdX � w?��c�d���,Y�i|�� ��'�"�'��O��}��.	�^�L�٣�P	g�RA�o�'B�Ym���M{t�x��t��{v��3O&���)v��yBG@г:����=O(!�C�_��?�).�Ŀ<ͧ�?����&���I�l�9���`G�3�?����?y�����u+�ӟ(�I�@kbBO����)5��%%��Z�[u�-��I�x���ēs���*��.^TLBF
Y�OB8T�'���)�/�d0���h��p0f�' ����[+@����4�V�z�L����'O��'�"�'q�>��I$la�A��OR3a4 ���H�3h�h���M�*K���$���q�?�;�����͉`s�8S�Y�@��?	�1����-+_�V����w�٩G	�d��qJ^�ʒm��@0i���4V��&�x���$�'�'wr�'Mjy�'�]�9v|}yW�Q=KK�d��V��pܴJHXB���?�����O4r=�" ��t��mb�h�.-�9��M�>��i+�7]v�)�S �rSF�	�ڭJ��� *�`��O�1o��Rb����O��9I>�(O�-�Q� ��8�J\�U=l���E�O����O����O�ɬ<�i�N���'ǎ���/
�	0U@�=�p��'R.6�!��.���ڦ��ݴgś�DE�{���k��Q�"��0Zp�@�J`�i���5h��QI��O(q���N���^U�D��8���a֥ާ{����Ox���O��$�O<��%�Sn����-)��a���.����	������M�II����K֦Q%�(�Ý7a| �wK��!C*�pT�����B��qӲ�i�0U�6-f�,�ɣy�ܝ;�a܂i�ڑY�IV9R����(�>r�]Y�y�O�b�'������ `��O��R�n�u[B�'��ɨ�M{�C��?����?9/���r��Z�����3 @,�����x�O@��1�)2�O�[t$��?Wh�Îʇ#����17�6��)O�	���?���/��:lؙ7 �	�0h�Pl^�P����O����O���I�<	��i5n<a!���{�XPQ�P>V>�X� ^,��ɂ�Ms�2�>I!�i�F-+c�n�y�a=V�d�@-tӼm�)s�n�_~���(n�e���i�=E�@�V8u�dͰDj]���D�<���?a���?Y��?�.���Y�iU"7ά�"͟%��p���Ѧ�a�Yy��'��ԉlz��p��7.1
`���8�s�ʾ�M��i�O�����霘��7�p�� �@�����@���	ѹ�� �3O Q�ժ�9�?9P�)�$�<�'�?�`��m�d
��M#��IբR
�?y���?�����dTɦ�J�Q̟��Iԟ$�eaF�mWz8K��	9?�@`�jOp�|G�I��Ms��i|�O���b�ƶ�2�â�݅1������p�7L�hY"��O.擗i^�Oҟ�ӦG�X=��.:����¡< ����O���ON��4ڧ�?i-�:$�	�B54��܉�D�"�?�A�iZ8����'pRJ{�p��]1}����ό�pM�p�ej��-
D�I�Ms1�iTl7��"iՌ6�7?�b�ǚ%X��Z`�F<K'ɇ�2�<-Qj?=��N>A)O���Op���ON���O�zwE8�D��F�^K�,���<q�iĂ��V�'�2�'���y�	�y�(�3�/�>cMZ�hϬh6�꓿?i��Dy���O�y8���M�Ya��Oc�f����g�HI�O�������?���#��<I���PcXP�$I.Z�̸Zg����?���?���?�'���򦭉�n]��t���M�()�@�3^���rw�o���4��')6��?�)OP����M;Y80�ǩA�:�	���"!��7:?����*��� ��'��{��<a����w�$|}��´a��<��?!���?���?I���-E>�l �hA6�m ��9���'���~ӺDR4��<1��izɧ�6���Z��i5�K+mM�)�ġ���?!��|JG���Ms�OEB�:tt��PkN\�ȡĬY�G2�?�PK.�d�<�'�?Q���?�fF�kјkd��#��0��M��?Q����d^��-h�gKzy��'��qI١(ԗm�:�B�E�%\���[��Il����S�t-��]A��w��?{�����d�y�5��)\��a�O� �?��J/����qR4أ�"L�tv�i ��" ���O��$�O���)�<�#�iO\4���<J:�)Fa�4jmpM(;��=�M���a�>���p�pih3�F�\d�تpT=,0����2Q��'�,@��f����B&U+3`�T�~���L��daE��>u�;�ƈ�<�,O��D�O����O����O��'l(�z�m\�V���[����l-���i�d9b��'-��'��O,��t���F�������D�v���g��u���d�OX�%�b>���̈́উ�7wuz�ɞ�C������2��D��LI��)�O� #K>�,O��O����(̅Ex<3���$~��b+�O��$�O���<�p�i�`�Ҵ�'Y��'�Y`F�R�?���z�NY�I(ؙF��y}B�'x�OD|�eCА!��|��ɿ$W�Ie����$\�*����r��Z�S�+�"��ȟH��mV�$S��뗥��f�xa`��������	ş G��'Y�����J{�&ڰ{�}8&�'oL6�3T�ʓX �V�4�4�а�3<��JvA�z �`0�0O�$�O �mZ�M� DlJ~2`L)r4�Ӈ}�����)� t!�ə��_,RL�8yЙ|�[�������I��|����H𤂏%ܠ�!C��y�ԕ���pyB�a��`z���O����Oړ�����"?62]+��C�Md�j�MN }���'�"�'zO1��I���ߒ�(���qp�̍x��������)�&��R�\y�[�C�V��3AF
�l��d�:!��'R��'G�O�� �M/����ɮG|�������	\�i=`���M�����<���M�ոi�Mɖn��?x�7��1
��ca��cd�&<O>�$IX,2ȳ�����?9��OYNu�r�Jsm�E�W+P�?b�	ǟ��	П�Iӟt�	O�����G"��eva#+T(� ]����?9�Q�����|���}���|��ۈN�~a���G�;��1��qp�Or�d�O�I=D�6�4?��-O�?G��
7ν Z Q�+
�-�yCS��O��H>Y+O�i�O��D�O���o�	�.hr�b�-5����B�OD��<qp�iB�l��'F��'F��w�Ф��	�X�B��vb��T��	��\�I8��S�$,��6Qj����T��37X�
�2@`a��x� ��O�I��|��!��X��ɂW�՝@*���͕�5�������sr�]:�*�G�4i��ʤ  @�gf٢=�z�tϞ��D�kB��G~�{P,
�{���9H?����a*˞���2�O]��X��l�����a [�̢B2c�<8z��/j�R��w�/Q�Ψ��߈uEܹP�k�"7����i��7��=8�F�/��X����.E���p�ԞYlAm�8�B\3n�9*�UaW`��=�>�چ��&��4���㖿+�f�z��!"����W�Z_�926]����aI � ����ǒ%N�V��%S9$�$E�\���Ke��?�K>�,O��x��e��PQi9ve��Kv	F:1O����O<��<�ɐ1PW���4�.2�2���F	>�	П��I�IP~B�S}�Ҷ�Hyz�oÄo�ʄ�@���d�O@�d�O��#ji�ǝ��� �F6�� �bG|�Y�h�6��7��OV�O�˓jP}�>�����%c&��W��������i�I����'C�e�P�<��O6����\�R)Y#}8*�D��W�0%&�P�'bR  ��T?MS�BT�X���W �J��CW.|�Xʓz�xT���i���'�?i�'��	�S,,-:��"s�x��f^P��7��<��h���OMZySf	�,�:��
q5� Bߴv��{��i���'�2�O�b�S�e^�gX�X���%E�.����M{V��F���\��ƳG(J%�O&�}��%\��qo�ş�����āvoZ����?����?��� ��a�����1L��W�dx%�Q56�1OD���Oj��	�����&�#	r5�Ѹ{VB�lZҟ���A�ē�?)��������J��)��L�d�D�E��K}��Ø'���'V��aR	��8r����h��̐�%����BH<����?�L>�)O�m�"��4�(c��~���CE
M�1O����O����<��IX){�	*��Lh-�?�����mX�H�'��|�R�x��E�>�W��0_bX�a�;b�P1S̄P}2�'��''�I6[�",iO|�ć�/Tj(URn§������L	A���'J�'��x���l���8�c�;`�H�p5����M;��?y/O*4�A�v�Sϟ���lʨ���
H� ��ap*G�A���sM<��)�tC,Y0Li ,��<�l�,�I. H���ן8�'��$�'_Zc&�#��Ƀ8��A�
:7Zڌ��4�?q(O.D*%�)��7k`Zј�Kc��j0%P1M���LW���'��'��4Q�0�O���p�
��M ��:]�کA$(�>Y���^���O� ʘۼ�h�Q5#À1˗�Z�P��6�O(�$�O�0���O2��|���~�<M������XU6��"h��#<����t�'��'�4�T&��$R� @7�Q��t�{��>��	H����<�����2q2tBR
 �\32��6gx{s�x�����O���O��p4zY��F6QRx9E{F�:A`��AM��xyb�'��'�r�'��쳗'�3�~��dV'@az`"��tpb���y�'���'w�I2V�ɨ�Oh��A� L�PMR5�⑭#���4���O*�OP���O����������JX�afҬMܦy+F�>����?I���D\K"A�Od���#����!�^c��í!��7��O"�O����M���m�_��� ���ln�QA�/�(H�@Do��$�	~y��C$z�'�?A��b�c��z�̍��*�x+4��[�VD`N<���?)� ���'�I�;6 ��;�Dͬf�X����ڍ	���V�T���Ջ�M���?1���:�X��X�+���"���u��{$F��{�T6��O<��Q����`�}�A%ϫI�"��l�+�t5!� ��QNݳ�Ms��?A���:@[��'H^��KF,n�+�Ůz}�x�e�{�n���d%��l�'�?y%˼:T���-9!��0�eI�Yśv�'2�'n���Ǹ>(O����l�R�_�Lv����S�$����6�IN	"�'���Iʟ��	2l�8 ��X�ty#��6Lx�ݩܴ�?���.��\y�'5ɧ5#��'C��ض�G�S����P>��d�7M^�O����O$��<Q���Xk�r��!{?8�`�ώ>e��ȃV�̗'���|��'���G'9��Ab��F����i�1��0r�|��'%"�'%��Ĵ��OQ�˛'Y�0�����8"��x�ܴ���O��O>�$�Oz������R�NK�U�w�[<5���@�>9���?q����䗕1�~q�O!B�N�0X����D:���Ȧ�V��6��Oʓ�?���?��d
�?)��Tq}B��O�F@�� w��^��M���?�,O���Ig�t�'�R�OZ>����:K�FUA'j���|E1�$�d�O��DT�G78⟼���
�᧪�ZW͛��F�O �oayR/^
>�d7�����'��4&6?!$�!!���f�݁]�^hzA���і'�db�'���ؓ��V�B���bR�r���$��.�MCcH[�GP���'$��'X�tf*�4�0�����@����/1�e�`ɦ}��,П���~yҞ��'�r�A�E^`h�e�?�j%Zqb��6��O����O.�"b@�i>]�	x?�|zn@st��fe���������My�ML�b���<)��?y��\L�����>L�6�S"��&��!C�i��jU�y�BO�	�OB�O�NN�u��0qΆ�}��,���$f��	�_�0]��U�	����'�2bJ7b�!�F�����p�5���1V�h�Iҟ\�?A��?��ߐQI �P�(SiD��䥊%g�F��b�Mw~��'���'���;..�ȟOZ�u �aeN�QE�w)�t}b�' �|rW�83Ġ�ܟ� 
�k�X\i!��b�l1/�����O��D�O�˓/0� e��D�Ti�җ.* q����:Ȫ6�O��d�<I���?qҢQ�?�L?�1$�U�IF�;]O�M��CkӤ�$�<q�{��,�����O����| ��>&0������xr�'�ίJ��eX�y��(�R��j���E�
(  ���i��2SB�4����������'w8��Ң�2�7 ���6�<����?����Ԑ�ܴt����@��e�b����5X��m�^9jD�IߟP��ӟP�tyʟ���G���p�V�a�J$I�A������K�	5Ks>b�"~����/i� �� !pv�%0'�P�7��O��D�O���&�<�O/�M	�L��8J�JqGS,U����'��ڄ:�$>I�I��	 $Ɛ�㭌^���SG���Yڴ�?Q�+�W~�����'�ɧugfŭ`�&����I���DH��� x��$!���OH��?�ӉH6f�(�q�ףjx��W-K�C��`k.O����O�㟸���08� \�+TOD�A�Qpiݎx�T�r�(_'=
�y�'�B�'/"X������4��[�46_ v�L��Bջ����O��:���<Y����?s�P&r�&�!��A�]��F9�����p�	�̕'tRPA5E:��6WO2�:�c�|D���Y)y;�DlZ֟ &�D�'- Y�'��CL�xY͜�\�\ ����lN>l�ޟ��'�r%�&J�͟<���?�FL� �&@5ʑ/�;7O*��OJh�4l�;1O��5N�Rl �"E�`�6%L ?�7�<I�0Eb�6�'���'9�$'�>��0�����T,hF�2�,\
B�8nZ�����0#�V�I՟̗'�q�4	 E�?���2w�H?Jŷi�ĔHqj�Z���OD�������'�	/(ef�8dF-I�y4b��m�d��޴�f���?Y-Ol�?i���#�਱�h�}��	�fE%WiJ��4�?����?���
�B���NyB�'���	�"u4���R6Tj��Y6&���v�' �	�m���)���?��"unm�pI{�A��R:�����i"������d�O�˓�?��6�,E� ��9V���M�'S�TQ�'�hʚ'����X��͟@�'�F���[���ȁ�fM�v��9@��P��등��O��?����?�Q%<N���ʈ/we�� �.S��̓�?y�#�\�{��?�(O�K���|P�718���> Z�ؗgYԦq�'��S�t�Iǟ\�	�%f�i��G���(����
[�8к���>9�"�2�?!����K�RM�OpR���k�\�h�*�Uk�p�$
�*EA6-�Ot˓�?��?)���<-���K�<:9"�$�2t �(@M�&�M���?�+O��1�h�]�$�';�O��D!w »J�z�3F�J�V��9�K�>!���?��w��Y��������Ew�U��)m�Е���Ţ�Ms*O^�떾�6-�O����O����e}ZwC��y��ѥi�] C��=��4�?��X����?�+O�>Qɑ�ɅKHJMz�@V�K��L�2*xӠ��bi���	����	�?�)�O�˓pL�- ��.p4� �&lN[�4�лi^졂�'��Y���r�h�0p�F�ӆ,�>0I��%���պi��'h�ᇧXE\듬�D�O��Ɇ0��Y
D�K���Εt7M�OD�l���S���'���'��9Ѝ�~ ��p	�)Ao ��tӸ�ğ��,�'�����'�Zc�K�5U�|��m�����NayO�<,O���O��D�<	T��@�j�%���OHP��N��_�n�ʓY�\�'��V�X����|�I� HBu�L�ܑ9eL@
o@�P@t���Iٟ@���@�	Jy��݁B(�ӹ@eD�2���7pf潙�"](�(6��<9����O2���Oj��G7O҈p�(��>���g	�I)�q�C�Y��M�I�����<�'�����~:�I:P(G�5T"$s'�P�Ƭ�3�iD�W���	ߟ��h(��i��(F��(���H�ma��u��6�'�]����'��I�Od���8�uKA$l�2��e���3F���S!U^}��'U2�'>̡���'��I %}�c�D�y��#�JM^a��T���d�݄�Mc���?i��Z�Z�֝�h58�3��\�Km<52��d�Z7��O��D��PT��Ol���O�&�X��֨6E:}�#"ΕR����4Y����i���'���O��ꓫ��Ú[�H�Ks� '�Uc$�\	f0o�9-f�I|��I���?�pN���$1�E۴3"U��5f�'.��'���f,�>1)O
�������Ux�F��E�CXz��2��x��D�<�CM��<�O�R�':�	�(Ю���#
Z�M������'D�H���>)OJ��<���ի�]F��*�A=K�h�P@}�AP�y��'�B�'*�P>�I'&�t����g��wo�y��اEI���Ħ<)�����Oj���O�bSb�28����N�"�rl �B�	D��O����o���$�O��{�0MS�>���R���z��!e	!!��������O�ʓ�?����?��*O�<�RhőMM�0Ձ�1_������>*���'���'jR�Hz��<��)�O05i�#��k�<]�LV�-��)�b	OȦ��Icy2�'y�'����'���O��CO��?P`P��W�O���J��i,��'��	�L�E�������O��)=�NĀuC҂P�&<�`DL�cn@�'�"�'c�+�!�y��'�Ɉ1N4�i�{E0-Jł��.?���f�<ԛf_�Pi��M��M��?A���dQ���"P^�" ��T�0�� �j7-�O@�$3p}�Vm��'�q����Ǝӓ.!��8s#S�vgJ����iNT�r�Id�N���O$����Ƅ$�\��7v���a��ؗrB�����,\�dp�4�ܜ�������O���(�BER`��L`\۳!��bwd7m�O���O��B�Ql�I؟(��g?IF� j��=�'��	�����ҦE$��[��h��'�?1���?�  �%uQ�xIv@J�AZ=�P+[�@���'9�ԡ�'+�	֟�%���gT)1"���5�Pm�ƥA����/Y^$�����D�O���O�ʓ{�h�z�J1=iFyq 	ADl�� 4i�x�O��� �$�O��d7��e)���1A�u@���.hs7�d�Ol���O,�=B\��=���Dˏ�u���faء#q u3��x"�'V��������$��x� ��� �a�`* e �jc��=����O����O���L�����h�<Q�R��A�8̐U$K�;Q�6-�O�O���Ob�a4O�ҧ� �A���8i�� �a/�@ɢ�i/��'W�	3ns���M|z����K��X��V���'�d��n���'N��'�6Dz�'��'-�IR7@��IX3lĞ��:4��"��X��D�
�M�#X?��I�?A��O6��	�77�U�2��
���"�i���'���c�']�'Tq����t�B��	��虁X}����i�\-�pu����O������&�@�I�K�V8���V#qeb�j���0N�2l��4A���c�����O@�i��/#4j�.`n=;B� �,ho�ȟ�����)t ����?����~���o�l�z�f�-�5i�\��MJ>��K44ɉOQ��'PR��r"�W�q�N=��H�~��e0ǰi���R>'��b���	g�i�y�Ə�>{����J�1P�Dü>�p��<�)O����O ��<aË[Y�xx��܋cDڀ)p�˻�dAP��O��O�$�Oh�(��;'(��R2
��)�s.ҳz��<����?�M~�����<��IW<%N��
C�Z�y]^���\���	؟�F{2[��I'b��C1�(I��]�3	�7UZRŠ�O,���O���<�7�ܺ�O�P{�!�����q�L�"�&-85�lӰ�=�*O,�2}��£<�P�wʉ�� ��4d�<�Mc��?���?�Ŧ؅��ɲ<���Oy��[&�[VPbqJ�i���`��x��'��	�@�#<�;i��T W�b@��%��2'���l�^y"�[�	��7��O����O����r}Zc{���`�\��� ;'�!Vi� �K<���hO�'O`1blѕ#
�hG�-G��@Qܴ�)����?��?��'�?1���	�� �n�V�,cE,�{V솷Tݬ��'9��Ѝ����O���KX0YJ��0�j���b̘ڦ�IП��.;��H�O���?i�'D +4b�)N��9
s��u�,�j�OL˓k,���D�'z2�'�
�X�'RvZR�k aV/5������y���D�a���'Q����'PZc|���3l!�zt��C�`�#�O���"2Ol���O��$�O*��<ᔁ�= �I��(r��i?*���4R���'5Y����ݟ���,%$�0�R@�L(����G"�QD�c�L�'7B�'��O>xa��(q>�g/YU�b5R�^:P��DH�Fn��˓�?a,O����O@�$؀P���: "h�A���_�lY��7m�O ���O����<Q2�ƯxD����ؽJtĝ�%��8�Z$hue�m��6��O���?���?��G��<����?Y�aX)3��@�"�Pt���x�:��?�(O@x�3KL���'��OBfh��Ɉd���:�T�p����ͻ>���?��)�T���ɧ>)���� ��5�TAH��x����
�
_�7-�<i� ��1T�6�'�B�'����>��P)`�!�.�"J�2E����uoZ̟`�	$���#��9O4�>�c���pEJ	2�C�8 6��	Dt����Ο����ϟ�	�?(�Olʓ`�+
��Bp�{q�#���� Φ1��*g�|%�����;����$���|�h�
�"�;�$�;�i�"�'@roY�~�z�����O��	4<�#�dR�hG:�JQ��A�@7��O����8�S���'v��'���hՆC�Yi1eõh�y)�cp��d��4,Va�'4�ޟ��'5Zc�J�B8�G� '6�`� �O,h�;O4��?)��?�,Ob��G�h�H�[6�η�,�A�AXɌY�'��ПT�'~r�'BR+�x���0��G�;HNl��aL@���y2�'�B�'�削(.)��O����@ɕ:�lݨ'±~zA@�4����O�˓�?����?I�<	C�K�U���1������A�M�#���<~�����ݟ�'����S�~r�U���@.9w3�LK'͂�A�Y��iz�_���������0R�"�O��V�W'��ш�+�x���ٰ%ۛ��'ir�'0�)'.��̟���?=:�NO�9��eb��*� #�ē�?)��gcR�Dx�؟Z���!��)�$�����<{�\��[���� \(�j7��$�(-0�e�G"�#����dNQ�G�!�D[�-_�ؘ�dQ. ��UCӨ%����Ŋ	aX0�@B!�6S)��ҨX=}�H�ǆ:(����A֦9��ep����&�zc�.��Vb� DܟC�iˁ-�+@�Z9:!��|\���䭒�
��h�+��~2�u/׸�~x��eZIr:�i�!�^���	E#�uy� �(D�R��O���O��d��{��?���o�
�A� X�.���
�+[�NLM��0d^���*>�p��g�'�tx�/7A����JB�Q�2Y��	�O�̲�ơA���sw�ޝ�����@�?TT�3�@6:t���O߁~���^�$'"�'�ў �'���27,UB�e$��'F�& �'u~8Ѝ�)ci�<I6H��<!$9�8��|����	�u���n�?��ii�D��޾����/
xH���ٟ����xx刔͟����|:v��`�a�phR�evL���D*6�fa;��7��S5AJ��<�Q
T� �^Mb6C�W�1$Ck(mK�M7'8Ds��M���<q�M����	 8 U-ږ(�BP�p��h�l�D{��I?�0�pF��>?1,L#��ԏ`5��!�r��4�#L��gX:�$KL]��ϓF=���'��4�P<ꭟh��|�q��A.�`jGl� ������O�o�Б����?q��qX&�U�1~H�T�J� �*�� H���kZ)xJŎC�GѴL���ɠ^���Չ�Jd��C�N�֟�åk[�\��L�	�T0ʣ�_"��J���,u���O0�?�IG�P�T�Y��^��jx�\����`"�g�U-o��-�׋�%+���hO�A�ɏs`�	d�8��g� �V�I�s�����4�?����	A!��$�O��J:��k�A�3l|`�+�70��
2���|8�J���T>1�|�	�y��|�H 69���B�FW�&;"`�̇��Dܢ �V0	�)���*�Ũ2�ČW���(+QN�.1P�Iğ���'��B��<�BI��3'^7-x�ȓr�V��&ő%ɪ`ˁ�ëU��IGxB�-��|"��x�W�X=Ti�fh $J+�����?�S���y�A���?���?�v��<��O� f@̣B�,��׌�r�nӇ�O���$�'\��v)�,���!5k�0I�'���y�x�ȔC'�7]�����S�4}��"����[������-&&^x��)V3?lX���+D�iS�$tR 5���5����AH.�HO�)2���2h��mZ3
���`�E\15�~�#g�؂$��t��Ɵ<�	����6&�(���|��	��]��.�lWx��'ݶb�:�`���4�N�e�'���d`��,�Q�G��B.A��&�"<I:�(E�B�Ev��ĉ���'0f�����.K&}�6�Q1Nh9�E�@�'�x�Bυ5�"(�ì-Tx��[�'�� ��܊y<z�$߯au8x�'�06��OʓYTB����iB�'F���l� l�M��jg�Ԣbϰ��ņ͟�	��l�D�Yz�X�̉�FM6��S�t�ےK����%���0��)�_�(OVYy�A�j�V�¤��(�B�o�+� �RQn�1'Nx��@�\`�<�1�� :�Q��C*�O|��#�)�OP�4&HF}�ه�	h��I�O��"~ΓLֺM��b�w�P���<����'-ў擣��T��;DI��j2�ແ��?��M�<�ꍠ6�i3�'��S������П ��&]�e0��E�Y�-��a�S�P-·f�M��<��O��h��(�攻w��3FP)��Y8������O�9����]��$��W?���ce�� .����OB��?�F��D�%:�"�w�\Hhp�8�ϓ�?��C�� �����74�k"N�q�'�:"=�O.��$E�x9���0����"&�'j��؉"j���'N"�'"�wݕ��Пؐ�W�}�l�p��2��������?AŊȠ7�H��Ŷj�n�3ړABTq�!D�H�9�ň	�kBl��b�'K�Bb��i��P�5B�fF{�+N��P(� Д6by��f��~B�B��?���?���U>�Qf��O�ޥ�f��v�l]r2�0D��z@HZ�ʹ���	:\z�P-��HO�	�Ofʓ	�0a�i��C�Kˑ>��Ջ`,�=1@p�Q�'���'��e��	��'�rLħ9+n)B��F'G䶬��g��Bd\P��*] 
M4��]������=F*��7tSS���/�\�DH�u0�J4i��p�F�O
�DE�v�D���N�F���fݞsS�8l蟘�'���4������v�B�S�N��̒�+��N��!�I�6Q4չF[�S�1x$���ئ��ܴ��'�r�|�N���Fg��Zj��4�y���s�jP�$�Ƚz��Ǣ�<�y�m@�udXMRCǗ��p�#����y�-4L"��������.O�y�MC%���0􄄧KP�S��y"��$k]6��v�Q�r�ra�t��yR�j��̓r,϶zn4��!�:�y�!7l�9BU�t⨐B�LV%�y)�q1d��ыH�r�J��#i��ym�erb������x%^$)�W;�y�`	�W����Ǒ�hp�t����yA�8���[�,�d��wcM�y�GC�&�d�;AndZ��8�.��y2L���� "� �i�V�n���!򤄓Ay���C���8�T+��t�!�@�n�7�k�H- ��Վm�\B䉁X��y`���m<ZW��r\.B�ID�z]���
�g� ��D�E���C�	�^�3v�p��D!*�,7�B�)� ^}���E37Y���$:<�T�G"O�d��.��T-���!4"O�(:4K�-)��P�TA�!,�t��"OR����/��]q堛�u��+G"O쬈�aE�1����҅�+H�DX�"O�k�偞8�|�{���5w� #�"O�ѫfHʹX��l����=qP �"O,$`EfH�z��qBoB�$��9�3"O�����L�ck���L\�tנن"O���s�f�D�gLYP/<%y2"O0�g㘉TYJ��m�;�"O���a.�:K 
��!nthb"O�͌+qBɣ�R+5��;D"O�:3��=v��EB��Ci튤Y�"O�%�m�CO�(�Ge�3}J��'"O\���c�3�d͟^5����"O�q��T�2����E����Xj�<OX�i���X���`��"~Z�$�?�<�SE�W�	o����n�<����,\O�g'��"3l��Ëe~��OMv����0<9$C�)}�̙
�
J�'�hh`2��H��Ypg�#�^ �ȴgd��c�-x�A�t+�
�B�	�vi��K��	+��!�K-o:#>aS.�}��aabD}̧3�|�%yn�@��EӚS�.D��D�Pk`	�=�J�J���ky��͓���èūp���秈�Ft �ė�&� � I%��L���'7VT@s�� `������ߙ&v�y��0Kj�zo��9d�����I,���Ň�9猼�gدBF�?QpjN\��[!���e��V����է��	0D�0 HH(��C<9� #&�:��@�5|x5ؤ��uy��B�t��'O�8 D�Qe?�|2�뇠)�a�􇀨G�x�1� ]�<y!��F�0E�y����e�<!t'�
Wl.�	4��T>���`�|~"G���r6�/L�i�-[��?Q�G�%��Aw�K>e��T9E2�T���b�>9e�˓ :�A&�n�D+!_�`���K+<�t`�5i3�x=��3���>�BkӤl-����Īw�~�Z�m٨P�,�hĥ
�8�P����@��A�����X6�}j�19Y�ٕ'Rr��w�Xb}�Ȗ5,���S�',�q����(02�Ȋ���ąȓ�2A���W�N�}s�GQR &�\3sG	Yay�D�����ү{;02�΁��?Y��@��#K�A�ܩBW	I;1sv@"� !$��+B�U�w��D"�`�2B��Ȣ�&'��S��R��1��� ��9�5J�~p"q�L3*�H�D��#�~"�,v5f���? ��R���DJb`�X@H���5���`L����%��'g*�;���.q��@���&�y�#�?y�Ik���U�tS���5�~bDJ�DF<��3���IF�`'?��7���	��ӟf�rA#�	�$gvlD�kMV�DB�ɝb�bx��ǂ0�5X0H�?��x�E�s���Ѣ�5g�?/��I`pF'��4���L=,����e�j��)��	�V�2���)�䎇��Y�"
DJ�-Jf ��B��yZ��Ӭ8v�)�(J�P�F|"K���4��=t�$���1ᰋD;���7�  ܁�"O(M!���?Tݢ7� :��:O`���K�:ZPĩ�n�a�ā�7.��a+�E�� 0�F�y�IX;B��4k�j�C��R�l��w�����dY�$��'�N���OjLy��Q���]A�B���M�1�'m&КSk�+%�^�R&�.G�H��B_([7����%�����ɫf�Y3�	�f�.���OִI��#>yф+ 5Մ�X���O.�!
��V�J5K��R�(�J�'x�lJ��F�|�@iӓK�t����ن4Jnu��/	!6<��G8+��m�S��ߡYegOTt��a��׫G�Hm�U�;D�Ĩ��ű	ZL��3a:'TXŊUU�d�4Ψ���O�p�AF��?a��'��H4�q�� Ku�K�&�ƕ��yr�[�fƔÔa����O�š��ڸ:x��3�Z�x1 L>~���y��G}pP02w�E��ģ��Č8 ��!6 �-yX���C	K��h�8"��">�!۝!6x�S�? \�G(@?j�=�p.�:Q�x��U�y���.OD��d$�\��V)�c-�@�=�:��=y����O� p�4}�� /L2�gM��R�ܐ �)��<�3Ɗ87%�8�%	�9���dE�!N�ĉ!AU9u(b�IB�� 1Ve�x&�:CI�˪OT�Q�*��T�D8	;�щ@i[-{��s�,�z)�`��>��
I6MtR��
Cz�(l���1OL%*3�H/,F��G�_�C��I+$�]��D��f�O��:����&zL$(7�X4o�F��C��ަI}½��� �3HV��!#G2S�l��/̛�
8�Z��O��h͟����g�:��1;�O�� 8W�ޅj�v�����;$�WPa���U,̜iyz�0GN
zM�B��2OfL�ѯH�2��j�@:_�t�o�N���A�+��YՀ��\I���䅮Y��h�F@�dz`�r�G����S&�ӲgD��j�\�Uh�ɷE�<r� X�F�P�����˦I���	�'.�(�d:u�x H�j
 #�ْ(����s̓hh���"T����qB�,�<ySo�F7Υٶ��-0B��C��VAiv�T��M�J`Ctq+���Hn�I�eK]ܓBBy �mZ 2A��@L�v	)�(�'2Y� ��-4A�Є�Io�~E�&BC�|RVX��H��G��y�u�O���!i�e8���Ņ�|!�Y"�%
���c�#,O�(�F�%+
���Ð'}8�q9u(G;f�6� �[b����:���ف��L1��8���4�� 5/O��Z� �$Z�՘c��� R�&�Mn0`#���6�G�Y��EiҨ
�)� �@���.�c��/U:�`��O�o�:�b���H�@9�� {F�9�<�W�߽ (���-�d��J�$V�Xu|�ɿ,I�%�D-G
fq"ĩ��N T�"<Y���1�xI��Ğ�s@�yȀlL�U�
aD��J��">qvX�?�_�Mq�S5A:y�����$����P�8R���,`���D��}�Y
&�T:������S7@�4�'�d6��] ���*�s�֝&I{�d!�Iب]/�͋���"����J$lOڠ�Q,ƒC\����C�"�Q�A�X�@����Z|� :�#។��dӼ]m?{ ��V��y�gd>˓P$UQ��+��	����G�pe�>i%���2A�PM�<�W�擾9����2�F��d��j#8:6MF3�f�*���O\� f�'8 �J��[��p��9�hd��R�t@s�����S�	D�W���b�w���+����G��a�_�#3�f�^H<Ѱ��?L�Q{C��%F8�Y�@�K��	�w$JX`�'m�iZ����Z�4^����ӌ�7 �(�+��pg<���I�t��9�!ϟ��w,@�qO��B����ܤH��!�>y��'nF�0pf�t+���e[��R�Ez�
�3w#~F����4~8�=B$�M%�HԳ"�Ǹ�yb^S�,��LU�*-mbRDF6�~Ro��O�>yYgH�d�����ԧ"Pp��B/8D����/� ]�$]�T�s�\4�rI+D�X��.Ѐ��l�?XM��(D��J���b��]l�57����"D�<�����:l8�+�4A�l�D@,D��X$�.(��dƊ �{
����?D���ѡ�:�m��L�*G� �k=D�Љ'@N%�V����Au���!��7��@q��z"��we0	F�R%{�$)�C����=��M���?9���s��*��Ѓ%H�&.���b���'u��v�0\��5`	#C*8y��dI#��,e�>պD`(��yx0O7".C�I<z�rG^J��=CRb�NGV��ӡ�O�U�K�<���Oָ������D��#������"O�1��(�AS�� e�4C��'��-���'6�I��'6x�� ��z��0aN�x=F��ߓ����y&X�@K�q���լ��Np�ɶ��y�#�0��p�l�6
��;3nҌ��Ol�p�<�'p�&��!䙀Iϴt#�j�H��ȓi7�A��t�����<d1p	�'�]x���Ӑ$�*L��4v{�S���#�HB�I��qR`�O�B�qW�'k:�OR�1�-LOĴ�7K�Z�d�9V I;V~�lsc�'Ԕ��K�t�|����ɲ+���GD#!��͡��Q���O ����F]�\Bax���7�OV�� �V5TR�����*CP~�;C"O @Q��68�mԋQ <5\x "O
(SH	� �~U�u�ֺ\@��"Od�A�T1�\`�藸y�n��"O� ����l}:D�"��"OԽ�EX�|�bm���8	��(!g"O^���&l��,x���-Ѵ(��"O���Z#dl5K�c@cD3"O���d�	{����ȡB�rq�'"O��2rVH��}�6�W�}�,X�>�pmŭJ�O���C�g�l�b�A�N�����"O��8'BR/#\�Dģ�,�F�ɤ��FX+�DÓ�����*�����D����y�襋JF�b��=�s� "i���A�R�|�tB���i�ڈ�*?z�����ˆ
�f��d�\���Z�yү\%_�03�L3a��:����y"IJ�y6IÑ�ә#3��
�b����ɥ7Ovȑ����E~�R�B x.@i�h��NU!�C�Pc�X�L(����\d@qO�X9�
0�0<�+
�F驡	�a����a�P(<����@��0,ԑXQh4�:�D�p�%�0��O51��Ra(ڗW���� O��`BJ���'���"��>�~TǨA�Vݜ1��'$�h[nQ YyV�@���P���I<�F�9��O���Q�%���4�h2�:8�:��3"O��A5�B�*V��b!XG"O������)'�,���
�И�"O�U��
�	9��Sˍ.9�4x��"O&���#�-c�� L�w��1��"Ohu�tgY�\^B�ʐ-G�.���"O�	�c�B�&��\��BZ��̊�"Oa�e�҅O,�0�ϥ0��	'"O�}�#�6u4��p�uH8��B"OX][�9��ћQ�-F�`��"O�M�EC�>V-R�0��ɳ*�h�# "O\D��Ct!���,W4`���"O��hS�&i�VJQ�<t0��"O �ۢ�>Zp�ꌘT:<�r�"O2��a�$���GI$Y,*���"O��ѱ� �%tux��B�I-��"O6����M�,r��b�Je�`"OV�۔�Z5
d���%2|�Z�"O`�� N0�p$cRgН,!s"O�2o˸¦a+����P�j ��"OJ|��؊%2��n���ٱ�"OBU�E"�LT`vm_4X�� 9e"O���D�_&\���A�H5$�JА�"O,�cG� .D��y���'zRE��"O��#գˈ;��cFC�h>!1E*O�u���09a*`I0��E��'s�H���V qS��c�z	��'8i�@b�5�p��R�Ba�&i��'�(ț1��)G �7H!p��I�'�<���Oܮ�D��F�'}G\�z�'�b$xp�D]�ٸ�fR�G�@��'�������<@�
�����5R,t�'���� �^�^A0�"K4a<e�'%�,[	�!�H���
%hd�a�'v���ǐ�omչP��p �� �'v^Mѕ��H��1{��VBB�C
�'vXd)Vm\?`����F��P�9��'e!rEY��ɋ��ݻL�~Hc	�'N�ZS��"t�j���m6��@z�'#�h�Ik)$S�T
9��yJ�'��!6 �is���F�
E.���'� ������w>5I@/Q̔B�'h(�����^��K��(JW��p
�'8fU{0�S���\�协j��uQ	��� �	�2�̐8,٫2E�4h�vQ��"O�3���#��`���(.�"O4�ЍN��ؕ(T��s5ք3�"OB)����W� Ir�#j��H�"Ozkv���u� �0
�6U.ر�"Oh�k2m��4�|��"J� X�=3"O���DBy�@f	����"O�Xh��ɪD˒��֧<f(Yj�"O�C�G.e�⹀�)Z�P2���"OL�ٶ��`�X�H�h��	�b�rc"O���⊁g%'([JtX�@�"Oؙ��+�����i ]!�D�6F���@*��yjl���[�P!��H�!*���v�<Nf\�a�F]I!���ޱZW� 8,H�9���x-!�d�K�|ݙ�ޔ _��`�c�#1!�"��Q ���n@P%����y!�dB-�@I�l�((�z0B�r!�Ă��p�"L%�B�����&&^!�DS=8
�kq��ȩ0Bоu\!�DHb��=�1IE�`@t�V�;O!�@�HDS%LK7w����@K:S!�D��CJL����� )��5�`_�^�!�D�Fhbx�P#Vؘ�X�/Y;!�*����x!�`�� ,�!�� 5rPa���j␴#)̬
g!�$B9��ݣv$�IzЍy%GQ'gX!�D�v@����=1��a��f�<u!��Ȕ(]���de�D�$��Ȇv]!��9W�H���3t��!&�ۑ?X!� �_������ْ{g��v��?:!��f�9ULжE9֨P�G*!��Į	u���������&(�� $!�Ė"e��೤��C�x�r,OQ!��U� ӊ�3���Jm��KR!�䜎?��X����"L ���CB�!�$����hZ��Y+�$�UB��u�!�ۙ{�	��n��r+���!�xD!�-��=˄�C�����@�=\a!�$�;I��� ���!�sN�,`!�-:�"̲q"~zxL���˪s!��;x��g��xڞ���-�<r!��<5����wH�?^󠍜���~�P��4�ЇK0:h2����y��7D�肐"�67�Z��F��-!�@���+D��"Ѩ�`��'LK��#��5D��J�b�h4;q�ĉ*6`|�q�=D�d�5A�I+�ڴ�OVl�{��;D���v��,z�L�1�Ωmr��2�E:D��R�5�(��̔�И铫9D����(Y�yqh���M'�C�H6D�T vC�9Y�q�#͖<G���c�2D����V-�&�X�@ʓf�@= ")%D�0�S����%!o�!S�6�Р&>D�X��aP&r��v,��rq��6D������q"tC�@�	J��� � D���ǥ
,�Q�a��wڪi�b:D����D
;�r��P�@��!Hb�4D� `�d�'V7lk�iA1jr���N1D���@�E�e�~���[�H�$�lp�h��I}1`D��	�)Ǯu���j	C�	
7*�PЇ!�.Q�u	��F�0��B�I�@C$��mZ�s��je"E���B�? ��5b�M&a���Yk��"��C�)� �Q�.�5.s̱sы 3e�"O.4Z �VN�ig��9P���"Oޑ����Vl!')�ɳ6"O�a�u��a��c��S��l!C"O��a�j�4.�#+�Ȃb��)�y2�Bv.B�%M��d��↛�y2 �R-���TEP��8t��M���yBCS�g'Ty���Dt��ި��%�O )�-O�pߘ�x��]�V>�s"O�h �.��j�t#��!n$>i�"O�`�Ŏ�>D��-�"� 	�˗�	n���)�[�bI��,]A �;���"z!�� ��Tj�B'e �ы��L�<�!�$�Rv��K!�4_F4)�$>]x!�d�x(�0�䤞?J �l�B�->q��=E��'��|����.�v=�����	��]�	�'�Z���	j���J0V�	�'�h�k�/ȏPppa��`~�X+�O��=E�$��+iQ����ɡ+��ً� ��y�\j���O�)7O
ɸ��L���IGX�`3u)�+]�r\���
�XǼh�J;D����حR�69ٰ�&������:D�laG���^lz�	V���L� !�8D�d��ݒ7��8���2dj��D3D��B΍�	�M`w%��6"i4D�` ���[�̈�6O
�aN&M��*&D�̃�+�HB>����/Z
m[�nȼ�hO?��[+�0�I��! �T��lܪ|&a~�Y�dS�F�d�N��쐈1|��8D����5�N8y7nPsRhaE7D��ʡF�7�@i��?�T���*)D�� ˝9���&��yB`<�Q�1D����7��0�M�P�^h!1=D��h&��n���X�E_�,�bq�0D�����֠G��y��F �C��D�b�,D�d���(tF���3 ��4 ���>D��h�f�z�H;t��>z�a�n*D�X %D�c T��BH�F���{��3D� ��#�\���I�#|�ޭ`-1D������"�؁�E�!0)�:�)D�8�C�!�>�8bL��e����w�2D� � ���`��@����Δs�@1D��0'k�38�3�.�f�}��$"D��!T�Q �5Z�NO�$�ne�G?D�D�T�O�(�����Ad�(�b`>D�H��䝻e�<��/�t�"�
�;D�����N�/��|#��t96�E�9D��z%�!#!�%j�n
�%~4�b��6D�p�ص}9Q/M
�6)��5D��z6fќ&�4�KS��T�����0D���ˆ.x6dA�`jקS9�`B�(�O��<ЊȪ�ꭚ�)X5!i���Z^*m0 $;�N,#���'!@���]��t��X �1C��1�L�ȓ�Fm�u�-i��IH��*��ȓ4���h�NZN�)���ҽ 7nԆȓ?����"&I�~���Xw�5a��1�ȓ)�8�[y8 �&�_�(�h��ȓ�~x6�D�e�*)�s��H�L�ȓH�D�:�b�/EV��n�[�Y�ȓjl����	f�6P�3�ݎC�d��r��x�gW�L:�%Au�B|⮰��tgh�����:�XI���
C����ȓ�]U�O�L0ݸ�e[؄�S�? 
�`S��M�Ј*d`�8o�"�ٱ"O�����U�Py�u�I�H�s�"O���0c�7co���c�o��b�"O�1X��b�8�C:u�.�"�"OHM�*�%�<D�Ԙ5���"O��HT��;G�`���7J�`�"O\ D�z� ��&��D��iR�"O����\ l�$���ۚ8���ا"O�XJ��X.A�5����/��E�"O�,1�(ZK׺-J�×�k4���D"O&�(�k�L R�I�o�y(�"O�`(q0I1���q_�E	A"O�������U����!�PG�]�5"ObH��bϝG�$}�T�#v( "Or%Ӆe�*|��Ĳ�+��U0�"O�m��� a�ܩ���A4G�z Y�"OJa	�(2$x����;��Ih�"O�(�G�@ &lZ�E�3q�ڰ�"O�X�NM$.`�����-z:A""OX��r�\?�.e &��=9�Uj�"O$�+��E�\�"e&F�",���"O��#�g�
+� Y�J�5 ���C"Ov@���O'd9�E�HY� ���1F"O0�1D���N|3�,�7Y���*�"O,҇͘�2wZ��k�-wv"��c"O��K�W,�1)��=-o���"ON��֪߿03p	sQ�5}m��'"O�(���Jt-�R��.KZɉ�"ON�Ѓ��\|��o H-nG"O�0�bk�/TT�a�K�o*�H$"O���W�]�Ҍ��E�fun(Y�"O�i 0�v��p��	 `{����"O�s~�M��'�z�J��%��`�<Q�Z�\����g���&��"�EO_�<�Cg�h��8��f̳����`H�Y�<�u�L�8@�<AU��8N�a�Q�<	q��]C��X�*�,�Ġ3I�T�<avo.l���H�k�&O�PШ�ES�<�w�ϯ<P�@x�'�#m5��q�!�K�<!g �%z.I�
@(~���P5C�I�<�`�u�P�Rs�-Z�����M�<Q#�D�j����؄G(&1�ee�<�R+��"�9���[�>����c�<U,�j� �����d{��v��e�<9�B�9(��u�A��kJ�;��d�<1���m��T�v#Rlś�K^`�<��P  ߸���l��;p"d�c�<�A���V�"=��� 
�&�SU�Js�<�"�R�W�1�g���k2&I��+�m�<����U|&���G2
J`���Op�<i�M3[��|Iv�P���R�ʁa�<��^;�`�h�ā)@����+]`�<q���f�����f=?+@+N�C�j�R�3���]
���D�P�2C�P� ��ݐ0��h-DfC�˖�ӣx�^h�G�Y�FI�C�I
!�X�͕11e 4N¶^��C�I�0a�="F�Z�����L��
�|C�ɞh�@�������;��A0 �FC�I8�41�'o�:h�h�F��0��B�	�
mh=�p�L�p,�]�7(�#��B�	"�ح�BխCZ���p"
�96�B�I7l�@`س'�S}rȧ���*B�	)^��a�@�c�2�����+VB�)� �<Zp[VFy1��2O#����"O �n�PC�@��ܩ$r�D@�"ObhJW
ܺ/DxR���$i�tp#"O=iӃP�D�jG(ZJQ̠�"O� �e ���"��T�4!�s"O|�9%�S.;YJ� ������y�"O�4�7`ؕ1�\�2�᎓2 �4�"O��j���1rL�󧁈�1�D�̓"�4��R��#�M@���F�<��)ߐ��P��� h.ua��6X;ȓT`�(Ǭ$��X����'(�����+@�x�Sp��"s'3@VD�ȓK����4�=C2� (u��x�B�ȓP"b	�h�"	V���)��Z�ȓ'-�!�3R2��D�0�^�ȓ<��i���7(k�АƏ�	�	�ȓ`+�)�p��SNB��Ubߚ2�|��c1@1n�3,��ŤU<�^0�ȓ$$���EDV�����:@nA�ȓbd�4
��ɃU#.�y��<�Ņ�I�~�	H o�j%y���]0��ȓB�(tMU�*9�P��
�e}4фȓ8p"���]Z
9�Ы�
D⪔�ȓO�YQ��a�@h��i�=��4��Os-Be^�k�X��ЅèT��ɇȓoex`�D��
$3��3,�	b9)�ȓ5T$�"QOG��6���+y�tx�ȓC���Cު2����-V�e�A��6 rTXU�QU�j%�ԢB'R@�ȓh��}�f�_H�U0�h�$rDr܇�|(p��S�f��% �W�.X��ER� bД��ys4#��@���ȓx��P�X�0��p��&�$,l��;LIx���l��U��.X�I後��;�0�#T �)3�.���X <����NI)�f�%����oʳB4lцȓH(���I$W$�����
~-��b,�J��5,U�f'�Fژ �� �q�����Z��rh���.�ȓA��J�4m�l�j4���/��ń��B'�6q4$`��M5�ꍚe/�G�<��*O�r��2��+�����\{�<�A�D&[	ZYIQ-G>J(�����q�<�����B�1���3D^���k�<�7�J�αRS�ڬJ儸�b�i�<��D�π=�fȌ-j 2���A\o�<�Ł_�h=2!x�@1,�Вt�F�<�����Wk��pf�
�<��t�r�JX�<G�	��Å�ͪd@hB��V�<��B�2��Y a��	T�<I2�&�Bx�FKz/�x�%�S�<����b��i©̚$a�(�d�P�<�0E �uP�{!	[\����"L�<���w?�٣��n��j��J�<eΛ*#d���@�U�	�I�<Q�.L:Q �b(��o[����%HE�<����)�L"7bD'=HP@(�u�<�0�fP`�M:�"	3�i�r�<��C\�jb|C DV�E4��t�<���6�%���	�_w��)e/�s�<�fa��T
������4�x!��z�<Y%F�R����� y�cPw�<��d�"q�41˵.0fqq��N�<��Ə�
�9��~�|�ڕ�Ea�<� ̈� �]�u%�)�$�-u�C�"O@8j��F8w��K�)D�hc���S"O�pjc.�^����ɴH}���"O6!2/�2z�M"�4n ���"O�4�!@	&;B�I��;�np�"O�e�P�3z�y{F	/dߜУT"Ot��d^!5�$k&�M�x�z)Ѥ"O0�$Bo�p�h��uР��"O���L٭�~(�A�ȧZ6�W"O������O�@ "��!P"O衢ϯA������H����"OZ�0�_�~�8(k��֩zY��8�'#l�c��ER$Jw�P�9��1�ȓ�ձtM^�3�~�9ԏ�	p��q��=O�B�M�O��Py"o�,8�Ć�����Pk۰v�$A�$㙩H�ȓ;'Bq����.u��(M-*���ȓt@`0d�p�hY8"�̭_��ЄȓkrR�� v3N�c�ʛ-6ˠ���m��͐� �4��k"�_-~H2x��B&�-۶�
9o�tm�0�Ʌȓr&������<���L�l-�\�ȓJ�\�%���	��s�!��. �U�ȓh�~qZ�Lۆ�l��V��H���ȓ"VJE���0G���j��\/m����ȓ��[�x�ਠ'���v��ȓ!�>B��7!@{'���t,��:�b�sƥ�.ah2=�#�O:�U��HQ�xk���2�~�A�\%n)�ȓI�y�vA��*DS&��Cx��ȓpS�5�@�]N�s�"P�L�v$��e����֖huP�JG�ǌ/v��ȓj�f!a�!6��mz�GN�,gJ]�ȓ�~}(�;k��Pj��A+~�ȓi���� �5tOf1�BC�&n$���$�t�&k�� L z0I������V�:����)�D艒n43� ��nv�d��.��a��/R��H��C�����)X�-�r|��C�o��}���Pm"�l����9�
�+T����ȓS��q����^<��i�^(H���ȓ'�BAi����+�؍���Q�`�Jфȓ6�ʸ����%1���J���%�,Ąȓ\� �����[e����&��L��n���SlߝZ�B���nR��ι��2?�x`�&E�V�q�KǱr�8X��x��rN�T�C"�18"ࡇȓ2m@` &J˻,�Pl�G�ѩ#�:�����p�G
�@���%^,���i�(����"a��ۧ�� QrX��+K <� ��:E%rQ�
��O��ȓL?5�¨�$A����be�t��-�1Ɇ+��k�"Pe�l��ȓwhx3A������\�&��E{��O5 �5 �o��U��_�v?�h��'��E��H�8��!(M��k�B����0OD\R�b�-�0v�(�b�HB"O��(�e(�T�A(WL(	�d"O�\a�D9>�8��P�V�j���"O$�a1m�B��(��Ј�`% �"O�}����=�<�cc�.l���b�$�O����O #|�,O4���K@&��ÚJ�<a�8[[�lSm�
��BѦʟF{��	\���hڰOF�M'D���T�05 B�)� ~l)���Ĵ�� �Q50��"O|8wϓ�apָ�AȬ,PB�"OXh��]�ȡ��N��A���"O��[�j�� �Hɣ��ˣ�8��w"O���w�'�D�2-G�N�q�&"O,�s��{P�\X��!n����"OPd��U�@�1�$m�5{w�J�"O4ݪ�뛤>i�9!�M+FZl���"O��@�Q�1�0�̙<R��a"O~��M�5ui�=c׫K	qG���U"O09���v��YF��>|8���w"O�	S�%5*���P30��a"O�ES�ЗR�D,�p��,�T"O�P�eb��(7�m+�!2����"O2���2  ��*�@�((�S"O��S0��G�i�W�֣>�T�"O"9�eʔ{��l�0��M�F5+T"O��A�ߺ&~]C��T]������4�S�I��l�(�8S��!l������ͺ�!��[>�^�3V#PW'X1�� � �!�DD�P��͓1� *4!����[�!�$��!,2�Kʗ�rT	g�Ɵl�!�$ٯK��m��n�����oM�	�!�$"/K��i��[�@�!D�V'�!�dFZ�`��%�Hh�BV2�!򄜗sLd�0��,bf��B�o!���g�ę�� "_4J���-<!�$_�($4y�I�q0����!�D�#%(y�
BG�Z` "�Թm!�䁦A#(�"�Į\0�#��<!�R�!+��"/����ވ.��'9ў�>��6/H�x�D��e�B�w3H�R��*�O�扙p..5X4&�,S2��P�v��B�I�8�,@��%^
F ʢ��:3�B�3�117�M ]�4<��T� C�I�3�X5�+��n(	�6�TC�ɜ��R" 0Tˊ;T��u{(C�It<QVe�GZ�IR��.*��$|��AQ�/`�z�����6�<).O��=���!b&�J�]4)C���c�!s�"O�� 1*��H��գ�c?DS�T��"O�� �_��9Um� ��Ubt"O>)�B��6�^l����4dF, "O���A��)AA m�/,t��+�"O@U�$�ޱ����D�S������"O�Бr���0�IT�G"qzM�5�	f>ə��e�H!˵X*��Qf0D�D#vş6e���� s֬��`"D�0`��G�0e���e|����%�<�	�?���N wtyR&gF�+j��w�6����T�u��ʎ9�u��X�����#ϔN6����ϋ0�����a����8񀠤A)`h9!�(�m�e�0D��(�M,\]�U����.[<�@���"�	Y����''I����
A&,0#t-ȦC�$B�ɭI���ywe��.6��c脂	c�C䉍a�֭Ѥ�� ����+9
�C��O��ْ��-Ez�fĸS��B�I/."�x��g0�E���_���%��D{��DGT�wa�P�V�:&��``$�?��'����w����1⬋�v���8I>A����5_`�����=5�0�!͓S!��� �z1�5C�"�5H��]�!�$�J�"����¹p2l���J¶d�!�� PT�EM-p\��b�C�-�q�@"OTruc�/�:x���4O1���|�P����W�R�!�ߛ:�<�%G�;Oz�B�I�{fh�z��T�d �`��4	�<��D{J?B�J�c��
��Io.��B��&D���Bm�_d�����E
�4�&�.D�P���4��%"��C%�8h��:D�(�'ި����g�ޅ*��h!VA>D�슳�W\ 
M�p� ~�x|+��;�O��m	~e�#��$v��* 	��
T:��ȓ>�b��Vn�����=�}�ȓX��$����5x�6�PѯȪ{�����l~�׍\�*)���T��m��&�/�yB(J�xz�h+�Lj$L8q"�y��hb�$�Rn�P%���a���y��@�S��E�d��M�d����\"��?��'^N-�Q��%�F�A�	=�\��'�x�2�M�$=��y�Cg�(N꬝��'�ы���3Ȯ����
�E�����'�J%�u���vY�N�JK�5r�'� z���D�d�@�E��5��'�9�uC&QB�"�g2&�db�'r�p�k�/)æ�+��  �~%���*�	ӟ(�	�!�����(?�~����?uri�ȓ0`��A(8��u�Q ����ȓ&öP�D���24�'�"B��؇�	�<	�J	�����p�M�u�<��VNMLpp�!�1f�,���K�o�<�o\��V����n�K	o�<�a�_#f<&�:b��-	3BY�Q�p�<i���-%�X�h��*ܑ�D�We�<1a"�3*���;�|�aU)c�<a'�}����v%��ssR`��lΓHEX�HL�.LI��EL~ P�IP(<�g�Q�U�N��L/i~� � d8D��PB��W���(g�)v�P��u�5D��Y��_y9(���-t��B�e(�O|�"����eU�t\ҥ��NO#wf�˓��'�ў�sdJǯ;3�&�4h�d\�dPH�<����v&�P��8	Q>��b$VJx���'ptѩ&��g;�8"�(Y��6]�	�'Ƞ��'I���,cG6��qO]H�<���
T���k� �7�jbq�Ah<!� ͔g�>����}�)�tm���x�����iÄ��y���
�ўD�	w�O��� ��®`b‖+szƬ
�'�p����/JO��F��r6b	��'C�܀�I��L~�P�u��g����
�'��b�O�XG:9Y&ɟa�|
�'��2Gʖ�GH蜠⇀*m�<Y{�'[�E���S�
p��QJZ3e��Y+�'Bݩ�E��
�h���̞-
(�'q� ҷ�:|[ Y3p�S�TS
�'&^h���O	8~pu�F�L\4^q
�'�`TX�g� <�L����YclL
�'-��	`E%n(� eV�Z�x��	�'����]9Dt��g&Z�&+~��
�'�.�	S*S��5 @�˔0��	�' ҹ��d #�`��'<�L4@�'Ū}�P�ä��i��*�34�T���'��C�(m�.�9t�A�/(��p�'���+Dh�;%�bx��ŭ||
���'e��ƈ!x��5����hh���'�X�1����� �b�c�F����� ��9b�\;
�����*Y�&��%"O��AW��_��I�aJ-d���7"O�����xin��6�ˋ*oV�Ѥ"O� ���Kn��t�21;�p"OL�:B헭T�� e�dG
�I�"O&|����R����4$Ƽ>�b"O���-��J�UR��G#�I�"O���oG;U9Dx����K����!"O~e+ �(B(�=�B�_$gDB�r�"O����Ў:����ąC�{B<�"Ǫ�Teئd�����#D�P�Y�"O����V�'�tY�d�
ƈ[F"Oy��b0%�m�e�"=��%��"O|��aH���t��ȄNZ��["O�L0�OOb�T�B��޻!H$�"Ol	�r�GO:����	��$=��ڳ"O����	D'1jy�'"6���s"O�8�朂)&�� �
fr$!0�"Ox��@[y��ա����6˪�a"O�D�#��,u�z)CW阠p�4�ӡ"O(uh�Q%�&�q$��)!{LU@ �'����%�� ����F?� HZR�.D��;�&3# mz�OʓJ\���
?D����c�z`0�[ �`7��;�&=D�r�0t�⹡hRX���0D9D�8�G��+Jb��i�g��uh��2D�$�&��73����MޔP�a0D��ARe�&[����$L��X$�./<O#<���f���s�%C n���" ��X�<YF�+g�Y���سSnPt���X�<��ˇh@R�$bް"�\��S�<�W��&#��H�k̓E��`�G�^y�<��ƅ	�(���� i,����y�<Y�oA/�J���U�#ZX�1'c�w�<�֥)/�P�;��&���� Mt�<q֤�$b�QG�>p���ɔH�<ih��?��(�E�^��J�C�<QR���6�ȅFO>cZUQ��Mf�	t���O��З�0,I�;R�F,&z� ��'����f$�n���j��
z
�'����E�Bl�>�Ȑ#.1����	�'�6|ye�7dt
P"ޑ+���A	�'�@a�4�/���C-)�}��'Ϟ�����$�DM� �2&r��0�'�!ԅN�N=sqe�m�>`Q�'���&�ZlH��E�0yZn�P
�'�.��C�ˆ���9���	u��@�'Ԝp��
l���CAcS�斐{
�'�bĳ�i���x�1��U�訙"
�'5�ui���j疉����hwx�0	�'-�mV
I V���kSN�R�����'��D+$���jP��SB�F���	�'��<� �68�ICh�-��:�'/����V��\6�T�.?(��"O�,;+�1mb�s�A&X�$�s7"O�� ��$}N��G�mn E�q"O�[0�D��8"�F02�t��b"O��9��_�e��9�d$��X�$ݙ1"ONi��N@5L����E] 	:���"O0qis���+�
��ópж���"O
I#g��8/}�� ��t��*�"O��Y���&@v�[�#_�z,��"O�����'L.�THp���Ј�e"O<�"'�L�p��a�4��:�ΑR�"O� �\0@d�)@CJD#7��=H�@Ăf"O@�3�����l���B;�30"O��q���8���+���X*d�
�"Oz��!��Y�Z����[�\|�2"O�!1�(A�iH���W��=��X{�"O@L�a��:O�*���G���.!�"ODAs�fJ�R��7��)��}�V"O�����I�ho��1�o���h�"OH�C"DӘ2y�!1@v�ȅY5"O
h8�
&�$ě�KΏ�>��"O�p�R !}��BK�*�@<�f"O�8�t���Kĭ�S@˓p|�P��"O�0Ó)�%����a.��#o "O�He��h���3EM�{ZbL"O649�c��3#���� sI�m9�"O�d��`�'!�ʨ�f���_1x4��"OV$��lF6fH�|h�")!�"O�q�����?d�hYdW4� "O,%�v��*z�zlrCc�,ZƜ�"O��Y dT�M���b�D��"Ox��*�cJJ��䀅)�x�p�*O8���ʗ��ȗ�*o�i
�'�T�-�l�t$j��?kz:
�'�N<CՉT`�L�"'̍8a9�y�,{�>����٨Z��qr��D��y�lc�t{b\�H�r�È��yR탵t¤9�@Qqa��pA�y2E!��`����iƎls@�̚�yb��7r۰� ��$[[nl) �u��ȓRO���P$W�n`�%�#͒�;7Z4��f�F��L ~5p��oO 
D�4�ȓN:v�R�k�3ʺ�325}$��ȓOO�yh0�� ��ō. VRp�ȓr+^8Q"�n,�A�[1	K.-��t�R��ங����TrU��0s�໡bP�����n�t
*i�ȓP�<`ꂧ c��C ErM�4�ȓ	M:i���ɚ�!F��,� ��ȓ>P���An��2����uʐ?PF����4�+w��������P n��A�ȓb�d����J��j�)���0��=��Tc���F�8XΖ0�5D�*#�d@��� ��%��0#�NY)����6�����J���� �H�*X�8��B���ՇȓE���
7aзl}`��v!,Їȓ@D���W�Vi�<�EΒ
�D��3�M�Uȟ7Jxs�(F�	����.�������a�v�CэJ;������D~Çt�ةR�dJ>�P�z�)T�yRϋo\�c�A�?�=�V�I�y�l�8�(U�f�P�#���V�6�y���)f+�(�5D�/#���2�A��y�-��(�H\�smO��L̳�K��y2 00��ˋ�u.8�š�)�y�c�0V�@t��U���ˁ��y�"Z!W{PX�0O�F�Q"H���y�	ϣd��g�O����Q�����y2�ʔ_�,�[��ݥe��RP�E��y2�ǰZ>d9�̴N�Z9`Eϣ�y⍇��"�i��ڞL>>� "lD�yBb�{G���)�?-	Z�yA ���yK֒\��@Gń�^d[QhD��y�h˻L�"����*=Q�0�N��y�� $Q��M/�.�I�����y
� ���� ��$�ŋ��2�����"O�9��@Q<��5S��J�i��"Ol�z���,���Ђ�Z�4��3 "OXC�^�]���n��І���"O����%�.�WÁ/�X$���'��$q�G�[t&4�v�	Sn���A=D��P�i	�84�r1#� G�L���<D��AGh�)��Py�/A�vR��z@/D��!�+OE��r��12�R�rm1D����'ӨuK�L@d���X���h0D� �p�^j��!�]�{.�e/.D�T�A'ǥ]�|!�%��j�7�-D�p�f  ����J'��0�6D��	�IY���4��f��{��tK�!5D��Ť0unf抩O)�Y1�6D����̶[�d��U�V��|m�b�3D�D����v Kq�_9'�N����/D��*�f1p��ҏ-,n��QG/D�pKV���G������L�:)L,�֮+D�x�d,�`<��JU��'�p�$�,D�\�T���:���@��1/�A��(D�4��!�9/PaK�!j�mp �'D���c�4Q��M�eC�l� �$D����<G픥�c�M�"����6D��ҕǇ\0�x#�o�CYxu8�,3D��c��ńP@�4"׬L!&�Hu�$�.D� K��.m�~�CU�2ve媶O D�� u _�=lh���ʋ���D�=D����N�|3%���F���8��<D�� g	H�?y�q�� �bi�%��5D�L�B��>u�1O��,b5�#M2D���k�"TٮD����@eD�@֏#D�)E垕6�=IV��c��*6� D���u�ފmA@ #��^��h�"h:D�T�`��F�Mk�j���|�f�=D��'&ߐyQ
��U��$Ttܔ <D���oC<T��D��K�;P�� ��8D�(�	$BI�D�D,�s�ܠ�a8D�<�Ǭ�_l���ɘ1x��4D��#��,;**L`A*%bP��2D����T�,���r��Go*��0D�l�P���u.��xԥ�}��Q���9D��$�Q.,X@c�!$���
u+;D� ���vA*��匀U	�����4D��)�bT;��ف��Ы	,��8��0D��ȕk �b�J`�Ϧ��i"�*D���!MΘY����J��u��2��5D�\�7���F��ŋ��2��\�uN(D�D��_"=&,tj0J�?e��|���$�O(�y^��+���<\�`���,߄V����{��sw�ӹ�� �����ȓ�b�I" �Z3^|�� 4����nJNP�V!�qC����%��,������x��ϡ.T�3�|C<t�ȓ#�P6G_0�hw���z�Ή�ȓWT$9�7 �`��������X�����Pyb?O2�iE�N�eܤ`���H�q����|��)�S��B��c��&(`�!�
�vRB��,z�JT�H�	��́1�,|.B�P~�0��m��a��Y`0AA�8�B��)Vry��R�=`XYa_�GD������x�Оf*������l�!"O�@x��˼h=��j"��k���Cs�'R��'��	mD����	���;��8(��hG{J?� �ԩ�%ӌZ{��kѵ�X]�"OxЊ��o�4���+zʾ���"O���FZ:}@��s!�36��(��"O(�q!�!L�LA�A��h�PI��"OR�*���V�� 2!�S��`c�"OъF��D�$�#�4t�9K�"O.`I�']%4x����|� L��'=0����C��L�i�
R�M��'��%��*�$�0ه��L���:�'��ѭL3%r`p'�ц7���
�'�x`b�Ù�Hl$@w(�~�i�'+b�P£En����B4q�x��	�'�FM�g�ɝh� i��ƕ7��a�"O�űAm���2ck@�s�$�r"O��J[�����	c�|I��z?�'�ў��<�k)%D����.Yb$�I�c]J�<��dLn���S�"3B
e	qÓ|�<q�K�1>H��7#�/����p%�s�<�t)��E��A��݃+��h	D�s�<�?;��(��P����D�Xx�Dx�CW=}���r&��/_a \�0�1��;�S�O�0�窝�	�>9Eo �~۔���'� �C��K0��)≂�(DP	�'��Y�E��,��	@�ϕ;��Q(	�'F2ŀ��@O�~a{�*�)7'����'��D:�a��jIp�,^�.y*T`�'�8={Ae� �������$��� ��O�P��J6$bųcj��Hc򜑤"Ođ�J#Y?f]��"I
^�M���$�O^�}�WV�D��� uwpQ���l�0��B,t�2�
a����ҍ\�H�ȓ��A�������@	G.,u�ȓo� 4;���.��e ʜsg!��
��薉a�t�7%Į1VĆ�H̓G�p8[�8]+���(۩F� E&��E{r�dГ*S<� Z)^ũ!�	c�!�S< V��QD]� �J � s!��Z��ء�H뤅���hm!򄀝du<��6<�V��&�>kd!��>k�h����;<�i��\�kc!�$L�4bLO��
�\|W�1y!�$�hL����h�#Y�Е�bހI���`��ğ���O�b�� -b*��R.��9A"O��頫�NŦ�:�*ȋ7ల�"O�����N-M��4`� ~H���"Of�Q�J�.Ը���.���,�"O�X�Ul�$�`�F�ߡ^��[�"Od���Li&v��LV�Ss��!"O�l���X�o�Q�ËWYd�H "O�{����I��@�oCbD{U"O�y$i،mE�$�ֆM+���	�'6�����!~�����Z��r3�'��<[����~*�+(�/yr0��'v�Ȃ�M4w@�8���s�F�s�'�
�Ai��$����!���)��aS2Y���	6����/TA���Sc��z��B�I*�^���{��U$Y�����O\��B͖lN�C��׶)J9R��&D��ID&$4HL\C7�2{�@�h#D�l�#�A�W:	��.0|HE
f#D��_�B|�H�ĖAmbQ��!D��HED�H��̒F��<.���C?D����gʩtXf hTʏ/>>2E�S��<1����(��
�i�2ҴeQt�3/���3"O� �(f�ۃ��YK�@��q�"O�a �E�=�B���_>0lb�[�"O���@�M��J��A�ȡQ�X�[�"O4@��a��Vg����\#!�|�s"O.ͻ�ꄵp�h!�+��#�% 6"O�<�7(�
>Cah7��%)S����^�|E{��;f�cf�z�z$^�!��
+��!�`��nf����F5�!�d�,1^�gi޺8o�1j4O^;Y�!�Ę2��,c�J�M�
�P�H�6�!�D�(T�h�䊄&�<4��'[�@�!�䍇m��P���{�XypG� ��'ў�>�˵�c����
�J���
���O�=E�A��аi�@��UX����!�D�:��`��(r���
�4.B!�d�G�Zq��䂈;/����	�!2!��vj�(v�ѪHX0s����.!�d�/.�U��ȉ-4l���j	�F?!��


K���լ�8�$�Jg���==!�$���y	c!�$	�l=c&���U!�ę/ٺ�1�� �R� 2�ۄO<!��[�BUI�M�g��X� N�!�$[�7����荼YUv[�$i�!��Ѯp��{�O��(��'MP�>!!���k
�Y� �߆ӈI�N.!�V7���Iঘ�h�\1�kRv!��q֔d��L\�hľ��%*�-H!�Dn����QAϜ:�|	�G�r�!�Jh�F�R� �<�@P���;,!�ΝI`��92J�����	Tϙ+l�!��=#|�k��ɑ*���	3Y�!�䆺"cz09P��-!��PU��*8!�䈷2��cԅ�z�5��,i*�'a|�c�n}�(�)��]��r�mײ�y2�X9@�8\�cW'׎�X���yb�Z=�Y#�
�ڤ��Q�Ѥ�yrG�pX��v�K�V�ٹ!�T�yR �,�d�*௓$QY�� �#��y�%@11�TX�ToV'X���8`���yr�c�x�#r�!�J�b'���D+�O��6mךhO\���e/`�	v^�p�?	�������uD�DDf���՗6N���"OF� SDE
K�J�re�E5��"V"O�@��S�	�(�H�d��E(��"O��6��7<> ]��I��-h��"OT-
�Z5dD �񩒇7�@A�V"O��q(%{7 Ԩ�Yh�.���"O�5�b/��W�Q
�	ވ�H����|��|��'>�q#l풉Aì�>6�=A.)D�$k$#���ƌ4����@�#D����/��|���1$×>�fX��`7D� c�Me\1�qg: ^L;�:D�<��V���{��P�B�3D�P���?(��KZ�A4�Ԩ�j$D��#�f��t���ْ��4(h�*'@.������I/ Ǡ�����	v�
�'��u��웚-%f����1�25#�'
ʄ	��#�*��枭l�$�2�'{t����g�\�Cf�zS��#$"OvЂ3��#F��(��J�(�H�3"Ol˒��)[HY��
"t�(A(D"O�a��.Խih��0�ށ��U"O iSe" %�h�V���4$�%"O%K�n��\�n�3��W�+���!"O� t��SƽS���:6�>c����"O��X@L�G����M�[��a�"O��P���,H� �V�NHYG"OR|y�Ҏhx�� 7�K�Rz�I"OЄ�S����pq�
�
���1����� E����CA���`R5d �����y���}R�@�c�.|��X�9�yrNѥ4h�ʑ<V��1�ב�y�H��8��!�
5+�d	&+Ҧ�y�MQ5i�D�it��	}N�H`�C��yD�!Fm�|���m�>���e���y&�e�x(���k���c����<���_�K��z��L8!�8t�	Ø"U!�A�#�̹�O�Fb4R�1O!�$��ѓ�Z�H6�]0�|C!�ԄeP�%p�b߃9���[t+�>!�V�J_���WǑ%ߎ��D��7!��ѐDr��O�U�Xx��(�6!�D�{dtD���&�d Q��ՓJ,!�dC����㊂[thb��!���ioܭ{1&S>u>��"��< !�ę�Bm���^�5y��Cm!򄑊�(���� �Er �S�_U!�^
 O�}���ʪ{[�h����DT!�D�#%�ͺG�nekP���!��#A�@�V�UÒ�ӊQ�ў����/l5����ͫ8�\p�̞�Z��B�ɱ���VB<v�D����	�C�	���)YŤ�������'!1�B�	�o��p5"��@bT�!aiۨ��B�	�1~��@$�W�II h ��׬eZ�C�Ʉ|[��A�"_8����BYպB�;��z� �}��y�`��3)�B�	: t�hk�k��d�$�ՅKcZB�I�Fh9�PF�
}�<I�tj�y�NB�	�$ a ��@/*m %	��PC)BB�ɽR�t��4'{]-��$�o�$B��#b�, є"�
vX�!���VR�C��zK�UZ4�8��|ieE&w_�C��:2�,�#�>e�xHcMļB��*}�H�x���-�ՙ1-V��C�ɕx`���5�Z�܀s��.g��C�I������M)S(��B�K�z�C��1<�.H�fJ�o��y!�J�.j�B䉙71�������r=�զS!��B�ɯl\���eBI�FиTbR���B��
�8P��V5u���a��',;HC䉶=�*`;U���?"��p��>RW�B�	�)q�(wJVY��S�;��B�	�jE�X#�A����hPa�R2&jPB�ɼz`�MH�$�,ߚe*�"�2&fB�ɐ^�f5)�oƃX�X	�,��M��C䉲t�p�U 
26�n�2@J�{��Oj����" �M8%K�d���	��G�ўć�S�>��p���!��8�#�	`4�C䉚.�����. ��Ȧ)B�o��B�58�m�#�j���8QlR'	�B�IG�.):,�0A7Ψ�e�2|a�B�	?z�p}���e� ��M
�FC䉔��@9@�
	���b�D >'3:�d:��0LO
�*�d-�I)saP�C�D���*O�A�v���)P*���@Y4U�Z���'t�V\�[�z���e^�<H��'��D��� �\�4YR��� �U
 H�Q9�UA�^~��R4"O�����"^8�(D�Ӧ��R�"O������"#�z��:A�.I8"�'.��'��Eh$�N?G�6y���f�tU�	�',^�	A�$x:QR��+bFM��'��ݱ�!Y.m7xus6b�+R�ְ��'@Tt�Vt^�����PP���'8K� ��k��p� ȴ
����'[L��ホR�f��ĭs5��'j�y��TU��z$eA�jm���'���G�L|RX��s�E9��0��'?�d
��_X{��cG�p�B��	�'4�!q� �40 h����~li�	�'�,`02��2s0ѹ����P	�	�'j�L���`�\d@�m�
�j	�'���-8;Ѡ� �Nǹw����	�'�P��� ��, �G���p�'%��0c�ա`���aC����	�'����!��As�ݩq�������'ÌI�@L��r:��*HX�'���Q��/;�R���鑦"{,��'�.���l�:=�Rq�ܢ ����'$T�2Un�UɆ����T �>]��'kXAy��
LD��I�4�x�'l��i�8C��]�ToV��9�
�'��pPV�V,�������"A4���'�PԨ�� �iE`媳ᛈzx���'�� ��MK�j�����*�.K�d;	�' H+��[�>�i���b�t���'E����]��\*�c�"qX����'�JiAe�f�$q7LZ�ev����'Ȗt���Q�X�f(�T�Z���H�'���ʕB�7M�>H0�N�f���
�'$��@[�{(z��ۣ0w��c�'C�� �J-i����L܌R\ƙ8�'�0ɘP�:A�zT!AEB�M5��'S� ���%_�:0�p�#>u*��'��y�:l]4�G`C,H�@��'�"�:�S�~uBD����<�4��
�'J�z�E�oa����6F ���'0xxA����*�dlՄ?-�8u��'�,	@C��=�qow�:pv�<�� �1򘝐�
E�kH��k�@�M�<�c��e%��	�k�a�ԡ�ǥ�I�<�fg��N	�u��;bz���Ǎ�m�<�E$ňf������L;Yz��jRj�<yg��'<��Y��X8�r�Bf,g�<��I�R�2�3d�:Q��Ӊ�n�< �\-\P��b��9B��A��$�y�"�81;*����q��ؑ��e�<)��ɚ���"/͠,f�+�a	B�<��%ɱw/������%C@��Bh�z�<A��O���B�/ٕU�� !P��N�<a#�ͭwN�bg�Ԑ)��`"$�N�<q���(-s l6`�
>�(��ĚD�<��Ι9��qAU�VRZF�C�<!��?clNh�4KH�:�m���YY�<�6x}�I0�\K@�@U�<���^�j�;s.Đ6��Yr2��j�<�U*1º}��e�I�=R���a�<��R=ՂS���"B�r�	��H_�<�� ��W� ����	�fVD�1��]�<��E��4I��$B������[�<��V�N4����ٗQ��A�GC�[�<� 1�kö8:��hG/W��ӆ"OZ8�Vf��8oF�����B��Qg"O��ض��|�.E��<U��+�"O-���	��D�B�
S>E �"O�,�F)�)f��4a̛FQ̼z�"O>Y��)����q%�Q0z5�!'"O4��	�^���(�C�4j�Kv"O~U'�U�\8,�0�b�8%�Lz"Oj٪��ZҨ�a�!�l=�W"O������m�C��*���"O8��7K�5pգ\<t ��@��y��|�N\�@Q�i�|q����y��	�"(d=���Q�f������y�ψ(�H�S�E�W���F��y�#[1)LY�@i<M�\H�u���y��%����C(D�pU혿�y������ ��h:|
�� :�y�o�0i5(�"DG�cf �Dlŷ�y�+�(r�8\���2V_"��SM
�y�*�,�Ъ3Y��M��-�y�
	F@����ּNhp҃Ģ�y2�Q
l<^IiF���D2*�3F�y��ˊMlP��t�D\� J���y�
����x�f����S���yF !
���N�b��b"�ߋ�y�(ɑ.ݦq�b�ۦ�1B�O�y�
̰>
���1hX�\S�#�ybj	��k$,�Y��3�y�F(q(���=�J$P�LN6�y�#I�+W  �fЮ<4B�����y�KM 2B��S�a�Hؗ���y"IL
`0�q# �`:��i�g��y"$<Zu�E���X���Wƅ��y�<P�LA;O@	W��Ű"���yLd�u�!I�fnb�ڡ�I��y�N�&�n�)�h���j���y�g0{�)���4����T�1�y�$[��������x֨%�c�Ũ�y��&����Ώ�x��Х�(�y��%ڨ�ʖ�Ҟk&�� ����yrƏ�(�(TT+��^=�Y���$�yFʌ'm�%�7̩l���`���y"n�:ê�C����b�\�a�'�yb�T�c�\�E��F���mП�ybM��	�����
]�y
�eV5�y"�W[�,`bD�L� ����1/C��yb�ƢF.@�����p����AŃ�y"�L�0U�6�ʱr�^��p�[�y���;�*���NI�j�PH�o���y¬�����e+<�S�j���y҄��k9���EԞrk�%"$P��y�σ�r �6.������1kԣ�yR�%��	�U��@���y"B��H!F�W�<�0���y�,b���S:�(��@�ۆ�y2M��)D�åR7/F�!�LN�y-��m�h�p� ��xD#q�M�y�	Wu\�b�)x���@,�y�I�xR����m>�=�Q���y�#I3z���kO'a���
O��yB�У,O4}Å��T��䒓i�*�y2�_-X��k�Rs$�Ht��y�&��s��h�d�=ISvt�ù�y���<2���q׾H��X�)ʺ�y
� �Ds�3Z�fM�Dh[Y*���"O|�8��/�� �FfK_���ɦ"Ov�x�G� Q5<��pe�0��6*1D���!D8�������� ��.D�!�B�$&Ƥ��eJ*N��|#7�7D��A!�J�<j��
$����`�g*OXH��<h�mt�E�z󚙹�"OdՒ# �b�,<1�3��d{�"O�g�	%T�0���Ė��@"O�x����6�$
�焰S��y`P"O¬���	^���֨;M�
��"O�ɳWB�9�~��;C֖��v"O� ��.����#'a�@_��2�"O�#E���j2b���@��*T�PG"O`͓�h�D|lKa���N�y�"O�h�"����=)M��<��Q��"O�l��ٽ%d�{KE�k��:�y�K;X�1�U�G�����y�U�G0��=MlL�5�;�y I�=Z��f�A(.��i���F��y�HP�zA!$;�uB���yRX$�ԡ:$H)�d��Ñ�y�	?��p%�q��a���y"��-,�h���"�>o��y��a�yb�ݗ���˔f�.14	x!Һ�yR�S$6���0୍.Z:U��ȁ�y�ÿL���`�E+i^�k��G��y�#�)Pb>����צ��*�+�y�f�xk���D�*:<Ÿ�)��y2���	=��IuLԧivz��2-���y�L_�
�TEe&0�f��A�O��y�oJY���hW�"(���@ ��y���@�f�Y�h뀊D
�y�c޸�Jpa�(w\���� ��y���Bx���mg�#{PBlC�'��E8eB���y���N�n2��
�'(��4g�>������{���9�'�2\ q
Ӈ}��U�5J��yqT�x�'=ў"~JB���K��`$�\'X��#�"�l�<��@9<Ƹ1�aID)l!R��5b[���D+�O�-s���A�,�)G��)<��Ğ�<��	/x� A�$�N�o<tk�C]�y����D�<y��O�~��03h����7ޣ�y��˩n�f�	D �y����F��&�Px�(�L�$'�@qZ���^��~եO*�=�zS�	x�!�c@�.�fU�� c8��Ez-�"^R���[ �1XD�Q9�y�H��<8ི�d�#N]�ruA����Β�~Ҝ|ʟ�R�x�b���>��S�V�������n�N�%�w��!cB�t�Q�u���>�G��4K���G�z�<�C��;$7č���V�g�1OOF�?�*�'Y 
���'cj]`n�i�OR(Fz���mZ�%���y4dB�6i:a@���d4���t�D[��`qyF	!~���ԍA�!�=Y�~�,�H�
J�?�P��-Ov�/�i>	�<aC�� a�T=��x��
�q�<	1S�@�r��P�D0q�IX�hFy2-V"57����I���ί�yBLϨ|욦�<��9pTD�y�ǜ�M����I�H���B��N�y2`��~�P��9WOKQ�2��P�!B���c"\�т� 0�j��ȓh��I�/ɜ�Pً3�Y����UB\0��E�ML>	����l����S�? �d{`M��}�h�ȶ�T%^C�,j�"O�)AvJ�2YbB�`�E�����"ODkGl
��>��2" �bm�@P$"O���%N�/Z� �@�^dҭ�"O����@�	J@ޑ@UȒ��x��)�S�V�D�S&�H"�Pi�Ʋ,ȆC�ɢ=\���%�X,3�ha���yrc�t���-5D����ߠX+���5l�-�2C�>-�8h�E �"���r�H]�._��'vў�?��ۆK��Xk!�ɲ]&���j?D���4dێo4����z��囁�>D��� i�.�T��6��� ���"�)D��`Ɯ�:;�\b�*���m@�E$D�Xh�l�4]�`�p��`��'D�x
PFL�t �1Sc�2���bC�+D���n�^�.ŲpF����")D���@�LD�<z��G��#f4D��3$A3��\"�+@�YI�(Ö&D��ХW�\p�֠�f�����j"D� ����h�\m��a�b���I!,O��<q��O6I��h6�$��t�Q�v�<i����&�f��3�]*oI ����n�'�qO �'d.�4�@Jܹ�d-�6I� �4]��E�>X�AK�Ƥ�EL�G�2�ȓK�a�D�4<�� �CHPێ���iW�,�S��)8�ZQ�C�6]T`�Γ�hO?� �[l�qZ%_/q0����/�O�2� �K����jH] �,�Aᘡ�ȓ%\جS��loN���K������XQ*�-3V�0�S��Aڊ	�ȓ:����2g	�\�F'�c����'�ў"}J�F�-q!�u���x,"$���]e�<ia'F�v�K��0kVM�G�Qk��"�Q�t9�y���@��q�b� �Ѳ��ߒ�x2�'#����Ή
���s�@՚0�f����'M �x'�H$ ֐���@�36 �)�'{�Q�T<^�� 2F��5������6}��)�=�FAj�G͍\Sh1��ʼj_RC�	|��D؇ʉ0f�&O^7�C�I%� a���$�`���Z�h�̣?�D�����!"�ܸ7B�Q�e��(��a�O4��l�(�x-�bB��o�mzvC�N�<�u�&V�1uDP�Gp��{�K�J�<�La���:��,N�>����S_?��g=�S�O4	(2k�%5�9�4�[7y���[�'��9�E�	$�p�FG�8u�M�J<	7�'�����*ݸn���25�G�#(�<�L>��O�#}��O'���t�E3�f��%K��R�'R�\P�l�J���ݖ'5�90�r�'wP�aRnӣK.���l������'��PJ�/���I��ќ	]�$��'����Ux@H	D���,>̹�u�)�S��?��D���L�����3�l�5�T�<�wN��� �^�CnVqhcAڦMne�'�Q��P���	 Y���ԫ;�>���@+D��Z�B>V����Eϝ�d� F�<���<�����[U�|�t�ޗ{̀L��� �Q�!��
=9O�y�e�I�t���ri��o&H6�'�S��yߢD}�1fM�A�F�P$@׌�y2�U�QY�M�@�,eJ��0�y���/o�!�앦Yqx�������0?�.O�!�Aj�Kնy��)R��6�3�"O�U�j�W����(��lܪd"O��P
�lcb4it�����"O� pu���%%T�� HI����O6�=E����Ψ� B��>)$�� �L��yra�=_-���S��#�N�(E:��6����a2[�c��c��;0MۨF_!���Ħ)(ȋ	O��@UA��T�V�x��?D����8Dj�9  дY�<�Ȇ�=D��JS��s����ժ�$K��8�'D�\ڤ˕�C�
�K�O�+�4�� %D�����$Q�@a���
�H��<��%!�X�ΕE��D�
	��;K�+#`&�8�����'Fl���C�puc���];�(զR�'�D]"ef�>O�<���'����i�>H������(��ʆ#3��9��'�$�2A%_��I#��E�0ך���O�U�L>�rg@��u7��^�XT��|�@9�3�&�p?9�O��Z�"��mi�.��@�a0Ƒ��G{���&����r��qCP�+%�4!��;ЖT���R:|��0b"F�z��'\����ɴ8(�(Cŕ.i����'2�=�çHL��'�C���d���m(����aPNL#�c��\�X��ˆ_�\M��e������c��$Z$�Ĩŝ>��M�$�,�O���On�Ӥ ��YA0܉��#ކl0�"O|�Xf�4&���� �$&�	���'�ў�ڐAӼ3�x�kck����L���!D��'�ǲ@���!�@���i� >��2�SܧP�|�T�֨L����&�	�$k�i�ȓX���`���U����mO�9B��oZH̓�0=��̸+�­�4��6���Opx��Gxb"�?8@�*��g�ҵ�݂�y�	�'b,�
�F��W;�,�GB��p>	K<qw�ԖH��\�u	�-3�H�
T%�d�<��������PENS?-u��pO@�<���S��Y��M:�4�e��g,jC�6�l�6��.<���K4E��t���Zz��4A��f[�,s��ҚjH���v��[���;lg��g%��	`B ��cl� �J��x��$2&��8�0 ������H�	���0��b�PCҁ��-<�C�ɥkf�CW��&ø�C���6P�bOf7�,�S�')��= U-�g�mY���2{V��Po��p�m�
^Iҩ[cD2�� �ȓqF�����@Y�n�(-1���ȓH#�|3Մ�sr�D�7��#k�8݇ȓH��B��:�(� �^°��V�kg$�2��p���_j�ՄȓQF���!�m�R@C���nyJ9�ȓ :3Å�k�a0ժR�5C��ȓ7¦�Z��$��=`�Q�2�M��O��b�IR����X�a��?`}Ys��dh�Y�/\�p�ȓR	���cǾuDTKS�_��ȓkkl�2$�-�cV�T�d#z�ȓZ�h`�P�K�4�p�
 H�0��;ֲ�"SFI<��[v)�+�B�Ir�XQ�� ق�A�T&��C�I�������TlH��J�C��!4*��)� =v0�Pge�&�fC��,>�$"�ŕ7MV���"	6l��C�	0%]Ph贀ש:&��d��6s�C�	*;9�]��Ѵu��Q��/ռ �C�Ɉ/��@�Jh`r�q�ޏ?��B��)�"���Α� -�(;1JQ�B�	�XQ�a�!B�P�3@\lg�B��--S�A8��=a��T��ǟ�/�B�)� ��r�R�/%�U��c�R��)pQ"O�h+��L���#��:Ш!��"Oq1�L�PT R�a03�����"Ot��#�P�&��)�B�Y�e|R���"O~���f^�U� �K�j��
IҠ�g"O�(�(�ap�J-TH�!�!"O6� SlٸM)����'�@h���"O�#hS0Qj\�����Z���U"O�(cA��S5���%j�֮}p��b#��JG>x�Z���"6a"�	:0*��j]�f�>r ��K�B䉔Arė4tN�(�j��1�� ��"O,�����J�	nz�P��"O>��p*�	}�Zx�v��(9u��"O
�QcC�'45A��(���2"O�u@ꔜ2�T�$�]�f}d��B"O�Eb�`�"Uv
�m�1ʤ��"O����@ Gޕ@"���3ʸi87"ON�[t�[��4Z��Vb��ѓ"O\���a�wBx���	���"O� �C��E$�b"�D A�<���"Or݊�)��}?n5R��
�0�V�c"O<�Y%�q����-i��!p�"O̩�� QRn��eZ+(���r�"O���qJG�j�tQ�1�)�JX�"O�u��.СK�KҠ+z*A D"Ob`y��J5Ө�K��;���b�"Ob���\3�X):q �.0p4�)�"OV�9��(yVѓ���<s�$h�"O��p'��������ʇvh���F"O�TR��B�!��� U����"Ox����fM����&L6gc� "O�T��Ę?%��S�Z��x��"O��!o� a�ݠs��5^҆:t"O��*���4�ȥ��W�v�R "O�p�B�� Pgl��-�/i�M[v"On��lת\l��g-�%^��1&"O������W���フ�1�V5"OT4�����;A��h��ܦ@��Yʡ"Oʰ�f,�tT�J��B%,��`"Ob����נ{ˈ��F�_�i����""O�4�Ȟ9�^��@lW31�D�r�"O�0��4?����q���>l�,�c"O.EJ�i�%�B�;��sK0�t"O��Y���-P=i�$H�R4m&"O�}��	�'^�ء�NL��@�"OH��b�X���-�g�� $�S��'�!`ebP6�&J�2������+O�UL<��E���p=��M7S�Zq��J�f�	��Mv�'آi{�mT�W�k�Q����'x���{���'1�hԂ�׋�HC�	A�RSe.E�u�@�y���w�n7��
c�¹P�.����$���@�S��\c�����`�<^���(N�lM��'G�x83!��.x1a�E�A�����'�NH��+��  ^
�Oҁ����'���:�)K"!.8���a����O�0+�k�_�(�v�-m�L���)��T	@���2?��������])���)��h\�� P��hOZB�J$'wđ��O�� �NԊNA*p���P|�8m��l��{��E1�',�v%֏-4]V�E=wĤ��4b۠�qG!(ŮO�M�����:��{�2TS���(8�~AB@"Ofhf�\hx�Q򨐢"���_��h��@� 	���'�q�G�B�V����#���Щ�
 ������� @f�7y�f�h��W��@��;4���@�,2��p,<����d�=7�z#=����% Pp��w�#����>$�o�=mhj��U)H��2C�	" �r�I�Y�bK5����P7́�S�2�!A����)��� �w���?߲��CH�v>4	�`"O�82�����ۣ(��1j�P�_���c��#Z�@��I�n\��ssތY3`5������s��Tx���&��k�nȼ^ r��㧗%�!�֌H`*�XE��K������[�W�!�$�5n�X������?d�"��b
!�D��=G�
5~�`z��uS!��^�b�
�#���K�ب�� �{\!�dߠL�̔�P�H�g�j�ŏ_�t�!��<2;�<@�ߤn���GnL�qH!�D�*�u�A`��e~�u��5f!�� �*��f]#$XpC�?*�!���i��|���M?� ez�

�D����B��(��I�o�Z����w�ޕ�"�-.�$B�	�:֌0�r�ũdf�H6B+E׊�C��*tX�Zv�'"� ����Ά�k��$JDF��
Ǔ�f4v/E�A�.	��k���_9!W��W �X"O)D� �˛o����盋*��1Cd��3R��	,]|����/_�FE~lZ��O:�.�z&`H!�Z�BJ�Rᘕ*�"OP��CcH��$Y�J_�&��	�ş:6�H  ?O�H�M]�#��n" ̛��)�)8|A���Z�B�r��>�(O���iW����,b*T%�Xwa4�5��tӸ�d�� �P��b����7,�6j��c@�-�a{"��=,�Z��vl�H���R(��!s���m��dGn�[wZ��ؼL�0�wEЙG��1v~: ��ӥ.9��r6�r8�ȓε�q�E��l+�4c��иq��:�P�;aAJ�7x�mk����¥��>�x;7����;F㲅xR��F|:uY���y*"��ɗW=P��"�D�f*S�4��c%�F�����*�qa�?:�1H�ɔ�mU��XwgH|8�`os➬��C�\Ʊ@��D�GF�l��O%��o��8ѣ�`���D�EB���/h ���B39e�Xa��� �j9�����8��F��3���!��S��x	���'ĭX3�U-"j��h�C tA���������[PkS�
�B��'J�3NL�sO�����;�h�/^���u�R�U#Ҩ�"O�XB�(E�W�� �G�:n���'�X�!k\�sJ���J,g�xz�ER��!P��z�1~�x#�L�#?�xi��5����O�C4:��`0�M���yLm����f��y��U2/W���� ��)*��A�n��yzH'>1�=ա
�bI��.���4H���a�K?J�ztJúbc>�24
ú:�����d�Lx�k%p�\u�ӀR�<��Ѣ�&J5�U�뉘�LX���:t}�h�c�'�����E�n%N�'�L��j�H�`�(>�����0k,׋,*�{2m�*U�DT���A!�$�+XJ)J@�M�F�)�'kg;9T#��ZD�Px�f�[��*ZD1r0AͯG�1�V�Q��ܷ`AL!;׀��9���'�'^��1tU�9R�X�hP�0R	K({ڲd�%ˎ ����F��������[��b>c���v�O2I(�i�%��X �/�Oz�ZCI��?��Q�cb�7��l3�I6S2vUY#�=@"4P������m#5�'�",r���f#�=+�a��?�d������~Qx�$[�7�@D[*�1x��09�z��a�� ]�착2H���5"O�����ƽk����
80�����"K�
�b���M�<���#H�?,��G��2���w��]�\�G)`x���q"O깸e'��}�{�
�c���)���[u
�(qGιS�X%��R��D�I�0R�x)R�W���P_ i���$Q
��5�0���Mc�OO�aU��p�j[e�PS&�|�<i�CM;H�� ,0�J���}������'ds�"}�$Np䐴�%k���3�Ig�<�U�J���p�r�Z��τ]b��P���|*铈h���H$*h�# "�'h �$�59!�$A��%	��H}$��O�4 <�P��%�5���RПD�A�O�=I��� ���Qe��k�y�CN��%��{�f�6<�j�j�TϦ�QgĽ=�� �flK4c�ܹ��Eܟw�N���jò��27�"iuF�_0��$ƙ���<#�\�fjjA��u�vܡGM1F���q�:����̠9�tH��
Ǎ~ĪC��5}���,M�&�PᗙG��0��ھI�|�+A8Ov�!�Afv�ų�����!�J Z��	�P�Y�.Ġ
"O^Be��T`�o���v��5ԢQ��i�q���8q%�g~O�vL�<��	$A".� c` 2�yb�	:Т�억;�*h�5��QT���m?$�`M��S�? ���5jE�����Vg��`9�%��':��!@���iL��I�j^�m�@��\q�b�B����C�I	�a�Ci�"I�$���ŋK�c��`���E&0"ڠ�ٗp�BD��@��H�l��va�g�<Q�� �`�R��1��� ���.E`�<A�U'u�j����_VD	c�OK�'�Х��S�sfzQE�?��*��J��\�eH�In�,h�!D�����%rF�h��h��uyǩ�>��U�Hk��:L�j����9�V�[p"CA�
��́b�<��h�O�hl�2D��B��Sf܆x����'�D0�pʔ?>`�q���O�u"QJE�b��(��cٻ h=#��'̀ipw��+r߶q�#8���hV��`�m�-z(���'N������H�ãg�{�����J=I��Qo=:v���go�~�"�9Y���sf�M,0h��Ed�<�+��\��񱢆��ࠁ�gMg?�%m3�L�8���=m�6mˍ��[ 2Ѽ�9�+%X ��j0q+!�dӵc1022�ؒhu��q篏##�.mkf#�#"�%�&Gq��$b�ߟ#=A�-�4|�\Tˠ�J�:ZR�;�t����b��Z���'�]�F��E�A>�q(GG�X2�a�u/E�.D\D�>R���f�R��$�ӂ�R(W<f�?�*G-{�$y�-$E%�QX��$R�z������ �&����8"��܇ȓdw�)�a�5BA2�y��۴Ha��j�M�fAD�ӛeo�Y�DƜ,�H�`�#9��ҩK��H�%
�*P�,B��!}����@/�
]�*n���B!|��ை	[׺����ъ.�.�	?�h�uxf`��J�#Q����-|Oʅ��L�1��T��4fr1����o����P�*��8��e�~�[6h
)
�`ȡ�3N�\��?q���~�$�p�,0�'%��rрL�=i�E,���ȓ{Y�|��ȏ�`lF<��ʚ4dL��ENI��(�>����O�j���%��K�D�:+Pۇ"Oz�!�Ύ#7eL�u��YL`��'��,B#��Z�L��I6A����1�N�:�x�I���.l���ןWXȈaF7�MK��T,r\�S���*d_"�'�B�<񕀜RN8��HV�Nn>�b�v�xD�&���<��"}�Ë X���n� <��|��Qv�<Y�C�2 h$��d�c#�q�]79�����ML铵h��D�@&��RiNLVD9 ��T3#!�$�%�v��5�ɣEB�າ�
K*��׻[o�
T��n؞#tl�6v��{4OI;R�B���B#|O��un�	J 83�47��������O��xA	�Vy��ȓL�PقV�
xz�-¶�YIN��?Ai	<�Z��%�8ҧ�l�R#&��E��&	v锱�ȓAHH��"C�ЂpKr���D0O5�):L>E��'G�U�g��Rb�|QƞM�8�k�'v\HY���CͶq1c�Bàd��'��z���Y�L;r�ļ�xt���ވB|���6D����d
'���pJ9&Z�#��(D��D-U��.�cS�ʴ �\i�2�)D�Lၡ�"T&�3�g&N::��$`;D��ԯR
@#8���������B��;D��p���\��t��*�&�`��v�2D������)]�Q�� à�j\�A3D����&��8��o�-~�&� ��7D�d��d�-��]r��t����4D�|1�#�YJ��&��/2����6D���C�H�,��Q�NA5F�����&D�0Si�М��" ]�/���@A�&D� �Z�'�Q��ٮUԌc�g8D�8����#1�NH�cT-e�8��#D�$�	<ŪT@f��X�+� D����
_f�@���pˆ��w!D����a�1	��p�� N4����3D�!���&%�ȧaM���d�+D��I'�^t���!��1M��l)��:D�� ��p� 
W��S��';�m@�"O4�ڵI	��p�[�e��˅"O*�s��� �n�r�V.�$\;T"OL\jCĎPb��`)��-s"O$�d�Qf)(�҂[6���"O�ҁcɗg�����@�<��pj�"O~���Ea戋�ɕh`�R�"O�`�7
��(|2�X��w���"OJ`��,D8kS�L��Z��|p�"O�U��a�	R�1*���%n^N<8�"O�Iw�Og݄�QХ�u��4yg"O�y�LR�~\�j��p��C�"O�u��$��>�,<��d�7���11"O��3��$ݹe�/��À"O��ȁ��0�!A���xx���"O2ܩ�l�@����d�]yJ��u"O���Dɝ4v�����$��H{b��a"OB�b1b^6�j,�wb�,E��e*�"O�M�wk̻r�\,;p�B�g�F(�W"O^��f�ü2ha���i}���"O��iV�+Z_J�;�
�md�x�b"O�d 傎?4� �2#2B���"O��6j��~H"@�dh�n$�#"OXǎ�i t(��Θ�N��}r�"O�)�o�::h�z��;#��,��"O��"so�X��,��U�z$�"O��գ��j\R�'N��:�"O҉�C��3�4�� �#j�p\��"Oܥ���͙�%�Ld�t���])�y����a4��6S�,$�Sh@��yi?C�𹳲�T:c<��T�ƕ�y��V�fU�⭞�2AB� ��Z��yr��(��)*9^��6e�7�yrI�!
v)� �-x�t)�녙�y�� 	��:I
�j�=���ں�y҇]�-KSc�붸�0Q��0�y��iX�yT�]�f�z%��CS�Py�#� #���/Z-�]8��_M�<�b&ڧ�� �"�D�6:��ICO�<с��P�\ܐ��Y4e���4@Ml�<Ɂ�E�R�ȼ�榍�K�l$��n�<�rc:^v�;�'	O$<�F�P�<)�غ����K� u@���%�f�<i��]�3�$,� W�P�2�*Q#�c�<%b��s����4i�6`nHݘ�P\�<��MC�p1���N7 ��H��N�u�<QC�g �8�'hF,k��u��$�O�<i��ñp�搻� @(#�q�QJ�<5L��RHvĲ�/K)f
��af�F�<)P`�]�)I�g̩2��T:KJ���eŁ�F<@e�
Ъ8r�
�1x�e��#D����e��A�����ܜ}!3�?�~��a������DljGjl��k�ڜ\x�: "O&Dx%��6Th����<~eK�i�@e1�f�Z����O?7��JтR��U��<�R_�v�!�M�C��i�"NC5~�p9��ֺr��	s��3%kI(M��y�M\͸񐔌E�JΘ`B�	�7�>��Ɠi���Ы��$Z�}6@Z�a���2U�_-U�>B㉩u�Q:�C�-86e`1L�c�
#=�(T�<�0��q�6��xa@�H�ኬv*ő���!-��B�	�I
",C���1R�!�n��v�6fi0ep��+��)����.�.ޤ}���S�I���A".D�̓�l��&�A� ǒ�,��@Q�-�>���B?��L�7D*<O��qC x:ʰBd%No���u�'�
Sk�?E?d� ��H��]���ǌ*���3.?4��Ke�/�9�WL�B'���!ғA�Ғ�����?�I�H�$*�8�!挙�����+D�ԓV�C�ki�@p��аQL5�E�k�Hq �M�H|N�"~n�-d���K��F���3!�%�BB�	�sB<�#V�`�}�g��kǒ�X�������0=yC��r̪̉ ��#P�6 2%�H����vFDX@�Xf��)E���c:�c�ՑN=!򤈌?BP"�0C�> ���
�U!�d�3��(�E�/�6�p��{�B�ɊMW~6��5(���F��C�	�A��qq��R$���@�%~C�ɏ5���%!V�x����O�+ԬB�"*)����BѲ,�2��,V_"�B�ɚYB�t�!�b��I'�ȩQjB�	=w���:W�!��[4AI��B�I�� YP�bҬv��U�6� R�B��%)��T�s�O�Vh��g"�2_P�C�Io ��` ��4G44����:��C䉺gO�(����p���)d9
C��P�j=���{���H�M��B�	*pz����㜪`���3"	�%��B�ɐx��D@*S�*��ɋS��9l�B�
���ф� Y���뇫_(0C�	�'�p}���'a�0���<	����&#~�΍�Gg�EYAd�H�P%���@u�<�#Ӷm�" @�K�1Zn��vm�>|2:y�f�����S��y�#׀=V5��JV��t�#.�(�y�$	��t�EB�H�2�K%�?�-��B Td�4lO�[���9�2(&�^�F�d����'p�]*t
�?)��o�[��rg�Ŏ{�:������.�C�I�5Ȕ�9�ٻ$� �eN�3-�����D�zg�5�S��;��q2�]�cv �U`�N�vB��$�,�IQIQ�v�b�g�:8j�X�qO���yO�E��'��A1˄�2AcH1�l�h�'�
-2�B���x��,e�H����!v$L���<���T/<rb���B83��/<t�{B�27�Ղ#t�2K$�[:�8j���
V�,����,D�L�����p$��c����y�-$���#j���6��4��>9�Bhְ{����%��L�6�$D�h�!LK�*�Ψ;F+X�
i�\�F�6ƾ��2��z�)��<A�`�Q��U)ҭ��]�9D�BA�<Q��Ҏ �<\ru�jVD���IIv?�ġ�z�����S?Kr��K�-��qkPE�b�H�Rl!�ğ�W\�p�`�߫|"�bnֵW2!�䄈"�Y#f�����I��|�Q"ϓ'Jn��E%�2�����o��Q#R���{��p�1`�$B�LhB�@��$Fx(SF�<u�P��i�\�`Gأ+��=;QJ�x�C�?z��OH e�j�xQiы}��+�Gס��ZN��E��'GJe��,S�UT!�G) �8�����'���$�[�vh�4;݌�Z�MV�� a)�J7����Bx-� ���v�dd��Ðaj�{"�9v(<I�&�ݦ���J�t ���Iһ\���F-D�����	"U���1Oܖ����'?�I�}���K�	N�F��>�zR _:u>8�� �00�T���;D��;� ο��mAD/��'L���!�8P�̋PK����e��~2��"\hh�ԬMl��A�f,���y��+OU��Q �>ol���/��MR��T�O H:�ѳ��O��'NQ��EybK�jla�"�4j`�ȥ���=I��F_��U�@kt��[��Q$�f����ǒv�D R�!�0Q����)Za|��P�Z��-y�b[<j�BI�e���O�}���A�"�6�d�}�ʙ��ۅ{����k�f���N�a'.����P<S�!�D� u�HAEn��l�8R ��L�TBɔU���N� �h��$�D�v�Q>�� *���"�(h�'/��8�"�I"O���'�!M�� ;��p#�حx�8J�����J,�g~�+�4v3l ��Ԧ"E�y!akR��ybiD-Xy���'��QBT�P �q�L��%g�)|�X�	�uּ��1��;"����e�ڮ���	�j)n��ƋC�~"�V�A�Z�
s ڬ���0�S��yR���u�v�bP-�x�X T�˯��'���+��ȟ����_�`=z9���x���d"O�`�2dL�M�l{�iI�C��i��"Oz�#HMi�J��7�W�
��� D�� 4_��;q�__w.��O�,�j�͐�� � ��~4�d��'�n��$�4SH�HӤڣi%��O���"�$�Y�(އ����1���x�h,�DI�F~��z"OjD
��z;^��£'Z��E�A��H����/9&m��H>�g�M�P���P7LV��"��`%��	<Z$-�ֆu8,�+'c˨��9��X�Zpu'�C�v4����I�Fv�Q���)iP�J[��;d#-�Cx�1t V�cH�*�Կ����%?%>�I�)��:��c�K'�!��#}���)C���jQ��1T�]�s��d�	�Lh��G�L�2��U�1�'fy��[`�n�\l��ꈭ�,���}O��:g��"�N�0U�]�s�>��7�J/qU�(:�H�V��Uj��I���d
�*C⠒&��? �%��H�P�a|�n�F?ʕʷ�ڗ$�\H鶨݌W��;t�oq������k���H�+)�O�����91���bv&�?#Z>(�O���?6%)W�1V��������6�� �b�NE�<�+rf!�dM5��؈c��? L�,b�A3Hd�L���<`��+�dK"4% �DF-�'�y�EB�7�"�2���/#,h� a��y�#֘u	$!B"
>U���#?f�AǠ�$(�����ӕ|��A*���O�x��#r�n��MW�=颙��'�~�SΛ:%N�poZ�k�x��\�P�]@#���]spB��nߚ���oͭ(�I��KXp�z� �r�_�Ъ)!7�z䌴z g�Wrb�A�l�&u��C�,wa�u��S�H��5pi�9"V�B��ޕt2e�L��F��'�,�!�CZ!b�� �� sJY*	�'�\[��B�{�H��p�ɪZ̡�%&��WoD�����Ͱ@�I �iő.bɒ���\$�{f-]�N9�%�M�h�F.Dy���K.k� 駦?D�P��XA�b@s���O���xq�:�I(�i�M0��>��`��e��3׎�7(���G�;D�����
�v�ik��D� �&��LS�<���	��ڷ��	f��~�*����!g��v\XE>�y�b��`i��Bǹ,M68@D�X��?	P�4z!l��$#lO(@��eK�O��A��-�%/Qh���'��@��ŗ9L HmڪN�$BC��4��y� O�DB�I4�L�h�kBTeh,X5m�}�d�h��/_-?o������,� =)�l^�w�d-b���o�C�	%J�z���K�4~iQ���^�zU��ǩL���'�"~Γ?�13�G�+z�p��v#�f��C�I5BIl}0RW�����g+u:�ɑk��-X��'�"UQ�N˹};tXJ6�-O �0�'I�IA4fÌ[�"H@�f�$/���
�'3�=�(�9)��ak� f��d�	�'�"��x��pT�[�f?��:	�'�(jqئ!�$i��l��\K����'hİ �O	��dx�f�,X� ��'�������kI�9��7u� h�'$z�����{��]��Ɏ�kL��z�'x��ǌ$yy���A�"3װ�(
�'��v��{��U�f"�,5��	��'F��;ժ�f�(�!���,fժ��
�'6a��/�Qm�h�G ,]�4�'Oڌ���s�%:�L�?-�I��'P4�kӎк==$5���Q�^-�'��4;P��J�.:���e��s��� \h�	�$'~�1+ϫN���"OT��!%��l���*��P�Ӏ��4"OP`[�@=j�б�$ӟ�� "O@0���?�PV�-4�V �"O,�ä�"��{�C��7�\��V"ObĹ!���W��qeD^�_dL`��"O��z�"�"MN�<c�����Q�%D�lX���0nF� 0C���Vގ�)�"!D��D�P'V�l� %�ȡPB0؁��>D�p�1+̐x��ekU�S�6���4�<D������#Y4��)�̣��=D��h�d�Y�8k���$Fā�w`7D�LA��G�����jT�r�Ѕ�#)D�d
�	��R��;#G��<>�1k��$D��C�M�5��L�!�,b�d����0D���5kѤ/�� ���0��(E.D�;�B���I�� F��<���.�g�Lt:A�� Z0� *�͓ꈌBW�A��D\��f�?�u�ȓ�bb7��5)]�53#	!��l��i�$���W�vB��V-A�I �ȓ?)��C�L�1;�}��ׅ'����B���㔌HSP����
ǪhXlp��eN�1C�ŏ)����B(�7o���=)�h�7S���A�Z�@}c��9$��I�P�B1N��IsI�����,�*�'zC��v�ɊZ��JF��9�T5��n6���Uk^j�)�'!�����옪o��x� �a��X��#�/Kˌ��i��<&�i�|��}�S��I��gH���� @������Vs.O�zbH39��>�|�h�	u�Xx7��wA�l����d�w@�h���T?y�;�L�pKØk�1����9�,}�'�H9j	�Y�S�O�<5��&Ŕ�C`bZ�k�e �'�*�iBl�|�	�ʈ�`�K�&Qudͣ6�O�8Ɯa�,F9DhqX�O�=�h����>	�O'8p�b(W���L�%���0� �:d9�'�v7m���>ɂş�Rg*)h�Ȥ>4\�B��5[Y�F���O?�����<!1��r�	#w��Y�k�<��ύ&4�p��� 6��HF	H{�<�R�"v�
�Ξ�TY�`���C]X�h�O}��nOb���"��M8����""O��Sa��?M���B��
�2]�@"O�y�̒8rk����B=g��uq"OxP�A �CWȥ��؞{�4y�4"O�%� 9o�2�Jw�L 9�RQ9"O؄soGE�������K��H��"Od�[���,.̒d�w�_q�h ��"O�$���)ʊ�j�O�&��Uâ"O�1���(,��)�$!(��5�G"O���OB9��:ƨ��|
l��"O^H8�I�9(9x,����4t����6"O����r��=%k�C�rH�t"O���mCP��K���<�RЛu"O�	�C��W}N�S��� ��"O�i@g�,zA�1C��!]����"OLŉ$瀼m!�	@�T ��Q��"ON}��E�'��t"�+݌>q�0c"O��ڕ�I2O��`J�eR��k�"O�A)a��"7?b��U�B�~5nxؕ"O����jm��;�D��;N�m �"O(��B���]�8��GC��48`P��"O:u��ɗg�:$Y�#c��;"O��@�E�7i$֝Ya@�  >q��"O���LQ�^@ 0`��E(Y���A"OT�2��C�)�2icG�XsU����"OJ9�t,.}M�\��gY1;�0�F"O�0!G	�e.��ԇ��$9��07"O�!�®\X)��Q*.�y0�"O� �8kcł�E��4&#��"O��t*f�B�e�="�3U"O:���%t�x�	$����MP�"O�u��g�=?PQ9t#	,sN9�"Ou�s�t�����<l�TJ$"OM��P�+���@���QjE"O�����.X�pjB̒&��('"O����悎8��Cl�#J��j�"O��z��%	q<�3Kհ	D��%"O�hR6�V0Fs�m�-�(9�Ր�"OV�7�
<���R�V4b���7"O���j�5=��`�,z��	�"O��8�/� Tz:*s*Z))ܹ��"O|<�H��<jL����Qx�#F"On�	�i�h������7pݐ�"O��H��2x�^U�EMXG�|U�"O��o�W^��2�D0a��4�"OxM��D��-�\�'���U�R0��"Of,���"UM�Y����j}���"O�yY�g+K�(!#M k���"O,�r�Ê�$���FJ �����"O;�k�&U<}�PI
V����"O`M��'�"e�dI����^�:m��"O
\���KL���I����D����"O�qP�7<>�X ���%�L�W"Oʵ����k�����5�<�
R"Ov1�����" :a���4p(]Г"O�	6�Ѡq���t&~]N���"O(@�D��x�z��@j-?T�q"O�U��K"r�zX��* J�̛1"O�}�3aնX,1�*Ŧu18� a"O���m��,�\�S�@�N��=��"O`A���M;N�V��)?1����""Oj(�d
R QrL�`����m"C"O��� jD� .�ݠPi��̺��"O��+t���J��0�'�8f-�r"O���V��?<Į�9���[H	s"O �����h��ubeG	H��arS"O�0!�Ȓ�$A���))�`C"O<t+F�1k�f���D�8�Aӂ"O�`��ҼqD<]��qn���b"O��07A�wh���mߙA����"Op�j�ʌ�%����]��P��"O���b�6��$b���.i.���"O�T�C
�@� �a0�-	s0:s"O� R�����p�!$P-$Uj��"O�uA�La�$�if��;aG���"Od1v]�n`�ac��p���2"O�|��ኇy��4�2F6Y��T��"OV ���G0XPsw�o�pi"O�!`��1ح�����7���"O�
7��an����
�x��ȥ"O��sU��
p�Ȃ�͟fž ��"O�0gJ̶1Z�Uڗ([���!"OQWD� x���WAφe��)!"O�y1" 52��)����/O�E"O����ʶU�j倲/Y�D4(B"O�h��D�@����Ѝ�k��R�"O��'�L��1��M�R����"O|}���ͨf䙻5l�&[���SF"O��Y��(�Bm�R��q[��&"Ob$ZD�$8R=6�ZY���"On�eJݑ.Y�e��{�H|�d"O���sΔO]4��s�/ �8���"O� x���H��C��DAF�҃S�ڕ "O�Yy���nf�h�������"Ot �k˕xtv�@�`����C"O���5���vu��)S+sDH,8D"O��� �lː�I����hA"O�xy J�%DJYZq��@��"O! ��l�
��eCK3gsZE:"O(��q�G�5'��; `�3F
fl��"O�{���[h��n��8ڤ"Oνb��@���Y6��3�l"V"O��YR@��id�{tɻ��XYC"O*H��İ�p�t�T�&�A"Oҙ�%��2���֯ۃ	�n�� "O��2QZ-�|)BTO?�H8��"OZD�u���BeY( B�
�%j�!��2I��U0�%�-N�!�N���!�D�p�*=[��T(I`��֣��5�!�[\ƌ��W���!��'���Z�!�D��U\� �F"��1��jU�_�P�!�$��4�-b�,ֹJV�Z �dY�'.pI����8�����χ%��Q�'u�
��	�l0w��&gN��
�'�\�x��܊(����N�E2 �
�'Ƹ�Q��*�l�v"޿0^��
�'[$I�!�yW��f��z��
�'�����/c=��3� R&$0�xA�'��i�-/�DH���ӠO�-Z
�'B��S�BR�~r�kgȄ'��T�	�'K�96��޾�a�Q�t���'��}�"٬�a��#���#�'VZ��cm��B��l� =+nf���'��k>]��K�Z�����'�ls��(d���nO3���2�'T�Q@�MB�~h�Y1�ض��'xؖG�l��pC/1�p@��'�<�"���l�>iR�aU1}pA�'�T�����K�2�`���8
�'8.��£�+53@i1� Z!6��
�'`Bٸ��X_l1�0�C�;�A�	�'�8��Oъ��D1�8>�Y�'�"�J�KB�z�t�(!���7����'(��l��9:�x�F�0/����'�)���W#�,�A���'�f�*�'���ЭȲ5��/��T6�8
�'�nH�e�p�ɅZ1vՁ�ƞ��y2���C��ǐ�b�d9w�ݟ�y@��=J�)P�H|���Y���ȓ��ZkT'M�,�Dn�
?0,$��O�La��ٌ(&�B�i� �B��� �� #�C�S��s�)/^�����7��{t�]�!����V�]�L��ȓ-v0p��@6$v\ ��.���ȓ}�5@%��V��:��U$x�)�����!UڥU���6�X	1�N]��e�04SSJ^���e@���M�l�ȓ%�X�JB֑TR�iY2�������pf��xB�	�1$����"0	�l�� O��i`���@�}�e ���̤�ȓ|�*�Q�!u��<���O�Ah����(��-b� /t�Ni�
uW�<��N�][CJQ�q���a��-HŌp�ȓ#z�$�ªJ$)A��9��gu���;,���Q��&h�a��K(9r��ȓoy\%�vj�Z�P	b�i�y�\���S�? �|3" 
!A��a�� N+=L��w"Oػ&�}D�X��
 ��S"OAj��،Wd��S`��;���	"O��y�@L*ע�C  ^![^���"Onu���2_��	��I�$ �x��"O��Xϻ�9��OO���z�"OD0.�Rh듇�>O�����A�3�!��M��ूIX'q������^��!�7"�����͝Cg|�b�ƕ	Y!�$�34�Z�����?EG 8�$�(D!�$D�[��\x'�ͦ#�bFa�W>!�$�~]�)�g��-U�8�f`1qM!��֛|�5@�-�	3E��,@!�$
Z��*�1�,��AV�L
!�E�@M��3V	��f��K�a���!�d��XK� }����n�%,E!� �G��#7��u�=X m!�D3Bւ�r�,E�h��h���"!��҂{��#ԙ9�0����;�!�D�dfB/I�*��P悭9�!�G�L�`E+%@��Lz��A�V U�!�D�)ۊl���*o��	��?m�!��ݫD�ޠ ��=�������'Nw!��2%u�%���ҴH��c¤Z_!�DN
4Ѝ�g&C�yX�D�#�k2!�ܒ��ꂠ��tG.�(�۸K!�$��~�@s�S�u=�̻�/�?v�!�$�tN�4ض�#,�i3��9%�!�$�X��8q�I,8H>@3Nv�!���p�X2�\
h�\h�J/@�!�R����S%Dsƨ��)] `�!�ė�@�BȺ�-}S�k�Ζ��!�D�26}z0۲�
R�Fpm��Xs!�$�gZ�-�nO�}�&����Q!�d�[?���G�%6�=xt�@�"!��5VR�����랥��o!�d�:)
����a��{�f]4��!�D΀ �ڕ���R��.��@��7�!�Ĕ�>K- `�9�D�$�L��P"OzP#��	��9x�m��m=���2"Obٻ月2��Y�l�X&<X�"Ov�§�!^ Z@	�,+�tXz�"Op-��̘DrL`ć̽@�P��"OT)9����8y6�/����"O��(��"��`q�)ݭ"��%hD"O�icՉ��j�ECN��X9J�"O���q
 
  ��   �  �      .*  {5  "A  �L  �W  �^  �i  s  Zy  �  ��  @�  ��  �  T�  ȥ  	�  M�  ��  Ҿ  �  W�  ��  ��  ��  V�  ��  @�  �  P � � � @! �' �- �.  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%_�Q���m���R Q�t�A�,�Or@���A0��, '"ѽv�d��"O쌩��9al��;P���u����"O��d�AR	�N��>����3"OTP
0U@F`�q-�#D��`��'�I%y��]����Q�}���7i���$�>Q��ۑeK,āc��/:TR	еO�'���,�r@k�� c�x�x�iY+bB䉇KxHA�ׄӏO�jM�6��TK��	��'"�>�Ɍ[���zA&��D�Hq�2BQ<S?P̐�'��L)��?z�(�4[0�`��ٴ8!!�4��'�
*m�������q)�{��d��\���䚀r�V�+�;<��{��)Z��K���ѲBKG�,�4��� @�<��B_y�NtCD៙n���S��զqE{���i����j� ��i�1B\�#
ϓ�O�zP@C!p��2�"��yv>(��3O�E{��I;Z7��@'�4r}c�N�W<!��6
�\������椚�2.�P<">�J>yPmS�e�f��N�(3�v q4��H��p=�!`�=Ԝ�J9$���� ]��hO�'
Cn�HRJ��Y<��'A����mM(<�p��=�q��ǹh�����Z�<	���y�>�1�L�8`�B W�<�ЄJ�H�m2w#��x-�%��P�<�ތ��̀�ʘ.f� TO�N�<�#�	n��(�%�֢$Xd���$�"�hO?牝��A4'��Hh;@�*`u�C�	"���(P�"xyv�[J�Db��n~���O�Н(���O�^,
c�Z{��AI���dE'�2x�%
H�ض�ʵ����'?���'��x���7:R��g�'Kn`��d��?q�'ȰY쎄 ��G��n`��'ή����D�p�!Q�P�v4� �'�H�b3�Țe ApQ�\��{5"O�M3`+�`� � �^�4��g��Ȅ�ɖ;��2�.�2ye<Lڔ̒�7sF��d!}��<-.YS�%Ԁ	��l��L��y"��!!X0�Tc[O�2e0�N@��y"G�:?���D��I���RD��y�hHP�m��ȈF��Y�#E��y2���}qx�b��R�����'��?�����1Vj<CƦ��?��0�2,7D�dhAAڒ ��@I����Nx�	D�3D��9��4WS�ț���	2���A1D�� �YCu���~ۘ�!��t���zA�'�!�d�j$�8��1���c��sp!�$���`���ݙ^�&P�&IҮ,T!�%d��]��a
R�J����[�QF!�dZG ����]!���&@�>!�V?�N�؅	���H�-��O��8�S�Oavu��䎘���N2b���8�'-����<2��:�'��M�~("�O���I��<����O�7k�ڔ��0���>A�`ٽ����]�c��p�uj�ޟH���vx���F��:|ʢk�rΔA��F~���]8�E�C��c�P�*�'��
^C���i���9�A��T �~��)ڧ&�q����1��P�W,�4F����ȓ2�\LA`�W��<ё$O�<��)���hO�>�xe`��5���s�H�s��p�6D�\�r�H�<��u��؁B��g4?ɫO����!V���sЖ�hA��:��~�T�l2��Az�y��'ա77 ��%F0�IA�����&��@�y�&�U$j{�dA�d/D�P����� <Y��(TZ���A�?�IS�az�h],8T"(A D�?e�Y�B)�M����s��x{�f^&�~�*���?Z�ZY��"O�X�T�L�.AV�ZG�Α����1OH���df���5K@��B��Z�k!�$/Ei�M;�䂅}��0XUfܢ_!!����AsE�e����߅!�ѵ
]f�ȕl����3/�!�e�V�
�M
+����B�"�!��ǟHH4Pɱ@D�d���QQ@�y!�Ȗy�~��VA�tI�'mӳ>f!���1L�0a��3J��(���k�!�E 1<�v�τW0(��ѳV�!��$pӀ�b#��K�pl�-���!��%~�H3�M�&�N� Q��I�!�D�"Ap�<i��+p��aaqO@#\�!��³m��x�pk�.vV�)���x�!�d��00b���J=nY����U0�!��6C���l� �� ���$�!�d��"-�ixk�<���ʅ��+	�!�d���̺��
X�����CJ�"}!�d��G�U��}����-�!���o{�e�$]�d���1�wb!�� ��2�2R�`D�m;�]-@_!�Ę�D~�1�t$Ϋ �>�{�Ãw[!����Mp��>#�
<i2%°l�!�����`��7�$0� ��2t�!�ć���2*�B�l}"� �,�!��=F��n��Ҷ׊F�!�$ӽSq6�x�%%au|�o\/X�!���
s�� X�nQ�� ��-�#!�D��;.��q�#�4����"W!!��͏��+S�P�|��кBQ%R7!�d�����A�m�{�ݻ`��&!��rC��C"J�j^6ps��6`6!��@���5 )�����K�y�!�Dޙr*���&�m}h�����!
�!�-u��ar�[5:>���d�D$]	!򤘩~��l��`�!����7��!�!��~�8á,I�x(q�G#�!�D�y�hcB�ޅc��	b3 �4�!�$=�4�x��$�B�N-i�!�D�E�!���E����2�R�7�!�dB� ]Ri��GC�4 UB��K�h�!�� ��aY�X����H5� �10"O���A,M�x�x�O��2�v���"O��W�	-m���^i�N�2"O �bQȃcY˃��gf�x�"O����T*�^�5�`T� �'��'or�'}�'��'	��'@&�y�@8� U�
O��N���'8"�'���'o��'�R�'��'jMe�L�0��o��K[�� ��'���'���'f��'r��'W�'���N�.@~��p�6�#V�'��'���'��'��'d��'��t�$��hk� K���-~Pሳ�'U�'���'"�'_�'R�'g.�B�_�^��A��49�ae�'��'�R�'�b�'��'*�'���Ӽ�ⱡw�k��S�'_b�'�b�'u��'�R�'FB�'jV�1!N�vw��I6��+��lSd�'���'c�'S��'S��'���'�V ��Dޮ�B��0�̈O�e��'���'x"�'�"�'R�'��'������.-np
�G+Q���2�' �'c��'�R�';��'���'.d�P��C�k�Y�0�*$�"3�'3��'xb�'�b�'$R�'���'=����"
�{r�@)�ǎ%I~A���'2��'b��'Or�'d��'C"�'<�e�B�K�%���M 2 � 1Q�'���'�R�'"��'M"�m�����OR��DR&��q��#0Pt�u'Mxy��'��)�3?a��ibA��ӄv ���������;��$K˦A�?��<��#E<W��	At�����-,b�3��?y�k �M��O��ӝ��M?��7�O}�C�ޱc �B�� ��Ė'7�>)����80P b*-'�:���)���MS�@F̓��O�B7=J��̌�A�� -�&�#�f�O��dz�֧�O�l@�V�i	��ܔt�x�*Ħ�A�8��-�J�v�,�(��=�'�?�R��" Sх�%h,��:���<�(O��O��l��0:.c�Hz�
[|y�"R�%���$��d��?��	ڟx�	�<ɭO�!LT;i�j���|������dM8�*擁dL��ݟ���ê1e�]�f�/��X��Hyb]���)��<��� i3�,��"�sxiqF��<���i &���O�(n�g��|򥅖nP�<*$�L�8m�t+��<����?!�K0)2ܴ��m>т��ZRȕ*�E	)���Ӆ�<�ީf�<��<ͧ�?����?a���?��-ƴ͠i�V�t�)�/����]צ�tN��\��̟�&?Y�	�1b =���S-:L�3NHWw�TȪO*�d)�)�����R�>t�xf��JU���3�H�( 2��'!*�	�B�����0�|�R�L�S`Iv
@��&ɏ>\���;�L%�OlQnZf�VX���s��Y`�&B�%����t@�P��@��&�Mk����>���?ͻl2A#�E#F��[o��_e���'o�<�M[�O|��/A���D����w��� c�G�@u:��Ee[2�B�Q�'��'w�'���'V�X��=RI�ht�޷~lL�A�J�O����O|�o�3X����|B��c'����O� G:m��ɇ��'�X�L"�'�צ��'���9�kRho�� TH�4)��$;V�
j�"��B��'��I����ԟ ��~����`M�l(+A�X/}�!�	⟈�'�46����O���|�QCaߖ�p��a�|a����<I�Z�I�����r�)���
�t��Ui��k���U_�x�0���P4����,O���?Y�:�$P�a.<:!B�V�q�"팹*?j���OH���O���	�<iV�i��-xဆw�T���Xa�<�8���72�'��7-2�I���d�O6�z�A��8DV��IyT��Jvm�<����M��O�	:B$T��Gű<�3-�3�������4�^�!T��<�)O��$�O��D�O:���O2˧a�4���x��AX���0� x4�in!�%�'
��'��O�{��.�s�l�$��-I��H�e^:�R���O(�O1���up�&�8~#J��!�/>5l��
�����ɹ|.��c�O��Of��|��rYP� G'o�,p)����!����?I���?�)O�pmZ�j�X�I͟��	��,%�$	��l�v(#���6�68�?�uU�$����'���P)50x�b����"�X��-?q��[	9�!2��B�'8��č��?a ,00#S*^9��8�+ˁ�?����?���?���)�Oz$`�j�<0�\y�3ɊA+�/�O��l��1좕����ٴ���y�)�$��Q7�#���f�2��������ןh�v������'^�iYTl��?eҀF��O��K���9+d)9�" �hi�'�i>��I��Iß��I��60���yťIH+�����wyrcp��3��O��D�O�����$�l}:4
��
.N�l���QXS@��'�r��P:��B�7\,�FA��9�^�*�nԬVV�ʓa�`3A�OPY�I>))O�T�4��<�F�P����qp�?rr�'8�'��Ok�I+�Mt�[9�?Ie	ÛC�.���ݤc��5��P9�?Q��i:�OM�'���'�r��+oXa���G*AOI�c 
 Y�j����i�	(Pd͠��ORq�B�� h���O���&�#'��d
��I=O��d�O����O"�d�Ol�?e"����^�~��&Ҙ<��yC�����	͟���4s%<��'�?�նi/�'5��KC�(2'����Ԥ\����u�|��'0�Oc�	�@�i�	���$�)B<����"8�*ч���5���<y��?����?y�����7�փ#��|3&:�?A����D��Y`W(
ß���ҟ�O�r�C!I�_xN��שȅm����O�u�'O��'ɧ�)�*V6��C'�X�j������a{`e�jN�xѕ��<ͧpm��V6��c��BE�(&9b0k�F��q����?����?I�Ş��d����g���`�$�V}lD	2��+LW�����A�4���?	 S�<�I�e�`Ӳ�ĕZ�b��t �<��������HǕΦ��'۴�81��m�+OB(^R2��"S�X8^��y�Y�l�	��I�����֟P�O�8��gn��Q�Z���e�����M�x��f��Q���'������'ZL7=��Am��OӾihר$Pi��E��O6�b>�ib!@ڦ��t��g�H<%�\����ۖQ&�E͓y���+�m�O�mQO>*O����O�@���Q�F��9��CK�A@r]Zqc�O@���O����<a׿i�tU�a�'���'X�%�IO]��C�d\����D�M}��'R�|2��M4�A�Ԍ��"�P�85ϛ<���9{E੊�o�7|1���y����:n�t�Y���9\�	��F#!�$D�W� ��g΢h��DHF�K�sZ���ma/[ܟ|�	��Mc��w�D �0�8�@`�m� Q��'#��'�©�_����h�%��G��i�Ds�5:��ƃw]��T%o
��O�ʓ�?����?y��?��sK.��툓M�A���~��H.O�o7������x�Ig������W~z��G��%Qeh�ZģU����On��5��*���C���z4a %�>A��I���=1l�˓:��M�e�Oа�M>�/Ohm����8R�
9Ip..�,����O����O���O��<!�iP��s�'R�:�e�18:�;��5UN�7�'�R6-'�	�����O*�d�Oְ�����.�"��ȯz�lӐոe�6M=?9��F62-�|j��<��?Tj
}8P��
W��Y1Mx�$��I怹��.;' �!�
&iQZq�	����	��M���k��Fdӈ�Ox]�	��[Ԓ�r`�G=0����7�d�O0�4�^��Iz���^<Dj0%�6+�C�(���ZZ��$RZ�Ip�IFy�'?��'2�J�+lJ)q���V�LP£���B�'�剱�McFF���?����?A,���SHQ�
��i; j�)Kf8��G����O8���O�O���.(���g�ZY�L@�
U�q��]�2��f��]�5�&?�';�
�$��pq��Q�m��2x ��������?����?9�S�'��Uצ�%�?O7���1� c��x�)Q>�����<��4��'����?� oًqxx��!�`��q9�GL��?9��P�iܴ���v�Jk�'���-U,4�a���6{���r��3&���I_y��'�R�'X��'�^>��`ߐf�屴� 1*��9���M����?��?!K~�tݛ�w�R��ro�YT�GlB�Z��F�'7��|��D��v�V:OL��QL�{���a���
��]2�:O0-`�N\��?�p�1�d�<y���?y�������z��"�	��?a���?q���L��&)Mß�	�����J	5Ym*����.�8�@��Q_��Rr�	����F�I=.ȝ�+�_6r1Bϧm�� �0�2�b��Mc��� l?���[��I��ӷ�4�¡�K�`�|B���?a��?����h��܈5�ѣr@�u��1kgo�1|���D�����lT�������M;L>I�Ӽ���� �"j��Z8��S���<	���?1�]�FpCش��� ���(��On���w������j�8n�&� s�|"Z���	ԟ��I�(�I������>9���a��-d�z5����QyB`�8�1���O����O�����Dʺ_�������v��4�� T�E�'���'rɧ�O^�$�����Na���(/!�&�6�h���O:�@���?��,�d�<�S����M�ō�8�J\�Qh����O���O�<�`�i�l����'|0��ɛ)^|�yAF�S��+��'�7�*��%����O����Ops�eB�&�ޡG⒓i��$ˣoRH9�62?1���>ݔ��(����!3��Pp�d�!A*A�5��8�Ek����ԟ�	��l���������1#�<�0`ע�Х��j�?���?ْ�i,�Y��Oc�)gӦ�O��`�`S(b������dZ����O����L`ݴ����m�D�e��k�����]GP��e͔�?��a �$�<�b��1
5����S5u`��b"�1�O�4l�.�*��I˟���I��ߚ!�0�e㚛;�@�NG����V{}��'~"�|ʟN���[	�^��'�_���\#�������2fO׏{ul��|JF*�O���O>i����{�F]a�B��Ta�~<	t�i��]iǁ�4%���`ЂB^>\�פv2�'�r7�*�I�����O�V�\Vz!S1A�(vn�A��$���?���pA�d�۴��d��~�|���Y�� ���rΧ
ɢ�Zti�]'�dCd6O���?q��?���?�����	ǧoI���T;0�y� (��"��n;[بP�I��	L���`�����GJ��`p�*L�c~�!��1�?����ŞdY���ٴ�y���i+U��3p๘B�F+�y���R7�E�	�)}�'1�	_yB �(0�@����%<��Y�MX��0<�c�iך�Y��'���'�|�@I0P-�`�%E)��z���SW}B�'���|��--����	W3�F!��Ǯ����F��2�|�'?QQ�O���Z���Snݥ%�ʠP���*,���d�O��D�OX�D=�'�?�o݄�`F�Y�C�j�5��4�?ɓ�i�P�c$�'��x����]
'4��c��˒��0%������ܟ,��ʟ�s�)_ܦu�'*LIA"�b����I���� �}��6O؟�����OZ�d�O����O����)1�E۔ �CJ$���BEH�ě�"٠(�'����'�0�%!׆"+�d����pđ�7@�>Y���?�K>�|Z#e�|>`(�0oÍ w�h�@)_�4�����CG[~R�R�p~���	�6�'}�ɥS�%Qi�vÌu�'�O<vV����ڟ�I韨�i>͕'�7M��*��B1~,����B�r�ܐkS�>B�*�d�צq�?�TV����ןD�	���Hb�E\���¦��A h$�ǩO��-�'5���G�?1�}�����5:�CY W�E�q�!�N��?q��?���?1���O0����+r� ��� Z�����'���'��7M[([\�)�O
�n�`�9%�\k�� !I޵�cތYp�`$�4���擄V��lb~Zw��@G�G�\`��,[�	a��1��uS��s�	Ny��'���'¦�<_�.H`���lH�9���G�~"�'��I��M�f��/�?���?a,��$��� Z����l#`��US����O0���OF�O�S�9�.�ya텅a�N��ɞ�4����s�(\�>(8?��"�'��%�P��(�.2>�q�ˇ-���w�D埘�Iǟ�I͟b>}�'��6���"F2E+���g58� �l"1AqD�OD�D�ͦm�?�P�D�I�s�܀�{�� �#NԪ{RR�'h���.�����-�Z2�)�9���ࢄ�Q�"!1���E�ľ<���?����?����?A/�:(C��?@1�*�;X�.�#�ʦ����_y��'�Ob���Y�����Ү��n>,�5�^ ZJ��$�OʓO1���B#p�Z�	�4rBi�t+�`k�`�_���'�<e
�!Z?�H>�(O���OPjҭ�9t~���!8j����gn�OT���O���<1G�i�:���'@��'�"���߸[RhW4{���7�D�}}��'��Oha{�n�:+� �@6�i6�� ��D��o�!�<�(���"���^�T�d�1��e�w��QX��A^����Iݟ4�����G�$�'��yУ���$�ڼ �Y;.������'� 7m�1p��O�Do�e�Ӽ+&�.V�LE�B˸d|�Đ���<a����D�(�J7�;?AƧN<2�).�����8$������)bE�K>�-O����O����O~���O�|�$%P�_'2�	�ʒ�W.j	�a)�<��i���{�'[��'�OZB���@[%`[;R!�y��L�Q�N��?	����S�'/���UDڜs�ݱQ�ɣ_n�[`k��E�Qx-O&|isN-�?�F�<��<9ӭ��|��@J���zAB�K��B6�?����?����?�'��SۦX@ٟx)f(I?s<9r�0	�j�����ן�"ڴ��'9���?����?iS�Ƥy7�Ը��Ζ$��͒Q��2+H���4��dF�hD������Oo7왺��t����)�ꑀ�y��''��'���'��iZ06V���C&�%G��@���F���O��Ŧ%��L`>��	 �M�M>��N8DͲ���mR�Z$yɄ	<�䓮?���|Z�[9�M��O�NE�	�&eh�-b���fC�=��P��O6hL>9(O���O���Ox��1���=�n	�ч�|��e����Ov�$�<AU�i������'���'��	��4���G\�DXDo�����J���ß��?�O��h�g�Y�T�a2 ;Ą:#������HU���i>Ợ�'`V&��0D//񃧇��s�F�k�%�����I���	��b>I�'nT7��p
b!��.�x����c�@��!�O������?��^�����5��cÂ;_�b�v$]Ey�������Ҧ9�u�Ƃ>^���$]@y"��Yc���q ��eܕ�JD�y"V����|�	ԟh��͟��O��l���_�h1�m£Lf0��mlӂZ�K�O����O2�����Ȧ�A��{wf7$��i�-�<{���I�P'�b>�� ߦ5�=Y�խ��Ig�ds�bC)]�đ�^�vh�dƬ��&�p����'�:̒�oNg�����G��9z��'�b�'�[�,��4;��I#��?�����1L�?���"�k[�0PI>y��.2���x�Is�I/Q�P�")��
WZY`����\���6���ͽ*�x�O~��i�Ol��RO\��c	�b7�}�!
)�$����?����?y��h�D��ِ~�
Q�d�܈�<)��Q�S��������0�	��MK��wό�����H)�P�	I�\=a�'KRW� ҩDڦ��'�I�D���?��� ��r�g�8/���Z�f<�!�%��<a��?���?����?!QO���Rd�6�B�9Ƹ��B�>���禽�i�ޟ��͟x'?�	�!�r}1��@.���i6u��e˫O���(�)�<)M�a[���Q"fd�%%"�:���e��'�� ��lʟ`ל|�\� CD��{�T$�B�_#"��2�E�����矬�I��SEyrm���0�x>iA�1� ���K�SD�u���O�l�B�&:�	�Д'yz< &D��F���R�)
K�&m�T�� `(����,�ԂӜ
�4��d������3#��������-K��*rNr��Iן����I����U�_4M4��&��AZ �� (� �?Q��?)f�i��i�Oc�(jӞ�O��K ,`&���=xI��G8���O4�4���ĤaӞ�Ӻ��V��B��
5d����a�uF��cM[x�މ��o�Ym8p9dY�5`�l��T�.���YB�u��/�I�b��3��%ymJ�[��
**�����D�sA.7���F�a��ɩ�B�]%1OXx��c�-�~Ї4kpy���(=��JA�Ƃx$�qˆ!�~_r )B��D|(���z,:�A6� �<��y/�<�4�c��<L����ŃQ�j!j��&hn�bg�Lvl��)���0"&�*`B��aE���E��ݸ")'U|�:�荛i�^��a�S����b�h�,P@%L
0I��a��iAR�'�"�O�Ũ`�
0xM �N��x���Q3+&�$�OT��Q"Yb����s�X5��8��rf
F3'D�m�ayB�S��6��O���O���DX}Zcm� �c��#�
X�CC��������Id��Ix�S�'c|��Ϟ�G��1
j8�m��j�����4�?!��?���|��Ixy��C� ��4���Ӫ3�v�0.���Żi>��0��8��ǟ���+��8�����T�aG:�MS��?	�*�@��U�<�'�2�O�5"�NW�B��m��"��dQ"�J�i��'3⁲�'��O^���OʩC�dPo>���H?�Z���
�	��;��8��O����7�5����@q���4D��M{P��1w�lM)�W��xBM���0�'B�'�X�����X&3G�9�v��vx�@��ˌE)�O�ʓ�?�K>I��?�����W��(���zQ!����6�jM>���?����D
(��ϧqjK�`�,d�����fUuiҝo�byB�'��'�R�'�,����O\�I��R�z(��M#'p�P�\�T����ByR�ƚ�맇?A�@A�NL�t��5}���N�rś6�'��'�"�'�6�Z��dŁ�4x�q��'iN�P�R)d؛�'o2]����������O��գ�`�)*��ؚ�D8� Y+F�	r�Iɟ�Ɏ-�(�?y�O@zu��:����im�����MS+O�eؑ��E��۟����?]�Okl*jtܽ!�J��:�>�9w,�5g��V�'�b�Ձ��O��>����ǚ8��Q�wØ"5Vn��o��@�g������՟����?M"O<�'M?\� 'c��S�h)�(^)�>����i���'�2�|ʟ�D�O���1� k��M�4G
1S�)��&Qܦ}������ɚRdڄ�K<ͧ�?�'�ภ�̏;L]j�
\*]����ٴ�?�I>��S?�I�x���4��#.�h%���!���$&��M��FB�P��x�O���|�%f�4Kt�Нs��U���ӇY4�O���,��|Γ�?���B�l�"Ƒ7&�n0aQHI�@T!(O����O�㟔�Ip?�0��+�:��$��B] ��T�����m#���L�'��f�	d��)Р�Jqr��^>�@xV�Jڛ��'�����O�ʓ5%��mZ�(b�ˀf^8#Z��#��0w$pO,�$�<�P���*�|�dCTNJ���/(�R٫5�#`���my���?)/O�$Px2C�k��
D�<r2�q�끺�Ms����OD��0l�|R��?Q��%�X�ϼ|�G�Rb�KP�5� O*�ĵ<�a�L��u�cļTg���gG�.�
Af厖���O"�F(�O��$�Of�$���Ӻ��F�Q���±�
.�"�Z�/]�����Ry�.�O�O~�i	$D��@v~��;�4U�������?����?�'��?�i�E�$fT`ɡ"UJ/�t�K���䔱jV�b>A�	$¾���!�/<B9��I�`F0@�4�?����?)�"&v+���D�'�2�҆�,����T~`�$�D1iҐ7M�O���<�\?��O:�O���7I�/J��Ĺ�![_u�`�P�i���8V�	����+�I�I�~Y��G��	����7,S� ���O<y��Y~r�'���'��O��,	�!�#JN����[o���&�(���?A���?)+Of�$�?U���T�q^d�h��|�CfDeӀ���<���?���򄕃C�\�̧ ���2�L�C�,����נGZ`@lZsyr�'��	��������a�(+�
A�l�ޥ!gi��*c�ǖ���O&�$�O�ʓd�`� ]?I�	�l��4FjL�Ajܠi�Ώw����4�?1.O|�D�O���W�Kz��O �	j���q"��c󀽲QD�5:b7�O��D�<)P	5 ��S���I�?�v�Q����̀�
OR�
����O���Oj��C�?5�'o��7]���/@�y��=U^��S�tz�H�M����?����
�W��#��)�%N�&��i�P#ѥU
�6�O��D��2H�Ifyr���'uD��@�J�N�
��f�23\�6����Z7��O����Of�i�k}R]�H#
� �9�P�F;�N@�rk��M���p7�i�vi��'T�I�P����� *��	!=�z]a�o;r@}A��i<"�'�bKC8/�V�����O�I�$F&�!�NיU�xzD�Z���ܴ�?q/O��0�4O�S矀�I��$I^�j�@Ð��~t��0$C�MC�pp$P�_�䕧oZNy���5FKS(�K�:7G����H>Gr(��'��1��'��	�(�	ߟ��'�|�V�P4g�%�1�r���ʀʀjM���$�O���?���?y��X3F�1*V��m!��ƣi:���?����?��?i.Oॠ�h�|"g�8Rd6 �h��`��d������'��Q����Ɵ����?�l�<n	�ƀ�N�`�2V�k�J�lZ���	����	IyBJ@7xXD�'�?�%`� y���Ae� �0�\R5!&h�6�'����D�����Oi����M�q)ÐT��S�4�����ͦ9��ğ�'�����~r���?1��C6��C�S�s4�уD�������R���I�<�I���"<��O������>A����$գ���Ѧ��'eR�c��~���$�O�������קu7��е	6IY. ]RҥX3�M{��?� ��<q&^?��L�'
]�����%���2�]8��<o� 6Ri��4�?)���?��'qx�I{y#��< `�!�׶xBhl�� &|^7�T�(w�$(�d$�Sџ؁�(S%n%0�s�㎫;���;�k�,�M��?y��/��P2S���'Z��O�=�VL�"��x�HƯs��=�i�RT����x���?����?�V�; ���bHB$�E�����ش�?��n
$ez�IKy��'��	˟�Ohą�%c�&�H:c!�:'���6�����$�O<���O&�d�^t+şR�L����IeeVu�#�M=���dyR�'i���,�	ş\;Q��/^y��F3��z��/����ǟ��	�<��h��'%Np�e�f>��3oI��x��*P:k��@դy����?�-O����O��d�1l���*�(AQc�O>P��j���&�oZ埄�	̟���Dy2Ƕ'��꧌?��<��� �M��ic�����Q~�o���'���'�b��,��	����)�P��M�6��Q�v�!2�yӤ��O$�}��p��P?i�	����Ӣ��Uq�֚ ���숀Q�Tyr�O��$�O���*%��ĭ|Γ��t��[�5����=+�XqӀ̂�M�*O&IP�^ۦ���ן0���?1p�O�nC=<�����_ds���/ӛ��'�2#�,�y�c�~Γ�OH�P�G �<����&��
 T�{ݴ&��b��i���'���Ot���'B�'��Q�ҧ�9t��`��"@X �Bf�uӶŊm�O˓���t�ߟܨF��̠�p`#�7\}��PQ V��M����?���7����T���'��O�MZ6,�|Jp�zfk��[\ ��X��'��x�O���O���O���/�$~�r]���W<��C�������I�_!T���O8��?�+O:��ƞq��*
:b��i����Zq��[�,�wFd�$��ğ�I�����y��Ӆ&�"Q�6�U�ڇ>�vQCA�>	.O��<��?q�m���2��^�b�,��D���IjƘ{1��<��?Q���?!���d� �A̧9~�M���=��[���1#G�}o�syb�'������ş(Ѵ�g� �4kKo�t��L�o��PQ%�'����O���O>�EʁI�]?Q�	oZ�`�ph�
Il��!N�F�6`"޴�?�)O��$�Op���=ZY�$�O6���^�[���70#^]�d-�����n�ß���ky�l����'�?����Qo����P
b;V)QElT�v��	������t�W�j���y�ޟZ!!w��b&ʸh�f���T���i��	�z�=�ݴ�?i��?�����i�-`eΡ1�t�b�0B�Z�I�Cj�.��O>�9OpH��y"���P������:-���(W2�6��W<�7��O���O���x}"X�h�E�k���q"�d������M�gA��<I����d4��џ����W�"-X҉ �,^H���k!�M����?)��_9���3T�,�'���O��y�B�nՐ�bU�V%6����i��]� �p�c���?���?q�Z�w#bQ�JN?_0Pě�!��C���'����gd�>y,O��iU���"�heAPE˃w�h��w V�#���HĨl�����O�d�Oʓ�$$a�޶J�n̋��$��l
:(�InyB�'g�	�t�Iş|��_�u��_.TMVi���Z��������蟔��ٟh�':r�� �v>�[�/A9�0��A)�%|Lx��g��˓�?1(O��d�O���)7���^�����>@�ZHX��	/Ѻ�l�ݟ��I؟��	wy��שY�"�k�Ι���)�H �*�&� נٿ2�&�'��'*2�'l<��G�'��,b�����@�E����,A?��\l���d�IXyB/ʟ1'��������[C���!��i�~�L���_}�����	�~՜��x��ʕ�Ȇ%���Bɋ�Q��m�Ӧ�'�0� �fӨ<�O���OJn�W$p�gŏY$̹Hpʦ��ğ$ �,a��&���}�$"��N�@DA6��
�Д8q�AȦ���k�$�M����?A��R�x��'��T񴪕�!ܴ�0��n�6�P�o|��{���O��OT�?��	�V�L�B�kC�Ec��6��'H6��޴�?���?�����l׉'�2�'���E��~Y��^��.8SC�HǛ��|���6����$�O���C*,?�0x���5N:*�"$ɹ�-n�П��kG���?!����� �YB�oD�t-N���M�k�`��U����v�P�'���'�R]���5L��dM���AK�5r;|��Ǔ2/�xQN<����?yJ>���?iu�]�FŸi���α���j�p ��͓��D�O��d�O�ʓg��@02�l�!4��8sD.\���=`����$P����ПD'����П���%�>��/B���� %�*#gB���{}��'��'���.BK�dKM|��P�5�ib�!P����+���%q����'��'���'���'d�P$����0�1���1*^n�՟H�IFy�m�(�v�.�$�����O��0鈩�ա�֑ɰ�\�	�I�K��-�Ip�I~2����XAb!�J��V)Z��U�'��Y2l�"E�Op��O���4���{�%�z�h�P��PEto�ߟ��I/[��O�IMܧT��H�qN	* ��H;�jT'@Cp�nf�eZ�4�?��?���0��'9�G�6����˿<�6$�Տ�Z(�7�O�*G��4��&��˟,��i�(brvE��h�RS`�i��V��Mk��?��]en�j��x��'���Ob-�t�@!E4�L�2�@0 "A@��i��'c����)���Ob��O"]@!	ǹY�>�(Ď�/��t�Ԧ�Ŧ���B�ڱۋ}b�'�ɧ5��!$�4T�"$�&�a�� ���-*���<	��?������	<@��L��嘃a�2G�v4����T���h��}����l�ɚG06e��l�M6͇kĎd(�τ����?���?�.Oްy����|2Rk�=�ˡ��f�B��,���O`�O���O��)� �O� �@�]�Uop`�R��h�U��}B�'��V���ɳ~on�O\���C[�����u���°A��eĚ7M�OV�O��d�<���y�I1|�N�#�.S!4��:r�J`Y��i���'�剫}�� M|:���w���c+h�y��˖5?pEq,�d��'j��'��) V�����RB�(/U)ݴ��� �'�\Mm���i�O��
T~���j,���B��N�RO���Mk��p?Y���3X�0���"��.�0�)��ʦ� �Oӳ�M����?������x�'�!9wm�4.W�� ���
�a��g����	u���?Y����
6iz���q���O�� ����'���'��{S��'�?�O� ��A&ƺd�L��f���h��-�	�I�,��J|2�d£O�R�!D2O�ŪB�� d,�5���$.�h�� "O���C���6�J�N�R��F�'İŸ� �0a�9�g� k��� �f]3h�B��%ϒZ�vӇJZS��c��B|���d�U5w��Q@udX9|���J� Ąv����L�G�J�A��Y8�@���х1�6Yu/�^U�us���cF7J� ��5�*��d�Ѝ�F��$:L�an�.�Ԓ7hG�A�r���ES��q�'�RjنP��'x"�y��|Γ?a.H��q�,!,�h)�p<9�H��'�H0�G�W�wcP!��%-z���@�td��c�V$��񄃅S���'ɖ�C��jw��=
�fE#�\&PVj����t�	R����O1b]���Er��ݫ�A��D����'�D7-�(#^
c�J�AJp���86�Pm�Fy�	R#���?	(�p3d#�Ov丢�O�xm�\I�8w+#ˢ�?���3̑���Õ&I�s�e�<8�*�Dʧ=�2ZS��3�z���*4o�lѥO�I��o�=x�bY���\�v#}��%����D�쉎V�,���WM�D�r�'G�>���$st�19k�9�R�{dL!qC䉐:�΍j�ʜ�J�zUx�&����E{�O\$"=��"@#Yx���V-D�-��L�ą[1_��6�'��'�����!ҽF�r�';���y'�%1��e�vΐ�8�.�����u<�RKR=]����'$ap�[6�|���%pm��f��.�J�KR���NTD��$�kh���=.�\z��T�Sf�������°}#&4���Y�������ą�(�O�ўx���*]lh����n�x��j2D���%�
�2��EW���֮k�D�	��HO��OZ�z�rX�G��Q��h���� K��U�@l���?A���?�G��F��OP��c!>T��E\�a�iZ�2����#���>x*(a�����=Q'��V[�9y�
��/P�;Q�� mJ�V�X�d�����'�l[��+s�l�٢D
�Izg!�"�?����hO�� c��ޯ<Ȣ)�'�
�SH�Y�0D��b�cV1CB��� �]��$P��.�	��MC���Q�_�m�ß��I�,�U�fX�%�"� f�K�H��h�I�4�"�ɟ����|
�`���$�� 'ϩ�,��L�L�n0�W�,Ox�33��DE�h��-4_�Lɑ�#=o}�x����?a���򤀡V�1��G�'��ac$�@y�D�Ol�=�)§1�dQ�4(M�a
B}0"��93�j���N�6������2h5@��f�غ"S����ߡ�M��?�-�|t����OT�h��7v���@f���������O���H�8������d�|B*��U�ꉬpV=0���
�j4�ԝ>��j�E5�i�O>�� �D8�̎�\_��I�!�#��Pub:}�U��?A��?�����O��]ó��e�dѠJ��j�ļڎyR�'��y�̝�S�:�ٵ��<Qx��խ��0<�#�Ɉ]Gn���K�4`��v,I�ި�ݴ�?���?ِ��M"|����?Q���?�;G���rF˗�h��ٻ�>��@§��P�|�8�{- ��Щƿ��	:�ɾ=<��c2l��u��it�,gk�X�Pe�#��=�!ךwdܣ�f$��3<S �j5O�и���"NN0�ⵍ",7&�@�d�O�nZ柈R��F���>��?I��U�
S����ʶB�X��!���=�I>�d�\E�Q���hT�`j�F�<���c؛^\��|��
i��P������/g���hX�t�bV	>D��"� � `�@+Tj$u�NȨ�I)D��j���o�<(hV�N���ѩV�'D��H,'�  ���Ez�5C%D����._�'�[�I�fCx�#��>D�<�T�X���qG�ŪF}p��'>D�����#X|�4$�hL��D$(D������@k�`��/>o���w� D��q��(jүd��d�V?D�hX�S��rED���rUn=D��K�Ė�i�,�A�#A��Yx��<D��J�Y-�!�;-� �(.D�T�e	p݆<Y&�#��(jw�/D�\p�j�F܎U�a�ùg���3��9D���&�ۓ/�$1"��Ý���ZP3D�4�V�Q��lZrI�5W� l�41D��x2ϔ$>��$p�f��p�� *��:D�0:d�ؼ m�X8c"��D<D�L����0(����	�� ���<D��R���q��qM��<J���8D�ܳ���Kc�\� ��q��dm8D���Am� b��4y���=`C��d�04RŤ�=&�h��s�"C�ɪ(M������4d�͖�U�C�ɛj;��AE� 6��WA�>J)�C䉇S|��Y�$�/��y@ Z�dC�I(GՖ�
)��L��xv���B��8u��+�kR1���ħܯKV6B�I����!�&�|(C��+B�I�d�>��!��/,4�Ц��#<�C��1,\՚k��c�āZ�M�C�Ɍ^K�E��K�8=�U��$��y��C�ɯI&a�+�%��ђ4�fB��04H�cȪ_��1�6�C�	�C���L�〽!% *i㞰R��p<)6$C�R����,��`�h�](<Y!ϏM+�<yg �}!jX��E��t��ܘ4b/��k�B�)��d��JC�y�P�$�0O��k�)��'4��;"@Q']n�u� ��}�&]�
�'��Up�'�_�h�)�,$qmF��J��2� X<L�qO��%٥�Ђ#䖘�!��׶Px�"O���Ζ�Cw��ف!�,tj��[T�D81A���>�!j0�Z20�&�ܖksj<��� �8ፈ�.K�<�	�=1@�Yڶ�^�֘B��0\��%�О
��x�ȝ3q� ���<�I3R�� 	�̓�~��A�[�O��B�		^����>l<!3�!&/�B䉂 � �J
��r�ܠ�S( ��B��>Նܹ��g��6� �yҋ�������]���&�u�<��eȣA�H�V��z�؀��e�<a���Y��@i�E�=��E2��^�<B0���B#1�y6&Z�<y���N��1m_<F�Ay&�QW�<��[*y�
���8b�0=)$�R�<� �	 iH&D�R �_�,B,���"OF\ T��%-�!���#L1�#"O>�k)�	�I� ��l�z�"O�I��T�4�eJ֎ۙ���D�'IN�)8�	� ,����B� ix�!�R��cC�I�3�����GY�g�yfϗ")��:⋉�?��f��c�l�)�矠C�lL�X��� .��G��HƎ+D�hK&M� Kk�q)��cfL*�Gk�����Ba��,��M��H���q�X�U�ȑK1(0��&D�B����A%t���4u�H-!�iÒV�(�CcB�e�2عd��F�&B��$s�naD@
 D�))��A7y�"<�"G� 	fV6�- ]����J<u=&)��&� ��&ބ�y2G�	H�D ��!؀ע]�y�ę� EЦ�r�4���s�(�/%0cT80��ő:Szl�� <D���CY86|b!��4xp1��}��a�/F1"i�f�*.���i%�!�-E�7�4�ٵ��
�ꔇ��&c�d��W�ik�0ڰCV��X`A���<���2@j�	3t����v�^�;�+H�R��- R�Q�k1�UExr%��jmJ��I�:�������g~� �n�~1�L���,�y��[�+Ӳ����Tp	�`��ܼ�6%�~�ӺK�e[���5�͏V�܊V�a�y��f�y2��>*&P����A,O�(I�FՂ�yb
�k����?��큣��'��D��e�,�Y$��w�
"�Y��PR��2���K���L��{�V>�[uJ�=�Ƞ{���pG�Ի��f�N貃J94o�XB��ٱ:7�ܲ�R>��>�%�ƖU�۵e��J�#�ّxrH��m�%u�'��OK�>�M�u,��>�!k4��6�� e����]�2 h0��>vl�!aၧ�����N;�dB\c� ���$u�d:�J ,������IP�FƁ�?�փ�m� S͗,�9��$*��=�x������bǸ,�<ٕ扎"G�-I h�d�ģ��/��'.��2�Ɣ7�t������fKN8W��Mgg_zT|��ț�q�䄕O���R��ZFؐ�O�I���/&Qtۦ�J�'9d���i�H�`MW�-:��{�K
��L>yΟ�rD`}6��!�ճ	�ع�Gp}B�WqnL���_b 8 \?zl���d�
�8	y��?O/$�*D혜���������'���Q:$��k�$�U��.����vm��TD�����:5�����/.W�xJA�;�|¥ȫQ�j�!d^%6�&��s =E�0��%D_��?awcҿy���Q�'��0��;�~�:�����'6�FlҕC�-\h`��NB!�y��H�B#�`������ʕf�9OV�S�\�
��3X�T�(tlb����ʐh� �"�<��A͌ћ$]��:�Q��kOl#���苓�j�����`��2*N�9{�V�/ZЩ�v>�O��'R=�;�)O1���s�	/~hD�'9
�aG��W�hy�E/�^Ȝꐫ ?6�qO�%H"�
�urmc�i)Y)ΐ`JK�db�A�T�|��	2��hJ�@5EiJ)���9v�� Vʒ�Dj�QP���l�`�ac��!%qO�	Խ��;$�X`���ͪf9~�v�8 &�ym+LSԵ[�$׏��v�&�j��
C�I6=)�$ˢqܐ�#
y��c���'(9�Չ�lób�q��D�43�19��)h� t�w�[�
�y��	(; u�s�K�J��Hq4kv�ah��C1�t��b�+��@e��<��'k\�B��򄊎@Z�'{�\�D��3���⴯�x3���L>ᰧ�78���� ��%T*=�t!Lܓ13f���ND�S��(#%�(�j�7k��XjD�{���2+��#<�$E�(���[��L�~;Ph�`mN��R剖�Șu+���5�)�de^���1�cB�u���(�Λ
y�)�DiPC�&�Y#�Ϩ"i���I=P�&i(fŘ /����� S�]Zu�<��C��tqg��"֌�>牁&Q*B��Q;,�*A9�FI�����AlE*@;�N?	|�j���7R��B� }�$����A?���z'�	T�p�#�O��JQ?��$w�1�O�<���aF�_3� ӡ*t�a�r�|�
4��`�v���f��1�ݸ'y�������?��ذ&�BMNL�O�����'���$Z>�Gx���������)G-v���%[�`���?]_��p�j�H�S�)K(�5޴a�:8�a%��^�0�#+Y�v�b���X�R���Ui��8b��ʼdc|)	���Qf�@n�M���Df.�)b���W���g�A�/�^�ʅ�.�~�p�x����)Ƿ(�d��I7��Iۆ6��L���� @�q(FD�� �lj�{"MG����o�%E%�W�S��I�Hq���`,F^��1�U�'"��d�?MFb���ujp �I�2�����'��豈�"oZZ}�Sn�~	t-�ÇP�^�)�ŗ{ev8�Hǒ����O����	��!:��9�	�ʺE��b �0�0����#��!+���S�.Q&�!%Ï(��$�4	EwD�m�;���`��\�OP��t�Pt�S�\c?ppA�9?���	�gS���{�y�o6
���=�|2���8̤�gN'�hu�T�	?gpht���d.�3zq�� "I0��<LݰI�aQ�p(�,�$cY�%��R�)�ӂB�"��OB�a�"�M���Z�I�B+ě�~�gڷ7�(DE7���I2cSZ�9PAڈc��	 ��8Rw�$12�վC���:��OƐ����O�s��Z�J��'ٽCό8��-q5�P���T�=�Q��9�Ę�^\"QS�O6\��e*C|}�7#�#m/�ܚ�f������ fܖ���gVZ�4�Ѐ�[�
�l���� ��*#�� E���('8���fiPV M	��Z^�@
�&h�	�?tz5zŋ"i��I�R�P��W���)GD�{�,M)Y�3&@U;:Ѫ�p�H�wHҕ�'*�Ћ��$ό��xc*h�� �8L�AG�<UL-�3����sdB���fb)Fx��

|����A�~7��W�)J��ď^l��sܮp�쑰�g�'y��j����O�&l9�ɀ7y*��B��DН1}4}c�n��.�7/��8��cݭyƒ�YU H�AU�I�57�I�nE�`�T�nZú����yo�(�B��8��M*`,9}�b��<)d$
=(bܒ󮛒k�ȃ' �D̓>l���Fc���"����ş��'��2���jf�� �6��t�H��s�����Y�<xe�`䀨
>��KBЩ>L���'�G�O����+8O��
_d�}K�-�PLV�QȀ�1�,�nښ/ɾ����
�
�1Na>#>	�'ћ�U��(p����`8�|�Ra/�1O�!V�\�x�8dC �S�$d�n	�p<���r�L������U�qꚫ��Q��ҝR��)y�j�X���+�b��G-f��u⊋Z�D���Ի"o�	x⫗�1%
 �<y棇�q�
��A�>@�)�Ί`̓z[\�`��Q��ɡ �=j�Ԙ�?�C%�:Su��(�ɀ-&#���GPB���1��#���:����D�%��''bH��7 �n�az2�81q��C|o����
�FCވ���37�>%��n���X�}�z��,�N������Zm�d�=Y�`�����ɑNlx�� ͏%-q�,���F�����'���[rܧGt��/P��j�'ȄJ��+!�����Pۓ9� %�����mD�yٜ$p�Lt�����63�\#<�b���s�8K��<nh ]�1��A~b�D,\7Z-����gS� )q�A��'�.9
eʎ�8n�X���N��N�0��a�X	��b�.:I=SA�x�&���Ț6n2�A�l�U��������BӅ^^�0x����x�gYt��T�1��'^أǓ�>�y�J��
�|!
0n� 6�"w�����9�*�����(5��+S.�L[���p��<�^�Pۓ:���/���1E�H�gE�̐��1I� �#5?�%/�g���<����+�:T�]e��hp���R	Y������=�k L��q�-n��Y(%#�1U5�͓[�����1��2��ܨ�r���*1!X��A�h��ɍ7�Q>�	�)��`F)8��i�Ԍ~Ű�I 6�d���ɿ�@��S�iK��S�'�����.<��lQ$ƅl�I��_p�;Bo�`�.�b��'�p䃧��;d�S�\4�0�aW8:�����Q�}���CDk����4���� ��)_�Pu;Pn'&�!��9�p>���C�߁+$�b>����R�V
��܀Ҙ@#��_�_/(b��3�	�s @L8Ğ�KD��K7�^��#>aw�Ig�ّs���4i�p�C�?�kw���,�PiҀ@�8-�� D�xp��l��`�XE5ٕ���Xj`+�$+��(Ơَt��F��������
�x�JE�v�X,�y����s5Z�
W��;^�$7��y��
`�t(7�J���Cm\��y��f~�Y�'(C(C�<�Q���2�y�"�#"���˅'6�� ���yR��4���"���hq�T�y�B�?�� ��B�b�1p�!?�y��΃wڔ�T+Pz}!�n��yRd��|N��TM��&��32����y�	�1x���%%�XQ� n��y2GM�?dƽ8� 4J	�W��yrKE%tG��2 g� YƨqT�1�yb,�&���� ��F%;�y�O�7w%��r �Z�~U��+�_�y�]�q�����DD:@qSe�ٟ�y���<��P+1BN�;���'J=�yb�_�V�B��*O8����ą��y�"X5'}��C�m�0�޹����y� Aky2��q�L�+�J��(��y���b�ɐ Ā7r6�l�`.��yr.K�(�rį!g�:E���y
� 8��A4��p��ͨa�JQ�"O��0!�.R�x3c�����d"O2$����1@��Ua7!@�'�h %"O`��և	�gx*��m�����"O�QYW�]��D��u�.�`��v"O�(���&?*�+�e�G��9�"O��y��p,������)d�`���"O0��[�I0�,���,ζT"O��xn��@�4�:�އE��R�"O�9񶃒837\���΅�D̖�!�"O0�k�2K2��4.�>����"O.|��$�턔�K��"	��"O��	q�Z7.�T�{`��	T
4�W"O�ؚ0k";.4iA�\=B�\�ɢ"O�ܫr�@<<$��r#ـ8� �x�"O�!Z%%��|����S��E��\��"O���$��7�IFk�5D̎���"OT���F+<'�u"��ڮd��M��"OR×�Ԝ�U����G����AJY�<�2�P.ɸD{!�4&D�@I^o�<�4�^�,�B�+��L�?�����B�<�dΈpI�`��.K�/.&=�ψ@�<9�`��="�sq��y� -�G�q�<��K�7݂��DK[O"��F��o�<S��>q��X
4@V�蕈2b�h�<��h�c�
9�C�]PB�T��e�<���\�@��$�w%�u�䓷�F�<񐮋�A5DQ⏂�L�ZX{�@�<�5�D�f�%z5BJ�I��|�aj�B�<�N�4w���(+M厹�n�c�<і��	i��H��c��{� H�A*�j�<�G�D>�
ؑ� �<N^)��	j�<)F�\V��B�I¡]甅�r��k�<� l�
1�&Jm�vyJҁh�<��A�|s�)�"��2���d�<�w�B�������X�����\�<I3.�0T�|�I�,�C`@Q ΏU�<yAJ�EY�`MA'h�
U����O�<�aN�6b��HXp��#�♩w�N�<�u�T+_etY34	T.5� �3G�K�<�F�*bFLі@�!Ƥ�Ȣ��H�<q�e/?֖�[F�ܢ<��40��B�<q�i�:8d���*T)���B��~�<� ��"oX �N�"��T�ǡ]E�<qb��[���y� �"����/_K�<Q���#��вNȈ��qH	E�<�V*E#"y��Ë��I�<��AO�U�<I�.ܷ/-|���%Q��ږDO�<�t�ՅjX���ܷU�>�{�E�f�<W�So��I������ @C�X�<� �,1r QR�Kd��h��U�<i�k^�mTr�S	I(֜ s,�|�<�q�+5)�b���mX$T���s�<�d�X�mLu1���&0�-���{�<Y`F۵j0�j�/H�d�0��D�x�<�h��L��q��86�ب�"j�<Aĥɟ+0A;�� o*��!�d�<�q�S�R��U�# ��2Zh�bE�z�<)�*�RYp�LP.[yY��K�<Qs! ��"4�E#^17.e!DH�<���	1B�l��Ů��H������L�<P�����ӣ��		>���l�<aA/@�<�$ c2n˓} ��/�@�<W��6��5�#��GH�����<� �b��B1cJ��Ҳ� �4��b�"O"M� �H�IXތ����5v��(J�"O�1�
= |�а#�)i�P�"OIЅ��0l���$M�Y�r��"Ox	�	6O��@eŇ?�:�Q�"O�}3d��~b8���Ē&��1��"O��1��ĥ)�������g��p�"O�����߃3�t!LW�1	��"O�|A!bL�y�.�ö)�\��(�"O���a�Nwی̫�G�d����""OPY0�ӭf%Zd��*�`�2�"OJ#to�`t�\1pBN�4���[g"O���H&"�pu�v��X�J�h�"O6d��f+�Ԩ��A?m�4Ȓ"O��2t�ӝP�ZU;E����$(� "O�D��O��&�:��I�(����"O,�q(#@�n� ���3��9s"O�9�ߺD?d<�������]�3"O�TK'J����+@�;
�h9�`"O�m:�N_�w�9#�%�%U�i�w�~����Һ)5���E�2L`Xb��Z�n�!�D����	s�:BX����BR�c�!�dI�3h��H��sYp��X�x�!�DݦV���U"Y�^����vE͊e�!�$��Yu<�!��#��Q�MO#�!��u��eb�U�V���Hb�_e!��n1�0��&Y�� �,��:�!�W�.��@%͵|�Es4Y3H�!��Q��B$�l�¡�d��!�M2(�����)O8!@��W�:^�!���y%"x9�n"S[��qU���^�!�_���tE��kN
l���گV�!�ċ� {Q�([1�lepT��	�!�䋯��'���Y7�DZs�Hd!��QYQx�Xw��(Ҋ�qc/��!�@0|�����9V���C%�N��!�d�./za[0�}��!��lˏ$�!��Y�t�De�(ٗ��pᶫ�?=
!�N$4Ǿ�X)��}�bJ��C'���,����k2�� #D�%�ȓy� ){���L������'T"�"���s���"��?���"F�d�t��*3D�T*&�Иt>��O�MK`�Xu�2D�|�(Uv d�b�@�g���U	1D�H�5F�)�́R���*.3���*ړ�0|:�(L�K�,Tt�����#�pB�	�r�,8�	��
@��"ܵv��ʌ���O��0W ��z^:I��ǒb*���q"O�����! �̬e�@�,Z��@"O�h;�L�6M@(�хI/H��UW"O.�aD�E�����ҸQ� ��"O�(Ձ����dBJ��XH�"O8 ��㊆�Jq��H��0��"ONm�J�x8h�qc�{�@�� "Or���LV�L��5!��K�%���i@"OX�HcIZ"R)nAQN�
ǶLR�"Ob�r�o�*��\PC��6
����"O2)��E�G�|�ӫ��II�@�&"O��ED�v�*��L,���w"O �� ��:��j��z����"O�Xk�&���,��T�W.tp��"OrjB&P85�d�:ak�h@fL�"O�I�u�7�8(Bq�\2VI�q"O
Pbd�.<:^4���7.��%�"O� ��ᤉ38MR�$����*�X"O��(���Z"T��!�E9(��}�"O��R��_1��6��[�N�@"O�x��솩j��R�-����"O|͙�,b�)�%ŏ�\s~�K�"Oj��b�Ǻk䜼)���z{�tb"O�� �A�"#�́�ȇ,���I$"OV�;B��g���h��G!Ј��"O��c�	Veʁ�a��|�x���"O�aCoԵMt�˂�ͤd��mA�"O:����`Ů��vFH0U�����"O�´�^Zp���z�(;�"Ot�h�'�:{�9
���z�w"O�����	"��htę����A�"O&x�Qb�t���q��9}��H""O8t�`�! �9�@�N�.�r��"O��� �S-v�� �&�?	�v�Ò"O����n0Cmh�AS�V�w>^���"O|�F�?7�D�����gF]�"O`����/��	3��[�d��"O0P�C����� ��\�j��d��"O�Y�ĝ�Ӿ��vnĉ/�1�"OlD9��9���ђ��  r���"O�Qp/5mDkЧ��.����"O��y��٪XJ-�F¬s���7"O"�PE�(lP�3k�[Aʬ��"Oz����s� �Q���p0�X"O��JA Z��L�!r�ɟ!���"O��6�>x/|t��( Y|5��"Ox�I��X�Li��P�P�H�|k�"O|�gDG1`�@�!�I����@�"O&)�`'q1�	����%�L�v"O����d�5��.�r���F�>�����S�@�@Č'LF,M[ ���7	!�d+�`@��	�dKfհrN�'!�䒦3�P�2f�,�vt��j\�S�!�D�^qh�a�;O�$�'gK��IM�����EGmt�i��O;D��"6_-v=��b�^4�339D�p95n��Rt���t��h0ܢsM6D�8��[N<��#uf�W-�ͪ2k1D�X�eOBpX"(x�P1( ���0D�\S
B�0E�`�E.�&7��eI��0T���5�� ~CʘS6HЀ�(9��"O���S��	<��12��h�E	#�'Α�Jbȅ& 0��Ra�!1����0D��Su�̴q�ܐVE�:_���aAj3D�\8S�ݨr�h�H�%ڵ>�^� �H1D�`eÝ0&H�����;05Y$C1D��B��Q�e6��q�)/�Ż��"D�(��Z�TI�H=x���� ,D����M ��n�[�0!���!�a/D�(��L�*��e�:`HѠ2O9D�,yp�>h��peCO�D�Q�T�5D���c��m�±G� }'��44D��dC�MeL�#剭f���#g 2D�l�� ���������PF.D��K��R�y�ހj�kʨ$Er� a./D���sW�9QZ�$K }�F@!��)D��XT��3V�TmhRFJ4 ς�c�<D� �7�ʘN��ip�\=S5̨��>D�(A��	�<�xS���1����>D��r�혬Or��nK#h�@�	7D��*�$K5���a�ȼL�2�0�4D�� Չ���I6\}���[
�����"Oi����K��0�S�E�C�X�1�"Oԅ��=f� ј��_"q����"Op�ESh!��rRMC�U���H�"O(�MB�@<��:�k9)�  �"O~��b V�Uߦ�B�ȜB�$�$"OT!)��� �0� �(X�s\43�"O���GF�+, �F��2��2�"Ora+qb�9m8��ׅ�4����w"O������p�GoԞC�6�0�"O�cA�
>�n�2���e
R"O�! Ҥ��Lgh���Ѳ#J
922"O4�)��>?��Y�b�x0�Dsr"OT�'�H�W"������{p��F"O������%8Y����u>48F"O�L�bK^)(r�����PPr���"O*�B�˘|n0#��DJ`�bB"Ol�!���+�Q�"ՅH����"O�-�&�m�4�Q"O�8>dv"O�*#�dܚـ��'�H8�"O�93S��@JxCA��ƥca"O���͐�9�x�p���,1�L�1"Od������t��ఓ��b{��y�"O\�#���6lxCD���wg.1Z�"O*Y�ժW`��L炠LT�l�1"O�Q��O@�T~\8�c�Ƅ��#�"OƝ"�?[��rD��n��"OL�ju`��*�ǣu�b1Z�"O���C
�+t�l�"C���B`"O��+s�Z�h-��q��?J��4i�"O�p�1�[� � (ـ"O$��n��M�b��OO�Xd`La$"O��P&A�
[����.>^ܰ��"O�"�Z%l0��C�ϣNN��zV"O�(@s�ƾXl$4�6Β�f�e"O<��eI"6��3͆�L(,8��"O�;G��O�Z(�Q�\F�	Pg"Ojm����]�~ /t�qE��e�!�dZ4 �(��Gȗ6M�fe�p��b�!��A�y/��g$ȽS��xgM+�!�P9 P$��v���"$�91��p�!��W�_9�|��×�?7䛵��0�!�d�=���P�|/&K4K]�"�!���9b�\�W`�,&s�J@/S�!�oԊ�q��O�4�u��T!�䊻	������/��M�T`\ WO!��Ҋ,����k� a���Z6R�R�!�DO�d�ꙣpc�%�~Q�*�F�!�D�<����)�(q�:�'��!�!�d������&H}�a����$�!�$�%w.D
s��$%Tf`ȥɉ"�!�DĴ&z�M�xIz�3��@�zR!��%@�vd c808��QF"��y[!�Q�D$�B��,n�n1���E7mO!�$�u8@���&Q�.��p���kF!򄑏MEN�Ҵ�!=�b���`W�!9!��̸+w��Z�o��_���U&y�!�d��"�ˢ��J�9�DI#s�!򤌎GA�Li�φ1B�Ed,[!�$ԝ�,zǊJ�*#�\�CL	.[�!�L��С "�a-*�@��X{�!���u��9��PI�*ek!�dɌa��|Ԫ�	jM�A��>�!��[���b$�!�� �CL�*!�� ʤ��M��$L�)PX�m� 8	�"O��p%�6Mڶ|� .�0<�.��"O�I�A��(氐W'k����"O4�� ��>| l����R�^�@T"O|���.u� ���5;�M�a"O�8i��޵[!~��d��y�v�ҥ"O�t!]�bӪl�TI��>ڎ`�e"Or���LL�H�P��j���T"O0���L\,^�9�@�տ:��p�r"O����m�5:���$��e�v� �"O�����9��xS$"�"Z���
"O�Њ4��'���@`&��b����"O �[Jԓ|�xD��D�w�plI"ODD��)����0�D�j��ط"O$���]�%`���~YP`�b"Of� '�X�d	P�!D&hc��ɰN0D��;#ϺI�=�Sa�<���6�9D���Ŋ#�4ݸq �u�����9D�t`���?_4\�ꀷ
�ε4�7D�d��j��?&�8���R�}]f�#�o3D��a��ȡN(����l�`�i��2D�r� ^
I����a/Z�}�<iTk1D�|z�!O�vT�ъAA˯ml
��C��
`�4,� $(oxP�#�@���B�	�r(�4�s�ȣ3�x]3��HM�B��	kt�����N�`z�/�MyBB�I}�5�䉙�u=�c�(S�B䉶p��SPmU��9"s�Vd�C��A� a;ᅏeXdy��?G.B䉔{ \u*����Z�{�'�#� B�I�>��"��͍FG�!�k̸^5�C���kTE�ogځ�@e��H��C�I ��P�_�]A�T;�˗O[VC䉏F��Q(�

Q�|��	�'��B�	3mHnmk�na
-��fՎ@�C�I��Li�dɋ�]<�R�Э�B䉉R�Y6ɀ	�(Q ��RM�.C�ɢ\��pM��:�
5��00z�B�%H�$|�/�1-�(��e ���C�	��X�s�j�/�t'� �D@�B��*t�(���ճ����Ph_�:0B�	t>E�� R��H�%�.&�C�	�77���V&`Nz��L��tF\C�I���i3ց�v�`�cf�J"�B䉋b���NX�y�2蔱!�DC�	�#���(�"� A��\"cᔩ<z�B�ɺr�P��e�Ǟ�"��j,�B�+d{ 5��'s��h衉�\�NB�I/\r��hE�x�U�S�]\*B䉺h��	�� �H��t�O�ge�C�ɔg:AQ��4?z�*��\��C�k �Mb���B%z��5��C�	&t欥�V���R��`� h]�jpC�I
L����G��	�A8��r�B�I�:`LA��(;���Į��C䉗qa`���%�Oj��@�  I6�C�ɱm?~�k2D֑7f��T��%&��C�I�+�bP�v�RLA4ap3%��X��B�	�%)�i��h�]����ةhf�B�	%*Ѐ%P��A����*f��B�	6,�J%��%��q��ÇK
/A��C�	�vu`�B�*Uh2���b���!g&C�	+%�,}��-Y "���I�/�]�B�ɡj>�1p�A8F��H��\3ӄC�)� ����j����`!dY3m����*O왺�MQ-��+QZ3E@�|��'��v$ƭ��x�q��!��m��'ߺi&�(��y1ɒ�{����'D�8�$��c���0(�q4L���'(�D@��ͿC�x�'�+l%��	�'
�+�I.-��]v�ůw���'`�%�b��2��5�H�GV͑�'v$L�t���X�k��h*p��'��l q-��%�^����	Sl����'�tC��H�Q.��a&���N��i(O$���̓x>��(�9)^�i`NԲ0�!�d����#'EʲLF�Z1螑�!��#+��i�)%��IB逐�!��NP5N�	B�'M�uq�S�@�!�W,R�H�� :[�B��d�51k!�L�kS�Ƅ�� 3;#XAR1�+D���
T�8�X�G:d@�����5ړ�0|��DA�(.��H��(S�\y{��\f�<yRJ-S��}ׁ��G�<��t�JJ�<!����nG���G��hϊ	G�N�<��kʞ�v��T�K�n�ـf.M�<���2Uu���7��B��8QN�F�<�b���L�|5 �A��?�0|�q�C�<!D��3�^JA�Fi�D�z� �j�T��9��RJ��Y��H�k^uՄ%D����Dy~N=Q$�E*R�&1�f/9D����kѠI��		�m�����Sb�p�<��'SR�@SO�K�5��Tm�<1�cP�1y"�i��ݨN���I�DHf�<��e���5��4(�IfI\M�<95Ǘ�nޠQ2A_b�X��a�<!͢\� q��D�1���WGQ�����8>/DRf��i?�Q96BI�}dD�ȓ5`�b$,/��(�gΦ̈����2�ɵ}b�m�t�]�ږ�ȓ/N4�1  &d I�b��*�^)�ȓWr���.^V��qn�o&���>��D�D���m@��rFQ"J�E{b�'��(!��5�`��h�vW�+	���y�#�$ke��2fϴ�h2� �yr�kڽ�g䈰Z^N�p��Y��y��?���PÃ�;DB���UC3�y�A�-
Y��@��G�7�z������y(Ɨ����(>!%����$ 7�yR�++�l�eIJ;��Tꖥ�y"ko��L�bǝ�~{���ǘ%��?��Y�����"Cv1l�R'L�6���y��xRA��g0*�
�蔫j��=�3'T�y�Ͼ+��Y���=e�đ3L��y85f x��8M4Qg�?�yr%����5��Z�J�\���a���y�ܥ.�h��\�?�Ȥ�3
����2�S�Oa
���wL6��ʏ?W�ey�'!��#G��8����bo�����^'�!�䜯s#Ni�&!�33m\L�� H�Q!��2�^]a@+G�vg8U��ϛ��!�d@>G�Dy�pNZ�(���� �!�_9^��	��!-6��	Г�K	u*!�ѻ~�����S:�TT��b�<d���)�'p�Jq	��2*���#�
څ��'Y���*�f�� @�/I���(x�'��Yh�JU�P�F����D<$ƚ,��'B��x��	�77z��d��'\=��� :rqi]%[������\�*�1"O����Wf��R��*{�6��0"OBЈ���mi�ep! +t�3�"O�%̔j�*�3�E�����y��'(�$V�$l38oe$vGm2�M����t�T�<�޸"#f=]~y���"D�$�Mǯ=�(�e�3W��aV�-D������$� R��F�lgz����=D���E�1_bX�aF��t��88t�:D��@FY�s�$ՠ�m�O�a -D�,*�.I) �2��⁚,Ĺ3C�&��'��|��O^�� h��1(`�4�:�ZQ�"O���aH�	����؂Ԭ���"ON0q���P��y�-���Y��"O�X�մUm�샱+Z
5�"O6\�⢄�UuJU����$=*�"OT�k7O�j�����R�e ��3�'���ܓ0@@��
yę�!]$��O��$;�g?16�"*j�L*�[�i'��xA�q�<ဤ�-^
�K�Jн}����k�<i��(oC��)qG�=\O|�R��c�<Vi͜4��P�=Aѐ�J�nCi�<�A�ܲH��@U���h�
ezu�i�<��O�F}�@"��z�*Q}�<�E��g���d�M
�#�x��0=�S�В����a>x`�8���Yy��'O`q%���\h���(���
�'��P��' Rh��.Cd*�
�'B�[g10 �<#���6�RE��'=�AHK�K�J�
P�^!11BX�'�Z�{�@	�e5�t�G�U�0Qԑ�����C(s��	
�Ś/��j���0]��'��{�L�E6�a�RK�a��يp�ܱ)�!�D́!(Zɒ��v��4y�CR
17!��{���I�$�x�������:y	!�Rf���U������GJ��!�Mm2b(8�C��Y��	/;�!��֭L�x�� CՎ;3��s(�;k��}����aţԏ��a�Ǣ;��9�l�<!	�-�,��&��_�]�@S��5�ȓ[rf�����W�>�EC�#0\ꬅȓ@e�3���Zm6);��_/�Ʉ�G�*`Ӆ�ۉ<>�p��Q}�a�ȓ\$2$;q&Ǹo���� ��*̆�.��MK�_'�雳uL��:J<��@��*_a�`fA�d��$�����R�E^�f�&����͆o~���ȓ\ϖ S#h>�Z�� Aʙ5��d��\'�d�����F�����<#^d��,��8I�O�}�(����a��$�ȓl{Lh�l	�$�Z$�s-��q����*Mn�xV� |HH2W��
t��$�ȓa��դD1/������	M+8i��,2,I ��
eF��ȇ�k���ȓ?z��k�OG��V`E`B�nc��������a�ˢj��x��ʓ�2��-�ȓUV�!L�bd	�#� T��<���p�� ��@���CA.�Q��0�ȓP����fYA��i#��C�=z��#@*�ك�($���"V��7O���ȓ5�`�t��*)f�� h��7>�E�ȓt��u2��ޠ��l�Ʉ�9�ظ��-^��3�@�_,�3�P�tN����r��P�����Y�Q-<b ����S�? .<����\��Fg�O�DH�W"O`+��Px������	�@�'�ў"~z�Ӈ!j����T/J�́�ơT���x�b��6�ĵ3Q"$P���RP �!�䁗9ᖁY�BX,%{Vл�J��t�!��G5L	B�х(�Ph�d
�p�!�+I��#R�֊�(�srdA�w!�d	,�h9�R<B��L�Κ^Z!�ĝ#��˥T�2~��J�"�8��'cў�>e��خ3=Z�:�aO�%�	)�-4�O���u<4]��*�) xԀ���u� ��0?�!�
�9�|0�bI�`�	���F�<��Q�b�U����+G(�H�$]y�<���\�k�Y3я�$s��T�W�Ms�<y���oЪ���H�f�Pq0n�<���s��JA�m9jh��"O�	��
k?��A���?VN��	����L +�R��F
Z�9]vi%��N�!�D[�X��	�,��sB4#�J;�!��,V2$���;�i�o!�@J.�d���1`� �  	�W^!��ބJ�(�����=_t�U��({>��P��(� �K�㗡,{@�9S�H�>���V��0�IŖ	�6I�BXV3�!�����q�\�ȓ�X+#ʓ�b֢Y���lɜ��'�a~�dL- Ȃ:���&�jpZ��H��y��_�Y��C�"��^l��B��y�IN��,�2�,ܜ�q�[��y���1|Yk�/]1u�2-�  X;�yR(Q(Pb��B�� Y��C����d(�S�O^��Q ������!#�hȀ
�'�Y�Ŏ����IGa�#X�}��'�R ��H�@��逖S���
�'�6)1�##<|~pL��G=��
�'c��H�йbq�<zSC�56���b�'��p%�]���x�U�+���	�r�|�ᓯaaF��e�Y:_����m\�a���0�Trg��0ڥ�[�O*��R�3D��'�ִ��+D�ĆA~��&i-D�|1�⒇U��H��ĒQ���"�(D�|�0��F��m�B+A�C�P���'D�>��ᗯ�6��M�%��(n�C�I�w�F1Z2F�֘(�(0gU�C�3�N`�#_̀�1v�H"58�$!�S�O'�k��>0h)�%�������"O����(P�(���j�%�q&��'"O���W"~Ђ��Dͷ(���W"O�I�w$���x�@���Ӹ>L�B䉷q�XT�e�P8_��YSf��Mq�B䉠�^����� d��Y�@پ"��B��3C*p���	|�W'0��q�ȓB��H�%$l�" ��A�M��=
��+��}NRi�ec��E�(�ȓ ���ŭpNf�*�%� ���ȓ-(�����}�tjW���mB��V/NE�D'��<� 5����mfj݄ȓ��1�j�7�̼��f_�>�tфȓJ�����L\�԰��MTy��-�<8���&�z�2C(��N^r��ȓ}��03a�ƣi��g�ߏu����IR5+F��c�d9R���dI�ȓ	�p�D�*
,�b� 0�(I��hN,	v��'(⠻kU�0�ȓF�4�6���Na�c�� �X��S�? �ف�m�%9X��� M���(��1"O��,L��8LIfK0�X�3�"O,�¥N�)T��� �M�v�BA�d"O$lS�e�����|Nލ"4"O��[�e�(ڑ��V�B�M*E"O��A����d�>�x%I>=:v�S"Oa��C��i���'m̽,@u�B"O`p��KN�BP�����D�W"O�zbL� �3�cT�=��"O��[&��D����R�ܮ*y���5"O|Q�jJ"��̩�@���a�"On�! �Z�	�V]��a�g���"OT4��	Ļ���f!ύJ�"��'"O��4(�2����v�V2m��Q"O
�F�6�|�1�0'��uC&"O���ĢG�B�ؕ0�bAd�q"O|m`P	�?m�����	�$Ez�QT"OB���-"�xvg��B����"O���BX� ��=a�E�7l�H �"O��k!���vOx�b�������4"Of��"��TL:P�N,?����"Oi�t�"d�s��.85�@h"O0��(�&0�hƺ,$ �f"O�YYS�L�fWv$����6��"O xCc��ix��p&�"��h�"O����Gږo"�K��F�"��S"O��d4M4�cg��m����`"Of�+��M�i�3/έ%�0L[@"O���ѡ��wR|T�@B�����"O^���N	Bx�aO����"O�D�C�ش!Ӟܨ0�B�\p67�!D��"�'8E���q΅�z��\s�c?D�0Rg�=x}��h��а1��"0��C�I�<$|H*��A2�0�A����C�ɺm]����')�ղV@0}&�B䉫K^�<b�L��X�#Mq�B�I?DA)p��(?��4��sg�B�I-]�"%qrOZ�H!�U��$L?C��B䉽{�p�T]?Yc��@�Șf{�B�p�N���[�G3N�y1�E6)�B�	oE�РgoS=�ꄸçY~��B䉭i� m�FM7X�%�%L]2��C�I5�y#tՋ�)�V� C��B�	
<v��E-A�t�Q�� !j[�B�ɗ%� y��V�DeI�.����"O�-�T���\T��)�&G�tL@�"Ox�z�v p�P���);�֔H�"O�=k�-M��|!��*-P��]�e"O
�ЄEM���Q!�GR�4m��"OD ��V�,��Y�O�� �TY"OQ 򤕾[ d�Bo��R(�P"O���aj��-��24��Q�.H�T"O�e�$aI�*
1�F��"B�ŋ1"O䅺7��s�`K��T�[B��#"O��3�F�=	��ԉ�'ے�"O�<��S��v�z��*M�� ��"O��ar�B0'q�h�����(���"O
i8E�I$S��	��g�"N��)�"O8�s�E<K���3�H�(:L��"O>�S��Հ8j�Q�01�M�u"ODh�TXȅ�vc�%*�9a"O�h%1D5(娃�1)hx��"Oh �3�/z�p-��y8ڔ`�"O�Y�B�d[�lq�e_�$��
�"O� :�ȧI�<m*]�5�76{v��"O�-��d�81Q띃l�lYBR"O���`B9Z6�-C����cq�I�"O�djuE
�<%&�9�(�Kh�V"OL�ғ���urRx(�b�\���
�"O��ce	ʰ�p�@C��`&"Ox!2�Z�$1 ݑrG�$%��{R"O�[���&wmV��vɴ��UG"O�tzac��{A��.9b���4"O�`P��3�|$;b�� h:��f"O�=�7)�d�������c �U	�"O�!�1,ʬ�J9K�i͟/�~�`"O)��o׎���(w�b�B�"O<I!rCHd�Ix�#¡l�ʨ+�"O�	ff̉;���:�m�N�+�"O����A�)��j�09��!e"O���v�W;S+�=��A�l�:4��"O�y!/8P�������\ S�"O29�焤n��t���e�(��e"Oh���M�R2%[E�^�m�:�G"O�<Z�kW��<�AG�mR8��"O�i�ޡ`��u1!�,[>Y��"OV�SRÀ�:��TPad�#=��p�"O}ۢn#>��PQD�<�콹r"O&eIf�_9rXd��"N�[vJ��"Of�!e� !NԊs��&J|*��!"O�]��Ya�e��;�t=� "Or�xb'Z�
��h
��O�`=��"OV�zŬ
�V��)���9�J4�Q"O8M���	3C�����,Ӗcl����"Opœ���;q�lɦ�S�<z��"OX�*@)P�dS��Z�L[c���Q"O.a�U�S$D�j����V5J�"O�l:�(F�� `"��I^��t"OXxr�'7MFNYb@C6B>I�p"O�<yDI�J(�)SϏ-��"O�)��	%'l��&N�4]�2H�"O�q��ݿv�x��jF�}�P�""O>1���<]�>T��)�mkԡ�"O�H`$'��0�<̓�(D	�f��"O��v�Aֺ-8�"��{�U�s"O�	ȅΝ	*�ȴbU�na���"O���A�5xPi�`�G-[=��3e"O"y�a))��8��1o'p"O��*����V�%)\�*&"O��Q
I;FF�
��Fy30-� "Ozr7&��q�X ��&J�O)�%�@"O�m�􋀺�uz��4<����"OB4�b΃�qh������$I���%"O��&��/Z��4�4Fi=�5;�"O6h��7zf�\)�/
+\+�\�"O�ڦo�V֮�x��(�ij�"Oxl����_Rt�g��s,��6"O> �@�Ǳ"���ǐ��D��G"O� P�f�|�"�F�S�:���3�"O�A����Dy
�ɴF�j�NY(�"O�ٶE��EԠkq�:o�J�q�"O���󻤈y�! d�-M(�y���#9R�4�2"��N�Zd`��қ�y/��QI�P-L��X4���y�d�!_���:b�הI:�d�_�y��\=>LK0���Bo>0��)��yr�*q�5y�2e�@���,�y2�ݲuB�0���12�H,�݆�y
� ���ӭN�����T�˝(8�c�"Oz���*B��,T�� ��|���R�"O�X@Qȗ�u�!��!�!�ĸ��"O��0/�������9u��i1"Ol9��E[�2��y����G�l�"OL��T�!Ȩ�����b�<��b"Oб!aG�u0��,�G�lyyg"O�C2�Ӯ7Da�aƍ�p���qT"OV��Uf^�`��D��!S5�@s "O�$P���:(�����K�.�C�"OX� U� K���P��ޖ~C&X@"Orx�Cg\0C��������1"O�����#��Y�eD|�  �6"O҉3��>�Z�'T�F�"O�I�uf�N=� �S%c� ���"O4ԋ%������Dm�F�d	A"O�0Q�#D�S��O2ޘ�"O�zf��zΖt���̙a�eR�"Oڵ8�K��Y��+��|�P&"O�X�6e�"V���P$�`���"O0�3�"A�D���ߥXr��!"O��x�?c�ҍ��lSLT|��V"OڭRa-�&28�� @J�:�"O��@�	Nd�h9�jN"d5sS"O����	Գ!Iu2����|b�"ON�H�WW�i�)�S����"O���᪟�X�����)�
ў "O0=����bB� �犰9��6"OZ-:U牻7[�I:�� �z���7"ONX�D�Q�Z�V��+V9ʘ�W"Ovi��_�?.
m �%S�=&rI	"Ox�rp�2/��S�n�!
�x� "O�0"�N��di���/�#�	�c"O�"��;P��M�c�G)7�6iP�"O���د}�xq	F�ˋ9�F��"O����I�:��2�0��=R#"O�`�#- 
f=��M!����"Ol@���7y���O�$��{�"Opٵ�Z�jW*�i���tR!t"O0Ш�n�4�D���P�X&"OB\ �$H�O���X%̹SM�Lж"O��8�N�1~�mIE��,TVPU!"O�A�R/��'*"h�\Ｙ��"Oz���E�I�V {����n���G"O�4!�!�5�����S�N<�0"O�����ZT�V�h�+	,���&"O� 
��,f��d�'	��l��d!'"O�X1�(Ω�b����ȔQ�
�`�"O��W#�2�pU����| p�"O@i�s�̭��(��,�{���K�"O
�tLӧ\x�
���l~p��b"O��б�N[���1��|ڮxA#"O���[���� ��b}S"O�7
Mm�
�8�Ėv�
��"O�@ �nۀD����䂾}��	r""OjM�� �(k�m��b�!�ȸSw"OH�q���3\n�����i��t;`"O0��u�	�Vj�K�J�1g�NiB�"Ov镫��B����#
�˴H��"O@)�F.C�S�a��(��(�9J�"O�P`�-ôg��=Iw� �p��"O���v(��o���!�gE
n��Y`�"O(��a��.��� �?�D5r4"OBIP�,͗:����k�1ɖ,X�"O� 0}�`�\�4�����i�b,�d"O8-�/� o�r8Vh�
}�lr�"O�l�:�nx�� � oh|��"O$���F7Xa��j�o٭-�2m��"O����POآ,�1Owj� �f"OhQ��nN��L�N��8c���G"O((c��	�@o�D5.&�|5r"O�}(� �:�Ф����/����"OFT�aΘ�~4��� �4��"O�8Jᩖ1'ƺ�b!d�8$�r@�$"O*\{��	�,�0�$�s�T�4"OA!d������ �N�$Nā�"O2l2���1T�(�z�Hˠ59؝��"Od�����R(��Ң�Ԅ4��"�"O܈bC�<d,��;@�W��D`�"O>4�Cյ5qt��2�#Ḍ`T"O�|x�C�����SaN4��@X"O|쩡*X�m#�DSrG�F˞9�$"OB�)���Y"���G�N� �H�"O��* B��TR�p%T�t89
�'��=ѶR�a[�i0E��:Q��'
����i*k4��5iSa[�'JY��.�-zRe���ۧ
��M�
�'���COF
萨Ğ|�\Ղ
�'ML�3�����닑zs���	�'�8L��h^�{D�(����c����'��i��&	�	�4��,�����'~��A��B���H�ǋ:%O0�P�'i�5ʔ�&w�Pʵ/J�1��(�'�`�ٕ	�!Հ5�q�Q�]����'G6���/0�HB���j@���'�$0
fK��+��1�ώil|��'�by�C�L�{�A�0
[�p�-s�'Y�%���^,l�{M=�$U��' �Z⌉ZG���q��h3.�	�'���[dc�/,!ny�!�P���A�'bT��i��D�Ht�ڧC��c�'��h;BF�q����Ӥ�;���b�'lQ���-cܰ�G".8��9	�'U2T�wJU�~�$l��`�4}�x��'t��IC�ܴ��AjZteV�1�'��\+�@	��*��_"f���'[��Cp@T�,R�,��#�"Fv`�
�'����M�++�MPդ��-c��:	�'a���4�˞�*-Ig�:7���(�'x���vղPr)����5V�x(�'��y�Ț'e���u�?%c��
�'�,��_�%��Y�t�ӹ2��	�'�V������kT����ʓs:����ک}N`x�k��E`ه� <^���jR8wv�2! [	<7�D�ȓU.pa�EeI7$�ڽdT�L�bP��L���Eć9�ބ� ���m�����9_`D[V��sw\M���pu���xT�c�H	�N(Kv�� z���
�����(2f�����u�чȓ���A��*e< �
��	
(��k��	ɢ�ˮb�րrpJ݋uF���<��"iX=1b��0�24a�������)rP���i�?dr��ȓ~��,Pe�?ٶM�ť44� ��bkP<� !@=�87.C�Po�ą�
��h��*�5��X#�Ϋ'>�ȓ���Ə�?"�F@�ZY�tĄ�S�? -���
�/7��3 V>����"OF Z���?6�ZQR@��챰`"O�}[�\�,��� ��/�\�t"O�(�Ad�f6h�vnV=��=��"OR����l^6	��HA�>��3"O���G:s�I��L�r�:�aT"O���W�4��Xb�؁J�
�p�"OdL�`��QU�Xi�
GS�6A�t"O~�h�O6��-%�Zr���k�"Ou�aL"<�`+Y����t�<a�䆠W@�8�\�%�ꨪf�Y~�<��偮Q��� ��"F�ݒ0�Tt�<����,D�`�¢ÛZj��
�!e�<1gNN�D2J1��.��$;Q*��u�<av _� �n�Pr�Z�_��=J�M�|�<��B\�&��ѓ2�(K�b�� �u�<1��Y����'P&q��!H�n�<�����^(�Eͪ�=)'��g�<��Ӻn���P���� ���hY�<� ��#J�|@���'Zs8,�r
T{�<Y��C�6�*�GeD'.=hC�}�<I�FY6)������.�@�(��SO�<�w@�>�%��c�]�5`���I�<!A	M�b��V	3���i�E�<��@�U)���KѠ�&h�rf@�<����8�:0��*��I��]*�(L~�<���<$­)*w�dP��.JV�<��oI�d*��r���|B�KL�<�"ń"I��B"	E�[Bڌ�vf�`�<�w�0B+����~Ŕ"���G�<i��۰o���
@D�b6�x��GB�<A�IV,Ă�9E��O7��{��\A�<���?<�i��/�s���҇�A�<�$��.@'�-�P��R�,P���RR�<a�f��<�|�%�W�#� !��W�<Q��ǝ�H��D�7e*�WbBP�<1�G˒j��A��*�|�"|Z���c�<�7�!]�r�N�R�8�а��J�<	�"p�v�(�L�m<kD�SE�<aFFv�~!�6��I�V����
C�<��	G e��ip�CZ�T���CT�B�<�q��\G>hs�#Z/˚�@TB�<�1��MҨdif�ݪ<��hv�D�<��4oށ���Q&n{�@X��z�<� c�f�� � �H#0j�:D�w�<ᠲ�,X��̀9�L���G�0�>B�O�q0!��:X�0f���[��C��>�pn��9�$��V�2B�\��ȓw���QÛ�K:J�1É0;�~��ȓl(p�j�,�\Lm�ċ�-]^��ȓa�����@�H��m�`��\J<|�ȓ#�n�J%H�?��Y(�〣.�~-�ȓ4E��� 8N�jHH�a��P�ȓ*���{B�,�"�B �̅@���?X����ʦN��<�$�M�@��}�ȓ8^
�҇*\�W��H��} �x��=b�%��{ւx8t%�aUv��ȓF�Xd��G$=*|�C�
�at*��ȓ2b���֦ɱ8q���d�doL��=z\=J"
�@~rB�Ńub�ȓ��bE�Q+v\����=-�L���Z����!����� �3}�Ȇ�q�Tk@hǛg�H19�!ٷ+��l��A��y"�U08����#��0O�6��S�? ]��E�k�6A�aȦc"dl�d"OBL�ȭK�����M �3�"OґZ���-����������"O 4�u+$&��dESv�� "O����|j���������u"O�S���&�(@�$v���0U"O|��C���^]"U ��D<-�@e�v"Obt����"�6bv��G�ʥ`"O�0��MÝJ��rI��l����"Od��B��lb��nD,�z��"O����LD)%�h�b�ڂ8�&��"O��e��L	�Q汲�!bCi�<�3F�)e��!���-"؎\�0$d�<���&]w\��4��l�e���b�<q��_:��h4�T�o�j)"��W�<�u�V>+����'�;gX�y௓R�<ѳNA�Z��U���Ĝ	6Th�G�<�a��1{j��GK�-?l���BCA�<����eҙ�I�\jl �z�<���َj�4��C,\ Zk��#��s�<ivA�W���10酸"�|D�U�<�T��8�2�閇¶]���m�S�<y�h;F�xPe	zEh= рZ�<a�Y�uZ�]��S��
w�V�<Q0"�,T��1c��
uM��F�Q�<��	C4��hq���H�,��F)XP�<!F�K�:$4�l�>%(̐*&��F�<�Q >~H�f��=P��0�6\D�<q��§v����6�l�Yfa��<�V�J�p��-���O6u����|�<�v���Y�d%�H��l��D�<)'�T:��iʮK�
��E���<��J[7UԲyq�k^+r��EVF�<9��O�g� :Ц�U�|��D�E�<�kL�S�ΐ�s�Qq�z�puj�D�<�v ��1!d=����/�����Ng�<���[����35 =��'A}�<I��{�(��ԫI�E5`���Hz�<��K�5(B�+�nրg�ʄiY@�<�"�X&ƹ�H=Jz�s��z�<QT	S�3��-�膺H눤q��^�<i�� $꼙p�6n�^�8u��Y�<�«Ќ_�
�%�[�b�����'�S�<��R�f�t��e-_��\���Q�<9���!�������'T�峁GJT�<i�H��PD��ʔ�]�\'X	K�L@Z�<%�̗bF5 ���>Ax f�U�<i��?�T��Qs<R�s@��F�<��l9^%���I�	��+0L�Z�<�� Ŭ@e4��c���v�Ƅ���[�<��Y�v8B�a0�Y:d$Fh#��ZW�<y���[`��868[��z�<i�,��f��K'n1^'�	a��r�<���?�hK'�E) 7R��a͒q�<�S�եN��-�%G���D��m�<����@]�Y��HP"	��L���]c�<��ᄢd�>4��i��^L���d�<aqd޹ފQG�ٖ
��8c�a�<���<5�j�b��a;4�b �\�<��̎wD�!���l	0�"�T�<�q�B�*��1�
79�V�� �Q�<����O�L��@JPL��ip'Es�<q�j��`^51�ғk�ܥ�Qm�<��+I��Л���'4���Oo�<� >���EO�%��"��M� xӴ"OT�a�2'XRܻ�U�K�p@�"O�-��N�6���#Юވ9���"O.�*��3�JT Q��T���q5"OH!@āهR�`�S��ҫ=��1��"Ov�b�Z�z.���
�)d�$��d"O��8a-צ��a��:o�Z�K�"OB0K�ID�LؠT��A�*V���C�"O9��ܞB��+�oʸa��Q;B"O� �fŅ#�b�2 X�.���sE"O�9�	65�\T�ծ�9�(���"O��]%$�Du�S��?j�!�"O�E��%�yQ\�Ó���]��"O��Y��[�,���*ROY�b�LɈ"O� �D�ŉR�JP��8Al���&"On����]Zj���	d���C"OJ%���� �LI6��hU�"O��#��ܧ{���\�dl��q"O�P�aN�B;FD����*"THr�"O�mk���|�Ɛ��L�Q�jX��"O�i #(�c�.��ލ?����q"O���5*�]?�ءf��4�(a"O�A�#i$h2Bd��	�^ʄ@ "Ov����{�X��Ƅ�=RT�``�"O.`�G�L��x��7Ê�FCd`J#"Ot��� �*,����=0ZE"O1@5a�[��*�B�<N5���"O�P�B�\-�ԡ)c�K+.@h�"O΍rW�V��܉���9
.�qf"O�0c� 'W_<�� ��nx ��"O�\���ب��A���ȋmn&IP"O "*E�0"�*cG:��0�d"OV�p��H�Rq��ˀ��� ��"O�|24�4�fXxvf� N����"O�1͏�X�v�r7���jXqb"O�⇣�/x����AѤ/�Ti�"OX\�g�!����!�Bf@�7"O`�x�eO�&���P�L�qd�}8�"O��Ad(Α8paawl�#af��D"OhY[��<R���a�vI0�""O<\�����d�q�� =�`�"O�Un!B=q�N�	`4:eb�"O2B��>�@����$||!�"O���Si�J~H�iǌř[��z�"O�]3%��$Gu �1ׄG�O�WLw�<�Wh\E�~]i5�͒P�~#�Up�<A��_0jJĳ�M��ZsX�
b��h�<�*Ψ,>4�b�l5�j�
���i�<9���:�J�3$�V�%A(����O�<��'/jZ�Y�F	LH>���E�<����W��E���'����_l�<)*ܲ-?�}�ь l��AH��RS�<A�4��%(B�йf�lQS�nR�<�Ռ
�-&�y����}iz #�	�c�<ae��zܨp������@���B�	�L�6��q�,`��2C�
 ��C��b�4qsT!ɤQ�ĝ���H� �B��8o��)i��;b7LP ���Jp�B�I�+-(T��U�TXJ���.:C��|�`p��_%�lQp�^�-�C�Ibq�ʅ���2�&8��HY�1��B�. FY�#�D��0��0��B�ɑ`,��ᴀ�C��M��3OĘB�ɞ=��\���?K��c��E�n�lB�)� Θ�SE�bj`��cQ�&�ta�"O���k�4����� >�Qf"O
=�Cmʠ}J����λm[<��"O
x{��2�@�i��P7W�x��"OFԳU�Q!_��`�8/&|��"O$qɗ%��(Yc �!� ��"O����՞H�4@�+I�.�m��"Oj92���r�x%�f�+�`	�"O0ly�+F8e(f( 6d��	Fi�"O�!��%�1�íqc`2"O�����ÔD��=Us��x�"O�}H�E�N,��"EA�B��A"O��!��y�8|۠ꇄt]par"O��)�`Q/*[�a���h=6<�r"O`	�f'R0x�\��	�,Q3��a�"O�X�fF�e)(}�R(�
'�m
$"OD��դ�)��JR��`��ZD"Od��AM�JxF��E���p$��"ODL��cê7����a�X�����"O���#�_
=+��A�an�;1"O�Ȫ5kP �Q���$4��Ip"O,$�
��e� \����D�6�j "O�+�+u���4F�l᠜��"O���M59D�)��X7�=["O"@�V��9�	�1�T�`�D�ؐ"Ob�I����B(�E�0�L��'"ODhH��B�x]��`�?���7"O�1:���-w\Z2��
S��%+�"O�8{�E%(���.On�D��"O2i	��P=��(�J�;}8��"O<����6aB4Bi�,t���"O���Ќ;�.���!�H_��2"O:�k�˴�4l�p �cJf�"OTx(�!�����^0iv�(�"OJu�$iM����KH>#B��I�c)D����C�F��)��D}��U�:D����CtmxP�Q��m���N7D�\��&үM�Qҷ��;����)6D���uˀ��!����L���U@3D�XX�E)�X�r����G����>D�,��ʀ	%*1Q���
l!�!1D�гÏS������-LZR�A��.D����Dt���A�B�\q��-D�H3�[�i�j�J�_�G�H��,D�x�U�O;Nk��Ȣ��Pt	!B>D��B�J�o�X���)~Fj�;D�\cg��)ꐌxb��)�2�{�A-D�ܳ6�@�W�X᳣���<[ju�ծ*D�|8#@�4��R�D9/��xQB;D�d8�G�3e����������m=D��c���5> �A���~���Qn<D���!�;�vi�������9��,D�d��E]��؅��1A����7D����2 ��� ��Y�"�֠:D�(A�Җ._\,���Ѝ�T@EO:D������nN9�T.M"�4I��$D�@+ph@����A�O�]1�4�q�"D�H���O�����76�6�I�";D��(5�B�(��e��h�n���8D�\�$�^32J�c�mY3H=�M���5D�`j��M ����S�2��u҆�/T�H
e-]�|c�u��N���<��"O��#��״hƪL�+�,Jʸ̈C"O^���;�Ztj�(
B��(�"O� �`P���i�4I%!��^����"OI�R��)|K�Ǝ�2C�Ȁ9�"O�P�6b\�tT�=���K�'��E��"O���N϶�C ����8���D:LOL�'�)UG&L��@�jĄ��"O88�U�D%h&n�(�jL-
��@r�$4��0*�Q��ɇ���Eo��gF�>I���.��'"٪����k�$�"I�Ce����'��x�����؅�A��7A���K<ѪO���DG�4(��S�V	+!�Y7&ւ	x!��7Uf� ���7�l��b�?#q����F�(d��E��b��������e�tM���qܓ���Y�Aִ|x@ ݪ%<�	�'�h�����("`�	b�0��r�)�$m@��|S��F>~@5�2&��yrF]�u����%\�y�VT �hW �hO\��$͂P�TBFB�:��5�2F�3|!��G�*X��#� >�J��w$��
 !�$��ԥR��8,H�*A�2�!�D��7�N8#�L^-c��Ӈ�T?!�$CB����q�M�2F��g	6	:!�$�$`y�s�S 3r��GG�<�!��ӻi���"�m�y�&[���D1�S�O~@�P5댄Z��8�ck�cx��'��,pr�	�(��ux�'j��܀�'�
�S���5W�2p@���Ԙ@�'��a��(Y�:���Ay)���"O�}0$l�(Z&���m�7[�X�t�|��)�*#���a��ӌp2�U��%& �B��w���$�Z��A��(d��6mU�Ity�	?�B���C@�w-<�f �!����_�"��Y/ƪFM5`נގ[�tԅ�QY��;'١?���`\#��>yU�)�I��b����ߣ0�:��B�K;!�������M�~N %YW��n�ў�'��а�����.�!��&kh�0�:D��%�μ���+"�Z�<�V �S�7D��+�g/zQ3$ŋ2e�;q&5D� `�C�B�2X*�e� vA���/5?��d�|�b�{��$񆅗
@�\��t%�x�`VI%��ht�[��P���|���acB�o������������As𤟓wb,�X����}e��ȓ|����� �&f���g�11���ȓi�z�ae��9���@��;;X�e�ȓ>�Vܲ��6TD�cwOT4e�D �'Ya~�jW%0�`����&l߈����0��>	�OJ���;!��eIcJڍn����"O���We�09���@��ӷ3����&"Oj(�h�>�D�U8m�J�e"O�%Y���#V�$9֨ <��ر@5O��=�~��'Ð���mǇ40`=i�%{-���	�'��
gJ�2m���'��= � �y�V��G{�OO4u�s�̮/f��p�DB�<^D�

���> ) �@'8]S�i
��'T���$��5^�ޑkq��.p�x�3��vL�O�O�#~R�4�$x��Y�a|����]|y��'�8�@��-Ƞ, B��U�Ɏ�D�r�'Tt�'3�\���n�r����$�-K��-�ȓV�R�����Wm�qE��|�taie*�j�	c������[�u�����	Υu��[��%lO��pP�mڣBB�pj�� �Zs�ՙ�"D��z�ʏ�N�H��6� �~���9��!D����3E��!��*Uġ�"�3D�� �y����5ҊAsU��
7����'=ўD�"܂�6(�w��zͤ݊��*D�����I�����aD1?x���<ʓ�hO�ӓ<��EmH<6��lc���$�����%?�N� M��`�%Z�	#n���nH���'wqO?7M��;�d����'�����9lў����'�L��X::����`Ah�M��}�%��}�!A��[3����NÛ�HOT��sI0ƫ����;a�S�h�c�'0�xb�B���ԌQE���'6b%�ǧ����{��Z�xC�z	�'Ĕe�2Ɛ&1Z�su���p�2̨�'��]i$�j~��!U��>V��p���9�S��oͿl#����C���@�]��y�Ŋ:h�aG%��+F��`-J�M���s��9Ӫ��y��0��� ?�`,:6"On�hB��#7s���iG;�P��U�O��Dz����� P��sG�� �͡�ޤ�!򄝎8 Xע�X\H ��_k�Q��SH>��Wj�Zɔ@	���􁆃$L!�D�����cf��V�XР��K�T1!��$�~4�'B>_�,�{u�Qt,!�߶$pb4�`@�#�8��H�"�!�$C"�)�5�^8'��Y`�5|!򄕂��4�%}N^5kS�L�L��C�	�y��3���7z�=�Х�J�C�I�
� q0�
f̎M�W�օkhRC�ɢR�N�s�U�W��p*�ȑ-L>C䉜��١s��\T�)Ad�3Y�C�r`�a��׀db�[��Ƌ2�RC�I75`�p��o�^8"*X�f���>Y�b
%tE�����.B���K0N �<	���Ӄ6E�u���8d:u�3C6J�҅E{��9O*L	SFE�4�t�g�~U4�R��4��I�P�(�=� �'�H�lj6-'���!��x_mLn��9��9D�| U�X�	��Y0(I�I�٠`f1Oj�=)F@7��!�d��M�����^}b�'!�� �'	G�ΌQ"%!Kj 	�O��=E��dH��zā.�"�L��$϶�y�m��B" D��ՑkTX�����0>��Q+0�,|au�[�Cg�ģ����p>�H<�wbM,��!Q�O���v��<1���O��I�B�<!(�(N:m9���B�5D���� 
�H���e(0J�\E���5D�8��4��)����S>�P'-?$�܀��W�Sw��G��
K������y��_)���Ra���J*�1x�hF1�yr���3͌��**l��i�'j4D�k复�Q��x���%lXp	a��1�@+ؠ��3����f��� 2ͅ2j���j'k Z�!�&{9$@��O��m� e�a!ڤlS��<�
ߓ?�e�%�.����!�)������|Q��*��4ȠBA)
����ȓ*f� ��IIQ~�c���<����=a��'�*�Y��)i�!��ѭB�^Q{�'���'�jH�lx ��^`j-)Q$�L�<���b��A;ێ�8`d�<Aӏ�� ��d��ί�^t %i�Y�<��G43���P�XO2fUHQ�[k�<A��~4B���� ;8�fx��O@�<y��֨g0Q�VN�34�.�� a�<Yr,ٯ2! �h�`��,4�M�b�Y�<rL�Z�F-f)��!i�y����<� ��3��vHxJ�K�'Kt�q"O��3@"�5:K�(hce��f��"O
�A��K=Ap����)�p@��"Of��d�;�P\��v�h�"O�m�'�8S����D�|�b0�"O�l���E�@���C5~�v��"O�ui����q����H�=^��E�"O���fkXA���Ӱ�,g��&"O�����B/Q���@@L�L<|��"O��(�e��7g$и�/ʿ۠�I�"OhD��-�P������J b��{�"O<���#�Z$G���m����"O\,)���R��#��ςC����'"OR��gIF:@����F�&' ��"O���"l�;y�T��F��#Z�b�"O0�!p�]�]X�g�8�D�"O����3P�@��S
2���Q"O*I�U�є�B=�'� &|A "ON��`��O&A ��?�����"O�P��	��,i  [;l�"O*����8����CQ�}��qa"Oܕ[��d��8C�&dv��:�"O��a@)��2UnH��Bе;v�e�v"Oj�y���1����7)C�� �"O�����&h��!v�J6F���1"O8���ē���-x���&3A��� "O�y��d��E���GI�z�v��p"O�D�T��:�.0��h�,^~2T[s"O�y�Ɖ�b�֤�e�-^�k�"O�[����dj!	�.S�� "Ob遗���i��``�H�v��x!�"O{s/ٙ��Ɂhɯi�X���"O2y���
}�603�h��	�`�e"O��
��̮Q?�8s'Æ4�`(�"OH�6�Y�X�6�1�*�
囲"OȘ
W*+����V<r�v�Zv"O<`:��Z�Z��Y��$�2ɾ��"O т�B݊$�@I�FԸ#�V�9"O*�5�.r��x������"O4�(��;P/D��%�T�R�F���'O$� �^(0��.P�s �H�'�l=1��[�F���ꍣb/��C�'��M�d/>Cr�I�Q��6R�i��'��M�򇋺6#X��1	U�S�h`0�'Fֹq�I<\H	p��M�|
�'���@7���Q�(�ehI�D��͈	�'�8�k�p��A��a�)4v����'^8�)K��
U��' x1�'غ��f��O������Z�haj�'�*hqkY����'�a�t�[�'��XCD��	d0��1K�3A]�Ņȓ!X����I$NL<��N�0���R�TE�!��[4��Vm\?[f:Y�ȓ�$Brl�D`|�1��֭ ��ȓ_op��`�Z�?���sM�B~X�ȓ3���+'��@���!I!G�v݅�Pdz]�EąI�6HpK
e>���6�� j���9X:x ���]�8�ɇ�Q�Azwe\8V�P���r�<l�ȓ7����FcAb�{ �Q�	�jq��%$��"�?V��K�o��#Ct�ȓy�������w2���ү5�����m+�钋 X��p����l�t�<��&�]���0��Iwpj���. s�<� N��3�  �M�g�.ȫ�"Ox���DĔ{��(��=�@X�Oz����0H���q����,�H]�!&��+xL��'�PZ���8�Đ���Q/m��Z��D�>H3�|3c�/�)i�x��'�Y�a8�HB�(��VC�IJ�:�6��>r�v)(��[� #8�y����ƫ��N�PӧH���B& �3cG���4����6"O��吰T�օ2˅�W�� (b!}B�
A�Pu0�$���M.-��25-�!2�"�:eHZ�`a2B�YV"��r�!7`��#��: X�p�Q"�-�F��I�C���b�́�&pȒ#�>w��#?�'̔�i���6��X�4C�Q
kӂRp��C��ўp�!�D��:�{!��1lh18�`�Q��I�+��\�5�I�"}
�ʕ�i�P����2���KVn�<��eD�r^NtiCJԎ*��,��/̤��	�S	�Gޙ��g�~� �U�7�U�w(µk*l��	�L�(4j�Z	-��a�wn��+���Oؤ����'����5S1z=ʉ�����F)��WN����/�SW����/.W��P�aB�#M"C�&]"�A��-莜
�n��(���nY�)5�=�)�'&�v�C��ԕz���uG(-�5�ȓx�J��QKG�p��t�pDA+q4�\��#��`�2�>A�q��!)����/�uA�KHJ��y�E��Re��"�"�����n����eNNF��`���������	A#P�h����}�B����D�,y�IЋ
q��U�r�r��޷;F>���B 	����ȓA���uE��X�H����Zq�.��ȓR����s��v�.����S����R��ѓ�Ⴃ<#h�傀 �B�FɆ7H,Bቆ-�4d֎~�dx�ȍ�5�v�?�[>�1J��4�
�]�N8�Cf��V�h�bR+�y"$��0Θ$V5K����C+����"��E����y�ff΍D�Ԯ�"E>T3!lR�H���C˦�y�-��f��s�I�Qx z�띶&ܛ��\�Vu�9QJCE%f�㖔�4���s� $���J�|N�:t�Pu<U��	'�q(pǊ�m*����S����	?{���F�ҪN�>��kK�R�����H<Z��'�<uZ`�Y�h��E~bB3*і��	S
��U;���l!T	�L��=as�]�wp����0A����i���ȋE	��sBͣ{���]� b�͟8f
�;T ��n�6Az��������$��2������Z��-C�O3�y2���
�eҮ[���2Ơ�h�a	�� _6��E��-c�l��OW��X�\����>�1,ǩ^�-��c��"�̰�Gi�_؟��c��P��h�׊�F� Yz��?F��b�ȗ}���P�ѧ����r�
ͬ��O+�V
,��p��f���Qz�+[�'�ָ���
-��d��&���M:3k�x4~��� V0��toC�g���Ңӕ5ۼB%3�O�X֩�"^jb�`%����E��g�<�W �d9p!��KX� )��[`p�Pu ����w;dU+`�ٌe��i��`@>Jl���'������	AJLpB4�w&zl��-�(Oy6�@4��%C�\Y'�ǖ��$A�&!45
`7��6�)K��k���h�,���է%���yZ��Q��R�i���G�ig����NH�4�i
���=�$A�6fY�_�ȃ�C��6F�a��I��u�旺#�*�8g��Q�	%I����gO�+��H�D��	E��'V0��IF�9�,��IV�W��i�K�f��!�2M�h� �I�?$Tqt���>k���f��5z�P��cF��æ�=l�ay2���+�@ F皮k�D���s�q�ҋ��cq�7M*��MBWN��[|�X���7^ܼ�RH�?y������IR|v���SJ�+o�����5�D��$�h8蠳�Jκ�$�DjC�\A���'|��@`D�M�O�aU�]�|*��
�#}��� N�2��T�Q#E�XU ���8�j��'R�@� M2�=&�
7?�`�g$~�n��&��*߬xo�Qଠ��]�]�-a5b��"�ᰅ	L����M<�G�P�3��-`PH�6x�,�!э�qy� � t����E4_���	ĪLp�&ϗ$8"��R6M#W�A�s��,��˅�̍2���P*�8����]�Z��S<,O6��e��p�H�1�_���`Z�%R�hVL\(�t�B����KŮx�MK
�T�*@C����j#)�?)��ѩ
�8���Ӏa��9pJ��p?A�dO!BwJ]	wMүp�jq�ԍ�M�I�g��r� ��Kپ\�Լi_�ڪ�ly�̟���b� V�htB
50���fګ$�Z 9��I	+v��tck��tb)��es4`M}SX�:���Y�D"1OԈ�GE��Snb�.�� �	̾(/V�b�|�/H�r���	�t�&��1i�����¤j����JF�,��?�lZ0��:שפO��@��-K;p���kp�_<�x�,��	2�!LO�m��� ˒��e�@�c�D��%�;����a�N��ț�T(���O,� ��K@���C�i�t���'Hi�֌ÎmZ�E�7	�$H��
�dG�i�<���D9�dᆚ6��5e4f�8��b����`��p k�g7.mꩇ�c�P�8�!U�Y���B%�.4<rD��v��%�"Q�RW�	��'"$���g|b@ Pބ0H��j@�V�l��T\�9p'��Թ	Ü ����ȓ}W�0��iFx���!
f�����y��8J�@�>Ulyk�kڃ4�����r�`lK�L�Xf��D�&�!�'��D�@$�s2Y�.K*:H\���'��2u�ә ����l��:�����'�"�0��	-qV"Yp�Ό�7t쌃�'��%��Y4l4"%����,Yz�']�8s�^� .�������!	�'�%Z�%��	m$	S�ɀ+�����'1	��ŕEE���Oݒ�m�'M��Z�'~ݠ���bL�	�'�đ�7�ݾ7]�A�oʗH�R 	�'���c�QP�T'[F��ƁG�<)���)-xSxً���h�<�2�){+���#�8r��;bBNgܓTP�!�3���WɅ.߶��T�9$��la5"OF��� � T�D��w���4��9"���B�O�1��3?Q��* ���ge]�+8:%R��_h<Y�aX�!��Ҁ�104��`��	,7��"�
ˡ����$��F���S�:��aˡc�F�y�`Ә>��I���OY}2���2ٌu{d�˘W�r�j̎�y�n�ArN�UFBYN���s ����XK��볠-�#��e�#v�^��EF�2y؈���F�<y��0�F�+@X�21p�H�d=`�����>���I$����	=t]�"j�W,��%b��У<� O�<v�}�%��*�|D*��1yy��0�LmG怂�N�&q�>���P:nh��c4n�,�pp�	���֦�Y>�O哏{֨����@�Id�IEz��'���g��|�'�_LBC�I�_qJ��RdZr�z̰��"�r����/C�9W-�Y�4���'��	���O���s�MѪ ��!�5͂�Dº�ߓY� ���Z���6�͌"�|������]����2fY����'��Y2d\>�z��p5�_�d�|�acs���?�3.Q9$���*(ҧ/`8Q%�R�ɂ�����X�b��WX��ɝ>x��χDr8]��GH(qblȡA�@(��hXL��D��'����sb� ��5z��7&��p��'���[�	_$.sJ����2	�����m��'U)�N���T5DU)��UmU�q{O_��{r���c�0��u,����˅��1�x"�d�7J�99�J6D�P�ua��;[Vy��_�%�ޙ�L5��;2t����+�0v�>=[T��S]RĻg��1M����i9D��C�S�(�V	����(��{��8%M:q�R-�p�)��<��FS� j��J���:��E�]o�<����Q0
��N�-��ar*m?�q(ذwt���DO�j;r�IQc�w\�C�Y�]�!��/N������W'����@�f}!�d	.%
-C��B�4�I��@
$Y!�$��^ظiʄe�;ځ�N��J0!��9=^�x%H�6F��Ip[77!��Q�[L�0Rd��~�zu&,^�$!��݃��!��n�%�hI��)��!�$�/��-K���7�:�R�\6]�!�� �Zdє<H�q�Ԇ\�F���"Op����W�F6|���-� �Ű�"O�!���*a���+�Ip���"OD�c)
�7�*�hADR�u!""O��9� C;yTH�a�J4(��G"O� ��NK#g�L��&M�80�b�p�"Ox����ZoǜXxT&�|��XyQ"Oĵ�w���0U�	�K�|`h"OP��v�Ò5""���D�)K|*�0�"O�0!ЂT'}�01CI)89���3"O�{�M}a��B7l?��YR"��y�!�$���@�+�c�Rt�&�S�!��U�aW��/�ddr�	&��5	!�$Ѕ{Y��a��;Npj�q��,#�!�$�5| �����>{�$;'�*K�!��{���"[�0b���C���!�Dω!Z��STOI�aP��
�Â��!�D�&& ђ�̶3�x�x'!�7�!�$�%R�`t8q�$����G+`z!�d6D� ��2*C� ��ԃ�'E�Y!�ɑ����h�U��Ir�JB!�$��;��yh3*��fypQ�J
�52!�dӧG��e;���Jh�˖I�!��B�!�H�3 �͊rB��P���r�!� �
4B�K� �2DM:dA%���!��V�$����rS�-Or���j��?�!�&s�����.�->��Z5��(T!�$F1:tuk�H�;< ;6f�;7M!�ѱt�N�u�K�q�Q��O��,!�$G�e�21����#N� -�"x!�D[63�L��S*KW�pp쒑n!�-�\dQ�eƦP�
*
o�!�D��# >��GO�8nLX:1��Z�!�D�1�R	Bo�q��"��L�!�l3x0i�o��<�(g��9`�`C�	�sр��匯&�m��,B�nlC�I&;�xPG��5��pˡ�.	>B䉮p;D1��P<l�<⯜:��C�ɂ^�aQ�m
�dB��Ã�� �C�;]V�1A2X.��Q�Y�C�ɋ5�h�Q�	�A�\9�A_"+rC��/r�n�[#���M��xY�d��iG�C��1YD�|�0�9�I��e�C�I�-�z�(Ӡ1)�a���BlB�	?���6.��D���M̡q�C�ɬP�^��$��("Z�0�U`�-c܀C��9p�#�O�:��=%��C䉽GMNI8v�;�`���li�C�*+�A�1/�&9bX��GJ
j�bC�I
z��,s OY� �j����F(&>~C�ɾ-�� )�O7T�(���<1�B��:?m 9�U�|'��$�TG�B�G�0y@��a�ѱ�ո�hB�	�p���(�N���q���ռ0}RB�	��P0U�V44���!@g����C䉯'ax}@�A'2l�
@!�%7ߨC��b��B�Nڽ
l�� (��!U�B�Ig7�Ɉ��+zR4y��ݑ9ߊB�I!9m D�k$;=��0�ۀ`^C�I�NF���\�e�h���[�T�C�ɺ۞,�q�Ǒ�� ����]�C�ɇ�!�o�>/I��,d�EP�,D�8��@�+*�B�iV$K��w�*D���eS,�lQ���Bբ�Y��4D�� D� �� �f�.9��Τ%H:=;e"O�MS�'�#�4�sR�R�125"�"ODR��8El�@���u30��"O�(SL��HWN�벢%.��S�"O��$��JCB�sÆ�'&� �"OƄ�G�?xz�9�B��D�
�'b�����9W: �f�μ�a:�eS�}T���� ��όA(����IGJ
YD��1[�в�	V�0¦�p��?qP�y��\=4
!�D�>V�p��L6K���Oއ+�I�e�E�@��~��S�O� �x���a��`#a�[����'5�H ���ĕ-Q��h�p�>1�c�)^�n�ᢑ��}��D9O�t����[�����?��C�t��)�D�4-��Pr/�&p��2v��H!����Ǝ B( Ŧ�}����ZΑ�92��1����5��$A]\A&i��B�_���{s拄�yB�NI�%1�l�Il���
��d�d�vx��KT��)�'I�d|�X�Bn��쏐S�
��}�$��O8ZY�tJ�S�mBH������%��y�L|�>���Mk�v=��N5<ih��c�^؟t��7��ѕ�Цt�����>���")\h�RN�3p!��QP��=1� �g����O�F����b>�U�:�<���xi��!��)D��`���=g{����$!0�,�3b'?	��H@b�"|"q��y^�8�&�؅�r%�4��|�<y����?PtQ���͢|�'`�~�<���ϝ7x>i�L�@B$����z�<� �H*-���V�G�\���t�<��BD1v�<`�ñ4R�p���\�<�G�ѭ|*
��R�4U��	�c�\�<�L�Qc�}
��,m� BJ[�<�Eφ�i}�ae� ��a)rEHT�<��L�,r#�i�r/�b8,հsNU�<idh�κ�Hg'�Ut��$�TL<aD(��^O����%�:Q*܎f�@zM�B�	�g���1�+E�'�Nt���9yc�?�FT/ܖ<3��D��my>�rd�o������L�<I�c��1�n��F��Y0~`��NCO}b�7I��Բ�C�D��\���g�%Ixm���fC��7P�����+]QP��.S�\E�O&� �<X�f�&>c�d�A�
-/�,�O��EĪL//�aB$��X���T�|����7*{Z9���8':4�*�O�{O�0hRI���
�!H(tx��Iz4�9S
S$6W�Oa�\����$W�a�%�Or
��'�ʈ�@ĉ�c�v�E��-2<A��O�3�Q,*��y�I�"}&�Ж`RXU��/)����$�T�<����f�)��Ɛ�4�r��!�)��	!aoz��1C����g�zy, ��U�Rf�Ւ�W
N��ԇ�ɝ{��D8��ѝk�j9C�l�RF �q���@ɩ��'t҈���������H& �Q���䐥nvր����}�𬣌�4��>YK�`A��zJ,M觌�&�y2E�+;����̖9Y6(�чJP�eR0���m�_�h��EÂY?E��'&�+�D�9(*����w��(�']X�"��2^E�Y3�͢v�25`Х+��<���4qn���|�L��k��ӧ�R�� ^!��ǻB�D�� �D}���{�C r*�XP�b^��M#q���_������'gZ�B�-��<��ꑪhzL\["&E���4���QM)�D�9���0vC�-/.����
!I�[8ZTw��A�8X��GW���S�*�(]����i���!�i\��/??J`�V�O��`S B�t��	��B��C#N��.ő�DݤS� mո<8����i3���$�ہ.��*_ky���'�L�S�t�`��	s��b�n�+A24���) �O�m"�Mұ <y)�&B.�L0ab%�� ���'��c�� b�$�$�Ǝ0�:Cĥ�6\ ���'�`џt���7�@y�f�E��!�����:S�0L�:���R�a�)c�'G*���B�L5>m�`�	P?ͧ{BM.R�'lRD�l�[ښ�YvnQRn�Œ)Oj}Sf�غCCP�����$�M?�Z�n�0%6�� ��H����3���!B�hK#hQQ?I�'#Y:�%)�;,ODc��2I�2 [��,5U���2"�
8�4c�f飥"ǢLz�8F$��`�uP�';}��O� q�F�P)��;�1�j]�L0�O�,+d�/WW����
�:� �3V����%��Dm��!�~RF֩��i���'|��d���d�q*�F۱^������� ^�GiP�o�~ݖOݤ�����5�ԁ�
��;���H�'y<sïc�:��S_��S>t$��&�����JU��##
T t��hz�H�<y�.�Sމ3�����(�\(�"��8��pZv�~�d������x�N��01�_�3az�kL=��p��Hc\�3Ac�g��'bX�Ý�Ϙ'@n<bT�Qٚ��炒!>���
�'69��$��(��@ݺ#0Zi�'��_N�e���I)�)�Fͅ�td.��'���ȓ�y������S�="'M��C���'?'�6q�¡9G��P�ȓ�L��6��9J�Lre�T9�I���p""g�����z� ���4��:�&�5�ћV�`�W�]�!�(�ȓ-��x�F�Q���S��[�P=��H��#�g4��C�/�I),�ȓe�Zy�wÔ�=ô�;�d�~�:���r��}�'+��oZ�X'F�f:�5�ȓ~)�3���g~�1��/L�	��8���0�Dӟ&���JdC/�t\�ȓn���s�
 �B|�ī�qF&���l��	qDÝ<�vb���GB]�ȓ-gX �%иN�^<Z��2)���h.���J=��0Ď�x @���@���O`� H�΍'W H��Tp�8�	{�p���C�RGR��,�f�S�
�&u$D3�GGoJ�ȓhF���m�4�>ȳ@frn���ȓK���a�Ď!50��\[�T�=i��̮,U����[2zw8�Um����!oU!�s�r�PWjD�:����G��8gS��
'��^8eV>�)��l"u�:Ɏ�ʵ�� ����M!���|���Ӓ*[�8 AQ�Q,�Ia��'�O� sɋIǖ�mIT3��zv�'Ş�襽U#	j}r閩,&2��0�A9M"�pJ��yR��L���rw�A1jR`��P��� o\H�pk�04"*A�@z"H� [���ŖA�<� �P6��"���H�t��UE�,Jm)ő>awK
����&]ܝ��A��h�����Ɖ0h٪�<���
&_ޣ}b���2��;��؀U,̱��J`Aө�: و��$
<>�k�CT{�r-����6F���cAû:F�O�Ss�e�HO�4��������b޴a:�,ȳj��Q͌B��!]�D��D;w����FJq t�dԜ"_N�K���m�*�(g�G���	މO���Z����G��{�ޡx�f4
	ߓ6]�=�'-G���6mS v�f�9��Jf���P�!t�d�O�( �3?�p�\!�Rh&��*�"��r�Ao�5[`�ea;?G`#}���8�(I�s�0��o��Q�t������0?�8"d ��N@�C��és|D�k�Ǔ���h����$1����*DM`1�ȋ�!�d�z��h ��ô	Uc���Im&��v@~؞��uf61��t�7���j��s�E4|O�Z!�>"QHѱ�47!�-@��ɱ!���K��?�H���K.<�+�ļI�İ!�ׂSÀ��?QPʘ��R` w�?ҧW��)9э�Ss���ff^�cll��6 5�C&F7�\�/1"�V�hC��8ajyK>E��'�`�	�㉏`��Iҧ�ӌg�"���'p��"�LJ#p��H�&��/���'S.�Sz��%�HP>^q*F�^�nA.̫�	<D�@X'�*:�<�p�`&
D��c<D�[B��.��p
]'HǞ�U�(D������L��Ʀ�B�
&D�� "����L�DU\dӒ���"O�TqΏX[�A9��I"g��A��"O��HP� c ��E��~{zh��Y���aT�ܢ"Ez]��˰8�2y�ȓ>����ԗE��3�L�nX�ȓU�"�ˣ�F�q^HC5,�m@�q�ȓx��Ma�iI�wd�@@ &֫hcF��;�2�p�-G�dU��ʁ������ȓD9���ŃN�А�$͜1shP��|պ$�un*^nz�:���z�Ҁ��+򜼉qA UD���@MI,���ȓl��h�D�A�x���;U|����e�Ȇ�Lm&���0'�;9�6���v׆,ꗫX�(-�SF*Dw�A��8����Z����@�P	
:�Q��<N6e�pmB�L����s$x��u��KZ�ZuHB������C�e�I�<��jB�1�x� �+����gF�_�<	d�սN�:`sb��8=��M@O�Z�<�Tf�"$�@q���3R4���#�m�<Y2ŕ�?�A���}��3dQ�<�doD�,�"l�P/Д���&��R�<���n�>Dh0���wji���d�<A�0����U��'��l�FOf�<I��y(-��f�T�<��gÙ`�<�f�>~Ԫ�Qa!Rk�.P��o�D�<����,�;A+�'cNy@��@�<Q7�8m�i���ޞSB��7��v�<�v�4)"��`F�m��@�T�<�	@?&z,\���V��Q�G�U�<��뀋1'ax�R�i ��Hz�<Ya�ձQ�� .�h�FpP �Zv�<�rEJ�8��iH�'�2AW�}@��Lz�<i�M��<���X �P� d{�<Q��]%F\�p�gO�/YJ�Y�&r�<��Y�8ܒI�v��|�����o�<���Ć7r�M�&�6���6�~�<a�CA�\ш�g�_0�J��2�G�<��ϳ?]�pJ�������B�<�W��L�=;À�+y�Y[�.z�<�Cb��ʬ!��Bً%R�[�w�<�D�Z~$�!->sn����J�<��C�5R�l�T+��^�؝�����<�gN��Y|\G+�9/L0�R�PC�<1�H8�"Q��5"΀���a�<QH@}��I@�H4R (D�V�<9��U(#��#u�Kd����Nv�<�a,�Ă
"�ҹ�4'EW�<I��ݱu�
�b�,�M���nNw�<��]l� �@�R�38�J�<P�B]F����,|U�e{���k��p��J ��	;�Q'��!�l�FW�C0�(�I#+��%�?%?]�6��7}#L�j��!
�d8��&}ѻB�O1��	�RnV:�H�K/k��i1��d��@ �$���O�� �{J|:QE��\�]"��R/� 2s�	C���2t�)�IRa>t�9#�}�T�P��^�&S�'�p�Dy���L�#p�V�01��	P�	2�J����	�(O�>�k�<d2LY���^��x�7�k�bɘ��N8�_|Rى3���C�k��I�K{T4�bI�
�0|Pb·l(�j I��
���@��	v�
���H���ą�-�ldzrB\�/=�����E*�yB�F&'&������S5Wh�a��U�:���닦iDH��ّ�\a�C�z?)R��k⓺A���4�>A�\4&Ujy3H�G^T�q���P�AkB��1����˪5����Y���BG���ӊN("���U�a�T(��O�&�"~� �P8�H�7&iЦ'\�.C��ʑ�K#��"}0��4��B�OՊ���$L|�f,�I�޺�
ç#������XnU�L�`��]� �'�H���?�qO����"��6���+�ဗ\bȐ��S����f���S�>�g?��ܙ�E ��KN��b�*A�@6�|r�H�@ b��>��gʛp� �	���#�tt��#D����H���H4A ���7�!D��h!cɢ(y���D�d2x��?D�$�쒗��%�B�O��P��C<D�
gƛY~�{�C�r^( sS9D���l�#=�R�U!F2i��2�6D��S-II�رX	��i�y�s�9D�t��������O�"(>��BT(8D�`i�$�k��ո1�-p�,rr�6D�|����&\��� 
[�'=�PD�4D����8p���e�3'U��� %D�|��D�jK�LÃ,�561�<�a$D�����JJ�m���B?H)��&k#D���d(&N, ���4p	�P�&�"D�x��P�]NT�{�&ʝY�|$�7,!D�Ԉĩ�!f�<�'�%uy$�C^�y�{��8�֕(m�%���&�y2Ɩ�Y0�mC�#=x�tC��+�y�hW�_A�Y�/ �N�R��G��y�b'Ƅ��Y;�XPU&R �yrO�,����g��^\��D)Ӓ�y����&���@�� P�d��yR.�K�(��W��9
�������yB�ь+�8P��˔�uܜ����y��ןL�zM� �F�f� B��P>�y��NWL\x��\jNɹA��.�y���5���H RN�۵)��y��?<����ꕣ>�6��4����y��+sL�W#6�J��tΚ#�y/z)pr��lЊT�R�Z�W�j���8e��c�qTD�ed�4�lL��^�M����&�e��\:"��ȓ	Er���٤94f�8�C K�h��\�^MҢ��kf�HC
�-"����M9>�RQ��/�����-k�R ��Ftj��� =i����F)oވ��a��`�C����=�t'�.T1&�ȓ:�ڨ�4�_+r\��S��.T+���~��Is�E6tQ��iGc�$6X�\��?@�ı�MD�7�\�9��"] >5��4�t�p�c�+R�µg� t�`��FI��
��þw�j<���#x�hi��AJ��"�Ɉ\����2@TI|����M��9����Ri^�y��C�RՅȓAav12bQ(V(,��.�6{�lT�ȓ*�Z�I���f;E�.G�V�E��Ne� ����q���$���EѠ���9�)��Vnl蘤BA���ȓH:D�j/r	�E�Z (�J�ȓ/� iv+L�wG�9�I_:W�لȓr�4����A��2b�6*<��ȓy/*��Be�P^y��a�)���ȓ�����1���3���A��y�ȓ
�(҃١;�:�c�G/R���ȓ �$�%��$��Ÿ�D�O񊄇�a��P0L�-5>b���G��Z�d���}k��@T�U�,Ő��2_�Tl���e hi��ف�����Y G�D!��'�n� 
%B��u���9Bg�ͅ�S�? 2�����2>R��FX�<v����"O�]�$��
J^h� �!H�}Z�"O&8{7�Q�Z�5c��ӶM+Vu�"O^Y"g�[Ac6�yV��&!$4��"O�h �ŵ~�h�%�I/@���"O���*�B���)�癬T2Bq�$"O��02�F�"�H-p�� �"O�!��	�6�"�ig�C�k�k�"OŘĂK�:��j���g���E"O�(�I�\�h-���C.G>a�"O�Q*�� �P��q�]�1��a�"O\�2��6`[��VH�����"O@���*H�A��@37gףF���"OL�˂�ڄ��i:���eg�=��"O��+@OXK� `P�^�7b$ͩ1"ON��a���Vڸ�bu,A�w�}�"O>��&�+����\�, S"OT`1צT93��(BI�nb���"O�]JF�͚A���#@b�M�V"O&�pCR�4��qIw����HD��"O��'FASV����U�,Z���&"OdX� ��5:̪�G'N�t8z���"O��p�5q|<���fѷ˦AK�"OL�d捚 X�h���'L����"O�	Sm��IE�sM�m!�3�"Ǫ2uÓ<�ѫ;,�֨�d"OА�@�u|��Ib`=��"O��cÉ�<f����fp�;�"OB�ò�W�>�)@��;bS�"O��aAJ��9�W�r�6t��"O�ٛgV�8�n�h��a�l��"O�S��%��$�t��#��0��"Ox�1�G;I�p!���ߪԺ�"O�����$�=���L=T��&"O���� �� �d�I�O���T"Op)CE]lw�8��q��f�>�y���%g����Vk�,���0F�Ԁ�y�#ڿG�i:0k�!qa�Q'�c�<yu���#�&kD�3o:������X�<9�(��7�*i��L�d
Δ���X�<��M")Z�T�DHH�Ms��uAW�<��M�J�2!`E�:�Z��w�R�<�"$�5����,�0�"hB0CXw�<�A"|dN0r��-J<\J�AVj�<�Q*g�t]r$��N}j�h���9�y�Fd��Y��O?���`t�P��y�F�`{�\�@�*2����+��y���3*��,#�*[��l2U٘�y�!&�� ���M;��Q3����y�K�?�e��ݚ%Й*$K �yr��[}h��FM�# �a�GF"�y�+�?h�pa��O�)IfQ��Ͳ�y,��y��&A���� 6�	��y�P�ri8�p���F�
��eh��y��'����Ĉ�,�*}�u���y�ğ)J����1+߇���lJ��y�i�/P�����`ȪX�yB���y2����iŘN��9��b܈�y��b.4Ţr��-J�iEI �y"��/F�)�UC�G�h��E�3�y��?0��*�iR-9wb��d.�<�yb�]�vp��3)E5"���5�'�y"�ܴ ��'��� ����yRf��8�y�D��-¬���J��y
� �I�1�Wd,�ԡ!eƎJ��l0�"O{���`�u|
�2�ϝ2Z�ܡ�ȓPb�њa	đ MX]�$��:%b>�ȓ��p��E���KӎP8]%��ȓ{�r%#�,i�H��H[�9׺��ȓ/����� �c1H���E7.���ȓD&f  H�5H><X�#Oɰ/V`�ȓ(�$��e9s�! $h��5"�ȓ|FF��+�36'�0����'Py�8��o��H��4MT<ii�,*Tt��s=f`�Vŕ>��� �>�ń�=�,e3e]�8�F��b�� nl�P��?��1��AH7�����]k�̄�/�v�@$��eL"HK$ꟊ5��e��nB�rb������fϭp�0�ȓV��;RI��~	ĥAcT�o6���0�}�O��J�fE���B������"��6U�ByyG��MGPu�� �V`;��Ÿg]����c��΀P�ȓ��xPD�۫hh �*�?�A�ȓv��4P�&\~�p���g����ȓ�V�h����0j�rU,�;,�e��ah8�k�l�#vdzԇ;� �ȓe���*q��_A��a��?t5��ȓO����Â7d�fQ���8+�؅ȓV����
�i$�����F�^<ⵅȓ/d��B�?�x%���H-�H���o���N��]|�#��Ϭ-����T�� �3���V����D΂��݅ȓ/�P���"Y>������m��E��I�i���X%y24�E���W�N��ȓĢA86,GJ)��F��}T��2�\�U�}�|a����2�Ȅȓ&> �	 ��!
����1��M��p:����13tLB"�G.bP��e�~a���f��udb?b+@��ȓZ���	`�T�A��'��3#� ܄ȓH"�3q �Px������Y
���ȓ9�MI�KѤnRqB�!�r�p%�ȓ]�r���o�#@1"W(N�%�r���:��BF+R�wZ�IP�ߛ+pԅ�#8æ��
Ϥ�8En��V��Ʌȓ,�mM�t
	�jH	5h`�ȓ`'FQH����0�4P�&=�l\�ȓ.�PJ!���c� 8S��:��=��s��1 4���#�BF��D��rzj�
R�G$���J��T���
y��-	�&��T+���c3 ͅ�G- ��  �,��5�B��g,�-�ʓGpH����>`v��ٱ�[�@��B��4pƌ��hIm-���j%�B�	h�y"�nL�mk
�,�(l�B�	� ! ��[�%5�`�d�D�'cxB䉨��	����3Mk���#�0�&B�I$"qVe�te�5j����ã�cM*B�	�(6䑫m^=;.��n���B�Ih�t�X$)n��8�'U�B�I>���w#Z�<�!��/vFBC�ɤnJ���c�x�8�'�&z�C��| @���u[�(kqK�^�DB�=Gc��ۧ�* ���X�NdB�ZcRڞ1.|M!��C�_��C�	06��MB0$t���j��>	
�C�	'w��X��ϓA�P5[��\�g��C�)� &�`�dN�?(e&,Da�A�"O s�ʞJd��Rk`%�DE"O�Ի�I������^��8ȃ"O\+��C�_�����'!�����"O̅�D���qa\I�,�&D���@"O��;�I��U�P���$�.<��x�V"O�ܢ�K�a>�}	 �+�f�"O<,c��U�(V�Y`�Sk�ڵ�T"On�#$��%�����/�*ͩ"O4͹'.��i��l�a�ք72e��"O�u�   ��   �  �    
  *  V5  �@  �L  eW  ~^  i  �r  ;y  �  ۅ  �  b�  ɘ  3�  ��  �  0�  r�  ��  ��  ;�  }�  ��  �  7�  y�  [�  I�  �   � z! �' �- /  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%_�Q���m���R Q�t�A�,�Or@���A0��, '"ѽv�d��"O쌩��9al��;P���u����"O��d�AR	�N��>����3"OTP
0U@F`�q-�#D��`��'�I%y��]����Q�}���7i���$�>Q��ۑeK,āc��/:TR	еO�'���,�r@k�� c�x�x�iY+bB䉇KxHA�ׄӏO�jM�6��TK��	��'"�>�Ɍ[���zA&��D�Hq�2BQ<S?P̐�'��L)��?z�(�4[0�`��ٴ8!!�4��'�
*m�������q)�{��d��\���䚀r�V�+�;<��{��)Z��K���ѲBKG�,�4��� @�<��B_y�NtCD៙n���S��զqE{���i����j� ��i�1B\�#
ϓ�O�zP@C!p��2�"��yv>(��3O�E{��I;Z7��@'�4r}c�N�W<!��6
�\������椚�2.�P<">�J>yPmS�e�f��N�(3�v q4��H��p=�!`�=Ԝ�J9$���� ]��hO�'
Cn�HRJ��Y<��'A����mM(<�p��=�q��ǹh�����Z�<	���y�>�1�L�8`�B W�<�ЄJ�H�m2w#��x-�%��P�<�ތ��̀�ʘ.f� TO�N�<�#�	n��(�%�֢$Xd���$�"�hO?牝��A4'��Hh;@�*`u�C�	"���(P�"xyv�[J�Db��n~���O�Н(���O�^,
c�Z{��AI���dE'�2x�%
H�ض�ʵ����'?���'��x���7:R��g�'Kn`��d��?q�'ȰY쎄 ��G��n`��'ή����D�p�!Q�P�v4� �'�H�b3�Țe ApQ�\��{5"O�M3`+�`� � �^�4��g��Ȅ�ɖ;��2�.�2ye<Lڔ̒�7sF��d!}��<-.YS�%Ԁ	��l��L��y"��!!X0�Tc[O�2e0�N@��y"G�:?���D��I���RD��y�hHP�m��ȈF��Y�#E��y2���}qx�b��R�����'��?�����1Vj<CƦ��?��0�2,7D�dhAAڒ ��@I����Nx�	D�3D��9��4WS�ț���	2���A1D�� �YCu���~ۘ�!��t���zA�'�!�d�j$�8��1���c��sp!�$���`���ݙ^�&P�&IҮ,T!�%d��]��a
R�J����[�QF!�dZG ����]!���&@�>!�V?�N�؅	���H�-��O��8�S�Oavu��䎘���N2b���8�'-����<2��:�'��M�~("�O���I��<����O�7k�ڔ��0���>A�`ٽ����]�c��p�uj�ޟH���vx���F��:|ʢk�rΔA��F~���]8�E�C��c�P�*�'��
^C���i���9�A��T �~��)ڧ&�q����1��P�W,�4F����ȓ2�\LA`�W��<ё$O�<��)���hO�>�xe`��5���s�H�s��p�6D�\�r�H�<��u��؁B��g4?ɫO����!V���sЖ�hA��:��~�T�l2��Az�y��'ա77 ��%F0�IA�����&��@�y�&�U$j{�dA�d/D�P����� <Y��(TZ���A�?�IS�az�h],8T"(A D�?e�Y�B)�M����s��x{�f^&�~�*���?Z�ZY��"O�X�T�L�.AV�ZG�Α����1OH���df���5K@��B��Z�k!�$/Ei�M;�䂅}��0XUfܢ_!!����AsE�e����߅!�ѵ
]f�ȕl����3/�!�e�V�
�M
+����B�"�!��ǟHH4Pɱ@D�d���QQ@�y!�Ȗy�~��VA�tI�'mӳ>f!���1L�0a��3J��(���k�!�E 1<�v�τW0(��ѳV�!��$pӀ�b#��K�pl�-���!��%~�H3�M�&�N� Q��I�!�D�"Ap�<i��+p��aaqO@#\�!��³m��x�pk�.vV�)���x�!�d��00b���J=nY����U0�!��6C���l� �� ���$�!�d��"-�ixk�<���ʅ��+	�!�d���̺��
X�����CJ�"}!�d��G�U��}����-�!���o{�e�$]�d���1�wb!�� ��2�2R�`D�m;�]-@_!�Ę�D~�1�t$Ϋ �>�{�Ãw[!����Mp��>#�
<i2%°l�!�����`��7�$0� ��2t�!�ć���2*�B�l}"� �,�!��=F��n��Ҷ׊F�!�$ӽSq6�x�%%au|�o\/X�!���
s�� X�nQ�� ��-�#!�D��;.��q�#�4����"W!!��͏��+S�P�|��кBQ%R7!�d�����A�m�{�ݻ`��&!��rC��C"J�j^6ps��6`6!��@���5 )�����K�y�!�Dޙr*���&�m}h�����!
�!�-u��ar�[5:>���d�D$]	!򤘩~��l��`�!����7��!�!��~�8á,I�x(q�G#�!�D�y�hcB�ޅc��	b3 �4�!�$=�4�x��$�B�N-i�!�D�E�!���E����2�R�7�!�dB� ]Ri��GC�4 UB��K�h�!�� ��aY�X����H5� �10"O���A,M�x�x�O��2�v���"O��W�	-m���^i�N�2"O �bQȃcY˃��gf�x�"O����T*�^�5�`T� �'��'or�'}�'��'	��'@&�y�@8� U�
O��N���'8"�'���'o��'�R�'��'jMe�L�0��o��K[�� ��'���'���'f��'r��'W�'���N�.@~��p�6�#V�'��'���'��'��'d��'��t�$��hk� K���-~Pሳ�'U�'���'"�'_�'R�'g.�B�_�^��A��49�ae�'��'�R�'�b�'��'*�'���Ӽ�ⱡw�k��S�'_b�'�b�'u��'�R�'FB�'jV�1!N�vw��I6��+��lSd�'���'c�'S��'S��'���'�V ��Dޮ�B��0�̈O�e��'���'x"�'�"�'R�'��'������.-np
�G+Q���2�' �'c��'�R�';��'���'.d�P��C�k�Y�0�*$�"3�'3��'xb�'�b�'$R�'���'=����"
�{r�@)�ǎ%I~A���'2��'b��'Or�'d��'C"�'<�e�B�K�%���M 2 � 1Q�'���'�R�'"��'M"�m�����OR��DR&��q��#0Pt�u'Mxy��'��)�3?iU�iK0�RE�!)0b@��EL�`r��7� ���d�צ��?��<���\qp��QaW�^�l�@!�[�)������?�vd��M{�OB����N?E�oA5ձ�̀2x���J0��򟬗'T�>=i0L�+q[6 P�� +J6�)�(���M���F���Ob�7=���%)�S9�H�e-��젘�4%�O��Dk��ק�Oa��v�i���f�(�:"��@ ��z��l��+��r���=ͧ�?y�:F[�I���o���D P�<i,O��O�ul�`�b��N�:��m�4D��pЉ�P�3������I�<��O��JP-j}R�{e��G�&�Bќ���I$ڈmH�b&�S�$�Z1��l�t�Q�D��79����_��IUy������d�=(��$�!��2��@�GĴ9���㦥{b`>?��i'�O�o�}���I�u�<�A2�T�*�$�O�d�OX�ↀu�����d�ꟾ �A5u�eCL�_|~����������4�V�d�O���O���Iu
[槓�V�}�t&�'#�\�h��6H43��'����'�Hl0g �m�V��# �t�Ԍ �-�>������O
ְz�bT���P	 �}�,��bަ0]Fъ�]��� ���x�+e�	Hyҫ[�9nN���h+{GJ�I��Y��0>Q0�iK�<B��'��xx�!�!8���nY�f� �1�'	7�0�I����O���OT��n��TA@�Bpj� x�� ȑoɉ��6�7?Y O>_���Z��ߥ���l]2�&<q����w�D�I�L�I��(��˟���P�ו)�>DC�I7t� =�eE�/�?����?�'�v��OP�6�4�$6e1�uX���\���7��(pJ1O����<�r��6�M��O�`�#9���3�J[x,��U��X�Rh���!�&�OV��?I��?���be����O�.
��4�`݌
�,����?(O��oڈV������D��D��k[�D9cr�*d�����y��'����?����S��.�|���B��$%2��oVH����g�_2�ha��W�擑>"��L�	�yrL	C��o��kP����!�I����	���)��ry�v�N�q���aNX�F펍v6.�Z5�N�gX��2�V���M}r�'��Q��QA�>dPC�H�	S� *%�঍�'>�t��?A� U���7�(� 	�Ŗ��X�;�d���'�"�''��'���'��S�lc���pl��C�,@S��d���4q_T�����?��䧂?�F��yGj� Cӌq �_�Y�aj�٢d�2�'Uɧ�O�S�i7��@�k���8���H���#&���t�Z�)�'�'(�i>���4�H�bk.6JPq�0�F�n��ȟ��	˟(�'o(6���^���O��D�{&�=��P�m���Y`kH�F���lA�O2���O��O��:���?r�� r "���������C�����&擝�"��џ�*PI� Gb�4!�%W��M�%��t�	؟���ߟ�F���'��$CA�0q��E�ŋ`R����'5r7-�q�.��OmZN�Ӽ#D)�[��0��J��E��,H���<���?��8��4��Dб%)c��A<�1��9?�|u�iJ0]|���G.��<�'�?����?����?ARG�&>�R4�6o��.�fu�FW���DS�52 ��ן���ݟD'?�	�R^tA.�*��Y��(,^o�@¬O���2�)�SJ&� �GĀ2b脽�!oC�Gg�8a&@	{A�	�'`EYs�������|BT�H[����5�F+^>����W���$���\�I˟�ty�Ik��ܱF�Ob���ƉJe0�q�hBt�V2O@hlZF�'���h�I�̠��1����N �.T:�
^)J"��m�A~r�D>x'����Nܧ���  L(�c����UF�>j��L�=O����O~���OJ�D�O��?e�� Z�^�I�+��M`�A��I��۴y�h�,O: m�x�ɥnN���e�Bh̴Å�[�yxU&���I��S�e:��lf~b������#wP�|HFU�7c@�b���YRjHy?	H>9-O ���O��$�O,9:%�S?�(��kQ$N^��G��OD���<��i��cZ���H�D�z���
��hr�n�<��WE}��'4��|ʟ2P��n�$/��� �>5�0�J�l���5)^
(���C*O�)]$�?�W/ �D$(���ɦ��\벴:E�	�h�D�O �d�O����<9f�i@4`���-;��4se�G�<��͓�p,r�'S 6�!�4����'��C*D�U�&A����BԡA�b�'זm�t�i��ɑ �rŲ�ٟ���Ћ�)��BIɅ@[W��͓���O����Oh��O���|�"e;=����C�@�\dAC���&�K%wB�'c��d�'p6=�\���A�X�c�H@v�q��OD�b>f���͓SĊxPEh��[>��AE)܊o��ΓU��I�ţ�Oȭ�L>�-O.��O�h	�a��in�����'@��!��F�O���OT���<I�ip~\Q��'�b�'�Ё[�e1o, ���8 ���B��p}��'�B�|b�ʗRͨ��߁[#�LE�����tPu��|1�fp��|�����j�;F�ʿ�D3�9^C�ɮq�t�j4%X�|M֤�a�����[޴^}ƨa/OFyo�~�Ӽ�%ǚgLmpag��l�|�����<q��?���w�}��4��D�1(����O��[��к��@�Z���|b[�8�I����I���I���+�BR,O�<%��������P��vyB�f�f�{U`�O����O����Ɖ{���c�%O��0�.��?�Ph�'�'kɧ�OĘL��q�l��F/txH�@�\�8�)�S��!�I�s�\�	IyrH��S���Va�6d����q��,`��'��'��O�� �MS�[0�?q�-X+'^41ō,_�b�0d�Α�?�2�i��O�x�'�b�'�"�\5o� a$ń! �\���V����i��I/Z:pt(g����2$H_�RaT��@�
/�H�R�w�P��	�pe<�� -*ז<"��R�F�8��'��Lp�*%Pԙ?�J�4��'�P٩�-�;�$h.zʲ,�bOS����,�i>I��L�ݦ��'N���cY�c����%@]$����B>=-�e�������O��$�O`��|���ψ�WO.�P�X[���$�O�ʓD'��Ʌ/�2�'2\>���ؼ|��]À��)���#�6?yVR���	ݟ�'��'@����Njd�����lS�=�) gF�	#��=��i>=9R�'q��&�����
%t�,�z�͖�On���@��֟ �����Iܟb>��'%(7� -iv���'��J���h��GB��t�<9ǰi9�O���'�b,Ԃ��]�Π@^��Y#�� "��'����i����y�T�c�On�'R�	��f����E+�nG+9�Xh����O����O��$�OB��|.U�����,��l��aks��l�d�YܴN� a���?���'�?�P��y��ƸwVtږ!Z�)�fl�6ib�'�ɧ�O�z�;��i���D�QX���LS�QP��G)c�$	b��	� ��O�ʓ�?��KT>D�F@1G��RO��y\�X{��?����?Y/O�l��NЙ�����	�ʍ�q�[�ez�2"�v]�?a�P���I���&��B��SyNhh��
�"vT.!�%�+?�@'2 %�BݴИOIw?��mY�5`d.��k��<��E�_�8�*��?A���?��h��������^� dFS&�X�$W������D�I��M�M>���s��Evvy#��<)�\��Ƅ��<Q��?���?R��ش��$J$7c�5��O��,ITJHx�r�Q��4�N%�0�|�[��������I柄�I���#g�O�:6ĹK��}�īB+�ry2�qӨ�ye`�O��$�Oړ��ɪqp��V�p,�$:3����X�'�"�'ɧ�O�hT�ӥQ+@���s(�^(��YզT���OTHᱤE+�?i��0��<��ۀʨ���ȀX�nĠ�D�#��D�O.�D�O�I�<��iR�Py4�'�	���1/&���H�/&Y�Me�'��7�%�������Or���OH|�fOV+��<F�W=QA�A�����"7- ?I�ҋ^���+�����х�}��t(׉[�~�����q�|��ϟ��	����Iϟ8��䓧s�X4�cҗ^-�m�u�B��?!���?ɷ�i��T�O�b�`���O:�T��}�ite��i(����d�O˓j6�,xܴ�����[�ҹBC�E�Fn*!i��R�&f��E#��?A�;�d�<�"�ݐ@Z���͒]gJP�flϪ�O�l�0 y�'j�\>�PBl٨�����cY�s!tmp��!?'Z���Iן�&��'q���S��@!p����jTI��q Wn����U �	2��4�>���#��OZ)
B�����2k��~�z8�0C�A<ǼiS�):�ʟW�bQ%@�2<DD�0�
)C5剅�Mk��@�>�B�^]r.Ҕh��T<�#���?�(\��M��O�����4��^�� ��i�j�_���ioV�iF�� >OR��?����?����?����I�?ib��$�ʒ ��L{R�B�Ij��nZ�;܆L�'r����'�7=��� ��j���������#�+]B�'Bɧ�O����R�i��d�s�>A��N�$[g40dZ�}<�D�@��yI4�O�ʓ��d�5sdqQGm�&R����hR�Q4ax�Oc�f|0e�<��?	��Zb���� Y�"�b��鹋�>Y���?IJ>a5l	�iFUؑ��S(1���k~�#YNhC��iPȓ��0�'��aݔx��9�܀HQ�U�`ł�H8��'
b�'v��SƟ$i�*�XĈ YW��54F�� �Bџ���4@o6Q����?��i'�O�N����!��@��F9��{UoT�t��$�O����O�p�hq�B�+��ջš�?���,�2����-X T+��LY�	myB�'�b�'���'[�-��n}��6��q�woW��i�oZ/>���I���X�s��"T.nV� B�ߧŰ� �������O~��$��F��QB�g%|*��n�k���r�%Q��I�5��US�'�i$�X�'f�����Y��1x��U_֦���'��'3����D[��Aߴ:X&q#�o�\��vn�/pY����.2��%�fڛ����y}��'���'�Z г�_���]Y"�ګ��\��� 5C�V��Rs��(�4�����aQ��W�0�� �N�{J�;O~��O����O����O�?]��M�z����k�&U�
�10�����	ȟ@cߴ@μ|ͧ�?!a�i��'�5%�A�^ �rT�ŕ|�FÁ�|R�']�O��Ah��ip�i�]�T(�D��C)�)F����IJFL���>9��'E�	�����㟰�	�N�$UZ�Ax�؜yA��O�X�	�0�'ϲ7�P�L�|�d�O��d�|^ұ�Hԙ@�j�q�����?���՟��	z�)�d�)�8��#"�L�jf̗"K�P�
�Û4-"&5��D����dj��|��!O&E�5ȀV� �HI�J���'���'���dU�tڴr����@B&���,�l|�!
��׹�?���&�Ăs}�'/�0��JW�<��dom�6�:��'R�[؛V��T�2�յ�q���1�'��s������!$cT�s@7O�ʓ�?���?��?a����%<Z�����Q)�pj2լ-�b@oڮv��8�'������'�7=��h�CfLu!V 8�)�
5�� a��O��d$����|7i���&��
�PX�F��D�� �r�g����Eh�$8�$�<�'�?�g"�8�� D�6)��@�A����?q��?i����d ��	b4C[ڟT����L�W�Х'�"Ј'K�aR����f�e��3���ݟP�?@�@���Ӈ��@Wd�`��`~�8:9JD���C>H�O7NP�	>�G" R�y'*�)8Њ ��-N2R�'�R�'���SƟ\�3�Y�:�uF/����(�r��$u�<��e�O��QѦ1�?ͻ>Ê�����wܜiQc�[�Dϓ�?y)Ol�iӬ�5�ԅ��nៀ�0�c�$Qf*���E�>�.��F�±�䓿���O�d�O���O��D�8<в=#v��F�B#��m��ʓ&���I�)���'�����'@�45a�n��!g���B ��%�>���?�M>�|5��/�T=3ք���$	��m0hII#T�򤂷��-1�U1��O��DĄ��E:�츰*C*v �h��?���?!��|�*O��o��P,�Ʉ�pم�އfLzd��KI�	�M��e�>)��?��}��Z����HX��D�e���gÈ4�M#�O��z7�^��Ҏ���w>B$p�,
U���r��g��ű�'���'���'$�'O����`AHzh��V�f �ti�O��$�Ox�lZ&A�,�Sџ��ش��o��`7G4�̋b�e��@�N>���?ͧ?~)�ڴ�����L��jm���ź"��+��F�A�*��׶������O����O`�dE�aa�,˴·9z����le����?)O��lZ�N����Iɟ���K��h���0���N_pTc$��2��DHp}"�'�O�S:�D�9�'[�Q��4�%�>�V!�3OT2W�d���Qay�O�X=��6G��' ����.�/$�ܼ���/(CM��'�R�'P"���OA�I�MS�@�bQTsӅ�U�]� @��>���?A��i�O`T�'�lڇFB0L�W�P/MA���P�N�AA�'���t�i��i�%�̐�?Ղ�Z��)�%�6Ѵ�6�c�����~M�vy��',b�'���'�2P>�R'������kY�E����M�'��0�?���?L~���dݛ�w\�V�]�[�( �Cm
�jڈE��'u��|���UZ��6:O���_�l��	q��>;b�PHw4O����ܐ�~"�|r^��ٟ�ە��Q��t�Ȧ,����!����I����	xy��|�:L�c$�O��d�OD����ӜV;2H`D�U(��8���4���O���'>��'��'�v!KWR&UH��J��߄3l���O�|ї���#8�kR�:���?9R��O�*��]n�u�#܀5aBf��Op���O����O^�}j��> �ҥH�1����;��(�����_t�B�'H7�#�i޵���\��E򰈈�bux�S�i���ITyB��	������+6�1����&� n�����r墰�Ӝyh��?��<����?����?i��?iPŚj�h�0^'�0 ����ۦ!ZǠ����I̟�&?��	�BZ8��M�z����W�qíO"��8�)�S�I۲ i��/�=I�K�B�D���-]�F�l͕'�
91fG��t���|rV�8�Ie��q���R-YБ������L��؟�SXy��n�|�gM�ORU�2�K��0���GB�����i�O��oZF��+������'�,���BD. 2HmCc�E�a�b {U�U�曟d�a��$J����^������������a��3��F�r�(��ҟ��IƟ��	͟��23h�72Hx[�]�t~�xـDb��'�2
gӾ��8���D��&��g��(H&��S*|��M�%�k�	��L�i>�BF��Ц��u'�iƊE�b@�>	���^�I(~�r��W��Ƒ��I�fZU�gDʲb�V����U���gU.dr���'�R�^�ΐj`�L/S	��REk-$��`�vj�<�$$�V'D�v�<�[�&w�l��nE�vC(��<Q��J�(D6E2l�<S�}��@�u+���"�S�'����e۳i�,���#H?$^ 5��Ӵq��;�O��a�$+B"F�[  �qg�W8w֐Ss��H��F�NIz��!0�"�����%I�oh�D0��Z/f���	� `�$9�&1�S͇|�s���,5�0�1��"���b`үANY+�*�Ӧ��	ӟH���?E`rj�'{ j�(@����r�/�����?���'H���ӟ䘚dg�4��s�@ #��&Y��#�K]��M���?i��ʇP��X���$�&�D3N���I�:��6-�O���P	#����;�)�ӹ.N�@��u,*���p�6�T�o3�|m�՟���ǟ���#����<��%�?e��Xe�7=��@#��Ƨ^�6�Z:��O��?���2I�ȉ�+��b��G�E9	/�\ٴ�?Q��?�uL�/#��Ky��'|�$C�%8bx�&n:X�\��f蛦�|#08�� ���O��D	h�,�Ҏ�#�T��
Q�\^�o�埐�rE�+���<)������`��.�@�$��	,�`�)��Bf}"���e�"]��	���ty�B
�CS�q23 ���4X�v-Y }3�I�>�-O��7���O����^KR�s �T?�B��%@��x\Z#b5��O��$�OJ�l`���F9�n<30�ԛ9^TkD%�'m�Xt�d�i�	ß�'���Iß��&Xg?)q��',�\��u���ͻ&�m}��'*��'�剽j��4*��J��ҧ=��I�Ԫ�bv�AI��[�@�nZӟ�%���	ӟ��%e�@�7�� "Xp����ʇ�n�p�n�ԟH��|yY���'�?����"(��L�UM��m���
7}�'"�'ܱX����?� �Ǥ8��H�@�� |,�*�ho�b�v@���W�i�R�'�B�O6,��Ck��!�:��gi�,H 6	K�٦��	� �`�g���O� �$�ؔ0f�A4`�;�b0:�4�#$�i]R�'���Ol�O�I�$�!�#��2r�O��`$lZ����	ퟬ%���<��s����U�ܭ  �	�ц�!	������i��'>"��S��O�I�O2�ɗA�9�4H� j��I��\�6-�O�O�%��yr�'��'���/R5q,��s�	$xs�%�Q�i�����kw~<%����$��
h*X�zE���V`ڔ�ē�?	J>�,��D�OVŚ�	�o��0q��w>c�@6r�b��?A����'	��O�	00���F0�sQ���ꬻ�i��-)�y2�'���˟��&B�}�D��L�,�8&%�/B%NxZ�*�ަ��	ş`�?������^�0���"�.*Ȝ�b�_M���
5���?�.Ot��D���'�?�EeJ�rT�H8��[^� �'O� m
�F�d�OJ˓!_�$��)F�٤)T�%�a��.H�P�@�t�p���<	��Z++���d�O��Ƹ���GI�}�,i7�]`�X���x��'��ə@�l"<��gj*i��|�q)b��-G
��'�R���k��'�r�'��TQ��]jwN,vF��l)��SC��#O�7��O�ʓ}Y�FxJ|2qg�l��sU���=��	���-8�˟�	�����?����I�-��4�eKl�%�Q�N��'�훌����O�4ڰ�=+��MJ�J��v[$�����-�������0�@N<ͧ�?q�E����t��]��Š&�R]��i���'剜��I�|B��~#]�m��1�`�:2M0E�$?��7-�O���"b�<�F^?-�?���TI.���ďU��&.Zxȉ'U�}��OP�D�O�ĺ<I��)m.��HRG0a��p�s,�=�p��ђxB�'w�'H�Iݟ���j�p0��Ö(��;!��� ��n�Д'��'�RS�<�e�֭���ㅎdE~9�rJSv�&�ڴ��M�)Ox�D�<����?��tɐ�ϓ�<J#-�,Q��OW(r���c�V���	����Isy�h^�J?���?A#'�Bi��&�F��@�<u����'���ǟ���˟X2�nn�p�Iz?� �-+h�����9fM����Ѧ������'lBT��f�~���?a��KP�L�6$M�4p9ڐ�[����S����Ɵ���0C0��'��$�?uidi��$���hƂ-�޵�e�q�.˓3<Xh�¾i��'�r�O���ӺC��-Ek>\{*�/|�����q��ǟ\xp�2?�*Ot�>�2��f�ĵ��g*C��{�arӮ��ƌC����I��p���?��O��C}� 0�ӅI��H|��7umlL	�iu����'��؟����E����`�
4� ���P�+~��`�i��'�r.��������O�ION��'B�Ow�0�r��qD�7M�O@�aǐ��S���'���'NN$�T��4m�C��ʷw�r�ەp�(���sibP�'��	�'�Zc�hL;f*ׇ;d�Ecg�N�[�����O��1�>O���?A��?�+O  �T�2E��SH	6NgZA`u�٪3���'B���0�'C��'��G��Z�`�sb��*2�Pc��cc�5a�'��'�"�'��^�АT�آ���S3T��3�Eڃ7���S վ�M+.O����<!���?y�;*� �'ߔ@�ᆒs���2i� ��5��4�?���?y���D�	*ET�O�R �	��krŢ8�v��
?8
7�O���?����?����<A-��vΛ����Tb��@h(Dí�M���?�)O�i �͟K�4�'��OZ葓�ўzs��p42���@�>����?��e=BPDxrݟ��c�%�m ژ��I@�S͒	{5�im剅J%hap�4�?)���?1�'p��i�i�"�8�L%��k���^5y&�sӆ���O^�"�5O�p��y��I�gF�����C�[�,�RI���f"	9RI�7��O��D�O,�)Vz}�U��3rH�-:�	@�B*yF�5��Î�M�����<QM>���$�'���p�"�OI
�ۃ�]&��y� k�>�$�O���Ȳ|��i�'I�	ɟ��}2V/�i�P[B�8a�Tm�� �'r�Z�����OV���O0#Ҏ�	6����߳S���'�ܦ���5� `�O���?�(O����FMQ��M�,��0���2�.���[��(i���'�r�')V��q�M@(��¥C9B��9Y���-Q�T��O�˓�?1,O����O��0i�,�p!��Y;T�9��7#�|�k�>O@��O����OJ��<� -0+���){.�t�1��m�4�a����A��_����gy��'?��'��dk�'�\0� ��ǒ-����"Nuƽ��`hӢ���O���Oʓ3���*�^?�i�a����gv����.V`�`�Y�gpӒ���<����?A�%e���Oy�6�1����)����ULV��V�'�2U�,�t!���i�Oj�d�X����8��}HƢQ�3���gf�`}��'��'qNUj�'��s����&�U*��k��:��+w�Ąl�DyR���^7��O4��O���k}Zw�������D���5 �|�l=��4�?i�Bz�|�d1�s���}*#�ʙ��ģWF��*������BC�?�M���?A���"�'�?����?qs��Q�>Аb)&*^� ���1��V�T�S�U���������$�]j)�h�7xJH��#)ʽ?�nunZ�� �I�D��G���d�<���~Bě�fF��S)=��)&C<����<���U~�O���'�r��$&aΑ�".I��epqaB�@6�O�Q���c}RP����[yB�5&/[�l@�J�e�:Pd��T������c���OT�d�O,�$�|ΓX�X���3<��T��~����s���fy2�'������П �e�|�Ь���pMU�C�b�I����I��l��ן��'^�[�p>��m�;�&�9cB4w�m8֠oӤ˓�?�(O���O��D�(S��ڴ�0��R�Ѣ~QY�E�	$��'���'�2Y��h7���	�O2�����GY�����}�@P��-�����Vy�'���'��t��'(��'������,b	�%�6�F=F�j8� �p�R�D�O�˓�� �P?����d�&����
R.M�@`"׻� �ˮOp�$�O��	�NI�|Γ���o\?i�X;�/��!ʀ%9ӂ�&�M�)O~0il٦��i�7��O�i�Y}Zw���e��5s?a�b���5l�9��4�?��S�V̓f��s�l�}�5mP1|���B�=�Y���H�e�/��M���?1���RX�ܗ'��C��N2�C��Ɍ#�@q ef�8�!�=O��<Y����'�l1���Ė�D�1ǥ�%�*�A#�oӒ���O��d��*i���'�������3�(��Ъ>��x
��k@rUlZß�'����i�O"���O(!5�O� E�1+�-�*Լ��W������ɒa�eH�On��?Q(Ol���Z<����,j�.tXS�K"}���QgW�D@�$e���'@��'>�_����0�|rUN��6C&��Ǎ!0g	ҩO�ʓ�?�,O����O��$́ H<��am_�f�T����޽Y���E6O��d�O��d�O����<1��R02��R��̙�$M5��(uؙbЛ�R����my��'���'���'*�|��E2X��ɹq�X�V<�-���s�����O6�D�OXʓy�0��A��\c����>Y�q��C�Q�ݴ�?IO>���?�s"��?�K��EM]�HL�wl�G��x�'w�����O�˓� ������'�DL��!�ޝ�ǀyH0�IG�A:WO����O�1@�3O��O���G$`���S�d�.)!WL�R��6ͨ<	�D�
���	�~����j�����V����BXIa)�����!)kӈ�$�Oh��R3O.�O.�>	�W*Z3`aB"�b)6�C$�hӠ�:����q�	ʟ��	�?�M<��P���4dF9JUv��k�o����$�i56��U�'��'��4�Ԑ�D����� ;�n��\RHd$g�0���Of��Ė9�r�$���	џ��C��p	�U�)���lܻ5b�l�Q�	$8�bI|*��?��� \�uS�ͻ#J�������
*0�%�i�r�F�8@�OV���O��Ok� ������8��%Qć��*ι�R��y��c�X�'>B�'�rU�,����Y�A1�a-И��*=��Y�M<���?9N>��?)��Ӌ>:�Y�$n	+]R�+�K��\hhX����OX�d�O"˓Ǡ���6��|��	ۍ
Ė4"�P�h��-��U�@��ȟ '�D��ȟ��D�>a�G�� {|*$�R�*^)ck�X}��'�B�'B�3k����O|��ɂ}���YF&�>G�r���ĉ-囦�'��'Z��'����'#�,O �iaC��Z���[�	��EoZ����	qy�S'x����d� ����4y����{��\z ��o�	͟��	�-�*��I@�	["`&[ez~m�e*E�\�� ��a�'︔��#t��|�O���O�D��.,�UH���r��(O�j�m�ş,��2#X2�Il�Pܧel�sb��Ny>A��`�	m��8o�^����4�?���?y��j3�'i��B3ĽI���"q�X���
��6�<c���D.�D&�S�8��+쌬A'�=�ʩ�I
��M��?��i%�MÔxb�'��O�11p��"� �d� f�L���i �'���%(�	�Oz��Oܱ�*�2X����A�n�Z�+U��Ц���0�2ٓ�}��'�ɧ5��ܗ:���D,\'tT�u�%�$����_�8�$�<���?!����<%���'��Ho��[b�A6>0N=@C�Em���O�����4(�jEfg�"�S5sS�C��Wk��������Ĕ'��H$am>iҶ��t��"���.F�����*�d�O��O��D�O^9�֊�O��!�L�gB�]�[AEt4���{}�'��R����>W��i��Ο��:�tȣ��e2�E �(��h�۴�?!K>������}�'���DS�*�d�&u��I
۴�?�������/Z��%>m���?���*�(��Y1�n��upu����;�ē�?�
�<z֙�SjM�!|�X�T�K!ڔn�zy���2R��6��`���'�� +?�4��tyD��w��h�)J^ۦ���H��\���'�Ґ��M�k x���NmӔ`!ᄉڦ1�I������?�JK<I��I>�͹��U =����֯]�H;�ɁǺig���6���,��F�4k�D�0���r�~ aC�ˏ�M�����D�q\�S�����F0�f�d(ޡ>p ��F�ܿ@��)�<9��%?Z�O����ΣvX�ɦ{�x-XV�#�Έ��e
�J�xB䉷+�
���� 4
qJS�H�pr���C�C����"��ն�Z0�(%Ǡ8k�,�4b���rZ�8x���yl�E�W�<@���'��=�y��\s	qb��+*�9����g/�lB��WO�X�BE2d3�����+nu6����(7x<�#w� }��摟?�4m����HSP2�GB�wld��%��H:� ��N�E�J�����?	��0�?9���?���?�L>i$#��\��@�n|B���\8�Xks
ފnp�=���-=��d\LVX$� �ߩ�FYce/�0I�x��0�?I��B�����NaԦ�8-�y֥��T�f�	П���T���O!�T)�Ƅ=@������sOj���'��6�ɾH�dY��l�(xG��J���p�J�o�ay�ȽO=���?9.�8� ��O��a��j)b1ڢ"O��B!Pdh�O�$7^ 8���U�l% W�Ɵ�'��)V
v��}��,Ψ5#8*dkف{�y��	���09fPCș$�H��iK#��4��@��BR�m�v�>�Fυ�$�I|�O�bJ�v��� )U�$���yr��6�d�����ăĐ&�ў�S	�HOv�����	���4LķZm� �@�Φ��������dl �j͟���|�i޵R��;�Ѓ��)P�F!p+܀���rE���?�7�
�5ق��|&�᥉ܥ;�0	���Q���a!N�m�Xɳ ���?�vjK�P�>�k���F��Ę�B8���c$�Iw�p�g�U���$,?٠�ȟ�T�'�44����.�<`���-��)��'ܚ�p"!E{������U=���'8B$%��|B����� �<Ɉc�IF��2�([�	҈=$��F�����O"���O>ɮ;�?1�����ŝ�>=LMe��)`�(�hѪ;�b!� ٌf����=lO�:̒�F�r���O�z4n9p�MDd��iE�3=�$��퉿#��i&AC3M����6$����OP�D8���'Krȡs+ɥY&��m�	<��3�'�L��C��3�.�XUo�i�B��y��sӦ�d�<� ���F�'� �4\�`�A��H<sV�HRV��'���r��'hb3�"��'��'���$��sz4)x�U;���;�=�.}�?!@�P�:��(��'�V5��R8���s��O��$�<��/��W� ��7�ջ <i�f��<q���?i���ٗC�`����^9<��5dH�!�D�WM;���CRkA
k�D�c��"\��v	ȵ�M���?	,��s���O�������@B���U1"cN�E#�O��$FD1��""IC�|2)���{寋,k/��X��ϗG�Z=7�>Q3�ƃ�L	�O>�� Bm�'�Ǘ�Z|i1K�-\Ժh ��>��bş��I���IJ��8���'�G`N�%1�J�Uuء�<I����<	��]�g�(�J`���Fr�*���H��X��d��4lBR�ϸ1�d�E`I	�TYoZƟ��	៴1�
؆#�:\�	��H�Iߟ�ݬ�PY�5+���������Xg���I!��}��.�l�t��ɡ>�S����̼w(�WZB��0�ݫ&�����L3s�|HB���#xY�%ӛ'��hh�(U!F���	&��3 �����'DB7��O(�z �Oq��	��ٔ�:#����F�~�ԕ��nU��\$��z��˔P_���׼Mt\a!��c������M{�i[�'x<�%�O��I V�	C͟x5� �k�/M�B�I>B����ꜿ6r+r價-�C�ɂT��q4���7:X� l�J��B�	���,���J0HC%�̟e��B�=K|�`��%�-�$�
 ��k�zB�I�lv��
�!�;%B�qa��C�	"+D2ղp̎�d��1�^����0D�Ģ�ԔDR� pAΎ�.����/D����cɭt��,ZS�R�u��ؖ�.D�8@��zlL	JQ�W�aPg�-D����tޖp�#� :�䓕�!D�$ȲbļA�pY��B6^\��[�:D� J5k�
��=8O�J����9D�t���ܓ^�=ط���4�Ȍ9'd5D���k�`��)�f8�����&D��#�b�c��|AF�L,���7D��)ްi� #�ےQVjp���5D�,���ۅ.�h�ٶN 89�a�s�=D��CW>k�@�X�Z?��*��=D�4��d5�D�g�էxĝ���:D��X��%#0P���$���b�7D�L�@J?=�4��@�t�pP�l8D��X�#�	U�a+vIʼT��T: �5D�4�تA��q��.Q�T��n0D��mՌn���2.	4�D��/D��cq�[GV�%3
*r �	��)D�4�TO
�[�r��i� TXsA*D�K7�J�<$�2��Z�vK�@ꃁ&D�0���PqXDB�kYN�6�Y'M#D�p�l	�O3`	u��2|>,x�L6D�@�eG&f��Dq'MǍw,���g1D��r�gV�x�V9�eǔ8^P���
+D���D��:���褋�%}��'$D�drT�ϷB�Q��ɋQA�()!D�p"�eM�s�n�v�I/1�`�=J�1�-� ̲�V3^VŨT
�>��Yv�"��ӎiV�� �ג2k�m���E-6D,C��/���F� 5 bD�V��C�6�����Q�yRi�g�l�4̎BbȨa��<�y���*@�4��q������I�Zae������1-喕+A��Zd^B�	߷\�!�d8�L��W��	�<��w��@]qO��{D�W��0<��']̸��e�zYP�cS�Tg(<I���7g� L�V��Tu�T��ij:]3�#���_5���g�\j�u( l/|OVb���o�<J���X2HA0�X1��(D���2&�w���j-v�ek�)"D�<�e��9i�tآjP�C8D�?D����n����@�+�"\� DْK=D���C�f��!C��L� g	��9D��*� 5���8�D	��Y��c*D��آ� L-��*�==��" f(D���2,�8|�S7	��d�1X�-&D�����I?K%������"q  D���f�\���G�(�T��g=D�� �<���T=�Z-��G.9����"O|ة��\!��P�
6Ԙ��"O���q���2qA#�Jۍ+��}�"O���R��p	Ǜ=��L��'yh���"�	�q�2�AAG�'	o^|S#撥P��C��=����ڝM�Xh�����s�^��?�4��$���)�矘Q nR�j��be#�c�D��H0D���m��:n5�g�L0'0�TIc�l�H�'�F;��f�.a���	c�f��k�O�ޡѰGĸ)�l����}��Ls�4g�v��٫� D*£i����bӘ,ԈC�ɦ/K]@hn�]ӕO �*#<�WmR�ߖ7�U�S��� �,�ऑ���-C�D5����y���->4�S3�ɵ6w8�P�����Gk�ߦ�V����s�P��%Sd�Хp��&]�HiJ�!D�����S-PP����UhR�s1 k�� �-a�6
L�p&@�ታ_l��s�LPhx׍�}#���Dӛ.���ݴ[d�A� 6��͸�M�E.:��f����B����dPza혋�r�R�CD�0"<I�`&/�����3/���|��HE�<t`;�,^�{7r�ɒ(@�<	����6]b@Y���$�Թχ��Ij�-6�iݱ�P�JN�� �ޥc����(D+ظ"�Z�<���	��m���&f��:U%C�<�b̈́�N⟌ِ��K�=�D|xTf���fHX ��@ԧ�V�se��	��RK�Ov��(��-�3<6�t��.O.�>9i1�i��A���V�N���Gm�g�&,Y(�:b��3 v��S�[�d$��yPBթq�PqbC((�D%��K�$��7���k��G�Y[�ab@άٸ�Ц�A�>T�$�!g&a���(��;�|J�E���y��XL	��Ԏ$�������?��(д{H�J�����4H9
%��O�S,1�>48#�<j>^}`�ÉxQ��<a�ө8���S�s�̡��%��'`�Q	�dZ�`�8Up���� �4������'~�S�*9`��I %�����"��5�U�b �ݸ�E Ux�ij"��^4)�έ;�� P��h>�O��'ZCt�z�Nŵ��T;s,V�Q��|%�T9w$F��}�1LW�jT])��8�"BM:�H_!آU�(��$��)�%,��3	��O��}��+Ϡ�(cJ«lrcG�Q�e!����r&$���(6��ʧ*K9@�w�ZyaP쏳H�|����$z����FE�9�������=apj	�_�B�B	��0ӧ��Ԙ'{�2ׯ��'��A�Aa$*����	V���9��і�V)��)��y���FV(��'in��b�3c Ijd��w���W�Ԡ01���V��r�Y�;�E5��'��S�P�^aȧ�����աOe�x�O���ѩ_7%}x4A��<Jj�����9-|�g�@a+�dC�0h1���ʗ>V�'��>���!.���J��P� ̂aO�^����꒮</4	��XvqO�*e<"ͻqY�AP�60�`j����5l��c��|R�����=9rFˠjf����b��@0 WƊ'@1SΚ!B��b�Y��<�6�����\�vuq#C�Rx���� 0%vts'Kɲ-�l@�#N��.G̭ȖF�, �X�N�5~b4�v�̪,���I0R��<���7���P<פHұX���ٳHJ+�t�O�۷@ZMtT�wE�]{��8�d	�	�(�"��I	Ni����	�w2������$�3od˧�Or��P�E�D� 1�ES�R����%%G	O5ZEI��2�4t+�{ʟ���!�w5<x`�㖙R�cC�
����ʓ'V�n�+A���z��{�^�pt�����F���!�1OF���a��	C����y��=Buo�?Zܠ��A���<Aqg��ܡ� �Q��Mm�(@*�d��$���*,�Ƀ�� V�A8��OQc�6�剤���O��U���PS!ԉ(�ʘ�4�FMsT�|��tFLqP�LN�3J���'Ȳ���A��~���d��@�$[z����'~L)�\>1Fx2X=p:܌��`�,ݣ"�\������ݸ�ȰUH�]�S��L��5�4mj`҂�n�]��%ɭu(\Ң��!f��0�B��E���P���2}1Pb���#��%�"�B̓c.�$�*;�)�T��f�m���Q��j�/�#}vֵc��v�����6���ˁ{k���`,���mO�U�9�l�;g,��{�������O�.�bd��؉���8U�Ы!b%yF �&aF����Z���d2(�fuⅉ�E�����ɸ'�V�S�E*�P!qԣU�KW
�I�d���@�R2�Z��p������O����+���	kc+DXh���B_�`�HQʔ��t�FH�=E���M�U��}�W)��������Xm���Z�χ:�	x���/
.��Ҳ�U�5x�|�Q%��wZ���'ΆI�rdR�(�>yd���d�PQ�9���`� �)�ʜ�6,�&$���9�ʀGYd��?A��iC�M�So��s��O~�C���π *9JTmV!o;z�+u̓�K u	0���Uf$�@�h>�W����Ojb�*]a��%{���k&���~�ɏ8\�����D��ቡ_7�4�2`�=$�c��[���q_3o�6�Q��O�ܘ0�ϸ'0�LY����b(jch�6*4�`�PDԼ|:��'��VF�mD}BK�I�D̩ůSk?ɢ �+C'�\��%W��8��枥l���0pJ?���f������:pV��`�y7��#��䢢�Z.#0{���'�0y��<R�x<D�����0�ND�o�r�3d���y���7��d�p"_�Q�����<m�j#**�ӟ.�Q9GK�b҆=��ͷ7������34d"�O��{0���~���'�HI�"a�+e0�]���&@�A(���d?�'ᒭ{�� �VZq������YF,����ȨV3�q� ��*�ȩ�a�Zy��h1�
7N@h�`e�ϸ't԰�CB�<�m3�����/fH}j�E�6cU8�*
�~�H|h�M�U�6��R"Ix�T"`@7%v��A(�OyR��!1�ܕڑ��(��,��L�Ո��E��M#Xw��QH��3����hB�=�}
��ʠ��'��|��ڀh1�-2�b�� 	&�؏y­�E�,� .ܱ>��ɊBř�?Y��J!�B��c��(�ԝ�ĥ�E[,�&�Q�9O͓&Ю�,�c��
s��U�A"�y��E�R��2���y��E�Qw�E�1�۽C�t�%>��7���&}�q������;��X��2<�P
S-��S��#Ok��pUb��@*eغX���$�R�P��	M�<�fU�!3
�H��'�&5�hZ�5��*�+�L� �nռC�1�&gC���4��D_CH�Z7��`��)٠>��`�g�)�&��D�M�y�+�7[�H��<y�#�`H��f�8J�$mr��	p̓�\$�(,4J\{�Rmj��9��a�S����i�TKŦ$�� ��A6Z���S�>��þa4Ŋa��c!�њ�K��l�8�B�A�8���:�M���C��J � I�9��,@������q��B��&����I�5����O�/1�ԭH�ϑu���Z�{���<@��5y@�Ѡ�E
U>���CH��Az��R�$,O|�Տ�"w�]���|X��Z��R�BT�@��r�~��'9B!AP&�/~װ8���]38ΰCS�U(H:!�\�x0��I֛\�p�c��\#d*"Q�pJ6?��H�wF��С�#_�� z.�^� O�$ۗ+��o���s�S�>�H�OR�:E��+K����AJ%���B�)E��x�� C�+��U ��	dax� �݊T�@c�L<⑩�o^�W1��ԥX5H�����+�zy洇�I�$�,={g%�92�&逦�¯s�tJ&�"�7��!�b"扛v�p=���0� (��(e��kc�'��  ������ �nV8-� �",%�X�{���y~bMH6|�8���y�g?y���0hf�DB�x%��z�%�7x7�Q)�'Q@�'HI ���/���je�%�'a���@&n��:�N�)&��Xa�L
e��#�sm���p��|Γ0�2-cG��. �������&a20�64�� �;\I�ib(�pb2,է�O��}k@�Ԝu�2h*�(<���'%�ѐIC�lD���$O�%�sɝ?^��X �E@�Sl�4��*I2|���1ɟ% ��;�Z#L.�3�i>�K��T�2}H#O�oNڽj��D�d��|򢅖ҿ��jZ+��+VnA�5�⸛'mȰ.������"e��>�g�
�dZ�ؐ+8�	��Uo��)E|B)δK v��pA�(�EQ��3g�8ٖg�]��FE�G�<�cH��@B5�M�qnĳ1%C?� �9튍�t+��iI�3����/>�>,x���7*?�eK�ȇ�o�!��Dv��\���FpZ�([GB^m~!���&�"�s�h"e���G�	!!�dѻ5�X)+0��v�F�[��9Y!�Ͽ9��LHA��-B�)CÄ[�B!�$͸~�@���GH�O$" :�Ð�d@!���`u�Z��J�coԀ"ւ�V!�D݂FӘ��1ɛ�,j�:���=p�!򄅲O��2����6WF����P;Wh!򤝀4TP��ǋ:Rtt��o�� �!�ؚ>���3�*
�g�!Rq��6�!��\�1���:!I ���!��)�!�$��<�W,?l@S�J�,r*�u��"O�Y�h�����B�7~�t�q"O�q���� i[Jh��Z	sϐ�HS"O�I�E�4��聃
R;0�VB�"O���ï�36��cI�"vE���"O�a���N�n��X�eЛ,0@���"O��G�ϤUk���/�f��"O��3��q�x��U�)ҷ7!�d01�Ҕ�aZ�6R��+�+Y!�� B��ri-_qԴk7�C�{����C"O҄����r�0��  &����s"O�����6C�n��'�� [��KU"O�  f�I�==L`��Β>/�T��"O*����D�w����d`�2Eu�p��"OD$��&X_�(R �	$?VT�)�"O�eh���!
�4�3(٬Za6���"O%��,�(��I�$�� �C "O|y�4)�]P�3����#Q"O�yb�A+��`�b[ep�uBv"O�3�@R�Fl�����f|��B"O.���G��_f��ף\y�(�aR"OF	P��T[$�S����� "O��*5��B[�k!�80�|m�"O�=�4f !^��Xq`�)xd��	"O�I�u�29�f���m�N�K�"O��'CՄd{�볍S5F��J�"O��*I�O�t�Md��h	"O�-���Rn&����Հq��"OBg	�T�9��ʅtl xD"Od���H��F��0"H dq��:�"O� {���w<�@�)Z)�7"Ox�+v�F9Py��
FςW�f4��"O~��T���w�� #Λ�l� ���"O��h�˄�$	�m{!�07��{a"O��+��܂{��V+� L���W"O��`��6)�X�A�٧))�<�0"O0gG��M(L��
	�
�i�"O���G�XbK*u�0O�1���U"O���E��f���C.�=��uXf"O�x��E���a��,N0�@��u"O<=��,ܛ[�&5�P邺3���c"O|�A���X�D��R"�7�V�4"O>Aja$ȴf�ؐ�k}�@ ��"O@v��B��:a�8q�*'X!�0&~p��
;�����Z(+g!�F�H�М�#���.�8�J̼b�!�$K�K��pO2f�@9�c
f�!�C?f�,5��B`���7C�
�!�B�s$�2&�=۰�����9�!��� rC�(^n1�v�A�1n!��`���
Ӧ�7@N|D����.u_!�$׊Wﶜ�V�Z,A,! �mص
/!��^?<�Rm�	K�;r��-�!�+V<
�����k/8"rL�.!�d�	B�~��A��?)x���˞�!�DB�v����Z.���Ȟ!�3r�Dɑ���1$�����荎[�!��Q�.<����O��Nਵ落|�!���,�ZQ��G�~�fq�ve�AZ!���'�k-�:t��⤣�G>!�]�VO8tУ��(DL�b���G�!�DR�3(�U$-J7�]��`*[�!�ý�h\��/��Rr��,�!�J4#6� �wBX ,Ha-
�q|!�d��>0�#�CU�4,�f�pn!����'zf�A2.]']avPyB�2^!�$JO��v�L�>G1�E`�"�!�$C�7���� ڃ+�&��(a�!�S�(���dm�5R �ъ�
�Q�!�$��@�bFlǌ4�L�)�:i�!�$�-w�rx��߿^վ�s�Hź]m!�d�;d�Q(�Q�tQ�p(�(L�!��=�B�$!Ψl��y����a�!�� ��iV)
H,�8V(��T"O��@r&�	ٜQ1�g�'Fܸa��"O�t˱䘚P��r�_�P�ѳ�"Ov������+ų�$�Z���p�<祖�#4�d!�:>��1�p��i�<Y�CI	/*�\1S��m�$}!�|�<���҃'�1?��zH_B�<�ĩħd�RPA�á��`���{�<I�h�5C20U�g��+d��92�Yv�<YWl��MQH[��T1"��e���o�<iwCV(|F>pӷNV�2��h��mt�<q�@�QZ�s�Ѳ<�n�jp��W�<!EGMjUY�M��F�
�Xn�<�P+X�2~����0NpY��%	p�<�k�op"�1��)т�����c�<��=�	��HL�K/����c�`�<�Չ�@�BE;�h�S�ܡ�`��Z�<��h�7NF��X4j̗Tջ�kT�<�����s�&0�g��k�H�C���L�<���V� �n)��$�2yA�D��eF�'Hў�'+�*I���B�Mf�ib"�M,ҽ��P�:	��,��Ib����fʾb4r}�ȓ,�,Y"�*V�2n2d�0MľM�ܵ�ȓ�LU��	�`; �qc&��1���R���h�ABR6���Sq����m��߭.�NY*���0w�X}��4��𭊌hnV}6-Y�*KjE�ȓ\<�!��#�X�yAT+bg�$�ȓ^��!cJ�$$�Ҭ���*gH��J:�TH�3/� ����+a�N��ȓ	���cX���!J+�م�E� ��󦍨�h ���~�ąȓ/�T<��/�h�L���ȥ<9p(�ȓ:f�<�F߄L.�8�kܦ7�%��w���yՈX�l��|ص"��;X��ȓ0p<��[�����Bƥ^�\}��J-�Y�����&J8���I� ~ e��"%�Wd>+����J�P@����+�[T�÷
R�xqoݯm��ȓ!B�x[FHđW 0q&B�)�pP�ȓYY
qRV$u
0�A�7� =#���s�)�� >>Z���ҬO�,�;�5D��p��3w(�%��3#�<�UK2D���Ӆ�H��M�!��S�tب�f<D���*]�K���c7�Ҍ_,��G=��0|JVH�]IB�Z�B��JB�A�u�<##�o�4����T>P��0Nў"~�	�.� �;2�� �1ǵ!�B�ɷn�n�
�#��OQ�\(�d2 �B�ɛ!�����đ)'� ;�C��C�	�7Xj뗄LU�ܝ#�b��s��C�R<�Q��'v�d�q�jʥmF�C�#ZE�۰�q\�J��ǺB�C�,vɢ�s2�V:�J5�
��
C�	�=���5=���B�eƎ��B�eH�9��b.U���X"ٜr��C�I 7�X��
�~����PƮC�	�8X�A���r~��&���q��C�ɨD�7둖y��eɲŬ	��C�I�T��18�$�ZP����0B�	k�ٚ��k̄����C���B�I�$p��H�!W���uA��-��B�	��=�ì�1M��H0'���B����h:#b�7<�`	�ëO#z��B�)� hE'��!���#��W*Z��\��"O��	K�L����C��&6��"OF���/�4J��*֫N8qr�"Ot���l�*>�@�I��p��� "O��C`Œj3E)���V�B"O:-��O$m�s���(��"O<��R�Y�C봭Pw	 U�=ѐ"O�0d��7`vB5�'�M�d�R "O04Ă̮t�i��KL9Q Є��"O���b�>-�*}�qI$L�PYr"O�!���"-xp-��Cw�l|q6"O,q��&�&7V5���ފȈ�ӥ"Of�ӄ�[?�)��B�E�F`k�"O������Qۦt�C��Esz$s7"OH)L*-\�#4n��pF��zC"O�����6?���F�I�Q�Z"O�G�S�EbJ����^2H���"O*0`iM�o���j4럐[=���@"O�������$����h%�,@"O��6�ÕS�Q��J�G�Iؗ"O&����D���"у��_!Z�z�"OLX�L^�.���w�� 1����s"O*U8#J�l�T �.鶉�U"O&<!Q�ڷi��0�k �@�a�"O�\i��G�ޭS3*G?^��;4"OZ�P��5"l��.&��
�"O�(J���
w�$�$���i��ӥ"O��`⑖e��\����7ۨ8�F"Op<�Bހ9�(��0mW7%�&��'��z�њTz�T��aK����'vt��dI	�v����D�ƃ�4��' h�Ǩ��x�m��{A�y��'��,JT�j��ͰS���S��mY�>a����C�bm�DPAH'R@rDj��7 |!�d�%F�𑂆�ډA�D3'�5�!��;���¢ǘ�m|1c��I��!�d�w�3��mh�gS'}t�	d��h�U&S�;t|�p1���>��Շ)D���"��##Y�e�b����:я3D�Z���~K&i�#�YE����l2D�T����K�Ph�A$��x8�q�0D�H "��0t�X%���e�b<0�c0D�h�P
��_��P�@����[��,D���2�ʵ%��Ѓ3 �4D�� TK*D�lz*��Gr�asM��a�"(O�#=9�A�5�P, �`�Jň��`�<�E}8uSl��H����_�<	�E�Qn��'������X�<1����&M�Pa��E��!c`�V�<�g:�Ԭy1i# �vq��f�<��J�0m3�}�g,�W�x��`C[l�<A���C.����L9�j�\�<��흴>�.��@�C�{�@x�e��Q�<ѕ'W�>���
4�Ά�$� �[L�<���(f����1�Ƞ)5�Ѵ21!�D��m���î-�ȕp��N�=!�DA�{�t `s�;9(�))��^?�!�d[3�ܵ� �۝Q#��P�حr8!�l*8Ȑ�2Aꀑʱ�Y�7!�DL0��9S�$��R��1CVŃ%!�$�;f|<)��_�sx$X�s��")!򤁫B�, 9�!�rsV̳t���!�$E�|��xZ��Y�l��"O��Q`�ݡ*��lk�ثlRf��b"O� �����YM���#@=уS"O�i�q��:Yt�31�]�b��3F"O��Յ Na�s�߂���	"Oj(K�cK��j)��R�n�bY3"O
U�g��1k}�᫴^Ft�x�2"O E���35�&<�sB�FG*�v"O�x�VKL�U���Z��O4|WR�*s"O,�����U�ؘ��AU�<�z�"O����.8V!��|�n<�"O�UQ�Eܷ"d���޼(Ւ<h�"Ot�c����~�6� P�>�J�"O�K�f�sD29ql��nZH�c"OH��`g�h�V2�i)9� �4"O� b@�?]^vdd���t�U"O�-rH�x�1�ܒ	��D��"O�Qx��#_��9K]�~�^Dy�"O�T0'�ƜLP�
ЪZ*��e��"OٚTFO ���"p�@��"O^@Ф�	0p�r@���D&�]�"On�"/�:U��x �`*�Yk�"O�����6~"|�S�ʖln���'"O����֟w�DI�ժA��FMs�"O�I��P ؀��#N���x��"Op̫b�Cwr����	�Ji"O���ЩIk-lp�'�I�r��@"O�p{@�Y'Ne��¡�_5ld��B"O��ssIM,P�H�dO�6Mft|�""O`�b�N�
*2.)���v��P�b"O4!�RG����kҬ"�jDK'"O��Ӄ͞y�Bȳ<YyL+�"Obi ����iA�ʤ�y�F"O���?e#�<�@Ǫk��|8�"Ox�yF�Կ
��g�Q��W"Ot��d�S'�ҵ1�@<UY�x�"Ot\;���	BϲT�UM�/!H�(��"OP���'�%7���P��x= ]�B"O
X�`Ęa�U�V�ר_���"OX��Θ6cu���능cfHrg"O���0`Y	�XU���H�=�`Uٵ"OKӻ]r=�BꙆ>g^�HN���y� ��0���;/��԰�F��y䆃(� zQ�2R�@��]��y���0"�L��j��C"(�B�K�>�y�(�"�YC���<@X���P�˘�y�ϋ�PAX��$f1��-�T���y��zY���G�
�"UtAJ$�
�y��O,ҙ� ��[���"h��yd�R���Y�e
Wg�9������y��`ˈ��t#�W�t�q�Ҧ�y��ðz�&d�2j�M���('�yb�A�BPؘ��J�~}�7@�*�y��'|4��D�.,qf1G�Q�y!˱q3N�V隰����n�0�y2ʑ6$̀HEĭ	sJ�c���yr��=14�թ0��5��T�ā؜�y��!l�P0� ��-b
�iD����y
�4V��Ӈ�؁.m��Y5gӆ�yR%�d
L����:��b����y���5D��e�FBH|9X�r!ײ�y���:K�� ��q'�yse�X2�y"g�f����`�Q��5��&��yBG��qm.̈ƪJ
zN�ٓfV:�y���Fx��Y%ř t�\yÉ���y�'ͪEYJ�!g$�d�Єk&Ш�y
� �՚u�ۯ_��d�׫�"�x�"Otm{&dM�*@��x���+��X��"O\EsѥC08_x��RG�:{�7"O�|b�
'dP2钂G�J�d1e"O�d�4�-a̩h N�q�P�v"O8Lx��m�RD �,���X�@"O�u�SkI\ ��,�1����"ON�� ���"�%�{��L�e"O�p3TJڢc�n�2aeD3:�<��"O�E3Ȋ'Rvj2�ڵ�~z7"O6�j�BƭeR�u��I�.��d��"O@D��E�t��E���X5?Ղ�r@"OP���5?�>����T�X���BR"O�1˂ ��x�VL��HQ�H� Q"O��2)��B��c�';�B��"O��ab�Xe<1Q[�Xp	�k9!�D�y��< 0�G8d�@ �bֆkA!��	���*Δ*>ČE�5���Z!�T1*O��X�����xh;q�op!�d��EiL�2��E�=��}���Ҩ�!��|��P`KU
��5Cw�I�!�"S��ѷ+�=\��p��X�!�D�{������v`��t�+G!��B0�t1�*�!	1��Z���T,!�O�!3<B�i�6$�,\���'!�$P|ڜ� F�.��Չ��I/�!�d��R��pC��7�&��&�n�!��ʪѬ8! \2Glm�Ah���!�L5%��t0���dd<C�G��7!�9G�<P8�y+m����̗�(#!�䒒l�V۶�bʎl1�H�;;!�D��:�
a����N�T�8�+J)l8!�d�$���t̎F�����F"p)!��\�8�� �X
�|J�ʙ%6�!��Z�ȒZ�"����j!�!�$ۅ*8� ��B��P�VI���!��7H�Q��W�'n���S�8�!��5,q� Ӯ�	;YbŹ^�k!�O-�F� J�,p����eJ�n[!�$H3i9��X�A8|��p) CJ5*N!��n"�M
�l?yb����aM--^!����!I���sC�D3QK�D!�D$�&���Vg6`�jD�-7!�D�)���ѯ^0?��+��Ճ\�!�O�!���铌� ]%jP��-�=�!��U�GHބ���.$$H���A,0�!�$ٛ3Jx���W&�=Tc�I�!�+DD�1gk��	C�Z!���8�0��)T�~����ĎK^!�МP��ab�$HK�$A���dI!��_���9sF];1���(��D�r)!򄘪 >.�GU�d��yHd�Q 8)!�D�X�BMA�E�2=a��Ɇ��N!��U����Rn�� �")�o��!�(	�� �A�D�Hn�J����V�!��� #
�<"��>6��a[�0�!� R��C��"`��!��:��"P��s��a�1̍�R!�d�jx�Q�����n\�VK�5o4!�䗺�"e�U�9��vJ�y1!��R��F��@�
ejUpz!��+��  -V�[���z@	�di!�"�x��Z�t��8*
C&	O!�$�'7�
����2)�Y%)J0!�� D�Bp� �T�����*wr��b"OH-0F�؈d�ġ�"��7Bs�p �"OZp�� ä:&Z5K���qu"Ov1�M�/.t�xi��'��e�"O�qa��؆i��<"D�MЖ�8�"OtYH %��J�hDHv�N�XD"O��1�&V�PF>��lU1���"Oriɇ,�$d�X*암5+B��"O��AE��6o�E����-|�(�P"O�*%eY%`ՔAJU��9����"O�袦'\Ϭ���\7��a�V����I��j�@0���T6�#� C�MB�B�I%ut�:E��$c�@١&"��
J�B�I�P9hE�ԯV$�3C^�"E�B�I^���c�_$t8m��@'	�vB��>��4h��sa��F�
�I'D��� ߩ[�A��Ɔ�)���I#D��Y��4<�a�d�Y�)���qg� ړ�0|B�J�����+�~��+ �_e�<��o[�2������gIB!{�(�^�<��ĥVi>1����;kи��Oo!�$�g�0T���OF�R�B
�B�!�DK���2���*��r��Vd)!�d�Q��<�P�T-_�^(YQ�S�!!�D���i�2��Wɬ���΁7|�'�a|�N�%i�Q1�cZ:ah<�-���y��
S)F�`���^�v��! T�y��
w���t�^��ei!k�8�y��ې|�H�a�+�Q�:E�O�y�a��Kn(QhU�I�NT^! [>�yJ8@���c�K6NzH5k����ybH��`*���H�6f]���%�y��K(u�Z�;&��A<�EX��R8��?��A��o�=F����ֆ��z&�2	�'����h��|�.�i��"y����'������,-���b�b�%^ ���'MhՋ���ktP���Ì�G��Z�'Tlk���y��P�SB0z���P�'�#��

2�H���ځ)� �	���1O�y�뜟A�&L��f��4*�����'e���ix�I�\Y���8v!�$�2�z��䆜�w��$�S�΄D�!�D��m�4�y��X.p�Z\!4�ˁEA!�Q4'Y�Ԡf�<[�XD#t�Q:5!�ݮ���Kq.S�?�bѠEQ"O�)Ѡ�,¾8Z��.���9�"O�4����&4J4���	q��'C¥U$#��@�J��s	�H�&��Op�q����9��oG;rQ,K�"O�9��IԖ���A����37"O�U��2O�zD'�&,֬8e"O����H� x�Ĕ���$~��e*b"O��v�ְT�UA�4�<�F[��D{��iG�cg�h�Щݘp"���G܏�.�� �� 1�L-U�,T�G�

3�e*$�4D�zQNG"�:��֨
�>��q�3D���#AB�:_~��$�C1^a�w�0D�t���9j�3慜 u�J�˶�.D�02c&��Gi<PN\�V(����-D�H`a����%@]on��Ök�O��=E�4���+�P|�Fc���Ҍ�3$ !���	r,��e����D(N� ~!��P�0�-��-KSo�S%-L6!��"g�p�H�I�8�� JZ�a
�`��S�? 4�;��"b���C�NÜ`�"OĈ����$2��;�m��Ş�c"OΔ0�Eȼ2�(���.��tՐq�"Ohh��I�a�
E��Љ]��%�D�'d�Ξr������	�H(T�C��P�aV�If���q�ɻ�4Ä4���e@&D� Q�[/0�|ٺ��R=\T]C**D��z	�9	&ayD'�H�`$D���	�:�b�=6�p�"7D��a�02�\=��b��@�z�?D�� �L�pW�t�
�<�6X:�&=�&��|R�O<��Q,w��$i�)�C�"OD���]�8>�S�Y&<�Kf"O���3V0�5G�{�ީ
�"O<A��P�V�܁���5��8"O�m#Bg۠]��uR��ɔ%>�"O�ċ�#Q1x��\X�n�p��J��'���K<b��0;so�DҞ�[���0��O���1�g?1T#Ys�T�d�8��A���i�<1�$V)d�'k��ڜ�fM@q�<�2�a��@�))������i�<�)�.��B%	&;��� �L�<!qi֮z�PU{�LB#lkp�|�<A�整*Ғq��չR<|��F�c�<9@dہ.��l���\�R��\��p=QWl	l�8 �Ud��_� �;Gf�<�	��|u��������TkL�2Y���ȓe�hђ��U[���6B$=��'�0d)���h�H�&'�C�:L��\��l�r�Z{>����{�9��m'l �@��*K���ѫ�G�XM���f~�U9z|Ey1+Hn�Ԡ#hM����=13�.dl��Ѷ��.T%�FH>�yR��E�t���U�I(�h��%�yrޅ4L��4c	)X@=j�(	��yb�F>:J�O�=�XM@Ua�(�y@�!����e��/$%e%��y�-+� L0gZ'S�� �*֠��>A�O�A��њ7	�}� D�P�����[����ɗEDB�q�g�]�� 3Fǐ�i�B�	+J )A�KΈ# ��#�Y��`B�	2
��mi"%����8C���NB��'��7K<�$��b�-'�C䉼A\�mo�\s�����F��C�bV�"UL V��`��&R�B�	j�,�EI�'��;P���r��B�	}��$�ĿI&�1Р
�!^�pC䉾^��9w�QpL�G�.QTC�ɑW�`a1b���V�~hW��5,C�	;h�So*z�`������FaNB��,	{�$�#��?B�H�OX�:9BB��!�~lhpG���6d�5ZcHC�	p��[c铹��I��%�j/@C�� t� �2��>A�a�b �6p�C�	�b�0U2Ea��Aw���7+�3רC�I�R`X���*��l!��xx�C�	�!�w͚�[�����7�C�ɍ�� +C;n��X���� ]C�ɰz+F�
��V�j�Tt���40�B�I�z��m3Ê�"~�4a#���ml�B�I�B���ȢBi�(I��Vet�B䉢=3�p�ш]++�9��h��fB�I�nŊ鐵�x�9�"��v�PB�	U���ƛh��}��O�FB�)� �U�1��&a�P�k�k
t���9@"O@cd/NW��H�)�+M�*����'�ў"~��M��b�I��Ae�٥�G/��x�.l����!{w���0D��!�d$0<���7 i�׃�?�!��?�P;v�ǹ;L��ԃ-K�!�$�03�$`w�S*슐�`#�=�!�BMP�P��ú��`r 㜻3[!�DE�S�<�r���	;��(�bR~:�'�ў�>-@�+ջ7d@T���Ĭ:,8`��&�O��$��Z���$K�F�	Ï��%�:��0?1�#ЯJ�00y�G��"4z�Y�<i���N�u�M:P��%%�j�<A��I��
�' �F�Hd��~�<!�G�/%���2d�L�huxF��q�<�Pn�)QV\�Ae r԰�Sb�p�<��La�kG���&��`sV��dx���'
�=�	[u����m[�^���
�'�!���~����5@�Xɺ
�'{�Y"dĎ&J�~�²�F�%)�0��')2�1W��8�t��q���\B���'�1�o�I��I[���	z��E(O��=E�-جE���
Ƞ;^�S�C(��'��ONb>� �[e���u�T�d��ua-D�HS�H �VT���3<�9u˪<�
�O�.���@�f�jŘ��H$6�r���b|�*Uo��1~\ܱ��uH�ȓa�H�®�?>�Q'H��+$���M`�� �OW�vf&$h���9����ȓ#��� T/*z�hSv�+t�^d�'�ў�|�CKƒ�Z�:2���9~�ͻ`(�X�<qW�'9f�Ċ&���h�-�F��y�<	�n	v�4D1��2��L�K�y�<�E�ɰf���Ձ�L��,k3��k�<1�֏� �����[���`�q�<�#�W�+������4�1��H���䓀���kl_�zec�eޫdN*l0��'�!�Ą�|��@3�"YMj89Ԯ��!�D6i��l �*M�f�`��~�!�Ĉ�^� 0�f�4c��\�E�;:(!�P?��P2��IU�A5!�$غ2����W>-�L�I�F��{!���,#z��P�#$T��k�LC�`r!��ޙV��J0�Y3_��c�%:���)�'@n�Y��(�~��6k���Ax�'������t:��4e�z��d��'�<c��Q<B#���d$Ol��P�'J������%���.ڪ^�L���'���Ƞ�G�3�za�s�'W����'_���U͂
��lJ�.�2P����'�PYya�=*2@���ȎS����D"O��9V#Mf#v�:�	��:�&́�"O2E��(��1�.V�Ja&�@�"Ol-�5��(OVxb���C (�"O
��'F��y�nG�F(�c"O��è����sΞ7z�V͈D"O>���ېnb<hF'��-���#�"O���D[xZ�"u��?�d]�"OVp˲i�t�9y%B�R��0�$"O<؃��#�neb�#��+9n�sw"O�}��i�-�P�x���'3���"O�h*TC@9�UA�Q?}T��	�'Gfd0f�ܑ�I�UB:.�i�'fD���Mԋ�)8�@ݔ*HdZ��� T�H&�o���2� dsr"O�u��+͵.����^�^ p�W"O�9zaH&mz��ȁ"[ʔ�5"O����)�� [�	*S~�j4"O�����7��`IS�ʍ8; <��"O����lAM�f}�&+)�dr5"O@-Y#ā,���	ȩ���"O���I�8E-�	�Ch\�R�	x�"O���,?q��R�g�':��i�P"O&�23c�?n1"���d0N<<�"O$l�1+Ҙ[v�M���sB����"O�c�A/�b9 ��6=Ҍ��7"O@�[U,���-�G,j�6-��"O���v���(���j���;�X�4"O:�y�!�� �rD��搊9�<��"O��@M �.ܢg%��x�h�:a"O����J\2\��kC�;(��d�"Oz@{I;|�=��>w�<[�"O�\�da�,@*�˔�ɍC�CR"O�44��.1.�2l��DI]qw"Oڼ�cִ �!�5O1_�d|�T"On����Nab����������w"O��HGٱ]P9��ʍ>��	�w"OXxbađ�l�*ܘ���a�}[�"O��[� k��Y�D���a�dA"O�;��	�\�j�'�?�~���"OF�ѓ)W."5��L`�\��"O��V��E��	j���^�� C�"O�V.0�0�4�V�B㋕l�
ņ��
�{���F}�a�[�Y���ȓql(��#)�8�BՃ�~}�ąȓ5��8�C�	�P=��%��;P`��p������2�~���.R�wSRU�ȓ`7Zm�Vkۍx�l�kV]J�ԆȓX��hqPn�%�VQ��D .w���ȓl�R��gA��'xݚ��Y |����ȓ<.*}{���,�v��	޳
g���ȓF,�B ѳF�L�t�Kc�j���t�6���H&>m�4���Ń=��0�������2�j���`�>[�0�ȓ 4�PC �}~@ț7��~�l-��/�f��DAΝC|P��s �(y;�	��b��1I �M���+�޻;��ȓe m����0P�,�ӤU9�z�ȓ~h�%ء�3; �c��-�XD��Z�$Z ܆N� ���$d�d��Ą�����$b�\�r.Ԗ����ȓ4d�r���%
X�Pp��K��1�ȓ!��AZb�L�c4�E�d/�
L5���ȓ��l)`��y�<�:pcW��(͇�1�\ј�Aژ]�Ɂ��TZA�%�ȓj�;E�(�d�	�D\.wڕ��Zh��hqm��TQ8���ee�e%�B�<�%!�"1|(�gkZ�Rdd�X�"�e�<iV@��6YF�A��A�6<r�)��Wb�<�u.ӗd��!(Gm�!X�3��	b�<1�ϙ~<��I�9,�*�ti�[�<a5Kq�4ᱪ�N���AU�<�5fA�4�ԔZϙ����J�Q�<��ᎏ����c��x�`�r��X�<���P�fdj`g�(&�ye�l�<�$d�c�:q��"C={������i�<�d�ҹ`��9K��#�N�d�<�� ��I�<�`	F�+v*�C�E_�<� &��`n��8v����:�"OZ���A�]�¸���9K���F"O��[P+*�0"�\^��!�"O�]I&%BMMt)�cNG���"O����NHł����)�ʈ(�"O��sG��D�b���eu���"O8!&��;��D�d!�2Z\TA3"O�\wJ�YPPy3�W�-I.��t"O�$�"�	L�$��<C2�!�"O��#2�?'Bi�e� �=���	�"O4x��Θ7g�L�-M�}ܥ	�"Op�aR��-g��8�6�F-u�"O���"���0�7��=`z�f"O<�+ԯ!��P��߈`D��"Od�	u��<}c��R�sG �Yp"O�����>tr�Qj�����k�"O���.�:! ԋ���nph� B"O�ypb��⡩�⍯��@I`"O�4��p���Ñ�|�fe��"O8mYu܇);�Mx 4�Ld�"O�Ԁ��͔|H ʎx�^��"O|Hz�F���ɳ񋒱w�Ȉ�"O |K����@��h&�X�i|�E�"On� ҡ�/aPd��I#
��Y��"O�A�p�G� �� �Ŀ+�T��"O�p b�d�ޠ� �T�6m��%"O�t�AHX�e��|�.O�l����"O�|�ˀ�#��C��ORhDQ�"O��#�ܩR<9�̜��T5x�"O��'	�w2Б9�mF�o�@Y�"O��q���=��4��
��
&"O4�B��׋I��r�@�ײ� �"O���g���tI���q͔�kA"O�l���/g�5(�$C�O"�sS"O��y��@���ٺ��O�~* h�"O��0ܶ�"��P���t��͚"Of;��" ,BE�̔6Jw$ɴ"O���p?�$�ϺGc2m�w"O,���_><���JFP?+%"O"Kt"\�=�����Bd&X��S"O2h��Նr	Tr@�̨LF�`r�"O L��!.M�0��4���?!���"O.Ԣ�[�l�di�î)
XS�"O�a�@ #yE��V[�j�]�C"O��ԠR"3����쒵(�vA��"O�ف���>Q<֠St�h�P<8�"O���ah[�Q8�-[C�6K���"O"��fm�%S!Z�@
��2��� "O(�%B�_lT��L�NHR�"O�m���)М���/�W8�r�"O��j��D�V�Ԩ����9$�22"O���25�Z-�T��hXݪ�"ON���G90Kr\�B�:i_,|C�"OX@� �3b���3�-BWfhB�"Oj	��Ő�Z�L��숞o�pH�"O�qӃ$ԑ9u2	pD��7�ndp�"OL�p�� ���9��~��0)�"O"iu�ߡ*��`�eO}�� s�"O��Q���/!���q�2h��]Y�"O@���T1<j¥��CG����[s"O�0ì޹mxܽh#l�;r>Բ�"OԽ2�]'_pVhi
�8Xҥq�"O> бH�>���#��wB�i�"O֙� ���
��XR��Z.`.X��1"O� ��+�톪#;F��O�/�B�s"OJu��G�;u?�Ī�M*4�ް��"O,��v���1�v1˲̅�&Ĩ�'"O��!Ƨ�;�� �0xd�a�:D�,�g��^�J�a��$4CN�Ru=D� ᣉ�|��۶	U�?vz�˧;D�X�!O	dT�0<�}��9D��`gO	3w<���DLu��9D��(A��2!Q�-�U��wg�X�`4D��D�ۛ ��j����l��l�p�&D��iE�/5���:"�]��h��eG'D���Qm�XgVp��#H�����'D���`��t-�i�'�x�$5�c�'D�Pvn��j}�����1D� �@��$D���G im�����/"���Vj=D���ƀ��=$���U�_��4I�<D����7�����Ϣ4�Թs�j<D�<�i��i*�	N�����w�;D�ę$D'� ��"#�<�n�B�;D�����A�-� @!g��#�F��W&;D��"�$I:kR�3���$F��s2�8D��KF��+bZ��mGY
pg�7D�h �]�{����D����c l�<I�Q�:8�!@oՁ['⨡�	�i�<ar#߱|���H���R[��ۦB�_�<qr�M{W��E��<j+0Lc�ƞC�<11�MXN��v�]�J�8�H~�<4H��6���[j�c���h4H{�<�f�ʄO�����;��谦�~�<�r�V7}�~��扌��Y BM�P�< �"6t-iD+��/�~	`���L�<YPʟ��T��-�$P	 ����S�<�gL��;����ٝ#бs��OK�<ApnH4"�B5�����")WK�<�E��>}`6�Qjܘ@ Zm���D�<9�G�p�i{���m�"$BG%D�<q�/H<p�,LdD����������8��2�(q���ecX�ȓc�L9���=M�`HcEg��^���=�h{Ҍ��7�1�ӆ2H�q�ȓ%<j�c�$,~��n /���ȓ~�Ƭ�a����:��Cz���}�t�ru�(]� �J2�ќi �"�4�{��	������^r��ȓn�:���C^p�)�IUlN@i�ȓ`�y�G��.D��H�ٍc�̰�ȓ1D��(�f��D�p�	
:y��S���R��֕QV1(�[�~���2Q���U�XFȄ)׹��B��?D�t0gj�9��e��;8lޜp>D����f��WC 
T�:��Љ�
?D����R�5���e�N��D� >D�ġ節<z��cށFN
��<D����o�Jc&H)mx�E�C9D��@��RU8�J��=TL��I�"D���Fa�0Ҧ���%ސ��5k?D��ʰ�Ɗ9Fl, b��l=���;D�pJ�� 1B)"�+P���3��2�/D���aͨCvE���N&o��t8	-D�@i�_!}���cdL�r���J�B D� :�#J$��|)� 	6p�j�2/>D��U���_JH�� d�2x��=D�h�&�9U������E�w��4.:D�di�E\:l�q	��C�4�=0�)7D�� Ȉ�!"�������,&��L��"O��#aF׽l P�w!�B��K4"O.�YĎ��9E��q!�?��;`"O�� �~"H�r/15��X�3"O a�)�l~[w�ώ9�6�pu"O	�5ʞIn��i�L�1��)��"O�����T�Y�Θ������"O|���F	 HK�Q�M��x��)2�"O�dےI�(��܋�gƶ�d� "O�iԀ�6S�b=@��	0-�Th�"O���鉢R�\J�D>|�a	�"OD��&l�+:�)BE�0r䑱�"O�� F8x����ȧ
��h�"O�8�w��4�D9z��G#/=�p�"O�ZU��?/���R��@�m2��JV"O�98�Y� �\U��&BL!���"Or<1��ڃd'f)b��ܺg��I2"OpL@�H&?�HL���;��eڣ"OXI��)Q�F�L�0��.m�F��5"Or�I3�ڎNLfu`�+Ԗ3�`�@"O�T�,;�0��%س&<P��"O,5�V�Ϩ���+œid�H�"O�(z��N6kn�D�G��
���'"OD�R�ھ�蔒tB����sB"Op��ƦK|�D3�'��2"Oh��S#�0����I�'a~AZ�"O���V���LWL)@`JG>��� "O�I0�A˂O�2ղ�kC,�Ad"OPy�i� � i"��AxBؠ�"O�a������쪃�`Xr� "O�Q�"�ĆYvQ�"�˘rI��Q"O�\�e>n��v`�![v��"O�%yd���}�(y:3���mS���"O:����Qx�(�"��A8�0t"O�}�e�Y&%� h���g�h��"O�Th����H:��Ȥ��/�أ�"O҉���(5�r���[�\|n�
�"O�0«R
q���3���PvP��"O}ہH��L�.��V<�.-�"O���CO�H�d*������� "O��Z���=d�.49�E�A��"O�|��G��	�A��U�M#"Q�p"O>�3B�C=5,��@rCМd�D-p"O�ܱ�o׆I�DPF#I�P4p"Oj�s�X�KU�b#F��d��%"O�EC僑�+(Y)��3���"O�Y���+ׄ>���� ,�V`!�ֳ
X�ȲƏ[+d���
�E�(wn!�&��Ű'I' fBG.ĚR[!�N|#����,��Q�������<�!��m�FXQ�5)����er|!�$;}V*���l��Q/�/c!�$D���)� Á;3Ѩ�ct-�J!�$�w�P��	rb�yQD��d*!�$Y>=�$��pJ��iY -	�bF"]�!�d#S���E��,Xs@1b�'N�.�!�>[N��Ы�]�(�Ɵ.A�!��҇j��(:�ʣ:$j(���Bb�!�$_+�VY*�̆�BC�@�1�]��!��ڥ��`��Ast�ȗ_αz�'rQ�Dɶ;�HP�
��T��'C,�ϗ&�J�S��B�'�EH�"�2Lp�A�Q�<a@�'�4\��o��y�R�j�	�Q��)��� ���u`�]�"��ф<�0Li"O d󇈑+m3, Pg#N�ph�#�"O�y�v
�1��á��3`F ��"Op�����b��T�ƌ7�ҙ	�"O��s�KV�������OTA"Ot 3�I�<��U���ظ_mR�yp"O��c� �8��=�V#�3��h�"O<<�TK�h�����@g@���"Oz���I�i;��qՖj1�P��"OiR"��3.eh��,�K$f�Sb"Olu�S����������h�"O~3���$�� 4ᒀol�Di&"Oj�;Ҩ�$X*�D���&_���"OPl��'Ρyo�d1���	c��b"O4)C%�oH�����`�"O�p�S�n��l�Q�Ý |H]�Q"O( �u���B���A�I�{l��k7"O�@�O "'�0qUb�c���"O��ㆵ8�8
�M�)NzQ3�"OR䂁�]�v�$Ӡm�	f�BY�w"O>l��h�3g��4L�	[��H�W"OdU�2�
'���p3�?T�`4� "Ob�6�7��H9P@�0��1&"O����ŉ�piB	Cျ�$�W"O����NʓD��	�W�g�P���"O�u� ^ B�J��0����5�"O�IWΏ�����u�Qby���"O*����G�ؼS�@��R�ܙq"O�ih���� !Ι��EX2>])A"OL��K8	�zԘ���|��A�"O&ɱ���=O� �7��7�H4��'���rW"�4dy^��`a֒X�����'� L�0���H����X�6���'HfXk@G$8�`p�ζWᶰ*�'j��(�	j�a�X_{�=�'��C�MG�%��| �,7W�R$��'�*a���
wB��ʈ [K�� �'�
Tr�G�R��� ЫLw\�*�'f�q�CS�~�
����OV�pl��'
.�@��J�4�x1��5T�:Ř�'`:}!�(C)0c�A�:#��-	�'�N�����UOąy��%�� �	�'�$���BO���Q���q�Lё�'�n���;1<"�y�(B�b�ua�':�Dp5	-8n)(��b��h�
�'�� �c�h�̋��.X�&!��'8�H��W�*=��;ԣW$��@��'��]���P>�h�`ۢߤ���'^���n�T�8d���R$�by��'PP�ჩ��V|��i���|��'����͊?::��VbO0	��'�6�C�L�~��d:���(X_��Y�'M��@LC�K.�[��Q��U�
�'ΦU�P�I�z�� �b��BE��S�'��c���:�����$F�栳�'i���ef[�kʔS��1>S>�S�'�FL�r�Q#��@A�6�`L!�'p�0q$�GiZ�}��) �%z@ls�'d�උ�"����k-��)
�'��ȣ�)��Wh���7�����'�d��Hs�@�q#���`E���'P>���<p� 3Sl�)����'�4H)!];~t��`�W4(Z� �'[��H3$N�,��JvG��&������ \�J���1�Hcs��F2
H{P"O$�s��ڳ*6�ՁU�=8|��"O�ĉ��z�<�ö%́2_zl�"O���C�( ˰���.��9� ��"OJ���I
� ��v.	� ���c�"O`��g#M�?�؀{�̪�0x!c"Op�w)�w7����jS�Kf\��W"O���I�:E@��	�OČ b"O�I�'|���0�V�R�Nk�"OFa8F� 'xXX}ȢAV��px�"O$Y����9
8x���{��93f"O
�)�ERr�y#V ��*�Y�"O�����r�x�kDj,�L"O� ۶=�()��ޣu�
-K�"O�<2%�ڵ3/���G�<MZ���"OT��a��n]��ǑF�J�"O�p��EϮT`v�9gV8]���#"OH� � */�f͡S@M	�Z�`"O����&��%�� �u��B�2��V"O�,YTMK\���Ţ�"h�p�b"OHL:��X\��PdA.��0�T"O¹¤ 
*�|a���#6}�"5"O^�Аi.q��q�?+̦T��"O�E��DѵHsv��N��D@��"O�Ғ&
%1T�8� �=J���Y�"O$$�3�IEq�ՑÎµc��M�"Oz� ��Ie0��� n��~>���"O
�����	��%��"|4���XX�<Aa�	�.�A�!	Ok���K!`�y�<!l�`����$�A�Lr� �`�t�<�d�C����)-J�0 P�hPU�<���K� �9��?
����ck�Q�<	��.tͰu�B�R�3�"q�q�P�<�P^ϐ�s���:X��G�L�<	p/�4n�� �k��YYd�r�O�<I$�½&cpt?�*���K�<Y��H9�*�5�N�=�Jł���a�<I�C�ZH�`0�J�҃G�g�<�Vd�0{�R(�W�ų3��X�%#�\�<!�Dʹ7ze��L�	�%����T�<��¹,ȁ�UI�U1���3�P�<0��c_��[3l�	
ƅ�&��E�<!AnR�h��9%&����� 
L�<A�h�	5��Z�ā#,Z渱jBo�<��E�Y��@�%�88��qG�i�<᧌ۀI$B�3��5K����PTc�<�$�&v4�	��%L�?Z�9� k�<A�L�#P۱�үE{��d�<	3g�=�P�'�0"R H�N=T���OV�&C8Q�a�հ����+D�t�B��D�����ҲJ��;f�(D�HK��X�;�-;�E�?r�Ȣ�%D�X+��{���/��^44t�'K9D��Eʛ�Q@R95$̚uF�d;�8D��9@bؗ6�
��a\)y.���f�2D�HЗ��S�8���ƈ:�x��,/D�Xjn�Z�����F�&c��kf�,D�R@��F��I�'�Uo���� ,D�p�qb��3��=�h�'3	p,8��>D��0()�r0���]�e0�vn'D��W.��`��p�0P#���f%:D��$D������2;�� �5D� A�X�0����R����I���4D������N�w���_^l��=D�� (	�$a��P�i]�TH��"Oxk�l:Y�t$��[�r8C�"O�����	J������E1�"OV4y`b�@�h��F
�p�r�"O����kD�PC���-h���a"O��b��� d}6�U�[��,rT"O�	1s
�)9����d��%��k0"OX�1f�/G��YW�٨nl��p�"O�y�O���b�Y�0=����"O0]�&�ѐu,��rg��I6V��"O,�H�E/�*5p���;GN)PV"O2��`���q>8yXg��,p,��C�"O���H�"�jqj�O�H�(�$"O���e�<[^�t�M�i��I""O�iS��)�Q�Ǚ|p��"O4�k�
'!bx���.^2���"O��Z��^7�����W&XF���"Ol�&/������҆	�j���"On<��Ig��D�B$����6$�x�<�5�H�c�ٱ�eB5�((ICʖo�<Y��тq�.$�p�W4Yu�	���s�<a�(W<bR6��&�聠5�Al�<q�  �z�v����tx@b��k�<����:mRd�*D�Z�X� ���~�<1ti@�f(��{}�� L�w�<�C�� M��EY�m־R�l1{`��v�<��)�5R<p���נK��t˲ _g�<��L
{~������H��R'a�<ɇ��.e+$��Bl��a�b��B�U�<�* @����⯗#�r��$ �G�<p�ʄc>�u�2H�6C�����A�<�&�F(���Zq�ؑoh���m�t�<����>�1��k�|1�lyr��s�<�4�@
���#�C� \|�k�W�<�2'N�g����m��q8�Zr�Fk�<���ҡ�4䙁A}���	�e�<qq���s}ʈ�4D�l�0� �GM�<Q3'�Tp<0�]�M���yG��E�<9�ƕ�6Ҟ�k�2�F4�T��V�<���T]��q1�gQ�y���2�AG�<	���o��z c_"�)a3���<a�ł�&�\asc��V�AH&j]a�<��gA,О9ʒ�I!G����e_�<�s冩Iȴ���W�K��㓣q�<�W�Ŝ��@X�����zU�G�<y�N�^�|�`��^<K�X&�h�<��됣u?ƥ��L�4n�B�Ko�<qӋ��\Af��N)���" �i�<��(A�)2��e�[�n�r�![b�<a�'�@�=���P%?����f�v�<���.tS���w��!&�Ft�V�v�<yT��	1-�����\{�|Ӱ �r�<q#���H�� pA��]X���Cl�<Q�����m�&f�8]����Эf�<ɱ�\�yvl9i1-��ݸFE�{�<9@>796�b�eG.T����C�P�<�0��mm�؋R`Q�PJ$2s�KV�<���݉+�t}��D�'�:@Z�h�N�<��Q�*[BE�%�3	j@����e�<�����!�G;�v98��G�<�!�ӆJ�T-6��66+�Eà`�Z�<P���`�,�P��I�j��Ms�-R�<�t��
��2�&űc-�9�sOH�<Ae��l�4�g�-~��a�(EB�<� ��6
�D�@�C5j�\AbQ"O�[��_�m��A���!��]��"O(ŀ��I�v�f��QBN<�J̚"O��x0�C�fDN��gˇZ��P�G"OHMK&GG�N���S(>	�+R"O�J2!ڈ+���YǏ��i4SQ"O�
R��9%|`��P�S�����f"ONLc��df]I�fޙ>���"O�
�YQ��1f�n&dL26"Ol�%�S�DMI�e^�ڼ��"O�hR�'�Z�I 䡜�r(�ԩ1"O���$�;6�@!CA�74\�A6"O���CƜ4A� S�� {Y����"O�ɫC^3N��h���&?���"O�R$��t��i@ �(,H����"Oz���h�C��T `�ϥ�L���"ON���H�`�'�H�i�ء�"O����	W�Q2P����.[P��B"Oܰ׮��m�);/ �=b�"O,0`��I/qtxYb(�_'�H�0"O��*D	�)V*ԀA�A���9V"O�5�4$J)�t���#��)i^�h�"O$9##%���hѢ$w]��x"O���fG����e����&jF>I��'Y���}x0���of`I�	�'w��A� �("�0�E
�f��Z	�'�|��a�(�<��'i�1�� �ȓ�nQ:���<����cf�9uB�l�ȓG_~����Ҷ(�傰f�7�8��|��$���Y` ��elZ�i�b��ȓ
nN��l�"��B�`� g���ȓI�
�e
<d)��ۣ���G�n���H�����
���"C�>���ȓG����ͣD���P�i�
����ȓ0� �r�(>v,	�*U�̕��q�f�V&@���A�"7#6Ї�Py04�@Gڝa�)�f�[	pGbхȓ.�l`�'K̗G����≞9"�,�ȓ>U"���<RH�d��f�:����m�SNV`4~�h�/�{ �t���,�����vRD`pWlFݤхȓ0��a��BۘL(��C&ɡT��D�ȓo"����I�6�B�K�O@nt^��V,��� �/{�. ��'D\��Ʌ���X�B�ֵ��5��b\�`*P��sd�X��ʕ#!��12�<J$@��݊Q��L�1��ȹ�Ҹ<�8���N:����ɨ+p��E��:GV݇�g�����(�`����8T�����$��� Z�]^]�UC64���ȓ=��𫐂7T#\u)RK�2Z:��ȓ\D���$
w8�h��6O~\D�ȓ�:����v(p��b�4+�"���N���+�5a�p��C�3!�hU�ȓH��ЃA�L�*�.�0�산V�$�ȓ$�96�?e�d��N�CX�1�ȓ-疘����G�L ��W�'�\��_����5�Ewn����+G��伅ȓ�JXf���p�T�Ä��Y�`d�ȓ2��4���b=�FD"DɄȓW�FI�Ł1GC�����e��`��Ez�d��'��kgf�˵��:H 4��$�=���ʟo�洐�eї9��Ň�r���Lߝwb��Q��.�(���S�? �i��*��R�J����-��Qy�"O�lɧ,���D�}����"O��P���2lJ����2����"O�yR&k�>?�{�!�-H���W��/LOʥiAdϒA��Q�@%&{�@��"O�l�Ӏ�9h��R�0(�,)4�$0VCՌ)�M�]��)!��>����ڿ��'�^ QHF8v2La��c���4(��'@б�R�}/�ɹra�*{�H�cM<I�O�����.@��HB�A�AE�M�")H's�!�dT���D�iM:Ҁ��!-�F)��8�DIzp�O�Zd�Rr͍�k����O�r��uPKL�Yfp,a���B?�Ls�'�0TX�aY�~^�4� '@�f;��ҍ��)�4�VW6�%�&��zA&� Ƨ�=�y"知@�4y�*@l���ؕ����hO&���+Vfla���"��h��޳_�!�[-^H�DE�;�Z����\7n�!�D��8���oߩVyN�����J�ȓ:3\} ��;u�t�Y"/�+H5�ȓ+B8�#���_��� �$h,Լ��R�D�*���~��]�T��}�T��L�/EUT��W�܀��(��hO?KDb��v=s�
k��= �o/D�h�IV�7�h�(E�U��Q��g.D���T�>o ��+��cSc94�軣/��s���b��J��ȕx�<i�-.�}�2l^c���1GVj��q���O��ր�5b`Na�%X�HE��'el0 �cA�z&�+��7tU6u�4/��'��I}�'�����	�1a��+�`pa��'�����M�yK���I�ʥ)��.D�HЉ���h:3�O�_$�� �9�ɚ�HO�O�z ��[�ʮ��6n�/����
�'� i��A�n�q0���.!�M0���<A���3T��1�j�7c�I�#փ5�!�ԍf��T̑�y��t�у�-y�!򄊷@��<(�ǒ91����<,!�OJ((��ICI��ek=n	��Bx��C>��8�2��#;��Ja D���G��v��(�p�i�Di� ?D��aצ��)^L��@�Ը_>x*�8D�\C�T��M��+�3j��TK  6D��
�)C.)XL4��ӉR6�@�uG5D���'� ϲ�H`iPW^�� �3D�ٕ)�=m��iA��(O�����ǯ<
�fS�Q��,n��$H�Tu��!���D~E��;�C���:ul��Вe]'�y��÷%t�İ@Qn(2t�WV�y�J�A������.4�@͹!Y��y�g�[6��R$@I��&�A�yR�)��O?�o*��ea��Y�Z��=w�I�<�C͝�w����]�A�>�0QMB���d&�S�g�w���U{8����
	|�&��AOP�u�0�keB\.(� p':?�����'��O ��m�^̔D��J
,4����|b�|��kV�)����<�N�sj7b�˓�0?���5 �v푲�� <Q,���f�'ޢ<1�Q>��劖����1.�O=���1D���`mG �2��@늾|S�=UbN� ��O ���i����я*m"l#�D�a{��d��r����N5]�R�J����~�!�Z�#fA�A�V�F �+��\�!��
\�M�OٞJ��%�l��5�!�� 8x�d�08�����m�[���#��'Zў|4ę!|n8F"��s>)�a�,D����N��i��`	�'�
Rxq�e7ʓ�hO��>J�4�)@�,`��/�J��d!?�qfG e��Y"��R=�ֱ��ڦ�	�'�qO?7�V�2�Z���0l¢����2OўȄ�S9�~x("G��L٘e�@c�?�LʓF��}��=[���@HVO��)�J��HO���	*�X�[����H��(�?u!�䞟�Z����A�k��"C샌a�!���(#^�A�s
��T��hr�kS�!�$��w�į�h��Ͱ F%P�!��
�,�Z�Nτ������$e��D{��0ɓu��\Ȉ�f�[��azg"O4���̣8�|�El]�Zf�t�iў"~n��VD|)�M��ke���bO�.�C�	�U4�S0��"^�z(X�G�%����HO�>��!�J����(�[~��j��>D�H0􁘒���&ƞo�U��O����'��h��"����k�
�`'��"��;D�$�����f�򢃃�W���ɴ�3D��ksk�h����ނq-t��2T�z�c�D�BP/�8V��L 7"Ohl�G�+��(1A@�8�DpR�"O�	2��%0����e�5 �f��"O�L��C��P ©�v��>|4�"O�a���DVf��׬��;V��kT"O�	�dlʕK�\0��lW,J=��"O�=�r�G!N�D� u,<��6"O���T�����U�"t'�EZf"O����f&v�d�J���������	G-HAr�E�
Y���@�&f���v������v�K +�ԛ�gS8q������<�S��yi�+���E/?,�Da�$��$7�O"�t�Z�'>NX����!��òi���$M�a�6�����*"x�}#�灄^�!�D��)N��ۧK(WF)� �ax��I�7����ܺ��3`�Z�h�z��p?1�&�N~!��$�d����Tml~��)§e͘h��Ȟb�8TO�J����ȓN>�BWM]�@F6�CWG߻H��9'�؇�ɉ^����矮Y��y��Nͺp����	k�I5-_<H
׬I�T4�P!Ƶr��������K�24np�5o��e ���d� g�!�d_-?v	s�[�\鎨�cdV�N!��A����5����\dj��U !񤜪$J	��O�G3��c.�X����o��9"gc::��	�k��zmЄȓ����S�4Iw��<i��,�ȓk�A�d��,Y��e1�̑85� �'�@���A��|&�d�G*�I��ړHǾ���Q//$�pK��ʺD�p�	O@�a�Z=�g;��'��{BI^'c���f��%=x����5�yB���1ж�i�/�=nİ F!�DO�~' �'.��~!�	vN�� 1qOF(�뉝+t��q�!��l`B �6P�[��C��:,-�R�N��>��"��1@X�"O�#A5W
Y����]rt��"OP4��←7�P�%��3n���"O�����]f��#�"R"PH�"O��`!��y����.gK��ha"O� ��n7\����\mAj=�"O�q���1X�亴�8)��i	�"O��'�*����� |����P"O� ������?~ƹ�q ]:�ܑ"O��RE�If�~�����;�ޥA�"O�Yj��_�DRC�	t|�aB�"O�E�"t�HC$�l�<1w"O�	�u/0(<EA��h�Y��"O�5x�"�(a�x�q"�	�J�%j�"O���Gw�Heq�hǎ%�����"O�MI��W��,	��ا	�
��"O�0�. _�L���֍S�����"O`+�e7-�^�j�!�5;lزW"Of�k1�]A�:(Xs�� b�ԁ""O�$q`ؙB�P����EU~XXW"OB�x1d4+�u;�>nKbl��"O�����	�ă�fU�.ZUj�"Oz �%�̲"lF�@�eł45���"O�Xp��On�7�O�,���+�"O.�2��*h��<�6�[�'m�i�r"OH��эT�.a��Ŏ�u�2�J7"OЁ��!N ��(��d�Z���k�"O.�`r�38��	*�_�h���"OfD��GB�-�n�3��</w�!yD"Or��B�:s �rV	88�k�"OB�@���Ǯi��Ҍo#��6"O�槝�;ܽK�F�ə�"O IBTޕ|�2��'���J �l��"O���!��E�>mkd�1���P"O2�b�O0F;0��-����D"Oz$���%Zi���QI��E�"O��[��p��(��"T��]R�"O��TL�X����0#�K�PS�"O©��BC�p�Q�B9]��d*O�t�Ƭׯ'M�H��Μ#Z�M��'�r �o)7�*	����wsڨb�'b��"%�QHrax ��\��q{	�'�"l��TBL��L� S��r	�'���y�n�6R4~��t@m$���'͂t�@C�b��]�R)�5k"��'Ī�G��7�l�3��4�����'j$�(��))kd�1�J�YN��:�'�}"r�Q�M��(rs,Ҹ*��e�
�'MB�k钍%�L9e�<8�9Y
�'��c�B�n:8��V	��a
�'�ɪ��-i(Ⅎ�*!�� R�'͈�P��"<�����L8��'	r=�Gn����i�Yc�TZ�'�,Y�`���nDJ��]�4J�'�d1;P�.���7$�
O���z�'W��H��HH䑑�._�9��T��'֬q V@Ϯ|À�!���+30�'pr�c@DL1@��ظPH�]�|P;�'��H�fΧ�⧤9X���a�'��I�5�۽�D)WkC\w��s	�'� ���P�'��|0d��d�"d��'�dU�dG�:7BѻB`Jfgn��'#B<X���%Q!��V�� �Ȃ�'�xh���5�����:6�%��'�&]P�� L�pJ�)�16�)Z�'�nܢ�Oܷt�V���5/���'�2@������p���#}(�[	�',�������(	�CE:��S�' U˦a��<�U8�b�WKVı�'���Te��YQ�NF�I����D�A#�JNI��DH�>�5�ȓhi޽�qΗ�t��A���D�\�t��S�? ��cg\�,��t��(�P���@g"Ob�h�J³^w�tJ��/`�����O`�x��'P@�(��dg�(0��)�ə	�'�j}��K$M�84!�۸1d����$L�,�>���<�S�rj���vG�aW�MzׇR�!ChB�Ɍ*X��G��xi�BJҬi�t�<>hP���P�dӧH�jeQ($�� �i۽�N���"O��BaF�M��hǧ��T�py��+}�ς����#��D\تa�C��"Df����� a��@�
������J���a��ǿ__� iuc�;e��i���":��LaQ���;�*�B�MqlF#?�'���l{�9�.���j��|yAf&�F�8�o�<v�!�DJ�CZ��IV��za�a�����2x`\�k�ɺw��S�O��x2��14EP���ɑv��m��'1 uy1��)J�%ɲ��$`�`L�6�>YҥSLʈ���}2N�:^�89 o��/XȱE�֙ܰ?1���,s�uB&`�_��1#��>S�Ĩ��ئf ���d��`��`<4�����(D�
�џ�#I�Z����|���Q1��rw��DNG�A	�Ņȓe���n�\�U�B�L�=����'���6��Y�S�O�&�A6���޵)�L2>IDe�
�'+��G���r�6����A94J����'g\����Z�ze����6r!��'i�c� �I��a�2�B�t��e��'���Ѱ@��1�¤[�$݊ț�'��M�e$�3L&�"R�]8v�:�S	�'�p�g�;Ʊ�� N�)$���']�}����J,�A1��E�s
�'��E��O�
�^��0	԰�(��	�'�~9��fQX�����l���TX�'�z1�v͝!E��0g��}�����ņ<�؅�
# �K�W��S��:3�X)EZV�l!�`
��OK��)�&	��������	�'����c\�>�2�HV�n<l=�O8�q��31x�'i���!�_�OO�q�@M�"�$a���u� �c�'i��2dF8CGL�1GXjm|�h��i�ȀW�H�b6�,��팭�O�h�QN<)�L	�'BL���yY!4L�|؟ �'��(�B ��kG�	��:�O+6V�ij'lőN��bbª~F��f�+@D�"���OR��Q7=-�LJ~�Ԁ�-� m��+�P6�H��/UD�<�V�s�d]��IƏ9�84K�B�G}K�J>f�Y��j��S"C���s�녽m92�&�)�<C�-���PD	
�<|�`��4l�ѦOFiȒ��+lи&>c�H;�0f|d��h(�s�"�O�X���sǎ@q�ƴr�ft�㡍4T�` L����?�q�X�9X|�#׃[>+����ME�'��\�Q��8\v���~�'�8�BOL%W�RM5
�7������
��*�L�υL��;`*�*b����2���=�^�)��<!��1x��̡���{Nt2p�q�<â��o�x�ꄣD(U�� ��

(1-�q���/L=B�B5X��S/�4�A�>�S�Y�( ����4���*LA*��$G?x� �')��$��n:Y����rJ�)js��A��I,��H�N�#4#޴���ԃ�;D��'���D�N�]�\��S(ӡ'1��K������@HlDyT�_��إ��̘2�π�%�L/2��[�H}�q�d�)mz$��v�`\�slK	%����N��,!ǉ$H���(��X��A��ϱu�@nڴ�H�+^8�N�	���R}��?QZ% 1b�$�8�jͫL)��Pe�D��d�5��X�qPtG��+d<�cׯ�"	˼,ٍ{��~2T�P�
3��O\<�SR�	()�&ώ*�dh�t��5!"0t�Ț�<R�l��SM��΄�%1R҃��3g�^Ec��U�2�E 8s&�ԇ4a�T��|R  �r�:O�,Z'�˅D�䕳�)WQ�9�v^�h�'�;T�Hu)&8>�ڝ�b�~��,�uw�+рU�
�\�!Ǖ"�]!e�\\���#?��p��K�+�ayb�A�@���AGD�6�������R,
t;t��uE���26�̠��JD�n���;�P?�'�]V:S�Վ,8�A��Y_m�'ĕ�1��~���R7v�
���S�X���'�2断EX$�1�,��0�f5�OvK-�)+� �h���CZ����ߌ,D�P�a�I�Ai�O}6�1*���4+D3�&4��kC�Gn�\1O@<3q삒�>�ZĦ�<�'	On��H>�!�ÆKO�!�a�_^4=�A��|yZ�0���+'%?�8��򩎳x9 x�pLҷ~�htp��F8o�UH�͚���q�>,���'�"�hs«S�I��B&
G�U�М|��B�B�E����ybW04�q; �M=j�m	@*���Px�k��2�:t*�퐿e����� W�L:��g<�5N��l�����5%rHL`Qf�<���G9n^	z "Mx�<) p�E]�<1s,��i�n�C�œ�b�V�<�5�ۗ^. ��ɊA�`!C�K�<�t��iH�3UK�PN>����W�<	Cg׻I�YAR�U%=H�����W�<�oF2-Y�ɻ0��|��؄mQ�<A�i�:Y:H�+^�*�h��V[�<yA�ݲi�b�Z5Dי}Pup�k��.3�>����'�D5��FP*���P�~ݘ	�[�j���A5�5�7���"0 G��*�
�с>��
 AU c�D]���+�"��e@0ғ�B	�ઐ0I�(Ԙ`">�陕o��|2 ď5P-<��Q�.1�!�ē�t	`u�a��N���ƵJ�<�Z�`V�C&$�t!�-olX�)�矴)���?���QH�6��0�n/D���
�5MDF$��Ȯk�h���Ȋ8�?�t�D�y6���K�*[���3�S�6M�ю��
:�Q2H �5=ڵ��ɒ@��١���[�6u[FA�6AN�����H�xj����f�dt�'!~�h���(��H�S��)��]Ȉ�$޺	N��A�3X\��B'\��ӸW�:�bdM, �0@��d7-��C�I s��-j$��F�pIB5#�('H�B�-"�-
S�(@[B=ڧ�yr &V@ D�ÁRӮ���+���y��)%�j�P�FN�} `!��?�J�J�(�Ff��ǀ�z��`���%�ўTp���r���X%�h�± 	+|O����	5��` &M�a��(C�>+�����>=`�I&�L�Gf��
�Q��P�g��O���x��V�M|��?A���.�n��R�O?�-�Qf
�g��'V(  q ���WB ���oԶ7ڂa�ȓ/�<of�hXpĒ8{�N\��!	4�p!F)� M8�ӗ�E4-Q>Yϻ<{�M�&���a0�#e�I��A�ȓ&���L)y��1���$�@�"�K <�ƌҷK�1&=B��L��?���Ʉ61K�+K�h �KTp���S��8:'"���T��姜'G����`F�>�  �g�.��P��!�/SS����AsҀ�B�'�2�"f�b�����0I��Qj��`ӊ�0X�lh��)��qSR�",v�資�R�u�w�"M�D`� ;�,|"R�!M��u�	�'�ԄC2�U7�����^7������&�X���ti�c	��քKNՀ4����1'�~�]QΤ�4h�#r�4\(�iU�D�Ṗ�I��F�$D=S�V��'��qBf������9#0PX`"a�%`�AP1. H�p���hO���h��I�4XXU`Z�A�j,����fN-P���	��@ C6��q%`�G�H���_K�P����ָ>���GD�>B����7������Κk� �`v���Zc,	/D������ ��F<U��yC-�����S��'��#���`�fX0.�o�<�V�6i\�����	�D<�H��h��%��+^(��m$}rmˠ0T�\`�;�ɕ�Y�f|��6$�jD��h�Z�{�-ƕ����5A��}X���b�4,ڒNX)�Z&�=��0
+P�)ϓ<����I�G�NaI5�ߚD�@��?Q����>~����2�'{��k�E�1)f��A��u�><��!�\L��" #�p@���:NR��BN�.
8I>E��'�N�(�B�t
8���N1i����
�'�F(�3,��͐ �KC�X�]��'�HUx�D�d���f/�.vk8�02g��j�  'D����@%�D]
���|8D�P�
/D��X�d�	���b���5����`9D���J�6vHE$T,g4�V��h�<U�	�x=Hы�(�ƀ�$�g�<�����^��t�'�.5���{�gZ{�<i��-�@Y�̀*i����Iv�<�f��9s�8)�ħҧOS�\�T�r�<� ����0�ȡ"��sE���1"OP�0�Յ5L�����!�XQ�"OV���E2i� G�f:�A��"OD�!��V-��ѣ	�4v�1�C"O =�B�R,�����,	RuC"Ota�s�֨~D�Pq�Rm@��"O|0�$���[V�\�C�;*���KA"O��C�M1>m �ac�2I����"O�uۖ���)��
%aމs�~�2�"OJ4J%j�qv��	 �ښl�=��"O=��� �D�R��Hń��"O��5�� T͋8���Z�"O�j�ņtF~��ϼ�T p"O�%xBEC���h�7��,�� bF"O(�k�@�^1T�'�L;;w��"O6x�/��
)��F��Q�2"O\�P� ����#�F =T\�0"O�����N<ԘH`V��2NCDy�"OT��Aυ�3T��P0�xt�g"Oj	�&�nlL�hU"�`h �Q"O�,�eL^�V8���
q��m�"OP��圫~�*�*$�`p�A��"O���JY,�B$F��Bidi"O"�� �I�f]�,��L+Kc��HV"OrY�tI����ap�Q5d��1�"O��J�	�ltU�ԛf"H�H�"Ox�)pa�}�$��fC�O, Ca"O��8��. �Ҙs@�Sw�՛�"O���G��gjv�7iK� �X�"Op�@kMҴ팬Z�4-8�"O��C7�\ѡP�&0�⌸q"O�@�Րpn4��L�0�4m0"OV� a#�>���3��<�Ƒxa"Oj(k�;h(��/���.��S"OH=;�̜�VX�KGo�(��0��"OL�c�N�[�Ή����r����"O�)6/X.���ȵM�d��"O`�a@D\"~=��e	=a�$���"O�k���E@� !״6x-��"O�ԫb'F( p.�7E�&�"O��*QGS�p`>��fl�/%�d�a�"Ov@q��O�U*l�q�ñ?�J��$"O��3S͊0b7��}�� �$"O����/m�`"'�P�G'���6"O^8� [�R��hac� �A�؂ "Obuk�k|hBb���Vd��"O�Slr�n���ˡ�\��$"O�P	�$ �`h	$EQ4��qQ"Oj�87	ʊ]���K��E�"�0��"O,��`�|)���@��yJ&UJ"Oh��.��A�`H�H�5s#�e�"O��BP.A�̶��r͏%��x��"O���
�{I�6�ؔ@��lU"O: !�*ĦZ��c,�	f��"OZ�B��;,x���$9n8t�G"Oݺ�C�+pr����֞ tb��R"O �B�-�&�h�I7�  ��jf"OpQ)�r�20��C#�2]�e"O��ŠX�,�kԉ�0[���!#"O���Ü�mv�	Q!�*B�tmJ�"Ol�ڠOʛ3}؅�% V(Fql��"O����M�~�"4oߩ�}�#"O��!d��M,d��/L�o��Q�U"O�y���<>k�H[��ĚX��"O� MYҨ�:�$�pS�-!(Y1"O�dID�Ӝ�8	S�,�����"O��zŧ���c��]!%��]��"O�LH��) �%��
n�j���"OPq1�����x"M$V�N�ڃ"O>I+ҧԓ; 8�L�%0�hI��O<A;�'͂�,��M�;,P��)��.��$	�'�H�!TK ���8!j�(E�Ja����-w����$�ӎb# ���e�z�d���ZK�hC�ɜ-z������qPy�2a��X%~�u^���*�NҧH���X#��W��\С$��:�+g"O�9�^U���Y""��9�HQ��)>}���y&��v�3����$�55Ѫ��/�O�<1zB�'M��TDT�]ٶ�� �Չ��A�QC*�$����x��<�7H�5s�t��!��t;�R �;�pE���$�������*�uAҩCDB��²U�"O�����T;.�L�R��7|��d0�P��X&��dY����>E�tJIb�^�i��N9Z2�L
�����y��e�(p�#O4J�8��DKU=}��i�ZQhCɗ�y����'F¥8%Ah�yQѠ�0Ne
T��JՆ�sJ
���뇳 ��c�1���:d���Ä���O�=0H˶g��_rNUd]x0�	ָ�q��\̧n�仐���'��9%���h��
��e��!��GnXM��E�:����'�ظ����|�S�O�����R5"T��QB]>Z�b���'<���ϡ6��}���P'.c��
�'�xQ��G/J�)�!�@#SP,�x	�'�!2�Ά�*�x��	LVCJ�
�'�6iB'F�s�ё%P�W2�'�\q�_:>0d�y�ǕC˴��'ǆ0
� S�t���NN�0��5��'������F�v���iO�5���	�'0b���h;&��ŉ ��ب�'�:i��-@*�hQR/[�SVhi��'�>a��mY7-�b���ΤNc�ܹt"�
Qْq��;&�P�q��OfPi�!L^����FR��=j6�Q��	�b��@r#dD�l�=J���$�!��܍#�^���77�j�h� �L��I 6���9'�2!�S�O�L���J�[^��6E��!�J�H	�'mPQ���'��)u��6h��aX�>	*��h�
%����}���*?�8Q@G�!�n= VOD/��?���T�Y�%�5��� �hcn�K����ހXv~���B/O�X�9?��D!���a��p�C��#��噦���_�b�t=� ��Z`�����G?�y2�G�5t���v#��R���#!J���DE7�l���^��)�'E�I ��<�.`����("�e��D�ld��ƥe� �!��M�U�\�SL��#J�����O|�>�ǭ��<��PZ �I/���"x؟�GO��Jj�{B	��r��#�J*j���0צ�&��B��4^^��Ҫ�1B�*,B�B�(O"L�f�Q�^V�ڂ*W�O�I��iU�ܛ��=I�'�RT�5g�E�$�DIJ��T�FnE�^v��@��N��`�S��y��K7$��x�C-;��`��`_��y��E�{-z1�bI*9����W�[�^ܩ�"�B-����<�']H�`��.}�'ee��3&�0P��� oP�G�����I�z�\��hL!G�p9;۴2r�p��
;D��5�v��YΓg����0�X�S&�h/O�i�a3L�O��[E'�^QJf�I:��Ä�>�����t�zT�'�P�p��u�L?�b��#c�Zc��ٺq�,� �B�]�ƙ`�27��d��2���Un�3��<��C�Lx(�����&�������-z5��D�SۛƄյ8V<��/�4��p�qP����O�����T55Mlx[c܃^�F��$+�p?A�ꎂP����hT���?	n����*�I��z���5��AǮ��Z� *�>)�xu�O�C�ƄF��ĩ�H�8 �":�[s
����`��"�X�ѩ�����L؟t�P�&���,3��k��D)��+.v�&�xz�OM�/L,��a�#���P/�<�4n[�d�X��n�?3�P�{��+����m$���� ��#��?`vH9�a�A`y^�+ԥ�x?�* z(��>,O� b�'Q0w�h�fIL���ƃ�"RzS�`m�(#I��h1D�Πe����'����O��u���Ѽ[
���c�(S���9�I8�O
m*v!"��|{�ِF���FI("��0A򯎶61�A�
A�~�I���ɑ���':�J![E$�k�+@�fE:1�h�\�'����͔C��䤯|��m�Sa4D����Ņ��}�$�1#�UC��J^^���|��Q>��T?*U��oX y]�MG��m2bT�' �a�F��$3���A�ӌWV��D��B���#����1��4�a0�a��y`/"LO�xୄ� �n$Ze��P�dY�l-�$@�R�py���$��D�J�,�e�t@c��_����"V-H쓗�5"�f��5�P�7��ܻ��D��x2�P��a�
HP���q��^N�`@��+\ψ���ا�D�ȓd%|�A���_=@�� _�#L��n�`XE���ī^�c��݅�,�RIH��(m���hV��o_�C�>}4,ݹ��ɀ6f�yZ��@�|C�I ��Z�	��HP��q��C��/Wӊ��A�_�T�rg�
H�4C�	o[@ݐ#H�0�b(��:sq C�3��$�W@Ȁ�.����v�C��H*�k�M����Kx)�򄈁B.-��Κ�^�������j`!��B>|��1!	_�Q\��s"�R9b!���<�Ah+Q�[Bv4���lB!�Y.U��q2�D�$M��,@,<M!�W<7|D=`'�+�x�>B�!�$�/����(�qR|���
'!�N^
-��L���x��E���!�$K`�0j��WgHl�X'�\��!�d,`9r�T$[>6�
��uM!��ZU`�L£�9#�Z��/ɻ;EqOe���]�0|AB�=נ�{R.��O�v$Ig��j�<��!�0`�1kt�$;q�(�)����B�JUF��O�UQC���p���T�\:N��9zO����F��#���&�O0
�>Aa%��>i�%BL���>!ASð� ��] �#'A5LOL��A|ҁ��O��Qf�']]��AU�zj�I��"O��q��G�<-z���Gn����|�`VBb����LLa�O=��rө�%Q��W�]p"Ii�'T����Y����6`]�9�"�X�eN9/J\�'qY
q��>�@�UEAd��U�״PR ���`�Z�'���`�A�O��T��QK!�1��r� x�
�J	d�J�D�bX���,��Y}�IQ�Ve�)�LZ]Ę����Q�|�#�E�
^L���D�>Y��D���AI_����w�)�yR�R�`�1K�}G�U�3�
6�?��2����w�ܔ8t�xw�2}�Hx��k����64̹�7�P=o�~�����|K��&+��M�e#H#7b�9$���;(MHW]3�<zK>A6�L���DZ/��LH�'[��M���3�O�9�ㇷX�����I9Q�T����33��\�$Q�7T�� i�a~R��=[Tq���������p��ӵ�Ԓ4���'�>�I�r������l�B�2���2�C��+V�f�0��=pIvL��K�O���$��	&�c7�����=iwb��o���p-�R�r�����L��� %.ƹ9Ul�HW�i|ƭ�bŨr�f��A��1��=�'W\�v��5�x$�d5n�a ����3砤�Rs�O
���'�Ō3��zI@;z&lL0�'�\0P� ]�RU���1vn�i֏��%:E�|��9OJM���HL���X� !��"O� ����7NX��nY,A֜� p�O~ܨQ�Z��0>��[42R@r0�Y�w|�����h�<aP�ӄDQ|��hɳE}��dh�<!$���w�1�7_�U��8�.�S�<)0��I� �5Gb �@�v�<� �l�e�N�[�����W4@��d"O��Xs"Y�xr �e��SjZ-�D"O�9i���y�<�`�g�t"��d"OH @��hI�hIe S�]�0p�"O,Ak�hq,��CM�7��"O�ѩ'-թ��R��E?#n2�"Oq�S�[��-���1.���"O"��0�|�7H��"�-"D�|�ϘI���)����F\(��gG#D����)�")�x8�d���u6l���m D�\[SL��,���a��$��H�tn>D�t�R+�4�iq��Z$V�XQr`K9D�L�F�O�B XDa��ٽ:�L�Id+D�l
�LD�R/����Ŗ�$�#$�:D�Tu���A�l��i�'�#�<D��b�H �P��c�ܫ&<$Б@6D��F�J�\�Hm	`M�d
8`2��8D��3�)؍tTp�'#Hg�A�&�4D���Ȟ�U-z����	:-2
M��(D�X(��E�'()1bb��k�#*D��kRD�>~>֬�½cj��B2 ?D��6@��a�]<a9��Ȅ�;0�!��`��藅�2A4\]9D�[�%!�J*��U�՘o�����/w�!�DܹQ���S�U�R�:�s�O�$4�!�$
O�i��6
�`{Š�P�!���*�b,�լ��+�Dh����r�!����v�2"�'��=�&.�1$!�ӗ]�@0F�E2������"X,!�$�
-ʰ
���.pF:��p^�F!�d@:39^��fa�oGθXV�!��\�G�4����5vYD��6k�!�$��^y�91%�*��8�,��a!�$�|K�4k�J]�j-�bˌ�Z�!�$H JġZ�P���9�KՇ	 !�R�\�t�H�� �|�S$)�#�!��+�r`�V#S�|�|�""B
k)!򄚪5=�3��5=��"�b�3?!� "���j׉J�65c��M�-�!�"@KK q�d�P"A_���s�'��31'��w��L�1*ԙ-p0LY�'ώa�v
˒[)JY1L�,U!
�'�&�#� G�(�Xp*V�ʀ#�'o�ᘁ*�¸�����:>hTZ�'�jܺ�'�$���'\5*j��)�'�zX�G�GUY�3�(�-ceZІȓdM�+/��H[%�Φ����ȓ9��(�#�P$~�t��n	.����9'��!愉S��`��݁_ʚ��ȓ/'��4����b��T杦R�D��Y0PJ�f�63�TՊ��D�M����	+x�f�l�px��V�E�~^}
%ӱ�h㞀���I�S�ӄ`Z�)g�ѿ^��	�'�Sc�'������D����K�Nȃ	6��N��<�B)�=d�8�ON�DP*ȸ�ħ2��9�BA�i�pL Q��%T�Ұ%���I!K�Q��fy3U�M���rB)�T�xf�x���x���Oz��rG�Kx�.�1OZ7n�dEP�O��C��铲iR��rA��-s$`r�Y��6mJ��'ˤ#:w�;��lK�*�p�:!�&�M��'Ҧ��	�'5 
5K���,f�:���jT�	p��<��J0����Ow���΍����2�cH�Z�vL1�'��H���^�C:�OQ>�HB%�K������k��+P��O ȸTLޞ~��H�zvv %>I���~���H?6��V�B��u��(�����C� 
n�!��i�4�
U�>�͟剞v%J�hlܷ�����A"�&�V�����o�)�g�? 
)J���[ư5ʂ��>�3��"4�"}:7�6Ԡ3ȃ
3�ms@m�![�aۇ�d�l�����S�U��0�5�Ӕ<�vY�U$N�o��O�������O]��s�M�-<H��T=�Y[�Onm��aڏ��	M�泟�O_�:u��֠Q�b9s@k����`={P��I��X/�aY秈m,8��s@ҧ�!��Vm�S03d,+�B�f�!��$E���ڴ,� �i�]�?�!�D��c�����˜q�J�+"�ݓ|!�ٕ��b�	',��tX�n�:e!�W yxXyt��q�dX���	Q~!�Ĝ�B���1��:O߼탗!]�+g!�$���\D &l��/�ȩ��=Wq!�DK�D�Z��Sb�P��ј���6�!�$ֺP:��p��z�\B��V�?U!�DݹF�l��e�@ ?�f�S.�p>!�dK$OXi8�`P��=h ̓�I2!���.oh� �/`)�}ˢ�D'�!�dI�{vT`�ȗ�q��%]�!�D͵:)�����OJj^tQebP��!���B���˶�S�i`� �B��!��:���Ճ�	C������!�d�3P�Zcc��c<R��0���J����Sf�W����clΜs{J���^�y��.��y���aI4DR��ȓN6���H�M�� 0��N�v����A�訕bM�"8S�	/f��q��=�$]pa��?ƸZ7��.`����<ငq1/H9{; ��q��h0��~\0�6�20 ĩ��;o��Q��X�<��EY�T96 ����vU,|�ȓ|��P�e@�$�2A$ϵ�ć�#��㗉ה;���ɦEƸ!�Q�ȓh�x���׊7rZuyd��7JJ(���С*�)X����~h��&�rx%�B1f�T�J����I�z� 
R'7oB٘��_v^���� �yQAU�/����G8d�4�ȓi�C�R��� ���'C䰆�<7�+��M�f4hF�I�P�ņȓ�T���D͝E��s�$�sX���0B\t�E	^�lZd��� ��t�ȓ<l�U��j�o�f�s�j�xv�����4�u�ѝwڼ�y�cD�M�����Q��M3��|vr<�� ��d�� �ȓg�&�I"�ÚC�`� ��A`��ȓ1��F�/x̓5そ6����ȓs�Lh`a/@wf4�Qd��-N��ȓ�F�k69]�̅R���,,����O^	���2�0���$b5��N�\����%�<:c��!a� �ȓ.�^��K�-���Q��Šyx΁��ضL���>>�zy���b�.�ȓ;P.9��"T!OvT��p,	-,-���ȓwҦQ��N�NR��R&�'09.ȅ�&$i�@Ň�q���'-Z�6��ȓe�v�@¯K���(���t��$��G�F�8wh��[��� �H�5W\ل�1�J̢�Ɨ�|Z �Y�,�A�� ��E��	s��@32�4-	�ݫP����ȓW	֥��"�9_&���"�zE�ȓpV��və�!�FM��Ģ%d���m}ƹ�t*ӕx�B��M��1� E�ȓX��� ��7eB�sC�xҚM��S�? ���.ݗ� ��'n�>PqJ��q"O���P�֍x(����n��O��*D"OL�Pꇢg�}A�ؙaM��("O�X�������KG�TBa"O�Y���X8v��2�&0���"OjI�c��M%6�1�i?"�yU"OR3Q��+}r��N04�(�C�"O^�2BM3jq�=�0�5�\�"O�M�6B�4(���@�a�2iC"O�	�D����v&�b�Ma "O�mR��Z����v��6e6j"OHL�+¬^5C�ն,��X"O���	L�	H�p`�1]�^9��"O�C#�V^�&�K%d*nʆ<�5"O����Ӊ#H-���јx��"O~li�mL�5>n�ht"ژ`RP��s"O��xB# ,"ƌ�AA�$)؁�"O 8' ' y����[)^�	g"O�T��m��z�",�q(nɑ�"OZ��ĩ�G��(���<�C"O63VA)0ݚ}Q���.Qi��pG"OV$E�	�:AL��7�;tV����"Op�CÓK�-0t%
6׆�r6"Oj��WEY��"ah�U�#�}�1"O���"HCO��� ��ȗ ܌��"O��+S�q��#Bm`pR��u"O^�� �z����F�r�<��'�0��/��x$6��B*�r��'��A�+N�r�-�p`��-#B+�'��}��`��hj�Q���BrS�Z�'�	i��$)��
0�i~P��'r�=�!߬p]��X��՗t�y0�'�4��R��;���F��m�����'��8*���n��< ㇎4b�2�'����G�Zo���7̄1W𾝑�'2<� (T��5���5ID����'a �q�͵"2���(J H����'���S'AU�6�S5��B���9�'�~�S�M�,y��# G�(>ᄉ��'-D����)B�\e��!
�d!lA��'B�x���X��i��ᏽ`���K�'� 9Yp�,��E��	�Ē��p�<A���3(�����(ڟ3ef���O�i�<yMË?`�yш�3�>\���c�<� ��
;QR���/?0�5�l�[�<yBO�}z�����6/�D])�U�<�q�C�RJQ��1}���І��R�<YV�M�?8�Wj	�u`�I�d\G�<Ѳ�A(F���I��,�yK䣃F�<q�hƄ�Vف�\�wIkō@�<aa�Je0���'���R��t�<YB�;M�v=�p��1�*�Â�s�<�3�B##r��0*�+B�z�ʦE�r�<��f��S[��HW��r=��I6c�j�<�!	'��Hj��ܬI�4̑ �]e�<�VJ��<���M�B�M�t�]�<qD�B��e��
�1�<<�'�X�<y6���_�⁉�l����RᢍV�<�УH�����C�@),?�ͺ�.�O�<��I�&`!�)��`�
���-�J�<�C�4bF�`Ô�ͤKi���RD�<IW��B���Q ��KFm�~�<��Ӱa}���ѥS)�I;�|�<ٲ%�+Ql�5�v�ןO���r'B�o�<� nL)h�[�dM���~�^A��"O�T��+�&-��J]G�`�P1"O�PB#>h��@��D�^�v�z"O�� #](��:�N�7+!Ԕ��"O�YٰGG:@2f0�M�'���F"O�l����8E�L<0�KՏ����"O���fū*�#ª��+��`S�"Oj�h3��lF<�`�+H�a:�x� "O��Q�<V�:'H@�Q(�!�%"O`Mq���,Z��ec��H���K�"O�hd��>F�y��倄D� ��"O���1,F°أ��M�,���"O��C�IȐ1��k��z�v-��"O*�AgA��TN��w�>Ji�ع�"O(�6�ގl�t��� �Tl�M"�"O�L�R�V&?�(�j7� � 5:�"Ol�ч�U<9!\+ƪ��Ҁ�C�"O ����%.��В
�%�j�J"O�0Xgٱ=�T����9v�B�I�"O:q�(�G󨑊��̡H����"O�|�5a�%f����j��Z���"O~5��CS��؋���4A|���*O��q�O�C���
���,T�'),�zg��%�A�w(9��'e���,Q�rE��b��D� �+�'O�-� ��31��z�kH0��'Дx���%I�h<��L�W��yr�' � ��E�v��� �����'qڕ�#Y7;�Q!��֖���{
�'���*s��C�f�ҴI�6w�,Hc	�'9p�)E�J�u&F탡�6Z�E��'X�0$	7/� �Ca$b)�q�'ڜ���g�hS�e�E �O�����'�n��eXZ��}�%�E�Es����'��PJr�OB�c��	c�]��'.F�x��)t��Q@�+��	�'���@2��/`� 쪠$�+w��i�'��)�d�ʔ12xH7mUw�F�q�'"��s)B
R�@]xQ䝩g̮��	�')��˦g[&->�0�u�C�YL.H�	�'�\�� 0=3&8@��g���Z�'� ��B�{���e��tǔLR	�'\h�1�Ęb ��#g��X��'L$e�&�ʈl���Q��X�f��d�
�'�*������Jٚ��GB�n�.	S	�'��1J�ʵ�I {d�UK�%��y��
q��0��#�J4rb��5�y��(A��DzJ�#u,������yR��P�� i�㊜h�!)�̓(�y򎌞!�v8Y�ډS#�s!+H��y��KR��Y�=3P��0�yO�;j�Ā����1SN�݁��؆�ye�8 .1�UNS�O�4A JN,�y��L�r��i���7G� ��d���yR�_']4@&@͑E,$���3�y�<?��]C��R�6��-�"�0�ybI�
	�M�m�*0������yR��,j��8u�V�/��p%�Py⎙����ym�(Ѭ���Cn�<`�).$��)2t�"l a�<q�ʀ�P
 b�P?o`����QB�<�%Ƅ7�f�Ö��;X���Sa�d�<A@�B�b� �*A�\����RM�w�<���G$+��U�"�Ȱe�xGq�<� D�2t�T3A�IR`���I� e�"O�Y0i˗tk@equ(�P�4ly�"O4P˵*J /��Z7���.�>�"O2��t����Q�D���r"O.�9R�g��H�Ҍ>%*�"O����k��9�rI�@$�& "�"�"OL9��k^3�\��"i=%Ƚ�r"O�X��[ʀ\mܕ\J,b��2D�y�"�0`	s�b��=���I/D�����'q��Yk����:w�,IƧ,D���    ��   �  m  �  K  �%  b.  �4  �:  ?A  �G  �M  T  IZ  �`  �f  m  Us  �y  �  �  \�  ��  �  #�  f�  y�  `�  L�  �  :�  }�  �  I�  ��  ��   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ��N~��\	?Cv@ӎҿF��(8`����y�DG�|�mYDG1E�>-��'��y"	�*]�MYԤG,Czr��v���y�M��ۗU�~L�S�Q���(�'j6�!�j�Sy���(�GD�A�'�l�`���!AnU1�V�GH���'8 81����u���Q�J�5o|��'�QIE
�8��Ё�۵4jxq��'��aj֕yn~,�0�]*� ����$�O�}jǪ�/G
xs����r�h'�h�<a�IQ#gq�Ї�5^����D`�d)�S��4x�H����V������[��p��!jN}z�ۘ.�K"�ۚ-�H��'9�}bmQ�4�R�YP�Lx�����=��#��F/X��e�%��.)�$�7&٢-�!�р=�D`K����А&%���E{ʟ��ߩ+8�����+|i��pF�*D�� S�+Ī�ɴf�=/��ۅ�#D�p:6���PY�f��n�Yä� D��J��]�k�FX���6���c�K+D�P�Ro�#�X5J�Iu�h	`�=LO�� �6�_4U�4	K�#�&�,�9��'D�@�&o�Hy �� �(]y��1�y
� X��,�	��̒��P�$�Z�`""OlD��+R�..��ǯF��6"O��{���6W���"I�)m�t"O��91)׀bP�̑@��<w���AJ-4���4��.m^��	��Ūm���[�@1D��ڕ��9�4(d�^�2��q�v�#D��+�dE�G��q� ����HE� �ɻ:�Q�b>Ar���}��Z�o�5^��{��1D��8�Ӑ|r�3�	صV9d|&.���]�㉣X+����o��)>(Y��DQ.C䉍>��d�v�	4iP'�7
��B䉣4>��2�-*�ˀ��@<�B��;�hT�uK�#]W�� ����]CfB䉗z���bJ�K����7c�B���qà�$xצ1�"�\$C�ɺ�8���&��-B�u2q-�B�i%�	�E�Vǜ�aEBت�r<S�'���h��� J%�^���R5oK�y"�N������\=����.ֈ�y����8,42�I>� �d���yk�QЀI��#S�B�$$�y��	(�v8��g!}O��8S����yba��'LAs��[o��e{��K;�yb�w!XB�6���@L��yRτ?~'xu���ވK�̘�a��y��l�,#gE���̒�M�ӈOZ��E$���Kdǅ*5wt��^|�<����9�n	�I�� � `���J��H�>���g��Ѓ���V�����-E����]$���N	"}�Թ`�,��=�ȓ``5pcF��bq��u�J(MƆ)�ȓm��HZ���;��un@�7�zԇ�kÌxаjȾKwα�q�ɑ)*�l�ē�����92yK�o1b�؀[@"O��R��*k�pI��M�f�HA'=�ļ>����O�A!%��[.�P����.6��qR"O�$�OG�M�2���� |�|� "O��p%�1fU"%M.tV����'��'�:�jW�@)��\�jJ�!�����4<O��� �F�GoP�c���sBl0��'�Q����)`@ݙ����P�$D�p ���5��y8f�Ůb�U��7D�t�4�F2`1�	Ĭ2��X�A�1D��x��D�����< ���+�d1��n���ӌ� '�-Y�_�i�ł��0D�LhUDI5D�VHh0���v��1�f/D�� G.6-N cuc�;Y򒙀3�9D��ä]�&'�qFQ�HmLY�a):D��I�8r�R��
f$E�"@*�h���OdD̀���ػ��ч,���	�'n�t�g&�Z9:�����rzvR	�'b��5��0YP�x�S�'B�I� �20�!A*j�H��'H��y� e��y8A�$_�ݨ*W��y��y�!J�Oj�����F#�y�h$4��۹@�,+d#���'Kўb>�	����a�yR0h�'���-*D�T+g&��u�L=��ϓ(��K��&D��lObi��b�#M7���ذM%$��ӏQ fnM!�@��$G�T��b��y�E�*qZ�h��FE"Z�P��K��y����
��q���;��HI@�U��yR�Q�O:F�����51VX��/Z��y"D3g=BI� "�H�K%A+�y
� ������H�$��G��&O�(��"OT�r��צ!����'�<�T��eOޠbI��(N�Ya�'�V��x0:D�ۦ헣X2�q�˘�+�@� 5�8D�<2Qo��{^����8~F�{��5D����i�)W@�厇�A9���9�@���O#|���Nd��@̎�(��'%��X��E�k��@rRD�?s0�u��'�t��o�# H,���Y��x�h�'�6|�V�q���&�ř�Lŋ�'V�������f�ԗ �<=[ϓ�OQy�#԰~��8�,]4�] �"O
���b�/H ����( ^�z��|��)��j�N̘B��8�P)9H�'KXB�ɪ�B���OE2J��H����f�C�I�U�@��E��Ph!�c�y�C�	�"w��&�H�s�z�XVDj�B�ɝ]9〈sl�
$�
�(�
��Hy�B�I�7U@8��E+G"��h�XNB�I3A�({"h�*M����#\�4�XC�	��"��4�áAJH���&_�B䉺j��,ZW�	�2�T��E]#�B�I�I��iǂ��]�`���5t�6B䉸B����ɑO
�i@��z��C�Ɉ`�xlt$в'3؝���3��C�I� T�vm� v�Z��;%�C�6-ƞ���(�2V_^�J�JK.�C���8����ۢK�h���/�x��C�-n��p��숱OQ|��'��w��C�ɺ]h�sgF^�@.RU�&(E�sZ�C�63��:D��?�0�ٖ
�}�zC�I%X��sg

QR�L6y��B�I���-��E�c����2�P)�B�	�.���Y`��3J. y�!�elC�I(�H��%�������c����hC�	$Ş�+3�Ǝ6���p�#�B䉱~*�����Y�|��%�r���w9�C�ɥ]���fd�?nv�!�pÌ'غC��'6"���r�Z�0���!�!X���C�I�_��mS��#8��EI�"W�,�*B䉳Y���T�P��
e�eMPB� Ĩ�Ѐ
^�Zjq��n̩=RC䉖��D���г	��k���X"C�	~�z��F�F����f޽FC��$����W�^'�\{��/h�HC�I�+
�ϤE� ���O��C�I<R��k� � ]N�����O�2B�	4k@,�C.؝&]�3Ċ�B�#XNԒ�S��j��Q���!���$ZND�h��/Č	��F�e�!�G9i�^yP���6�"�A��v�!�$ؠB�ڤPtJ�9��x��;"�!�DЎQ��@��a66�ɤ�@�3!�->���P	n{`�9N�+Q!���m\5���C�2]���mJ�Y!����+5�Ҟ5F����mɽf!��R�Lx���g^�B�m�4J!��Џd�����3B4}�ek4�!�$
��8у�͋i����1HO 7�!���7N���B�J�M���
\�9z�'���3#��x�.�%��3C��Q�'�н�R���V����EK/=9@��'r�a8��O���dT�/�X\��'㞤#5M�ښ��P?%x�:
��� z�f��5R$9B��^�(��R"O��K��"9@lAAh'u���"OJ}A�#�9�͈4gHsj@�c"O��/*�8P'�pm���7"O��ڰ��p� 1�f��_ObHYu�'���'"�'�B�'�b�'P��'�z�(dMKo��I)�l��(K���D�'�"�'���')R�'��'N��'׬�d��d��sN�W
���'��'���'���'[��'aR�'*a"�b��}�ش�S�çR��"A�'1R�'~B�'�B�'�2�'��'?�ðK�!Y8�10�i�
$�� ���'�R�'��'x�'N��'�R�'��hz0�Y�t����"ql�4�'L��'���'d��'���'��'B�X�����AA��\7����'B�'�"�'JB�'�"�'=r�'	��E9��qC�80�}�W�'�B�'+��'�R�'/b�'���'���f�c%�(�aC�Js(Ju�'���'�b�'���'��'y��'��P�Ad-������33��TZ��'�'���'�b�';��'��'��▃8M�r���l+)��=$�'R�'���'�2�'���'���'�i3Î-K�����G�J�,�w�',b�'#�'���']��'���'"=�Ea�mh�kwƒ�

�Y���'kR�'��'���'���rӔ���OR�ԥւ7� ��� XAd)�ay��'b�)�3?�T�i)5�7�U(I�z�kP�N��X��2��D�䦵�?��<	��G�P�ǅ�#��tP�&�!6-ZHy���?�����M#�O��S"�O?I�Ys�d4�6�̽v��9�b+·Ԙ'�r[�$F�H�2S�t����'?3B	`R%�y��6m�9L�1O �?�C����6�'x|*���C��d�ڭɅ�ނ�?���y�Z�b>]���馡�I��:Ǣ�M��M�ĉ�ZwJLϓ�y��O�Y���4�&�����E�*��a�ܘtK��Z�'���Q򉩿M���N�:��s`�׎Y^�� �OP�%�0�����>q���?��'�I�_�>m����A��F��<LP�?!O6i4�,�|"o�O�,B��[e�����R�%���3��u�-O�ʓ�?E��'��A��R f���'(d):Ha�'D�7��7����M+��O?X)�rL� @�2#ˈO�
ਜ'��'�rE<Q�F����'9���J)D�|��	W�K�ht�vG�^`�C�ɅY��<����d�!8�
I)(��C�IR0z�CU�Z�2P4x�ę(av�p�#=Sj�q�3ā�_��a��]/:`Sd�!wd�81Ɯ<Ip�4 �0M�S�`m��jߏx��xу�ݹa��`�J/v�΍h��7|�-+��L5��hڅl�����
r�@���v�yr�P=X��S@F�A ��@x��@1�D_�~?��9�P(1�e0Î<D�H�S����+G�3cY1 ���rC,i� I�;F��h�V��qH�F����m���9wqR��q��n{\�:���S���3��'�t�0E��y;đY�;��P��DYE\I�v����P���3�$�F��e�)�d�\6V���c��ȟ?dȶ狚(u?:�v�-OX;׉�������h�	�u��'���8lގP�I�p���Kv�$�~� D�\-�����)`h���dT�:��Z#�'���*�o����d�n�b�h%�ӹJ��؅�I�!|p��V	��%�QW/�(5����ɭl� d����M뷶��,O^���<ª��iuZP�#@(2�|A��T�<� �"�2ɖk� ,�U���va��I "���T�i�9��@�2;b��3���U���2�#D� �(�^m$u{�E�EQ�0���"D����c!� ���ؓ#x�H	6D��)�/ժt�r��7W�'(�0��n D���Сb�\Eh�UVi�H�+=D�`i����g�d,���/H�z ��;D� �&,�07v�)�(�+;�Z<��`4D����=8D�S�j �l�X��qn3D�0"Whʝ�<Yr��H�����,D� ��I<�e��fR�>��I�$7D��نBV)"xB��4��g�&��A4D�ↈ����!3��
긅�g/3D��b4��:>Q��*R'Z�[��-D�̈�M܉,U��s�(a2�y�9D��c��D#".=�w�B4h����5D��
�T2�P�i�����s�.D�4�f����ՙ3�8���Q�D.D��	`�4<oZ� ����@��,D��re �)��!{7�I�f�X)��.D�X⶯�K(����<gN4Q��H8D�� ����<I�Xc�9 4
�"OVp�r��5Vv��$ቐ\�&y�!"O�xcՋJ�=z�͛Q �c�"OؔC�+�`�Q�թy�\K�"Of�O,S e���"Xcx�8F"O�  >L���̝Jb�5j�"O����~�$�/�q]XE��"O
-Q��
KrU0�Z.=C��a"O��0�)bJdTy�/F�ӼeB�"O0D�#�O�"�ȁn�*Y�vI#�"O �� ��zR�HP���0K���$��5\O��B�һ`#��@�+ɺg��h��';��F�S*MÐ�D�n��q�m٩6�:B��A��󏛆<]�ast�>��#?��ؿ?\4��~��+|�.��.p�.X��)�S�<��W�`�D�G.ĦK�B$�A{?!#�N2�6�Zvh�b��2��m:���2��xM�i���ǣ�	��l`D���3"�@PŊL<'֎Y�N��^�&H>H*X�������ቇa�f��E��;i� �#c�-�X��䆠 �<�1k�c���K!���	f�)�'��8 F�3���T���͖U����.��;��͎f��1D|��ɒJ���c׍�9gR������4��,?@���)X�m�>���K�1�y2aբ��oJ�I���0����Gk��
gZʂI��CM0��6ił�h���c�*SX��Ë
�u�ұ�d�'D� {�(+-��] ЋDw���Z�E�'��޴K�z�
�O�K�i�O�"<�s��V�,���N%C��!��XX��JLq�N�ue�F1̴9׈�1F9���A`�v}c�\�3�-�.r�f�$?#�9��)C��uE{ҍ��8a�غ�ߨ/�(�G�������L)oW�i���Ӝ8�\t:#l�9�y"�"���v,�<8k�b�@��y�f� *G́��f�D`[% *�#��5PT�R0)���UNȦf�,��
����a��+��L��#�Q0��dÚ�[&���̻)Ur�'"���ቒO�z�q���ef`�5�O�	X���$�$l\�}��9 hX�g*^��&91�B�x�0���:&ℇ�	�Bt���GƂ�OS~�c���HN$#>AV�3w}�Y��aڏ1��Q?���	�.7���3hСKĎԫb0D�l�"ӿ8��{��K�r�zx�@�l����"��w��u+���H�m����$"��NR;I�y��S�b!��$Y4\�g&�d��9A@O[�`�0M�AI�O� Kr��3Dt�t2�?#<YuFGET�DvjX�-� YQ#�2�O��g�Ҋs�:=��ՐLl�%g��`Bĉq#$�3 ?\B�	�|i��ɢ��:0�D�!-Z1t"=aԈV�tI�eS�b8��O��d3�8F�(�x�N��\Xn��
�'A�'��C�:]XP�����شvq�Qt FG�S��Mk��W��+S�_�@�Q��@�<�"�ۜ |)jEM4!��kqNw}�CA*��Ih��ڕ��4ApLe풦?ɜ���������G7"xᓭEe�����Ͻ��C��CM��z̬$�i��e[��#=i�e��f�?ݱ`��dD90m�D�:L��-D���c���?&�cB��~�L��Mx�,�����$������f���~�����	�l,�W��y��ϯ/�| ���.az$1��aϦ��� Tv�'�'�$���NA(h���2f�a�Z��
�mB��7���Zr��!P�򱙔��7N���"O� {�&��$�����d�k��ɫ��."[p>E��C��i)&��IF�9t���wF%D�H��F�Se�}��<���ەH�>)��˿o�`����/}*��'媉�␾D|*$Ӑ�i��Q��'e����-L0Ry�ك�@���,�����J\��e�X*v�'��y��ϧE|~�	��P�aB�2�-�>,����0 �7a��m��#h��� ũU;�M*�'A�M����Kcj��5��b�֙��O�՘�c�S~2�R�,"|ڒh�Va�yRr�!P{���X�<� �u���.c�����o��-;`I9E�Op��Ĵ?��m�C�<�Ϙ'�v���E�2#�����0#s��Q�'Av��e�8���KT�_87�����ך'v~�h�n��'�'��P`h��z��5��h�EӐ�:�#\�a����8�L E<!�%.Q(j�^D�$'�;<���b���	�q����J�0z��f˯��^��H5��djrG
�u�'F��N=����4�4�a�v����'j�
���3	h��Ye�F�B�L��TŜHBWG�>1!�٢���
+�x���P#�Ҳ`-��9�&�)�\�ٶO�Q!�gN�{~�@S A�#>�@��a��t�v�_2(� Iz���S!2Ms�&Ӽ���	%"}8�+��ʹB�l������?�`��jg
�Ě3�XQ�G�X?��49��A����c!?�5�C�^�s[��E�@9�0>	FE���i�D��10y�Y��W}E�rd���ߴU`�|BM�:H�I�y�O���#�ö�X�(w�Q2}H$	�'袕@�1q� ���Z�W�.�р&J9A��� ?��9O��?nϪy1�r���6�~13��? ������6/����D��I�L� �G	��-6ㇹ+�L ���V2@��� �~��&��YLn$��K,Dx"��` �3D��.�|p�E���O&�͈�<yc�mJ�ϓ!�����.`26I�u��/(��ُ{k��"k�T�C�#_\Pu�%��o��HI7�>ᆢK�h��DZ�y�����~"�i��4��њ�A�6���䀈&<]Dxp"O�\j�)Ź|�4[d;tʞ��$�܅fR�͓��A�4O��T?�O�K�0���p�� �ΔPc%Ű?��@�p�H�Js�U�j2�t�OC3�|apQ:OX�DYW��LUd#<�-��=t$)Ո�0O��I���l�'��7(Y�|�yx�Gҵ��iD�H�t`���3�dK��Z)p�g�f��$P�c�0��(<.y�YB�o�d��<q�p�W�"?��" '��O�)��4J�	Wެ#�/!��Z�*�jL�A@E#Y����닢 ��Īv���<���!l9�)����g��K���(
G����C��B�@��p؟�����djF��0*�|y�� �̅Iu'P�&�S�
:�(O��!AV6t��Q�e�+C&��q��	,I2��a ��S�X0%�~�1�ͽl��Q3Wg�L���Ñ�j�<ї�t��Aq��x�A����fy�}���a�-�6�ɋ��L�N�$�P���wK�|!C��E2!�v@��Cf��	BFl,A��c��`F� %��a��Y�8�tJ�5�Թ��"U�\p#C�<D�8�1��5z<�p�٨y��9�U%�O(=3T��M����� k'k�;V4Ĕ��G#^��0��IHq~5�aG�<�'H�K�hQ�D=װ��Oj�<aU��*���@��N�!Cj�|�S�ȑ�"�E�:�?�ib�0D\��*ܤl6�Lb=D�h�2� �?Ǧ�2���7q��j�a�mcQ�wd:�D�x�����  �d	E���ݳQI
�6�!���[�ƉD*&Bɺs�O��HX� H��d�'�u��@�% ��b��p��=��i`�y�5O1���$X�.�i��V:s٦0K�"O|A��l�`yh]�R�^��P��I7T> �q���י0D�Yrs@�o��<��.-!�d�@�n�`�D��'�F@��ՠQ�@�-VL�c�"~n�.{���`h�G�̬A��Ż[&�C䉙30�"�	Ym	>](T	G<04�H�iH��'|f�i���:E�h��AC^+=�ڑy��B� ���O\xB�]�7I�,��']vk��b�"O$���F�R]��X��T��&Ô�	�\�H�p%a:�'=b �
�CC�CM�8ɢ	ۯ/��d���V	�G�Y8)T��39�l�
a9h���/;�)��RE+��<�2�,�3p=$4rd&D���c#
}����ˏ�s� 3��>��)��=�����/(�a� Iυ��|�'-��R�a}�GBae��	�]�8���1yh���,ת'fC�I�[>}*W�W��F�|"=��/ӺM?�eΜ3J�\��@,PI@��� 9D�`bf�F7aIiƄ�/@av��@uӬ�� `S�S��M� T�jd�B��-�Տ)����"O(!蝏E��C$
]8���UX��n�0>�$��m��� $�֢���#��fX��1�K���y�m߅0*���X�C��x��V�yC>Qt�� AOAh>-��j��hO��Ӈ�Ӧ-}�!
J�n���#&Zt'�B䉿��@���a��Ա���sGXB䉮,�z�L�
Y�|��L�e`C䉖Z���L؝p�d|�RMޣmʀB�I)���:�e��}~��e��5�dB�B�6)��-�U�t ���+�C��9�j�@K�\F��6Y�BC�	21�~��&)��d� `bsC32�lC�IvѸu�*ơc��!K�D�4C䉋X���k��C$rO��3�#�L��B�I
�D�Z�̒�\�\��$��$yI C�I�|��À�9y�y�'uJ>B�I1X"@K��� Wq��	@c�C�:t��+�R�?n��P��ނ,i�C�ɸX_F�0'�=ۂĚ��X�.��C�I��}8�`A�c5 ��7�E�C�	1z�lI�٬�q���T=3��B�I�F���+���t��#�E�<�B䉳 ��ā&\�.��XQF V�B䉠5<@��ᢍs�����&:�,B�ɁyT\q�_�&�4cU�X�B�7u�\!�E
�)�24K�0�FC�	��Z,��+9U|q�K�6!(DC�I�K�|���Q'<�͔+�C�	�(J���Q   |8� ����eB�I�pt��$i�
O�L؊�IO�)��C�	:51F�s'�.h!­Q�rA�C��!v�̐)�P%\��"f��q��C䉃6ʸ����Z�8	­H��
-9l�C�I	P>��)�OI�4j�D���=i�C�	�eZ������J:JH�ԉ�1j>B�Ɋ+�⡒6 �UB$LX7�Q�B䉣��� ����/4�"`ʇ�B�	�dI�%�	L�-Y��.�C�	�1��#�!ȏdV���@D�!"�C�I2[�4��*46+!��XVC�0&�l����Cs=4�
��9�|B�I$?&�I�V-H/3m���¯N4li|B�I�oX��`�A�;R�Y�C�2N;!��Z�6�4I���zN �zG!-Z"!��ڑ1�%�B㗕C��kD�[��!�g�����Ϝ*�p{���8p�!��H���ˇ�5"�{4����C�	F��5E���<�1G,O�#WC䉞)��� B$!&�{cHF�B�	�p��H�@�w�H!)�=CD>B�	�w�L�c灥<"�2��M H�B䉷P�p����{wF=�1·o|�C�I(��@�oV8I�4� ֏�M�C�ɨB����dIȶgVI2�IK�K4�C��=1�j�Ss��2S��k�����nC�ɆSMl�`QlK�UwĤK���R�B�I�cȤ�;$m]�_ߒ��"HT3>2�C�ɟ<w^��4%I�a�d@T/F1M7rC�+%��C� rBQ���C}�4C�	�S��*���6 2 ���4-2C�Ɋ(�>�sDI�~�"��>y�<B䉴�%Kۅni �1�	�4%�N5	%"O��1*'�� ΚU�7*D�� >�鐻4E|����	>����"O��a��I�:Z2쀆t�dA� "O�%�r�G6GG��;��E�q��"O���
�p�0) �hܲ)v��7"O,;��IQ�q��
�B\�8a"O��+��K��\Ҵ��_|m*�"O&��d(�;T|�"��e[�	9�"OV���֪)L�,{�5g��y�"O�q�v���Q9��y�㎟q���"O�̙���`�����jn��"O��������Vo���1��'���
�dƖlz�ӺI����	�'6H��$��^)1W�P\x]�'���5"R�k�t�qK��M(�y�'�v���k��R�����R�Do.Ű�'�����X�~�1q0C��B��:�'Ơ�ZN�/d�(YՇ������'� hFՐOw�x��
V��r�'�������?Fb`)��&$~d��'��(����L�z�C7���y�jÁD�� �эS�>�R�0$¦�y���:CI�MGLX�P�,?�y�L�:2k�؈6��C	���n�6�y@���[�M�<�֝�am^�y�c� e��cϥg@�ifJ� �yR���gƐ� ��Žf�e�Ug�yb?9I���F��)Y�D���
4�y�$�� .��uj�@����f
��y"�O�spV)����&:_�X�lD��yb�ݽ��pXG��;3P¨!E�4�yB�9>�K�m; 8��d.���ȓF<�+����M�"h�pծE��W�0��Z�0Su�ߝ2@8�ȓfL�ӇH'9�]��N�KEfA�ȓ<ZЛ�b�(�"RB [����ȓ�h|���;DT���`m�Kj�ȓ\�q�bė/l%�p̘�? f���FT�ydE [�m����$Z� ��>����e���<�c`�K�'�����o\u:��G��G#N<�1��g�"��a���bPcW&�n�48�ȓp D�"&��2f0��Jrc����ȓPd�2a���mB:���k��Sz�9�ȓ �nl�Bh"s`�\Z��K�b� ]��J3Z��%H�m���g0u2�4�ȓ�:�r�XZ�6��׉�+ �J��ȓG�P�I���5J*������EuDцȓ��[��R���5+�����a�������`�%���2���Q����j9D��xҡF$Zu���'B��P�F4D�(��*D�R�2@��ϲvK�y��,D�P�3�ʕ�z�zQI��y�֐���*D�T� �4]l�$1��5���*O`e���
+**t3�FRx�D�� "OR]���O�|�R���˒s8�\Z�"O�k������ҫ��a`p"O�����7 � T:uC(^d�"O�I��%��qi*8:F��d���v"O�x���� `�y�O�fHЀ"O2�3�ϋmb�	����3a�H��"Oڸ�#.�BU`�.�Ih, S"O��8$��tf�)C �*�n�ib"Of\F�X�9\J@�f�.q؆ݘ�"O� ��(Ҽxj��y�$E�j�@	�"O� ��R/X�0%�31���,	)6"OND�a��dJd���&��%�T��"O�k��9�0��E�P6d��4�"O�t����?,c>9S"�"4���9�"O���Ɓ�Xl��7e���a��"O���p�\d�L� �X�E��"O����WK@����-�|9Pp"O*1��m�,OP���#ah*�S"O�z1��l������Y5pe��yv"O�1�ѩ�_FHUH��MIY��X�"O*�����?O��Á�vN0`T"O�����=s|�ms㆘)}\��"O^��SOAQ��0�$���}��"O�h�â�ZÎ=�ge��~��m�"OT���T���Ȕ�Oڢ�����yr
�N��Z��:H/v����y2��?,�V���-EZ����܄�y2�
h	t-�� �V\P��D��y�\�'<���p��`ryj�h�/�y�l��()D�acLM3�!*t�+�Py�g�~1�p$=2��a!�]e�<I��-� Q��%��4���/`�<y�)wj�|A'Ǟ�d�$P��,^�<y�c�7	*��b��z��؊1D�U�<�%΢�*��T�O:8-*l�S@KK�<�b�Χa��]���Ӱ|�@0�d!D�<$�:c�t�2A
�-�
�x�<�ҁ�.�ި�� ,��U�"�k�<A��ց[*(xI�k��.~�yI'!Gg�<Q�]$���F��p�4��@O�<Y��_���C&�K�=S���f�<1���m�������8% [��|�<Ab����9Ƃ�n2~�pCA2D�� ��r<4���@�wF�j�0D���#8'K�4h7k\� $D�	�,D�ġ�ƕ����,�1[��]��(D�����,(������34ʀ�a�&D�pJ��^�1A���B��r��a (D�xxsM�����B�B�0C�;D����d�:GĀ�JB�߳Q:yP��-D�(H��o��\Foܜ>2� r�>D�T!�	BU儔��-K�"D!0�=D��A��X71C^�!v!�8$L p�M0D����H��|0ܑ��]��Q�A!D��B�,�̫@HP:^r�i��?D�p����#
�و�'�43���3D=D�D�蝹z!���2ݝZ�V�k��9D�P��[-xrZ��BKի)?V�B� 6D��+Q��`�~�S��ҮWWJ�I��4D�<�"�v[��8����h�Dp�fM2D��2J�e4��:��Κ+�*�@4D���"hE�QN	�b��mdD��2)-D�[V���ΰ�;&!��2�xY0��,D����TXL�m�掏�G�,�Qe7D��beC�A�T�S6�v�4X�u�?D���E��H��=iT�������=D�Xpo׷f\q�@H�}���h"&D�4�0��	Z}�Y�U.E�$�dٚ@
7D���(��S-��Ag�A>>LH���L:D�@�r��52�
���ŝ;	�.%�Q�8D�LA�nR�"$R��q�\���x�b+D��c�*X�r ��Si���l��d4D�Ը�-�&!��jS��-�n4[�(D�h��ϻ7��U���?pA��f%D�� 4����P5+v��v����yZ1"O�P��ҷX�hɠ
�>5��@�"O M:��6'����(��LΨ�r�"O�X���m��h6H��m,�A�"O,���Δb�c�fX>�JyJ�"O��0�aS
�B�k����!�"O���kR)>���R#P�4 ����y�l�K��h���< 1��
�y�K.�ֹjǭ�μ��`W�y��RI)p�0Q��5x�8�1vF���y2B@� K6�a�'���r٣Pϕ:�y#D Mհqpd�= >��z π�y��4�p5�tKA�{��1�@�H��yR$͹+H�h:��1 �ع ����y�� r2!أ�ߴ��t�r�1�y2*��p"�A�M�I舠Ҭ�0�y��	�I�p��H��{�
K��y�R�L{D�L�x�\����H��y�cQ$��m+d�[�[���N��y��HD:���J�X��٣ӣԇ�yB-�"J�`�B肳HX���o�+�y�e��z�Jb�m�p9 ����6�yr�@'r�fU ���`�l��G��y�H�v�d�1F떬���D�yRC��G�"��VJ�;l0` "�yJ̦	���� �43l ����y���ę�Ae��<�@���݊�y���dbdHGù9/�Eɇ��+�yrfZ�% J��e��35�|U��,��yr�Տ4gN�U�91�b3�k�*�yrgR�b�*�!t׼"X��֨��yb���
TLE�ɉ�/�p 2�&ג�yB���o�Pq�0�ӏR���+B���y2�<v�b0q�/.J�<�(b���yBH#*�!�	<N��x� ���y&��)�0�%ҵ;d�r����y�a��N,:%� C"๋qǅ�yr���d�+�#��h��9 6�T�yb�F{�FRG �2D�+Rm��y�h�	U-�qJ��##�1��oL�ybJ�i�h������]c�A���yB�]u���A��>D��J��yℝ�&����U�XQ��S���8�y2�Sw�8p��'��|�9�G��yB�����B�ֲ+�� �����y�r�,���R�䠸 EO2E�C�	3v�:�j��)ŮT���:Q.B�ɐ��i�VCV.(W��S�a���jC䉇 Z�5�H��*�h�L��FC�I�s:��u(��������F
�C�I�B:�A�@Q�C����be��tC�It�F��P
�F'<t����;oC䉝h@(Тe��F��)a��0h�B�I;e�����b�6i����Ԇ��A��C�.<��I;F�ޠT�X��YU/6C��1zuD��	�}×��*sm�B�d_��˵�̞5R�M�W�
��B�	�V�F�q �L�A�����z�B�I�t����"�:��$%Z3X��B䉏d��)@���0�D�ڬ6��B�I�s������t���qB�����C�	}�9��m�=(=�pxR�©A�C�I�.Wܤ�``̱paVK��C�	�C^j��K�C��1R��'L?|C�)� ��:d+�%[�wy���>r<�A��,����NFN��Y�ٻG����ȓ^d�R�ǕIfȍ1���0 e�ȓ3��8�MP� �@|����_��<�ȓY���ʪoK�|��g�]�����䨔��-N=�й�G�|���ȓG`�D�#V0[����E�W�x��ȓP�~�F�����.]�,��Y��m\T�Q��T�
�Aǌ�=&��T�ȓ:���������$2$jG�u�!��g�&���-(��|�`+2�R$��SHֈ�a��MjX��&�P 1�<܇ȓs�L]�#ɕ�j$�1�o;�:)�ȓbDvQ��+U�4ܠ\�2�̵y����ȓd��ȢGr����ɳE���7��@���d��� ��հ�T���=,�х��*XhiPuo��"��ȓ~��)�7��Վ4 ��A�ט���p�D ����(O��1`��޺-��E�ȓ
J��	A�?����&O9l~�����p�ٵ�֮�f�1��L��4��m�ːK
 �n��K�\�tB�	6MztCV�LM���U��o��B䉤^:��4E��|�`4��l�0v�B�	x�=4�P�xO�Q��@���jB䉃z�ey��NYZ�zu%�1�fB�ɺS�B���Ȇ:�n��I��<e�C�	]4>��'�ݠB$P�Sv��U�vC�I�8���B ^'�����v[zC�	�|G�8#C����!��/u4C��.s6M�@��5U�X�y�H6�C�� )a�� �&B�$Z����C�	�k1nE���"K�eÅ�:U��C��6z�~��)	��"��,�zC�
r�� @'}�J���ŨHlC�ɥL��`�WI��w0q3Rg�)d��B�I/Θ	qM�hfnS���&P�B�ILD$H��j�/[�j4�#d�a�B��/n�<�;d �����*DF�C�ɣr�!�KW�32n�h��5<�C�	��UUi�*df9YEI�*P��A�'���p!��bJ�����6|A�eX
�'|6�1Ԋ�-@����GV�l��!3�'��@xf�	���a�P�A O��p�' �;���F!N��gቸ^�JEb�'0谂fO��5�W�[�Q!���'��y{�Ã�n5Z�A���=Pͮ�b�'��\�,Xs+X�s���*B�QY�'o|����Y���;ZQm2�!�K*D���A�#�|5)�e�5@�X�P��5D��d,�PY��2%
�^[6��S@!D�H���Қ#�(����J�n�2��"4D�Rq�����I��	NmH��7D��s�وB����Z9l)��s�+)D���V�*'?�]h�#X�L�� ��K%D��3V�BJ\9@6O��VȔ�a&"D�XI�IΫj^M�V�5A��ٷ"D�<kH�8J�X�����FdD��ue<D�xR���4��҆�i�\%8�k8D��R#���U����.��J���j�j5D��+��Y�z�hU��'ױ�M؆�1D� �u�l�x��c�Ƿ}S�����/D�h�è�(�ٔ��ɨ�9@k-D���FK�)�i��E"?\��#%+D�� 6�����8:v�;sb��(�|#u"O8��&� Ԝ8& �-��M*"O: a��5�A��Ё!�<�8�"O8�Pw�WP0x�*��lQT"O���.^!{^��KAoDQ�2��"O
�C��
#���v,�OV�	�"O�I:���"�9�k��x䞤 "O�]s��L�y~�l�u�ܟY�庵"O� n¸J�*E���h^�i�"O��Jc`yr��e!��~7���"O�1��Ʉa��L���2
��B�"Oր(P�ݔ6����2m��zm@E�&"O���2��e���u���p�D$q6"O*I��.�^�pj�I̚z
X�&"Ob5!�)e���ে�6>c>ͩ�"Op���M[-el�K���hS���"OL\�����&е9�Y_p��"Ob4SP@����}�2%[�-WD0c�"OD%�CZ�*���1�c_�Lb���R"OR�q&�Жe}���f��\Ɛ��"O�ՠ�d �[�gT8xC��[t"O��Q�d��
_�aYC%	,x*~E�"O����őR]��A$9-I��D"O��s���~K����B9?E��R"O,�e �%;�� �F��c����"O��G &9��Y�K�5aK�a˥"OB�@�"�aod�`��V�^J�Xr�"O�(��P�&hd+G��PN�A�"O����	��4�haI%h^�MD �C�"O�)�����f.��!*�I��"O�Ԃ�(Bn��Y8ǆ@�j@vy�2"O����H�C��eR� 2�hS"O(y����"��9��E��;'��0�"O�vc��+Ь�S�Q�9��('"O,ѰPI�t��x��eO0$Z=P�"OD��$�ʹ0MR}3v$���}3"O���才�^���0�,;2��9r"O�8Y�����x9y��cw E��"Od�k�I	e�5�cbu�%b�"O�t�!Ęm���t�ͼ	Q�p��"O�T)��ƒ̉CO�l(@=� "O�Y3��
-&��1ar�
2T��"O��2���O�^�9&�W��>��"O�A�q��
}�t�X��-?�2� "O�ӵ��,3�:�8�K]�3���	F"ORh�DMP�i��F녚d��T)w"Obx8�ߧ���dcQ
v���Ie"OF�SD	!c׀%���Õ �0���"O���q��=b]RD��eH In�@"O��Ԅ@@ò�0uC� 5��!�"O�x��̄�{�|�*TC��Ij�*�"O�hr Ǌ`!Q����m2���"O��J�'�6KghT	�gĖ|K�%�$"O�Jv�҈P.�b�dT�8��yu"Ob��� ��6@])f� h!n�҅"O��8F�X���	Ӆ
�Fy�Ԫ�"O h�V(�G�$���C!kV6���"O앰B"�D�|p�1O'S�	��"O����X�0�~�����ON�ܒ@"O8�q#��j����b$I�52Z%"O�����!6�����B�} ��{�"O� �pDC.T\���!!F`�*8�"O��'�zkt���/Za焥��"O�mz��ėeI���$��4���`�"O� L��꟭I��8�'#I�G�.�8�"OB�f-��D �%&�\/`���"O��K�
 �E*P�ч��`P�Cv"O��J���N�Ȉ�!Js:(#"ONĲ5�΄\�4��o��qmZT��"ObP3��ߩ�-1h��4|p���"O��b�n۔Jv�|�2���fR�	�"O@ �A�.Hzj,�&�&(W��p"O��A얰wJ���%g?�%"O �&M���,(W��8�Pp�D*O���H�b�)A1G����'"ы���'
f�҂
ͱ7�<y�'���Y`���!i괚Q6e�! �'l�-�(Z����o�7{U���F`$D�Dagd�)~A@�/ ���ɡ�� D������'q3�Dj� �!5��њW  D�`0�ƮY`��6\�
�b?D��!$�sͼH1��޷[�*�Z+3D��a��С/��c0��
`��M ��#D�H�Q�öP���aW.5���D7D����Μ#�@�z�ր/	 �`, D���t���s�lЀ7�H8E��!HrB D�,�W��+�T�)q@S�)�p�C;D�\���-g�>\�B���bhYc;D�,�sM�&j�xU�(�K��@J:D�������F
� "� �,����:D������n��Qc"�p$:D�0Z#L)8�*a8��_�W�x��9D��H5�@8($x7`?\אy�:D��h���W,6��GI�8i��7D�h ��)�Ȑr�>\{�`tC4D���f�q�X��f�U�X(f`�c.D�����xb��	�~��k-D��Xr�����%IU�4v㨽q�)D���3�ʻ��i��c�7{��z�J3D��ۆ&[�G3�KW��]X���),D�� E�_�K&@���*n�Xq1��)D���0Kϵb�&����A�ص#�2D�g�U�>��HxÁC�˪�a��0D�x �Y�0 B��#ύ	4j�{F�/D�T ���5h�BX��G�8��%`"D�0��J�Iv�k�l��b8 Q�l>D�dS�`�G��@���ɑy��š'@/D��1r�T�TT!*�
ڋ]F�ܠ�G0D�\VC��d(�Ps�%�kGP�h��,D�X��G |︸�Q��.�����+D�����Wa`ȂR)ŪFߚL!RJ>D��At̛�y�U0o�=BΈ1s/<D�0 p�g��p� 
C��)��9D�x�ᐫ>�$�4��x�{��8D��d�9'��H�=��a1�8D�p�ƆD�g
��hY�Vu���K;D���B�:0��z�I�8L�L5�9D��X�H�A�@h��υ+t�> �Qa5D�h��GS�(��7w�6�A�0D� {���,eФ1�C(хy�쐠��,D�X�F�/e����gMZ ���)D��������1@���u����h*D��K����;��ܑ�"��uS����-D��
%����h@B�9<��))Q�)D�$�"�J��
�IR &O|Y렄+D��j���=ol�SM�<EAtg*D����/��g� !q�� 7�Q�@�5D��!�h(N)(t��
�>#��Ѡ�O5D�� ����J@ܨ��%��$	`"O!�6��'V��yS��ʷ-�.��"O.ª�:��5��ԐX�bPQ"O��+�'�39�r4C�`S��0a�"Ol!Rd'N�y��d��N@�m�"Ot�Hd�]�*ޜ	�Ů*)�Uۄ"Ox���̧" P�F���I�C"O��@�r!xe�� R ;�Z�1�"O�E#��ݭ(�P�aFH�P�*�"O�Ժ�/��%�")�˕3>�� �"O@CC"���.���<%�"�*�"O~��H8+�����ٌ1k����"Op�����*V<��ӆ�lp欣�"O1�%��(Z{L�5Ywh��{�"O�q+�#2��y8�+��Y`i�F"O�dr���&�hEJ %����s"OX|;��3,�IFiK�v��E��"Ob\XB/X�p�X�*�'��CݮX�"O�eBTNP*v�(�Q�j*���"ODDj�fʭf��=82a�	���P"O��C_-c�FA�K�{��TX�"O>y#C�݅����	1� ��"O��"��/<p���hI��x�@"OjQ��
J?o��5Sm(/Z,�"O�i��6$��5z乓"O��X� �8"XۅI�lxe�"O�]�B̐P��E��bޓVL�k "O�є̐�i/|ܒP���L
�ly�"O
��֫ſe���Y�I�Y*�"O�=����Ψ��4/��:�U�@"O$#Ѕ;L��0�͖/f� �Y�"O��3߰D�d��So4�d��"O�]��ʇQѺ�b3d 3Sz�c"Ov�9c���!�� "v��> C �X�"O�qK�31����˂;5���"O����I(�ι���_#F(��p"O���g�#p7�< ��ñ7^��F"O8���Nl��J�(�g	��"O�,�"%�;����$U
�IP"OJx�����VA� 27�řfנ�7"O�9 c�٣ L��4&�
o��Ih�"On}���L�<��5ر��"q�Ơ�"O*�*s�TYb�9W웗zf�)a�"O���fLW�z<(��S-V�Ia"O�)0@�9� R���;UW,ؔ"O��ɒB�	1�T�v�E�VH����"O��I�*F	~Pcul��zF��"O���G	�p�" ��C;��s�"OtH�RF�C�.;7�B�Cz�؃"O�q�a���d!6��@�H�X-`z�"O��8cP.-T����I�L5��"O6mD�ΔS���uO �mb�Xq"O��BE�+C�Pc����ՉT"O�rf&�v���Ⲍ�'a���"On���I����*�BE�D�Lò"O�t@��)}�UQdc�ʤ"O����^!IЀ���-���"OBxy��?d(R�xѡVc�4xa""O�DX#Ů!�VPu �!R�b���"O p�@��L�=���?�:���"OT�B¯U��	0���qѠDQ�"O���k�s5�l� �U�2d\I�T"O��vצφh��A� v�"OVm�$D:&U��9�DY�3M�m9!"O� 6S�\�0t�5�%��q=,��g"O,�i��:�읣�R�'�2��"O�0��`�^��y!���Z���A"O$i��&W�!��$���RmZ���"O�ɘ���?�]p��:{�Ly!"Oʥbո�(u1G�>�i�"Op�"X387v)�������%"O|��Â�&G��X��V�i	�bw"O�t��L(X��P���!"O�])S�C<0Z�Ԣ���&B����"O��Q4�(��4�6.ƺb����"O�P��.��Z{P����k5.�+"O���6�9y���xfK@�~@���"O蹣t�ރT�6� ak^`0�"Ob,�B��1b|ɸ��ː6)�c�"O��y���1���	0%%�U��"O��g��4�S4*�$L�8(T"O�|;do��X�|IČm�ʔ
�"O�-��0D~�z6�_�`4�Y� "O.���i��w	D����T%�H3�"O8a#���
��Hi`�%-E���W"O�{�Eח`D�e*�D�%"6NMs�"O���T��?��ñ#,\2�ܛ�"O�$Zc�V|�����Ŕf&^)P�"Op�YaK���XP'�:K��"OH�J`Z9�nH�g� �U�Q"O���ɔkX ��G��3�B�"Op���#�)�.��g�e�>uG"O��$Ε�d0|!A�]� ��"O,ز6�-5�D� .��?lV�!�"O�����ĥ ��ࡡ�x�xY"O��ˑ.7X�G�����<�"OJe�J�/I��5��˖�n���� "O`����)h(dX`�Q�B�"�"O������F1��U�
�v\	h"O~�w�J�^;$(��4M"P�)"O��Ccg��`�5ۆb�X�
H�@"O�	:&��>J�<�!�\��̂E"O�4y��^(�0x٥�;ݺ1�"O\
&�GZ=C�%��)Ѕ�q"O d; �
D{iI�c�6ȓ#"O
����8c � ,��1a�!"O� hLKC-�`Q�K"��E"O&5��Qy�="R��K6ph�"O��iu�ŴKV�y+�M=a�H�"O��yW-�w%�a�5�ݤ��؆"O(���Lm�D\c��$�����"O<lsŮ�y�� Kޒd�0� �"O(�H��LAB��	w+;a}>���"O�,zB��Kݐ���9vNݰD"O��9��72]��Hj����"O�1P�F�]�@�� .����"O�q1E��?ؘ��瘤2�Z�ZB"O���W��Y���ޚW��uq"O&��U����磁L�+G"O��!s)�&g���l�.3��Z�"O�XZ5/[�3N:8���[9����"O85[����h;D!*	�8w^j���"O�� ʡv�H٠RA�#b����"O��P  U�C��=R���~5� �"Oܸ�e)Z������P,4H�z!"O���$�Y\բ`���` �eC�"O��(�J��h�bM�� 7	VY�"O�	2Ag��h�*�8�![�z��5zs"O� �q���g�p�wn�Q�.y3"O(0���<�<�C�F�2�s"O|�`D&��)K����w�\�zd"O~�80g9f��5�S��=��@"O�����@ߨM �g)%��q"OI��%�'u>�cg&�`��X��"O����()B��h�GB�o�ȕ��"O��N�p���$�f�P��"OB]��
Z���&��
T�:L�"O� �G��6t� ��KO���v"O���&9�"-���,'@&��c"O���1o��q�tn��P��J "O~5�B�T�W4��5n'V6�z"O8�"�[�T���L�3>�9�"O��I�̋*^IF$i!b�}��ذF"O )�u��#d<~M�M��"Q�R"O6�X$� q�6�a�K
�V�S�"O�]�tE���9��V1Ft��Cs"Ot�KK�)`� �dC,ZF��3q"Ol��V��t�H���Z�0�|11"O�����	%	4Mh�E*R20\0�"O��@�F�H�yK$Y�g&�Q�G"O�ie�Z�%�d$��P�fD�"O�l��FF��t
��ͺ��MЀ"O��� �N�Yj�#ب:
d�ؑ"O��k��p:dɢ�� %\>}��%1D����@(g܀Hps� 6i�n}
��-D���AEQ��p�P1�/@Y:Ç0D���T�X>Uxl�Y��:g�<��Ch$D�r��()lh���/(U6)���6D�|��-�}�1b�֛S8&{%�?D�4k�K�D�T$֍�!hA ��p�2D�\3�# �갸���7f��ܫ� /D���F��.k� �K�3� .!X!�!KX�)�Y)��2�c�l"!����R)j��́0$P��eDO5E!��%f<p�$j߳O�x�ڧŚ��!�N��d����B#�{T �S�!�䄱jO�(���S?z���G�Ǣq�!�$;�&�!��a:���F�t^!�D�0[���pG�ֆq#�e%M]�3!�d*Q�@u 2b2~(�q2d&ϵg����,||��_qaDz��R>RB�I�v+��Xč\��(�3�f�-:)�B�I�sʶᓵ��\��%pe�G"��B�3b@k�����=S$.��cl�B�	V�X���ԯJ6�Yir��zR$C�Xlp���#_@�+UdS�hZB䉤f����$�P�"� \���s6*B��@�t�Tc��<��#d
S�Jc(B�	�	n��I$!E�r�fp�S ]3�^C�IB�>AHΣq�P�
E�Y�C6�B�2,��i��F(pNdˑK#o��B�	Ts��{�jZ3�I k5-3\C��>�dID ��}�`���ό�� C�ɬ$�P�f.Q� ���!FʮLL.B���2E�gk^+Q��Y�ˤ;"B�I��ĩh"�8�Αq0O��2l*B�	m��8)�W�}��F۶n�C䉁Y�� ""��Q�TL��)�[�B�	�J]t�{� �:�\�@
,sU C��.�P�*�[�)q4��� 	��B� 4��`Ү	I��а0n,M��C�	�7�܊H $����(U��C�)� tY�`��jn0�y3G^%�Y��"O�S'�]�p�f�*p�"O����b�F< ���[-�L)��"O܈kt���7.F<p*(��L�!"O�-��')��M-!3���.Ƚ�yB�L���`(�#*�J 8#�_��yR�I�w~d��A�NҴ
��y������6AB�	�j���!�yB�R ڄͳBΓ�n�IR��G:�y2���6^0�c'ʇ�b=�PV舌�yr�@�? ��!�V��a���"�y����� ˾M�VH�s`�#�yb|(H��d�D��ҭC�yRHB�*��W)ٲ8$�e����y�jS;9\��FG�}�x��R�y�`O`�ۦ畀v�⃦��y�
���i���| r�jF5�y���V���*�`Q�vM&�P�L$�y2�G��|�E�;j)"�>�y2�͊/���鶥�4��Q��G��y�$۳f���zPF�9t�P���)O��yo!���e�� K#�yRE�EuN��珎<_Z�:��C��ybBU�u~���4�Ί.n����4�y�a��Q�'A�N�(5��Ļ�y�K��.��ј��D]�����y�HX�*�
�'� 4��;���y"�Q�21a��'��0�Tn���y��!cx����P�D1�sឳ�y�.E�6���O��F�Y��jP��y�LZ7	��X�!�$QΖ�w���y�dųN�xK�G�Nn$�V@���yRH�-Ur�ʑcW%M	B����K%�y¬��u�DY�s�?T�4bb ��yR�A�",D��nP��~��Q�0�y��ڪ	e��ђ��SPa
1�	8�y򋑝|6l�p��׬rq�졀ň�y2�8oV��6*�5n�ĩi�H�y�����`r�ޅg�:!O͛�y��с
�°����ZK�0 0&ݛ�y�UB$��Z?|�������y�ϔ���ݑ�c��Aj.�;���<�yR��]�H�@�B��3���GL���y�&�X� �y�Z7W��� ׊ߑ�y���+|#�C��WB�k'�yBCݧ$ ��&K����IZ1�yZ�0���?T��Y���?:���'s<h��D�����go�=��9��'��9��͔h��8��'�eU�Z�'BH�s�4�C�dܑF�V�'sZP���:��T1#c�o���'�T��1a�?��}h�k�"���'�V`R׊E�$�Ł0&�p�� C
�'fVY��DU�1��ܺ�l�a�N�

�'�}dL:T���qG�K|�aI�'�h�u��49�L��%��&E਀�':ഹ� ^�z�sb�����'<RЊ�"�_�Z�P��$
�R��'�
x�ϝ�D_]y!F�Se�a��'9���@71#8]�� ޛN����' i8�I@9QO��K���ZuP
�'J�A�/�(3��y$���V-
�'�x�ÇZ�<��y��=Ӿ�	�'�2@@�oRc"TACHOQ�B
��� Ё��>Ԃ{c�}�b�9�"O�` ��
�6���S�P|��"O�(C怿EJ�����|�b!C"O(�KG��#j-\4���Q�%�1� "O����N
�9T�Q��2����"O�� �JɥJ<BԻ%'=y����t"O�z��l8	ֿyX��R3I9�!��I�:�)F��M$BmW�a�!��<.e��!6+�91�V0r���:p!���"p4��A&Ɍ\�P�q���H!�Q�~�1A.�.���
�f:.�!��c��@R��<@�>��ڻR�!�dE�`$��NYG}�h�R���!���h�&�QpJJ�Y�LΥ!�!�$��	����`C�T��\��J�m�!�6C��q6��z��Q��W�!���5����LM�'_����F
�!�!�d܉a�@-
7�
=QT���?|�!�$�<T�1BQ`�3c��d+ĞW�!�dԷ?N�XpM$bYթ��+����3f,�Q��0'	�Y�'��y�&�?G> K�@�'"��0�
�*�y��ef�<C򋌏V�C�e�y�k��ylXt Λ�~Z��T���y���xgeX���'�ԳvL�/�y"��&)^���!���6�:f�\��y"��������f �𩘁�y��N+,tp�z�jM�8�"E�g@G�y�E"~��"�>)}2� ��7�yr�U��ڐ`�#.xf�"�mʝ�yR�A�LH�d�;)b�8樍�y���<�s���?-���B`�K�y��� !^���%�O���M[<�y���/MI��o��:��5  ��y��8��(yQ�R�HyB���J��yB�݉NF>tk
�9�������:�yr[�E%<D���[����ԅ�y�k�p�;E�4Vo.���N�9�yrOO&fA��s��!H0���Y&�y�1Ut�Ƴ;PހЄ�0�y��ܜ:��xB�ǁ-���W� )�y���"ܒp�©$Y��G�.�y�,�)nWP���*���d8w��	�y� �1k���� .�
� Y�C�0�y��u������ ���Ce���y">J��-�
��th+��T&H�ȓ0��u:Q�L�%��1�ַ	
�ԆȓbU\ #�
�Z�l���<#�	�ȓ�Ha aL�blt����6MP�}�ȓN���@�e��(Z1���2sf`��&^�� G��xj`	��Ey����p�>�	U���%r�B����$��gv,! �^��-�-��m<��ȓH��B'�7O�ɂ��11���ȓ;�Ta��"PoԸ5�"��*B���ȓm�J����5(Ȑ=x���CJ�l�ȓKP �# ��i(�H�3Ⰶ�<t�Y�ő1��� �*^=Ԇ�f�ȭ���U�k<L�D!��{(L��D�x���į8���AfO N�ȓ+���Pm
 N�Qp�Լg !��m͚�T�׶= TԘ#C����l��ty֧�}�2�#��"xrA����o��I�h�Ă֝F�����l<D�� �a� ���6@�d
Tg~_�D�&"Of� `D�	�]y� �B�E�"O< 0�l�is(M���!?ja"O�tÉޭ0���� �/��R�"O��"�)��PU�g)��E�t��"O�P����X���gƓȖ�bf"O���4b׺j�ze����(�b�"O�	(֡܇���2�4?�,탔"O�i��OJ
EW��s�(D�+��uyt"O�����I���#�!�k�T��`"OD%`���%q:�ur`'	5���k�"O�Qx�E�Y��@!4�{ߜ�+"O"�JF���%e9T�l�3��?�y��D�!
����t�XZc�Ŗ�y�����V�)�g�l)Н�����y�$�]�:�ge��5ȑ�@�yn ���qC�G�X�2�9a�#�y�L���x���ؤQ��ܳ��M�yBI,~��T���d(�y���L,I�V-X&z*�X!I��y��� ܤQ@��_��Ű�e^�y���>n��hyB�z�tqP�盖�y�*J%Z0���c� ��G�ٍ�yR,�bU��8�C���1��M�y�F?LRDB'��Ͱ=Qܐ�y��6e�>Xx�iZ����6#+!�� �e��� �'i��dB��7�!�Ę	N����D��5�f݂D"OZ\#`�+4�t\R"'@�^%$�QV"O���vl�����ҋ"��A��"O��H���j��|�j�5�F-"�"O*eR�i�1>4)3��I�h0�G"OB�+'�HNo�TJՀ#���"*O�%І��HaLjH�<e(��x�'��0�۹k�
=J��ڔFg���'�XH��Ѱ]W�#i��9R*���'˜Q1�▟�n�x�Ã �`�@�':vL�7DҔm/z�1��K�M��
�'T){�� 9����񠚚rG���
�'{�5��̌\�Ȑф�[�fT��'9$�H	�"m��I9���@a|���'�r�#$��t�,���L5�J ��'-�,���N�h0�(Фy�@���'���薬��|�䙠���r�1�'�� ꁧ�����du��s�'�x�k�E�&�,�`R�b��P�'W����'@� ���"TEr�{�'#��d&�� �C�p���'P�B���&y�
� �������'���ƃLudt�j�j�rP��'�� X���	]Vx��B�0-]
x�'�Ź�I�7Z�X&KD�V�����'�D�h���H�F�z�-�#P�x͒�'����j�v�0]ZT��O9zp��'F$��e�#X��)B�/
�v��X�
�'��h������Ԁpm�g%N1�
�'$��{ N��U�B.�X1�9a
�'}��3�hHF��� ��T(U?�s	�'#<�Q���p�"��$dL�A���'px(a�V�ln8,K�@·+�L�	�'�.�{�B�A��YƄ��mh�d�	�'�ح#Gd9@-��s�蝨_�N�	�'�@�s����e*AJ�e��^(��)�'�&d� �/f�$ɥB�:N$��)��� ��z��މb�\�2d�>��!�U"O�����ޱ_䔅ɰ�<�9r"O�a[�A�IH�17#j��"O$��`C�R���S��	$\	�u�"O&�8�Jʿ99���[i:���m�!�D��e��\�W�?XƲL�D+G<(�!�t�$��u��;=U"��ӫ_�!�!�B,%@���g ۉp�B��W$�-N�!�DϢ�b���������#�	�!���A��PIB���B��5�W[a!�d�g�"i�fH�N@B0���5D9!�D˪ ������+��!��$�"���I� ��Iu�̉s�!�$�/6��:�-Ǫ6뢌��I# �!��V�2�0�ܽ��� \i����>b�,J��JMr�g��p���ȓ�F��%��Z^l跠R���X��K�z���	<�� ���OW��c�����ŉ<�L(ÖK�7 �h�ȓY#�ذRd�^fr�j�dɥ2���ȓB����-O	A���n� h����ȓJ=�t�OY�[��*�k�=�Մ�BsKʿ0y�!����,�� �%?D��+g�U&>�Qy��J�;l�Pԋ:D�0ar��oS��C�K�)ax�(�6D�<��N��?�Hqs���;q~l��6D�a��LBj�ݣT��sp��e�3D��C&⌳=�L|�SC;|.���0D�X��� <1��#�ī+	�h�ǩ3D���7.�'D:��d���h�Р<D���En�$6�$ڲ�8&��T3h9D��c�ꓲU.�(�q��'cBEk�	$D��;B�b���㒈�=(���C#D���p�M�
�$)��͌T�e�+,D��&�Sh�y�sH�
P��rJ/D��Iǎ���9��&��7�iPI-D����̖`�  Zv,D�DOf�t?D��G�V��8��-(r6 �=D����^-��*���
��h`#h:D�P�T��lJvm��\P��YBI;D�\�"̌�/2t�`��dX>�Z�.:D�d�� �J�<��bG��io2�+6o6D�4#�dO.jP���)F��St�4D��s�Z�ZC �r�鞝u�`��10D��d��
b��d@3n�w$𳢇-D�T�R��	r��ń�d18����?D����ʮe��ʃ^8��m<D��ɰn�"Fm��D=�6ъS/-D�� �� $$�\��.�/X�*�ِN,D��"Qi�&L� a�	A�4�	Ȧ�*D��Ȗ����LI2�Y�#�$D�X��nϴ=���SWꊻM`>�� !D��q�S�PBQ	���w��� D��r1Kξ�$8ٴ�?^g��82�+D�(ᕀ�w�P��@ E�:��4�(D�(���8-1b%[�9�
���d,D���!A�(x�ł�
@p�?D�h��Q5R�f���a�@o<D�L��e�/xk��	���#=�"�hb�8D� ��D�0.�J�3�<je� !�#8D� �d��r�>�ӕK�������7D�<
�	�e�D b�`�,��5�*D�d�kщ0�s�Ȉ",�}�R�-D�4#!�����Ē|�x�@��>D�� ���G�M7���C ]4z��Y[�"O��3$Ȁ<�"���f� ]��"O�!�"B�M}�L{U�B�h��T��"O�B�O�8R�l��̂�||��"O~q�p�S7:
]���șy��)�"O���q�H�8!(�����xd��[�"OP�ㄪho�����&a^��r"O������
�������&.Snq �"O��b�L4V�RC!S5JNUi�"O:L�;�UZ7�ǩp�[�"O0ijA#�.9��XP.ϩR����A"O\qkрR�I�P��m�H��/�M�<�SH֠8_�q��+�~P ��a�`�<��?c湲�L�]�9��YV�<	�ѽZF0�`���m�,�C� w�<a���_�N�B���V.Ƹj�/�N�<������H0vt�I�&HJ�<��F�a�J����N�Y7����^�<1�G��N 
d��{�P�	s��S�<��k̻���ւ)��X�e�LO�<����X�Ĕc+��i�Z�NB�	�f֭��-&E<�2�Q�csDB�"�(��	�&`vA��j��B䉊mඬҷ�ݹL�j�7��6$C�	������Ā}/I#_��B�I%!����¤[�z�Q7G-S�B�I��4��S"����Z��*��B�W����Ǜ�JM��^�eU�B�GHDȓ�Iܰ@Pν���$QږB䉽z�~�	��̑9��SuY�C�B�I�}�"xzP:j��0�3�
!�vB�	�z"�`���ɤ*DÐ�R,��C�2Y��Z�B�6_�Xs@@�%B����O�{�fM�#�˟�@Y��.W>t1!�������R&�ƬY�Áy0!�D@+"mEZu�Bhj5Q�,�X!�$٬}g"�"N~�![��v!�D�2��\#w�LT������+b!�Ą4>���e�(x����+��PM!�Jg���Sb�Z�*����K9�!��	�<g<���!���;��&3�!�V
$���s�[ t���c�!�$��h��(�蝱D۾��mQ�X!�D��C�2�H�d��.�y��#8<!�$ ��졕 �>��8�dN�x�!�7Yv4q�����9�R I�P��!�O4bz8<y�/�;�LL�@�K+T�!�Ę	&e&a�g�S�WO����b"w2!�$R�u�2��cNӚX#(�с�X�fJ!��B����7F��֝��@6�!�dҤu��0�ؕ0H���]�!�D��4��#g��8Z�Iv�#�!�d�a|v��s �
]n|���7)�!�:�@�:�nN�|U؉��F��w�!�$�.y�A#�f;FEx9[�KK�#�!�$�"8s4 ���)��}�Ʉ@�!��G]���Q�Z���v��<�!�$ш3lQba�B�1嫜?X�!�d�?#�����N6���3ʋW�!�A�*E�ѭ�%"#t�!��'93!��L��m�BJ�9st$E��I�T!���\z�4�刕�
��%h��?�!�$W>]��Xs��6�~�Kf �sg!��9R�Q�2�]����! ��!�� 2I7%G,tc&��O�^Xw"O��ҭ�e#�C�&�N��ӧ"O�$
�H�z!��ȱ�	�T�2�"O�Q���1D�S���
c$��%"O T˱i�D�x����Lr�=��"O�ȉ5�S0:$ţ`����i��"O����O�x�銐8R �"OV�yU%V�&��0M P	☓d"O�H�f�
�Z`��2ThdĂQ"O�A�����H@��N�7`Z��3"O��*!n_"P\|:�B�)r`r���"O(���D�*%��pb�ͶXV��"O,��V,.���H���/���+�P�<��S� �T�0櫍�K`<����N�<C��R������F�XP��N�<q%A�[ ��fI��H$��s�<��,R�1hq�qeŝ.�5�Ӎ�J�<Q���9I�Ԭ����>@��
�^�<A�K����К��9���F�[�<`#R��4Bv��^ 䳃�Y�<��dT&3?�Q�BhVi�> �D�o�<y0�Җ>�Лa.�._ډ`��i�<� ɝ�>�
=��}��Ȇ)�_�<ϳIzz�R ��w��h�7ϟc�<��>�L-�fD�0]ɠ����^�<y�g�s6ht�����lƌ���NVW�<�ucУR���aD��Y_���R��x�<ir��5g� h�U�WV��(���s�<QsP0Y"Dٲ�c��x��1�w��D�<Q�+��|�
��͊�(�d�iZZ�<�	3v�I��]���CC�R�<���
*/��� �V�_nډ[�F�v�<��i�>r ���!`�sq�y��n�<�@�R"�ٗ��\/�݉#�i�<) ����DB��ɋ?I��Y1��}�<���g�~И��zl0���
o�<�բ�6f����
O�0]X�K!cLn�<��u�t��cۑ*�P%K@�<�ׂ�t���A�BK�H�X�e�V�<aE.Q�n[���ώ����xg�U�<Y@b�5(��`A�I����h�ʞP�<A�lķ$�����l~x��p��Wa�<q�ƾ=�h�ZWÔ>�|��M�_�<A�ȑ�bh�m�E`D��$��^�<���̇{��H��Dń2�����E]�<��� [�D�b K��ytܘ�Tk�[�<��OL�%aba���P�������B��;�ڕ��f�=��Y�pc��B�	P��BSH���¹!#k�)36�B�Y7��e@6����C�n�dC䉐A�V!`�"ڶ�x=a���,\�bC�+������m'Z)*�&Y�~�,C��1ZHBa#6t2i4�Q? bC�	�j��x$��l��O�.nC�I/Hf	2@eA*%��;`$�!vTC�P	��+��1,���m��&��B�I?E@��:�,@#0�����ϖC�	�}�)9��ǥW�xA �I֢\�xC�ɴ
s�4�0�ۂ'�F��O@�U�vC�l:�j�싿�ک�RoH�/k�B�	�_��R��֞h��d�`�PR�B�	?|�P=X���*:�i�`a�'p�C�Iy.~�s%m�7A��Eҵ��\��C�I�a-R-X"���v���C~vC�)� ��s��R5�M����4	is"O����E���5!!�7>dAA"O�pK2�H?4�ޝ�%��-g�HH%"O���A�]�hp��!���d"O�Ը�cͧ
�RU"֍72Y�w"Onp�S+�5�� ��Y�P,�!��"O�Ě�`��l���+�6�i�"O��9�ׁb�ƌY3��Ꚍ�&"O (!Sb�A�F�p�cR�ް�%"O� w�K�
�]�E��(�`A"O�0��,K(L=�ᱣ_�O���"O\D�Bȏ=Z�@=�u�A �.d�"O`�Ye� �;Zq�Wˑ� ��h@f"O���i�6w$|�bj]�)�`'"Oб��N�-7���5�����%�"O9�C+��jM>�P˔�H�2��"ORY�@k-F�Ah��V��{7"ORء�hA��*��מ'sNhf"O�Ĺ"K�U'fÇ��Aa���T"Ob�*�I؃]���v��4z*q�"O��t�׮�^�!``^S�Ą�&"O��҅.I�\�]�a��W�h��"O�h� �N�]Z�M��Đ��e�"O� M16h(9Q����� [�"O�p�_�15f��֭T�V׆�e"O��4DH)tt3l�T�`�A"On��bGJ��ӷ�Q�t�N�I�"O�ؑ��v�Qp���]f�0�"O�p-t}�$�+qu��T/�8HL!�?ֈ�)�㉋U�,�b$_!���/���UG��T���$$!�6	�t��u ��A�
�ʦ�	?Z!��ES���F�z&�Ͱ�� !򄐿"���i��|�
ӆ���!�SiB�Q��+f�@��C�\�!�ބ2�`1mP���qr㐄�!�DٴBԢ�JOK�d��Ѣ�5�Pyҥո9�QrGȞN�� @���y�ίn���s�mF.v���!l6�y2�5XZ��H�o`�m��EL��yRa�7�	�R�	t�Q)#O��y���,�m��Ҟdx8�t�@8�yb�{�^a�V�גtQl��R�T��y�E�zM�;գ�k:������yBȂ�-��Pصj�"o�Б��(ǔ�y���֑+`��ֈ���mH$O:C�	4��qp��sf-��)��XC�	Q0u3e�	Cl
6D�0#XC�ɕV(�sB�;X�P��W �.UtC�I'{�h!�OT�F�DX1�J]<As�C䉼6��p�F	R=�ly�b(Y��C�	\Ǝ�1�W�2��0�è�9�*B�	
�ȘV-^'x,���蛅{ofB��/n�(�sK�^�z�C����8`B�I�]�x�ҰIS
b�X���*�H^
B��$f|�92�C�+�R狝�MB�ɰS�Z�sƚ� �3g�� �C䉔h$���L�b��� ����XɪC�I/7�܂�f��B��!�ŲBǈC�Ip�8��� ,��-{fC��|C�	Lr�0� ..Pd�P@� �#�fC�	�T�D�S�KG�|�B�2 ��9A��C䉾+o�ĸ���	,�����'"C�� d�Z����qsءto�Li�B�)� ����ͯ
�J��z�r���"O(�Ve�#nL���$�z��8`"O���k��V�&��̩���9$"O�0p掔���� ��gHn���"O�0I��:V��Y���,V>eK""O������`��@��
IE(�1�"O
L�b�/b � � ϗ�3%tlXr"O��xu���#Q��)Ch�!M!��"�"O��� ���5z�H�����S�"O��aB�`�Y@���k�ܰ�r"Oz�s�o�*��䨥�y��y�"O�*_#̈�1e�V��9�0"O���N�!\�=�"%��a�T"O
�[ǊJ� ��h3���!()h"O@25�r��X�C�2h�(�"O�4Sp��<{������z0IA"O��Pî���ęҏ؀n&��i�"O�xk�FE��pQ��O�$n���"O|�9�H�&P9Z(�q(�*W^�5ce"OxҴ#�49�+d�2KxT�Y"O@��B$M�~4|�!RAL�'sĈ!�"O�U��I'�dms�Fr�9��"O�h.\�E�BZ�ڔQ���)(�!�\�I�p�z�n� Y����Jtx!�䝬� ,��膧c�<#��	H!�ċ""`��	+�9*�,ǯu!���-	LX`t *L���t�G�L�!�G�x�H��#�8y�D���)�,|9!�$ݲ$�(�!P�_�Y �LQ��\�!��ݚ\f̻�$P3i���Z���n�!�DR	�A����1�5�a�D��PyJ�/�mS��ƣ�<e��Ҽ�y��r���@�O��&��&��y�� ��,%+�/
�� C��y�A��7{t��*W�^=��KD��y���@�"�G��P��T�y�G="E����N�WnF��D#I��y��w��؆���T?�TKS � �y蝝X�Ի�lL���br�\$�yb�I� � mk��ԠL���Bb_��y�d ���@YF�OJΈ��G�?�yb��EAp5��ӭBWR�')���yb�S*[�*������?c��Ƅ	8�y�A�H���D(��C�P��	���y�HV�\'P��E7;Fh�"���y�$\ �@�I |E�Ր�H��y�!�	d��H����1v1�`s�"*�y2&P��	�#`V7Q~9:�
I��yr�N&*��qh���*/�<���C��y�E�x^d�R�*�2+.�P
>�y�,٠<,��2>.����[��y�fN6Wj���B�D�4�V&��Py�j�9Z	�]�AO�r�vuːiRc�<�U^��|t�F�ЖuG.��Gt�<Q�cYw��rQ!ڪg�6qAs�<Q�"J��28��JQ�@��whLo�<A`E�W�HE[��"ݤ�"���l�<1���1c~�g͝"dԾ8�`JN@�<G-�ib�E����I�4��R}�<�U�4�J����=�� ��r�<)Ջ�	� B�S�O"��I�f�j�<����d��8�d�:6IJ�)�hh�<G�ßGopT��R�+?���z�<���U´Y;p^����0db�<� �����3r���¤�U���"O��x��B�q���p"CD=79�"Or<(��C0UV��r��!�0��"O&�����m���)�f��M�"OH�L,OS$MYL,@�(`ӆ"O�� )��j�HYwoF����"O� *�	ղ/�%�b�Ǽ(���"O�9�Ј�5R	��֥
5[f�!�"O�����͊:RBK�Oe��S�"O�(S0-Ą#����K�1�"O|�$�Я�U肇�;sG���@"OF���	�G�|�bF��Y3��"O�ݓt���N�d��TI<K0,��F"O�$���*F��u�(�2l ��"O��R��jf<�@��P�*���P"Op��4q���e� �p1�"OjѺ���6A�T��B���F�r�z�"O~hS�*}�k�+L�>Qr"Oz�#I�Rw>��5k��q�0��!"O�����cB��t�۠ �؜�e"OȜH�+۬I�h1��Z�̬�A"O�!YU�śHx*�i�L� Ty"O���r��w�(�R��$�t��D"OV��� y�&u������Pz�"O�mH�H�`$���J�E<,K "O�q��`K�5�^Jé\�&b�b#"O���! ��Ud��QbD"Zj��%"O����]�A��yQ�둋"^�6"O��bàI�E��8��	�7ZF��"Ot���c��\zW�Q�W� ;C"O�ĸ��9x6F9zC�����f"O�;��@���S�e���p"�"O֐X�'Rʸ\
��±�c"O4�K3�#}��c�ĿV��"O��Yn</|h=x�f�$P��Ac"O|��B�U��zJ�fCDf��R"O�h���1	h�0*��%�r]0'"O���&e�K�Z$%�:�e�3"O"q�Ԏ740 �r���I�-��"OdIc�-H�fS���6�е=�i��"O�@�̓
Gn����ɻ.�*���"O�p�a*K/f�.�3W����L�`"O."�H�;��i��lT=0*�"Oz�It%Q��ҥɃ"c.�K�"ODL��o�8,M0��	qְ��"Op9(]��h��<�6���"O4�B�Ä�}��3�N��r�P(��"O�!@r�Љ~s���χ�x \��V"O:�3���;�1� �	�e�2"O�+���-O�U�+�0� ��0"O$�(�D����+E�!�Z��s"O�9��{B��*Uɀ��"O�J&�h�a:@�6��""OtE��E+$��U�w�/o�H�"OD����5�2PB���@\��0"O��0F�;��Ԣۭx��=9 ��d�<AW �~I�u��-C"0��S�Z�<���!(�޸2��C'91���`�X�<Ɂ�ӧ= ����o��� OB\�<�􈑲aB�(��B�F�&Nt��	ux ���%o���;��յx@*���b���l�n���{q)��;)��l@�; %�>"�z���-�r�X����
TS�iN�Z����Ȓ j� ��S�? H��� G�..��CDV�/�B"O��RwH�.y���W���:�p(&"O�H�� ;:d��kW�[����"O�8R��>w����
V� �)$"O@xL�	l��Q��F��-��"O�ء���-G�D`@�au&)��"O�������w�Q�F#�cDؠ�"OZT��̓_<8=ڥ�]D���26�'zp%�"Bh-�)P �,5����!Q�I�	�'��ZQ)Ag��Y��kAT6�\
	�'#���#�� \�x��I�R�Y"�'���@��Wvv)J�)ː[#�1��'��9�A¯������T]՞-��'P]��Ô'cZ*!X_�K�z1c�'W� �޸-tP�P�j�3��0�'jR!��G)S�z�r�$�����'�r`�* &78<aƪ&q��Ai�'sJd1�EClꅎ���Y�'+�t��)�?8O55��W3N�
�'�6��hW��\��Ԅ��L=��K
�'sh(8gJ��j��vΝD�P�	�'m\M��l�0�@���W� �)�'��h����\fxPG�RT�h�'V,a��J�M� 
S!+f���'���#r��H��iD���a�V<��'�X-��e��R�erD�V�U�&���',t�(��U3���a�W[8u�	�'U������P'p�� ���H-�%��'�� ��f�xQ�ç������'E���p�:Q�����/1�t��'$$9I%���'K��AD�Ѭ8h
�'V� �tF�*K܆�����)#DEMR���!3��L�:w�A��L�o�}�<d��c($�r���#[��(:h��ƙC�/�h�,�%	O��0?��hR6/��:v��b�t��gbFQ8���cHXC�5�N�<!5aL�t��g�σ2[���Z�<YE�[2�(�f$M7\F�����V~��H�m���a�/��"�2�I�gM��U��|:�
0HU�<�����M؊���"T~���x��Y(K��q���x�`��KN�3⊡&?����K�<"
D�qb�eN���D<�O����K�<6��!���2D�L\ 	��V�x�;�h� }�r5[��'r�p�DLM�0��c���l#�tQ��d՜,�2c#�����[�-_�I=E 4t�t&P�D�� �։m�!�D�7O��4
�`>'�a#$I3B��I��D�\�סj��1ֈm��>��yZ�1��۔���&H4�C�I�ʞ�h3�M��ɇ�S+m�d��1��5"��
ڑ�(��V��?����L%YYA�'�/�n! ����6Ma|Rk�~K��QFR-(�4�0W��hl
=�*Qt,M���t~8��&Ps8���l[����>ۊyc�f �	�n(�X���O9�	�7��0{;�	�~�����X�(t��!?]+��ڒ"OV	b$Å-n��T�g�Zm-�EH� աE:H��6��'{ݺ!�&�� Zr��	a��p�O��5>�U'��u��P��!D���n_�`����W3h��i8r�ޚE��.�遇�E�n��]P�E���:�	?/�^Lbq�ݜ\�,�s�ǳ`���^{��� F���yQ�����$���w�܋3Y�4�O�y�N�#"	Hs����� T����т;;��B1�X�~6qOb�8�Y����&/�K��I�eW�����,��u#��B8�1p�n�1�ȓX1M�J�^�D5�tn�9$(�X����n�*q�%�� O�إ+"��[5
c?�h31�Lầ#�7G�$��>�,�"O�m���߀
Dd#Ԏ�<��]����>��9��$ �E�f��H �e��.��(O�cQ���4�Z1�� ˺Q���'�4B���1i[�1D/&g�Ĉ��-[@�6�YP˕�m�pev�͛lӠ	04-#�O����*-�ɒU�]&&�����dEN���0�0;V.��r��Cn�EL���'uРm3�@T?;IL�	W��0S��]��S�? &��ԡ>D$���9
���(→#dV)��ēU�X��0�J#n.���#ڼK�����Xv��C�v��eU�<ك�V6f: �aMG-l�Z�>nfaCCQ=e��(t�*fW�ٓ��e2��@���:<�D�V�B�6^<#��(\O�Y�pC��h��˥"�1P�"27j�ʠ�2 5�m�Fb�.�1kC�'��z�瓥0��_l�t���}2g�'�(e�C
�L��Th(�~r��'F�2���� +w�,���M���x��LT��(�e �d���$iI#WC�u����aX
HxvNJ�N��<b%��g��~⤉�)aЕ㕬¼o�R��Ǐ�yBƟ c#��$�_(Z{ڈ`0DV�yBȡIV���M�0=��@�	ZV��KR�+q�mr�APJ8�p�I@+:-d"K�Rp�IR�E0��5p�H�*{!�\�
�Q%�"M�����e �r!�D�>rD(���"-2A�c�!�d���	s�aѴ�v�OH.r�!򤁗H��b�-ڞrJpJ���!��8T�-3�H�\&l��-��&�!�D��qʴL��`;���r�ġh�!�dZ�<�Rd�w'� }Ӵ��a*Z�!򄉺}�P�&�l�Z$�B�ɔ�!�@(E � V-Y�2�X��b��Z�!��ڈq�H��WZ�2�h���{y!��g5"�& �l�Z���AN�mJ!�d��(��������A�z4!�W��t�;5)�7y��$�!�$�<�X`�#���b��:!�$�x*�q"��63�R���(	!�d�*E��3��6���K�g�T�!��^�C+���6jJR�rD ��{I!�$��A����=t� pCG_!��t E�r��6{@H4ǜ7�!��
Lj,9
��)N��@
a�!�DH���1`T:m'40H�f�D�!�d��m���wn���BяK�:O!�D�dc�Aw/��O������Ɩ"'!�U-��mW�0���2���n !�Ě�_�>e���H�7�����!��[�!�d�2��`Tn�,תd�s�U'X3!��ؽ?�ؙ8�B�\�bt��$:!��K�"
�X�V�mu"FL�b!�)r��2�ȅ{��s��z�!��H����H��_�������~�!�D�3z�  ��d{�(��M� �!�Ē�(�B����Wi��;��C2~�!���[�*j��I+6K�<Iq.^9A�!�D��zI�Hj�f��|N� ��O���!�$P4��P���B̖���MP�2�!�D�=�:9ш�,]�N��`�;Z�!�D]8p�ށqQ-��9�\�aug��!�$Z� �(�#"#�	�ћ�&�-`!�+s��y(�-�(��
v#R�l\!�D� kXTظT���-���q��'V!�$�!f/�MKqA@�w�is�ʾF!�䂗tޠ�zW �l@�1g�:n!�D ?���K���B��X�	7!�U&�������&�(L�tG	w&!���(T"8gi��l�C�ɋV<!�D�"f%�E�v��&͐�� I�J!�d^�x��1H�%-G�I��VS!��.v|�\�UCڝJK���� �zc!���[F~ �"�����Q��ϛ R!��D�\z�����H:r���� �R#QN!�ȅh��iAA �3d|��#�,	V�!�dՋ���Kpe��Lx���d�<G�!�� �,;�Hgм���*�U��"O�:��������K٢B�a�"O��Pa�)@���*Di̜)���ل"O.�8��(�0��7u�rej2"O��	S�00F���Sَʹ��"O ��e��G���*[δ )�"O�AkH;e�C�	�U�|�0�"OB�.ܢ}��#P�K����"O&@���Q!O����EL�v���w�'��$�YpX�hJp&
�E��/�z�jZ5�2\O���1Ş*[�RE��'�0�B� G��1�D�:޸�Q�'�]Ҕ��(}��j�ū(Q��CJ>a�+)U��c��%L�^"}RትOlF�A�+J��$A(��Ue�<��LI#xj��	!��T8V��#,ɞ �W!�1JS���b�P,�~&���ao.|r%�f�E���=��G.$���d��t"P��A)_�rP�7f�<be{G╛��A�q@GE��(�ŦR��������![:�]z�-O:�g�?`�|��	��4�d���*��S�60�aɛ�P&D��V�yR���,vlAg�Q�P�5	�n��I#U�S��\$?
x��e�,�>p�	# ��}�oFwǲu9�$"D��)��ܺ���+G2d���pw�'�ޅ�am]��v$S�+ُt�,b>!'��"v�I2<@�Тrb��H#��:6AݵH��5����0�H#4�$�E�Į�1~��i���@7���ɊL@�BL^�G�ج�bCު)�����`���v��Na��'"�q���U(�˖�G�*�
��G�04�L���C-9��QT��
^�iC�=?��(΂y �h3fI�? Q�u�^���O=� ��	 $���k'%�0�A��'�^����D4�dX3)F=y��a�H�	&l�4�N4�dĻkO���O��'.Q)-Q&� �qf��=w1d�k�'(AVk�Zd��)"�O�c t(����86������ɟ$��yf��y�o	2�(���_D�9
�!���0<��&�v�(�r"���	xdy�g愋h�<��n�;��@����VҪd��'���]q�Hg�ظ� J��a�nT0r\���4b�|������,b�O
��Es�߫FYzB�I�cY,�#�C9>*BXv	8e�`5ze��;6���TeU��{�6�3�䈑'b��6X��8�!�L!��I�*����E!+���$*,��Aٺ^z�B�s����D^)/2���A�|�f����ay�OC� �@�h��_�v/T�;�E��^6$�В#¼�p�@OP%F`B�	�|1��E��vk.��*�KV.�O,��J�IR&��'#^ �H�4�%�A.V��r⟴�N���"O|��G�45��1�� >ArT�����]{�DCs�>�Co �gyEʑ�l��ʎ�q̜y�V*D�y�'m����K�jC� �E��?�F���&����+B�0���6�P5����o�!���uV��� �\T�� �&a�!�D�L�ҡ�uU��3�o�B�!�䐒)�`�ӄ�Ì6H}YсK!��u��)3.'a#����!�!��f��uS"��|`�X&�L�!򤓸,��� $9}����0�>E�!���>C�p�Pr�>d�<����a�!�Y�ڕ�E�D�`��mJ���C�!�	Q�H�IA��
� ���U�!�dļ`�0HFH�d�ؕ��	�!�d@�H$��G�ڟ��}�W�Y!��̓}���s�v�B�P�8X!��=�4��'������w'Z-#M!�!�V��U�׎ ����F\4V�!�WRJn c�gY+Z��Q���t!�$�'HP�GUZ��獓Ge!�����q*��U"W����F��-o!�E*khN��@ �P1s���>�!�d�8<F���#SҊ����.�!�� b�����\8x�у�H��p�"O���qj�W�x�3B
���"O^�S6�[0�&���� n��t"O6D��n�:	V.�:p�cS 1�r"Od<� ��?g� p6��DqQ"O���CˬP
�z4�K�}5p��R"O�a���C�U: `a16�W"O�A���Q�3z�h�Eg�G?zI�b"O�a9���;'I<]�ch� a�yn!�� ��`����:v(����:}E!�DC�v�Jт �r��i��K!�d�a����!GH78q��$@	M!�2��� 	&�x��!]�6؇ȓ<q̰�"BW�]`��4c_T��I��6ATP�b-^V�ir���yu.���Uİ%��/s{�i�r*��l�ȓa@h8�*opp�$DOYFB]�ȓ3h��'�N�ԐA�b���1İ���0n��b��++hfS'���z����"��5��+Ng���d�:;�"��� f� �D��ja�ʆō�T�"��xޘ���H�m�r�V��C~����2i���F�˚U4�	f�d�i�ȓ1�4�pa�ƣT�8����u��~@h`k�\�A���1�\:	��2 jxgΕ6�w(�N����b6(�{��Xx��0a K�oDDQ�ȓ0>r�q֎�|�H���~ߤ��ȓ3�@�r���AZlݩ�\�{Xa�ȓT�n`�Uđ��*ـ& �-��e�ȓG0`��3ı������bJ4���O^���fǘq����0��.�~|��O�#r���)+nT�)]X\��NO���p�N���P�7Y�H��ȓ+5H���W::|$p���ѷd�$��ȓ&���)/V)��f��5K�{2,(��5I���O4*E�Ywa<ݸ�e�<c���B�ON]2E�X�	b4ч���L
��abڀR���� A�S�� �v����dRH	W������ O L�É�!"Vq[g_���%ЛZ�f�bEI��gN��q�?D��R��S7Q���ʒ�	�u�Zl�@a<?ѥ�M�e�N��pA�9T��?	X�]�p�6���EI�#wR,�0$/D�U
M�<Eʥ�F�ya|)�QׂT�ܔ�C4Oh<�w&� b��qO&i3
�,��"��3:�h�E�'E }3�,G�G���@��4f ��a!�8f�!�(��@k��&�N�/��[R���&ɴ=D{�G�H����rk�)��"UfI3��Ĩ�+>���C��H#nRnD��N��y�*��}����E�n����'���MÂO�t�P�P-��Q��[�#U?�h�k��Vg�`�d8���Pt	��\�!�$_���8F�)R��q`��:z���9�Yc��%%���ۗܟrGy���,±̀&����/�0>yDؑ�rŲp.��"�MA�"��U�>������D./�q)E�V�:���8��D�#��F�a�ؼW��O|��Jկ?y�u�$g�~�6�aR ��{���ʐ1%<X{����U|4��G"�x!�X:Z��aK�L�'@"�#D�ӝtT����	�4!�UZDG��E�&�'�X;�����v���1���^Fȹa@Z�TC䉘� �A'  VZ ��U��k�0��u"- u���^��Y�6���qW�	�ٺ��b�A;L�4��u�ة	����DP�q�@4c���:�I9�,�,c��M` G�r���R�)L�|�Zfitt��d8.e�|�� i����`ҹ"mqO��*P	\2 �MQc��7>t�%,-����B~��s�#�@Lz5��:F��Ї�L̜�2�R�儑fJ�1����'b�flq��H�r2�ϰ"����2��O����;sTڕ�v(��o��EJ�ć; �E��#vJ|1��܃0�Jvk @�p[���#������"c��<x��3#tBd	r�=�S�? N��U��'Z��=С�t�����'|���!]�A1���-d�h���B�.杲��#��8!/�9l'B����^i8�d�P+?8�^�b�j��.��xI�%��KM��"T]���F�ՁSr]��d�*��t
��Fa�#�%��v.8���k���yr��8b8&Qb`�Z�}:y M��E�ʠCV�S� ��AA�҅��[4�x�' ��NʢWwJIIA �R%�,p��ʹ4t!��C��1��֧+$,��e��&�f����1N�~Q���:Z�ftJ ���B��Gz�/^x0�e�=7����F!�p=DO�.dx�u@�d��@LqA#ǵ`�M�rMB�*h��P2~D#��\Tx���'�_�s�: �Ь�C����V�1���0���AD&_|f�I�@B�4v
M˟��2V�Q.�(�`�ǱD\�
�"O̭+�
�:�A���M�V&|�6��; ��Ⱥ��X[��yE"�hA�>�ɢg&a��C�KtD�����ۼC�I'�l�QD =+�li#�Ƞ	F��	�D��O��S=����
/o�rA�/��xƌ(��0��|�$T�
I�L���-5��c�B�2���*���6FI��a���4]�th�Ab��3N����H3V)�4oܜG@����'_����`��`2 �*{ ��h�m��
���!��xA�k�o���Ȓ�Q�l'$�ȓ']�u��kV,��x��-y�\��ȓZ2��{t�/�l��hɮ1�ȇ�?��0d9��3�Ǩ>�$��ȓNv�q�!�ݡ:h�A�񫒳%�J��ĸa��(��:=�QBQ��*�)��B�HX��
�zɮ1ڴ- �8�$�ȓl;�x�� #Z��ˏ3*B�ȓ>߂t���χmEVU�NB.s$܄ȓ�`�{�S�eZ��(�'}�I��۬�G�&Z���煘m�p}��9L,��O���� �T�ZX$���@;(�r��$@�X���:+Ҩ��wY�l@��՗z�2\�E�M�`z8L��$k�		�*.CD	�S���<Ԇ�G��S7FA(as<t�5(K%`%N$�ȓ �@�zcD�G2FA`A�P!m?.��ȓ�^銃��h�{����>���"�^���LL�NZ�E�$�ݒ5( ؄�m�@ c$��5�2��E��pp��?H1`F�6<���I�!́GN܅��ΠP��է-l��F��{E
e�ȓ*S�P"��8_�)�tCǻk�͇��ְ���)��4�Eh�)f�t�ȓJ�6�V��4�RA��(a�<Q�ȓq��ᙐ�V,u�@պK�&f���ȓ@�x��G�|�qS�'~i�̇ȓZ�:��fDǂ%�t���鑶t?��ȓ@J*��d((8��WL�7_�R��p�zt��	Z�"(�e��/{G�,�ȓ4`�B�A �@�wiك8�T�ȓ7�x�zӬ2�@�K��I?Z� !��o~v��nܷy��}���/.�r��ȓE8��Ҥ,�\6p��{"��ȓsݔ���5�r� �x��ȓt╉ؠB���%j���<)�ȓ �v�C�C[��@d��)�Ni��(�!���HNȘ�I�0��`��e`�Q�o�,tr�X�`½b	�͆�(��(�j¡�0d���7�����(��j��u,�xF��	ò��Y9�L(�J�2gހ�pb�*�����
Y�ӵ�]��,IhR.L�71z�ȓp!T���W�yHA�H�1�����k�ҹ�tИpx~�0Ҋ#w����S�? �u�ud�^�Pq���F����E"O���I9i�(t�P��H�ؤ*�"OP�٥`�%b�*A׭� ?���b*O!#f�*v�2E�V����'"(�83Eƨ*{P�$$�9�`�i�'hl�˒�3�ڱJ$�ֵ	��R�'��=S�C[=,���!L���{
�'{�[A�D�Ś���}�X���'®��Cݬ�NT9���N4��'�Z0���[�f��<JVB��(�"с�'J�9�mP-�H ��3\b����'��i[�ȬzҀ�CW��9A�����'�tU�pdT����{�D�QM����'��Ps7lQ�5�9���Hq����'}��e��,4�E)�h4G�j�:
�'�$���m�H�qq	�%9�^D
�'�x��u��59$�� ��.߰$��'��=���0������p�1@	�'@����1�`�f�!Gn��'90��4ǂ��~�Q6kK�A��2�'��v��!Ό��`�ތTR�'�r) 9#c`�8R Z9`-��'M���B�`���J���ҡ��'xօC&lы8�2Qu����v!��'
^d21���:�V��v����'�^ț1��7RC4h G�a��0��'ה���A$x��Q*�$�;dP��'��Q��� ?��)��n�2w�^A�<��Y�Q���1GΎ�[@�Aª�|�<ǥԚ.*n�i�T;y��(�%�A�<9�$�A�<�P�܏?֐ЗG�<�X+M+��� 	�.9`mh�I�y�<��͉�z �q���]�w����H|�<if�[������W� �����}�<���.U��(�&��;��C���}�<�S"�K�D��Z�56|�B�Cf�<����ZT�X3����1�e�UO�<A�"?Ox�0��){ɹ4BGs�<��@�8@�´Ȇ+��m�f	P�i�d�<��@�'>�x��D*l~Q��.[[�<�g�����Qר :=�J�!(NX�<�⮘�ݜ�[���0y����n�T�<�SO�G�a:dG20�B� ��h�<df�á)�(Q��@���]�<��]� ��KK�&=+��S�<�E�W *f��˳�H�9����a�QL�<a��Ęt���{Fǔ�b��9�'PJ�<Q�F��h��Ñx	�H:q��c�<�Ac��d1,����J�mc�$rGB�c�<�1O� L�� OW 2�u��X�<�P�J,Yz�"G� a�B0K�ʆW�<6	�EKxi ���[r�!�N�<i�.U1 �̀Z�F��)g��2�L�H�<�ČX��8�S偁�}!*��nb�<���I�
�J�h��ݦ{)�Yҧ\�<Y��Z�����"hT5Y�*�[�<�BV(��Ȁ ^4Wz��`4�X�<���B�Ohj�����;�����W�<!�_4Djb���F
?R�E5��k�<��@\Z$�\�Ҝ⠝)���]�<�DM_�y��h 7�ӑmʶ�����Y�<ia!8�*��s�O�P�P��l�T�<���ël��á� -S$H�a�n�<� � �d���F�X8���"�n�<� �-�v)#
H!��ǭF�n�"O��i�)�K��TGF��2���s"O��Q��F������-D���#�"O�K�J�^���bR�I3(�@��"Oh�Ѳ	��(@<̨��L��Z�"O���Q�X�����#��&HSܩ��"OJ����P>q�	�s��wV&��"O������"�|8sp�P6���@g"O4U�䔍T}�m��X[���"OD��I�$AR՛aĐ�lKm	�"O����28���$LY�"OA��ʃ�Y���@c%a�3"O��: ����uj"e�&FI&��"O.�#f�:
�3�ՒN��l�c"O(SoI�1*�Љ�؁2�N�@"O�㧈ڑ%bu�4��Q�I5�'V��b�ټB�t�9�͘�h,�� jW�W�B���i���'���۱=�>m9s���!E��HIt~�Z���3v�l'�����Qy짺��w_�h9��G3q�>�	 �ԙ.���p�Oy�`�)3\<-���v�xi�U���=\�����0b<t���t�s+D�zӧ�gy�)��xU ���Z=4���1I���?�G%��A|��Kӛx����5��4�T�ٵh1tD9C�9�X�Rc�	#IĚY�N��x��1O�,A���Q�8cP�ˢ�Z#F�4c�,�ƨ�d��|�'͘�"�oú#m�\��c�X��O<��������OW i�!$5��C�^.�<�vEA�?�A�I����4��S�go���I\�U�h��dD�B(����(q���'�RL�ᓤ.T<aF�5�x�y���M�R�Ñ`��#�|6��|r��AwP��$f�="�N��C��}gxeɦ��W$��9}�����,��!#$j��3UXse)�pذ�'X�Ixb���k�.��.[a#���)�*K��XZ�M��D}N���!x� ��d�%5ٶ}I��*[��nz>��g}J?}�拊7=]���R��9�N9�󉒇h��|�'�b�mڳ=�*��ɏ-du�=� 32�<
 �����?q`��#&�Oͱ��LR���DPA�+�BV��C���CT��>�|܉4C�0�4�AV�z�h�`�@�D�(�f��?i��&&�4 !$B
�Nاľ>9��AI��H��$f��G4x�s'���e8rm�оi��+���ӰS���c,ϢL�кC���F\	3��d��Gx��~�ڕ�`Yg�0s�`����}��O<��1�)�$	Ϸ/��'�X�Z�HH��y/�L���!�K�U[�a�^$�yb$�3h�^-���γE%5#��9�yRl�<3��E��@3���0E��(�y�ȓ)���CQ�H��4�Ф� �yb���(������K��f�jTb��y")�mz9�Vi�}H�@S��y���s���ҏ[
+�R��cI�y"��[��B��I�$�E����,�yrE$ja��H��H0F ��y��V8h=���Ɩ:����M��w:�4љZ�P�`m�?Z;2���F�x��e�#9�@��Å:�Q�ȓAm`P����R�lA���(�}��X��MQ��#k��]�s�_�W����r�8��
�"M ]�U�C�`ޤ��{��K�˺z\`��J������{14��Нs���9��� ,@؅ȓD�	/�M�)���"#o&�ȓ7�Q�b��m�a���
��i�ȓz��]���^���P��㜛E�لȓ���B�+�F� �ł�i�<Q�ȓ-�[4ehD*GKR8�Y�ȓ5�X SG_9W���!fʌ�KIt���f>ʽ�$�@������'9�@��ZBP� .W�a"�38Sre��S�? ��dh3~�P���()�1�&"O�T 3�8p�:P#/͗:�А��"O@�B��(<�a�6N��B��`(�"O�1�nN�.N��3��J�����"O�݈a�21
6��i�3}�$��"O��P��bBP6��2&�,T��"O ���N7s�hlB`ǥP����"O8#u�ޅp�T�-� @v(E�"O��a K!^d`���"+_����"O����HG)��=��a�wr���w"O�0IҢ[ 	J��NpZ��+"O����8#�ఠ�3-b��*3"O�T���Z4\L���Ň�dM���e"O6����`��K۱zYJ�h!"O�ɚע�:j/bлQk�A>�ř�"O(���)g��$�H�6"�1(�"O\(i�(�,z�б3�l	���"O�̃�l�
m����@�t�-��"OĠ2щ�7L���1�ؐ5�ts"O��Җ)�>��Eb�`�
��!{�"Oruj�N��H�z$�@�\򢍩D"O�52O����/ӣ�$�4"OFq�0'�3
��m���	���'"O��ܩA�|�*�M�pdTi�"O*�K�dۄ+��р��R��A�"O�Pxem�5u�N�"���8QےP��"O��ϰ��h���
Y����W"O.Kg��1�"܂
�`����$"Ox����@7s͒yS�h��\- "O^�:u(Md�!Q��*}O~5{�"OzP�a�P�H^$0�m�r��	�b"O�\������V:/�p��$"O
�Y"mH",�,@XS*f�.�I"O�e���ףm�>�[���cq��I�"O��bhO-I��XH�
M�I����"O��1�+Z�FɊM���.C�8��R"O֘��L�u~qadfeʂ�9"O�I��Ǘ�Qx�ͫC'�sV�d��"O��A�CJ�}I���!AY�b�(�p�"Oj8u&�\�Љ���~ƔT�a"O��(Ї-N�&�:c��.���f"O��`���"�T�D�-n
�=C"Oj�#k�1Y[zlB�*^�C��`�"O����eګ����Hـ-W�{'"O�\ 3eV<`��qB��c-���'"O:	���W)AKxxIDO�����4"O^�)�JO�?�H�PtMZ���x��"O�я�	S�^��6N�I�J=)"O�(���u�r-!.��B�j�+U"OrŪ�hřVҘP��ӟ�,�p�"O�U��̫y<H�3�� N�����"O�9�Mދ%e����BWS�vQ�%"O� f��?K8��`dCQ3R���X�"O�8�V� $:L�����?x�^�i3"O�0���iW�A!cM8�R��g"O���D��$�T�L�85� d"O�i�������k⁈�s��h��"Oj�(kN�)��:!�,�L�#d"O@4�S�Q>h`0��tP�"OB	�T��_�@�Pl�5qN ��"O^y�L���0�2�^9o0-��"O���FIm�h��*�"]���"O|,��
!!�� P�^4`}*!"O����&B�H����c
��3�"O� �H�gG�M�H����d�#"OQK���#���f�{��31"O<�2g�յ}�r�Y�Cլ#~� ��"O>ăc�(�(�C�CW.=ӆ�:�"O�ҕ��fD� 1B,��V(-C�"O��!����v�&P��i��8~4y�"O�q���2��	��
ǜB�A"Oj!�u,�=���'�V"On4�U-6=ݸY��Z9th��'�l�5�Q�   P� �ܥO��K�'��5�ė ���C�M��q	�'�dI�Pn�O+�d#g�K�Ir�8
�'i���ϝ��IG�Wc��-�	�'� A�,Qm~��u���Z7A�	�']�A�>J4�YU�X��e��'��!�g�T�hKt|A5o�M��!�'��+ՆN3$�p��٤S4���'}J�
��3Hr숁Ɇ>��ɛ�'TP��l�Gy���@W���h�'�Z j���'i��m���h^Q�ʓb�l����B�p��U�!��?z� �ȓ3?Z���8<��`��B҈!�ȓ,�L՛pJ�XS���لZ���XB\�B�=>�T�a�c	\�ȓ���b�E\�t�ӥZ7�z��9.�p`C�v?d��KPf�ȓl)���U�ڥ=n�����
~�jM�ȓc�dC5KOю���c+]�Y�ȓ�(���+��  ����+5׬5�ȓR��hp nD*K帘� �)4T�ȅȓE�Ū�$��~~�넡Ү\������)���!x��{��B'� a��b7PtZŦٷ�֨�$�A?6<������,�|y�4*Q�Øgq��ȓ iT��P���I�,΋T&�͇ȓ@���PE�0da��LXs ��
I�\c�(�;>ObAWL�3�p��ȓ$���c������%� ��ȓ3o4K�%�?=w^�cɝM����T,X�!J�A��D���Gk��Ʉȓ0FD�+�^(��������U�ȓZє�W�'Bmh�@�Ȅȓ}�ph`��U�
��#P&	�f�x���v��	$�ש;Ez=��j>T��4w�-�A�ߎZ�\���lۇb8@�ȓ��<1�IC�0l4)��	�p�|��ȓ���.$`����8�^L ���~�<��I�42�n/ĸ��߉K>(���'\r��N����s��4E�*��'∡:R�F�g�"� "E�5�n�*�' ��9����1h��/P�	�'�l�;4A�����]�q��|	�'?�D �Fͪ1���!*�j��p��'!Z��T&�
����O�`��,�''��)��ST��+� [N$p��'�T�z�o��N�9��Z7TOd�
�'p��b�):?��BRB9����'�*US�	N�A$4���l�90�zy��'F��CW*]N����.\�a`�'���:�HY�B� Mٱ
�'�����	��O��!5�R�c.,i
�'�,I��oӿhԸaC�
d�8�	�'P��p.ȱ^��m��aɸ.wtH�'TI�3�X��,ł�O�J�2��� b0�Bh�jh�b��A5@H0r"O�!q2 �^��^t ���"O��A��`��9 ��#C[�li�"O� ;1/J5g ��s���0KEr��"O�f��t�jȈ�$��Q&K3�yB��Ɋz��ݎi�b�#pND�"�\B�#)�,�� ���Zm��hÌ�C�I�>x��;#��W6�� ��+R��B�I�ͺP���6u��Qq#J�m�tB�*7��hz�C �2q@�hfB��%�z�s�'�>T�"P�X�2��C�;9ވ�hҡ7���"�6^p�C䉢J�pmcæ]�`���ڂ�3IjXC�>j� ��k���A���	��|C�'Є�h[�1�ĩc���7[|C�	�q�"L8�&�7QJ�q���̢ErC�I)1O,�k���6�4X�U�ɠ$�XC�	

x�0�G=�i��h:sPxC��$U�Ƶ���K�\�}�WTKPPC䉢킅8W��B�] !猿3�&C�	�Da>��� $��q "@]�-�C��,R�M�e�ۗ6BH����F 5�B�I�;�8��p�F��[�B�x��B�	_m��+��_��rHZu���FA�B�	��Zɲ#�X�V��\��	<MzB䉀�(4q�kK9(��[&�G�bB��;9���[���2v�z���M�6A| C䉎o<j� ��\$����'�U�fF�B�I���T˘(��1CD&��B�	�:>i���k��+GgS6R��D�(H5Ƽ�mF(e*1���N�Ts!�ę�u� eQ��:4T�x�g��!�J+8��T*?R�5�g�;!�DE�AG.d�!녫[bN�
R��T!�ШdLv��Ǳ\&@9dO�9Q!�dЍyOdpz���U�1Q�h�2+!�O�>d�<��b�T3<�!*�,r!�;^XZ�pׂ��W$���g��j!�$��E�Pp��X�6����'�tW!�DV�)g� �2!���1k�(1W!��Q9M�ة � ������Z!�$�7��ĐC�[�-��Ez���V!�dS�^�V�3e[�!�*��%��c!�d��r��ś5�	6��%�c�V�-Z!��	�P8��S�쐘^{�@�G+=!��0;� �  ��   �    j    �)  z3  �9  @  �F  M  HS  �Y  �_  f  ]l  �r  y  n  ��  �  a�  ��  �  -�  n�  ��  ��  ��   �  ��  )�  ��  �  ��  ��  &�  �   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k��'�O�����;-픬�ª�O;v�92"OL�p&�V�Ae�Uk��K20)�"Ol�:��a޸q�JA>W�(I�"O���*�'SCF���� k����"OZɪ���w�f1b#�?��
B"O"�S/���p���{���3"O���S��J��:�oBXY�I��"O�iq�,Ц^\l��Ψ���P�"OT,��˓>{��x!)D
z�^	(�"O��B�=2t��g��?͢-Q�"O�|�� �Cʤ�A$�z�j}�6�	Dx��"g����ب���_�b~N	S��(D��aĮ96`�+#���0� �D'(D���d/�g�ޤiՎ�?>x*C�&D����S)*��C��Hg�a�O:D��t�Z�}�T��l��1PQ*2N9D�X�rدr^��0��R��L�`	"D�L(C���O;>�"\���$��>D���`g7?�Z1#���Ĝ�zp!<D�H  닗W���uiX( \jAXE`4D��cbB�*0L�AALպ"RQ�4D��W�8=�T�+�(��m�����<D�\*sœ qt�w�Z$��!A$'D��y��_7F6��u�׆J����'D�и6藡u[0�r!�W7WԕR��?D�8y�拁&4�A"[3���#�=D�<c%�ǖ-�@�q�E�Y�v�Xb�9D�qc��G��H�ƭY���5D�(ّ-�"�4�+�صWC�}���3D��`1��Z��s�*�!l�M��G2D�Rcb1"��Hu���G�����3D���Ȃ~`�Y�����i��#D�Pp��`ɨGǋ��M��6D�L1s*�9nޭS��G(�l-�Vk/D���'#�#�h��Bj��iq5ԥ-D��c@��.�"\��f��A�=s�L6D�H*aKO�j�Jt"W�ٗB6vm҄6D��{dE�${�u�&#�}�7�1D�H�˚�/��S��S�p"�����$D�t�2�=�\�j��VN�v��E$D����#r��x�+�tAn�Z��#D�t"���g6���g��CX`���#D��J�5��cMw�V����4D��I���-!|hŮ�_�2Pp%�8D��U�F�G;DqI��
4zoH��ԅ4D�H�����2�t�c�I0.�}{��2D���7mF�@��d(��G�k���@r�2D�PpR��U����CX=�\ٱ�.D�La⠕;o����+V䒘J�.?D� k�ev���X�'RP>����>D��e%��@kdـrCE&��b D����I�]2�*֍�<&1ޤY�l<D�{�W�,ّ�L�b�h��A7D�� �0�/G0q1��hv%͒S�`�"O�=B�ᐺfPLd	���|4�"O�4�g�6��I�$��/���#�"OR\8�d�kC.��"H�|Vn�A4"O !R$��(au����I�@�CD�'Hr�'��'C��'|r�'���'F�<Bt��Udē�A�<���'H��' ��'X��'C��'R�'F�陥k�c�Ty�A�� 8�A�'�r�''R�'v��'�B�'*��'�
9(&�J8"Z-X�ˀ(�I��'��'�"�'V��'4��'���'F��f��|>ě�Ԩh���2�'y�'+��'��'
b�'���'w� JW�֕3yM�ŨK�M{���'JB�'���'���'o��'q��'D|���¾g�J�ʦ�k�T0'�'���'���'���'���'a��'��zЫG�Y��8qH
X+]�!�'���'���'Ur�'��'!��'��xc䖺6"|,���W�D�"�R��'���'���'���'���'�"�'��dA棋�@��^}b� ��'!2�'{��',B�'b�'w�'/)h�M��>�Tr�GܨC���
"�'�b�'C��'e�'=��'���'�B��C�q��W��[5�V�?)��?i��?Y��?	��?	��?Y��B�:��P�"A{��m�9�?Q��?���?)���?���z��'c�l��F���o�x)����KI8Ud��?�*O1��I��M�#�/��� `MP�7�*�&�B�g����'�B��<y�	|�K��B�\�@���A�y������?Yp�ń�M��O`�;�jH?�9�瘯gJ�q��[ -�)�r`#�	��,�'��>%�kV�I���J�%�� }����5�M�"��^���Om�w�Xa�@�\/b�֭���F<��ɀt�'t<On�S�'Jy
���4�y"&\���+u"2(<��#!���y�?Op$��<Cў��؟T	�E-fT�*F@�'R8P�V.d���'��'6���1O��3B�@[B�a OJ9��`�@/�IVyb�'�r4O
���-a$��,�;�˰3�Y�';rE��wkdc��te�ܟ`c��'��!���tP8%#'Ąr?f���Y�D�'>��9OD����Q&C�S����8O�mڌb�f��?���O�%a7)\�e��)j�o�I�,���'�r�'�B���f���ϧJ�������j ڴ�[�/�MP5��V��'�H�����'�R�'@R�'ih�CɃ7F2�hibCO=+�z̻�W����4'�]���?������<���!��qa��mͲ�@Տ���QͦEr۴�y��8H� ��T�$��4hu)��|�B=�"/�1Or<�O	L�{�M��?��8�[y���I��f�p؇�Bh�pX`�'���'�����t[��j۴_�4(���8�J�c`K�:�`6��#R^�"�'���<A�i�X6��O�  �7|�����C�f��=�K��u|6����9��3+��@�'��'I�� �17�h�	w��H�<x�ql�9|�b-��?����?����?i���O�<�xU�_�F���f*�Cq�'B�'XJ7M�.d)�I�O ��+�
�r�^h���iܮ�01�F2��%���ٴ
��O<z�a�5�,?��&
��-����1#:�$7#B,4�y��n�O�;J>�(O���O����O�tS���%��(l���\���O���<�@�i4P���'���'�ӭ@V⑈��WqX�w%+\�����O7��t�|��� Pq����ƕ<7��d�JF��4���tkt!��4�	ş�B�|R 
0���I���!�����!#�',R�' ���Y�l�۴3�\���~�ՠ-	*78Ʊ�3m՚�?����?9��Ho��Y�t,#��]��2�*I�T�ݴa��nU�|ԛ֘� 3��]�~��d�~ZP�\���4��8�.��`��<�/O����OV���On���O`ʧR2^�Z�#V�nj��K�;Ec����i���b�]��Ih�'�?ͻ@6쁡�*C�E[���쟹S�@�	��?��x���,��V���<O�t��`��(�4xV'R�F��+"=O�Y��b��?�`�;��<�'�?	�!(
���ō9��@�ևݨ�?���?����dMӦш��F՟����|�ꓤ"2�i{�D�(�6E����v����D�Ot���T�ɱH5��3�)��O6���%c��<��l8WO��A���|�w��O�1�L�<p������J���� ����?!���?���h�6��U'�Z!X� �[��w	ߖrH�D�֦1�c@���������?ͻe7�4s���h��h� �Hh��?��5����8=ޛv���a�o!�䧙&@�����B�Z�f��N�z�l&�������'5R�'��'?�tٔ��[�nxAu�̚D�N��RQ�L#۴[� ���?)��䧋?�s �4<Ȋ	���xzX`gL<�����E:�4rs���O�J�1D�M��7�E�<5hE&��Bؔ��O�y��*O9�?�A� ���<�a*Vv��8�F@�%���������?)���?Q��?ͧ�����Y�L̟8���T��0� �(�%�1�S��ß���O�����O��� ��%Bs���c+�̸3�ҳ8߆�J֢
!]��o{~�+Y�*�Ԉ��Kܧƿ� �����#�z|
��M).�� �q6Ob���O���O��$�O(�?}�V�K�X����hxNI�aן|�Iɟ�ܴ/h<h�*O�D<�$�o�������h��%z#Ĕ6gQ�A$����ɟ�Ӽ#���nJ~"N�#o��S�+�u���:t��P����Qg�|�]��ٟ�I��xk��>03$	�5
P	U�#&����d��{y�rӆ0kRH�O����O��'1�&���c�*��)�$�]qX�'��֟����S���Q+l�$[5F�Ay�1�@{;���A�@zt��O���?!�c"��+FG������>o!.�
��K'Z���D�O4��O���	�<���'��Y�&	�Gk(�c� �(`,�qS�M�5�?q��?9�T����4s��$��l 5Ny`���%=�8M��i�7m *p+l7�e���I�g� ����O�,�5��q ��$���"`��R�y�0�'��'��'2�'�<7�*��`_�Y����0�?RD����B‾�?1��?�O~��?ͻl_�Q �И
��3���[Xx�˦�'�61OX�S�S7m�n��<ٵb�by�Ԁw��f� 8�.\�<a���`���� ����4�X��k`��`���FA(�Ȟ�"?���O~���O�˓\��v��A�R�'�b��v��X�ef�1m2pȣHP3�ODʓt�f.y��l$��J�f�S�"Q����\p�Qk�e(?�2c�"�B� I~�'&���K��?I���%`��Bwj5��	�f����?q��?���?����OX5)��޹8�rha�E��T�UCA�O��nZ�'���	���Iz�Ӽ+���Xy��q��
�Di��@�<���i*7� ¦1�5���E�'T�B���?�XC	/EL8�L�#dnH���D�M��'j�i>��I����ߟ����3�Va��H+Ch��P/+y.ɗ'[
6�x ^��?��Ԉ�$@<���w�1K�8�I5��.J%��������S�'H���Z%̔H듩��]�TrԊ��w����'*�x���Uҟ@{ё|�Y�pbńS�#�"�;VDO�G&�@�@����$��ݟ�Siyr�{ӌ�q���OF �Bʕu���뤌Z"t���4O��*�IiyB�'x�Ba�(�H�i���Yp�9f|HX�`�x7&?�!aC;@*X�I'���	���dARÖ�5l��;���:G^��	������������f����s�E_�C<XQ�An��:�N���?a����雨r!��˟�$����%�-r!ntӗ�?
�2�[7�۫���?���|*#ߏ�M;�OH�Kh�6W�h��Y�\î��'<&��d[�T\��O���|����?i��B���Kc�ܺ4�m�gl�1Zy����?�*O�Xmھ{_�!��ן��	Z�4'�
²q�1�^��6�ʱ��$��d�<Yu�i�6M�v�)
ԎcD, �!��B՜1a1R�(���*ݓ����Df���$!A�|R�P.@�0��U'�&	������\>b�2�'VR�'z��dX��޴��x��+ͺ/��@�3��.RX���η��D�O��ȕ'[£Q2e��I��M[7,`R�H��&���}��9CBh���L�DB���p�O�f��$G��:�2%hKɢv>\��'v�I쟀�	�����柜�IP��j�xQ�	���"V��3#�ϥ��6��"���O���4�9O��4��ҴHK�k�~lpTm�=h�R���
�@mڍ���?��?�����6� L����L���(Z�yq�=���<@�N�O�œO>a,O�	�O��JW�șN$�c ��VD�m��O����OR�d�<�C�iO %���'�2�'��l��$ղ;1�غ���:�p�$5?A���M;f�xRGF @�4��`ßQ l��i�5�y��';6���H���H��Op�	A�?�&��O���&�3y~lKש�:b����"�O��d�O*�$�O��}����l��(٢q�fJ�؍����6ޛ6F�@J�I䟤�?ͻWz
�ȤU0Tz8���� �A͓|(�Icӌ�ldQ�(n��<A��<:P�����"�`��͜%p�F
��i&�`��#
�����4�����O��D�O��d�.J7R8!P���1��BF+**�ʓ9u��gK�2���'%r���'����[�n�}���ǜ/i40�[����4n<�#��)�"H�J J���H��x�D�1k#
��pb �~4��$bbF`��'�hX&�p�'ؒ$8A�@-._�ܱ�hM�H�{��'�b�'����dZ���4f�9���o�N�
��� �r@EZ*a0�%���?1��^�8��ПX��4Q	�K�b�j���#�(/���{B�*�M#�O���������w��b�4|T����݈X�l��'0��'�2�'��'E��9�Hۀx���%��^�b8hdl�O��D�O�]mZ4B���'��|Bc�;`I��iӄg"���o�a2�d�<a��M�'7g�=�ݴ���ǄV�@�K�e8���0̄�Y�^�Ӧl��?�#(�$�<ͧ�?���?�N�C�$�wgSl.x�	���?������ç�Ɵ �	���O���Sk�b�D�l�'{��K�O���?I۴�y���<\�(�s� �R���ct-N|��E�h3^�h����)�RjQ�	��<YE�9W� �FV	|����ß��	Ɵ��)�Vy�Co� ���B\��"7����c'�],��O��?��iy�'���K!aET����G�u��@�'R6�P�\H�6*?ɐ��F���,�� �x�&d��X�"�1�$�$㔱��2O���?����?y��?A���򉅞��)q��&Q5Г�ڹ>&d�l�K�����p�IJ�s���i�-j���$�s)=.�t�@#,�ʟ8��;��Ş7!0TCش�y2�֕+;���@�X���t	�7�y��ڿ��!�	O��'��i>=�	�"(Ш��Br]`ph�H�{=4)��͟��	����'(6�X),1���O����w�x��a;��'P�kw^⟤�'���'��O�0� �,8�8�1j8����0?O��Ą�2�xq0���I�I�?��0�'��I�  >��KÔq�L�R��Ps�Q�I��8����T��b�O�2�"/ҍ�Q"�Xl��j��j�bCw�r�h���<������yW$�6��)��~(��[�⇶�yb�'�r�i��\��	m�B�	쟌p�j����c�;X��[E�
'o��=b�����%�,���D�'�r�'��'%D�8��Z�cs29��G�	k�`�yV��Q�43�F\���?����'�?�u��"`D ��5���ʒ�)��$�O|�$�Z�)�Sn)��k2J�^<r�%�"4*T"԰&���uE�T� �OƩcM>�(O���M2H#�a��,��X��Y2@F�Od�d�Ox���O�	�<պi��5(��'X`��ާd��IȰ
#b�|x��'�B���<Y!�i'x6̀˦�Z1iUp�446�2������X��Ymh~�B�^d�S}�'ݿ+gf��9�ġi�ʗ�9> �/�<���?����?i���?)���l�S�z��c�Ӓ7��*"!\��R�'*«a�TQR���<q����R$eȃ�G4)�L�ya��'y�� ae�|R�'Λ�O��!K&�i��I(&2��VBQ�@��-� V�q  �h/)��T���BAn���i�����b���?�c�	��@b�K�	N��E7�E�TϨ}���?�'��R��M�<����?���i
�OW��a�Ў��B� 3Ė�7���r��MЇ�'���'����?q�I؟@���xP�H3Jm4�P�.`��`@�z���A�4?)��T���-��2_�Ԡ�ᐳE� �����Z�&C�ɵ|�~A9�h��c�A��L�"&M���$J1D��;�-C�b�	�غe�����Ӽ �t�戊(���F�n�P+��I�z����j�-t�xA&�ت$xr	d��2?�~	S�A�Rƌ�;%��5W4�D��;�8EEϱM�ƍӄ��\��P3D�L���Q�zh˟2J�QH��VZ7m�;�����-#��ѱWǐ�,$!�0X#H#k�bE�$&t9��y���%3�$���V�IhT�)w
/��5�r��h��BQaN�Ax,����B���+�c#�5��A�΅�! �+�Q��N���A�hR$n����lj0�ҷ��
i�\ai��pT!�E'g7�o���a�`�EQI|DedC�LԀRϒڢ�x$#ȼJ���q�D�/t��Y��ߘd�.�h&C��?���?ɶ	o�
s'�z��T�O��.���ן� �gȋI>�]��"�]ر��ɪ4PŅE�YvHًT�\9���'�X|�U�&)��]v8q��~�r�yb�ɝ%v��$%ڧH�f�+��[{ܜD���&pI�݇�S��tbr��$a+hM�J=�]��I/��_}DɁ`�"q��s�.K�"�f�<y
�	$~��P�;�����E̛H�ȓ3�x��'��T�];f�.�@e��6hQXU��'*7z��5�y��ȓ=��e� �-t�$�"OKP&��ȓG�.�
@��6��Q�}�DP��IM�	���N�8���C:�`�ȓG/�mXE��| ueK�G����ȓO��4�[
,�2xu��3~(�u��-d����({4��D�M6!�ч�;j]���0�"����Q����ȓuoV��E��3p����Bo�7���ȓ:��)SrF�/0���2��.Q����eR����T��Ub��.!�	��:�	�<�t�S�J+�P�ȓ"�T��"��?
~}B��x�^%��G�1��O�Yx�"���#lv��ȓ���J3L�l��q�:E@rه���8�(ȉ�� �gy�����"鑳�/_ނ%	���f�A���-pq�5��� W�>� A�ȓ9�D��&)x��;��AWkP��ȓ[�V`q�@�!���#��ӊ$�8��[�t� �+B�i�S�R�KTчȓ��l���T��J�00뺵��#��!ʦ��;�nY"GKa����p:DLp���4Q�t(�A)L����S�? pT�'�U�g��L{r+C����"O
H�3Ɲ�b���Ã
�6� �A"O�|z��D1�0�3�4��0`�"O<�R╞YR��3ҋ�"��m�Q"O�ၐ@��Dd툧
rp�A�"O�a�6�ʫdrX9�E�[
!d<HKG"O~i���գش��W:MG8!�"O�������H�H�*N���"O��l�6W�<��2#�2/��Bd"OZ��ሟ,np�H�(�]�a�"O̔C��[�*���΂�Z2�Q�"O�@E�4W�������:'VjY`"O�љ�DW.C\�Q���hL�#�"OV�!B#̰r�*�� ݭ`b}��"O4�@F��!G�"����\�6��"Ozg�N6��Pzg�?+ʵ9"OS�h6�6ظsA�%�q�"O���C.�6ŰPy�M>i��Q��"O��uH�\���I��:�
�t"O����Ȍ�}L���PÉ�N2�8�"O�ʄ&��q*\����5n��s"O����,X�n�f�RA�#�9'"O�!��-	g�Ȫ�j�5Y���P3"Oz)4!�`}.l�E
�,|m�"O8�Ks��C��[�T�p�9�"O�L��Ee@��A��	;l 1�g"O8D��n�Q���r��MDZzqx�"O�yQ��)Q��ʵJ��}@�p)@"Ob�+��h5t�0ѦO<X*�"O.�p�?<�:	�GkS�,=�i�"O���B�d�f�z��]�����"O2�CW�|t���jj�<���"OTй�K�42r�H�Y��P�"O�t�eM�r���tbȐA�hx�"OL�I�'��aP��4�Y	F.(!@"O �W�?J����;S����"ON����>~�6�T*�:�R�"O|�ӕ���:�!6�A
r�PA"O�1C�'�Y�Æ�l���Pt"OLq����;E�xp"��#���C"O�;�J���(���חƽIp"O�<i��4� �hW'Qt���v"O )ޏQ�h�!�V�0�i��"O6ԡ'�	�a�Ѝ����� X<8�`"O��sЊC�bL�#� lJ�L��"O.�:�O�X%�`&$� 2D "O����H�+�jѻ�Ś68X�@�"Oؕ���K�����8MJ�0�$"O�i��MA'5	X�H��Y�FԊ1Qp"Ob��0h�(g|�S���d�qz�"Ot��5�����A�M�O�PU"O̵q�7a8�@�a��.�l컆"Ob�r�i�V` "�&\hiBv"O����5n�`�ϔ7%�*�iw"Op4´�F�r����M�h�vyc�"O�E��G0 cԢ�ŕp�٘E"O�����W�xD�Ts�+VC�@<�a"O��G�+P�X@̎�@���)G"O�@��AB�fz��#&��sw"OqP6ˊ&Z`Q�DАX�X�F"O��ɕ/g�\,����Mp�}��"O�\:�/��9[N�!�7U\�\�v"O(��qKJ#P2��M�d& T�"O$Ũd"J1]՘pI�,ˇ\����G"O� ~m�hѨ1V��G�Q;[�X�q�"O��V�A�(:���1��H%f芔"O~��u��]�č�g��-�$ip"O	3�c��Jq �Hf��I�b��C"O�� ��!I��D�c��	C��x�p"O���lX�qz����J�"�x<�"O���Wʌ>+��-2��[H��1"O�A V��A�f���[� �l6"O��"��3x�Ԙ��FW�"o2���"O~IGAY����7�� �p�F"O�YK��M�N�2|c �	�^jRHjc"O��0f�T�^�~(��@�v;��""O�U2��!m�����m�0*f��"O,�2��9�|%���ژ���"O�	H&j�+}+�),�t��3"OBH�B;$�@��?o��$"O0�� �G�X�(��ή*%"O��g!v�N�
��!�"OE�3D\��PMdmS� ��
O!���.2"��T�%g�.2�!8nM!��,��
�=��P����1�!�
�j3����C\�hH����)1&!�Dѓ�C�+[>\x���/;!�dB�2Ɯ�2�=u���c�V�	&!�$��ʈrQeT ����+��K�!��14�FyCࡂ:9(Xj�5�!��^�0p�����3��ڹg�!�$�p��IW�ȇ- ��rD�A�M�!��
,�R%�q�K<l(���D���w�!��e���k�(�*�Э�5�E�<�!򄕵L� MX�ɲ��<Z��V>V�!�DšE;��j%@�6�� [��R+j!� Jq]��K��*�xS�蚔*g!򤍛ޚໂ�L�9Zs�P�,}!�d�Nj�w�@�x �����
�Oc!�d�+f>$w���vIPY��"�M!�d��rH:��Sϙh��X���ϰC>!�$	2�N(���M�Yi$Y����m<ў�JF�ӷǀ��#,Ľ4#Ψf�SnB�	/2�L?{��M�i�%(&��$S :���"~���c��9�G�A��)R�k ��y�f���tX�oDT��$:P)����Ӫ>������0}XX�vI$O��p@F̶k���Dܖ]���I_Jq�6Aѱu�����LxrB䉡C#����lT�"��5�
Z�=ie�ȸֈ�>$�7!�	u&�$�Nު<JV��#"O<�@W0o����:16�ܚ�'�t�p@(�)�M@�CA��T(�w*����'��pB���*4��@Ax_�X��OpD�P�Yg�a{��19�A�W����-�7�Ս��>Y�gT�{����N�H��<B@�ǐA.Z����ϒU�!�$�&��BÇQ9�eQ�ߐKF��\0�l�������!�0}v��4k]�9GdM:d"O�u
�$�N���1�ă6A.�`��i�����/�)��9ǋЍe ��Sæ����C�'D� (Vǔ�S�*���l�B�"����>�R�ħ�p>�b\�VcB��F�G�<1X@�a
�pX�����2�y҅  w�@���l���8�#�yRBS�o�­ìȐ\�"�X6f֭�HO�rZ�|D��C�3hrY;�AL�h*Ĕ����y�k	�U��*e�e�*��J��M����>�O?7	:>j8�Y��1�
UȣI�r8!�$�}��M#Ԧ��9�:8�cKI�3�I-��|2��o��KcA�M�L0���W��y
� <��cٚ)L�	7	��H &}��"O�g��	Zz�8jQ�n�h�"O8DK�.<��(�-\���IJz�<��gZ8q;|صD��dڒ�x �Q�<��J�2��0����OVv��T@�H�<)�L�J\��ҢT3h�@�%n A�<I$hYp�x�%�PWv��Ю}�<�iF��j��+�"J3)9��Iy�<iw��_�� &�$�I��Wt�<��4"�^Y5O���`[ �
p�<�`��1�Ό�a��n-SU�Zo�<�k�_��1oT~�
4� �j�<����qdx�)�&_�(�a2p��h�<�"?��Հw�]I��Ċ]�<�O�j?��X�풭CD��q�X�<�l^t�l����/|5x���j�<y6H�%Vϐ��e�(!ZB��3g�<�f� i���xq�G�Mzt��
B`�<��5Jr�D��B�v���!�G�<�Xfa f�'��ivfD�<�	�o�6Pk�+V3Jq�9t�Bj�<ɄL��V՚��P�{\*E��)Th�<Ѧ6T��E���ͅ<�Qr��l�<�e� �|��4�� (Y�IRɆ^�<�b"��	�v���F<�`�`4W�<��	;1\�t���8^��t0Ӣ�V�<�3�YG����&�6-���II�<iDK�hn��E�ƍ4j�*�$�M�<aM�!�����JZ�d܆��3NI�<"�G��<v� O=
P3�H�<9��_23[4�ѱOtxD�G�TV�<���v��H��;h��sČCS�<�b("J�p5H6Ċ�}�]sT�<��)I�K&2 X��P�eU��#� T�<! ,E<&��)���)p?#��]P�<�A*�,>����H��`9F�N�<)���-��iy!b��B�0����n�<�&�l�� 3bȠ ����G�Fg�<!Dl	3~t`(0��h�:u��Od�<q�S�vw��⠉��5�Bȕx�<���'�P��w��	(�Ae.{�<)@N�,NW:l��(���`9��Ds�<���G�$��\%���J-�m�6K[X�<AP�ޥ=֠��.�wE�`!�_�<B�D�r��`��		��pvF\�<AgC�c+����-b0���dK}�<�C��Z�(I�GގXƒA�1�S�<�#e�
�ه�ۊ3~CC�s�<9�(�)�� �K
}��5��r�<Qϝ}�D	!'�V/*"�d�z�<I�m]2�؝���Ǎw��Q��Ot�<��lD)Y�H�s1��0!d�Y�$o�<!���8)��[s�� ^�L؆�m�<�F��"���pF��� �l�<���O,M�` '��C�����@�<&�'RW�!ЬYh�aH�n�z�<�S�	�x�A�ͱ?�dL�F�A�<�7hɢk�����,:{�L+@�Gy�<�p����-b��B(t�[�R\�<���(/��I���$w�x2'nKN�<9�ӷrG��K�"�+l��9
�'��၁IS��*����ڔ?^����'��|�$ᖤ~:��q��=c����'�@*�H�;q��hJ��05�Ő��� f @2X/JYL	���:NV���"O� S�ծ9Y
aq��-K^^\� "O��f��b�8U�K�c� 4��"O�A5F'</pP(��g�Hѳu"O��� ��
R�A!U�Y�lpjg"OBx[C���JIz@1A��B4"OJ@3�>y^��⏆�ؾ��U"O.0��e\YZq�	X*���"O�"�m�df<�P��W���r�"OB�R���]Hlm�
W	M6M�5"O���)��uؒm�HV�gC�(�D"OJ�c��\<Pْ������B��*#"O�����Sm�x�g%� :x��"O�I�E�X=�R��7Dܥ��"O�yW���_�.���%z�P�K�"O�����/"����d�h "�"O=�cj��x�&�H���#m�ق"O�=�2�)h��X�DBE�|P���a"OF؈��T�؂�����,}`B|�f"O2� �C�,P��y�!�
N�53�"O���3ߖ!`��&M��5:"Onqⶍ�(3��,{Rˏ� (ɠ"O~qR>-`�x1ݟC;p)�"O.x�%��;�D�5*�%1r	�g"O�3��Z�'[Xt9�iҨG�(`9�"O^����UH`v@[�H�gZ����"O�PÒ�&@��	r�,E��b'"O�4(T0J�R1;CoX�r�8�"Od�@�#�(Ժ��c�SÚ��"O0|���2a�t��QT#�<���"O:���^R�4oC=_I�q��"O��qHTQC��#�ԐD"Oޥ��ş1�h0B��݄a}8<�q"O�0#�� j�d�F���UPv"O��aa 9����`r2!s�"O`�����|$� ���J#L��h�"OXuBu)� .t�q����8� �"O�4�b� ���JӬ��<���0�"OJ���lƻ>���0�ʻ[ؔ(�D"O�]�e=n�n�"��Ù�Ɖ��"O��Y�MJ�hh����Y�)��2d"OFu/ٚH�L�q��D,w�yX$"O�x���f�|�!d��2���"Or�8ƉjW���f��l��p��"O��Xrfɜƪ �ȯΘ���"OD���&[� �氻6��;`��A�'"O�� �iض��Ss�\A����"O����/��0���.�:���"OZMb1�)~B>II�+�����T"O�e�C�EY�0�`�6>�Μag"Ob�۱ƛ�;�8�VkI�I~"	[F"O�]`��H.Y��U�gպ[b�U�`"Oj�"�I
j�X��E]@�`i�"Or�q#G�c`���s$Ͱt5�L�S"OPp#1��j��E��iNa7�t��"O8Lڃ�h�H�P0��n$B���"Ohg$ܧ����`�@:?��5a�"OVܩ$P("�t����jJ��"O�����@�B8�`B$��4B "O�Rc�UH�fJ��c�X3�"O���Uf�".�9(C/�5HS"OȰ�O�N�~pBZ��(ݩ7"O�t���1. >��C+��'ͬx�"O�y{C/�i;�3���9;��A"O� �ȡv� \/�œS��jD�;�"Ol(�k�f�{���&;��Q��"O�d[�b��s�\��!-&p�*QI�"O<�x�#�8�\�ENV�|�����"O�A���L���X׬+F�H��"OZ�д|oΕ22�N�:�8�3"O�Px�J�0xr��0%�n�r"O�X@��%:��%s����K֭�yR�λF�X�	��V�6����N�y`̱z�Jł�%Q\Qԩ �X��y�O+��a�s��* 
F��1�,D��KGd��k��`FSw�p�:0G'T�0`a��/è���)�i N��"O@�bp��(B��"��2@	Ze"Oȥ�u:C����� G".Ļ�"ODU�E�I�&q*� �╇O�XY�"O�x���TF�[⠃�]�X�
�"O��H� Q����F�����'�\X���d��9�eJG&J���'��}�R!Uey����ε�	�'�|DY���T����"���^´���'þ�	Q�X�V%��Q׎��u�H��'��x8��D.�֍I�KSY0��'�>���ǐ�����U�~�|H�'u$=s�AϹR�"�ئ���A
8���'0V0Ä�K�Dgz8�q�%���'���2�kȃ(:��d��%=T 	�'��u�
G
w�����QI@0B�'88{p�ٝT-����2,W��q�'�t"�a��Q�<Q%Ǉ�(N<4��'��L�C-�&��2%/ޜ
�" ��'bxӗ�2ބ(�D(���:	�'���[Ç'r-Ơh�f΃|�w�y��O;D��r6k�42�� �dҊ�yb$H	c\����&����f ��yB%1��� B�"�b��v�=�yk�/o�]�7���Q�#J��yg�u����rD[�!�0��B"��y��	�F��_�f�&i��8�y���0^3�H$t��=Z҆_�y��������f�:�@��ya�$vL�;��Ip%Q��L�y�J`2��j��L�=��i{c�K��y��Y�l5"� �NK�#Jb� ��y�մ"��!	C�\9LN\�D��y"/ӊ9�$0��؈N y��,�y�H=;��:VE	1��ٙgn��y2�%�RԨ�N�� �t��_��yB�?�,���z`��ec���y"�8*�\8�liD
�iD��y�@N0����/~`y�0��,�?����C�T��冲$㺌p0�E?X�ȓp�theA.:���A�- �cs����x�V�9cK��g�`���)M�9�*���2� l���ө1��@�g�|�
C創~�pH#�CNHd�c#�@�B�I�	��K��?k�`��] x�C�
10Rh���E.?t��x��.O�C�0hu�E�WG�l�����Nu�C�		1�M�1�m�a� e�':DrC��#hb�(��o}� 0eL1b��C䉚\]>9�%�(_�N�����Xl�C�I #��h�c�׳<������B-)O�B�ɬ0O�����r�������,+a�B�)� *|BMS�Sd}�s䔯���;�"O�`�T����z�yщ���2�"OCu�V�(���&�L�O��"O��v#�kF�:GT	vhf�i�"O�|⣦�5>��b�썝2�
�SW"O9	q/��.�"�Z�+�4P�H�P"O����G5l�<ٻ�����$l�a"O0�A�
Q�l�,q⒄ڎl�rܣ�"O �.C�d)����j�4�"O�е�Z,��٠�(��$�1"O( ��up��7NGc����"O�$���>����ȪQJ�8�"O�9b	M��8�1��@�C����"O� R!�(ʊd�#˦M��1�"O�az�LO'�)��C�f��iA�"Ov�hW��n��lH#a�|��"O�SӤ�94��f�ȨY}p�Xq"O��ӣk�PȈ��T�S� �V"Oġ��Y�n��� �L�K\�p�"O�m��cP�q�h�1�ɡk_�u �"O��a�U��s��B���3�"O�Ё�݃h�ޠA�"÷k�����"O�@ �,Y�E�Z�<�([�"O� 4�M[��|@ �Ⱦw�D��"O�LA.Ð���W-E6d،��"O�xSŎ	
�ڑ2gM_���x�"O�p� [�b�pa�6/�����"O]��`@4f�q.O=�t1�"Oڠ��m�O�\ ��;
o�k"Oj)P.0tD���C�8m��:�"OԈԤīN��Q�q���{U�pP"Ol�E%7�(�&��6k�����"O�؆�L�x,���J�O©�"ON8�D�.k�Ye�To��Qj@"O
�b쒧bi���`E*���{S"O���P���FX( ���C#:���"O4��M[�g[�m�d�,2d�$��"O�pr֞ڮآ�އ\Z�8	�"OUh%o�6fX)��oY�-B���T"O��s�.A,4>�����>�|8"O:� �j����O���2xJ1"O���*����ݲI��a"O�P��/�?�ni@ڈ2� "�"O�u3��G�Q���"�.�h���#"ONBb.n��4ˠZ�yz�1a"O��zd�MC'���=xL���"OP�l���9�#�ǘ(��`�"O^=��/N6|B�A�6��9G8���"O++�%#U+7�˓@�@���c�<� �ǆ[��M���r5k5lc�<��L�4aP�Z I�)�D�C�z�<�q��@U�0*ab�+bh���H�x�<y�,\❸!CL�<�R��'�u�<�A,�:e�1Y��B&8�p��2�W�<9r�	�4��ub��h �9�S�<�l�.Ge`���f��2�~m���ZU�<Qǯ6sΘ�Zgď�/ (����N�<��!Ѕp ҈r$��8��r�RK�<�g�al��RӢ�	�Jň� �I�<	�)R�wXкA�Q+�bpp��JI�<�6��5
�mq�ܩL�T@4�DF�<A3���*���a%b�.N�h��g�<�֣��t	ʄ�UO��<(����`�<Y�/C�I%�RE@��
D��X�<� ���ЁGg�.4�4�/����2"O���6�H�Nh:�����n�t��G"O���d敂E\����`ڼlݖ�`�"O�ܹ$�'O�����Ϛ�6Q�"OnM�Ќ�XK��ל]Ê$�f"O*�	02F�<0�.�h��ɳu"O�q75~A␁!�Ѝ*|P�t"OH�� �<<�~}p�fڵhQ��P�"OL�#�"N,����˼3d��bP"O����E^�gߤ�@��]�<r@"O \����.m���'	�	�,˔"O�]7	��H����eQ�p��"O}B�D�(�8��Z�"t��w"O�h��x �qE�E�dVԍE"O�I�`����ŝq:>�+�"O�d�����>:���A��$XM~�t"O���4��u�g8I@ɰ�"O�\Ä�N�R�J}z��!EHq�"O
�1�4��d�g��BG�|p�"O�@7.�&J�:lZ��~Z��'"O��+e�F":���ՄF�!�LU[�"O��cٍt���1�9d�@Y��"O:d[Pؖv'���֧�uвY��"Oĕ���>���sUFU9N����"O���w΄�Wd쳗��<v�i"OZ����Z�2�°g9�E1�"O���e��&��Z��� ;�9*O.ȒƧ�e�&����.+҅3�'�ԴaA�_�B�BC/�8ohF�H
�'��"�$Ӥ=I�� q��Di	�'� �G�̊n����OV�5�~��'b��r�T?F�v�!%+U�-�J��'����g�O!Ӟ���)x����'	f���d��"E����Ɠ����'q��R���q���3��Ӣ#+.tZ�'�v1V�ʨW�DQ@�'�N%0�'[�,��D�F;6e���F�(��'M���^��vmBJC���'�p�;�I� ��H�0�+ ���yB�p=��#S�Z�nʺ��K�yb��6�n�(B@ l��hW���yB��K��2�
c�P�kZ�y I ���"ɦZw�(�dȏ�y�_=<����RK�cUc �y"��a���r`�4L��1cR.�y�M�)�h,�`L2E� � �#X�y�@�~��-Ku+((涤Bp��;�yҏ�wF��bed�<I�8�@�y�j��.��@ĢSP^�lQ�c�yң�Ja��h�fM�W~����
�yrj_�!;6�V�W�Nގ	�����y⮛�*���E�)wC~�u ��yr>cm���-L�t�J�9�M��y2�R,�ؽCa	@r�a㣛 �ybM��H������iF�4!�숕�y2��9yb�2B�ɤ,Ӝpz�!�!�y�͎�q�X8ee��"�%�f�"�y��2W��ق�ʝJ�qo��y�ѯ/��c�+�3xt �5@���y2m2"Rj��D�±~7>}" hI;�y2�Ή(���K�{�]{WE��yR���$��A�5��3f�PM�E�+�yb��"/�H�i5�@5Z^|J�H�7�y�D۟-'Čzg�������]/�y
� ЙQ���u��]�c@�t9��Ȃ"O�Q��)X�C�b���׎@�ժ�"O�mH�D
0��qA�%}�А"O�l�$C�?3Ԍ���G� m:�h�"O�͓�g�q6�����'}�P��"O"���0�`�Ǡ<o�|{�"O���)N7��+ �"ac��K�"Or��&!q}n|`��ۺ&Q&��"O
mȑ�S�������	%��I�"Oĩ!4��M�-Y��Ɩ`� ��#"O^�`�79�J�=_����@"O4���E�qҤ	���{�"Y�&"O�9q���ޞ4p�d�3p���"O��Ѓyg�0��e�*G�lZ"O�;���aX��5ʗ�{��X�"O���M�2u���0@Ƽw�e*�"OҴp׀B�W���?j�P�d"O6��!@�E3Qd&ǧS��A��"O���E)
4��P0+�d���D"O=�"��tq^��E�ҩ$�"��"O H�N�D]�����&�� w"OH��5Z11REْ�U�}%r5"O�)3V�4
��*qM�&��qs "O���F�>(h���S֗o�}c�"O�4(BfA	
k�	��d�����P4"O��s��:
��S��0�o=8�!�D+�K�惋v.DI3n��Aj!�߷�%� ˠS<�I���k[!���3�<��g�p��`أ�P�N�!�$��,g^�*W�a�� 
#GԻ>!�s�8�e̯�@�1����(!��\ɶ��'S��&�(!��,j&����P�
ڬ��7�/z�!��R�Z�l���'�6g�ݐ��Pjq!�D
;Y��CR�[
w~�!(6HU!��ڧ#��]a	w�J�`��N�!�D��¸�&��:X�����G!�MKn]���BY��I�G !��&lȌ��- ��B�Ӝ(�!��A�!ӫ�?)T���A0w-�لȓGt^i*�ïj�����琑Z�ن�n�r��dm�%���w隋od���J|��
`. F�ֹʳ��?�ֵ�ȓ)ո�`tC�*ikL)�'�	� \�ȓb�릈Sj��*�"ޝ^��U�ȓ.�61#�L�A�깂pC�>�(�ȓk(\M:t%I+��rf��H���ȓo��C�G�#�X�U�֖̀Նȓz���H�k�,���iݒ>���ȓs�^��U�̍7�Z�0#mմG�	��e�F�p��bzdx8�	�6wpD�ȓ 66��Ra��>���Z�n��!��cr%��Fᗸ!2�x���H�;�!��-oS�mj҂��d�	����.�!���I<hgCe_�J���m�!�n�y�1Β�FX�p��M�!�!�$�&ez�{V兿l�䃧�D!���a����$0}1�*!��+BkB8�B@�E(d��$.� !�d�(C �8g�� ����v��L]!�d� ��|s�M5i����BT~�!��].&7F�B���K������!�dť%��᪂���|�*"��e�!��B�~\�A�_,�ָ{�N-Y�!�� ����3'&s�Ն���ң"O�d����B�f1DMZ�m
љ�"O�9gŅ�X��sk��U�p��"O��˲�95-Pd+` ܥY�^�x�"O���A�E�.W^ �ӮV�%�����"O����24D�CW��m����%"O�H9�G�C+�Z1���?xf��"O�19��/��"S搟cg�9("O69�*�}.$0��´�3�!��kͼ�H��Q\�1��nJ�z�!��"f���u��cn�"�.ɲ^
!��0��hiԫ�jMb]�s���f�!�$L�+�K�?>�sPD��r�!�,>ZX�!u�:~�k6F�)P!�$]-f��OE�w"i2� ܭa�!�D��l�����3,`����F�,?�!�$�k�~��W	�
y��A�E�P��}�$ �+�&(P.�a��H�U�A0�.ړ�0<qFoβ�LLH�\iZ�	��+�W�<�� D�J� ��Sj��dx�Qh��O�<1AD��`�U�ٻ-h��!�GO�<9ArHEC�9g4xp�`�<��N�}��Av#�A���˓)_�<� �#S�RxJ��C^a���U�<�U�֗Z��h���	4�Z#���S�<��g�.L�Z��15l�,��f�<�v�5�V��1z�~ �bi\[�<9��Ԏ[���0TcR0Kt!!��Pp�<1��D�m=�P���ԮK�ɰc�`�<y�`�3q$�Y
��҅і���l�_�<���i�P�D�O�9 , 5�QC�<��.ĺ#�02��P��T�-B�<�CaԕRp|P9�J�pz�V|�<1���>aPb��JP�+��{�<aQĎ���\I�����*��1�Oo�<�W"=?세+�w7����%�a�<�쁖sM�h�3Å�2,���Y�<�b���HI�Y	�*��m=.QRc�Y�<�D�A(hI��ʕE߰#�$-xS�}�<�p�%,t� ����Q�v(HF�}�<�G��9 �yS�Ё47�a���s�<�fŉ�rg���A�Gx
l0� �Y�<ᰄ�H``��
��$��}	�F�W�<��I��ݨ	^�	�zLA!΃U�<ѵ�G�\�>P�%�_�'�ܰ�sBT�<�CĞI�&���gu�t����O�<��̊�t��p�J r�dQ�'@��ȓ���S��,u2p�>;�h)��C\�0��B!`���	f��h�2u��s�r�!��[�U>���o��U�����]� Y�2ID�H3ܩA1j�-	�b��V�z0.Y���zTH��7l�ĢE�2D�pɉ�F�� 셅t��@�N1D�4�����qȀ�§0#t�P�!4D�$�dO�
]�e��>H>���0D��q�F�:=��S�u�Pi.D��W�E0��hԍMQ۶����*D���p��3	▅�B�Q�bh-D�q��h��BC�X�fފ�9��8D���!��i���fK�>�r9��l3��o���@�nN J��%O8�.eB<D�pb5#��F�(}�*25D���3*R#f^�ӧlW9?z�C¯.D�<�sH��Pl)q��տ~Pi�F!'D�� l�����>��D�Uh��a�,,q�"Of�R�딱v�N�q�Eۻߺ�Ã"O* �S�$+���W�nx��"O�0��]63߁/�ܑx"O��pw`#`z��� ��i+�"On�sqC9�`�d�8��!bg"O�h�Ԏ�}ֱ��&A1B�p(��"O�a��6R2T���V�DIC�"OԈ�-\_6�1;�X@3!�'W���B�|�Ps%H7y (9���`�!�$	%;�vha,��;�ɲ���if!�$6|Ԗ�� (9��)����?T\!��U#G�~}�Ū�1E� �*bP\!�$�=\@'	֑R�X|z�b�H.!�+nw`4�`aРI�h ����M!��KY��͖������Hџ,������|Zp�Ҏr�b�
��])]LX��N�<9 �}�8�q�ҤC3�Ec``K�<0K�c�h���Y6&$(#w��b�<q�G�5z�>����d�4D¥N�r�<!��R�+�y��Q�fCu�<���7KAܴ��-�2ao4��w�K�<i�/�$�Eb�̌�N�	��E�<y�&U�|*�eëG�֑���X�<�6i��8΀a0��~� 0"�^�<2F�S�����s��	åe[[�<�� � .�r+c�P��2��S�Tl�<yQ/��n�t)�G�j� �nVh�<��R+rjL��0�D�$��L�<��E�����&]id�
��W~�<y���I�
ģrm݅_�hiBa�ET�<�dJ�f<@�⢇�N�P٩a��T�<1��	w&L)y�B�v�<���^i�<�#�Y U4&�+�F�6�hH���f�<i�#��"�,���jβHXөS^�<
��P4C�m_�wA��dv�<2���G�lLp1��qH���'�s�<D��0�*-��i��kf�s�<�c�7���cf/�ETT��#� i�<�paF�QP �JPN�iD������e�<A��L�$;�`�9A��skTx�<�u�� �Q��	2~V��۴�L`�<���C�wk�1قN\�t{$��F�<���ͣ}:鈷鉑 ��e�6 �Y�<� &��C�n|ʑ�H6�eQ�n�<a�ޟJ�ȶH�8(,��jHi�<��O�]��R�C��j��H���e�<�rG$BB61:G�q�$1�.�]�<1��7)��`@��,F�oh�B�	6hCR]���߃W� ʓ97~B�&\Ƅ�������8d,��&ѦB�	�chV����S�Y�T͘���2504C�	�w����(��IE��(�4B�Ih��i��ͅr��\x� :
��B�	 `!���w�����ϝ�5K�B�ɳ\6H�'��1)���*6�� 4�B䉢I�H�"  ОWp�|�4斔,�B�I�9Q�Y u�	�czhZrJ�uJ�C�I�`�hy�N��Q�\�!d
'Fp�C䉵�(�@��U��QQ�C�ɫ�>X��O�!'���0$��2s\C�ɵjZT��$a�)I���A�G,C�	�J�!���	3<7Hb@�B�N�C�I�zI
��B�(a2|s�eK*X�B�)� X(�b*�@��m�]5T���"O\� �R� 6�A���<!;L��"O�X��2��)�#j�t��"OJD��ċ�3��x4��4�u�"O��:����1#��8/�6`�V*�"Oh�p1�� �ȧ��aĪ �e"O0}Bt�Ipr�� N�p�{"O��[�J�g��;DB��A!p���T�L��J�S�O+FEʦ�*�n�R�#Ѡ�n\k	�'�n�q��S/]~�X`�&
u:T��'�|�Aq�ގ_�	zd%		���'/�2�A�
r����lE�y��k	�'�,!Ya��,�2EX�JZ�t�Vii	�'�5"%�\���V0+��٢���y"�MJ� mˆH#3gj�(wC������O�⟢|R��*
�<maR&@�&�R�2A��f�<�`ۯN|�U"a@/��	+c�a�<QG�
)�09�cK�@���*�T�<i�)Ծ+#^`q�D�&��I��k�<i"<bQ`�� �޻3���f�<�u!V�̓Wd�#xm��8�K�<��Iׄ�p�C��b�A��p�<�4)�$t�t���aP�,`�"���n�<����VX��e�L�4�8d:�f�<I2`��_n@��ΐ�vV<��Eo	|�<�P�֚`|�S�%~́EIy�<�R!O� ��E��̚?mU��{���t�<Qdd�?d܀D����%�<�SQ�Ok�<y�G_�+�hU�-P�G��{�"�L�<9�I��
����(�4#�>�R��r�<7lB0|
 �A�T�zS��r�Z�<�TlO-&��+O��t��X�<�b�Z	�y���0L[$(Mk�<��'�*o�軓�Μf����r�~�<��E�&h����\�|S@3t��z�<1�Ѥd�R��ת�D�n�Hb�t�<�)˫���"v�Nr����l�<�0�B�h �M�ыÞ}�2����C�<����8$g��3��(���Y@�<��I}���j E�pZ����_f�<)�	A� r�Y	a�RF1�D$�f�<�"�A,?o
��C�Rv^Q�Պ`�<�)ə;V�����9��p��_�<9��� ��C�DՆK8��d�<1wGڊ&}05��E��(�(ã�I�<�3&T-/!PH���=k^��@ �F�<��+[3�L;!������L�<)%a�b8 1� �-rT��&�D�<Y��T�[`%`@�z���u�T}�<!�H�(AW^x�ǋ�xAؼS�D�<�&g�i먩[#ٶ.�D��z�<���4Eelٰ!n��<:"��ѣ�m�<�&�Ô2�Vm�g��fW����i�i�<Q��<'b*S�DM�8̺��Gz�<IS)Ч*��IF�Mx�����[�<AT�A�]��5���:=)
v��Y�<yF+߶
pb-(&�YL�-*�(^W�<�$��]���r7u�`�W*I�<���*"ڬ��	����95�n�<�Dڗ
�Ւ��7m��H�V��O�<N�+$$3��Q�SʒIhc��B�<)���
	.� T�9J@ֽ�wH|�<C�^�`�2�C�O����x��vx���'��][��I�_p�H`ŀ�I�F\��� ���9�b1��$�&^�h A"O`�`��C4"V��у�'Y��x�"O�(sr�[��(�Lּ!K�A��"O�u�e�����d�.5���"OPc	�c�-eި_�@5��"O
��Ġ��dP�z��[�ڡ�Q�'"1O�%Q����Qj�sq��M����W"OZ�ths��|s��O����"Ol���wZ���A�${��"O@P�� ��-��C��>iC��b"O��)��֔P.�� �C��%�!���T
Apa��A�I�D��n�!�dC6z���;eL��77�4�'b��F��}���a�셙o��!��n��54x�P�5D�(��R�1�9�Ӡ{�<��-?D����O�)�:��saTv�"�>D�tjsIֆ�j��p.Q
&-^��S�:D���"̭�\�YB���1vH��$.D��*�ҳYɺ��P ǿs�$���8D���E'�$��!1J_<&}���*D�d;P'�2켄�DK�$-�s�)D�tz@A7N�����$�:�g�"D�*�"�z�T��G�#N��8�� ,D�|����8�q�d�Ju��n.D�*��$1����%�eRm���&D���KI87m��'�X�@�Z�/D������G�uӀi�3�l���b D��R F��(ٹc�ˑI�xMy7�=D�4�D^lS�W�� `Tp���9��O~��I�$1He��8r�[��]8I��򄀹4Ă�����|�"!�Ң��yr/[���֣צ>)ބ�B�6�y2H+|_Ș·�*>x�
R��y�F��bdZ!₆Щ$r������yR/Gze<�� �S:Eh3c(��O�#~
G)�_~rAa�
|�~��D�b���0=qb��4�LĆT�XH�7�
G�<i�F����3����e4T�t��@�<�W��z*��ǍZ�daZ�C�}�<)�jEdX�I[�&�R���F�w�<��/�)\P�C���Q�А����W�<��
�S����)qe���I��NP�O�$)���C���0g}�Y�%��	3(��f"OR�P���V�lA�d�8s-���c"O
ݱ��K�7z�<�T�W G���d"O�e#�?�J�b�"� �tIB2"O:���-�O x�:1�W^��CS"O��W�T&�	Q�NW8����'�1O��,Q6�V�\���T#��Iu�O�2d$r7�ᚱ S?K8��
�'`���M�0���xA�,>�~��
�'�Z䁥M!k�`�[T���gJ,�:�'#Ta0��?A�!�ca�4]�`���'u6�R�G��]�>��#�]�\�b��'�� K���2ZJl	���@�^�R���*�'yAz�B���^�^�֡�12vE{��'e�4��E�zfz)���M��Y
�'%L�c4	P:;����È���V�a	�'�$�p��9s���ŭ,���'���#�8�BT`��:,�0z�'V�pa砋�E��}�C�t/j���'�X-��A�y�F�j�"٭[g�ϓ�Ot}�vk� �>5 ��ڋj�`��3"Oj��e�`�$�X�h�)�^�{�|�)�3� ��ڦ���녧Q��"O����N �;�<�фE(���J"OL�r�H�����P⒩6$>��"O�9�F)�-rN�EɆA��Og���g"O�A{�+E��I���TBp(S"O<�&�;�Z�� X'0`m�"O�!��5xj�8��F3Ј�W"O�e��0��	�Ӗ�`	"O&-8�J��m�\R���;j��ؙ�"OH�2�=U8��	�k�D"O��H�厷A�p�B�ܫO�4UA"O�ir'^�Gj^�g��[����}!�ݱ!�t �U\@0�g�7f!��D�.�z�ZB�fHހH�i�>8J!��]����A�W&<G�!�rɟ�L�!�W/c}�}!�$ -r��d�݄K�!�D�L�N�W����ӁЩ�!�$�5`;|0��h�$U��g
	��!���P0m3a��9lٸsn:�!�;p� @�cN�t-~$q�c�_�!�d�	/T� �
�b L���ɡ&!��J<��W(p�����U�&!�䁙`X��K�LɁH�4��R��[�!�䈺/�a+��D��P�b@�y!���lXr4J�A�,Rq�8�F]�h!�d�#�E�����``�a�TE�G`!��Õ\)�P�F��op�љ���E!��!\�Q��kVR��A��45�'vў�>qт`��v���g�2�8���d!D���Y!oo��g����lp��>D�K��*v��cX�p��q')D��5P�C�����Z�H�����"D�d�3��2U�p9�e�XA����!D����e�6gJ�)�5�&{�D��k D��a���� c�T�n���# D�@:�O���0I�N�_�Ԑ�F?D���G�9:��ɓ�@����G�/D�tY5�^*x��!�Ci��v_��B�9D��E�=�
�R��?���[%�8D��K���E��I[����> ��(D��*ʃ[�^���"s�ءK�"&D�Щ�a�.&T�T��S<��h�/)D���s�D�pɊ�q�(�7Tf�qU)D�����2-����#	E�s��(�n'D����L� &N�\����	 �<��0D�y��x?���2%Buq �1
$D�<������虢�
��cE�!�OX�	7|G���#�B5~yb�F@��C�I���	�F�X@Ԁc� J�jB�+/�T��O�t��D��$ܳ#�VB��.<r�ha��ۗGu����/4tC����r�&�������H�T�C�ɶH�|d��Hۻ�D�G[bC�Ɇ,l�i O�}�FLR���X���t��;��2�����s�T�#Ƨ,D�8�iR>[Pi�a�)u�"�u-*D�\q��W�=f��$��Dd�;D�P�Q�4pZ�)_ 5j�+b�;D� �e(�	o�~�Y6� 3amL=���9D�� K��>�t	�/�O.4I�7D��ҵG��wk�}�
X�+r�0Z�6D�$�DN��P8&akWl����A�8��O�����	>;������ih�D�/<!��C�cd�U�G�M�F�V٩Å�+�!�� ���u&V�v�j�UCR05"Of	��`�$q@��ҫ[�X�"O���&៖q���1U���*�!�"OL�1���i�` r�=ur�lj�"O=���(%t�٢���jJ@�Đ|��'LazҊI%?ʆ ���Q3Tؾ$S���y��P��5���E�S�d�S�֎�yrψ�dCH��uK�O�N@�rk�(�yrkS�"�q��#]�R�〬��y2m��*����b�_fI�f��yr"A%3��R��KR��B��
�yr����0���>F�)�\�y�HY}���� �<=��A#���yr��#:���Ѷ(#�IԎ���yB�4Y�8� K��$}BE�$ ��yr$�%@yv8�OH#29�����y"C�����s�L:-�H1�@���y�!�3�eQ��7%�>9�C��yB�O%'�h��sE�3�,j6BW�y�!�F��9Y�藢1���@G$ș�y�➶cD��U #D�`&�2�yr�I9�U��.$�=�$Ι��y2i�y)6�� a͖���1��Y��ybi�/<�v`��d5���2�ʔ�y�hR�)z>ds%�5QP����y"�ʓ�8д�1Y�0
�㕡�yLC�SݰUI��+�X��Bd]��y�/��Y%��C�cv�	[B �6�y��.���
��˦k[�u�A��y��Y�x�<*�EݧU��\�d˙�y��<yb"�)�̷<�l$���-�y2�؞�m��M%i変(!+R��y��U�GUZ ��'g��tX�o��y�ʇp�P���Y#`	0���y2J�<W�D��A5h�Z����y��-g=^�Re��^���#7H��yR,N�G��Qb(� +,�0FA��yRc�
P���O	'v��"�h�y���X�[��]�u�P<Q�n^��yb�1
��Y�v@�V�f��ѥȯ���hOq���2Sa�����r���'$�\�G"O���d�C�en�R6CƇ6n�"OL�C3*кvL����\�l!��`�"O�u)!B�����rwc�x��lq�"O�!I��8/�,��b�]��CF"O�Xveٷ�b��Q���+3"O��T;Ԯ%�T�L�$���s6"O2p���fz	X��\��&"O\e	��A�R@��
�.X�u�$"O,�QW�����7e�дp2"O�A��jؽ7v� 9���e�����"O$�#�^������+��qD"O0���
(9�L���dÔ8���1"O��b�N �B���"���X��"O�@% #�^����ʶV�*s"O�D�U�̧"-����D>4F�-�6"O
x�7GWlP�G]"h�e"O`�s��C�D[�F�-���G"O���❱MW��F�?�d �"O�1����A��EQ%�>1y~Esd"O6�-Ye��W"��[s�ȳ�"O��N������ŢK
���"O�|�tıJ�,))D+�sU,8�t"O
�:s��M2�|�v��-eLj�3�"O� T���6E��>�ti§"O(��צ*��[���-21�Њ5"O�Z��ʐ([t�p���;���Q"O��r�dFW����?�P��"O�,�CR�	QA-�3WNI U"O��ڢ.}����l�&J���S"O��b)8)^�sB�XO>qѱ"O��u��iNJ8Ҥ��+
���"O�u�AE�&��i��U�T����"O�Ԉ�C��t��A�`�"8q�Q�e"ORt�@��5*�@��2"��GL:`�"O��AA�H�Te�1(4�:I0�8�"O�)k5&7��A ���PTb!"O�QP�K2}DTt"v�=rp�"OFE*3��-0�m��f�"S`�@A&"O*�X&k�<�v5 ���-UJ��g"O29�F�O�{Nxt� 7?FyY%"O"u�73P��A��-��	A"O�i��@>lL4-�������"OTe�g�Ơ^TD f撁'�@y�E"O�z�B�#Oވ��Q�\�P�"O(H1	��d���e�*�
���"O*����Q+����,P���;�"O���1$4�9 êV�4
,�+`"OhU3b�Bg=`Q�Wj�	?���B�"Oj8��^Q�T����^��"O"�	@�, A �N=)G�l�"O���҅L�b�p��י=4y��"Op��P�TE�@ڥ�A?Q HMS�"O���!
B�^��X����-洉0"O",!���E�}
��D���r`"O�#7@V�l�f	�E�u�@i����
`�b>ej�CF�/-�]�l'�b�Z�&&D������;
"����A��Y�ظ�)D�VQ�d�mYq'1����D4�yr�Ph�pc�&Ӧ5wXyYF�	4�y#�!?���g�,*\@�����
�y�U�؈�����QX�%�����y�kF2d-0Yi��N���������$�\K�"|��'^�#�����J������u�<�p���(< �#G�E�Z�JSp��t�<�p�ؼA�j����Q
���*r�<ItS����c�솇i;|Y��B�l�<�G�3�l�A �C<��`a��7D�T��Q�)2e"�kW����)D��7.�Ĝ,3Q��V��|h��,D�\걆ך:��釩L�&ބ�1�)D�(�`�Q9z ���Dǋ�\r`�ů*D�,���ʿJ����� ,X|�w�)D��*�+`��u٣B��Z8�w�=D���dG��HY�����(.8��G�:D��c��;4��QIRN<!�p@2�8D��Z��\^�0���<!��A{"�8D�\�O�3��)���v�I�/1D�����͍c#*	wL��%m`�	�G/D�� W�M���qjbF,���h?D��i�aW9\�����F!v��R�H<D����N��A���G���x�R)>D�����HR��0d�(�|��Q�9D���b)�b1~����V�[�3B�<D�4�7,��
Y��x�K��䤀�<D���"/[*�ND:�N�5)� ��8D�`;2�!stIc�V�%Z��P�5D�Й���\��YrvI��Rdh�5D�!�� j���h��y+8ڷ�̱J�*�4"O��ueĵ������]�1����T"O��G�Ѹ �|tA�JO�����"Ox�SW��(y�[� �ehp�YF"O.�b`��	�Z�V�`XZŲ�"O�$#X��ay��_�2;t���"O�Ux��5%�J�Ia��"#%T�@"Opإ��bs�U�D"*�B�"O@���JE���a���s&��[@"OZ0��͐�c��e���z3�9��"O��!Ak��m�2�!�	J-���g"O�����P��8r�βq�$Y�d"O��[��]r�k%a�;�R�Sv"O~K7.(Dʢ����S=�"M)"OF|����7D3v%#�@(d��Y�"O2(�c�( �)�e�+M�`a"O��%o�4X,$c��
�(1�"O���͍ZLR��f,�b�Hx�"OiQU��;M��KT,� |���""O���M�.	rV�rb+�&Sy�m�c"O������.nj���ɞ�_`�tq�"O���chӚuZ9�2"�<n��9��"O���Ei�����[�t\��"O�Ъ�FM:� �h�1x�9p"O�8I�I�����1�.ukB��"OV%(,��\����:eil)�B"O�����=f��xa��MgD��S"O(-��O	V�EbT��Rg�ti�"O\��$K�_�$-�$�#Y4-9$"OBu1�� ��'@�S`��Ѓ"O6]8�ýR{n�a爂�E�u�w"Oj(���#:�����V#Y;��PA"O}pG,ҟ ��a4e�'"�5��"O����ę�:^X�s�ጜ7	RQ�"O�X���I5�d7�J�ޭ§"OVl��#�0��]�4�	���`�"Oj �%o̵.������%L�����"O4���ۖӀu�ql�ty�Ț�"O<�w��-��\�@�ޫ�p ��"O����5~XQw�]�z}�j�"O��[��?�:<��I�3Tڈ�۠"O�$�B�ܯbMD���H�$%���"O�y�t���B��=��W.0	�hX�"O�Q�A��;R*��a�%�j�ya"O<ř�bفQV�;"!8��J"O�ɐbҋ*�Β�I�� �"ObPRK�8%.��TGѪ|&Nm�"Od4��"AliZIaP� l�(�"Oވ��%� * wD�5tUs"Ob<�%�u�>�C�#�,�$CW"O�����}������ٿO�F5�B"OzE�P`NNG���!�ʭ%�*�J7"O�aC��
#��{�ϓ6���'"O\�ʷ*����W�fT�"O��p� ��p����[�ȁH%"O�������� 0��E J�A�"O\�6G�0#8Y��!^>��1�3"O
x) @
<
p��ef@c�0��"O*�1dB	 
�������/E�e��"OB��̖�$�&x��M���	�"OjeD��!x0�4
F���Ҥ"O.A�!�'�4�d�b�(�"O|T	/�.[Rت�6'#T-r�"O�T��ܫ�((%M��\G"O� �Q�&�D	!�ph36�ؕJyle�W"Ol D@L�J�"ܫ�+�#DwF�� "O��QA��4$�pF(��8a�]��"O���E$�(y����yD���"O^�#2ထ]#����EI��6��C"O�L;�+΀=DE�d�jx���Q"OԌ� ��;FzD0#Dx�)cr"O,Y٠��;�VŸU`C�(��b"O��20`@b�x1*��N���C"O�P���s4��#�qh&�0"Oz���L,[�!@Ԭ�(Pa���"O��`KX8]�0��B��"LO	��"O�t8R.Y�� �`����I;x]��"O8���"-c"|�7ƅ!Q?z�(`"O�'�Z<8�21�Yc$"O��u��g�Z��3�W<k�ИI�"O��H��^����1���HPh�"O��	�����7�D�*�y�G"Ov����P;2����aG�+M2="q"O�4�e�Bn8q��K��3މAQ"OD()�G�J���3�+-.�9ZS"O�H����/�fy �	-F�N���"O� iР�u�$�k�KN�Nq�V"O����U�%|�9y�Ǻc�6���"O:Eb���3B�r'ʳ縭��"Oz��(\�mqfE�E���:�"Ox̰���k+���E�vȌ] �"O�X��Ey�H�a%
رS�P���"O>�`�X�<�����)I�.�� ��"O2-�
�;����p��y�"O����Q�4��+�K.~İ�"OjU�N�z(;�i�,j�"O�ق% %Px�L`P�Ŋ#�$��"O�=��"K�kn`�3��V��K"O	䠝�<Z4h�I/����"O�qXr�!
ȥA��
0l��"O:�s��� �,=� �޽XuH]�f"O�`5�^�!NR��U�ZxW�t��"O�`��G3�@"s��kP ��"O�aH�o�+U���A�H[�l]~eiu"O����ǃ�S� ���/!;ƙ0�"O������(\�H!#u�$-��B"O�!4@/i�� x���<d���"O�4s�ƧWyh5Z���7�>H�"Oʅ3�۔L�DY[u�J'hĻR"O�|�h��Du3f���p�r"O��Y ���Y�5��G��P "On��n��B>|��i�v�8lA�"O2e�fL�e]l!�d煈t'�p�"O����%1���f�[�Ҥ��"O&����2)4 B�e܂����"O�X�u��&2>D�cd��vL���"OD�3��Պ�ڭ��b��Q��`XT"OP9rE�Ծ1$|-ȶ��5����"O� @��F�t�H�&�,ytBUأ"OL���b��J�Z�"���C��!�$M�'I
�[!���e�`�s�E��V;!�۸V�&ȫ��;
��P���!򤏿?�8�ڲ�^�"��s���P!�DT�r@��O������g��wf!�dV�8^4�8p�0K�X��g /3�!�D\x�`��MU!Y�G�!�$DC�rD�Dk�#�� ���D�!�ė	j��Pc�a�<�����"A�!�� ]�U��D�r�It�׏N��U"A"O��Ђ��	f��hC��E�>����"O
�R�ޜ6VdS�-�_�~Չt"O���b˂%x�;�,�K��e)�"O^�Y�� h$\A4J�2K{�Q�#"O4$:u��!Q� Y���t[�D�5"ON�9g��:��x�-�(H���"O���ӠM�=���R��ߗVC�kF"O �x������u��甲4'��"O񣔤�c)(�p�� �<��"O������8d�\c`ú~�S�"OJ� $��b-�5�T%rrI+"OV�*b�����!Ꝑu̎�y�"O)���`%�лI	
D���"O(������H�j��@/,���"OtA�@ �6f�n�����pp�"O����ЬF�T�����U�0p"O`��%��[(���a��,�B�("O���ӌJ&j��DYPaj�he��"O*��E�]�Ǹ��bT�d@���w"Op��DFWp4@I3�ÁY�U d"O�IR6ő�c+�0Q�͌,lSZ�@"O��Z��;���F/ �:1�p"O&��􈄰��H�T�j�~�+q"O���v��+$��hC&�	ۈi@4"O:���,��HJ��W":�=˥"O��ڐO�o�49Z����0��"O�l�u�I5aRl�:Ď��F"O,t�E$-Bj��읗  ��2"O^�W�?	��D�V	le#�"Oj=����
(BL���a�� ��؊�"O*@���=�h:#G�%���2�"O�h4lA��ܐS���!>t 8�"O0a�U�N����5��?B �e"O�ez�a�'1�=���\	�� ��"O��1!Om_H��O��ᩅ"O�p����W�rx�Q�߉X����"O�3�
��"���r��Q:܍�C"O�!��P���쩥h�x)$䒇"Or)X�M�HϞ0�FL,u��ɓ�"O�8R`�ڼ���;L���Q{G"O�!��`�*��1#!ۦ�h}J�"O�,"WA�E��"�@�y1�xzS"O�
A�8� �-(�`�p"O�mR�$ŗj�8d��oЮ 7�q"�"O�Ea���a�`͂��SC6�1�"Ol�E�NDU�+��KR"O����A�WB�:uQrY<�j "O�����{.F�	e�� C�ۗ"O��V큁w?6�S"hUq6Vq��"O�� �B]	,�Ԁ�S�A?S�f\1�"O��@�_*�
�� �H'NW�e��"O���	-�.qHͯv@��"Oi8��ш @� FM[�(D��"OL�I0G��7������0h ��"Oj�*�M׍�.%���Va1���q"O���((��}b�V�D�V 9��2D��S&�^Z
	�Ц�m^ ��2c6D�\1FoA5%tZ�k�փc0Hd8r%!D�X�P�C-X��@LP�kt�I#T�>D�9D$�2(����3G�1���!D����$2nŻ�NA�8ۀ�>D�����]梡�D�^�����J/D������xa6f��:��F� D�� ��D�߄_@d��ynP��S"O��d��'"�ĠRl-rO�P�"O����V;yd��`�K�UF��"O���C�PMP�퀱G����d�g�<YVF�3��]+E��THgo~�<aF&V+A�����VQ.�;g �e�<a霛v:�RӆΪI�̌�u��b�<� �-b��Yt�����Ð`�<����.P/)�v̭T΢D��]�<�A)D�GЦh���,/���C']�<i��¾Y�jC+ў5��Uk0c�<Y�F�4��$��͝[u΍e��H�<�w�� *�ޝPpMV z�d�w�FC�<!6�Q�8� ȲQ�B�2Q�T`��<��L!!x�&LSb�JDB|�<iDӴP�d��i�
6�a�"U�<I1b�GK���E�=+��y�<�4�C�PŒp@rN��m��=�w��q�<A �|��|��f
�W��顦p�<�$ǂ~3^�H��!r��'͘w�<	6,F�,�z��GN��5W}�<Y��W�ֲ�A�)L:v���	�@�<�'��8��h9��:(��x��{�<�!�P�zl�!@+J_:eh$��v�<� K�
��	p�����Qek�u�<�@��S�	ʅ����FV�<��Z�Xu+��>&�9ӑ�i�<Y�b�N3f���Eӷnp���\c�<Ѳ��&n���S�K�s�^Q0���]�<�!�ņLzY���b��:E��[�<1��1V>��`�X�JCЧU:~�!�.`f� �;R,��g�N!�ˀbA|��w�1P@����/W!�U
�Y*&�Z;m09�夕�	�!���O����T�pLA0�� q�!�d�G��,�f�υ%�,pNP�j1!��W�*M`"�0 "�l�L�R"!�Ĕ('ఐ�KгO����2!�Dݓ�&)��J���D�L5l!�$Q�����RNF�&;�}���4�!��B5�!Ϫ`�l�l��s�!�����K ���͉����}�!�I�'Ul����@��:�Y��!��Sy��Q�"M�B-R�P4�!�$Z�Y8ht�f���(ph��g�ΨK�!�d�)Q���5�:SUdɱ�J�)~�!��}y�-��Z)9ڌS�U
:q!��?�z�acM�5\��
+k!���Ҡ�Я6�����S1�4�+�'z�Tp�Ѫ>kΝ�`��/"�	�'h��F!1��X0��'��<��'�lQ� F�x�Ⰰ�"� �j�'UR�+��̼\��a�Jٍ0t{�'����r��6S�i�E.�)�Y�'늈�ǯ��P�lŁuiJҶ��
�'���hl�y�TZB%֫3c��
�'��X��Ӊ���z�葍U4<��'��R�rI ��R.T�f��'f0�;��ƶAB���m�Q����'=|ݚf�&{�ȨQAقA-"��'XM���=�hi�bV�f��= �'�,zG�q�Ȕ�ï�q�N�#�'��X@�I
�*D��㣒�f5D(��'����dK�/�
��o�>X$x]���� �9cAW�Sj�T����{0�Q�"O|��d��D�D]�
ГG��I1"OP�2��S��KH��V$r"O~�!u启3�p�gǒ4	ޠ�"O�az��Ş/B�% V�e���`"OdL�Q�ԲDP��!ʵ1��}:2"O>x������@����w�9�"O@!���Դ��L�֪J����"O*��1Y�4�6|H�Xh�t(1�"O&D�	˔Z�S��8���"O~���'�b�� ����$"�$�G"Op�K�$��� s�h	-lX��c�"O�]�vi+9:p��F�>w7
���"O(�F��`s�-�3Ô
	%tpp"Ob�(��ɣZt�RQ�ɆEi:��"Ozh8���;s�M�a	�#)2@���"OV�(#�_���x�G(���0P"O��WKN�Hn,}!�N/6r�"O���&�o�
����I����"O^�[jN'T�҄�09�ൡv"O`�9R+Z�2D�f�	 S@�t��"O���l��/r��M�<F%����"O){�� 	��k�d t"O��PO3���I������"O@�e���a��My���9U��Tq�"O��x� 4&��)@ݸ=xA"ODL��,X�]c�`�3�ЅD�콘�"O䠃g'Q�"Y��Y��(��"O"�M�/$�>T��H)u�"p�&"O����݃'��l���ħY�ȀP"O�	C4�rO�U���-v�4d�"O�ԡ�g7�ڠA�V's�>�h�"O�y[�k��AB0@j��]�#�
��C"Ol	�����`�I$P�j ��"O���Y�+�JZE�J5T�6�g"O@��&�p�����(��ᣲ"O͘�Ì$}�y��gE:T��Y�"Ot(�'�	v�ε�a��l��8��"O�TJ
�����u�H�C���Y�"O�Iʄ�D�#��P�@j�;
"X�&"O�s���x��y9E�)�b���"O��3���iel��C�cp䜑P"O �js�*��y�,� U�=�"O@�6�=}}�X9s��<JVI�3"OP�Qf��DnX�`#l�>����4"O�i��,Y��H׷W�f��S"O�T�m�,1��h���B"Of���e�}x����݈Np����"O�Ik�cE�e�6�3U cq,;�"O�[@��'1\�R@D�Uchl�Q"O,��ԫR�$�\ɰ��)HJ�Q"O�aREY4X�\����ߍ78PK�"O(��)��96�I��_6?ֆ-�Q"O^�sw�0Y����(kǆ|�"O,�{c�0=�r̩2A�@�t�Ђ"O��ㆢU9��0����3J��e"O��Ð>Uj����.HD"OV1ည#<�� =j6HȔ"O ����x�hT�#o��v����"O�0�#�b_p
 �0J�(��"O���`�%UM�0`S��"��L�"O�`�Ƨ��x�V�^&5Ӹ��B"O&T��X���1b�-,⌈�"OEJ��+��P+w�"pI���$"O� F���ǌ�D�64��0_*�$ �"OTy+7�P G��9��n߳<j�"O��P�R%5F�5�q����m
"O��;���l�d�Ӏ��i0.0"O� �Հf����S�`�f�A"O��bUcQ�S׸��$�CN����"O��Ѳ�� P� Qz���ib�x�s"OnD�t#;��1��̮xY`�"O�  M&Z`p`3��<X,�s"OJ<�B*X�34*0P��8?>��"O*$[7蛭ye4D�6(N����0"O(���$۔f�xx@І΍Fi�(��"O6e�߆$laH��ܪPֵ9�"O]��j_E���E�*d1R	�"Od	���Ť�HEQ�ā�}�hAD"OT첔��Yc����Q�p��:"O�=�m�#U"�h�BϫP|��I"Or�2���]�5�$Ǜ9lv�;�"O�`�eF���Cm��e� A�"O�Q�_�\84M�)up�"O��40�źQ���s��\��"O���3K�R3D�@N F��"O���
�>=���7���w��9�5"Oڤ
��pĒ&8?�d���"Oj`0��O"X��c��w��*�"O���V��d�:��T�I�;p=21"O|�yQf���V\��g��+PR$��"Oʑ"�@�,�vѠ0AF3���"O�p��9��FY�Tz����"Oޕ�6��p��m �Νlt\���"O�X��V�{�hd�A˜no��k�"OT,��g�r���	���d>q��"O��@�Խb����AçJ$���"Ov��6e��͂X�FU@�@܉a"O�$X"iͯ;(�|B�G^Z�X�"O�1�e�2Y���*,����"O�|�wB(:�"��g��D�"O 5�ǧ�7`Oz�{6+�t���	�"OP��n��|����i����ȓw"O��3)ʷ8�^h�h "I}�:�"OBY�#�:p��%��>2��#"O�A��m�8~F�ź��Ŗo��աp"Ot�z�"�$���c�d�RM��"O�Uf5o85��)2{��j"O ��E�}�fiQ8\R� �"O���fJA�aAzܡ��E=P%�K7"O��#�A{Q<���G�U�Vmy�"OR�{u�+~FRiZp�Z��W"O"!�2�Z�Q�� z d�0���Ѣ"O�z2�ԣK*���A�`�Cu"Or�3��љHrD��%�n��2�"O4T
"J�	fnfQc��Z�r����A"O�� �߯��1�d��>h� "O������i<Lɴ�۶8�8��"OL���f^��(�ҁ L�҇"O��5�Ė�neӆ!�	AO��"Od͐�$�O����jլ`.L���"O�e���B��гj�"v��T1'"Ox�$�G���a���Q���"O*��׀<9���.�/p ��"Oڵp�G"m܎x��c2��y��"O�XX�HҧP���B%�9ؐ�X�"OB��sC�'G2�1��	�@ў<��"Ox+0�Z)[J�4� ��>Î�0"O� �`Q���%WN)�#���C�J�s�"O��{�����4	&d_1 z���8O�2�	�gM�){R��>���T�I%\J5�"��"=<,��v�M�t�B�	;(.�`]x)�(׽w���"O�u�w/Z�~��EK4���xcRL��"O�4�뗓4Nj%�"��fv�[3"O`�!	# ��?7h��"OF+a�O�u�D���$�XE"O��z�R�[������Y�Z��I"O�9ZA�(U�H����Q!&�(�2d"O#��I!g.�Ҋ�$���"O���V��.;dܥj#(�0D����F"O<���`U�!.x)�`&�e��I�"O�e�u�/q8BC���R.�c"O����Ꭿ���˥#S���)Ѓ"Of�����)�~5�B�G�$pP�"O>���cŠMf��` ��JTJ�"O���%�g0�3ƅǙ]��QP"O���M�{~��J�d�<�$���"O00pq/M p�8�0`�.�����"OٱP��N �B+�f���D"Otd�g�Y+ �X��` W��TI�"O��$K?U�����I+\����"O�xr��q��2��`q�1s�"O(����`xR�����"3ݲ����'yP𩦏����I<�M3��A�_~��{���>��C����D&ǈt}\�I6H��E��O��0��/�NA��S#5�\0��՗P{�P���eK�C䉀LBb��o�8�8�#��.�dDl~JG�n�E�}&�P��ŗ�J}�r�I��J���-�X��HŤa�@)�թ�m�w
5P�P"�*�QWR��	�~$���7>ӊ��V��nD�)E�`�E��hc�Z�8�Y�O��0����s��y�t����d)�'���c4���{4Jݲz^�	.OvT��P�p��Uq��ئg�Q?������Ҵ� �M�;�ԍ��2D��KQ>!�X��L�ww��B�됒��3R��\@�(b��g�'��Pz��*��q���\�8��
�� a����I��u�G�ۙZTt���J^��lS�ey릱�5�G*�p>i"�ru��z��_�hM6�k�(d�'��PBB΂�qs��"ge�*nF$�[�h�?���Äjj�ه�A,1}�]X�-3D���p�	����Wl�U����N8S�(!J���}2�Q�k(┋P�sމBO�=���fW6٢'�1D��g"����0��� �D�ĥ�{/>\��K�G�:�H�m��GS��	C�	�Q�$S�`C����B�^�,��٥i-|O�9�"X��U �b�j�ƽS��!��D_�Is������(C�n�%�'�>����&�PK���M*�@ی�Ʌ�k��Mru)F'K1�i�f���H�X`��O�@� �B˹f�����'Lێ���'��!�����H���5:c���t�P�v��L� �Cfa��f�O�����9�N0,u��@`�ITP*f"OVM��� R$D�R��@Pb���T&T�p�� �(�0�r���6�VI
�	�(O��+U��)�5��hK�ء��'Lv(�C�ӵs����sO��b�n �@Y�U8v9Cae�1��Q6��6��j�#7�O֜�sL�6��}�mӐs�81Se�$ȸA���RdF�dM��1�Z�h����	j���7��� '�1>ʐ95ÖX�<�Aa��8�1�V(]РȪ@ʘ�0i��I��t��խ˯�!�N!��9*e�.L�})�@�U�C3�����
n!���w��{��V�E�4bG��*z�W��b�t���1%}��灋u�
�#��$��Ր�8�P��ӖR���	;L*ͣt�xt�m�eN�"��<33���D0��_ad�]iB�α0�`�H	�ў,�e��
GKUh��]�]�=aҧA�*�T�F.-Z$b�H�2%x����`�	#.Ti9�4;��I^�tUz�"O`���N���Ф�1�j$x���iY8�q��8	K&�+�mF:d#|B� g�Ŋd���wb�lb�d>��pYA�)D�,��S,#�:���PEV����.�?�2��HC0iN )hE�h�J��͈O� %�tċ�!|��s�բNV��j�'(V=��ݯU1�D�σ����Q�_/ (��",��48p��9�p?�3n^٠!�@J�,��ibV�I]�'ά1���! ��M��iЎod�U���X�D�Mc�I
Mn!�$�<��q�6	�ǐ�7*Ѽ���3ϝ7i�t�RH<E��co��a	�4�����?@�T̄ȓC�F=" b�^�d���k��l��+І��3�	"�NY"�&�%�U��͚�PV��wx��LL��ȓyy��^�qN�˓�0}��Ͷ�`�&�'d�ȑ���AEv`�ȓJ��I���@���!C4-cr��ȓ����d^�f
�\2��1}���ȓtx��sS���a
ء0�ųv"x��5L�Q� ��)�̉+ʪ}��7�F؃��dM ̣�Ů<����ȓn���B��N�J%G��Bu�`�ȓJ5t`{�)�{�h�P�#�<)��?Аp8"�!�H�m5>r�ȅȓKg�� /mYj٫���t)!�ȓHyL��"���H�.�'��tU���I�0p��G�3#N`� �fp:P�� 5ʽpbbD"'o~(�i�=b����Oj�3�K�?H�@� &;���ȓk�PM�u�BX�� � `v	���<�b��%{D��A�C��y���� �`9cB�4�l��@G���a�ȓ8�,�X�%�%mAԽ��O(-���ȓU�*%Cbf�`����!�!�T�ȓ�(�p!#٦
���8��V~I85�ȓsP�ł�I����"��-��|Hh��`�v�pJ���,o�������i�72J,:��/!JU�ȓ�栈�#Q!��Щ�a�%f> �ȓm��0��'	�c�:���6h@ܱ��h�~��-N7S504�È��:���ȓT%>l��@�xH֌�V�Lv�@��ȓc΄���7����P�u:���f�`��+��vRjEC�)a���ȓ&fND	V�U��<$
�	C�M+�ԄȓQ�4UIM�0`�����>���ȓT�ƴ"G"ݡRc��K���(�}�ȓ>��;�h .�̡�h�&����_M�G��u\�4n�=s�]��K��s���M�� D 	5b����ȓ:JR���X<K_�Fg�,|�Շ���' L6}@�գӬ��(��ȓV\�#AD��Nᴨ�t�x���t(UA�&҇h*��8��Q=z�<��a^�;�F_����H�8J&`�ȓ[MDq 怼mH�*� C�M&���Wf��pB*B0Q ��
�+@�g����33���C*j�t˵�V�>ن�+\�o�9�h�Rs��[JC�I?|Bvm��/ԝf�$��ī|p(C䉨1�@��C/2�Ԝ���h^�B䉱g����(,�!��N��B��U`��4�͚;i�A��44H�B�ɩcn�0"#���������B�>W>@)81c��|F�@��$*�B�ɜ[M�B�L �gv��E��� b B�	`��ѱcǆ(� )�¢��/w�B�I�L��@��	/�8 ��w!�B�I>2K��"b��#��ăd��5��C�)� P� �)�0�����o�-�.�ja"O���k����S�R�����R P���Y-#�ؼR�&� |�rݚu����!��=-��bDyƜl�s�+l ���B�*)G�W�D�|�',6@��
鈠�eO�N4��	�'�$B�&ʟ��U
]%+=�����%m��ɡ���P��Q��/h(�S$D˲��"5�E^���ddHZ�Z
"���%��6@����*$��T����V� �ȓ5RvȪ�%x��qh�-j4�`&�$�c�-X�f$�Ԇ�[��D�t��=�&��r�P��(�(���y�78�t��c�@��D���;�A�H��I0&(�	K B���L>i��',3��U۬a	,l�DK(<�LӒ\��Ms��?P� m��f�#|x9��n�6�j�C%Ȑ�Jh���ۋ<����P!o���h�H�+_ax�F�E�YkDυ�@�L)��M�Y���R�P�C���C#�[�u�Nyx7O��)V��A `�b��H��[p�� �e����yv`�1̚e�rhB�'q�iy@��~[� ѥ�~�b�ȓl�}�,F�K�<�B�,D�u�����v��TO,$�ڵy4.�U̧��J������=9����a�?B��d���J���B�� (g��k�OW�>��s1�|���`�0Xx��+�z}����	�B�X�S�&S�Ws@�
�]+FP��D\�4�D�ʳ�;1�B��h�\/`u���� ��YpR��ފ��'64�H���_5	�I[e��1���P�#?��J^hk^9#� ӄUd�������O���нXh���܁V���`A�<�`N�9
FF̊u��$	d(���� ����d�[��A� ���-�|JJ>q�ID�xs���')ɟ9���X��CC(<�����I��2��ES!�֙ZJ=j5���I��{ï6eb����0LO�Ic��>Cx�I�h���Qf�'���]�m���q7�ټl�\�GC�<� 
K����i�+�{�<i�!a�:lC�e�(&����Yq�PHѓ��3a+6�B`�G�O`$����H� 1�O&�I��'%�#�N���kd�����<w��� ���Q!����ē_��YunR1q9Q3%f���#�:I�t��O!�	�Wi���İ��S�K� ��T[z�d�������#''Y�t�" ����zR�ɖ&ްX�.�<a��~-�j�eq���7(T��[4ʋ�z�Zd�Ѝ(����n-�ɷ}ܩ���Ӗm),��ӴH	�����
_1xC䉯#x-�դ��yDbaQ��2"fB�F�6�s�� �7$X �@^8�"B�	ZeހZ7�N�Kr8��O�<B�4"Pl���:6b|��.@�C�I�� CS�F��Ll9��5�C�ɵ�,��N(�h�Rޜ��C�ɦ.@��''�<�P%�	pxC�	H��h#�K�/c���a��%"s|C��v�0�l�_��v�� ��C�)�ʤ;�L��qe�	"kb&B�I,�4�⫟4s: ��D�DXB��\\ ��k��'�� ���P�NB�>n\~�p �i{��rV �	lT0B�	�l�Z�H�#V�
� j�\�4B��$Me������1~���p�o�"3��C�4F&�`2�`���x9D-܈��C�I�R�<1���N��0���k|}���'b����&Z"��A$�^�i��)�'�8�#�$�L�n�R��A�I��5�'��H�U�y"H�8�*�Nd\@�
�'���bAH:T)�9��ñEd��	�'3-�ph@� �J�h���1�'i�(��@L�9@�ۋXa"���'%t�(FP�[����T���Y��'\�Ѻ��P�T�d9�S��${��5x�'�Bm"$�d:�$�L��tV`:
��� r���ܵ��RӎM�e؜��"O|��h_2Q����( ��5s$"O��	Y!KV��c�h��- "OTI��`��I.��B� @����A"O�a�-�k��x��[�It�41D"O�
�'ʤJ�8�Zs/�k^��F"OF���1^��r1��=@��"OB12��E�_:.�A���7:����"O�8!�B�<Q�U�K[�l&p��"O���ۏTR>���Ӡ	���Q"O���#�UM��Q[g���zP��"OJ({2㗌E�0�6&V�
.�y�ϛ7�` ��,fK�B�y�� �2�y��������һ�y"@�&i��i
�Z��8J���y�+:�DiRS�U�T��1H�N�y�Ə;t�!�MO@[��so�=�yB@�T֠L\&Kk���E$�y�.�.>���e̮Mx|��.��y�A�'М���`	�:�
HPG��!�y��Mb��%�P�>��(�l��y�6(o�A"�i�8�sv���y��%Z����O��>K`0�ef݃�y(�|��H5B[2�R��,�3�y�}=����Ҭ~2aY7�+�yR��Y_@��MϩFH�b�Ѝ�yBC�)=6IK�&�H��%Xt�K�y�A;X����}���@����yB'M�8|p���'[� �pV�Z!��<y��'Z�"��O� 9!a]��x�:�!3��(�W"O>���Ōd+X���	,p�N=Hf�x���Z��b��.�|�V�E�w���"��t� }�"O�)R�cL�a��`!��o�r�s��#G8��!���(�3���] Z(d@V�W���a��*4o!��_�IP��2.�ia��rJm�V�\�f���VX���G{c��JS(G&g���+�J,��|7�qV
#��i22��j���73�9jB��Z��Ԡ�M�W�<92&�!~�6��1O^�Hq �Ly�˚�=�(UPBD�D4��A���
�b��!	 ×&1�R\��O�f!��N�'l�%"ժ乐L?L*��� F1[�(Rq-���ītR>�<)���2d�T��*H@��a3�EX��	���>	��!��T57���9�f\�l�Vm�zDTi��J0i�m��	V�ِr�-K`Ŧ*츣<��[	U����ϑ"0��E�(���I.�qSBC�)��Taua�Zm!�dS�0� �@��+~�Mȴ<[29�새C�ăZ=��.�`D��w�<��
ʕ"�~�q�B{��	��'Q4�dh'p\�q�@'s�Jl��%��I�v`z��D�3�Tz����T�f�'�*9�2G�	q��ya��
�m�>�@ߓ6���6���1�<�R���u�F!tf�ҷ�֩=����\�
An�a�'WtȐ�I�| v�j�۫I��j�)�=C��@��~��%��5S�6��O�R̳����j��L�'Zf�\:�'�J���l�?�hqfMًRx���eo*ǜ�ch��`ي�PUg�\�B����;�U*�X?URj1@eD�j�b��"O�Yb��ͦ"SVjŤ�/��̰��'s��`z�#QC���2��<��]z�
��(O��D�+�8ӕN�0]o�m�0�'�r���sV8��Y�72
����P|q�܍!E"��C��Y��(�O Y���/-��1Y��6�(Hs��If����	9(�`U�5m	/킐i&�S�4 QT�+6�]�	L�|�2�PV�<q	̋�7�����ڞ^���H�i� �dC��z´ى��Ld��b?A{�3�ٲab�OIE�儉{�ə�"O�Hq��͌3��ٙ��W-I��q��a)��hSn_N0f��tO�R�@Q���(O�� P�A>�*)�A�ĐLV�K��'HdH�D� S�HիB��A�M�ɷn�F�	TCZ3`��S� ��u��d�fM4�O��4KO8-�앪�ǝ��֙���d�P��m
� &\q�I9O��=�zm���~� `���b��ZT$�x㑰�4��"OD�w�V-4�8IA��:��(�&���~�
����WGL���L�jE@#|Z�h��s��vk�h8��.ڦ�K  8D�H9 L�=-�d�3��Ažxc������b���;�)4l�6D�&���O�]۔$İ#�H���ᖡGDb���'h	R$��Z~�I�����H��'n�8?W��DFnn �����p?�G*W�DIh��:\�<�p�OFx�',��('T'�^����ɗV��-Rd��P{��0��n?!�d�(Tw��D-��F}鑦B1 �f�JU��L�6UI<E��FX�d��釽'�z�c��b��Ԇ�1a$01  !�(��o�pT<h�� �����Uc�I���y(��1�.!��{ D[���-�����:L"P�ѥY�p}[��Po4���ȓ5��-�Q._�2i��MH�kE�M�ȓ��b�FK!M�dE��H=�0��[�C6��,lm�C#J�&�hd��V�r�d��_�$y�Ҥ�M�L��ȓO! ��B��t��j'[3e���S�:9��/�&$ԅ��tO�m��Z��[���
�W&L���0D�$(d��K�¬:�I'�8��tc.D�LP �A8
�&���ȅ,)DܻqG,D���0�Վ9	���"h�Ь*D�26��(�a�v�$aO2�f,D�t����W|tD+a�Y t��;SB(D��z�V&�8��wBU�.8��d�3D��(WB�8�FT�SJ(��͹%.D�����~���&�h�"����0D�:a%;w��|	֬�LS$4�$J/D�x
R�0����
�����IcbC�		k_$]`��ܼ+�k���6C剋=P.��ǋ��>k�����!򄏑*�t����+2nٺX)�ࠇ�B|{�������?}����ȓ434�;v�+�|0���y�虆�X�*�[�&��~!�)��^�Q�ćȓh��p"/�z^�҅O�<ל͇�j����W� ��j��=Jn��ȓ��ѳ�N� �>�!"�VXr%�ȓ7?j0�2Fؿ/��XrB��q��[�	H�ܷ%�H$�\>% ��ȓH�@1���:�j�;G��4>��,��gܜ���k��˕ŏ>:H�<�ȓH�`�p��V.}~� 3G�"�-�ȓZ��:�'�/i/B�k��*!֒��ȓk&�I�שQ�u����s��:�L��ȓ����@/�ڠ���O�����ȓ7��D��(��A{�F�"Z�h�ȓH#@D(�� )N(��X�����ȓ`Ĭ�`�4@>��bݗtF`t�ȓP.:*�/�2i]��i�LM�X��^�q{��}CH	�s���Y�����YJ�eeā+�|4���7=�����|��i葥E9jrѻ���1`bv��ȓ.f`t#�jN��b��a�A�8AV���cH~�)�I]�+�4�@)�O����Qf(�j�9�Ȁ��CMOt-�ȓ��)�cŊ5lh��s6�
�c�Tx�ȓfo�(���;e|��%�v����U�*�󓏋�[>uۅ�
�8& A��{��yÅ�S0��ǥy��ȓ8v�� OK��~d�`'��P�X���i`�V��_)�)����i�����S�? �M�� ��I��`�g�P�d-Щ	�"OT���̢Z��ĸ C�6���"OИ"��E�	����磗6L]�9��"Od-&K^�L�� 0�kA@P��"O&���P4I�dA���:;��T;""O|E����;`4���\+�H���"O� ����8u��<8�M�z�x��"O����պ:�F$@e%Z `���"O8��r�њ�~pA�N�O����"O��bVe�#i����Ղ�5�$XF"OJęC� �6���H������4"Ov�@��O�1�[#��1�"OM"d ��/��:��
�w �k"O�:5$�=���3 ^=KGP-"O %�rJ�p�4����T�QK"}��"O*	s��(؜����w7&���"O.<� �9K�hZC�Z�>&t�w"Os�-��c��MXT�@�t�r�"O�|:w$N)
t������dRm�"O���G�$md*��g�ܙ�"O�(�-��Jw����f�k�
]��"O8�!�O� Q� ��ƝNp@)5"O�[$�չc�Eb�G��pX{`"O�):
��ܙ`t���0��|��"O��r��]Oi�i�w�
�� �Ƀ"O�] %j%?���ք��c�,E	�"O"+�� �vZVhcUȚUr�p"O*��� �f����O�B�Q`�"O��Y�#W�8��su��3����"O�z���v?�`�re�b=���"OZ�F��$`�t����` �:W"O��s���5)�2��@�Ch��c"O 5�a���9�,8�P�V�v~��1@"Oq
�ڥa������]�%J<�R"OFH�4#�Zm�D���x���1s"O�uf�һ3N�聠0;��{�"O<Ԋ�Ć�h��u�2f��	�"Oz�ӂk��M��5�RװYq ��"O@4bL=<8,�2�,�D���"O�uK�ýN>� &�Lmb���"O�3�6_MX�#ӊL	���Z�"O�A�َ$��Q��S�q�B�*�"Of=�q�Yq�"[� Pq"O��z�GJ�q�j�3b�$��"O$d���N�LDRT ���kꜽPr"Ot��OΘ@�n��Џ"�r`"O
cf�P���4��i	�q����"O
b�b�=��0�J�U��Q"Od�����o/��Re��)犄`T"O�ܪ�儺C�A�t��.y#^X�C"O^=AAJ�z�n`!T��<^$�"OF�j�Ğx�Y����/L� !�"O0�s�܋3KH�rF�6v��J0"OX4p6�6~�Dd
R#�= �<��"OZIr��5E�8\Y��4���+�"OND�2I?�ݘl<>�P�p�"Or�ѵ���E����˟�,_���"O��j�#U�MX��0��"R�9@"O�1ᐄ[�N��;�	���4�"O�`��)I�w�:�hW~4��"Ot$iP�'{�u*T͋�(��"�"O�t���B�l�
��L�K�2t��"O�	�AB;H��C�_ x�~E�G"O	��-N	A׀|��o\�J����"O� 8 �mҒ6~"z�Ο�X� A`�"O��a�߰Z�!bv,�K!�ya"O"�Kr#�
U�T� ӂ_��"O�)�ʟ�{NY1ԪB���A�"O0S��S�s�J!0�+OU��yA"O��{LC3����+ȑ6��� "O�}� -�hT�y�T���k"O�Uم��8�jt9Щ����"O�h�hG��t=� ���Vr�"O��K#'ц_|D�PD�kjTah�5OQ�5�ՉbO
��V��QQ��3��I�u!νSŐ�k�H��aɲ(urB�f��j��P�e���B���N�4B�ɒ"�@0ū���L�Vi�;$��B�I>�N���[	���Y'݌Y����$=?�v�Q%l�L�fEg1�����<1U)̭�X�h�Lߌ�Dtm_R�<9�iQ0
��Y��A!c!�*&HPQ�<A��R,p*���I�>r�Jb�s�<!��-��`��
ٻX�`h*��k�<���5��h ���3^��H �h�<9F��e��x�cŋ�e��8���n�<)�$4�r 0�O�>���A�O�<����*�X�YfRi�6���m�H�<IӈT�\��	VbP��r"�i�<�4a�`��$Dċ>�i(E�Q�~!�����H�&C<y8����%\�dv!�d��?� �C�!T@�D��"eM���P�x��]�ïIS,�¨R;c}4�Gy�gS:�ȟF�{4�ɦv���b�D<g{�ls��%����s?ѴgF�y�D���菷l|�I�c≟o���?�~2�	
'��+$�;{�4P]}���O�>�h�,�I/b�2�'%�J�����Op�����S.P�(�2BՇA~*���@�U�8ͅȓ>��ȷ������c��1>IU��\�܉�K���ԃPzb֔��8�"��C�N	��@ϕNL╇�srL���gֶO�ܳ�D�&��ȓ �n��v�����B�-@>c8,��2
��G�]�z��!�"i���ȓ'�*�# �k�^����[6X���ȓ �v���dJ�N-��Q�	�?g�L�ȓq��,��Aϡ~����S�\9Fຸ�ȓ&��`i��<}��T��5+�H\�ȓ��HӀ.0o#R���'�4=$�ȓ�
��c��:X�n!xPl_O9hц�?4�mh����ko�$�0Qk�2��ȓc�$!Qf�"����6���2�J4D���%��,��LaE�&*vH3j1D�P��^�S��v@Y�u��8�ua%D�<�g�U�y+���� (_��0`��#D�t	�߫bB�x��?L� K"f D���7,�RXB�ܰC��L��(D��Z�	]�o�z6��qQb��f�&D�������2e�f	U��ps�#D�t�  ]�~���{vG� ^��1B�,D�����ב�T�� Iu��Ġ��)D� ��H"0�z��ui\-dF�@c�&D��)����=}���喴M �b4a?D��ð	�	�����.�:bV�!�%>D�LX��� ! ,Ƞg*ԟC["x�ũ:D��p��� .�`�G
@�����4D��x0*�>�.4�CH0=А�f1D��C7.8AB�E_�j��7�3D���C&JK�L��	��b����'&D�� *Y�Fh��������e(Q�"O�E�>bp�D2u�N#U�	�r"O�q �D�*u���'D�1���"O܄�T@�3q�I2��! ���yc"O��R�6J�#�3;g�Kw"O4l���˱8�pœQ���t�8+d"OL�{A�3w`N�� 
�=v��U�W"Ox԰�� 6̺)9Djx���"OZ#Ǖp�T@��.[�*���"O���S(Qc�Q�m�/�R���"O:��TfàkJ����%j�F)R2"O��`-��P#�|
F+�[��X9�"O�u�&�+F$�*g��;vR��x""O2`
V�@�/��#5�֑R;�`��"O(����(|@���	><?���q"O Qp4�N�7-B���>�"])F"O�xZ%*K��.%F�N�$uڂ"O^��B��?�R�ݭ�d���"O�x����><�Đ �E>�^5�"O��5�C���Y�(<8De��"O�b��U�j�a��H��Q��"O�p���'�(Q�GL���"O����W"�vXh��I/����7"Oʤ1ch�(�,���$]r�AF"OZ�r!j6��T[ƀ��@@tq "O�E۶�S�bJ�銶o�H�����"OjV�ߞ�Ъ�LC%abT�"O�IK"c��ܬ���@�1J8[R"O0�%�$#�nAηh��y�"O�܃��ۂ4	�ԩw@�-sp˓"Oh;F� 5�
�aT�P(��3D"O�,� 	��j��ى*@z�h�*Ov�r&�u�@�y�ƚ�i_"���'$2��p͌*A�HU!�q�F��	�'�<0@șv�j����i�*Ʉʓ+�zTӲ	��P�~})��T&���ȓ���dg��\�ty�#W�W_�<�ȓ<����`��e��A�6c�@���p���Oܡ ��5�&A�V��Նȓl���	���\�ʕ��SM���ȓ���&��Sb�mj�l��xՅȓ`gl �7�9u|��5i2kҜ��ȓ9��\%�ߴq'}IVǓ�Jl�ȓQ`d��rE�7���E�.v%�݆������C"R2�����&-A���ȓ��ؠC,?*�;$"S|�`��jTj�`D�4H������	A�"21�P�UA]��3��A�[���Rv�qH��	�v�L8`A^�&�E��/NP�� �O�G���:�)ټ^[譅ȓ"7pRopܼjucC��a��Q��!��C7l��aҠI�/'��مȓp��Ⱥt섭,Y`��mHS+b�����`*�_cV�X��(X�MX�]�ȓh<�1$eӘ:��!�6`aeڠ�ȓZ!J0iԎזNH(С� `�}��p��P�#d�?HZ���M:����ȓ�T��j�6.$�Y'NI�Y+q�ȓe0||iV�S1x�`'J� C�I7��H�D �)SiFSULT��B�I�!!�,*���-�H9��U?Xt�C�I�A�jXS�n��W����˕N�C�	�(��)�)�Yșj��ɵ`~C��/h�V
U�E����9Roȷc4xC�)� �9�W�gx �q�+ē)L��"OJh�����k�*��0�1"O� Y�Bį���E��8�H�"OtJs�ݒH0Tq���L�V��"O�R��:8����D�W#�a��"OTu15#O�k����ViH�h��XQ"O"m�b*��0�%�׆@��1"O�mR։[�)\�[1f�6&�!ˢ"O�4�#��U��]��dN�F�x��"O`����K{$e���ڑx���"O4*
�MkĠ	d�ѦbnV�"OȀ��Y� jàB	 ^B��D"OB�"�>��s0Ӏ	Q��j"O\�y3F�t��B�++h�T�s"O�yx���u[R��!F�/h���"Od�,ԛub��Iޡh@�"O��!4*\�'$��"J��?��<`�"O6�ӣ
 �/��-Y�'� c��"O`]	aN�1R��6��<#2���C"O�yWj�
&�5�f%O�!-l(�"O�2�A�^#�����ֻ-�Q��"O��Q�K�L��Cpc�3%���h�"O~���X�`7٨���$u��"O�}kW�׆>IF-KQ�¤v��Dڒ"O.����ZYʍ�$��?)P��"On!�`Z�ihyA�A\<f;�W"Ox����¢a��|�� ��#��"OjY��Փ.qN�JV�}�r0�D"O�u���1,�n�{#	��� ��"OR�Zj�X2�gR�q�L��"O����	\�,��Y�q�51�
�za"O"���O�vM� FD�i��"O�9��%Gl*���Aa\袷"O�)H�k
�s
�%���|g���"O2!C`'%	�@�i�#�[�j"O��7�F�u�()����	~�Duڴ"O���'�PL2ʴ�C�>�@dZU"Ò���A��������v���"O�ɋ6��68t�k�)*�n�cD"O�x Q,F3m�L���*Q�X�"OSVC��{��Y!�fյ*5��t"Ofi �
h�|�p�]�fä�1�"O�P���%^�Y��	�n���B"O8���(�=a5v�HrV�O�� ��"O�9�@�G�]D	��M�V=x�c"O�؊@&�3|�ؼcr�Ҥ"L���#"O�����+G���r/�-X�����"OB�+������pB.��\��4"O����E�r�Z���ݥN���i�"O|� E��5�H�8S��=v��l��"OЅ���* ����uΜ�m�>x�*OLd�0��DN�E��>R^ԙH�'À��W
a��$ ��^-Ch�H	�'?��K���Ү��k-�y#	�'5�V��`�F��V ʧ�.�H�'m��U��-�<;�M���Ը*�'2�LÓd>-��,kS�M�W80�'�I�d�JQ�ޤA��+8��)��'�~!R �Q%�T���;4|NE��'�zxT��?@5X� li�'�1#wiI�`l�0��� �Ab�'v�p�[�^�*]��/$�ܬy
�'PB<��J��j�:�eQ)�Y�	�'��+��O�0"�S��L|O\��	��� � ��ȭn��H[S�_�j��'"O00(Uqz�����t��IX�"OX��F�@h�!�B��ҵ p"OrYb �
K,юͭr��с�"O�=��J1fQ���m=� ���"O\�Bb-ȯXr���b�
t��5r�"O�i���!]�����)c5��A"OzyѰ�E	+1������\�PB�"O]��n�'��� ���bdʔ"O�x@E�[�<f�f
P	�Rp"O��"��%I�$��qD� K�\�ȣ"O�͋B�цdf>�Y�cL�L��"O��br��Mx'lF�iϚ1jg"ON��̂�e]�-��+���lK�"O@�ɗH_�B4*�4r!vx�5"OĄ g�U9��d�wD�J"8"O<� 0/\�*��x�'n�<�V}[q"O��B悜a=��e�/��|Ѣ"O�8��O}ȈĻơ��6�d�"O�A�6���5�Hf�!�.��c"O\�k�痞W�UB�ϥ(̔(�&"O����l��̡��J�	ێ9�$"Oڦ���j�P�ʘ�W��c�"O��CF�Ôh���*�q��"O�4cV`�48��u�a�#@�ppc�"O�mZ0M�y[��8���1��d)�"O�[��.������E-�6"O���ӌ��'т9J�"D:Oy*0h"O�٣����(�X���
NP�IU"Of���/�0a�$c��N�Z�E"O�h�4ϔ'[�&�i�`h� � "O�Q����%oن!*��^.l���"O� ��7���Y���4y5��ڳ��B�<�1n�8 (�X;��8g�Ps�Ș�<iP���w�RA��(C*.��i0!t�<9�㌈z{�M ��N��t�W�s�<9��ԭ.e>��&O�{m4@&�s�<����jJ��{1Ɣj5��Ѳ��C�<��֔Sٲ��ԯؒIV
�Q�ID�<�&��"   ��   #  �  �  :  +  �6  KB  �M  �Y  Ue  �p  h{  Q�  `�  {�  Ν  !�  e�  ��  �  ?�  ��  �  ��  ��  [�  ��  *�  w�  ��  �  � s
 � w �! �' �. �6 �> .E rK �Q  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*hEz"�~���n.�h򂅵,�lq�Q�<&��;
��ʰf��-ꤡ�A
L�< !�6I���JŢðP�65��K�<�)@�,N��d-�*��F.r�<��펄o5>e0���2h%��
c�Kp���'h\�I�Ažc].ekeI\�P�E��'}|����Vw&5[E�ғv���'��8�'�H�aj�أG����'���Y����Z�,�A�:\D��'z�Ѳ�*%M<�hq�ū7��a�
�'x��YGd�1+�-0�V"+��A�y��r���[��̧
ǀ!1��A�DJ�d%D�hy����1�R��`��=jT*ԥ$D�4�Ġ��e�P��FG�	Q��*D6D��:��2%P� ����"l !�䆳M�`����7H|ٙ�D�
G�!�Dg�
D��NЈ�$2�̅�!�YJ< �Uo�G!)Qb�l��ɧY!�}�°>�#a���DT���>!�O��S1ʋz���`�����c>O����V�Oh]� �0�<�SŎ�
gkў����i�{*
��T�Q�B�X�� �u!�D�M��PĊj��.M�6���)��1�'o�$^A�hZ3���B���@��=D�$�wC�M�VM��m�@`J��D#1D�d�� �h�b�wh�1�"RU�.D� ��ˇC��Sgٛ �M���+D��IsቁC�|�`�p�Kw�)��hO��SŌ<"��L7a�)@�P2qK&D��C�� T�E�B��24�ZW |�����D�"�B�8fBB-i<z`G�ܕ�!�D�O���`�l9ܱ�tO/]g��.�p?1!�W	}_�[t��>G2��!.�`8��&�� @鶃��o|t�勆��� "OJ�`�,ς-)����V�5��e2�"O`q20���O����b�H���c�"O�ڴ��;x���G
Ǫ��p�"O���W�V�C��5Rb+O�ZnY�"O"�h^�^��0�⬒�hG�\s"O"|�bM/12Mу��$>@��
�"OV�c 
XR��L�0L�T?I��"O�t�RŊ�k��j`��b�3���^�OCD�t(-�H=r�}�lX��'Xx̀���,��e#%��:n*�T��'�tp�L��0S���N�Z�'�-�n�*��MӃ�& Z-Op��b�Z�[f�ÓPQX�ˇ�כP�x���IB~r/9:h��J3�v���9�Y��y�$�!��4"F���n��ATI��hOh��)��?5L��%-D�q�Qc�T=y!�Ď�z.zݑх�49�L b�mL^��)�'U���IHj/� �իe4����'���A�ã�$��#ʗ�b0�'<\HYDkTq��|�"�1	WF���'��5sJN�HL)	����	��''d`�0!Q�JCN�Q1�Ő4p8���$�m�O�\M���[�B�ւ��.I��'3�]�F��+F��`:�F*?\l˝'"ў"~��L9fac+j����B�<YtG�A�*xA�Ų?j��PC��U~r�'#|��ƃy���E�_�g)6Ib
�'�>=�d �<vB��:ŮU5u< x	�'��CQn�� g�� ����0����	BY�T�2/J�����\��C䉓F,��暼~�|�� ��fV�>y�����3�H �(^<.�8��Q�I!�D�&P�,8��XV�tS�eU�]�!��([��u���j�X�R'��!�J�F�aG�Rd�4�����~�!��$��H���r�@A���[�=!�Γl
�`wW�Mǒ �rJ��!�d�>!�u��J�t��((q�V�g!�d��h8P,a��E�
�e��!�đ*؀�Q��D�2����Љ]�!��)W�J02�I�$�fX��o����~
���?�a�Ȑgj��(׬
�}�'�f�<9P�Q�R�A�.�Qb�%��[x�'$�?�Ys��&æŲ�B�-l$�(�:D�(V*��U�H���J�yT�2�g3D���`Q>����9 u�SB�2D� �6C��E^\Yؠ�A�c���j�"/D�$���M$R�$TH�
��XA��,D�`S�&:n�J,;�CU�R�b�+D�0�H�.�dZrd
�g)��G�'D���w�Ӧ8s�����L��\�	+D�dzC��r"ջS�� �֨A��)D��rg [H�B]�G�6Z�l$��,D�XS�B��Ak&iJƤ��G�vY�e�)D�p�(�=�(h)v��O�F]q3�&D���T
�9=��y!)��=1G�"D���rc��iQ���,��d�1�"D�<Ǐ�y��ā�i�
��@ C,D����]�Je�m:�*R)e�p��7i(D��9W�ʑ�d�c��P�^��"*D�pb׋!�RU/����M{�>��0<Q��E�(��L��̢��tF�L��\Γf]R�a���D2�uʒ�yw����S�? Ƙ��B�)k��h��ބ=9��3�"Oi;m'_D<��UNa{�"O$4�E��
S�p3K�8"��a"OHl t��.B]��Whҝ 8��"O���Bʪ-�|��fUC+D #ґ|R�)�H���/��U��p@� B�	�|�`�pF�	�K��y��G\�k�C�I�-=�S"䇅Wu�[��؀K�C�G�dyX�e��P.6y��&֒SZjB�ə�M��K36������>Y��C�	�c�j� 6C�n�(
����B�ɵ@�=)' �Y�8�y�H�'d&C�	�6:ة1�A�%ư��ʌ9z��B�	��~���Z�5͘�A!��m��B��6�:��1G 8mgpx��$Xn��Tw̓#��a�	-j�~� u/ձH�}��%t� {�,X�� 0�M�q= t��$���2�G�4��<:D�ۼN�x=�ȓ�@��Kɻ`�D0RRe�����ȓ����H��X8R=�TC�+�\9��U����Q�N�X;N=�|�ȓN���C��D��ٚk�����m�,4k�EǸ7�6�իצ!�B�ȓOla%��:`ƌ̛Rd�#IF<��w�Ha��Iǰ=;�NDS�̄ȓ#���Q�M-0���+���=1�<!�ȓQ��d{G�mJJx��H�a�t���
���S��b��=���7}�V|�ȓZ\����Ç��Ke&4�P}��+s�b���b3���E�T�$�(<��ZG��B�C��({�H��+δ���ȓ$a�Mq0o� ��)��ڨ*���ȓ$���	�(;�R�P��j�t��F'ܐ���2k�����O��ȓ-alt��(��(�^��c��T�K:D�xY��D0���BDO�4�����>D��#k "|�K�dA�j�|H"�H7D�� #�)8�p��ݮWtV��%6D�8�����p���!�b�J�*O���P��]0��I����%�ʁ�1"O�[`��)[���O6%à�ۅ"O�I1���Cc9��̋/zZFy��"O��"'��XG��#e�\�RQJu"O����H�����}�Е��"O�pp$��*�������t$���"O�M�V�g��I��A��j� "OR���I��5D|�ʖ��<+n��v"OX�CeF6�U��#el��V"Ol�pE,�<�@��9����"Ox)S0o{�b���p�8��"O��(p�ǵ �(���K�=�b�:"O�{3�Mu�l�ʴ���o�<-�"O��[4��Ub8!(��0äACQ"O,q���B�X�Z��B�;Z��I�r"O(U�e��@2��ƺE�T�H&"O:$��/K�,	��Un �Xt"O�|��oZ0���g &�j!!C"O �� �(#��;A/�=Y��i�S"O�<���x����@���I��"O�B��
	[�	
w�-��\�"O挡���0�`����,��a��"O ����
��`²�[�xA�K�"OP�4) ;��l��@�Q.4l�"Oz�y��OT��h����	�$(0"O� T��dK��4�1�tN�3~����"O�}1�dA�=�r��L�jx*�c�"O�P��O��_�k�Bl��3�"O�}cs������h\��9�"O�c�@��+�8i8R��'(H Pc��'y��'���'8��'�"�'BR�'w�hIeA�=gD��C��N�84+�'	��'o"�'V��'R"�'���'v� Tb��$&(�%�E�����'�b�',"�'���'��'�r�'�&i�#B�-L	��
wň�OT�p+$�'�R�'Y��'e��'���'�2�'�V%N�vo�8��aO=�(5R��'Y��'��'�Z�M���?9���?1dK_4f?�!�Q��bj�I+I �?���?����?���?q���?��?�Faٓ(@�8��8xZ���bC�?q��?I��?���?���?y���?�4㉷F�=S0n�w���Z�)�-�?y���?���?y���?)��?Y���?��FM�Gj�!p�"T�.�8�A���?����?Q��?Y��?���?���?Y� ë>�ʩ+��+GԈ�0EH]=�?����?���?I���?����?����?�(��f��v&�A���st�O�?����?����?9��?!���?��?��)ùG1Z<�a"����k���?����?Y��?����?A��?I���?�#�&hjH4�$��&(�S�BH��?y���?���?���?a��C���'��FSg�y�"�Ǩ)U��k�d�6��?),O1�����M�w�P�:C<h1��N�rr�$b��/bV1�'��6�-�i>�	��A�
�U y�)]�f���Ѷ�PΟ���K�x�m�D~b2�l��l��N�",|1�IV>n��A�F3]I1O��d�<�����K��ar�	9bJx��J�:D�	m�l@c�T�Rq��y�
�X��dJ��$ ((FC����'��Ĳ>�|
�#ŧ�M��'�` 8���lj|˒f��h˚' ����i�i>�ɞQ�t� �C�
y��)U�2���	`y�|��e��Q���Zg@�a1J�����K:⟼	�O��D�O���X}��׫o�,�6,��6!ڭ�	�����O�Уq)�1��ԫ���d�//p�c�W)�#T�Ҏ\�ʓ����O?牋ZE�]���R�\Z&�3����M�B��R~2�t���S>?�F�ل�[
$�|�P�N�W���˟���ʟ#��)�'&��?-�`H=[?��\�!&�a�I4�' �i>5�I˟H�Iџ��	�A�a�W� �q�@] �ݕ' �7�LT����O&��/�9Ox�j!�(y���vG՜/� \�p,l}� o�ԕm��S�'9h`ڔȍ�4�rX:����`^P�Cc�P.T�������9�ł>8O$�
]w���'�ŕ'����T�bz8��-
�m��P���'�b�'������\��z۴C���3���g�߲�k�����1�v�0`�4��'q��e��&g��l�<#+.���^C���Uj&�<�����}��[�Ƅa���",�$�~�D'���/[�P�lHҡĳV�
ْ�N�<���?���?����?ш� ��4^�)S�Ш]侴�B��.?��'W�+l���:��<	!�i��'�`1r�g�8Q���")�D�[�'�B���D���;m�V��0�u�$Yd��h4��;�)�r�Ӎ9�� �5�'�(d�'3�6-�<�'�?���?AӒxqX��EI�/�J������?�����ͦ��H	��	՟��O�nE�6��"�f �"�wQ��	^~�+�>���i�h7mM�)J$ϛ�+0Fp�5�͋D�P����F�x��jO@3��'��ם�U|��by�w(<�3�\*g�Mj!mQ4L�<�2�'Q��'���O��I�M{�*¼Vt`��@n��}����ϑ�}��s-O�nZ�x��I�AJg�#3~hhk�ߋF��y�s���M3T�i{n��i��ɠ2�hs��O��'�,���g֢+h-1�G�8^Ԓ!�i����\�I؟��	����I]�t��!�@�[DE!~�\k�Ğ�L?7�ΡvJ��$�O���-�i�Ol�oz��D�[���� ����;锽Q�C� �M�W�i<�O1�~ +�j���IOf���;Ғ=a�-R�y��	�n���S�'�"��'p�7��<ͧ�?Q��ѳS���3�j�.�zJ9�?���?a����Y�� �l�۟��I���['IēC�F�xUlD5f
9��Yy������M���iݞO&�J%9+]&L�^�U#pX����X��-F7S��V+6?� ����_�$���;�<L�u⑩g(6�ضgcmy���?���?����h����^"_]摠v��74"�0xхD�'���$�Ʀ��Gg[y�hs�V���#x��M�ѧ��0���H�L����4�M���i�&6MI�[��7�7?�7���\���R5=4x�(�o*ܹ�5a�1Zt�+O��lZoy�O���'�2�'JRb�P�����Ĥ?� �U�	q�I*�M�`c�-�?����?�O~��aߎ��ghJ)&d�����)��Q��\�0;�4J���C1��IA�I�����
�6%�.lK񏙜��m�2"�=��I�9���â�':�E�'��6M�<�%@ӲcX�Y;�.����{��C�?q���?����?�'��DL����D�$��- l����9��u�Ƥ��hPٴ��'gp�d����O$6mϢ(���#��G��R�lĂl �|R�e`�6�P��X�
@AI$��E�r�)����� ¼q	C,BV>豳LU��F� �>O2�d�O6���O����O\�?E��/�**�B�Ca���m�:��Z����	��d+�4}�Uϧ�?q��i��'����g`���u��@�$[�(0��ݦ!���?��p˝�)�'�I�Ul��J.Bh�2��J�t0�EV�]�`��	�(:�	��M{.Ov�d�O��d�O�4�DR�� �8)]n�Y��Op�Ĺ<yG�iC��{�S�0�	o��Ļ]���%I�:�L�o�n��I�����٦*���S��+Ѥm��\"��P6jyX�$Y?R���&�{��H�W��B\w�� �	�d7�i���E"ejD� H�CC8��!�����	˟�����b>y�'��6�ͫq�5�T&�3,��M�&�_)f���g�Ot�U���?�6]��l�4[�N<�g5T(P`'��/���4z{�TR��6O���ٞ%˼��'=d�3��}I���h�K�-�<H[c�i�	����֟@�Iʟ���Z�t�7��)2�	�x�[���&_��6�?D���O�d6���O�nz�)��5��
ɂD�"�(��4J��x�O���OF�e*v�i1��I��sS ��V� �mӯpF�0*0<9�g٤˓4Û�Q�L�I��V�";�� ��yӼ�Q䋆ҟD�	���Py�i�0�qu��O��$�O��2�XQ\�� �5?��h�0������O��iՉ'L|4zcgG,w�]@��(i�]��O��k���%}�V9봃�<�c���Q���K;���)������K1�}2B��r*���O����O�$�'�?�!�fɘ��eNآL�@b��?�t�i��S��'.�b�(��]̲�"s�(�x	t�9%E���ٟ����-w�ɦ��'\�B�.��?����M��!iŢ3��\@0�
�Wg�I'�M�.O��$�Od�$�O��D�O�иT�̩=_�h���'U<�!�	�<1��i�\$���'Z��'��OY���M;�$ش,=#<J1�B��(�,�@�Ə�O�O�i�D���>ڎ�Z�,Ҕ0������}�U�A���p��˓m�u�g��Oօ�,O�lZy�}'B-�\�(���#5�(���'��'�����S�$
�47�T��;{�@��V�a��!@ւ�]I@��3�v�dKH}��e�� �	ަ�s(%;U6��Ĭ��3���Ѳ�|o��<	�!!:�j�lZ-O�l�;����@� `~��REgՀ��MZ&e��<	��?����?���?�����_����cd�w�\Y���^���ҟ|��4"����O=�6��O�����!��-j�8�oAQ���r��|��i�j7�ퟜ��E�|Ӡ�蟔ذ)��$H�
Y ���cL-;bq��'��&����4�'���'���A* �3$��O��'^��q��'��W��۴MU�����?�������<���$~pp�$��I0��$�O$��9��O��T��	,��WIT���}�`�t�0�x>D��U����x�D�E��0|�L����dE�8���Imޝ�Iɟ ����)�Gy��x���O���@1�����a$I0�F��O�mZ_�8o�I*�M�1f��%bŢ�DH=aо1"���ob�6�dӞTc��q���&r���d韠1B-O��G��1�h���c<\x 4O���?����?���?����	ʾt]6�5 �<+�d	��o�b����������?i�O�R�h�󎄣c^QjFFV-�FY`��Zyz�0n�;�M�%�x�O���O��-���i�D;� 9�B+�6r�t1YV�[�@��Đ.�Hyk�bU$�OD˓�?!��
����*g���1F� ����?	���?�+O�oZ(z�J	��ܟ��	6�����':���Ƌ��?��R����47,�Vh&����k3�C�E���£.E\/��O���	_	��e$�<��'m!^���?񥣕�Z��� P�4�8�rw���?����?���?���	�ORc�ְ@� J�F�'L��ł�F�O��oڣS5ބ����P��4���y�A�3{�xU���etv�9����yr�w�Xnڏ�MC�jA�M��'Q�'��CB �S1{�n@3!�,-P�*Wf�6D�}9��|BV��S�����П��	���
7�� )�d�[�&[� � �%�~y��z��4A�O��$�O��?�붨��H��'o]�_$.�������D�����4\���O2� hŞ=����Y��0�, ��t��"�D~�&|+H���	��'*�ɤgA�a"�͓�$8<��U�s"�����0����i>��'�7�S0 ��K��F���ŏ��:��%_n������?A�^���4��Veu��d�S��z�Q5�t�Dy������6M-?9�m05���i'�����C��q��0��Y�h{����c�L��ßx��ӟ��ݟ��2ģB2fG�� -Z��x�!DH��?i��?!��iH�x�cX��޴��IC��ç�M(;�c��I�����x�`z���n�?!�Ӧ�Γ�?�4D�=9��4@J�[84@a-��E����O�T@H>�(O��O��D�O��is�C�}�4�8��^�(zp�a�-�Op�D�<ǵi-��1��'���'�哊,��`�Κ�Tl����&���}��	��MS��i>O�i�b)�(H����T�̐L֭�+�4���+��L�	�?	i'�'�8�%�T�o����i(�D�IwP��A�ܟ���ϟ��	Οb>��'6�,��0���I)t5|����[���!�j�O��I��u�?�1^�0�4_�|�ƈ��]m�}�*��.Tb�i�7�J�	w�7Ml���I6GG�r��O��S�? 6��QIߨD#�[
��x���x�>O�˓�?	��?1���?�����)ͥzY{O^���Q�C�]0�b�nZ�x����I�����Z�s�H������d�J�p��/��%��Y3#ݱ}O�Fu�0�'�b>�h��Z���ΓY�.iP߀F d��8g�6�5�Q��Ol�{N>)O�I�Oܑ���i���H����M͠Y$�O<���O��$�<1F�i�^�H�'���',�qq�h,<��1���Y�)���čp}r)l�|�IU�	�2��|4�,#�Ǆ�rr�XJ2
{����&"@L��V&�$�b��'��D/�۟����'��QµJ�v"���)�t�|�d�'���'���'��>e�ɄU�v�9��0�8���&(�a����M�_�?��7��6�4��ŀS�P��Y��3X����0O��o��MsԼi�b�1�ie�d�O~5��e��J��B?m�p�W�I��p�$�V�"�Ot��?1��?!��?�dr�lۄ�X7x�)�)N�c��,OP�lZ�	wx�'�����'A�yz ��a���1`�E>#�`!�c�>1Եi�X�.�4�T�)⟈9;F���6�;���&� }#@B�*vD�'h�<���y��ğ ����P,0��*�* j��ԡ�����'Rb�'�����$V�0{�47�D�1�:*0`��ǥ}��Ike�V�uX��ޛ���syr�'t��g�r	xq�A� 
��Ş�wH������6-l�X�I4sP���O����;�츋D�ǹi�89�i�r���?���?����?����Oh4�*��̪G�V�b�k?ZP]�V������M�aRh�d,g�ȓO2��(�{qz�b��
6�`��u.Rn�I�����?�Z��@��Y��?Ѵ�] u�Y
��&,8֜�aŶ��B.��?Iǁ)��<ͧ�?��?�&(K�P���S���8%@v�J�:�?9���$N���*U����IП��O+��x���	L�<�/��
ri��Ob4�'�"�i�ȓO���O)*�Xt"-g����v�ƩQ9��8��ҫE"4�Wo�����$HP���OZ�2��ƹI9�`�
�f�5J�O�)n�/k�2A $�O�k^��+�)�Dxh8�f�ğ��	��Mˉ���>qw�i�������sȮ�!�`ч{V�
��n�DtnZ���4o��<	��4�(�[7�� ��(O���e#�!p�Y�]B��Pq:O�ʓ��=1r��Z�SSB�*X0]1T"�=�V��cib�'��i�ͦ��4~�"18��߽gh���ɻ\�|���4vƛV�?�4������}K��eӮ�ɑw��d;�ဗO�^�(���'��ɷ��D�'�n'���'�前p
pU�B�, ǚa�ǋȉ0D���	�	���֟���Ο R')��<� 
����x��A�Ŗc�����MC�i��OEࣄ��f+���� 	:��!ez���	&�P���Ù]t�'����ҟHѕ�'�l����@\<R��C~VU��'�-��DJ9xaLQ'O�V}2��'�6-%fk����O9oZE�Ӽ3,�"8�.,j���C�|MYt��<���?i��if�r��i��e>��7E����Ռa ��zeǙ!k�(h��h�Q�'��	ԟ��I˟ ������	�	-�L��K�	i�ذeS�q�"<�'�7�X+�����O0���Z���ykw��++d�)2�fܾWw��+�as}��'R�?�4���d����ڑ�\�ر
�EQ�xRp��`I�>H|酘�� ��A�kx�Q{��Wy���*��;�.�%�����!22�'�r�'D�O���/�MCB
��?�a���qɌ)��ґ�`��pD3�?���i��O�%�'Y$7��џ�ozᦩ u8� �+07���6��[�f�nZ�<��k�������p�+O��)��U��/M���� ��[5r+�LV;O����O���OR�D�O��?������a~Y�C�K(d�$0�&�Ο��Iן���4jk���'�?����'�p�+��,�A�Wh�y�Ļ�`����MKe�iH��A�g���5O��Ā@iX�U�B>[1��ʶg�"Ee��F� �?�#5�Ĥ<A���?9��?�Tl���AA3Iɗ9��CcP�?����$�¦�q�g�Ɵ��˟ԕO���$rg��W)�7Vv�!�O4L�'�D�V���$��S�?��T�?V8����Dݰ(Ej�SrB��L��2�*س?C-�'<�d��$$�|Be�Nm|��Q� �1p��Ä)
�f2�'���'��O��A �O@�	��M#v��*3�<��e��q�ce�M �����?�¾i}�'�̽>�ôi�=� ӄ{iےdl�*H�'Jqӌdn��Zm$���y��'2�h��?���Y��1%���Vu�s�k�1x&�}�H�'o2�'7��'��'F�ӛu�����0V ��Ь���ݨ�4�0.O���-���Oz�lz޽A�"x@� �["ٙTً�M�S�'���T�O����۹qߛ:O��U��d��#.��w��kE;O�]�G��?qG!�$�<Y��?��K 	{�E3�mJ<\����e]��?��?a����OѦ��a�kyB�'w>`���_$v�S')X
.Și���]}�"�$uo�&��RP�QK�>�:�:Q�_��0�'{Ή��,�&r()���d��&q�T���n<�:e�1斞T����m���=�Iß������ş�2�	�I�4�'�g��'6	�u��a< ����'�6�����O���O���O�EnZ�|| ����%������WtZu��n�� �4S��u����LbӾ����`��u�����?ۀ �e�J�K�<��	ϽD�����#4�D�<���?����?����?�TkԖ#V�;Feطn��q	���ڦ�bs�͟D�	ӟ�rPᆋ;�Č�v#E5VS��&�G�9��%�Mc'�'�����O��4�:���\�m��(f*F2�����*ؚ4�	���R���K��'�zmә'�Z�M��*�=3�0sѩ�5�ؼi C �?	��?���?�'�������.�͟���j��Hb��-I�y�Yy��|�OO剰�M�µio�6��)k�r�ʇ@Q��JXj@�$rf�1��f����ݟԁ���4Q�ju�e�ry"�O���Q�z��|)@σ ��ї톚�y�'���'�b�'���)�r���2t��0�BA��]*�����O��D��qr'�z>}�I �M�O>A��T�UkR
R�m�h�Q���0d:�'��7���m��V��o�<Q�e;8�(�ʔ$g��th��ͩ�B��� �6�X�DJ�䓷��O$���O��$A�*p��A��(�h�Q/��|yx�d�O�˓4x���؉"�'�S>-��̪ev\`ZEP��Q�3�:?)�_���im�r�|�L�`}�:���_Ԕ=Ô�
�,���f�J8lz�/O�IZ�?�Q�7�ā<K�ݘ�Þ�c���p��Pz(��O��d�O���ɨ<�¼i�\}��^����*R**К0�р}�剷�Mӎ2*�<Y�4R�	X� �1!�ֹ�v�ЍY�<��i#6� M��6�+?1�`±-����1�$#�:Q&�Q���>q Z�b�g��yRP����ٟX��ǟ0��Ο`�OiPx�g�@�\�$���E�3~rX �b�$�ȆK�O����O���d�ʦ�ݲ>Y�f�W�2||���_2!;��A�4;қ��,��	�2��6�u�Py���H�(���hS}N�Iӧv�$�4��BD�t�I_y�OH��9��S���J�����ҌR�"�'"�'�剪�M+hL��?����?�jÀcP��5H[�W$�+g��#��'���3Q�&@p�2T%��I�@�$�ҸY�#���jհf�.?Y��T"^Zrcd��G�'RY|�Đ��?£�%]��u�-:@M$RD,t�������8��Y�OA2@�":�R���#>�A��gd�@��Ǵ<��iz�O��;
y	a"^uʦy�B%B��צE`۴m��V�S�9,�&��x�ļK���g�-A�]HF'y9jA��D)tD�$�T���Ϙ'�b(���#&5��H2ݮ6�|j�O��o�.m0��������IO�'��}���nP���
�mZ�Yc_���	Ο�`K<�'�?�'e��$aˬX�>T�FY�d/���MӖ_�,{qd@�9��6���<�Q�27����,�u�Kk��?a���?a��?ͧ���Ҧуb,G̟tӣ��W���"&'^QojQC�`r����4��'\�6��F�qӪ��I�$��ѐ�*�_ڄ�G߆TRq���bӆ��Q�P#�z�JN~"��FO�h�R/u@�!���&����?��?����?1���O�P�ڷ�ڂt�.]-�%8ҕQG�'B�'��7m�6w���OJn��'Ŭ�(шO�	�̱ ��]�9T`�*w�*��O����0is�y���	�|�����B�Àb�r����5��&_^ڝp�O��OF��?���?��	�X؆�B�A��hĎIl҉����?I(O�Im��..(�'�Y>�p�ᙈc�^`Pg�	��\X���:?)�_�X�ٴ3훦�8�?EXQ�ܸ
ߊ}ʕ���O#�0@���z��V�\v:�������ɟ���|b��,ek�xȱD���,�'�¢_�B�'_��'���dZ��K�4!8�(CX�UX��N>z��2��β�������?�^����4p�,\�]�Q�*o�	�Pk��V�y�6�ZP�s�V�	�n\9�柒	�*O��-Շ6;<�s`��+��52OZ��?���?���?)����jGv���.M��؃�O��e`�f0�N�O����O쒟�d����ݿ0`(���"0�Q@�
d���)�404�h"��F���7f���b���q�B��*���b�Ol�����-�"˚|�Py2�'�r�G�5�T����tS�PQvDҎW�2�'�b�'Z�ɒ�M3�,��?����?�� �7���0��9:��z�i���'��������H<�gJ�0	��P���9VҺY�ȏi~҆�s��D%Q�g��O����g�b�Ǹ*����b	
lM�5K�kya��?����?���h���D��`�� '����6i���$�ɦ�8���П\��!�M���w��p���4
��` V�1���(�'L�7M�ߦj�4]�D��ٴ��$PcL���'NP��Ҟ)�N=��*��y���u�,��<!����ې慗sB�U����)D�Iу��Z�4���[��?���O��y+O(,8��ô+1iu`�<����M�3�|J~�d�X�`n١��@n�r�e	�L	>)*@ �����!i|5���[j�Ot����bĈ&6���@�G������?����?���|�,O��oZ9?����+pr�H�fBb��x�RD/J��	9�M�����>�i��6�����X�g�q/n0Zp��'���,��<�0K�7�+?������	���'��c��O�q8&�ѓHP�q��;1�D�<��� Ū�$N+fl���1�N�_1�h����?��5]��HF���)�ߦ�%����D��b0����R�nX��e ��W��f�~��iO�b5�7�)?!0/
I�? ���B��A���SAJ6d! �
�DL
�?a��"�Ĭ<����?q���?b*�:Zat��ˁ��|�����?	����զ�8�C���	̟��O��q�e.�5�4|��,��Q�jX��O:!�'�b6���SH<�O�H쒲����eJc�(u���ҏ)�0��"��% v�i>����'� �$�,���އU��
t"]w��L�VJ>�LzشK��Ȕ�߮�Ӂ���-:%�ۛ�?�����dOG}r`� #�	��� F�۴P��q��)�4pB�!��4���ɀ	رH�'WTʓ��Ź�.����3��:-i~������O��$�O4���O���|�$� �J8��k�mP8.2ε��g\�uN��'����'��6=�r�5&Y����a��Q�ܙ�$�Φ%ܴ,v���d�O�t�Ȝ~��f2O�$[��
 ^�hQ�������D9O� :��Յ�?��	1���<ͧ�?�-B��(�%�G�(����%f��?����?�����ɦ�RYޟ��ߟ�1��ݿ� d��Ŋ,�TZrO�[�tY�ɗ�M�'�iXO.d�%���a��Q�gE.HJ��+22O0��55f�9�3غ'J�	�?�k@�'E�X��p�� y��Q�f�Z�;�v	�V�'~2�'���'�>��	�)���T����5�KJ�u�X�ʵ�'L7Ml-����?i�i�O�Λ�{�����Di;�n������%1ش|؛���}_�6?O���6n�5b��~����a�`��L��H>=�$����(�d�<�'�?���?9���?���G�K�z�CϨ����3�����ř��ȟ�	矨%?�	�Q�2�3feǫ�4����W�^@LU��O=lZ�M�x����ՠF�!:�D��$U���� A���5�-������h�DN��O�� ��I���ƭrY4�+s�E�G�l�R��?����?���|�/O.�m�n�N�ɘX�ؤ;gHY97C�up��˥0�b��ɧ�M#�"�>�Ǵiw�6-���X� �f�hRv�ܲ��lb!�W�+�Lm�M~�E^,9�[�'���f� i���L@4G���GL�<Y���?����?1��?A���#��83�7-�<�k�!�.>"�'X�	d�4�j�5�`�ąئa&���%�5w3���E	�d�C�I?���?���|"v@Z��M�O�yC��]���A�$N�l��%���̱��m��-@��O���|����?�t�.xh��U$]
�f�ׁh�|03���?�,O�n��i�>D�I�<��u�D�6�L}P�%�*}߮��Zg���k�Iҟ�	���S���	1���!r�ñu+� ��E�b���Cѹ-қ&h�<�'4����J�	mv���B��D ��6̎�%ˈ��	ڟ������)�Sy�|���!�>u�\� ��BF�왗䋶^C����O(Xo�Q��4����Q^X=	I�V�m��A��֟ �ݴ ����ٴ�y20�b�Y�Ev�)O�N��iQ�kȑCB��
AթeB�<����?a��?y��?1,����B�ߗJnn�	@䆣p%d�j��@զh���̟���ϟl%?��ɓ�MϻWC�����0	YR��N&jez��?�x�O���O���ɱ�i���&Sf�����=�`�J�[��$� Oo@��'��'�䟨��:;8�ਰM��,c\��l��*dz��ȟ��Iܟ\�'zV6��t/��D�O��(�e�f�		D���wiʨ�d⟸��O����O��'�@ːH�� 0����?"2� c�@c���	�XY����Ҧ��,O����(�~�'q���6nQ�m�<�aW�ېE4�`�'���'v"�'B�>��ɽJ٪1H�e@�c�� �"���ɗ�Md��?A�E��F�4�^EQ�	m�H��4�
�O�v A�>O��l��M��i�Tٵ�i��	�`>� �O,j%�AC�(h��-�<[�`H|!'�̔'�r�'Ob�'���'�H���J�hm`��ql�6Z��}�uZ��pش3�������?Q����<a�ԁ,�0�H�B�f᳥�ڡhk����M+�i�rO1�z�ʶ�� *g�ugF\ 	�~��L���|��@�<���C3t.r���������
�1Ƅ��+S��@X��
A����Or�$�O��4��ʓ.�D٩vT�@�ؤ\�$�A�2���§_�%
�
h�t�L��O��o��M�i) =Y��Ag��R�nY�'z���d��Y�v���yR-�BG�d��S�߭C瀤v$�X�6�?I�|�A� q�L��ҟ���ܟ����@�z�C�"C`bԺ����-�q���?��?�ӻi8�Ms�\���޴��(��=#�� �c�̓")��A��x�n{�d�	��$a��?�����X���-R�B�k�A4`�x�äf�(xj���'�@&���'�"�'��'����`G_��h�ei��&|�}���'gB[����4<�&} ���?�������&��AQ��0rӺ�#uM\}�	 ��D�Ѧy�ܴbS����?Uc� ��L]�6uZR��
5��ڴv�,�%�C[y�O_�1�I,�'/��$�� +#�ɠc�$5�����'4�'2�O(���?q��Ɍ8�|�1��A H���G�
h����ݟ��4��'� �U,�(\(b�&��p�� Æi�g�	�x �7�� �"�Ħ}�'� ��?U�gX�$h��	Go
�I8�A��I{���'8"�'+"�'���'�哝f:&��V�$8Ֆ��b�
y����4H5 }����?�����?)r��y���=�N}�vD�>`�$���F�>_h�7��=�N<�|±
��M���� )q�L�%�i�U��P}��5O¤�V"��?mm8���<��?A7/V
WР���D�A�UH��ب�?����?��������K%��䟨��🰘q�5LQ �)�.�&W"��Z�f�I�a�	�Mv�i�ZO��2���S:��@׈�)��LSÞ�Tq�Q3	��U�V�B�5���Pҟl�f�=А-��"N����h�N͟ �I���	��<E���'���Y�'�,��,{�'.���R$�'-�7-� n��$�O]mZH�Ӽ�"�M-��q��"�k1�U[����<���?��i�d��i���5���k4ٟ�A���6M#�eP�m��uӴ��"�ģ<����?Q��?I���?q��V��" Aн{P�|�˖��˦}C������	�$?����9fH1ƀ#���@eғo�L	�O��$�O��'��ޟp��di̅覃��lю��'c�i�
my����Ւ,O�H�V���~��|"T��������yC�b�%ee�����������۟�Ty2�~��Ԓ�i�Ov�Z2�=ڤ�FK��*P(�O�am�U��IJ�	��8���M����0��xC,��XG�Z?�P���4�y��'��I
��Yi:)Op����$����U�`M���Y	c��i�1O����O6���O���O��?���H�$��P�gG��}�� ������	��L)޴��'�?IU�iR�'�R���E)CW�	8� �Cº@˳	5���O��4�$��kxӜ�M�X�`#��G�A�w,Uy�!����;Q���n�I]y��'���'`BgʐU��䄏u�����X�'e�I�McĈ��?��?�)���e'ju��BG#ҵ*��<�N���-O��DgӢY$���򟖵�m�.CT\��
�')����Q+Iۤ�T#������?	��'4��%��R�����3G�TC�(�q�Z������ ��ٟb>��'��6Z���X�'#�2> ���C̗�z�����<1G�ik|�ɼ>���,0�� ���!bF���&Q��z(b��r�V�D�+��6O2�d�s��Y0�'F	�	�&���8dݢC,,C��Jc���Ny��'RR�'-b�'��V>�T�GK,�u�geK�*�m�f��M�dE2�?���?)J~��3ϛ�w����	��p�����,܉w����'�(=�4������ps
nӸ�ɀ*�܉�砊�8�\VRrF>A�'��y��gN�  w�|�W��џ\@�O���� 1���$*B��<�I��$��}yrt��aV��O����O6�[#P�T������J�@ᔯ#���O�T�'�6mɟ�&��{qcD�X)#��PP�I��he�T�I5"$a�o�"����'������0�'
�)�	�/� ���Z�����'��'3b�'�O4B�A�3�-�0[ι��h;B���0��D�r {��AQW��O�D�$� �i�ɩSI�,����PMG
t��k����Mð�iF�R��i���Ol�S�J>���营)"P�!��/i���#��f4��O�˓�?����?���?���Q���� ѕ��)�/ ��,O� nZ	���	����@�s�P���ARt�@.C�B������R����ǦU	ܴT񉧘O�
D96�l���P�,˿k�a��C%�D�e]�����նdZ�!�e��wy̈́�q��<���6�Bm*�.��A�2�'	�'��O��	��M��j���?�e%9b.��J���,������<�ųi��O���'�^6m����ڴeC�|��=+g��8�KԒ���Q����M�'&��0Վ��8z�	�?5���n"4%B�M��H +�K�:@���	����`�	�����Y��I�i;��ݽ8=�!����������?���?c�&�	��	��M�K>��AH>H0-cC*��c�RLrFf��H�''�7F٦]�8	���o��<q��J�����2�R�w�I�V% ��E
��!�����OF���O��Sq�*���!�B9.�)%FE%)����Oh�9��Aʯ�e�i���',�:�;S�	�A�
m�6&� in�@��� �Mcg�i��O�i���]�K<FD ˷"r6Z&�u N����Gm(�����O��J>'�A%d�T-�4�*�����?���?a���?�|�*Ovqo�:zP+�D&K�,)Bo�s0�i�3�^�>?2�'�B6m'�	���dJ��a��H�!]����� ~�-W�W��M���ib~�kQ�i���O�0'5����<���VX�l�R�Qk�Z}Y�	��<�-O��$�O����O>���O��'c�`@�2�߈�` Z�,t� q�ԼiR�a��'-2�'��O/R)w����4@{"3�Ŕ0%S�����}�]oZ��Ms�x�O��D�O'ډ�i�3h/��6G�)L\5�v�	t�d؍s ���k'��O˓�?��'�Fl�ӹ+À�P0d\�d"|\q��?����?,Otxm�/�\��	��	&�tq�sB&<52�GH_"`���?�']��۴<z�֠?��*k�L����\"�)��/2%�d�Oju�%��.v��Zä�<��'�����?qq��r�a2U�?��Pe���?!���?y���?���9�}*���+a�|%y��u�~��O�EnڡT*��'�7��O�O�N�$"xa�	́&� +�48�Dk�vlڿ�M��߃�Mc�'h�:Yw���ӑ��Uh ��}j$��Bf^'K���I��|V���I��IܟX�I����/J�EW�����3����CKy�e�Lh�OV�D�O���R��$kR2� ΋�\�F�� mY ��>�i�7-LZ�)��?��� ���q��?\d\�BG�ZН2c��)� ˓v��7��ObxN>�/O "�1F�DuM��̤#��O����O��O�I�<�&�i�l����'�P�)E'ےFA|II�{�Q0�'�7M�O��O�d�'ir�'�T7mɕ�n��l�u'�X��K�2�Di�`lc�P�	ԟ�UCҗ*<��%8?9����c"ΎS
RL a�I�DM~�B��@�<9��?)��?���?A��ġ�7MЂcV�>uD  K��@oB�'���e�t�c�=�����q$�8�$-Y'�TF�q6N��#���ᛖLg��	P1eqD7�%?I2�E2'�Z��1B�`���+f\�R��O>�L>�*O�$�OX���O��%/�!n�6\�ǃĖP�P���m�O��$�<�3�iÆ��g�'%��'+�Ud�iNЕ�\�K5e��)������MS��iFO�I�\��[�Kߴ�Z5g�H��P�&Ƶ|�JQ���/R�˓�i�OViPL>���=�ڍiE�&7��=6gΑ�?���?���?�|�+O��l�8�V\#�,ߗ&&.�
c!Z�ΤrA���t�ɲ�M��b+�>��fe������V�P�:0	G,�O��m�Iz^!m��<i�O~69y@��?U�'�z��5�F#\D=Ƞ�F@��;�i
�j�@d� �ׄ�Ȝ��&�e���G�C)t��!�Zx��k�~i��H!GȞԅK�\z��V,��C*NB�m��b��ç<��6V�E'�1���)\� *3�)cG8�9�@�	Jdl"�ƭ(7t!R�Q�Y��q`ń�HV�(��
o���.��'���C�85�)I0G�;j��y3���d��h� ��G��g-%�Kᤚm@�JS+��� �A�59v�b�ˮ=�`=�ٴ�?���?���<�Igy�)��zJv�2SO����q�zm>7-_�/p�$����:;`M�઄� <��g�5#����i,2�'�bQ9X
f�����OR�	l\mA�!�e¹�0,�}d6�<���1��$>U��˟��IW�X�'>�]��[�kXl�۴�?����o9��Wy��'�ɧ5&&BH��ؓ%�
��8�c��	�t\��O��O��<� ;޽(��.8�4q�-�#x�ʥq�S�ԕ'qҞ|��'pb�ˬ\*�`ŌQ�X�!U?}�8H��|��'<"�'��I�]���+�O��q�b�&:Xx�	�i��L8�޴���Ov�O2�$�Op��d��d8�CNM�d1����%n,��d�>����?�����lp���OH�CN'O�� #6�^$������z[6��O`�O����OB!U�$�I�u!��;��Vta���W��7��O��$�<i厒�dM�Sǟ`�I�?p�.Ŋ'/6H���*c޶@���	�ē�?���������䓒����-w�t��g�(c��@�eϔ��M�-OdQ�Ĥ��Y��쟼���?���Ok,R"��AiツBΔPZ���%�6�'l�NѪS.2�|rX>�L>��!�D8�J!����b��mڃ_,��Sش�?���?y��	�	Uy�U�xœ�Bۍh/T����J#6�t6m�.�R�<����*qٰoT�x�,e�PGٮ}Nv�ۃ�i R�'����s����D�O ���V$& ���	R��z%��*T��b�`:"/�a�؟��	󟔘`$S�Ϝ�aE�5A���� �Mc��k���PQ��'V�|Zc�X�2AK�N�>�ڗ/�5_Z�;�Ov����4���O��D�O��;H>�4�8U�P0jL+,�8�D;$��	jy2�'k�'Y"�'� <c��/a?�hJ!�ק�������=��'���'��S����G�(��􊗟1���R��	� 5&\XŠ"�M�+O��&���O ��
����an�k�
�-���*�����l��?����?Q,O�R�EBz���'o���N�'H�^�be�܁zg^A��x����>�d�O���;4��OZ���F�/?�D.� J���0#�i��'���.���KK|������`Ӑ�;Cl�%�F�"��$�(�'Tn�F�'��O���W��ܫP��S�i"g�A���	ş�K'lS��d�Iǟ`���?q��u��՗r�ڤA��\�y���M���?92���0�&��<�~:�n��vB�[��8Q`�l��,VԦ-�#nH��Iݟ����?���I��}��X4����(E�a���l��J��)+��=�)§�?�`�W�?9~H��ȝZ�2隵�U6���'�B�'��|�!�&�4���$��L��?^n�1�2OT#�T�{�Ge�J��-�ĊJ��O�D��$`Qߤf�H�R7j_�q,�A*x����طX�D�_���a�2��y�q��>m:�A9DVly��x��]���'\BU�8�	F8�f��C�|px��u���� �`yb�'��$�OP��je�L��gڰF��B��0+��t�4ybs��l����@�	_y�Y1VJ�?=�Չ���=k5l����-@\���?����?�*O���|���|�!s*X���rQ�ڋt0SV���	ğ��'eN�[/����9�#��O\fH;$d����gnV�M��B�'r�I�tvOR��u�8��(r��_��~�7�i���'�剬5(�|!�����Ot���)O���"s��#� ����>T���'�'q��R3�y��'�I~�EU5�:qz���^����c/����'$��
��u��d�O8��埊�֧u�,	)yR4���,Ӯ �HS��)�M+��?����<!����7�*{��{c���Z�X0��듋2�p7��sn��l����I��0�S���ķ<iu� �ܣ%��6���Y��B���d�i����'��'��J�d��[&i���B:p���3HɡW���o��|��ҟ��J&���<���~2'�57{�MZ�K.
1FԂu���M����$C3*��?�I��h��
�<L	V�G4�����j�-4�n�m�ǟ�H4@�+���<������Ok,ȊINH�)�Dqs�i�Y��2W�8�	۟����X��˟��'��,+5�Yz�D�2�_3:h[�(�2R������O�˓�?����?Y�#Ǎ- ta)K
�
4r�@��c�͓�?9���?a��?!.O�L����|ʲ��4T)r"I.E�Hp� W¦Օ'(rS���I៤�I���i �0I�Fs}�ej��|�NPش�?���?����$P�:�R��OZcO�(���
�p�LD�G,�s�Bpش�?�.OJ���O��Ĕ���O>�$̤HnF���㌂�<L��a] i.��o�����GybOD�7K��'�?Q����&��J�H}����fŮ���@!
����0�I�4���i���O-rџ(�Ȣ�N�^ZE�לEm ӾiX�>v��,q۴�?����?���Ym�i��%�C9U�:	�7�Q�d���1e!y�f���O����8O$$��y��I�i�P���7T�8��#�D:���J�j��6��O����O��I�W}BW��H�ϔ,=&��f���EA������M���Y�'a����8��-�"�8z�dԫn�do���$�Iݟ����%��$�<Q���~�E�V2��˕��>'��]���¦�M����$U�?������V4l@Ǆ�o��BKA�@�4�?!sh�7	B��LyR�'�̟�
?���*�0�
"䀊X�2�bA��?)��?����?)*O��p�fL+�P,��K,O.ꔐp��7k6��'T�	�� �'UB�'�P_��]�
�t%N�0� Z�f�q�'�B�'wB�'��Z��h����t����81�jJ�D
( �-݀�M#-Ox�$�<)���?���.��MΓS9��I�Ƈ7�ib���+݆4��R�T����P�	yr�ϢM���?AI؈C5�e��*ޓ)$�����[�f�'�����������@E�b��OH�Z��Z{_�9� a�+/$4���i=B�'��a�b�㪟6���O�i�w�%i� �A�dءk��U�Q�'�2�'JB�_�y��'���uRS��qe�?q!�Y��
�q�'FL���r�,���O���韆Y֧u�)�b���T-ȗv�2�KE��%�M���?���<����?i���OA��Sů�9�P���#M�C)�0Z�4X����i|R�'���O��ꓮ�$��31D�׍�&�0�!o iz�	o��a�H��F�Ih�'�?i����c� :��B�ao��3K۫Uϛ&�'�"�'r�ms5��>9.O&������n/9�Tͣ1#)2���>.O\x������I���ۗB.�,m�g`�Ur-rf�)�M���I�(1�R���'�RY���i��c�c��D��0�#<�P��&`�b��ޚ*g���O����O����O�˓+[n�0���d��8�>���#��O���{yB�'������Iş�(7
գ`�M٦���c,Ԑk���/��Iԟ��I��,����@�'���+��k>��  V�UC`De��HJ�`g�Pʓ�?�.OR���O��DG�\��$�5̞-�ƛ�XKV����
�AjD�'Tb�'nrP�$�Jɐ��'g����t)�U����t��3!�n��W�i��[�������ɫV),e�	P�d sdH5��r��u�ǧ&�f�'�B^�D@�"���ħ�?I�'{d����͕3r>t�""M��ic��ŜxR�'�������Oj�ӵX���h���7��g��bu�7��<Q���"��v��~��������@�iJ9�
���[L��Z%br�>�D�ObYR�O�OJ�O��>)n#��U���g͠}��эtӪ���Iğd�I�?�L<���Xċ�� b����H%E���"��iyh��V�'U�'p���B�(���2u�=ȃ� 	���mZ�$�	�s& ���'���O$h��˟22J�� BO�#�J���i�'��5)�):�	�OH��O&�R'�O"N�|+��\=��brk����	�HU�}Ћ}��'ɧ5���;sR�$�p-&i�d�"����'=�2�O���O��d�<y�A�v��IɆ��\ڶ�_�91�V�x��'|��'��
�
��6cN�`/Ph`я0e�h#�'5������	�Д'�Y֧a>Ɂ6��8e�^�'���l���>�d�O��O��D�O�@{4*���9.ҽl4��{�Ag��3�G�>���?y����4��'>���B���t!%m�$%2W�Q��M����?��-Ǧب����F�J|�r@�w�n�1����3�.7��OL���<��&^#=&�O]��O�JTR�/9:����f�y&<�%	%���O��dP�0���9�d�?��I[���Qcm�6 �,��d`� �x˸�!�iV�'�?��'g��>���&���uv�<�Α0��7��O����7����5��.���������V,���iL+L/�7A]��oٟh��˟ �ӎ��'�ܔ�5*Q�9�v�{ƅ;TbH� �xӎ骵��OȒOD�?��	�D,��@�#�_��D�3㇠/��@�4�?����?Q�B��g�'���'��䕣B:��iE(̃:6�Y�J�f�|��M���|��Of����s@���Q�s�҉�4�ߍ}��UlZȟ0��W���'e�|Z� l���mI(FB���GC C^9`�P�lb�'�؟X�����'Z�J6��
 �ذ�D�%��8Fܑd{\O���4��?i�}~��we�)�a÷��0Zk�Q���?���?I���?�.Op��6��|"�'�:?�P�cF�h�s�MZ}��'rў��I$A���I�u��M��	�4'�:P�a�3G���O��ON�d�O$�Dۛj�'�?���	�,���.Q��0�SƐ�?����'��'~��'x2�}b͎6Y���O��u*�M����-_��Z����h���M�^���i�L�Vͪ��p+*�!�W�&�e)PgI&Q��4`����5n~�� b]�TzŬN��9��gU<����J�AತH�h��!F.U�����(.���
^�y�Tݣ�2V��+�Eү��9���&l�Vx�����F��S�U��b��8B �k �q>��"ǖ��rF�ż|�K3��
�1)R��/^�z���O��$�OD���O੭�w�&d��Ǜ��0�&*^�Y�]
�iO~9+�ӷT���Ѧm�-��O�<�'��,{m�Ai�`3�CՀ)�y[���:1�j�t 6a9*	����ոO��������o�$At�`�`dҢt#�p�3ϑ柀�'�@����|���DT.0a�;j��w���=�!�D�>'g
�Q��υ4�j<�P�E.m�� �HO��OhʓJL�q�펠Z��b��Ѻr�V@�#LF�I�	*���?���?���h���O�瓤.��� i^�
(�8�@m��B�D����7<�8=�&��:�Z�)��'�.���h�g$ϟ��8a��
����C'*Xx"��V8��@��`�(q��v�Zm�Ď�3B����O�=a���M�T�؄`�5q��8I��׉�0>�N>�.:r�&	(��Er�i�"J̓���'�IZEP`X���Ā"xI���1�K�4�#���>:�N���O:�Ci�O���h>��r�����I"s�B�
�R�o"�j�pա�1���K0D/n�z��ğ�H(�3�͘O�du�efd�t���B�&;���VE�8I�桋�D#_M깻��I:
����O�˓N:�܁�<�%�]�'$t����2��P���T��w5[B��hb\e��N2�hO��Jߦ�$��4lP���o؜�(UmX��?i-Od���
Ԧ���O�U� �'Ǣ�т`�V8���D����v�'h"aO�WH>aK���H�~)ԧ�ɲ|.���)u��wnfИ�ϡorX�'����t�����=�M��i��1�����&\�p�Oa�q�'���S��Y��+��a��E,�l��,"D�h����(��DP��7m~��b:OR�FzbN	a�`�#d[�6���Pb��5�7��O����OR)#�Ʌg���d�O��$�O�NقI$<�G�I��xb��
p�HWI�?V���SB����G���O|@�'&���׏5�txg!�m
���d$[���Y���A��JB@�O��',�@�*G�>���f�dY��'��	�36^�4�N�=�� X	d����"�+���w�<�H/<Z 	I���� ���<I�;�����Ο�'���aO�.��9�$�=}�
p�WBߚ",.m���'b�'5Bo�~�����J�	^���qb *�0�`Ňel�AQ��$'��ó�0=A��O!��\�D	�`a�y����T��@���
w��� 7#��fH��ǽ7�J�<qé,n,��Dk�x�0�F�ilv��I��,�	Ο��'�b��-u��� �s}�X
�BP,g,a|b�|��H|���i�"Z2@������R.Ø'\7��O8ʓ,м(z"�if��'�8��š� ��  h��m@B�'�N�����'��I ��(!"�"�$�	o�R4��I���EQ���gE�x��<3��`Ç�ȝ[B��W�ײmf�}�[U�z0�D(�h "�V@�'#jY����w`�qB�؜��s���7\�8]��im�ȑ�Ki1Xy�GD�> +��������N����Gۼ>0�|	��O�cA�b� ��k�#�Ms��?�.��Ta��O:1Æ�E� �c����e`Q �O���˰	���`k�L���A�ʟ�'��i(y�f�`�^5Ucv���P	7��K�hK�/Һ!N(�3vI]�H�2��c
�:l��.t�Rȑ��>@U��Il�H�Ӳ)�X���׺[��("^�F�tc�0��`x�h�@�q��� Ü2���ё�!O@uDz��A37VQ�d���r�U���%�6�O�d�O
�f�1n�d�O����O�C6g	>����Gd���VH��]*����2��$��{li;��|RG&k~�H�! i���(غ<`� Q}�%ķd��}&��k$O�3�0,h@�C�p{�Yp ���M�P�iB��h<��,O��d �l�R����_R�3�����	�'��`C��ջX���І�?OM�T��O�Fz2R>!�'֊�2�5
xT �;F�<(�	�'��V ��*�귀07�f�@	��� ���򈅘C�mjd.K,$��J"O�59�-˨� �f*�1.D|�"O���kÕY�a
�J]V{@"Of��@BQ�d�tQ2�'�C}���"O��jGR�6�\��am�*N_4��"OxQ��݊OC�(STnI�R�qY�"O����I�ԝ�㞷5.�(�"OT	����,�0�d@;<��aW"O�Rc�a�b@1a �e'ȼ�"OZ���B6N��C���W�M�2"OFU���1!v��`A�8	v,��"O�����A0���`�)>���#b"O(�y��Z /=||����#���z�"O���!�פv,͠`O�-o�i5"O��!T
J�Y�̤����Ga��3"O��+�kϛ����7yC��`"O���v��3m��|R�M��6���"O����mq� ˣ-�(�$���"OH��/�g��`)�#�|�!"O$ձL�.w�X�ꑃK�<��S"O�@��g�;qpdفvI?}��ԑW"O"8��#J�><y�ATu�R��"O�U���O��D �M&H�����"O���Q`�5E��R�._�r�LY��"O���bO�="�U[�M��� �"O���Ӥ��_��L�@)�k$@��"O`%BjO�f&Xt�`�K�d�z��'ML��@�޷V���Q�*�D�H��n��qq��-3��x�
�>��x���1Q��$#'!GIS����	�$��9R'�8""�$�6M�q�ӶWKZ`���Vh{� �b�E�-�B�ɬi�80z¨ܠ"�B����ȟ.� ̘���g�(�#�ly��ԉ˱ݮ@�t���ũ�<��c�P� �T�.S y5"��3G4GK�(��L��ȩ	�yڠ8X�N�$jJ
�!0ړX=fD��nJ�EE�k�!�!!6J(��I�i��w����*� F�Y�,w�սe���SQK�%k���5m�20WZ�Y£*�O�m��șcyp({��S�0��c�>Q�B�����&�M�� ;w$n~*�>e�Ӎ�&?+ҕi`��Iۮ���"OҹQ�V�n��P�C��*���-�;upl����K(���S�'L�TTB�k޵�R����<��L�a�:����6�T����z��� ��:�����+Q6�d�D'��3�L�]\���a��ў�I���#�*b�J�=-Lq��I9O��TD��j9��2�%N%��ac���O�b��K��ځ���)G��  jJ�����?X�p@��G$�.m�2��/F���D\��m��&��#.H���&��*Nl�BlO7(R��r�B�I)V
��
_�d�P�bF�\�T��`�@,/�dHR%��~2����4)���;n�H �_0=�����0W�̅�K�n��wd�R��u�U�� 
^��ucy��F�� )z��� ���(O��i`����4@2A*E&�Ls��'D�슣��y�R(0�n����52�Fðm8<�A'̗0�����o��p�4�ԎӣY��}��T��}YC�ʈ>����i� �
%ߕ1,���Wg��N����r��2�\Ǌ:�ԟ�a0��ϧ3�\-:�/!@�=;"�'�^EAEK	R~�,݂Hw:����S�;l�8Rꎌ	I�,�p��9x�>D�O<%>�S��X�{�&�b^ޡRU �D<�,�w�42K���A�!�?�#��M73�<��b�q� �.���WK،t��7p8r1��9A��=��R1��d�N�vFDB���j$0c�ȣ�6�L�TH��{��s�z기�PD(D0���M�<I��P���\��@ +9Y������a	����Z�#-�U���jj8Y�,xͬT;��K�~ �򩖳%���Ӕ>�O\�sunŞ��q�P��&1@��ד~T.4p%�>�#ٚ?��ԃ�@�[� 9[7팑.����W#YhAŦO�O7� p�f�9�yw��3Y�l���K1Y� <b��֓��'����(��|:�6�pӁ_7e,����Ψ1+T���N|�+g	��F�[��� [��G{�RC6�m�0�+���CBC�g�8�>�P�x>ٲ�	�0/|��)I��D��� �߆|*Cɑ>e�TL��Q�J�$1;�e؇r��I�}*�8�iϾo0<�֢�!��t�'��j�����	�+�*-�^�9���"a?}*�� ���"�/�r ��ϐ>4 �(�'�0�s$,}�ȖJ#f���gȕp�
�ȣi��elآ0jF)m��]C�@j?�}*�*��qʖ�	�C���
�` Fx��^:�8�(���ا�'od$h)��3(�Z�ztM�xҒI�BN��b��1���W$��N� �εa5��;!3ڱ8,�8r��I�}���]��獰�m��B�{���WJ�N��ւ�E�nUQ`	љ1�4�2��'��=ҧEƿR�0s#���w��}����!yRt��1eT�qC�k��s@�4]w������D���`݉{�A�w��>~��!jb�'��}94�>}R��;d� J����(	�A�9%��AЀ$��9o!��T>p��|"t���<�uD�i]F��3	ChA�՘ńEl�q=������IC�@��*D%t4\�TQ�(JX<�:�����J��	������UM~��! ~B�(��Iv�)�d�,��<iU`K�`lj P��9���1 ��}%�m{qT*O���A� 8�S
˖W@d���'x��QD�'c֌���״r���rC��19�h��Ol[��,�r)�dgܺQ����R��Op����,�$>��ؖ��\T�`�-�*k�!���=�^�*��B�&���HҌG<RTH��w�ŋ�,5k����&x(RDZɚ��C�zޙc�$� UP�Z���)U*6�4��a�,W�b�REB�Ԯz��:#�]�i�8�'���qN��rS�pJU�F�H�h�؉�"z����6(j)p����0<�G�ĵg�@�TC�;'���J��(�0�Q�,1(t�b�ēDK���� �<5Lb�VHG��=9�d���C��B'�iB��:�Z�N�рX/jt�A6om�C��2�韲����IR̪"D:ۺ�;s"O����J ��4bܡT��1��~������b�����g�m�!��ǒ+f�T�RM��lE)r�-$���퉡T�����b�m �d�%����4[@Y˔CZT�<3�b��R�V���t�I�BQ��f�x�@�6�����'���T.+#
X��X6?XB��Qx[b�9BN�.`?�j�/�10�ó-ֽcd$��' p<��	(DQ�CͥF�ّ@-�>tI<O�ݱ'�J�=h�y � �5!(¡����J<X?��0��D��9��̗�|J���Q� ��I#m��f�7pHt<���	^< 5��H l�x�L�����	��{�h���w�2\J��a��C�*|,(�x	�'�ڌk1,C�b��ȗ)��{d�Ia"�|�!��;��h#��ܚVC2�)r۬��D3��6�¬~�Ȥy��%4�zT�����y��tzU��	�R4.��S"I�]��AT �P:e�fD�V��ś�A>���C���$��#=��
	7qk��mނa�̥�i���!=̤�a�;5Z �"f]9y-&�֝�}�.�qr�Ðk2��φj�B�o�|��	Җ1E��3a=�A��+�@��%e	3�>q8N�X�O�O/4��w�0� .Ȋ"�إ @a��'rH��'�0�cV�5�谹�Ɩ���ٰ�>aw��a�.,+�i&2L
ѢI}�-�y�Џ��	Y�Q�`��b�牟I٨	S�h�;Nb��6I�d��yJ�F�1�,�R�M�u(��BR���@bp�gÂN����Fy��U�^(��r���jH֬�"��U��[�mU*H�2���պ��Q�O�	�"~#�rB�#�����k�I��؇�	�Ȭ}# HSm*M��Q
 ¡i���B42Ѯ���T>�	�Ca����;�|�ʛcDX�u�*Gs����a_�S��_sd ��k:v�u���Or�!�X����½�Ĭ�Ǽ��A��Ҙ�~�+�jEg'��+q8lȂ��!g���2�'��qڔ��NX@�mP#'�Lh:����"�z��gCC�2���@Ɋ�c���h������O&
�4X��\1	��3?���W�H`��W�`�-��˚U�ɏ@��iY���k��u@��	)��P���h�0HY��h����%����'F	��i½v�L��gER����d��pX$�Ucp��q��/���:�U�����(7< �}�-�"I.��A��!�p��\: ol[J<a�%�"'�e�ȓ|0Hۇ��-'S΅PG�F�u���3	��=�h�p6�L(U��X�B@�\S�Hڅ�����q�~�(W��a�F�h��;��C���['�V-te�`��9Za�W��J"C�=7�$��"�\Ő�@r+Y��~B(�ui��)���;	b$�>a�j +�R��bj�:�����̓R̓z����ă2F/��'l&ց��n�-�u+K)z�!{���7
� �ծD�p䑄��#2�n��K�F$;P�ςÀ= ��?oغ�j@*�C����?�	�$�U� ��yG%�-Kr(�1�:���2���yb����B���iã�	x�jس+O6���'p�ձe�H�Ch�]��c�x�1�C-;���D�3Q�:l�%H
d�~��w.[�KC�y"@/$.~��s&K��4=AD^�!Z'ܶr�����%�Gڛ��Z"k��R�'s��C�@�N<,$D{"�Z�0~�Q%�J�vq�I1� 9��m��f�26�QI
�v*�O��4��s���"\/ڱ��
_�2�ib$��g.,-�	�S�? |���Ȓhw�ZeMO�;ĊB��(��-�roI�V�ӧ�L>��|�E�'o	�3�h����L�$X�iB�-$��YfA�Vi�1�RߍV3�IX�AS!�~��rx�'���H�'�Z�"i�&�X�I^�^PP�I�B_�4�c�h�f��D�$��5�k�$( f�����!v�A�t`�A��q��A�P� �	4�&���
�d��6��">W�@+Ōx�0�
�::Ӆ�|�	0D,:	8׍�1��VĘ�K��㞤R��P�Q��UCvn:��$�W'\
�
�����*���y�JUTq(�	�e̪=��	��`�7,T�B�¼�ƣ<�ӊ}N��ݰ�vt�J�~��tJu��!v��C��#ʽ����^���J��Y�h��<Gx�Ȼ'�F�y�)ޡS=ܜ��$���$��US�`�UNQ>�z��c�k�a{��H�`�g�LW+��b`�[�q���R+D�B�K��.V�y��	
�;:,�@�%D�T:��D���=6l�{� �
�Rqz�Gե��'����p��)T�l�*��!n�\��H��9�圱cr�=�@튂=�}���U��������RE	�2�8��c�Z7�fYi&E�p�� E��y��t5c�u�S���\�ph��΃�h��h4��pafy�ȓA�y��O�N���F��f�K�лg��O�̰+�Bt�Cd�-p�D	�'����g�Q��E�/ �B�t��
�,��m;��ؾ
H�������0ZeC�9Z�1���>��qKU&����I	���O�ӠGD�
~�- ӍQT]2Y���ɂ;��jV��E�0ȇ�[Kw��	���AL <��P���G*q^4�s�eM`���i k]��a�/9V�����X�Ʈ8�|ȳfč�P�
�<�|bP&W�,�6�RFD�W .���_l�<�AN�2e�Z� ��-po���� ��iX�DLU ��4pt�rM?��C,��kOJ(�%G3(�X9�9%��2�>+��l�� TS�
�#Q�U'�fq��'ߖ�?1�PR5Xt�b&<Oġ���+��5��!  ;{j�1���
N�����@�O�����?1�B���f�t�F%єD�44�	"�N��xC
�g��	%i�>p�A��B���ɘ=��I�T��zb�����(P2��ͼc�:A�@A�"���%"O
<���^)n-����E���r���R6��<�"�X,5��;z2�kV�OX�<Y��n#�8�N���&M�3N�W�<	C@"�|X�gI$|�L	�`�W�<�&�\�zsМC���-1�	�rM^o�<��)�#F;J|�ă"�"�AM�k�<�%
�
D~ � �
i��i�<�Fmԧa����@P�Q�a���h�<)Q85�Q d+ۙ-i��J��d�<A�!�� ���gJ[�#�c�<�ŋBic�qK �@]�ҩ+��]�<�g�>G��}H�AAڠ<��B^�<!�l�/�p`�	)T~~͚�O�<!u���4�ㅫLp���TS�<ل@O1iFtڦf;����_P�<٤锪9���	�q
��Df�<I�F��!E��Ф�!	д9���K�<Y�h�xd�F�:M�q����<��٧H��3�Y�SԤ��N�<�$K��=�XU���z��Q�4g�~�<���;��\�㉈u�z����a�<Q��Ѹ\�M;���!�H��%�Y`�<Q�)Κ~���U.Yr��X� S�<���?Fg���G����4u�<��O5<(���[#{k�8��͑G�<��k�<}l��x��5����ɝB�<AVH��	0�T��`��u_9�'j-T�����Y#
��)��+ˢ|&%SB/"D���R�P� �`�bA�^�d^�q�
<D��hB@P���E_��qH�:D�ti��I�N�|	3��(���aaC:D��x��@?on��q���2B�Q!&:D��R�oK�#��Sp`T�6���7D�x�3��	X�y�lG3@<,!1J6D�� ce`d$�q�e�ЕX����U"O� ч��7�
��WB�{wd�HD"O����)	��|hHѠتLe�u;�"OR�XTM�jx&�ڛ$O��E"O��"��$�R� 6��"�"O^�$(˙���P�����"Or�N�; �#��^� �m�'"O��p׭��7�b@Y���3L
���"O��I�̃R7��M2H��"OL��
}��gk�>e��5�S"O��9�k�//�h�b�*�Jt.��"O,4�C*D/p��4s��-�Z�;�"ON�����{�������	��]�A"O8L���
��c�����(�"OXU���
$�~|�᧛�"�2MK"ONt�`h>�Z�qQ$`94"O�(�`a
<�v��U(�t6
���"O�LP'�D2�Q{��շJ�\ :G"Oty���<|��ֆ �t��TÄ"OX�#i���F���DC7�$��"O�=y�;*�l�S lI8�"O����([)tܨő��'@� �1q"O��0���:~���:0��15�!��"O(��웜պ��bk=Uߒ`V"On�����!4�Z5��?Tۆ�!0"O�t��L��t��]�La�"O�\�&��q�|�yr�nT�}rg"OT���)`̘���-L�49�]`"O��KH�n��	�c4@I����"OR1�vd+IG>L�v"�8_@�D"OXHHV�M�@8f1S�P1"ODc��*_a�{ա����-8"O$�as��k@� �B��g��܃S"O��r�K3�$)VN׎�����"O@i��H2��"���=r{��!A�'Yў"~
�"ۮ^�x����= 
Ԥ��y���F�0W�ءಠ�&g�<�y2��<P 0a�c�i��-G��p>�O<�b螐qP`,0��xT�)��	Oc�<qr
S.:R�q���*��H�Ec�<�B�5Gt��@�L;ZV�s�(�I�<�����~E~a�	#C���D��i�<iT��^��T"�!;�`��Bp�<��O�:
>6���CQ ����2*NS�<9D*^��tz��Y�2'��G��S�<є'Xx����.)��	S�G9�yr�]-����䐏a�n�P�",�y.LM�A����a!:%bV) �y���( /�� %Z�f�čÐb�%�yA]�.��pMߖ2b�I�#Ļ�y�g�&���A�-��D��� ��yrk�n�VYCЫ�%��0o���y�B�?"��5 ���_-�y��6	�$�aeJ� �^��$�yB@�s˂�H�mT�'�Œ�
̈�y�IHԂ���p�D����Ȳ�y���`	�}�"��a�:1²����y� ��.JYx�E,
=�\���J-�y����b�$	�Ĭ���ɲ�y��Ay�8��:����˻�yB ���b9i�&��tb���O��=�OwV,��CF3#&B�P&hъ?X����'k��d�L� nh�2Ȅ�5�F���0O��;Z��$z�C	���8��"O� ��k K��s$�-�փ�|��9�"O�4PV���?�����*F�ٔ"OR����2lFx��GάB~��"O��2ڞ/� c�4F�=j#"OT�BcC��t"�%(��1��(�"O���r��*�� �Lޚr��5S�"O@�r]�K IV�M'�͑�ʔ�yr�ŝ!ʤђ�G59�Ds$I��y"`!f�4 (v�^�2HР��L�9�y�
5��y��*�="�zL �!�R�<�R"Z� @,����2��iR�[H�<�UDB.k,��	D�ګ=���� �B�<�Y'��1#�D�0d���y�Ђ �>�[���r���.���O�*����qFx �v�K�Kt�k�)�f�<��">;���r(�;+�4�+�JHz�<qA�^�`'�.:Z��X�B�w�<iWL��	�2C�� ��l�U��l�<Q���7i�*R$��Se����\`�<����r���rE��'P�,��`�<��-/:�*�Y%�����M[�<�FG�蜝� �h���ʕY�<�
΂#��i�7�X�V�hYrԢ�K�<Y�� 2��Y#M]O�)j�cR�<q��N�8Q�a`�	�H�iCJZQ�<ٵ��>O�Z}a�!A*V���B�<�����p����Lp�5 t�]{�<QCae�BH�Q'C?(�10��Pu�<A�
+� :6E�2*�܁����o�<1V��� dq�E�U,V���S+_k�<��ƏT�V���F�x��Î�q�<I�%S]��E1p
Έu��hbD�E�<�'��!X}zV�X-!R�a��JC�<��_�~p-��DЅYliyU�<ɶ,!/"ڐJ��_ csjѩ��}�<Q��0u ���Ij�"yI���x�<���/	3@�* ��P��)YE��M�<9TbG�C���X�I�!_�*��~�<���^"(�@�(��S�>���}�<�!�$MJ�b��K�Έ�+�'�N�<i6��3_:�V.�}�,m�L�H�<��J	�K5059Iʺ�~ +ʓ\�<�'Eѥ}���Z��N5!\����W�<9�A�Er��Z0g<�Ƀ!V�<��ΈS+
�е.ʖv�Ydd�P��2�O�Q*ٻ!�~�t%X;~l��ф"Od"��	�d]�t�_c^��"Oܘs�I'�:M�3�ۘ ���J �O~�=E�$��lU����܂Z��ip�E'�y"��N@Ԁ�@�Zu�r��L6�y�̙�S��V,�h݆�P���y��@��jvO��`�(]Sʐ��y��?F ����ϖ�0�v�#��0�O��"�^�|��mՀ#*�6�b�"O�})������H]'2�,hRt"O���e��>C�@��ӧ��=��|��"O��r����|y�Lp�)�dm0�8�"O,L;P��}�d�B#�ٌ4`�A�"O�,Zfe����#��\�.J�1�"O��i �EU��a�o��W.��q[�PE{���ӃU�a1��-\���'�NdK!�D#k�dS �X���C��O.!�Ė�U*ȍQǈ�
6l�{Bi��*!�D��j�x��$�C�f�{R�� [!�� �h�v#	$��	��gJZe�%b"O@��g��1TPb$Ϣ>~���"O�M�C��8�ת۶@Gz�H�"O�|c�o8W�:5��M�M ��3�"Of��%��g��䳕(Ӹf	JIf"OP����9ր��'8�(�"OTl@�MA*{�KY3hJ� 7A�6�y�mB�
�)��[&8�Ca�ǥ�yB��8q�&`ZGƃ({��[�̕�y�Q�#8R�wbY�$���y�G
�yRL�	k�q��n������y2�n���*�ʅ�5 B0�$�yR+D�C���$�.R�(s���yc���vLU8����&�D6�yRX�|x<Q��X"2�(���U��y2�?"̅��=v����ujV�y"-�=0�X�J�(['@�`��d̄�y�L�P-8؃��țK�*ň���?�y�Ť]*�#�*G[�i�fϏ��y�@�-�6�Z���)>h���@�y2'۩b�n@�BD�~�ڱ�
�y"�P��N�
$H^�u��x��]�yrnO�X2Tl9�#	�E�4{Pȃ�yr��4���s�*�`P���W���yrL7EV��[b�*�JdBD`��y©ѿn��{c&Y�F���ĈU5�y�Ȇ�B�6�0�K��n�ԍG�y�(�0T�v���f�>	c�HrVm<�y����J�$���Y�-T�k#V��y��"7����\/rBH��K2�y��Hyp�	a���TAV��Tm��yr��C��i��	�!Ki����y���{�`�B��o�:��E
!�yR��<5J~�b��&(�!����y���d\�����	�\!ҲcY,�y"�]u������~�0��q��'�yR�˨F��4Rw��:,߸0KfF��yb'A�*I<)1R�R�Y�Q�5���y��O_��D�E�C&��`U�-�yRk�*$�*�����ZA��6�y"鄒5DP��g
��y��D�k��y�
�Ѭx%&K��>�Q$��3�yb���$��]��G�w��X��ރ�y���Qr*t���٦p���Ai���yB&�#�X��ffΓa�� ��=�y�A�<G�e8�&�D�X i�
�yr$�[�
��Ԇ�{(ѡ�e��y򪆤f�X�H�g޺y��xc-��y��h?f�	��ԩ#x @%�y�(\0v�~5��/Ý7��B���yb��<-BX���_%!����!�[��y�GH=S�Ѐ��Yِ1cA��yR,Q�\�FQQ��_�}�f�h��ǖ�yr��&j�P!�d-Bݖ ���%�ybI�1���Ը<��� u���y�@� l1����
ڣ>����
9�y����T�(�Ka���3���`���y��|D����.�zek�'�y��3b�i�K��$�*�k����yR��]X��	$K<y&<� �N�y���u�`�qC�~�����J��y��!~��3���:n��0�ɵ�yB�V�)Z Uak��hC�\�&�'�y�ƕZ����IL#_�X�0����y
� @��1b��5����WY*9|=a0"O}:'�Y5J�K�,��Р*Ol�Q��?o"y����%��'Ǵ�2�<=��a0����jp�'lH����5���&#ku��(�'e��J$nH ִ@��OJ�^�b�'����چ?* �(Z%h�����'kX���\���Q��G�6rq�'���5$I,
I��敉DP����'!8�Ȗ�-�`�a�K�9\���'D���聙?!D��!�U6)��L��'YH������M���<��'/8�s�e̶@����w�؇f�� �'$�TI1E�C�9�m�R�c�<�
ӡd��IĬl�na�r!c�<A�k]�y������휟^!�d��f����(G�	=�Ļ��R�6U!�N���!�%M.��hicM՛F�!�D��!��S�&Z�f���(�&S��!�$�f�RD�N*g��yAsD1J!�$U7S;ʱ����M�n$Q&݁y1!򄚊m(�pAKH�Ep�i����')!��O�=k���=R4D]�"�s!�dR������TL�0���Q� d!��T.��z�<d�*�!���!�D�,-�&k�C\�0��T�����u�!�хa���bL�8T���2��&k�!�K6H�*�F��-$�m�C�(r!��U�D�����[3,y��(N��!�DQ$�ѡ#B�B.聲aܮ�!��(^X:��Y�c(\����LX!��L�%Z���aDA�O���6
�:5�!�Q|Bt� �%�P�iոp�!��M�j��lX��'\�pA��� {!�DZ"����Rǖ
�f�uNީ`!��T�8b0�<O����U�!�O��515(�� �N��[s!�d�N�� �%�셹5�NgS!�řH�쳢�A�P�݉��E�+I!�_���xq�[A�T�q4��:!�Dݠ\t��rǇ��|+�^�s'!��0��Y���~�ɺWMD*Y"!�ā�u��i�eHO�ʪi!��S�h!�$% H�K�̈́\x�b���o2!�U�I>nuX%�ѡ�PA��E�&B!�dW�%�I���SE%��nT�M�!���%I���#jV/6a⠢�͚�Z!�ЈE� �I����L8ʕBBl�1$!�$�|#Z1�g���i%�5��N!"f!�$�N?�Yk�e�02����7i!��8�
G-��
���'�=O>!�$P=��v�T�.	\0�2&J&6!�$�?�1��H|�d�Gj�t$!�X�
]�,R�A.Z�*��/��ko!�D4W�*u�qg��\�x�u�V�0V!��f�8�7���>L���F�!!�[�{��r���Z�{s�D�s�!�� �!N����zmB}0p!L�!�ڵk?�S4�HT�Q�/_�}�!�D�ݸh��L��2��1�!��:�p�����ΤPQ��)�!��,w��.�	q�4��4��_�!� xu2����u�����@�!��]�u\�� jX�^N9�QCQ:F�!�� �L3��B1���!�&NrL���f"O�Y3��S2 ��36��O74���"Ov�4�����8��! �"OV5�u��a~�!�^����"O�Q����\M�d� ��2t�zYz@"O�9x�&�?:00���̢H�5�f"O��!A"�f�q�B���f"OZ�J4��oT��� $~hx��"O��Ѱk@0����	!
9s "O`�)G��)8��M�'�&�rU"OD�j���+%���B��. ���w"O�|�3��:����M��@��"O�E�c��z3ޝ!�֣��A�q"O2�(Q�z%�����^z(�	�"O��C�,��z��=�1Q�XW"(��"O��P@�ǖ���6'TQ��y�"Oe@�ԕ5�᳃��661�"O>0zf��bP��J����r=3�"O��#&�V!s���b��j┥�4"Oq��O!w휅�ӆD-E�F�*�"O��k` ��;�8��Œ�kG,u�"Oh1e G� �cd�%I*\d�F"OƝ;�/�,f�4�e唯=���6"O�l�fc�62��9U坯z�NIq "OP���fؕQN�00�i��2pp
F"O�<Q�	�O��#HU�;�>y�$"Ov���쑑}���G�(���"O4������@d�M�ef�zn"��U"O`+� S>%I*�#�V/`h
T�R"O��&�A.�z�a�$�Pe�"OJ�ْ���l����Ά2��)��"Ol��ׅ�� �*%x�V�J�E�"O
=��!�;n�%kM0<|�s"O:��A�����!9W�H�"O�Cdትf0X�e��x�\��"O�q�A�[�j�T����|8M�D"O��E,J&z7� �$�ҷZk�ia�"Op��c������c bF�D"Ox��'�ޔn�����
Zn�BT"O���u��A�P(Z���Z$�Z1"O4�z����2d
A��O��[�"O���`�(Y�n|R�
�:(�y9�"O0)��9/F�X��A�Q�^�;$"OV���>t>����ߌ3�
P	�"OΘp�ą#9l��CA�l��l"O��P&O�8f,E3E"��+��0(b"O��oԎyq��y1�>	u(�"OB!����+F���*I�B�A9�"O�I�uD�7����$L2�h4 �"O�Q���.����2<��jt"O:���Y>m?V�*4��x�@ �d"O�uR�$���dQ�	J�� ��t"Oȁ�0]6sSXe���۞Kj�!��<}v�*�-r�*ٲ�E�.>�!��#�D���
��f���0��L!�� Q5
hSߧrа⃁\�=�!�ā,����t
� [�=YcǛ2M>!�dԼ*,9�vb�k=r8C2F>
!��!Q#����0I�
���K
5�!�$$uy�I#Ўߥw��ؒ��H�!�^�|:��%[����M4 �!�T7XnP}��k���H�kDY?�!�dZY�����@��f�l8��:R�!��*�h�� �S�kn�R�.�1
�!�� ���`/T�3����˗�?ٸx("O���oةr8��I�$^�"["Od5��@@y��锟Y��r�"O�L�C��)�Z����hPy�7"O��Y̸t�\a3�A�7��3""O��1`��'t(h""�� 쪅�C"O��AW�I4 �t\b�炥b����O����M�>��R�9i����-�!��
�3����M�bJ���� ?����9�g?���"�(d:��O'2��TI�<Ya�[%]��M�ej�'3ŐMc�A�<��X=�F�z�
�.T}QrW�F�<���_
1b����,N0*�ɣ�I F�<a��޼d	��RO��A*P���Yz�'�ax�!�6PV��1g�eዛ�yRl̖~�vp��(�)d�"a� ����y�C��+��4�&�h⼨�[-�yR��R��:�̠{��m15�1�yR� 5tG.���M�<+�|������y���tVa� [;�6��RD��yROC�~I��d7�ʰX�끬�y§�G�f$��+B`�(V�Y;�y�H�x��� 6:��5e]�yR����!1P]�hgXh�d ��y���B���5ش]�X��t�@��y2�ۉ�0�hs $�0�D�͉�y��ȭ9u�	���C|�X!z��y�+�=�>	�"�HK6���IB��y�C
.V�1@�g=1��� ���y��K�Se&X8$X�vO�4���y"d��Q����#�0$6���F�0�yb��>c��M�a"_�w|��	���y�,�(K\���  �aD�Г���y�d��ިK2�`v��h7#F)�y��G�)��Q6A	�V�u�uF�=�ybe�{�`i l	eJ�<�wHI�y�i�
&]8������k$,y�GHN��y�S�[�6��`� `��A�7��;�y�a<3�BP*�\�R]����
֞�y��G %v���7L�� ���V8�y�Ț39�b-h���D^�̢��Y�y�˫T$e���8gl�����y������g�C�]�u��gN
�y2�;=���9���ר�"��#�y����v�P��EU�C�\���!��yR.<�}��'���^aC�����yD�>������R���NX�y"��>h�����æ�V�C�Ց�yr��J<%�� �x�.����y��T��LxR4!ƀ}�p����yb���)�Ai҂
# ET ��-���y�o7Ki��1����qCp�@G�D��yBLM;j��847`��SV��y��G�=1t4 �0]p]���y2�6{Ô�0a��!x����	��yB�ڕ.D���6�N<?��wd5�y2Æ�3c4�bSÊ�d�ē6�ڍ�yH�,)��ڣ)�i�&�ۅ���yC�P4�[�a?x�H��1�y҂V�IdE�vKD�"���j�m�y�mІ+����B��"�튵�D��y2�܋C`jm�wɊ
���[=�y2�ذ-b<�7�L< vD+���y�!��N�� ��	�j�fV��y
� ����G+l��Xj��J�_M�	"OV�A��; P��� S�qEH��"OH�ڢ/Q:��<�P/ι.[H��"O��cS�B��r(;��{;�mR�"O@�5.Y2|~>(!���O;-��"O� A�
��w�ZY�����`��"O���ޒn����a���I�<�ʵ"O�J@.O[�Y7Iΐr�: @�"Op��rFC�Pj�V��:���T"OREJ�bē��I����T8�"O6����j/&Lr�v��b"O潀Ơ�Dͺ�S�#��)^�܃T"O��#A��@՛U��Gѐ�"Ozp�ƉB$�,,J�&r�B"OT4���[+*:���	��a��"O�0�I&�JI(C*lxy�"O6p(�,R�dB�zc�_[����"O���^�^�Z��6A��O\�AZ�"O��@�W��:`��1e?��"O$��#� 2pNJʖ�#L����"O��#p#�-.�йP �E䅻�"O��EÔ*.
a��!*mH�"O��KdB����ƌ�h���:�"Oȯ"Oc�i��f�b]�����TS�<���,���Iv䗐sv�a��g�<)�%٘~���b�H�N� �K�$I��G{��iL�m�|�1mZզ�A�+�t',C�Ƀm;^����٥àT��F]�l�C�(o9�iwb�\2x��"�Pʣ�9D��"�&P����K�,(�,2D�$p��ޢզ����B<R�;q&0D���G/��](�U�mk���@�,D���%`٭i٬eňۉ$����@�O���(�$�|Fy2�6P�`�a MPy�d��y����#ƨt����#j��H�M�y�ą1J餬p���*h �h/	��y���=w�eJ�"!-j1�͍�y�j�3$���)�┻g ��QF�/�yr	.��M��B4Ȯ�0(���yb��C��Ѡ��Fw�9Ë���?����0<i��"9�zո@�X>WH�i���L�<�֋D�G���B���96���dɊI�<Y#(vY���@��cdjl�<ic��iD�`���8Z�q��6D�����)Ɔݓ�Q-��+ŏ/D� �� ľP�ХB�a��yCd(D����!�
�Dm�t��#5�Hho%�Ip�'���G��:E��K�� '�ԩ]C�	�BD�k3��Q��$��˒�WB�I�<���ꐋ��"����4y��C�� )�2���%J�7R�PrJ�$�C䉺~F��re�M�<l3���$#�C�	�^�@}3�fF	�6��7�Gq��B�I�z]��	��$y6��*E�Q���O���U�c&�vՠ�s��H�"/ڽ�ȓ�8���%�4����Ջ�/A��D��ai���B ����G��(>#�@��Q�֍5'�2�t���C�,H�t\�ȓx�����N6Y��A D��)V}��ȓ&�H��	Ə�$�`���%(b
܄�O��D���RHp
pG�U�,$���x~@�
�^i���ރu�p9BeG���y�%����ma��;<�C�E�y)Ġ"0]���/�.�꒢/�y
� 4��7�A���k5��97"O�I�q.�,�fd�у�,F�Ӓ"O�Ȋ4�=;�U ��:_74�s"O� 1+�F�<�Z�RJN����]��?y���?)*O��ӑY�X@�OG<�� �̆%h�~C�Ɇu�J:%m�Q��b���
PC�	3Y#�)�)0q,���o�oQ�C䉀6h �$ �%��ђ�B�>bt�C�ET4b�,M>tڽ�O$żC�	#4+��C�	+��¸M/�C�I��l!�Fl�S��ue��?��I�hR1�2��&`�f�L.@+!�d�l頱{�V?5�(=���|�!�dX�w��!@��
_?�	��ԬK!��?f|�2х��O�y�)<% !���d=��2a72Dc�(�:q!�R li\��+�r� ����o�!��X��ęź0�0i��l�{��'Ra|��a��r ��R;��Kv'��y"��]��e�i[\*�{M֐�yR�0[8X�õ{C�@A��yB��0Ѳ���V��������yBԤy�h��Ń�#��iʂ����y�#��Z �9�Y+/�&E�vbĤ�y)V9	|r��b�D�*���3��<�yrm�"Y<�����W�#������y���Q�r�30�Z�K��5YA׳�yKV�7�`��6��t�N�i�%V&�y���%�"Đ��=n9� �h�-�y�'O) e���ǬR�{�x�S6��5�y∆�s�"e�gb�m���U-�y���*����+"n�Mi�ǒ4��=�$6O�m�℈�t����L�%:wVlqc"O@A)��UO@<h�dJ͑g`�A��"O���UE��n˧SyN� ��ǚ�PyB��g�-�h�#R(�����d�<IծY�����ץll`j+�E�<�r���P�5��d�8�h�ɀ��X�<�q�߉;�*�[�Ө\N��T�<a�o��2\��nQ�z�-�!��S�<ᦋU8���ߟw��p�J�<y���$��|���S�sRU��C�<��D�Y{��Q��O^n�pc�|�<i���>\����E,"hU�P��N�<�U'�&$��D�4F��98��b�< %��9���Q�)���F��`�<)�G�S�q*�KV�)�!9@$BY�<q���b��E���ۣF����R�<��FW�+���j��
�
r�@2��X�<��f��(�U��ɔ�}����i�<���\� �Q��	V|x�B��M�<Qd�\�1�(uf隄hB��I�^�<�!�#�h�y���E]v�I�I�s�'���>�ƽ�*�!%�e�&�x�nC�I�2Pr���' j-I���,�HC�	�Q[�x��1D��1��)]�*C䉝%fuzW�B�;�^-��d\-m�B��1
.�<��i\�hF�C��z�B�ɠ	@>��ŋ�;�4%ȱ��v�DC�	�i�D��Q4*C�@@Y�~J�;�I��p��}�'Q��P;�EQ3����.G`[��0�'��1w�xLa���$P�����'���D� 
�"�	�����z
�'�i���ۃ�~��p႔(���x�<� ,E8��R.r��E+uŎ+c�R�Ц"O*0���&3gđ�g��px�"Oqs㦟��Xyb%�� 2���6�'�\���ȟ�'?)�OnRxCE��J�l\Ӱ���o�@
p"O �i3 E�U<��{���0F�a�"Oz,qݧ}�L��R�۶5Q��`�"OZQXJ �M8J%��|H=)3"O�5�RG@���d��ש}0��s"OP�iP�س36���(M��@w"Oh��+�
e�DEt�g���1#�'��'�2�,8RJ�Z�l\0	UP�9Sg\?6L���e�ީ��EE�hƭ��?&���&�\P�/��X�`�	�[-���ȓ] �"`�޵{�fE!�g�6_�q��@�D�X2h��^p�%�7XHM��aV�:P-�0p�T�s��/\��ȓ0O �u*�~���X#c�$��Iϟ��<��p�X�P%�2N�d����[�<A���x���~�V�� jYQ�<y����V��XR����r��S�<�ei.)o2���*N�@.���Ij�<������H�xw+-��)�d�AB�<�W�E�Nu.92A=L�9"�Ȇz�<Y&�I�F5�����j��yx�x��T̓v���RlM0"�Ƶ�Ŏ�$� ��|���ևW�1X�a42��M�ȓad�cS˕+	�:�)T�Aقe��ck��a�UO�2D�@�Q�P8��%Ȯ��B�ԔKYB�)�懗��ȓe(�Z�-�{��ei�P5���ȓ���ȴEZ-)l�:��{E~!���韠�<�4%B��c	�
�8��Nh�<QJ��O�`kŁR	'�XR �QN�<)��C�W�p�E� ��xL:sAR�<)H�R�R1� +޿	��4���D�<A�������c ��bL9ˁ��x�<�PmJN}x#�)˵n] p���~�<��-M��q�p"=�X�`�)�bx�H�	y̓L8"L��f��l����qoZ��ȓ-�0���JX�R��h{2�>7`���ȓz�tE�1�0��0ӳM�3{��Є�}�D�kQ�G-n���a�(L�qh��ȓmN�و1�߁}�Jܻ��̰G4h�ȓ
����) ��Th�26��ȓe�-����'b�4ků�	?��4���M~�+��$��咫[L���H�#�y��n�<�.S��qkɅ�y����n��=���@j�������!�yB���..�) ğL���X���?.O�O?uIԇ���(;1��"k
���NL~�<ђE\�k�
��� M�`��	�6�
_�<1a_�	�>��B��i��Y����X�<��i߯Sa<mQ�ƛ�cǈd!�X�<��
�hrʹ�,�v�y�Ҋ�[�<qbÇ�C� ؤ���(�փc�<I2i�l*>�!6��a�i����D�<	��F�aĐ؋g*	S�0�2�C�<!�eИZ�T��NAXb���M}�<��}�rp��� `���1�z�<a��.��T�� F>?~�����k�'���'�>�p��<�,q�W,Ҽ.f���(7D�|{R$�,F����:$ �U5D���A9l��Ph�\�_	�5��'Dў�>�S�2c  �Jc�*%.��D<D�� ���󂌐E��)@�(vid��"O�)H�-�"h���̃�na ���"O���+S�(eD���g}�=16�������J̧bC+#؁j��� ��vf�0 "O|��E�Dv�Vճ3I*6L�3�"O�	�ԥ�1N08�摪W�A�0"O^xⲠ
"��K����V���+�"O�8�փ��JF� ��O�fI��"O$�YtK��\h(�0vl]�z ���"O���")%H<A�#(YPGT����I�M�d�g!Y�Qb(�h�C߀%�C�=��� u�E�-=@�i^v�2C�I����v*#2�r$B#K�#D����hOQ>���Y"!_N12U2zW�}Y�8D�`q�$�-(�b]Ç)��PW���W""D�l��#�!9��A����tn�iw� D�Ҳ�3[���j�� F�
��>D���䏒yf@8�~cحpA?D����,6d�Ԣ�,]{Pz�/��C�	yR�%8��B��bP"�F @��C�	�P��}��O	*��<��%�#0��C�{�!��jU"F9ZP��E� G�B�	!�`�B���R�d�W$D�E:B�	�i�N0��C\�Q.�3BW���hOQ>�p2f7?���� �#c�f���9D�@�� Ĳ�ޠ�U��&}�bB�$#D�4hd
)�$m!��A)4e�a
#D�D�@9p�b�ؼ �lA�a'#D� cp�S�i�-k@f�kJP=�2"D���W��xI���d �
�I�>D���7&�XE��ʖ�1���VJ'D�+Ĉ� >��丠#�3y�Q*�� D��j�Z�~Ѓ�d�	Kp D����k�65|v��2�8/���Q�(#D��� �Y�Υ���S7s�`p�e� D���q������0�((,,Ĩ�D4D�0��,��؁!�,�;9]�s�K1D���#ɔ<K�Z�*)�%lj�L�Pm/D�����
S���!�S�Y� !R..D��yeMΣ5����o�,-}&eSAA6D��@B�$K�j�R
"�$��%�3D��GnT�K�$��,YX�RT�/5D���'oW#.(�SO�;x���2D�<���D432 1X�T 3���Sc2|O�c�����X�~�[ �^�F.�@�E2D��b[B��Z�CɈF(�F;D�1�ۂO	sUo

e�x0�7D������j��$�e	�Im�Ec�*7D�|{⨔55J��M�<x��h�M3D��A�̄I� QQq��$[\����5D��[ʍ���uH�Ѩ*d0%p�&5D�pbë�~�X.��Y� q:�.D���t���vQҤѰ��Ӹ�a�%-D� ����4*L@�b��+^�Zi,D�(��h鄀CR�� <��a+D�$���hl��7	[#4�85Z+'D��6���tD|uX��>/}x@C&%'D���2�H�q� �i%�|���hG
$D��kc)!V���AF+b���@/$D��2�@�����rF�n�|#f�'D����A�n��}�V%R�,�vT�%+1D���t�A�#6V@Ĝ	lRh� �/D�ԺS�գV�>�yR��9�<q�,D�H�q`�;�%�c�?Gp�8aM&D�� �dF(��Ud�H�#�"��#f"O���Bh�C<>��fl=_�صK7�'���_����#�)1�0�:��$D�L ���)
�|���\0TSh ҖM!D��b���r��"M]6"� �+D���v�� ����g�]>z��&�4D���a �YR%1��B;6�8v(1D���T�͋{uz��$/�60�0%D�tȗA��9��b��C�U�a�Q�#�����z�k��N�°2��'���"O6���h�9yu0�"��@�[�|�`"Ox��R�U�d�$z��4{�R�!�"O>���k�mgJy��C5<ta�"O�d��k��{�<�;LZ��"Ovb@�ʾ$J���KΪeH�!"Oz�#�b)U���s
�p�1q"O���%ć]>��Z�ō�:b����"O�Q��#��I�6��X ��v"O���"��?%�4�@w�4+��[�"Oi�Bg�<5�P�bA	 u�"OJ���ܠ[e8��b�O�p�H�"OPђE���42�Uw��(�W��!��10<�,��
��p�- �!�5y��!U,�9AF�Dq��]>#�!��)}�좥b������s�VQ�!�䆳
�$�k�Wx���	ɖd�!�
�شpA��-g��QTG��!�dG��e8M���M�ѥ�z�!�׼h��"�S��P����S�!򤚮ca�m�3���/���q�JҎ=�!��_Y|c��A�:�����!�$�vzI��O	"��ă֨�T�!��5n�x ���V�YSЫ�&�,E�!�D\�np( ⷠ�+&b�9��*޼	�!�$P:����%ӒV&��`�#�!�dТ@:�Xȁ�O�R�52��4X�!��N�%	���E��Ā�d�s!�č�)�z���Aȍ�p�+�b�p!�d�)�,�(qċ&@jL��a3J�!��cB�\br"C<q�����	�!�D�x|H��gۃUs>ũ��X�p�!�խ �.��uZ���i^�"�!���X��d�"%�p�FgC��!�&>0�0seLʹ4������X�!��ۣ0�X�6�]h�����׉[�!�dR�k{�A�ElWlZ�h85 ]�!򄔻 -�д����F�Pᥚ<I�!�D�m3.�RɝH�ച�T:!�dT1KN:��g�/���[�H]�!�d��N�Ѝ���!��愷��{�󄁴n�`�8��٘q\�[�̵2�_��%�"~��\$=v}�҂(83&1�`���y���1^L���.���dD�B	��y�F�3ht�he�٢��}�*��O��!E�'���!����d�����-oTL��'�T�qU�<<f!�ǀJ*�ź�'I�Hx�d���5�Ǒ�H��{�'�̑*�C׀4�p�����	�nY�����'
�>��v/4��̣?&�� q�f���#D��/9͌dZ�
ւe?��!�U!�4l6�Fɚ$EX���aa�[1O6#��'�<���5.P4:�◅`���'Ѐ]!�nي7�Tm�@?h(�i��'%
b`��"dQ�7�d���y
� j��Ă�� ��Q�PEV�l��c�'ў"~bQ���r9>
�iΠ"��3PO��yR�W0�l��#ҿ(P�� ��;�y���Wwhb��#S�,�H��Q��yr C���<�'b�+Qn���̖-�y"h�5� �ZR�mℇ�i��ȓkJLuH��T��!�JC������ǟX���'�d���Qؽ9���rq��rjfz�* T ��1%�CJ�ZT������􄎰C�	f�j��ȓ`2��b�i!L(��cGbȅ��I+�
��D;�!�0��qA���ȓ�d�f���C,a��O���ȓ}�Ubc�5"Uzx+R �@�.�Ɠp���&c�F�ZEhF�*j�\���'��Cw"ά��#�Z�P�'&\Q"��u#lXTI�_���'"�B .� w5rӁ��}�:�'������M� ����r�,ElJف�'�����ÝLq�u�1D��&\6���'!TT�\M�5s���f��'�
���j�3�&1��Er"�' �E!�O,6q�c�	����=��'k��ɒđ$�`
�
�5Z����'�0���a�3W��逵�� )�S�'r�qQ$��-��}�NI�}Wz� �'����b�G��� ��q�2D��'�Ĩs�m�T:����	.dY���'�,�8���<R�>P2s��q t���)�t��/2DˆFJ(���{��N�y�OSτYc��W�*U�i�g��y�hG�8����Y#mxi� ܸ�yr�E�x��f)�*`��V�y��b�� hSP���A�D���yr�>�j�(�@^�;�L0���ܵ�y�Kŝ.��C�+قK�л�I����?���(0��a��C�n^4�Їȓb���ĕ2W�����n8��/�Ġ a����fTU�H�ȓ�� @ޖTr�H��nٜeLh����L@,$��0�ˋ����ȓ'��D�!ɚJT�i�������m����*[&_��$�,g��ȓ8D�b2��H�7��U-�%���	.�<�3	П	cT9�b,"�B��=�I�uA0|.�J�L��L����0?ѧ�ߧPN��rj��QX)i�G�<�n���PaC2���J�0�ĊGn�<��C�X��P�&.4���;�Hl�<��e�p���3���/�3�"O��
�
,!����5*�r�k�"O�	����<0>�0��D茀"O�)YR �1Dd�a�kC�U�h��'n�	
ׇ�L�� �d�q��'q�Xb�BX2,d����KӜC\�H�' LIe+ǭ3���Q�[n��x�'��]
��?%h�C��Xv~]��'L�jv��	._� RC��:h��x�'�xu��g��x�j�Xb*�5=���'�䕫EƧwy�%���[����'�<a���^���a�Y.���'ch�kC�X+D�|�#h��S�'m�!{R
S� ��S��ZC֨�
�'��m��A�i� �#aS%P��a���hO?��  a�`Şu���0�!(~�� "O�sa�2d�d�sǏlԩI�"O��#ULZ8<��jd�K�6�:iZS"O�|�e�R�A�bS�O =�"��1"O6�*`O�z*�y���5-�\"O�=�Q��+Q�ej�ɞzqA�"O|��EêI�� A��ik��0�"O�ŸP-UD֔Y�wO8X\��'�|��'l@�[�G��٠gIƤ�
��'^�;Q�Ŵf>��@7&ӥCqp

�'����½{;��c�;`n�	�'��xK2��; 1�Ia3Q�@�2`�'g��ڲ̓�;i ؓs'E��J���'E\a���_R����m���h��yRϋ+L��a�סޤ����/����O~�d6LO�����S�Sq��.a� ��"O>5�@�މ_E�T@G������"O�����b����&E֙2�x9I"Ov@i�lP%�>�9oM�c/�)T"O8zc�ČA������_�H��"O�E0��<{���WbG���J��'\�'mTI(G��f<R�+�PRX�*�'��t���$5�H;i���x
�%?D�8���F�K�2+@�O�|�N�Y�1D��j���2��0X��ȃ|h�Y��`.D�<��ɏn�.i�#GF����P�H9D�\��A 2|t��Ą .����@�7D�xك'�h��}��@��m� ����*�O�I�/�Iz�	 ,0?�(��N�=]���O��d+�O`̚����^9�'
�"Ơ2�"O���G�J�1+��'�Cy�"O"}jtE��j퉑�*G�V	&"OV1x��W� �#� *��4X�"O��Ҷ	z�^2�� 6S�`���"OX|�q�G��I�ʚ��1��"O���ũ֙C��,�&N��ɀTQ�W���Ia���EF��3�J�O'Rmp��+D�A�]�X�}��XKd��i*D��
���k�D{0'̴t~8A:@�)D�@�S�� ]���Sd�e[ܼQ	(D��p'ō�:��Ahs��/V��9D��[�hV:ttx���աZ��ჭ8D�l$��Y�0Y6�V:i���p�$D�� �����7�S}H�q$D�x@I?Ct�0"&!ǆza��1>D�`�6�O$!H2�F�51:J��`G<D�DqC��+Z#u�R�\��A���&D�0z�!n�6ې1��c�F7�q
�'��<��HL�(㠒�D��	�'6��B� +=dr��� �O\`��'W�h�`ց44��$&�3�`��	�'�p�Yq�9̲�����!���X�'����3� �,vЩ�#��<B����
�'���9"-��_���g�?�I
�'?n�Q��8/��Q0�֘=�N� �'� b�n
���[���0��
�'ގɂ��7n�ҤHqk�61)ְ
�'>�( R�'g�L �G+A뤑��'��8�6h[|��J�#S	wR�)�'M\a ��^gw�h���P�y��Xk�'��D)�
k$��i�*�x��i��'�$�p#ѐa�
�Jf�����=��'T,���U$2Y��i��T�v�P�'�F�h�O���@�+�I{���� �P�A���"`����`"O�ɤ�E�)s�����9}@���"O�$�Љ�T؁�S��4U�t�"O��R��<�1F��&_$�P!"O@���NS�;%��B�ןN�H��"O��^�N2n�� �'U��|{�"O�Y�Ӧ!K�f=2�)L�'�,��w�|��)�ӿ&�\�3�ΪQ����3R)�C�I�X�>zT����ڀ��l�%"$nC�I�F���	��ͯg��tH��L��B�	�n$f�@��	�
P�qQ� xC�I1�:```�%`�*��7����B� ���R�U-d��BmD"$�C�I�_O���Ń�&^�v�E��;Cy���hOQ> �ӊU�H�D�	*�{�$D���7
�<7HL=�v&�-V��h�3�%D����
�Sܢ�A� Ў
'� D��Z�E��t�'%[�����)D����̲9Z�b���<V���l'D�L �)���ꝑ�!/`\��0D���!��/����!��BD�1�)3D� Raֳy��u�R��Td~�{��0D�`+�V)�l�p$���D�´�#D��Ȅ(�?f琸�P�_�B�ó.?D��@��E�W:y��N5CW
$��=D�@�M��%���[֯�7(������1D�X�`[V���w���}ȵK�*D�$ �eZ<A 9ې�S�B~����)D�Ъi�7�(��'G�,�P�'D�p��`X��a&��[EfͲ�A$D�S�@�'5���-ƗZ���q(8D�ث� -�҃äZV��7m D��j�JH�+���Ȁ����� �#D�@A�/��*��TҀ��-#�r���#D�Xq�I�%�b�'aY g
*���!D�����P�OphB�=5�J��QF D� �����lڦ���DƴQN��*�,*D�Pȣ��(wx"���(
F���J��)D��0Q�E��hYSQcH����	U�'D��ǄD|����3�r=�gK&D� A .R(A���� lL
��U�")/D�� w�_�SxL�"G�h���d�9D��3Ŝ�\k��U�e�o:D��2]�ThT�!���:X��*t'7D��1�ޥYr��t��S�R!k�+D�lh/*r��c�U3m��t�;D�02V� �v���#����&ak��;D�H(�Ĝ�"��83/����rA:D�����I��*؊�Β%<��j#D�`���4L�&`p�D�Ǧ�iӧ5D�8�գ�-�j6I��"���@�3D�����:4�h�q���;��ق�h0D��H#�R:L>ܩp��}\��D.D�{@��8pJI�#f��i�l � "7D����մO����&W�R*@B!D�����PP� �\�6�z��?D�$b"g#
;�:�g�Z��7<D���CH�3C�@��꛽e�
��;D�(���Ё$7a0'��]4��RC�8D��sT�E_"#��9���#	l�<)d���!T�DP���%[��RpAd�<��VP����ơm�0����`�<Y�GW�<�|�:�C�6����e	[�<�%��(=pB�AGK�D�V����Y�<� ��h�ƶ~^Y�f_,�
}*�"O�4��٣t:���U�z�\u��"O@���k�|��oɞA�q"O�YYa�I!<Z`��'霸��i	v"O���N�>(��qt�0�����"O�ĲB,Xe���K�I���6�
&"O����ѿn?nT��ȁ-7��:d"OĄa��H T�Bǚ�x+`�S"O��h���F��H��/��L���b"O�ڰ��f�F��גC���a"O�����Q#O�V)XS�Ց3�\�C"OY� )̱K�)�Skڅ #�$ �"O�I)c�V�g�jp�D�TΉ��"O��@�.\3y��w�t��1�"O�=)��̯eu��C�N�;�zQ�"O�xuC��~_\-zs���|�*"O�h#)Lq���P≇>S��4� "O��XQ�)+ٴ\H�i�:M��|0d"OT�p�ڱ_��(@���F�
y&"ON�T�� �x���UjԼA;v"O�<+M��C��y	g�� )�r"Or�p`K>e~TQ��D��X`��a"Ob(
�E��f����Ӂ R��	U"OFud�!#p���P3�(��U"O�A�GPpm�<㐭?Y�H��"O�-���?;�,l��L�+ns�"O�@��+�&Q��8��J�X��U�"O@L9�� ����*��-�m�c"O4�St��CfQ1�^�(�@;"OnAC K�{���S�"[���
�"O\\Kǌ	�p��V"�g��4k"OM��h�2D��+��l{���v"O �K%dȂ>�t�&g��{`�,0f"OBP	�_;#�<$��bVZQH�"O���@j�./��X�Be[��ڦ�Hm�<��/S�/�`Ȼ1hP�$�L4���Vh�<!@�W�?������P� �ɀ@��e�<1���E�������"9r�*\e�<����l=,�F	_/%���E-d�<q+R��n}�s��;O�<Pbm�G�<�������1&��}t��b�TK�<�īYVP�Ъz��[�	RK�<�P/�aA�`ڥGU$~�mC!b�<���x���f�K����r0�ME�<��)�T��#�)s�`z���C�<���Ȑ$%����	��}�y� B��<��C�O�V�ٲ�Q�LA&��2(�z�<�,
Nh�9��H
@\yCd��M�<�Պ��8�BH��j`�AP��J�<�&� VYJ�����7a��^�<��/�*M��S3g��sdT�R5"R]�<�� ǉs^F���0yBuB�Ϙq�<�'�G�7�Y7@Q�:di�eG�o�<�g�$6^���S���*l2�P�a�h�<y�jX�!)5��T&d:�0�(�d�<9W	��?=��	dmZ:��#Ą�`�<��j.
Q|�r�j�&�tAh\\�<���R�G*p��CA�%bxm��"Tn�<� �G#o��5c� ���59���s�<�Ш
.S�� &�9.���Fn�<p��+-8�@�Q	�ƨ�^�<�F��zO��:��ܤ9�%
Ċ�T�<�`�]1?b���v�O%u;&m�EUS�<Q5b�\^�Z�Bׇ0�~�C! RS�<� ���%N�	Mv%�T�	9��<�%"O����K�g[ m���C��!�"OB�2�.�#uBԥ*q�Q�f��"O���F��7]_l�S��q�"O� IT'��H��c��*^����a"O��8W�V�w��� e�Z�a:����"O�s4��$��b�
�Z&���"Oz�r�dGh�~�S��R�	�q��"O����`��=�iSp�з%����"O��#��(MlxQlӄ7�&4"�"O޵0eFдRDH�+��r_�(k"O�@9�'Θe�>1��")vPu�'�J�x�����O�'���Z�'l���d&�3d�j)�N&���"�'mT13��-��UH��#�HX	�'�Թ@ǥ}r�q�e���^Mb
�'|>�2d+��Q���A��=���S	�'ʂ,�a ՃW�85yGK�0��ձ	�'�����g�K,��A�/��"�y �'� p�2�B�uU��ꕋ)6nI��'F��5F�� C Ihv�K���'wbXy���Gn�!��ˆs��=�	�'~�@�׃�9t�Z��� �$�}��'� ��-R.(��A�;涨��'�$�p�Ñ'2$8(��.�=Fq�Us�'�ҠPflٳ\��av� /�Ru��'�<EIUNX�v��h5�����B�'��W'jR����膐s<�`�'�(�Os*)�%�O.or!Q�'gfR�FYad�b���d ���'8�F��z�.��V|����'5����n� |y^���.[�@��,��'_�ի���4J���$,x�2
�'��  �,�HH�2�X!#Xՙ
�'`�IJ��^X��s�L[3M\ �
�'\���jY�i��8B��?�R��'k�9�7D�bƌJB"ĵ1��x[�'�H��]�u�N�2�W�y��j�'7(��s����Z�`��"m�����'�aZ���8#x���cGf
�'���ᖡ�9p�x��lڰ�b�ȓBG�\A���5h�Dɣ�b3q�ȑ���8�A���t��x�"�-Nfz}�ȓjN�%���+p�L�5��5z��ATȔ{r��	uӮH�#([�6RD��ȓM|�e�ġt:�8
&�Y򈥄�K�:0��ϸY^���Vv@Q��g6L����8�bl1"M� L����ȓpU$,���H6����h<!��ȓϘ	R��?��җh��!�P@��*+D	�Ծ`g��Z�g�3ck�)�ȓf�`:fe����O%k{x��5���!��.��M	�:A�H���F!��ǭH̔���)	�6GBԇ�E��4���3B��P�ѥ2�$���|���:��  Q�0��J 2�H���^�ܱ�I
+x��i1�E�gz$o�a(<�`�1x53�+���PӅ�S؞P�=�'E����K�z�0�ӣ��D�<Itm�{����ř*S��0rN�i�<iB�`:x0�E��Lk� �t��d�<	��0l�d�9chH�ޤ2��K]�<��ƥjZ"q��Ɯ�J٦8�f(X���"�O����>L;��I�N1�2"O� 
x��oܤNPL�r� p�����w�O�z8jo�+Nf���"���C=�1�'����Q6y�E!"J�+H�d��.O,�=�O��'l>�+�G�'���� �r��H@�'��Hh�B�+Y�H���b,��A�'��l��g�RQ��]?ֈ9�'iV��e��,4�J!c;[<qC�'a�ս"��ؒE��uؔ��ĢJ��p>�M<	"j
	�B�"U0;|�!
��Vj�<��ɁZe��$G�B�@�3��i�<�w뒠^�(�3���&���#��f?�G����'<T�	�]��(
�����
�~��nQ�9���8U�%��Abڡ�>�%�)�I�hdxp���7�i����!���8\<�0V
[S ��2��	:>B!��13X6M	�!�l�Z���텻}!�$*<���� KCOl��,Ω?�a|�|�DX"\�l�s�Ço�=���W �M;�'��Ѓ�S��ՃcF�k�@���'����h����鱢��]DF(�'ǚ0���>@��q�A��B����'�j��6Gt�Ш���8U ���'�2hy3h=�r���Z�b�(�Q�'ex�!B���D-dяT4Vz�Z�OP��dՁ`L�5E� �}d�#�(�8��v
O���3hY�`}$��!��y�-���'���\q��v�\�f����!�<D������?���y�Bäa]��6D��Y�E�j A��y�TР��5D�\��.��Z�JN��8��fL?D�� +P�8Ƞ�Si�=L D�J �?�O&|�Q��9]��s%
v�Ɂ�'S ��C�X��؀"�(�s��2n~�C�	.G�*��G�#�
�� ���0���$Ie�'� �B{U���3��O�&���'��6+�	�(����WiJ�rpfJ,B�PB��G{���"ZB����&���8`s[*.���?��Q�!PeȈ����
3HƷ#��ȇ�_�!�4�:i��e�ef��[6*A�ȓ��4M��-!#�Z�Bh��?�����8>܉o�8={t ��)� B�f^���e��#�J��R�y�B�{'��Q�0V���'�D�">	�{"�~Br�ByT(@��iݢ�kF�U[�<A��H�T�����ב<���(���S�<O�`T:���B�)0�X�pS�X�<�I	�,i�ScJ+�ph����<q���hO>u�q@	Ef鈓���He���*D�����J 3֘$�`Q�I�2K*��G��H��m�4��q(�ܴ~��5!�A)}�)��$:�P�+I�������цB�I
/�Ĉ�Db�'6Qf%H��X�i�B��!a���%�Y��#��}���k�� R�Z��Y2� �6Mj)r�5D��	Gȃ#� �2� (/)@t�-D�p��w*�v`jxB$��Bl�:�=E�ܴ!x���7酣��p:�q;$�O��=�|:�4~ݜu��	z0dlj��@����'��~��O�;�8}[�j�I�=1��y��d�>���S�g�ي�e5*`�qcE9Q �~�V��q���8S�
p�v����v�3��1D��d�ɻ�x(e J�}#bH#�/��ȟ��� %.�@��UM�*s�U
R"O����Z����@��5�� �$7�S��ހ ���rlB4S�����ۈ����"O$)DI ��J$��:xPM��	ux�|9�(H�&��l��t32 1D�hQ�H��c��	  fؤU�,	@��/����%2����r&�ݪr�ld�@"O�)�mV`H�e��V�t�#�?O��=E�4`��W�=��ۻQ�n��Ԋǎ�O��=�O"1���(t6<��ģ���\���'6ꠣd�E�,�B���;w~��'�\} ��E�'�0�P�H4RH�	�'W�����§C���0 H��~`/ؼ�E{���iE��Ǭ�H�©Ȳ͋�u�:8��'� ��fi�!�r1Y�DpJ�R�Ovi���=D�Dp{3�"<�tNځ����9�DԱN���	�i�t�"�T�(R�!��A8'f�#&	u�6|:�H�h�!�D��H�0������!8Od!�d�S�z=�Qh�6c���!Y�8�!�N��J�P�(�TK�=���C�i�!�$ٮh$���"�O�E:x�)�@t!�䐍�P��k�:u,�AgI�}c!�dR�0��{�f�b����%)��s���4��d�'��[�.��\(pǈ�981���(�S���q��u�q�M�VК����y��,�rS��¤(�o֯�M��}�=O?7-%� ajb�1�zR���!��!N0p����a��}Ӷh�%�!�dS#~����/�PO�h�' �e�!�d5��XT�;o?����T*e�!�$[�j�\b�+��Y!Z��lM#�!�@Vr�͆z�03C��.	Q!��P�E|ur���������՛��)���x�B�S����N��<n�!�M,D�0�bG@*4ͼP$�߾]#Rm��*�>���3��j�$�9o��˴���Gj���3��rT�V�0H�g�3'�]��?K�y�AA�&�R4���'fb<��Z%��e��LT�=�4A
�1�h��;*V�JS�4g�j��S�" ��'�����pE;�@�_At�u銠!"�C�	%j�r�H.Ș(6P�j�g�'HO�C�I�r�$������9r���+�$Ϣ�>��8�h&���K��x�@�_��O.��d�G�P��)۱!�a�&������N�Q�������C�<S��P(��;W��d��EྌI���>�)��Q�8$� '��F{�����K�J�Т��z,�7 ��y�n�5lJ嫶f�z���M��=�S�O��u��l��)��UlY`��'p�$�1`11�ɓ�ia����y2�'o$H�f�3h�����05�|���'�z��C��J�RE0��>�2mY�'�t�B��[B
AiG��=�yb�)�S�2���Q��u*w�b1�B�	(s���
�������ɏ(��B�	3a�N�HV�����A ��1N�^B�7g_R���Q+=fl	rC6�:B�	�"��Rfm�R�cM�$92�C�I�����F�f�0� �����B��!w����,V8�R�XF��6
lB䉌?VVa�w&N�}��A8���zjB��6WT(`��2K�jbll B��j�b�`�����H�0.��k��C��*���$˓RP
���	#i;�`���� nQY�!�+��)`��A!}Ð�H�"O6Ps�$�FO��A7a�[��ty�"OxB���V���a���̔��"O�ӵdժr`0�9�$<@"O�C�F�:Wp�)v�]�M�"O�1"ȏ�f7hh #H#)��	�"O��˱m:d��1Ѷdԛ	)�"O��x����V���C�P>]_ �@r"O�h��#ղ%kzM ���i��"O�I��(��_ʪmk�� �\�y�"O����d��B3|�
�'R%	bDa�"OJ�)DA�c7"js�$G:��"OTY��?�x�W˦&76��S"O6�bb�UN�Y��I�x��"O"T!d!�u_�قq���d7p�X&"O���v��@�$<���@#|��"O��e/�;A �y��G�?y���E"O}� ђJ�]R1&�G���&"O:����X}8��qd[7v���"O>T)�k�R©����+*��L
'"O�aJ����A�	0"�^�4�k�"O4�I�c�n� ��_�_PZ$�f"Oz�sR�U3M8XIc��d:,���"O6�q���c��SEf(��"Ob|�FI�4L����$���j�"O���aJ)<������<p� ���"O�XS���0�zP���p$@�"O`]ۥj�;�r�L��uŘ���"O�)ae��b],�V���{����"O,q�#)��w�ni@ֈ��5���s7"O2AX��^�^���A^��1��"O�jA�ՈB5ʵq�	LbDf���"O��+ �$a�nY{�W#��:�"O�<1â�HF�b�m҅gd���"O|4aV��1XMP4�VW��t)R"OT�x6�>O���0B)�:�D���"O2�"�oL�B�Q<C�
)�ܙ'q��D�3_�T���"H��P&�W4�yb�0#�~d��N��y��ygR��yB�SN��G�6f����R��y�oU�%�>ɦ	[7H8��IW��yR%�q�"E�Tb�9O��%Cbb��y��,yx^�&J�ļ����y2�_�]OB��) �K���UB���yoƫ	r�� 6iM�L��z�@��y���oP�	觉_��� ��%�=�y����Aǲd:�`ۖ��a�D��y��?��{B� ,�� ��yR��2N����� }�*a0�	��y2H�/���!ADT�\����" $�y"�Z�`L �)T�\�_t�������y�f+9�Вs�E�����)�yҀ�<�⁹����,������y�Ŋ�Z��XGɛ�-�ZycB���y"��N��Eq��%�$�i"����yo�"������R�`R"���P�y�-���ЭH<~]p��̏�y�F�9fÖ���iȖ�Lp��$�yB���7���l2�~�`M*�y��B�L�<a1���ph�`(��y���Up�a��Վ��p���J#�y��e˺ՙ��>=��ږ�ߦ�y��f� �
!�7 ��IC���yb��T8�p�%S*�>�r�D�6�y
� �I���<���C���%"�"OtȲ�P�f`̸���q���`�"O>y(G�'��1���*}̐{ "O�eQcm�)���Y�W��W"O��[��Q�u����&Y�X�i`"Oڰ�S�1K���@eآh�`�"O�����9B<�̃�M�d�rp�"O�����64q�����Q��@��"O��[5]�D0:���(7aI��"Ol�l@�k��B ��.eJȩ�"O�0�a�S����o�0@�dQ "O�m@��)���B��K.&�[�"O�S��\*�yP�a.8i��"O��S&�TV����B��]5��)�"OΡ�å��wE����7P^2� �"O�h;@�%^�܉��]�bG����"Oh�Ç+�Y�R����c/d�c "O`�;���*�� D�-1uZ�"O|IK��pK������$9�d�"OH�*C��=p~�I�Z�#�d�&"O2q	��+�8k�J0G�(j"O�La"T'�|T@���� P��"O�A��Ɍj����kW'�Z�@@"O>����;���i��^H�"O&�"��y@JЫM�?U�(8�v"O����D#�m�C�ˊ"u�A{@"O�a����;!W�~Y8���"O����A�n~�8�!�I�G� R"O��ʓM�f��HHu�bL�b"O������n�6 �_(C� �� "Oƅ��*K�r�0M�U�n����"OT����_Y`PG�'���:�"O�8Js�X#�ι)eۑ��1�"O@�酀%V|�f�59�8 [F"OV�3���D4	���$�ı@��IeZR�#��S�Q��(с��0y���G��j�B�I q�]��U�%?ޝIB=]���Qg�4	MT�&�"~���H�4B�.2I�2Ǖ�R�ȓ6`\���.S�|�3�׀T�J���%d��
E΁�<ba{2#M�U�(e�H��=�f(i�[�ʰ=��gP!�\�4��ڦ�p�E�I������J�W/��7�0D���b-]�s�P٧�"������+�I�J@�Q en�X�G��cW��ظӊQ8W���pq���y2&!
҅b�MM�M� Q�U☪k6�xR�ܪe��ʓb�V�|�'^��JU�@�	����-��_�^T�����V�"}�a��qsPѺ�	�N`��@bBdBJ���m�t����'�~�P�� n�����܈P���I���s��ԟ��2C�V�<�b�����4	��a*�*u��O¨���'�FThя��8�PQJ]�*M�La�O0m��ջR����q1C�<i��~�ҧE�]]���k�
�TI���Y��4���=)���ɾU��H��3r�L����Y#?Q��k%(�t~��r���J�5�����>Z�jQh�8��XR��Q>�B%�~�\�'
݅F谉R�T �h�W-;r����$(6.0���*�E�~ě��~+4�D�;)�lUJ�{����Aφ�x�`�	3|�A���[^\=�D��,B0��aX	N�"~�	�>>$���j��wخ`2�� ��I��U�tƑ D��=��l�SфE#?��M��0ev�8z��'L\<��n�<�T��ɘ�^Yi�G��z�(��
9H|���dD�<�9��x`Z�r$ҋjEK4醆:6������'�y� �1��L0�O1���2QN���1���:1Λ�|
3#�2or)/��  A�!҃w�}1��ׅ,�t���J�)�mƭ%��ɵ��t٢bś��n�b�Y�_�V���'W�y:�-�m�g~��U�� ���������������O:tx�Hʓ^���I~Z��D�-]��Q"�KO6�9A.I6��ŀPL�s�f��� ��{�b�!���V.�ҩ�P�O
9� �5�~��O���G����q�:4�N���r�ޚ*�	vaOR��98�O��Y$�T�_EB��䏽K~�;a�>!�퉝��h���:�V�r��(Cۚ��W�Hr"���?~*q9�!Z"�|@����6'���D�&i����`�5A�� �G,N�:�������OLdcT�̠y��,����-m��q�t��4��'���y?����,L
v s���0A:�>��]L�ڌXW� ��� nH��+70�]`���2Ck�+` ���
Ds���9��1O`�� l�rѐј"ΜA�8b�Oʀ��Gt���H��)'�Y*���q! p�t��Pl±��|��B�p߄ �e�j�.S	�'5�,�q�=t|��3��j��1M�|S_����a��U;��ъɼvx��v.�l��9�OFj	���ģtLr=S��E7(�p
�L��:M+6�FT�H޲�B4I�,Ѭjޑ2��Ek������$�ٚ������'��	!ꖥ��B6��#.I=G&�?Q�bO�c6
c��KƤŬ	hNi+���D�8Y� �DOPԢ �4g�j	��
w
$���I9f�P�����/A�Iٱ&���>���H/C�U�!f�z�.�SֈՈ>1$�p�R(ho�#A#0�N���'��p�bIB�� �U���d�PM���֝b�4�C0E�70̬p�吮����V��R�[�$A�\k�nV$ؤ�K�<�Ԁ��`�\1j��6G�]�d�U�O	���d��m{��K5T��� �?b�T9b.���/dφ���-������H\8k��/�����ܸ��ɄdJT�(��jXIG��8��DP��P�p$9�Uu֘��$D$ˎ�f�
�MN�iU
_x�'OF�)�J�~JL�'4<!A'U(~q�1)��a��̨��� i������rFF��F8�p��	=�� ;vX&5t pD#�6}�Mm�d��ho?��'���� 9�t�&�
�=Dir�e�hu�̑PO� S!�Urf 7.܌!9����iC3BMI��F��@IA�&�9�\:�KD�m"b �
���N����#o%v(`2J_/����B��(ѧS6.4
9��M�	b�C�	��H��s�S�Y`���+$ܒO��BX.,аى�i�2~Xq�6�MjtX��̞b[!�d^-���+Gm!��1J�d��bp+�a�D�V� �?�'��y'IB0O�E��$$dπE��'P"�a��k��aÍ��+��8e$�&����'{�x3�FK�~~��#F��$��	�.�C!'?9#��=j����@ȕG�u��O�<I��$}#��Zny�X���K�<���ޔS��HА�6)�ժ�*�y�<y�M�;T��xS��`Sȱ��jo�<ҋ4d��%���[ 9l�sB�Q�<y���H�&�3@�!jC�H�<yV��a��);��&tTZpYN�'n��c��R�g��mc��($tP�WdZ=m�ȓ@�|�3��[�s@�a��=" D8�'���+�	
]�a�)�g~@N�g'�сdBR��~b�����x��]L,-ۓz��ݣ���#W�Y�$a@8�W��i�"�!b�'՜�pQ�a��)S��Z�\/��R
ϓ`�����O��bҍNB����,dw���T��:��\ra��+�x���#�X�w�~�� 3�_��y��xC+�O�(��D"|P����bE1G�0�Xwd����3HM��y��ya�ʀs��y��ا9ԠM����O�g�^�}��i�3M��Op�	���g�d5� 
_4F�X�B=4�(��I�7i6��*0Cºh�z|��k�^�j`�F�'1.��V,�n��Ą�����.�vX�fm�:J�x����u8��%a:�p���L�:0Z��+���Xb�"��Od�D��hq�MsU� �|D6"0�	6O1Le�f��5Vt1�8 ����!M,�9H,;����"OX��g؆=���f�@�:�BذfP��Qt�U�1 ��%�"}Z���;��U{1��j�60S��Tf�<���2X�d�[D��P\p(�t��y�I�Q^t �d�'�5[w/�H,�$k���L<��	�'qvU��ŝ�"Q�,��N�5��H
�'�E��EWz�kd���	4q2	�'n����ޚ9l$�BFM�+m*��'�x�� ͂4O����"�95"Ts��� P���su�8ؠ	ڈkN=  "O@tv��3/]��SF()����b"O��1�^���1iP�0�C�"O �(d��`��tbC�I�/�ĕ@E"O�8�GƔf݆�R�˞Vے�y"O6 �"�"jhX����,�>$�d"O��5㏶�L��C����x�x�"OB�(� �a�[D->v;(��S"OLH1��>R�h��L\1����"O$�q�)� ��XGJ[&Aʄ
�"OT���O�1>��xƩ�x�ؗ"O�HS�@@�pRP8!� �	o�xʷ"O�$��(� �:�#ń5+N�!q%"O\��gcV=*O�����_+Q"�M�c"O4 $�N�(�U�&D:b+�찆"O"��^�9����7}-05"�31�!�D�(0��Qʀ"�:| �($��x�!�D�$�h�C���J������?FV!�$�1SE�X��Le���#A�F�]�!�d����DeK�s�4���T8)K!��{:<Ź��О��Q�D
�yS!��C��Z@�A��� ej�0�!�Lc`8ap�.�
U&�db@��4 �!�D�2a�P���HR*S��}��(ʣC0!�D��A��ԡ��}�v�
S�T�#"!��R	�|��	_:�p2��U2g!�D�+BL��jթҬ,a��	��P�!��IW�-2����gg.�+�/��_!�d/JH�"��?MC���TN5-:!�D4;�8�e�@6�)�n"'H!��[��`-�l�ڑ� F�r�!�<t�l�Š�"=f�y��I�!�+�2��G��/g*�SW#��=�!�D�p�^@���[,
X�kS�BU!���'f:y��	��B�(��%:6!���L�8\��SB�!�5�	y*!��
�S!��JDA��9�@�s�E̟%!�d�1���!8�x09���t'!�Ă�wN.�z��� �����PyүI!{����ņAHbX2S м�y��$[:a�f�RR#b���yR��lJ�R��P�(Yp����yb�F�&
t�KP�K�Ls���,L��y�E�cuܐ��<wEZ���b�;�yRe	_� y�'�&�$�8ǈ���y2ȋ�{vh����\�
h1 Ƭ��y�L�;��Tre��>k�v����	�yr��cZT=+�Mոbb�4�1��<�yb	�/�tB���;41L\j"�)�y��&�v%��!�y����L��yB��&C_2H�&��CU����y"GE�Ks����Êg�<m ��ܤ�yR��:Z6	�k$�B�B�)��y�O�z�@�kΔ{<�h�#h���y��|@��!B	j��|�B��4�yr(�.kx�`M��D��!�<�y���r�L<�����$�a�4Hδ�yҮ�(�T=��I���Q��kׄ�y�aQ�tx��V0�T�A���y��Z�$d�/ {
�4�ʐ��y"�\���إdн#@LCᥟ4�y�,ݛ:/�4|=Ь�dK�j ���l�j��L�F<A��_�)�!�ȓ/�Z�@���1F�P��	J����S�? p�"�]��&�N�23�<	3"O�2%��:.!��z�gU�~%�Y�"O�L�DCO!>|�ۡH�m��M(�"O4�Q/̎n�Ԁ�D�ːmLrp�"O�8��˒?I6�A��8؈��"O<�� ��v��ŚS��N'�82p"O��)@#S�2�Z�KL���Jv"OԌ�s�S�u�2��`6o�t��7"O�B'ʑ=�X���+P���D"O�`�'%��W�8�i`�
��|*�"O�!��ͮZ������Q�p|��"O\�!��PBȌ����G�lXZ�"OF���P9b]�ĢT,�c���"O0��V(	�b6�a���:���`Q"O�ق�P:[GnuB"�0b�h0�"O��᳤�So6�3G#M8Z��࣒"OR�K��G:S�B�����sǔQC�"O
�ۅG�Y���Q�ѱ/�$7"O��㗭ʹ4!���	"u�^5x�"O�q�rEγ:�b��FG�=qe��a"Ol���� �>�X:Æ]�|tT�j�"O,t�u�r����d��.�$P1�"ORdk�gI�8W4�B�fT�(p���"OvD8a L�4�,�%�Q�옫5"O����$�~�a�5g�h�:�"O��`�͂gߐ�W�.~��$"OH���,����5�Ci�� ��"O� ��<�����R<	�u�"O� /�8n�`jUf�)��ms�"OXD�n�;��m����=ބ1�"Oެ;t�Q�PP��w��5�@�і"O^@`�1N�p�rP�H.�a�"O2-�Y�xJ��bO�7��R�"O"�9���a��En]�!L��j�"O�� SeŒJ�v�i�ā(+~e�"O�$g�S�u�>q9�i/�`@A�"O2���LXH|��!ɕ;��c�"O����F�8 �����b�b�2"OP�ă@;rʤ����9Z�j��� M�T����bj��k�IB�qX�$��ꂮúB�I�n
���ͣS���Ŋ^,ZM���&  �+;�8&�"~�w�r0����2��i�E#y�N�ȓAr �j6��Q?r�ys�@�U�>����g&V, ��W�6�a{�#�%P�����/�)H��P$�����=	���x��B�Φu)��9��!�+^��h �'Ĺ�yR	��DĠ��hUډ�G�L�'�@� 惷L��9� ��	ɴ	GŲ>Y��+qI��z�XC�I"-�ׅqIP��+)���qr=|W�5/O�����Y�4�1��]��(���8:��sD+=D�d
ӈK*&�䂖d��=�vD]�1������M-nCİ	ۓ����iH�
�⹢h�F�m��I2z��1���x�2Ho��t#��J��;s^H�B�l\�C�I&X��т�E�j<�A�1���qO�� �B�\�<�"&�6ҧ��C��"��䠞�7�p��pU�h���)|	"�i�*<~�2A�E	�����O�u��Y�Т���8�Hi!.˂uY�� �d"D� ����ci��#LJu�h���"�D�	�&J�2����d��0�ȤKB��QN�)�b�Ra{Rcʈ0 T|`��O��Yш9yX�[t�_$l� ��"O`,s�"ۤZi@1���K�n�h���^-���P����8.��Y"��D� ��CN�Z!�d˅��M�p��t��P� �F&K!��w��lA!��?R���F^!�$S�L�R�A�ۦV��U�D'�0]J�'��]�dg�pX�� ��('EϪs �i�a/��FW����'�ܣzJJ�pQ��%$�aKF�Dv|���
O�z��E%}�l�#�'��+�$!�ɪfRH���=#1��1c�)Q�p�j���ƃ0��9D"O$���ªEa�Pu�3<��t�OR=:S��6����L��}z�̮��,��M=�QA�M�X�<!�ƥF�A�C�>ԉ��^Y��'jMȳg���0<9�	G�[���Sׁ4S�T�F)|��Xbs���ʸ8` �w\#eM)B�1���M
!��ͮk��0�'�!��*����6�Q����uv� ��� F��jJ�ۤP��l��"q!��J�sZ`�Hq��%���Jӊ�)���E�P.D�NW���)�'nI$�� �,���z@A �D��!��"af��g�N��:�Mг=��O:$X[!d}�u�	ÓY�܀r��
�jK� "���Lyt����.���)Uʉ�T��4Ƀ�ǎ2�Z U��������@�l=��A�>1pʁcޅD�DAL ��~J�,j��QA�
�uж+6�D�<a�hRvx�łY*0��(��et�<1��L�x��䧁�%ေ#b��s�<��	�bwJ����)D{�t˵-��i�ą�=Ѷ�7�gy��Q T���Q���AǶ`� �[��y��[�;�u���Gw@�Q�gS��Փ�Yh�}�ȋ�}�J��UB_�F
�y��W��<�u�� E�Q�Ʒ>q�&��m�z���/FG�4�y�C�<1��١�8��mY�M)�)a���ey5)� 8�?�`G눤0���ɉ�&x�m.D�J��&0����sk��1KD�(⪋�b��uK���!�TT�g�d�yJhb�c�l�T)�Һ>,���G�}��'\
!왠�N�"Q�j�Ah�*�1�(�O�Xhd�����ӯO1��Hr�'���/N2��@�'캨2�	ʥ[U�P�S�F�Gd�$��'��w��W�(K�I�=�F��K>YS@I�8�R���1�'|i��a�	-
����*�ْҬ/D�Tth�1'N����ǍLt`�ѧ��B��{J���Bc�l�g�dfG��� �\;M��UK��APZ!���<���cQ��P֜����mA�����Y=����R�	�hYXUGV�f����Q%/[�z$D��$�'�X�Q C�Q��R �JА0�	�'p���A�
�Dx����ftC	�'�,J�&=���i��V�����	�'d�8��ˍ.y8�D�UF�y?�Li�'�T��튓�  ȖF�4X��'�~�')G��T��2��tٖ��'9tj 'ܘpڋgH���O�
������OB�@a��&r����kˋ��s�'r�� �T#wu�$���݅3��I��O��S�A��,�O�>�S!"6�p��7��--� ���,D�L�T�ڭ)�5�Y.�`��Ԫ+}+�_DݲS�W�8�� �'6,�{$��|W���)�Oz�Bb,R�6q)w��_"P` K�� �ڱ���x�D��j��y��Ɋ�f-0���O0��&�M�a���(��To�*�Tt� �kh�U계���y���h���Սd��u��0�~b��Z�ps�h�n�퓂+��I��7 7 �
�放kV�B��.-j�
#�ˠ{p��1L����'���e(NY��ɦZpt,�V�3FU�,�U��#�����	&�~��F��ed��9��^
)�dl��ʄgX�H�'Wqb���O���0q+3~�|���d��t�6����X���O���)d��	*9:1�ʹt�jЁ�'i�tp�׀[��(�p�[�nq���O�R�呇I�ȒO�>A{�(�%���a"��G�nQQ�e?D�x�E�Îy����C��Z9"�E;�d���^1*
˓aN���חb�|!�#إx�Ҕ��S�? ��JI�G�ժ@�R;
Uq"O��s	��g���&�ݦ4�� ɦ"O��� ���{a݃,�h�
p"Oz؂D�܏Q�,dZF��usHPSf"OPY��ͱ�2Ǩy���"O.y�d�ۛs)�|��C�� 1sQ"O����ʝ(&Z�HcbO1
݌�5"O�Q1P�lR4�G���,բa	e"O���h�=��G ѕN��䢲"O��
�pi�!��!#��s7"O���fh��hƔyS��"+�F�6"O�T�1���2"T�c��8[&x�8�"O\]�RF%S� [�Q�B����"O��� ��B��pS���	_B��"OL �6��$-<�c��4�f��G"O��6�D,;'�ċa�¯C~B��V"O�!p"�]:;���K�YkH�[�"O������GPp��-�QQ,,5"O ���K��P-�g�Ϟd@V�h�"O IA+Z�1kp��� !��U"O��b���?��՚S囀m�TĐ�"OD�+�/��Pf(��b�E龵��"OR���I�M�B|pӁ�"��"O ��C$�):�x5oZ'h�H�"OH�+��/'�hb�>$le`�"O�1�ՉZP2�p�T-��%(t=3�"O�=ۤ @�� ��֫O̰�"O:��T$B /`D%z"bQ��:�"O��c��M.Խ�B���� �"O�Q3�m�5M4%ȠKS�y;�s�"O� r��>]/���I�)�`Ȳ"O�A�ŋF8���W��:��"O�" ��5N�H�@��=w�T�"O:�Ж&.E�X7�Q�D҂"b�3D��1�[�,�|I����.��iY�'\����^��z�E��0|" C�;�ݸd��&�u(��1Vx��'��0�eτ-C����	���𠸧k�*]M1%d�E�b��{�ĭ��e��SC��XD�O�$�	F�[�P}��	Y���ـ�4<�
qC�bC2%C�T�<E��%�.n#F�����" �D��Q�ɿ^�����>,
�md��#	�'y��� `釱�&�p��	��,�w�_��|��'~L�uF!�R�S�D
B�ӄ$ߪ50\kRQ*-�!B� ��<Q� �5&4���>�D��%�;	I��	�OƓ`ЊE nd�����0�f8��"�����~"gF�gN1�7�!qev@s�S=ordPQa�T�|R2GFG�gL���̺��_3ۤ|�Q�\��4������9�m���ȡÐ;O��~�L?I�u��*+�zњ���+w�~���ƄYv�����W-y��ר�h��i�n� 0��g�V�5�8<�$�&�@��y2ME�P��Չ�S>qG���A$7�|X����a�&�H�%��;@z��j�\�VO$[�\�	�'C����v�]�4Xl�za)|3l!�=ތ��&˭\..�c��Vr}��)ЯT���V�I�Ġ@޴]��䌼a���HiL
��I�5�)%�	�{HFI��`J�|�!`���H<RD��D�4o҇Y��~
ç!��Q[Q�W� �Q��2
P")Y5�~�� !��T� �"���r�],�8���\�;��J�']���IciR}y�83a��ދhqz����	X�Ĝ���Z�����G�?��D��o��^	�������`����bX!u
��G�T=[ V�x8�ƕR�}q�i�3q�>ŉ�'f�Pd0 �c���;ċ̾<ziv+�1��8��I<C��6�/�(�z�/�X�Q3"ES��]�5a^h����E�5"P�9E鸟�R�$��se�����iuC\�K��y�p���W�ޤ��'�Y���[��O�1��٫�X���D�A��Wvl%��'P���"����s����)��[6(Ԡ�Ϸ9�j0!w�"fb�B�IH����ע{6�]a2(Õ<�B䉆+�.-���Q>4����wa��H�C䉅�� ����m�zt�b��Y@�C�	�+@:�*60������6K��C䉈wͮ����g�2T��5y��B�)� \�a� �Bx�`��@�;�T�J5"OZ�Cq�IJ��a`Iy���J�"O
u;v��S�&�H�����-sS"O� G`��W�Z�Qt�i��b"O�93�_2˅ 2f�Xr�۵w!�Dյh0<hE�Іs9�����!��-��\�n��*U�� �� Y�!�$B��t���(�2��ܴ`g!��=b�0Ak�	'l l@���76�!�d�7��t+`,�)����6�ʿU�!�$GBx#�f�#4���v�_<�!��y��ǡw
�ȑ�&��h�!򤀚PR�UIQ��*$Z�z��M��!��0V}������#"���$ț�UY!�d�-a���f*Ȯo/P��U�SS!�$60m|�l�Y&ډ���m�!���FhA� �{�%�s���J#!�$�T��E�a$G�3hl�Iٮp�!�$��-%����6L�F+��N�!��ة-7�-�bX�\�d�SIƀ7�!�$�)F���(ٍ�
,(2g�;�!�d��;�pX�@͞�S=�jb�ٿ[-!�$ý=�ŋ!*B�E�4�;�!3�!�$�7p:t�Aw�V?q�i�uA��Bo!����h��㙰!�H�s�J/e�!��<<�#���pn��"@�,$!�P$Jx�H���7DP8E�c�S)c�!�$��F�P슉'5t q�i��~�!��N�>��
�2����h�]N!�D_�+3��ÄŚ�P�,��5G%,�!�d֒u�^�@OϾ'�l�BR� �!�2��I9c)N�BƲ�'��!�K�<@Y`�ձ���!�!򤈑�8$�B�2�j�b����R�!�D��?�BA�`��)U+�c!�W�dvL����M�⤴z�CM�H2!��"}!B�2��³�*� 4�]�f%!�D�",>(xT�ª#.���)!��_��z��N�*NȀ'aM7!����s"OF�	�ɐ�ܟz�!��<�$�k� ���u���ę$8!��T�4k&]�g� (�t��#�/W!���r�h�̷f{����ǖ�!�A�q`%�$eTt����?�!�dH��|\��E��f�@��F�	f�!�K 'X������%&ar!��²'�xI��ڸ�<��vB�YX!�$G50�q�&n���Q���*!�!�Ď�5Ӝ�w.�-��$���B�)r!�ď�����%�P�����+}0�14"Op������\SNx��I�#bH��W"Od� �t9�!�B	-M�$�1"O�	����P����BbǰQ�"ݳp"O���e���k!�Q@��j,u��"O^1C�ɳt�2��3L6{[J�I"O�5q�#�d��\P0��yY�xS"O��F��Y��)e.�-9��#�"O��ié�W�\ ���ߞt����"O�h���ΐv�r���M�%f�0
q"O��ԳR�
� ����H�U`"ON@���0x��gG���5"Or���G?_\�rV�J�Dڔ9;�"O�P�S�V�3��ـ�C1 ��Ƀt"OZ�2u��#|�l��+ -G昀"O� *�t�G7��u-Q�RBL 3�"O�,��n��{����3>B��b�"O���Gc3��e��ݬ�
�p�"O�p�8�j�blӿ����2"O:�!ų Sv�@�;m�J�"O�x D��k[*Lk&��,kGPl�3"O�m#�'�P<�-S4�81)�]�"O|Ĉg�P��<�fH);�:e�"Oi�N�-v�H�rƂ�%W�0"Om�TE]�PK�+�S`�c�"O�����˯��Q�JtL�<��"O�,i�N�3 ����"TEC�M��"Oڱ�E�G�P��\Is"�w#��(A"O�%L��bސm�E�� pJ��b"O�P@�h��HP�hݫ����"O �x��<f�1q�M��[a�iB�"O�1P ��-����b�~�4���"O0��5c
1���qB� ���Q�"O*�`Gݻt)"5����!�̀��"O�ev늌,~}����"���b"Oԙ�,ނ�a�a�z�8���"O
�HĆ��3�Z��K��\��4Ѕ"O,D!)�9i�`�f�$4S���4�y�F% �>Rk��C�̫�T�y�6�tD���w��y;����y2��'#Y��#c�� G�̀���ޏ�y�I3��@�$L�2�Ys�@��y��iɬ��G5z?Ԩ�I��y��#����f#�)H�����Y��y�lM�]Z�m�����2�y��]��X����*#� ��/�!�y��Zl
���hӳ"���t�T��yr�3b���Q��#!B¡HE,ˌ�y��ݽ� E
��j�� fO� �yj�!�9��|�v*�y2�K�}�ӑ�4GRyk��C��y��O"Y��X�ƀ�*}�ѓE�D�y�!�0BRaI����Q���4EP&�yR�yؑ O'%��%B�&Y<�y��	�{�t}��;T,������y��>n \c���j�E��o��y����p.6�"�Ύz����!�ݰ�y��3T3X�9S��qK���p���y�@|lF�2v*!��U��F��y�Z DՋ `� +�n1�)B"�y��L��$�����0�Ū�*T�y"�*�j5xPZ�|1v=�7�ʆ�y�@ލ4�ܬ;��H�";� 3���yRn�=QB�,���bU�B�ۨ�y�P�f����Ϛ#T�����yr��:V�4b�nCPP���7�<�y��ټf���Ha�"\��-h�!��yR�ĳ2����,ʊc��su��8�y��b����9Fw�) 2	A�y'M)2|IA��LA @����?�y��O8h/j�#���<Վ`�`ꃸ�yr��(��y��N2@���è_��yR��2Vt�6��#a�dqb�GT�yB	�!{��ԁU�Zn��󍔿�y��59s �a�$U�`X
m�yb�Ljl�8v��M�� ��
��yr��^�^|���1N&��`\$�y2�1����^�dQ��K��y�� V��O�5P���iD� �y
� ~%�d����Ɇ�G�Ԩ��"O�=��-O~qr�X�b��Aj�"O��yG)W 1�$�'��
C	�.�y�/L�'�ʜ:���,u�^T��5�y�f��R�x37*�
o�"����Š�y��J:5����dӴif8A����y���9R��  "m:_/�<)�U)�y�	8|)�q��$� ���A��y�G�j �PɥIC�(����� ���y���� #G.�Z<l!d�Ӵ>!򤅪��tA�.ZC�I,I�!�ˠ��bE���t!^�qr��9J�!�Ă+U�5���Dn"I�wo��@�!�d�G��#v�N
'u0BQ)�P�!�$�֐���x5��{��W�h�!��� QX#��������@`R!��Ȩ.Gz4��E�tl�e�c��'qF!�[r��Hh5�̋ e�8�H!�!�dY?v��dػJ؅r�&A7)!�ǣXvĺ�C <l�h�o�9!��E;+wְ����0eG-y�nɪWY!�D�800"eH��=Q�N�G!���a����t��1Qd�6�Ԫ!�!�$W%'���aj����x��Q3F1!���`�����F^�6�nH	���U(!��a��AS��'n���F&�?5!��ԬA�����E�L����d�T|F!��P�Ȝ*�K�Fȇ(u4!��t�
�3�H-8ۢ\I#�Q	n�!򄘰'�b����+�� .X J}!��5)LZ�ɀ�,�b	H�#��}@!��]Q>�I�!�5�4CE�t!�dҪ�")QƘ�[����fϐ3&!�D��zD� ����%����Va���!�DӳHy*�!���av<����p�!�d�!Y[d�@��W:����M�b�!���(��h����%m�:T���Y�!�dV�3"���Ɵn�p�:���:M�!��bcd1�&/@�{rN�ض�ޗC�!�@	ad��AU�@lp���>�!��J�=��cw�?&=l̪���`�!�-v���-����\�GG�!��&�PŐv͆�-�f��R,?�!�V�Jz�Ё�,�/�Z��ǔY�!�dj�@|�"h\!/��pj���'v!���	|��=���q�2�qq�5�!�DE&a]�\3�Գ~'��5%	�[�!�D�9v<�0UDdIJ��ÙN$��'WPT�%��27n����7Jr���'��QbD+_%S
��X��Ɂv�dJ�'Z�=;6�؂	y�@	g�;t�<�
�'��4#sFо5��,���Y����*
�']VE=X6�ٻ��-m�1��n1D������11!.5j��=E$D9X��.D�8j��p��\8�C��B����g(D����� ^2Y�%��_��Xb&D�|�W*��/N�@��O2�"L�D%D�x�!
iw�8�B�EҁY�(D�� f%�\�Kׄ^�9�A�8D��C.� {B<�X�o�l�VE9D�ty���"4���Ab"@fx�'�#D�t�`�M�=���3�@>v����%D�x�aHZ���E�'K�\��5D�P�r    ��=�f�H��т3t� �����C䉭H|���Z#D(I��֡*�C�ɴi`pYy��U�(r�Jվ`DC�;�(�Dϑ� [N0s�V>9C䉍,p��K��H�T0�Ei��<1�B�8����� �:lB/�C�I7
=Jq�Ƌ)98�es���7BC�	;k�0Tw�5s�9P�fB�g�^C�ə����qb؄q�j-c��=hRC�2l��`ҕO^������:�tC�	;��@{
�	�-�ţ\1\ZC�	�P ����*)ät��A�x� C�[rX)���4 [�0"H��/zB�	�`�n�����Wܸ!�"�,"��C�	:Xdi1u�G�h{���F���:��C�)� ����S.n�dH�G�,Vh�s�"Oa��E=� �q���=OX+$"O�ي#dG�AC�tѐ&�7���Ȅ"Or�x����W-�س&��I�$��F"O܉�P#
�8n��!�Z�!�洲"Ox�����.a#��9㌇^^�09�"Of�`�Sڌ�(��,'iz��f"O��VO�8d�����M�}U,��Q"O����������-JiK���"O�����Y>S����	��0Ry3"O�487)�[ �r4o�;��8`"O�aЮ�.#D53���x7�'�ڦE ;P
�]���a j.W1�A�� ���;减�Q�qO�>1���^���7����j1�E$���� +y�c?���*Ս��t�P
ro�8��'�<��i��UGα�Ì>,OPH�Wd��tܐ(�q�ڮF}ƥH�D4~G �`���3c��b�4��b?1��E�%-��ↄ)QA(U�U7,�����*2(mL����QVx���f@5lJ���+j�*Q�Cŗ:k hI��;i�n��F�%<Pv���� 6lF���'�,�ͧ���/�@���*��?%b��	 "��	Zq.myD�x6 �2���Q�)y(ؓ���b|�ىuJί3�r���
H؄8�'px�D���l�౉.Ӈ%���pʌ�{�ƴ�OP8�A��.�A�R>3;�A����s�O*�R��gFR�Ņ��/�Eb��'���S$�<^V���X%G*џHB6�Ew�b���-�0!
`�a�A�&`�T�9�KW�=�`,3����%�b>	�@�!�x��DU`z��g���8j��
��7�daE�|\�=)�$�Wav��S�X�p���2_Є��SJ�
=��A��<������?����s�X�Z�p�#)Z��*X�?�(�
ݥ(Ty4�E:��tDv�X��!F�XL���>���$�����#�7:���B�b�8^�NQ@A `���f�vղ%��B�A�	m����\�?�O���	��"�~4�,y�,l9�.]b� �(�'n�R��e##?�1��/K�Α8����4G�L2�fx��3��K>w�3�!�kN�	C�Y$s��o�7`�0d��m��g�2�d.A�l#JF?����q�s�6ʌ�i����#H3�.P�%Mr���̈́l����c	2�<x��]>�cr˛�u���%Z�"�(�
۽���y5�`�t(K�[�Ψ��a*�S�n*^�~�4x8\�����4i�z�zQ+�_o��E	2���C8v���o�,1�bT��Em����[��B�hǇ-�L��֠A<r����[D�@:�i�ym��E�ٙT�\	�e�H%P�`�wN2[���A�O(��D B�6{�����+@��r$H8E�b�u�۲{`��
@6��6-�a�]���[zD	�f⑑r��(��7d��8��G�h.9i�Q�FIz ��C��xr��)w�Fbƨa�O�̳�eL;�TZ��M�':�}�qO�<8_̜��iģ0a�&8`��ed��O8�X9%�NI�tr#8_B^����LP5�T�T��&$0v�����
N8�L��Op�H��F9]ADt�AD����"C9-�e�3AE;H��AQ,*4�Ò��:N`��!D���b"�/�Y��9��K�+�������M�W��$�]�7�詢0��+	ڜ���L'��+S+_�����y��-^66���ɛX�&�+.O"\���O�]��"�@��]k+�t�����|/��q��^��ft,@Z�3��,�|e�r�91.��s���Afj�jn�)��;ӂ;?��@ܭV(37������*��8����W�ŧ��e��f��J����Y~ITp*@h^me��� �:����'�ĥ��m�fFZ!J���kXcq ��#	D0�W n!@�+�>i2=�D��w\?5R��D{ ȱ�"E?aw4���#t��U3�4,~�qBD=L�B2'�۷6bju�R'�-N��tiĢu��m{3�'t�q���I�R��Am2Dj���*g�Q$O�
���'���"D���6(: Ǆ�� !K-O��nâ t�����P�>���c�]�u���t�2���S�]<��	�l@���I_�i�^�����C�s�浹ơ��U�A�	3p�(a��n�$� !&;�{��u���hu\��F�&�ʍϻz���K��H2`�]�"I�e��o�t� 0�L�HT,EС�'������P2 ��`�"�P�{q ؼ�~bh� �p��\������K�*��yP2(c$Ѕp�_�;��H�@Q��b��Ђ`�ɉ��'2D.�#�
 ��k֕jdh�"^gr���H��(~6�ҠE�!!�A!F���:����r'B/	RfAIR�U�	/P`MQbb��Dٱ��M��Ph�d1R�lOr���&H d�V�r�C�*?�^��@aVj�0`Ɗ�/%3@�
��ćPr�к��P�7���^�$�ZXXu�M�:�1OX\HU�,��'�TT������;!�(����D�6:����N?1,�R�(
K�ZH�q#����s�R)�����w0�u�fAϕ'Ժœ�/����'���jD�.&P�p�も7�lH��!ЫG?*����2*$pS�|�Z�#R�#
F�8p�5�d\ᇁ��,���M9s)\��
W�N���c1,OP,��k,<�� #	��GW���ϋ�_JH�����Xrm�VF˜|����ę�Z͓�@w���G��.q�$�"´Y��\�|Q`��O/����~W@�wON�O8�12l۵8R����A6{�� ʔA�4+���EEQ3(`8U� �gsdA��
*ܰ?�T��/��dy��ֿU�B$��c˩N� �ʂ늖}�_D�?�'aǭ�8x�.��v#�.z#:M9�'���Zv�V<2�kV� 0pːh1i��f�b��sc��g�L	���z&6?6yݕ����`D�Σ+�6���.H�K���뉯L�t�"�R0$f�����hx��%�7n��P6bBl��V�׈;RDq��9O$��1�z��K��g�? �@���:��y���φfD�̳���H�x����Z�w���Ba�ȂD�WmA�?a:��G��N��$mQ,	Yf��ϊ&2�t@ !J��L�˓�h���O�aXqÕ�Xv
i�7����X����0PU�gP��p�s�+�e�}ҝw���S�!��LRc��o�h�4@v�pBR$�JlQ���!<Oh r�ay�"�@�<�PW���Y �C^'M���$�P��0���T<�e�$N�?J���G�:�;��Z�����EH^�9�-Г�{���Î:i��)q�ըof Y�ۀ!E��7B�b��y��&ѷU��-X�d�!z'�E�Z
e�.Ԡi�8Q�h��%�֡�E�Pm���4�@ru��	�J�S4 ?��?S�-�)R�g��У�Զo*r�so��<�	�	�Ӟ�H�;��_�j�X���j_�~B���l�=5���̓|��m�����B�í���߼�"t��RC�I[��M���[��ʪG���r�d�7 a��� �ɹլ�
$K�/QD�]s�&�����k��K�h	���pNW:p���ף�b�Z�����`��G
�5�1&�	�c�^����i�t��E��
4�@m���N#I��A��.ZM&�(�L'��(-��V�d��UDC1�^]�!	�I��I�i�&4Aw�S�`c���4D��P̊�	�S�YS6M`��L�+��6��k�RAH���Bʩi�e]�x���h&KR�9A,-i�=w]ة��o�a�0�����w���[_w���#梘.Mj�$� �&y��Q1N��p|F�@��T�����Ś���a����T��a�Î�iI��B�ݝJ �+��T�p6�H�f�^/u�ݩPH�:mnB���~�f�Ч�ȃ� Æ&(0�����};�(����idT�J�!��}��q�t}�k_[���¨A<�D���ז.��m��	:'��YDc
��dY��4�0}I�а �fH�ЏQ�/Ws��\�$ |cH�hĺ��"��16��Yb@C%	0�����H~�@�Hj8y'�ؕRt �&�3�d��=7�P� g]-7����ÞM���c��ŏr���RS�_<4�?3�F�p�۟�ؐ�Oͥ>����\�K)B�U�z��� �T�"P"�+w�օ�t���Xڑ#Ʌ)%v�n97������}:-F�@����Ō�+LȈ��S"Z`�l �R��	���R��si��2W6-۩[��r$ͫ�E�
�V�Z���#D?D,ѣH�!3��X3��++B(jD�E�:��$Z�iJ6T�P�����A6Z���� 2�����gI�|mb����Q3[P��Øp��7�*h
��%�O2��@G�yfz��f�0?����=�ӥ�3�$� �F�J$�B�\�8_0�AHS	wc�X�T�C �)����&� �&	K>�� �0=V�����{w����8�LȂb9Oz��G�� K����I��hON�E���Q���__69�-��Du�u�QAy��	"W� �HP\/�vL�#��?����@�>�	W�F�9X�ݳ7Ȝ�m���Пs�0�#Ҩ�:�V,��o� ��O.x0$�ٔ�<�Y�_�~I�'��DؐQ�Pm��BW��i�K�ą\?pBIk��_0:H~�#��v�q,�����؜'���3i��u�k��jܓrD �!�\�r��l#��8;wh�S�����x�K7g�����vC��'r��tsv*;9vd�o��"��a�50*:�˕�[�y��T��(�RTL+�S>]���䑢<�yvD%y���)�0�\�a�Y�a@.�!��K�r%�KA�y
&�"pШtI2�x��D%dJ@�*�A=]�Nu��+̷D�(-��'���z��
�Ym���i�" �~��0�@
9�TQ��0I��x�f�y�������D�d��7o�=�����<�|!�ıH�)\{����ƭZ�!��J�N�F�*q��'�@��i��%��A,Y�9��J�K�R�Xq��
�t�ڻR_Z0&��.;�* ��nX?t���3�ŀ`�6�S˂��0=e�GN8�6%�]%����-U.�M� $D"kT����"�#gl�"%��EL<�;$ur� 2h��]�B�xG��E�PXK/҈T�ij¨�V�X�Rm�5%� ��Q��'��Ec��O�RP["��U�hD�ŻK�/o���c�h1V�u$]�j��)?2��9�pa�TC�ѓV��m���#sH_�F�C��i4>�)�$�?Z�ؐ�B�ZcF�:w�CJt��͹!/�c����k�8#*�E�e�T�u;"�Q���1D��xB	$E4vi��h֬4�l�	%"��h�� a�X(�6mʳB��prR?�I�jU�B�ED�L�ؙ���`2Lz#EO~�a4@b%ϾZP���j�:WDh�@6��5W��{���@Q��4�/FGb��D�F
YhUT�B� �R�ֈHAf�����5AU��;�Bo��B�X�
Iy�Ι�w]�(��Z���|S�@1r���s�eK|�� ��4c$	wY�sU��gNZ:���X���B��FIz���D�d�RŨ���%]�H��|�H `f*T�~7�x�ug�&EAj<�7��'�@|����	(<9���!p'�̠�섖+���`B�Rf� z�"���t�uRR
MC�F��a˙�*X
�&	L)�F��HG�~��sՉ�d��>�R�������3ғlㆡ�DH��IzJ���
A\BM8Ej%z�%�s�E="�� D�W�<Xr��0=|N��"K�G^�?����
�	�b�K�Gx�ȑB���{�j����<@����򮐜 z����._| �{��R�k����4��	�%F�=-w,]�Q/(u,t{ ��_l4��ҥb�����?�
s	��>�4�@sA��h�����M@�;X�!�2���~b�o������"Xf�� ��[Y�ՀV -�x	ⅆ�
kIS�I� �J�ꡨ@'k�YT�M7b��r̔��P��A��CO�@{�Ȯ&�T����%��k �G%�`�~!21'	P2��� }^��c�V q��Pe8n
��ge�:b�jJY+.(t�����v�#� װ>���Dg�.�qC�-_�W j9��9K~V%ɂ�\w�'	�}S�M_2U��d��X@��VEl��}(��i��s1˃Qٺ����4	̂%q���%A�~U��2`Jހ^�:�pQ;Ѣ"#�����V��㟰`�*�<3v���B�&ANPQg�O��p�c�G�<��Q� KZ/1D�:'#F8"�X���K�����d�(u:~�KB	��9��7�׶:Tv�P5FrC>��g� >k#K)%�l�����o��q0b�04�Ήj��^�ٶlN�(.8+��+�?�5n�i��4YP��	6�X��M#gb��"�O?���� b�{��Q0?3�YQv�^�]ϐX8���(Qf
%�cU�I�b!\	I$�VI��/(h V��gBV�m�fc����	�\�R�,�+:��(����+�a&P�y �
DY�����n�PXH����D� 4%؟'@��E���'�@����P5�`��ѕvL���N��tL�P6�N6S3Ui�D ��$K�@��`.�\{��rA�����J�X���P2Q	�% ����<�J�SSb؅�|U�<Ys��n}R�n3$=�3�U�7&�U��h�$$�|5y���(T��2(0���֐P!lС��D�L<�R��d`~)A��G�y�89S��D3*0���Q"��8�JK�@���zc�%}ȥJV��7���i��1[�h�����f5��(�ꋚD�����J'yƹz�̏2�� (��Q!�6Rָ�႗{'�x�B� As��M
~(p�Wb�.2�D6PԼ��"�D�b��ǡ�O� 2�������FxFi���Oܕ�'�`��g�T'I�4c��z����AZ�o�4�bb��#��-ه�-I���_^I��d�'�t��<�5�<$�`���iT72���)�LT��f&��]�tSP�#|��)�d�og����oV� m�qB�IR��vf[9_�l!#��џ&v�e[$.J'?�T�Ca-V�{�`}1f�;�	�z�jaq���4C�@���9�ry��M�c��usT.������bv��ra�z[nр[�?�y�0�Of��B�H�E۞��I��':/������J�ظQ攨-��I�c�H�i$�5��@K�l^��Rk��{�C[
d�>�R_d	��w�`pH��3����G�2U��ٴ�5�c�0�)�禭�����=~��TmӟZ>�H1�E~t��s��2H�6��� ӈ�^���'ǋ8u�<��-R�_*�AE�|vl˧��).m�0�w(P�$��1*�>LO�d(��q�!��oZ<A4rɂ��8,!(<����c�tXt��/���"�/l��y�nB�bղ�����>Af���\�4�"��wn�YCU{̓vd��h�bK�ըC9"瘅ig0�T�k�@ 1�PUH�j��U
n�1�� �N\�K��f�� ��Na{2�C�C̈�yQ��"!�iKm�h+(,`��V	Bb^�UѠ��^w %��SN���mT6, ��� �Р'��T*q�Q������+#XC��I��)S�`��o�L�26���}<l؁tKX3 �����D�d}�'��L��!  �j�\�v�Q�|>n�ӻ[��aA��ĖG|�� ��Q�]����.F�0oG�f)�w����n��b@�Ce��j��]�6�P�"0�G�(�%!dF�,5t�E8c�4��{b��4�ðo�>0DV)���G��'��Lѷ�O�p���ᐠ]F��r��)GK��8o�E��f�v����q�4��#��cUIg ?\O2}� V� ��S��+Ѥ�z�BӶsj���m������|��'÷
��|��M�,����\�Mf�@���
��hH��B�I*68���rI�$s�\|�b�X-v�6�H�.��A"�&+��:�Ҩ20���R�i�&�����
A!8-�f��*u2�j	�p>�ĉ��$1��	)rO�Sf%,��h�KY�k� �rWdM3a��A���'��%�f
1�3�dD$�L�	��@�X��eAC���d�&rƴ��G�
1�*�kg�33B�IB�L�;r$�(�/����=���>@�ոChƯ,�ܠ���Bx�Шs膮/�Ҽ)�da��&	̢"r���A��M��]8BM���y���)J=�2	��9hn*�OG��'ij 
��q^hU���ӨJV�l��bW�M��p�P��S��C�ɝZ��LY#K��N� �!I�M��ѱ�i�4���'���G�,O��)���V���p�FS�iB ³"O��Q2m�D�<�s�Nߢf����'�D Q4��{X����֦Tx(#�X�}��8ەA4D�h�t��Q ,\ˢmٱH�L�g�>D�pK���[��q*�J�]���1D��ہ�Y���,I�h�"� �.D�8K�T�5wZ}h"G]F7�j`O*D��a�쒌��Ȓ���  �����(D��1��"1`m*BM��V�~9b$k'D��𡔅�j`��Ǔ2�TUt�9D��{0͐�
�P3pjN�S�\��/4D���ԁǺ.�t��Qf/�
���@7D�D���G�݈��ˁwKX�i�i7D��YC��m*���ߴS�@$#A2D��16�#��	Y��X�@ �0
3D�੆BT�u��M�9Z+^T��0D�H�`G"N�}pЈ��F����.D�T�Ŕ'�D`	�C��Ql,D����Y���C��Z�Ĥ��f*D�H��oK�t��,�f�����B�4D��Cp��0f�*�v����M��4D���d�h���C��K(IF��*7N3D����#K����a���S�n0q��%D��JUh�
BZib��!��A��4D��	Q,T�f�.\!&��'[�D�y��4D���Ro��x�j��Qˀ9�@�c�0D�d�e�;s�P��f	Iv�=�(�ɎNy��@(T��K�T�6a�b� �戏b�4 �CG��,�bQ��.4}b�ΒX�����=���8b������tD���
p���H�W����0bM�)�'Vp��ծ�^w��ʅcçDH>��w%�.\�H$�e�)���/����u(V)Q�����$҅:w�5󢉞�^�`���?yN�Fǎx>�rp�@�!4���I�mK�����ڭ��b ����M�V�PX��3� ��BӏǆG�nQ���@I^�s��4�zhp�OnB⢈�0|c�2N3�u�c]�y֌���S�1w���ȉ��F�$�P����!�"L�=J�ٷ�C�75�$ɗav��A�>]8�%��?��v��*_���kFFD,	�ɤ������j1�$jI<E�$�՚`�܅k��W�C�ly��%\rZ���8Hz !���"��	(�m �Wo���MǧBʜ�*������d��0|���+@�Z�:��޿B��U��@��
D�E-s���3 D�^4�����ӶP��&Ծeo��j� ˚z}�u�!MKxn@�S��)�?��'?������yOP����%�\��5��	k\Bd��$���HX"��	^�a���RQ�&���M�X֭���n�,uKҘ[�� ��@��a�j��ç�ȹ"wd��b"~p"�ūr�� �1�|{F�� 6�G�~R֟�8�a�IU
��4�x���D�"c�VQ萐x�ɄE�a�䬑�`.T؈".:����ۂaω'u@���#J6�a�d�$)�1MЍ�
<X�E	LN��'6j�"�@�%92O�OO������*`m+!������4MҲ��a�O*\�oM/�~
ç��в���Ʈt�`�w�čϓ-��M�p̪��35n<���4�ܯ#,���-\��-YsnY�@���2�'��q�S>�Y����$)�F֧����`!e=�	��~�����<�Oe��c�f=I�d�#r�pU�s��� v!��ِb���RL�k� Q���	�6I!�$ڤ�P�F�4i�ڤ�ͮH�!��'t�^�8�K�,Nڈ�7�:z!�D(1���h�O5PAPm�3F�?o!�J.@�)O9H�|�f��'kc!�d�<���y!NX���p83�R�_�!�DC<���2��3
�,9[t�L�u3!�$�<q��A�/��=ߨ�����5K2!�D�*��bbET:��PΐG�!�d��1�F4�P�@�%�B<�s�K72�!��ZP�@C�e8x�!H�&��#�!�d�s�HD
�mK*e��[qf�'�!򄞻_f��L�?+YQ�״"!� e�2�(��6���c�N!�E�P<)�c�D�@�^��Ǟ:!�_�cbų�M��:�T�@�!���!���Y=��Q��&az\H�G)
�!�DѮ{�����z.��.��c\!�d�Bv�P ߀i����Ԃ N!�Ė72�"D�u��,~qA�H)�!�䚼O�,aɐ��
wb����	'j!�T�j���'%j���c0.�O!��E���mΜf�����hU�C�:B�ɫp��!s6-���W��hB�I9D�40���s�H ����TB�I�M�����Z$f�x���"�rB�I8p� �]j<e��*ɕ3�jB�	3�$�[�'�'���шF!	�(C�	�?X���Eҧ^�c��5V�B��)V�48�� ��L�a�*��B�I�Q�>u�H��HV�̳ma�B�	L~���F�x|�&Kw6�B�	�NĐ��%�1H�X �%ƛ-\:C䉋'�!ȖG�W���� -���tC�ɸ!��D��+f��r3 B�8k��E��ĘY�u�-Ha��C�	�F%	jdm@%��Q�  �;y��C䉋qi�02v����Z�V�xB�	X�v� �C�5Mp����WRB�I��I	�A�'<<�C���$��B�I,h3�4������=��J����B�	�Q��q+`˗�f������ 2 C�I�B?�������Y�����tC�I�}�l�0�ƃI*h�� Ɖ~��C�	�z$YS	[%I#�{@ L" @�C�)� ��!5t���>a�8�"O�][�iwv�x�΋�PU���"O�<��"�?l(��]�GF�(ad"O���Q��t��]��K�1F��H"O�0��&Ӄz�8���ʏ�I�@���"O~Q!�b�E�P1CD�`�$��"O8�rԈ�x�N�+bjD��S"O�0�=[ ��L�xƠ�"Ot!󀌪y�f����̹!ݢ��v"O8ݒt,�0`9�p�A�M[�.�9�"O�9�s"� (��5Q�НD��-I�"O2] #��#��������f��"O�s6�<���sf�ԭv��xp�"O���A�E�tZHD
\�4���"OV��ġɔ#�$��MP�c~�|��"O�EpЌ��mHtA� LĄ x��3"O�T���6�j�YB,�S�.�1G"Ot����K�U|�P�*<i<�Q��"O04ۤ�ƟA��(�oHGT� ""O�II��^�K2Bm�N?D��"O�p�G��`���IW�Ky-|8�"ON�s�BC�e4ҥ��Ù�"F| "O���G�ޏ6)��IA�=�8q�"On�[c��&IUH�Co�'2a90"OT� ��;V�X�q!��m�1a�"O��E�I$ބ`'N@76 &"O��3��=Hs���wLαy�L�2B"O�L3WL�2E����Iu޸��"O����!��c�M`cH��9w6��`"Ol5��$�7�-cr̎� N	ړ"O0�Y��߳J'lZ/R ]��"OT�5�<6�;S�/e�M�!"O�	Y��A�$k�j�)U�L�F"Oxu���5,��)93��;S< ""O�Y���M�i�FE�'��;EX؈"O�<�cF�o�`E��&A'E�XA"O�8H��J�!��t���65$ތ��"OD40�%
?x3�)��I��(� "O��s���:�C���г�"O�ȸ7��xzൊ D�)]�FH
F"O����E�h�n I�c_�0��B"O0���jROy�Y���� �%�r"O��@×p^b����E�@��e"OrUj��Ԓ,j�-a���"~�0�B3"O�x&�Q�aX9͹J�bT�G"O���C��~�
`��o)o�ٚ�"O�4IB�;LB��P�%.qZ�{P"O8�
D��tUtx ��V7"Cʌ�4"O���v��n\���&���_���!G"OT�@d
��X�"��Y�k:T"f"Ob@���œ2���:a��#���"OX���]5;��0+��X�]\��P�"O� �d�p-��Q/���3A"O�����եuLp����sԔ�s5"O�L���S�H����恅|�ܨ90"O�d�w��Ff�3� �<�!"Ov�`īN <\8�B�P���	�&"O��j��ۅ=���Ibb�1$g����"O܅����o^���0��fPD1�"O�%xB!�.,�(�2dR�.Bn�a"O��c0�v�L �J�wN@�"O�͛��Y
%�R⨈3l�bX��"O�E�s+�)a.��1h���S"O,9���>>��ɴK)s����"O� �]IA�գp�~��q�{��9��"O(x���n$���E	/?�BM0�"O�`��Í_���r�dF2|uj"O }� ��N~��Zv�B={�	"O��HG�H�uN�<Bs�g����"O��EV�y�d0"�N�/i��7"OH�Ӗ�*;��;�F"2X)"Oह�&VW@ 9
w������+D�D�4��-R��qzr�μ��� 4D����̄�ZQ~5�2�߻- ���)%D��0��֙{Ȥ@��A�1R�L�"a!D��9ul��`gV�j�'�P��9��"D��y�T�".��(ۤ#n�q��?D�@��ȃ� Wn}���/�����(D��b�CL<�2�ە�
�?�q�(D�t���ǯ-�~��Q
3K�Yk�1D��3����jyl�؅�F�v$�i*��-D�dCqK��q�hI��~��@ D�4S�I*_���d�}�p�2�?D�h�E�A-|����C�	ez$���0D��X�B>���Z�lB& z|�B�+D���F�ԥ�����Z�(@pP
t	7D��	7�8L�x�b���34��c6D�P)�k�"�p��W�D,j�� D���d�˥?zP�iR+h><�9p� D��Ӗ!�_= 8���3N$���<D�\9��.,�>t�MP<zb�{#�;D�,�� W�Z�Qֈ�J�>�b�%D�h�!<ޖ�G
�+A ܛ��"D��1UF�[�>Er� X�p:�i���;D��Xd۬(C�� 1�Ȋ���,D��Nʮ	v�P�e�C�Xm���8D��0���S��P 5�UE݊:� 1D�x3�a��f��*�ҹ!�6�7d4D�`P�L�TX ��N�3�� �"-D�h[q^k�N�$-�N�����7D��C���	w�j1Z�B�w��d96$;D���c# p��xS��9Q���ul#D�,I �	"�(1W+OF���C�<D�x6O�>?e�����H���
�7D��i�C�K��9�WB�7_X�!�E5D����D��H�4e�b�4���G1D�����)	%�=�0 T�r�8(Pl$D�|���ˉE�����O�(�W� D��9ry�d@1��=P���@+,D��z����ؤ��Q'���ұ�&D���5f�f�ĊS�ц.�,ee?D�h 4I=]�6��a�N�"��`)�#=D�؊5�кp�^X�T)�&?l�� �<D��
 0�`��	!D�P��2�=D�p;"�`m�5gO�E:D�T�&J�<�:=��T
-����+D�<[G�D�9Ÿ�82MH�O�ze8Qk-D��R%H\�(.f��F�p�zi���+D�Ȋ!�S7{�>�bũI�p<(���<D��ZC�!���k��1��C�*<D��zD���+ﺜ8�.����(�7D�Tc�g��)9�V�m�X�{�5D��Q:XsH�A�-j�8�{u�5D�<3֤�X��hyAAӃ�(���j1D�� R�Y0mGd���{��	��A.D�4a� �;Ԕ	j�؝E�v��E-D���R� �
�������f�Y��,D����c�+$n�Bf�߄|Bɢ2�)D�� �Q	ui��F�P<I5���b��ak"O�2��������n0|��"O��1��a� ��@
 nYH�"O�@2��5Ɏm�%'Y2�x��"O�	P�Qr�v���	��Lzy "O������nx��c)[����%�Py�NΕ]n��k��Wp|����X��yr"P2\�$��@n�la�аa�I!�y��N k.�O�	fBz�Y�̠�y���/0w��b���H�J�fJк�y2*J$y�V)5)�Fu�(�MJ��y"�B�w����'�n��(���ynڱa`�1*�.�<2���E����y����(�&�Y�9>�yDf݃�yR�X>	b������0��D�R��y�ƅ2e6�uA7��h*���c���y�(/:H>\K��ٰb3`q�q"��y��HƝIB.�^�~QRԆE�y"���U�D��(V�f�i�-�ybF���x��n�a�@�*7�L6�y)F�
�ʅA�f�3$��������y�Q�Z�\{��ėQ�҉�p����y�J�
h��L������yA����Ex5�[O�:��gG�y2�I2 @  ��     �  d  �  �+  �6  �B  �M  �W  /`  l  rv  �|  �  m�  ��  �  4�  t�  ��  ��  E�  ��  ��  (�  j�  ��  ��  ��  ��  ��  ��  � � &! �/ �9 X@ �F �L /N  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|`I!'G#\���%�T��'ItcbꀀK<�k��̥:O��'������Ǝ8�ݓ���"J�S�'y`=c �d���	%�BPiV��o�<)E�I�M��c�Q'��I���k�<Yb�`��s4��/~�����M�e�<Կ��رD�E�?�t�Жgd�<��j�aZ����Aّ'�F�r�b�<��"���e�ďfe��ѣ
�[�<Y �{�<Ԑ�[�0�Rѳ6aE|�<�ǆȕP�,x��H�o���ۀj|�<��\��!G	��lhP�qI}�<�cێ�,����ޣ��@�#��x��G�<��Fъ��u��Z�JQK�%v.1���� ׋� ^:�Bэ]lr"�&���I�-4��Bbʴ9[��g.A�$&��$@?�vĥn9zt�&D��v�����Z�<�5��@e�
I
p%j�a�L�'�Q?y[��Ph�d:�
�Z�bg/D�$2��q�HÄG��R����I�r�����䕘!��8r@�P�Fi�	� ��!��̲��u*4%#\l􁦪��,�du����	�j�����
���k�h�7EB���˃���.*����u$ML�BQ���C���C�I
|����d�2�y�e#Q�B�	�� R��g� �t��B��1�s�Ee� "<E��'�����?l�i�|����y2�6�Şw}��̞�� `�d�ǁ���a����dE�D��p�i^�;>��S��%+�|�L3}2jN,m��+�lRu��iT�y���>�����Q�g�عQ� ��Mˌ��%��|ph�9IV��1�!�;qu��UA؞X$�>�XR��V�ԎPԜa�g��:]&���d(8a�МA��řcYx�h�G��%ڧ\�ƠB�!3]��`��G�44��^�Ȅ�-J�S�d�Ӱ%�'
<�'Bў��$��Fa�,ʕ0�i�9j.!�$�!i�;��@�f�I�Iſ+� �牰D�-�Dk�;�Q���c�C�	;<�4Qd �
����'�4��'��Bm_�K;�HاA�H5���|�����Hȸ-&�tbr�Žp#��v�/�yb(Ͱ6��9�L��o�(��^��~�!�S�Oaƙ�gh�[8|`c��e��e�'% �;?ʡ��� J���
�'��s0i�3y�Bd˖��Vy~9�	�'�F��A�^_8@�D_�M}F��'����7�[�Y��:C��JF���'�*ex��N�d�B��9;� b�''��SѪԮ4	�#"K��7cL�8�'����d �el�0J�g#����'�HS��Q��*�р�	����'a�|@0l�9�0�p�A|�`<��'/x2���93�]���:%���`�'W��P��҈4�����)뎨2�'R2K����y(J�0�D�Z"m��'�~���j�$)ԡIg�0����G��O����^�E�� �9rdx05$?��{rɚ��I�m#��Q��Lm��$*Ǹu��ʉyr�'q�x��H��t��ѯ���r�H0ND$��=�3U����"��M�霂���.�69���ȓAR�L��/�B��ǭ��-����=���?Q��Ӟ6 ʝ)��^�%x"T�&��~�<Y���7?=f` ���4~D|9qM{�<����J�Fa@o�`Ѡ�sS�Q�<�[y|�d[� r:���`n�EB�`�'F�|�ڮe��)҅��F��b�O���	^���O(���b�>�bI����O��p�	�'eF�Js��#y��L�Ǆ�U�
yK�}�x�鉷4��9{�ɐkL����N4Z�rB�IlZ6�+l�	<�ؽ���Pdֵ����'] �cV�`����jG�%��9�'jX-���_�"�ba던�Da	�'�bY��R&��l�� ���$��˓�(O��5,��N�R$�7/T�j�~�J#"O�BS�]9af�K��G�Y;b�s���=lO�A��ydVEk��ה:0��"Oȑd<$�X���$Υ|����"O���t.R9ǎM�1���S
nj`"O�:AJ���,������eh�ha�"O\�!��שn=Ҍ��$�	'�<Y
�"O��#@E�U��C��W�9���"O�؀�J��}:5��k
:�P��"O�D�G@فE5ZA�Cj`D����7O���df��	Y0i؀}�~��)I�5,�,���'���ɉi����AE\���z�&I����5�I�|9������?& �S &�T|�B�	���0p#� ��� �<}��B�I�Jz��5B�% dY��T�A�6�F������ ��A��ƛRTV�BpH�>���6"OL�ke�I�Z t�A��V)(��2dU�p���h��Q#w��
T�� s!�F�H�ZC�I,A:� Iv�CQ��2�iħX+`B�8P��(��_�!�l�s�H�3
R>B�I�T=dX�!��N�ZAz���._B�	,$��rVk[	l��-q-�)
B�I�e|Lru���Z%��� $��>r�C�	0����ThW]jP��-B�6Z��#��c%O�>�ȉ0�F.`�����4�O��$�QԅƪuJ�AK����>���0ƈ3D���� 	F��AƂ�5�a �M2扃5���?�|b���b�c��$��iIGhd�<�0�� T�4+	I����a�`�'O�yB	Q�$�� ��>;L@�cc/_1�y��%&�&aYF.đ-�E �Ј�y�C���v�Pg:��P�7J<�y�n 'Ǻӑ%�0�؍qbC��y�ώ?~�Pt,(t������	�?����v\8���,�H�Pu��!i|���ȓ@��-Ӥ@+n�P�Sd݃B�v,	��O�����!3��q9�(��D���fcҖ^����)"?��,�;�2%��۷�����(�f�<���H��z�eZ�j�
1I�<��l����v����¡К3^lm��	�!n��M{�O��e�k�!�"��"bN؜�"O$Iǣ�W�$�����w���S��D�O��s�{����P=j��1���{�|x{V�D˟̄U24�K4�ҔT�X��CDP�(��:g(I�&�ݱ*�������>�rԇ�,�*I�K�J��f�3��!�ȓ%�M�adT/J�������n4�ȓ�Jt�0o�zB]��j�b���^=�P������[Ôpc���ȓSܐ�bɇ,�����ODN�ȓ&��MJ�� m=j�%)F@�م� �]Y�Fѫp'T�C��J�[@�ȓ?�,�B&@�����1FTl��b3�Y��N��z�	d�.n�B�ȓ9����[��䪧(Ų!xPl�ȓI�@��Q�(]�r�I�Z<��O6�dұk������@�]�(��׈��H $��<1ѧԗk����n�hU�ݢh"69YŨ�<�\�ȓ[�p�Q��L�r��a��_p&ȇȓq_Mb�o˗%�@$�+�# �����<_p�+3
�h�F@�3$����@ua���7���9�'A.S�\�ȓ:����<%�.��P)��(����|��6�Ѯ#���ޠg��=�ȓ-�E�� '��ߓ4�� �ȓ"cr�@�0!{�	�fΈ�
@�T�ȓu+�,J�$��P	�)+vN6Utz��0܅�P/ٮr�\��v!�h��x�ȓ^��`�$5)x,�N8�f�ȓz� 8��O�]1l�RT"�39���ȓ{/������-��$~(�ȓi<ش!ĭ�_<"c/ק!а�ȓi�Y�&T�w�^��n�%4P��ȓ*�f�K�JB�$
��R�ĩ�ȓx?�W� ❩3 �.��\��`�Y Th.���)˯vD�ȓM��R��+�:v�Փ"6E�ȓz #U�$ut�A��7-�4q��S�? ���*E��t��Ś���(&"O�"&H�8��U��e)���u"OnQ�A��r<x�D+^�@:8�W"O�h��&Y���k��N+/���"Ob�p����U ro[�[Ά�[��'��'��'��'&R�'�R�'Ӡ���J<OT���ʗ/p�4���'���'t��'�"�'A"�'�"�'�4�Q*J�$BLc񧆈aR��!��'�"�'HR�'��'42�' b�'���D��'�� �1�u�3�'��'���'���'���'���'h�v��k��<"#��>2\�E�$�'���'���'vB�'R�'E��'�Dm٣��"D*����Y�r<�f�'���'���'>r�'���'��'&����
���`}�&�ȐF.Jp��'/��'���'e�'1��'��'"�����5`�P� �R�F�RC�'Z��'{B�'>��'ub�'�r�'@����k5c@�A�*�-5������'���'�r�'e��'or�'���'��)�ը���e��Ȓ?'�=�F�'�B�'�2�'#B�'7��'���'_dQWhV gg�0S�M��˂�'���'%��'��'Q��'"�'���AЂ��t��!�,�W�'{��'�B�'���'���'+��'u�� coK==�vlz���f�R�*s�'���'��'���'R�a�����O�Ձ��	{����rrgjm(*O��D�<�|�'dv7��%{�l�ƀ�M�hX6�	W�~����d�ܴ�����'���FnM2]i���5�T���*G;��'�:���i5�	�|*��O��>et@2`�h6�IC��s@��<A���$)�'~K\�9���[Uz�	6iǃfc���&�iW6�J�y��	����]2T����l <Px�G[�s�$�I���ϓ���i��6�d�����	P^j�p��?6���S�lc��̓"I�~�����'����J*�h��q�
�#�Z���'~�q򉗤Mw��N�	�|��(_-��h�c>����>���?��'M�I�F'Uc�M�7h�X��E�ԢQe���?��۰Y�Ȝ�|���Oʜ`�z�:��/F	������G�&Ѫ/O˓�?E��'�bi��	Us�ZȊ�#�O�xi�'�b7m��r�I �M���O�P�Î�3x��Ǭ�Gঁۛ'�"�'��$
��v��T�'h���O?Z��B�{��	B1"��;e��'����$�'z"�'���'N4��� B�U�ȑa@)?�9IW����4e���)O�� �	�O��R��T�Ttʓ�̽6}60 ��M}�*s���oڇ���|��'��2o�S�]QsF�Z$"5i" �6 #�հ@OS��� H�Θ �B=֒O�� r5�E6��#'mF�:f���	��M�ЄV0�?�$Ѡw5 ��6��&�"���I�!�?y�i��O���'�7�_�i��4r��(H#��aU��*��Y�4ǔ���b���MS�'�"㘥8���S>p���?��_cpv����P�����%�z�����'M��'��'7��'��O��1;�'�0X��f5V��].3��=��'��Af�˖�3��I�T�	Uy�AѠ)�8�J�,�1��B�#7Xg}¦|ӎDl��?�x��Gɦ%��?���^h�P󐥂�Z��U�ԡ3P�wn	�Y�������O�n�?���ߟ4�� ):0 C��up�1��]�N+�heN��Ok��ɤ\�"4�CM )UC8���џl�	�M#��&<,��X;(G�s�`V�y0��ϓ4���_��yB�'"�f��	Q��]k���OP�i��W�Q��s�i L����f�G`,�xW�8��d쟒x*�D0�O��R�K�J���prCT��2uc�D�O���O��D�O1�
�l��J�l>��#�/Y��ԑ��A�/������'���o�,�R�O2XoZ%�t"���-���Kŉ��SX�)r�4P���MS�IN�f7O��$�!0T(%��'A6�I�<D�3=Ƥ��plԅGfJ}���D�OZ���O���O`�$�|�̏�Tl�x0��ڿD�⑑�É-^Л�dT�d��'>r����'�X7=��P��ǇK֩CEOۢ�f�Bh���شw鉧���O��Ԭ��s���>O�	��-���T��Ân�bpw7O�Щ�-	4�?,.��<����?a�兎l%*ёP��'��i3wl��?���?�����Ϧ�*��S��t��ƟL��(M�h΢�3gCQKG� �����'����O�ToZ�MKR�xr,�'Y��(v�$^����Υ�y��'�N��0�(\l�$:eX�h��r��!�i�bҦ��c�_6N�X[�J0D���'"I9 �Xa6/۞RTD�(�e���$��4�a����?9R�i��O�N�xC�!��ك���?4��\��۴U��v��s���2O�D^=&iX�3�'wC������.���.iW�`(r�&�d�<����?y��?a��?aD
\���	0��.{��d��?��$����FMЂ*���	�?���PyB�� RL��s)˨Y�h��[�d]��5�M��i`�7�K���?��S�n��0�'�%m�TC�'�/:���ք����N>dvčA�y��O�˓l��L�ER��tnV.j�ƈ��I.�M�ej�?1��@�a!Є���Z}L�����?C�i�O���'U�6��H�4x�r;���,x8b�N(V@����'�MÞ'�2�
�7�>��S Y����?��\� R�;��x1dn�	6��B�6OZ��$��(=���цܭDϠ�#�)
c��d�O��D���e�� J"�i��'��ęf�ŧ
d*�A�	�7H�D�G�*�̦��4��g�M�'��ʈhBF�2E�x� 4(�lA�=*���&�����|V���	�����ҟCcٗ^����r�=:�ؼ�㈚����	xy�,m����O���O�˧k��5��$��lА��k�z��'���[��v�p��&���?�g�X�L�h�c�	$1t��Sg�qΌyZ#�V�tE�'\���Mǟd��|b�= 4m�06�$ ZIO�?�b���O.�D�Oz�4������I_B�S��ր�lZ��e�ײFٶ���D�o�8!ȆU�(�IB����$�'-07�B!v�
�t��[S���Ѧ�	%�nڰ�M�&�E��M;�'�
�37�N�_���H��'"����ύ>):��DmM=��lb ��d������ϟ���^�4�t����6�ش�����3`�ܙ��i&d���'7��'P�O6��~��.��Jpn�W� e��J�ɏ�7q�yo�5�M���x��$��5qƛ�1O�D*�&�2.�j�ЯՈL��%(�0O-�S�-�?9t�2�Ģ<����?Y�a��wʄW�:3GD��c�?Y���?����d]��eR�/PyB�'Ъ���[�SgƌB�F�; �a�����Y}҆{��mZ���[��4��ԖP&�\��lG�^�`p��?�d"I5sYt�1�΅����q���n����j�Z�c�`Vb�@��Ѕ��H����O$�D�O���(ڧ�?aTk�"Gǖ�2*�0*_\�:��?�?y�i���f�'�d�\�;�4��@�b	6�`3�Ԇ��x�<OVpoZ�MS��iw�͡��iE���OXa���&���K�;��хe��k�c�0�O�˓��O��� �8|R�Ȼ���1��D�P��`Y�4X	:8����?����OZ��@c�_3k T�K&iHC-���w�>��i2�6ͅR�i>����?	Ǫ�����='j���/D;��b ��Myb���	K�=9�͎o�Q���b���ܖ��A��sdyk���5N��1��8j�X��L�4m�#e�Y��<�&��__��*G��&>	�f�&*}�)5�^�}N�<iu �a�Y��.Ò/�����Y
-��R�=P��B����ɒ+B"c��t�_/It�0���S��}s�a�3�`�7�L��h�Z4/�2-
Ψ�S���r��$��
���j�2ag�Ѱ	K��C�#��x�)u�aF&�dh��2��. ��i�5pH
9����"/򽢀�ty�ǃ$���R�F�*�����J��x��#��t�!��r�d��O&��<��O$�$�#]���J}8����pc��r_��T��>����?Q����,�y'>��@��X���i�(e����r%X�Ms��?-OX���O��� �,W�.48��Z��VӳϏ,!$��oZʟ���jy���>d����D�k��Y���B�	�^�1��G�6[�4�	Ο�P�h)�Ο4�s�N�3�"�PH�E%h��A�iy�ɰ_o*�I�4��S����!��D@�en. �C�1�Icq�J�@u���'s2���x-�i>��	�?O�<	��ܥEYl�H��M�Z<�E�i+\ŲTEk��d�Oj�d��ze%�擪%FznmC��M�MGz�R���M��JS3��D�O*���1O~��W�8}F(�v��zO&	�T��)5$ml�ß����*d�����|2��?q��y_�,j�
�;}k�� ��
;�	����ɰ@�Nb�D���0�ɼ/^�I� �,�����.����#�4�?�֫
R�����'�S�Ln��]���z�Ǎ�q��
�K��M���=����<����?����D�N��9q�E�"Ih�M{e�ۄi��J��ES�����	˟l�'�r�'qH�	���*U����0�P1dT,��'���'�BU�(i�mD*��4��1\@p�s��^a2 �������OB�D�O^��?��Y���O��-j��̤@�N�3O�D�n�Y�Or��Ot��<�@Ɠ	��O�ژV�2R�*�u�әZ�ޘ`6�gӊ�d>�D�<��s�'���K���5��&�ӖFČ�lZꟜ�Izy�&�G��0����k�G�+"���A8ig~�wD��G�&P�L�����I�2���4�s�� �q���J5 ��qF��Z� �i7�&A����޴%���h������<T�U ǯ�+GdB��e�Y���'�ҁP
5"�)b�g�	�kk.�
�fީO/b�d-	<R�6-��u ��o�ޟ\�Iԟ�����|ri܅��u"G
Ʀ�2�~h���??@��ٟ��I�?c�\�I�}$�ՋD
�^(����.r�P��۴�?)���?��Y�v�����'	"*��;�8�S�պ9-�X{b͛���?y��F���<���?��'�ڡK�&�j��h1�Zut�Pش�?���З���O��$�O��ܺ
;~&p����8�Q��>y�JF/?{�=�'���'j�I˟�*���{��f��-8H��і�i��t�'���'����O]R�s�j��1e�ac�k&��А�����ԗ'I�М_��IJ�`�X)Ec)W��lK�K�e����'���'9�O��DU2HSj�ie�i)^YQ�ǐk옼+Ђ��U.JT�O��d�Olʓ�?�hR���O��Y`jY�^���I� xѰ��%oݦ���O���?���]�.��$��@AÔ�u����t�^�^d���v���D�<)�;�B��)�|�d�O<����'��	H�oʃyS�x`,S�?����>��[r2��ώA�S�T%�-"����dV6ũ �����D�O2����O��$�O�$�J�Ӻ� T�c�� |��ː)Y*a�#P��I�b��5y��<�)��3
6Mr2(�)m1���Q�'��7���IO��$�O���O����<�'�?!��C6!]\|9��B����s���:��(کآ�s�y��)�O
tRGFO�����"Xy���%�æY�	؟4�����`�����'��O��F��s9�J��~��@Zwe�n̓M��u����t�'��O(��t`�(+C�ub��*��p�r�i�b��"P�՟x��� �=�eج�� �R��i6]+U$B[}"J)n�����O����OZ��?�n3n�Ti�B�Т]A�H�G+V�5k.Od���O���;��۟x��薍I��l���p�����Á�u��%c��7?��?y/O��č0 ���Rע1�����W8hp�"L�Q�7��O�$�O|�`�I�2�����Nk�pa�DJ����]���8a%^����ş��'�a�;V�S�@"��R�<����Dߕ����5�M#����'%�N��E����O<����2&��!Q��@�4�Ȥ�Ʀ-�Iry��'Ɋ ��]>9�'i��L��S���@)ȵ�(��&X�R���<i��x��u'�:@_���)���T�`����$�O4Ha��O��$�O��D���Ӻ����uQ�	¨}N�{%�Tx}�^�`Q �/�S��>Y�=�WnbqF��Ge��s�7��J�z���O�ʓ�b-O��O�3�㍶�f �����2lQ`�l�q}����O1��$�6$j�MS1��)\'l��6-E�R��n�����'A ��V���͟��	\?!�k�"3�"5#�M �8����MD1O�]�-�]�S˟��IS?Qr���Jp�FP��(;�J����I�(r�L�'3��',2���E�.mZ��&T���(2F�`�I��R]Y 9?!���?+O��dP1	"p�� �+�h�����m%p�0 �<���?����'X��Ͷ��4�5	H�RK���3�5V�� d������O��Į<Q��m#��Oc�� C�:D��cL��)�۴�?a���?��'����W�'�M��C-"$T0Q3�b�3�U]}R�'@RX�|��� j��O�¡V
|�pL)R+�/2�(��P�Q�6M�OJ㟌���n�dYW�=�d/h`5`�@���S�� ��F�'5�ݟ�з#�W���'��ONШ���V�K�(�᪂??@���=��ϟ,���G�%��b��}�Z� h��i��G\2�R �'j�g��>���'$��'���[���Ky��D6A��X0��\�B�tꓷ?�v�F�y���<�~�U7Р#'�Yb��袀��Ǧ��F՟<��ן��I�?�����'<�bt�X
	�F�y��=I��aӆ5:G��E�1O>���
b��`��(W��ܴ��6v)�|��4�?����?�ˊ��4���$�O<�ɴi���@!��)�`�h���*��`�y��*�~���O����mJ� 
���y%�G�m6��OR1x�C�<!��?A���'p�kӬǚN�P FK� eҝҨOL"1�G�%��I�H�I^yb�'���*����:#f�'u5ʁS)/B��Iޟ��	����?���<��h���U�no��kgC�p�F�y҅�=D��H�'���'��	����7j�S��IŖ�j�04'��<"�KA�	ۦ��	쟀�I@���?� "� X���m��"	Dͺ�m�_>xa���n��?	�����O���«|R�'��h��H�6t~6�ڠ�ZhcLd�ݴ�?Y���'�Ȍ��\�����hօ��"%�w���`�H1o���'l�$R�[��柼���?=k��̊��gB�-�=CR�α��'�B�2�̅��y���A�i\�p4��a�� 4��Gp}��'��$�'sP����@yZwF�P@@]+=�`��ٵB�HS�OX�$��W�P�a����I*&&� ;��V��3��&x���f�`���'{"�'�T[��S���1QH�K$�aQw�o)��6	�/�Mk��N�S�`�<E��'.5BD͇
QpT�Ά3gyL�a�jӈ��O��$۞\;���|r��?��'Hl ��H/r3�A3�ɽ�`�t+9扼6,� K|���?��'a��a�H9B�P�6�����4�?A�,Z����O\�$�O����;Q�����\�4�j�	gH�>�Q�+�Y�'���'��� [rD@3GF��[�]!uI�䳕���vGp�'���'���D�O<2��G�`���g�]�1-	:!٦M�������ԟ�'5�@�iH�iץ.����%q���c���&zțF�'�2�'��O��	
W�� ��iW����\�w�b{�CT�7E�� �O��d�O&ʓ�?i!�,���O�L6GߓV�㓊�\zƱyq(JΦm��N��?)g�Ů��&��P��[�(�S� K1]Tr��S!c���İ<���P�Ȭ )��$�O��)F�]E��c��H�Ƣ�'I>v��>!�7�f�����p�S��!��|;v���dɣu�p|��N����O�}Y���O��d�Op�D����Ӻ#�/�2�쑪���3}xrU�O}r�'��`�/L����O��uiӏ-&,vu�i�H�"��4����i�B�'�B�O�����L]n��0���<.����Ҝ}��$mZn2\#<q����'�H�K#hF��V�%.� �F!��Af�R���O��$������'��	���S�? ©G�x:$TX��0����i�_�T��@f��?���?G�٬ǆx;�G�"/Aޙ �� ���'OX�QdJ�>�(O\���<�����h��|a��E[�:�H�}����y��'���'o��'��Ɏd�䐀T�d�����0<D|I`j���D�<�����d�O��D�O�d%,ܡ
pR<���V]��E)�b۵�1O����O���<�H����J4'̺�H8>�9 $��0ěS�t��dy�'���'��D
�'6N41�o��T�v�� �>�@ [Emx����OX�d�O�˓Lj��7Y?u�I�A��̺tN�b����
Vz���4�?Y-OV���O���D��[?1�㘨	�&����
>����¦��I͟\�'�����"�~����?���k�6��$�y_��2��m�.O���O6�����IXyRݟVt���Y0��Pp*?�bR�i���{�V�R޴�?����?��'#��i��A�L��dXIU��P�XREzӚ���O���d<Ox��?1���U?t�xE�G
���@ɵ�V�Mc�cR�/����'X��'��t*�>�*O����'J�'��T�]0�
)R����U�Bl��'�H����;U>X�B�ۥa���k�ɧL��ݛ�iz��',�0{�$����O���2'��80$NI|7&�b��=��6�6�䄖2K�?9�������-0w�����wL�=C���WN�A��4�?��cϰ��v�'&2�'yrb�~��'\b\R���)rT���'vR�O6I��;O���O����O���<�	�2�0JOR���<��d�0z%���S�L�'��\�H�I֟PΓ]~�}�B����~]`�mB;w�aQ� u�h�'���'^�U��;�����EL�pm��'�2}d����M�.OR�Ĳ<����?A��-���n᚝#�4b$�x%	у���U�ia��'�2�'��	']�p���~��Ɛ�sg�L�S'�I�4�	�i�zu�w�i�B[�H����8�ɑ)Z�Iu��<`	�!�`��F^��+@���AG�&�'T�X�ȳ,
����O�D���%��(Ggr�I����'r&��Ћ�u}b�'�"�'�RQ��'��'7��2pڬQ9�Q"�lջQ�3>��^�����=�M����?1���zP_����ZM(p �!�Xs��	�:7�O�dœ`��>� �S5G���Qd!�F	D(XGMS�P�(7M+)��ioZȟp�	��H�S�����<��'^Nk��J�-��?��(҅�yB�'��N���?�ॏ&p���ш�	U�!�kC�L���'9��'�а��>�)O��D���#��O�r48����
�S�6�Oj�Kbr��S�T�'���'k��Y2ɑ�-{��A����囕T�&�'S@IW��>	)Od�Ĩ<��{`�D�q���Y��R�V!�@Y���T}�K��yB�'.��'�2�'E�I���e`(0��˶@�#X d��۷��$�<�����O�$�O��e�X+yH��!_�^ä��SHL��������Iӟ��Iiy��B�,�5
,Zp�N-lHaR���
�Z7��<i����O����O�t�2OkV�>5Xf`�?K�&8C@�&/��V�'���'��U�t��˟�����Ok,�	��]Z�N�It���b���)��6�'��	՟H��؟t��+g�@�O�%k4���s���p�kƕ!2���"�i�b�'o�ɉQ�����D�O��ӴL~�ċ��ڥC���@�lP4p�'���'ҁ��y"�|�џ6�+vn�@��)z׌Sl���
 �i��'�h޴�?a��?���|��i�UP�#�������?=�T`�t�r�$�Ol�Yb7O\���y��	B��X�8ք�Qz� a�
6E��Ĉ?d�6M�OV�d�O���SS}R�`xgAʟ?��X�$n(l����/�M['�<�K>��t�'6�TRU�B�X�0�J��R�w�r-���n���D�O�������'��	���������`׭	S����N���QnZ�'���ٟ��i�O����O�q��7�ы���4N�]�AȦ��	�Ʋ���O
ʓ�?i)O���8���N_N��˃-A�w�}E�iI���y��'���'��'(剗&�@p�ݩojfxaf�I8��-PP���Ī<Q�����O��d�O���*§xnD�gh��0!��NY��D�O"���OF���OV�@Ԅ��d4���&�E /�6L��:.^�+7�xb�'e�'_r�'�.���'�d��sĖ�Q�`�9W(߂ h$8��>)���?�����)���'>���n��(	�6rT� K"�8�Mk�����?a�B*A�>9�脍$�+ �.2D�j�a��ʟt�'vLA��&���O��醍V~Z�i�m��b��Ÿvn�\&����˟���˟�&���'op������\�Ҝq����ml�PyB)�C�6��F���'��K/?1�ŝ6P�*jǖW���;Aj ٦��Iʟh¤��$���}��&�`�@A�ã�io� 4Cͦ�fꒄ�M{���?1��R�x2�'��<����J{�i��3l���2�M;��<yM>i*�V˓�?�p��,�rdr�CE�R�u:�#yٛ��'��'��	k�@;����l�"���Ŋ�0x�h!�F����>	֫|��?Q���?�2�Ɍ�V�G�`N��r�b����'�����)��O��$%����0� K1b	�e!�c�Q��\�q]��xdŏq�IƟ��	����'�b}�c��%0$q��c;�(�pcZ=?N�b�@��W���D��ǀ Vl�p!ȑ��R)�t�fuSQ+P�<!(OX�$�O������M��|�S�T' `�'MΞ	�7�TB}"�'B�|2�'�H��yB�s�0s�L��E�}�b��;0	�OH���O��d�<ѥ�נ[\�O�\�b����3�-	$	R<Z*`�"�$#�$�O �$Q�Aټ�d!}�՛=۠�3�36�9�D��M����?q.Od����^�۟(�ӟ=����A[��Yk�(+z��J<����?���^���'k�	T�hz� �4+�:�}��Kh�]����̓��MK�V?Y���?���OD�)G�@�	��v<�~�K��?��`�������OӪ�#�[�$�ҷ)�#M\rEi�4g�pu�i���'S��O�:O���=���ƁV�cL�-�
֤jŴ�l�˴��I�Ė��*��_�$�4y�dl=3�"F<M���l����	��d�c�����h���'���U�pH���f�.e���s��U��Oxa��d�O���O����G���0%��d#� R��A}��A�(k�	zy��'{�'?j��4��`b�IՁ�>`�
9pű>	�/q���'�2�'��X�#�_�	��X�e�0P�2�;����.���C�O����Ot���Of��
�Ƿh��u��IH7H����ri	 +$@'����ԟ��	��p��6���I�h�J�""E�+v�"XD����h	aڴ����O�O\���Oe���,ڛ�˯S��|ru�W%lKls׬(����On���OB���O�P����O����Ov�zSf�ɀ�ֱF�pY�M���d�Iڟ���.B-�!G �$��I*�,�7eP�>�bu���ԛ�'��W��c�Ϟ����O$���f��'��~����!�%7۪Uz�����?qRl�"��'��\c���!�`Ͳx���S���F�ZQ�ie��'������'�'�b�O��i��2��
l��!"C����/yӄ���O��z7�C�<1O�����M+f�d(��A�ibr����'�R�'5"�Oo��4��n�\Q�!G-{Ŵ���Ɉ1l��6�F�8�S�������r%A\8�J�ʅ�'�0�r�V��M���?��"K��Je���Or�I,��$��	 J8p _(oc���+0��ݟ���ӟ��ȇ�u�$�˱f�'�¤�C�_1�M��Y��h1S�xr�'�R�|Zc��)�#�0a�mqP��l�F] �O
�R���O����O&�)M��r )�#+�D�p rr�	�I({��'?�'��'>�'��80����Q� r�k��0ܐK����'N��'�R�'��H*D��	�� c2U�E%Ǜq�2]z�h�(���'�"�'��'�2�'4��:�O�E�`鏭b٢����/>;�P��:��K)u�N� cn��<��e�g�+���4+v�W4ct��thR�7��C"O��b�[8jJ�p��d�
]
��O�@c���@X� ��hiw, �Ӭ�>2Rh�D�p�n��E '�X��;f�I2O;m��P�c�0Dn ���9i��@2��85O>�"'�%*@�s�I!Y�t032f�&h"���b�H�(l�5�G�-c	��ˍ �����RDĀ4��%� |B(���ų(�HC��'sR�'��H �c�2SȔ��;P�N}�ǝ@J����nQ=���S����'���gMT{NTW��I�@D3�A�O�d�ж��)GJ$�S��?)�L�6��6�s9�wfћr���G������ڴb����"|��WL��4��o����s�@��̇��5.v�iW/ƅr��pA��1#<���i>]�ɀ{;ލ`4�V4
�(�!�,Db:a��ٟl2P�XY7B$�	ʟ����!YwX��'u(�f��a�1��)[�% �	+�a�O�ܹ�G��]�~�1�Ө����$��*ot��S*0ehep����Н�?yq!��l��@�����3ړUN�ҍ��JC�Q�����D��|�m�d���˟�F{�[�t���M#�Z2,!��q���%D�4p�Ԍ8"��uf:~ԝB�	���HO��Ny�\7mD	��KabN�5���2���ef���O����Oh���@�O:��d>�K���6)-���?2T�A��G"}4�цL�@��t����Dx����k܁w�Z�2
54��Ё7�C%e�p|�!�AZHj�"PO�Dx�`�!��O���Y\6��@�.~��m B���-:(�=���3U24����0f����^�;!�$̧v��sw"H�t(��Lƚ;��@}�Y�lB�
���O
ʧ1�ม ۟d��k��άGc$@fN�?����?�4�9U��a@��^�.�����i��L4�X�̇�R��4�4�˙�(O ��#�t��+f�,4�' 9&:Ţ#��R�`=ză�3Xt�Ѣ�(O�,#�'����Ł+��hl^*'n�ԲC���I���Q���
3a�_d�C �Ⱥ\�6�3p
=�O(%� ���Q)Z��U�WK�zt���y�P@�J�����O�˧:�da)���?��^���դ��,kv|�"�>j$U�`�4k"ع�`õ��E���	+��O���k�b�NL�A"܇!��4��	�TZ�I
l�yQ��
@�:@�Pl%���q���I8�=���¦KK�۲��x����Iߟ���'��h�V�	�hJ�|h��@lH�2|x��S�? �4b�%\J�Hd!ߟ~���I�ቭ�HO�8�t���˛�u�l(�F�%T^v���2��¥d�>�	�� ���<�Zw���'��H�5�P�@�􁰍=g+.�R�'֜�k6fZj�R�o;O։�q��^d<�ӔcQ"���%�OXI�p���(x�Yv8��H���emܟ>gJ��E�����=g�r�'TўH�'B�h���M�'�F�;BA)�nu��'�d�2T�%;|ΰ��L�� gX"f�)�S�TV��{"	��MSu�Rи�"����p�P���?���?���b��Px��?��O�`�bu�i�B�A7?�Tk��L����F�L/�p>y�!W��dΰ@��)���פ_ݳ���%A�|b�
'�?9$�i�:H5!�yC�l�2��6������s�"��<	�������'u|���b+�IQZ��
�!���;n�a��)>~1*�0 �̕1Z���I}�Q� ɂB�M����?1*�X���;� �F�K(8X`�J4+8���Oz�DCPOZ�ڒ?�|���-r�n�����
?iRe���Yb�'�F�c�E��h��500�*H.��Kbb�6�������:��J��b�4�?�*�:L�ӎ�6(�!��a-�]H���O �"~Γt-�tåw0eXg*�D�,��	���X�s�����l�i7%�R�� ��+!�i���'	�%xNʀ�	��͓O�f )0&�>���`�L@�Dy�.)�6m?�|Fx�,B�L���sg)�� %���I'yϤԳG�2�)�矼�D�ta��eM�#����B-«_C�Y�	ǟ�*���'���6jͲ��4k��E�8a�౟'���'� � �h �x*b*va���Q�����:~PD���ڂx�(��ߕ>����O:Iɂ�
4B��$�O����O,�;�?!�!��P1��̨G���"a�I.G>P��� 	��e �T����sdU�P���z�(((� Y��FJ�#a�����?𾤁�R F��h�'�*�B�$˚xq����O��ԟ�	�<�'�:MGJ�g��A ���
�����';�y��<��A�I�4��B#�瀅	���dͤXf������Pu#��?��i8��4ܚ����?����?I�b�-�?A�����4I6ܻ��i�м@���cm<�p�UR�����vO�=�횫�M��B$oj�	1���MnVU���{8��QU��O`�lڷg.�F+��QḆ�a`���� �4�?1(OL�� �)��M�M�@es���x8X+��j�<I�	���Q��Ȕ"�Bآ��<A�Q��'`�A"Oc�R���O2�'j[�$j� �5���@���`z��!�V��?1���?����z����D���ݮu�І�<_�S�\����@ 6����>zv:�<��^͢#��$���gQ6f�(i�O��di5`�� �#wY�@����$��Qs�%m�T	n͟�OL�0JAdΜt�� �3M�,	��'i�O?��i��)��aI�Z*���E%'cP���O�I�sf�LX���(-�4���E�=�2�I:�D��RN���L��H��4!���t�I����1a���R�����f�&ų�B�"F��(�)�3Z1�hQ��&:��i+���0т��5�rxy㕙%��4<���s��uVz�����2=,L۰/�<-����EE�*�*���)!J,wި���:e1l)�猒A��qDx���'�j�s�G�qu�cI�)��%s�'05	�$6I�áN+��b����F�����'�l�6fF��`�v�BG^0��'BrO�cO a"��'�2�'��"l����� c��׎����]�=i�,:S㥟��O=�Zx���&�ȓפ� wV�t.�OA���/?X���n|؞X�6Wt�3�O�Ƅ ��V���$�=3�t�'�r^�x��I�LZ8�)�*�~\��%�+D����J�0X�4y�IX7Ű�H�Ȓ�HOT�'�򄝆+Yx}o�%N����9y�e0"��V��<�	���Ip�����I�|" aU<B���4le�)��CւW���
�Q*t`����*}���0
����5���v���Q� U*�:�OP���'
n7m�B��`�Qhӳ1�J\9UF=cƵmߟ<�':��?��Њ��>���dF��ER�JbO$D��94�i�H��!Ϛ,#����a��j�O�˓����R���	}���H�!�y������A�$�jb�'#��'��˳���7�b��?0���T>mhq�!��a(WQ�`�e�=�x� �iX��(�7+L�3atX��c���離&`v��3�W��2M���H��Q�8Ѐ,�O��m���O�`t���>e��T�K!vl���'��'��a����g+��AD�N�qz���-���� ځȓ%�7M��u�$���}118O�m��o���	��O#6eH��'���'�<tr��>FD�A�+@_��#�	�w���y�b�b�0�ņ֐�������Ͽr#Ͽ'5!�EEn�%��M?]����iDW��� �Q��������X0q��4�Ͽ+�S>���ںx�(Z��D�2���s���?Y�O�$��O��ð�F2h�`����Eh��9O|�$(�O�Ұ@�0.�W�H8&�	��HO˧}.My򧜓vJ�@��D\	dtR��?�GI�&�*���?y��?�Ĵ��d�O�|h�,	e!<Mz���?yl�3��O��O_�$�,�@�'|:1���K hKU�AjW�}X�x�'܈*!n�B�hR	��:���$$̥ ��@F�REZ��H:��I��~��Y�L�	by^#z��=c!�c;(�b& /�y�iR�+P�l`��-]4���6���3`�"=),���O�N̲���ã��2�ЊU�W�u!�$,�JaY�D�/��Y�ċ�'��Ј�ݭz����@�L>�	�'r�ՠ�d�'�$Cv�,HX����'9�[��ۻ7tҴ��A¦�r�'t�R�Gٿ'�����ɪ��L��'�HL�#��X�R�8c�_yZT%"�'��,豧L�p�4$S�b@z��#�'˪��u���!�s3.@�EM�9�'@ͻ�Cǃ{�j�s�W��HE��'�2�h�*z��r��	_��i"�'y�*Ǭq+��
��^z"I�'eL4ä�yy�L�ыТV�����'$�4(%�L2�)�F��i;�'@ް�g!H�~'
��9<6���'ʰP)�$���,�'��/�Ƹ��'ib�ˡO��v\ 7���/Ɗ���'f�=5jSpK
���V#��L��'���X�+$$ykF�0��d��':F�ir�S�$�H(%�ʏ�de�
�'���a N�:7�����"� R��
�'�<p��IŜp���;�
��B�ډ
�'}�P`Q�1����'� 8��	�'��pz�OYP��7��,ZN %��'��b�U>5�6�E�Pr}c�'T�!贩��@H��3V��Nш�'�b)��V��E� Jb��'��P�Ǎ�@���a�ȭy�p���'��:lˊ&�(	�1k@
�,R�'�YeZ�Q>�A�ں�H!��'�Be����LA$�À��qO��h�'sL��CC�+)v�0�>
yR�'R����L�;H��w�3/����'�֝!��۲U�4���oOK��*�'쌡��a$k9�D�1���K��	�'g�u�e�1o�=
6���mR\$v�C����*�� �"�E�@�6�~*4o�$W��ݛ-ʺ�b6�E3u�T=��Cɯ�B�ɻmJ:������h[�Aa��	�wi�ۯx��ic�X�r��E�G�p�
��b�"l���D>_T�6`�%g��b4g BKax"�ʔaˬ88b`�y�`YD.�a�|Q���A*
hʜ�EH1}<�A�5Y����܉>��{B˾;6MJIH45�ҝ˕i����(꺄x'�N xA��lߖ	��B�392,�������rR@<�"咱��;��  �"O�!�!�1+�yr+�:NiQ� �*f�BZ�n��c?�mࣰi�$XG(Sj��g=A/���wl�B"�/Sv\A	U� 5�TA
�'�l�@E��58L�����-���6H�(�?�A@�('ΘӴ��-ԭ����\���u�d�+d�y:s�S&%�p!`���Maxr�é[U��S�3?���k��*v�����oK5l6$�!DI�X�$�y"�ܭyu�u��nSZ��{���5�f$1�GPT����4��(��䟀@h*�eQ-5��pA��®`��)H"I�2��A.�"mԍR�%@����I�����*�"O �1JL�����Ɋp���x��|cD�i��A�{�(A���3&!�5B�|�&�P�޹λj.�b����*���c�5+�����x��R�^{�X{����+lCD���ڿ��GT
�݃GK]9x(��S�ӎ9��d�$��<<Ĥ��x�:�D]����K\
=p� "��T� -�n��F��:oTɻv)���O����N)4꬀�J��W���ԫ��^�KQĝF��Tp�&�
k��h�Q��P�@�k�@�O2������Z����~ʟ�y�f!'@���jM�L��r&���;�"�>kX�� �@NO�e�� ��%����FNd$�ӭi�bZF��M:N��GB�W�^ݘ�'ց%�X�ڠ딿8���s�D�R�עE��=K����<z��dI$JU�,Y2#ƃT�.� �Q��c�|ҖO?}����u�uI�
8V���`G �y2�KD���
OfpF}� ��Xb`��I>'�2F�\�B$���M��!��\TQ2b���R�J��>ͧ!�-���i�|`#4��(ZPi��6y�0Q#�V�'��i��M�6=�`��b�k�@pg��S7
�(���Z�\��"<i����lá�O�)̧ �esn�>@���3���<6`�	p��J����9��U�`۵"�����0�%��8��O6����G�4�����d�� q�'�I1�J��$	�[��b�D�����g>}r'����G�V�
	�U:#�¡i��+1���b�}Z�O���B(��y���) ����R��O4 �6c�+�ܼ FCO��O���j��?V !{�J��zY�i顉��
��Su���'V�:T[��i�N����@��>�[#-Κu���p��H�'��)�ÞuR�[�񧿫THW�t^��筙^����e�'p
�ϓF����s�Ox`�I�!��Бd��w��鷧�|�p���n� ��$y��r���"� 3��|}���=y��%�T��H�(�NY
$j�YIz�IH����'����2O�*ap E�2',I���vh_ g:����_�Xd� V:/�批N���&�p��/-�l��׼\o���RCYZfe�+�p̉q�H9k�0e��m&O�-@�h��(�ޜ�E��S!*���"$�ى��ݩT�	F�O� 5��fp��:sBϪgޱ�P�R����fb��s��~�;}R(�q	�ML��jǚh+P0L<!/ĮuQ�D[+>�g?Y���i�|�jφ�\<��#H7;�l Yp�YH�:�ꑄ]����cآ+LB��cK�
U�F|cq�	(8XQP������5?���I<Q����/�n9�JJ��'[�5�͂9#���%�����J����C�+t�@T��m�>�X2�h4�	>GSv�#�i��3hjhF��X�l�B�:���6 �,1�!�'�����#�����D�yشS���p���3!�}І��o�P,���<�$.�	YWʤ���G�
L�z�R>
b"B�I�D����ɝ�$,�d#�G^�m��I "H ��?��'��$�K��5U��;�*��I���\'ga}��ۙ��ᣢBO�pW�h{%H�/J�T��b�y�������:a�u��B�0yޔy���5}���P^��"�vqx�j�K��hO�%@c$�7E㰄��M< Z�Ђ�O8�(	/b�e�+i�t�8����p�1�)֐I�ƽ��A�hX��y��*9b@d�2�J4*��M/?ɰm��N�hUr���uO��C!Oh�T>�Y�f�K9l5j�Nɣl��Cc,D���eY"���#��,L��|�p�V�hٖ�#v��+x�x�䧘Oش���Nͼ��	]Ė,r��Yn�����[J�<&�(%V���+�"0��NN!�P�-O����@�y�1�1O&E� `L%|�F���A�r�
��mR�M��U�CdD+���"#�_?M���,h���sL�1<�^|"�)[b\Hˆ�~G$��	S"�j���"2�\����H5E*a�5-��V��, ��9�U�T�"�&����,Ox�	���	UW\�x'Q�#�kS�'	�\e�H�J<��W#Z�RZ��p`��=��a`�G����'��A 47O�t)��;J����&����W�'픰��G�e��z��,Ą������p��(c���PK<���$F�m���~��s�%$@�L��E��<%���G�A @h�4|�D8��J�?>���E{��2LHl	���L
��� A�i��!"G�մ��� �
x�e��'�Hm���+�����O������0�1h1�׫c;�h��+��&�,�/�OJ�C�A�xn��W�3>��s �T����:l�d��C8�ɭ|
��qp睫R�`�7O�
𼋵f��:���M�u�4 P�D�Dҩ[�Bڧ:��a{���:|
�y� +��a��H�Po�,϶0Y�G�/�d�7�Q̱;�(�"_AL�Y‏8?@�"<��2|'��#�@�A���0���<��*��&oT4�L�g�;V�|X�L�O�=Hs�'x�ћ�읪܀�a�dJ�HN��2(2�l�iA�H�D˦����)2 ����̎�I�4O��6 Hsl�kE�O'!�u!� X���)d;�aے'�;_�R@Zj���@��'�"#�<�P:��˺
K�����yr��g3���0����~bLI~�����`�0� D�Q%�|��s',?�O���2��9eqP:�d�	j6�Q6A1�^���T'�&����O������^���DQT&���ˆ8�����j܎Q�<eK�(Z>{s�D�cg�/u ��	��ĚY+xȒ`a���O�-B�-	y�Dri�:a��8��E�O�m��� :.YIʷ,�|�#�V�V��%�$��J�@��3�e�+�� ��JY+2�4	���<�R��X��%��ZQ?�4GV%� ��Ӏx�Ĉ�9elAq`hELBX�;4�'X�W�t�'dA��,T�:�F$�vɏ
�<��I��y2jU0)��x���ہ�~�_}�'��@p �M=�4�K�)B�Z����$G�y�! &\J��"�&À D<�C�#v�������Y�pE�y��Y�p����'�(q Dξ?a��G��N�T�áU*\��=b�Aѳ1���R8@��P H�P��;D���cr ڱ%E��!RZƊ����Ǿpx����A:�"���ٙ�h�i�/_L�����<�vL�xJPQ@�F��e�@D�4#�-GT삣%$�tHZ�T���ي�9�
���_�d�'�X�^����x�H�������: �
�?� ��3~BX�a�V�Z�v�a�B_��X8�/��X6l��!e��]�*�ϧ�?�O3|tcKP��a�׆�p|��X�N��*d��a��>��y�F��j��ҝw%�9��%6s�CBگNN�S���\�Ra1�'������d;-��q%4w�A��dƘ� ܪv-ш=bt%���O@��0���<A�Q�J�Q���H 
�|�B�.C(�(�v`�2��5X�� ���p ʛ.�6(�$N�EɈF��P���` �B5��Qc']/�H{A��y��(P��<u��T� ��W.�}��'ʔ��0�ԃ�#��8E(Z1�LY�M#H<z�I�8uz���NJџ c�&�o��XFN̙F�д�Vi�0��f[�%dĝk�I�(K��]z?�O+$s��T�dvn��΄;i����s��;gl�Ke�!jn�xB�ߩ��&e�咀EL�Q.��G��_����(^I�����O��P��� qbi���W�,p����/�i��X��k�Qq��P��;ѱO4U�%�^��
}`��B��Fă�J3��J�5����m��)�B�ծ�4m���Z'���OR6�ؖ&��*Hъ�<Q4䆣3����U�n�9�� �2�n98��	@ZD�2ȏ^��,E��O �Ka'S�%���j�	ְP�À
R�T�2dY��[�6`	�G�L( �?��d��`H���9���s���#/͖	����j̰0����G��<���~��$�p���MzI�T/K$	T��{��]%9i>��C�l4q��爠2�k �(VK@��b�4Iq����B���n�H�G�/p��'ڌ�"�?�� ��9'���Ks�!+^@��t*�AȱO<�@d�?o��xg'ܫ�yu�#�T޶%���5,�`���A��e�lY&��4���D��	�*Cr,��Ot�I'�$�B��-���f$�dgr%rIX�k�z� Ti�:.�r=Br&'�U?���йV�ՙp���ӣ�$����+^����1<<�FR;`k���dI�F��9rV"��oy��Iǀ�9��uh���#�rI�O�0����Ӻ�I	��H�� 1���A(T�D��2ʝ@�UX��U�b���$@�.���3Q�I)@�x���/,y�����6}���I����#��d��'̴��\"E��秘O0������e�k���4<�ڕ�jCV�6%|����%F�� ���Ȕ2R�EhK?ٛ�j�H-���d��3�p9�㗝)/��'��"v��|����V�t{J>au���:�0���WA	 1Xq�,w:��B9�l�S �U����|��O�T��&x!C���lb�x e�?%T��e�4؎�"��' �&�����sU���h5A�#Fxv��g��b�e��� �O�T� n��	��DpMJ�qt��D�
(��-�B�4��f
)��%�:Y�L�*!1�ё�S�6C�������I>��4H�
�?��>���&,�E����#�"�^`I�k��4:~c��X�!��@H@3lZ�0�Iy�-�N��{���1�� )f�EB�(�M���D<�s�@���	���'ڞ��կ� *�dApH�>f���噎}:��C@��eK����ԟd��D�%8����Ї9v��A�
��ɧ~��ʵk�l8������O�TI�p��|q��M�_��� D��H�����<����]}"��=� Y��ɄSw$�3�w��̇�ɉ{���������%kL�;oNV�Tx��
��~Bϑ8�r�'�.�S�s�((����U����S�ǎI�Tj�F9D��+���<Gi�Ea"ǐ�hC�@9'�$D��2����#s�! ����֭"D��J�a _Vn8
'���;�Z�3�H!D�D��́� [�hB�G�&�PTzfI)D����� �|��aÓO�$y���3�H3D�D���W=}��ء�*�m���{�!6D�8H�*�dT�I�B�� d���5D�$���f �i�1�6>"U��B3D��zb-���G$ֽk5D����=D�\1DB�7A��0���֨k��S��8D���p!M %f0%�U!p�$+�+6D�� eD�i���sl"^,
yP�.D��29HB8X�h��
���q��*D�\a�Ȟ�~�"�����L��f�>D��Ö,��h|��b��R������;D�0Ic�Ǖ�@JD�Ҹ\�<����'D�T�2>�Z��+�d�"�ԋ'D�0��@��>�X�!�3 T%P�%D�h�ĕ� �� �eM�[oм�G�=D�`��0h�4��A
2粄J�A;D�� FU&�QZ�\��eɋtW��"�"O�Y���X�y�*ɒ�FҰ�q�T"O|���![�=����6E>~� ""OlD9"E�|8�+�#�p��Փ�"OΡ� ڙH��%�爖3
���#"O���n�*U�ąsM��y���"O�L�uK��.��-�j�d��R�"O�$�n��	�H�l�4�"O��K5n�T����kP���<�"O<�iU*$&��!���F�y.d��c"Ob|S5�������ؠ/#Rl�t"O*!TE�)+}bl� �x��c"O�`��F]�f��c�O�Mt�t��"O�H8qaB�xG �a�?!tl��5"O�tg�	Cl��Q���2Uz�"OZa��!�L��@�ћW�r��d"O$�bs� �����vyZ$�"O4��B�I

��:�EC5�u0d"O���5͜�k.p{�B�[���"OFIٶ�]�V&J�2Q�ֻ�(@h "O�-�@�0��բ�8��#C"O�9�(Dp�
�ip��4YmʀY�"O��h7�u��Ta��ݐ;g�qV"O
��'˪P�$8���Ī&`�� "OX���c�\�~U�	ԥk�ȡ�"O�Xhh���P��ʵ
�t���"O2	��d@�,��BP�I�;� *�"O�Р��̆ � ��c�3/((�T"O�h ��;7~���K�8:�0V"O(,���)#n<����u�'"O�1��A#N����KJ���4"O8�e熞�܉��n�<E���s"O&,"���]N@C���ВE��"O�X$M�?H$���:�3%"O�@��.�Tj��_�J��q��"O�\��A�A�Z�'h��p�d"O0j�	�#+��f(v���K�"O~���mD�\���SA'p�h��V"O�8��-��4�����F�	� с"Op�p� �\ �h``U{n"`�U"OB��ɦs�.TC�ɂ�V����"O���I:rqV�Z`�T�87��ҕ"O.�ɑ��~Ѫq�I,$��%"O�H��H:�| �kP�v^p�"O���Zd�و��t!���E"Ol�s���9
9~h���+i�T�S"O����˖����q�D�U�b�q"O��[pG�7��}���[����"O�E��׶..0�$�D�X���"O����A@Z����4 X�ӊ T�@ ��G�����F��	:f��psB(D�Ȃb�_�U(����`,�*��2D��a�BÄ)�V�b/��ee^]��%D���� U?x����ԍm� �*O�����.]���QR(#�^l��"O�xy4N�B~��!0���x'"O}�ra�e4���`��xV�,�Q"ObIZ��s��t�X�j���@q"OJ�1��F�����ԥiyN��Q"O��Zc�lC���hH�DL�D"O�p꓈�50y�Vǔ�:��s�"O6��3�&TJv��� �"O�q�d��;M�0ՙ�$B+7&|�(�"O�Z�`�?P�B�b �?��� "O� v=������>���� ���{�"O6ȸ� L*�f�Jw-'��@�"O歐�iP;2�h'�:^R��"O4,�!N�mQv�ad�<�X�"O.x�� ,�6�D#��@"O������b����[�.�:�h�"O Pa�Щv<�h�A�;���"O��4�6�`a�����e2b"O��� #�%NuxXYe㐨��la�"O䩢b�]b-\��wO݂D$�Q��"O�p`��J���H��I6L�3�	y��$x�2�y6���W�Y�f9$���0���{�D ��T{�ڶJM�y�E�6����(�
Gֆ�MC-�y�";���I܏M��L�%��6�y�$�=|v%�1BʟKT�`%�G"��',ўb>mcB��j��8BUm(W���� D� � G*��0�K��4���F D�tˣk֭"�����o�gȔ<pwL?D�H��
j���z��|fpRР!D� Q�IB���0����y{8 ��=D��(�b���I@$�Qur�#&<�Ir���'zA"�ᗄ�
�\�3���f��\��y��0g��Q�`��F��i\ ��y	*h;qG�<d�e�Pț�@�ȓaƆ��Eϋ�^aV�*P�"l�|��s��M�gg6NeP�����Nu�i��~�whN%L7*A���DsE��������Q�)M�I�t'�<����H���R���`�A��A�������b}���,hjn����Q<h|%��o��y"�ģ������
�x�B�@���'���ډ�����s̍�#xr�(��O�oE�iv"Op})V &�cr* 6���z�b8�S��y"��_���C��Y��#I�&�yr	��0�\M�%�Ʋ���IB���yb�[h����JJ7#\ɒȏ��?1�'4�ږGC�Y�ސ� o5N�>x�'�Z�Js@�;�b��WkT 7�Z	��'��%2$�\. �廣iJ-EGN\�	�'M�Ab�Eڸ�P0��ʦG�T�q
�'2M2҉�&$Bp���6:C�4��'�(���OG
� QʤE�4��,��'p��&�(Mj~Bs�-,:�T1�'��5��WDm�x�'�S?+���"�'ԑrDJ/ ����V�Ȏxc�;�'٬���-!�v�*���0C���
�'��-�Vn)/��h�E/.}N���'��1Rh[%P�^\�`� =4P����yb�D�K�|�	D���w�8�S�b[���'��{rFڐ�d�,��i�ZQ�@
,�y�H*�D�AJIgY�]���� �y�F�"+�]�fc��Q��ŀ��g�<�͊��0:�X=D��̈b�N�<��&U�L���dƼ�U��h�p�<i�i�&"�����V�{^&�ZG�p�<)f�5m �*���}���[�%h�<�p��p����7Cn��@n@Z�<�a�M���,�} ���4MZn�<Q$�ĜNc@���� `��A�f�<a�V�{�+b�N�fX��A��a�<��/]�N@|Zү12N(�Dn�^�<���F�'L)��Ӱ|[�����@W�<�RX������Y0B��M�dh�i�<� ~�e
�(�:a��Y�}D����"O|�5k�� �\��H��U�}S�"O(h���.�4��F��6պu�"OT0ÔZ�	�@�+�l�l� �"O�x����;n]T�8W��8h���'"O�Qr�@�]&x�P�;� �`"O��:��[����[�I��k��`�"O���E�4��Ti���S��E�"O�x���#_ےu#5oQ�4���"Ox9Ʌ�Mb�����JM$��2�����ɫc�:�����iŤ��3�ED����-��ñ��Q#_��b8�W+B�<L!�$K�j� k�^�(?��PCː
w!�dI^JraQP!�"U& \[ظ~]B�ɻ>,$� �
;��� �'g��C䉛)��is��	 ��Ur$�M.@�C䉴;)�]�A�0)H֩��aF3+!�C�ɓ M��)>^X3�k��9��C�:>h��Ơ�9! 4�"�o�bo�C�	�:�m	X� ��r���`ש#D�Dq�i��ʌ�tO�[l�"�e7D��SS�Kf�ɻ��
+Zb��Ӄi!D�w�:B���S�1Vn��a=D�T��^;a1�e�r'Q2}q�҈&D�`��k�>X�40�a ЄRR:���%D�|�բĔ��i2P���E������/⓷蟊08�JP?EЅ�s�RqF"O����?F�̑Q�I��.�ɶ"O����o��dH����-Z�"O\���ו: Z���@�hձ�"O�h�F�O�c/&d(��t{[���'H�k@
45�D���!�-�H�[
�'V�=S!�>3)�aRuc#T�I��'�.�Y6�$|��X�sJ���i�'Q����*O�.I�����Gh8�'�\�pd/�:8�2��# :�{�';����x�,8YU��Hy0��O�eҲ� V �Yu�L�Q.��"�:\O���SkW�>��K�	վH!B(1"OJ�ZVD[ .�"e�c#ƥ"4|I6"OD�k�nA�.L��hEn�F*OF¢n�,*����M�|�pp0L>����߹a4�R���Dv�@�f�Tf!�D�	��H�ªN"yp�؃I@�"g!�D��-Dx"f�/+�ndـ�<\!��$���]�{�hp���vG!�DC4�A���	{�*��'>6�!��!j�=c�\�f�>]yCa"~�!���H=�ɘ6���"��i�%R�A�!�� RF(�r��<JP�8���h�!���>G�.�i�M^��S���^.!�D��p��Y�����V$�#J�6
!�L�_�0m����y�����&^�!�$�+�`)�A�6m�A��
	�!��L;$�d���I�W��j7� !�D/��m�G��E���<!�$�#4b��H� n�L�N�/.!�D�(v��1*�%$X�a١�R%+p!�D;r��� ��A�c��	��Q�fY!�dP� ^�8��L"R�� ��� pT!�):�m#�F%nǾD���ɑBT!�$%ր�%�Ѕ.6DI�o��V�!�D, �L A!ď8��A�7^�!򤉶_7^�J�ɣ$�Db��7!�� T��C��<I�L�Fo]S0hܐw"O>@;��Q��έ��˴,�-q1"O@hs���|�����%�=@洼q3"O�X ��� ��#����\�)�"O�[��[�"V���
��e��"ON�HU�Y)��THЅ���V��"O�@���6&��:�D����"O�� Đ ���kC�;5<��e"O�ěe��L��A�k�5>� "O�Ƀ��V6(Y�p2� �~0Z�"O�CH��ڹ[���5��A�"O��a��0yy��2��%�d\�"O�5@TlV�MJ	�4�
����"Ol0Y�`˥|{zL���4e��;2"O6�UA@$p���V.Y1O���"OF��2ɘ7,nPl�<3���"Oҙ��J߻цS��J�'}��"O�2�s��1'I�c9��"Op�A�QA+��%ܞ!L>��"Op������I������`�V�y�"O�� �!"M^��R'UɊ�P�"O�	+�U
*�I����![%���G"O
����"VD��Z1Nȿ|�T��"O���p�C& Ѣ!z�m_bl��"O z6-��> ��B�R
)8@��"O8hQU�޹f���;Ao!Q ��0'"O��gk�$w9�-+B�D�欥�G"O,IX��<�h����N�r0"O��#G"ԧ��Űb�T;޸��"O؍��cFj$�ъ��I�ꀓ�"O\A����3S�f����ơ)����"Ox,�UiX � ��֮-%l��"Or���O.���*U¶Em�"O�9H�F�h9F�c P�H�FxY�"O$M� ��	��ur�@���c�"O�0��'źP*�8���8E�,2"O�$�4�̒A�jD[�@������r"O�ر��}n��2E ԍA����"O�}�ޒWe���& V>0��S�"O����K�faT	�j~,���"O`�ĥY�X� ����-OO��"O�h��+R��ft���t�B��"O�u���{��@�7���~���A�"O�l0�ˎ5�Qa@�1jg���b"O� �� �!Զ�S0��)X^=Õ"OvyꉐG.����A.T`�E"O%�q!,K]>���C@�w�.�W"O<P��$�m���Ӣ�U�x�d"O������hb���z�X��"O
!3�'Bh� H�(��a�"O�`�ѕhv�Q ��Z�d��X�"O�X!���`���(�D�#[w��R�"O"�@�.��ݶ��ʺys0�:�"O2Y��#ح�bPyg�D���d��"O��	"��dy0���	~�C"O��Q�q����d�E??p���P"O��#��%gP�<�!"ڸV��!�"O<`#&M�Y*Z�X�+���ԑї"Oج�7�3���ь˖k\�!�"O�!��п[沈)��H8v��"O�d�T��JԸ-h-kaB�[ P;!���ge��Xu��9�8P#ÖE!�D��qpv���\=O�����"�P�!�]��:ġR,o�ĠT�#�!�� �@�`ڬ|'�$Ё��I�n���"O����ޘM!
��0L�>z�Fؙ!"O��g�� '�T�DB�
�
h��"O@���I�O;T��i!Kk��""O�����B�cȄ��Ađ���"O��� ���|���@�.4���"O:�zE̜#�*l�S�F|���"O��	tiO:%�p�cn:�d(�"Ob�����D��U�$AF�b"O��rӌ�b�h���,^mZ�\��"O�`r�63��U��63> ��2"OT��r}3jq�j\�i���c"O�ixtNG���J�Iɣ'��I�f"O�=�F�9_�(1Ί1rz�+�"O�Ѩw�ǩ2Ϣ��NA
0��@g"O�5�3�w�����G����"Oȝː`�|�hĊs��ܘt8"O&uA�%f��x�NJ/RqĬ��"O�\�sMÃ�dB%΋�m���"O��׬�0%A�l�jpF���"O�sr��lc~X�P� EdN�"O=;I�)/,�����,# �Y*"O�(j��O�l�+���	�'��P ֠B�a��!�gD�k�����'��m����B'�����	jX���'*�$X��V�h{ (�7�8\��	�'BZh�Ǆ�!|�"I����[����'�ʹ��` �!:�`v��M�����'Dh$iԎ�^�^�U� �[ ��`�'�f�
�l̑>��U�T!%d]�X��'�v9�(ͯe��0\��!AF��y2BP�"yY��PBV�L�S%�1�y�[�,�*�g�7P�p�9DD�1�y�E���&�t)�Ӟ��Cd��y�PE5��������� ���y
��Ԙ��i����pUL�y��T�x<�����wRz|ՁӅ�y��	e��肓�]�޶�H��_��yBbT�k�,PK����E"�t#�"*�yҩ�d��l�26~��A���y��K&e����k�>4�V�
�E��y�-�
���B�ɀ�)���a��y�Nڣ��E[�S�q����yr�K��	#�E^�����׋��yR֞$��Ó�"h� K.�ybkR;E$ʉ��	�9SZ4`#`ś��y�l�$,U��1�mȍG�3rO���y��Y�	�4*���;
*������y���$Tl�`�D�06��z�B�6�y�Z�r��c�)6qn��4�K��y���/6b�#���Y���sM�y2���jd|��ςIqf9��)?�yR�WW�	�veQ�*��3!�6�y�i�&c�)a$pEXgʕ;�yR�S�	ɫ2B��7I���,�y�E�"�@�JF�4�uk��y���kR!�*̾ 
,�KӉ݉�yr%%T{z-�r� t9�(do�(�y"���
S25���'؂u������*�3b���j&��thH4�8P��3xYbn[0kv:Ѣ�ojh�T��3�hř�L�t| �AAA�B�d��ȓ�tQ��$)�pk�T5:ҝ�ȓ,�XyS��B�8��5)1���S�? �H[�#��,�m�C�T�(��
$"O��)�N�n��X��âH�|��a"O|UY�#�)=5�̒a-ǡrK��� "O��ZwÆ#OJ9[�␇W�db"OР�׎ِ6�0��s��&U
�"O8��C)ۤ��E�a�턘��"O\���NK\�Nak���ky�,��"O*Bq�{�pȢ��5j�!��"Oꉲ֮�#-t`�XZU���P"O�l�0�N(P���K�D�A;̡�e"O�ahe֞�8��%J�p'����"Oaу�<>vL�Eb����"O`�kM�M�
�̍g$� �p"O�	i��ݙi#qҦDC�u0B�h�"Ofy
�N Hy��F.�ry����"O��@�˛\���a���#:P
�"O��3�^G��\@Q,C/+�r��"O&<��υ|�N8Y�k��T��`"O�d�gD��>z��4쀷A���aQ"O�s6�S�
��AZ�4*CNt��"OF�I�+�.S|D��wD$>�W"O����J�\0#Û�"S�)R�"O��b��Јy�lҪ7��L���2D������e���P1a��C��4X'�1D�A@0.�ɊP��b�r���:D��)�$ҞA��$���6f�+g7D�$���T�CĔP*P�K�_J,0	`4D���Ă��c��P�aD�P�$�8'�6D� ��1S6BT8�N�>D�2`n5D��� �B�W� ���$��hqh.D��{G*��1zc�Ҧ�$��T..D�� �)=T~�xC�N�O$�M0D�d8�$��{9~Bf�t�c�a-D�h��ʛ�w������G�Ҭ���5D�0�W�J�n�$���:��rW>D�D����#8L���# �`�C�D=D��L�-Y�� �Q@!G0*\�r�>D�Ћq�&o=>0��ˎ�)�^`pu	=D� �����LI�KN/h��0c��7D���G�q#~�����{��0W7D��q�Թ=ϼ��D�K%t[� 3�c5D�8�QZ�H�ᣡʛC
�t���'D�����7b����͚�	n��`�%D�Dj�'�VH �
ܝ,p�` �k(D��ڐ��B=�Ex���=Nr���h!T��S��,�v�*���}XN堡"O��r�`��N�Z6MHN�cc"O�hH�(��LQ�F�Q��"O��E	�?���
D�	
/6x$h�"Ot3�+�i2�qK�N�1 (���"O�xɒF����#m��F���G"O()��l"���W�\�U��"O\�W捰�s�*��講�"O$|��ab�<���1���%"O��;r+^~�D�bX1q�v83s"O Y�qo�H��p# ��"O���`*R+c,F$���K+=^a[�"O���f�"M����I,�i��"OP,���W�l)��� �]�xb�jF"O��ҥdʽKX��b�4o���b�"O�ꖅ˷"S�i�0��K���;f"OM*��*1D�#�!J�q*1B�"O�"E�=���c�*�/�iC"O�c� �9���P7bfuy"O� xm�R�ϽN�!��#��e>@u"O��sEьMܤԨR>I(��"O1����0"d'���"O�UqnW�x����6sF\3�"O�Ti'�%L��{C�7c��l1"O�a )D�_m.<pGÇfʹ�1�"OT5�
�	FA(2h�M!�AW"O�8�-Eb��uJ���g!�9�yR (O~(C�_z	�)?A ��Y�pp肎]�d�Ӈ�'�q�ȓHXL�3c �<T��k!��:M����ȓ(���J��t`��  /�Ф�ȓ,�=aƏ��J�q��=�bp�ȓhti0��L9�ڄh`�@NV0��j���8e��&i�������:)�I�ȓQs*$	�i��jn��,�
6nN���9��)��R�*L�q ���1��e��9����2'�H�L�y�`�k0��>��XH��{Vj+U��6�h�ȓ`�`$��_va#gL�<��ȓd��y@BC�XM��r�~���en4����[|�����id��g$<��#�'B�h0A٬ ���ȓZuD)ذCZ�غl�ƥ#Z��ȓ]�1[sDW�jC��)$C�si��ȓHW��n�0��5��-+xE���ȓb�2��Z�6I�󮑪0\⠆ȓ{��=�$ڞ`c���j�%^��0��^Z�jD �j�T�Ɯl���ȓ"�Aiɠpq:��R�%��q�ȓ�������`�T��� &��ȓP*i��/<&��w��$c+8D���FѺ
y��P��F٨���'D����g�%����ϓ�#v%�s)$D� �be �+R"��e�V0^E8�(D��BPC� 	��|�7��\Q� k9D�(;G@�f읻�'X�Gx@]C7�8D�P��7q����&.B>L�t��e*D�����@SHn�a_�N�~Isub#D�
�ǟ+g]l%P2�GL���D"D��e��;*�L|��+�}6K#H D�� ��T6-u�htQ��3�2B�	%3�a�a2[$�X&���j�hB�	���rV���Z���`tKA�2zDB�I�j��E��q܌+���s B�	��x�j�N�C��hU�U%C��C�/HV�P0j�6c�PÂ�7w�C�	-6��!f�WrR&�"�gM1i�C�	� ��i��MuZP��Ǌ�Rr!�䕯F��p�g�5)>`XÁ�K5F	!��*j`6��wΒ��´;6�Y>!��
�	Wʽ#��N;[�d���J�d�!�ی�#�M��D\�'�I�!��n~������q��p��!G�!�LRα�vG�/�ȍ�w�^�#x!�dT�j|23+±#�m��EE#a!�Ę�?��ت� ��Z�C2�� 4!�$'+����eJջy�n�`DR�!�#
$�=P�Cة ��@��+T�!�(TNp�نG��=�Iw �2v!�D�?e�-�E�^!$��%�ńʢn!�K2�4�0�פ/��$K�D�MW!�d�ZWLI����+\�c��&et!�L1�>��̮<��4���*a!�� ܠ[qi�M$x뉵6���"Or|��C�UU(9�R�Q(HPIU"Or�i�-H��ٵ�^�D�����"O���W��x�z�E!�(��p"O���b,�R������ݠ "O�u��O�%@��J��,b��}�"Oj��w��;l|ށA�mC&�x5"@"O��0}H�\��� pu��"O ۇ�1yz����Pm�H��%"O������mi�<;�!*�|�R�"O�``/ɇy���C&`��-v@9:�"O>x����,�%z�n��Hp蘀""O�ʖ��vh#��cP,�f"O��r��(T*�sg�M�b�qh�"O���gH�1n`az�C�2G�R| �"O.h`�@J�*�XAl� 4���'"OЈÒk �%�Z��e�P�xf��	%"O&�J�+B$Lk��	�hd>��!"O����F�#�j�P5*[=f�`C"Ol4�P+=<^��Qd�"}�^U��"O��z��,s�4��"\�z�8R�"Omk�7�TuA��4A��	Bq"O�ٙ��R�|������O[>1�"O��@�K �l )T@�6=2Ԕ+�"O��ƭ��S�<�Q'&D=Bb�"O(�0G6zE�X�� eJ!��"OB�tz�LDQk �Ax�� �"O��X"�J�%4�U��*�kaE �"O�|�p��s�Ω�I1Q�	�"O�1���Yh�H��j3��*w"O������U"@�X���h.�=z"O��Ȥ� 29��y�M���"O�{�@Z d�x��ƤA��"B"Ot� &��z��#�AB�#0~d�"O�P�ui[@��6��3��D��"O2 P!��Q�՘��?`�8�c"O��K6�Y_ր=+��+~��]�P"Ot����ҰC�W'�@T4�D"O<e*TD�X�t�%�#�eX�"O@���LM�j��ݠ!�4�"O��H�/���;� �>�B:�"O �����2-QP�O c@L�#�"O5�f䕑C��A1A�W$���p"Oh\��L�e�l�L�(��+$"OH1�6`����r,ċ-1^��C"O��#���(/����g,�r>�Be"O��	��K4*���ؔ+!e���#"OZp���%�nP�Q*�*j��B"O�9���p,�%�Z�p�2��"O�����gH���A��
@(�"O�9���H�V0g��
�`��"Ol���HA�Dd����U:#�́��"O��)��/+����[f��e� "O,m	H��6��x!�"^�{�����"O,DB�C�0B���RH�!'}�"OJ�a�J�u	:2$��?�%�"O�I���<��J�]�6��"O��'mM#BT� 2���8���p@"O4ɠ�6�*qq �҂G��T�4"O���$@ &7V��h�+%��"O�]���j�I2�'ӕ\$xy�"OtHx2��;l��s)&�,xG"O��R���↺t2�p5,��y��hB��Ȓq�LA�D ҄�y
� D(
��R�U��@���J>(���p"O||�	۬M��!
W>�)��"OZ������b%I���/ ���"O�\���	�8�&\:�Jǜ �ه"O� �V��(h64ԀE��FwP�"O��
#��\�⸻��#A2`zf"Oa�F��+�Y��J4X\
L�"O̽rІ��-~Ԉ��B�'U�]QC"O t����#	�TH`���T=�q�"Ol��#+X�vgnx�u�́5C���"O���"C-���Շ��|B�"Oeb�bԼc�#�ʓ%��Ke"OD$ v�R�Q��:�-ˍTTA0"Oz��&�r���cf�Z([V��@"Oe,��EJt�1��Z�lX�Hc"O����L�Q?聴f��t?|<�d"O��	�*+�=��F�{<l\B�"OT��	���P0z%��D��1"O�|�v�D�b��	���9;�Qۅ"OjeѲ��p���k�#V�L'	Ya"O
\��%T�%���P�L�'LL�"O�9A"Ì�1N�C�t�d��"O��Em½;������I��R�"O�p��L�3'�)7 ���"O���`�&��d�& Y;4B<Ҧ"O�ȓ�ψ-#�N�Ғ�Y�T �г"OT(�7��h�e)���c*>��b"O(�p"��1#�a�N�:#��@�"ONq�6���
D�4,�0Ph4Лu"O���R��:!8��pJ\-&R���"O�� +S��F $>� *1"O<�8�R
	� ��Ś�`F�Y�"O��Z�I޴Y@V��$.!�����"OZx�RFѠrt�N,7D�t"ON�uBшy@2��B�0IH���"OP52���1���� �~�hhy��I�<Yce�	_S�:B��t��� �G�<�ƈ�;Z8<p O@�Vj�a�m�<���K�M`�S�Jܟ#�6+��_b�<�+o*�Lم�B�YI�5h3��a�<�2gU+<=��`�c�l�S���D�<	'��RG��x�BP�).44�A�<YQ�U �BUPp�q6����Ji�<y��ܹ88�sIP2�cejLd�<A�I�9�"��g�X][���/�u�<��)�	_
]�4kH�	�l��`SI�<�&�&B<\!��LBvH*���J�<����3GD���f�-ЈA2���^�<�ǡ�<XZ�Y���O�B,r�ŔE�<���%�L,~��#��K; B�ɡ	ZR Y�+(��iEm�740C�I#u��0�e�,;�����j�RC�I�j��T'L=qP���CD�#T�C�ɿ9���+RG�� UH��F#"s�TB�ɚU��m`��G��0|"b�!�hC䉽S����w��?FJI��T�
B�I.�h� �n��+f�YuEߵ^x�C�I�D�50R��r	�`a��$�`C�ɟ`��)3�H*"s�-ha�\�ZpC䉇ac�ۄF�n�he�H�JC��zT6�Ȓ��EL� �W3�8C��?�0���7!�ʗ6	�B�	"NP��$f�� pR	5ttB�	�k��9����[* �� ܦ�4B�)� ����ʖ1���C ����hV"Oh�@�NۆF�ɐ�$��%�* 0!"OP��䇚�c"�2��ShЌm��"O⠐��-0�}#�(/���Q"Ol��eM1��2&��3F�*���"OЩ�QG:4�l% 1�?d�F�	U"Or�U�^�ҝ��LU�Y��D�g"OP�QT=P8� ���1�ֵ��"O��MŧD��4C�jM�K�x��"O��g�^TF2MzSCK�}�x|kU"O6�UL��d�0�	�k�X�B�"O8U�p�	8�:��NV\�["O�Y���fw�[-A:kh"��B"O�\qGP#9]]{��'gD��v"O�}��D0A�,6��;Y<F1�"O,�a����X�!�F �~Y��"O�}� �X�ب�Sd�0%���`"O��	��<?Kv�Ȯq~���E"O���F�	�W$Q�҂��0D� �"O�H�6.��cιz�B\e��HF"Oh}���Ex�S*
lbR�h6"Ox=cĀL�Q����V\p����"Oީ#���oꮜ���Zp�]�'"Om�R�/T���g�#=���8�"Oxh��Ps4��/�^q @"R"O�(476��$c5��,s��`�"Ot��)o@t��-��|xeZ7"O�MaRL�~���٩(\���r"OZ��0�ՠ*���Рb�>���8�"ORx���eJ)ো!@fB{D"O(q ��@�Cܼp@���#+�)S"O�:g�I�0�@�����,�8�"O0�{C�	���HFCϗ�<�PF"O���"@4{�t=Q�O0jϰ +�"O4͑@�ikTZ�$Q�=�t��"O~x�W��u6��:�\Q�ޑ+�"O�c1L�_o��qEB	:4�"O���4���8u��	g�j}	"Opٲ��W?K�r���ו@����F"O����b�6B�N4�iĄey4�Aw"OЕ��X5q����W��k��k�"Or��AG��_�����> ���"O�@2��ڪ;,���ϊN��ib""O������v�Zl#�M�Cά`c�O��@���C���!�Z:`5x��O��=E��h^�^��RW
�?6��Щ 嘠r!�D��^�D���B��;��l:Vĝ.&�!�$�I)�p0q#�d���%��`�!�	��<3�'I�q���	�3:CrC�IpL��!G�	"\gz4B�'ϦbrPC�	.|�af�vǞ`K��
�P[VB�I�O�� ��9vo�`�dȚc@B䉺L�9H�G�8X�α�*H�@��C�I�jRm��L2Ҿ-ZT���} �B�I�	l8�GiN+, ��) eO�ۤB䉄3�*�0Ō�vl�AsB�L��FB�	�o8�x��}q�-Z�˖EB�I;#%�h wgP�y�\3���:1�B�ɤN���el̥U����GI�`�jB䉻D>��ir�E�2��i� ��d�zB�	�D�r��Q�mB�(B� C��&���(@�M�F!�i�,y�B�	6p���M�	�Ţp�ǒA��C�ɷ,TІ�Y�R%Hh�QjC�>-~C�)� 8$��-A8��})$�<W��h1"O�a�� \O<ģ��IoQ yK�"O���פ�F���bK�%��˶"O��1�[2k�P����s^�(��"O�U�Z$^��J�&y�IQ"O�A��d�2��Q%1l4dI�"OHᩳ�_�\�� ��3n0�	��"O0%`�*��B���+$b�O��zS�D���L���n�z0�OC�ɦKцDLC2S�, ��3�C�	�$x$Bf�,�t����s0�C�Ix�̸�J+&�m�u`ݟevHB�
���ڧ��^+�0C�nΟQ��C����mc�O*h�����?R8�C�(P_x��IB�6��H;�bݳ3PC䉝47"9j���S�Z(����"fC�I�)'ڑ[�d�#h�:�c��[(q�"B�q��`�/Kb<dL:` �B�	>vXv�P�	AX<��d&�2,~B䉊u�|,bS� 6W/��i%Kg�C�;[a�92�piة;%�@0.�C��<e�$����-j?���Ff]�B䉜QQ���	c��M��I`ŮB�	]#D����ހ�8��D/�B�ɒ�T�nĢa�*d�p#�=s�C�əF��,��!�⬅���L���B�	�C	R�A5������F#��C�ɼ/�6�st�O/t*�e�G.�-O��C��,�@zeň�8qn��v)���C�	"M؊a�@a֌?�2%2#N�:g�C�I.���7ɖ�\�u�䑥V��C�-kyI�NȦz)�`��	�*iG�B�?�69H�
�[�@�Ѓ�F��B�	��H�a���
���v�H�0רB�	{���§g��w��)�AELg�C�I��8e���6�q��&P�Ou�C�ɇw��Wd*d���ǁ��:���"Onq[�(����k1&I`|��JE"OV�7�/s� tb%Ċl^�Q�"O�癎hh���Tg�*Uء(�"O����,��Gz�Ձ����2`��`"O�xA�/׉]r���LY���6"O�0�Aq �)q�a��{G�Y*"O�ݠ'/�>:�T���H�~6*��'w�	ß�F{J?�i����n� ��j�,��cg�!D�T�� f�:6��8Z;���3>D��e�4fL����uz�z�;D�l�0�Ӹ@���W���Cp�f ,D�4��EA����-e�J	JAl*D�p��"�7x�#�IL0%� j*D���B�-�<�ءa˝`�%ID�(D����,�(s����
�V
�Őv�'D�,��]#p#�48����7���i D����+*�A� E3i�@0Щ!D���d	+�`x�+j�Fp�£2D�8hB�:�Z�{ !G[/��K��6D��ju��q�(!�D c���Y�6D�x�`F� n��8��A�T�f��M2D������B8����A�4�H�E 5D��x����~�CF)C0L�f��e�5D�\ꓮ[�[u�0��+-�e�ҧ0D�����T�UF�A���&7H����k0D�hp���uOȵy��G�#��a1D�L�:D8��`9i$.�e!;D�� �@;��X~�ђa!x���"OΌ��/\ _��`�Gv1X�"O�����(k�L���/T=��"ODȻ��\�y J�Q�A��0AB�"O���
�M��D"
3,{�4rS"O�ĉ#�M����*Ƌ��
��X�<��%A~&�i�r�� T���)y�<�`�@�z#R\y#e�'.x�!��E\x�<V$(X j�:$��[ʀ�BN�������FJ🜖�(OFX:(�I�΁iA/Y���u��"O�9鱢�6:g�����Gq���"OJ-U�T4B���#Nu�!b"O�e�̗��`ș�'WҠ2"O��H�NY?�8Ě�CJ�b�� �u"O�� F�e��Z2���w@�8!�"O��XBV�&���S-�9Ƥ�u"O
E�6�z�B6Cƍa�R��T"Oj�v���~nZ�Aw���H�t"O�i��X��ۓ��#R�l��"OZĂwč�1_�E M�uO4m*�"O ��r8��%/>�d�U"O~�@tǖ�OKJsUY�@m�)��"O�M���( ކ��lB6$V.5z�"O6Y�6ֺxn���@�ڎ��!h�"OB5���" �hm:�*��#�bh2#"OZ}��	�Bt�cu�(M �[�"OL9��

7rD�8%j]�7H�8�"O��fF�1�HQX�J��I@Հ�"O4�E�(�N�0��T>f1$H��"O������ZNe+ �±6&�غ�"O|�Y���.g�شz�K��Xi�"O"��"eT������%0u'�2	�'G$P���6V����쟒;P)J�'e|p�e���pBd��tS�'�jYr�O<>�< �s'�'H� B�'X�"�J�(r��K�%ح=�j��'�����ڋH�ru��m��4�e�	�'�`}��6 �����:H��t�ȓY`^���O׿���q��M�[ ��ȓJ�ڈ�0E8L_P����Gh<�ȓH]�U��<I��-h"��*掅��O�Ԅ$�5��q���X
����xh(����!R�m�0>�ćȓOq�`�Έ�S$(局)S�^vPل�e��m��/+q6Ĺ��޶>�2!�ȓ!���q�l�6c�2�괣Up�L��m,8誄�:"n��R��0���ȓ� �;����0͂���(Q�a�ȓ"�*=�eHVx|���S�$$�@��ȓ���Ñi�'��P��X���`��-h0��ʗ�� ����ȓ�Ȫp�W��$�'a�F�z����걡��̀��E`G��#�y�� x�����D6'��@�_=�y2�CTpQ�Є>56�yG*��yr��F�x@)CÁ�zFD�2F�܍�y���im&9��A�:��4�"D*�y��0l4�T�(٤���x@ʱ�y��6�\4`p)����rl��y��S�%5~Q3"�آ�ؠ�fGG��y�OU�6jb
ط}�l��ڄ�y��=f
�i�H��}�v»�y"���852�*J,�- а	�-�yr'��*���ie��v�2!��ɉ�y
� ~�J�fF�rդ\*f�E� (m�p"O i#�j�9i:��s�Ԁ	l�k�"OH���fJ�B`�Q8�fյo�a
�"O��9��ÂD���i�T��!�U"O(e�g��;�.5��cһD���k�"OE�2I@A���α@����"OXQ*#��޺��B��<yq"O�F(�Ll��D���
"O�Tۦ���De�|�&�Ȓ��$"O�l��GJ69�L�3k!?�Z@�b"O` rs_-6`������6��CG"OQy���_�NpPs�՜Y����"O<My�ↅ6:tH�6�ķi@�d�V"O��3��W�5���tOl��"O����ۜV��yR$�\��`�"O4�Y4��Yhb"b &���"O�x+ n�W���Wf }t�)*�"O��ړ,[�:v��pdօ=frp��"O$EO_�'��R�J`�t�`"OV%�e��T8��K4HPb1h�"O���%�8u����+Z �<���"O���o�����@J�m���E"O<���<Q���w���,��|��"O�\3�O
?/�)0��G�@|�t"O��%T���3F�R�wA�4"O�	�P"秃�0	�����17!���<rH�Z���m��	q5ρB�!��[,e����?U�b�#��g�!��uO�z����y���W�N�`�!���^Q61��I�y
)@1�R�6�!򄏓S����a�M� �q�9 �!�ִ]a"iJ�X">ʍ��F�v�!��S��Ҝ��h����K��!��{�|���J&m�
�d�8J�!�Œ_����' � J�ޤb0#D�Ar!�D�hX�H���  ��0f��MC!�@�X`&k�,� �{s�U*s?!�7[ ���M�R�$��a�;!�d@���0	Y�WL�(����%V!��ٳrt���U��"q����47!�I����7l�?1����5w!�D�y-����
��)h&�Zlh!�DL�]˴(�b/�2�ƅ��B�&"Oƴ� kC�JH�@z\$<�u"O��(�Q�d��`�� �`�"O��C6�B�ݐ��=�$]�@"O��@2"K�/5*���K����J�"O�%�fm�4{����k�d���r�"O:a�	��@b�[���c��2�"Oz�3��z������C��${u"OB�Ѓ�]�8�Z *M���C&"O��)u�ݷFd�YIR���=�!"Oh����))��+&h�)�0���"O�\ȇm��W���hdɿ��YJ�"O���I�?^&^,����R��3�"O H�V��;K��|�t��"O��X��F1e�pe3�'ݜ;�Xir&"OҌS���/!>%�0F5_�� ��"O>�2�=�r���BZ�K��)!�"O$ ��ϕw����0 ��?�<�I�"O�륅_�t8�,H�n]2t���E"O�If�~��!W��y�:\1�"O�y��bK�@�����A1q��|
�"O(�+�i2C�\��"A��$�
�32"O� ��� ��G�Τ��"J�Q!*�x�"O��[��!M!h<����c4��P"O�a���g�t�$�'%�P)�"O�-��C^�`���Ġw۞�8�"O���1��j����N�	��Y�"Or a���N�X�ʢ͍�_OҜ�R"O��� ��|�@���.FV|4��"O,�����z2�@�>a27��A!��Ў����d�/e�0�øm !�$N
}����!�� ���箞?2�!�P*y��(��ȏ�o��!u��J�!�$��e����K;j����J^�j!�D�!{�����.ʹbb}��hEA�!�ޞL�T��1"�W�lbN�T�!���9Z�4��՞X�`�`&�7|!���7������sm�����,Fa!�Du�dGS1[\���KR�$a!�dN%h�0;V��)3s���֠�?;D!�$�)i�޼�SM�|y.9�4���j&!�$��t��DƀM���@G��!�d۟.N�y�ň�.`��)� C�3!�䊉��T��ڸU8X@ѯA�V-!��"��Eڲ�[)b����
	y�!�� yByy�i��);R��6�._�!�ĉ�ac�	BF����Z��T�!�43�
qA��B� ���!���!�DV�;	$��o�6��|Q R�!�1�h���&]���yJ�L
�%�!�@�sjt�y�a��+�6����!��W�&�±�K�Z4 ��M'3�!�$ _xpx�j��i���y��߭'�!�E�PPa��W�Z�`5���8'�!��ö_�<P	��):~V�R-ڸ`�!�
w���PsE �zt����Lխo�!��ٜg��E�e��;]u���ťP�!�$�3`�9F�C�8��Axe c�!��ք"�04걤���x(�!�$�)q�ac �h�(�c�����!���"��	��	�)S ����[n�!�^*NTtZ�@ �>�����N�!�U����7�M1��PJ�8T�!�$S2���se��A���(T(W=I�!�DŇ5|x�qwM�.��t �f̽q!򄅲\��ڤPol��&�'qY!����Z!����pT|�p�d��+��� "V,�d.� x��dNO��y�)d_֝P���`�\刡`ҳ�y�O\n��
�_�<i�5�y����!�t��&/A !v��IE$�&�y2 	[��e���Ɠ�������yb��12-�b�N�q0!�HA�y"�Ä?�jyݴ2%�u��*!�d�:���� *ܰ����"�!�$�n"��<wѤ���f!TO!�d�)5Ka:�b�<}�0a"�U�E!���� ���U9IȁH�$Q�Q�!��h�aqpbR�pD�92��e�!��N��ؤJ̰�H�fGp!� �+�$�XÆ��޸pt ąXU!�$����2�P�*�µ���¨>!�D�8�ys�g��9eL��HK�l�!�$A%ٮ���Y(X�Y��G"M!�䊌'`ÕS������Q�!�"��1q��1A�a�r�B�!�� �X�*��4Ӭ������n�\��"O>��`�N<f��t�-������"O�@k�*�q�2�8�,��6��A T"OX��ჴdS 1˞�Gd�Ӥ"O���D$�TYhRj�I5r� r"Oj���`׫X���؀)]K80�$"Op����-�����M2&��"O�u(�dS1djTD���ͭu!���W"O�u@OC���J�R�j8hb"O���ƀC�y�,IbBnN�vr��%"OJep$�0S�"!m�-VX� ӷ"O�,0s�ĶU�@#q�ȰL9�E[�"O~EU�@z���q�ɛ87*F0�"O���C�L� �f!
G�N14��E"O���2��l�
���W�-�LR�"O��{��͵/�
�(&#�$�ъE"ON��n\����Dc�E�<�w"O�ejN =��Q((t0���"Oj=qf�@@�(˵�-6"��X�"Oҥ�&�N)&+�À�������"O��p&',���� F]�c��u8�"O�`�����1� �=�L���"O��H�	����F-R�8�q7"Ol7!�U
�t@!KR8;�pS�"O^�0��("�5� ��5-6RC�"O���u&��/f�M[ǩ�9�H\14"O�:��R9S��&�ܓ/�x�u"O��p�쟑k�z)���
�7@Es�"O*�r�2�6,AbI�9|Q&Ep�"O�Ԑ��0MV�PA+�<1�`$��"OD	i�䌣	V����?�p�8�"O@!U��2A3B��A�λoq���F"Oʭ: ?��mR��˕hmD�"O�X�넪q>���q�A�U�#"O����N�0_�$̑��I�ҕ�c"O��5�W>���#gLP/V�� "O�x�@i��Z `R� �9ZG@uR!"O��6d w��8�7o� t�tY�1"O�AoL�.P���㈜�m˴���"O�I��"�bcgՑ�Ft�"O�ix���
Z��7�E�4� e0b"O�֎ �#�L�Y$F�Z��ñ"Of����+��8��E-���&"O��W�P��:q\���Z�"OLa��a$��1��b�%�"O��X5/[l��8C��-w��-��"O�/��a��L4/�:��S���!�I [d�r���X�:�-Z�V�!��,D�dE�J� oJ�Cv	i�!�Ćt����əgk.��_�!�DΗU�8iS"��'F�J͘Ӏ��K'!�d������I��_?-C S�'!�$?�F��Ǎ��aO
�'�V>U!��ɁX����g6�:����9�!��+�(�aU�ǾL�'�ͬ0�!�ĖW�!Q�i�>}��8q��,�!�����t��g��T��M�bÅ�{4!�d]
���.F%�����"6C!���
fcI��ڸv�u����M=!�D�t�x��3�Y�.����5!!�u�� @V:���,Ay;<��"On�p��K����]�@�J$�_��yr�ˊ%���``�L���8��b��y��FB4.<�`FRj�������y
� �<�r��{vbT�&�7�z�"ON2V�֐U�֨Bb`̏��SP"O�]��B_i�v�bp.Q�i�x""O�Y�a�>3n�����<&N�YP�"OB�۲�T�+�`dz&		��<P� "O:蹲L�}_�飀� X"l0�"O:�	�J��0#��y�f¥#����"O��dL!H&
�E�F�(]9�"OƱ���
��Hu��V(#��{�"O�Չ��P3Hp<��@�n��ؘ�"O�hDCز~v�<bjӓ^��d��"O��s�a̮KiP�RI�$k�b�H�"O�h�GR���]��	�b"OZ}���S��(s�J�"��i "O�Eᓈ[*�ʘX4(ޟ}�(��P"O������3�bm(�g�����"Ol��N�M���V�̍r��"O^���j 1�x afS+QT�}�v"O�uq ��b���#����x&�0p�"O\�9R.�3'D��j��$=i�"Oz�*��*M ��3j�4t@ܸ�D"O"���GI�">�ćX�v�2$��"O<]���g�.�6G[�r2a��"O��r m�>B�+�g�+Y�h�"O
<���ǨGJR<���'E�|Y�"O*�P��[\�`���^���A�"OP�k��L�p��y��Y���r�"O�apD���xiN��떦_�z�P5"O���a�¯xЬ�鏼�U�E"O��Hk�m��I�@Gԓf�ԥ:�"O��b�֟-������$��"O��"/�=x/v5�o�5o�����"O�S�"�(��qh���)Ȧ� "OV��&o�k6������}����d"O�I�H�<F����U!���"O��h��ա+w���dK׫�v���"O�Q�q%бr�H�%+�P��trQ"O�e�tj��.��@D�S6m��BQ"O�p"���+*^<�bh�Mΐ��F"O������vN�)&hޔ@�.%*�"O@�b +�8Sd���"�2�C "O��5I
$\�Ha��/[V��i�"Oݓ4��-�X�9�CZ�X�~���"O�d�@��z��U(�Dy��ye"O�}�^<6 ��B���gpp���"O�J��20���ir�4iY�����~��s��F�&&�9�E
Tp�!��Dkm�+P-L�n�Q7	�H�І�}�Y�V%�|�R�ǧ>U�A�ȓ)�ڕ��,c�ar�/�4لȓ0�D�D��+*�X�y�FЍ0X݄�>V����:��퐄*�%@W�<��3�\�z���O�J�!� �%��qҠ�MˉPlI��L�'�ȓ0��1UP*!��A!�?/:���%��	��*���8&+����h��B`.����G���1)�y�����&�j�% ��ՙ��5R2�p�ȓZԎ%�g�!�y�5*/ \U��v��z����B2��b��;_F��ȓl_���+�+f����")�Q�ȓF�JH����T�v��#�>�@L���<�cAbJ�i�z���m֮fK(8�ȓx|}���L=l�d)]`� ��S�? �t���Q�vtIѶd�I�I��"O��� L�꼃".���p�"O�8ȁhيD<�U�d�D�j�TP�"Oh�rhW�#R� �'�=qL�t��"O a��rcNU��H.���"OX(aA�� ��0���S�0~���"OhVJ��(P���!`F%����4"O�L����u����������Ԝ�@*T�)�'C��A��ǁ$6�����n�1i���ȓ"�^�چ�R9j+�8s�b��H��|�ȓ{��Y5�&db����kș����ȓ:����!��&X��B�)X����%;T@>��B�\�F�ȓm��ܨ��
��ȫ�݁"	"q�ȓ4K\d2%^|Ȥ+c�OA
���l����Q&2Ga���D�� �ȓ�5ꒂH"A�S��R�`�$��}C�����3{�ĩ�7@�(����r�'u�ֆ.B��|2uH^�wcv!�'��2f��	��f)1y��j��O6��'VAZ�� ��*} D"O:��V�ðO�y	���H�nM����?|O��Kf��
>���Ь,T�T2��IFx��8w.���da�Bi/+Ӳ|�`c-D��%��)^��C$�Q�!��ajSE.�O��5���`M��Df0���ϝ�D��u���J�';|u�e�H :|���$ߕc��
�'�����Je8	�)`@�E�	�'PYꕉQ+;ܜ�9���&\70��}B^��F��c��^��y�c��r���0���6X����'�@a֎�=*�t���=^�@|3�'�ў�>	�g8O\�Cr��|y($8�$E_�R��&"O��ˤb��بƣ�%WF��W������WL��`����>Y~�� �K���$?!��V����J�D�0�n�S,E�<��M�%x�4D�AF�1b��]
��K�Ą]���t���3���.n��Ƨ���t��C�<�I�����vQ4]�a	GG|q򥊓&a�4�"a!<O: �����xK�-K�US��3
O~��R��!Z�,�w�S�bn����.]��O�'�Q>�TC��٦5�qZ-N`��Va1O�eӌ�#Z�>��QJX.��4�t�%+K!�( fXa�d喵,���"�^4VF�'b>��=	��I�(E��L���"-# �q�,Y�E!�W�D�VIq�D�jJ<q��]	�!���c����&��ָ��T0"�!��3.�t1����J�B���KܶO"�&�Ӻ���s�dp���B�G����+
&a{B�<�I�R��B`B%�4�0r)��%#B�I<0�H��a��h>��T�<s�"?��	ٻWg6��(A+n&��\�@��4O�c�Є�xy^}'AMU��!�`��\4JC� F�q��W�Z`����U�pC�I�:�tB�=�J�L�3Q�B�I�Y=��"�X�������=��B�� �V]"a�]K�xX"��$�B����m�q�;]�̚�Ӣr+C�I��9AN4#^�y&����<C�	f��SN�-*V ��� �2C�ɨD���o��"�
�H�C�I�� p��³D<Ri��A'@��⟠E{J?��� 00(�AWMS&
��bgC6D��I4+g�$�0:ّ��xg�������Sg��{
r��r�I6i�*�n�8=��IVy�L7��� ���sɘ'~O��gnH� �0�"O���G5�4x�Ǜ%2�R��Q"O�A���ɽn�)��4��i�"O|���(��b�v+d�B�+"�Ɇ�hO��C�sd���4����oY;�!���3#Cr=�u�Qfet|YQO��vl!��S�;���R,1eZ辉Pq"O����� �`q�TQ�ե(Ŧ���"Ob蓧d/}�	�`��-Y�R�:eQ�|�	�qO��<9�hJ�
�d ሒ-|��8CX�<)oBzN�s��+�<�ÁS�'Nў��Z�i��L'1�~� w��=<��Ԅȓl��%�fd�W��8uo�:���ȓE�pP#�iQ `�:���nN9"��F|��ӛI����Qm�K�^�j���i{��IT��P���ػh�ԘP�b�6f@̨ 6D��˕#��wD� �U惣V����5D�$K� &ɒ=�D��}��s��h�4�'��' �	H�i���Y5$��X�!��$���c��"D��{�d�>'vT���M�I�$�֥�������E�fE���&s*^�У�#���?a��IL+[��j�	ɐ����R!�$iO.D�q�V+��7��8����c���l��kZ)� KV>�~�i&��!� C�I�W�Bh���F�&�fX�]��4"<ɍ��?Ej�`ǯ4PJ2tB��78�5�%4D��	Y�oF���F*S@N�� �)�<��哛!f80S
A%���#[��B�(G��h��ز$T�|���� v���Y�IVx�l+�I-3�m�$M�??�8����+�O�r��P�v
X���q`���N��ȓO2���"E�/$���G'�Q�^�mE�������yR-L�#�<��W��=w�eAa�yrON�{R,\X��JG�vd+4'Ђ��D"�S��ͪ�\9?�f�a�m\x� Y�"O�@j���p/���5̐?P��=��i�P���IG�� �S�̴���lH�r�F"=YN<���-��Y�h�@�o.xL�PbW/��Z�*B�$�ͳЪǗ	���z�c�=1����?�	�B��y"���"�� ��	i�B�(Z��B�J�9f~p03��^��B��15�,���
4'��H�>��B�I:J	�a�nCV��R�*G�02�Ol��$��'+�u����22�%	B(�t�!�Նh�^��l��Y�ظ�IFR�!�x����ؘL��80�hKA����'��O?7	>-m�R��^6���&�M�V�!�Ϯ�������{yPyJƦ�*�!�dʡD�y�t���<��S�ʎMa|R�|�h�2W~��Ȍ�;�
��cO������p>)%ۭaJ|AD)�THr�j���1�OV���gQ;<ul,���2{�c�"O^y���=y�9��E�V�Z�E�xbS�$'�b?��n�_�P��,A�]�0m�6$D�l¦��&Gd�`��+L8I���"D�I�AB�;��K7!ʩ_����%h2��p<�AJ�3-�m�G
��Z�.����x��P�)w��JLjE�C�
�y��
��Ļ2�@˪���熛�x��'�$	S�
�78{̸���H(G@��B����>A��$̘41�j�:� ��Z%����y�l?�|�����%�0�x�N�yr�9�h4���?�T���א��'�ўD�'S@�B��ߒV���Cl�5~0h
��� �<��f(/�9&'�
����G�Iox�d7@#��xC�@�Bf���c'D��Q��T�<̈́�h��_y�e�$�#D�X�a)�9>$r]ru�IoP�)���5D�L�@̣,4^�a�LF�+m�ca3D��3���	-h� [u�E
ʐ-��l1D���g/A).�����'z�����.D�0zQd�'=� ���@�8>�����1D��tk�o.HcĬ8thf���A.D���D�I�XVC�"��)��o+D�(jFJʗ!�D���͖�f�d�)D���!�Y,p+\�W͒�$��k)D����Ѣl+�@����J�{DM(D�,H�n�@����˺.�%���&D�"-�� ?Z@�Wh�c��pH��1D�l�M��h��6sɫ$@#D��[G
Y�b,�h�r���^޼�tk>D�,
�g�;yX)��OJQ����1D�@�+�Ġ#��҇��
�0D�t%�H�6��\���3C̩c#D�,@�hֵd�|��֎]�pp�eHE?D��cPoի2={d���@ Lm	�(*D��а%V�d�*5�a�p�I;�/+D��j&jOl�r�J�,��g�(D���g�W.0U�����3��@���1D�\СNðr�ޠ��Vek�|!�k/D�D���^��ʵ�E�̼�'�?D�8��F�*Q8�k��M{XS� <D��)��H�N/9�ʓP��)�U�:D�8!������IqP�Ǘ|Ct��W�8D���/�g�p���8m��@Q�8D�(���o�z`X��C%4|��9!7D�l����ma�1���
M���n5D�\���8
�QѦb��nйwL!D�蛃N��l2!���Q��8Sg�4D�D����`�N�B$�Ͻ?���z�L7D��H�
�`��E�E�Y�wҜR�!"D������q��<Z��Z|x��"D����$��]�p�m��`�Z��u(+D���) �
P�#��D�5�qL-�O��@V��#I$iyHQk�4<c�*/_z�sq"O�) �A8?q$��3�ݞVz�I"O�p�f8X:��FH�"v"O�X��l���JH�I=��	��"O A��KT�{qP�Q��;|a�z�"O��REbP7'�� �a\Ba�4�1"O�ݢ�C	\9��"�Nto(���"O@\ ��B)�h�c4���6U���"ON�ѥ�7-�|D2P(D�Jn�1�"O�[��ݪt���a�A��;8�y[�"OjS�M�MHaP� W�-�x��"O����p_?8$H)�G�
pν�ȓ�P	j�ĉ�fF)ۢe�%M�nȇȓ`����"޲(��XCt�Ŝ"�Y�ȓ,OI��&�/=|��r�M�3A~�ȓ�}�æ+S��� b�3i�=�ȓS�x�1�L�1������*<�L��e4��ө7b��i�I�N�4��Ku�A�S)3	���k>���wL�R�J�-R,�� �lW��`h��1BZ�6}�hD����~��Q��&��I3��3Q1�L`�Ȥ]�q��E�����&B���S�O�	C`��.J녁оFT4�p�'w��Xf�Ǵb Y5@�8��5�-OTp�1�(x�;�H6O� �1xP+	#����ǌ"C��6�'D�X1���
`�AW�I��rN�;��c��v��t��I-2�Q����n"�}ᓀ� -S �<�e@�/ <�i�Dl&�u�K|
���,��3��N,? H�x&�t�<��,e�H+i
%f��|���1/#��b�̀�V��p"�JφȎG��'��I ׆	�/�D����B��&��'	���*Q�I	�8R�+wSj�0� H;������!@D��"��׊a	��G}�`T�C���b�E�5���BP�+ڨODA)�H��(gX�CsJ�)���E UFS>���UH�:��A=y|ȕ�ZMX���I�Xb�`���2	�,@$��=�4�VWS��2�`H" @����C�zSx��%[�7�8`�?���B$1�|h��e%��unU}�<��☨P���a�n�~80�BA�4o,��Ju)���w��.��U�O��h��D��z�8�O�(+`�R)e�,�Y%�N����b��h�a��6��'_D�d�%�ـy�te�`LѮ�uz��)Y���������z ��&�~t��;_\��h��p��<�CX�f�(�$�.:�`��
J�1�'�f�)�
K�{9�)ZFIDHf��M��w���B�X�.���g�bU�5���,���R�?�I�^[�CgJ�'(�����E�Rf�&%+��;2�;����F޴+`�I�>'K��c�^�%c�u��&$ !��/@����y(�" V�)�#4Z-y�*Q�~����Nt�����W��D���D���y�h��/e&�;�d�\��y�Jʚ@�l1�r�ED���k>�a���1+o0�c$D_��YYt��AĜ�B"LYD|Q�i�M��8t��`�b"K�I3ȕ(r��`���-�,�`���>�A6���J%�G铟f�d�XT�,au��j,Ց{�&�9��F`�fg�+�T��)�<a$Ƒ�c|���r�� ����#��e���.Mj(x�L����Ϡ���q dUȈS���Q��ŭ+Ed<�!ۊ#�����3]e��� �)C��(�
�IT�-�FX:�?9��{љ�ń&-���C}�֝�����m��иU�\&�<��SÒHE-���Ϗ^]�� ��Қ>��4�D��o��ذ͟�N�'=����Z�H����)�%l԰yn�s_Phs��y,ݩ����TN�iD.IJ�O�?��]ϻpc4)�ȄHĦ���Lwl,uK���Ҟt��,�N���1���|:���Lξ���h�pl0IK��A#Pt�y��ek���!�|$��nZ.0�qЖ�P80eJs/��_N���^�����ͿId�r+�"[6yS�'�^��Qm�+�,��S6auFP���о��!jR�%W.MC�'E_
��1mK��"�IR�(��U���i���Gh�'� �hX7Nl%�'�R ���� d���Z�|��1cID�KE�4����0�1
ԯu_�����o$���HkڰZ5\�ŇI8 �X�P��w�ܟ H��&b����>-l
��L��WJ�r��>k�@�R��N��u"1%��"a4��fi�?/h$?�ݻszI�XY���ҒU���P��34��ԑ��]�R�$1�%��?C��]R�-yeK�]���
`ĔD�-7Ct��eI3 �m�P��B���R��X��(30��?:�GV�%�r��$G��dx�&�A� �0��А�:�0�Ů*��I�=	 -�7�J��b�E��l����%��3�ҕ�#��O����r�[�]�`�gX�<�Mⴊ�,s���e�6u����-��H�������U�P���Y�9������M��%�􈗁6W�,Р$Z�y��A´j:�d�4�������5E��"����L�!���k�[�@��
¿� ��t�[+K���ňU>6�6�ې�C-Jݢ��T���]�T�Cê?���weL��OE7zӆ4��i����(�Px��AL�DA	kdN���)ʥQ�N)����?P� !4��h�ir%���
�f�+��P�A��qʶ��L!��.G>T�	I�i[&m��\�'����OZ;{���pa����6w�x�"�i�u!QaB����'d�N��|���#n�Dbv�.*����$'�	bL�`�J��,K�H�Q�L!!D�=b����ʃemI(�A&7�,��P�ʈ"�̑���^. [3CH�8
8��x��I48qpB�$�Rұ��#Lf��4#��p?�R`�=�� �'��	c�LL�͆,����"��h�H���rаڴXqx�Y�o1���"cZ�y�͘�QbfX�p/ۭY�v�8]@0���[r��"쑃=��E#�HKN"]����/�1���شR����d![z�����8��ecU�
K4i��p>�����0��Ί�"1�Q��I�n�ǥC�:����H��#�C�w���,F_t����	�28(.T��g�E�t���͏L�%G{�K�`��!�4'�?�֠��.��'�д���̬"��YV�#Ktb���(L=����Qf��x���]�tS��� M Q	A�%|��ak�,�O����I�@�X�G	
��"@��:L�@j�Ġ~��tK��6V3����d$G�@ ��)�� H3�3�B�;r�y���P��U!`���1�"O���˔�n#��읜L����oI(Y�L��F��m���$������u�<k.�5��\N��1��Q�%��)^�`�UL��H�ԙ�Bn]5Y�~��%�K�YǠ-��l�9)��U�����FM�`��mq7���S:�kc��.4��� MN ?�����13N2�"��
��(�c��p�8�D�m�'#���a������ˋ_V��"�)�l��
،ؼ�ȥ!�>)�)�����A-�	[\��_�-�L�AÂ�;<�|� ��``J���lŚ1&�`��/�~�`()�2�L�A�I�8u!aݾE�e`ح_����A
U8��-[�Y����A܎K�lZ8ͪ]�&�A�Y�(��Q�Ɂ{>qȑn��*���H�iH⬴)I>A�	�J䢨���Б���6�؜�DnJy<yؑ,�$L5��*]�{)XTJ��޹��u�q��8����w�ĦB�𭛀l� F-����y-^Db�韻��7M�0J��\�d犟}���$Eخ0=)�J�7N~�ؙ�/�)NW��z#CP1I��T�$G����T��.1>�T��}q�!�e		A�j14�A
=�H4��g^\��0T�BK���hĂyy�<��'��kZ��ab�\��80RE�9ZS�D��U)JM��΀%X������aL���TZ����Z:[_�|{P�#d8�Ԡ0��x��9nJ�-:qᆂI��<�� �1
�
��b	;hA�Z�� ��#Sώ6�J���B">�ۇ�=5��L����Z�|Q34b��[��4�T5��+״@$.��
<6��(��I�Ҩ��ꐇ>�v݂Ēx�O��ub���)D�#_ �
� �0�F1� ��^�VtyR��,[��Xr"�E[ у�Q��\ɪݴJP�q�ˤ{sf9�5B\*]�J�;1����S�]!��	:j���C$T��x� 	̷xOn�ˆ���8KXu�q �$	��Xۇ9o�����6�P���̷zFz�N�L-��-�0\��ધ�5n4��t˕0(� ��+�/xI�P��f�Y�'�Zi�b��k~�J�3k1��+��)H�����"�j�|
�H�B��|���z���qÀ+di��iʤ�$:CP^R`Y2��'>�-x���"'���꤄�h_()a(��f�� 1$���{x�8р�W�^�*)��Gj�a�@��L5I%ĩa���D�6sl�P! �R�P$P0ؐ"r�E��ΎLL"�bA/0�����d�e�ߢ �)K�1�p��1��Y$�b�`��x�P5��%��!�j4[�ś�Qի���貭@�m4��(h��V
X+��v�9�	*j,f��ҨW���;���=ҁ�Fb)�be���8p�������i*n��R��'��sghX�>��N
C2����ٱ_f)BC��b����P$+< �1�`W 7�����r;ʝ��&� JO\吰ף��	���i�1�tD�
[jbA`r>�����"NEJ��شA-D#�G8a�H�[
��
��'-��h���IQPɻ�)�6b�9��B݉.�}��Qc�1 ��#���r)P�[��IQ�sx�̓(�y�u�O�3��ŉSDd�T���6^��ԅ�	�@4J��@nqON(
�)N!4\`�9P�E�-��E�$��"P��zc%G��ə�!ڂ/��L �ჷ9��3�l}�2H'�8�N�vu�y��`�,qO`�1� X#jN�}��%�&exvl�7#�"�)��d�|Z�hR�GG&}0b୻`��)I�!7�����I�̼�w��ZcrX���]�1���%P}�~��e�Ǵ\�		�(Y�S ���<��:�bX2Ҍ!���yV2���ՠv�������	��yӀ ��xT6�!`�*Y�:)�E�:TGfH0(����%���p=�$�C��f�tbB6����eb|�A�� -2@��Ȁ<_�7m.b7&����Dl>��c�1��&Â�]�B�8ز��a�������a�)��}�!O�(�&���͊?V�a��C?�α���.���`T2�"X�/��{�N�2��:N�1�=�̵��mD/��A�W����D�K�b��58��:yّ������*{eFP�t�3i� �����=m����,E&�V�9rc�=X�8�c���g�T�0rjD 1Nգ�o�9BtNA��E	��O��;F�@=A�P�{��=��Yy��O�bG�#4��?�Q�Iܖaf��v��=C�^�3��9��MQ�=gN���b�o��l�D'O0J���S$�%�����-�OJH��L��	� ;��O�7|hu�VŇK�=���35g��j�7mAZPؤLP� +���(1wz]��4�%,Ž!�h�j�f��cc���'�hf{�l����,d������F����a�&�rs,��[.6-��gH(�A�l��S`��kRo���a!V$C�1�fe5F�O��bো�&jX+P�K�A��)hV�ɺ��De�N�d;Z�����a�p�Pl�U	��"�A��d򕫂�)�
%��J�z(n�yM$Z�2����X���ׂF\�'�!:3mJ�]�6�Kl
Լ�2�`Z#0۲X��B<�� �mJ�%�c
6^�"�#���ܨ�J@� 5(ݨ2"�8=��mj�G����I�v!�/+��˓�'�����_�1�*��Կr����$)�x��Q3��4H�7(��N�����4Ko�Q�qfêz�	C9�8��,� 6�
]J�Nq�fuV�' ~�3���2TC�TV���F���`1hE�G�NST� ̈́
3��$a�Wvr
���E���\�`��c4nQ!W�H^�h�%4�L�JUmߓPFfd�FGո�O�2�)�Ncz� %꛼#���`�Ϩu�}�􆁯6�XLh��1��#2lU���3h��0uN1cѨγ'�Fuip� �0��PyU���ؙ�'�3r�v�d&O�V�d%p�	�,t�cnֳKl�t9%
�����R���t�b�	(U�8E��ѻW56`�5�
7̞Q�e�)D�kE�'SR�ѝE��ɒ�3X�aC�� �%�
�9��/ar�!Å5#Y @��ПB����FV�7P�y{�w�NRF����aH�� +'Lə	�L���E�7��}��b��~�PP Co����5ƴ[ �I���U*ĩf�XJtd땂\}��t �@k�����O"�Jb -jxU�4oL,2v�(x� �iܓ;m�` i��bEàK��}kr��sf@��\❏-�����<y��yȔ̆�B'�٨PY	Y���7j�O�j@"��$��n�{� Y! ��R��Z'5h>��Ӎ�6��2��wn�Q#���<�r�s �"��j�fZ%0c$��c��5��}:���jB\�:���)�҄�o\g�'.Ѐvd-apP�bZ�8�A�Z1�Z� ��W�y@⣌ ��%���Z��A%݄#<����۳�V���R�YB�m��I�/�s 
5���2!N�"�<!�$�8Ƙ 5L��%u"}����-(?�1�F'
�r�q��]�5lj4�"#�"r�`h�������cf,5�zǮǥ�h�)1��1dd�	�' ��)��:��8R�mH5l(ȀBb���~r���nD�A�6��"�ǟOJ����6gDan�l�Z$a�"�N=��	�$>g�I���b%
���T&U�#&_�hڱOKR?
֤�*�'Qc�M1a��hAh��O�Wv�p�]��T�Ѷd>t��ӏa�qq�JE�kHx�s!��R~%�+Ť_ܶa��)�&�Pzd�3b�^X��-[f�\,&ϥM�1I�#"�\bt(3c�X��4C��xb| k"b�`�� �
�J:"��G�N�rT�٢,,@����	6��qi�E�����/p<���)B�|���㆙�0�ʀp񅝀��D^�5�l�鄦�*� �$a�>s���Y�lW�JgB��	E�Iy0H�
�^mr�C�#�ܖ-{��h�$��x�*��N�Jj����E@@p�w�S�p�,�4�@-��l�[�|��'ꆕ]X̴�A(̿pKN�*W�{�hH��E����{gd�?�5
/)m�� Ħ�:&��rUK@�WH���Ϛ4dX�fÏ�6y��@E?j��e���ԣm<��03�QB��<!���[X��?V�)�+Avj�B�pG��Z珂�E�������GE>Hp���(u�<L	�
.Et�;	�	�ªܽ��qSMC1nIqẻ�jhX�Ia�_�@�$�H!�6�	4A�(� �×�R̎x�����a[$G:��xr�Ƅ/�6��MO�}z�����ud\�B��S����qA�����@&�,�&�!эxp��� 0�k0�ˇWR�U`E�f ��5P����
P�"S��Y-��!(`�B)
��b0� �R�� "Ā���� @�*0�E*H�@8�dr M:|f�0Hj��_��DhT#ʧ"���K A�"$�5ʈ�C=�h2�i��э@�r�4���!ɥy/�U9D`�� �	�8|�h���F�Ӧt�<<�T�D>/��&�e��,���ىt�r�{�m��1Sh�y�#Y���(�n;3� ,A����d��4�=��#M�^KVt �BՅ�n��6�Ug@�RRd�P(^M`p�o+L��$A) MZ`����l���b��eF�RB��U�ʍ��gۡ=c�M�"�@��x��]:+v�	�[�b���hsV�\�@b�;�J�*'n�=;Q�P g�FU����N�..I>�ۣ7wb�qtň��������9R��}K|uaB
»8��Ӧˢ�t�5�l$�2(�� �F�'j��P���C�Ҥ�ٕ}�zm��ُ`\ɘ)������\�z�X���V�`s����n���GJՈ9d�I�V�V��#}�w��9��96[�D",�:b���+�Kq�Pt��I���,��M�~*fi���y��I�P�����ߙN����K�H>�l�!��i����`�]� ��ψO�q �m�4c��4cV�[�����q���ٳ؄Ƞ�̟���s��a�Y�t��y���=h�)F�� N��q�`�*m~،�����=Y��3r���O;�@���P'>��P֏�+���{�/$��V�*���s�ı~)
q&?�م��b��낦Ѭ.�Q���(���+�G�6�`}�O?!Р�0��v��$9�~��C'D��0�>d��Ha�6�3�j�<�I�P�
���,}��	�4'��ؐJ�K0����@	Dr!�d�q�>h�5B0��tÖ�I�qO�e[�d�
�0<Y��T�C.���'
��S& Rp�<q�n��c��E�6���?��L#R*�r�<��/Gvs6����y�)�J�m�<���ՅdAV�����6$.8+D��d�<90
�q�LВb��:�E�f�c�<�-O�T��.��=/2���#t�<�B`�!��	EA�VF�+�#p�<��h��!���p��S�))(�vG]m�<yS��3J�|��eS�FE�T �@�S�<pL�eF*0�+2G~
��㧅I�<���	�EP8���T�]�LACE �J�<醇=2"~�0�)��P�a;���^�<)TK�-O�v��$Ϊe�����Y�<y�50��ȩ�铩\��&b�P�<�Wj�h��<����'1$�����g�<Q���NRbi��4ɂ�Q�a�T�<��ձ.�-[Tc�|ih)qPK�I�<���,#�̰`%ώn_�bd��@�<CO��Gz��W�ӉY��@�1�F�<�de@(?�`��!��_֕	�C�A�<ArkI�*YH��r�K0II� '�t�<1��Y�yvE�����T��~�<AB+�k�~p�!�>�RL)�L�s�<٠�A���Y0��2O�ݳw͝h�<�'�ZqX@�!/��L����gMk�<��Z@,�
f����2 �x�<�'�V<I
p�RR�V�j��T#�O�u�<�$�W��r���F@��Y��v�<y3��;M$�[�LF�}Vty��Bn�<y�%9g��	�$�*3vP�L�<Ar�E�(��U��J���X�I�<�â2��4!pf��V��t��k�@�<I0�C�/�̉᧨����)FB�U�<)�R%i�݈a�	���{&?D��"`�p���s)�6@�X�4�<D�����L={�>��3̈��lD�B�8D��a
Rr�h��7j$,�� �6D���	�xxD� t��?���2�2D�t��j�@\9V`��J���huM:D���A`X�;d5��+J�f��܋T";D���$Gj��1X�a��Q#�KRG$D�3!��-w4(jҫ��-}8q��+"D�<ÂB]�74�00�F*��e�7D����V�D��r� TT!,�9�&5D�J"�>���R�ԗ�{�A6D�� 4`Z�'��%H>w\���"OΈ�eI[�u���R'�	Jn�x��O��ˤ�: Nr�O�>����<����"՟m�V�b�)'D��Q#i
*�fp����G>|�2®<��!ʶOK�(�	K��0<��' y��P�@�i�b1�/cX��r 
�D:i�k�s��d(���5�r�"'Dӻ%���+�';�9BG�J
k���>G����ߟo?�2�9L s��;��ra�J�7;��c�L��Cg!�ěM����!e�yPf��7mȼAɔ�Z-Z69Їe׾Z��򧈟�� h"��q%a�):���tD�?�y�\��K�0/����HH'{���`$�~(��BO�)��\�G���|F|�B0GL]���,1��XB��*��O( c�����y��$7������C�B�64�Bb��`ࢱ�X�#3���OB�)!0���oXt9�� +ClL���G�D��ŗ����F��M[S#^	;�<���BP3\�İ4�3b��Z�M��p��͞����I�!�yBI�u����%����Bá�� V��b�ΊX^ɘQ� �5�5��N�����lp��p����ㆫ��}ȃ,W5
�$�"#�ɚD� ��)��G8L|0I��F�ΤrgÖ�4Ḵ�� ǧD�Qc�4T�j̊f�P�А��I�i���Ex"m�?3��X�Ƚ<5�<�%g�V�5�!��Dӎ�'�<�alY @۞��#�΢Zp�V�M���H�!l�x5�M��39"����W-O_(�P��VBڢm�?!b([5ObxPZe'�/��)/�N�Y�%Q�k����\�\����O�qQ͸ F؟o��ٕ��(+�Z�	'e�
l���џ�O�k�����6S���LZ��V�|����-L	m�h�
�'EЖ��7-� r��}1�CJ�c�$�Z$�~��0"��q0��b��|��!v��QQw�g�,�B$-I�#�����%�Bh�ЄɈ�<���b
�z?Qs�ON,řE%����'�8-��'�RK^ag�֡{c�I`�R/h���o��x�b	��Q�$�فbֻ8�����KV�{b�IR�y��{�p-����> �����V%
��	�pg^/E%��C"o	a��Ix��`�H?#t�A��B�qC2й���1����paD�I�lɒ�J�i���`��F��$l֭�d�ƇJ�����	M�z��@j �jz��i�Q�Ė0U�"���+�yC�]9bLC� KjkhS�~���ʷ��"ěd	�`�I
7��_��s��0�*�qҢ���I]�Y�,�GK���M� �Z5X$��k�b�j7=��A�BJ�v.h�S�l��y'EO�2��x��Q�!���"*X�)Pb���MbB!N�*�����O��l9@�P$'三�*,Z�k�P5&`EQ�F��'�2A w��M���,(�丂��$���#/٠i<J�w�2����?b���`5 �,�>Qb�	�U%�K@4R��rH>A5�E�Q��"���%�Dye�1V^\c��\�x� ��^�%�H�0�4�`�2@�t��9�(O~����A�=�M�wlÈ'�>���c��zΎ-	ŉ_�5˴����	��x��Wl�V��q��H��[�[���Do�d[��w��x6Hp�"XkLH�|z�o_ e��EQ�k÷R�~��4�������[����%�]>o�̤�f�0<��ŉE��
Y�����(��ksT=��/�����U�ܼj�֐򶧕28���ɣ ���05���n�8���ɶh���D�k�BU3G�N4+K�I��yb��(C�y�D��]F�IY"�N��Bq�eN&p� �`�D[� �����^�@@B�ÎeJ�iJ�����]�̚d�b�J�M$tY��ʌ	��10׮�h��������j��В�@���@���w�R��F��I�d ���v�������CH�a���
Q�x�Lΐ
�>E"�<8q�dl����Y_$0`�I&�j}�Dg&y�N%�E�� 熬0�,�N~|\�lԢ_T0 Ү�����w49Ku�A9Q�> �֮�e�����T%���o��ҧ��R]+F� ),l���7F����̜6d\ �q"Å:���r3d��\����� -&p�s͍.2K���%�O�����X�:�Q�뒯Xf���>��W%^� b��}{�*��͎�0�<
f�:Ov&�1N�W(dk��
#g�����'��@��!C�cT�$j��I�!6�p ���6R���"ޏ>���c!oU����A�N�ƈ�A�׿�n�a�E���F�:�NR!jb�^�r�h����7GF���	�  :w �?4�Ź�װ_�bM�P�w�A��#^{f9���W��MԎ�)uzȻ#AN/a�ɺ�wD�ɰ�)ʴ/�d�S�ٙe��+�'{�=�sjK� 6�8S��Nb	�vg =��\PK34K�E���2j{�-�j
�<�#$��Kv%���'��z�77�,��b�,rw��BӓQ@pqEO׻=�f���Ա=��IsJ�-ӛu�X;b���AҸ$gX��"�Z:K��&��s,�SR퉂t�T-#�i�?W3���%��3�Db���Aŋ�6�^ 	԰a�H�3�#,X�cE r�N}(��o�ִ@�I�E��L �f�����͋��>�u	��bX���$��Bg��`c�P_�،QV�YIx�i��
1N��	�dU�%DFo��hCD�߼���G���D���A ;�H��X�<!�
1�V�3f���& ا �%_���
�9cJ��h�|�P)%�	5�@0����,<�kA#R���*l+�@� ������#K��Җ 
	�b�B��������)��T:5�G��,N��k�Z,�����a�a1����#���
�)мWg.�P� �e�r�R�	�.��Gz)�$ٲ��%
��iV��X�I�6I:���^�fԂFŐ/|.����$L,�}+�+U_ݰ$�u/D1�0��st�M9g�OQ~ȋ�Ϟ;?Y�Z�g�y��4�I�(<��Ҽu{�d䎏�.%�q!��ٲa�0i�ǎ�7k�T$adB�ք�7~�T�n�@(�e9شc̎A���l�ȥP�D�/ X=!&D:Stf%:U ^�-�$��В|B`��/�(���b�aE(�5��Q ���B�B�	.\91d�ɲ�� �]���Co�
2��� L�?"��!��;7���@3A�ʺ��p"����#�؈6��m:� ��Y�G�9h�d���ȼT� T�A��at��N�����{�oC&W�i�'�i�n�@H�=V�,P�!dx6+$'ȄS���F�H"b�¨ �JðDy�lx�Icp�<F+��:k�')�Fx2,+�	�%H�`&�1xLIx��14�0�1�AEqn�-�!�f <4iҝ!T� ���OPqhv�3������p�"���M,z�>�;��@��
��c�Q��#V)�$dt�[7��2aTx��ͽy��;3+ ������T(���.��6��E �
.l1�>~��<KëY�!����f�P ��Ӈ�� '�T�G�ɴ	:8����$�ēh~lx���,O��{4�X ��ٖ!FE]*�ڔ�K�BFz�+��͏zz~��b]�S�ԈĎ�����/�F�sA
\���ъ�*����R1?���A�OᡄI�/+���b�lߨ�,P�M���*ab,'N�f�KL�����."��z"�iڨ���w��݉�J��~,`T��@�Ff~�S�
��K��bǧX]xt�8�£>�Djޭz��i���-�zS��%������ta����^�,�7�1Fa����/J;Ǜ�g	�j�36Kȑ^�f	�BcC`�i8�H!��<6%F� ɖ���PD_r%Ybk�&"��U;
�ldB䧈
��=���C_Τ�� ƦC|��0�\�'8����'�fxD'ɍ������H���z%�<5�,�Hs'R0H'�'k�Ib���e�Z�S��4�*�ϕ�6�>��S�K"��ɔ��H�2p�� �-ұ�V�7YAynڇ�PA��O��V+��J�LI�P�ɀ'Zb���R��O5ޅ���{�ܠ�!$Ũ,퐡��c\�%��Wk͈LL��2�x9�an��E �ۥƅ�".,0z�j��vȗ aElZ0������h�j!X��'R�y�($h4�L���� w�̵� ˋ('�Q�fK~��)27	܊����q�_�j1�P�׌�"r�¡l�W<J��d�D��9�G_=<�����e�4������$�۱C��'��OPF����B;~�$��п)E���$���G�� k�MRD���'P�h�����t��!�X��@�A��$.ކ$(r�҈��'B�`�D
K��rt�"y�D�
�B�� �-{�J8j��^��rQ�#�|����7�i�~O�-Z�^5��B�)ܸ'n�� � O�tBf-��UH�ˊ �MȄ�G�f��hSeA�1o��]�}4i��Y4;�\MX l�����Ɠm̢��2b�%C���:�h,�
�-'�U:���! _���dRɒ�rK	77���R�H�I�ZN��A%���]�dx�é�?�Ŵi�����	Jry8����ebF�1\vL4
'I��i�0��kf��L /Ś0Nn��*�;G����7e1�����,�!���K��_�yR�6Ɠ}��A�>v���Sq��!c0y��G�ywm��f֤�AL��4>�v����>	V�Q�=�@�Z��!LM�����R��:@!/!�&(�T�ɋ�,I��m� �<�"���IA���Aj�8Xa����y���#������!���z���HO�]X�G�A�B���Qvw|���u~�q��J.y��T� ��`��9h��\g����ˊ_f8毙�r��9@��Kl�'ef0�fL�L��\Z3�K �>�HTFր2k���d�
$6k�4
�O��Amh(�&LN��x
��
"�4�`$f6���r���nx<���h�"��z�/c� ����'af9P�E��,H�զA#`Xu���W T�mؑ���\mL(B��ij%h@%�&@��f �&iLY��w8D��ًctT\S��P�� Gx����6y�D 
3 ]pb�̪Gdb`�$��J��iMȩeH͏j�^d*���j0h�p�]W����V	')�b�+��P立 u`��V�"�O�}ki�8]> c����$X'�_5@�\`��� ��C�U�XͲ��.k�.ts!�C�:�J���J�_��$�F胶>�=9DL@�qp؝2�h�-u"�s��ĢB�XX�眪���
����B�Vb�L�ssҁr@��s/�34N�E�p��&��^h.`J��	)yv�zehA�?`�!��F¦��>qAf׉4��Âɟx�ڈb�L�&ih�8�ʀ�*��б�)fɠa2���ʦ��%��=�f�L���y���L�x�"���#������0>�u��\�n�"4 �<�θz&-J�Rg�./�fe�Ï�+f׬�ɀ�Q�r?XԊZ,͉���o\�L uhл%zY����ܟd��&�J4���#��a��,1,Y�=���8<2�D�'�MD�2��#N�иև�O��H�gǼYh.�ґc�fs&���J�0qf����-1F�Qv�Q�'��T�F	X�V��*�L�c*,:��Ll���;*\�w��z6b@�F��H�&�8U��1B�a������xg����ȝ$ϒd�G9ndܺ'�}�a~�O�90���$��3/�p��q��/���C�!�
L���B.����Q�"/��5ର��0)�dԐ��'�yw/�-g\��d�#�|�aaV8�p>��i�[�>��+�|yB|@c�5�V��HK�S�^�g��!:P�q΄����pE��<~L`xrc�7�B,��苊��D�O����h�uF�����0,6]�=I�%ؖ�$l�d�D�F�����6 T�Y� 郥Nܐl��c۬b�f�'�=���ɴ;0��z6�{��)I�ِ��O�D�C^�$�p�����i"�dω$��Y�
8\\X�V���J���ߒ#�`��u 5j%�J�Ď
"��9i�L�s����"��=T)���`#�l��D}�J�;/W��k�	�7��)x�0��A�7H�L��Ė�2��� nHۄ!H&+�FX��jS�}����6I�@�����$睨k����%Ƃf�r�Sr�ľ^#�˓	��1�	 �p�h�:�'PԚ��g�Ux~�*�����I��h�}��a�'�2}��1q��y�*���nߛSuh�rs'̜��a�W�����0�v��u7��c���7�2Ty����q%�ؚ��ͧxmp���J�P_��IQ� �S���	�5
��q�b��,f�Zl�WJ���@�����(�2����{��Y@	Lt�/GD:�-Q>L��ݳ�!�3F��J�F�	5 ͓�*ٿ~=Ctj �!R~8��3����a���B��R%��9�Ӵ*ɕ�� :$�)AuDݲ�d��@��H!"B��DptF�%jX9�ʗ�&��< �D�G�6�5O�GZ @8�#Lv��9kR^�FA*d��%l8ʴ�˞�&��O�CR0`xrR�N|��a�ӎZ�>Hc���oG2��q�E=����Opq�I� ��1ň��L��@A�6!������?u�`-�c��9�(��9�4TҔጓ$F<XP6�@�c�4�3/�N�4!��Cg��i&( :� x�DAM�!N2Lx޴
,�q��#�-�p�����}5D��`bڶ9t��_�2����Ux¡@�D�F�
t�L<��}8q�:� `L��Vt��T��#S�?�ܺWc�Y�f� 'k�'>5&a���.~?th�e�O�<~t��H��`�q��n,Lb7�8^My�-�%~�99��@$q�p�c���e� q�'��-�]0�Nd��5#���qV��2������-Z��|XR+b-�U1��ܞ`+�qas�M<;�xĊ�(�&��ɩ�%ӇIzU�Rf�q6ع�%/ZV*MX��+mv�Zc*Z�Y���Ffm����t>ԥ�E��S ]�VdP������!^�c�TXr��A}�ߖ�J9k��J�@3bh�E[�M���Գ`/*=�Ot�"��Xg��h6��#8��X�EѮw� �������UH��.۴]a��D�!f�1�#��Y�2���G���%тp���tn�=g��I%-*U5(�!��I�2좓�R�����?I����32���Y�#�!���k$� �A�Ɨ;��X�!]0@����2|X�H^P'�1�%aCT���`mE8h�-�o�/f��;de���[1��z ��� ��6�e�e���%��`>m��A3O^<Zd#�Λ1	D��p�^�Ș@OISp1�ई�T+2�i�}�c�NV׍��L�d�1	E��p�lM4#�Yd Jh���{SOR�1��d�`�јD�ЈF/
�5�*�X�,m݅ �fpɓa���	Ѳb�L�C�jG$)��ǟ)��	֊DJ��O?R%B��f�h���͉&&8���O�Y��1t���D_&�KT.�$L^�T)S��/M�iQ�!1E�>!�;�Ȣg"~�R�/I-�Flxp�i�ȭx#�N#P ��eSɦc?!��)DƼ�У�k�ʷ � V��/�>>Y����[�$B5���"�(��g�'�����!ZW@�P�A��J�aY��~""�;,
8�� �C�9O<`������W�P'��2k��ȒF�F�%�U?Ua{"+۹f�.��v �p���"�L0f.�@�e/h ��1��M�I�h��!���-`� ;H~�d�+]u|@ NN�BU��j�h�'�\劣@C�sw����~�7+�
"�I*ċ�i��r��	A�<1�$�3M�GQ
b�1C�ty"�_�D*��B�Ll��S�z�1��C=(	�9R�kÓV��B�	�L7�e�H�Ղ�`\�r1��DIn�9Xax��ٕ|P0G��U�
��7�G��y�e�8ohmP�ήJQ�ZրY6�yb� 3:��� �=s���9�$���y�-�5.5��7^��jb-Z��y���
��h�#�!X�М��`F�y2ㆄP��I1E�G����'��-�y��M��m �G\�;�x�X�ǒ��y,Z�g���!��Z��в�-��y��0?� �V&eޔu#�,���y�d��	WR��'��X!��(����y�f��o(��*rOW�P��T�$���y�O!M�\�A2f��8�l���	1�y2�<'��h��T2��u�A��y"8�s2�2'��	d�΂�yR��k��h��+̠�À��yr��7��B�W�t4� ���ȝ�y2A�-���3��=�,��pNM��y�NʅK�n��_�8H��� ��y2��8���qw��	�L�k�/A�y���[����doؓ�j}�C-�&�yRDȯb |��m �p[��#Æ��yr)�"MB�a�^#{�h�s��#�y��A Z�P���d܇&y�!{ C���yB�͖b~0��-'蕃�I�y�H_	f�s����X�2I��0?�T�C��t���&A��2����{��R�GܓR[-�Q��w��1R-�1Uq��ٰ�
�	�� .G�a��$J� ��ı�4A��  �D�����$N���т������h

�H�4%R�c"5��Pm!�d�A����:T��KȚ+S�8a�NV�8�Љ#}Ҫ=�%��蝔1���3�*T�@�p�������'��&�)�IƗ2�qe��M���t*ܞ]��'$�LGy��d�B�y�TA3D�T
n�H�t"'��$ڡ�(O�>͢!�ԀLO�D��o�h�����bӦ������J�%+��,	�e�>sR@���^)lP�*��>�v�O�$�k!��U�2�I%��..���@�k�9��USs������0|��DB5�n���)B�5Ub	y�!�{O&�X�8O �RC�����Op>0�֌]]�� E��Q���C#h����ŪQ�P�)�'R�H�P�耮qP�%���E��4(�����O8�a����d��.h��Tz�DΗ>���2�,�zw슖;O�6�R[G�KE�~֧�S�P����KD"��
SDC�A��`�>��@���0|�$���u����~I���bN�~H����'N����3� Z��Ȏ!#r}�3��+Q����O��'�FO��a�S2Lf�����+:��T�T�C�%�t�OZչL<E�4g�%l;Də7f4��Չ��y��v��S�|�a���$}�"5���H������Ҟe.�OpE�ߴKz�c�b>� �$�KJ���h�pe;b�3?�)qӢ�ʍy��)�<k@�ӱ!�K���@�ƾX��$�������56����d]`Þ�$'�>O,R�xL���y
�'��0���2p.���N��: (��
JS?yQ-w��	��?UH�LY���C��?��W$ N��a���y?�)��?,�!�y?J�X�܀ܑ�*D|!�DI+u.�:�	CJ'��*���!�d0s���c��~�x".ϊ�!��F��@ڴ��[�(�B�g!򄍯|�1����
��@��(��W�!� I�>$�V��|��e(Ua���!�D��9:`q���ɯkm�]2� ��^�!�®9����h 26.Ec��BC�!��R�v����,d�f8#��Y� �!�d��>"�Y� $1&V�C��Ճ5�!򤜯
*X۳��#K����Sn^��!���%B�t+��>�Й��l��g�!��S�7�z�ݝF�P=�U�ѩq�!�D>d���	(Ԅ�*&�499!�d�ti�eKɹu�&���YK+!��[,Q�d�g�2@������<m{!�d	,J����#�`�(�,Uo!��'��ňE�_�qe*�������!�d�:M*��T<	�T<0 � �l�!�$>}�	�C��*g�a`#ň�`�!�d�/&��Yba�5w�j(�)H8!!���-��QX�!Q;)��A1� ad!�$Ö`z���j�3���v�Ʊg_!�D�:l
��U�0Gl����^aN!��u�jʖ�R�cX��P O�Ge!���#"�f�����HF$Mz�����!�$ �AG ���S�:�\���3t�!�� �J�`b�ϯ1�.u�Kߓ�!�R�rW`��6 W�{2P@�ˈ�L�!�6K]�V�z<��K
�!��w:��R�DU�W�\(([Q!��	EG�E���	Cܔ�
�A��!��$:���Aճk����c�"!��8Bք\��T�`&/!Y!�D��2��D�c�ZN�� xU�I%�!�$GiC���&��u#��;�"K�8�!�D	�T+,�` ��d�����x!�&4��p�#�	G�`d��nžl�!� *� 
Q	�(<H�%�՛'�!�Dطt[\\(��(K-�������l�!��9���!�ʎLy���ܡ@!�D�'N�0$�?Ll�A
��_)!��y�� ��?*�y8�ǃ0a!�d�"&�ڦJ��\B���C'}�!�d�5ta�gM`*��(C"�hz!�d�6:�´�ׅى�(|��N>�!�$A�V~�,B�JϗO��	���w�!��3vf�8�A��yvp	P���0c�!�����S1M�)F���B�aW�l!��F:k��(1e�P�4�"4[!�M�pM!�$���IP�F	}�\)Ҁ�C�!��b���i�l�(L�~���g�>�!��#F���I0�	�4Y��2(�"V�!�D��z���eoݡ��Vd�'�!�dE��tJ�b)���!eb2*�!�� Xlu�>B��s��B �i"O�e��BQ�|�h5T�ͅZ�`�"O�:���=/��r�B?P_�-�a"O(��íW�d9d�#5���ib"O�8��Lj��*0������"O���f[	��I�7�TbZ򤺂"O,CT��g
@(�#[="	�"O����cP�o�(���%J$#�� �"Ofu�b�X3V"�`QS*Up���"O���/�8dr�5�U��+� *�"O�t�b�йtPB5�T�+	�mI"O�M��C�d<f�+�4�8X�q"O�L(`,�(f��KN�}�JՃq"O��zb^�o�pP[�*�$P����"OV�۲Nʏ��  �)�Q� ��"Of�rĝ0A�0�r�°�^l�w"O��H�E�xA�i=.R���"O� :�l�6��x�i�1�റu"O�HV+C��00��QE�� 3"O^ah�E�yU8u�'��`?z��0"O� 93��kh&�8�F��)�<ؔ"O�M�WBM�W$2(��/E��蠤"O���%(�e��k�n8��Yٴ"O6]3"֎�N�sH3㔡h�"O�%�sCõ+]��`�(�^� F"O Pbș^έ�`��[Į|Q�"OPzs��k�A(�M�AS�"ON`P.�;8)�f��Y�V��"Ov��S�X�"U,	;��8�t `�"O4���.Ο3|����"�(�"O�{F��ry��+��ȞK��XB�"Ob5g�	�L[��X�6�
�#g"OFpA5��eʤ�g4�����"O ��4'�(j���Xæ�K��a�d"Obu�c�� ����gڶ^�z��*O2YЖ�Ӛ<)�E���+]1ޅ��'������"m>���	K
@�6!�
�'��A��`]q���D��7�% �'߬s�M�֘�(݈;�r� �'H���ƍ��%�E	 b���'�؈b�\'W2	#��� .t=��'A8a�!g<Kb�Di�r�	�'2�@`��v��	`ǝ�#��!#	�'	���6��3[CD�;�L- +�I��bN�Ű�a�a ��άH9XI�"O�����5R����d��֝"O������J�R�Xc_�Y,a9�"O�C���P�J��!I2"�ʄ��"O�-H��
:	�.��f��h>h��r"O8-�u&Y�O�x,0r`�����c"O��zWG"��a �bx���4"OJ���>C��	Z�E7QA^؀�"O$$�3K[P�AF΁	�A01"O��0Q)�M�J��r�R?vSz�Ӡ"OX���P肝���	L5���"O ��&�{��H�F�X)5X��"O ����9.���z�c1PP�i "OF)3u/� J�(@�oR,J0["O��)`*G�����-02�٫"Op��(PL[F0�-:��4(�"O\D@�E�9x%�kl�T츍J�"OJ����6?�$�	(�FX�5"Of��B�W���æ��t�N�"OT�r�]1�|�c�dV�v]�	�"O� .�j2Ȃ"�z�`b�>�՚�"O��#Ӆ��l��U+��!Hx��"O��q���2(���@�>5/����"O��+�������%o[� .��g"O��S�O;lY�8b�=_����"OX���BRv�n$�k�+*(-�"O������8H��e�B낈�L��"OL��EĘ�H=�	�'��e	&�E"O��B��],N�\9h��$h�t@h7"OHՁ��r�܁`�T�A�>�Hc"OXA
�$�=����c(��A� �)�"O2ث#��7/(0ِ�2��z�"Otq�h� *�L�U�@h'�La�"O)X�+���qRN،���q"OpUP�.ҝ9���Ҳ,\�r�(���"O4剂nΏN�~�I6)R��:��"Od����ޭ%����(M:D��,�&"O,L�̝=�������\��K�"O�
#���V!�"���"O�x:Cj��a��낄V�B�� ��"O:�[G��Q@��0*@bX݉�"OLpR��d��8��H-_7̘�4"O�8S� �&�#���r$ftA�"Od�X!	C����A3�ۡ!$:�H"O:@�6@C"�}a6ƞ���"Oވk�/	�GkB ���7w��B�"O�����@�	�x`�T鏟?$q`t"O6���gV~;ɚEc!�LE�"O�,��˺�<m��\�*�L@�"Oބ���R���D1g��<�B�qv"O*if�B�pVx@��cF�4�sB"O����B(�c���|q��"Ol1*�(�m��m(��� ��h�G"O�ٻN!4��[�dG9�� r"O��6eӊ?����)�� ��Xф"O��WGV�(OD���a���aY�"O��jբ9 Z�ʀǋ;�$d�'"OH�(wc�"���FG�O�(�'"O���3�\1a5Rac���SC�Yb"O�e�u荗L΀@S�^%V:�Z"O��P�#��v���c�F2*�H)�"O�-A��ʈT�:��G�t� ��"OB�cb�k@�D��y��+"O���=V��Eȶ坦#;X��S"O��戲�
�	c*tѱm��P�!���1\�`� )���Ye�-~!�Ğ���:V*-+��
��ـD!�ā/������B�f�r����%�!��O�x���a�b�Z�S�^�%�!�$Q19G��(`!��@�~�ɕ�J7�!�d�*B!�\�!M�lP��G�ǃ'!�d :<��Y12N�F��*��}$!�D߭�����(�R@�p&�<`!��!t���gH=q��pѥ�28�!�̙-�	W���
a��K�8�!�6-(��]�T9�!��$˪,�!�D�8,i��)Ӡ�X/⁸R�@�*!�F$���󠪎���0��Ⓓ[!�d��@@G_�O��9�U�f�!��̚s���ذ���5�@��'��!���0~
���V�R#w�,���A=L�!�#a�Ћ�bP�S�X�nU��!���f������F����k�(!s!�ę�d�6�AE�K?-R� E,��5Y!�� �1!FFI-<`Lm��çPϖ��"O�lj��ϊy!�
X<,��0p�"Ol����M�ڐY�J�3�^��4"O���+X�_j� g�Z�Y�<���"O�1y�l!:f���CB@�1�"OhTrB����L��aT�j��@��"Or\rU�ˑGp����N��ز�"OT��pn�J�4�+dDű:@D�R2"O��r��.��ys��!V2@iʐ"O���Q��o��ܡ2"��*����"O4��.)|&&�E1�� "O�(��T�ҸMc�HB�Xa�A"O0���`� Ґ�qЍ�2V�2"O��2   ��   �  F  �  �  �*  �6  fB  M  0U  >\  �b  �h  o  Uu  �{  ہ  2�  ��  I�  ��  ̡  �  Q�  ��  ٺ  �  e�  ��  �  ��  ��  ��  �  �  V O	 � �   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R��I^>�Z�l�)N�HI��S�6�CJ.D�Lh!Nġ ٳ�fݒ!�҉��,��T�I̓L��@|� ]	r"O<��w�R9{&m�7 �)Aj��P䘟�F{��i.[�����N�&�6��Х�}�!��U��0C�/��10.�`��s����<��-�|����G�� 3�iC�ą�IH��?�������O�3: � � D�<�%L���.�����%*4�U����h���� ��#��]C��5'�.��"O�у1mF�1�dIU��'i艂��O>�=E��܆5�>=��ҡtN�pH���y�mX�~�vu�g��G491ŮK��yR"�0A��٧�K�E9(ʡCI��yb��!G��p�$��i�^����P�y�eɯ0�<Y�(LO0P�3��P�y2,ئ ȷ�ɼE.x9u�yB�G�6�vy�*˰Q����	٨�y���TN>aJ�������"�!�y2+�e��[����,�ű�hV&�Py��G3h  i"��yD�RAXv�<AU��{1��s�-�P(�A�t�<�4 �xA�!A���O�hH�V �n�<�6J_�\~������Q�W��t�<1@�]�)p�bI؈k�FE�F+r�<Y�[.i�T�9Q%@+||����.�U�<�1��i4�T-�dym����v�<�`b�� �����*�K�y�<0��7qz��ekM y�p�#�N�K�<��:g�����+J#^��)�a.[F�<���ׁR��!�jI�\H4!x�<Qb�ݟ]z��۠�ۙ	H�P��w�<���f[�%!j�?���cl�<����E��iH�
�(fU��Ti�<	�!]�hRU����, ;�N
J�<��ÿ[�F�:a�#u.�G�D�<Y�l�&w��J"ٝL�H���A�~�<��M��(P�\�*�1&����/ZT�<)�����L
!*5c��q��N�<�S�]9�Xt��+F�yFiSH�<��E��y�t�׆*	Y(L�É�M�<1RB�VrȲ�.]�L,�`��N�<�Iƽ2����C�#�^Q�H�M�<��jr�, ش��uX|<�)�]�<��#,�<��嬌�roܵ�u%�Z�<Y��V�-5�i��Z�Ҳl	BœV�<q��2 �d�k���T���[��O�<	�+��>e#f	ڽ��z�L�<\�"C�|�AE��5�F�n�<Q0�|���`��T�*�����@h�<9�.K$.0�hV �BW�1ؔ�m�<��L�*������Y(i��j�<�A�s�"ء�ɐodA0��d�<� ��*c� m����T��+�I�j�<��m6$�4���6�F(�vȔM�<Ʉ�ɃRԀ��DO�����j�p�<�U�ǣ0����Y\!T�����b�<�6E�)b��m��$��H�#_x�<!�Ə/Y��j��@2`f��2D�v�<�F���PD'�-?��dX�
w�<	���%&TKw�Z2G5�Y���s�<y�Ņ;ra�i���­-,�*Ԍ�E�<� ���vcV*w�Mkf�G�<:eY "OXU�B����4\�ǭ�M 
}��"O�T;UaN�I��q� �R�D�B��r"Ox,BKW��X��
M(����"O�쒅D������!�����"O�YAd%ϥ^ jY;IGJt: K"OlDx�Ҍ[�<�8e�M�@\# "O� ���@*`���I�?UM��8�"O�E+��	7z�y��K�>M�A2"O�ڠ��>t5>l�4FȲY1
dx�"OVT���H�p���#� �I���"O�!�"�~��)[U$����C�"O0���Р0��ϟ
��:E"OF-�c��p\�娥�=R��(��"OH85�N�n"���&�Lk>�A�"OlmP�j��i@�d��*d^�j6"O����(G��@����.R��2�"O�qKeđ,����n4��`�"O8dbElًf��0���N	0�Ā�"O�ubQA�7��}؇˔�_/X]�!"O�쳲��@�D�/)�4�*"-��yR�ùF-,x@@�!7�,������y������1Q*a{��4�y�MS��H����V�~Ё�1�y�i��+<!��\��|q�/P�y҆� V��(�r����ƙ��ѽ�yR��q;���B�܄��͉AѴ�y�珳Y�H�Ҁ-E
�B-xQ�7�yb���p��U��\�9&�{���!�y�O��r�:vj˕ 1"!��j��yr���P��F�F�yA�-�gV �y�#S=V��a[��9r@:��g%�$�y"���!�֔��ϫ6����	�>�y���k���״0����K-�y2	]���`Ɗ]�T�2�A�m��yB��4�4�;�ǊNhy��8�y���>^}��8�[B��ųt���y�l	S��ئ�McꚀ$���yBb���8��۪W�؊t���yBʇ]h<e��K�0@9��+E�W�y��
<��=���C'_�yB�֡3��ȗ6��T�CQ�yBB]�=İ��ܢK�^������y�I*OM�$����H��-P��J��y�4R4P;c��1��}�a�5�y��=������|E}I��V��y¨�X�U06D�iEr-�Q��y�)Й3��|x�K�6g���p�I�9�y�k͗)q���qgU.1�F� ����y���Ȁ�"�R>7*&y��%/�yrCƆ}'`��M�,v������y"�L�jd��C��;!�q��a�<�yrLͯL������BQ0��0'�3�yR��zPY��Ҕ@=z]٠JԀ�y�*�/j*p�+#5�jP�[�y2Ȝ'��Y�.P�(�TI�F��y�aQD"`<*��7LF�̢����y�Et 2�lU�D\�Z���y�'��d�,����]�@9]+ʍ�yrD��~��Ň�:$"�֍���y2"܈e^��Rߍ9j
��Vg�y�/����s��1"pP����yb��;Sr��CA�$Ѷ}�$�ś�yB���1F�.1Ȁ�x�*YI����S�? ��r�/�;.�8m���
��lZ"Oj����e@�9B����X��v"O��ȶ�J�DVb�x���ABx�zP"Oư�e%��2�T�O��J;�dC�"O�ð��%'
�:�A]=#���T�'���ş���ܟ��I��h�Iʟ��	,#6��B��gb�9��n@$�����8��ݟ��Iܟ��I����	؟��	>,D:����8�;�N8>Am���,�I����	ן��	П`����D�	� ���0j��F9
X8Q��	 ���	��Iß���П��	� ���8��,@��Pb�OG�Y�&U��`ƌyf��������۟���ޟ�����h��ߟ0��9��S�e�(���)2MO�+�44�����	ʟd������ퟔ��՟�I-j�J�C��)��p�b%%� ��ߟ<��韔�����	џ���ڟ(�I�d�ڐ�S�I���J@"=ؐ-��Ο��	�0�	ӟ���˟������I�egpa����knA� b�X�N����H��ʟ����I����I؟��I*]��)�T`�Q�U�s�[h�ځ�I����ß ���@������џ��ɦB;�QAέq���JE�@<�Nx�Iן(�I㟀�IƟ`�I�� ��۟P�ɔR�*x�E�8r���j��_80����I���������	����������3,X0�;s�, �0�G�M�{�2x���<���P�I֟�	ß�ߴ�?���"������Y�_(��7��'/�W�jy��'��)�3?aG�ii:�����x��Qi�+2���Q�Ǉ�������?��<���U��X��ڎ3x>�KTe�%�2�Y��?���W��M#�O$����L?� v��5P@���f6���ä*��ҟ�'�>Q�g@�8வ��-m�Xke���M�%�u̓��O�L7=��<#7�f<Ѐ�1J@iٵ
�O���b�ק�O�xC�iW��֯$=�hĔT��\Z 	�<|��$j�LI���=ͧ�?�q�x���*Ō�3����M��<�/O6�OnuoZ�7�c��� �C�p�|�q�7�<���Cl��l�I韜�I�<��O��Y!�N���9U�������	(O�34�5��(N"�U⟔Z%'HjpB��ҜJ�"�X��iy�[���)��<�u�:�pP�'��h�bb���<Qұi����O>�m�R��|:ѪR'B���#�;ym�4�+�<q���?9�N
���ٴ��d}>��'JI���Ti��p�	ӎ�$��Pӄ/���<ͧ�?a���?I���?�wi�\�u#��J����A���Ħ�jp��I���&?��I�GٶPJK����5� �r@!�O8Hn�2�Mk��iQ
#}bDL��E�nˠa�U�~���]I�p��4/�~bc
W@F����'7p`�O���-O�q�pd�?�(8[�-��3���O���O ���O�i�<1V�i� pA�'휤qU�IK4Z�:�O3�X���'�6�$�I���OT6mӦ!�b/T6X,̤��%� rø��PM�_w�9o�f~������3h�O����7��&#��w��ʃuez��T�	ݟ��	ߟ���]��U��Q8��&Rw���ȑK���x��?I��i���D_��T�'��6�:�ĒI���kEK*F=!4cL�i(E��}}2(iӆ\mz>m��
��Y�'�$8�N�
up��EW/
�)�PH�X�.����~�'��Iş��	���I0Pɴ�s����}��a�6P�P�I��'�7,U[*�d�O���|���
svT��h]�N6�P���z~⊰>�¼i��7�\ݟ�~��&:h�����=� I�8i�h��jC%`P�Y2*O�˪�?�gi!���"o�� h���k�
��A�v���O��$�O���i�<QҺi¾5;7��x=ĔУ���@�L�%�+s���'��6�4��-��DV�=�E@A�SN�Q�H�3U����;�M�@�i���h�iw��RWJXq��OK��'�X`���`Y���/C>��ə'����(�	����	П<��I����]�J�{�bH9G�h��h���6m�K�P�d�O��<�	�OH�nz�5H� ���D�v6"�	*E@��M��i����>�|���M�'���P��m5ԉ"���B<��'�z�����8(4�|�Q���󟘫�"X���A�ɛ6��=a�����Id��UyR�b��|���O��D�Ob�0FϼBT,ɘ4-G�Z��i�6��)�����ٺٴV�V�T�qh�#�Np�5� ���aVd/?���1	8ʼ:�lˡ��=����!�?�3�19�*�S4�͸Xb�㱩��?q��?���?i����O8��τ�B[@ԁx禁P ��Or�lZ�>� �����Đߴ���y'�\&0舰��� f�J�P��H��y�Bh�:n��0 � ���q�'�J�r'�H�,Ǌ��	R�L�U:'
�(v�<K'���#��T�ܕ����'��'���'ZHL10	U�
�ԀG��/ Dn��T�h�4>7~1���?��"�'�?)�4n&�Q�!�h���T�����SDV����4<���"t��E�d����j"�[<v8��hf钸A�0o�X3�I�KE<����'�b�%���'�)��!< ��T��I�
�n=���'��'�����S��+�4x�@C��#�d��F�1Z�]IC��+k*Y2�yj����[X}�Jh�,�m�П�#�L[�!�`�3����q��˸tN�5l�o~b�	�,�
e�E%BBܧp�k� ��#O[1����J�1YV�-�R3O����OV���O��d�O��?�6ޢ/�L��j wA���B� ���I�4qZ��̧�?qd�iB�'® �J��4

��Իh!R�� ��O��l���e���_:`>�6�+?Qv틹f�ˊ.�Z����әr���%���Z
���{�Iyy��'C�'���97/����D��F�� ������'h�	��M���қ�?Y���?�/�Jl�P�օ=tZ�q�Ö	 d�Ǖ� ثO yoZ)�M��'x���L��;B@�����
2o�@@e�4��DK�C&*��i>]������v�|��(�ԅ1�,�*T�!��	1(�"�'���'s��4]���4R���s��E+U�L�[1�ݏP�8@�FG�?�?��;śf�'��i>��Ox�mR�d:��k�ą3�Q= j���4K��&o@
Y{���t*u�m��ԦmyRm̀b��9�7`-nb���"��y�_����Ο��������ݟ8�Ob^�;���U�`PӇG;IX4�*@a�`���
�O���OԒ����N���:$�(9!��D�f��!s�CQ"Y�	�4gM��8O�S�']{n�Rݴ�y�(�9�=���WA�w�6�t�|���TAɶq��x�kQ�	vy�O�2��� (���m2ت��Q�B�'�b�'m剠�M��ʂ6�?a��?��J�-}����F�5Zwڼ8Q@���'
�]{�m�b�IC}rl�('@��V��^,���Q���Y�q�*��٫F�1�P� V!y��2��;ڔ�1�b�;ADBŲ�'��p=̉.�M+��?����?�J~����?���h��B!%�7b�x5s�ɓP5*��5u��+L/f,��'��6�-�4��n��R�|i��
,���ӸI�$L֦�h�4-��v ��&֛&��D��-w������1p�-��l����}�����'f��Oyz�4���T�I�\�I:7�Qc!�	Q( ��I�!Rq�=�'a:6�1�
���O��埀��=���I�fB� k�j�.���jl\'���'���i�6��p�OȾ�۳��8�Vl�A;F7<� 5��C�>�iDX���p��\&�q�wyKK�L���ʱ9d���C����'���'��O?剃�Mӗ@��?0�}+Vű��Z�y����+D=�?��i��O��'sd7D�	�ش�6��/HT�9%
�.�X�E˱�M�O���.���r��*�i��s���4�F��J�=P� UC�h��<A���?���?i���?	���'E���B o����GV�dl2�'-�%k�V��<����AʦM%��+�ܫ6���vDF1�~MX�W<�?a+O���e���
+Gw�6�9?�W��83��Q���CE	�2o�.�,c2+�Ol(SN>q*O����Or��Od�O��%s�lw�؜LB>�V���O��vћv�
(�"�'��Z>��Ъ˲^R����4��2Ģ+?q�Q���42��L�O>b?z&_�V�lx�2f�Y��#ܣw<����1O�����JПDі�|2+�*H�!F��4�0$�
�2�'+��'Q���[��3�4$ؤ��@^U�@m �NH@]ޙ�����?I�r�f�$�{}B�aӨ	Zp��j��9�cn	WT*��q���9#ڴ]nv�
�4���D��)��'XT��O�F�,U��ݫ�[���Y*�`�\�'8b�'�r�'���'�哎^��%ô��-m˂A�[J-���ܴT������?����OT>7=�Р���!�2Q�P)�)ւX���ۦ]�ڴMW�Q�b>��ŖڦQ̓`�ұ�BK��+��c��N��<�+� �3H�O�đM>�+Of��O�Ż���x��肤q6�=�ׇ�O���OL��<AҲig��[D�'�B�'y��`�&:�P!ӢL(�����TC}��a�&�m���M;�P����挲c:��d/�	Fҝ(��:?�C)��u��[P����'b���$��?)ţ9Y1���jB�`�ԝCO]�?����?)���?	��I�OTHq@�r��pi 1Mw�*���O�0m�1{|,��ן��4���y��`e����	ۢl2�j�Ʉ��~��'ݛCo�Z-�%k~�z�z⽹%����e�>F�V �KJ�p���H>	-O>��OF���O��d�On�)�œ�l�\a2FJ\Q�2�+dŲ<A��in:3��'�2�'��O��Ƈ�*(藁I�r�D	pw�Ł#@j�LH���t�j��	M�OT��0q���6Q��)����P97l��)�0��Q��C%	\:S�")T��zyB"��{D0@C�m�NdYcȐ	��'��'��Oi���M��C�?Q����6*rC*.ǈ�k�ჾ�?���iD�Ox��'<�7��Ǧ�jߴ?�Q��P�J�1R�9z�ī�ǐ�M��Ot�1���J��=����[q�_Ҏu`�H�oF8ȫ&�F�<Y��?����?y���?A��>|C��U ʄ0���í	%R�'Bjo�J8�&1����֦�&�HC@��1�. �U̕*?�P����?�ODEmZ��M�'L����4�yB�'��yg��f!dKu*]�&C�+v��/p�ĉ�I�T��'��������쟄���oL(��e ��{2*l��ʛ6U���០��P}��j��g/*	��ʟ���$�M�'H�
�+BI�$���b6M_�@]�|�'e˓�?�ݴ#������Oy�fKY�/J`���͒�(1�$D@�l��!��g��Uv��?ISf�'XV�$�RW��,C*�Ȗ�RpE�e����ퟐ��şD�Iߟb>Ŕ'��7��<iVƑ:��!EWn�2��	*']���u��O�����?�Z�t0�4��A�{���X"����yV�i��7m	#t"�6M`��@o��nT�|�'�O����?� ���ũR?xr�#��XY���g�i�2]�' �'`b�'�'e��%���9#@[�n�E��IIOHYb�4?v�l���?����'�?�Q��yg��='K��6���&�:A�a��95&&6m���E8���4�0�iꟜXs��v�,�3���%x9x�r��;Nh�	/1,��w�' ZT$���'�'1�)�`�P]�!a��[,F�Ne�@�'$��'��\����4P�V4"��?��	;
,zPJ�1
(u 2k�9�hͣ��E�>y�i�66M���'�:P�`'öٸ�o�2���c�O�mSS�"Fq@M��8�I�#�?io�O���.O 8�Z��F�*h�m�CG�O��$�O����O��}���d����*!,i) ��[�Z�!�f��A�-B�'��7�&�i�1��+�0FCPQ2�Ŭ�� �V�j�A�4
"��b��+� o�Z�\�eA�m�JEA�$��	��P�4KʡH$u��IX������O|�D�O|���O���R:�����Ȍ�(�z�j1:Vl����Ζ<�'�r��$�'_ܹ�7�
�TTb1dE$H�� ��>���i�\6��韐G�d��s��4�#�I�?�q�P�^�	n��gϴG��I�z�"A��'��&��'@F�C��6XҰA�s�5|�pU���'�r�'�����4\����49�lq#�~�t�#G���	�uX\���-y����\y��']��/`ӄiy��^� ��`vmB�?'�7M"?����u^��	�;��'`[k�e3~�{�`�`�8�����^���O��$�O����O"��<���쓔@NDUisfI�
�I���I�M�%H�|�����6�|��]�H��`�\4��t9u
����İ>�Q�iG� �'g5��4��$ԻD��p�'0D�X��U�b�$TD`N��?�$�(�$�<)���?����?��䘊F�ތ���i�L-Z���<�?������ަYBjE�P����0�O](8#���<nv�	(��*��D!�O���'Q�6�Ħe;���O	�[�+'mv�p�M�#X�s��$,��Be�	Y��i>��`�'9da'�P���#�(21�ԕM�D4 �mGٟ��	��	ʟb>��'�7��?j��8��3j���h�U;�����O��DKϦe�?�cS����4|:.)�����8���A')uPM��i�7�P�=�7-,?��,��iB'��d^y�T�� H��W`
Gc��r���<���?����?���?i,�F՛��ܶI�12%F�%3j��$�����X^���	Ο�&?��	��M�;N�f�͙�&��p� �p�t��e�i��7mAɟ ԧ�O�~��iC�^5)�!	���o%r����H9U�D�~ڤ���B�O�˓�?���L�8:���Ϯ4�� ^I�,!����?a���?�-O�,m5`4��I����kTu9&τyr��`5l-a�F��?ɔ\��ܴy�����O��a��9�1��G5�CEХSd���'�j� �(�P������4���|�$�'�a����qr�9���S�Y��'���'���'��>��	e�BT�Rƚ=8�ʽB��#r�D��%�Mf��?y����6�4�P8���Q�uL��m�>����A�O`��jӂ�l�\��Tl�]~�rFv��s�y�*BW|:d�1�\4i�X�Su��	����d�O ���O����O�dnQҵb�_^\�EO�}�V��PU�d@شu����?1����Ou�آ�n�004�)�U�-��ڀ%�>���i5�7���@E�D�G�W}6ԁ֊B�0�\��U�7��R0d���I?H��J��'uX�&��'�B�Qb@&2���@B N�{�l����',��'+�����P���ڴf&����vԄG�Tw ��dЂ8M@�s�`����A}"�h�"%m��MCa�̝�l}����.�Э��I4gD��Aٴ��Dъ	� �J�'T���Tܮ1)ASt��-  ��2N��u̓�?���?a��?�����O���[��Q͞�fc@b������'N�'|H6�]���O�m\�1�dT�A*j>bx(esv����������|j�X�Mk�O���H q�0�T��;ȑ �o���`��GeғO���?����?��?(^q ��E�u�P�s)M�&D�����?I.O�m�:T�����R�N'QZ��'�^�pM�X�ɲ����y��'v��E�O�c?���'D�� ��&+ǵn���`�N F�"��n��m��������*f�|d	�6:�eR�a�?M���qb��\Tb�'	b�'z���\�`۴N���2��b�����I�T�`�D�?!�-T�V���W}��w�4E�.	�n�(X���9R�X7I֦1��5�oZ~~S�O(.-Q�	�V����D�̑����aB2�/�:.��<����?����?���?�)�ح"�Js��p�FBYk>�y�pI㦉�F)ӟ,�������W��y�_�X��Hȕc��6J.)��T.�7�զ�����	��6�j� ��n͔AD�Cw�[-qIDePf�}�x$��2u�r�FF�ry�O#�{�����ǡ+���%� t���'���'5�&�MS�ϐ��?���?a%�4d: SQ�G_�~j#���'@R�``��,x�b�oZ��D�4F��9P`�Vh�<ZP.O6��	�#�D"a�T�r2l'?�B!�'l2l�	<o�p(A�K���4GF��GT�l��Ο8������u�O�R��*<=H��FL�BJR5B��I(8�g`Ӡ)	Q��O���ߦ��?ͻuO�A( �1�Q�1�G1p�n�̓A��6�b�z n�5hT�nZ^~RИc���S� �Pxr`	��ܬ�A�çA�X��#���<����?I��?Y��?a����7Ht1� �3`���EP��� ˦x���ퟠ��Ɵ�¢�M,M��q����A�:�����M㴼i�D�8ҧ8\>`��.($,dċ��n��h!D�I��q�-O������?���?���<9�M�9�ఔC�-F��QF�?����?���?ͧ��¦I������l@vE;${0�(V�^�֤����Ɵ0�4��'��H����v�0,oZ�
��P�O�G�DA�q��f<��`ئ�'6D��� �?����tD`�1��@.cU�=��,�0�n���p���I؟���矬��埠��aA�6\��Rv��c�a���}���?9�*D�V�U#����'�7�*��կL=�<�D��8t6<� �X#W�^���Cy��'���O�>�*��i��I�_�~#� ./�����dOY��]���` R��N�{y��'~�'��bV�Ҝ)���7���WVR�'�剁�M���O��?a���?Q*����*@��2#%\�A9И���O�m���M��'���v�P�H�56*-UE� ���ZsaV�ؤ��ۢ^����|2���OF��M>�&�Ԥ����S&/���2�듾�?q��?I���?�|Z+O.n�|��%JT�\j|����7_��K��x�ɯ�M��"I�>!��iĝ���?8( ЭQ��iJ��|�2Pl���rӖ���� ���ݘ*O<��Ш@�_����go��> ű�8O��?	���?���?������)f92�z�昽6P��� Q�q�nZTL��	��IA���r�����a��Z�q`B�Gx�T�জ=�L���I^}���N^��:O\-3F��*i�z�r�B�]����>O
�rD����?)���O^˓���Or��P�e��	�į�t�Z��v)P�`�Z�d�O��D�O\˓Z���R�n���'�g{Qr-���/s�ԉ� _�N|�'�bm�>���in*6���]��O�-I�#՝&}$c�l�":�d�×�d
�ʙ�&:(���n�S� .r�����+�+PU�A��j\BónO���� �	��8G�$�'���Ï�E�9�׎��F��<@��'p�6��6�����O�Eo^�ӼC�N&BSB����Lp�h�A���<!e�i�^6M\ꦙ�s�O����'�R�����?��܉#�\	WeQ�k;������]�'9�	ן��IߟT�I̟��ɨR���rD拻�;���o��=�'�X6��5lǘ��Of��<�i�O,i����3���06�Ҕ5���)�lWT}ed�jYmږ�?����<�|�/ȸ{����`;w��Qȱ��n ʓ=�d9���O� J>�.O~T��m_� Q�i	��O��XH�L�O��d�O��d�O�ɺ<�`�iK2(Z��'��tj�+�[��yBi��tOnxS��'��6�+�ɬ����립��4O}�F���1�.P��x� �C���0Rq�iZ�	��0���OaL�&?��[c�~q+��,;֑x�k��z�֨)�'hR�'���'�b�'��%�ENݏ@T���eR�X���<9��+�*�.����'�7'���GT�3a/H���!���T^p�I~}BbhӪ<nz>IYp��Ц��'%>H{`��(���o�C�p0��Ǆ�3��y�I�x��'��	쟰��ԟ��ɾh��Ae����hR��ðK]nL�	ҟ��'�`7mC�d���$�O.�$�|Ba���4����: ����t~m�>�Խi��6������~�F,ae.�1���6��ԠB�En�ɂ�h;.��+O�Iâ�?�sl&���� �s��; �<)ĉ0�����O@�d�O��I�<�1�i����f��~�P!��C����&#K"@mr�'��6�3�	4��D^צ��b�!�Lp blU�e��<�B��M��i�Ҝx��i���� �H� ��O���'���[�SXi��$+�!�'��	��h�	�0��Ο���@�Tဟ���E�̢8�H�Ra�GS@6���@�D�OV��#�i�O�mz�=Xen�j���*W�����2Ѓ�?��4Z�BR���д��"���	/*�ة�q��*�R@�*�扈+XU��'+ P�IoyB]�T�����Ćȡ7O�z��:-��u�S#�՟���� ��ly�i��5��A�Oj���OpU��(�&Z�@Y*.~���5��3��$G禽��4���l�>Q�.Nb}�0i WpBⶪf~Ra�Ӣ��h�42��O��@�I32�RB~a�0A�o�{�ఄ�\�(	��'�"�'���Sȟ���8P�+�㐖>^ժ��:�4\�����?AG�i��O�m��Q�fo�-l��J��I40*�Ħy�4*��������f��p�UI��jn�DLQ�]�:�z�Ȼ1�� ��	�Am�&���'�2�'�R�'�B�'=&�:X�F[�,�t�(��RAG����Šu'�ԟ\�I��0&?Q���F=p� �O��)	J� �����(l3�O|Ym��M���'��>B��B)"ka��#Q�CT���"��#R'Uyb�o�V\�ɚ8�'�剢+��\r�哪ZQ����V
�ڑ�	����� �i>�'A�6���U��$U�Z+h�r�.�Rq�x ��t�T��R�Q�?�%[���ش^���nӢ����:L�٣�E\W��$��hςe�6�<?1��Q�|����P���i�k���[srebPK� [4���鎋aQ��O��d�O����O.�d?�S3� s&҇�Ɯ�blSa�j$�	ɟH��(�M��,M�$Cb�B�Ob!�J2��VBA&]{��hAa�� �'�87mΦ�#:���nZv~���� ��( �Mu���*r�e���\;���`ܓ���'/��Pʘ�?�dH�#!B�k���B5�}A��h�<����79`�W�1F\��>),1Q#@��2vf�q�$T��t2�#ԒbIB1��!Ө�KPB�!P��G��)0��
X�.��SJ_H�7��YIT `�k��x�Fb�{�"�qU�l����AsέP��9smVLkUFL�~]�q�:p��$B�b��o,@Y�"�/%��T�dDܴD�6��OT���O|�IO������ߴ'��a�@ě@N�	'����ȟ�(�
ԟ�'����sQ! �JȻ/�ȅa�iP�4�U�ش���_�`�x�mZ��i�O��HZ~�.H����! G�68r����ġ�Mc��?�/?�?	L>q��Tf��<�rtS��=?�p2�
�#�MӠfHa��'���'z��F,�Ɇ<2F�ф-�@f^	��ݔeR<(�4l}0Ő)O��D�OΒ�����O�h�@ɟ��й����~Ǟ`0��䦁�������;C㚀����O�Ӈ
�JHɡg���N���MP�S�yR�ͲQ������O���^	u$&Ac����is��qO�_��`�'U>���'�U���	�$h����ѢǞS��@ZVo�up���O��q���	˟��	ܟ��	ٟt��dвc�Aʇ�»
$b����W�Ce�I䟬���P�Ir��T��YV]����a0l�cb9�\�����Q2��?����?	��?��ы�?Is �q��c�g>:�=؆k��s[���'R�'��'B�'�,z���!�M+��.T�>�PA�̹d�j��w}b�'sB�'|�ɍb-�0"O|2�+�O����36�������ݛ��'�' ��'X̙��}R��	ш��c�^�����!�M���?���?��
����O������c�v����n�%�6��3���&�����0���1<��c��F,j!��q0���'n�nZß����8�r���Ɵ �'����'Zc.���<Z-@`e��+J���ܴ�?���������M�S�*���C��2�`@�cP��6 n�(vD�	ǟ�'��4�'"X�$ねL�h�|��4�"]r�q��^��MsBڴDg�l�<E��'����#�	�B��ű#�Q%M�Jy���'<��'3��'(��c���	m?qtJ�:�3�(��B�y����p}��'<R��%#H��ǟ���Ο��{�nAh0H�Ũ<)������n�Yy"E�|�)�[�a��N�D�p�h�F�.�"Lj�Y�x�pM���$��?a��?�*O8�cKN�S��Tg��prx�6% �4y'���I�d&��'7n��S'�"`�`X*��b�E�ͱ��'��E������ݺ<?���#�8½�d@��y�)��U}Zh�e@�J��C�$��'9ީyƠL����⊬����2e��m!!�n]-n|�WaH�M$\���E'�Vl���R$q	�d�������ò��Bҵ��gE�%5Լb�J9&����_>*��Ȓ��e)��)7d<0�S��)�@P���Ԝ��r$ϭ�"@��.��EAN5p��
� �2��z;��;4 �k�d|���ĜS�������?1v.Jkc�LI���=FTA:��Z���i�Df�@q��R �$#��"��V%��Ɍx4ĝ�F�^�Zy 0�R.����S@҈F娅�Oހ��暧7�"��.1`LJ�X b�O"�lZ�H�6�)���X�iG1A(����Vl*�B�	�r��c�χ+�FxcE+UJd����g�'��xsR [���b�o�-��rej���O����?���I��O��D�O���WԺ�FfǜorT9� ���bfHY �	]6�E��>��3�h���L>��J�(���QjQ&�t�A3K��p�a�/�&�9�J�ȴ�}r##�Ty�f-��Ȑ�v�0�Pe�+�x%�	{~Z`L��S����	���cA��7-�jJ�(��i�ȸ��~h<�q��-T��h����,&n�Q҆�a~҈4ғ��	�<�ń �m�vѫhh�t-y��E��dT�	��?���?��h����O ��p>}�.S�c�mR��r�*}�"���<R����?U��l�>|R���w�I�m���,�zȆ(���^�iE��)P�X��&����æa�6�D,w��b��T#���K>q���(�Y1����]I�F�B���#�M�Q�iTBV�D��F��[�$���)�����cH ��U��U�B�ؗa<A����B��K���<�#M���$���N|*G�>u����\)/2�|3��O�<	f&05��d+�(N�GLār$��K�<�I�2�8$@	�X[�u�Bc�~�<9�-������.π`�Pف' R}�<��F�>���Z��˔<͒�)�kB�<a�%�NJ�I'MD�ka��C��|�<�5oثrĸ]����(�8(jU�|�<���U�3b��� Ȍ��pLB7l�u�<i�$��M��&Ԅ��T�%�y�d�	h}L�J�΀,2�r��W;�yB��)z�R|�1�2Ft|��0N��y�B�X%v�����J`^U����y
� ��Y_�gt����T,��}r'"O�L�òA'00ZA&ؔ0��}"Ov�����f!�Ef�(8�%�"O:89&@�`��=Hv���7� �V"Opr�a�j;8����ۏ$��"O@D�@+�P�t�0��~b� b"OT��dN9Y�	{u�1��"O�q���8�H3@ڍ3�^qq"O,��āB�aXX����ȞHN�"O,`h��*����#��)��"OJx��;%Ŭ����8N�x�"Op�#��ըB�Z�B���	k>��f"O���Nk��8rp�\��
u�"OB�2/�
�XSAҍXK5H"OL z0"A�&(A���:K�0"Om�`̈�D
2q��@ۨSH���"O�=0o��:���SVo=���t"O�� �+qެ�G��)B�S�"O��"��:�~��Q�Jlȣ"O�������g̈́�z��"Oh�P���<�X鳔V�e��"O��1��e��  KA��zI[�"O�񺰋�<���I� � gܞp��"OVh
���d�I�@n�	:ܤPq "O�8ڃ,Ĝh2�m�����k���"Oj�B7��3�n��6�1|^m��"O$ ��U�\M��R`�f�4��"O�SeD��	��D+t�X�t�1"O��@��^�(t��@^��"O��R�18' ���dK�WI,��Q"O<���Q+�d�Be�HdfAyf"O����&�D���cR'pVXHf"O\$
��XR���dF�h�p�r"OL��!Ȑ4�ĩE&�zaF��"O�,�U57@&�"2�R�)�LM��O��2�$�Oԍk�%M�4zɻ`��q��L�7�'�ƨ07����	$v��c��-N��P"�?D����Z#SĒ����+{�%"�+�^q���)+�ar n�t�	�a�U�Rg�C�	�~[*�b��	t���J��Ҵy��0鳭B	v�1Oģ}�4��	2Fl0Z6�q¢I;
zZ5��)��Y���d�fi�s�A:��)K<ў't��W.U5v�Xڄ��L�|�J��1e�'"������<�,U���b�����|I,��ԋL�XpG ��v�Y�7F
C��Pː��!7��I�d���=�����/j�đ�h�;C��×�4r��'����2G����		ָ1H����Wnp�i�� k}�%V%��DB䉔�ʴ1#���	��LK"/�I���\;Q��h�xN�%�'�Z��O|�`�Q�A���/0NHP�Cѭ{ vĻ�N?D�X 7��8rz�X3�@ X���kD�%�?�!�_����A����4
�����j�P�M�sɎGY�ѱ�+�o�
8��Iz�p�C�%M!'>��+��+2�!���8MdV��5��:`?-��.C9B�̌�Bj�^���h�#��t����tb刐 7�	��"%����t���a`�?�7-_�dy�5�_&A~�h��ʟ5<���钑�!��<���ę .�����F&�\��1O+L��*\n��Uc2��%�0Q���yW+kpP�[Ӫ�WD�( L��y��8;�����MN��81����l��ADR?^-^���#�3�<�+^w`��҃O�w�qO�8�Q���`D��(� B=JTh
��'�A�Ca�*vXsV�@0Z͔�z���
o,X�{5�eK`��D��G�ب���݈7��zR��l(�A������G�ֻ��'>�Ъ��O90�hJ�D������:/~��'۞z�=�t-Ŧo��yx�%<}�C剹|��bI7�JY�`�U3OI����g�v�r7���j�4����=��aM~�<���z',U#m\���
kPR��'��@K�c
�:?�1j�G_9 5��U�����@.��	p�a�r3l�S����
�1b�0�8"1�>�I��-q�P�VY��� Ԉ�<	F�X�M��,s�	;~V[������ �0��H<,\9TL,7������)���q�ʅ� E��q�.�8��O�G�<��`�Uu�=l�4����K�gp� ����G�I�3�I�䁀�@W�t��}�iɾ@�2�"O� H��݃t�"ق�͆��\$��/�$<�6�F��O�a�%# W���ͻb�(A�fmǓj��5b֧j�jl���0�f|���ֆ"H(@0�L�=`����'bN.}X��G[�	�<���ïv���"���>@b���q��W �l�%靲#Y^���7��+RW �`��޵u. ��`C�%ǲ�?��%cC�J��+�`�},B��co4D��B'���@V^ ���ʢ�&"��4��	`�"l	�-xtf� �����C%F�-^�b�zFE2UȨk@��r�<�V�H;z{"Ay�c�3-�~Њ���4(��	�W�68�����M�S:�"�<�,,h$�ϙ72��%( ��R��ô$Q!=��
�R�<q8����%���(��Cm�f��/�{�\��	�*eh@4h{�ʠ��"؆ȓ ���[_-����A,P`��ȓ�@+Qa��w	Z��t��?^Pq��w�&ؒdE^����[��6$��	�h���*=J� KN�"0��ȓS5N$'ϙ9|�8�6�@/`M$!�ȓ0UF���ŎH��@�/w\�@�ȓ�����Ûpil���U>U���ȓ.���{0��<���i��<	L ���h#s�ƺ6���©��{��ȓ\d:8 ��˥hc��!Ū�	ܩ��{���xӁ�+BvD`"���Ze��ȓC�\�K�e(PtǁE|���mUԙb�E�Q����Df�+rjՄȓx5�Y8!���/r���*�
8ھ݅�vA��Dg\�e}�M�P��xd����	`d���dڲ[�F�Zr�74x��{�|e�gg۴��yr��ع3�깅ȓk0*�K��]�>�:Ub�a��q�ȓ �-� ���c���6�Ӊ"�����T����<BGRi�&��+�l���k�|��	�%}��J������C|VL�G��	^���q��əE,<������7�Ƈy)�� k؞��-��-������N��܁Q (��)��s����S�DliQ�Q�gaɆȓ4�2�![d��@WL��j��@�ȓD< �S%6%�p���//����ȓ#|PWʆ�|U<���S.|�Q�ȓz\M��m�*-��P� �F,�J��ȓy� �'둑B�e�w)
)t7Щ�ȓ��Qփ2/�n#u�D�/���� �&����Y�'V>�B [� ���ȓO�����HE Hi����P�ڰ�ȓ7���qN��VN�I{�iH*p����U���&��D�(ň��G:�0�ȓV���2,�:�^����\$1K֭�ȓU�[ê�N�قI�$�� �ȓ��˵	EgB���ˡ6�9�ȓzL4Ng{2���$^!�t���P��rF�&vb\���kѪ��ȓFpZ1����*ܮ��򬜴!x~�ȓz��	�`̎X�q�0�D�A��S�|����ͥ"2%rW�̌t�걅ȓ�n��p��3H!e��	�����9�$���J��o�xء�H�>9C�͆�`r��'�M�R4�4��7\��͆�D��PPG��c� #E��)vU�ȓF���R4�Y�V,
�YF$)��
\�0aiI�H�(A���T�̅ȓZ����Q�h�RE�ʑL^�A��S�? ����MR6��j`�9B^�"O|͸mRyW�YHEIV��r%"O�@��NZ�DRh�!��'@,|Ԩ"Oƌɷd[{�j)���F�T��%"O���茬F��E!�L�HU{"O��˴c�s$���B����xh�"Oj�b�G�0��M�U��G�A['"O��ٲ��ej�I��!S�άd"O�������ʃgݎj�\�ɥ"O ��Ao[�hh}�f�/� P��"O���rD��S��s�#H�#�fc�"O��+6-�>X ��@M�8=F2��Q"O���[���JD̊M�J��$"O8���-З߰1�
&@���V"O�#�\~��R��/l���A�"OJQJ����f	D1'(�G}��!"O|E�2����JxSǦ�rn�ٕ"O�\��B9�d��M��hc"O�KQ��59��0ze�Ֆ!4i��"O��`f��=�踨f�M�a%"O�Tk�l��X8����[�]J�K"O�P���K�o�2%P��XR,�%"O�L��O�R��m�JǇ:W. �"O���Aʶ,ʬ�hjOtdhQH�"O4x�u&
�=���yԨ��n\u�"OpX���#�*�Ӷ���n��X 6"O\5)p��#G���p����qe"O�	�a	kQ8�)G�H-~�y��"O�#�
2S�"�r�(P�R�"O����A�/:+ʈ!�^$!�\Ah"O�ٹ�gǸ',��ñ�ѣw��AH"Oh�*h�q��P��(t�@"O �ơ�D��t��kB 	�~�('"Olhy��6:`J�HU�J�t�"k�"OP1a��c�t�Rj!��"O``�&g�{\Հu��C�b�"Oy@䂥u�쁨f�_U�t��"O�M�-���*�p�GV$CF��"O�:2�%��PP�_�i&
]�"O �0��\'R���
_">hh�U"O�qS��Q�(�Wi��L(�"O������s)t$xPHW�_��I��"O�|���(_��d���S삜��"O��sV$O�}ƒ��"�&|� ��"O�h��
��zd마v�r��""O����i^�f��L��A��X�"O�����D[6Nс=��={#"O��D���8K���������Ye"O��{Z�K�.��.B.	�c"O>����G��葶��$>H�"Od$C�IEq����!�6$����"O��k���h⬄�fKV�R��3"O���PK�8 ޥA�
떵�"O�`�I�Lh`5��R���+�"OP��7@�)�dEK��Ė�l��"O��B+�-2�l�a/R�6�8p"O0aկK�����B�<�T�G"ORl��Ҁd�
�͘$j��EXu"O�H@��,my�@��NRSF�8 �"O��ce� �,��D.�j��HU"OHE���\9���kY)y���U"O	��&��a��!X��FN�X�*�"O�t����7�`,�h�C�:g�!�$Ԗ3�̒`��;Q7�偒i'�!�� ��رE��\�3��7{Pu��"Op+W��uI�u��%��$U&$"T"O�p��k���z�E�$C88T:�"O<�c�) �p@���O<�M�T"O�:�
W;j��FD3j�@��"O���«�#X��"�c�#h�(a�"O�]s�Q.B:t�ѡb�Gߞ�JA"OP�jG'�;)]�H0 "]�K����!"O�`PeB_�C٘51��_�x(x@"O��jGAZO�>�S&\�H��"O�1i�
��� P%޹	)��b�"O�]a��X%(��|a��I�8Jp�"O܈j�É�4MK�>KL�e��y�\�"7�m��ΏI���uh���y��"ꈒ�"°�f1�䄗)�yi0����
Y�x"�mD	�y�%ˁ2Q�l
4F��Y޲��S�Q/�y�ہh�N�+t/YQFnqV���yr���9�,7JLKm�L�5eI��y��S�]�Xe0� �2�~-Y4mJ��y��̗G(����H��%�ӫε�y�mG-)� Q��t�
d�c�ŭ�yB�-l�\e!��pG�x2�ⓝ�y�"v%@`wǗ�9X��;⍈��y2dR�$������+���;T@�y��L�\��� ��q�{f�Y��yB*K�n�6�r�����!�ܘ�yrH��|������ԛ&��p2`��y�Fl�䬸�d�~\|�sF����y2CH�$�@ju�ɳ@!�8�թ��yb'�o�Le�+��2��UFP�y������Eлz�Z�G@K5�yb���7�=Ӷ��q�
 ��B��yb��i58 f� :>H�%)��y���J����]�,xN鉵���yR�#hv�x��� 3������M�yBG!�.�J�$(��=��ۉ�y��M����+�)V6��� ���y҄8v�4��`�T�X<s5��y���u��!i�}
D͛�cD>�ybZ�V�KBIzl�*C��y"��
T^��PCa��	�ԔY�f�	�y��WXfL�
�����k���y��&:]�d %�9y�x��4BȔ�yEϢZ�zĀ�u���˱�э�yR��7��������,� M#�yB�X kx�8�%�\?v�6���I��y�j�9<.�Kf�­?��űe�˘�y�EX>��ڒfʿ��䱳���y"��N 22���
�����W�yR��
���Aj�64 I�)���y2�R�QY^�[�̑G`�RT���yB��&�u����=f��4�c�K��yr
Ӷ�4qva��YH"�1@����y��ȃ|�uكf�z��[@�Ӹ�y���+;*�ၣ�?	�`Iٗh��y����Ab�������|�,� �C%�y�G���yq�EJ|���1w���y��[2>D��P��&l6�G(�y�`˭X���4	ıS�fl�v戛�~��)ڧnU��[�LߦUj0���կ�8P�ȓ�搃F�N�k�L�
�)Ozy��iІI ����h���%�TY��me��Ӣ�?�f�#��D�mu|���S�? ��yTA�+C��H�L�C���zיx�.�D���O?�Tq�(" ���puk�2Oj�͘�'|~�;4l�av��	ÑF|��a�'���zsϒ�-#�$�@m��E��TB�'���,�,��( 픥I>*X��'�콱wƋ�LX��-<X^���'pd�B�s��0)�@S�~$B��'��l� 3x3:�
�R�x�pZ�'���@AԀ
��]��@�
G�q�
�'f�pC�;j�V�e�͡C��uk�'Į��Vo��]d��Iը6��1r�'�!cg����L!̩2�p�9�'.i�nA�B���K(tyԩ�'#��s%�/jqԴ��aA�����'��9ҩS7P���P�R�xY�	�'5� h�A��#y��&�ׅ.����'a@����*�~�x��/}n�U��'d��Z�@���]�?���k�'�X,Y�E h`Z',Ėf+<�'g�l�c"ڧQ\���A�,�f�+�'؄,�rLՠ,�lz��
{C�d{�'�B̪w
O�I=:��#�ĩcqŸ�'���y,P$<"E�SmĪn���'0~A7%��ze|tɢ@�Q��'U�{��=tK���QbI�"A+�'���Ae��P�X�y�n
	H��'W��(��ϚB�� �%G�3]:I��'0���!�a2 i��^�(~P��'��x!EϯY��\@���.Nt�
�'��T�Aӳ=��4�Q��Q�ث
�'ZB<�U�$bྉ�	Br���'����-N�'�F�h@韾P~B�B
�'�Rm��E\�H�h�P�a��I$��r	�'�$�`���n�tK����d�	�'� z#AI�Ma��I��B6$��E��'F�$���^<Y\���̽+|���'ִa��+p�](��I�!��R�'�A�5�*3�=s�Wy� B�'?d1j�<��=I��K���'QD��+",��ű�+I)jچ���'	2H�o�m���!U9\�m��'@�s��:�}��e@�K�'�ԼBB�W�Z9��~��1)�'U�8Y��%�ɜ	x2���'-����ٳ*�Ő�c��Z!�'�\�R	ۙG�Nq(%���jx!�'��ڋ8'&�3�f  D�	�'L읭(U�ְ �K�&� ̫�6D�z�� j@X��(��!73D��a�ń:>N��C�/�6H��a�1E2D�,�Ec�V���.�>��|�%�3D��	!�ye�S�ܸf0Hz�a1D��y��ߘ:�Y0�BN�$p@��<D�4����
T�@��T�+Aʹ�R�'D�y��JT��)�O-q��-i� 1D��Q`,�4��1A"����0D�0��Ɛ���E�v̵1�k.D�pa�XÖc&�*����-D������Y6�lڔmϊZN��A?D�� �eX�Z�D��cLVjIC�=D�|��)�*B��P�Yx���?D�0ir1��=Q��"�p�C�#D��s�aH�tY�1d��4V,���<D� 5�
�CHv�CA+B�F�Ց��'D�� ���2@
j�dTR3���xqp�)�"O��P�'
lƢ�S���h�"�"O� ��"aiQrB 0#;���"O�!+A�Q���Q��S�c"D��&"OJY#�Ƈ1I���O»U��R�"O���+V6**��2�$ab"OdܫPh��h>t��d��E��h�"O�4r��S�����I��T���"OQi2ȉ�n2�	Ua�j�t<�"O��s�L͙j"�Ep��ˠ:���`@"O^���K�@�P�@�M���U"O�������y�j���M�y�� �"OLu��n�;�4���
�ra��T"O����R6k��PBgJ�wx��� "O��g.[�{���c@�ur�`�"O�xj�0�Z���3P�9�"O���dK����j�/O��"O}A��/5�p {� ���4�;u"O�3��1k��@�-K~�u�s"O<�yN�x�77��EZe��c8!��Zo߾Ĳ �M,( h4-�1
!��Y8}T��G��m�@��,
C�!�$Y�|�x�jT&Xy�����!�dZ�\��i1��O�-,��ˊR�!��˜n"M��ѼY>��fh��e^!��&8ZW�ɝG�H�Q��TS!�ă�?1Xc3�C�4�&�B��S�.J!��D"��M[��I�ld�fB/
=!�Đ�%ļY��jLq@G�!��z��M�B��h�>\{�ċ�Qd!�䑡^�@�@� ��P�a�!��r
�c"Y�;���x��M� �!�]�k�H,dI#�n83��?G�!�DD�t����+d�dM[P�V�ny!�UC���k�5fܢ��({^!򤒶"�~�$EWyxl�y��;%6!�D�7F�p�ۢ*3�<����_q/!��4zu�x�&�U�u�ܐ`�煶p�!�dUj�Nա�i�4Uܬ%�Sg��?�!�$�-F�� � Ή���RťS�-�!�$!��q���J;f���S��r�'V�����y�2���Gŀg��C�'�xAA�ňKI���©�<[#�T;�'�T��!��bHJ�Rg�\�XJ
�'
r�@��ԬX�b,b�!S4Ym�lr	�'��@	�T��CG
U�tl��'�6,I� �1buI$h�2_=�p�'�@I
���)Ed�QaT�B"�N�1�'�6�g��;?��[�oF	�jm��'�8�����8�\�1ő�φ��'ި��`f �K���+R�H,��'*�{נO��f��P����k�'�&��p��6ļt#�e�w� �j�'�l�37�FD��0w��F��%@	�'�l���"1VͰ�����6E��#	�'޶}�MkS�L��e�9r 2�'���C�T$NN�Bɑ�.V�z�'���H.AN���C�Z~)�'��T���W�t�T���G^R��e��'V���Cl�^�nh�#�s": ��' ����v��*����h����'P�푥l5!i�|���T�M�8D��'��-)�EY#$����A�xx"T�
�' :Y�'Ԟx����
kk
Ph
��� - abZL�%��c�=2���c"Ot`1�dư	'�͗)Y/��Ȇ"Oj��&��+Tɫ�k�WD\Q��"Ok ��"ř�ʁ
4b-�5"O&̘�FH� ����C�TX�b"O�9��n 8PX8I�"#'�p  "O�y9!NB���ć��5���H�"O���띊E���zw��<8^��s"ON�"ĆP�"��#��!B/X��"OBl3oܔ%�dⶁ�e����%"O�]��I�&��I���~4��"Op�����&P�6U�WA�x��,;�"Oཱི�A!F��qcM^��Ve��"O��b��Z{��˽&��k'"O� s����R��S �
1�$"O���5�A�Q`����Ò"F��Pj"O���].T�XM�BH������"OP���h5�ٓ2-�%w(�k7"O��q�aC�Vd@\@�!u}�
Յ�@�<D+7�<��!�� 4h�"�O�~�<a�ÄZ�� ң�&�B��!K�}�<q�553�q%�<E3,�s˒e�<!��ϊw��W��R A����G�<)šW4O��mؕ˔ u���2�OB�<у��E�ZM� o!��s͂d�<�ѩQ{؆��DX"$� �c�<ЕIt����0fб�%�^�<��匝+4�g��h��}c�&�q�<�v.���<5'�
?��9�Kx�<��"xP�3"$�L��F��z�<��/p_ԙB��zơQW��v�<��j�J���Q�lԞp�&�D�[h�<	b��c\>q�h�6��{%�|�<1a�W�,".y��Ά����t�y�<�פ�.x r�I�L��!�VP�<1��+Q��"�
4��У6EYJ�<�dG5_Lx\3�#�G�i#��Qb�<�'P�=d�SC`�g(����c�<�W� 8�i�;2��T ��a�<�t ��$`x 	<"��!�g�<�׌�"~@b]4��:)�x�i�!Ba�<���,nR�1���(��!2W�M^�<I��=!�9��Js�� jE�VP�<�1aK�Nc��q�X�E�ܨ�#.O�<���Օ)A���N��9�LK�<��hO�yr�dmێ#*�ق��q�<�0&�!_��X��0z��x�̕y�<I-��{aѣU�,<�5P���r�<	'@��x��ţۦ�:�C"\m�<�bј(��
�&Z�<'r@�1hm�<A6d+�=�a��<]�!P�ă@�<�fL��N���f�8H p�lh�<���"@<4�S��57��<yU)�]�<I�a��\L];EŖ-2�H\k��D�<aRm�3 ��R��+Gd��R�%A�<�t�1l�j"�F+Tm���F'�@�<	�lL
?��u�VJ_'Xp��𶣞{�<�W��1
��R�_V�$$������:\� ����&�H !�+�Xg�l�ȓ/8F=�Ae_4����BeݷF�4�ȓ\Š����Ӝ&T�ċA�ɵKR��ȓ�|%�U@�otX�Ԭ��
ْd��2����.;l)P� K%Z���U����$ˋ&TZ��!�8�~$��S�? ~|�B`�7�Y@4��:F�y�"O�	yk g��	�7��)�.tڇ"OL�r�g�oЦ�����%��DB�"Op��@���s�M���:�"O����AR>Q�(���摼R(�)�"Olث��K�&Ʉ�5��5{[4(a"O�X"Q�
=咠Rp��&h�����"OL� 0_v����<X�B��"O��h`��Č�� 
� ���9�"O����hN!2������'�΍�%"O���j֡|���
e������7"Oơ�RoAV�Vp�NWu���@"O�tIթ�tҥQ��Sj�Ъ"O�@�m+uX:eHsc�)gl9�R"O"EI���ډB���u�rq�e"O���ǓX  @�C�%�fbw"O�A���w���6�(��4v"O�h���Z*.TȦ�		eX"O�{RL�3�|If�6Nʼ��"O�E�F:("6<cӀD/r8h!"O캃iL$?�y�5������"O�e���)��刀eM� �|���"O"�A
U�)-��r��D'�d-��"O�Ӷ�m�"��!bN*K�p��"O~h�Qg�+��c�ʟ��~ ��"O ���E$Ay`�G��9�MA"O��i�Ϝ)bb��R�-VH"�J""O����D��o��(���.5�p��P"O�M��;��KV!G9��y��"O^�[%�Ԛ~�&���!My�Q��"O�a�g��ل��P�@9pV1�"Ov����K7+\t��,�''�(`�T"O���#fC�^�����%��/��1"O���� ;�KĪ����rE"O�l��i��i"�����z��)�"On!h��yMP���^a��U"Oj��) �/	�"#(�9?,� �"O��k4��)~:�𶦃�-vc�"O�� s�Y;-2 �4喃RD��"O�m1eKP�c4�B�51��P"O�<�6f��LW��&�%lV(A�"Od�Z�ї`�!C/��:�a"O�t��o�}f�1��ğ�j� Ёu"O�i�Þ #\�TÃ�F�H� �"OX���9��Z��PN�+�!�D�@k����d�� �rH�C&�!�dIv�M�����}��d,[;P�!�$Ե	�����p �E�y!���
����F�R�A��bI7J!��D
Qê���	C���!�ۤ�!�D�$`f����+>h���^t!���6��"N�GGl<r'��^!�˘f�`(q��_)X�)�VcZ?!��<6m��p��/�j���Ò4�!���P�Ag��t��	�!F�=�!�ʶ<�0�!J����� Ł�m�!�Űu!�	h�gZ�~c��CO!�䙵<h�Q
�f�i����܆�!�d�$?���!���cTl�(N�!��N 
�h$8P�Ɋz�UX�M\�;�!�䃆*��أ @ྐ4&��>K!�4@>u�d�hk��@r���!�U"j�U��$�L��
"	L�!���.N�`���X�L���\�{�!�� �`��Hk@�x���[�Z�"O����-�q׈�:gJ�-�Ԅ�S"O^�v�̂&5�R��ͩ-���"O�\RR�OXRQ��ܧh���Kg"O>%]�?���3A�Q�/��U`�"Ob-�4��XT�y�	ڢ6�0	 "Oz��G�0"Qh6O�39ߺ�$"O���B�͛T�����n�&͎uBu"Oz������y�:ّ��'	�T�kp"OV���ͥvb�C���f�����"O�]�tZPy� ��%W!�)����$ړ����_1����{R�Ц�o��'|a|�BA�(��كE�+2�@e���y���k촄Ig�l`���B��yr��.\�*�:D��)^Jp("���;�y��/a�:� 3��Y鰄�O��y"��̐��ȀR/����H��y�.����-J@�I�?56p���S�y�b�	o�J}b��S=B?l�t���?��'�Q�g	X�`9 �l	�4���c�'� <�f�:N�҄���
'��1�'v�3��'v)��XC|I1��_�<AAIȲ6!<${%/C�9�|,[t�v�<9��11j���[�� �hS�^�<d㍘?��<+�]5�: �G�u�<�ҥ��(��E�U�ӠXr.œ��A]��0=a�FO�;�t<� ���p�˒E^�<	F*�-O�. ��� ����X�<�0#�.�������H� <ӳ�H�<I�%2z���PcgU#1�����A�<� %�(���b�c�e�n�p4"�B�<��!��/���W�b���05M~�<�u�� _ ��)��V�{ ��3�eHQ�<���'�p��c
\N�#�K�<IA��0)����&�!�1��_�<I�o$���3�V�6[ʉ^�<��oW 5�*]��_|<���@P�<���^] ,tX �Ur�6�J�RQ�<ACLQ/l�.�gD	U�����L�<Qq떷���� JQhj���f�Q�<	u���3dIat	V�Z>ʨ�`�[K�<���B4o{\;�
 �F����FA�_�<	EV�$8�����xk��]`�<q �V?�̽##f�>I���˲�f�<�@K#3��	�W!��v|@Ѳ��G�<��Κ?|~�y��óP`��hpc@�<iWBȼfXa�U�줰�^���'&a|�H�	�Ԭ�3%�wp���)�y��N�$��a _�@��Y��
��y�S"&��E�ʹ~�X�.�%�y�솴1	B
(�l��P���y"��l
�t�MO�+���7  �y­ϖr�H+��XF�{O_��y2M�	'�\���W06�{a���y��� �b�0�]�G碹�!V�y�O��U��4*x�(�w�E�y�9���7�БKr���/��yrM��M��EU�-���JY#�y�nK%ZCD���I�9BV���Mڲ�yR/ߘa�Ԁ3�l\IŲ�9��y�$6��"6%8I��U�u���y����v��X�8�"�φ:�y��3f��I�f)B�����K�y�`��{�P,��D_�C)�I[�͐�y
� $����/]dՁ!��J�I�7"O�������s�F�$=����"O�ez��B_�1����$ui��'C!�ªEA����y�JhQs)�)c�!�D�.sZ�A�B'G6lc�T��W�g�!��T�Hɱ��X�-D�H�'0�!�d�B�e� F�)����f�Q�!򄆭��q�%@�ycT�
W��9:�!�䓿)�$�0Q�[<;��%.K!�D��k��C HO"&G�9;BƊ�-i�O����$�`σ]dГaC�2A����
�'�|l�"�.c""�˰NV4(�d��
�'�lpc�^�@��D���&/Z�	�'�6�����^���Kc5��M��'7�\@ ��6�E��2�:��'�P���,_�1 i����S~��'h�#��ײ(2b1K�mҗaj���'F�<`��El�R�y�O�*���#�'Yܰw�Y6/�ꌳ&kB�'�&�
�'(遥��T(<bVBG��&U�	�'����^.v�zI���ܝ=0��2	�'���a&� :z���6֐��'�젩�ʗ"��<B#�^+;���a
�'��\p1���h��Mӳ3o�=�	�'�4�p��ck��p�L&Y(&$i	�'�jɨ�''�xaV5X
�+	�'�.%�^A��)�J��E&�5�	�'�riq/F:.�
���X�R��e�	�'(���wb��Ii�02���G�8 ��'g��*��}@��ݫC� � �'�qpc޶-�
��R�J�0l*�3��x�ѹ[����I:� y�=�y�Y0^	T��pOG���&��y�P��9��P!T�P`E(���y���jٸe�qc��{\�	ɔ���y��W(5h��r�bR0{�"�����yҤD�n:�<��:w����W,���$.����'��p@����	W� =�6A��'�z}�g	~��\3�K�'9����
�'^m#���Ńb`�2 ��!
�'��-3���l�n�HY�)�(m��'	���ʌWn�|��8;��)�'������5�[�0���iR
�'��b!˚�򀴀0�WX�Ԩ	�'��tc�'@�c�jLn��H��	�'�T�"�A>(�t�XW#�{n�Y�'�@���,�?eS*�����|�r
�'���pM�uY�f�J �d�	�'s�13,44� � B[<��'�<4�2!(#E�sB�q32�'��ʦ�O>e=(y����iCZu؎��9OvM�%�������!P̼%jW�D�Od�D�O.�$�O��'<�N$�Z�^�9�&���e"O��H5+�$�Ne�f��9�� "O��IC�4>�d�+���U)v� �"O��1��<9v����;\���"OXhx�#�tD��j�
�pz�"O&�@��ǋatPUŉ 7^����"O�lӡ�» �Xy�g�G?$u��P����ڟ��	ğ��I�\�IG����=1������F07�d�����y�.�1*<n˓爉c�h�����yB�T�w��鰆�b> x���yr� mZT����lߜ�s��+�y�mqUD�O�.b	d�C���y
� L��bX��>�`�K��rU��qq"O�=�M�<l�AK�2%�u�7�|r�'b�'�"�'�?�7#�(B�yz�kU0]Y$4kG�%D�\�d� T�h� ���B�R�$D��󰁌4�����@:g<�QE�7D��F��_��M�R�\�"�4D�p�'�֬x�T`�N�	F�֭(Ҋ7D����ߚ=9��gˆ;T�U@D)"D�t����e|�1�B'�.�ЂL ���Ox���OR���Op��4�D��Q.�dk���9�h2,��<��Ð.|�xx�k�wդ��0��p�<Q�K�`���p�N�@Y����GXj�<��"
}8FjZ��n��v	AN�<i��#�A��^: �9x�b�F�<�'Zx,�(w�܊R`*ы �	yh<y��� [�,ar���7p�
7�_����?����?	��?�����)�5�F4�5HH�B��Q�ѡQ�!���}	@���J�@���ƪI5�!�ɥ�nݸQ��2$�q�K�,V�!�d�;>gz-��d%��(��&l��'q���bF{Z\(C�K��w�p���'��*��eR��ql^�i�p���'��T���U�s��2��$B����L>����?���?9���?1ΟxQ��S9HO�u�pǞ�_�ٙ&"O�����D�K�e��c����"O���4�X�� JE�><�J��"O
5cFN֙%��8��	�.�X�!6"O��E���zP���0!��	v"OH��gB����:!M=P(B|�P"O�eQ�/~�]3�䄋$�|�'Tr�'�b�'��?	���B�|��V*K;Y�졊0�#D� �0���*~��	���?���a��!D�|��-�~�@8���9*�\%9l!D�����U�/��e��n�s��ץ�y")B*J|z���pg�M���y���M�L4�T�� �N��#@Ҩ�y����v	�,ׁq�p��թ�y�V��f�/q�pt�u�X�<�`$�#�젲CZ+g��ڠ�[A�<)t���X<p( ����/q�$��j�\z5ϊ.kX�e�eS �:4�ȓN�v #q���V���$$C���T 0�Z��4���G'$�Ԅ�F��CJ֧Bdn��g)�%��0�ȓ<&�10!�9,hI�艕B��m��-�>��S��?���ʤ"���q�ȓN�M
צT<QD�K���6s�`��R���0S �f�R ��hʎr,Єȓb����u�ݒ<����h��<�n���o_B�6ȝ�!.�!�O�o���'�џ��<�W��$��p��M����wn�ٟ������w�[1����M�^b��ȓUa�j�G��yBG(�����*R��?` �����p"Odi�"�^�b�Nu�d��dB�X�"O �r��8%��p�eK�7(�`��"O.II�"�?	2U�L=?!XD��"O6)�V��;K>�k
^�{��-+C"Oj(�K�� yEC��0�> 
"OT�[�IC.,ɐ�Y��A5[b�}Q�"O��)�΋�0a��(��utJe3�"O�aC��ܲa�A����"Ch^3�"Oℛ���G������<���{�"O>��f�-�<�&�N�f	��:"O� �B$w�� '�=(�dH� "O�8�-:�N�a��S��T"O�@��'���~�kq�9U�D` v"OHM�Ly����2K�����"O��r$��<H�xٳPn�����"O$!�a,��ED
�0���c�L��"O41��']Y>������w�\�!�"Oֹ"6��s�씫��<��B�"O�Śh
>�x]a`��tL��"O�yq�% s��:�OF�!��dp0"O�|���D�r�D�CR�ޝC)0��"ON<�$�@�j���إ0����"O�I�Fl^s�f���./uT�F"ORT���ЀQ���Y�s ��"OJ|9V��-±�glQƺ �W"O�QRq&~��p
�ʐ�g���4"Oz��E��M ,�8�ʞ/
��I!"OP�ۄ�N(���� k����"O���Q�;$qI����$���X�"Of�`�͇$g��r�:��yI�"O�C����w�\I
P"K2v,���"O�Tr�I�ZqfUϕ�L\(R�"Oč(��^-T�P
E�\SM,t��"O�8�qk8[}l BnU6=��"O*dBu��4x_�P+�R�tdS�"OU��(��rZ��0���H8�"OxT*�ŕ�K>P��'�J�O����"O©A���2#R�x����(�"�"O��P7u��Ö[�Fovha�"OX�26�	�`#p�P�LF�,A�x[B"O�����	 �\A�W�Т:��h�"O�hy��V�S4�C4�Ƌ}<�[&"Oڝ���@�`b��8x)��"O�]��!bN�Y��9r��y�a"Ob)�2���Z��K��m�l-��"O�!ie��K7<$�5�j�5y�"O��r�[)Bw�٢���4�2"O�(h���4%�H���r��,��"OƝ��L���YqN� /�n8��"ODE�$�E�O��c.�(Y��UA�"O�Y��~\�-�4A0�P�"O�M��$(T.h@!�P�
��a�p"O���!�I���;3�� MD
���"O���!�
��Ttd�B�� c"O� W��J�X��W䎽T7���"O��X�@C�w�l��Ë�<�pUz�"O"�q���)5G�2&�("��t؃"Ot)��ӊ$�NP¦�\26��4K�"O�� ֮��]�\�@��B.̄��w"O�A�4�����(8Y�v�s"O�L�@�(@�����<�R�0�"O�	�,ȿZ���J�)f��}"O��$F�8a5hѨi�,Er��"OJ�3��֒dt�����?��(�"O\P���'^5�UIc1@����"O��i�`Y<�s╶q����"O4 X$H]�\�0�K��˒ko�d�"O^֠ �-˰�x�bЯ;Y���"OPu�;Eh���|F�A#"O�%[���ǎ�@6�!I�"OVɱ ��$��2'�?%�	z�"OB��%6dB@�:<��@�"O��Y��2G�Z(�1�6����"Oj�B������F��&<R�sc"O� \T`�HS.>X҄�Va77x�V"O� b��v�@J8.+Ra`t"O:}��/?��pcB��".��F"OD8sn�3E�p�)<�:ѯW�<ђΚB����*�-ext9�Mm�<yf X�s9S���B�,�2 Q_�<I�(E�A�x��ʩj^<�H4��W�<����<� jSiN�2~����o�<)V#�p^\0o�9E"�-����a�<I���#��}�*
5 /�i3��v�<q!��T�NQc���/'�Ӵ��yr�O`d�s��áYۂ;�"�y"���|�F-#�j�=O�pS��H��y��C�|����)P�E�}i��/�yZؕ���ɄB�lڳj
9d^��	�'��A,Q�Dʲ�ѶK��e�	�'�@��!ͨ��E��'vBܓ
�'Z�zӁö^s �3VEC�ͫ"OlI)����R&���r�ޅg@z�bR"O�#l��rYqr��5:�"O������9!$�9�d�2p!"O*�qEY.r�8a�b�J*�ن"O�Y0ԧ	���#SA�)v�eH�"O:]�2Mk -�5�J	��(w"O�t3�ο)Yt�;&&3zLN��"O@���"N�/�"��R8j�9`�"O�ժC�&o���B��H��"O ��S��+~>�ys��1��̳�"O�!��t���H�OZ�nm�p"Of��.#-2iz����9����R"O�UY� ��-p�qq��,�\��"O�Px�M��SV�jԨ��&�1Q"Ob��%��V<DY�m�
u���I�"O<QHY?]C����DXNx��"O���K&Lzm��A�S�"O��v��;Ո�ô��kX�"O����(��'Q�h��kas� ��"O��"�ϙ�.tIҪC�6_�QD"ON��b&��Lx������+%t�23"O<QH�fy�Q�A[�AW&���e���y��+R��)b+H+0��y��W�y�%�%5̦1�)@0"Ӥ�	���y���M��s��ڬ�g��y�Yz��h���� �I�'�џ�y2(��pM@����Ȟ�������yB!�!�T�Z�'B��#����y����HŻ�pL�" ����yb�*�@%��T6�(�Р�Έ�ybbʎv \��ֵ~r������y�L'P��eY�lW$��>���ї"O�5(rKS'd_,�
S�	�=�(!�"O��#��	-Fȳ��S�K�����"Ob�[�D�-�A����\zB���"Ox�����k�<;�VY���kB"O�(�s��:s��K���O㖅��"ORy(t��>\�PD�c��	�8�*�"O8�cn��(�XЫBN�2kԨ�p"On �gG�hK���#@�Q`��X�"O!�#�\�[]�廗C��=�L��"O��R�j�O����ռ�͙"O��uNKK��YS@��q�R-��"O�U4�&YUȑ &OԴp�H�0�"O�E�'	�wH<���Y��(Ja"O ċ��
�o��YXvL��ݘ"O� ��q��628��rRk5@�j#"O���aG�>�ΌB�*� ���� "O�1Q��~�����(�}�"Oe�V�Ɉ��1�M�O��w"O����72�ԩC���B�p���"O� dd�b�|1��x�xA��'.�੡f��9��Q�U�O����'�D�s�jIwC���ț�C(*���'^0�@A_�QJ�m�#ى>�q��'8���T�s��`���"Lh�C�'v��; �T>g���捻����'Tj�bR"ǽ���肢M=S"�(�'4x��"��13��9�'��D���'ܒ���N4�f��Ү�,�X��'��!�l)��}T��	�'�^��s@׿��P����1G�I�
�'��9��?u(0�DR1��'jp��1I_:���$c�x1L���'-� 0�	� ����&/U�pp��Y�'���Q���#�!���1#N���"O��b�gO%l��� F��/��3�"O��P��T��=��g �},�!"O���Q��&p�`x2r�R;Q�i��"O�Mc�	�Usn=0o߉6�P�`S"O�d�T�[Ot��d��4��ڳ"O��p!��2o8��
A悪!�4P�"Oܰ;q�B�l{6aq�E^�T�c�"Oh��HJ�}�J4�&�לM�Hِ"O4=kË?�$%�'��5�:�5"O�0�)[�4�<�&Lɐ{=Z��%"OT!@����u:lJr��w6&�YP"O�(R��<G�=��$/���F"Ovx*�#�/c��`p+M�2n�"ON�[��%�*(�Ϗ�;���ۖ"O �P�"^�D�酥B��D�t"Ov������(��2��aE��V"O@�ٱ
P:k�YY�*D;�l8Q"O��#�eI[t])3�Ȧo�vMzD"O�L�0(Ԡ�z��	IX��2"Opi�Qf�.W`�m�� Ut����"O>�+����	���#�a�"O�9$����h��D�eX�]3�"O����(�,p$у�¿QKFtcd"O�`G锗&�I˵M�ZIp!˒"O0�H�Ұ!Yr�� �
�=4n�F"O��I�BL'm*f9 bKW��T"O�9����Uy�q����&
�x�"Oz��� _�zg�<�BoЩc���k�"On �V�<���ӳgP��tq��"O�蹔h# i��'��X�$�(#"O���(VGjV`�oԐ �hD��"O9#�r���P�n�nU�ib�"O�=��d���DB��֙L�rs"O��P�T��)���+,*�)r"O��qP��*b��@@v�H�T��`��"O愰'EE�06f,QĮ'��`�"OB�Iw�)5��B@�H;@�^��"Of1I��P�'�P���v�|i8�"O�r�L��|��x����:crn��6"O�h��ʄ5�01���:I_�y�"O�L����<��P�BLA�XG���"O�m��Q�����%�653��y1"O�M��ݏS,�T��0A!��"On�����rGD krn�>u�� �"O� $qC�I��}���ږo r>|�2"O��aI�T{�hҒ��K�&�#"OtmY�U4�<��ؒ9���y�"O��$��y� d�7�
�^� ���"O^�٦`�1%:@���JߦȚ�"ONܠ�O�v6����S?K�Dq�"O������(����U�{���8 "O�QK��1�n]q����D��"On!�E��@m����B=�"O��q*�'"8f%8J�
J��
 "O�Pc㪙-*S���$��#)�F"O���`
Sd��XP�R�,�Lĳ"O�ħ؏c'�y�@��>}B*�+T"O��G��F��%,1iHX�眬�y2���J�8�&o�n<:��Q"�y�I�_��[g�!l��ջ���y��)Tq��E:�V��A��y��H�~9��"��",��`�JV��y"+�>�P��T�*g�X�@�^��y���5T���c�J""��(wiB��y�/�|G�y�B�K��-Z<�y2,�
#)	��?��1�VDǛ�y�À5��Q��ؠG�|u:S�д�y�R�N�*hkc�	�I�
i���yB�?h�@�!È�@T{�	D5�y��R�	�ց)��V�f�z�S&�D�y�kB`���\�/��2Ɲ,�y�h�2�!3�g� z"�)��W.�y"���n�x���.s�,��q%��y2�%l��v���m����P���ybF�Md�L E-׮[)�ف��y�*�CT�#Q��aĜ�
1jɸ�y�/M�Ru�Y�W���`��ya�(��1h�z�>3������^�z0�؆�%���I@W]8Zs̆�b��<��[��@#�,]d!���:N�\��ȓO�tX�$��J���b�d�4['���ȓS���D"E�F����Vc�+$P����~� MU�+A�5�,��-Ĵ���qd�I���H�
+��SC�ݪd�ʝ��)�������(�:ܓ���Y�^M��x]RP�R�_`d�3��[=�Ѕȓ���g�՟Y-$��`	?VO܀�ȓfx *$,��$(��� 8᪁��1�^R��V-��0[%m��rȆȓ���IBޯ~�P�%�R|���ȓt���)G�^��� 8S��,|�f�ȓc���eLŴ)���r��Q.L���#����e�W_ްqE^�@X��<T�-�%W�*,�Q�	�'0߶i�ȓyJ<IG'C"N�����8�ȓ.�0ׁ�5W'~豬�d�L�ȓpȈ���ݮO�0��$ ڔ.TlՇȓW�^8#��;�I*��	p�>��ȓp�E(Wcň"o�!�bG�t������
a��� y���9�K�w�R��ȓ*���I��W���A�{�f�9D���!O�	L�-ˆJ�y.��06D��kUk�%*�ٓ��"MR�r�3D�s�nYJ��0زI7h�Wo%D��s���UF�h�E��ґ�-D�[ʋ�`�fĊը��Ӝ�P��9D��Q�ƃ�n9L9���1`Ә� �8D��������y3�, �e�aD*D�� ��r���+Y�8�0�� -�p�js"Ox�����)t�̕�d�Us׶XD"OB�
͢u�6�1�^�d"b"O	����OH���Y�Ă�"O�*�n9N��P��U��|�R"O,�b���5��uj�A��S� �"O�4zbk
�&]�T�`����"Opj�.�O��X*U��4�~@��"O 2�'��]O��9�iƎy��X�""O}4&��DP�$"4c�!%b�9"O�����)h[� ���Ň$��"O1�%�\9�vݪ��;?�@�v"O9(6�MuR�������&"O��8��&|����CE �6�꤀�"O� ��NV�j�H�CR�Ytb�q�"O����\��t���A��aY "Ot��em�	^�)0���H	Z�"O�ͳ�B��v욇b�>:R9yp"O��J�&G?\\�{� @ 21��"O����؉$��F��Q4nš1"OV�a��1�R�Z3��#O~xs"O�����(���#F�/7~h0"Oꠘ�ǿ!��S��3y4H��"O"��!�ǜ`(}Z��?b�@y��"O�(8�
J�
�����T�Pĥ�"O��#s��s�"\)��	�d��"O�p�Т�bk|9"(�H��h "O4�ѱ�ι*w��#wg�>7�	R�"O�}��狫1r�hh�K�� ��"O0�LA��n���_�:�jV"O m�2��;�ܡ�&
�9\�=a�"O���l�"�4�dϽO�va �"OZ�0�٦6Hj�ru�]�7�V%YT"O
�b�:�"!�@�X<f���0"O��[v��J���9�0-��"O\Q���	�d\Ȃk�:_�F�(G"O����՞��|��G�t���"O����bϪ7�F��J�$&����A"Oz���*�Ti�`��0B0�)W"O\D�ᯜ�#L��)�1c����"ON��"�^���0#���0Xt�AG"Or�y&�j�PZԡ�_��"Op���AƏO@�q׉�%:��e�'"OD`5d�j)2���$K�p$"O�p(�t�E�$�=��p"O�)�b��	0��×"Ԫ	z�P�"O̩�D�
6-�sSaWb".���"O��`��ٿM��5y�O�Dr��r"O�h��I���\)֡o����"O��r������V�G%UR����"O�l��X�
đ"��$7����"OX5*��֦v����g�;%�}�"Oh���.B�`�\)���J�E|�� "Ob!��E.l1�K�Ay�!��"Od����WWv��Y�h0�(%"O�)��M�p%*A�7�ɩ��;""O��yE�I4{�h@a��]�jpg"O���A��H	da��<s�j��t"On� W�
�U4��Zu����t��"O��1�D���y�7��_���3"O��V���=��M�&�2P����"O�ȣ�
���T@`��q<�F"O�� @���I�&l#k2y�""O�4�2�� >�<LI�J�4)a�EC�"O� ������`LD:4��`�IP"O��vN��D0�w�O��X�
C"O���Vl],�&����T�bդ)�D"O4D����ܙ�ӧ��x@�"OP�d$�%¤qA�B=z.%(�"Opm���C,h�����dM6z�hrp"O\`9C��'O<�;fC"���qD"OP��!�F��8t�7`G	roe*p"Ob�K���p��a�s��ɼ=õ"O�p�F��v!3⇒O�z=�R"O6�Z׊�m舼5a2&yz4��"OZ���j�y
�X�Ѩ����"O4�����Xq�c��m��A`�"O��a���p���CU�"VA� "O~� ���Y[�P�¢Y)A���"6"O`k%�6�\�r�^�A|Ƹ�""O�dK�fغ��=ӡ�!M�Y�B"O�!hqĕ&��£`҅1� ��"OH�q��;���ӎL�e���kd"Oh����	�P�`�<L��@�"Oj@�CM߅D}�w�ȁ+��4"OPa� @=9"Na{�ΐ��ѹ5"O�e�S���V��(�P�.� a��"OR�Sa���vQ&�ۗ兩C+�1z1"OzEY�LX�E�����A�����"ON�:`�Y�5��ջV�F�"O���EޥM�x[�-G����b"O�xcq�ˏ8ِt[ cΒP�lы�"O����g�''7N$bBƠH� 4#g"O�Px4có$dh��f�|��`�"O�|�ag� ��\�1�\�S�"O 3�∳/�l=X�
ӵeF%�$"O���u$��5��si�5UHa�D"OX�i��!"z�U0�,6�$�� "O4�����3l{^	�s
��E�9Җ"OΤ۲l_�`��#	A�Ro����"O�I�.�'��j�蜆�� �"OrJ��"��
3H�.QZ�"O��%�xT8IE�,Z�e!�"O��C��	3b��D��jҢ$q
���"O���"�,'4@QƩ¿Z]@�"O8�Sa�BD�l��.�?Y��4K�"O�e����8s����+�(C����"OȐ�G�''�F�7��?��9�`"O"1�FP�nh��b�F�B�"Oz8a�L*�n�" b��L�jW"O����`F\�i[b��O{�Y:d"OLiaR������}pl��"Od�aÇ-Y,�x&�::ilQh�"OJ *� �;H"�)����#TBP��"O쵈%DC�_��a!�Q,@�NX*C"OҘ���4����(Z�^BD "O�4ь�<`�0�g��L.��"O��Iaę�{d~�05&K�%��ڇ"O�i�$�-s��A����/|Г"Oе��k��|B�Y �P�Y u�"ONP�R�T�)�BՁB5*��:�"O��BR��$�:\CS�	����"O�Pj�X�%=`��Aߥ�NY�"O>1�s�D�
F�x�e �#{|��w"Oΐ�#Ulġ`���'`�%��"Oz  V E<L����6O�0KU���"Ou`��P#H��:����X=@�W"O�u�NX�=X|��P�D�$nXs�"O� J����V��hY�4��1"O@�g�[�@�vh2�ē+��;1"O��0O�̑S��=͎�"O��9R+�-R����e��@�F���"O�a�҈<U�)Q����)�"O�I8����I[t8�0�䍲v"OB��g�3$_"�:Ƣ�9W�L�"O��zw�ΊPˮb˟���x��"O�q����/�V���X(5�pQ�$"OR�P�� �a�r�b�v��"O6����@�^(����[X�1Z1"OI �'G4�V��|F�h"O����IH"8�TL�Ag�wP��!�"O����NЫ6� ��&�3]f��"OR��A���`����_�z��4�"O�4���ߨA�R�pw$
+�¬ d"O.�hC@�VƲȨ2ɇ;��6"Oؙ31�L<Wt��I�MY�X���"Oꨱ��L4�*=a7zؔ��E"O(D�B�G��Uf�u��0�"O�h�w�[����� �I:䬸G"O�����tK��s��+\3tQr�"O*%��+�1(D�JP�D{���"O���o�"��l�aE��&"O����/�5$�D�#l�P$�L "O�|��P�j��q+%	�D
��'"O��H�+=�!�bK�`�*p"Ol��u�ѱzPDժ̛=i���"O���"��#Ħl2�jC�5��xI�"O�pP���q���hK�|JL��"O"�B���P�
��#��j�l���"O�� ��װHWv��"��H�&�y�"OZ��T�(g��ĳ�d�<�h��"O�XRd��>�0�s�;Ȅ�["O�q�r���0f�̚��H�QerȂ"O���E�X�W��8�柃[
$J "O9P�_J�@�Z���,@�-�"O�Y���'p�iZ�,��g�.;�!�d�Ms��;S���6J���e�C�Yu!��'@PIfCY�6����2FO�5i!�ֆ�qbV�1��� Ug�Y !��V#x��-����~���E�b�!��E�09���-vF����ɑ!��R�}ʝ3��Z[��0��H!���X��e����gp��)���P�!�$Zy�9@g�P� �,�"/K�{�!�';�8l���56�t����!�DS�a�F��ޞc؊9�����Lr!�)S���aI-s��,r"oӎF�!�䌃$+��CУ߱E�B)�T�U"�!���O�>��E,{T��9��X%�!�$�A��{'�'YH.��!
�B�!�$�({�r���.H0Һ��p%��!���;#��Kv�E���p��-!�$D{��$Q�ǀ4	Ÿ��a� !�!�D��]�Qp�G�[����bG0S!�U=&�Nkׂ��y� �!DD!�$�i���qR�+N�8	�@�a$!�DN�g9
��Vi��jq��'�!�dh*�����z�D,a%/��c�!��R��\�̉0 "��d�k�!�$�f�X�P���5c5�|�T��%�!�7!{�!ɯ'44�V��7�!�]	~�|ى1n�<x@~�)#B��!�� z\����s�S>D����"O����,�w�d�
wn�(����"O����C`F
�렇%��P9�"O��2����]h� ƹ�Ф�"O���@
=x���C�
�^g^��B"O�(Z�̟>K�v{bD-r�\�f"O��i�5\����͇b�\�xq"O' �,T�tT��6��5j$"O~9�� @�
z��S�"�xA"O���
�ii�r���-����&"OH*uGR���<%�9i��s"O<h S�SV�H,�¨	�� q�"O����"o��=��I�(��tqG"O���H��LQveR�JU�`wNU�"O���3n��#>�P��[�o:�	�"O�D��C *B��[VĜR:���d"O��K���&�	ғ"^�Y5@�13"O%��(ğw�E���)����"O���F�?���� Z0}���F"OȄ�Y�fU��S��AKg"O��Q5@\�A�ܜ8�$�r�\��"O�]
GI��8��`�*�;B�"O>|Z���/F��9ei�7~Ӥ��"Op}S��]ULH�r�^'[&��A"Oʕ��B� ˂	�"�$�&"OD��gk�v�ީ3sV��48{%"O���'�;R�Y�A��\�04K�"O6l�1DB!��1��E��'��I�6"O�P ���R�8�q$	�2x�"O����0�M��D@ {�Ҩ��"O4,Aw�ӿA>L
�ep��s�"O̐x0'��Z%��q$�<�@١"O����2MX��7B>$���"OĘ�C)��q]���¨�\B"Oj���nt�<���JHXh�"O(�Tٲu����AV�&:���"O���$`\]{��CO� �u)2"O�܀����Uъ|���pu���"O�k ��dx5���j�5b"O�3r��9o �]xB�W,��b"O�0K�l�1do�(Ksᑩu	Π��"OH܁cb[�
b�y�`��L��)��"O,��@�n�>h3g���(���"O�$����^��ȡ�m�8B�ܽ��"O��#��	#���C��
0"i�F"O�q��*,@8<ZQ�#�D��"O*̉w��)�H-�J���"O$J���1Q���5"�E�Fu�x"[���<�~:��=����  �L������f�<�RB�z m�1�ֱ/��M+$g�_�<�U*� "��僑�����)V�<I�a��.lL��ǉ+��d+��U�<����*�da׋�0�"��4��T�<i'@�3]Z���Mv>�Ä�=T��i6��[5qՉ�c�v�a_<!���6P�U����*|�.��R��\#!��ԧu���
t�E����vAW"U!��_5g��AwH�=zL;��?!��'z��h[��/v���Wk�!��F��	ےEX���;v���!�䂂;�<Q�AGت�~x�IPA�!�$�4k�����ȱn�NE��GV�s�!�$�4h����I�F��`8����!��Q��%/�,ovT�s�&0�l���� ��2D��T��=�e)D(H�J}(C�'���>z�1�� �)���@��W�X0		�'�d��_?�~0)��$VP
xˋ{��O
�}��hl� 3FY�pGLtZ�耠*� ��P}.�YыP�KZH �Q!�3��9�ȓYz&ؐpJX�x�%�`k�+Jޔ��Vmb1��nä!�p�҃J�T�ȓ���ڑ	�M�s�ܮ"�X���`�&� �	+d�I��͒�@�ȓ��d��a�z��uB�5Kb.]��	\�$� ^�2e���.�ahQ,ãJ1!�D��$��r�/����7��}-!�d��z^���3�[8L���B�N�}Ҝ��%�S)pTL���#�Ch!C�#%D�h*F�[�~tp�'m�`���%D�T���68��2&Ԁ�VQ���a��Cተ|	�Eb�^�*���KmҪwTB�I5I��L�6�/.nڵY@��8�C䉪CT�P��͡L�f��D��/N"C�	�r<� ��4wL	6��<D��B䉏!BB퉆��~��y`ELWMU�6M'�S��M�AKJ*W�B�b���S^L�2�
XQ�<9\�J�R+	�4)�$2���N�<���o�����ƍ6_�f��fMJ�<�u�v�� 1�P5�
�@�G�<Q��M\�[�"�u��Y�Oj�<��,�
�T���^�̤0/M��D�<	 o�q\ƕi& Q�Z
��T�ğ �!��Z����y�k��3ؼ͢S��~�|b��L��Θ�>m���YQ�TY�L>�yB��8ZT\J���;���hc�.�y�
4^XA�  �2�6 ����y�ă�	6�M�0 ���d�8�y�LE&rB�h5�W�(�Aw��y2툀x�:�
���J{ m�G
��y" <uh�aqf�F1�%�v@���y���`�<�F��'0t8���;�y�N �9�&���Φ3�� ���D�yǘcѶ9���Y:[}�5	pgݖ�y�N�L�\��C܇W�j�Sp�Y��yB
�,��a�‴M���Ԍ��yR�@��`�`E�(1WI��ʜ��y�E��8�T��2���<8
��#���y�D�5n5ڸ`�&԰�����	�y"���<�PĒ7S�>�˲�?�yҠ�1$FƄ���H�Qаn��yB�Y�L�}:��&)�[� ���y��"ytPU�ui��4���N��y�Ŝ?{c���ce����צ_��yrG:A���"�K��~����F�V�yCs�Z�2@,��I�M+�ʖ�y2
�(�X4`��2tT8�'��y��ϡ�����$1��*�@���yr�b�JuX�!1�6�*Ѡ�#�y��]92��b4����q�W�y������
0� �J4�u���y¨	�r٦9*��J�fW,"r��ybE��]K��;Y{hi�A��7�ybG�O�䀀�H}� �����yB��{�� S�����BN��yb�H�&x.Y�S��p
�)K����yR��O�4��bM�l��Iz��H�y���9"�p�6`��+�%���y�c��A^��i��F�nT��;U�8�y
� ���5,�9j�k�̧I��a��"O ��f�5�� �S�����y�*O��Thö��t#�悅/�����'=8�*q�R?UUD�rN_%�H�'�jy�g)���䂫!���a�'�Z�[uJ�)� #�-��=�x �'.��q�*�: �%�^)~�����'���@#�ܦk^��^4^y�UI�'�Z�Rf.�8U&�)�����	��m�,)S��F,'Mb��"%�]<h���&�P��=F�A���۴D�]�ȓ`�Ī���9���+�Ă:E�5�ȓ��l�7�Ĉ~J2 [���m�؁�ȓ.�L� F$*h��I**���l��xp���`��@[�K�#���ȓ��u�
3Ԃ�ʴ��#N:؇ȓ.�d��2��?3�lIu��*I70��ȓC�t��Q�K�8t�*��.t��)��L�d��$N��أ���(y�r��ȓQp�+v��,k(L�b@
��{jV��ȓA=:d���-	b�N��T�Q�ȓQB��Xw��O0B\ф�O"$a�ȓV9�Aɓ��

��m�Q>B���(�P�:�.�F��Ԓ6	�F�Ą�t��a`���0xAf�츄ȓO�����Z5y4��q|,��ȓ����0/�IkJ�pȞ�9�n���s|e���<$�M��@�/���ȓ &q��ۣo^zc��.P9�ȓrX<�R̟�~`���	�7��]�D0�Νx��]b�FF.^#����*@��"�)�hJ��֬8K���ȓ,f~Y[#�J�洁�Ș�8�PU��ZY P����9c��7��i�ȓ2,����[%(h��f�`����ȓ���H��oa")76�LH�ň�b�<y�E6]�\���6 J���5�Y�<)�N��!R��7��봁�y�<�7�� C�6�X  V�L3e�&�<�2J��U0�+E��0^�R2I�d�<q"�	�N��,Ђ.Uе��x�<���A*��	ֵ�k=l*�)P�<�d�L
~��S�3t�z�)4��g�<预>N�	��C��$)LYdI�o�<��'V�!���"�b�)#\����j�<A��ڭ-Q�`����N0�!�a���<ag��;zv�3�49�xG�J�<A�D�2{[�y��؎'Ȥ��Bi�w�<�v��w�`��a5�IS���N�<�DQl D%�B8D��P�`n�M�<93���!��4d�ƈ����m�<	f����Y�)S�y �K��f�<�u��� I�����+:?j��ˍx�<����
���0E��n��Wn��<A�X8h*� iOs�a�T��|�<� Q�uq2JU=f^zc�A�<)�`�Q��Uqv���V� �/�s�<9�X�-S�4���*9
�90oMr�<Aҹr�y�&�X�X0ţ�7B�!�ʌ*�q�b�U�d�^в��<�!�$��p�N��@���Nۈ@�W�-:�!�$	.]�x�φ���AA��S��!� *w�d�R�OM>Ӏ�y�AL��!�Ԡ��=��
�^z��GK�!�� n䈱n��HX��ޙ+m��S�"O��Y'J�)]*���
�3�.	��"O�0���Xl�����B84P���"O�)ɣ�ML��w�:Tm:�"O򬹣c�_�3�˛�~���"O((�"�FK�f��l��g� B3"O$L�3G\��y�-ͷj؎=ʗ"O�\��I?&���*V�T�U�� �"O���"���J��8&U�"O6��6ͣ�FL��it��"O*a2�R-(o|u�R�H 3��833"Of�N�/\�QG��
����"Ot�xv�H�ue��`@ǟ�%n*虧"Oj�����%jlX���W��,�f"O�-9r�=<���Aɐ�L�ݻT"O�ᯔ�s��Mh�ِ7A8]5�'�8�;s�	'�����]�xk�8��BӋ5Z
�P���O�8Ei�'���s�E�
����u\d
�'�vmHEoɈl�Xq8GFZ�ZP
�'~�)U�oCb���!�]�I��'I�%2��A� �~�R�3Qǒ(J�'L*b�P1���ɂL	J�����'i���E��Z�B�G:9��ݹ�'s\��� /=����-V�>��%��'���7�z��{��ܲ�����'�ʍ�pk�m������ $�z�H�'p,�Cr���]s�Y�q$�
�"O���P�bӆ0�懘
�m� "O$ݒ���V�z�h�f��5���´"O��KC���]�M!'\�*M���"OH )#$�
e ����E��(�>M��"OH��ʅ�_�*��v$�2t�R�"O�����ˈ{�ڰ�W��3]�H@:1"O6!�eF�1����@�ʽO��6. D�����R= <��"n	��HU+�$<D�d�4��wPb�	�P�K�=��;D��y҃�@���`
L�V�@�B7D����1^���d��(c�x��j#D������:'��11��7/�F�{�!D�8�Ba�z��Ĉd8s=Ne�r� D��A��8)tx����~���/=D�t��B���81��.T�}��@(�f>D�lY�ĄlʴuC/!TɈ��"J!D���t`�5a8UDK�MT��p�(D���E��,����j�a�h0� 3D���G��pڑ�B,�%C��g/D���F�Xr���([�EveI%A!D���!�D��H9bd� ׌�V�>D�4:j�px��@1�[$ y
�!� =D��vN��$�P����E,u�2 �� ;D���	F�"Y@�8���7&��c
8D���Gɿ�	h�e,V���SI*D�H�� ٬:� Y�8B ��jp�/D�ؚ�e��^2n�����&M]��3%,D���#b\0��Ĺ�"ڱlC��d� D���&BؖS�Y;�/č%yHA8�a3D��sH[0|��C�j��}�:�Qr�7D���iϽ|�J�����1)<��Ǫ3D�@��B[�a���&S*RT�$2D��t�@�:\�k����qz�Ƞ�1D�(k�C&�<4h1嗌f���'."���d����j�v�b�eBި�ڵ�J��,�<ѕ�ʈ��].q��K�?aI ͘�^8��J��� i8��V䌿�ƹ���Mm(<I��B�<W�IfᕸH0��$o\9v*�����Q���Ȧ{���kP��(��<��j���d����� 2��A>����!�Z#/T0lpO�)k���H9cG��m[n4�L�f��=rѬ�25|����F�m�Z�C��Ӟ�b&�Oڲ�X�O��%K�"ӪtC��� K$����'G�M�&J��@t�	�3�t� E���]��1h�*��By8 �Ҡ�W��`�u�i^y��N�EY�����",N� 9�yh'��k�h XrM�,8�OX�xd�_~����0�M��N�ם���!��B�R� 5$\�-��"Ц��l��
uӀ��*O���WcM�U�f�
���ѨZ�Vx�'�T�(l��a%*rK���)�OHѳ2A�*Yr�RG�Q(X�BH�爕=*d��aE��M�1La���B&Ɩ4�ȳ�k���P��&ʈ,`j|i �I<z�t��$�S؀��򩊐izd�#��S�?��	9u�I�)���W<w�:)�C���M�1�Ҕ"����7�'Ev,q[2
Z��꤉r�-	�4X��	���T��`X�ز@L_�P�R4�'��ɒl�H%6��*�{5���c�A1;˛6iE�WB���5}L90v�ػ�Np`Yw�|ɛ���P	���NC�W���P��JC��3���Sհ�%�Xs7��
<��us��'�m*3�4u2��S67�u��'�����OzW���3�R�~5nD���+���w%^(:�"����G���"!��'7���1%X�RLb�W:33"����~�"I�؍y����?݈2I�,B+,�4�ܚ����X(� �E���D�y�!ӭ�rt���Y��ad)�U4Ն�	=^����N�� m33�!5!F���<��	�{��y��_�b��yH�B��W������Q�&��V�R�;����d��wU�a�W��%',C�I�0���f�_�et��z/ѫQ���Z��^�or��CG�s��ju���5��&��jWҼ�Wc؊{�A�E�M�p��q ���w�<�u�ʹ[H���t!{�0���Z/[봼�E$�I����O�����e���XO���$aK������"
Q�F��c�+���	�So����E=�~d34�	e���U�E p�<���-g� �@O,ZkD(R�+S;���$�&1,�Y`o�n����
aj�e����d��vX|0#��S���G��5H�ص9�%�20�8�iA�S1�܈ ��Q��M;��|�ayZ�p��͋f�O8sAbʹOQ"�)k�8#�.�ŭԁt+�d����� ����3Y�V9��̷IU*�1��<�t��S܅pcmS�Q����?|L~�Pb�U�.ߺO���$�*S[�}��U����oIH.��۷
$��"˝7i.,xᓣF(�,M"U��3.��I��BB8;f6-^%K��0fֺl�Dh�b��	Q�'�<+��r4CÎ8ɼ�b�@�`X�S 5; ��L�(S�4�H�t> ��i�A+EJ�f�l�ƯO�K9:%*ED�cV���lb����4�R QBNA F�'���9��P�	�D�C�	M��H�#��%��)��4��hɔ�	&};��mڢd6�aF�-�j��O��>.�&�
(o�)c0L��j,��a]��<A��(I*�pʡC�O�D9#�39j���.�v ��ze��8�8pc�F��M���D�[�x��2���nnؠ�'�Nԛ5J��*t�Y�f ͈����8���Z��H<�@�_���HV�?)���-|"��'of�!��A�aH�U#3`͠>�h
E�߂X6|�s 	�52���!�?�E�G>��I M�?�l
�{R,�^�2)�F��&�nݸ���3�"d���'�!�׏=}ưkSl��]�*�� ��uWcΞ3�^c���	tC_?�V,dV�(d�mP��A4���S��@Cd��� 3�����߾|�)��ɭA�|1#�
I���;Q�Q�'Ӑ�:�� �6��l>!�js[�X���F2O�xfH�YFr��pÉ�QخE���'Gv�� c��P��䛀2��.�=Y{R�Y!��.	&� �Ё�(������B�0��T 1GX�|�f��.,Ѹ�bfh29Hg�f̓fj61XG�<�d��6���M�&s��!�2ĸ#*�*C�yz������[�P!�VI�4�ڒ�:z}L�E���%h^���~r�B��U%�@�0fȢ5mM�*a!���P|�ᒒ!��P�)��؎-S!�G=@U��HS,��;<e*���23!�$�I��h teňo�$m�G�|9!��_9�y����/*�(�AE�'!���k��%R��u��s3DT	o!��@�Z���� �0I"����!�Y�α+�������ɲTp!��3W�R�R2nL�#d�@X��	_h!�
k*H豴�Ք8L;r���!�DKH�D���{j�yr*[p!��""*� ����4X�{�jE *�!�D+F'��s�O�� �n�k2)V#!��
0���7�T�p�~"C���<�!�$�#^��
B��
���BӢ��!�D�FV��2�*D=M0�,�g�v6!��:Jv���-?ZXV�gr!���-!�
Hi����2���3"O�]pf��34���R���2�"Ov�rʋdѺ�x	y�l��"O6e�%~4B��_,+$I"O��1��U��i{��e�Ð"O� VȂU���U����*['`~�d��"O�D�u�7|�TY� _�FSFq�"O�P���\�� {%�3?E<e�a"O��X�IT-�����^2����"O,,�q��I&�LzdK��\��"OP���!Y�3�V�B#�$B��q;�"O�h��	**���G�9�"OT����V-s�hu�eO�  Ny��"O�
Mn�B4cđ��QSS/D;m!�6R;E�aGK�n��pS1��"r!�d�
���sӴ�,��m!��֏|Ӽ�X ��K�j4���3�!��Q�~Y8�v �d�"̺��6-j!�R0|-�$�R&�?�@�IvÀ�MI!��?�����I�E#�ɹ��H�B�!���Cl��C�g,
`Y��S�!򄛥fqH��]:)�5�h �!�Da�>�AECޛhͰ��!�!��P2)��h�oΥ�t�?y�!�
�I�a1�Ŋ�^<|ò��(�!�$H�{���`�܀1����ߑZ�!�+R���T��,5n��Bo�v�!��U<9�X��934��3��)�!�D�#��HH���W� uar��/�!��H�z���S�X5�����!�D��:nH�f��	r`���
{�!�ߕ�A�.�?�Z����M�!����.�����ȋ-}�!�G�/��@�`�ɨo�葹�i"�!�?^�B��̈)Ƙ�XRS�|�!��o�:H���L�=/���>+!�ڟa�1��EԪ,�QTo!�!��G3p�~�!��1X�5т�9@c!� �����6_������-x!�dL�+�)�O���w#C�$X!��8&Y��0$��-���V���!�"&(r����S
zM��^~'!�DY�qF��c�˅$����!� !��WsA��
�*��m t��P!B��!�D "H9j�Łub��s�� �!�]�RC�8�ₓ�n�f̓���Z�!�d�.�M�%Aڎ\�5�SC[ t�!�,8�ғÀ!�
�g�
�!�D� ���;P�:/��2A`��L�!�d��yE� ��j�[���+5Y*G�!��n�`i0���Rժ��KV�R�!�X=S�M��M1?�-�6KB={�!�$E�y&꨸��O���h�2�PyB�TL"=C� >BV�ƙ:�y"�|����ƥ��GPr�Bӭƻ�yrH̅c�AK[E�0�놋&#�B�I#iL a#��T@�V	x�A�n�B��e�v���i�8�>}��KzB�5+�paAɛ��ԔC3	��@� B�RƜ�B@Z;~��S�`L8,�DC䉴n�����.��AI4` @�M�-j^C�ɱ:1*s'H�l�v�'�K�
$C�Ɉ7zʼ��ɛ�|�8l@C�8��c�HȮuC��`�呲BZC�ɡX���9u�
1H:HL��o��C䉯0�v|���J:�9��׵)�*B�� &8�<�'ꖌ= �9G�Q�ErB�IFb��r3�N���WHȑ/�JB�ɝզ�A� #��9�A�?�
B�)� ����@Ur%���̴<����0"O@0�bM��$�
�s��� ���"OX$���S\��(!�>*��R"O�� O�H�))6m�Bjl3d"OP�X %�C���c��r&؄�`"O؝ŉ�%+���,
�^�^t�"ODp"S
��&�%�*�L��A"O^���Ĝ�)��`i^4K�)�*O�DYEl��9H�4��A�#�'�pp��j,u��s�e�B%�
�'͔��iƜTJ��K<XLj�
�'�:<B��]�\�H���#�^9�m�	�'�X3g	?�B- v Q���	�'�vM[�/Ir�|u��O�U�x)3�'a�勱�� ?²УጘO,�[�'�J	�炱@�D��2��>;���'�}3�aƱj�zX��>+*�z�'�܉��,TMJT���P�]��'���eZ'8"I�MŪP<\K
�'����� ��l��૛?O- �a
�'q}1&��{zH��Èx�@0�'����quN@���w� !�'�=���ݼyk�,�2 \�[���'@~���^�h�D� ��Ӑ���'�\�����m�n sb�i�T�R
�'Ԙ@ �V�&w��ZscO f4�@	�'s��h0�
*q|y겈@Q<lAA	�'�n=WdC�jFP���H�4J�Jq��'=��y����Z�,�.C�0�0	�'�m��'��(r`�Z4(>4���'D�-�Ӣ�a3\)@��ҀY���h�'�0�����m�Ri�!.��_A01��'J������P�:��1ꃢQ��x+�'8x}��J�'�<a@�D�Kh�@	�'/�i�9��]��ܘ~l�iZ�+&D�Pa�"��/TY�P�4Q�Y���$D�xp!(�s�|���Y�f�HL�e.D�pz�̔4"�	Y�│+� Kw�0D���A�RFz4�;V�1Z!�$D�h�R	����:tדC�hU��n/D���&��]�9�Vi�;e�^��� +D�h��Ǒ�#��L{��F�{	<��u�&D��a\&8�U�uH��ux���'D� ذ�޾_�D�8s���4��D���"D�|$FDH��
Q"Z��<0�i#D�`�Ƕ��;��qqn���'4D��3$E�jf%+r��7iC�2D�$�M��X�`\Hd�?�aðG-D�0r�@�yۮ e��nUu+��+D����$Q ?˦	�@	M�X!�,QÄ:D�\�4�F��<)��	F:�<���8D�8��S<\G҉���a�O6D�THF���*�Ĺk$ R.PB<X3��+D�dY�_+yy�LX/ 7Ԣ�6A4D������<� ��#��"~NH��.5D�����Cl~�x�9^�p�9�7D�h
'�/;���%N�8BryW�5D�xi�)�=]�t�)@(�4YJp12D�8x��E#F��!5(�*C��@1�<D���1H� ���j׸C3�ŊL8D�|H$Wz�@�A�&׈��d�*D�T8!
]��r��L�*K��W�>D�|i�ІPt�(��<a5!{e?D�8���_H�8钖��(���"6�+D�� ����=iSLD�3a��"��H$�|"!�#�����	96H|sV�0Z�Fʔ�"c�4J�J�
��	9F
T�؟.M�pgF|1b��U�i�MQ�ƫ��)��1���q*�2�n���� 4�� ��î���(d���ٟZ|�(� �j�B�Bv�O}����� �����!hF�-{ȃ�qP� !O�1�qI5dGT0����#w�9r�>#�H{6d2h$jyr2�� 0r���iӂ�p��OF���Ol�A3ճ^5��Ȃf�OM�!*��'�b��1EL4p��L�	�:n�}��A�r��T�ǭ"`2v|�%A�^d�
׼i��	��ǍJ�,�ቐ��kd&͙=�f��`)	4`*Oٸ�ASn�@ �c�Ys�Q�[(��2�,��,L��!$W.G"�U��W2$Ѫ���@v���1n�
	l�xxs� 6�",���П��fʆ�0�`{���1o�,iӎ��o�|h[s��6�<�ݻG�H	��f��`u~�.M���C≵P�}s���;�n����  <�9� [4Q�zd�#��#}�>s����!ڨI?��Q�'M�-` 	L3ݦ�p��#�J�؄�[%
��Tx�l�mX����	�Orщ��'慃��81�Q��X��l$��"C�H��f�4�t�bXG�ZpHvI��tj�Aa��I�L&@�8�-]:\m���۸.!O� ��6r[H,����s�KP���	Ģ>�F�*�ʋ	H���E�HC�q�����P����A�n\���	)L���J�it�Y3�烊�R��ᴟL�o�?T���O���c� �8�)�#AZ.�n��,���&�rTc��!򄓕8>�MBd*r�" @�]x8Q�ã_���Dсx��вsi���	"�n������Q%/����ݡ7�^�w}cw"O0!�d�Y/_~�Qv�\P�i�
��M����%�>��5�gyrE �*�����H�{8�Yz����yr�1'96�#�5i���rژI�[���jX��W~�|�1
��#�p�P	��Q扄�I�$� |R�m��{ �$�-e�0)-Q�Ul���m۞q�!���;u�(��2�ĝ&W ���
A��Cg����DI/\H0"�G];��	\�� ���Э��K�9%H���E��-=����%�'I��C�,<��Dռ\�F�+��N-�ѨA��3�IE�G��r�fh!3�� �L���?���L@<@�}z�Y)Z<�����$�$�3P�v\	!�	�?ᡧ�=L(�-e��R��e*ف�>�yG �q��q��"���X0O��r
�AWj�q�@�K�f`������*��h(W큦��Ot\��"	^I4��V �Y��,;�Ň� F7m	�u��2'���@u,�;��	1��98B�I�!Ȯ,a��ڈ��q��� }�j�K Q����rc��yr'�"pɛ$J7�2�i><J�kt�Y�#@��VMQ�N�>���ՀJh!���'��a�玘�6�����c߾�pM)"�DQC'T22|n���2���i�N�����p���QA^�<!"��X%�)� D*Βh��� r�V9���iB�fF2�9 p��c�Һ�0��98,�^1ܖ$k�lG�H��i0V�W���-ɲg�t��$ <����S�l� ��H���c��O���VI�-k���Ƞ+�����ؓ�ؙn��[!#16��;w�NTKE�ʳw�>T����J(�����~�{��B�:��G!��t`c闺D���)D�`�qPK��5�t�C�4>�dq�7
n�Q쩈P���Y�Gl�'pf���$�r�&���@���XW�1;���C�D���͆� �Jţ5%_�d(D��:�`�B�'Y����^��ѻ�cתc~�X��y�#W�b|�\�'l`<kg��O�2�2T�  �'W�w��iڵN���Ӊ��Px�"����ٸ�%Ҿ̴�S@���O3u�@�~��!���tܺ�5�ƕ17�SB�<y���/(u@�e@�5�$O�Q�<��+�5BXkG��(Cd�C��A�<�V�׶���O_�>���d�d�<��G?J���fJ�p�s7cFI�<��H�>?�|���
��I�؜ʐ@�E�< �ڞ=��C7��-��;�)^�<vNÞmuj`[���HR� ��K�_�<�V@E��R9`u	X#l�h�)��C}�<�F囗^.��Y`i���	�B�A�<���M&.iZUAӛ&#,5p*�V�<�F��07��r ��(�| ЦIV�<��"�	X�$%��J�>hj��B�V�<!���S#�<�`��-\���A�F�<�/�>�V���*o5��*g~�<ɡQB�I�f^+4���iԦ�u�<��a�4>PvܻэF"~Ǩ����v�<���RI�DA1.���(6�
r�<� �􀓥��^Pqˁ&��(g"O~�;p
(�x�k7j	j2�L�E"Oܼ��J�'���B+�S�@�"Od�I��މ��CT%�3���p"Of ������c�4C�"O��9w��'�е��̀Ƣ�á"Or�d)�!�I
��ڹVB��S1"OxAbe�+xlT�pо�Le�"O^P�t�� ]dN�n��ȸ�)P"Od�����@��	WB�$p��e��"O�X1R��:p�Bg����L8�"OxN�eO>|��H��,���"OFT��
ˢv���C��=W�Z��&"Ot�#�
^�i�zq��%�Vm� "O`�+��M3z%�y#�R��pyU"OV�2�)�83Jy������u�4"O����H�/i�����ԺE�e�7"O�u�-̙n���Y�V�
e*"Oġ�ÑF��d���ա*��lQ2"O�AB���$/^����]pCw"O�xC�,�_�@�y ��Q��"O�4+6HK;jf�tLp����B"Ov@2T�^4Ddqm�0�����"OĘ���0Pj�e�`-	��P�5"O��X����ry�=H
�[��,�"OdM:��ߓ.!�mȑ�ȝGr8��"OJ��D��4�l�� - v`��"OX����<A(ٱ�o�4|,z"O�XIm��	b�Ы�(�gT��"O�Q���	
6)�6�V1>@I�"Om�� �X[R%A�Ȅ*.tS�"O��!F�`m ���g�4�Ɲ�!"OJ���l�B{�X
�݌7N����"O��P����ъz�(Wa�`�K�"OlYÓM�)}b���d��ݒ�� "O���QZ�%�H衷��E���1"O��{��@�Q��\�X�b"O>�`�m�E�Rm#E)�,�i�"OЕ;��A-!�`$��5����P"O��s����"��`s ��"Ox���
�a��5��"�>x��ɻ�"O���2�MR�}�PC�-mĚ�S�"O��pwAE2*��jw�ǭ*�����"O����m��W�� �B����"O�AK�X+ ���K(b�0��V"OX�r֠F�uk�d��@��
�|��"O���6n��z��p�Uۍ^��R�"O�@"Ec�/\R\���Q��(�"Oj8�1�IIi�`�WK^�r4iy�"O�Y�/�-_}�eDX�M��� �'�4	�eҐ� ��((2M�'�T�[���1A�<�J�@Q#D�L�c�'�f��&�F(�U`ajзl���'� :棕q��ܰP�ׄYP�Y��'�D����˫;<t�a�K1HC�Ip�n-Ӏ(+�2�c�lC:�BC�����\#n	2Y'�$�B�ۤ�Z�-�/*|1�m��`.C�ɇO���� ��*��4@څQ��C�	@�@Iz���3���Z���n��C����|*dI7;��t(�cY{��C�8B�@P��7$w��[��5��C�	w�"� �.3[�th�F
R��C䉣V��2kI�w�m�F��}�C�)� F �dV�a��H��L�z^�!k�"O��"*C�O������?51ڤ"Oj���E^�
4�|����=��:�"O!��1xU�� ��rZ.%"*O� ��ᅛ&�tZ�)W�J:���'+*Dc��^%k
�h���/B.���'�@� PKU��$d��Y<���'jrc��Þ|�J0�F�)"y��'���3(�
���h!%�ZE.���'r�h+D���;1V� 5��r ��
�'���SՈ�f�"�"��
iFA�'���zP�Q2X�m���AP�Q�'�ܫS��B��i�D^�I_>���'��
�ˏ�|P�J���S>����',�գDJϠu�(���!LAx	��'�U�@-S�VĵP��$;�XiK�'���p���\�b8��l ܬ��'Yt<�"	ډ7���օ �w5��*�':�dr'�z��(VL�)y$*�p�'�B	"�(
�\}�h˝瞑�
�'W6ѹ����@y���ӡ���B	�'���	)��b�����/{Kv)k	�'-�p�B�l��Y"����iE���'GlaGM�C-(�U�i��U��T(�1�7L�4�C��ҥ~���K`�	K������4� @����<�$C�73:�y@A��c�d]�������ԹM�4eS��Ύx��y�>���g��ħ=H\�P5��LrU[#�	jN�'�ࢦf.���|rre�S��$y��6����j�P�ʩb4�dl��L��%�ܪFR^UH��O��-���ԤV Y��J�T`ʳ院�NI"q�@U�bt��蟈�įK�	�咦��j�����L��0� ��i�����0|ZV@�C��h�sc��_7���q��e�-9�+�f?�,�{nd��)V X������vH����%S�F�`nZ���]��.	���`B¨8�LȲ�g��9ᶂ-t��x���� ,*��yF�ߓn*��JW;Oa�t��YA^*�ňD�\ � G�8h�%��%?Ia�q�a��ח;��4�g���|u�gƎ��yDU�)g�@���U��<(��ڮ�y�O�r �Qزc(h���#��y�DB�-T�$��ι
�^�����y��<rT�!�܏x�~��!����y�C��F8��8E�6��+����9�S�O����@I@23d!@:[_|���'3���i��B�$�$�G��
q��'�4	�)�@[@@
�,+�BJ�'Fl�)T��p����eG����0�'=��𧩌�e����C�3�!��'k�q"$a�Q��a1'�!�5�'�f�����%�	� �
�2��Q�'�&e��n^2hĨ�:U�'��y�'����υM$ƈ�G���r�'��x�L͛-t�]�1O�%<i�'��	����11^:`)��Z� ]���'�v=���633fq�dK��'��� ��'����7o �PBR��	�'�,��*�t�zw�W�0��	�'�Ȁ#��7Tf@�SmL)1�΁�	�'��t�4�K�P!m��툩q�����'9����a6�2�11�ɐV�Z���'��A1�J`y^ ����T�V���'��i!4o$tzJ�0 	F؎���'��v��$;��U�'�ѧDo��P�'|d] ���6+� �C�+����'��I3��cIf\`u+�3�X)�
�'�vup��2.�R�2������  �!ਈ�/3艻�c�]DF%k"O�,Ҕ�J����QC� 53����"O< �HǂlX���Ѡը[)��`�"OX�ѣ�k*xx����yY�"O�d9'�ܚw�"�B�,A���"O��U͞[�<1뀱5����1"ONE�5� �xT	ny�I
F"O����a�v�PH$ȅ%=��ȃ�"OY�bN�-M;�511��&S�H,�"OH��˒�d+��`��\���D*"O���s*V$9ܼ��D�I�X�ʉ`"O�Xyӆ@�yJ���B?�N�J�"On ���#r������r�6�Y"O�Ɂ��sNN(@�H�ݰ��7"O��3-�3@��#��I�y��\��"Oj�r	F��q/� h��`�&"Of�H��ʑ33���.�=X{m�4"O�p�'/]�]^�m�R��J B"O�]"��� ��A��l�8yg2;�"O����?�V����6L93"ObD�c�� vµ���ֵ@�] "O6"��Y�{B�e��AI�qr|w"Oz�hlZRȢ!�e@-k��k�"O$=@�.#�8r��  "�Y"O�z`��{�贫�̀�g�J���"O��ѣ.��3gf@����"OhJe!Z$tr��c��!�hq�"Oؕ���#5�IL�!���"O��y���8XY(P�P��2����"ON�9'�K�V��,`R&�<N�=�"O� ����gr��j�'m��k��!��~�����nhQ���ѦtN��ȓ[��yA傆0���S!�&�����_�����"�����S��p��A0��%'_:P�ER���#���`�Zg቉V���Q�i��p�x��A2����J+V�v聳I�K.0���gl�ٰ��%g>�cg̔GI���h�:�Έ�G�VA�b���I��w���e�*fId1"§�:&U�5��N�n�3� �&a�2ɢ���[����Q��b�Q���I�o�<y�ȓ]=�� ȗBa�	q�$V�9����ȓJ��;�&��N����^�@��]�ep��a�Ȁ�]�j��a��FVH�%(�>`�X8�64�n,�ȓ|B)b�K�&�<�IU��X�D5��W�f�A.N�f�)�6?�4Y����L�x.Ե���0n��ȇ�b���Sn�?Ch�ԈW�cy�]�ȓP�;3��&�h9j�֧)A^L�ȓf��P��F�a��t��5�T�ȓXzx�h�J+���a(U������!X�Ur�d�u����~�L��8<`#uċh�*j۴
�j���\����6$ρg4M�$%�J�ꁆȓVSh r"U� �V���N�V�8��ȓnRj�KrEٺ�8���Z �ȓo�,Y�s��9ǒ�ˁ��>n�H���]���֢H�j�����lɽP�ڼ�ȓ?�e���g��)�ֳ\��T�ȓQT��!�J�n���S�^P��K�t(�pEͷW��1 �!H�$E�x�ȓRc��(�N�;$`���^�jх�S�? ���gdkw�2�P�tTD͙�"O>�I#��YpwG|8L0��"O�p��#�xtk0���{1ҁa�"O�hTNM���hD�SN`s"O��a��Ϡ#����C�=��e��"Ont�0 �D8� "ƒD����5"O��[4n��"�F�P�H�4u &"Ott�K�/F����ʛ�h,˦"O�����[:^n*�	M�@�=��"O�M�ᇛ�A��|3���
�^�� "O�!��C1V[�X�H�/g�ݸB"Ohy;Rc�h@L���FQ� af��"O�H4�I�_�F*�N�=`.A"Of�ڣ��Rb.k��@lG.i�%"OX;�N0��- ӄY��B"O�]�2(]��Тd֣A�4�
�"O��˱�N,���!����,��7"O�Y�Q��֤�b%�$�L��"O�����Q�9�ҡ�� �X��"O��1Pc̦.�lkAT%7iNA��"OZ ��ݸ0�����'RKf�xV"O���jU11����T/��A0�x�"O�h�p�02�&L�#ɖ$<8�&"O:uP��o�m�.	�x�(�"O�;f
 �/��]�c�Go�rt"�"Oޭ�`LM7}�lC�JE?��m 5"Oeڐ!_	dzi�`i��B�x�w"Oj�:R(W&k�f�H�(G�AhV�!d"OFYzE�-t�d�g�;DQ��G"O���r�F=zh�"lG#=ܫV"OX�� ��*\cP�5� C|I"O���GN�$���u(�|�8"O��J��H(j �c�οs��%��"O��i���+v�XE�N���AW"O��gä6K��ڠ,;�.�#"OHXs�h]=^:���#iۿ��xR"O4L�a��(���Ć\�F�s�"O^�)�/�#$�,U��/�2B��ؑ�"OJI�1�B6^INܑ�m=!��;C"OD�j�e��s�f|{�L�G|�$�"OL�R5n��0� ��3|��bW"O�԰�8l$ ��B!a�.��"O<�C�+Ux�a����<F�D�z$"O����T>� �ҥ˕�yo�,+�"Od *��R�6A��´PnA9�"O��a�����8�R��٩qV�E��"OV�
��q�^��3h��Z���q"O$� ���c��G�y��x3�"O��U�ĵb,^�U��(2�T�s�"O�cjɼ|8l���՗W�dhv"O�8��V,g��I5�Otq�s�"Oq'F�6Mh�1���C�r���"O�@ 5��:p`��ц&P��X�"O�,*�B�792��1��بF.��#'"O��{��Jzs(K�n��yplAq`"O�A�CJͯ �;�nZ3FF���"OZ�a�E��9n\���deZA
�"OX��gM�He�	 �=n��"O���w�Q,�Yғ)�\� �#Q"O�0
&�<=�X�UiH�X�t�p"Oju�C�n����HD;?#F��"O�)��H�+2���ȼk 
��"Ohj[�.|����3)���"O>���].5��2�.40튑"O� �ŉ���1yw�� #O(j�"O�@��@؜M"(��.H�'0i)U"O���6b�~,��r ��.v�kW"O.dR���R-;u/Ph�T"O2��7/B&U�1�t�\9r���jF"O쁣`�
�L9�E���
oz���"OP�W��0����4o��Td�ՠ�"O�t���͍0�A�dl&+QraZ""O⽉���mT �t̂�=B��D"O���EA}>��&��	{��܆�_w8��uj�=�q����<A���ȓM<�0à'�k}f��Ө@�>y�ȓ5��p��� g�*|�uI��N�ȓa�6u��n¶Ƕ�3���F�,�ȓU�8t�d�-,^�K��E��^���6qЭ�򄗷<�p��a�6�&�����L�#� #�mc����/�i�ʓH� G@�%`��� ���+dC�ɗk���FN�+J�����U^\C�I�@�& BJ��D��q���#r�XC�	�V(�ck�x��m����U��C�I�DeD	e�#YI�ips@ScY�C�Ih\�X��^�X�ဲLQ.�jB�9d��(�SFR% ��iT�.)��C�,vO�,�V�
�fS�)�7r&B��??l8uG�#q��U��AX��DC�	>�L��N� �U�!��u�TC�&;dB-������e����p�C�		Q��٪���V�<Es�k�� C�IAv��L��I�:Q�bc �B�	$<h��#T�
�Om`ѹ6eY�-�B�	�[c�U��׆]�$E��?�B� DD�c��D��-�
M�K�"O���C�w���S,�7��� "O���	ί3ΰU��ζd���"O8��D�B�#*�Es�KR$*���S"O`��$��T!�UpD
��<�&��"OR4cc��y�´sg'̤i�p���"O���wH��n�n5A%J�O���3$"O4%!��O�l9� ��A�3d��1i�"O�:�.�z��:��_/��h0 "O��KZ�x4�Өs7*��"O�|3�=�,��!���m;�"OP�"���:7>qpH]�����"O>�X�D3p��$*7	϶f�,���"O1ɡ熖y|R��P�b����"O(����̂9&��a�$���"O$���˙�FV���e��5>�M�2"Od��pĎ���$��K� ����"O�ͫ��+�hI��� e��"O$q+%g�$Ƽ�^-��mk5"Oz ��NYs�@�h��"J�;F"O$l��,/^��[*�S"O��S   ��   *  �  _  �  �+  �7  �B  eN  �Y  >d  9l  �x  ��  ;�  ��  ��  7�  {�  ��  ��  >�  ��  ��  `�  ��  ��  B�  ��  ��  i�  T�  ��  W	 � �! �- = G �N U J[ B^  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d�?��+�сg��:�h(+a��Un$��F� U��yz�rMY(P.؁�'2Q�@BۓRLx�b54�n��'�Л�O��@k�b�P4ir��g;D���HB �𸡆㎨5�6���:D�ĉv�%ΤqQ�-׻q�頑�$D����-:*��Yg�к/F�`BR!�II���'\+��0�e�=��d{f��S%��ȓnydP��La�Fe��6E����ȓ�u��
O* ��1��@��Z���z�	�F�^ #���L��"O˭o��x޴��?a0�W}����(Y�J�65	f\�<A��%9Љ(Q�ˋS�X��"�T[�<�/P�	U-zQ��'�>�J�,US��>`Dx��$�ߦr���(�Cu�ځ�yR/�2���"P��9s��i���\�y2�֓zwB#4��4�驴M��y�)��GX�@��9c�}z�2��#�O\������j��<P׊�$Jl k �'4���y�zm��f�"� ����ݼB��	t��JA�Ȋ5be��>[�>��U�"}�'�O�	/?o�*ny G²M#�)����9���D��/r���8zn���	J�2�qO��	8��D/�T?��ӊYʊ<yF�֤f~(�*�K"�dm�H��HAUĘ�^�nQ���Ή.�C��/�f]c`�?4LY�RoH�U=�C�)� ���iP�7�e�diE;٪̰�"O����m�$����>A�<	Y"O$}@'bU�TV�ȅ�ݠ?��m��"O�K�M|��	��P%.�y����f��i��ʍ��.F�:�<Q�����<��`5 ���N����z��:o����ej��4/M�t�4���� ox�<��	c�oPL�QgA&0RdIg�J̇ȓ��i��۵O��(s�\�9D'�r��X�S�'q����g�����dXU��ȓ0���1ed�xZجX�$�f����?	�BJo���I�12u�匔�cDԻq��XZ!�Y�� C�[$�LeH��� lH\����s�����J������ځnw��Z�,D���햨J��	�k���$xP%~� ���>2`$���f_>c�`��QGzB�~r�_.�����q�T� �v�<�NP+$����5��!E�\:%�s�<q�^C;x�ʠ�� }g�z�"�e�<9��]2��<�QDTLz�$ٖ�c?I�:�؈c��@*,���5�Ǣ`�~مȓ3�^��[48E��B'�ꐅȓǫ�b�ɾhE^�X�"ܱ�X��ȓl
Y��)Y��艈AD/y����ȓ>h9bWOQ�W*��n��_�@y���+�S���ٹ_s��AvK_{�D�e�\��y�i�7Ze������ i���U�A<^�Q?i(O?��?51Ȑո2�˷�U3W�����'�p�㣋7on�Y�g� �N=��3�yB',lOޥK�Kʊn��� �n�$��O��>/&1 F�:~�������v�!�$���|DCAj�(yq�4۔#VnџxG�k�O�0J%J,��X�N^��y���!�\�����hXW�T���"�S�O��Q��wp�tB�d�>��]��'��Ȣ	�uL0Q8�e�J���	�'�R����"Kp�% ��u����'����y*�;&.ֵs7�d+듹�󌱃��$S2��3w$4$e�#>���I��*����kGm\��V-X38+!��rH	��H0.l�ы�-5$+!�Ӿn|Ω��0\Q|x�-̝�!����*P�F��U��W��hʉ'gb�Γ[��xr	F�x�1�[%fc��h��,��d'O ��y���fh��D�
T��a:f�>)9n�M؟؃��E#�\�A��T����8�ə�HO��2�7@�r{��f+,r?`цȓ3��Y�«٬/SD���D1�Fz�'�0�Y�M#�骤��~8����'��U��@����P�fO5%���y��?lO��p�≒�TYJ%D.k�h@ "O����nL�>�0�kt��=-^!x�"Ot}Q�N�EYΩq �т'J����S�On�M���R	V$���v�ٷ����'�<�e��*; ��"�}��b�'e�#B���8:��"I�̉�'�
��� ��Bc
ι
p���y"�'`����1�6�bFP�
��	�'�*嚅.�K�b����8%����' L����Do��C�>�$�Q	�'�"!���*p��Y�/УF��ո�'9p���hT 5(���Ԧ�m]�q�	�'�(��(Ǟ��=%�j��0�	�'אYд.� "�Ԅ�kՖZ74 ��}���� ���ʟ-'~��{4эB�MCp�'�'fą� Cb�����&��b��	�'/�ծS-�&Y+R ׫`6) �4�Px�L+*��P�+��_�4�&)���=эyB�T�������mB����H�oDL�<���Od%�%���9�R�U1�2#�"OpXsD�A�41���޶lʑ"O�X�P,�����"ēc��Q�K4}��>%?)�<�_rƖ��4�A���X��''"4��Hլ0.�����}���m��I�O��IM̓ڸ'�,
)]�^l�U��87��3��y%ъk�h�q��� B��(RcK#-�qO^�GzJ|�u���D
V����B��=z'�Y�ȓ0�\5�I�H6 QB����\����'��x"E�Y&���F����X?�y��F���m����*ϴ,7F��yZy��[dԷ_�b �ƿBB�C�����͑�<8,ۆ���8��C�I�#�q�hʝ;�2��`�	>ϤC�I"I�H�ѶGƌD4��z�C�.{�C�/yQl�����s܊e�&jZ�C�Ɇ,�qG��'%XL�����0~C�ɇ��}�L=!���R���C�
1�䤁6+��O����"_45iz�'�ў�?������	M�1��$uTr���H7D���sח9��B��<*5�%1D��8���i��A��&�����)D��y%�����B�+Z�s����;D���Vŝ S)e�7I׆n�~L�a�:D��"�����b��3W�-b.�`:D�dB7� �9�5/�"3g�w�8D�09$䎐_R�w�K�(;C�*D��x�'���4�`�4>o�dR�'D�����6��RHR}-���*D�T���E �mYc�Z�:64L��n(D�����X2EQ8���N��b�ap�%D��;n^�>�s�=v���A��(D�x�E��?�X��E�V�'۸�pFj<D�(�F%�r�H�vē�H�~m�G�<D� {��D!��`�GǅJ(ZU�f�;D�\��+H�G0+�LFN�*�x �$D��q��T"J���E7���!D� Ac��.f���F)¥G��$��O+D�P� °i!���#�3.�<ɡ@*D�|q����
���pE9R�t�`&-D���d���Y���2�E� ����(D�0c��FE4\� A)C�Bs��SE$D��Ҿb�m
�a8QV�ɻh=�yl�Vz���ү�8�$�:��J��y�%Ya�Aq#���J��̍��y� F�ҴBVn��1�4� �nT��yrj҇U84-)��y�����y�Ɯc�l(ʀ�M�7V�=�+Π�yRN
-��qR׃�2�>��7f���y�ḭ{��X���0�t Q����yB��U`�!� zi��'C���ybm��z�����x�BL�3�6؆� �Qk��O���'ZD���ȓ �Z��NA�I%t��*�7�b�ȓEw�$��ڷQ����󃟇8\����n�ƕ���):hЁ��e��.��ȓ+W2����0ބ�d��4�2̄ȓ�����	�%24i''D�(B&���y-�����x��*�;k�Q��S�? ��TdM�+�=�BP�(����"OL�q�O7![��Ƈ�&FB��j�"OT�ؤ��yL����P5IU"O���1��-���C哒0�2��&"Ov)�U;�@��ݏ�J��U�'�B�'(b�'/��'���'`���U�nЬr`͛��шC��Y�K�՟��������ğ��I̟�����	��H�	99�(9�WeUa�`�R��ϟ��	��Iݟ$�I�h�	����T�#מ2=�T:t�X�I�^e�3hJ͟��	����D��������$�Iٟ|����N�r��sIα���Rş����	П��Iޟ��I韘�����W�@�v05$ڊQ�е1u�ܟ���ٟ���ȟ�I����	����֟l 7EA.Qq�@�j
03T fK���X�	Ο��I֟����� �I�l�I��K���-���0"I@E����W����Iџ��	����	����	ן����D��%�&Ex�8c���൓!�
��X��՟|����	�H���H����t	sM=fE6�cƈ��~��3������՟|�I͟P��џ �Iݟ������k��J�(*~ ��P;�:�C�$�����I����I���������˟��I���.8�г@&@=U��� �!��A��������I͟��	���������Iȟ��I�v��u��+U��h��R
�u4�$���0�	џ���㟜��ß ��4�?A�0Y����R�{��0��+�R�|�q�U�l�	ny���O<m���ZD��l��x�@��=�n��a�)?AԴi��O�9O��W����; �3qB���uL��i"��D�O\T���g������l��|�O�>E��hO������-\z�qX�y��'{��c�O!d]�֢ç;���&[I�5�r�u�:!�d�$�ӧ�M�;` �x�OF!}|�`�p(V�� ���?y�'E�)擦%��YoZ�<7@�4UYn K H��(�$�,��<1�'���DN��hO�I�O$����a@(�����lnj�٧;OZ˓��}�F
�'��ѻ��@���
�O֥1x�{��YS}��'��>O��z��H@/�:+��E�ʗ����?��K=<�|����O>i�ol�����ؚ1�0H�l	�Sɘ�.O���?E��'m
� ���*$�⊓F)�'V�7m�&\��.�M���O��С3a�{��8�'gN�I�"��'S"�'gҢF�<қV����'	o�T��n<���'E�_������e_pu$����Ϙ'U<�` ��8)j��q�����Oxmړ�8�'����ȼ<FV�3�/
�g $��&�M� � 	�'�7M
˦��N<�|1��0�������#V; T����}��(�X���D��F^����dQ��O\�g�ɋ�a
��|k`�B�,�����ɖ�M��A���?'`��&�EAы�05�����<�t�i,�O�X�'�6���47�̋b��7g��<X��K]�x���"�Ms�O<u9�)E����M0�i��Dc��	�Q�:��-�09O��OT���O���O��?��� �9Zh�� 9[o�{�/���<�����Jݴc� �ϧ�?Q��i�b\�ĐD>.�0,�m<+�B�Z�G����HR���y��	� �7Mg�<�	Ip9뵆Б'�X���.Pf*����Ի_b2��x�I{y"�'r2�'�RK&��m�Ԉ��6o�(P(�F�r�'���4�M���Z�<���?y,���;�n l��fV?.��I���`�*O(�d�0c��'��!�"O�f��%��:|�(i0G��P ��3��4�TxҰi���&�D[Q�kX���@X>l�z��������Iԟ����b>E�'�h6�	u�v�R���I��	1� :���On�dU٦1�IZy��'����M+�n�9`S�<��l�h��*��F�c�`Tk�Jy�T�Iٟ��P�����gSty��:QU&؁��4"4�s���yBU�t�����	؟0�IʟH�O`����[�|��M�e�ݾe�{`�xӰ๖o�O*�d�OВ�(������]<F���Yï˴�T���C-;��EpܴIi��&����Qnݩ�4O����:ϒ���Λ=(�z?O� 9���?�� ;�D�<���?A���*Y�*���C��^����U��?a���?I����D���ma��������""B�AX�	F���d����S�j��	�oZw�I'g��/eL0<jc�#p؄ꦛ�Lx4�آs�<�5lAG�q�6���?�0� ] XѲ�n�1���#dѽ�?	��?��?����O:9���ٙ=u�0iRKK�o���C'��O8�m�)v�je��ӟ,�۴���y��4[uإ2P�VM�8[��Ų�yR/}Ӫ�n���M��%H>ݦ�'G�pJ�ƅ�?q�E�(#y���@	�\[r���
WX�'Y�	ǟ`�I�������I.f��Ӱ<h!isB�(<��'<�6�45��O��-�9O
:r��7��%GA�ԭ mJ|}�lp�2�lZ~�)�S%RP��'��(NxƠ	�a����"
Z�y�z�'7�;F����M��+?�Ģ<a�K^RȨQ��)*��q�o�*�?����?!��?����DJͦy�Eu��{�K�	��çnlv@Z�����T�ٴ���|jQS�0��48n��'<��$�K @��!�(��L
�XR��޶VD�3O�!;�)I�FH��Y�O�`�d���$��*��� �KA��^�� �� jD�	#:O����O*���O���O��$��.�aμ��'eRJ�p�fM~�����O<��ɦ�
�r�t�I:�M����򄝑_*�G��vH��� k��O�pl���M�*�0�B�4�yr�Q7z���dN';�L����#�v���gϊ{b�Dz�4>��ʓ8zV�+O��$�O����O|��h��h���Wb��+nk#��&NrnDrA��<	��iQ��`t�O�b�'3�T�wF��R 
�;�	#ъ" �H��'�ȼ>Y�i��7�6�4��SH��P�V��[�|�`�K8�:����� %|�@§>���f�}Y��g�l��-O,�:e% ܫ��є�l�d' "M����O����Ol�4�����OH�/��v�I�f1����ݽ~�p�4c�%c�c�'^�l�r�O�)Zy��i�bQ�E:\4qc�u����Tow��d�#E�R7mk������pP�~�IP7S�$��H�'��dڧ�[$r��D��C!�M)O ���O����O����O �'v�ڥ$b�76�͸�#��[��$ҥ�i"<���R�����?�s����3�Mϻr����� (����Ղ_e��)'�'���O����'!��HS�i����<@�� �T/��X!/W\��
 �%�¿i<��'[6��<���?���?P|�S���>��0�u ��?��L5~�B���d�ئ��`k����ɟl�R�`��1��$ɇ7ߪ�⧇d�	ǟ���O�,o��MCH>�D)�0K� ��V#��k�	��#_�<��O5Nerd�*?��(O2Ѭ;Rb��nZ>b��:]`6x5�^(r/�KPET�TO�'��' ����O�n���j�QD��;����"A�)�l�ݦ��r�w� �I��MO>��3�/P�TX�8�@\.c<tĸ7`�\?�ڴ%>���'8��2��i���O��#�ہ;k��S�/~�[�nO�d�.L��!� � ��.O�1n�]y��'j��'W2�'�"��6��0��
ܚ?R0���J�ɾ�M�T!�Y~��'�񟎘a��6s*�Es�&��Uq*�E}��zӒ$nZE�)�:ZΝ����$�3��I>x4��.�=HXЗ'V|��q�8�M��.���< �P"�D����������?!���?Y�t�@�� �������a'�k�U����,�l�
Fҿ}���0#�՟�ڴ���|
�U���ߴj��'8q�ʁ�2�S�A�xE�V�	3��9O �$�� $P���2�`*O������%̐4����`(�j��9Q�h��<��?A��?����?Y��Tc&$��t�P�-z�v�j��C<`6r�'��d���z <�Z���ڦ�'��)�o�/g�b��Z�e��r����ēD2�vluӈ�	��S6�l���	�b��$���E8�5�Cܥ`͈l�BD$:h� ���r�'j��ܟL��ğ��	�_�ĸ�c��S@Z���Z�a����	ܟ̖'c�7��c���O����|:R��<pZ�
 ˏ#3�ۡ�_~rm�<����M��y*���QB,V���*@��ʈ7����L]�F��|*�+��M� �|���1]eP�ɲ�э�C�%���'uR�'����R��
�4(l��bG�}Q�tK�&���P�	 �?�����V�|��'�n�E��� �4"�1b)C&鶹��NT�&��6-��!��Nצϓ�?A�̓�Zh�)���	gm��G��PI �뵅��o���<	���?���?���?�.�>�ӵk5*�I��=Q��5�`(����������I��d&?��M�;?rV0@GU�A)���gA+@	}�e�i��6�J�)�.eB��e�l�G���QS�������uJ�Ir����r�t�IVy�'I�d�*���#�����Dٔ.2�')B�'�I�Mkq 	�?���?)U�G��H}��W�'�R��SIY��䓦?�V]���ܴi���|2�M4]���`�k\H����y��'J��� "�#��!83Z���~�6���?�J�w�L����b�J��S�G,�?���?����?Ɋ���O��ȇ��D>4�r�ݭ��!��J�O�Em��c��TW�6�4�μ���W�_ޤ��3��Q�9O��n��M���n���b�f�F~��O� 40\wMVe���}LXX�jK�=����`V�	vy���$N^XU��νu��Q@W�M��X�P����7��	ǟ���iǪ+��}� ��t� �B��4��I&�MKc�ik�O1��Q� O ?Lq	0��h6r��&	P�.��H�<���$Qf�ć�����D�1XC���s�Ƭ��K$�p�[���?���?���|�*Ot�oZ�)F���ɮ\�h"B � |�H��%��ZI��I��MS�2��>�ǻi,`7��}�u#R%���:��o�굈�	��#�~lZp~B"F3<x��78��O׊P�vM^��ׁ	�F�2�Tj��y��'-��'�2�'|2�i���5Kf�[2y�x�+���b�����O�����q��|y� w�ԓON��5��8~�A��M��	q��Ї�K��M�Q�i���-�,b��6O��U�v�j���l@,~v(�ҥ�JPj-&�:�?���.�Ģ<���?Q���?�Ƌ����֋]���@��R�?����[��k������<�O�0��@U�W���`�D�F���"�O}�'�6��Ʀ%HM<ͧ��'� ,�l�&�����	u9Tx����'��T(O���ڟ�?�S�)�dA�x�n0��F ���m�r��O���O��	�<�b�i̽!�I=QB���Ʀډj�����H$r�2�'�H7�O֒O�T�'��6�H�ZH�cg��Cd�@�.�7�0�o��M��g��M˚'���/z8��)t�)� � ���'/L\���S���9U>Oh˓�?���?	���?a���	�|ה]*��[)]Od#2L0LŬ=n����t�'#R�O��S������"/R�D�Hz$f�	OAԙ��d����.c��%����?��S�X��)oZ�<�r�Éj�%�ѯ�c���+����<�� �2���>����$�O��d��Z��b�%R!��Y�cүG���OH���OT�0r��E:�y��'�rkD���MÖ'��~RTӠ$�,��O8��'�b�im�'��#�
ĈtMf�S�hY�X��!z�O��Е ������ �i�����_ោ����J���X��y���w�Ǒ�?1���?���?Ɍ�9�:Y��"��:㴀�n��c�,�S�O<Do�>nZ��%���4���cF��I�DuI�/D�@ܶP��O��Dk�d�䄟 ���s������(�b�]3��Rj�2撝�'b��hܶ��|2R�`D�%�$@m� F�A֔p�ٚ���F�}Y���@y��'f���3K��>0
���F�:���SƔl}Rjt��o��Ş[�u��m/&]QI��#�x`P�nR/c?v��,O��s�aU;�?��O;�$�<�k�&�Z4kM���$Z)�?Y��?����?�'������xӉt���a�7��\���͊P@Q@�p���4��'��e��F�y�.�$��.͈��G%8O�\
&�{�yC�)��x���9�>d���qݽ����4�w��@J_+xE ���)��q��'�'��'���'�I�p��-iybɓ� ^; ;z�9O����OZ�oZ�-8�3��f�|ҍQ2,� ���)Y�O}�����#C�1O��D��	ÓZf&!咟Xcth��YwZ�f`��L0=�&}�ڬ���v�0�[K>Q/O��D�O����OnM:hs"X�"��$e�)�O���<�ipfdT�'���'v���Okp8���S96�YS@m-t�t���'��>��i�z6-�g�i>��s��c�?� �镋HL�JeR���,A:�p�Yʓ�F��Oz!(J>�Tb
%+=؝Q@��4E{����?I��?���?�|b(O��lZ�:[��DM�2nA�A�ب']�!�VJ�џ �	(�M3����4�2��'i�7�_*C~L�׮�.�dЁkU9y6�n��M���\��M�'�� ��w�re�ӗX��ɰn��"��I<E�ֈ��e��+�N��jy2�'J��'���'U>a�fI	%�Т2(M�M�&Ei�叓�MÇ	M�<A��?�H~ΓCܛ�w�^�P�$����0G�=���Z(�*}ӆ�O1��(��j��~G���,�hu�#h�fm{!N�LU��)xV�@ѼiQ"�'���'���'�
hV�ma�5k�40g>����'���'��U�x�4<�~����?��v�r��%��X��tŎ B�A�����O��'�6-B��m�H<Y�
P�p0 �� t:�Ðe��<q�l�Hp�jZ?UYh�9,O���*�?�1G�OX �J�8|-��rWOFd�(�`E�O0���O���O,�}B�"R
�����X���k��@�Z�$�J�u��B���D�Ȧ��?�;3 t(�c"�zN�`��A�Sr>��.!�F-iӔ�䁃|քб��	YFٙ���H(���E����s���4��`q薰�䓗�D�Ol�$�O�d�O��$�8ٌ����)���Ќ0K6�X}��� f�y���'NR�Oj�$�'r�B�R����T�܍�� X4Z&��M�u�i1O�D�O!#�e�|���"� Vu-�nO1y-��XpǇ"�򤓺=��a���'�ı$�h�')���P�.�}l +5�"!���O����O�d�O�I�<�6�i�jy�'<`9�0͛� �J�X���_��3�'^7�6��7��dIަaJڴ�?I��S$�*�Ñ.�:��*�@�z��5!��Q~���8!�AbXw���&?%�.M�L��H��MS�};t�_�Lr� E�4$�,8��ٺYS��(��G�d��#�K��Qk��{��Z�XZT�ۂ@�ezx�[�A� I�l��F�o�L�fԻ_
l��]/,m.��8t�!Ĭ�
�@��C�� �n!SG@k^Mzt�L �X`W���ȩug֣M�A�Š�l���y`�5KC���P�� ֋	�	��bݵa���Z8h��PΠ�kb�#t��uAҧv�a �J��1��-,nᘥ!%�#�Kd�2��Ƀ�H�	
�(�����x8j 
�E3Bdz޴�?����?ٱ��0̉'���'r��NSr�����E�v���3rEߺ��'�"�'���vA=���O��D�ON�a4�Ȩx`L,yO�1���/�7�O0�S��y�i>e�I韼�'EFEiWI�Jl�%�5�A����ae�.���?�1O~�D�O��d�<��Dƈf�*hZ"�Q�J�I#���c���(��x��'�r�'j��ڟ�I�q�ak�Jږ2���*�&F9GԘ)���<�� ����h�'�`j&�>]wC[M6�8 ��w�XU�@��>����?Q�����O��C ���Ɏ������.��XH6��?y��?I*O�$�ca E�S�# Xq��/�p�� �<^����ش�?����$�O���ԋo1��x���3�P�����I6�U
��S¦���ğ��'\܍�š9�I�O���ư�x4���P���0ዐV��y:ҵi��	ğ��ɛ,ߘb>��I�?7M ꔘ@0���$�b��'8]�P�0����Mc�U?)�	�?I��Of([3��2��\:B�W-7>����ij����S�D���43�ʬ��V�O`�pa
��R�dn�)F�]��4�?	��?y�������d͵���*��D>D}��!0)\�e��7M�%�V��?A���<	�e���;F>lM<��'�ڂA�0��E�i���'��BRnO�I�O��DQl�? �]r��r ��4�˾M,41��_����䟐�3�(�	����ߟ�TI�v��U�MO�L'�]Bs��%�M���>�8�顙x�O<��'���v�&�Q'
3'-@�i���W�1�4�?W�_e̓�?������O�w+Ɉ'���ie���X�̔:7�P�^��ʓ�?	��?A�R�'Q�񰆞?�
DX��P2c�2�)�ҷ�8�OP���O ˓�?�uK����h^�!f��f�)����)	�Mc��?)���'��iZ�q���aشiĘ��%�>~2}pd�-o�Bl�'���'��Iӟ��f���'I� (����#R�����`�����y�V�D(���d�@��}�O������L�#`\G�$��iB"S�<�	�?�X]�Oh�	�?X���B��)���[6L���q(T���'`bG�S��\ �y��vi�R���b����g�03`��7U��I�v�:U����X���4�QyZw�4|��	M�V:zePC.�h��4q�OH���GW>�������~��H��l�l��%-/�6�ۊ)S��'�2�'��$T���֟H�� 0̈́8�sM��)��I�H�&�M��F��P��<E�D�'B�ԩ���T"!MåH�:ѡ��t�����O��$�">���|���?��'u��!�MCR��Yck��;@%��4��=UF�H|���?��' �E��e�8}^��j�aٚ9�jZ޴�?Y�&@���O��D�OT�<:dK�8���/_w�-8�E,[�ɦS���CT�>?����?�.O��Ē�:�q��	�r(Z������ ��<���?!����'����/-c���&&pr��BD�l�2Ԃ�����$�O��$�<��2�.`c�O�؁Aqk����'ڼ(�����MK���?����'���+���شD�yӌӖ�%0E-�7��(�'�b�'_��ȟiңBr��'!�'
Z�n�����,44z�F`ӆ�$"����DC0�LO�"Ej�b�-
�j?�t���i�"^����4%��O���'��D��9X,�#�4b.y���Z���b����
JJ�F� �~�D�E�X>x����X#]N�i�u�b}��'�F�{��'R�':��O��i���7��g�Աa���=\�XlˇD�>i�UN��k0��A�S��s\X9�C�!Q}r�$��0��7-
�$1���Ov���O"���<�'�?����(T�6��D��?O��ʶ္E��ɚ%�"<�|:��H�<�چ(���r�-��=�"��E�i�"�'�2K�3��i>�������R��-��)ҴY�h�`�2d�j����U=���&>��	����#Zv��o�;[� �rj�R .�n�����Z`y��'���'�qO�A�p��(N}*!�ĥ\6%0q7T�Hi�F�Q���?������OR$1WFۜQZ� ���X�S��}���BКZ.O����O��d;��ݟtX��n�t�����=��i��8*�Z���8?���?9.O��DȈS����#Z�t�r�h� a��|�vkA�|.�6��O���ON����E�gi�l��B��j��`;�!JedNc�\�������'XB�׏l��Sɟt!® 8���c�IG
'"�(g��,�M���'��&���asO<Awhȱ&�¨9S	P�j4��'�֦��IUyB�'Ś�2$T>%�'�4�ش{�l�Q��!��l[��U;�db���ɀ5��YhE*9�~J�S���:�ߖG	��'O}��'|�AC@�'EB�'^B�OE�i�aITMN���x�g�Ia*達�>���^L�ꧦ�[�S�k��L�Ɖɕ\-v�ЖkJ�}�F�l��:��Ißh��ʟ���Zy�O"�d� \E
9��E�4^�4���mY,6�ёtCBub1���ݟ�)TBK�1pYav�ݼdNj@) Ɉ��M{���?��t0�/O�I�O�佟9qO\�Qؐ�B�V�7l�(��%�.�'O�m�!�3�i�O���d� �߀'U\�ل`��B��;p8 7��O
 �)�<����?!����'}��3ÂѪD�艒�(f�,���O�ݑ���+;�������Iny��'̐(�V�
;���U�ـ1��X��j��	ןT�	��?I��xɼ��Q��!u�^�C�	K��Кq�_)a*b��'���'��Iڟ8�e��Lڔ&�"i�R�3v���{��4r@&^妡��Ꟑ��\���?�� j�Xn�XX��9��z$���$C,��?)����$�O�E"P��|:�/�hQu��F�k2��s�I�Ѹi���D�Or���H7=��'Τ��!U%eS��(N+�����4�?Q-O���̣dS��'�?����EC"�(�V*-����JƖ[V�O(��ȑ]��r�T?��e*�#u6I�qI߾l�L�pǣ>��M�a���?y-O��I�<��`~�UZV�V�8��ǫ
�@Y�'�R�%Jb��k�y����H�r�l�2�Q�3��e%֦�Ms�,ڍ�?i���?����)O�I�O��#pb)^~�(���O�VZ��#����-�����e�c�"|��c��)�F��l�KC�
�Tq��i�r�'l��A���i>�����+)����tD�jրѣmi"�Je�Ěg�m%>9�I�����2����.C�[����ՉA��8m�џD���Ty2�'N�'BqO|���L��?�0�� H<,�83�Y��G8x���?9�����O�s�kD�o����US�r����I�d��?����?��'�(� � x�'Җ?���� ӄb8�a�d�Th�ܐ�'�"�'��IߟԳP*[fZ֫=oE�x��^�g)"Qr�)U��Q�	؟T�I`��?��4+
hm� :,La:  Uw�ziI#�к��7��OZ���O6���<�a����?����~�ϣU��� ��	x��cH͈�Ms����'�R�̥���O<����
a�h���
����,˦���Oy��'������O��ꟸ��4eC� >n�ɔ�-V�8aC���D��?���ErJ|�<�OLJ	SW�W�Ǵ,�TdE5-V( `�O`����*����O����/O��D�d�����e��|�A���I�Y��I⧯#j��b�b?Ӧ&W�1��@A�M�P�BXs�'{��\� ��O&��<)�'��4����H.K���RfX?\�l}�w��5�0o�����p� �)§�?�7D^�(�P���Wl>��0c4Y��'���'O:܈vR��럸��M?ل!&M_���c�mG�L����/2�1O�X��GP������	g?�v��<WE�P��J֟h�.��,�I}rj�U��	��p�����=	���g�(�� ��"��9Au�F}R�5=����O��$�O���?�&-�`5*g��Urr���d�|�ꉉ.OF���O0�$8�I��s�l��FE�D�r��`��MiBn[�lhՓ��3?����?)-O2�d�\�(���)�� u�Àh��)qm71#�7��O��d�O�㟈�	�1Y�p+P�u�ȝ�JP���%��@D�T�-(�]�|�	���'#��O-d��㟀`��`��+��ݩ��H���	��M+���'$B��iX�=`L<I�
T�|�pؑ�G[�L����Q�Q��[y��'{~aZ>M�I���J��l�Ǽξ���\^g�H�D'��ٟ( ��3Hb��'L��GnZ�[ ؊�Ҍ}�8�l�iy��	pj`6�O^�D�O��I�L}Zw�TDx@A\�O��������X��4�?!�!2͓O��۟��}bG+� U{�|����F ��G�: �G�?=�87-�O����O��i�g}"]���,Xr� �l"YH�Hcᚹ�M�4'��<����D"���� �O�&@@
�����YRd��M���?��c�E�\�@�'G2�Ox���_�Y��a�F/"/�^H��i�"[��3B,k��'�?����?��R�+8�3���}�$�*B֭Wɛ&�'� ��6 �>!-O���<)����d64���I��iG�$YPLn}�ǆ�y��'��'��'o�ɀ#�L2��İDv��"�dVF��a'͚����<Q����Ob�d�O䈠���&cz#AM�.̬��e�)�d�<y��?����Đ�RYv1�'/¹���
sg\�B�[��$mZzy��'�	����	۟��dx��s���dOĄ���R�l�0PI�	��d�O��D�Oz�-�X�]?��I�dN�!���C��������L�9ٴ�?*Oj���OP��Ҏt��D�|nڮ4��b�Ze]�x�҄�?��7M�O���<Y����՟0���?�C��3d����Ìt��hT �����Od�$�O�-a�6O��<)�O.-ل"�s����Aܾ@�����4���8+�n�����ڟ��������Zy���[�0H� �G�0�8�;»i��'���;�'N�	ß�}*��8P+�����@xLh� c���Y�NE��Mc���?����A^�Д'Ođ��*��R�8:�&̪7�d���t�L	�?OڒOX�?��I�|�bE�C�ʁTR�1k��tv����4�?y���?`3*���Ay�'G��T�AN�����S���)Oܡ	��F�'w�I$���)J��?��AN���N�5? )�B�FQJ�R�i�,��e�듯���OR��?�1X5@l&�%)D����@�?=%�'eŨ�'b�'�'�2P����=�
iPd�ƪ0���E"A�r~���O@��?+OB�D�O���:5����.X�̌+�^-���0O����O����Of��<Acm	 Ni�	)$G��+@�E��r���{��6T���Ioy"�'��'�����'G������;G�Rl�C�)K��&�v�����O��d�O�ʓ*����E]?-��>Bo����� v�-#C�*';�}��4�?�*OT���O�$F�Y�1����ʬWj��)&�I5=�N��B坾�MK��?�.O��aek���'$�O�^�!�I�k��L5����7@�>Q���?	���^u�'P�	@RӂǠq���q�/h$H@�\���'DZ-Hc,b�x���O�����|Hԧu�D�p�p�X7�DEˆ
���Ms��?�7���<Q+O���/��a�d�"�_wpt���ؒt�7�8&X�8l�˟����S�����<	� �/p��HceG�A�D�@A_�6S��B��yr�' ��x�'�?��*Fp��@&l�"2���q��@�PG���'��'V��+��(��On���d0�&2����Mو/j�hrqb�ޒOh ���O.��Ok�] h��qҥN$�}�9u"�F�'�^)��L9�$�Op�d;���zs)�][�E)��^)�\�!_��q�a��ʟ��	��'��|@��� �`�O��^u0�&8$��O��D�O$�O��d�OJ�1�#�T�`��$^�2В5�؎]����<����?9���$��&�X�̧�  �.� T|���#V���%�|�	hy�'���'sFI�O�ۥ�=~�� 
��
L�4��5]���I�����oyB M(@	��t�2u.�L�̓AX�db���A��p�IßD��z��	V�� <�0ChV)�r����K)Q-�W�iB��'8�ɨppp8:L|����C舢fx̐�M��M��躢��C��'�b�'t@
�'��'��I-~�6�o�#4�����Y5Gw��_���e�@��MkuW?���?UC�Op,��`(lh=h�̈#����i���'���YC�'Z�'lq��$�><���Sk.{�Q�ǵi�:��'�q�L���O�����0&���I�,��R"��L�^�8�kA�z�@�k�4������Z>��'�HɁ<P5�&2sI6�����,6-�O���OR���EB��?��'��<cVdZ�Ԝ�U���@�(���4�����C���'��'Θ�;�U�Y�%p�"�H�c�&t�j��F�"ϲ�'���I՟ %��/��E� �ð<��U�����.�o�����d�O���O��pV��Ñ�$�h���\��-�u瀕�}��'t�'k��'� DC�"j�6�zBn�pcd�bK�H3�_���I�����y2���VX��S6C�>m��B�@�b�b�c��듆?������?��\t$���D�i �{r��:�H�06G@U:@^� �Iɟ���Ayb��%\��� �D�Ǥ'}޹bsH"?���������E{��'T�\r%�'��i��0"�F"���b%�	|p=o�֟��I]y�,&|��v��kLɹO�W�
�G}���T�?zb�O*���8�b��5�T?9�V D&t��1�@��'uϴ�;��g���O�l����O,�$�OZ��㟌���Okl�uJ����á? 6���	Gn����'���#��3�y��4L��P �!-����NZ�H����4�  �]�ŉ��?A����X��OBB���ޢXSn�@��Ѵ
w�1� m��Q*0+(���?I%��	{@N��$J�{����&�"Iw�9�ߴ�?����?G,�<�?!����)�O��	�J�$,5�Q�D��ݰTM���jwN-�ɯ���H|���?���c^e��Ս>��1u�����ֿi\R!ߝ1��I�����OH�O�����L5��:����/�u�5�Sx}2�OT��ك�O���O��d�<q��T�{tP����z�٤$C<|(���P�������	ǟ��?Y��[�h��<"��W�F�(�!�C��gl8JN>i��?����?a�fo�;�OϪ����B`��^��A(�Ϗ)�M#/O�� �$�O��d�mv�����iT�q+fH�.�j�`�I�"��Z�O���O@˓�?���?Q��?�V��l�2l{��MޒR`��0z��'��'���'(�l�P/�-�ēl#`��0\�֨Y2蓿!��o�ݟ$��Zyb�G%��:����@�F�mD%���;%��#De�R��͟t�	�Xj�"<�O�*����J�观�?a2�;�4���'"�o����	�O��i�p~��dm�� w��DI���ReE�M���?�R��M���OKxHȇ��KΎl�S'�#�v�Pߴ#���T�i���' ��On,ON��E�0,|bR0��!h2S��mx]�#<E�t�'%>���	�&æ)&#I@,ѡe��$�O>�$�;�˓��	�O��I�l����dDˆb�h��W�W���c�L��#'�	�(�I蟘�WV�lO���SA�!M<���!E�2�M��.-&���?y�Y?��	a�	�l1dP(�l�7���T.M�J�S�O��0�ǐ���ʟt�I���'L��ZA�\�L���7-˶W*t��c_;�O����O�D#�	OZ ia*���^����`t��`8�ğ�I۟,�	�l��*�w҂�@�КLZf��1#@�{2-_Ŧ�	ҟ��	l�Iҟܔ'ԕ��4T8�7=a:pA`�#��"B�\�'�R�'aW�`��j��ħ�qS��-�D��O
�5k�1�U�i+|��'*Bf  ��'5���S��
s�\��f�z��(ڴ�?����D�-z<�%>a���?���8.�$9Y�j�$C���C�S����?q�K���Gx��"@�F�S��`�IkwVةd�i��	������4V��Sǟ��S���F�H5�:��9�K�FC�o���'����O��, S�C�lTL��lU� EX@���iH����j� ��O��蟬Q%���I�J����� 03> �E���eb� #�42Ͼ�Ex��	�OZA,��mX"�ķ1c~���;^�n�����	ϟ`{d�ˠ���?����~��B����A>E���a����'1�Y�y��'��'C��y�B=g���`�G%Hp�c��l�8��ͮ$|�$�x��ß�&��X
e�X1���O��P�ޞ?��ST0u�=)�BG��Ja"]p"t��X�$����@yp�I���\t�	��BD�E���KUj����Ϙk	Z�:`�]PQ��tŖ**��6�D-��ňu�
?AC�(��?k�f�k�m��2��u��x� Aӧ샻<�^Y��@�W3���4�)G��H*`k�+�����D�(�q� 
�H�.Qz���%u��!��E�9�t��נ,�,����I��-"ǃ;f���s�MͼG��x�o�KQ�x��!�9�	��\�q<�1����E�t����@����=�r�a����X��4I�1��ɀ�4���7�W�)�&8��3�Q�B��M�Hhx�������9���/����D�#�`s��"G�J�K"��X�Q��5n�Op��!���y	6�sdGA"[lD��q�B�mc��I|����	�%4�P%i$-�����>�OB $�� �z���5͜X����j����=O�QFI`}��'J�;]=6��	ҟH�ɥ&�&H�B_i�h��˒]�`��̎갽�ՍϢ��q��S���'��	  ��(��)�1vK�x�oW+;kN@!MΒ%��*Tb�O?�D k0q��i����X����8����?I������|�cܩl���F��w���F��:�y�� }F�OI�g.|J��$�Ob]Fzʟ�8*��	&ĕbF�ݤ9`\m���O���W'G�8r��O���OZ�d�ĺ{��?�p�Q�
��Zre��[���DfU�; ��28:	æN��x
�U�g�'���"+'0���'\�/��t��OṚ �+Y5�P�ܓ����$�	a�%���'f��c0����ٿG��'�ўԖ'�$����Z�#ꪐ�t�sK���'0V	��6lE��n��qP���*�S��R�d�'n��M���Ŷh�Bژ3~`�rG���?1���?��o�������?9�O,�}�eh�+�L���	C[����J� ���ۀim$4A��'HtA+f�^dȡ���^��d鈀���B$MX .���A��'���
���?Q�eL5w�8�s1�H�|T�&f_��䓆?��������ȃ��8���:iɲ�Z���#�!�$8$Rڽa��)?�fa�!��Y6�Dd}�X���e�Ɔ�M����?9,�35�;mfh!����{?���P��/$���O����=J�����&�� QF*OL��'-��8 ��	���������dѐl(��a�Q��N�q�k^���)�);�p�Bnģ`v�K��
�Q�x����OR���Ot�$�|j���#!�=Bc-߅9��Eyh]��?���9OZ����,F�nq���W�uH��:��'BDO��дl��,����G��#;d}�E4O@U;��[}��'��S� 
���I͟|�ɹS��! ��i�V�`u�ثL4t�+J�r>�X1�툐c�T)S�%ɽ���.����4���^o������Ër�αb��#�:Ո��/)w�a�JзbS�F���V4]`�K�T�`M��%��p�i5 ��?iӼix��S��?�'�|Ar�G� ��h���?�m�
�'�20`��-v<ܸ�$�D�])��H�'�7��O��{1`T�+ީDj�(yP�c���O��UB��"���O,�d�O|����K���?�"�sBY2'�F�a��0gĊ��VhH��D>��b�fOD H����HO`���B�;��m�AkN7n)������$6FJ���ԍ+�8���2m��!ғ:$8��X�"��LR�J/�����c���Ɇ�M� �i�O�OW��$j̵Chjɲc�,V1����' ���×�O�04��zBf#�o&� ��I`y�Y�d�7m��݈YJ�k� ��`�[�H�\���O����O0�JSM�O��p>]y������jA	U�=J���Ǩ�oЭ�CK�R���H��ՕD�tD��Ò���J�$��n��J��ɿxR�l���;�j�@ƶVxX���	>NJ2���¦���[C�J�iŖ�IY|�huJ��M�"�"��<��Ҕ�T�����1�x���QW�<�2�^b�B��3�J?^~<Hx�L�<١S���'�F�#�e���D�O4�'kz��S��joj-�	�?m�xM���C��?����?Qv��)M�����POD����K�u3$x��c��p9�/P�1�Q���KFBUdX�qE��?m��$>)���Bu*nJ4��3l]4Jѡ3ʓ:��I��M+��i��Y>�j�@ #�$��]XH�#�$-�-��L�S��y⎁�r�ڰ	F� ������$6��|���x2�ü0�ܸ9wO9��6�,�yB��'X˶��?�-�������O��d�O6� f�91��DCc�R�P����W`�F��B)Z�E�k��M�Ou1�2L'&S�A �E�� �˅��)+CD�kq�p#�����\O%�1��>T�9���;.�<��K4���:�o�(0R7�ۧ��Cp���o�؟PE���i��t�Gg����Ya$NڨI���̓�?�	�^�2�� Y�,��@U�!,�Dx�k:�-,ҵ��Kc��ڡ!�<"�E�Q�������?�%�ML�Y��?����?�A���$�O0���h@��n%{�G�S*,`i��O�hA�����*�'��I�`�Z'l��S�H@�x���'�(� pbي{gzxϓ.k�M�D�M�V��`CĄ� �n���N�؄��?��S�'��X�pJr(�Y��At�Ո4�hpP�&D��kDn��Vd�xh֮V7�"A� 'F�HO�i�O��(9Ɯ!Ǹi��1�G��V���;MƼu�P�[��'92�'�"&���D�'�󉎤Cҥ!��'����`��u'���dNU>}ʼI�	�v�,���C��d� l�%nT��A��O�3�{�-&�O�8H��'c�+�F�u���/�0`[���E��' �I�D�?�Oe��)7�%b#D�D�;C�@a�'��袀`Q�P�s�g�8瀬3�'������M,,3��mZş��	j�� �#V�Y:^
H��̈�n�c������$�OL��� �h9�`L�lf��S�4��"�J�@ȑ�(�<xJ+�(Ob��	0ߘp����0�P���m��^�q��7 �Q�t���O��$+�	�O�� �@�;~��B�H�!��I���O��"~�Q~8��"蝄:MP��'��H]��񉁶ēB>F�{/ڒ\}�Hb0ڋ7�t�ΓR�dEXŷi
2�'���G�$��ʟ��I�Mre;��0  5� �/ZXFq0�Z�IĒ,	!�������|ZK~Γ�����O�FDjc��>Z������K����	>����B)�4"}���?��&Eπ��RfR�c5�Xb��H�,�i閧
���'�4���)u��:�*L�@�骚'���!ړA9�S�A@�Z��1(�#�.�
Ex2�z�f�lZj�O
����AӮY��ݹ�&�.��#���?CL�F�Bp����?���?�ն���Oh�(LHRX0�c,r�4�b�O�ԛ���Z����`�',O ���	�$R�r(\�V���G�Oఘ�/Z�z�h}�'�>,O�����ڈ����C� \���O��p�'�D6��U������Gy��-v0d��|Hčb�b[!�yr)�3Z�<,z�-�1v]�07�jh|#=�O��I	`nqڴ0�BvbQ��v��b�k�>Xx���?A���?q�����?�������=H��"�X9��l�.>8��*�r�6���	9wP���d�O�H�c!Ά]�L� ���;��aQ�'��l���?	�,ūDlm�ͭ*  ��
��?������O0��'1H��ku)��7��Xc�*>HWb\��^�@֥K� 7T��@U�	R�����	~y��1<F��П���W�d�Q�%:R��U�=R"�hB�Ѕ?V�)[b�'�"�'0����:O��O哵"B��Z�,Y�7�.E�n�T��<٧삮b-s��V�@k"T*0���~셈GA7D�Q�xK$��O�$�O���|���A���3b�v�������?	���9O��;���$?�����#Iߪd!D�'��O�����3[�d�5��}2BX���	Wx�x����1T.�5 GҀ'E.��� %D�d���o10�zBQ)T��x2�=D�,��݌E�p �d,Z �	&F!D� �v)�'f��z�J��2��`%D�����n��0:���*x�)A	"D��k7��m�Dٴ�D�c}(a�?D�|���կ<��u����4W��b:D��yw�57�
��`�k����c9D�*֪Z�{�%��H�Θ�0"�<D�軄��5'xe�p�I�W�p�*��:D�8�A`I&
�L����9*P�h=D�pq�`��#����%E�E�4���.<D��0��������3Lu��;D�h3�)�_��cv`�TU�;�a5D���ti��1�ܷ��(�4$9D�	��ѕHێ�J�\�hZ$�9D����ǽ�j(S3��F�r���(2D��[#�[�PfDP1�+�j3w�"D���N�L|X�׆��W�drdN4D����cL���l΄dw\=P�1D��b��_�w��[�7��y�`�$D����B=t��Y�CJe���j��=D��8�c�C̀��`B[�L1p=`c	 D�t0�[w�0��F.��'�>5��(<D��ȗ界b��T]HE�d�9D��`�Z|�b:�  3���W�6D� ��*\%��xQӣ���"�/D���Gd�a9��"T�ܫ"'�k�I0D��8���va $�!�ƁCL|�I��+D��1�K��P�.Q+|�QV7D�0�@/+] ��EA�fThDB4D�t*&�	�/��U�C�_�Lw0�1��2D��85J˾`�Q��[�O���@$D���Ǎ��+��@���m��¦ D�\Qw��k��E(�*�1W��("&<O����̊4F\�x���>� ���G�8F(��{A�Ą8�S"O�A��D����}C�T����Ց���(�a)��SãSH�Q?e�bb'r�u�D-@�d�vU�#k!D�ʃ.ӢG%� ;�F�
M��mҁ|h2,xP��C��b��'U��%87��ļ�W+���P
�K��q���'V<�S#��2g��+2�˱-R�����$l2Jt&������,�Ju(w�ܟb��&M+�In�Y�6G��ZDl�z���|��Ě�yZ��`�kő-u���'��9F�h�8@�D�����%؄�3���V����@D!��X�_ ,Y�K(�<9Ȓ�'`-ڐ�'��xp-�
HJ�#��%ck�}��'��<� ���!3��uEFx����&v�蔹�]q�<�l�U��JP��%�|"���
I)S�#��D5l�?�'e|`3�����|� c �M�;�\�s��fy�� V��Q�v)�i�'�UơU0��y4�C�9{��1����y���	5��,|�J�B')��<���0���A�T4���y�E���#�>C�:�
��h�'��R���6�0�1����`��x��[����JŠ܎�0�Jf�
���i%�P��	̟����S�6�B�՞SE0���h�$�!q�t�²i��+�l0��肁m�K�8�d� -D�; �*���{
�k1�X8Xb`� ��1��nZ���B&��d��)���	�X��4�J�ls�'��`%t,� *l:�\9�%���y
RJ�����
,��}y'%��Ms&#�=5�,`�D� j�h� �!'���2�4	�`���e���>��~����go���b��V�a�`�'��`��F�!`���/��x��	�D������V S�8Y��+I�/H̒�ݗ�� #��u�'>��6����|�)K(p¸Y�f�$vnUkW�%?9�Պa��!6~@���W�r- �I͟pd�4-6�UjU�5��Ԥ�A���b��]�֎��'Vm�v������9K�"����aHx��Q$!�	~�\ �,_;"a��Ѣ�O!x���l��k��h�(�-4�( �G0��'?�i�O��1��ߏ_��Հ��[�<�Aq�<����&L-���	cY �s��, М�O���2�!Ϝ�U���p�*i0���?�5��&�<\a��6�Og��<HK��C2��9#�e�NB�A�x��4�X~?5%0��-�@C.��D��$X���,h���N��eS��)%��+G������(ѨOt	[2m���.�v��K|�PQF�KV�����7�6����@��D��P`�o'XX��l�*%k#F��"cp|:�ƒ�-�\]�O���D���U=�%V�U:8I�ј�(x b[�`+tq�ԫ��6�UQ0���(��H6B�~B�L^"阇���8�x�H�z��5�c,��Y�܋����q$q�R?�A��F<�<��O��ʷ��X��2D
9s��Rb��<+����	��q�3� �/-��S�D����=R!�2o:wP�	A
�0��'�h3v�p��pd0���I-4R %�Y*��JT(��+D#� TaA�`8����RU�R����8,�ꨣ�ƙ4n8|+V���t	a�\1��C�L(�A��'N��ũ�)סO� ]2��7@��I�J�].�>�r���psV)F�n��a ���iE�D�5.����+�!�����5�/�1ю�Q�OM��1��֎I�"�ŗ�Y�y#��^��)��*I��|��'�`��KP>�"�[w3�,�B�Wx5���>�ȝ7됡[1�B�6���be`T-aO��{�	�U.ekG
�F���dE%G��#�U+	2=���9�0���P&Z� �(Ó\N0x���: ����
K_.TuĈ\�|��	L'[�N���鉇k��z�D#��#)��v�,{�i�j�)���3��'���X�dZ�忣'%I3�ԙ�N�-R�lp��酭����q�~����ԟH���郇W6&IK��W�^^��Q�W3#c�P����-#L#<Ѥm��^=�!ç
�&�����a~��
$V*�`@*v�RQ��#�?��P䦅��V�?�T]�@�ZC�)AfJH�ɔ<�@�h��];b{��!N�3J2�L˗D�v;ܴ!���[b=� �>O8MyR̈����vNʏ���p�ôgU����ݍ,g���5��IX��3�N;{���/�)����oEj�O���g5�Ӻϻ0�� C4)̖ê��dm�5���+; ����@87��"Uc�"��*�HL����R�&#=�;�D�Q
�z^��g���!��ܙ|��I�OZ����t� #N�Gf[�sy����H����'�B!v��7m�x�D��'wo,L��O �k��C2�<�ygi��	!��>�e�ݪ������gh,�ץ�-6ܬ���K?k�Ru���<���̈L���N?�K4�A�Dd�dH�ꏘq�t`��f�c�K@Y�D+���4�j�3��Ȭ �`d�0&�/J�<�e0O��HdWD?q�Q��>�a��C�n	��.�$[�PP0�5l)&1�R�'�$�����)g�`I5�ٵB7�CS�B���rť��Y��r�fZ�g%�	�6jv���'OJU
�镒.��S����MI�Og.IQ'�	��hl��n��|�O���b��"��� ��ij�8cQ���ЛK��|n)j]J0@%��y� �����M���� C��� (����0�	*��i8�		h.�93� B�C֭�@���,m|��b��'�0�8�iͺI��ɈR�+l&�s��O֭�'��H=3� ��M�ș�R�<d�QX֋As���Ѐ�)k��y�wy:h�aaJ6nU��ɓ@��k�r� ���_��$]��M��V�x���,�Ӻ�A\�
R~Pɂ��
{x4p��->i��@�d6OT�����<7|�	�N#��d��	]��l3�,(C.\]���=���D�Ob�p`��7�?٧]�Ql1�$*G&L}��M�� p&�X�Lʄ����ŢxŮ,(U������A��}Ъ�"�T6-��r� N��~Zw��!�p�Ѕ q$���y>,!�	�H\
�O����iI�g�I�1���A�A���x�烸J2�ZC
0��ɡq�>���(RI?��y��ü�w�[?�V�Ul+#\��n4w��qDd�E&�0�m�	OiF`B��4�4�F��f�3�I2|�xm0uCR	�t�	���DB"Iid��uh-~;�%�#��&��)DK�`\�RE�		����g���B峀6���U�fJ�$f�X`a�P�;���%Q�x��?>��i��C~2D>��$���9F'|<� ����^y�7�M;y�bP�ǐ2*Q�|c����*���%Ԣ���h�o}&�k#��?��?%E Բ%3�	�CZeC"���"[��B,Y6�)}R-UV�$�B,)��� Z�`�r%�
�06B�%4]�� 5o�h�B���� #�dX@�M_,s�b>�)�fN
/R[x�	�d��f�5`~]3#��m4��36�9m)��(t7��=ͻ�x��k�X�4�UjW40�H����8=�Љ�E��%vD�S�Y�L=��+@(VҰI�'�	��QNaX��"�P�R">1��!p
�H�&�1B�^�!B�0��ٺ�A�G	��uI��4才�T�s���d`��G�7tF���@I�9���%?�s�A4�$�#���Hݫ�(!D��9�j˾��X��C�(�e�#'��it$�U���xԎC�Q��'K"�t�u������
qb�H�'J2����(Z7[ma~���vVA"c
�I(j`r�T�b��@�!0�a����XDk �+0y\�S�I�'6�*�������p�T�8)~#>I���E��$�q���h�/ԍ@�|P�Z�f�:� 2pXb��Q���h
�����$��T�ds,�[�(����"U ��3PGFgAR��a��ٟ(P�G�t53�$�N8����$'���T��!<9<�Ӕ��2�HO�����U�ʪ̃Q� ���'Y�����@�d�K���"�Zu�A(�/Xqu
�߸ ����EG����5�^���>a��֚
�$q��O� f����k�Ʀ�XW)�nU�H��ȃ3���	�U�����8=`�X���d�yir��$'����w֮A��|2A��bϜl0� *�K�*hR���3%���p"�A�BL��'�l�+,�S�|	 j�2�4�������"t)6x`�I��YO��8����B���<Y�h�q�h�����_�t�vAv��7P����h;�tZf�U��*�s� �>m����I�%V\d)���3@ɓv�,��O�t��E����8V��'6����ԥ4��L�&��Nr�H~�UN��!)�0���/�(!��ed	Y�˘Y�Z�#��|�ho��?�'��1��Ϳu�.�k��T8�*�o�b�<����ą9�֕(�O����t�ك��A7jk�����%̘�c%N/��p���XȨhF�"}����D}? 
s��,%*�����6Q���I�+�d(S������!���_� ��i>m��a��Z�%�ּ8t�ӦΗoN}J�iUS8��KVX؞��e�}`�H���J��m�� \ *�b���	ܣT��0�'�Mԧ�Ob�����|�E��'s�́"*�,JΑC�̛}�'=���l^�y�D$y�M�2��x��'��M���%g�q�bKC�dTyb�'50-�'I�-��E�)����n�lhJ�g}�V4H"�]_
���I��yb�P�db���h���z�9����6��K�C�{B��rCDT����	�T :5y�/�(n�D5C�A�k���d�5�f�(D�ϔ8v(i`��� YQ�`6}��NMy2#UB��eµ�?�zm����4�]�`uJ(ON���	�/ד(#����Ú0~�×��B���b�|���$����f�>Q��>7#_r`>Ib��Eg���Hˌ"�@��	�NW@)8W�̟ �f�jp$�:'��\�T�৮J%D���p�cV�32^�'2�'xrhP���j�'H�1K �-m�&\��S��*M�L�tV	r����Q&�`����"�I�#��QЄAI�g�dI��
�e�"�O�� ��5K�y�`��L�0t��(k�]Pg������V�V,����V1+e�q��?��gy��"Ad��S<_� 8$@Wf�< �~ʒdۓ���\14t�!F� �l�$Y�}����KS'\��	��fħyF�(<)���k��H����4�xN�|�����Hf6�mQ��#�4���ɈO���Ė�m����N�(�!ŕ�
]n��"AĊE�����6O�U�v��5I�VE*6,��F7�n�50���<����$�^�@�:�X��A>g<j�zq�'���L��}Fv�	��>>�1�O��0�M8}�|}g���\s����I+'�K����f�P�5&ƕ������PxR	3��$�4�� ��<˔JF1��2�@_��bޓ)d�O�`�L��]�9~�PJ�������A�?�C�I�D�~H;@�6��#Cg*]N<�P����C�D�':��'X����)(�O�2�;cH�O�`(9�k	���H�`>Ā��؎�$�*q�4�6 I�9�d8(#���LWu�@b=}RN�A�9��'gܤ�(Yǐ����Քj�Z��'��1Y� 
�\�V(�[%x�'�hh&�(� �EC��Qvޡ��'఑yu�ӻr�@���aY�P�8��
��� hm�ъ�_��:�X�+�@ ��"O:�Ѫ�#y�l�Pkҿ7|��Y�"O�b�0�p��C	
xRN r "O&!���9r���pf��C�$"O��4"�/���A����(��ܨ�"O�a��_�T`V}`��~�ָQ�"OB�y��, \���m/2�K�"OP]�ԉ�!�`�P]%I�X\27"O~���[�B�̈́z�	e�V-!���Z�LQ�P�
t���y���%!��WZ1�B�@�T6`}3�M�,�!�F�(�T% � P��r���!��"a�lYQ��<3��z%m ]�!�V�@��p���� ��V `�!�E�����+ >�HڢOJ�R!�I�Z �������\�=��߆x�!�d�!X��c��.���խ�9h�!��AM�$yq W�b��L6�!�$Ռp��2��5��!�wK5�!�J�LQ��"0�^��c�I6k�!�D�y6y�f /"���CQ���!�D�ZbXD tc�=�4B��.t�!�Y
}���r�J&{ʎ�1��<1S!�0^����L�.��\��"��7P!��UNu�������#�"X�
H!�w�2 k�"Y�\��<���ƥa��DH�6����/��g���y"���o�\�0��>4��:�<�y�DQ�~���E 1<�(�A��y�畔Qd�뗆O/wb 
�Ҟ�yc:A_��X��J4&�E� !C��y�n�8J_Xuc�!���hЍG��yK?_載Xv�Ω$��Xxfg$�ybf��1���1Rl��dXU�S��y�g��Uh�5�4����z`	���yB��V����+�.��=��@��yB�P3S� K�m_nf�`�E摿�y���)3�b�z�':ˬ���Bٜ�y!��C%$=�kQ>���a2�[*�y�Q���䠑��8����cM8�y" ����Å� 1���-��y�C�%��1�`L	5����cL$�y���7Xƴ��� �,xff؋�yR�R�02F�����wH>��1�y�@�0h>����M�v�ґp���y2S4a%��%�)8��SUC��y�-�.O�X�%��,o��tγ�yR����<�;���&]��"7����y��T�K@���re�n=�h�����yR*�*�<�ٱ͇�m�p�f�đ�y��ϭLM�q#�Cm� ���/9�y2�Ҩ�n!x��.QjuP��[��yB���!"߻;H�[GGV3�y"! �E��m0H�1�H);g"���y��:V��'�0�!a�ɗ��y"4rM�w�ړ}I.�穕�y�X�k��*wb��#� [���yb��'�
08U&�"n`��!�yE�u��@Y�j؇-�d�;�oҨ�yK޺6k�1��-/�\1q�`��y�i��o%�48��+&K-"��'�y�[pQ����LH[�K:�y�AʢO��5s�b7<��xQ
���y��J"Z�x9��!.��0��ƾ�y
� 
���z`d:q.0B��0"Or�A�&ťMl�cB���$9d}��"O�Ձ�ȁ�!��a餀HG�.6"O����@ʨ�� j��y��*�"O�`�t��.��������t�q�"O��JE��j�=ªY�'] ɢ3"O�@�!�g�t�r�
�j|�@�"O�`J҈�{FМaP��?k�4�"O�a1Ҫ�k`rXq�)D�?K��Rg"O��"���7Z�꩙��	|5|��"O�����I�NXؑ�fH#M��+�"O��d���B$�9�ͮ~�r��""O�����S2l�A�@�O��Hi�"O4��Բ�X|s3OA8	���Bd�I�<Q� �+s��j�%��#��9I��UG�<�F��Z�(+F#�+Dx*qAJGH<acA��2	y������k�Ɛ�(!��2iƄ�d��Y�B0��U�"!�dұsC�ܫBf�j�Z!��(E!�#I�ddb0Ϛ�}bm����`,!�Ȉ�$��Q��3^R�,�P(ѯB%!��X�0�t����-$����	�U!��H�{��
���$`9��Gs !��7r��(�F�D�>���(ʴ!�d�[��� �:*F�(��D��{!��_�s'��Bk�ACHp���*�!� (=p�P�L�M/�С"Y�{x!��A7p��tT)�,)f! �|q!�d�M�V !Ӌ�0l���`!��RX!����>��0EW�	j��2©�<Q!�D�%@�0űA!�V���	�	�,�!�W�d~f,R�L֟-w�)Fִ=!�����@\j^v9+��/z8!�J0P��x�6E7�p$`���!�D��~�ҩU��6B�=aC�	��*�S�Ot�Pc�i��Ӧ�衤
�����' J�Y�Z TԒ�i�<T�����'#�ps��(&��␎�$5��r�'sў"~"7䏿R��� =#�.(�'QF�<9 I�����bO:r��@!�	Nz�<�E^�$d*��'�8pb�ط�^<���R��<�Ԥ�.�FE��d�
x��<q�-\O��Bb�]3Tn<����&.-�s"O�ZD�_��>ũ&$^Y�P�s"O�`�儼zW
 0�āh d"���I�O���K� )u2�!1�]�rj���'Ȫ�NF����p�GlT����'Jr��W牖!;���W�S�1I
�'e�X�R�V ~�bɇ�߼o���}��'��kF�_8Vݦ����';V���'r6�2��5�d��	܆A1��'��ݱ�@ȸlF �b�Xo8�ݲ�Oڢ=E��gN�L���ʕ 
�(pz%91�(�y¬[�}br�D2�t[�oͽ�yG��%@�YB�W	���ˍ�y�N�J�T��!�ƔA,p�$�ؚ�y��SZ�ty��%�0R�4��0�y�cZ'()�F�Z��Pi҃��yB�M��,�W�ɺVtDEP�̆(�yr≍B��3�h�yjш�X	�y� �<�r9���	:��`@啡�yB�Q&.�n!�5���H`��y�e��G Z�ڐD�"���7h�4�M����s�\Q���B���W���r̘"O� Zd3�]�S�8���: �F�q�"OR��L�*J�����΃,�h�"OZՊ��*sˌ|P�螪*D��O^�B�'�=Dl�AMO��2���9D��ș5l�J٫F�=x���E8D�ԑ��Z�9)�i��`��r�Hm��G4D�d��N�/(t�
6P���2s`3D��d(��*��E
g���;�`��9�!�dTRu��3$�X�g�~4	� ��QH!�D'A���A���0֨P����|!��\�$����ײ0�r "��ͅ)!�dD�mr��P�<{��my@`_${��6O��۠���U	Lh6�F1�ر�"O�HTe�F�0�݋��Y)��'2�DС+��QAf�a��Vxt}����v�E�0��a[K��F�^-�)p;�O�O�%$�98��y��C liR��2"Oxp	D˝%�fD�Ǉ�X$I�"O>�)�n�u�ě%L�c���"On��s`�*y���K���q�"Ov%h� G������] �"OE3�lŘVf�@��L�,��"OXI����1U$�,��
����"Op��s�޻DWZ���(Crh؝	e"O�$A�!ڔ&��M�#(�:{���'"O囃�>���Ц6����"O�)Y0/A�P-2L�l݈j�x��f"O���@�`�¹�7��36��`T"O�(����#tlJ��D�grꄡA"OL̰��J�u]��p!DMx���r"O* 1	B*?�0��I#g X�"O��	Q�^�R]�-�����r�"O܈�%c��S$��iD_<���H�"O�u���Z�t@�E��`�9�"O���K�� ����㌫-%�UA�"Oj��� M����W�R�N	ƙ��"OV���/[V��$fT����A"On�s�dеz
�o�S�L�
A��"O�0�v\D�3#�R��H���B�O5��"R.�)h�@P0�%JG>|���'�8���OۥI�T0¨T�)�(��'�rT����5�D���H9)���Y�'��Ճ���b��Y�I8.�J�'�P��#	 �Ի�K�O_zX������G�\A���6�0#a���B�!��+A��a�H�?E�N��Ao�,�!�$Y�xj�,��O��a�#p�!���)(ݪaꟴe�XUi�k��=�!��ه^��9"C�0+z�d�����!��G�|Qg�I��l�uK�}�!��B�=���q��4����d
�*�!�3SE(X���\2f��]�i�!�&I��]����x��b��-V�!�Ău��4�֏Γ ��@�^�F*!��=ּ��֙E�y��k�!��PeTX
f��a 8��!���sJ!�H�}�̉!�j�����Z&#�36!��A�z1{�E$+*2m����_7!��{�&=B�U$2�u���V�!��QƁ�w�J��"�Q�{�!�D���D��dLy�x�RU#A�#�!�d�6"�h �A�u�@p��/�me!�D՗VV�@K4K�?�������0l0!�$ق]���{򂀈EYh�"��B�0�!�� ���Çэh[����K}pT�2"O��0��Fi \h� ^�T\��"O��Hڴ��!	�(��G"O@�#��׸���aƁ΂: �QX4"O� ��*Cb�Hh3�J/e�h�G"O*Iq�D� ��b�kda��"OhS�(�'~�J�i!M�N\Y�6"O2U�ƊR	v���b�2�"O�8Xp���>�(�0�b��;���s`"O��Y���;MX�!*�`G�]��5�"Ox�0�NV8/e�T��n�� ���"O̸(wA�9�D��6�<W��lJ�"O�(&#�:�̚��­c�P��y�W2���K��^)!�fAM�y�EĶU�ܡ�%��>&P��r�N\?�yB쌥5�x 굢R1�"�0�
��yR@!	���Pe�����K�yRc�0�aRs�W��B��j�&�y�ƀH���A�.�V�����C��y'u)���P�G��r	� �L�y���5��}!��.�d��h��yr�؝G� pA%�df� S����yB��,L6X��l�O����#�y2��L^�����F�W���y2�T�f�Z
��@�� ����yr��!����H�, 2�{#�Ԗ�y�CC�S>�Z��!3�aK25���'�z%R�%�<[lU��J�2�*�y�'��U`�<��f����@�
�'�>|9@+�So�1�d(�)
e��'���`秙u�����ߓ�&���'��)���:���zt�2̌,��'����Gݭ~;�)S!���֜H�'�p��e�H�&9Z��`�$K>mj�'�d�H��ن"�5���}F|�q�'���	r��0�����Y6x��d��'���8S	�m  ���̀�:#���'찑M�)h�h���H�I-�,H	�'�Ԩ$��D<FP���
�w���:�'}"�x��Ҳr�E�F�U�m|��'�!�G@_0J���G��m���'xf��%i�~�bA����s�Bx�'�H���@ (fSE|�z��'��@p �>71�p#d�V�`bu�'����F�J�F�#����_܊���'�H��%F�8,�\�B�n�� 8䴪�'j�u����xo�Q:r�δ/V��2	�'�l��!�2���(��2=���'����Ƃ@�U�d�N���'o�D�U�/HS���6!A%v,Y�'ܜu�N =����D�D���:D���#O�&.��@u+�P�7D���u�сqiz%h¨��0ּ5crn3D�󗈔	Q"d9s�Tȼik�-%D��:�.� :H����Z�zĹ�P#D��po	6]�΄`�E(~R�)�!D����j�\h�b�;Th8�@ D�г�����
���g 7L�:�3D����'�&�ѡ�
A
�e�%D���Ge�/�>dsf�H�_�� /D���o36@@��F�q���Ҍ.D�H�!$�-X�xpZD��Z/`k��,D���<�x��m�'#�ăf�+D�l�Շ�g�R�{� m�ّ�'D�� ���񅟑abjM� �+�l�Qg"O�Ya&��z�p�
qF#]}Č+�"O�l1��?2�}k3�ta<Ъe"OX}�v!�2Mi��T�oHR=HC"OT�Hă��W��q�RfɪZ� ́ "O���"��zA鑯ǆ2�J}
�"Oj��4�¥H�<��ڶ<Qx�6"O�@����#ZpV́�&Ѭ?�Dz5"O�P�Avl�8JхŌ(%�8��"O��#���9��R҃v���""O��a��N�o�( Ѷ"ԪL�d�y�"O���"��߸�RQ��X;�AZC"OH�c"�AZR ���pʐ"O�@�F�����@�4&Ҝ< u"O�a�w�51и�T�U�G��U"O�ݫ��G ���(0�D�b�6���"OPx+��3X�D��҅� Hlp�as"OԬ���ߩ��I���v�t8�"O8�@��L��Ik�*C)���T"O�DpwN׵#t\B�	M��iE"Ox���@a�
ѹ�G�%rtT�y "O&��R�Z[E�H�s�]i`���"O��1oc�.�bD�>%I ��"OV�%솼T^�
�c	�a����"OHD3�=5��hā�+i�򨀂"O(�J�`�$]��,�᠌jN(�"OT�*�j�	YrDl#� ܎UA� 
�"O`Q�u#��Z@c�oT�w���2"O:0��J�M�d���8j�ɨC"O�(�!}Y�1GjìU�e�g"O\�q�	�v "��a)T<U>�ْ"O�ɹU,��4M�D�چI7�-B�"O ���*R	mۢ��c�){�]�C"O I ��G�	lHD	�"�:r�@0"O��!��^����� K���u"O���Qh%6Υ�� �䦉�"O�J쀿_��y���]69�"Op��G�n�0#�"����"O�I�b��aT�b�^�xt2�#�"O�G+@UU��p��ɼDs��Kt"O���*��+ ��c�
"U��S�"OE���X�7Oq���0M<�k"O��G�G*Pm2@��)X�0Q��A"O��!Υ<$�}[��­^���X�"O���E�͕��9A",G�<�H2"O�a2��TXؑ #D�}L}�"O�M�ƋP�Y"u�#a��W ��X�"O��	�H��K�擇'����a"O�hs'�ÿ1Y�ȁ�� �$�$l��"O�ݸv��
gr╱v/Ɇ���9A"O>M�䭀? 7�	*Ĥ�J���"O�LH�LQ1�aZ�D����k�"Ot K4fԫ+�VȘ
��! �"O��u���L�1�&{�(�z'"O*�q! !Tw�mi�+�dL���Q"O~���G��h�@�T*wE����"O�LbPc��J�Z�g���Y:U"O(�
���7A�?8\p!#"O&̚#��u,Ȕi�.��W���!"O��(Vn�=}�z���L���U"O�c� ���q�"S�""��P"OE��(����cU>c�qJe"O�5�s�լ�XS����wqV��"OF50PԨWh��0� �\�.e��"O� �Ԋ�	�5YhHA7��^�8Q)0"O�Xxbǽw�iق���u�]�""O�56
�$\B6���wBRp�A"O��H��	ۨ4��M�8[F���"OlHR�Ԑz���cӞY��X��"O��rAg�@���c"�&�9�"O��C�J#��p�fW?Q�Z���"O�P�4�Ų;�$���G���M�"OD�3�PL.�K�-�'Ԃec�"O�h���AE(Q��īV��p""OnM��T�J�N�@���P�@���"O��0&�\K̦P�ak�z!��Ӌ}��2��DSǸ�:��\h!�	3l�D���Ū8�X-bIE+�!��U�E�J�qg�	%�N��/�!�d]8]�<�ċ;q����0��>u�!�䑠k0�׋+g*�����ua!�ړJ�B���
D�C�0e�Wf^�o�!�DLv���K�ʗ	y�������tG!�$	�
QD�ӧ-	9l��x��ňt�!�D�Lg�K׬%h���L��Ds!�\=e� 0���=+2��bfI�'j��b�Cdޕ
���Z#���'�J4AC�<K�q�P"J�!�'����d�2u$pX�K>?H4�j�'Ӹ�I�'�� �P�P0�@�'V���>�a`�R|�L�A�'�bٙ��G?�01 C��T��
�'����&�ƞB�����>�Ty�
�'X8H��e]�F�=�6��*5&��
�'�l�µI�J������Ď2�RYP	�'���iЉPH>�����u���	�'^D䫗-Tu�dz���u�)�	�'��}�&N��3��0�u���s9bTQ	�')8%���J�R=�$��3�,\+	�'b 9���qp\���נ&�����'��@���Inl�󏉯*��EP�'�>�@D/�#ɶE�܍%4y��'�*�	P%#���u��,$4�i��'ZB�8Ҫ��Z�$e3$$ƫ)Xİ���UV�{�zL�hį�%C̪ j!�$w��	�R�O(�����҅Y!�̔*� �;�@]0ZO6�×�T�no!�$�!:
��26,u#�A�EV!�$
��*ɑ'��32�!�fֻ/.!򤋪`֍� G׊R �=�veE
`!�d�2>��1�f�>jo�%Q E�#.�!�Dռ'�v�AueYXv�3��:�!�D$N�����;>#�L#�ĉ��!�d�8~6���!A�t�"U��)�!�I�9��,J���\�2|����w!�dI&
�B�Y$�U�D>FI+!Fק!�!�<W}�p��Z44%�DH�k
�*c!�߂Y���u�8�QajِH!�D�,|��C�TP���)\6XG!�$ٰP����[���d �A�48!�dPB��q�)�N��q��EE�DT!�����6�YֶEp2kG�?�!�d�=��&.�W�0�ɴ�9!�$y� ����3�t�!�.OB!��X,�Qi޷��LI��ݕD�!�D�C:\��Ň�b�J8�B)�
�!��[�X��R�	)Z�j*S��
!��՟T�a��8�ƔI�@7�!�� ҽ����8��yh �	�O�p8W"O|�'[�UpVX����B�����"O(Izu�ҀTI���q $o��-8�"O���*C�'s�%��T�y���"Ox��F�:Aq\��F��
\��:�"O:�" /Z<�TEa�N@#[F�aC�"O�#��R�#{���Ǡ:	�;`"Opl�2���u�,y�#�)��dZ�"Ot���ɮ@P�� ��^0�v��D"O��A��֕FYN�{&�&;f,��"O0 ����� B�@[�
t���"O���r�L &�>�0��Wl	W"O�=x�'������ Ŗ>N�x�q"O
�5���q��|H�
82�9�"OF�{��h60��Cݛv�e;�"O� 1��"n���3��21��xs�"O��2sBZ+|��x�7��r���8F"O2�8�nϻ5Y�D+%�KWS�e�%"O���b�{��/Q 
2d��"OP�H�CM3�Ȁ��oy{�]#2"O��7@�(q�ޠ��+��y�h���"O~�S3!�Rx}S	�$�TLؗ"OP�̶ jιsq���"�N�sp"O Y �I�`4T%+A�[e2B4"O��S�!�,V���K�A�*fS4� �"O:��E��;J���\�$@A"OfP�o>��$ĥI����"O���d.	wOn�p �.��0"ObA�$�Si<�u"MD�lȎ�x�"O����,ٝC����wkR�@�=Q�"O�58��|I�!�	4rC��1�"O*�zH�-\Z�`��G��o?����"O�i����O�:� p��&yH|�"O�Y"�N�"i�@���1��p�"O"�
� ϑ<^�� S/��p""Oj��#��&4�0y�R��1q��ҡ"O �9����A	�l��s����"O�9��ʨ6��<�f��"#z�"OZ�)��uv���h� 0	>(�W"O|!�l�KL��th��|�j�r�"OXY˧AV� �����0Ϥ`;�"O@q�ƪռmt����;~Ä���"Ot��WE�tYr��X���r"O����,�lzU�T��iH�"O"8!`��Q�1���_�ا"O�y3d�n�Vtٳ.ӸSF�0;"OHa�DꌿL�BDpG�ÚUdе3�"O�M�ğ_F298�ɬ��|K"O6� 	�j��D!S�� F��ȕ"O-�1�Ĥx�����Ά5��!"OZU�P�M���1���`q8��"OX�ס�����(f�l�s"O�� �=�Z�	QFU� ]�= �"Ot��t�UY���[Uo��t���z*O�p�!iLq7jx�f��l9z�'F��+��М�HQoW���@	�'�0�BeS�J`�؉@s
$A�'3F�SFF�>��O[�Z���	�'?x�9��
4X*L�4����Q	�'��bg��,�Ȁģ4+F��'�r��h��y�q(Z�#.���E�<�#]�YT�α~��Z姊I�<�R�M8�De:���-7�6���L�<���P �Z��@I�J6�r��LI�<� D�Z�gF�W�"xb����gj�,I�"O��Z��ݹ��hqKY��<���"O>��B��
�(�ɦ���N��@"ORLsCCܺ}���*=�����"O�7�S�a����=s��"Ox�vY��a@��H>cr d�"O<�b��F;i�=���I����E"O(��T�	~,�Y|<�]��"O���1-/�6�!'��?,��{5"On�)�mè+��h�dh�$= l(sV"O:��.W�TАY�T�X�/���"�"O �	r�o�z(����s����"O4�;f�:5�1��'~��"O����g��A8W�]$k_��`"ON��g��̀b͸M��Hk�"O4aDʂ8F7"����	W��8""O�t�6O��,-ٳJN�����R"OVu5I��Ӷi*A�~���"OD�"��
4]\��qkW�bBL� r"O�uk�|�l��Ӏ� O[N9�q"O��2VnK*) �*��f>�1["O U�ƅ"&���Oٷ!'Z�BQ"O��Jchźo�ڌ(Q�W6 !hX"�"O4�r�Ɛ�F���bT���2��!"O� �A<=����G�3�(-��"O�Ţ��<k�e:�ǝ�S�|���"O��򍛻�+���{q���6f�Q�<��j��)��U��$.g�J��N�<�P�C�.~E�e�
���b�N�A�<A��ZQ#�&�/�-BR��H�<��d�5El=��àg�����|�<��f$B��j��x5���WIy�<IV��&X�KGɍ
/=�a�a�s�<�� �)j4���gK�2���H�W�<���¼hG�A�^�Y���2�(D�����_�9(�5
�� �����/,D��R���JH�!�A��J-|�{wo(D�l[�j�$4�B�CJ[:r�R��U*Ohah���3T�Փ��S>R��w"O<MH�PM!�-+0l0Ӥ��"Oh̛VÅ)D��kҐ"�l�Ä"O��k��� 1�B$R�L�W@9h2"Oڽ��kڛs,N�i �@��%�"O�ՙf�+Ɔ��CI��w� mir"O�9��o��l�4�����|Cb�#F"O�� �'È�zM��>)D%�"OΤ����E���XF/�=c,N!��"O<p�s̔	�,4���L+&�q:�"O�E#T`E��D駃��T�ra�""O��h����B&���$#	�t}�8�F"O`!��Δ�H3���gb�=:0�`"O�x��E�m�� ��#��Q�"O�|X	�RՆ�{�N���8�y�H�K�\�c�ɞ!����%�y2!'PN�Ih�U��l�!cA&�y��-W[�L��͠����Cv4C�	�0�~�hE�K�:�"�P��B�	sR�I&I�P�h���B�	�h�ryi��	=��0�QKA��C�	>��PAs.�!a��|�PkR�H�pC䉠+�R1����:pThqvfO�,�C�I�'(N=���2x1zw�K��C�ɳn�f��T�d��K��SR|q�w"O�{��!�7	�*
;����"O� �jQ�E�P�H�HЧD.S%^��"O@%�eMCWĸ�$i�/D�#"OX<5J8oFt����_�Z; ��"O��R��EKN���C�?ޠru"OD�pA���f����C�L�^ib"OF�D��G��z)���$�b"O���W�TRT�j2�N�1:ZT$"O�,�5���9|��ps�$Z�
�"O�T2$�[4@�:y�(Q���"O.����3p��P7G�\P�"Op��W� (m'd���~��%`�"Op��F�x9֍h�N�Y��Rr"O~��qF���/

����"O����g�KB�r�օ^�8��3"Oh�v��(mu�9�����EB�"OzE���n������CM�0�*O8ݹ�;S��2anĕG-�]��'#��rd��9��R��1�'2t�[���"nj��G�*>��ț�'�<T�TGI>ό��c���0�l�H�'�)*��pJ�@F��.���C�'����Ύ��)C�]*vd�q�'@�p1�3�5���8#�l���'�b����r���B�.L��S�'w�i�3�U�0���Z���hL��c�'�R��� lDn]�ACPҶuz�'cd����9Hk"h٠*�;w�|ah
�'�5@�CL8�����rF@�
	�'�� ��W=���O�V�ġ��'%�U(��$�S�#��F�h���'���!��)w�4ͻD��:C0ɘ�'PU�Wg_�Y�&����CH���'X�`@%A�==��S��&�p��'�t�cԆG:6�8���C�
��!�' ���K̸hX��RE�#X�v��'����� �@���Ҳ�(��'��&ʷ�f PA�U'����'����@.ɸ.=>�Y!$F�U��'C�0Pkδ^�ⱂ�܈n���@�'��� ����9HKS��R�2<h�'+@1�t��h�4��%�L`2�p
�'d�!�f�L�B!�1!!in�
��	�'l\\�!�˨<~��j�E0g��$�	�'Ev�#�c�=_��D@�����N8D�xӑ�Ы�R���l]-�^9aǆ3D��:U�-�2�15I p7���1D��k�H�(W2�ШS��J��A�+0D�<��G�t�93�jӘf���H3�ON���<����re��8����k	��<�V�����);H�D���
%�ȓ/����m߈b}���*��/��ȓkp�)R)ϸ[�N����:_����g�6	[ �-h�lk�&�4f�l��+�� ���$CW֑��O�::D�ȓV�б!r�B=>�`UҳM@�S�z%��}v����N9l©	���U�I����Yk���0��2+�2E����H
E	i*��	����	q�Ѕ�ȓCk�щ�g����S�N 6$��Htp��K�P�Τ���Gv^�ȓ7<u�4�d;��3���f��ȅȓ� �զ7gvHH��@�g��m�ȓ. YBJ oרh9��gU��ȓr�Be�e��"��ĠsO�Yü���S�?  ,�'�2� U��D��z��}��"O�L8��f��Y�� ��B�S�"O ���vrd Fe�2;�h��"O�P�4��m��HG�/sm�<
�"Oh�Jҧ�!����)����Xg"O�u����$쉐��>+G����"Oh���+� �ɰ�˺:ĕ�S"OZQ
�['"�ƹC7w���@"OU{��D5s�3�FN!BdbIJ�"OD��o�F{�p8���%���{�"OH=Xc��d�ؘ1T��)K��u�f"OT�F�6*�%�!;S�hLRQ"O�� ��_����U`��(��=�"OT]k� 	�dϤDIt��M���å"O �0��?"�������)7bI7"O"0w-
�V:D��"��4�bt"O֌�� �j(�Ikv+,P�c2"O�9	5'�=w*���)�n���p"O��	tnЃU4�������c6|�u"O����'�1sl��UR8��"OH�Dc�4��5�4�J) J`�""O��
v�B*��uҴl��=O(��"O:M�-1:�t=[�˙h�H�t"O��P�٢8�ie�)Z�p��b"O��j0σ���B�Ƀ�Y��@�g"O �1�
��d�ӈD<o��%!�"O��Iw	V��@]��|�J��G�IG�O�@���MQ�y���zK�/�(Hq�'���*CȘ,U�p@�C #��d��'����%�D�o_�`3&ñw��P
�'񂈫E�'�J�L|^�T 
�'�n�
�A)>*艣
�~ʭH�'��5 ��@�Q�ܼB��V��'�N��E%�@^\�u"��)�<��'&B$�Vg]�9l1�d�"i�y��'��� ��*a�ABt� M���'�(LɢA�׌�g�Ի����'*`9S�͟7r�h�	��U��'[���E�\�tL����,�"yj�J�'�h� b�����
��`�X���'�>�I1[�jA/Q�q�TE����"O~ y��<��!� D��S�,@��"O�A�Vk�X0q�Q�ny��"ObxE�&i'޸��ʂ7_4E�#"Oh	�P�"P7p`*���CL����"O-+�`@)�DT��(�2/�"O�e�9y�R}�0GG_Pvm�!V�0&�ȗ'��k�@�0��+��s�K8D�l����a `#s�� �JZ�G"D�$�!M��4 �̑rLA<xk>�@�n5D�@�]\A��7�fq��{��5D����T�Z��U�A�F7o��y�6 )D����@JT�>8rd�C	cʸ|
�&D��Hwe։�����A�1$`(aW�/���OF��>��N�@����@+ �V��P..�d1�Sܧ<�ŏS+��d�r��l���ȓ
�����Y+Y��,����>�����A��2�Y�h����g�K� ���|%��Nٕ ���M�TO���y�Ҵ"4�2����FN�%[s`ȅƓh��ۃo� �:2h��@��H#���<ړ�y"�.���v'�!x(�2�f���y�K:W�
��]�W����L��yB /P���+�Ώ:YbT8�瘟�y
� �������1,�!�А��9�"O|��׆�2��}�dT�3�6�˃"OZ�P%�
=iɰ����:t�j��5"O8\�'V�G�XxC��!�(�cQQ�4�IW�����U�Ü�"h0QkA)�2���i&�$!ړ��dS�G�!H�Μ�Ĉ�E��q=!��@=~�L�����Ox�х�01�'ha|���k�"P�Ʃ٬,���!@)�&�yU�9_��H�.�v�*���y��(@Q{ �׼�X|�]��y""q�P�2k��f�$�֥���yB��dC ����`�ĕ��J#�hOh�����xu
�HGNƪ=�>,A�hV�W"!�4��� �,��
����!��I��8�F���O
8�H�C!�$ݢU����ᏮAV����'Ɓ�!�� ~��c`��-���Ԇ��!�D�4<��v��e��T"�/� e�!򄀥U���s�G�@X�@� ��'���'���6�U�CA78���4E[=kx*T�ȓUr��8�D�:
�J& �H�,D��E�`��#h̀4�0n֠A�����A#J�,���'��_N�!��M���չ Jei�%�j��Ƥ�RdA�ƖUs �[�}�����0�tm�@ňtdq#�͊%ݖ�'<ў�|BV�F([Sļ�f�-u0= ��[{�<�G��HIR���P� 5��k���n�<����n �X�t��-"i�0�i�<!�\J��"ǖ���t0�Ge�<1�BK*0^��`�\��ݒ3l�b�<AdÑ3��-�0�����
xy�Z��'��F��/G�s2�� ȥ �v��Dl���䓐?�M>���͔/7F	{2K��`�r|r�f�!�D�`�PХ�#�H��M �2�!�� %�1�a�:
�vh���2N'!�D͈a��1���#� vʗ�!���:cd� 8 I�C�V��+ �Py�J2{��)`P��XZp�i�=�yr͕%���8��B����MX��y"��,B��9��Z�������y�L�apP,1#N3�&�#�L� �yb�Z d�&�IQN�&E(�{��Í�y��ߙ�0�˔�K�%^x�kE	�yR�Q5>͜U�P��Q���dnH��yreK�B��a
�MG8�J�qQ��7�y�j5L���e��2� e�'ұ�y"���*Ȭi;�쁗"Bl�3f�N4�y�M��
�p��"�3�B�	��D�y��V��X)J�`T�`
�HR5�۫�y�b�Ne0u�P��Hy��(��y� ^0	$� Ƃ�BV�+���*�y�[2�z$kAhP,~b�`�C��yb�Ĕ@|E�c�Y5& eC͍-�y�g��d��� !����(@��y�猼F��<���#�BH���X��y�oԯ� ��(U�ܮ���c��y�@ڬxx����Ix�>)2F���y",ƺYkfMB#�I6*�����W!�y�Q-G.���c�hH��B��y�
<d3rQ��aƑ~?H����yi����9����y��-)%����y�f�+5�0��C(��z��+�y2�S3f�^ճ4 I5 ɶ�r��<�y
�  7�*��$��*J 1@"O�(%�ӳd��+qBZ$/	��*�"O��Sħ
/�����[�X���۠"O�KU�$)4�C�F!�r�q"O.I��ط/V}����G��y���y��8`&\�B.l1�'�y2� ,>�VhY4�$�����y"ŏ�)z�D�5kv���V�J+�y��EP����g�Thq�H��yb���;\�ʲ��	��X��y� ����.�x�(�7����'f8�Sb��z�R�dC)�|1��'=��J�8�L�+D�0|��'D�(̴D7�@`��([V<(�'(�y*u`�4֤lk���E����'wh��"˺vLdze��0��#�'3❃f�8wT%	 ��9�Q	�'��U��NW����*~��j	�'���4mX�.B��u"�
&���p�'��������%#�	M4��'���BD(��;�zPkTA���l��'��PG�]=-	��ؐ��(=��'F��h%6DȘЀ�Q,y�n!:�'2͡�&߳qh�	Y�nw��x��'�i�喯f�J�h�X�n�B���'��ᷩ)t��(�K�c�9s�'.�����$!x�p��6Wmڨ��'m�r.�>:^�!�s�TJ�d�r�'�z����F sz��aQ0L, �'�����.@H��D&�"\�r�'��	�j��Lz���c�ͽQϠ�J�'�֔2V�Lk�v��g&K����'��r��\�`�씫THÊ+��Q�'��M��kGcK2m�CAz�a�'����'ʝ�H:��& W#_�h��'���P�ļ6�^�iE'�[�����'�"�*f�B����Ͻ���	�'_�Y��R�} ���f��O�a�	�'�̥*�f��^�Ș0ᐨ@����'"�a`�,{��� `E�-N^�)�
�'�T8g�V:S9$�S�@կEUX\�	�'~&0���V-#u)sM��'���
�'s�P�D��.��1�g�)Y�Q�'�xU�0�i��{�GW�� ��	�'���P �
-j�c�):�pQC�'����G/��ꬊ�I��hx�'���s�l�9i�`[����}��tJ�'�0z$�|X�� $>|&�d��'�n�;"���|_p�p�C�oeX��'��{��ɩ,�^��Wfǉ[�l��
�'*,8"��X�84
�
���$���8
�'��DP�ɑ)<բ݉3ΫM��E
�'
��ʐS 20���S�G�t�	�'G
 ��fC�"�K2�D:����	�'�(H����ݫ���:g��y�.�x X� �,#��xS���yb��S0ڹ�bN���>}z2�M��y+�7[�����N��a ��y�!��B7�փ	>����ƒ�y�)�&,�J����!y�J��g�1�yB�цg~������tn�a�7��y�41ER�h�Y``�І@���y2�R	:&�A�sI
e��	V��y2�Բ0��mӱL�Ej�����ߗ�y
� �� ��L�g�.|�`����HHa"O�Q	Q�J;�,ST/΍Bf)#�"O��;c,�v���Z�t/~�1"O�q0U)��)7��K笏}#x�6"O��0ChN=M2�uz�"
9*�"O�Qq2��b�� -��(��QS�"OxUs��ԑ��µ�!�Eф"O`L�$aN'��$��j,LF�<�B"O��3!Dҭ�1�	��B���W"O�,�%Aэ4B(+Q�{ѴeXU"O�p���Ӈf$<�qE�P�7_��""OR(z3+֩D,4E�������y���bE�f��3�����Z�y�EHz��(S��(2z��bF�y�͚2c�����Aq2�DX�g־�y��=F���]$n�ڈ�"b�;�y��6r��;e�
i����ņ�y��ӭW$���K�aՎ�"����yc8��@�5fO�R��4����>a�Oe�g�� qLƭ�5̛�#��Q[!"O��s��vŁ5K]��v�X�"O��Q!�G�P���ߌ+���Q�"O"�P���)q�^ YU���f)s"O,q�ү�W�t�c�Q�a
PT!f"O.i���+���;VO�!,\��!"OxE#"�Z6Kh^|{�Q"YVX��'|���<'���gk�&�fa�d�i!�dQ�4��+��g�0<#�-��Y]!�dʡm!6���ʘ�Ҫ����\!�$�8X��iU���}r�+�Pv!��3F�r�T��:-�~�+Uj��J_!���-?[� *D��=ʦTz�HʢG\!�[(2�>�T�� �0���gO:Y�yr_���'�T�`g��"oP��D�)c��q�	�'� �9��$o��8�K?���	�'�����Q5d(Lm[�㈟P>4u{	�'��`p4g�n8�9��<;%,A;
�'��9�GLC.hx��#��tg9D���e���k<�P *4N�x��$D��5N�J�R�2���&�6u��/.<Ot�D4�I*74>�xc� 2�^���
�V�B�ɕX�2�Rab�d�h໴"M�b�B��8|U�A�@��k*�$����`C��p8UU�٭Y	�A�%�9`�C�I�'b	
Uϙ� �O�lZ^C�I�o� ؀#�D�����L8s[C䉆A���AgɟT5� Ap!���T�F{J?}����`�0H1p�N���.D�ܘS��"el�8!RF�����
(D��E�$i�p`����N�lA�l;D��0�9T�M�Q���	Tn8�@�:D���K �i�:D���?<�&����9D��� �l \Mi���7.�Xi�V�;D�����]���N.(�.�xA$:D�X[ĈS�T��(��(�O�Ꙓc$D�y��O%
O�SV�D��aK�m"D��ٲ�L�<abǬ��u� ��5D� ���),�رʴ�+%��$*��0D��z��ʿr�]��	�6��ѐ�0D���w�1�*�b��]�UZӍ(D�pKA��t��s���b�~��J+D��	Q�Q�7���2��7~YxUD(D��St �!pj�36�^�E�'D��!����:0\j�����t�h�O3D�� ��)�ؖ\m����?D����"O��٣I܏�Wl�_�4�"O�L�Q&H�o�5����$��- �"O>�0A��o�$�q�2"��u��"O ��u�_&�Pqb�GPAP���"O~� �b!�F�C���[�"O��# �L�D~*G�֭k�h8�R"O�ѪcT�[D��{����&NhPx�"O�m����
��E����v� �S"O\��GE�v�!�φw4\��"O^l)t�^ Z`,
��_S�T#�"O�4 D/��&���2� Q:Ұ�"O����'B-9�`��`�ORƸ�d"O �"�/�� ��b�שX��� "O�@q�I>2�8e��	�\av0I`"O^9R�E

p�#�^�ݘ�"Ot(SpŅW��Uc��U*0�� "Ojy���4�A�b��< �9"O���M(h�(IH��Y
H ��ҳ"O	)�їj�0d �X�*�s�"Ofi�-�6$fĥ���C���"O�|��P+3�z��c���N��8�"OX\򦇉�&��k�.ALl�"O�� J�5:�PRB)�O$����"O�� =*;�Y+�
D� B�S`"O<�pK�"���gN***�ݐ"O�ha�!�'5��3���uyh�y�"On4j$�X}MVx�R�؉7b�T33"O���A�;r����فUY��Jg"O0)�'JR�m�8A�Wdlwd`�$"O(�T'�4�x����(RX���R"O2="'oW*Z�FU0����@<K�"O�8�����*�+�%6���C"O\ n��/4�92���?N�E��"O����'ZX���e�|%q�"O��J6F����qç���y��"O��2m
�&%��r�%��@�q+U"O����cPN�!pWjۉe��x��"O"ݪ��zۆ�S�E1?���	"O���'H X_�9�æ˺e�s'"O� ������0��"Z�!F"O���u�K�L�f(	�B�4;8c"O�8�qA�-y��}h �Ã_�B"Od��'���1���e���g�j�C"OLab�k�O�:pj5l΋$�R4�"OX�PR�
 � Υ/���"O���S��T��U��:�V=�"O�-��ު1p�!�7��N���"�"OfM��Ƈ�j��ɒ�m������"O���H�
��� CRu�r@QF"O~l���%WI�a�� �(8r@�j"O�ѳ���$\<�%0 /��ae�"OV���Ò�qJ���+R���S"O4`��"J�2���p��0�G"O�誷��;}q�D�5KL{	f�V"O�<�௅K;(\���~����"O&q8�J�H�p���P�c�R���"OT�cCJ�z�(��xzh�;2"Oʘ���X�l"��T�M$z<��"OMq�Ӷt�����OZjgV�"�"O"-��
��y��"��uyJf"O�ܠ��VX��4 L9Nr$��"O6� "D��8~$-ە@L�: zA�d"ON!��Nj ��X(?��#"O� �h�t�D�
B���s��)��y9�"O���pmߚA��H��(�|k��A`"O�|�b/mqĄa���P-
��w"O�)���Ǆ���jG�_�s"�؀b"O@�Q�o+$�j	�%ə�w�i�"O^!�@ �j�$:T�G�z`~h�e"O�UXPI�'Z~�yv@�b<���"O<���+�]�p�&�ɧA^Yp�"O�H)ed�"��x��CD??�ل"O��#�2ZJ���-4���'"O"Y�GÙ�lH�S��6}��"O$x��=[�}˳�X.3g8�a"O�l��C��g2<�� (S\���"O�lc�O�/V�PL�殒]RR��d"O��24�>�4�yum�TA�e�q"O��:��؆x�Ta!�Z�`0aa1"OlT"v�����@�f؅^7)X"O�ܢ��@�lR`�e��3F*�t��"O�`��(g��d�SFR�zyF���"Or]b�Ĕ zyH���ER�) ���"OR��A�>L�<a'$ל��mr"O��A�Mo��qд�@�|���sV"O�+#b�5>��P
�d�
��P�7"Ov����y3v qe�m}�""O�Cu��N�,*A�F*��P�"Ojhb���J��2�	"]�����"O2��D��~�f�(��T�s�B8"O�a01g�}}U���,R��mX"Ob�3u��"��%��a�~�H�"OD̝�k���� /+����"O(@�&N���H@�O5{����"O8��sM�2�lN��;���s"O��q�(�'��A�MQ�g{�I��"OlawhN�s������YAr75D��{��O��x�P'ï0&f�!#�1D��P@)Y��&���݄q�j�r�&.D�Xx�H�~�l�'�*sr� ��1D����PW�t(A�)C*V�rn.D�2�͔Z<��{�&V�om$EX`�+D�D㤁@�0� 9�������*D�����]~�a��̓��0�[w�'D���B�1�u#�a3^��x��#$D�T ��]awR91 g��Oh� *O���E@�t]���@oQ�!���ɐ"O%��Kع��-'[��� "OrQ
�l
�<m��ĉ ��	1"O��6��+R#n�{���z�"�a�"O�@�L�u���(Q�ɘ]���"O(1sT! ��@� ���Ըw"O�iC��T;�3Qƈ9&y4Ģ�"Of�h�dҩ&�$�e�[aJ(a�"O��R�#ãB���)*j2�� "OR��U��E@`�PN���1W"O�@;�X4E�F��,��|����Q"O
�z���7�tąH6��ݚ�"O��qF���\o�1�$D$M�<i9�"O�͑W�˘p������B�'"O@Ԙŕ�N�HzR�Y*O�4`�"O��A�cFY�,q��w|�F"O.@��
�w�`l@'Dg��	�"O<� b�\=t��ms�I�'vN4b�"O���e%Yi��hA63s6�3Q"O����Ԓ@m��bEN�V�m�S"O ���-O�xB"�	�D>"��d˒"O� ������iPDV�55�3"O�q��+�5|�P��B��R�W"O��� I�"r��5�N�BP��!C"O�0��g�b��zƯR�8f��"O�E�@H�(]�٩�,�i&p]��"O,%;��ٰY�v<[U+q��`�v"O��"%T�jC�@��T�B	ê;%!�D��Ot�!�P!�:Y�&LX���'3>!�WCY����D�9+��"�>3!�H$���0�A� ���0� ϑ9&!�d�f�q Z%o�يA�O�4!��0")�2�ν9�(��#�s�!�dЇo��X��Mњ8�r��v��~�!���bp8(s�"1�>M��*a�!����9f�Ö,�|}!���!��&9�x�����`�U�*+@!���4���⅍�)&L�v��/!��/j�lxx��݅qN�i�e�8!�d
�Yw�Dcb˒�.i��i g�Ud!�ɗdY
��ߡkeZ1����+rZ!�1xD����<|@�"�<T!�>��4Zu��63Į���٬ A!�'x�&q�G�	o,4؁!�
�R�!�U�+�D<�s�\}&��$�A*�!��h�0q��XN%Х(5CJ#G�!�d^�>�R��!g��MR����!��VHe��a^6�,�3�7[�!�Ď�)M&�ڑz���I�"��{!�D<
��ycOX
9�F��g�{!��бo����ƀ��`�3ÂӟD!�d��H
�}a���g����a��?�!��74x������3�	�woE�3�!�X�H�ꨛ�"B,oz��U�Z�2@!���S�P!��$�/3���CV	�jE!��_�Vp�1��vjY��G.5!��h���fnEaB�iCf�XL!�Ě���X2ϝQqv�
����~�!�dC��@3�2h��R�R�@F!���>�����9�ĘsC݀!�D@�,�z5�F�8P�=�p	�^!���s�����>L>�U;s�M`�!�D��R�2���5<7P�� �X9�!�X`�Q{!�$}�l�T�� !�d�9h���N>uz�L���ڛH�!�U��ta,ӂ�
$b���V!�?�N|��25������ՒBY!�dG*F��+��ǯ|?.�	R-W)@!�d
1W��!0�G���t�1�vY!�$J�?=�(���Q�v����n!�ER,�����|H��ڒtg!��^8W�ݩ%-�5b�р0L;]�!� *_��@ǲQ��XǀH!�dӓW� ��O	^�|i�e�7�!�S�
�TZ0��p_r02�O1#�!��͠�$���&K�$Y���c[?by!�DW��D�p���5ڪ�󑌛�e!��K���O?+���k��3N!��3K �d�%X�щ%lY�NZ!�dV2i�p��s�	�lK�xh���\`!�F�Ԩ[qʈ�+��P׈� 7_!�	�0�<�i&�W�z�V�Ȥh��_!�DU�d�+��2�>��*W�JB!���(zLPp��R�F1󆯒c�!�$�%x�
�! E�j�L�ʧ�>B�!�� �,��ݬk�\Ç�6ID�8�"O��h�O�~�%c�E�� c�|��"O��y �?s�&�X��=;t��"OQx�ߙ �ȵ!��ؚ2/"�!q"O�����k����N��U��"O^���M��Pٔ ���>~�fX13"OJ�H��Y1�B`jAi��+)N�X�"O��f�>����e�S$�ј�"O]	�S�w�2�B�g,Km��"O@t�V�G�4�t-h1��1rTNI��"O�5IW�a�Vu��1|��R"O*|;�/��/˒	�e��9�!��"O��Z1�l��{������"OVP[P(��RXQ`1+o�����"O�)I7�!���)��1~.��&"Ob�Ԏ]�7T&�1E��57g� ��"O��҆E�I�qcv(W��.;�"O��i%���T]�Ӧ��"��ts"O	�Ui�b3�4�'��<���"O�0�vG�v�A0�h�Z�P])�"O�@R���ЀhB�Zö$YD"O`�"B�F�li�5)�d�]���"O��9�)��bWd��@ռ/�t�#"Ofp�R�U�|�v���H-b��-K�'��'�剦G�� ��%P��v�(yTB�ɨ��Ͱ$`U�^��q�P�,B�I./��M+��sϲt��u�B�	
�6�{a���������B�	,_�l(�ĝ�+
�;P-M�+�B�	�q�VQ��N�2ij�(���1ۮB�	Q]~ɊR���Zà����J#T~B䉥L+dxҕ@���91��3m�B䉹 �Y ⊔���)�S�ɨ���\aG�)�iW3�Ĵ�@�^l��W$�!�D+u�D���շp�H���!�Dў\]�t�G=U����;N�1O���dQ4f����HL�5�� bA %�ك1�����g̓4���9��E?� �w"��(W�؄�mEH����&+�ā*��ʄ.p���{&��͚4�,Պ�P�&ܾy�ȓ>�����(�DH�kѦ2n �ȓR{Xx��|?d���"��<�l�=QK>���*>��tj!O��{&,:q��%!��^&K��@2�b�+_��R��(�'ha|V/�0P�TI�*	$���T��y��5���0W9[�qѧ-����D.�(O>u"+PJ�q��!��yS�a*D���w�r�ԽA�D5i����!;D���dG�2�hk!�h�i��F8�O0�	r��+b U�1���p���|-0B�I�`�+�O�X8�9�a�/'�nx@5���G{��)2B���J�
�/g�v�K'
�3�ay�(\@��h?p�C�.K�i��!��\Lv��I^�wUp�£)�w5,y�Ea_��	&�X�:�Hc��>I�JP�t�x-��N�D�8<ré.D�k�b�ٳ�����c�5ac���d*}�HB06̐8�=.�m�ClO��(O ���Ɔuxɺ"Jæ,^�,[��ׅ7�!�䓈Z�(b6��LI��)S����!��K�a_�;���C8��Calт
2��E�$�;�0��	N
�I�����y�	ե��Q�2"�/��Ip���� ˄�<��y2c�1J ��R�!Ș,��������>�O�4@M"n�- b�]��A�%�c��B�)� ����X�[!n�#d�q�	�5�'��OH��N�7k'*��@�_�&�x����y"�U�W��Y �j��Q�`��bJ�&��Ӑ��'�Z�)�ӶB����Tc�F�����*pW ��2ړ �.��A���Nո]Z�bQ�@���'��}nB�S&��y� ,�y�2o�_'�h2\�y�JA�1w��k����|%s�@�e¡�[+?����
\,Rja񄒫aġ�ğ*nD�@�A��~k�]�A��y"��[ȼ����l�\��va�8�(Of��dVTY��Ņ!)|࠳O�D!�My�R�Y���3m��0�Y!D�!�dӘ c@�S�[�(�$}	��� m����F{��������(q����ІF+�t1�%C�Ty��'׈�2pf��>N� �!*ϊ,�x��'L����G�l*��kȩ tf�3�'�DaJg���0!����"#�qДxR�7�� �3T�i�䢈�KO�lQ2����|�	���D��TmҼ�Ƣ�� �&)�Qa[4�!���T�YA����Z<Q4Aj�ay��ɾ=�&5�o]-2df����)�DC�wL�(�r�?Y�f����l�*ɉ'�*���aT%Rj
d��n~`-Jd�0�O��D�>�� �(޼a�˥r�<��D#�W�<��� ~Fl ���=�z��AS��?�
�'t$�R7DĘ8����$"�@�ȓ�|!⯘�n#"A�W{;O��0�y���'I0��1L�@
7��J\4�3&�'��r,ٳ%�X�W+\�i�L����A��yb(�$c�`�0@�v1�)k�#ٻ��>��ά<�q��S�Nj��D�9��=q��<�O�|F{J|�PҺv���sa��\Z��a�p�<іe�UF���N ;��q�r�\r�<)��h�UkNDr��拙d��,�'�tP�1A߳-��탴�"^?�ai�'����D}-��p����T�\1ܴ��X�d(�3�\([�*��N��j�`X"%����ȓU����wJ��2��G��o�����djܸ���
Y�J��W(��S~�ȓ_uP��Յ�.�߲^F��ȓ��}k�D4R8hTK�"Ֆ7& ���n����#%�ͩ�#��U=P���+��
�d��K�����8^[��ȓoP�Z�E��
���e��.��Ɏ]P�g\?�dh2Մ2�LK��J���	e���O���[$�W)`��h0%��Ya�8H�'�.�c���p��񷭒1L����'�u�B. �\%Y�@"s����'1��c0��Ng1`��Хk��t �'�l{��4o:��P�ϸ9��RH<��|8���!\=	@T�� ��m�l�ȓZ�(���K��=�Jp�q	J�P�H�IM<�$�ѵM#ܫF���@��6IWl�'S�?����zT�1IL�J��mZ�J2D����囅
VFq1��D���!q�<i���6i��(K7fԍ|���F��,>�B�I�o7<����.O<���	�N��B�>e�Z��\5)�L�����*V&���ċ�?�ѣ_�`��d�d�	0fJ�
BLIѦ��fV葐a�Ϋ����
�q���b��%�<�A�HG�$L!��"5<���"ظN�(}��H1HH!���X�F�@Ϝ.=���
��ӗE���r�H�C/�:p$�;��E�eHY��xX�����j�� �4{����׆�O�=E��� �H���D�ˊt[R�Ǜ.���u"O�:f-^"n�p��~� �մi�ў"~nZ���؃�P�#肰k�'{�fB� "g����K^5_U�2j��j��B�Ɇ�*�J��.<�y�p咽UH���2� mۤ�!��H������\ծB䉆 �0����؉*� H���P^�B�I�t��)�w�A�~�^��a�/c|B�I�lӔ����G�y�$�S�FFJ���7�	84�����bΖy�����m�B䉭m�X<e,�3
�A��D�M���'Jў�?�;S-�&x~��J#�X�5~`i���?O��IB�J��}�jB"j>�J�	�%ZO2 �ȓ6V���;2�:4�%	͝omN��?Y���~:��E�r� �{F`��	 ��y�`�m�<��Ӿ*b1��Y�(RT?�HO��}�8����	�%)$�I��I����ȓL�ݚw�	C��Pr�îI$�q�ȓDf�x0�l�(jP�R)Ln��ȓ,��\R��%a�>�I	��Նȓ�N�	���]A*�K��ehņȓ?���@R+S���'*�"�2���7�
��a�J}Dx�㜅duTi��Y���P�Eз;�aC$�PS�`Ԇ��$Ē���:���ׄ�`���?�bM"�m��*�v����>ͅȓ"�&����	G�@ J@�c�0��;P��D_�# ��0S㚟U�N9�ȓ��!Ɓ�;;�R�2�[���ȓd8\��"���.�b�2���%�ȓmð�#�D�G� �I��鞹��zξ�ځ�߳P�f���Ɛ3n���gpr��� �2-D���_0.�h�ȓ�`a7KK(���d2ʲH��rZ���.7'�U��'W�:�Ԅ�5����]>{�ܹ"�$� \�4��ȓp��lr!fQ�Nm�Egw�`��ȓ�d� B�Z �$Q�Q�%�, �ȓ[St
�(�* Jw�m��-��]��=����!��ԙ�Aږ~(�9��:^Ɯ��U�Mt-� �%sн�ȓqJ�(�d�
83Fr'Fٳ�A�ȓi�2أg8��R��/\�:t�ȓ6(�S��3�b�`n��
��ȓ1�)C�ŧS��!s�MG�,p���dL{S)�0�a��4�&��ȓ~�0A�-Spu25�Ţ�.n����yc4 �)Ű 伀@��� C��Ą�MΡ"!�^.Q/��s(��-���ȓx7����S��e"L
_h�ȓnw�x`0��+L�v�8�a�y!hф�	�Jp��jə(�8��YT��,�ȓP�hPy��F6�]P�O�������0����]j�f�kq��nl�ȓ'a$�էkG�EA0#ٚ��ه�51L(8T�!ƴ�G1��,����9��`̴J��Q�C+V>��̓�p��A3:&������G|��01�J`�P���`g$�k����y"mݮU^Y����6Ad��ǅ(�y�a�b�k���%��)���H��y/�3�*I��"i��,���y������H�CK8`$5x�����y�D�r��T�İa��IS��
�y��ˬLJ@���X:e��!pL�;�y
� �����^6�8��J�"AR��Q"O��x	 �衂�`?HCFE�t"O$����86��!�0\=&�x0"O<ȥ$�&<�DX�'�TAaqV"O@$��o�g}�@p��	�.6<�"OFE;�/���
�0���Y��Q��"Op�;�!V�8ИZ5�΋#�61"O�QeGֳ]���D|�n�""OY(�dӾ}-�p��\�wX��r�"OI�mI�Z�������Ip�("Oz\(���/�T�Z NP<��"OV�p����i`��D�8����$"Od�#�k\W NQp +�ip��c"O�Ա�	�@���!�A1i�H���'� r+�Ǧ3���<ɂ�P�_2x�T�\2��
be@x�<ـ�K�9 �.�?nӦ(RJty�@:Q��A��(��)�0lↁ�v�O����D�j`n1��"K��58�'M�5��h���3
�>�Nt�ߖ�Sp|��hY?"�����O���'��'K�P�3i�R�4���؃>�
��d�<�"�O3	�~y�g�\�&=���J6T� (��W�|���P��^1A���"8�&)���9c�0���Y3pQ� ��R#0�s&�xI�CG@��9�vݙ�LTuPS���jE�m*�"OnyYf�ʗV�DD�!�;*��>O�tIժD�(�A��8L�zQ�a��T�F�?�ke����y��Å[��e㐎;D�<[��I)h��y��Ls��Ғ��0P҈T�"��K䝉�G٩(È�?��3K>ym�!G��0X�:c"m�$�zc�ҍ��L	�N�#3ቨr��ș�J�8��%�7*F;^���r�-�,������f"=	��/\AX��f�H�g�Jq$@%m�<h���"=�w��R�@� ӵd �W�G~CH1#���3EΗ7h�5�P�Ģ,U�GyB�A9"����`��6iq�P��L nlZ���-�$��d>O�ʶ�T#+$��z��9J�dB4䍡lo^�?�Ȃ:�ṕB���]x��] �*�K���+�6L�w���"~��!h��U$}��FI�jm�Y���"x�La�aZ�Ed�\�V j�7�U�|�!YT&Hog���[���Uo����@�� b���I.{o�t�GM�R T �4��
a����e,�\���w!�:;`�e�b$�+r*�%	�~0�����/C�*�'Y�
���aS8>i�}�b��vt6ט�F_e��$B]6[���x`RAy�eQ=N �$��Ʌ�\pv�@-4�Є��#x0u�P�V�(V����,��?�� !,ӗsfͻ2���Z��<��/��"Y��W>.X���?���C�C��|���ZDBl 6�O+C�*(v�p?)20kxN)B��A�F��M3�(]�##4����v�<{�x���a�ǝ�fLR5CA++ψ<�F�]�ap��ǧR<��LH�h�څ�!�G�u'	U���0;ҠZ1�~�'X#9�a�CNfPk��N�Lt���e�ТE>��t�x�kE"C;�l���L�cE�����4�p����;g�j��M^�A.�)��@����[���M��{D�^3\� x���D� -7��h��F5_zh@P�:7�d�`$��`L�e Ƅ ���C�`OC �`�Xxt@@h�:6�L�����jd��� ޤy��Y!�Ҕ�^`A�sN�!�"<1��7(^)ăܚ�Jq�1J��K���
S�lt��-�-S��@ӄ�м��|���r%j�4F��K�aP�2�'��T���Mt��*��N��hK�q��O�PW�b�>-����>��D�95��,K7i@<@n5�5*V`ϊh�v#���`�e Ǹ^�d�!FI�n3�y#���!��*[x�1���l����� �x�DW3T�b��בݴYrA��/��2W�r�5O�QR��+�zU`�吩@Wl=�-��Q���ϖ6]���$��?8���3SWD!�p�M˶���{H.!�J��!ޡ�	P�'��0�s��D���c���Z��p����MsF�X�w�,9:�+Lw-30'%b���Q�̓�W�d�٤��w:]��*s��qHr��!&1vs�GFb�
����OV]��DȰ@Kl�2��F	��6Mӝfj&��C�Uu����%3=>�!fS~9�8yU��U��s��cc�����$՝e)�7��5��O�M �������-3���'$����]^n��C=(��qAb�i�/�	�����E��S�%T7"CKC�iRZ�mڐ�Mc���)mE�����W|��Z"�	p�����$I`��Aq�4:�Щʥ��"3�А'/��t���M(X�9�(�p�*Lrw+38�މ�%�Р0�܌J��C&q��	�M�(
� `���?hp�P:FO$u`b�:@`�.��v�M�f��m
�F(�h����8`QAc�9X��aT ��FW�1���5iؓ�M3� �g˜̂�֠r�:k(� yf�I��5�-�>RP����A��h!�)��⒞'ӈ�{�eZ`c�`�Ʀ]��Pw ʉNr�X;B�u����I?K�������"%�h���	=����t�^�>�)b�)�k4��ӱ�H=N���QC�!$�d��v3��Err!UX���Ɓ��էO�W~R�������^�)�6��J�l��>P]�IjBA�8mf	*�(�U�T��^:I�Q�C�עf��8X�
�l��y�[�,�9��2AR�ҷ��B�,�AZ�M�I.���J���R�5
�6�p"�@�J=&t�t+�< 6�M�p�Ϻ[��S�� ͚���v� 4�pc	&����L�Fo�E���n��!��/̂@h�F�S�tX�ƌ;~�Ȓ��O���lA'����H�6+��+�S�Gl`!bnX=?�`8��>�.�&�����3/��+1�S2Ei@�13��L� ��L�`�c��S*S��uY��ʰ�T�2.@:��%�K�^����,;�P@��V)1�
f�E�i�j�IrG�r�~�2q��+c�R���nF�!}Dp�LV�;�RƮDj�f�	�7�� �d����gP"AA����'��,��>���ǺbG�����԰��Td7���HE��U�P��ǈ�P������L�Rk0�H�ō�?���.����操P�@��q�	�T������l�B �v��C�qB���l�`����n���Q��۶�V�m��d�ߩA�er��Z�i�x��V��k���0𢅙;O��MR�#�ڍQ��]+R���Č�o�0�s2��!���p�b%�T�[s�J(�LQ0� ٗS>)z���7"�@�)�c�e�A%#tZ��SS"-�Rm@&@XV2	2w�	;2(�T�VJ1+�D�A���ecZ�rv�Gk�H�B�t�`P�e�#Z�����ŬZ�@�X�b8UnZ,�u _9I~��'�G,��{�FE [�Ӕ@�/��"I�ScL���8It���'��D*��c %#��M���5V\���2�IGy"��A�Tm����5%DA�ȶyPBi(T�u>Ic�!��0eJApǃN$F���Iާa"��F�Tq2�p�A�\��Ij^J�Ts�J�|,��P��H�*!{Qd	u?I�i߱l�Y�UFv8����p��Ӧ ��7�T�Qt�C;j��aI�	��o �ӏTCz��{�\%�!�P
\��a�CF��0�
Փ�g1���E�4=i.�R����zB�<���T���� uh'�Vq��X#&�X�&EI�U�4�X��ia�2�)��h^�)ƐC��L�l��O��p�R(BQ����lV�{V��e�Z�K�4E ��K8�Q�����V9@��ł[�H�2U��J:����T �}��y�/�VyF��AY,Lsa'��P��Iŧ����ڴ!��{��A�/
PtX���X�H�|u���$� ���!a�¥�O���P��"@=۶.�R������	�
Lb���0i��a0e�,3N6,���7��4�d@����C+}��qC�ȑOH0�L��5C, ��2�� ��I$[�)zW"Æ��FB�a�t�U!�#up�p��Ywo <+�f�$Y�	:�A�
$ʔ�`ϟ"��&�m�4)vJ�0)I��릅�o�Th��	 e��<�2��m_.�EzR)�6l"��q��GVf����T�}�"��c��*�Ra��W�(bJ�7�B�9$
�*�zYSj�>�u�'��P$ �J�N�aT�xa�Q�$�@�swI�>'U�lDzR�1)qJ���ҐU�୓TH�,y(X��jV�D�ႂ:f�SF�'�d����ڭ/��S�1ev]����;M��2h��j�1���&�v٘e��.��i�O�����$�>� G�mp̸�-Q%�d�
�J�	��G _��(2���u�B�����*���Rv�R�[��P���ũ-|���k_)e2��J�7tT��b'�
)����S?_��	�@<�����&X�1`�T�PX�ćO�JI1���L}hP@C4�4�T�%P�)
p+U �@l��^�L%��C�>:�z`��NR$j�,����U�04���5i�6e�V�K�'-n!K�I&"X�D�`Ӱ�@��/s��1���6\L�!F-�u�f�R�@H�#*d�-��i���\ '{�����C*Nو�BW�.WQ��8D` �^.>�F|���I7ʖ�-TH<j��[�B=��[X������3	XU��y����5K�N"&e ��$(��X��i*Q)B��>m��=BЪݐ��̖X�|	�kV�8�n%ٰ���8r`V�!{��
"!·�,���˝�%b7=XL8L��[}\Ź������4Sw*8F���g@��]Y�6-\f�Lu;G�Y���3�˜8αA�w��8 r<���]:�L�K�LE��S�G���đ�a�U9c��T9d
9#u,��`��;�B�#V퍕B��+RGM�f����c���țk<Qa����Z1�DR����+�B�G"�Û	����bZN�$� �_�G�$yـ.,�U���g���R��ۅL���9NP*�C�‰<���0""��n�4��5K� �����a��Փ�
�R�l�6]Q��LØNa��{P�=?��E��%�$|�8���F�?����'Qi�7�BJi��S �ڼ=��]�qeP�?�DQ��L�A}t9%ˈ�?mh��<)kH�;g~��3��r�@Yt'FU���C�W=�H�bh�k�� ,ю!�,���lȑ+�^P���"��X�m�Xǒ0�R�o�$ʈ"��0��A�e�üb�(��?$z��Xc)޶Y"�{F��{}��ǝ�3��I�E��=a���GP="z��(�N�*B�x��">C:Jx�&Ɲ*�j�bD�V�}.��#�'����ģ����i��,[Cb�b�۝J>X���I�p����d��!����4cĝ���)W��/]Ht�q�
�zNpYg��I9f��[�q��I�EDB�Y j@}Q�	`ae�:�L�*_�1,,$��.b�
5�+}#J��T �<��� ����VȚ������I:�KIގq���!�:/�,7�2,�H�[��QE�g�н��HB���I��@�"v�I!�
\�i�&��H�+
�:��AZ�[j����+��PL�?J���5�H��J���+�0����D��@��h���Ґ%��8�؅���!��ϔ�4!���	p�u �i�C��`�YwAx� V�]d`JfGQ v���eo�)��tH�	+�vH+���Q��4���� ��3�K�o�2�	?W-�iK�I3!�� ���"�b�c��Y��� CR�Nn�-J1I�T*��rS��idfƶr�����|<J��$�7�ȃ�jG�/F*�H�f��'�,�Q@N� � ���	Ba�h©���$� �!�x�:�Df�4$� �qp��!��'��B�իa;��r ⁪w������$�v	U,L)R�fpCE@�Q�!!ւT���C�J�#� �f����Tyaf�.;6�� B�	�j��͐�Dc��F~�^ 6�
�X�c�jc'�^�(��Q12@�)]�sv��2p��ɂ�"<�"A�a�nKG��-��iQ�f
%��EB�` t��l�#*e�xr	�O�b�Ⱦ�0=ч$�
j�q�`�e��)3�*K�{C����ិ�b|9&��1T��@��$ˈo+�D3��6o��RW��["?��ɲ�:"2)�榟�G�T)Q��'l�iH�O�w����M5)�A�-ݑA<^�q��8��43��0�1��vz�AGf�¸����"'Ș�q�va��$�8#li�D'[���z�'$\���(�ɴt:T�b�ȍH�0��U��
4�Ls�	�+#s�(p��H�N�	����b�&�*2g�Y�ݘ$ITR)�")ҩ v�$h�%��K�@��'�~԰g�Vdep9֥:M(�녏x>|��f!eW��ca��>[�h�觃WY?�2�]	$�Պw���V�D�4kŗ/e^�$�}ƺP�ʁ�J�Pl�"�,E�0��'��@��Y��֎[&B��t��dj�1)��]� �p���bՈM��ɣy��0��k���LDJ�䘱2ʀ �M h�� gH� ڨ=��c���Ty�Jrs���$���|� ty��0b�u�[�oZ� �35��{Xz��
�6&��51BA�3Wߦ�Ї��H��a{�ې'�![��~Pj$�t �y�HP$��6I��ڤ���OP̙B끬4�n� (�<k�x�ad�D�-��z�� �E뵤݉y�T�� h۸7�`��S`ٷYF؝����	���;3G�= �q��\�|�F���Ț;1�t���'Dn���_�]T��pa��;^�DZW���j7�m�!T��h�C�&pHx��6�^W̓sIp��vG.N�h��2�T�*:����Ufy���(+[�R�:TQI�Gݯ̈Obx�D�E�_��APDdI.g� ����IL��I���y"�ɓ	�tP�� � [��A �D,a� ���ǄHpU
 ���Jv� ,ΣG@�z��$��B�D'O1`bց[�49��ǉN��؞�m����@�8~�$ɤ�ʏ y�4Ȧ�)H�����	�O
�� �O���T@�:zr���DE��f��ȍf��kρ��(O������h�0se��Sd/AkIZ����̵$.���q,�M���2���a	�l3"�����L���6���85�-�3韼T�f���`�f�[}��9Nǰ��XS㊗9�M����>B��Swv��Y�k�2xٲ�k�s<���G[R���g�i
pU`�`�M@�*_&{x�LE��5��d��?��A�7��T|Ex� .�I���ia.���:c��:3��̈$����!�ɋ�1 ��c�)��M��Q�ٝ���*C���0��ܨ�L_�q�Q�/����� �<9)�HsW!�z�L���'(�@cw�;qp(i���[�� �A/� 6����G"�f$�U����R,"ȑ8:w~4Yr�0Y��<�q�ţ3���3G�5��!fL]$IEnUIt�GF����"B:�(`",�so�P��İ ܸ��b���G���J���L�@#�͛-+����jʭN�|٤+D1۶��"�NF���Z�4�B����3N�3g��/=�F4�go/g���Y�C��a�<�nL,]��@��^�02xx�tM�w�*�3�d�)C��4@�F Nߨ�i��'OЌ�*΁1a2)�̟�O��s�ʆ�V�,h2�lH����y��_�U�|p1elåv�q(_6,��c��iO���
튍]N��ҤU�f�N��tAơYۺ� P��,OX��d%d"��t���g�&����ÔZ�d�Ab&B>N�h)��yV.T����oS�R���@�^��~Zc�H���U�Cg�рdCُ[�n��
��v���k�{��Z`f��3r�I����v�.�S9��@Ȍr�*��c�$�T�Y����"}2���:�k��Rj��DMH�'KҔ v���>	�[���M�'��SmJ��� � �&!e�� �qy��\���)G���{�唩PQ��@`�:@���FY�6^L�U��'�C���~���K麻	M���"��bS�d1��	Z��HKp  �O��Q���""F��0��ܥ%EpPAuQ�!�'Ɛ�$9	��JjyB�H�A�'�X!b\W���A�G/zx)��#�Oxp9�C�!�՛���~�(DB�*�9@�^$À��=�x��Z�u�my�lMe�|���A��O��ZpG���.˅S*��5�u�)g�x�Ѷ"OYja�@�"�n1��ǌD�2�b"O^�h���8^`œ$�68���"O$b�� f����L�;J���"O,�90n�=_��X��	2C�H�"O����	�\����^ p�
�"Of�za��c� 	�d��(|2�YE"O�dU���R��H���2gi���U"O܀8��i
D��O>:F"��"O���âX�0��*�!_����s"OL��� FI��!
�d���"O����y� E2��Ҝ$Nn�� "O������mj~P��5%���E"Oڈ �&	2 ��⡒�G���S"Or|�P����亷@N	�M�!"O\�H��\!����˶D�n<�v"O��H�!L�c��Ux�J,�!��"OBw�D�6İXcm�;:N�!3S"OE'�2X�xE��=i!����"O��P��:�	R�L�<��f"O�ū���]:��Q,�1c���"O��ui��%bqf�-9��8"O���V��B�\Ȣ�&�K�>Uʣ"O���H8�AX���1r�
U�"Ox�j�nN<.��C�i�!c�E�"O��&H�"������
��0g"O:��� ���Zu���J�hQ"O�H`v�� PH��P

�^-�c"Opy{�L�+�Vt+n�%�T]�"O`���� 1v��l�o١s`�Z�"Oʌ��@��%�P�e/��rGVU��"O ]�7��,V5p�I�8,DP3q"OV�8V*�3u��TC�&��c��,ȡ"O�H����CL�-�u�ۿy���B�"O� �����J/�A�
�|,ݢ�"Oꠈ�*#fB�A�jL#oF9�"O��b��̏*;�)Ӥ1YTqB�"Ob��t!V9�PY3	O���"O8\���+d<b�B`���4"O�m9�ۍ]T��uc�""�|��C"OX��ԪV�2tT�S�U=u�h���"O@����ґ�7#L��v�H�D^�<�q!�+0)R!T7��a���^�<W���x�qG�W�\�>U�K�Y�<�`�ύ*��u�1��5/�l�T��c�<YB�_z��	�7#ۍ>y�]c�(�\�<	��$aR������1�s��NG�<�1�ۭ#1�PK��D�X��P���C�<��K�昼3�Lx�x���"�[�<��B�
t?�	�@��T�v�L�<IVl�&\ Q3v�	T>�����L�<�F9�ҹ�6�ɢ]E��I�b8�C�fZ�'�r-@����8O�!�T#L$���H��P#mp9�"O �s]3,�pE��]:)P�Y�`���@q(x� ���R��S�Z�d�i�+O-UǨ��`O��94C�(�����A�3 f�����&���2�ܞ/��!"�^)�x�0)0�)$��>`�"١E&P�J�v1ƣ�%q���dɜ:��a��E@%y6i�������'��;\
|h�x�N1PmL�0=	UB0b;JH��%U���� �B�''�ƣ��o) |R�Eۻ218"��
�q4�L*0t�5ZԄ\S}�u�ȓE�y@��1�2E��F=d,ϓd�	���L�r���fA�@�Yx�,P���OZ��FU� �JE��I�W\���'*T�� �qn$�[���}� Q��×T�Pw��9'�y�� �����M$qL�O ���טN�h5`Tϒ�W����>a��%@��#> Ä/L4|�R"�C���� .A��B cs��.(45Q���	�| ��2�HO���e旗��4�I�O�h2e��508{b��#�HO�"�B%
]*�� �	QA��/2K�2��Kv�p('���Є��1ʓq���b!��Ir�x ��$� ��z�E۝H��*e(F��y���-tR��ᄋ�(T�x��Äɓ��b��I�"cR��(3<l�YP&*�d��9����-��Zd����OZ|A3'�����@�I*j�*�Zt!1x�e��(*��ԷU�`��K9àh ��U!E@yK�IV �y,Ӣx�(�� L��&ԥcf� ��~b)�ce|1 .�2 &]ExA�%)�"	��.Z�d�B�) b�> �]� ҇,�i16��)��[2�$a u�bnۗa�V�y�"�<$�]:� ��5fe�W��Y�ω#prYUӽE
�aXui�P�'�(�!��K��p�������R+�,�w"F�r4�q"K!�|͹2�A�y!n�CM�U%� :�(�/������u7D�O8�%7�3T	D�1}�3P����DR��O���s�]�'�8((4gS���D�Z>��hB+@u21�ش@�V�5f'�f���d�|�<����,Sf�X:a���C�����ꦹ�5*�޺[c��$Ў�c�Q�֑7*���p�cΣ�05ڔ% y�Xe��	�u;�<q�x�%R�~�Q�T�E��$J��֨mP�)!��.,G�e�� с@��t���ij��$�)hT��(Ӫ#=�v�Ɉ0&�u����= QD� ���?����܆Nn�k�e��f�i�c+K�e(�E�dA�� VD��ƚ�<���(�Lz�D��C�V�nѧ�O11���%'�I:ў� �GU>XB���L=m�F�I({�Vt�W�;��9J%�J�J�D��G��x�f����ܠP��$�$,�*}�Tt�7K�:��*���N�N��w/�|Kh9�&�l�� ә*p
�'���p�'1Q�
�_�hB��NL &���Q+zF~�U�*#�b��AW,l_�쀰�8U�\�jb�׾-p�&��^��C%nŪ"�hŋ��.iV����O�	���]-y��	��ո1��i�En^ ;�݂W9O\�;�O�_��)�Ac����1ċ�92��E�Ŏ_�1ȸ�`l��*�I���+j��u��͊	���	�hB�0�*��.h�ؠ�P�	�c^RP�g�@�*1�#�0Y�x�e�Hx�('A}�a(vK"̨��υ'�YRT'\`��Vd����i���Yo0܉�kY������eܺ�F�]�'��d�C+3;<\9)F�18˛v��7�3�+�*[*���vC̤Z�R ��@?g�(���"�=k<�P�En0�[F+�*Z&���I%�5� ��k�H��򮄥����H��N�'���32���'<v��-�?Y�S�G�����*O�r��eFA2 ���N[
�L��Ҫ:RbPy�����y�p�'��#5��6
���P���\����aݍ�^�����՗	0R�0�GT-�HěF יJGPi� U�S~L��b��nj��t��
6^�xeǕ�(�DثV �F1ꕱ)B�1<�;��v���c���Z���� >�1g�Z�B7������z`~A�V�J�>KVT���M��Z�`�V6h��X�c���M���F���m�Lx��Ȱ�W}>�І9���ؓC!aJtF�I�hq��9�
	Q�⑤@�jX��}IP9�6���d�	�$ t$��GRƌ�c��!|���̘>W
���͋:�9HB���o�k e �KR�qc's�ͣ�l>Q��wЭ b��m;���vh��}4 8�Or;��Q01 �\8�肸�J``H?�����u(N��C�9kZ�'���f����d��>�������{�ziCF��K�����m@5���ֵb����D�h>���͘$hZ��q7�S�U̪	�7oS�.֖e�&�؛v�<B�L�2{�,ם�c��a�&�"J�J�f�<O�t� �\�֎�-!\��c4J5�n|Y1�K�j�N�ҥ[�G�J@�L��T���ϸ'V,\SW Хg�����ُ]�x�2���9u"fn̼hՂ��e�)F���c@P�a��ثfM�_�|�"� [;
 ��~���E� -S^�Ԡ7h͎3��4�gk�;Uc�"�}�ՙ�X]���_�02�(:�Dޭ!A�0ER����Js�.��*�D@�Y6�Gj�7�4Q�R*��WE�:@E�z������-��b�w}�8��Z�8�����M�<�L�h5��*0�09$�N ��T�~�C��o��`�ֵ�hN]�M;���DϦo��P��=f����	�6J�h�V�lW��#��]�H1��(ӄ��mԛv��"�v�[��X�Q��H�h���9T����]�|��'"�p�s]x����\�`�L�'����</:\�be�F6O̬���i�S]������(S|~@�D��k�
�)��	!8�\�y$D˧�`�h�F��vⷬ�EG�h�`�ֈe�d��@���}�V�i�dJ%�~�8FI.�f0�,@NƼcp�[�HHE劉���6k�Aj9���$�	-&���0�*�$p��M��t	�P�g���B�ы\�u_"iRCVxb�$A�m��U1'�&2I~y��fO�V�)�K\wZ0I��{g�@�P�ÑoF�m�NO7yz�2��<���ӻ?��A��k�^,P�P�[iX<���=���UB�
��a��c��=��lx��<h�A�%��;l�S��F:P�sF��_��I�1��?��p84AC�:e�m�0�����M��0}����,C#�̞��H[�6d��P��00���`��6�&]�!W>�{#�\_��P�ݎ*��\r�N��#��Ue��&/��h*!NT7!�Ƣ<��Y]ưp!��<J�֐h��Zu�R�y3-�x��D�2��� ���6��)&^bV�!��9e���f���8�[��=6�e����n��6� >t�Q��[Gˋ*9<�UJ7���h��F�<p�(�qP��%{��e��12��� �aJ�2\��[p�R�.���\'}���N3?�9rU���\ʔ��L���UFT�N �Ojl����,7�x ��X$y
Q��$_�J�cjƃD$������$f�p!�¹%7����־S@�:F��q�&�S2ک6Ex�S�a�k�\qwC; :��n�}~R�F8���"�ä�[���ay|�ˑh�$k(h�*�3^�Pqafƹ���Q�F�&��v3��xrÀ�*���i��F�2$CG��!=0kq���N���!���uE���3�eeQ�هK�Z�ʃh7y�\�p��
H�A��K�:�lx��G�$�:��O�Z�t�<[�.�<�0	�"/�]x#jƵrq����3Q��t1��K�>�A�c��=Rr��$,�*Oa�$QU�1�|�G���Y��0� h�.P4y�+��v[�0������b�ZU�4�n�w�N�\��ʰh�� aI+j� 5����{v@�D됅D��=� ��0C�$_�8Tr'U�T�P�+�
3.q�Eh�&xLeՉ�;Y]:p�!�l
�`g�k���E��:�����N�~2c1�[9]Z0d��Xi �0S���h���*I��#�d��|ܪv���lf���O>W@Z9ЎG/n�z}��Ɓ�O��s5�D��f̊6,�Ԧ1�
�a���PeQ"�,�$�*I�@pXF��_ �x2H��mMT�F{�
R��}8w�	�����r#I�_� m�	݅v}�D���-0���U�S�'��]`���$��"I��T*�a� �f�Hթ�2�k�T�y���0� �#���$ Cq��:�o�V%طC0��(:0��8Dt��6Ɠ�v�4ӰJ�!n�m���Ɵoe<a�AG�~b�N'3�X{S�?c�yp���#N��Y��ȓ2m1������m��	'g�rdY�o�,�jY!t��zY6mg���5�ۭ*�,�EE EԡvƓ
Ak�k���T1��Ї�M3�iE!5�"S��,-9��@�40�^Bs�>����/��-��(w��$��JΠHN���n���8�L!j��4�qdU�+������t���F�ϠEP�BVF]�$m�T��������V{c��0_�D1�,�~Q!"���9<����K�&[ �J��*A�2EC�!ڛ;�N]�]@=�C�F�6M{��Z�:�JQ�UB�|���D�of�l	�ؾAI2:���om����˄V8� ��T����V�C�VTQbb����1��51�Z�!�H����1B���� �d8�YQ�N���5����!FC�)�`��'[�o8�AT�@��Uؒ��'�F���Azr��q1撲DP	Ya�^���G�=zY(�5O�<��mOVC`��D��%~�1�4k�"��PHE��N>|M�g�I��O����՜�Ԡ�����B�+4K�t��m�>D����Yo"�Rs$N�ט�3�������VB�3E�u0d��x��S�	$x'޽a�G�G^��˗Hݱ�a|��P3Z��!��-{��qӠ�Ӕ\����dsN��'Y��>E�U	��]���A6'�/~��Y�`�Y�
%���Fk����Ɉtfv��3GEL؞I�y�����H$��`��iͥCD���k�
c��s���n��D�p$�x�2�&@<ئt�V	�&NR����
b��[�ʷk��5�3,��!c�O���a�`�$Ϗz�U�%��=��I�E��y�����/�X��������%~�,�C�ɞ3�M��GE�\^t`�'�<���ZvZ@�Ł�'y�"=5�O-w��҂�@LF��A��)P���2P/+s@���;^L�R�l,u�ם�E-Y��R�P=���7"x�0ۣ��bЌ)� �4#�\P҇�3=Ka~�d3b
W�a�1�d��$D��y�ƀ!q>n\y6���WCK�d�6m4jw�e� au�\9��;s�1�|E���ʪOq�Q
�!�+�0>�,��	F]@&C�X"8C�iǎ �rr�m�7#Z�=@�ð�l�P`V"c��d;��^� P2���zb�-n��U���c��"\B:�0/
R����:�B?�A�Q��:C��\jb!�� ���5|��3OA7�E�r�-��$0�%:1��`à�.o�=��L� FS|��I�Enݢ�i�f�Ñ�;x��AB�!֯~� 1��K�?r���gJ�%GdɊ��S��n�ӡGM�|��i:t��=%b� `"��/qn��Ʀ�1(��B����?��F�lm���]�P�K��&S�hz�-Mh�	8q��<kpQBUa�%P�.0�&������@�[�TY��Ե(�y��E�rp��PG�Z�]=�hhflʬ��9�'Ġ�:A@�wy��)U�>�;�E�u����w'�5D�h�vV�$��=�T��pʟ(C�����[�^����
������q�����v�n�#�e��t��l*�z�/�;���稒.����n�7g(�qM���L�:� Đ_tΜ"�&@�լ��1�T�qN�u���2n4�1-Z��@���$?�"�.�*X�@A3(���J*��,1`����C���r�-!�6T��#�,�2�	M�~11e�
�`���[��xy�z@
�:����`������� ����� 4�KG$�,�ɗ��0�L9�!#R<!�f, �l�~R����)D��g��v���J�Ԩ)BԒ�O���]r��U�1��|���A,(��y��2��L�@@/-���bekG�FJ����	),1,�Q`hϯT�r0R��<r>�������ReKǣDM��kgcȪ*>6��hέP����B�٩�'T�@FI��D�k�68)7�I�'��MۃO�*6����C�qSV�&�0&z��H�.8�u�嫄Xl �"�!�N���%Z�L$��C2,h�Ar蕭>�U��'���*
�l��CK�=x[�����Z�����W?9����EY;O���Jm̓L��5!����V/��4C2B$��84� ��k���#ÄR#A��<��!�;��O�$� �A+z q�DL�K}pM��%I�
�haD���y�G�y[���hA�E%` ad�MrrM���	������h��y�0#\�\޶Y��g���M��?O����-
5;�����&��qC�§�h�͙XO�MI�.6�"p�1��Lۊ�ᵄ��'��y�O�X��͘]C�q!��&���k�f��d�ߏ�(O����K�jbp*�/.>�y4KS�|8d�BfɍOԢL1e��<�:���G/M^��Є�˗Q�T�c�x���,���g���,��i���)O�b.������4�6���Mcs��7М K��ܧa׬e��哟2�L,#��0�ER�-P"�m�; t�2G�1c�F� �=2J����*p�+�
6�W�N��<\���*ғd/�]C��C��X�l�=V��Q�B��W'��qD�كw���3��`'�E{�Ξ@��H�LνU��qv��G��Ԓ� A%^�b*A7z�<y�i�/�d	t�'�>q�Iͯ)֦��䝻5�t�{�׭s&p��-{!a�Ό��N�����٢@�V��p����.��Y�؉ �M
�h04���'�,���˵M�v�|I��'�j��eKb��A���Т
ԝp�a����CAH8R�9�P��F�����8`���#ځH��ߊ	���[&�|�c�3��ы��;и�pvB��O�M`�(G8a��÷��t�e�Lu�f�c��S��)�B��_��0�����e�����`M3
���Pq!;�?2�K�-�x	㡠��D'"�R��!ఘ�"�ֳ�����D�l@�hܧ7.!Wգ �<$�iν]a��!�a��_AjZ��B������}�����yOq񡨋;|<]�*� �*y�g$��]���@D���	رL��yN}�qh
9�~Zcٔ���/��MR}ȒnM�1\�8��tib�����i�Vy���@�H�
P�B��ev)3c�:{��$��.�P i�07����H���0�{ܘ\�pf�4(.����<��pt��۔L�P�)�'Lt�a��;l�,����81�u�TW�����V�`���$?��fk��P���dn�M2���
��`��H"U�Z�O��`�����}�%��hb���r���B4�>-���J�7��� ��OS<a����)4:8�m׸d�x�'.J���a�j��)��S�� �B�1�'3���ꅑ
e@����kQN�
	�kSJ��\�@�u`դ�2R�Y�,ĉDT�� �9$�4�b�NWr�a�Ƃ�j��Rv$%�-'��d7�'}n��"���&2F,@W�KNB8�ȓ�H)���p�q+Q�������H���4��^h\�b�\�6�X��!��|P��%I|��@���{�Ҁ�ȓ̆%����K�4]�"A��n�]�ȓ ��4C�/;w�&��uΎ�U|tL�ȓ]1܀��ܐ2p ��ˀ!�Fq��g����✣/o+�Iaѓ`c2D������!��1��![���r��0D��)�ŉkܺQ0�O�!~+��3'B/D��RMj�J�V"�)}���[��6D�@���	M�֌KAL��N�p�Y#2D��sb�T�p�;�P�WdI��C2D�k&!P9SF<�S@�&Lxx71D����c�=#��Xk�nA4T�B�	�}�����Ǘ�r��(�D[�kb�B�I���!�/m�,P��K�h�B�	�u�ЈE�܎  FAA� ӄB�	�# �P�3F��;-<`֕%��C�I:=�Yڵ�^�!+�5B�����C�	l�<C�y��0�THWIQ�y�	
�3��뗋иx�V���Jդ�y2䇳f)�i�vaª`lX�8���yr@&R5�C�B< }�5 �	՜�yr�˞}Sz4K֥ڛ|����Qb�!�y��@"X`��)��h������	��yr�#!'�(3��N�k�N�;��H(�y�ˌ
+$̈�T�Ew7�1T��y����h����kͦY�6(c2@/�y��/Y���*D�)V��� ���y
� j��G �?o��:�D�(�Z�2�3O�\��-$�^X�O�d2t����g5b��Dki���@هvJ��sFF�J�t5xI>���t��V2��ͧPp�]�G.K;X�� �g�nl����{尀��%\�by�t+��X>U���K�a��L�.F�T�mqR* ���D����@�g�$�,Z�(˅f�H�� 싌�	�4���?E��6B��1�f��x�00�JK��M�VHS����ȟڵHB��)���qg_�E~H� �K�'���Ʉ�I� ��	m���Ŏ�;��O&h����O��;��w+<]�.\�q��c6Jěm�bD%�hs�L�7�qO��<d�A��k�N1I��E=k�m�^�X�d�	n.qO�>�礑b8A�6܅L�l#P�tӞ0Z���S)!����Q	`�(uAY�r"�m9��ЋK>�b��9���O��M������ �.T�(������:�@I>�зit*��yJ|*�����JJR+K�oK���G��f.`�)O�)�w�_��1{�"���N~24$�.&:(��&[h�z�Q�N���?i�c`��`�OQ?	�+g��H���؟z5�z�C�/l\5x޴	U�'��u��S�Ha��s*����I �ƿ|����ۈ���*Q���0I �OP�$�!���9�yK�HK"�u�l��S�$h4����2]bJ�`�.h��˓;�v����㞐*  !���ó{f���'JR>E�P'��$��R�*M�{*���'t�Ё�N��D��fW	cāK��x�6��1d�S�I�.��N< �ĹT�W����9SY�a
�l�@�|�Ѯ�<���~nZ@2��-��e�Є����9CׄߜrI�C��&
L��߳tL��!�䐾T�a��JU�
�Ydh��%\\��Ү�	�?Q���E�(R�兎-츙�çw�B쉀I��ERH�HV�ژ6;�ys7��a2ߗ^�z��m��Hc`<��Ȑ!�y�a��sF�@�-�"D0�	L��y�C�c.>)����nT�Ԋ���<�y�iU��q���o��*U/�7�yRXe9�E��g�m�(��`G��yb� YH���12}��NЗ�y�P��xA�T�g��a�y2ƙ9+(����1f�$)%��yrNԛjg�⣭�95�"��"�y��L�$�p�F�A!4�4��ZQ�pB�	�qM�p)��8K�T	Q�+\3gB�I��n0C�L�C$L�#��,�C�	�~�@)�怑�e6�Zt�R�2�B�	6Hsjt���X�u7���p@P�f��B�ə}ް\�ԫ�,1O�)J�
D��B䉉=�!z�!-l�m bʌMhC�	*K0b\�Ə -��"��
� VC�I��!b��9�`�*�	��>C�T]r8IA �yt��k�5�C��>����.)+',�*�	�5V��C�I�o�8�q�ǔsL6q ԉ�<y��C�I�s�^` �AO,E:F肨	s�C�	�ne^��(���ɢÂA (ʮC䉱1�b��T��9��T��S�_�vC�	�c�z`�� E2�@1�)�d��C���PPe�0��<c��͐#a�C�I�qX�H�/ ����"eصRC�	�4?z�e,�I	������pw*C�I�><�H��'���9&�F�, C�ɪ_X5��
ˤt�����IO�lM�B��8�#�D:b]�y��P5�B�I�^}.I�7m�a���8��N�h�C�I�w����ܝ�b�N�zT�C�I�qf°��[7ߦm�)M><�C�I�BG���h��`�n�h	�j�C�I>b/@d"w�^;� 5����(�ZB�	�5�6�ӳ��\ΪЁ��ǋCK�C�I�+_<x8��V�!18�HC�I+)����ħϻP�4�-M"c0C�)� x�j�.�x�0�_<Y�\0�"O<�a+^�rE��(���|�0l��"O&��1��&y.< �B���a"OJ��g����G�G|(`"O���&d9��������ʖ"O�i`w��(6bH��!�ߥV�dA�""O��坭q�
�JSf�N&�yb�ƃG����j��BԬP�taB>�y"�ga�-R�z<pc"	)Wm�9
�'�6$[�'R��.8��m�#= �
�'TeYt T�V���FW�)��i�'b6MX$��M���G�wbi�'�:�����g�xJ�,P��
�'�>�E�����j�Xd\�
�'WV��p	��r�6L9�W	��Dz�'{���	F>���,����p��'��l�
v�� �W� �Y�0���'`�T���l˴�X�L�W	����'�2���>���	q�F!W�j1��'�P9�@�>�p��C�)SG�u�
�'�H��s(ȱ�Ɂr��2 :���
�'�蠉ET�r�Dۄ�į�JI�	�'�N�C�NF1m����ť�
4�D�1
�'ېY�E�Z2�%p5.�%,dPs�'ڨ5���a�&��J߀) ��
�'ľɐ��O
zF��d�L�<�I
�'@d���f�5�\�R#�֬܌�X	�'��USO�=��1��U��i!�'���)���B���s����J�'��]�Eg�:!���iDA	(I`%B�'@��qGK0����@R�5��
�'cP��Q�&�c��\�|p<�CO�<y���3.����	�F[�����N�<�"��.ri�O_�H�sk�H�<Y���h�a"K{"�;�b]�<yA�W��&`��ܔ\�p�{��a�<q�Zf`HhѶ!�����6�\�<i�>vQ��yS�� e��)C�A�<Y,R23� ���]R�$h".h�<acH;#�$����:X���1�d�<��̜�9V�.QѰ�2�*Ĳ(�B��-Ζ��4���WbNE���(cXC�	4Y/���D�P&| �Ec�b�(�2C�	����5B[���jD�M��C�	<��L!R�'|����͋*a{C�I�����t'O��$Jz�B�	u�} re,|-��u�ȌX�B�I� ��U��EF*g�( qkǒB�	;"i�R�đ"+��T�X?4C�I�Yysϝ�5�����bT�9�C�|����QC��E�n�6���B�	�O]N���#���ʃ�˹i�C�ɝ\�ԡ�@ZZ�N�iv/Ƚo�C�#e�fy
���>�L\Z5�.QΎC�	�UG����V�@,�uO��?��C�*����'obԓg��W�rC�	8k��0���`Ll:�%��zC�2�rš�dن.J��W�!B�I�S�:, �L�Z%&Ia!�9��C�{-8$B���7fi�5�0��C�Z��%�7��&vRq� �=O��C�I�~2�:�՗Tz�C �"��C�	�)�Vh#����Oqd����ӴC��8�&�%%ڃ_��e6�P�Lh�C�)� p ��C�Fڴ��U�Ī{mz 
�"ON�JVn	2f�M���+~N����"OH@XD
�#R�BMH@�P(;g��c"O0Q13M�Φ<З�R_�:�B"O�Ma��[��VcY�=�ԛb"O �pacF:;>0p��OB����hE"O茱 J�ttr��V/�X�}��"OvL��c9P&=�n�SAfD�R"O���1��[�h*�F�n�"�� "O"�`�.�4��a�	^���H�"O$��E�I>, ��⎥~����"Ov��eI��8y�
�2p8Q�"OX��G�ƥzr��blii0"O4��N\86I)r�
�5]�$"O��8U`��>���Y,rV:C"O���S�}j�B��X���9#a"O�ș�չ3��|Xѭ�h�����"O�D�4e�1��Ta$b��
�0x��"O2ku��J�L�a���UcReq0"O�(�Q��Ō���.V�,��Ԙ�"Ob�����YB(�&��./	�`�g"O���٦dC���ɢ/�4e��"O> � /o�p�QfS,1��X��"O���@Y���3 eΧ�~�i#"OZٱFe	�n� �;2��z̴h2"O Q2I���<3(�
R�\H��"OAr�S�O����c(���q��"O�a@ɜ0"�d��F
���"O�I��E*+Gt��6e�l̄��"O��:�Ǉ F�l`�!�8C(��"O���e��,��������£"O����iRp���ԪaJ��"O~����#r�(rD��3-�P�"O �� �@+w�D�#ϐ��Eza"O��j�$Ɠ����U��!.	�i�'"Oz��aӕI�I�0#Y^�T��"O�-�C��J�4����	�X���"OT�85��>x���q���FB1[$"O���B%S�X�ŏ̴P;� u"O`���8:zp���OÖr)���c"O�$s
͸/� @� F�n�9B"O�"SO�+f@�İGE%u��a{�"O@���4NU88P�"�+��`��"O,��3p��h�!�p~��c�"O�� '�u��)�ª�/b����"O��+p��6��Ȓ%7Jj4�"O �j#"ݧ$�J��X�Yڠ��"O�=P�G�ڸ�&��&uk���"Ot�!ŋ.I5:�0a�Ak,I!�"O����l(|7���E�e.�dCA"O��s���.�T��P�O�q�B�#V"O� ����=~��2���dM
��"O��P�XH��b��a*`;�"O��)i��LI���,K�E�5"OH�Pe�
����M{~�;�"O�,j��'B�(4���. rqQ�"O���%�,&qr���U88��yA"O�t��}���6 AF-^��"OJ�s�A�2)�9v�X},F��'�bGQFt��c��=<+�'I�$XEB̥%���L�qݤ���'M�tɌ�0������fi���'@�B�/L�/v�z�. t`���'��Az s
��A��
�pt�
��� T���S)r��`@�W���p"OR�h�k��J,r��a-�r��}s"O�e��	��k'�� ���x�"O8TAp)���"&G�"��5h%"OVMje�k��E�G�j��C"O+�۸|��D�Rm��d܌{=!��M{f�Ir�G	�&Hh����7!�D�!J���#��q�lp%��!�$�g�b�q"��b(hyA�k�R�!�$�b��YD.��"d���O�U�!�DخpC��yW+����I�j��P1!�䐧#z�P3$�-0A�.�i"!��Vn؊��
_����� !�1�
�)�Ũ 
�BmN�I	!�Dǃf9��0y�|�F�֞_L!�d���L@"���`�(yCj�;!�@�tC�ᡑ%M�"�l��2'�%�!��#�6!�ć�l8��F��!��ο5��y
�虻\���9rf���Pyb-U \�St+�S|� [��y�E2yJ\%���E,���	�y��(���0��h��k�NЫ�y��]%Lq �ҵ��:�0@�3�ylƈnŴ�f���Q	wM[�y2����(5�N�+� �׿�yr�������6c� �dX7���y�,A��y��S,M4���.�y�Ԏp��eˎ6vV�Q-���y2��ML�l�%%�,m
<$٢��yңF<s�6eq� L�a�n��B&�y�ˇ 0  ��     �  �  �  t*  �5  4A  �L  �W  �b  �j  �u  �  �  d�  ��  �  5�  w�  �  ��  Ӹ  �  X�  ��  ��  A�  ��  ��  f�  �  q�    s
 � & ! L( �. 25 u; |<  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��Inyr��-qd܋�FS$��Q��Ԝ�y��˪=7&}�)@
HZ����2߈O�}D�&D�=��|{�A���تI� �yr
��l����k��I�a@�e}��)�'s�T�:g,�(5(�K�
܀$�ȓJ�`�6 З`C��[��84��5��2��yr1�L�E�F�`F�D��݆�n�,m Gˌ�ZQ����<����>^�䨍��Yt!�:U�ȓ_��!���8%Kڀ� �>tp��ȓkb	�q�+�Y��K���@!��czT*��}M
� �+�ifN�ȓcA�|�ҏ>	W����g�n�|��X��B���n������01s���gE�j�:���A  8��K�N�2G�U,q�҈��˅�/�<��ȓ^&N�ypgR�[Ěq�Q�lg����T;4)����j<̛��)�LQ�ȓ44�����gP4�&H	/e*��ȓ�hY@�A:�����
�az(���2O��z�L@*_u�TA��3�2���S�I� p*���&oB�U���J�~B�	$1װԑ�H#If�O�9 ��"<@�)B"�@$a	F���f�©h#�^�<��f�([803"��(S�I8@b�H�ў"~�)� ��h�.ב9���i����<�Z�"O<�K%	��6��%�g��&r"@<"C"O�ёe�
�3c���w�"���"O��B�&�$�F��@΁��H1)R"O�h#���'������A�
�W"O�̡���9��f��������"Oj\j��O"� �Yqa &ct��"O�Ђg�pj'���-��`"O:��F��Jɷ��Q�����E�G�<!Rl^��-xAA�����4�M�<	���*��cfچ��;�d�<yb��
'~hU���9Q��ma�<�g�L�K챁���*2�6�;���^�<��KݻW��U��I�#?d޴ˣ�C]�<���#@����fJ�w�ΐ�aO�C�<!C�,?PnP��I'GAT���C�<���Gi(���G���5���:&�YW�<�2M|�1N�w���!*V�<�n	�h��#M�u����%�TH�<)V!Z>~�2��䅉7[ ����E�<a��ԭJ�,Qk�B�1eoܝ;0�V�<��f�o�zE��,&�h�q�SO�<��Wa.zT��Ä~{�xkp��P�<�d?^���Jt��>s��h�N�<�p�1P<Y�'Q9k$0m8���a,B��=q5�X�R��,[�!��mU?�z"=���T?����%�}��ԀH�P�*�&D�d�%��'m�<���"�rFL�7f%D�世a��p�z���Ј��"Q�7D�D����/Z�DS�	ΕQs���b�Т=E��4n9�$���[ {Ѵl�r�(n��	���l?ɷ���UIڐU������}}��'fT�!	�w�X�����P��4K�'�P(8���Ԉ0C�L�X�&,[�'Rh���R�Y��$�b��XeU#�'W�4s��L���#����!oT��y"ˋI�n<�e��� �L)�y""W�k.�uS!�I.g,+W �	�yR�	�e�TҧA�����/H��y�Y'7~E���	�T���d��yb��kc\P���Z=j�*��T�y⇒�Q�2�c'�/].x���K;�yR��3c���r/��+s��i�'��y�@3�vYA�"B3F=r��3肆��I�d�a|�L�z���ģSQNd�ï
��0?��+�?y��7?������@��%���h�<Ac�+\�(�ꐤ�`�Ȭ�gb�'�l����i"�h�D&R�lQ�u��x�!�$�gɠ�k/�� �A��8��299�⟢}�� j���≽>����ǎ@�<��,ɡa<���
�8hf�T��b�dQu8�@��E xJ���XǦ���*O<��W��?Q AŴI<�9�"O�QP&D�N��Ȳǂ�o<��y"O����K_a��ǂ�$i�(�4"O�`���M����a����"O
���DЖA3�L���ߒro�p��"O|		�*&Ơ����C7n�������(O�O�� ���|��=��Y)=�8�!�'����w�x�R�dL�<ŴL[�'�
���/dC�5�*��@(z����x;Q>��e�E	nG��Ǡ~���*P.8D��0gC��X�������H
�ن`3D��9�&��|Xc�dQ~w�iˡd#D�� $���bX;"�@���9R�:�`"O���CVkdYY�&[���"O0������t�E>(�H"O�A�I]�<WJ�Ãٳ�J|k""O��A���?�p�*r��G�X�W"O��Pg%Z��X����&'2đ��&�S�	^�Gd	k4�N��ڃ��*Y!�dD� �����vw��[�8<đ�h2	�QڈY�T1�j��P*���L��I-5��9��� 3|���Z<y7(��tp���2�H�fHn�<�A�Qu��e��X�L"8��on�<�5JAY�0�C/� ,Hb�ѴɞS�<�� W�|�v��2;�^h�g@L�<�&c��TV�M���.u��ma�}�<S���!��djbL�n�\�C�z�<�!�L�^fĐ���Y�W����k�퟈�D�)�0p���҃0�,q�4�F(��m����y�ڎ`� գC�F��`����GX����l��ͺGLp�ѡ�1��>���1�y�/�E�0�b�%9d�X��H���yB��+1��Aa�	F���C._��~��'���+}��IQ�gX�4bÇ	�V���p�#C%�!�$�#C�ԥCfG�q'���h��B�Q�,Ǔ1N�YE�"�y��S�D�څ�ƓG_�<+ЌS @/z ��U�<�T} ���A(<&P����jvyH:S�r�<ɦ�(~F-*��J4�����*�o�<��J	.U��4��CP�+�\$bŏIk�<����N�f�

ן]�ZC��i�<q�%�G�Z�a�ph�l_h�<�!)��gOX��цНEKzi�2/�y�<7�3v�E�1+"�J��v�P�<���y�� �-U{��LZr�<� \�c���H��חGjv���An�<��J*p�،3�O�~�US�Nb�<)aFD����O��G�hК�IHH�<���%��=鵬�?�*�� i�x�<Q���G!�5�4�Y�%4�t.n�<	�%_�i��p'��79��ԡ��UO�<i���3��[Ã��VEB���P�<y1�\.z�X5�3������dFv�<�����6�![��0�{� ^l�<�4�J�Q_v�+Q!F_�-AA�O�<Y�%
�ł�ş�F�x�dFu�<A�SK^�zDl8�j�H�u�<�C��4GD���##	�
e��[p�<�'"�tt:��-�3D�6��.Zl�<)��3�0)(��P�6�Xcc�Kj�<���D>2^B�H�&;IH;5`If�<��Q�΢�b#�ڶ ��lÑ�_�<q@ˏ�QRry(
;(F=�G�^�<���k4rpr5H�`����T�<��C8[����F�����fRP�<�d�L�	#��
8�xԺu`R�<���P=�|�R�M��@X���O�<�6bV	w������Vjx�p�#�I�<�%��S��D� �_6zTPp��N�<���n��%�D��4���q2M@N�<ѡg�l�&X���]16��Q.�J�<��E��P�Z�I�Ҧ�)1&�a�<�'��������n�x��ZY�<QA�07bF�R"�C�RS����LX�<���4����bX�V�:RF�
l�<� l��J�&X�tȒŜ(pN�a�"O�MR6�T� Y�!2d��>d2��`"O<Y"��Ħ<����ab�$(l�$Z�"OI��!I!#lXZP4y x�c�"Ov�
v� �Y��(�6F��t�P7�'T��'Q��'���'42�'p��'6�}�fM�AX<�bugҺ� �"�'/��'GB�'���'Y�'���'B6m���N���b1�Id�V���'���'���'y�'�R�'���'_�$��̚.UJ9�j��nPJ���'�b�'\��'���'�B�'���'t�y[��LY��AGżG������'f��'
B�'���'�r�'�b�'�x�
��@U�戩�c���8���'�2�'�B�'MB�'�B�'���'��C���3yk�X�rf�8�4��'���'��'�R�'r�'���'�P��NƜ	6��s��GZ�@Ɉ�'���'>r�'�B�'*B�'�r�'����ӣ�(9��҅�ɃO�Љw�']b�'z��'���'��'�2�'|HZ�X�c֐YS�%�j�&�Cp�'���'CB�'���'e"�'���'�\,I`��Q,0ВG�DaNE���'9�'"B�'���'��'kB�'7����� p%l������*��	��'���'���'���'3��'2�'�X��)
Cǈ��&���tr�0��'���'	r�'��'yҌr�d��OL� �2Q�}j���E��)!�Ky��'�)�3?�մiЎI���E�$��Lp��|v�I��͕��d�Ʀ��?��<���<��� D<^�&�
�d
������?�Ǉ��M�O�>��J?Ͱ��><�vD�C�_�>�\�b�*�	��X�'��>s�Ğ|��z�߹U��mz�*"�M�����O��7=�.Q�F�Z^|��oţO�
H���O��$b�4֧�OI�'�i��$ςA�������0&��52���~���n�k���\�=�'�?��@_4v^Ԩ£>\�����N��<�(Or�O� mZJ`�c����`�x����%ێ��A㣄�x�Nk��ן���<I�O�]k�U���A!�K+@�ĥA������cG�iK��7�"cF�����K3NK�J� �zWIH!gId����{y�Z���)��<a
�6`�Ru�7��5�bh��<a��i����O��nZc��|����Rs�|�C�5�TI�ĉ�<)��?���
E$x�4��dn>5y�'G��}���E�i,,��a�'I^��� >��<�'�?����?i���?�)%h��ą� ��\���P3��$�؟�H`E�Ox���O*�����7�Μr�A���������P�'B�7������J<�|�� P"ԈcϛBQ|l��,@8��� ��Q~��Y�p>P��I�#p�':��>��%(`+�0!�8(#�m'8���ԟ0��Ɵ��i>q�'V�6�6���g�li�`��,k$�S@��e��$Ӧ�?�U�H�ߴW�6+f��E� �.kV�$+$�)]�t�Y��]7�7�$?���f� @��pܧ���@
S� ��X�e��Ki�-��<��?����?����?i��t�3s�|��,+6R=���L�I���ܴyˠdΧ�?��i{�'��V	I�>���B�KZ�6/�!��( ���=x��|r��M��O	H�ōD8L�#D����ˁ	[/� ��:B��O��?y��?���CNzY��T����v�\�gˀy���?9+O�oڱ2�����ٟh�Ir�d��� �E�N8^<r�OM<�y��'y���?�����S�T��M�#]<Q�D�Ӄ�8��p�t��;3��탒Q��82�
T�I<<�Q��!W�X-"��V+S> <����ğ��I����)�ny�x�$��"/]$L�t!��ěPF�4���$�O��lZC�i>���O�LoZ�%Wִ��6Aq�8s��\�bx�Pڴ �&�. �v��� !��>Cx��\@y�O�>n{z��&��-�<H ƤZ��y�W����ID�� c��O��⧠C����4h�rC.Oj�$.�S=�Mϻu|Υ�c��;(	LQbBz#&�X��?���x��$�J�6��5O68�D���	w�I�W�H-S���`�1O^rw�E��'��'������ɕw���q���%���;J��W����	ԟ���🀕'`7�9fP����O���� �@������/Z;T�Z�tүOj%m��M3�x�h�*8605#�>uҀ�;b`�1����?x� V�� d����`K��c���׺W��-{�,��j�����ݍn�!��R�����k�D4�*�(ޜ����'�6�2x�Z˓m.���4�o��j��@ e�U�<�пi8�7MŦ-p�L��	�'6( !ҫ�?�wjEsb$M2%��lh"��4j��'��������ޟP��ʟ���� �j�p���B�E��(ɂ�'mv7-�pAL���Oh��$���O ��E�Z�n��*��L�\5[G��k}2wӎ�m+��S�'i��TH�%Q��R+U8Y(��gyRH�HTRY����'V�	;4Ц�"�I?`�Ε��%h������yڧ*����q���T���P�.9sV�;B�y���4��'�R��?1���?�����S0������@�;�S,.��E��4���a��(Y�'I�c>�� ���cT�T�\"��5	�q��:OD���Oj��O��d�O��?MI"Aݢ	�Rxc2�T|�Yy&�Aԟ4�����p�4�4�*O$mmO��,aKU� �$���`�ETH�I<��i�7=�2e� ,x���i;2XBiJɪ*6C�=�MQAm/���$X!����4���$�O���׃oB5Ɇ�H1KM&�Rd�F:���O��#`���Ķ!�b�'2P>-Cd�٘������6k��yĄ>?1Z�|��Ꞔ%��' �@QC�.��cڼlb��*��� N�Ƕpx��J:��4�4��/隓O"a��H�dD(��Mݔ3���O��d�O:��O1�`�nf�&G�'�fH����;l�(��'��d��y��'�Bj`Ӫ⟠��O$�$�G���8�G�[� p��C���D�˦Q�C����-�'�\{R�B",O���J٨}��qT˂S}�Q�0O�˓�?q��?����?i���iD�HQ�	�!�/��#B�y9���Ӧ RFCǟ������$?�����MϻL3483�M(�pM�J�!������?�H>�|���:�M3�'�6���-S 
�����CG�Mʙ'�2mc�a�ߟ0/������O���U�?��((3j�*X���`⇋6-4�$�OJ���O��*4�VAL�^�'�2+\5dƼ���"f���Q.�+g��OX��'���'��OTD��Mb���@eP�d?��R��4�w��>`9�o�-��'r�x��ʟ8�ޘ%%���G��$���O4D� 9���q0�{"��9l��ٳ�ӟ,��4~h� Q*O@n�c�Ӽ��&E�9Њ�� ��=�sl��<���?���i	��xS�i/����!�П�\�O�d� yA�i;K\	��%��<y���?����?9��?����CK�� $��MS��xg�K2��Ӧ}˥����|���&?u�	f�2�0*]=[$b�s�)9L��ٮO��n6�M35�x���.����EIO;%ĦU
QER)[����FN=e��IIml�c��'�U&���'�>��6I��(R���e�J��L;��'��'�����$Z�h�ߴ\�0z��u|`�r0/�(�)f�b�͓����d�u}�q�HoZ
�M#�S"lg�U� 2#��V�
��J۴���XZX4�����O���?adY��*�ׂE�d�1�y�'�"�'��'+���pj���Ua^��2I�Y���D�O\�d\Ц��s�|>��ɛ�MO>���J8�ᄪ��X�b�(� T<���?)��|j� I	�M��O�N4"t���!����NZh������O8@SH>�)O��O����Oʨ"�-of`�X���ܩU��OJ�D�<���i���'���'~哀k�	�S�LY�tx��l��W>�����֟�	P�)�b���dI�R�U;l�P�So_�/v�i�䁃e�L]�)O���?au�.�Ć���k@�Q���,�"@�m����Ox�D�OB���<�÷i2�Eұ��f@�qʳn]%K�>c&#��Y��*�MC�rn�>���i��H��/4����߹H�p5;���zm����n�x~�ˈ 4�����|�I�8v�z9�6,�TG�dcQG�w���<����?���?�Ȧٕ�����80��������
�%;f�R6mX�H��O���:�9O*8mz�5Zq�lq�r�дM�!bs(E˟��w�)��n"	l��<�$$K�x�ɑE�9�����<��n�"R*�� ������Ov��ɤ8ʄA�w.12
�щK����$�O����O��V��	����'b҃K�i����G��Z�,0
�*;B;�O�y�';�'��'���sRe�_�Bd�D���Jz���'n*�M�f%q`���"���?i���'h���iO4H�v���ӕ9Tx8��+_���'Xr�'������7�ɟ9g���+�C��!�ß�h�4Gi��9��?y¾i2�O�nR�3�*�{��QvR|H�$���z]����=[�4�����!���4i�!w���FtD-1Q*=ឌsC)Ԍ!Ԫ�$���'(��'�"�'��'����h�2xmB��`�I	J`����X����4O��T���?!����<9����4��:-@�J��A�K�%?�ɉ�M���i�O1�"]R�(�'.DHa �[H�K�E=�|����DD� �t��\�O�`!��5�D��Ǜp�P5�Vh��������@�	ڟ��fy��{Ӑ�P�o�O�$;`P�WhY8�D�+2l)�=O�9n`�F��	��Mˑ�i_�7��5������(���b�Byc�Hx�JvӔ�Z<�9pb���L~*�;^�pm�勊�9����'b<�`��?����?����?����OV�� �ЕW������;{��zTU���I��M[�˟�|���}��|2�V�m�B�je��0��4��#>QjO�,lZ��M#�'u����4�y2�'Ul�Ж�V���9�w)�(jvtyb5.fQ�I}��'
����<�Iϟ��	���a�K,�����>i$�5��'��Z��Q޴0�����?9���'i���C���& W.��u��/^�P�'��.��&�v�-$��S�?I���*vtȔ;�e����R�);�~�k���T��'��t-���lI��|�IB��Xa�I�!60�Xx*׆=���'���'���Q�Pcٴ)��}P O@�Dz8�t�)2΄�Ya�����̦��?�tR�, ش[|��R<�QJ`���^g.���i��7m�	
ݾ6�1?�%�-��I�����  ����8����b���Z�6O(˓�?9��?����?�����K�2�4-p�K�&�� @j2
[ <m��{�~���ß��IV��ß�����k���!s#,0��M��hC�蒧ɛV�f&d�||'��S�?����"�(lZ�<qW�	�h?" h�Q,Y��e�2jB�<��#C�&|��[�����D�OL��X�(~��#��!�0�I3 M5y��d�O8��O��gܛF(��JT����`��Π(8��V��%�wh�-8[�O���'�v6���i�O<�� �/Ld �LG%-�Z�cYl~�G��J��,b7ㇳa��O���ɲa����4|�FԢ�n�;p��<��#a��'�r�'������UA�#6�YB�DX�^r)�5�ޟ���4�����?��i-�O��đ+
�Ųa`�/X5��C>4����즭��4W̛F�S��4��D�-:8��')
�p �Z��R�K�J2w+2�p7�#�Ī<����?����?1���?���Ǎ
��eC�S��ȹV�&��¦�@0d�ty��'��O
�!$x-�V�z�u�R%�z-��x���pӮ�$�b>�RŉǞ$t�<�G��S!�E�7O�q��H��QyRM�5�-�	�'6剀{� 
�Ιe�L� G�N�-�	����Iܟ��i>=�'<T6Mޝi���3 �(��'�F3oDHiS%ۇ�����ܦ��?�PV���ڴ�F�yӎM�A�C���F��G)|y07��7�6�n�@��;.fe��O�'��D�w����XX�hq2��b�\�ڛ'��'=b�'�'�����kf��@	��9��t�bF�O,�$�ON�oZc��'HJ7�4�D�&jXs4��!�~�{ÎтK��$�|��4V	��OE攡��i���#�.�P�d���(C�/D:K����'	 �dB�I�`�Oy"�'��'B��x?`!��$��� �K���%x���'S���M�eM�<����?�)�%f��9򸲡�؛]Lڼ1土�ȭOZ���O��O�S�~��"X�6yd��u푦;�Y��᝖p��lp~�O��������R�%>V:����\ɚp��?y���?�S�'��dM�]�⇕=����Eń�B��E����c||�i��&�'3�'�
��?YDF=AK�t�@�&F�ѕ�T�?��)�j���4�y��'����� g�9O����^�-w�0�EM��]<I0O�˓�?����?����?�����tu>���Zw� pbV�ǿ�tlڠ9���Iğ��	D�s��A���K�m�3����\y�ȥሼ�?1�����|���?a
��M�'�����K�<BF���
�>�Fe��'��Q"4�l?�L>)+O��O��Al� 6���d�5	.��b��O.���O>�d�<�ֻiyfxa�'�b�'��yjV��~��X���x ��%��IZ}R�'7��|�S�p�)��FM�sQ�PXu�҉������fY��n��b>I�0�O����;���� �8\ɳ���6S����O����O:�D9�'�?!�H̞B�.P�����a����$���?v�i��,v�'��&sӐ���?6j\X�-��X����Sl�6���������	Ê�ݦ�u�i�1�ģF�#�FL[�摨�\Ł�f�C�t�$���'%��'���'t��'�]8v�ЉZ.��1f�=RKF�KU�xIٴ}Xp�B*O���"�I�O(�s����=*�B�C_?zxN� �~}R!t���oZ)��S�'g���@S��n��1)��Szi<`�wo�S�9�,O䥱���<�?)�;�D�<)�jR�@�Ze�B딌C�X$��̅�?���?����?ͧ��D�����%�B���c�C�h�v���Ï�"�������9޴���?�]�������k�4F� �a�7c|R��LD�^��HA	���Mk�O~��P���������w�z�Ëڤ=�H��u���"�����'�"�'`�'�B�'��j��R�H1,����(�X�C��O����O,n5>��џ�ش��& ����(Nɀ�R��i��غQ�x��i�� nz>(T�Tզ-�'3L �QN؎:n&`ҡ\�Q����`ZŌ��	&P�'��Iԟ��	ȟ�	7��H�b����Icg˲v������'�"6T�{x����O���|p��4��QȄ��(.a	E�v~R�>	Q�i�6Mo�):e/[�sjpء�'#��9VI˰Q�"��DV*Ĺs(O����?9��(��ЅtjdQPqIN����'��3r�!�$Yʦ� $*߳,�͹��ͦr�>(x��A�4��-�'��7 �������ڦ��-�"F&�{��3W2p��c ��M�G�i��ưik��?"�&�ct�OR2P�'
>M���Βax$��I���ࠜ'��If�����A��qz�
�JK�	��ê�M�t�K�����O��?9����S��PC~(P����!"��;w�i�O�O��3�i,��1��Q��AG8%�dM�p7zX�'�(eڠ��П����|�Q��'T:�3��F�|m��'�"�ٰ	Ó[�v슉l}�I֟t�ŌHu� c�&%\dIp��E��
�	���m��ēc��˕f�Y�k���V�f��'� x6��h�٠���Ƀҟ̠`�'@ )YN�H��P�&O��X��'H��z���2T��]���]����R�'��7-Z�I���כf�4��5p#Ȁ(j���!�Ě�g�6i��9OL���O��d�u�d6>?��J�a��'2�� �:f��2��	�CS���Y6�d�<����?y��?���?A��'QV�0� .���4�4��d]̦Y�VH�柴��럈�2�Bj�$A!�AG�x� �34�	�MsE�i&O1���7A��)���V�vر���XR�!3#�<�a�C�r�������D0AO\u)`Ƌ� �E[�Л[�$�d�O��D�OR�4��˓k��0V�R����8���D;@y���V�UGb�l� �(��Ov���O�plZl�Z�q"�Ō>f���B�Mj�qC�E�}�'|4� @d�i�K~���v|����eP���n�Hy�d��<����?���?a��?�������d��c�1�P���O�`2�'7�h�D�,�<�óiU�'��HG�CM����G�G��m�Қ|B�'L��'������i��$�OV`�n� ��ل,�V]���(JM)�	���H���O���|���?9�x�  � (�)�41C�[xG�����?�(Oz�m�
r[�1�Iş���~�DL��)��d��U7�(% M����Mn}"�'�|�O�R���-� F�e�j�"t&@�a�x񅙤K9P	��O^��I��?A�+5�$��j`��	���2�D
\����O6���O��)�<��iU�M�E�O45zT9k�фMl��!"Y��#�M;�"��>���Q�<�7�¶1,
�qQD˝h3�ph��?�f��M+�O�1��N��J?A��ĵ(��He�� ��p� a�H�'u��'4R�'"�'8� �r�v�6�,�K�N	A�����4B�ش���?�����<�S��y��S?X�\;��Ǫ}vЫ�J��JN��'ɧ�O����p�i��䎭�v�!���T�a�A��4�$�:�r]`�C֒Ox��|z��"� Ppu�Ԫw@*��Eȉ0��?a���?)(Ov�l#�@��I����I2iX4��O�%�"����hd�?a3R���	��<a�
�-`�i�� ۩>�@TR�.?�taK�r���)�J�@�'{���� �?YPaTq�D�n7h�I0�H��?��?����?Q��	�O�q�Vkޔ~~�4���߿�h��qN�Ov�m+E��'��7�7�i�i�F+� W�%��,!.��1kz��I���4f���[ݴ���(����O$ha��
�`����axӖ|�V����韼��ɟ���ȟt�$b��k�8M�VD� D �3`Yy��|��`0��O��d�O�����č�O*�\JV\P���|�D4�' ��'�ɧ���'�2��<���P*4<H!������E'�@�	#RRlܢ��'by%�Ԗ'Gd�`�C $�a�6m��4v�'�B�'�B���DZ�8+�4:L�v�n!����fIH]�SB �gv�r��
��$@}��'�w�~<
2�9fU*�
��0G,��kR�X0�M��'�x@���Ss���?Y�]�Q5:m�s�YI�Z�R3��x���Ɵ�����l��,��D�'m��<2���{��3�h6~F����?��5��ƭʉ��$�'� 7m-�$Ϭ����	�w�T)�b��`���O��D�Ot�䖨=�H6-y�t��1��H3d̺O�������k�F�[�
��?���2�$�<����?!��?�:Q� ��U� .E�Hh��
�����OJʓ6�& ^�v��'(R>�:&D3��sF�6T�r=a�k/?a�]��p�4mś��,�4�����9�"0rׅS�H�����lb�C�n� V��D)�<��'iJ�$%��Gb��;@Fٺ/(���Ћ��Ԣ��?q��?��Ş��Dצ�%�U8	d-I��kz�Yg��D6X��'w�7(����D�O��k��ߎ)��pY���;uإ�g��O���?&�&6� ?����xa��>uH��6}�-Rs}�����A1��$Γ���Oh���O����OT�D�|��I�?y۰9�"֭�2��IЖ����۠�"�'P���'7=�D��Sa�� 8�(Ӄ�:�hI�D�O��3��_3D)h6�g�\� �N#���Wg��D}��(�Ni�<R���~pr�I��_y�O�BN�<g�qH�'�-�q	F`��2��'Q2�'/�	��M�쒖�?i���?IS���#mT�b��,+���Z�H@!��'�:��?����=�T��ƤS�c,��I�iT�q�';���Q�O��ps����ƟXs��'��i�5�հX���������\$�r�'���'���'��>�I�1�L�'iH�%t�C�ń6$����	��MK����ݦ9�?�;���X5 Ry3d��-���̓�?����?Y����M�O����� ��'�M�m�<܊�\�g�$����':-ܒO.��|"���?i��?���{�LX���=P`Zc�CD��.O��lڤAF�������I@�s��UmP��U┿�p���Պ���O|�d'���Ů�8��	�dV����d 8HB���#��	5�@4���'2�&� �'�¼!�(�5vf�T��'�z�xz�'���'%"���D]����4UA��K�z���@"�߳4���S%�i�r��՛����p}R�'R�'�8m�e�.z8A`gӰ'�v=��N�x �撟���M��N����I��ؐH׮	�lXp!�.��0�`>O��$�Ob���OH�$�O��?E���P�Xi�hG��9�r�`�i�ty��'r�6mA�h���M�K>�DMB�N#�`��h�DZ��L�NՉ'P:7m�Φ�S�y7��lC~҉��� �@�HM%fbB�h��2t�D-b���?�&$��<ͧ�?Q��?�c˸V�txt���:h"4��?�����$Yߦ�FA\Wyr�'���*naz�Ye %)�
���n��h�	ܟ�*�OLAoڊ�M���xʟ���D;b�40��C�Q��+�L�O��1�!S�D���|�S��O!�H>��4Rr˅D�=4����fÁ�?�Ʀ��	Ɵ\�)�SNy�`�RPX��ǚf�8��`�S}����.�+���M�"b�>���$�.�8d*�>b�����48�	J��?Y�K���Mk�O�:B���O~������$�4X�����K�'�����8��̟��I���O���G�,p(�өF�>B�=�0��(,�6�)Kz��O���7�9O^mnz�mf*�
l���"��lT�q A*�����I\�)�S3'}t�m��<1�Ɍ�
Z���`�ͤ_M 	���<���
���Ip�	My�O�rc6Vފ �2�����J�r�'��'��im9�4�?��B��KE�T0��B,H�nd�mʉ��'����?1����D bx��OQ�U��77Z� �'�����^�&�酳�~��'F`#֪9���xU%ܧW�4+��'���'s�'!�>�	�v�N0���.��|`3��.K�X��	�M��\~�Nӂ�杕'F��dS0/H�h��g�L�*�	˟�I䟌�R����E�'��a�s
�z�� .^� L��iY+v�@ի3�D�����4�����Oj�D�O����5Nn2e3F�Id�L�5.�$W�� O�櫗>q��I�$%?M��5��t"�F�Hd5�(�,e��{�O>EnZ��M���x���Ұ@- (B$-��\�ש�pK�)	��!5��ɦr�7c�O�YL>A+O�8��#;x"��5�ۛC�(` �'��6-N����<8q޽��a�fzMq�f�;-�������?�^�t��ԟ�I*S8B��$�Y'-	�x���
 @��Ȇ�Mۦ��'(�h(׋��?�pV����w��!��DN@$�B��AN�
�'�r�'r�')��'c�0�{w�T�;`x2�˃J����OL���O*�l�C�@a�'|7M"�D	�R���r�	+�B)�uOW�p��4&����ޟ�ӭ)
 �o�x~��Q�L�,C$ß�����"�3u��4��s?�M>�*Ob�d�O���O��쏙c"%�$�@
b�� ��O\���<aB�i ��a�'���'	��:D��:�'ٿ;�8=�4&�g��Y`�	�,��j�)��@)&���3��8'�Tت��Z�o8���'�<�M��O�)ӟ�~�|2@t2�Q⥖'>��0���Q�j;R�'f��''��$\�8!ߴS����GE��h$ !��CA�-���zu�O.��d�ʦ}�?��S��1ڴP��y�e*Ƞ=;���-�	�9	S�i�N7mF1Tq06�*?�u*Ѡ28����	��Č7
���!Y�<���� `���BƝ�k�fmr�IFP0aǯ�7P��[7��+M�L@5�|�B`���2Kè�$��c܌�t �/�!��)���1׬�%G��I���7�
Ԛ�	y�B)��-��c|��)F���pqV��/S�Z���+�Zt�0��4���y�b�6(���i n�.Gn�(p��1�c�oN�̞X�����9Q`�<<վ4��m� [FDQh�˙�p���AO�;�F�B3��*&f!�F�׽`��f�'lB�'�����>I+O��V&C��LZ���$,/�M�ԯ�����c�Z���O]�%��%~^�
���n�x��W�Gg�7��O����O�m���U}}�^���	c?qA�X-"������0�(����y�J�!�H>9���?��b� �Wf�Z�����ڤ ;ά꥽i�Rn�	B�����O�OklȆ$��%�4Ӿι�E�Z�E��	�O7��$���	����ny��H�l��Z�I�@�I#7�� %����>�/OH�d#�D�OJ���g�,X;a��}h}����WO� T��O����O�˓V��9��<��Q�G"6�q��R)9�*��6�i���ӟD%����ӟ�٣nv?9R(�,g.n�rR�"FPpZ���j}r�'���'���L��1�����,4��T�����*�DK��%m��n��ؖ'���'�Y�C*�>��'��Ah����J#_��]ۀG����Iڟ̖'B�$�*�~����?���4�����K2����E�R�V�"�x"�'�b
*'�r�|rП�aʚ�^Z�<�pe�WH�8ⴿi0�I�Y RTXڴ�?���?I��nH�i�2 �Thm�4�:�0;�l~�f�$�O��!���O��O��>y9 i� 3lX����P)����h��|�r�릉�I˟��	�?A`�OPʓP;�x���!s����U*VX�u�A�i�9��'5�'a��$K'rJ8&�:EC��*) B�n���������r� D:��ļ<1��~ҁ�n�f��!M`��@����'��4��|R�'���'�����F�oA&j2�'|�~�p��l���$�nL���'��	䟠%��؋7.aB6/ˉttų�b��~��	'(����Iiyr�'���'��ɹ9���qrg�rVD�̅�,<:�P�/N���$�<�����?��鶴��DR�v��K�AuK~�;U@����?Y���?a/O��hT��|ʢ!+"��<*�.�l��!�3��d}r�'�2^� �O��ʟ�`�Ɛ.��+1��5҄u�v�ș���O(���O�ʓ4_�����B&[�0)Ǎ�G� ,��fZ�`�*6M�O��O|��|����3� ���E��~%��"���d�"���i��\� ���Z�O>2�'��\c���3� �8F����G"bB��&���	by� S��O��K�H;F���ӀO��FM	#p8������A��@�������?]��ulV�D>�9�&��;��Q����M#����dc��P�B��q=�i�� ̇*Ɍi+��ix2�I��'&��'`��O��)J�&DO�9��bչ`� 4�c&��փH(�Q��y��I�FRPAQgGR�VP&	���l�䟄�'蠤1�^����	Ib��s���(A�����R4�|k�y�BƓ":�c?a��_?�VX=�)T��"��̸����I��x�'n��'��'���X�oM��)����$Cz���>��
�����'�B�'I"T�\�\S�;rmކm4��ӖB+n�4��.��O����O���?��eM��G�%\;�pBb�:�F%��"	�?�L>���?�,O2����|��aS��V���,��"E:1��j�A}��'�|�Z� ����ɟ�j���M�cD�' +j��`*�2����O���O��'�L��3��TaS��1���=dv�a�3��W�7m�O~�O�˓Ƕ�����S,\a����W�j��uI �2Sw7��O��$�<�oP�D��O!b��5��z�"$
ԭɂ+�4$`"�P��M�(O��OL��F�OD������ ,�T׿<F� 2D_�h�l=�&�i��I�l�����4�?���?��'j��i�	 �,�� NR@HtkZ3!y<�1�	gӜ���O�5�#0O,��O�B���v�VHBL�U�P@�W��V'�V��Iu�7m�O����Oj��p}�_�Pk��/V�±1�F?p���	X��MKG���<�����7�៨b�g����{Q��Z� 2&�Ѳ�M;���?�� \�0��Q��'!�O]:uO�0V��oS�/@ q�i��Z����m���?!��?1uς?j����Ň-|�T��t,���'3(��0j�>/O���<	��S�h}��Ż��O�I8����K}"����y��'r"�'���'���]h\�����D; ߞ1�� �p����$�<	�����O���O�;7�ʳtG���nA�&�֭�A��?f	���O�$�O��D�O�ʓ����?��8P�F��H�f�;���H�d� ��i��ٟ�'��'gR���yB�d^r��po\`J l� ����?���?q-O�(Y�PK�d�'_r�j��V=�6��� �3L�j%�~��D�<i���?Y��y�����i�B���^�O��i"E+�xa�pB޴�?)���򤀔L 0��O�"�'��fT+�n�k�bN(l���j�i�y��?����?�G�T��<��O��y;	�	�^4���\�,��I[ٴ�� �rhmZ�\��ɟP�S�����VA��Գ
|�je�΍ LXP�i��'ײ���?���?q����&XL�T�_H��z@�	�M�JJW����'��'��dE�>�-OF� A�8i�Ω�C�M� �;jǦ=* {���I���I\�'�?93�-j�@���H%]�{EgA41.��'�2�'o�����>�,O�$��(��1q*���/I�˦}��bӸ�O0)��;O���8�	d+�¥2� +��R�i ���M�����uZ��'i�Z���i�m��ڑ1��6`�y*f5����>�5H��<q���?I��?!����N�n`�অ�L(*�q�"
�n����V}�Y���	wy��'Pb�'Р P磅]�BEB�,0nQ�t��yr�'���'���'��I�JM>=1�O]��Kڜ�$����D��X8 ۴����O��?����?�'�[�<�&�L V{B}pSd��U�+�mY&H��ڟ`��֟̔'t��5d!��Oۖ��C�]	`�:�S ˝"'�m���'������3�ǟ��OxIK���e����.K.�9��i_2�'��	0֦��O|���ʀ���cBB��͍_غM��Li�'��'6:칛'��'���U3���/NS6�q[�dF�U�vV�LK��[��MPU?]���?�`�O>q��hF�( ��3π�`�i6���ud(��OU� `��`��r�%��^>b\ܴ8{ؘ+%�i�2�'S�O]bO�� /xyZg�ҘY�R�r�E*l>@(m�T��IK�Io���?���ոp��,9ql��B�T阵�6)B���'&�'�(=ʦ*(��O��d������הW턹��M���(��e&���7�:p%���Iޟ$��*_<|��ُD3l�@�>m��۴�?9FGʭ=c�OL�D�<1��+ KM�^�[��W�i��U�^}�B��~��V�x�	ǟ$��[y�=TGzA s�Y�
�^Y�5j��qJ&XJ��7��ʟ�&����ʟ��f��MS��U�F)R����C(7lD$���������Lyr��H擝Mˌ�i��R?���C ��(7�O��$"��O����Aj�$��.B@LR�)�2xU Zf _yy:��'���'��Y��q�ʸ�ħ��x��"I67�i�폶fv��ɷ�iv�|��'w�N�6>�>qA�ՠ 4�h��Z=
�$�RF�˦!��ߟ\�'�@#e0�i�O^�������K�]2�gJ6qx���d�Ox����O|��<�O��Ѣvn_+���P6��{���iٴ��$W�V���o������O����}~�Y��~� �ʂ
V6�Z�Nߡ����O^x�G!�O`�O��� $�a�!?m}��pI���j���iv����oӮ�D�O��$����%��.��Q���,"^���F�ox���42�P�!���S�O��o���a#�TZ��yVn	�C��7��O��OZ+s(�<q(���$��t{��F�\����6L2`�"Y@G����'�j!�H9��O���O2�p&DC=4�*�)��O1�@Z3���y�I?��2N<ͧ�?�����I#?�t�1៿7`��)�T+r�O�BD�<	��?���?Q�4�
��"�=P�-�E!s�2�+T�_<����O����O �O����O��"4�ǄI�|T
� 
�t=s�§��cӒ���	Ο���Oy���l�8�'~`�	�M�2�!��>NQ4��?-�M�J>���?���Co}f�%Wεa6�S�/z1���!����O�$�O˓n�"tj��d�@� �r7��3(=X1�Rd	"V�6�O��O��$�O�Y`���T��)*�l�t�a�&��(R���'B�Iß(i���A���'"�O�wD_%d �U� /�R̪��Qk+�$�O����o�pPs�T?5� )�i�H93t&C#q�Д-bL�Y���n\��M�T?y���?�B�O(�Y��<��e�2�V
U^�(���ij��'����d*��?���5�;<�y�*	8\6M7K��mZ֟��I���"���?`�R�y���s2�@�pR|C�B̭I�����O��?i���X)�yx%���
����@%\�`ߴ�?���?a���+���|j��~��0�r̓B@I�+֝�g�Ă>?tb���� =�ħ�?����?9&;Ue|dAU"U):Q�ᄆf���'ZtC$F�>9�W>�$�O~�'�>��6�F�Hb�۠	�?$n�@�O�Tآ��O���O��$�O
Xٰ#Z9,0H�6a��A5��X���(q;�˓����O��O����OܬYclRg$���
�8U�	Kc��$V���q�>�E�ʧtՠm ��JC`c?y�B��&{F9��@�!�,Պ/D�Pt�-_�dx��䓕I!�|A�A)�I9����Ā ~�b�#�-����	,P4XҀ��x�n5���:N��0�c#
�!�D�)'nT�?&��C$��Zzи��
�L���Z ��$r���$���Ph�H[y6ڽp�H�i��a��Y0B��H7"�8���1�O�F�x���P�ITX-Y�N܅]��rc��*�$K�k���CO�}��� �U6w�����O�a� :`��rf��*�}��|z-���`p"�;z|H�K��ޫR.�3�>Ae&�'`��e.�(`��H��[���DğTe6��b�pp�<����I䟸G���'���
 aD�3�nI� lIHr�M�<9��\D�QZ�o�YELe���H�ٍ��#c �(s�@�V�� � d�9l�ڟ8�	�,����	; ��Iß�����] I�>���"��h#q��<,Ƚ��L
	��	,4݀C �3�䍉1MX�$���G�L�  Z�pM�'T�,���m�g�!M9�9�/���ɪĩ�d�&��	o~"�S;�?�'�hO�!hӈB:ge64��F�$��Y�"O^�����|�.$H�+ˉY��E������4���d�<���oI��^,��.ëK�,0�ဏ�?Y���?9��n��.�O���y>qʃCH}/8��&Ӭ.�d�+b�Q�/�V����
;$�u�a��`x��ط'ߤs(R�@%�	��xKqN�+��%B��D|����B�����DQ��S���&%��T�� 5C�p(1@׮MǴ���Oh�=��b��2#N�p�. 1�T�GG ��0>�H>9r��.��衡^�dʠL
0@Rc�5��'^剱`!~ȫ������7h���k�Fl�������0�����Oi	a �Op��w>� �'`��e!��䢭n��A�(�������%�T����d�31}vlC�N���*i'�~��]��N���&
���+^��r�'�@*��;l���>qB�5���U�;�D��� x��?1ϓ_��â���d���R2"|�� 蛶
���ց9�-�*N)�Q�n���y�\�h���_��MS���?!/�⸙V��O$L�$j�.R��
���F�R���O���_<"u��L!��|�'��-yT���VM@���+�![d�QI��9a�z��Pӂ�,�=���i?_*�-�S�=ZTX%�b��2{�d�	���4�?I���NH+B
�x�"�-v�)2�AӘ'~2�'K�hP��G	p80��Q-V ���y��|RcӴel�v�I<,�� �,��:��C��qN��[�4�?����?	w�`بU���?����?ͻ?�L���A8as�X+W(ϰN�����H��?H�	5��i���/�3��G+Z����ܔ{��/8Q�<�cSF�Ty�O�Z��	�}&��DH)*� �R.I�;�(�QLI̟��'t�Q��S�������h��,�/y@�G��g���çQh<A�N_�}�)x��
4�2��!�@~�"��|J���Ć�Pe>ѳg�]94��4. 1k��W� V��d�O:�$�O:կ;�?	�����H�	'��I�Cbґ_�dD�Q*%��S�K[� K�N���0=�W�ͲsS��#�Y���j�({� p;'aL#�Zq����0/��,��iΫss"�<w'"� �1I���0C�(�$�6W9n�aF�O���$�!N4�An��\�`����ĽOSa|�|��M u���袌�'@��hZԧ��Ϙ'T7�/�D��=��n�ޟ��	�VY^aX�"]�u4q�W�O�E>Q�	D�!Lԟ@�	�|B�$s�D%���Tqr.�0$�� ����j$OBM8ߴVpv�Q� ��gW��Rl�b�d�P�~�@�� <��x�Ò-�?�����D��#|�8;�k�F�,��Q �{	��O��$3�)§l��se�N �耪�`G�R^4���~�����V�ڥ�s�xgI9�yB�)�UU�P�Q�Ժ�F]�3�P6Ypl�ȓ;,>�pK�o��2�(�*�楅ȓ4������~���&�_.	|9��z{$1�G�Tu:Yb��:t�^����V�.���a�%�o��ʠ"O2M�ա�w�"��G�dN9�5"O�l����<B$t�[��4\�4
p"O*�3��	e1���' �oT��*�"O�1��+ɣY8������	J��H"O�y��h��LCIM�xz4�R�<q�*5�[�-Q�`sf�ق�M�<��<ћjP'	!\ 	E�OL�<9�垬/~�<sAk�"3���`�EH�<Vҟ0e�-���B�}���U��B�<�1D�3(��a#�p��Pq�t�<y��X 9�m��ōe#��[E�m�<��O
��"T��a�H�@�<q�W0J���Ë-qj	�*�|�<aBM������	m�����t�<�����bf
M)dFAW2M���p�<�R-�.Œd���V41��l�dBX�<)�{���F��0�@Ws�C䉓c|h��HO�1?�\+Bd�vC�	��LВܥ}4��p�g	'��B䉺$-L4s��[�A��X;b.�9UlB䉤�2L�qc��t�p���n�|�@B�	(��t��_�P_b=���;E��B�ɿ;�v�J��
4��W�C*t���L�O)�\����&X5.�>%��=r1��:$$�aJ0$��k�.(j���32�Juf )����M\��I��3�|lA��mpȣD���9;�B�	%f���#
�+��R�.��bP`�I�|�ѻ��Ek��s�4ӗ��+H�W�ޙ{� ѓ�	"D��1CR"Y�f�t6����0�a�$�!f֯ 7�cW�[:L��x"�«+�]�� _8ȢX�R�p=��
�h�y�����K/>��uH�`�S���h�j�'�����/^�3�O0d1,-f˓�m�1O,,bÃ�-v�����E�qs�A��dD�3x�J2��(oB��T�R+�yB�Q+s�@�zG��u�l�:c	G6n�0SĉW���Y��v�,����3?���$?����V���&�T���e�L�<Y�E�Z����&�!��[�˒�e��8��@�;)�P�u�;\OЉ�#ʇ�9z����N�|�vUy��'���i#��&;��ۄF�?QZ I'�#(6��3dW�v=���'�
���o�'dn��Gϣ?�Ь�y�O߃ЭS���=}xD�Dn�1S�ؚÆߟ�|��L��yRO�,�"���9}9P�Ѓ�I���0� Bؙ�\�ʼF��O�p�-�Q�Ҍ����O\�e	�"O,��!=O���˖(R�A�H��f	Ѳ���񐥏�,	"�ד0���#kH�S+`���E�(�1��ɉU��H�&�O�Oq�3�H�
fN=��NV�H`�݀P�>R�C�IX�n��HM�0�nL3p(�� a|c�L1t Ц`�|����F� Q>�B���/Ȉ�� G!zɂ!���3D�(㵠�Kw����,�1*��ɸ/��
�p/Ȝ��D֕8�>�'�Eh�,Ϯ+�\����#dt<��8R��$�]���y"��&ܾ!+������ ��!�*K*gr@�F՝;In��2�'��y��޽d�F�1о(�Rg�$%:4)yw�[�k����ȓ)��H�B�[^��gf=��u�<cn2}@�t�v�.�b�U�p\���QH�+�6`�ȓ~�e�2L��|��=g+؊(�A��H6lC��'�64���,B�'�0�h5q 5s*h�a� D���p��+`ЀKga�`��L���]*K7�����4�1O�иX��' ��p���%�ӫ�7m����)7��Qe��v����4�>q{V�=�¡Kğ�\��I�3d�J�&�d�b��#K��
"e���<�<	&m	�P;�=c��=����!��f��l֨�9�>8�CKð(m���?7�I# �]�G<A��Q4��wK�B��f��XSf�2���x�;]'Hi���aX���⬒�`�]�ȓH^�X�`�K��xxC'����P�Ů������>�ɬ��л��g������ț$
���[�0=	C��R��e�ե�|;�FHZ$D��9ض�J%2�L#���'��d�.�,��	�;���v(_6sAȼ� �D��b����-l�ѹW���-��ȍ����:q�2�G=)�� B���D�PB"O��h׊ԕ��X�P�L�PdR���6-H\���$�*�(�� �ay�c��o�@	2��e� C�	�O�aB$�'E�ѲO2l'���:f�2|P �Kq�z��$�L=:�i�6�xu��9�Ms˓aZA�uhĥCg��;������4��(p�D��<︱�E�
�����4��0;b>-j5B	�h#J�	w�M9g�i��4�IT�h� �Ă��Q�2���0����~���Y�6�H�i���>n�
!�N�<i��ľV���n^�����*�5(DÝ�s$x�G�<.gn����H���x8C�ǐ>�N��6�'8���	2W�t��B�0S��� ED�q�D q�O���C��h���a"�?#<��I><�>����&|*}�	�ʟ��僿��i�į§/@���A6�|� �$J�U�V�\�r ��$OQ�8�H��Ju�'��+�ݐr��w�p�1uo �:�l0ZU�Z<+�N�0�kFN�2�8i�	��i�pwh��P��\GF�;�yR� ��F�9����� s��;Ϙ'�l�JG
P�	°��̕%b]
݂��D��iH 4�R8����@�[�0�J�n�4��� U���Պb�!8�u�B��P(EM�hVaz2ɴ�b���@7��C$_��yb FY�z}p+�d��+2ٔֈO��3�۾0����sfH;S<��kG"O���V/¶�`NS����J��J)/u"mEi!ړE<��P!14��̻d�:�I��V�]��.����Db"��{��	Ij%!��\�&Bx��T#�;?�:���J��U7*b����B���KK3a<Fy��Í�1OEIE*�9m���"� ٓ$N�����OLijdJ�&�ʓh)HD0����%y���V�ɑ~�������o����C ?~�냧��|����n�)����䔂6�p K'�f,z��2S��#9�h9�1oɓ^����tBQ$K�ў��!���I��Lc�����BҦ"�O,�CТ��?�i���2Z�L�p�gW�^@�Mk�DQ�V�()�Ŕn�':�����!S�0SP�
� I9��A�f���Q@�1L�9ӎ�Ĕ#M��I8��I�F�J�PD�O�8Ѣ��S���R��уŴm�t�����yr��5D����BOE�<�TD�6��'�P�F�x��}J�ǔ%�4��� u)��e�Է$��LX�M�O�R�N�/8V�|H�״e4���aӪ�:�ӒQ�ڍxi��<�ܥ� �Z�#!>,��ͨvy���'��B)���Ƶ���O0-H�`Q�=!Բ�7cD+)�|Єh>v���F%+ғ?|	�Y�X01�dW�>"d<�q�+�Oj�#癞���'(?�B�����0(@,�[�I��2��$�hMEzZwЀY���Y�>d�%�Y�������L�.8���B�4=��PI��O�>a�=c�;S�p]q��պ��W��J�%�l�Th�<i�T�ʐ�d�)jT�Ȕ�@�T�� �(ؖ1O��:GMƱ(hui��Vp��0F�S�����r�v��b.c��YG2�D�Ņ}�2Y�A��(}0�6!>�.4�� ���O9�(��,.�aY�k��ׯ,LO�I�"e��M�����B�P�$AѰ����!�X�0tˑ��H�ִ��M��HO��""l�;$�ܤ������( i@�'Bf�A��]*+�ɧ��'L�ܪC@V��1PT�!v�f��V��r�N��#��=Z%aab����#=�;�k 2�иC��#c�x�AqL�
r~V�9�B�*a�D$��R���>��O4��aak�clt��;Ox�Cu��X?��8�H�%x���憌+U�1O��⎜z񫌮C
�X�C�'n��,P����ͨEcr:W۫$κ���+?�Z�[6"߱S%0�K��'$���݈�r8SˋdN�� ٴz0���ɞd׀�C�F�*����	����Kr�!}l5��b�q����<|<��7B�#T�D�I�HQ�:z��ٴz��Mq�!Q��ְ>������64X����}��� )rH~h�#y(�'$� ���t�ɧ��{Q�����U�R[��S=L�xQ2B�N$R��1��	�=<(#v/I�? N����E(��p�N�4s�XZ�;O\eℚ|�ㄺ_��)G��H2�i���~r%I�|;4��7���[��HO
t���[�]ZH�����?��U��c ��2⤈$"@q���O��"G)^�x�� @� �O��!���,v��	#\��@v���jjb-���̦�x���P&ȝ�ڴ%7��Ћ�S��������?!s����nP+��IO����aAY�]IP�}�t�d�W��*�'E�P)��Y&����d�10�e1�#�1b^�=�g�֜u.����^���N��FK6�~���5�q�w�� !����[�t�V��l՜�@�Rh��wX�Hk��	t�'ΠTq�
��v�HD�!(��D�@ѵ�X�6�X%�p��>)����ʕ�F*Ȧ="��KKB��i�^��DKA,�@�����7 ���j�Ɂ�#�Dz��� �ls���$�`����~:�+��'��xr҄�S%���B	�:�zƦ�g��(3Q��<U#�7MF W�Ȕ�H>�q�O�T�D�H� .�آ��1r$�\��4����¬mz�!C*�(CTG}�fR�&��Ezk��hf/�+bpJ����	'�`��".���#��?��D�9ph��"
K�6n,��S�֬O��ۇ��<��{2E�ve󩒍�b��[�j&���-�TA�4$ ��DF'R���T?a*]_�T9����G�XйT*�pc(���	e̓tk8�A��a�����+zJdCf%v �<�p�'5
�Y���*�1B�^,l.��{�/4E�U@ݚX5n�bQa�1Jvb`�t���[���A���9�I�-�����r� 7m �e��p�dۈd�h0�0d	 VNў�XAƜ�7-�Y�ec�V���3f@�l�x�*���vPi�K'��ZE^���=��_��5�v�J��k��_J�-���M���>)���/X5� G�-~�FXd�F�B���i؞���@�W,0aAG� a)����~`����'7,�����>:n|hČ=iJ��U��'�|��j��<�XD}��T��LrF�Їk)��ׅ�!�?a�W�i#�4���D�N�9�i�^�W`^T�#7O��
� ޯ&�(8I?�Sb��>zN黐�w���ڴ&����wBϥl��Aeǆua�+��8�}/�tڶCG#_��3TGǈ[L��O�![c���Q7�	���[v�j@���Cup�A����^�\����8&Z@:P>4(m����p!B��`Λ>xۖ�+�)^�E.�*��Of�聳e	�b�:T�2ړ�y�$Յ&���xE'��Q�bw���Px��R�>�8U�6�\+op̸���
�C���ER�ˬ3-��3��Rk��p������pJX�9�jq�ƫ�U��@H��'B���P�]4�ȱR:7K^i:q N:8��S�Dϗ���!�ݕ��D3}��HG ��6����F�:qQ�`(�E]��^�ar,O�#�R� Ł??A��H�,�4��E�Le��)���k�'L�P�@E�J�����$HCV-*�Q�T5����j8�H�/X�+�0ڰƃL?�� '+��z�Ժ��M�`��$~��G���a��D�@=D �Ŭ;��׷\�T\
"G�>��U �χ��D�?Qu!�<]��iS	�_>j9�%Օ@�~��� c�q�I���%O^�IPE1X�����D�,E��-�.�?	5���n�4	6��CS��剚q(�%�p�,����GR�9���<w� 2TX���]V���P�a�I��U�z,2H㥊ӊS`nB�B+R�OtAQ�m�/a=��4�F|!PfA4]���+	��p>��ק#�{���PVl!,�`�z|�5
ϛG��y�h�&QBB�FzZ�yg��th)3�DיQ+2諀-ֹ�y�ΤL�j���Cԡ}�5!�W��M����j���Kā=i�4)�"�yg�A�'�8�eL��F����&	\)�y��R�u�ճ6R/(!|�N���y�ǝ�p��pQ��'ְ�e���y�n7;�-���6Sq��و�y2E_=����C�9� �J5Ξ8�yb�X!^(��#�ۏD�zQ��b���yR%A.e
�zV�M��d��L��yb��..�f��
��t�����y"���g��!O�5>ݘ�`���y�O���v�T.,.D���i��y��W�4d.0�mS�,�dPW��y�t�BqB�'ءmH�`��î�y"�H
IR�"M۳tK&)��y2���2E��]�l�$�i���=�yR�ޓxEi2a�Tar��A��y�^5�0A���� ��T�T��y��1xz��]�t|B�z�U9�y���,�>͋��l6�4	��3�y�픮aϠP�̪H��p�L!�y�.'t
�1y�l��9�ҝi�c���y¡}"�m�*�2�6Y�c�F��y
� 
	ĀB�`A�M���#^4�c3"O���0��k)�XV��'����Q"O4h�&P�XI �PC�-�p��T"O�� �Y�0m �b�vdi�"O�\��d��$x�(��
��qj��S"O�Dk4B�
 �M���V�pc�"O��; ��p
�(���|V\E�"O��qgm�: ���@�ZIH�aG"O�m�B�۳|�����Q��"O2����v4.���]�O<p,��"O�����j�čB�F�fC�Z�"O��.\�h%�F�8�l8`"OI{���%0���:��ڟ>�h�i�"O�qqPa��jb�9�䞰&�r!s�"OXuAa�ѴY�`�&ɠ��8�s"O��(a�"q��5�4��;b�~��v"O�jc#\�y�X�ŮP��"O*4���ەETL�	$�4h��{6"O(1Y7��z�V�2�]�M�Ī�"O����e]�V��i�[�JF�UZ�"O:�rS'��;渄)"I�m�>,00"O8t����p����`�|z�eD"Ol�
P��
�����m�>��3"O�
�,���{f�L9(�P#!"OtM�ԢY-Tx=)F R�)P�"O����P�n�&��,�٪ "O��������[�/\		eN ��"O�jB�ҷ'�-[��9eZ�dX"O��04��.�����';F>$u`"O*SE�(S���Q�"+3J��E"Ox,1���F�bLs�!��c"ORE�S X2s���'!�,fF��D"OL�(��g��xBPn��3e`1�#"O��ע��W`:�N�$qq-c "O�}k񈊻R��1�&M�$s��[�"O� y Cg�kVe�A_�&"O�d�f�%krD�a�
�S!j0��"O����!8z����Qju�"O��c#�DNN�P�R(ti�d�"O��#K��N|����sd:���"O4|9�bG	�D�A�0_AB�"O\y���K�dh�[�JJ#i����"O�}�����iC�}���[	��}�"O�ᐤF�J�ڌ��GC�m�0p�"O�pkڝa���ڃI�Uj8K&"O P�EC1��	d�FeB�!A�"O&��kA X�L�e��v-�=�"O�1���pL���D jKҹ�"O�+^1)/¨3B�X"q/~u��"O6�:䄈�(�rՋv�ʨ(�Qkv"Od@P�E�o��pc ��%o"�)��"OL$9V�_=@��P� !��=x "O��	��U+[��( ֦\�����"O"T���K�05p�A��!p��R"O��(P-I��`Q ��+HH�9�"O�4�0�U ����6`�g:�9t"O8�rGdʮ\VrK�푈#����"O�� �n�/A猜{�m̄{����'x�z���C`T��R����H�'u~:K�!��D�6qQ��# ��yB�S�U�6�P���EpI�����yrK��B(@G�ٝK^u��ć��y�&�^[������!=".��6� ��y
X�Icƅ�F��=68�!!���$�y
� DZ�d��0�~�QY�e`e3"O���O��R~ m��'�O;Je�#"O>��7ńG�0�b�D~)�y+�"O���2ˊA��M��j�2��"O�E#aHQ;w<q
��m��4i�"O	I�e�9��Q�a*�<��q��"O��B�6k'��xWI���t�""O�h�EM�8WkR�)&�܆��c"O�1	��Ǐ|p$�$��/e*D"O�;��M��4�8R��I�"OjX���	%�<h�bpEd��"O�%P�h؋Y���Q%!L7/��'�'�:� �`�4��o\6E8��'�ք��bHr�0�zteZ-x{@ �	�'�P��r�1_j�2���%�݃�'&έ:� (}4�"t��	���
�'?H3c�B�I"����*FI����'��Ј��J6�����"v`���'<�h���;k�9 R�r�x�
�'m$P������V�)Q�-s��E]�<Q��I�S���0��I�=P��Xtk�\�<a��ynxl�'z}�c��m�<� P+'.�[0AK?\�b�r���t�<QC�Ƴb�P���M8!-��CCEK�<��l�/_F�$���&X�5���W{�<9�剗��J�ʘ�_��5��t�<���6����>>�|("�s�<�g�$�~(�A��?Z�zPOF�<�2�ݒ]8!j5�C:����TE�<����3�"�i׍@'Ad�1���U�<�U�! 6��`��`� a�XY�<�@��S�R�+��Ĺ%�����i�<�rG����A���=_�$�
�<Q��� �na�ъ���ȳ�s�<y�R<� �c$_�2pA�_f�<���//�5�sFP�)䘜# KPG�<�RP���E�&B/.��=�&�j�<�4�V�v���#@�D.	�z�"2�i�<��ʂ7M
$�d�n �m
Θp�<���^� �ڭ�c*t� R��B�<i �A�p�`�S�),q�(�@�<1�$�0��(Z������!F�S}�<�%�ʝ	 >hb�ƍ
l!��z֢�w�<�E�#E����.C=��dRE�Ji�<Q%��:8s ��Q�75m<t�oe�<Q�m�/8	�<�Ѵ=��L���g�<ђ ч$��� ��LD���k�<��@�7�>�h�G��3S�`�g��O�<��NNIl���ہs��h�ʂI�<Q�Q�K������>���#��E�<�emX�nX��t�;	Tܙq���<���{*�<�Ў]�YZ4�PE�P�<� @�rCfQ����Llj�zbFAO�<a�/��j�k�2=�j0◇�f�<YĦT)2T�z P!G�|*���}�<�d#
!>0x�͊+���	7�C|�'R?m����7��[�n��}{jd��M;D�(�Gҏ lI�MLU|J�Ю9?y���+
2t��q�J\��0Fߋx֢=�ÓB&�l��j��o�t��ċ�अ�c�UBw���x�(gJ'm5����IR}�'&rvv�kT�I�a��AC%e��y�O����\�D'U�x$j�m
�y��T�'���+re��N��s"F��y
� 8t�q�7+�B4��SY�Y�&"O�l��#ָ}�d�Rq��uVv�X�"O|Y"G��g�0u�f�ǩ>�x�w"OJp�cҠf�]`bפg V��f"ORt@ƌ׺mI�������/�����"Ol=u��.�l���R7	���"O��@tA�bW��#�h��~<�a:�"O��KabD���D#��2'�4� "O �C!�,69�x1�I�5�8�5"O�x�/���N+����)�"O<�AQ-Y�Yh�դ0.�X�)&
O&6mQ�E[��"� T�.6L�f�ʄN�!��/�L<�f�&$IP�ȓFV%�!�đ=Wi����8D�l�$FM�A�!�d���P��7��C+��kTE�<|!��խ�༠`�$)��x��#��|!�DЋy�0c�`Q">|��"W&c!�dZ�D�J,��C	3
@�ԋ�
t9!�&;hH8���C?$#�m��JG<,�!�D��*�5-��knГ��&�!�$H!A�ddS�H˂"W�Ł6�V4%�!��Z{�p 8�Eô08��P�Fאd!�ȸ,�c�R7^��m��o�SF�	Z����I߀k(\�٢/�:V�WJ(��p<��D�8B�d}��&'��5�lJ�<�P�W�j����G�>$"��a�C�<�&�ʨppk� 2�v�Ɇ,H}�<�5�g~r1�i�X��CDw�<�ck�"U���2�@ J,��1J[s�<��C܅�\��k]�K.�����F�<)Ӄ����|{���
��&�}�<a��	�5�,���J�Z�b5 ��y�<�g��/Q�"�ȏ�zI�d�w�<�uk����X2*οo�^�%�)T�0�K�.z�b`���]t�!�l)D�(���U]$M�b]��B�z�&D���Cd�;�҈:3�-C��1�J#D�S���9�>����t�ʅc��&D���V�_�q�8���J�LTTc�7D�ೳ��-"�la�H��ab��y�!򄉎u�(����3�4X�aҁ�!�d�?3�E���lJ ��i��!�N x^Z "��A�vN�H��2m!򄀾o�T@ �-e�leR��U�!��iD��� �@�k����E��	M!�7^�f�"����<i2 "�z6!��Ձ&9FȡR�GQ�0U��!ʲ";!��O)"��-<܊�HqFF�w�!�D�"y~(Kg�Q�(zt��gŶ|P!�]$�Uy�I� �ᓭU% !�d�~)Z��E�=�6T��� J!�D�;M(�Z���u�.���k��!�� 
�܍`�̑0,�D��g*A�!�Dܠf]BD0��[�l��a7jP�!�dB�� hBE��P���çn���9E�d���GG��m���%,�6��ȓE�Z���f
��F�i���=y���id���S{^4X&�V�J1���W���+� �a�J��Tœ!)��͇��V�6' j�H�U��y?�l�ȓ7*�qC�I5z���2p�_�'�8��ȓ*�\����ͫ`y���M�oN69��r���k�O�*!B���Ɔʺ`�乆������#3м��6@kb���S�? �ݒV��/X��K�F�]�V"Od��R2%�,d��	�&��`R6"O��yT��J|��s��$p�4��"O��1��li�	+%�Թ+�>�A"O2�k�F@�5���1�%B?(�<*�"OH�����)"d��\� (��"Ox9�`� S�� �Їv���YV"O�	r''Q$c8�B#☪#�!�E"OR���
,�8��Aȴ�"O����Ą�	D|� ԏ*Y�B��s"Oh,�V��?J��Ah�e�hu��"O�H�����ӬR8�|Ũ�"O� �g@�^"J�
c�ݠW�Z �1"OT ( �=q� ر΋��f̳�"On��t���L�Xȁ���X��"O,�3��[6nz�M�U
¡b;��Z�"O��Z�I^46% ���ꄀ"9�0�"O�x`���>/�p@�S�?@ �"O���"�X�7�,#���[4Pr�"Oxm�a��ExN���3u����"O�`�Η+,�т5e͍�ݐ%"O�ˢ�/+Y�M�f�Z:j���@"O* �E��'Z��CO�݃!"O�yb-��RB� ��6"O��%5W�4 �K�c��)�"OL���-W	tD^<��;[���"O�}ٲ�J�h���pǂ�Ϝ%�"O֌��c��u�R1��&��d���
�"Op�#���Fc�Qb君���C"OVHb����j�LM����~��Q�p"O�|���Y 5A��P�"GJ�8�D"OZQr�B�?~����G��	����"OtT�EH�;o��Z�C�e�<�"O�}�R��5� �Ӕe�Ow\�5"O�����ϴz��4�Wc�� u`��U"OH��ŏ+zi2���ǚ'����"O �q$���nM���	1H����"OX�kaF=����.���a"O���"DQ�<S"o�N�,("O��p����1���Q5�
0,��Y
"Oڰ��/R�y��&/��*	��"O�91�8¨����&df,eKs"Ohx@��cp:�PAˋc`���%"O^eQ���"���
�b$�}K�"Oz�
c@�t.X���H|Z�P"O�0�$(9gx�� �_�8I�"O���ȹ{t� �QN��d��5"Oxe�S�X�tt)+矅.̖�J�"OܡCSGA؈��L�6�
�""Of�)��S�	.N`
�"RA�b "O�s�N N%��$�*0V|yT"Obxa�dX>+��PE����H�w"O���׌��Q����ëJ�C�v�Q"O��zG��f쐁b�U"jߌ��5"O�pC��^Z� �IϜ2���xB"O�B�m��%�xI�T(Ɨ��Q�"O���C@�0S���,�����"O6x��F&g8����#�V$)�"O @0���$YL�2�C�y�0H3�"OT�Pe�&y�A	��Qdw���"O,@�A�y��0�c��+v"O�-� ٕ}���3���;�� ��"On��TK	$%@��_,�д"O�L�WT�C�̑��.� r���"O� |���?(�!�3$�-S��j�"O�`*MZ$'V^�k�#�6Q�tY��'�����@en=#4�	�;#J��'�6����ɖx��e$�5�`{�'C�mS�Zg����/&�A�
�'@ �9����@b�B(z
�'<��2CCC)bL��L̚w(,��'|,��g޾Tc�a��*.�ؼ�'��)г��o�Bt�叫.פa�'��xCr��jr��D�Q"q��'����M�G+Z��vf�L��M��'������Cu���K{K<�b�'}��
0��d�<= T�� � ��'�tJ��*7�4��ά!��� �'����i{6�06�I��r��'��� �B�<�68�u�� ����' ;a��O֡z��#S����'`�-`�E<)/�KU��NR�,��'����mћJ"I���Ƴp�Z��
�'I|�;D�U�l�L���l�5�
�'XX�JR
�<8��%Q`h��MH
�'�Y�e�>=c��f�$�!�	�'\ZċP��+0��p3��
m&	�'sn���FĢ]V�j�k��g� �	�'Dn���*8��sO6jL=��'=j���� 
�4�
��h`���'����I�f�$�ƨ�\�<��'-�`�i��M��p�ٗ �V�H�'!!��n@u	 EA�a/���'n�вD������6Iݡ[��Ic�'�&p���ٜ3�����hɺ؁�'���o�#0�(`�d�)=0в�'���A#H�t��A���ژq�U�'pŏ�<䞸��H�j�fi�
�'��1��1�<��K�`��)
�'H���ə�.Nu��%W���2	�'��D+� ߝv�}��c�O�����'��D�1+�z]�$KdEF:�Y�'E�hZ��Q�:���f`í<�B���'�`�Xu-ћ1!��9a��7��(�'a�l*#f@p�hL"�h5���S�'Z��#`��k舍�0��/�$�(�'�lAñ� :lM���'�&d��'�a�k�L�Q��$�ٛ�'1hD���:׎ѩ�E;P�T��	�'>iI�S'� ���E���9�'�n�1�О?Qp���F8'�����'�h����0�D�e鉥w~�{�'��H��ǈ�{��iZ� ?k:p#�'P��X�i4oI�̻���_��`�'�`���B��3��%BQ��z�'ž9�fR�N��U�C��&4�<(��'������7T�C�\�+�v P�'�l�A�ϥ`E�"�Y�S�$b�'���H�#_�&v=�@��$I��;�'@�̱��D%i��;pfPPC�Q��'!��rű�xZ H��V�E�:$Q�'f��L�7�p�#�P�F'5K�'�8"�?V�$�` ��'Y���'y�i���Pne���ǅ���"%Y�'6D�0a�AF�� 1��`e���'OD�S'F��>ԆM�TFC6#~�Q�'@��0�)�&���i,�#�и@�'��D@e��b�I�T�݆ ��	��� �qsB�X�G!D)`�H�4�Uc@"O��j!�ْ;����0��h+*��6"O<E2��ț%oV�A�$^�]2�E �"Oƥ���L\�0�A`��*/Ĥ��"Oibueêapld�ٽ,4J�"O���1�,�HeN��"R��w"Ox��u�I�|���#�0��"O�P��@P<j��R�H� ��"Ol%	$(�.,L��� 4�H8'"O��p�*������i�7 �0��"O�`F��#\�Nl�R���K����"O��#��5o<rx���9@Ҙ�"O��q5i 8^����/�&�1�"O�;%�ߠ#�����j�RX""O Ԣ�k_ST�PdV9?�p�c@"O�$	�Fö]�Xp����>~0�2"OR]ӑbK�eV�jSdŇi����"OR	���d�|u��a�|V����"O$��e�ު8ڹ�bkB;F󨀉 "O$L9T�ԩY���Z<+;�)��"Oz��`��<'���⃉U���aV"O���f��&���#��;o�dg"O$䒧	��*��d��d�v��:w"O$�#NJ'=�TT���Ӧ9���pC"OXTBC醠8��R!O[�HY`58R"O�T�D�Ծ(j$Q�E�ӒB��(q"Ov��1�΄L�����[��@g"O�G	tL��&�O�3=( �"OU�aD�]fX��&鉌V��1C"O`$��>U�����N�&/m@"O.y��A��Ff��Ƀ)"�1(E"OT�+�fK�8h��)���?؀"O�1�O�M
jYp�W�4�vРp"O��J�/܊$��6h߆�~ �6$D�(�&�8l�̄#*�:O"� ��=D��!�C�.&�QaE�AT����	7D�����&��2�A)4МKg�0D�hT˛�a'V��01v�t0e-D��9��ƁX2AQ�끮u�v���&*D���uLU�2�I��F��m)D��آ�L�S���QŁ^9�4pc.*D��p%�v?�U�5��w�� �;D����m۹m\~��k�s
��[�>D�X(��#��A�Ӳk�z� ��2D����u(E��"r������+C�	�Q�$�s�@�h!<�Wדe�B�	>�ȉbf^ h�ؐ*�'�B��1c� �����7��03�e��[�<C��;��`�5GQ��� �I��(C�	i���IUZ����э��n�B䉏�"-*��S�9Z&��hB�hoB���ʴ&��"A�(,B��8 �,	��'!Y@�r��42W.B䉄eF���P˛�Q�xt�p�syB�əL@0������d3q"�Q;B����!��X��rp�&'̵}FB�I�xƹS3H�'1o@��!^I6�C�y�0���>0nn�a �g�C�	�D�b9��E��4����u�C�I2c���8�!��#V=�W,C80\C�I� X8�!a��+�b#�fV(6�xB�I��Ve���#b:\�U
�,c0dB䉍�uys��8N捙���670B�	=){ʉ)vA73�ˇ]�ZfB�)� ��@@,FaYv@�O"4C=�!"O�e@a�݆VHFAZ��B�5@N�5"O��9DK	/K�0*C;Xn�� "Ohl���!q��"�\31��� C"O2La����=�TI�b�5T�lD"�"O�`���@fQ	����H��
"O �a��0+Q ���Ϫ~2A.�yB	�8hКa���1��8`�[��y2��4
���	�;,W�����>Q��y2D�)<��ePeU-r~`)�� �y�%� �ꃅD;4lR���
�yh
�~D8a�Y�t�cҦ\�y�dY<{]���#����a�����y�˔�2t�P��L��u��q��yR�1:�%k�J��f0b8)ABƥ�y���P��Zc�F��
�"�� ��=�����ˏ3�$P�%˙	 a��P+�!��
VϚ	�0��yk��0���8v�O���dR�ZҮa�$�X�Jh~���S2?b!�$�nL�V#�6�:�"�O��DF!�$](cT()V�&\:���\D!�� u픸	pdY?5��!ю��!�$��4���+s�6Z@��C.]-c�!�d���8�#/��b��t�!��A��X9�MC���]���1�!�^�a��p�ҢA�x|ląȓt��w�ʉO�,��*�$gl~���2Q�z�N�1�A�w`�n��ȓ7�vA��*�5A�P��NB99���ȓ ��X{Vaہl�D=����/iv��˟x�'.M��ףMT�	��<T���'#�t9�K��p�^�h��{e&�
�'�0]�to��eILk#�I	�
�'AB�fe�x	� ΃G��P
�'��@�m�~��r��ٸ:C �b�'�(�qm�.~<�Kщ,w��q�'80xSF&�� �� ���ߓ��'�<ण�R�Y+z��(E��i�<A�m��N�!��AɿG�4��LGK�<�!�,s�&}�"tߢX�3��\���#�v)3&�G�<����
�;.
�A��Uz��B��?u�
&`�/l=C�I-hpQ�*@+z�z1ǘ
)��B䉚Y��B�n�3]���Ћք_Z�C�ɃK-v�QO�j�p���\�B�I�0A�Q�3�х!h8��#���B㉺]�4�Z&�L�.Ĵ;0��6w����'�a~�.�~t*|��D�+��y�
���y��J/3H��c�q�pەe�9�y�FR�d� -�Ҁ:-R��e�y���&��tI��;>�0Z0%��yR��Xa���@ٻt�T�$ȓ��y��	�@e�ϭn:t;4A[��yRɘaQR�!vy�r���	��?	�'�dJ�O��'�"�J�f�:4Nu{�'an���͐Z�6t DE�=+�2��'S,�P��3�9�[����3�' $�)u	;p�*!�c��*<N%#��$�<���)�V��'��f��AW�ߺ	�ў���J�O�Z�kue]��ҷ�G1kG�[���.O@�+���C���S�n�r��M�U�']!�dӴ:0�΍��l9�J
? ��w��yT��^h:�S��7#P��N<D����`C3��Y�I\�@Qjt D�� X�2�K�S�̨�挝�}���C��I�G�D욛�����-o�j-�T�����'�R�O�~IP"��qv�����8nT4��'�9{fOB%d�1�l[�cY�a��'��j�]�	�l:7��,Ԍ����x2�:��!��m�\TZ7�H��y&N*mI�6&�6Z���f�1�y"���-��X��2U�e���É�hO����N6(xz�����(`�PMݿu�!�x�hpZ�g� ;$��64��O���:�����}
DőF�Er�igO,\�Bi��ORp��t�E��)g�O`B�ɨI�^���%>JEt�yՏ�
 FB�I/�T���ؑUR ��P�A�"B�I;5��m�'b�(�(k�OY�l��C�IPL�!Y�l�0"Ǐ��Vt��鉲E�H X#�պU%8�)�'��pG{J?M3E��g�̹�mA�#�N�<4��I��͌j��,��'�5��jeK�w�<qU��/O|� c�	
M�B���Mu�<HI�8�l�A�n������q�<iV�_�uB(�a��34��-	��DA�<1�Gō�(���O�](�̠����<�`@ XTJqIVK�)-�8�ё��}�In���O���b�ײ�b�{w�U��t����'i>������xPg>-0�
�'@|��q���V�1=�*�{	�'��,�Ťa&��8�a
0)�q��'
=�!��2`�͵!��J�'�*���y�L[��
En��'�����X�y�LX+Ĩ3�ܘ��'��l�R#��[��e+"���$x��'� 8���m�>�fE�p �9���x�O2�~ؐBɅ�*��{q����y�ڢdp���C���$�Xeya�� �y��ӛB���R�[�#'l9�7,���xbaW�7c��w�F�,��m�*L��tx�l�'�Z��,9=�J-I���*X� H��'2�%)��ߥ5��́χ>G�MsM>i��?����	�k�╸�k"��d3�G8P��0?I�G��?��0a�bf�щ��c�<yV��y�p�0��R�J2�0��W�<��̓����6i�v`��	�k�<	���4�]C�
V/j�����'�g�<��B�'qL��G��"
v	K���?IK>���~�@��W^A�lƕ}U�q�R�J���͓@���h
=�����Q����C�I@����o
7!&���IE1$���bT�6D��x�+�n�i�#ą�Y��6D��fm��h���f났ni<�2D�2D�Ĉ ǃy���4�� `��.D��	�d�9��<�C&�B0V�)�	П���ӹL)�t#0�j�ĸW�-�f���O����y��M;�4�*��9��%�O&Ջ5`%��y0!ך>d���V"OB�c���N]�-�5��,�(M��"O1� �6Qi �� �>J��a"O�@���Me�����f���p"O��K�J��#�68R�%*�"O4x�&�K'@��5`���7|K
�bP"O����FU�<�vY��C�,3:"O��J3��5]u����
- �"O�|	5�Y6^��P�V�^|d��"O�;tO����r�m��#U~Z�"O� >�P&d�0F:�ub1�D
)I>Q	�"O p�qM��=Y�5"�ηk>6�q�"O�q��_`0�*�S�'NPG"O ��&B׀��m�Oʔ7�6�w"O����"��D?*z�� rԢ"Oz�EE��L)(D)�n��
v"O%�ô�´Rt��!9���Q"O���B��󅅌[ކ��"O��]�sO���1%�o0@���"O}��W<C�́��CJ��f`&"O"4+ G�;J�q毑�N$# "O"���Ըeخ|9�.�L���u"O�pk�'N�+ ���E21℅q"O2��EOL�Q
W.�VU��"O���CޣȬq!��,�xl�%"O���ω�|!J��J /�,�r"O�	��IH3x�b��E�EW�NI#$"Od���.��3���dGY�z0a�f�'���'��E#���# ��#�G�a����'Y��[���!���{�B2
��(�'d�����Z; �0���BV4e>Y)�'!n�@ƼaX��0)���H�'�`4���Ԡ.�<�8cE��0��'���F)�=0-�B$��Nd%�'I� CGm�0z��BD�;��i��?��i+��b#�@?'Gd1�á=p�5�ȓIu�I�
�qל0�'J7h��ȓ9Y�<S��v#�lܙB"�CK�<��/֦]
��ׅSء��Nl�<��'�"\����d
�m��ْf�~�<�����a�rd[+rl��Ĉu�<���\w,xT���Q7XdPyp� �G�<��"�5� �:�g�T�~�5�G�<�5��&@P�	��E�+:��!gz�<)��Zb!F8���P�M��s�Rr�<��kC�NZ������	Q^��珌r�<�
Z;f���މ=�捲B�Ue�<4�ӣA���q2'aܸ����K�<���:\�M��I�3�ր"*�L�<�`��p�I�k��:Q��OI�<i�b�=).M�5�l
���KC�<%�E.8��
S��SZ�LkEAt�<��^oƴ\skf���r��Vo�<� *0 q�����΁kR�����n�<��D�#KI.dqC��<�laz7d�Q�<���ߢ3Z� ����n�ؑ)���t�<�SH��P*��OE$B�.]��jCk�<��3�az��F���� �d�<Qp��&��X&��b�d�Ҕ�J�<q��9N�0����
�*�<	�w�C�<�r���H�:(��N�~�ܑS g�<����8�P1�@�S�Q�H@���}�<� �E�.U�}���R>������c�<a�	����5��#�tsB��e�<�A�L^c���f���=���Eh�d�<�B�)o<ڍȑBU�&昘Yǉx�<�hD�N����!ֶ\I�i O�u�<QV��@�6Q�ah�lF�xH�% q�<� ,�2eBsb̰�2�	��SD�<�e0p��AbS�mX�9(���T�<�g�h�4���KгW$�4����h�<���ʕ�� ����XEt��Qb�f�<���[�(�v�J�R,tiH��H�<ɐ,��/1�LC��9`<��ө�B�<� �#��(pLe�ч����{�"O��p�ĈfO��w�%_�HU�"O�J��Rk���r&�Q�T}�W"O&�F��W�Z�@e�D�����"O�)���Y9�
R��:�X� �"Od�2'A+�R�GP�!QT�[a"OP 1�C�����-_~ͱ"O�9�JK���Z7M�G���	�"O1I�
 SR���͟'̲�؁"O�Us�K��b5S��q�4P�b"Oj3��?q&Xt�3�V��f99f"OFE���UTC�,T-�r�B�"O�%Ђ*�5~��@3恌K���"O��K�S j~E�S������2"O�y��i�fL��M�	�px�7"O���gM�8�4b�,�	Vؽ��"O8����'m�v@�t� N8J�h�"OX)#p�]P�n<A��~����"OE!LE@c0�PV�<!�t"O��Gح.l|0�Gᅣ�""Ov���&Gp��0��I0Y=�m��"OΘ�T�C�>��=���y"O�y8�F�9g�v����
tX]qc*Op�!�g����]�4��&6�N�
�'���ö-	�u��ȑ�T��*uZ
�'1���c!�@n�8�al,A4ݩ	�'MR�GT��Fe�3��F�����'�h�r`�·B�D���KͲQ�ʓ}VX�b�	�&���Ƀ�E���m�ȓ�v<*ǩ
��5�P���!1숆ȓO�\��a{�	��!I�k�R	�ȓ_�D�ʓ��i-���o�Y�v]�ȓ0(��K��-%s,(�!�#p
�U��0@-�'-Z|�� �%����T��W�]��J 2�&QJ�e�_�d��A�xl���� Ib�
@mE��bu�ȓ'�r�&c�>�����H�G�`8��J2��1
��^�`����X�`�΅�����IW���h�<Liu �5>���ȓG�|тg��8>p��֩͜9�Ha���pD�5쇖,w�	8����vy ��ȓ.�XA�-�!h=昃w"4wc�܅ȓzM��y�9D�z���E��X�rP��w�4��c�Б"Ar��߄�����
0ٻ�@�6�A�k%��u�ȓ9���s��P{b:����(J����{Y��0.=v�F�0�)�~��e�ȓ)����v�	��KQΏP��
�'���Jb,�g���9�N�Oc�E�'�1�Ti�
r�|h�40y& ��'R���DD�4�v�ِ��04I�yJ�'q|42��n�����ƺ0����'�2��
*fid�)�+#���)
�'��XѢ�"AMb5���N"bU`�'����ǉ^4���&'KL�1�'�U "ǣ|���U�T�KNN��'�8TwfK�t�@���%�G��)q�'|L��T��3+~N����G�\+�'D��9�O�{'B7oE�l��'drC���f$P��2�R�2�'Ѽ���h#i����E�,v^- 	�'WzD��� <�2���M�0�h�*�'(屷�*i[�l�������(�'��XC��$Fh���:�z,b	��� :��j#\�l�2G�Tnt��"O�1 5�:{�(FD�x_��"OF��� <�\4��MCh���"O8�ږ �"��U�Ԑ<Ԍ8A"Oͫ�!�Rl⍀����#Ġl)�"O�)�ϕ�<h��yB�=w�"T��"O��%ϒ*>�>�!����2"O�I������mB�J02\��"O��;���	�n�Pw�=m�Ұ��"O2 ��d@����7-۞M��1"O�B�E��k�@����U�Ĩ<�Q"O"�	ҡI�i��H��L��:�"O�I��${a-��S�S����"O2�*У���CDll��M	�"Ol��
�"�$�Sg�
 �"O,��@ ,�����$��1ZG"O*�8t���q�.���CT2Du&��u"O��(g�:��|��˶rv��$"O���O�|�L�a��5
t�x��"OR�vmԜz2D��"jyV\��"O�l��A�خq9 :@q�̂T"O�1Ӫ��[x�𥬞6Q@�a�"O�1;����@e:�kZ�]���"OzH�N��J9H2��|�J�2�"O�x��	�4:t�	;��+ڐa�"O�A0G�/Ȋ�zEMx쬌BU"O�x&끑s�P��"� C��d�"OT�Ɯ7�tI��A�SSnp�a"O�aP��4<��p�N�B`,]��"O�%ɲ�$��g.��L0��"O�xH�"�5��t���X�P�T�s#"O�X��"[}@
�a�9}Z��F"Oȝ�5��m��)��YjeXii�"O`��A�8%`a��,��*��P�"Ox1T��'��%[�$E�L���"OV-1M	�u�`��>D�Jp�q"O��p��?e��90��B�!�1"O��0��%JO���j�#���b4"Oa;��\���C4* +��ew"O��� Ğ���5�7�$!9�"OM P��]���	����"O���jK4	~�S�pF��"Oҡr�I�pG���FĚ�Al8�"O�-���U�F��X��Bsd�'"O`QP��2Ӛ��7�D-]q��cc"ON��"\�`�-��`G�+� ���"Oаx����YRo�g��٘�"O��0�\pعb �'f^�ۇ"O��G���z�����o^9��"O\�%�PPp)-�
mP.���"O)�6#٪e����"YrBb�Z�"Oxue�^�J9��L�N�`ɑP"OYs�l��J���'�D�||��"O�U@&!	GR��u��\s���"O���5�ـH.^4g�=BU�I�"O�����O�T�"��ɜ_"e8a"Ö�����b�b�$\ 
4B$"O0-#Ԍ����ժclUQ�"O���6J�~_�X��A5�����"O��ysD�*���q�.�*��{D"O��;��2KQh(�R�ܘ]�tpR�"O�Bチ0F�f����*� e��"Ojp��іr���s-�./��IxD"O�,��MOۂL��:��h��"O� �y��ӴW�{D)pU�؊�'%�'�a|�h�#~�l��D�H\�2�o-�y��
$�܀�&�RzD��� �y�Z�m̻�Z�5�����`2�y�f�s6�cCE�>E�P��B+�yR	G�~}R0����D�D��R�y���%;q�L�L�8h�kV�T��yRJ�?��٨���x~���"5�?9/O���d��g`4�R��XI�D�E	M�$!��͡tS|XȠ�XC.�aA(�)p�!�>��0B�`F��U3gF�m�!��[C�\E�"E���P�f��-�!���(X��p8S��0���q��	R!�J�`�4QR7�#s�����CF��)�C��Ĳևݓ ������\����?���0>����~z�Ib�ί
��ڵ��m�<�w�B,`�J!���mJ1) �m�<�a)`�t`S�ǥ`B0	ti�R�<��Ɲո�0�C�Df<+�j�<�%@��3�[�)F�t?��2'(Ei�<�`c
���aF���F`p�j�'�a��dEX�Mrt���
p����y��|�$궫S��A�W㍥�yBg̕d��Ta"��JK��A)�,�yR(�=��Բc���/j0L�G���y2�(u��U�%f�Pj�	���߸�y"��3q�i�@���Hs��@Á��yRCK�SF�8��33���:C�ѕ�y2L�\>\����;wX�����yr����#`+��hV�M�y�ō+E�}9��װv#�R���y��#)�fa�⡑�A9�9C�υ�yb�3z^����I�P�ƀ��y�W�9�h��ɻG�2q1B��yR�͟i���G�:�t��E���y�F<R��;ED����$;�y�c�h�Q�����-�c���y� ��h�	��`#��M��y"H��sH�5Z�B�Y�X`�tLG�y2�R%`�4�HU ]*J�-��ǘ��y�Ęb�4bԧ<����e��yb�S9m�`�2e�B�j�������+�y��c5��$,�
A)�8�y���9%H"E{奞�Q��X���@��y2J��1��<ya�J �MIG)�,�y�'ٗ�5�vhڱE�(��6�G��y�ƭ�����4sr8l�2�I��y��~��y���dDθ{rh�yR��$je�ĽR�pxB����'�l<��/���L�IȫPl8�'g�-s�!ϥ��̸�LI(}E�Ej�'x��#�OL,Z�|I��ꆦ,�������˄g�X��h�z���M!�DW�v����2L.":�,�≁�U6!�đ$`�@ɱ,�,H
V,�"I.3!�D��`�0���̫�����
̘
#!�$/K���qDJ!t�ND����*l!�ވeՂ��A��*"�I"�\�X�!��Q �)��O��t4��$A�G�!��T  YLϕ%L�m��c٪�!��]V�1{��E	,���qD�т�!�D)Y8Y �i5ӺU�/G (�!��W�����N���:�n�y!�d�8;�>)���Ir��S�.R�!�� �I��V�T0���@�J�U:�"O�H�Uʉ�8�2��i�
(&"P�s"OИc���*@r�880)={��9F"O��*၃�UE��"��� �M��"Of��'��cX4�haF��r^�I��"O6����}s�5���$w�`V(�yB
��EO���Ӫ&At��EN��y��Q�WA���I��HF�K��y⭍
 8@Q��+a,��H�y�G�t,A`Uǹ�HI���&�y"�@�"DHSD�_0I�f,��Mq�<�0%E�+خ�{�ČnL-�^`�<1'�_;Vm�x�q"�$���w�<�r�B�?�=r"/j�.ȓ#�s�<ɰB��Ss���m�"C��m�2#q�<	�&LG�}�`0�6=Y�H	I�<2�9�ld��Y��`5B]�<���
u�6  G���soH��� X�<�%JM6,8V��R�S�l!&�����W�<a�Q�u�B��'FN�� �k�<��&��Q�t�zE�ԔRhDhh�L�o�<9��M��1v��2o>((�MOS�<Ie@֐Q���F���;O���gUM�<!󋉷\f���`^<ysx���AGM�<���5(j@YPF�7<~%�W�}�<q�	&~k��f�1�Cl�n�<��σ�ޘaBϋ~�ܱ2Il�<ɵ�'$%����.J����ff�O�<��ب+�l-�Ѐ�lxR䱱�Bw�<�QH�|��p�e�z@�LS2iQL�<q��8��w�F:O)T��g�F�<a��h��@P"��)�*lj&�D�<��ሇ.{�LA���{s����eRL�<��b�m�^E+�c�1���bHG�<鰇�w��&� �i_��x�y�<2�ޑ>q���Ѐ��)��@��w�<�Rm�|�#	�R��Db���t�<�#
�8*���H�)�y�&8��t�<�m�:7�S�Ɵ�DAk��Rq�<	/�X,�l�4.^�Tj*���Xk�<ѣ���g� )�쟺k���$�e�<����*!�����<RjL���\`�<��	�(�jȋv���@�"ׁ
`�<��aA�MPVӰ�4f>YR-�_�<I�Fɢn��]c ��3_�� Wi�\�<)7��
|����"Ζx�� ��T�<IM�_4H ���=L!�`�?T��ۗȄ���U��0<��]�wf%D��Rf��%$^1c!@�!p�/D���ѯ�) j�A@��K<^и��,D���Y�
DHqW�]� �j�g&,D�J7�L�ub:�3G�(�L����)D��h��T�4P0Qi���k $�7�'D��A��ڎc���T�hq���C2D�����z�S��\%`��)�;D�`BcU#`�R8�
��<�����9D�D0�l�f���IK�A
`�8D��n�	`�2��k uj�6D�@z� 	lA>8�e`ŷ ��N D����/��aIn-+e��h��a- D�t� l �#,��8h�����V�)D��p0Џh�^�y�R.�Q)��(D�8�%(O��4q�O��|���x �:D��
%��,dÊQ#��V�̠���:D�� P�83�ڴA݀��� J�y0<}2�"O"��b��=?z����M1%��P"O��c�KA$�]�g�s���"O��+pD��l+��u��T�@��"O�p���E��}�B$��m��4"O�@��CѸ-k��d"��*	��"O�K�Nɶk��,�,"��e"O�y��(��W��$SV�"۶0�w"OZ�x��ōlO�l�v/�l�2Ő'"O4t�s	�08�O;(��C"O�i�mŗ�Pp��.�_��1�C"O|��E�GeX��FY��ɸ�"O�-��B�>o{�x��V�V��<ۧ"O�-���V��G�K� ����"O���t����(�S��"O�Bh�w�j(���B"�>iz�"Obd�1ȟ=K�"�{U��o�*q��"OUA3�1u�05y�@,8tR�"O�L� �@G�,�z �Ұ-�X���"Oja�/TaAx��a��,g$�I�"OnՐ����;�LIZ $1_d�y"O�� �JW�)���k�G6Ova��"O@�B �\'����R�(��Y�"O��83#&tx9b�ƣ?+$=��"O�e AC�`0�����VDI�"OBB����0U�D�9��5��"O�=j���2sXذr�� �\i	Q"O�������&,��2@L��PU"O�[�g��d&t@��)�@���"O��Q��˿q��p8�b.'�"I"O`��B��5gcfD��C�[|��j�"O��{�
]�(�bbΗu��H�"O�� Î�:d6\%�� ��'g���"O���"gX�]�L@�o�'d|�A"O&���T�i��m"T�Ѿ@X,��V"O����œ(����̜NHȲf"O`mRQ�Y)t8RY�M�JQ�=!�"Oj\��Y��H�&�=.f<��c"O�s.\��8��^�k=@}�"O�Y��J�s7J�3�:/�1`�"O���m!��rTBׂ*vx-��"O�4��L�i{��["��6���9Q"O(���A0K�f�I�_7T@@)"O@�EP��hb�Me7tق�"O����A(<厱Hf$�,Q%�eE"O��mȠ9v������8$ay%"O�qx���Q�!� �%AV�Ѡ�"O��@�eaȐ02ŌJ�6oj��"O��b�D���4KL�6�`B�"O�|1���$)TYH�'�+ &N%#P"O�HRpc�,��+R���F0Y��"O Ę.Ŷ*>}�P��2GR��"O�AK��^Q�PF	?^�2U�D"O��GH�x8��wT�|��੥"O,j`ܻ6LrA��@P�i 4�C"O��(��T��5��a?J��"Ou{�f��
r�+��O2TJl���"Oj@����O4���PE���I��"O1
�� _CR�aց[2-�TTh"OT��'X4X�8��*<~t,�"O�pK��j����^^�MrP"O�x&��~�
yP�K�[{���g"O�E���W7T%*�˂K�xD��:p"O��9p�O�T$J|ё`�'��Hp"O� �5�WI�"X������v��ub"O�R�BՊ ����(4�tZ!"Of5��D̿l�ޱ��m@H!�	a"O���!"	6R�.�(Q��E�0��"O�� ��M�-��	iŌ��!���"S"O�@�g��0���ǐDK�"O@���!̠���� G��S¼���"O������>	��8���:5"OX�`R�!�Ix��L�c�&��$"O��� �w���\ }j0�iE"O�݁B<A1�\��Ɗ�_��Ӣ"O@�dԪ^9���E�yve(�"O�!�@�5
&�Y��-�b�k!"O�т�(�3 0>Y��U�N�ta�'`�h�G� }N�3Ԋ��v�{�' ��T%�5-i����.
�`�����'-J@��]��z�I��G��N4*�'G���5s�����-	�5�T 1�'/��s�;hZ�)Z�F�%?J���
�'��9ō

x��򩌅:-�`"
�'�"�����+b��!m��-i
�'�<D�Sŋ�e��ȫqmڴFx�C
�'�b���[�&��pBM��C)fh��'��T�±*��`���R�p�'�� �$��'C���EUFƨ9�'k��2�����%j*�Q�y9�'Ij�X�N�r���C7�ʶH�H���'I��@D[s��`��E���'\@l1բߝ��ȥ#��ްj�'F��a�C"pa��ŏ��`)J�'�~@2�Ƶ(���b�H	(���K�'��l�B&]>l�6z��Pu`�'Z=�+��w��أ��*}��%��'�2Er �۞{�{����ѻ��C�	��4�&.�1w���xW���C�	9n�&�h`�K	 ������j�C�I�1�0]��KȞR�.)s$/[;-K�C�	(zj6Г�%V�p��U��O\hrC�+St����SɊT�/΋NԮC�	��
��W�0�6114�� ��C�IH,�B��V-C&���n�K�HC䉈738Q��凍W�m��C5B�B�E�����LϦ���t��C�	��\hJ'\�2���"��C�ɫ`d񓔧@��ٴ�ؼ(��C�	q*U"��� ��4 2��;l�C�	#�q4�ðB�q,Դq�*B�	6{���d�݊ ��@P	R�0�(B�+i�d)i3L>�ڕ�a#w�B��9]*�wcϟ�9��MH�&s�C�	/ Y�3�"Ü��@Ƃ4��B�ɟm�l��U�X�8���2�C�I�P���#����n��)�}> B�ɉZ���w�V��DX�fi@�K�\C��)5��@�b��!�P�0�#L"I�nC�ɔ)�8�B��^�n���DK�X_\C��fk<Q�k͚�"���n!!k.D��i�g��H
�xҏE�՜�¥.0D��"`�+$�b�Άʬ����#D�|	 �#86�d�ףM;iˊ��� D�Đbi[�r�:i�E(͓`��@�W�#D�@OY"�� �
M�@�R����"D�<�1�N R����h��I�����?D���F�h��d����8��*D�� NY�� Z�0��钸Az�t"O ���D>,:�3dJ�	 � ��"O����Ճw�2���i��5�^��3"O,�y��
Cm������o���"OX���E���:�؅:��e�G"Oʽ�Q\[D��	�)�yL@kt"Oҹ���/���[p�]�'F�@z�"O\u��KW-G�N@R2$!�jL
u"ON�`��
��c�I�X}ٷ"O�S��;v��a��T��q�	�'�&L�E�N�o�e9��8!M���'�� ��c
i��&�B�Rs�'�t�)B�Se=i��Q-�䑢�'��T���ѱ/����$�୉
�'{*yʇ�(|d�v)�"خ)h�'ǔ���D��z~���@��@��'$�YB��H':\P��14D�t;�'2ڱ���^,M�T�M3]�0T)�'��4�pC�/"z��T��*�Y�'1�h� 9��]s��%{�ڥp
�'Y ��5p����a��"	�'l��s!��p������^��	�'��īW�=	n��BeY�CD����'Of�+"olHHD3ej\c�'9��jу�t��m"q�ڀ�`�'��@���)y�Ų�K���^(��'v�Hx�&M�G LȻw�ܶg���'sN��jE`P��jG�w�,��'Q�s"�@�h�1۱̏�>]PZ�'�B�P��/[B�I;�g�73�h� �'a
���Oܤp̬���+�C	�'����b��:�<a�oϩ#<ҹ��'�4��J%B�N(&C��I�x+�'��T�����iRBl-G{�г�'�h𘔥�#7�j,�ƭY�<I"�	�'�RE+ńZ9޸mIuN��B���'��KJ5%N�!3�\����'O�q:��&e�0�'��zV���'/n�tE_)���f���mj�'(���DZ��xم�&��'>���D�H[����߳L��j�'���*�	?�L�!	�8Ly$X��'�b���L��2�&e��NU�K��9��'^��k#O�2�D���ۇA�����'��I�Þ�&�N#�M�=�H�h�'L��M@�.2�|���MMBn�����Y�,w���Z#O.��
� Y��y"G��Q��!ᒌGjEJ�7�y�,��'r�ajU)�":������!�y��>_I�[�.�*������5�y�oM�nҙ�QMՀ�N˒�yr�}��	��/ڂ���h�jS �y��ar�LA�.�tl_5�yb`���6t�w��1��(P� �5�y2�s�0Ը���$���T1�y���0���!�ar�(A��y��
bzr�Jp�	�+H �!��yB�����d�`0 d��F8�y��2H!6�˂��h�٘���y�@:�X��\�r����ybh'S(��b�$[�
�̸�y2`�$V��!a�@��T�$��֢�y�kʅ7,����[u$)C���y���0Ip���!ì P��� �y
� ��!aQ�U|�8� ���B|h��"O�<����_���Rǹv�dw"O��#�N[�V��l��[?n�v I�"O�С�Z>tG��g��7:�~�9�'7L�!Bύ�z�ظ�Rg�C`�X��'�
�Q�E��j{4)��I\'f�^L��'�~1���{���k�
ܷ9t�0�'ܥ��H!8X:v�\�Z{�'�v�˰e�-"%X8P|8��'��A�!�@I�]�Deʸ>3^���'w�� ��&\h��'ô5�,(����v� q��5U$��8 E�i���Ez"�'{T�
�l
�.X�!N&U>�䨋�)�S��mF<�L���E("�q���;�Mk�'��(9�L�Se�0 %
�D.�X��'H��&�(��;D"��h���!�'�6(S��.bL4MbS�^�Z����'¶�0��;P�h"*{���
�'	�ّ�ģ<�����V�dh@�	�'?��� �ph4P;c�G�Jq�0y
�':���%&��_D��z�j�;����	�'c����&t�d9�H �,�v=�	���'�����"5�4Z�8M�L
	�'�v]����!'�VUS�d)/�,�{�T_���'dv0rQ�	�Z�v\��[<C�ܐ���̴D�1#�ٺ��"oO�����JZ��ϟP����pG�lf�e�ȓo�Aұ�X3t��Hڢ�ږk(�L��HhV���T25�
T�D��
k+��ȓ)@�z�j�Iw���t�τZ��}��S�4���ϻa(�+���,�T�Γ6Fb�<E�$�D�2aA�(�n�$]I揕��yRW�-�l"��"d�6�˔����yr\� =L�6���1��{� D���'�ў�zD$��K#�큂*Zj!�B���TY�� �����'�O��HX8g���`'�<B�C�idўb?Y�'���(R��8�Px	b��)� �'؎���� �r�4m��OӉi:"���O����T�v=qv��,�h(�w�K#�a}��>a��J�T�� ��"�H�8�X7Cg�<VFӤr�b��`��+&�"h�|�'�#=�Op>\h��A)%�(�9�C��!7��I���!O��B���2M�H򠮁jH$R�"O*�Q���x�SN��/>N�b�"O�Y���5�>4��M�
�d1Qf"O�-�b㖯5���c�� �xA��"O�����~S88���,{�)
f"O�EKUC.Zu��;bK��$c^��f"O�1	�kB w���!@�a][#"O!��-F45>*�����"��qSq"O*% �aL:E�2�6'J�@�5"O�\�Ѐ5@X����� �0��`s"O\ kr�؃X��j m��u��"OZ�Č֕Ub��:㬟�F�����O�=��V�>�"F8 �L���F�#U�����z����>�偍%Y��0`ʁ2��4B\�db��D{J|��ފU
�� !OK�4%�`��I�<�u���K��͒3È�c92TK���ɦ!F{���i��XR�H��60��
��d�t�p�'�0У�Ǧ4v�mчE��a����'�:�)�o˯sp8w��Y�쌐�'!�y{���iEu(s.,S��Ds	�'��a�H�ו���
FE]�#>D��R��(Z
��!M;!��V<�O��$�>� :0�P��d�ɰ1��'t_P2^�4E{��	{��P�poK0%��M��d�0K'�	ɸ'Kў��х2=��h5�&O��i�sjQ0 �|"�"}���{P�I�G�(1�H�X�/���p<!�O��'d|�qFEȽ
|f�#��:�"D����]���iV6ey����M\�أ��>v!�Dŏɚ`��F�'�a8�	@!�XI���e՞Р,�Ï�-Y��	6,#Q�"}z�݊!S��b4d� �^(*aL�a�<�&nP66NA#G�_&b�1��M[���=Y�\4
��kdF��1��b�<1 I9T��(&�U�l}�	Kw+�W�<�rO�Kl8����X^U;b�{�<�g�J,UY�`[�
�&%�P�!�A�<i�n	d"FP���	8x��KY�<y�����%AMн
�`q���E�<����>)�Y�^r���4��Z�P}�5�U���Iqy��I!H.1i؁g����mM��y���#.�X�U��=Yڍ�2�L!�y��&���
��%Z��B��<�y�.��Z�E�E���j�!E���yR�ĉ,8lTz�C i�6�ܳ�y"�̺�<����ԏO>i05nN��O�=�O���3�� �}����.�}�ĨJ�'-R�W�j��
�ܐ,t P!���7$F|MFx����Dn�)`��ƍN=�:y���"O2�=!T`�i�`�
����Av���D�I�'L�?MC�,(a�F�q��0f���:��-|O
b���2Ȍ' ���qE�0j�\Hj��/D��W��g� �T�r��Z�'-D� �t��=X T�# �gif�@��>��4��>�E� B�̙�ա�>4O�i��ANx�<a�*�>D@�4a�#	jqb/�p�<I���;�	���>DKk횢>����X3�\Y�B�эZ�L��GڣZ!�䚏]b葴� ��)��%u�!��G}0�E��I�c�(\H�V�����N`���چ��*V��ybK�7Y¸��'�3D��P&)��}c���?E��r�0D� �ec�]�h�%g�%<�ZIP�/ғ��'��'(�P�����A���"��{i��6N��pƉ�Z���)�� 5l���+�RL�S&�n�։���/{*P��ȓ6���2%D<�\	����H��Ć�Ld�Pǩ��Y��ɠƦ��i�N���M��e�$��+9�5Y�d�rՅȓ ��Qӡ�/.@������,3��ܭ!$hΛܬ#͖cc`Fy"�'2F���2:�3`h  A�'�0���v��`͆+,2�m�#�<$��P�/7K����!���r� #D���6ͽ"�6=14�݋mtr� �"D�H1d��X�r� F%��f��C�!���<ᓬ�e����T��^axeEP{�hF{�K[���$J_vv��B�T�j�n� ��I�l,���)�E�� �5G�\?�C�	4��������XZ�^�C�I~���FF�sq\\x��l��C�I#!ziZ����<d�jSXB�	�R��=h)���M���w�����\�k��%T͌U�R�^�u�!�_�`ܶ0Q��
�Xhl#$��T��)�'n'*Љ���9�p P3�S1%�V�;�'Yd�RQ��N��(`2�D��LI��� �)�1~�apQC��f
��8"O:�z����i�4�B"i���"O�5�����d��"��j�v�9�"O���g釉�l�#����M��(��"O����`�L3)1C�]�O�zX��"O|���vRr���k�?J�09Zf"Oz�X�cF�%��	^k`���"O�q
2OǭFGfe"rc>��D�8D�@9�+D;n�6MY�O�#m�r �56D�����Z
C��b��mP���5D���T*[�#P� B��a����4D��
`�N3���/J�{��M��N1D��;�Y�ƘX�+M�(S2d@�-"D�� d۠j� �i � ��)B�%"D�����i�x��Ȝ�b���B�:D���R8��8 p�M>�9�f!-D�l�`�����۝:u"�z�	\�7F!��pL�����Fr�L0&�I�B!���+X��;�-��c��8�R�B�o;!�d�48��d�$I�aA��3v�?2!�{r�j�`ϣ5�i�"јJ!�@W������,.!6L8b�M"s!򄟭\�4��X_�vCTAێ4�!��%R2�͊��H�9:#���!���(J@B#P5V�8IRdӄ>�!�D*�F�k�����.H��� h!�䘩w�����9�DcK _!�E�t]pI#;ˤ,pT�-S!��	y�EZ�MK�l�+��c7!�dD'��@�
ڛ!�(xR)D;5T!�D��KNt��e�(�I��QP!�CSduj@EƸ~��(�&Ρ)�!�$�1\�A�53fX�D(�#\�!��܀B��b�Č�:��@\B@���'�L!w�/L�0(��8n��	�'�)��� �#���Ca�~L@PS�'�fT�PK�O>�t�fڀxR���y�]��zF��&�ZĈ�4ؘ'P>�y�� t'T��� �u���+�'�<e���%C��!�M̆RU���'H�P�-�+�p�EA\O�8A9�'�<��Ǣ�|�t�i��A�r��8j�'F�=j�QJo�Xw���A�'�h'C�P��!+"�L<;g����'�̸�E�6?\Q����=2�m
�'�.�:DF�4_�n呀�7�l�C�'Z���WO�
Ŗ��fF�#p$���'���[
�o�lA���$	z�"�'
x�9�N�m.��z�ķruU�'�2ջG� �,��}�뚉�(���'זQ9�&Q#h�m�����Y�'<�S�?v�i7�	y�� ��'��a�^
$�Q���C?s��Di�'� ta�i�(P-�� �z)^���'r�u�A�ؠb
��U.��Y�,��' j�a G�'W<�T�ґz���{�'u �h��a��ã�#�0̨
�'���h�=1�(Y��ژ�Vp
�'YH!�5枛;� ��勇 x�A:	�'�j���JT�	,�]�E�Q5w�J1z	�'��<[6�L<TrTl����=_��'"�!��]147zQХM�ް
�'�L��W_M6$�hT��+�us�'�L��n�tԩ�C��;~w�Z�'�( �C[b�*���b-l���
��� ��B[�kB��E����6�8�"Oܨh�N�vH��U2�LqI"O8��1�N�j�=!B�����c�"O�ka�]4JK&� A�5G���e"O⁡���4PP[s ǜm�f)0g"O��#�N�
��yb�ښ0<�W"Oz�q���<��P �,2s"Oh9��.��I��<)(�5Z�"OLЄkP�Q�T����{�� �"O���CAR�j�@�`!e	O��ˑ"O�|�u�^�gaH�H0��Jݹ"O��{�l�6)�2]+��^�Y|�t�"O��֌@>]F,
 �G�#XTp�2"O�8�&��#5�v�s��%�d��""O,��E�"Pⰲ1L�:��Ts�"O CB�z`V,qU�B>KV�i��"OJ��X�#&HaBˋwJ��ZS"Oj�x�,�C:X��)��
��Ai�"O<�3��>{Q��js�6f����"Of�I5�ީ�>��G,ؚ'FŲ"O�����10�xtS)�X ���"OF �D�N6�y��Ѷ_(�$�"OЌ(��N����P�x'v��&"OJ��#M0�����'��I)�`�g"O�p�U�0O\*����ڲ1���g"O2A�7���vS�`� Y���ɥ~*6I��FD�O�| ���\ ��!��B ����'�}���� �ԽЄo�*Ȑ5+sܶ|�<"R�K��s���3�(|�\��+Ԛm6����+D�0��f¤���@�"'9�����O$D�!	ˏ7),i�c�>LO��S�fÞq#��kԨ��V&b��'�2���%�"s���s�ƀ�,�|=�%��hd���E�Ј%�!��X��A�X�KI�EP��ן`��O�³��" �-��/-§9h���jXI���*ZX��ȓG��M�0�)D�T��B��� RD�އ�.���hy����p
T��H�鵏	�W^x�qV+.D���r	�$f��&�Q1��U��O$p��mn�(i?LOr]Q����)d��TH�3c1�D���'�$s�#�?ebEq�kX�v�v��AaT�; �/
^!�ď*�xu{q�Q9
ST�+um��a�O���S�B�V�����&�'`�b��4DD>R��D�P�*�����Jv����1;�*���kZ�`�&0�Dg02X��C�"}��9Ol�hKH "��m�p��u�q"OD����Qp���y�oƉG��HѶ�O���ŅL�}1L����2g� I��-KR����2*_!�D�&L|�@�r��O
pQ��fJ�!�L9P�d�I�b\�1�إ���м\s!�$MZ��r"o�4'�P��l�lk!�dc�|�If�Љ<����q	�'\��$1jU�m[�G�%l���LA3�ޑr�^6uz PҶ�,�Ox���jߦ��3�I>Q�� ��'1$E�feT� K0�"�F`?t�%6���H\	[w ��aρ[�<�6JEI+�`�>Pd��\lyr�	�v\�զ֡s���BA��0f*:��6�,/Kj����ȽS��C��/@�By�d�	9��পI�UIn�R$mՓO��I	m��\
$6�����0$�|P�m��g����Em("U�rH�5(vE¦�\�j:25�J"7�� �V'iM��fc���a|R����AA���%IEm���OB§��dZ��g��7R�B�S:�`����E�r��aaG��2<8B�ɵe��vo�/~_H˥BN)_�˓��Uq��:�d`׍Y�)E�#}��"Κz���r�̽t�+���	!��+v.yz��@�,�.=A�%�����&uY��lR PFʰ���{��[����\���������?�#�$����4 �\����}�9��6+�RY3P�
{߆ Ё��c��� $�0"�4W���Ʉ�ğ l��e�Iࠩ���N'm!�QS/�.�A!b�r�(������JB�qjf�M"�yb!�8@%29��ƢOނ�ൣ���yBbZj ��m��^9����;F/<-����J�7��Y2���	~pV� a�ٿ]!�>p��J�"�
�.4j����X��pG��c!RЛ iB�dk�0�q^?!k1b�ɘ'h�D9���L���p �-,�[����;�Q�#TD�k�k�SR�����Fj���iS��p�+ue�h��0Y�f+LO`���ݟx���$d�|�ٙF��h�h��b{� ��dU~����W+��y"�,Z������MZc"O���7k�;���i��@Th�p�٭~�� �����R8D��@$6����+K�9�1�� ������9��Ug��	PF!�;6�����
Q��m\=JZ�K#���r�@F�f��X��N����dπ�"j�x�y%��-@ֱ�G��D���x�F�,��=AD�ˈTi4�"�ET�(0���H</F:%c⏀{��ģ�C�/�"���$R1 �̠��ĉ<H:�7�O=p�kB��Zܠ�+'";x��?�t�G.u��K�ϑ�8���WMLb�rQg9`O�͠��$XdC�cC�@'�`;���I0S�H���iC�i�*a���+# �"r'É>0����S�)��b/&p8�С��.j�&q����3���
b��T���Zq пL�6��1O>��-���������`<	@���Bz��X:	�����U�j��\Pd� "�� �>P���{�L���P��*�G��}�$�]��D�3���۠	���-�O ��灓&s$#��8W���G� 'I��-Q�n��#%O\�r7l b�d
 ��Oh3E ܨx�ʀK�ܤV}fuH�cMb�A!�)L9&<�Eb�OƘ��S�tCd���N.
�vx �il�Ӝw`��;u��%D�J���f��7�,5ˋ�D�v������Ɂ�:{b������a�|�q@��YW���m��P���BJ��u���;~n���,��`���<Y���@Y�W���,VP�X$�S?�"������t
�(\D�D��<1�"�D/V ��n�����(5Pa*6AA�ők�f�H���VD��'E,^��¯֊9?���P��e�	p*����'��h�C�
{�\��'�) �F��z��Ř&�������ܭ��j��>W��@��3~@\P�=��P	޴m�*�`�m
XtX;�O�MjP�&M	S�l��O�̸�m�$���r���i����ɍ*޸QB��:NT�![��ɩ
���	[9��Oqa�i
9�(�4 �Go�&:>z勣cT6�z�KWDÀz�4I�sC־8=L�x#�W�wM  ��$=2n����~po$��,ٻ$�����#9�I��a�8NȄ�s<O^9�n8����~
�2d�\�<!�LS-S��q (_�jr�l��@�C�:�ReH�5���f��'^н�O���|���i�H��
C�_�� �CO�=��0�&-/^�4H��܂>���#/��i�@�'(x����^�gբ��2�>+��I��۟o�+ �i�&I��C��� ��o��'��$��|�v��5j�>e������	RH��U���D�]���	�(��!��'����&{�7�'"*�(��*=dB,b2m�0z�����_�C���v��-��	�6� X�3��_|�!Ư� �(��8#G??2���h��1y��'s`��a�z}�I
J]���cC�_��?�I"��iڠ��޼H�:!)%��"��)��Z��?�dO��TN��>�O�����3>�m���yb<]�#dO�YI�%�lP���)�'�u�d� q�����fK1@�|	���"8j�Ɉ�=o����4r� ��qL�0�QCP�G	��I�q�J�KǉO��s�^�+�G���H4�'Q������&y��ܣ���D���K��\����OX p��&L�" ��g4��>9  +54�8��
�ȟЉ`Q��:m@ ��	#j�d�!"O
��+��
�M��쉰fX�X��H�=��ݔ'Þu1�b�g�#aYի:vǌ�g��6N�C�	�Fj�%xL�.�(�����+�5a�F%�����'�Ɣ����?b�beK����ϓb�fm[ҩ���$�	%�xaP1a�G ⤂�/�E!�d�U)$59�Œ�Ę+���e�!�$E1z�朡P��
�21[Vl�3�!򤂞v>l� ΂%k�:�jv�X�R�!�d��F����f��I��顲��2!�d�7Ly�y*f�S�y�x	����6!�D�;C|h��ǥ ���Ӑ�ݦik!���gǢ1J#�3R�������Y^!�d��W���iA�6"��"��&2�!�d�-]�0�IǀQ�a �ћ�ż"�!�ą�%���8E%D+nט��&:Z�!��({ߜ��,2 � ���q�!�dF�%�|�z����/qD��S1M!��%LgҸ3���� Eĕq�b�>!�D%��UQ�ች����K!�� �I!�I�t��"�Ι�{ X���"O�l�3DP*b(�y48 P�5D�0zȏ�"��)�(hs0����&D�����:zk�=� �F�+�>�+�d"D�`AI��p��E��)��`t:D��{�JE�0d��!�+|���Q�8D�8Ѷ��V�h��SM m:f�q%�7D�����6@�.EZ��LX{� /D��˖���X�1i
|	�e�S�,D�,���� /4l�&\f]�H'D��W��(0)@)��l֦O��؀�c&D���RkSd���0��=���ei0D�h�u�"�p�n����2�I3D����A؍L���rЪ% ����.D��q�O�C�h�9V���Bm4�20*Od5�t���?��(�@ΣT�`,B#"O�|�7Ě�P��jO�.,s���"O(a�YD��;�a�&���w"Oδ�E�'o��ź׮Ml$X��"O��@���<� �OU��"	�'"O�L�0+
�^���׮��<���"O�Ճ��&$� r�oš 
�2�"Opl��#D42�Ē��$��a�g"OE;� VD��5��:�.$�"O�e�W�����UAňEZ
� E"O$��@
0m�$ȇ�F�5�V�!"O�a�*��ȔJ�$T*��3�"O)��:��8Ji���R�"O��YąE�T����+`%>=�"O.�:�ӓ	_�IZ'�DO��u"O����3@z8�gh_ R�*3�"O<X��(Ԭ)h��(�� ��Q3"O(41���p�t���.�=����%"O��*�a�9*C4x
��Ѽg��R�"OD-���ӊ}`�F MQ��2"Ob�!��B�\\�󅏕|6 d"O�x fΛ^|��Ӯ�|�����"OL�
��%4��`(G�����b'"O~��I��h���[1���<=h\��"O"I�s,L3V1�!e�H@�IA"O��u/��l,�0G[B��5	$"O���!*�\��iH�R�P5�T"ObiK��ښ~ٴt��)�&��"Ou#֥�2�lTK^�z��p�"OJl��,�;M���94�W�Ľc�"O,��!�_&��ـv�UD�Α�`"Or��#[�lo����J�l��1�"OF�����Wpx���hŦR��
�"O�� ���?����g�X����"OJ=[��v9��QC�N�ri@���"O~�V]H��"�Y�QM*�"�"OL5��]���b��0J)�a+v"O!ၩ��i�*��Xz�ir�"OD�iF�ߚ"�2���.̛0m��Y"O`x�`R�D	Z���C<��"Ov�)��ֆ_�^2	�E$�4x"O�%��;�"��҉&-�&"O�\0��F:(�<�E�U�Xe&�@c"O��)/���� A�yH�"OKI[�1�F+K~b�B���ybo��%Ę��"��z��I@˅&�y�C�1rqCp.J-V�E:����y��N8W�V�8��[0o�"ya
�y� Ý13@&CZ@�p1� ��y
� �}�7f0�ҦJ�)JHK6"OD���  )΀��#��E
l�pD"O<�@�Gͬ���H�:>4+""OB�0t���b.����&Ï���+B"On	����W�\<�3�רmH�C�"O� ��+KNx8`&)�7T!���P"Oh��2Ϝ+5d���DK�)����"O�0ƅS�<1�#�͜v��(�"O�99�H��,B�4KQ? T��"O� S7@x � �B�|b�=#"O  su�@�,�2R�W-UjR�[E"OB�
�3Nmi�ǝ�`���@"O0I���$�8`�B�i;�)�"Oj\�.X�pƑ���8;#�]ې"O�P�)��T{V�&y�1��q�<��R�e�I9�,��6LX�h�I�<�M�]�\a坁:֦@Y��I�<I���W���fL�'T}�pp�AS�<�/�CYD ����\$�����q�<��^�d��` �͎c�&P��P`�<�F �0`N�8R�G̼����Y�<�Un�0�ƀ[��L Z��{3�JB�<@b^�&�h=��jǥlG�Ek'�C�<AӡCq3�!� ,ωm�zYK��Jd�<�1@�VƄR��,w���ĈD�<I�G�8W�N��dٮM߈��d�
x�<���46�`�vM��W���32��u�<���V�<hl���b y+f(�[�<Ѱn�rhvq���#$5�,#���R�<�q��.2UR�Xu�ӗem>Y�J�'����Q�U.3T�>��H'"s��q41�T��C/D�,94��L R��¦g�<�Y�&��Bgy�T D�S��yB�Dw��B�B����G��y2a�*-�����,���E�?�)H�s�.�poB��0=1�i>]�}3�F�H0�:�/
k��<���&�r��>6c�� ����Ĭ���W$rk$��bs�	@A�y��P�
D!R�n��?9
P/7��ls ����؉SC�Ha�l���_X�X3"ORab�̒N����쐜O�c��'%��� ��m��	U��~@K�K�5�gD�Q�@�{�$���y�H �lqw`;x�r1YpÇ:�?Q�Mq�����W��0=pk	4O�(f�:
�h����R��������.*	A뉴8X�"�nO:(��d���E0#;���ȓTuR8�֯��a3�X1�CG9�d�?!g����H�߿��4d�" �!�x�a$D�HvƁ��"O�}*��Ɯ#w�`闣�3!ˢ��v)X� �f�"���)��<I"�S4=s��ɴ�\��ک2e�WT�<qp��.�������|J�#�V?iP��-&�"(�ۓCV���ЩQ���`��-P�Nd�ȓo���zu�:"�f�3'�;}RɅȓ;��l▣�<ZH��&��2[�`�ȓ�db㦁$ÚP�щ�@�^,��l�걑�!ݤ-�� ��]�IZ��l������;M_��@�+G�k!~<[��?�L��ԅȈ��>qeʉ5�T�8U�݈H�Y0�ICl���䊇(�BTm�(N�d�$q\���@���VEG+	�!�ě6ވ���2�����7�剖.�XHf�L�Y�X����E�O4riA�'1p�8ԃC��pnR���':���d	�#�� �N1wK��Z#��#{G� (�� �X0#d_���g�7)<DP��O;.����$jl�I��	�5.(t��� }��i��6T� X�o�mP����C.i���+Mm`y���d��Z'�W�L��?�U��TT ���\;Y7<5H�O e:��}488�������
�'��y@�^��Q��v�`*Oh���F�}<VP���&uX���� ΍˓��3_�@y��2D
��I"O|�@�,�? � a�$_�vq���	1��pأ���b�Q��/�;�ϸ'�.܊c���R>�|J0��kX*�X	��$Ĳ�:�X�I�:
�0Q��Y�YHtЉ�j�G+��� ���0=�Fb�#_At���+���
Db	h��� C�*�|L���T"ATiq�QZh(}XC���.|���N�@B�Ieq:��v&ؼSB8�v�Q�EL^�'"��`v�ȣ+����b�O���G�D���x��Dru�^�$�mz4���yB��h���؅L����b��p�|e���^�[�Z%�H�"~���nV4:¬��` K"fe�C�ɰ]0伲@�5C��I��*	;��	�e�)���T[azb�#1<B89D���w<��huMV��p>��b�7\'�y@��4t����ɞ4]��s�^4S�C�I�SP!�ץP�Z��mC�	�pz�<�AׂU\	��0�'kxHt��`I(A0�D�3A
�p��\���:�9����p���B�,�CpS��pi1 �w���O|�:S�P$l��4L{I��J��y��[/������ [~lD�D���~b'�% :���g��@��/�p$U"�,�aE?�O�@�LxX���Wm8JY���Ԫ0-:ج�0/��y2e�j*d��L1.���h���(Ot��Q��i l����A�H�X3-اo��
d��h,!�Ė2q���$�jq:����AK�6nQ�Q���RG�|���i>��#�lΊ���f�̓w�̍�����xE��h��TP��GO<l(�
�I����d�=�5��'��!7c�� ��l�vaĳ4I�1!"�p1��O�E��O0�v%A��ͱ�g��}��)�//D���f@�Q�� �����4�[x��S
X�ه�ɽ0=4 `���5��y�2�Uϔ��M�b���Ň�2�y��RC����� ^?��C���M�B(�2ހ�"~n�x�ڭyEˇ:�0����PN➄H��_+!��������yt��8K����.�R<��A�O�Q����6rc����,i;n�"�G�H~b��"����v��,��E	�c>�8d�G�F쩋5m�kN���-B�����8s�|��U���BG�p�ϊ/|�,Se�]�(,lDAp��<�'�0P��%���&}ʟ�q�CT�Z�"P&N%+��ZRdF>�'��Jr�~�`L�O\6H�դh���%�(v�\8!���!�u˳�ЙRY��a
��S��M���P8)c� Z��֧fN\�˄ojd ��b�K��j特M��M�6�P�*g�S�ӑw�yЇ�C88�jX� ع[��	��.��S�G�b�'�IX�G+�+g[�,�����3��*,a0��r.�#+\*iH��|bn,�S�.f$���.#+[ �K倓�O��J��;`v}s��+}���}�ĪFnLv��?=
��G��ҥ�n�H �hP/�O~�*�i�*��DF�y�
-�s�W��)�Vcܨ,A�� ���F�@�Fҝm9ґ�2T��*�G"N{q��'��qc�K042 ���7Êa0sO�41�s�aCP����K�eR#v��TI�	6�2�*�$T�5T>	�� �K�@�� �A�0�
�DY�/z���'��)9�%A8��'��5iS�@>�~��S_������50�|���#T��
0�2�O�D�5 �%�?�Ջ!�&�.%��p�e�:ep�'ij����3q0������ɾ��S���"�r4"�i*K�,C�	2��� ��0,&�8����p��<��(�9���ؾ0L̑Ӌ�L>1v�eM��#��ׇ]Ӥ��DaXH<!&�����1�F8O���� �}�QaJ0�j����?F|����4?��X[W
 �S�y��Z4>��PKG����nD9_�����
s�<Fi;D�(��	?���k�d(���U`"D�t��aĽT[��DmȖJnh
2D��9G�^�g~*��3vd�4m'D�08�`YQB�)�O ��ծ0D���֬�GY�<�p�����+D��;0+��zDf�+CYfU$L$D����TU���z���LW� ¦�?D����bS�C���@�DCĮ�!;D��AVlK�V����$I�g�@M�EO4D�h�ԋ�!pO�D%�#�J%2�/D�� @�;S�H9YzZA&"�?[a��b"O�4��ƒ�6��BBCi�lµ"O2Es��?h�J������12"OD���Ͼ��3��[�Dm��"OL�K��&�ڔ.^�=�*1"OnY��%��8���-sZ͙�"OΨ2@Aۗk�(��1&se�U"On���p��t �.{��(�"O��.YC,�A�WcRl�s"O@4 `HQ;B&��QF-�
Y����G"O����X��1k�ѹa�P�"O���T�b�dؓ���
�v!��'��0�Ń�z'p�yu��6KJh��'6�U����s�>]�a��!s�		�'�� � U�B����adȬ��'x*��Y�i+j�ᅣ�N`z��'�mS�F1ej*X�9��Y�yƝ!�Pt���x��U3%](�yB$��&�������y�����)�y�F�sz IIw�?vGF����D�yR���	�~q�5+o�l�8p���ybN�"�~��K��gTN� B1�yr#&j��<����Q�`����yBϔ5���:����i�'�S��yB�q�İ5$�"���ԅ�y�-@�YZ���M'$*t9��
�y�FÜo�� ύ,&˚�iB���y�`νB���a���hk����y�	C9I�uQ�R�"Li;ӄ
�y��N��@��$BX�	v�s���y�H	2� =q"��
+q1�J��y�g�H�雳��H3 yP�\��yҧ�7!N��ئNވD����oZ��yb��BV�TС��O��Qy���y2bωbF�8F)]+@�����Ǣ�y2J	_?N�!��E h�B3�[�y���_���,��M%$���O��y��K/7'a(���Hz
�C⬅��yB���sS�HSj̀3CP9��h��y���V���׌C�6䘅)��� �yB'RZK	�#T�E�R�qwV��<}r��"�ȋՆ�8�g�	�]�ȓV�f�#� i�Ж��?	%�Ȅ�+�� t�*��PжdZ:�t ��8�V� ���E�1���ǰW���<�b#F�P���c��=]�U#d�ـ/7`0Eo�?��� � |�Z����z5��'�
�� �m�b��x�)§/ra�W�\�L���@jJ�.��|t�����0��S�O�
aY��͈n�l�Ն�
�&D��PU�ވ��y
�'kZ���
�kw&�8u�P���Q@̓u�T��(`���`)�5"��0x����@A<c�4p����ا�Od`�(Q ��Xn�M�B��V���O޴��'JD�S�ORr�ۥ��$6!�Dzc#u���'��Ij�
$�������Z� _� <�s��36��h���)%1��e�?Ep��0擆N�֙2ǋ	:���{�˙.�m�4]���'K�8̟JЩ��d	RS�p�2$�(�����\*��D�Q�"|�\�5��(J~j���k�<a@�Xq��h��4����%lc|��D;n'�(���:Q��壛W�D+֬IG(�1�F�E�'`�Y����:Lᥡ�%S�H�� K�I��a��)��Y�q��Ax��ϖ]w���P�R�F�-��<��TE�(u�P��s��M��u��Y@?y�b%��?�1�}� ��?�R< �
�*sF�q�[)Nm��
�>� ���<E��i��	_�vP���_�=��`Pg�Δ!����'�(��$ú{t�q]w(Q? ��9t�eA�"@�ew���e��̩�K2 �(�äE�(�a�� ��bU"2���Zq�=��M�bnۮV$�(s��/��L��O?�� �a�"삯5
��S�&� jς�Q!]�.�,�R�`��Tsç5�(�I�P�I|��@�FN��R3�Rd�
��'4Xt� 6�,J���q��sU�K,�bE�s�"D�L��+r]�dI�0|���@}�I#r��<������G�>��e��ݴ"FN����ٟ�|����2Foz��Uh�\cT�����3�B�	3)�	2eȕT�HIF��,)��B��3n�n,���2W�L�I��P5�dB䉴����q����E�O�8�FB䉠lE a��p'BL��iφt]B�ɦtd�XГ�٨c��k�k��v�C�I,h�|)�Q���v�u�,u�ȓ]Nd�DH	xŻ��ǜL���mGZu���͡Z�����)�>~��u�ȓq|�x��jX�A#|��,<*iM�ȓ	,#�,Y�Bq���� }�8Ʌȓ��{�̍�C�6m@ƂY�p��0�ȓ��Q�튿!HV�c���5R�:�ȓB��9��+lV��I6b4CEa�ȓ|ڲ��@��[r�) E��2M}��ȓ}�p�c�ِ]C��Pdȱu����ȓ\P��V,��k�n囤�-7��$�ȓV�zQ P�ْY�lc���&w?�̅ȓ]���w��y[��B��#*�V��z�@��k�mf u�E I�u�R���y�D��唞z��Z�l��`��.����rD"�Z���}��5�����B��b1�3��1_o�)��?ʜ�/z�2���oX�(��Їȓ VZ����0%�84�b­?+����j\LVb��qLH-�$�V��V��ȓn��e�hӹ&`x�*
�w�䉆ȓm�,(� bX��b�(	�p��@��'� 2C-�NGM`�LI&�Ԑ�ȓIن5�d�_����`pB��$�V��ȓ/?�gg�#����lǭsb��ȓ|��h�0	�*���h�(`����*�l\Ձ "%���r� wx� �ȓ#R���$�@3+X�ʒq�@\�ȓw^�L���1�t�y���Y{�-�ȓ'He��_.+5j4�vO:l8���b��m�AJ��w����G�=v��Ї�!� �Q.-|��f˂�.�`��oZ�x�R�0�S���4$����3&�|��hJf��@��3b�����c
H��!��g�\�3�#&F(���hf��"m�P��,C%��q̀D��Ig6	V$���������^؆ȓ7 ��xc!э64���Ϝ%�B���z��|(  �a���"�kܖj5�Q�ȓ]��h����~A��[ MP'��h�ȓ�lL���,c�h�;PM�YF���xy��	�!Qv=���^B:r��@��%�&��m�f�&�4Q��k�t���˓7��Q4M��r��ȓ�N��� RG,l�"h	��jI�ȓ)pz�������όR�P1��g�j���Ř
Fٰa��jZp�ȓ5:�5�Ce_	.��p��?zч�0� ��LŒvK�8�!�7[<���ȓ\��h:t�8p��͢r�X�� �ȓ{�,�h�bּa
�D�����%�b�r�C��H2���y|�����$hդ����ա���y�Ơ��S�? �D	N�%���! M�H8�AB�"OJt���L�A�'�M�&1��#�"O��2L�9  I֡�'"O�=�6A�5�dH�u�H9D
�Ъ�"O0�� #A�c,pA"�e¨[�0�*�"O�y��I�FG&L�5���UB��V"O�]��/�K�t�c��4�$�h$"O.	���C#)ux���
l�I�"O����$H�<Xc��%���{1"OD�qw�^"":��!� � �H阕"O,��i�6����Y�"���� "O2�ZPd%j>�չ"K�I����"O� ��葵P��(�@�K (���B"O�I�d� �����˽zc�8�"O"��`ʭIԁ��EJ�W8��'�^�ka�N�"����"$-cz]��'�\���i��Zcf�
k�o�K�'�nHx�.T�w�2���z�r�'�(〩�({��%�P�M��E��'� 1C���_�\3�K�J6�1�'R؈���qA����I��?8�:�'H��@�C� u�^�l]�h:���'����1��[-����[a$dz�'�hl3FׯRd�{%DA�O���b�'E�1��B� ����FS���'REX�+ P%~`Q�"I73p�b�'�T넉5�$�`3-�%0�@��'J����V�W"j|�C�(CAk
�'5�	�aF�7>p���F�N�ܨ��'���SD,ޒ�H��$�̀D�A��'�BȊs�	5$ЎF�&���'TA*�Ɂ$X�4�hƣԣ6���'w0����|?�!�������'��=�D��%:���3���Ƹ�'M�t�2U�^5�	! Oؿw��i��'6~�+��aa�Q���^uk��	�'45��.T�ܤ�pw��"@��L��'�j�I�H0��)���;���
�'a �����>^r)�c�18Wx	
�'��U[mՂ-y\�c AӮ: PY(	�'�*EZ�掻"hܹ�Y_FV�	�'k��c�MR�A��lZ�d�=I�� P	�'�`��ț Y��ҦNBI�v:�'�8"S�m��옶�M�G��'e�Bc�J�{�6�zv�D+Е��'
vɡ�H+ayvd�/ �4�z�
�'?�ԛ" 4djFX���Eф��	�'�F��Æ�M�p����R.}�	�'5x@7�܊sV��+cÝ�~�\��'�*��`�=l��3̓�D���'��x'�%fN� )���'C��#�'����	W:�5#���>8�X0��'/d��DFAxv�uA��2S�d2�'.F��! !u�	�$G(p@�	�'ެ	���
����O�q�r�i	�'r>h��U7,�x�5I�m`	�'Q�x���߲����
�X(x�'����h�*����UJ˩�M��'"u"q\�+*���ui@�x�`��'V<��"�/E�&��U�8e;���
�'��bI�.Vf���s'�X����'o���̚~��TT���H�'���E1pp�Q�T�Ē1��X��'�$��aa�1Kr0��c��	Ag0dX
��� H��/ء]��P�Lo\&8��"O�0�����aR,�Y8X)�"O�@�E�F�G������?���R�"Oҙ�#��nͨъC����y"O�t�` �0�h{���B���J@"ONe��Đi\�x�|i�"OؼB���56��Hc0�\���i�""O$������B�н�(U�d��!�Yk��=X��`�8�`u�ѯw�!�d��A��|��K�5z�D��@��%�!���z�ً�F�a��)��/N�!�8J��]�sHNOȬX/4�D�"O�y2��.�|ǅ��W-��1G"OWg�5H�\T��(�0!"ONq�0�I� t�vC�'"����"OX�΀�A�B9�T$-f"�=�%"O���g6�*�L� >E�"O�����"�&h�'�+p@LP"OdAӢl��0 ��P�#�h�~��f"O�-ivB�?	�����?��]ʑ"O�dhWd��CdM"S�^!j�IqQ"OX*q�٬���˲Ϙ�zg�(@�"O��[t����
W�/a.0	�"O��c��2g�`A0�P&
�R�[�"O��h'�	�h���`�����h��"O> Q��FkQ�P�g�t��\J�"Oz<Yf���.Isb&Q��Dp�"O�	��J'D�|B��&ȝ �"O�T�E
�g)Z�aD�j��"OTD��iڢ�R7�L&+�찳"O�=�6.�3[�Jڶ(`��=x�"O}���۽ns��37Ҿ���Y%"Oڽ�e�)E@��Ҥ�+ D�R"O�Dsp'C

�:Ux#Λ6O��9!2"O��gg
�:T���ZNz��a�"Oش�DM�3�2e�qk�=ex��"O��+deU>=��DS6��`���"O8���'H�2+��q�`I:�p˦"OF���dS8Q8�x� <0���t"O�}ؓ�Ay���qᡍ;d��c"O2<+ä܌Hs|!�Ca��tWN��0"ON�@��H����	�sL^-�g"Ot�c�k���[�FHl,�"O�3�O3C:�� ̏�.3����"O]�"�ҰiN��9ǁ@�e����"O`Q�q����f�A̰!�,��"O����hMt���L�q��A
r"O
8!э��Lr4C���n����e"OD���Ƴ?Lع[$�<H���R"O�Q�C[�0Ⱘ�ׯK!$���"O��;��������m=^��=x�"O����@Cc{@�
��^;q۠U�f"O(��DC�D�l��î�"	�����"O(�k�g��q�s�ݨ�M�"OșQ����5~���g��l���"O���_���]�K:H���1�"O�k$Β{�d`P��:Ƅ���"Or�"��f�N�
+ŌV�`Bg"O4�XF�+��y����<V���"O�u�% �$7�U˃�Z�1�X�3g"O�%�ˀ�:��M�6��ʐ�`"O��)+l�X,ʧ$O��"O�i���9	v�|J#�^
k��a:U"O�KgH����h��À=t���"O� �x��F�9S|�c���:<HM��"O��.A+�4���D�A��i%"O8�)�b�h�Jܘ�)ߚMk�ȉU"O�=���5j��5�rJ� hF�b"Onͪ�G�
\�d��ލ-?)b "O `jqN89
����� "TI�A"O,UA�N�I�b9j���>TSV"O>}!���k�D��D,h��)'"O�)f��T* CV�0X6|��"Oba҇,i�Vq�T�Z)[���e"O�P�	   ��   �  >  �  �  �*  �6  eB   N  �Y  �e  eq  �|  �  ��  $�  ˝  �  g�  ��  �  <�  ��  &�  ��  <�  ��  ��  :�  ��  ��  �  � j
 � n u! �( �. �7 |> gE �K �Q �U  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01�m�{�0Rda�#��i$��� NMӠNF�<(�������zVޙ@��	L���)��uv�8��� �	�"�Z?�!�d�2DT�З�J��93g�D�$�qO��'�?�p���ZD��+v� $�����=�騟�2��ӬCp�����k:�1�>O��C�)�x��a�W�	�	��
��NB��	�'���p���e,���T�L��M١�:}B�(�O�iR�F:+-��K��-9`�|�	q̓��U���T�o`�@�(÷k��ȓoδ�v�F|c*@�n�r ���?�ӓ@���[PfN86Rt�� �/$��}��ɭ�?馕����I.Ŕ�hD>�T���(-D��#��S��x!b΅3�F�і/+������}J~JE@�.+�Fm{��q�V1���R�<�0H��g���B�듽[ZR��'�FR�<i�#�?���5�7z�P���s�<1`�%JH��'���Iʖ.Qy�<9c�3}�\y�A+Q+G�f�PE�]����?���FE��Ă�a�)e�a(��Q�<�u#A����U��N0��;h@d�<�Ã	!=���A�g��-OTm�2kMd�<a�C�kE���¯ �`S�b�<y���8���sǮ~��%s�O�^�<��N١,�*!�_��X���PZ�<����}
B�+��6E�⬸�U�<���2@o����:W�VDVE!� J��źqoƨ5��@� �G�!+!��
�2���ŉ�����=1.!�dK�2z䱵��4��"	� 0'!�D�TӞ��D���C$BY(��!�č�u�L��䅮	�Ex7�:1�!��˫!Ɛ��#�6]Vj��L�	r!��DU]ph���>A�*�7!���6}�PI/�
7�5�R�Z�(!�$��E�x�f���g"l�P� $>$!�D��M��;S�юg�9�ӂ�>�!�4oBX�����l�Dx3�؂~?!���,ԃ5W�}�a���N10!�DP�g&��s��G/0
���b��x!�2GԆ`�w� �$z�����b!򄕊#������ ��XIүD(!��F��� ��R���	5�!���T|Q��P�*�jE*��W�!�D��l4aC��[�/���hB��!�!򄀑I�&�ؗ��V (�D�U0X�!�Ğ�3�b	��JI:(C4x䅘�N�!�d�+V�IS�F�\@:m�FC�L�!���(wp�j�N��E�a�qe���!�$6zĶ�k���~
p���"�!�䟃Um ��J�XGT�����I:!��+��ŋg-�=IFj$�`��/�!�@*����O��>Ľ��I��!�F0cUĵ�E��(OZ��:���/�!��)Q&1�զ
ih� �`��By!�DA�Xb�Å�id@xi�`gk!�$��vt��4H��0`V��"[�}�!�DU�z4:�ŏ��;��TC����^D!�F�W6�8��C�e I£]qE!��6x6ܐ&�V	!���hA!�P��޽Q�P	v&��R@��l=!��j����� X�l��4�C��Q#!��lkL�)��	Ґ�YԀ�?�!��K� �攚B��n�"YԢG!�%&^�	��ҳp��e)�$R!�� �)���]�Zy�]Y��Ɍ�M�c"O�Q:�(��t�����{�tuS�"Oh8���%q!�@#do�"_x
*"O(Y���X�7�`��ܗ-x=zS"O���B���2���H��v�']��'��'P��'�r�'��'SN�P2H�PTp@ �9E����'���'�'W��'"�'���'��l�`&Q2h@tYP��� ������'Y2�'���'���'�b�'r�'W��G��b��P!3��3&f�=��'��'�2�'��'�R�'l"�'���y�N�T���[ a )�|��'G��'���'�"�'���'�'IE�iU�U�0���윅=�����'���'��'���'��'"�'�Esi�qFȐ[2��+-֌�q�'�B�'���'0��'�R�''��'������{�F0x&KT@�`a�'72�'�R�'1"�'�B�'���'�`aQ⡌�d���j�$.:��p:�'-��'NB�'�2�'kB�'0��'��ʀN�7�,`�0�ȁ=Z�`��'���'�2�'U��'12�'�B�'R�|�`	۔H�@�C�P/�vIc��'wB�'o��'���'"�'r��'��hk7F��P����S�V}d��#�'|R�'
��'���'�r�'w��'r �F��e�Z1��T�t�j����'r�'d��'�b�'t*t�P�D�O����-/�����F�J@E��Ny��'8�)�3?q��i��`&�6����N�<,y�����N٦Q�?��<��Q�@Q�����$2�-\�y4����?b�>�M��Of�S��O?Q�cC�zD�#F�͈6t�!{�� �ȟ$�'X�>y����MY���(?rDh:�A��M�1��q̓��O�6=�` ۤnH�#f��S��%f����O��j�P֧�O�$�z��i��"!���a��ɇ�
`ĂG���|�x��A,z�=ͧ�?y�C65�.p�T$\&O��I#aL�<Y+O>�O~lnڷv�0c�P�Rm E�� pBU�+��쒢�LU�]�	ϟ �	�<��O.E�@�,C��-;q�K�z@� 򵛟��ɼD�� �K5��<E�K��|�V�K
|.z�qA��:e�����wyrW���)��<�쁽:�Q凃#k`��)�N�<!�i�ey�O9oZH��|'aD. t� �֏\4X�p�IW��<���?)�M��|X�4��$u>���'���9NS��tCRj7JY�"��:��|�,O䓟��J!���Hk֐pi��5S|dr��0ݴ!&\H�<Q�����z�<����L�:�f%����7f��?����y��$�'0"hY�t͒,K0��*�j@��Y-9V]Hs(�2��dÿ�bͱ���O�aL��Y���!nFJd{�k�6�<p�,L꟤�'�	j���M;b��<�qs�¬�O��Aad�[�<ɓ�i�O�9O����OB�$��m��4�&�X�5=&�t*LU3�1{�f�&�	�~�NI�I���i�?!��צ���ư�;�lM�ޕa��!��Ȋ5O��Ľ<	+O?�K��oÜ(�5�/%<l����4�I:�M�u��i~R�w�ГO���-ʊ*�]�!"[�����	m���'���';�RΛ63Ol��)�OT�C��,1&1h�]q��yc/ ��?YC2}r�>?ͧ���Oٸ�L�|2&%��iM9d��P
G?OOBXoZ0O�b�ЕO7�Hs+\�Gix��d�C�T���O���'[r�'��$&�i�Or-7(U;M,���iW��&���g�O�0z 
�����i��'�&�,�0*�:m�̀��]�p�&����Οh�IDy�Oy�ɗ�M��18/2����4q��V��2P��+O�kӠ㟨��O tl�31�z��ٴJ@��!8��� ۴�?��o��M�'(��A�g�&1����Öߖ��6)кێ���B*[��<1��?y���?���?	)�ȉaE
 V���#�� @zj�ȦA�6�qy��'��O=��|��@��u!��?�L%�%A�1��m��M�O>ͧ���Qe0�4�y"c(��u�P��9n���+�ybʟ	�����1��'��i>�	9��ܓ �[&;�>]#%�J�b�D��	��	���'��6m�!����O��DCA���K'	�Rg p�T�Cg0���O��o��MH>�B��>�4� �7��@�X�<���*�H��#T��'_�4�Ɵ#��'O�P�ɞ3�l��Å\�<�B�'���'�r�'}�>%�I:�t��pWw#0�R�柗?Hn��I��M��U��?��;���4�N���&®z��p	� V沙��1O��nڟ�M{�b���ߴ�y"�'�]#��?A�@�.����'�B�w��-+�%4�'��i>���şx�	۟�����ɉ�$��DEhp��[�vM�'2�7�� {�*���O��D,�9OJ�G/� rL����I�"�L��O�|}B�|��mZC�i>M��̟4C֎�ga���7Ɔ�R�R<ч�S!x)�yfe/?)�o@'X�J�$̞����D��`N�A�ĥ�V=b9�2�Vmz��?1���?�'��DӦ�Y�M��TB��0�����Ž09��ڰ�Jɟ$p۴��'���+b�� c�ZTn��$���?NS$t!U*ӓ|~A1h�Ԧ�̓#�Re�3��o/����y���u�C��� R|�J�s
2XS��+��i��2O��$�O����O<�$�O\�?eir�5	��	�DL	D�c��֟P�����4u�x5ϧ�?� �ip�'����A�2d��1�!�\�����l.�d�ƦA�޴�:�C��M��'�2N�*(+���\�����ļV� �.��h��|�^����쟼�	��\X�$�:���
 ���78Պ�Lȟ��	eyn~�@
���O"�D�Oz˧p�x|�j�4_��i���z%� �'���
&�`t�<�&���?Up1�Pav����ɓt� p�e-����SC
4�<�'U�BOΟ���|��� ������)�ҩ�g�\(W���' B�'���$^����4(���Qc ,KN�;rcY�F�`���d���?��j8���d�M}Ii�V��"���|�ʔ2�ĤM ��Q�'����4%=��۴�y��'��'��?	�R�T;�Ο;k�$�B�$b��s��m���'��'�b�'���'���:wO�-������n�� �Z]��bݴ��1I���?A����<٢��yGE@�T��C�L��U0�I! �g���i:�7�X~�i>�S�?#�+Gɦ��Xތd��*OR��c�����k�%A���O��#K>Q*O����O�0D _+��+jG?{�J]
-�O��D�O�Ĳ<���i�X� E�'�R�'�"���b�Y��;�#�(���a��DV}� l��=l��ē�B�Zw&�݌5�G�U�'�HQϓ�?q��]��X�P�W���$�L�{�R���B�-�*�*$%z���*�R�D�O����O��d$ڧ�?Y�ș�jȌ�$?+u&T��nJ��?id�i1u�W�'B�p��杲<zt�BdH����1�#ȏI&��;�M��iQ�7BM%&7mu���	�r!�����Oct�"�ҫ{�I�G�;jIV��K@�I{y�'�B�'���'7rl���1L�X`���V��Ux���[8?��ß�'?���e]��R�L�t=4q'�2Y��*�Ob�o��M�x�O���O�찠WJs?�`˱aS-C�Ч�B�"����_y��X�} d�	�{>�'�	:$F�Q̷ �,9 ���U��@�'�b�'�O@��M����?�F`(Gv��Q�{���a#�¥�?�0�i:�O1�'v7����];شeĘ)v��.�x8t�>�v�2E'
�M��'���(X����ۊ�'<���w��!�'ń��Ǎ�� ��5K�'���'���'���'��h���:8�� B'��S)�As�c�O���O��lZ�#x�ßx;ܴ�?�(O��F ��Tpb�
R�`s-�H�Ɂ�MA�iO�$iK��v=O&��AbhL��%����$ ɕŵ�?���9�D�<q���?���?A�@��_�B�*Ы��k�h УE+�?)������ߦ�:�c�ay��'
��Os�e�w�٭@��X���J����O6��'6m^���kN<�'�"�	�i�mwn���F���B���"0��#^�,x+O�	ñ�?���%�d�2g��}��_���|���3l����O����O���i�<9��i����,ש����_�m��!��B��,���'��7��O\�OJ��'6�ƤD�>Z*p��n��}���$B6��Ŧ�r�f�)��?�b��/2��Ц�������A���.��Ġ$�����<A��?���?���?�(��QCrFA�B���O�}��)�f���z��ȟ��I�D��B��'^�7=��icVDUV��`"U{~��zЮJ��)��4>[�����O2�4ˍ����?Oj�E��6�i�&@~U�E�F4O�0�#���?)W�0�D�<1��?����r�]ء X�_w$ј2&��?����?�����즭ֈP`yB�'	N�pc��9��<R�)�{o��)��'W�'��ʓ�?IڴH��'���p�nȸT:f���Į|�$]@�'��g�7*�:�z�J����	�?i� �'2��ɜ�z�ғ��q�����N#w2��矴������R�Or���S������.����Ε7~32�q��]H�e�<��i�O�8v�M�LG@�i�ꛏ��䦝��4Ta�恖7|������
SU0�T/ݭr�D�kDKڟpr�����bR��'�̕'���'F��'���'��`�ƛ=H�Fy�P�$E��T�V^�ߴr��-r-O��$3���Oj��PF��WH�/5�2� �얉m�����sӌ�&�b>�KrG�o�̘�j� W�2�`W�2�d��yy��]U�D�	�;��'W剣"��O�33�8H0��9�ܖ'�r�'��O��ɘ�M�5,���?�,� 2|<"u�ɦ5^ev�_��?�ճi��OPȔ']B�iw�7͙b�4�a��Y41T��1+͛f��d")o���7o�U�&����aL~b�;"2��0c�&����aB�w����?���?����?�����O����o�%eD@a4mZA{�qa��'���'�"7m��MT�}-�v�|"-�7p�`�sQ�B�J��OY�l�4Ox�l� �M+���d��4�y��'�2=y�W�t�:EB��I.�!룅��x��	"t��'��I����؟���<ddk��vI�%���c�&,�I��l�'z7m�������O��D䟔�)�NO�5	��R� ���J�$��	�����ON7-�S���I��wf������R�z�ȱc4Gzɹw��=.��,���<���<���8��5l,����$~I�"ʗK��p���?���?y�Ş����ݦAI��}v8%z� �į�Q�����,��4��'��0���*��cC�ǂ7��iQ$!+4f6����H�m�'���k�N��?Q$U�� �%�a♧C�B��U��81�9�5O���?y���?���?I����I1��x�T�֯a�-�3�I5_1<�lډK�H���� �Is��iڛ�w�r@�T�G�X誥��dC/g"��D=�Vig��Y'���?���t��mZ�<ɐ��i�6pB�A;��-H�<��o@�;���)����D�OB�$"D�
Dhd�b�@"��/޺���O��$�O^˓4S��τ& R��'�B��x�̕�$���*�~���[*h��O@]�'5�7M�����I<	�jџ^���ҡO"�$*��<��Π,�d��
�3!��m*����)�Rڜ!��M B'�!Z�.@!n�pS�.�Xa��'���'���ܟ�ぉ�.S�mx�Eב]i̭v"���#��(v�������4���ygAT��`�Y�����q�4�'��6M���=�ݴ��u��4�y��'�x����?͚�Ɉ�i�r�Z&iJ�@�z1��)קy��'��	��|�	�h�I���ɽV�*i��+C	%t�!�T2^���'q6-#)�����O��D$�9O4�J�G��v5J��3��ɗ�Pl}�q�Nq�	Q�)�S:?\&H
�(S�V8�hC��[	X+ ����U�`���'!`���ٟ$B��|�W��Y��	1�ۣ헆Y�(���ϔӟX������I֟��yy�&~��Y�u
�O�1D
�	$A;@M�,X���O��oZe��-�����Mk7�'A����B��i`
Sl^~�J�+�:��Y&�i=�ɮD��@��OX�'?���'.��b"�O�S�d��1	�Nh���	��x�I۟���� ���i�0�KSf��	�p��@@	��?y��?2�i@�%��ObOmӎ�O���"�0+�J �r��|�%�T�MO≇�M����o��M3�O���&�9;�ȥ5���9��v,�R�*���WC:�O,��?	���?��z��}���M�ȱ�d�����y���?	-O�nڻ*�<�	�h�	H�����	�����O�,�!�E�X"��X\}BNx�t�mZ����|��'18�)�O�.��q	���%,��iۂ���C��܊�I[��d�B���bM��OȠ��_�o��a�d܈�L�+$��O����O����O1�����e���p ��%+�<��Ȭx�4\�P�'���n��㟀��OT`l�%��q�$ɚx�8�r"e�5M��J���M+�늘�MS�O�UB�D����<�ѕ����OP�`��@�`��<�)O���O���O�D�OV�'.M��AMP0U����![m�)C�i�@�'v��'X�Ow�Bl��n�R�&�%�ǜmzD:�gC�S�v$m��?�K<�|�Ɵ��M[�'7,���� ��[sG[ot]a�'��pRmA����֓|r]���Iş��� � �:E[�aW1��(��Q�I֟���џ̗'6M (�����O���֣}��3��Q����G$`�x����O�o��M��x�-Ԉ��㯘�^z��]���$_13���{���;�������̖��`2� t���@�ڤ��,��B���D�O����O��$6�'�?��DFAb\��!��T̀��4��?�ƵiW����'���hӬ��<DԌ5�-� Tę �'7��I��M�2�i.6�ϜD&.6�:?I1  j�����6�	��<Č#��G,�2J>1*O����OT�D�O<�d�O�)��EG����Sѭ�3S���b4J�<��iE
��4�'�b�'R�O����qC½xR��5Qj�!	��43�:X��B��1&���?��Ӡ J��[#��=A� �h �.%���%��5�ؖ''������ԟ�cp�|�_�t	v���X�������C�Ɵ��I͟ ��͟�RyB�n�,$�3��O��h�Έ�R<��`� �6#�2�X%��O��o�y�%��I"�M�V�ibt6-6$�r� �XhJ�c�DKD�W�Ӏ�	͟� *��nG�'�Qy�O*���"�ܜQ됪+f:hB����yb�'�B�'/��'�r��;+˖Y!�C�e06)be��W
��OL���Y�Tnc>%�I��M{N>��#�cs�A�4䓊*l<�7#�]>�'u�6-�ͦ��Ә'���o��<���[=BD���
6(f!�E�<C lmb�T*q�d�������O��$�ON��E3 3b¡��s�jy�7Vg�:���O\�r�V�u��'��[>e ��ɐ ��p�s@�z���� ?2W��ڴL��vD(�4���M7��������y���*�ΕAe�41"�-�li��<��'f�B�d^<��`d�Pn�
J"�&�X�~
�����?����?��Ş��$�ȦY�U�Pa��Kd�U  ������1^
�	��Hzڴ��'��gg�6��NY�T�F�^+x{�)�s )��6m�ئ5^æ�͓�?�2�׷+�D�����K#|��0'J`�����L6�<Y���?q���?��?�*��tC4�q��QF�J��j��t��禕�ן@�I�0%?E����M�;�^푵�=~&V���5���!�i�>6_I�i>���?���]ަ�Γ$��);�#�6�H@�'��/H^�`Γ>"Yk�m�Ot��N>q*O����O�EpW�	i�R�S�M�:PA���O�d�O����<���i�j���'���'�Ι;%(�Vx���$���/$�@�\Gy��'�f�;��\�n1bĈ�#&Rp�Ĩ�'}9�D�O�`b$�5"�p"�´<��'Ӗ�D
�?)&c�+��$�JC�yB�7�ı�?q���?Q��?����Od��#k�!X��@A,� k?��`��OtoZ�F�M������ߴ���yw)�:�$���H�	��5��U��~r�i��6͘��0����?�䮄����]�? �u4L׺qYB����J�\x�0���<9���?����?���?��Ö�	�x�B��6L��B�(����$�զ��+��(����D%?-��*S"h����o}�4G�YB��H�O�loZ��MC�x�O~���O�jM�t�]�cgx¦��1���ÄZz5{7ʚIy"�u3`��I/kf�'0�	�#l�X�T+@/y� ��Wb�����ៜ�	ܟ��i>e�'$(�D�$qvr��9�d�ɂ�h�Xԑ原���w�&㟐�-OP���o�t��yG��&3Qz�P���[�1��/Pɦ��?��a�#�H�IY5�������3𾘚�Ȇd\���p��^���O�D�O����O*��+��*��y7�ޣT���@Ł�+hA-OJ�d�Ŧ=P��h>����M�J>yC��=;
n<��\�O� 9)Ìт5��'7���1_c�tn�<)��3�*�K��Կ	N�AG�K@����$�P�$�����$�O���O���E�5��Z�nW�l\�3ǜk�t���O^�Yp��
�Ot��'�"^>���ۛn�\`p���/Y��wc7?9X���	Ѧ��N>�S�?EY��U;k\\�v��&O�p��o֐U!X����h|h�'K���X՟�|��XHHE@ 	TCm�`� �����'}2�'r���O*���M{gd�ڄa��}8(��%J�S��\Y���?As�i��O���'�7��,	��F
�vZ���d�H�D���n3�M�$�W�M;�O�sV���rd��<q��<�
����8%�
�b���<�+O��$�O����O����O�ʧP���+'�H=�
Q�&*$�l���i��!���'�B�'���yr�z���,*�@�ň�$��'���S-��n�8�MsҒx���IZ�ZJ��3O�ŘV(�+�\,k��Ӊ?��K2O��!OƳ�?1��8��<1���?�7���l�k�c��B�;B�����?����?y(O�n�y�8�'���#^N.)�f�
)�X,�Ƃ� ��Ofm�'�(7͆�{I<�%cA7z8�RDk�P0�aZ@�p~҈־x�����i��Od����i�"GT�iqsb�L!ʶL���>d3��'W��'��s�=xb�� ���#@BֽwM���2e����ڴL��̢/O m�|�Ӽ��-$� t��Æ%?28k`��<AV�i�v6͎Ħ�j�����5�'q$x6A@�?A��)�V��ɡ}oh�C��&dT�N>�+O���O��$�OR�D�O��G�8OǌT"R͇�T�`Ѣ�<�p�iP�I��'IB�'C�OH2kC��n�B���*��TC��:,(����k��'����?-���kW�Ał��P�H�5 �	���Pr`�<)Z��A���O��M>Y+O�(s�R�/%伱�C�"k�\jo�O���O���O��<���'IL���r�|��D�oM�ip��9ɨ�+�"՛��d�v}ҊvӦ)oZ8�M����9ɚ���lK�	��sg!��\pɈ�4�y��'�,$�f!U�?M7W�����ߍ@�ۆw)��i���	R3|̹��f�h�I՟@��ןT��͟<�Җ�E=p/60*�C�e�Zy���?1���?���i���ʘO���s�>�O8X�K�md4鱤�]�]	Z0z�CE≃�M��i_�����0O�����k��yzB'F�
 �`�>T���@�&�&�?Y  "�D�<����?���?с���@8lp���xh3��+�?����$G��0�n���	����O�,�"���	Iȱ{��Ͽ~��܉�O��'��6�Ħi�I<�'�:P�O�M�:,�%	��$p��NA5��
���*W^���*Ol�ɜ�?I��#�E�n�܊����5�\Q�g'�����O��O��4����O�>+��N�5lT��B�'�N4\laB��E�4X�f�'v��eӈ�O�K}ic�X���Vs�@�DI��=K�tc��ZѦ���Wr��=Z��O(��%��4������J�a�8�2�$��~�^,)��m���'c��'a��'�bT��Sq� #&�;I�YA��'<�d�۴n�B P��?���䧨?	p��yÕ�q��H;7I�R��1ig�I�%PX7�ڟ�%�b>�3�*Цi͓U������]�j�˰�;R����l�Lq3�M�O��kO>-O��$�O�}��(C$Rd>͈4�޽�)$��Ov�$�O��d�<y3�i�&A�F�'���'�*�c!,P�12��ъ�3~��2�|B�'�z˓�?ߴ�?�,O�j�-�c�R5Ba���m�ȓ����j�� e�����)�S�d�"��؟��G��6-�%jd��X�p���ӟ<�	�4��ş�$?a��ş��	�yY�t�����铤�B�������M+�kZ�?9�g�&�'D�i>��8���k$酘�BЈ�'�Kޒ�����ش�?Q���3�MK�'b�#�(a� ,��\a#P�K��� �S-
XV�|_��Sޟ��������+ "
0|~\ t��3;C�	a �zy"�x�|�B �O����O����dR�P]�I�c��38�p��+̖Gv��'ݖ7�����J<�|R#�ɔ=I��R��:��q�œMǄ���$ʫ���Mv	k��'�V�Op�l=��3Q��7N��W���
��mA��?����?���|�+O����OZ��� \�r�"�aG�(�����
r�DE���?�%[���ަ�ܴ��(j�dx�T�1��T�����&�MK�OB%�������#6�	�� e(�c�*n�	��aU/V��@B?O����Oh���O���O��?�1�i^V%D��vą��eS1~����ON��D���:��o>Q�	�MsI>!�d��"xԈ��'>lj�]J��H�'�6-���S�-x�}lZz~�b��� Z�x���8MEn<c!��`52q���A�?!T�.�ġ<����?9���?9$J(n���u
F�?|��0�.ʖ�?����D��|� *�O^�d�O�˧8�h�1�ս j�͹��.����'���<���~�H &����?5�6Q�t���9���P�Nٚw�Rn�����c��D�'���Lԟh:�|�$�BҦsf��..��"OD��'��'4��$V�`�4��1�,@	�`X��KM� e��!�&T��?����F���o}BDm��aё��"�ךMX�(��P3>lmZ��MK@LX��M�O��b�˓�J��<	6��H"��S�Aw4�vR�<�/O��O���O&��O��'K�X��NK(𒀡#�3.	:ƴi�l %�'���'��lz�{��>�$�!A݃ �J�P��M�M۳�iI�P�b>9�a'B���/�0Je�F3y�,�J
l���V�D0�`�O��H>�.O�	�O��y#jS�CM��(F-؅1x�8��L�O�d�O��Ĩ<�v�i;D��'G"�'��};�lF-d�Tt���м!8!��d}�Df�Ȭl�ğ��'�����a^l᱕
N�xpy[�O��rsk��?��:��V��?��OD�d+S�?�B(3g�%U(n�Bj�O��O:���Ob�}2��O�"��b�	N��E����z�nh��)�6��' �7�:�i��" �D�\��M�R�A
�Eb��Rܴ���'^T�hq�i��ɗD����O�a2�cX�V&�(DG;jEaG#_f�I_y�O��'oR�'�R�lb$��=�ji�
�DA�'�M÷� ��?���?i��DE�#\��b1v!�d�	=˺��?�ݴ�?Q�O���O��G.A�p����H��u	⛦B^=3�J�����7F�d�J�.	ҒOlʓ{��p����#N�X%��-3f��L!��?I���?���|b.OrqnZ�/���Ʌ8����,}{ l�c�r�6X�I��M��J�>�շi��7-�ODĢ$�5
p\0M���֨,
�p��hn�6�՟4�d Y��B!?A����S�I��V��9�h�8��P�5��<a��?q���?����?���4l�9C����懎H/�	2�dվI���'qrgp�Z,�%9�Z��̦�%�T��d��5xd!�O�
}v��ڣi��\�'��7��ަ��	�j��qo��<q�H��H �j������L�'E�C�����<����4����O��dL�
/��*���)Zbx�S��f4��d�O�ʓp����!b�'�[>I��K�!�(h�͊�!�j�[�c/?�$X�lJ�495�&�'����W����ӥt)�y"\�q�uJ��
Y ����������c�	�%�l�0�،:|��"C�0t�~l��ޟ�������)��~y��m�VtСAQ9{�����7-gV��hȠ=�D�O�Mo�N�<��Ɉ�M;1�;~	0A��^7���t!؆#��6�'��@G�iV����"}�$�On�7p����X0<Pu͜sT����d�O|���O��D�O����|b2U���q�Â-Rh�2��B*Q��e�0l2�'"�)S���x����w�բ�)�KU� ���4B��F�'��)�W��lZ�<9�KL�?��s�薶D�P�27,��<���07�b�$֮�䓶�4���$��)�8��+�.(Z�BpED%�X�d�OX��Oʓ7L���̛���' r��0�lL�w��6�����n�f��O���'d6����e�N<�g�ZIߊdا	��[!zxg��t~2O(2ZZr�\2a��O{P)��5a���L+~�:�Q��2�$yqO�^B��'��'���Ɵ����h@-s	��ɾl���dKئ��IN�4����MÊ�w�T�U�2v���"�R���XB�'�v7��ئi��4�.�3�4�����np]��'�0i��TX�F��vO· ���ӥ-;��<���?Q���?��?���X
la�B�r������U ��@��|�Işh%?q�I<o�L�����?M�!��c��Sp����O��m�?)M<�|w��m���"�.ZB�9��(:ucF���H���Z�$��a�$餒O�˓[
�"�EM��[c��3e����?���?��|+O �m�0VǄ4��%S�<���(G�txS���][v�I(�M;��#�>�i�r��t�|Y��yV$㗃�iu�\�qC�'�|6� ?�sM֍SS>��߅��ݿ�'D�nȜ8��DJ&<��e��<���?	���?Q��?������5MT�{� ѭ�d��c����'��cӚ��1���D��M%��zOJ�X!�a d�A�!��&@��ēBA�Vh�O��fH�hƑ��z�GJ7Lu�% 4`өW�HI`F���<��'6�'��'��'Hr�'X�����>�&LK�G�q�ѣ�'��^�4Y�41�\T����?i����@	J$����9���`��Zv�ɤ����Ӧ�1�4Mo���)�=`�"	�2l�xY`@�o��y����VHH���@�d�<ͧ/f�$��|m8Ě�M&X�BD���P�4�`a��?!���?��Ş���˦51&����F}��;{m���QlEY� ��ן��ߴ��'��˓�M{fL�v�f��J�7UMl�Ƅ��Wd����ЅDlӔ��㟄����T��a�fy���W!��V+��m`RfiS,�y2R��	�Ißt��ʟ��O��H�)Ί)ud��Cу_s.�$x���2#��Oj���O��?�����+�]'V*�����3k�|<z�͘rK���`�n�%���?���b�Ao��<� ��q�� *�ʌ)DLOA�0�â>O��)ϙ�?ٔ(;�d�<����?�G���2D*�M-�20���?A���?����CӦ��p��Ey�'�� ��2?���0�2���;����w}҈{ӂ�mZ��ē�F�)��Ҋ)��=���n�q͓�?9�f9��A�&Z���������dM�d�%C�M��(��W`J����A�����Oj���O8�D-�'�?!d�Q�o,J�kC�I	Ck0۠L�#�?q�i�� QX�lH޴���ywFϋqTƴc �
#ĨHZ��G��yB�l�zEm��M㥭�6�M��'���"�t����q�$��$DZ�\�ȀcW����Y�D�|rP�T�	۟`�Iʟx�����2W�x���=f�	�,��n˓���	g�R�'���D�'�X���m�0S�E���*h$���Sg�>iA�i�7��P�i>��S�?�uJ��RV��bㄹg�E²C�=@")eF�Hyb	ˈ�=��b�'���5E36Q��F�7��mS,��:X���Iӟ��I��4�i>��'�P7�ï
u��DZ;~�rK4�W�9��Y��7"5�DE���?�e\����4dݛ��}�$Dk&��%�l@'
�?��e����iA�7m~���ɭ,��1��O�y�'��t�w�\Z#��
Q�y13(��l}��'s��'���'9b�'.�t!`"�Vfx�`cj�'R��e��O+x�n�$E���A��ny2�g�^�O���b!@�ex��x�OT�Ol��[���J≸�M[���:P��MS�O���fa�H���I��џq�p��%�;f�����3鈓O�ʓ�?��?���H߶��6�F%a֌g �K��Tr��?�+O��n��
�4�Iݟ��	d���#mТ�Q�e�;g�`ʔ]����a}��}��n6���|���]��!"��Dma�[�A^%K0@aS]�{C��f�������A�=��OU�lތi�\�S'��~�҄�1l�O����O����O1���k�&�Z�fA�A[?O~�����_�H�%�'�v���T��Od�n�;R�S�O�@�R�#Eޮ�Z]�شq���\5^K�6���K7nUB���D�~y��O_�1�v�Lڡ1���7�y�U�X�	ğ���џ\�	ß(�O��	� ̧ L
��恄���F�y�4����O����Ov��������]=^���)F.��m�az����������M�|J~��ǀ��Mۛ'd�"$+� a�\�'��=��و�'�"iƠ�Ɵ��#�|�P����П|�C�R�/������/*�h�lɟX���t�IYy"�j�<)[F+�O����O�Ȃ�P16�C�ʞ
P�ce�,�	�����=���&J�ICfۊnzT�@�Y#�0 �'��(�TH �>]�B�����Ɵ`���'��Hb1�]3L�=h$f�..�b�'�b�'{R�'��>���{l�IE	��n�V�[�}u�l����M�G���?��j��&�4���˳ B�\Ft!#=�r4O��n��M;�0�0��4�y��'�`�1���?�Y�)�2����+]tN��Z��U$��'J�i>�	Ꞔ��ş��	7SZ��P�BW�1^U	�L�/_n�'�6�ǟD�x���O^�d(��+^Ⱥ(�ANO!:8H�k'A��T�$Ę-O���}��&?��?y�I�o�h �/�R�����U)�r�*4,R�� R0�d��O�A	H>!,O��r��ʅx�m��jM�o����K�O��d�O����O�)�<���i����E�'*���ޜL�0Uل�	�s�����'��7�8�	��Ӧi��4�?���lH�@wG_�[�i���5g�bИ�4�y��'�"D��E�?��O��I���4*��]�VmL<*���\cv�t1O��D�O,���O��$�O~�?�	��֩�ʥZ"�O2A#�HrG��ߟ��I�|�45pʔͧ�?�A�i��'��H
�F �3KԞ�%;�'a���M'�i�)ȹ6B��6O��dCuӺh��$^��-0�,�,[`t�5oO&�?)E*>�į<�'�?����?Y���)Q��(�	�,|�
|p�hƶ�?�����D���VgADy2�'��ӘvBѱF�Fw$tpv��i����	3�M��'����O�F����̰S�K�;U6�˥I3m#BU&:�r�/O���[�?��o5�d�#^��Y:����(�D\�s�ޫ(�:�d�O����O���	�<yǼi����ӧ�1btNuYĜ�Uǎh!��=R�'��7�9�I���_����T#���)�0�|��H� �MC�/-Œ�4�yB�' x�Ç�C�?�k�O�I�rB,YU��u��,x^�|��5O�˓�?q��?I��?�������<�D��.T���:�fP*dX��nZ�'�ҍ�'�����'L7=�$5Q��j��R1@�/h�x��NӦ�ߴ�?�-O�)�b�$��F.�7���Ó䁜?b2��u�	�/�R�C`Jz���Cå^�R)E|��dy�O����6��-�&��� l�4]��'�"�'��I��M����$�Ov�ڒ�)qjD����١PY�5hV,7�I���O�7�O�ʓ^��1:��S�D�E�2�
�K<��̓�?	f�.1�:�#I~B�O{d��	�2��J�V0;C��!�DL@�5;��',��'r��sމ��ڸwj�$��n��Z�Cb����jݴp�\�j��?�s�i��O�\��ipԑ3��� sa_��Dm�lm�ڟ���j�禹��?a�C��l^�	ԿC�B䨧��b@��D�#E �2L>�,O�I�OX��O���O�I�$|�ޡq�m< ��tˀc���D[禁Y���Ɵ��	��(&?��	�)�� �B�V�}0��% Y-d��O��oZ�M��\�O��d�'��C� ���V ��g�h��%L�<�\�aMb�ɗ'n�����'�(@&���'����E�b��� �U�Pxh0�'���')2���T[��Y޴%�0�p�r�1�+atU�V)E�(��9����]@}B�f�Ԁ�������W"�@7�Ǉ#.-��
^-MeBIo��<I��v0N�C�g���);+O�����(��NH)�����d�0h�=O���O��$�Od���O��?I03��s7����i7�H�'.�ş|��ɟ�h�4i1B!�'�?�E�i+�'��U���B_^I�2Ȅ-x���/?�d ɦI@�4�Zuɘ��M[�'�o_�-�b�HPa^�n�^h��Iķ{?z)���ϟ��6�|�Z�����`�I矔xRn�5� 䋗,�ujҙ�����D�Iwy"�z�L2���O��d�O��'3���S�oх�$ R#�_�7md��'���'o�f��O�O�	�t��1�
�kؘ�3)�106H�5��XVH��*_�d��˓��q��O��L>�b�Q</�- G*���4�C��3�?����?���?�|�+OnZOkd�`�_��ၤ?N�Ԣbb�ɟ��ɺ�M�B�>��ip���gϘ�U[�W�ޞQA����i��o���m�l~���/UE�5���Q�� P�
�0u�U\��ǉS�v	��Ky"�'l��'c��'/�S>A�H�.}�<���U+t��Q�[�ME	F���O���X���˦�]�5�z%�­��W�,����πvd�A۴P���5����0h7md���2��S��EP���l,"����d�L8i^R#h��Cy�')$��V�L:3U/%hQ��D�	`��'c��'��	>�M�&��?Q��?�����/��$����7_�X��߼��'^��o���q�l�&���J�Kȴ�w,���I�Ш<?Q���x<2�R!�=��v8*����?	GC�s,�2��
12��Ġ�(�8�?9���?!���?	����O��Pw�0���V`ؘ ܘ�-�O@�m�v� ��۟�!ٴ���y�ʞT�����u�
}pp`���yb�iӲ�n3�M��*��M��O�:� ����
+�l��%^9�����w�O��?���?a���?���o��	Y!i	�a�>(hSH	N:v��/O.�nZ�'WJ|������	q���,aFƓ�y͠��6&�5��(to����O�6́a����	��ԧ��u퉦pH5�"C\�|1�AH��$�}�ՠ��-mn�O�˓F_8��'-��Ū�H&oef����?I���?9��|R-O�<oZVp�$��%9A�X��O��*��g,Ѕ�ZT�	��'�X�Igy��.}�	ܦq9��L�A609Ѕ��|�����̗�?��oZ�<��w���*"��%�r`2*O��)��\%�G\���P�f�-<y�9O��d�O��D�O��D�O\�?W[2K����#�v<�E1�+_�L]��'1��w�>�Ї)�<)e�ih�Y�l�Ì�~�Z{ ��F� AY���&��c���JeӲ���r��6-u����'>D�9iD�8���è,/֬�2��R�b�AX��Ey�'���'C�ݦN��m�P� �R��I�b �A��'V剔�M�E'�?���?q(�h8�rc�,f��yCJ��lq�="��H(+O���O`�O���O/�5jd�к1vӤ�> D�=C�A\�F����,\�E"�I�?�
`�'��%�x���㺉 e�U�ѭ�2���'��'"��$V�(ߴ�t!��
TWaVaz�
ߎsL�)� _���d�覍�?!�Z�xش
q�-�"5�L� H
>�pH� ��ܦ�B�4z�cߴ�yR�'�������?�W����OM�1W�σt�:EzeMq�@�'"�'!2�')��'���=������`q�M��MR��ٴb�zD���?����'�?	@��yg ��9�y3`�Zuܶ��e�<+��6M��P'����?M���R���o��<I�Dþ0&zP%��4	FBd(BI��<)c�[�&��E�����Ol�D��.]�Ԯ��]����Գ"����Oj���O�~����>PZ��'�bG�*�
����ͻչ�l���JN}�p�p`�Im��L�����,.\2ԵI׌Љ;���^�t�s�nĨ}w��K~���Oё��_x���@�P&��b  �)y~j9k���?����?��h��Ό�s�.i7g4B�<�:$	�������MʐlVgy��aӆ�杹9�p��T�u,�ɧ莍sͶ�	��M���iq�7�ɦ(�N6�-?��O���)�d�:P��N|,Ś��Y�x�luIL>�+O���O��d�O��D�O��y���=!��b�J4W �Qů�<�v�i�4�p�'���'���y���SB��4
�GC��C�!ݭe��ʓ�?qߴ�ɧ�'&��e�`�J�{�NG@��Hp�-4ZDX,O���C��?�a%8��<a �^�M3� 2���5ZxI�s�æ�?����?q��?ͧ��DƦ���E�P�2F?ri��퇼m�k�bΟpܴ��'��iٛf��O&6P�|S��baǴ	L�:g5~*)�g$e��z��8�D����X�K~��B��1{Uh��CY")��E�B���t��]���XU��ql̬�U��.V���k��_aR��G�VѢ���"^�fH�L�Xe��  B[�;~	;��'�e�Q@ɗ|�q�g0B��㬙�y��)�{P�C�ȼ*���x�I�ݲA��6"��j��]s�Dl��`C�R<��p"݃{9z$���۞wL>��4@�3�m�V!B90��=�gQ7lH�!ڍg
��3�ޔcdn�p�K
)�j����G�� �ɜT�<"޴�?a��?�Q�߇>ǱO��ĭ��;�KI%}��l@�F�%�l���tӌ��O����(�:�&>���˟��	.�� tis׆�=dC��bg�)b�p÷i����[~��'j�꧰?qK>y�Ƌ�:YN�"�V�H�"ٛ�o�Be�	�r����&!?��?���?)��n�2�U�9���ϮCjqB�0�?������Od�OH���O2e��V�A�Y����d/Yss��h�(�ß�p�����������Ɉ-�	��%�d�X ��A�L��wJҨ_�8p
�4����Of�Ol���O���f�'M��.��J�D{�'�w�z�Q�a["����O��O���O��ɢ|j�'B�p���:>����Ô,�qߴ�?!I>���?�P*��#��'� ���@����Eר,l�x��xӘ���O��D�O�)���|���?A�'e����6:�)��K�O�Ȱ��x�'=2��&X]��y��n�{&��7���@ L'�p]R��i���'�e
��'���'k��OH"��5IF9����`�� \���Ɉ<�M#���?1.��C����<�~r�Z�H��V)U�V�xy��ݦ�0$	��M���?�����b��Vx��1IW'.���`�+��m��n�#<����'O�s�E�*��D��Ǉ�fҥyEn�����O���=N0��'��	ݟ��Y�V��B�w�����$/����>I!̛>���?!���?QE�ބae6+��
�A�E�&�'] T��.�>y)O���9���ꀨb�B�r�E0e�G:s��rtZ���A*�h�Iٟ��I����'-�}b(�{����@G1�r��ϑ�I����OԒOt���O�Y�"�Ջ(Fb)!�3�54肯D]ܼHM>����?Q���Ğ')��x�'\�}b��-D����%`VN�YmwyB�'��'�R�'Z���@�'#�ldDCh� ; F	"n�� b��y��'K"�'#�0>�(ʨ�N��Fζ�Jt���qU�<���^n��m�֟<&�t��֟�*S*�Q�mC�A�@Fе�jy�,l���@��HyB�Bl��'�?���"�K 5r�H�AH
]��D��,@�	��'���'u�9�3�'��Ի�O �Ӯ)�p��Vf�ޔ(��{D
6��<$� ����'�B�'x����>��cS�a3���T���$O��\C��o�����*fT-�I�8X���OWzP��g@7VL�s`B�N��@��4N(|@ֶi���'�B�O ����\j���j��X��t�O�TA�D��Aq��Z�b!��y���?I�+�Eb]�v���x����כ��'��'�j�/n���ty��'��d/q�E���K5�X�MѱO�4���3�D�O��d�O�ı����o�%�!F�h� �o�٦��	�,8��+�O�ʓ�?�N>��:���x����u^��1R�Ϸc5�	�'���x��'�@�P�'���'@X���A�о^�=d�9+��A�gݨ���O���?�H>����?�A�=jb��"�DI6)��K('bH��N>��?a����$C�L�ͧ��L�&H["7��*����Bd�'���'=�'��I�5���i�A"BѼ<޸��d����C�O����O&��<YC�W�C��OD���[�l�B��`�����:r��'P�'�剑%E$P��z�INH/�iC�G
7���z@��-����'K�V�#0�ħ�?���C⤚�v�"U	*"fp�;�Sp�Ijy��H��b���ٟ����^-��9�T�B(C�Čs�i��I\v@!1ߴT���֟D����$\��!�v��v)QСj��w���[�H8u��ş�L|zO~nZ�o� UaO7� ��g�.xH6-�8,"r���O���O�	�<�O� �H�M��9@���i�	`�(#�g�6��2�ׇi�1O?=�sM�3:%n��S�\^p`���$�M��?��y���,O��l�d!|�̘�4
:������{����<g��*Y����Ĥ�Ps��m����Qy:ց3DDgӰ�D���x�/:��\�+����}(��өP(QܮP��T����+#1z�b����hy��'�PPtOE���}b���-.�|�3��E��П��	X���?	�l�|	Y��c/nQp0Ĝ�nQa�`Y:ò��<a�����OڈP�e�?�j!�^�Xʮ���,ѿ����~�P���O�����┩F@�7m�B)�]�BN��ar8r��Q&2���՟�������'�2��".��P�R9p!v��� /(�qq��
P7P�oZ��|�Iey��'�����ҕ~z�B	���(	f�Z�n�
0(�I��M�I˟\�'� �A!j!���O��ƌ�e
K	�B`x2dd�
e3��x�T��9�R�l$?��V`�a�c뾨x�(ܺbx�	n�jy��$EN�7�OD�D�O���z}Zw�6�B`��Iu�B�ƕ�j���0޴�?	��5N�y��?�-O~�>ar�*�����a �P��q �Dk�����Jئ���� �I�?��O>�JY"M��!	bxe�A�U+V��Y9#�i�p�'0�Z������ꠘ1f�cE�F@҉>���Ѹi��'�R�sQ��X��'���O�9	��a OX!^�=@S�i���'����/Ѧ�yʟl�)�O���\ -Z*����/�:aΛ<w�Hlş�ڵfU����<����$�Ok��U(��i���$���3�h�����a�H��������l��\��'CXض�C�`U���Y���𡎃m�<ꓜ�d�O���?���?Ѷ��	R��pC�d"����Ywt ��?���?A��?I+O�YB�C�|� F��0F�����h�����i����'���'��#��y҈O$�Z�`�3Fy2	A0L:7��O��O���<�	R�H���ß4j�"�tP\4*�-[)4+V���L��M����D�O����OP�Hs��x��'b򕲷MY�/U0�k�@	n&�,n����Ify��Ԅ1L��?Y���JWJ�Gjxʔ�R->R8V��rX��O0���O��dN�wt�|Γ����Y$�f���-2��!�KN��M�*O�,�v�ᦽ�	ԟ ���?� �O��Ս]ET!�$�
#�R8
�(�wW���'���%�y��|R�I�>i�`�0!ܿ{��ԘG�yH�6 ���7-�O��D�O��t}2U��{�E����єw�D!��M�׎��<�����)�Sß8@`,O�+n�x�Q����$q�͚��M��?)��`A]��V�x�'���O~5j6�%L�$\cI�p�y�T�i���'�4e���yʟ��i�O��� >2;'/i�T�q����S��mƟD���4���<�����$�Okl��.@<!h��)x�}hfDz�&��7X��s�'��	�?)��ܟ�'�jdG&܏;b�����©Ffp���B�q�����$�O��?9��?Q���
)��cG�
L�����)A ���'�b�'���'���%bL��OL��H�+{.:}J �O6��r�4����O�˓�?q���?i�#��<�G�A'Hf��t�� �4� ���'�R�']�R���7.^���)�Ok�'K�\�1�P�N��y	��J�T��v�'%�	П�����P��~���j?�e���vR|���K�ȀU����=�	ǟ0�'��;A��~"���?a�'n�ިjfm��~�v��_%$�y�R���	���	/t�
�N�	S�b��4}j5�5nϦ8BZ-0G	�Ϧ]�'�h� a�z���Oh�D��-ԧu�-��Fi�W��K#KS[B�`m�Пl�I�_[H�	��9O��>�b�cM�*�4��%��BA�&��6��0T�dn�ߟ�������S&��D�<1�F�|򺙫�IU,\ !*ubş|����Æ�y��'��~���?�%o)jd� S#R<#������ٟ<���'hr�'� .[���Xyr�'�� �5h���A �>7�ep�A�7>���|2�ݲ�yʟ����O��D�->0�iV�}�^y0���>�m�ǟ��@�ҕ����<Q����Ok��..,�!�(k��2��Gm�I�?����qyB�'�Ҙ�T+ {��a��ƞ�/;�U�Y� �g��>�)Op���<���?��R.�ꡊ	jT$$R�����������<���?���?1���$�C�r��'  �Qy���	�|9*aA@Z4^�nZuy��'�i�oZٟx��|�l�i�@'[�sA�4����4ӐCt���D�OP�D�OpʓM��A��R?��ɝl@�K���/(�j���i��,u�h�4�?a-O���O���k���O���#Ul=�VN�H"-�M������OH��<Q1@�*/L�O���O��8"���Z̙ �	_�+��!�d �$�O��6|��$+�ĩ?U�&�֫ֲ��t�	�I�a��qӦ�a1�I��i��?���"�I�:gĕ�'1�X�V*_�<n�6��O��W�e�H�D-�8�S�|Q���EgK*0y�_8"7�D�6��l�۟h�	ϟ��S/�ē�?�bH���d��$�Q�֌%�E����ƭ���y��|��)�OVp*���|Z ���B�2bv� �ۦ��I��X�Ɋ*h&�k�}��'��A�i:d۵��"T�i�*�<f��f�|2��j�\�����O��ӢRmx�) �^�89�%��g(�6��Od�����g쓩?�J>��Rg"��Y8H%, ���0ZNx�'�T)��'@�	�(��ן�'�|U S�'�쉣� ͚%��֟0�xc���	c�	ɟ��I.�t���@
�
)��Ax�:%�p�ԕ'��'�BW���"����D��(+Z\	��B�+��������D�O ��=�d�O��J3����Z�?P^��cV�c��3�VK��'���'�2V� ��*�+��'W�|�y�#0t�Ĩ1plR�R.��z��i���|��'��)��yB�>�H-.ո$[�?�~1���ؖ`#���'��W������ħ�?9�'@-�AR��4$����˄�!g�J0�x��'B!ͭ�y|�П�!��!��֍�}[��J��i��I�����ڴO���П��Ӱ��d�R����D�t���[6��F�'����Q��|B���	L�%Y��p�DP�+�oR����*$\�6��O����O���P�L2!CTA-"%&�)a� ���iV�ۂ�'��'��,�dUe!�,R��ș*�t*b�ʿI�mП����"I.�ē�?���~Re��8zzEk��R�,��x�g�(�M�M>��		�QB�O�b�'�r+��{<�h{p�5�p�+�,�	?jz6��O^	��ƻ<q�S?9��s�I&�\:FJ
Zޥ0���RV��J�O�8��Z&��	�t�I����'GPlp� �}O��3h�*(�"Q�&.�W��O`�D�O���)�	�\GB�co�#`oB���H�=�PŠ��$�I�T�I�8�I̟`�w�L⡂I���rL!^cWCA��!�'��|��'�Bk���D��4l7h��Wݱ9���1�D�	���'��'B\�@
�Ԏ�ħ[�>A�EJ1tzm@�	=D���i�"�|"�'��*��'A���v-�l~x9z�D��i�4�?��������h'>��I�?��� ���HC,�4�A�1��`��x��'�]�O��޽ ��>,�H���^��YK��y�9+�b�'?�@�+_�I�0��D�*&v�!)U*D��8��1β1y�!���ʸ�6��%�$��o˾�x�J�8Vy�;EGǙu>�	X�oM��\]���H�EX,���� w�"��A�]�甸�f�/����)XU�0ϋ`
X�Q��[��0��V�������9y�Oɧ�� ؔO�D���h�� �"�k�s���!+�8i0���O����O�Ȯ��?��_d0aS-�=��Pp�!��ZA����'�Q��+�P}����B_F{�� �tSj̱Q@��+�(�#�	���!l0�I^�Q<l���hO�t�&� �b�e��E���O��d�'���uyB� N���i\ hPQ:���9�yrM_9P�)�]�CǊ�af�)(
"=�'�?�*Od�#d�ަ)r�����<�E@*YԀ2gj�柈�	����	�=[&,��ܟ �'+6<��PcF99B}�ba�&t��y���=Z��DZ$��wF�{�r��#ǩW+W�Ș�cP�U���C*�iq�Lz��єNYma�jr���I؟�2�z밌��E�� �� ��f�g�'�џh�Q�S]��dDưo�����5O �=Y�JЋD�ɻ�䝐fJ���&a��<���i�B]���Ԧ���)�O�˧x����+8p�6�V�T��)Ȑ���?����?�u-�82qX�	�/E�p�F��򩕴����I�\bF|� OY"Q���f�X�4�(��m�lb���IlC��2��X�ip�!˗I�+s���/O:Q����O��2�Ӌ!�R�{0�L�BS�؛!	�pCJ�z��=������C+�MP�H�w��v����=�� @��aùV)��:V�����
]>�m�ڟP��R�4O�z��'��N,R�2mP�J��S�8��I
z�Nx���^�H	q#C�K}*�^c>�D
:o�0���Jʏ$�����g���(���zdI������O�< "��<l��,2`ᑨy�ΩJ�d�#��d�Oz�S�Sb�I��n���Ed.4�C�(-bB䉆i	&	���V�G�ʴ(�&�'}p,"<	S�i>m��=t� t���R)5�P�'X%j8�4�Iß�I��uˀu������I؟p�_w���'�r�3�!R�n�ȣ��ٔi ���VK$U��uG��gN��Ef[������i:�D&��aޥ�
�ʒ��5�ӿwڹH!� hh�!�ޟў��g&��kY@@sG��/
��I����X���O��D'�$�O��D�<)�� 
O�ʕB��;�lX�Үz�<q�Eݰ�B��@1�t3�,ǸH`�����⟀�'�� bf�s�0,�fE�j���:�Hc��xC$@�O����O��D�?<�D�O~擑V���������c�Κ�xF�Qie/F�$��(�tf2�O4L�`B�h�8�#��V�%Z�$�|WR� S�S�m��!M{X�����O$��V!^� ��#�@1)R�P�7�X�OD�$�Op���r�1@��/HZ�7%�8;1�����M
������|��_��IJ���O�r����K�A_Bm)�O�<(�<��'�"�ga	 ��l�t��5����'Q��c�X�Z0�uy$d�>=8��'��1��-5*вd4���H�'����HK�9(p!�Ħ�.5<1�'���JP��:R���pd�/>`��'���Z&�J〱��������'��]��ܟq8���v=�� �'��T��G�74�����l(!��'��$��I�A��sূl�,���'GT���BӪ$e0�b�Ԅa[]��' ���0���h�	XX��H�'�^� �խv��QD/	Q^����'�>�#wF�\FX����>M�z}�'� \�GAln��/��F5ڌ��'Р���Z�B[HEI���>dp�'�H�t�B����NE�1�\x��'���3U�U2\J١��,,i�
�'��hbȡBf%!S�)��h
�'@ ��#��rގIWjK/
��ٲ	�'�r`�g���<�M�uE4��'��RD�I}�(��5t���3�'2�Q
�����Qkөm� Ua�'��p�V��TA��O��I����� �4�w �>��E��·}^Y�"O^�b����>����1�z��`��"O�u ���5���0y��UH�"O��0�f��FBƍ���(��"O�u�7���RQ�M�5F؃r��y"O=y�j�0��}�5/͗ZS�1Y�"OP�� *�6w��H����O8>� �"O��Y��!mjT#���~��1�'"O�]:�"�Vxa@7�r���a%"O ����ˇHpN�b�뗽D�Ҹ "O&��,�+=�P]#���P���g"Od�Ui[�G�$�	)��Dӈq"O8����>r �I��!�1P"O�j�P&6���(��R���"�"O@�#�e�o�T�bh��v���g"O�!��璾i�4e��{����"O�t���$�P=p�J�d�l�"OiX��@��i�6���p�$�@"O����K��,a'��';�!�"O���!Ad����$�7�*�9�"OҐI�A$q�fT���t��XA "O�h�B����P0N��X��S"O|I�A,Vd���"őv��"O��1U�B��lP�S��$�(K4"O���CL��>�i�E ƅK8�!ir"O��� �	4�p���L,���"O4���J�7X:u�N�(-T]�U"O�ِ2`��lb��dҷ�j��@"O) �e�*?�݃�Y ��P"O�	ֈ��7J h�� F�u4��"O���j�8x�x��%M�aj@!W"O&pI��I�+/ź!dC�t\���"O�!0�)C�d,Ő�bL��J"O-@�D�-
��X�W��)��r�"O���A��*]�Y��ÝA� �q"O� ��F5��=�� �R��Q#�"ObU�-Pj.$s��3�H��"O���O�<u��k�z��E���O��Kg��n�S�O���ˀ
����*e*غFƶ�y�'�N�� �I�1�x@eb�09�DHH�t� ��$�p=y��ݞ��MY@آ�~��&�}��(���r{�	�c�"Z�f}�����:^�)"Or�nTxB�@�a��X+*���I3D�V����
�<4lgk�"(�
�j˵27!��]	9:
Ы�-Re1s� D)|��_�h���>E��E�k+�ƚt�۳�]5+�B�ɀ7���b١Hw~e	$����'��܊� )\O.�	֧ԝ@�� hS�i��1��'�J|Z��N�|��E#�	��M��u��чȓ>���b	?[�މ�����@��5�D�ZQ@F�(�8����H�V�!�ȓq
�y���*D�@�r2��9�� ��,�
�TDɇ�):W™&W `��V��z��9�zRr�5�v}�ȓY�bPy&��}�|�GjX�"F���'�܌����-�EB���M~�Յ�|�t8��DC��X� ��8Ԛt�ȓT���JR��1~�xr�\rW���r�t*��ȀVi����E�"�f���4?��K����9dV���!���y�ȓ,�t� �*\�褕(��g>p��D��eHN[�ɰx9f�[>	ҤK>qV�I����/Bx|��'+)D�Г�m��<8�,�-,y���?��Ɂ'ł�����K^�g�'��UaD���U��CцI:t-l��>�l�ծa�? LeC��9(�)z�FY�XҒ��5�U5l��ò�'��1�*O�p�r���wʆ�+��D6"
B�`�,WFJ�[a�?�c#NU�#�⩠P!ܟ\�2$�9D�T�t�Բz�BA�C��?q����#w���(=��݃��޸\0b����2����O�/�䰇/�a�!�$C-z����1��0`�T�%(N�k�"��w>O�,��&N7[��T���?#<y��"�K�AI!-�b�AQ��a���hC��9D5H��gF�>�d�s
�!���0�B9}nD���M'�O��y�gP�;�����/خP�D���ɝ1��,���6��%��
<��%7�ĸ��&V%]�v����g�<iC	?^�8�'�T E��"1�Y�<!a����X%�- -�����ӥS�ļ ���Bk �r@I�62C�ɉ7_���q&P�=(���"$�pT�8s�k����/J2 K�E/FxcՇfdF)P@��5�(Đ1#\��0?ّ�J0�.��Q�j��U���pi� ��G/nɊ���GK�B=0��򤗛L'��@�`�&<X�	&�Y0��2�� ��7���l�艓��1H��A�Ј�x�`e�'�@�*�O��:������j �БiXV�X�1O�A{��Ψ8=�eԋa1����i͹%���Z�#�"�pa��&J���ťG�R!�d���ƈIJ�@�ѽֱ��:OX��d�E D��x7l�X&1O �{10�z�
 
�&DL>�!c�3P���r�'�P|�SKD"�n��.
9�����������O?)�ӏy��W)_�r�Ћ�2 r)����S�
i�������� @!����B[#	���*��-��7K��@��&K��t�'�8X)�:�O2��dM
�h��JZ;�p�����i7���6�qO�#Nt�DjS�� 
P�+�Z(\^��@$C䉔"u�@�Ċ]��L�֋�,Ac�L�҃�l��lPn��O���|V�9��BS�$7��څ��M�'���؁���<��c�4��՞;�YѰiJ�6K�>*Vd��b��Y�4aSk�f(%��}
�C7E�n�ҡA��kL�"��� ��qQ�ݘ��M��h�5A���>v0ŦC,q Peb!.��b�-C&��|�\�?�KG;{�,[��P�Y��`���J��dɪ�~b��O*���N��?1l�����#9�|��seΆFR2�S�/��\Ȼԉ^�f�?ɤG	�x�~�q%�BZ�x�D��@#����ԽioV$@��R2c�`�3^�R��ɪDHp]Hb$�+��<�3"����|br��0�F4�!`\"o��Q���C�ɘ�ލ��A�G���i�x	�>	r����D�)"o5zj��\�`�
ْI���Q���>?9�)�x�䌠B'S���ܢ��Z$i�����=��Y0�K>� �"J���'ٱO*�X l�?�����~aE�)~�	�_����q�@��K�$_�Q�,Rk+=��%�
�)v�4����'�v�>�6��/�F���IiJ�q��[�8�T�_F�����I^��Q����#E���$M��� F>{�hH��.݅;<�G{"KۯMh��І�"�M{��R�]��h��U:V�`�`�j^�y�+>O�p���|9H�'����J>a1	�"����ץ"Hy��ޘ��7-�U�:T9R@<6-כ:��eاfO�J��i"%�7;�剛!�re�4 �v .)�`ـV����$GV?uAd�	�1����>9ԋ�	[�i����t�� BG�C=�ܓ���Z��I#�m�tE9����`�#���X[��@�1
ND@w�>Yf�4�0<Au�	�b���$Mի��pP���{Z��`'ܪRT�>��'U_��m���X�"=�d[�#��ؓ'xH��D�/ Ϟ�#�X�h�A��6>.u1��#S�`hI<�f
�Ǧ��jH�@؁���E��lm�c!Ԍ.b\��)�x1Gy�?Sll�g)Ĭn�\��	��JD:�o�?,�`H�`�A��U#Eр#z�����T�?c�S�M23ـ�F�h���ea�>qc��&L��D���@K��>	ǮBN瞬�㎌m�~A6mHp�	9sZ����'�.-2�l�4�"|J��)[ ͫ�����O����C�}�I�`Nռ����M�T;P�W�b��� �G�2<~�@CŐ��S>e[S!�Y�>���
?���6�7��Ip�~%eЏ,�*�%#ʇ=��|Q��/��mҀF^>Z+��rŮ��<q%�M���I>E�%V�T�H��'Ts�b�c��іE�b�I�I�H�B�2�$�<�}�È˃m� $��CQ'F������i������e��9�0<U���Z���҉?1��ɓ�ϷI �E�hA(��ˎ�|y�}� ��!\]1O���:�R�X�,�<"0]9"���4O���O�k��c�naTOL
$z�s�M�H9���a �F|�L�#�`�G�$�ԥ[���A0��_�����*[���u>����E�2����p�;�(���"'�M	�Ti�Z�v��"O� �X1��Ҁg�(I"Iʄl4����5s�,zr�<�BˀI���'���0f�-c�Q9�
�'��Y�(	�	�jɈ`ݢn�h�� ��~�A�d���Hf�,�
�O�j}� Жah
P�$��z��-��	�mC��VAXux�Y��'�x��(
U\�p�2j��tQ�'4d X�D�N.hS��;1�T��K<Ѣj�6⢨����,@k:�}:Q�)4E� ��4#B� ���P�<�t��<�.Q"b�� q�`!�UƋ��� �O��@���7����{\��UbѴ
���UM����t��y#2�A���c�G	`���Ǎbc���]&�MȖ"˻U}��d��5 9���g�-�BFޛ	G��A��3�\����0�r��
n!Z���Ԧx&-�ȓ�$x!�*_�{@��k�-E���ȓR����/�(lr���#��32��ͅ�JO��4AS%&����i:G��C�IxȀ*t	*~���G��B�	�l::���Ib�6��IW��B䉺K��ٸ�ʏ�zN��"'*�TB�	($_D�á���R!={-�%"O��) ��<�\�b
aI�=�w"OLq� �տ_\0x��K�1D��"O����<t�z��"��W1��"O�9"��H��z�Ȁ�C'|,��"O"(�k����y��g���� "ON5�Tm&d�>���$_n�@�t"O�L �DĈ����� ��j"O�y1�iJ���X���W�~�Hx#s"O�y8�û-�&ݐE!T8ը�0�"O�p#e�P"TM�&�����"O����#gl|x�'��mO��P�"O����q a˂��V <��"Or�u.�z�����"a�E&"Ov\��<h�t��McN��R"Or%��D�*}"A�l�0Wi~=c"O��
VH�$.Y0@��(`>0C�"Od�Ъ��q��k"埒FAnp��"O8]y&JKD@�]�!E���"O4K���/;� t�ך{�x�p@"ON9Z�(�%$�|���@G=s���"O�,bӅU�$@���A�%���Ї"O����
yv=h��A6����"O�X˳N!�T9�C�@=�x��c"OZ�*d
�3�tP	`M�	�r��"OR�B��L j���L^Xj��"O�����#bi��P��M�!�"O^��*
<q{�r�ɍ5V@���"Ot)�@΁�crF[���T�:\�q"O��[3 �_����'U�7f~�h1"O�xB�ia����q��~�R̋�"O4i�Ѭ�"hʔ��d���k�"O����R (������9�ڌR5"O���d$:*��K��6\N�Yx"OR��e	>W��SsH �AU�� "O�9鐎).��1�f��7V��E"O@X�/��m���0h\�_ �"O���s�L-�R�3��	���a"O:�H���#�򈉳!\�\�Ґ�"O"YA��,V��J�o��n���s"OqX�.�d��9@��m�� v"O҅RTŀ�^�&-�v,��:��w"O~3���-�=��J�f��$sS"O��hD醳PxY�A�tpm��"O�D�Sb�V�ڹ9���72�4@"O� ��p��A�la>�V��Oj�k"O�-q�mȻ(|���[��"i("O�p0ӮM4Z�Z�{v˝�+���ٱ"O6��EF�/1�pu���[�Q��4��"Od�0u��Xu��&��(h̀���"O�5��Z5;f"A�s�՜n�8Q�"O@=@S%J�8�4�0viP�w=�@"O�عW�2tF����K�o�8"O�lj�	F��l��M;�0���"O��F��$d��� Y�z����"O�%����&�&\YVE\[	��Js"OB�H֢����]3#��o�0���"OnH.w��*�c^5����"OB��"+H2q����f�A�6s��r"O��w�X�"RLx���=E�H$b "O�z�J���4����� IX5"O0��0͉e~,�&��e�FTq"O �Ȱ��:.TT�N��s���"O|�$i¯�h��'�V�=��"O���b�6���q��C�4�� "O���%N�<u��J�������G"O�B+o:��򗄙�r�Bp�P"O8��C�<����✨L��c7�#�S��yrN�,��"�_=Z���Q�fI��y���Б����Me>���N��yN@1)��"��ъQLRi��Jܑ�y��A�{��ȃ0B�Ok��bgL;�yrG�"�\cV�D�M�\Xc�FG��y�W	�ʀ�V��e	��@�y�h-_#��ig`#Q���HpgӁ�y��=B+�88נ�6��Rǉ���ydE�0`�C�2E,�`yAd��yr&C���H���!JKBy��fC��Py�~W-+kD 0���:Y��ѵ"OZ��c��a�t��.�/�(ur"O���*J������
A�] �xy�"O��Z@�� u�����n�r��CA"O�l2���)P�P�0fSd�HE"O�t��A�i% feV�fhX��y҆�:N�[f��;L�0�A5�y�	�o�-$'�74`t �΍�yrČ�c1��
3)D�h3����y��::(t2��(p�B��y�bP�S8���3�� +�\Ju)��yr���l`��B� �:u�'g�9�y"	�t����&����B�nL��y��ށM�J%���0�pb�nO��yBgB�8�b��45���%��3�yR�� ]������5d<a��L��y�*��H�2�s�^-4DX���
�y2̄!����HQ*-�vA�0m��y2����D�ų3�0�����y2%��)C(�A�.�='u5�u딭�yB�԰b���V� �P������y�c��|I�[ ��X�90����y�H�Q
ZMp#�N-�lY0A�A�yrj�	ĊUB�O]�>�2`h@��yR�Vg�R�R�G��[F<��!�6�y�!+W����A߶L.P}hv΁��y�H"hݨ�AoU�B��4��G�"<Q
�z�~ �Տ·aC�aå�%v�LQ�ȓeƦH	��3�~ �[�$X|�ȓ?�h����R��T�G�ߞj�̑��#���8%�Ӈ�����ǝ ����S�? �E��`S�g���ŮH�oe ���"O���� ,|d0�-�������"OX8��a�MnL��Q ㆌ{U"OX��SI[�T�䁛doE5K�A�2"Oz�Ф[�2�~��n�1 (i��"O����)�)l�F}��hTN�x�"O,�J ��m`�f�"���W"O�9s�Bfq�M����<��k�"Oҹ�ᗄph@��ph�2b�ܸ�D"O$ؚ�J�3q02,��˵K�Z\!%"O���L];U���\�9t�4��3�Ş	�&@�%e��$��pc ��1�h���`0�L�a�X�h��Sh���<��G����"��8h}ބQ1k��X���ȓW�y8��\�, 9��H�E`\�ȓw�8A� 5��(�" �1Q��hR9�`�Jz�0p@wn�a��H�'�ў"|�N������H��GGH:'!�d����F�աR� �c��  !�d�G���M�_zA�U��P�!�ĕ�n�JUH�E�5~��h+T� [!�d
|�X	3���h��(�Ӡ�H!��ڕ�bqQ�/�;�>����<*B!�!>�i�lؤ3�P�$T&y:!�;ubB�	�JWV��	T��hL!�$�*�ʔE�#2Q���S�Y�bE!��W�p�v��a��mH2�����9'3!�d	�x�
}`OM����3oGA�!��3�"��%Ժ4�����͍k�!���R���^u]R���N@�C�!��@.Ou��1�%0�%"E"Z��<��'�� �!��f	`����N$�uq�'�H,rs!�B����@E*��'M���Ū���dL�o\m��;�'�t��^�x�T���)Z�.�F,��'�.�Vg�=E��3qk�0��s�'�Z�	+ӗB������7�iA�'JJe	�������V2�N\��'ĨRbC5~�tT:��;V�@�(�'����"�S"��	*˘� ����'w�L@� ��+���.z�6Ĉ	�'��-yf��M�&�C�q�ҭ��'��rc�,ٹ�"R�eU@!��'��YDGۺ%���3��.ʚ���'X$,�ƒ=��8S�.�Ȉ�'ɆՓ�d��6� ��B�W�s=d���'w��"`�}P��ы߹j����'>Jh�k�h*˓�0`�,Y
�'�����H�F1�3CD-#�*�+
�'�)��J�;Z��L#bj�5!����'��`H�-�����A� e�|�
�'�~���K=sL�dS�f˔.��|�	�'u�E�l�1/-�I�P@R'y�l�	�'�.�n��91��Z�_�J��]�	�'��!��c�c��!h��
�<|��'Jў"~�� Q��|z�`	�T�̨��ld�<Y��)pkl�&��c
Ѐ�R��J��t8��QW��)	��Z�l��2�\�(�m!D�����O�6q[�+��Z�l8@�B!D�xRB͓PQu���!d(dy�<D�p�sA+H:Ry+� �W"4�k��7D�r�i��)P�8�Ċ'8l��5D��* -��7�@�&�ʞ=�h�A�4D��gdL�$�4�ۢ��6D�� ��YC��(u��	p�ײI<MJ�"OԱh�
`>�j�@ƺ��v"Oش�EC [jx���X�K�
�# "O����O(}�f��� ��D�v"O�`�p�dU���F��x�꠳�"OR�ЂBn�D����5%O���q"O��rd��~��9��閃75��s�"O$���AЂ�vc��/��r"O|��H֕+���〪j&��Pg"O��a1&�����θ�v�;�"O�K�Mɘ~:8��tG��"��l��"OF�A�K��<�b�Զ�����"O�q{3,K�ʨD2R ��t�̸�"O��PԤɂ�8YC��f�> �"Oz|9��-@2@0�''#��4��"O�ţ��1A=�=bǇ�h���"OĬB�d��O����&Y�l��"O��h�%��p�zM*]��aѧ"O��G녡8��%rc�δ]���)0"OV@P)^�5��3
̟^��Cv"O��� ��$A�ꬹ��<\��X$"O���v�L�z^r�����o���£"ON��/�D�x�*e
�/z �z�"O��p��A}�Pv	A,X ܈�"O@ș�OH��t�I!5P����"On�8B r%Cņ��Q^��R"O�����3qנt��03Z.��1"ON�I� \��ec�&wr�"O�a��k�7D��zf�Y�C*��V"O4H�f��:�mA�n� vS�m�Q"O(�ҁ ~[�09��*IA>�p�"ON4��Eo���.�
�Ș7#D���Q��78.��Ӂ�/^3�śq�&D�ЫeK�;sɲ�R2怞wVJL�T�&D�t���!>YʰX@gR-h��C.%D��t!�c��H�+�= 4�a�8D�t�5@X3!m�(�¬�~� ��!D��hs�Ut�H�� #�����J>D�����F��!� �l��x�$�<D�hS�ϖ�ȑX!�'j��ⶤ7D�\�#
�����Ō�f���`5D� b�@�����S�()��Æ5T�V�O��*T��.���!vWh�<�R�iNIj� V�2�̨)���O�<�A͜�a�4� ���P`�Qa���I�<�qė= B������\��D�Da�<��C�Z��r�n�3i ^!	3M�`�<��oG0t}�U�CД@�Hq�vi�P�<�H�M ����iQrB�l3�!TW�<���X�$�t�S�C�v�D�
��X{�<���4&��,;db����&�]v�<�B�+��t��&�5��%� �u�<)�#D;?���)I�22	�E��\�<q��
�A�܆IH�t��g�M�<��e˰L�<E��Q�2ɩ�m�M�<9A��+֖P��@�����TL�<y���)��Af�՘K�����'�K�<٤P�K{��S���U�ĀįGE�<QpJG0� C�L]��9��~�<�C��EQBԋ2W�8�°�s�<� iI`pTKp��Lh�l2�r�<)6͇���'
Tg���Iq�o�<�g�
�F��Y���9��(	A��u�<� �6^�����`ˌOi3�J�<� �Ź$�0(c�`�ˇ�5�8|YP"Oj�q¨]q���2b鐹֖�"O<�D�&ڮh�q蟣���"O�HA�ʖ��~}%�4�>��"O�P�� ��~j�g�`r��)"O�����#.H��kG�U	T�jH"Oș��`�&�.9S�b�<��P��"O�y	B-th$R�a�}9��`"O�;�@���
6Ɓ%�V��5"Oj��PM���ur�CQ�`�"Od J�+u�(��Ъb�UsT"O$\B�CI;b�e�&aO�S\U�g"O��7c�|�)�����y��%��"Oɓ0��:m��A� ��e���"O�m{�!��LPx}��Z����B�"O�v�L���3Pu�QR"OĀ��IϹ}�\�Y�$�	\;L�&"O:���[��������<Rv"O�z0�L
r�$s���.[P(�S�"Ox`��P ڑzd�K.���B"Or4����(7� 10�MD�(�q�f"O����m�1[^�����^T��"O�[�	�#*�0���[V-�d"O�=�"h��9x}����]����q"ODJ�O�?���)@m��hJ>��"O
�`�M�+}�ꭰ�,�� J�Āu"OĸҢ���(|�E�3� ->L�)�*O�3� 4�)�Pg�+)����'�&}�j��|z��K|���'��h�@����8�G̏:E�vs�']��_>M�bQz���?��5��'m:y[K��L>�E��
,3�ĭY�'C8͋��)c�ٜ)T��'����Oћf߈U��9&i����'�Nd �6an��r&ƚ9�1`	�'�l�h���P93r������'8�EZ��֭lҞk���)Q�x+
�'VR@�u_����po2P3 m�	�'��8z��?��y�A�\Tp��'��h �� QƲ4�l�<S�]0�'��c�;��[�YO	� B�'�j�;��$S��q��/�4H����'�8Aѐ���Z�F����:��0��'������)]N2y�ǀ�a<��'
dp�vH��ex��3 ʰ��Q��'�d�j�c�Bm��3�.Ԍ��'���8!�݁��X��&Y/�H��'�(��ve�8(�k&���Q�l܉�'�p�G�U���Չ�%Q����'Ϟ ���YS5H��LQIPP�r�'�
� �
�y�H��ė3-�(��'@��C��6r��#���2��c�'�D�I��ڂ&�|��WE�./?���
�'zz��6f�T�0��Y�.w敒�'.���� 6u�H; ���o@���'!��p�F8.�>���*T�fŜy
�'~T�0 o�m�$���E�b�0ez
�'j(4a�4s.�H��S�/����'I``���3n���3�]�#븬P�'	p��sH����ȕ��0OK�� �'(��Q��p�؁��LD��
�'5�D�q���|�c����x�@	
�'��{��P�f���CԊ�� E����'�z�1�����j�F!�8!���� Vt�c�;_�T�@C@"wK@1p"O�O����B�� �ș�"Ỏ�K�(6=X���95����"O8�d��jx`h��ؠi���3s"O(yHCO�/T��#��!C� YC"OpXK�D̠D:�2��N�$dau"O:l�O� W��!HCQ�Ig"Od̋@�_�"��{���<Fp�r"O
��Ae��A��a�E�RL�L3e"OP����	���T(�GT(*�"O�R��=�E9��,�j�"O��[�4W��&1C���0�"O2a3�2�����]�w=��rf"O����-��m5��2b�!�]K�"O򙠢��+NΖaBկ�����"O@,�Va�lC�U���D5-TH)�"OZ�@w�L&��DHũ3� � �"O��a��_�0�N[4I-'t�{�"O��h�c�Q����d8r�"O
|3���&�R��U�� ��%�"O�ذ�ׁw1�E`Á�k@�<� "O`@��#4�D}��!Y�}0̽˳"O"0['
"a8l�#Bwn%X�"O Y��ÖF,x��� ȴ�"Of����M�\�ɂ#E*+�R܂p"O�$sK?v"Fc��|:�1"O�3���n��fG]Rs����"O��j�a\
JK���Ui��X�0 �"OR4�u�M/;��᱁TB@՛�"O���OM$S=2�H�X�x̢l86"ONp�^=&�����
3�p��"On�avN����� "�n��"O�*�	�T&\���&V�nq�"O�%{���*�	�� ��Li��"Obd��А�
��υ���h�"OD���Ҷ8�Bh��� 5<�̪�"O����Q�5s��#U#S~���T"Oll���Ъ#b]��̚jD��4"O�b�Mgй*�.�9��"O�l�'�5E���b.�
6��t��'�1O�A�T���zL ��@-v �#"OD`��>����M?~ Py�"Ov�a�������bh> �$��2oI!�DQ���0�bG�J���S��@!��2at⁫� ?V��E�V�P@!�D�3Ы��!_9410Ǌ��y!�K#K�΍JĪE�d'�|�P�A� M�{��$P+04XȂ��-ii�H��L��7�!�W�|�a�iHzh&� ӥ�"/�!�ϙt�$�R�G*� I��

�!��*i��
����?6a3S��(!�$����t��%e�%h�Er�!�d�7̺�n���$�s��T@�"O`�	B�B&���[bʗ>^i����'���
���6`�]:@�G8��K��'D��Y�@OS��`A��aP�@�b�*D���bK�z��Q��)�P�Ԉ�gk$D�����ρ\V ���n��jB�#D�8���'�2͓v�
t����B�"D��f)Z�|�0A�,��<"�
?D�xr�����$r�b.°Ģ�	"|O�c��
g-_�r���O!+\� O?D�|���1B_��h!���cr+)D�l1�`Z�l�L`)�!�
]f �xe;D�� �H8go�������%��Y#"O �h撙F��D��5��eA�"Ov��v�Q.p�+�J̄_MF(C"O�RlO�c2F���.^:JP̂�'�	 hQ��!��M"V>ܹX�+���B�9'Y�m��ۣfʉʶ�Ds��C�	�3��HK�N[nЈ� w&æ&�B�I�C����ض !z9�b�E9uTB�Ɇ8X�p����e��H�㞽�|B䉐C���{��֔�c�[�.C�I"��ڐ
��8�h O�QG�C�I6R�F�3.��;6 �S�G�1��OF���U#=�b�o�46pm�G�H�!�Dؼ(Y��P&�5z��P�oTe�!��pU����.&�~��b.߀#�!�Y�,�%[0U��M��KB�L�!��&�x=C��pΙP�L�"�'%�Hc�PBn��i,F���p�'��	��!ךL�Q��=:�`��'}�M��iI��Q�`��* ��}z(O��=E�NʲlE��b؆{ �Whǐ�y��ד;�~p+�ϒ$" Q�����y�C��OW�\b�
��'�c�`���y�M=_�����J��0���^��y�c�u�Fr�k� �;����yA����=���юL��H���+�y2�˟,� }����u���#��8P�	ϟH��a�IV�'��gP:�P�s�M��:m�	�'��q;P�ܱA�L�������'�.�6	���0(E�(]�
�'�@P(�mE�]pXxs4iӴ;Z��	�'cΔ�b/D?�@t�Ķ[�xH	�'��	�(Nu�ec�bqb��'���g"̚i@6�p�gݛE[:�r��?�N>Q/Op#<i�  d��A�+��x��J�<��A�p'�K2�?��!�a/�����q�S�O�Z� �ᏎH2΍�Rhƺ#�F��T"O2$SM�f�ʍ˕�9�a��M7D��ʲ�W>J����L�I?�e���?D����U��4m��*sZ�]@ph?D�PKX�"�~�����t�Q�%M�<��
Į�p#�lD�8B��k��a��I�23�
ݗ5�2-�/�O޼�	����?E�$LPX��<Q3��3K�(YҮ)%�!��3�T�ZB�ɺ;]`�1�͗#U�!��&W�\\��瓪N�p���� �!�ēr �`��"��"u��7v�!���T�J`P�Ͼh� ���#\m�!�d��x�^��$ʁ�������$�!�Dǣ��)9��/'�ε���M��)�'S�n��5��pߴ�S�%A72�ڬ��'� ���@�8,y��H�zH��z�'��U��K� Wh��YW��<��0K�'K���Q;~�2�[�_�3=|��'ڐ�+/������H(P�8�'?��bT�'����F�N�
���	�'�����0D1pI8V�U#�F��'�9Y�b6
{ZX�Dc�tB��
�'���A��J)s�������qB �	�'��%�{����㊐�h�x ���'��:E"�>�ʭ�S�ȺP8vT"�'Jv�s!��j��}q"eǏt���c�'�޼;��C&U ��؂��r6&��'��(e@-qVʁ�FW�t�6%	��� ��b֛QAҴ�bۍS>�"O�j��t��QrL�(F�邱"O��2���/� y�2KŜ&4�i��"O�E�@��0u�X %�� ���g"O�D��͈W����Dب)k���V"O(xiƆD�iU����cF�Y��"O�@��(ħ7;v�r��Z $K�yѲ�D�O&����,"s��B@�_�&��L9f��=f!�D��S�A!�"p�Py4�9%\!�ĕ5���B�Z#'��}�&���>!�Jht��$��r9�} e#P*H!���8'���$�E�P)�5c�e!�Dʄg|I�5#_Iv��!�;BN!�ќ��0���[�Sc�X��BֲR��'��'�a��`A��J���X�w��@�e�2��'az"k@�R�=h��	|b���-͋�yb D�ِA��KYuݸ}�M��yr�[ZpQ� �	ss�� �I���y���47��#܈gc��k�	�ybE��I�$`
'�=`�A��ڗ�y���Դ)űPk��҃�F�����?�N>���h�.@r7��S���q��F,��҆9��:�O�ѡ��7K7�[#��,�D�CW"O��s�8a"X�q��Ի2���y�"O`9����i	��i�j�s�4p;"O:(2��R�s'�
fq��K�"O�E���K��|��ʔ�&��a�!"O0�:� Բ~������^�AkJ8p�\��%96���ܑ����#��<��LxF-�w��7z/R�pB̉�q�d���N&x{�V�,^���ņ�8��ȓM�8�uGN�z�������( }�ȓj�t�F��o�<���fL�Fr���9
TA��BˣA�:�惔SY�ȓu�iG.���]����>/E��J2��0�ʘc�J�Pg�;gEb����	�u�a������
��,ܜC�ɎZ�������D�҇�7�|C��/�@mH֩3������GJdC�	'4~L)*S�ѽ6��hh�%1&C��[�@5��M�Į�@�w��B䉱7� }����Y�8��dы��B�	=�Xi���p6V�Ѧf[�Z�B�Ii`daB2��30��x���Jf�C�<P�.cj��~�f��S�(Le��Ē�9g�qU̗!ZS:̢��[6!�#B����i�(h�tkZ�3!���=~�P�,�,�x+'��*�!�d�g+Ȇ�4
�(ɂɞ���	D�����  �!�����A$m��[R�,D�����78�(%!�NK i�H�j6D����F�'TJ��%FȞ9��='�3D�\���>{�����c.�Y*�*04�X��N0~��ě��D0=[��a�<�W&߸-?l�qK'o��<"Te�_�<�"�Ɓv��5�FV$'G$�I�@�w�<1qc�05_�`�U��`�.H+(	m�<���J���F�>e��X�q��M�<�1��Ǝ����6H �C!GL�<1f.وn*RI���г%:�����Hh<	$	R.N��l�͎&	�A0A�<��x2�͆U�V�Bң� ���S�!�;+;�1�Q`�?J�<aB�,�!�D��4�b6�+X�� �=�!�� L�s"!+mf\x�!���(���{7"O����H�I*�DO�rR8$��"O�z'Ś�$���ßG� ��O�Y��cND��&� ��&��W�����<�5�G.[�p͐)I�iҖj���D?�8��H����j�*x���g>D��s*J*��E;À�N���t�)D������"X��D��/�Q���(D�T�A�նY<쌉@S%��C�M%D��J�R��=#`n�?K�\fO&D��x�@w��RŊ��x`�P�*?���O���>��H� �,�t�H!D2PN>ړ�0|��P�;�h����T ��k��t�<��6D��=	(׉�jlk��z�<!R�ڙ�hi���;�Ȣ3(Z^�<�pbD�}r��q�Dػd��aJ��a�<)�K��x*F1�m^�\n��7Aa�<��C��R��EG�4���E��UyRW��$��|�珃�k���V�2&���Y�(�VyrY���	s>	z���v����?4��;�,D�\�H����Ms�"9���4W5RC��4+�2���n�y���6���K�HC�/���c��}0�Ё%�sW�C�	�#���ÀFAP���!�45�B��4�Z;��	�!������*B�ɩS}�hs�q�¡��b��v�x���8p	�@'Q|&�9��[39��ȓw�z���-رH� ��D��U�>L��{�,���P��{rAÅHR�X��l���5,ǯ�V�;���5j(�ȓA���r4��c�Z��'��Z�"��P-2����2��-� ʣ�ZD�ȓq�x����>���jp
!\�1��$�� Ō��7%����o"X�����| ��K�v��e��[�4t��ȓ\�z�ٰ+P�
T:�3���vu�ȓY!x����o2Q�fk ��lŇ���  �I�.��9���5Fd��A�`|	�fD?!W��L� �:��ȓ9_���(Ϗ5iJE�3�*m�M�ȓ@�رdo�)BB�r4��ȓ���R��W��NИy�a�ȓj�$�t�ҥ�.I1��D\�مȓep����[� Ӡ���b�o�\��ȓ+��	anX�AE"����Ȇe�Ѝ��I�<A��߳
��L���F=3F��8e�\e�<�jA� 6����V�0gfm(E��_�<Q�e�;�%�deډj2������W�<�`I�b�J8���ZWJ-�OAP�	S���Orް�G���l	!��S�s�iC	�'"�q��;Jdc���8M�xr�'Ɔ�"a�)
��1�Y���\+�'��q���3b�\�R6��_1�ńȓ:��K!/�"345ڰ��sV�͆ȓe���4+@1�třp
�=H�Ɇ�eg>ѱ�NE1���PfY�2W�ԆȓjT�֏��{����&�-Gl�h��#�
]R�f:
_ �pRi��sO��ȓd�E��F1�.��pÀ�7��x�ȓE� ����?.���K*p���ȓE�Su(N�>��@Q������ȓ"y��3��1�`a�S%T:'Y���ȓ+ĠMB���*,��,��VB���`3�U�0�[�=�L@��ɰ[p�l��S�? �<˳��S���K��{�h(K��'U�$(>}>�)aG��B� Y�4N�&m�{��$�;|KLx�H�V�V��!m�"Q.!��+ ]�H(P���^�r(PЬߟ3)!򤖤1v��[�,�0��؃Ҭ�8�!��8W�5�3� ~4Y���#�!�d�]�s�n�+u*�"����{�!�.z��e�P�*5��4�����!�����I>O�M���[T��01�Iٟ�IŞ[``9��L9��py�� ٞ	��	R�'D��thHl��xJ�+Ё)��N>�r�Ҡ[�)Y�p��P�ajPm�	��Ѕ�	����q�B��jj������18C�	\ �I�c
_4V���L�&/C�ɏ&�Zղ� V�Nٙ��ҏb.B�I�B@�V��oX"���-t�&���!?a#�k�$536��T#Τ�c�ux���'�fp{�刬}��)	�%)� �����hO?�`���*x-t(j�eH�I�fIŤ�pyR�'ʶ ��DG�^�ft%@J�M�HQ�
�'�����l�T�yt�Z36��R
�'�������K@���SL̤x 9a�'���Y& ��XsLR��D#� �8�'bJY(�F�'?�%��O�Q��'��:2��@�RS�A����?��y�OR
w�h '��:&��qp.��?��0?A��^�G�Ԉc&Dgp h��XU�<�Sd���x��G� �jٻ� FG�<i!�ѥP/X<��_2�XiAΐ{�<�v).�^=�pBΗSH8��k�z�<9�-��]��5��-�-sנ�q��X���O��T"$���]36�Jb瘿Z��l ���'>� �L7 fء��ZQ���'�|���O�u0i9DJT�M�F%�
�'�Pp�%�D=@**���6J0<���'"d��GJ�� ��7B��+,�@�'Fu`�o�?Y6z�Zddȵ(����'�6t����=�!h�Tv��(Oh�=E��ENZB��uD�5^L�Q���$��>���y��g���r)Г]�Te�#��y�A�n�.A�U�\�S�؀B�͟�y�̜>�	��,0w��f����y�[U�JdB�c:W�ƴ@e��(�y�^��V�1�#%NV�#����y"�E.���#�� ��P��%&���)�S�O��2�bE�t+�ɶ�F�1	�'�,��J".��#!��4x�eZ�'��쀕�˚�0e��ލ@T]�
�'Z�	dK�\6��`��e�‪�'�
�1�QllIk��\��H�
�'�
��`
������؀Y�QQ	�'�L`�iQ�k���
R��`�p�'#,��T�J��j�KI�4	f@���?A��?�����i�ODb��	�H��8 �\��B<��X���>D�0P�.ޣw���2,^��#ĥ2D��8�7K�Hԑ2=�/D�`�em���X�QE@-E�F�C�F+D��0�_�-�� �� �R���a.D�0a@3E���ؤu�����.+D��ȡ/��.`8��X	K�<���OP��O��$�O\�'�?��yR�99�y�hǹt������O9�y� \�!���Ch
�8!�/�$�y���F��<�&.ˆ(�R�O��y��!�j��7M6!C~����y
� �8��T�e��x#��s�6��2�'�1O�xwGDr1HQ�����Fex"OX	qWŘ�Aj-��[�y�� ��'ur�'�R�'��ݟ��<yen͒/�DKf���UHv�I�A�<i��˵�\��l�BK �c �2T�́wNޏ�J�)��TAQ���ph(D�ș��WN���t̑�^��"2�$�O�$�O6�ɇa��j���1N1�8B�'�h�S'�Y�B��"�:5�YH�g<D�L��Gԁ=ې�	��Z4H�r��8D�qbl
0`E�s��Q\��7D�Ȓ�+5�Vj�H��Fa�F�'D�T��F�V�h���g�C�PX{�$0D��
��7F�\dKu��%)�x�u/1�O�re �����`�D\hbi��|�B�I��(m��g�+;��T*�k7\����0?��Mԍnn�_{�t��J�M�<!aB u3r�3���[���HaEo�<!#��+5'lQ� �צa�� 8��Vi�<���I-f��2�K�-�mbGT}�<�C"ө�\$�5/���y��d�<��-^���A�����ND�I3*d�<y �=M�`��B��J*��ƖG�<�'%S�ZH���&��=���9b�L�	T���h�@��)��+G8������$D�h+F@�Iþ0�sHG�A�hSA�!D�к­�:�
LB��DG�aP�?D����G�,��Q�jͺH-� b�!9D�,p�A�)c�\#�e�L���ا`6D�<ʆ�@E���b H�)-���b� D�h �O�O��a��*�"�T�*Q�=D�C%�"Vȡ�MQ(�VEa�k=D�0��QR��e�7'�j-R6�8D�LK�BQ�EE>����S�tB��6D�\��KE��C���|zj�(��7D�@+���e:Ɛ3cH�6f�isD!D��1
['x�dQq7ʗw]�!0R�?D��5˃OW~�(w$�,��"�<T����KV�V��n��GCl`�"O�qz'ϛ3��
K��,�"ObU�"��f.�,��H+ԆM��"O�M0��<p~\`�@�h� lsC"O �0S�v���"i��M�<	zr�|"�'�az�ڬŊԠ1��lr�8:�΋-�ybh�F�
Tp�%c���ԅܱ�yr푌@T-�q�4\Z�)c� �yR̐�}u�)�bL�\k$u���T
�y���z��Ԓ�l�$c�4@���y����pB�����%/��yr�W�!g�L��3�`Y��hOL��ƅ+S��P�Sj#�4��$�!�8~��+Aj�N2��a��J\p!��\�b5,qcr�����eQ(i!�d�'yt8!��'\�6��,0%�G�`O!��?ʄV�Q|��;�Q	��q�ȓ_�(9��O�D�D���\+�	����1!ǜn�Xpy�R78֠�ȓ ӎ=K��tE��'��6�����Q.1��ç|ӰqR�쓨���~��ń�M0���V�I"G.���ȓF㢅3���X�ʼ�t��d<4Q���r���σI״5@QH_��̆�Z�rb��MQ�;��C8:���#� �N߯/��]����:r���S�? ��j�8O��Q��ә3)��x�"Ov����Uxp��,���x�7"O�I�N�/O���EK�1x��"OV�ڐ^�M>�J$�-U~�%"O�]���+5"���H�}��"O�ܘBeT�yKN��q�
�7��A�"O�p�D�A����`͵%&�*�"O�T#�@�t�B�k��C:�H�"OXt8у]<k���Ӗ��4)D1�"O���#�^���|�U�Ρu@�A�b"O�t2��]��V�� �աq'PH�"O�=�D�_�(t��ӝ5>�+�"O2�ZW%խm��ր	�=�ze�a"O���T,��6z	��A	�,�L�v"O�U���;m����Ca�f��%� "Op-����M�����`1K�f@��"OЌ20m�'4!�L�o��d��"O��B6�P�,�h��hD�s��01�"O|�P��R-*f���Ҵ�,�h�"O@Ԃ�o��.�R�ѧ�݁��$@�"O�ԛ��Sf�c����Ꝓ�"O�Z'AH�kn&��ĦG��p���"Op�xc�L�
D��ş�Y�jI"e"O�i`d��f{��d���""O�5aC$�4K�0�6�ÓM��b"O���ek̄:f��ъ'$�ik�"Ozm1�K� #/|-ZcӶO�q"OLh�&��D
��[���`�"O���0����b�x"O��7�՛@"O�Sv͒�n	��(�,�N'�8{v"Ò���J�  Y��\<��i�"O:1H�߷��Y㥋ҒK�x�`�"O�ѓr���e�d���B�X@���"O�����4-ȭ����!D��"O�ɚ0�[�fp���8�p�"O�`���Joh����.Ɇ_ДU"O�)���!*rM��ޛq�Rz�"O�[���| ��M�+z�ЕC�"O4��.�	@�qp�X3-�Ե2�"O0�8׬�d2�`�a�94˾���"O>A�Ee��z@���.R�V���Af"O �����,	�`���d�J���� "Oސ�ꏦ'���Av�H
H�X�9�"O�0z���)8rH��5�I�pr����"O�0��*�+8�j���H�-MR�4��"O�|Pť^�*8fDabn�l��l�g"OȄ!֭R(=?��ǍN�o:||��"O~�く\H֨��U�6�$��s"O����z�h�ȱ)B��8��$"O}�eK$+�1�N�^�@!�"OT��a�P�̒���,�6��"O�h`r��=I.�ER���i�h��t"O�ecã�y��6a�W[TtKs"O]�f?\��%@_�D��8"O���%���&�z�c�o(���"O�=�H����DX�@�%Z��0�"O�\�r��#&�Btxq�V/�$��#"O�p�&�����y�M\�`�@��w"O�¶�Gkp�c��`���2q"Ox����)o(	8F���v�����"O(uj��am����M�W�H��V"OZ�K��V7x���[wE�"����!"O�I��hŬ2�n�i���h:^="�"O|��G-�E0:����)l9�� �"O�  �������E�� -�Z"O�����
"�a{0f˕"�q�"O�(#��X!�@�6eLx���3"O|ADқR/aR�EZ����"O� re�I����:��֖�<ѻ�"O|�Y3�/pi�@
�cU	u�քy�"O��lÜ2�4�00��"[��A��"O��I9Y���b�0מ��%"O��+�i��>��@����
ϸt8Q"O�	j��8��ȅ��>�y��"O��裁��O�"�۱Ȍ�iT����"Ob��.� �f�%�'aK���$"O�I���زq�t'۸DD���"O����7fLL�匒:V$ x"O�a��6�<@���	���"O��PA�C�
ݜP�
�@<[�"O��$�[�YJ�څ	�69��"O�-�"�=�����\� xIc"O4}Ñ�� �q���0d��=�"O�4���ĄuX�)07D :XBqkW"OL�
�F�<^�]�4MG"{��M+�"O�%�d@	�9k�aۖ�M�M�"d��"OVrR�܎3~�uyï?<m��SW"O��Rw)I.0���ͻ2\�U��"O$w��1kJ�A�5'ݎXС"O�!��CV�"�P�U%C�f�8�"Ob�h`iD[�̔X�#�2D����"O*؋�	S��22m�T�i%"Ot��P�+@�"�������h}ڠ"O\P2T��
qC�0$���}��8F"O�9�!���N�h�e)W ^.�X�`"O�)q&`#2�L�'�^ez� 4"O6�K�e�Q0�-I���~� �q�"OD�p��	RD X�oӔu{̹��"O|��"!H�2A���T�8��,k"O*,��@�kt�� K��QyZ<��"O�$ᇇ�^{l@�ҙ|`��"5"O8����d|�pQ�ʓ87Ih���"O<UI̕��b������y?j��"O$��C�� �dP(e�NI>�02"O.e��.C<;ކ��VeC�i.��{�"O���ło: MI��E0 ҝP�"O*T�E�L�Y$��!@e�&��C�"O,�snߌ(`\�e�ו�
���"O��z@��d7����R����;��d8LO4��FC�U���Wc�%�$8��"Oj�(u3� E����<�R"O�i�0*��:�8l����*���"O.�PC�6P��[�◭N�j�G"O, bs�48/�0[T�C�*�:���"OXȡ���E�h��@�Q7�8\�%"O�a�E�#�ݡcb��,r,�"O��HN�7z�V�)@`ʑ(˸p��"O��'�b߸���.��-*A"O�4��R������P��%��"O.U���I�-��x� n�t���·"O �kV,Q?�#g���V���"O\��P�ƥ u���>"��A��'����i"��9��&`�sA�\�H�!�O' �[�͊��f��p.$=!�L�� H��"�@�p0�Wl�S!�d^,y�Td3��1��E�k�!I!�$&>T� �(�?:n�4ҁ�-Z�!�I�\�֨�4)^+wet�K /Wh%!�� �SpT�Zt�q��.قb"Oz�H6�MF؈��Cv!��"O $ӳl�6E�	1竃&a	�]�"O�<���Č'A��ࢭT�!�ʤ�5"O�M�e��<�<����@�(��'���~b��Y=N�Ӱ�֮���RtH �yrlj��BqKP�Q�C�y��x,)��m�5u�@hmS�y/�
6��*4��"l����5�y"d/s~�@�mǮh?�E�Eڒ�y��6v��a�VJQ�Z���ӱ���yrK�<��a+�ʙ?T�fբ�����=Y�y�Ő<��Y����S<����y��	!^�mxա@�Ihࠈ$葅�y�^�C	�J'
§8}Թ��	&��>1)O�YQ ��,�(5��?�d[C)=D��B�KaܒXh�b��ic�p�2h7D� ���8�X��AOR�3�O6D�d��CB����5fƎ2�V�p�C3D���� �$?�EjT���5�R��r.'D��9%��rTb$�bM��>V~lAsE*D��xT�N��I��խp���;U�;�ON�IP�tcÌ�n�z��%J Z�C�	�i4��Ή��&=��jB-s�|C�I�S�̔�Ҥn�P�q6#L'29jC�"0Ǩz�O?��9�v�KN��C�	yizݐ1���e΂TY&���{��C䉷���:��4}F8@�-(��C�	>:��u'D�'HD�(�&D��h��d+?�*]#J��T!֙i2V͂D�J�<)�$P?u�y�c��
F��l�B�ɚE̼)�AJ/�1���L4�JB䉸A� ͠������O�q6B�ɘf�"% �	�6"p��rk��$&�S�O�2���G^�2�����H&yJ�!q�"ON�C�o��p$fL>}>x��t"O��ٱ���C�tL��G��w��y8�"O��s��,Kg�ES���$���1"Or43K� 
(��Z���!pl��R"OdIBf"1_��Y���-[Rls"Ov����� M=���c+��DD(��a"O0ԙ�d�2�дK@�ەmC��(V"O
uۦ攏SQ<t�tʑ =8T��"O����J-f*U�C�BXi� "OP�� N�.�U�^'���*�"O�TJ��%�(����#GL$��"O }(�b5�j��2>�q�G&D���لl���'��4V8��$�$D�) Ǔ%~�Pc�o� <�fa��!D�,P%n���v��8CT|i� $D��A‒)���+	<Й��,D����A�[�P�`��D�R�`T�!�+D��Uk�2�
�{��
`H"u�4D����18$��e�@�[�"�k��4D�xB�)��;R���1��92xP��3D���T�J)?2�3u����X�7�>D�H`s��L��+�ᄌ`\��e<D�0���#6��`SJBɋ�Uk!��_��8(�2D�(	#��]i!�I�z��dJ��"2�d�ȃ"J9`!��G�C����(D�*�҅����!�DR>4����Ğ� ��b��$�!�$�Q%��6�I
4�*U{�R�P�!�ě!��̙�"�{* H��&Z�!�� (a�@(~r�2w�ݪ~�zXˀ"O܉��D�z&�a�떓=�A"O�E���ȭW��B��Ҏi�dܢ"O��ei�t�E�F�̂��]��"Ot% ��:*�XS����}����"O*�X��@WJr��HC$w��;"Op,Q�HN�.�������0�p��#"Ove��V�w:�%��!�2�Hٴ"O H#����%���M�U��a�f"O��x�'B�'J�ڡ�0����"Oެab'��+�50��Br0�C�"O�	�5���j �1��B���U"O,�(���)�
j�d�f.a��"O���4G�H��`xc>&-�X"O���-
����U�!.�"�3p"O� �$�2B�,�q��szܙ�"O����F0W�<seEǔT����"O��l�"ld��� �Ex��B"O�(��H�x�����:��	؇"O�P��%��|@�w�њZ���ڲ"O������Vj�i5�=a{f��B"Oܤ"ǀ�iR�԰$
V
M�����"O�h[�Y�s~��EC��zߔ@"O� Hf���*�ʡ:t�A̞K�"Or=�ԤÈ(�` 	���w��m�g"O� ���ђn������$v���g"O�q��mF��
!aFN28��X�"O��
�g�i=���g���0�"O�岀�A� <j!�#T6}��"O��륫C�@�f��"�;'�>Xp"O��RKӃn�Px��Ag����"O�H�w�#t�$|qj�9A�,}(Q"O�D���C�J�F)��ґ/�l�a�"Oʨ*բ�='�X�LڊU��Y�"O�x�r�C�2P�0��2�f�)�"O��F�ψ� J�mN�7�l���"O�@@CdX�A\���cO71�T�	�"O0@IP�=z��xQ���Ʊ
a6D����+Q�	S�$a���u����*3D� Z��B��8{�*��$�T�<D�(�7&�zp�I����q] � �	:D�L�	��:<��G�Rڬ��ǃ,D��87 ͛eWD�9�`^�]�꩒25D��薣ǡK�X�"W�r	�(Z"1D���b	8W��͊ւ��N�1%e-T��
օd��(g牘hTA��"O.�`�F�0�q6:RΙ&"O�8뢯A'FQ �aƦV�U����"O�t@�N__����N� i�ܱ�q"O�	Q��I( `���C��4����0"ONM2��Ӥ&�n�U뙐s[��`"O�Q�3-أp,x�i����L��X"O����`�?��Ёu
����p��"O>��C�.G�cL��m�8�k7"O����M�=,�R�ʗ�S�l"O�e�낚,�`���ۤ�|U#u"O�m����k�����(Ց]�2-c7"Ohy0F�2yQR���	̨Q��#"OLข�inP��h�2i|�)"O�	
_���S'ڒ#НK�@��yތ+ʂ,Y��\  � �22�#�yR�P%Ɯ�2f��@'��DÞ	�y�oBi�`)���51;���W᜹�y�ˌ=κ]��%֒)H�pS7�^?�y
� " �S'_� mYOp���R3"O�QX7eH�
�Q5h�g����q"O�9
2�wYD����\1� ɓ0"O��Y�GM ?`����@G��8��1"O�����h*)�P�]
8���"O���bU(h0� �<S7Y�f"OvQЗ�ͱC&����q�,X��"O��{R���H�,7eђ��Q"O�,"�f�,@%.��`퇂l��}�T"O�8)��P�y��8⡝-R�"OReI3��b�1h��'PBȹ�"O�a��:�БfaDW�H�"O�t��j˱�"٩��U�� 3�"O��XDꙮR9l�q�FZ,a�nub�"On���<uRp�i��"du��"O�4! 	'y���ɴ*�<V���2""O�4(�����X��IM�,��"OHM�Q���Jap�z���.�D���"O4�����`��M@�gմ�Lp�"OQ��wH�yhĴ*r�	�"O@%a���o^<Z�&Y�nn�|IW"O�j�c�5� \�`��?l��T"O��	�a�����X��|{a"Of{���s{.�ۑ��lפ}(�"O5R�Ա��Z%�� º��"O�� �!�f�`rd�HکB�"O���J�h�b9z�'䌚�"O�%"��S���b��?I�Ě"O" �� ^#B�
���(�~=�"O��1�N�-8���1���*~���@"O���`���Y�HL�d�2�"O>P��+�_z<A�̖6�8�ȕ"OT� �&2>�}��,%��b�"O��[%*̖1��Ƕ����"O�x�t�ի]�h<w�.m2y!S"Oʁ��X�"L0��7�˗(�f�"Oʠ��C	�]�V�WƘ��C"O�f��Gߤ��s��>�X"OZ���b�d����5$�p���"O��2���(R�� ���C)jP�"OE�B
�v1T|X1'؁�� ��"O�%��@ɢv��ge�o٬�K�"O�1q%�*p�pZ��;@�t=��"O�1�q�#��0���F�� ���"O����']�3'�yxr��f����s"O���&��+�ʵ��̘���"O�� P"�?u��q���?�rh�G"O�%�լ��������W�"�xU"O�9 �٤	&Hh�0��>z��Q�"Oڤ�U�_}�����[{��Q"ODu�4Ȃ�)��ݦ5��!�"O�l�3��B�%�$��_�xY�"Oty�ǂ	8��bB�+gtB"O����;~�$���ݨdY�lɗ"OD��
F�:��p& Ĵ!D�@X"O���h�
C��<�4��\Dn�Ps"Op���
ȓ>���D�W�>5�q�2"OxcAS1�.p�7�eI�-��"ONL�p��	��pˤ�ѿdH��q"O�=�7M��^�ܳE�]�c$��Yf"O��G�F79����Ug[3y���x�"O��贍ؗyR ÆWJ�N$��"Od�K�B9G�{�f��=�@h�"O$���[�����UO���("O� �S1 �)X�m}��E�3"O<i@�ӸJ�.0"k�N���{A"O��QɕLm��YF*�l�H���"O
l;EcЁ!�2���Ș�8�§"O����Ň�f��b�֠%zP{�"O���KN�m,zP�#��Dt �Rw"O�!#�d�'�Fh�cF�� �pY �"OD��Q�9߾�
Q썽N�<�*�"O���Ʃ	
�d��JKl� u:$"O�*2�M fY �	�ѻ?���"O��q�«R�>1��H�']�0�j�"O�)C� �5��iBɞ�[�p��C"Ofă��NY��ʷ&V)3X%��"O����x~r]X�˃�֭��"O4]��<L�n��D�P�<q�}�S"O��AH��D���iL�]vR���"O�ԱS���!Z�J�S�/Q��8�"O8��cƘ�gAL�V�Z-n��q�"O�D"c�9% i	dѵ"7�x�U"O��4��5$D(���5ʵa�"OM�#H�-!�Vp ᦉ�B1r��D"O4�R�%s4E�׫@�b�š�"O �a���2o-@[�T�^���"O޽a��1�|�[�K�H�(�h�"O�A����VU�5i��,�:�`"Of�Xs%�Q������$��B"O�1h@.U�.���T�orv@CV"O	����2(N����cK��pc"O���1�� ��M���
25�0��"O����䐏T�x�s��Y$S��[�"O�HسbB�>w����Tz$��`�"Oyz���!d�šQ��+�<1�"Oec���	w��W�?�&\YgGl]B�	�`��)˷&�hk�g�%^0C�?�����&�~�a$���[]HC�I�m�� �W
NBZ j�@:|C�I�u}8��'89�D��KQ.@�^C�ɞ#�l_���!ʂ[�rB�	]�0Mq3JғVw���boI*(�ZB�I�B4�聆�B����'�.Hw�B�	+-�Ȥ���	W��[�/��u�8C�	�(��C��6�H<�îK�y$C�	�=V�I�����Ҹs�bD�B�ɘRj�v�(1��xbt��0*аB��ąFf���ǩ�7'���Br#>D�L@A��;]��Y��q�Ir��:D������1=��|��*W(}y"��<D��&��2=hm�.߬Pi�Y3v�n�OZ�S��M[t'QGؑ��ٸ���'oIX�<�����,�
P�
�*+����s��Q�'�axɕ�;Hb`��/eF9S���*hz���>�I���X��J�hA놪ܫ	� �y�"<���Y
w�̋CmD_i0ۂC�9U�Oh�=%>K6F9rn�!Q�n�0�8 ��%�<ɛ'4l��Gx��#d�uȗ�^� 50`FS���O�#=	BY1T�1ٷ B�O�Q�v.�]b(�Ob��B��<��R�e�����E�T�x2��* ���+�_��Kg�	>
�C�60>��[����XW��2 �8C��<gPء�
�7����K�C�I�Yk�˃
�;*X����*A���I]y|ʟ1O*�#���@:�^�oR���Q� SA�)����b@W  �Zt������IxE�{�$��Zx�P�!�Ďg����,�(<j�X_���D!�� �|@6����Vd��ꃱz{HX��'�'wr��ɒ�F�i��_m��ݣ�фzlB�ɭo��Y��O�u&(��[�h!LB䉘XנL�.Є|�a����F(��=��"	�����q�b�Q��_3mK��%�lE{��4�܌6��d*��X��3+J�.�!�d��1��ÂݼnDv��a�F
��y��t� $�tn�;ZAd�����C䉨���j������ K�E� Ol�=�~�AF��}�TϠb(H���_�<����
?�^d EKV��0r"HY�<�1���h�'�
�iQ+����B�I�o�����IZK@����_�pB�	,}j�B�AŴG����m\!s�����O��	�<��sh�S�xQ4ۉAC�'cI�����[�r��ك�sO�C�I�nr>%*3n�/Z��$yTGR�hC�	�[� �.=v�b6���4z����'k��xr����BE�G��!h1�]����L��qTJ�=E��P�t���o���w��<l�v���ܰ?��j��`@v�2Ç#/$� ��m�=�y����5�f��vS
hj ��,�y�<	��E�#R���D�m������]�<vaT.A������$��nHX�<��-ж-@��r�N�t}r�L\�<IrG^ ;�P25/K"`�E
�*C@؞��=y��ݐG�n�z�bU�`a񆎏|�<1�d�j%Bͳ��iZ��#��z�<��E�S�"���A�V�L�`�jVz�<��G��^h|qvhMt��3&M�<�,S�IۆM��T�4.����
Jy��d��(��$���p�ǣ/9�t�P��ēr(�)���b��� $4�#u�F�HIec�F�>!��D4`E�I>!�}2�i6��Ce[�5j�1���8lغ�OzOԴG{"�'�P�hw/Ȫ<����j��#����p<a���'����a�-�"�Y�� �<D�V
O�Z�l�1bִ��B�{H���F"O�1�F��Q���x����B��;��T������TAD�0�b��3*l|�3- 5%!�Fb-�t t�\�+�J��D	ƅy�=E�DcŦ��y����$ ��t1�
��m��')�|ALφ1`��U�$��5 �zQ��� 
ˠX�,��S�N�؝�!6D��;���2�R]�$�E1�g
.�D?�S�'$�B��N398�ѓ�)(I^�ȓ�Mг�& nq��+�|e\y�ȓGFh47(ǫK�8�2���7�Zt��<5 P�8&1n�����6 ����ȓn�9[�/[/?�d<��A8�T���d0�؈�c�`���"`K2�X���T�f��u��-m��Jf��-f)Pa��r���i��hn�a�w@ͱK�ȓ#���+Ο$J���1GbǤu<=��A/��IC��z2x`�H#$}���ȓt�n$[ ��GO�e�j�xo!�ȓc�قȚ5,=�A���3^�d$np(<AS�S�hB}kr�ĩ2LX]��!�v�<��G�,"4�rQ.D��Yg	Eq�<��
�&S���ޫUC�1eHn�<q#��<Ap>ѓ�*�*2�&];$��N�<�4	Z�J-��e֤!�����N�<)UA]�iF��gG�]���4�]J�<! �H�a�0 cj\�N5��PG�']Q?l�
XH�MU��d���*�̘�W��B�)� B� ��P���h0w��w��5zR"O���G�m���c�ȹ��u;3Or�Ӈ۬n�B�g�]�"��`�;�#�S�;��`� ��/cX��	,���ȓXp����L�zf��oE�'r$��oz��'-پm5���%O�H����5[.ظ�Ԟ�����E��^�ȓ<�0�W�1����W��+P� �'B�}�`̑��rH[�T�iज़�yrG�<5�4���Pf�����	��� �S�Oi�ɩ�[$(�~�J��"OX�,�	�'�t�2���5}�Zph�B�M��<��'�$�����
7d��m�(ztL��'�����^�M	��*;�~�S�(&$��c�b�WO�a�W�÷)��l�E�'D���X�NM��f�RqZ�b�.;D��)D��0R;F5�c�%p&=�Q�9D������56R�ju�H&���a��8D��y#�H�B��Rj	,z�iw�4D�@t
Ј�̰�b'	a�ihf�/D���6�OPƌ�eɘ��lj��7D�$�o�	n��%�s@��ԡQ6."D�d#U�V6)��$
�	W��vl#LO���!W%P�R��C�(I���/ D�t����"Ӛ�j���95HX��=D��01���w�D �0��u�()j D��{s,gN��#�$�1c�0<R D��.�#%�"����� W�ash�VC�ɥ�v���&U�Qd�Z�(�>��B�I�yv}�#kF�U0�P��!ftTB�Ivͪa�V&N68���J�p=B��.�"y���M�2`����=Ĝ�<��H O�$�&*"��35!���M��"O�X��W���j���	�}K�"Ol\�ExV铡[�,T
4n��N�!�d"|����䆒âѐR�Z"X2!��7~|��UKG��h8�	B�!�DD�B���s`U��J�ZR��N!�C�C����иd����#�i!�D�+�j0������CA)���!�d�3eF ���T�"����
�!�$�-l
6.��(y0`�e`�!�Dї;&V8(���e�����]��!��_�vP�$ؗ	ӉK8��Tn~�!��;XK���Ae�<Fq�E-�j�!�$G�E�+�G�tfx���K�m�!�d�0�T-J&-U(Z�^1ӔM�� W!�$_>u��Q`$�c�z�PK
IS!�$N9G5�!�`�]0������_!��?s{�=���S�F�<K��*S(!��Y1JA	E��A^����CT#!��! �J����D/:<�`����!��V�a=������ZL��(���7�!�D^70АCg�
�4ЂK�1P�!�D�
� y�N.7�x�����(r!�C�R�,����);�$��K�@{!��*+#�(TID
��rf@`!�$F�`2��P�?�r�sd/�MO!��r�t��`�K�z�~ y��N(eW!�dۼH��V�DјD4O̐:E!�$ /��Ъ1a����}W@��1J!�$
����G%�78PL�!E��@i!��i��i.MB,	B&��!��
]��8`���`V@�*çM E�!�� NZ�g��T p� ��h���"O2Ţ!��F�3$R�IF4�"O���� ��DX���g��=	~�}��"O�Ѳ�,L-^���3k�=&�ۀ�ɴ]����#�9qxq�7��d.�I�b�`'��{�|�c6F�4!|B��.O��X�ƾ9A��kQlV WOVB�I	8�� )=x[�ɺ6�W�c�B�	�>4`c���zw��M�B�	�d��9���. ����R"v�B�ɇ����9��braQ5:l�B�I�	��Ys�ߋl٠<#3g��h��B�w]��� $���Dh
1�%�B�I �����Q�"0sS�/��C�ɨ:�E
6,�%_.�wB��i��B�)aީ󕥏�H����� --�B�	7:�.����/v�Ԙ!���vC�C�U�pZu� ��|"B/j�C䉒q�Ԙ���ݐH&��`�mӰe6B�#&��͒W�֖A�NjGg
�B�	,dޠP9�@E�����al�8A.C�	�h�䔋'.�F���a�G�I&C�ɮV�� � ���!��l�fB�C�I�k9BآE��4ڌ�@'
ėL��C�.hl�;GK
�'�J�z�W5paXB�	pR`�w�F�4�`�&FH���C�	�?��KVlńo�H���F�6H.NC䉠 ڬj ��e5J��
�]�vB�IE�|9��w �k��ߌc�B�Ɉ.�N��@ U���r�
��zB䉂Wb.t��/1��]#��X�C��.��#���k�"�41�B�ɗ�(�`f��[Fj�@@
�žC��G�n�aw�гSnQ(4�]!r^�C�	�]D�5��يf�.=���W�C��>(x}I�F�!	�:m�e�7Jv@B��4F0H�Q�喂'���1�Va�:B�	��P̚�E-ⴻ�A�w�TC�8n��!q��{"��5mW7`g�C�I}6�v�.)G��� ��9,�xB�� N��9D�~Mj5�a�}�C䉾A�,`Ʉ&3?VmJ���Kf�C�	�4��DS��"z�Zm�u���(s�B�	�i���@S-|�2e�@�B��B��C��{���D#^�2���C�'6�4�'gEP�i�
��aC���\
�ጇE+8�a!�	I�6B�	�kPP}s
�-@<�h��6@ B�ɛ"�� �� �k0�s�&B�ər)�ۧfە;����*N��B�	��@'쐙`���#'BLPRB�I1$y:0�u��R^0	4i�>B䉌;���%hÞl�هK/@��C�ɵp)��1�$).��C���
��C䉬i|`�P�_04Ct�� \�#�PB�	�3ڞ�9��X2&N2�L��C�ɺ'�������z�YC��R8C�I�9�HbGҮLlT��C ��=)�,9#������_�A�6�Ӣi0&�'�$&�!�����HZ1v�̠enγJ!�m�HF0!�d���S��M����;5��qaf
�	jT�<�bT�<i"K��i{��܀d��pJp�L]?�u�[��8{%�۰<U�!���_�sB��u"�L8��)��W�U8R�CHn8N4�ͭ"��T�e��-2l)�ēÆ��AW82��l:$�JSC�4Dyċ�Ϟ�����0���� P}y����q>�,�C�*͐8�f"O�M�RO�1� `)�dV=]�҈��]�+� �i��wNlݗ�����w� ��I�mN$�D����y��	��p��W:ct��b��~bG�9�ʹxc�ա1ay��9E�H�gI���؆�#�p>I ����ms�Qk�����ީ
F|�gK�OŠ�'4(�+Q�B3D D���!�c��d�D2&�!N1Fb?�9�nD�u�h0�ѯJ��o2D�,z��:��+Ѯ��[��mr�o~ӂYc��2 ��I�"~nڟH�T Q�d]j2���eh̢M���d�DL�-�C�ذ=9�L�(u�(y��׹,	*� �Fy��	�_�, 0��׹/

Р҇Q͖�Br�\�*�xc�혯ag��1 ��}�<�cfL�I�D��V�$/5X��ÃQ��yr��'-�΁�э�Oh���Ǉ����AU�g���S��T MU�1��g@��x�Ue����#�A3`�0d�� �=���P:\6�A��F�Arܼl���,5'�'�<�7i �gt��b�'<h�'�{�'e�y���J�hL$>9pd
��v�P)��J7@6� p�F�pWi��Ʋ<Hs��� լ��D��:=��M�JEzB�+f���$�z�鈜��Ӻ���իN@��5,�2���q�ON�I2pA�q)�>b�2�@t�W4��B�I.4���MF.M8Q��_&X�,�RK�x"�`�O���,2����ǬH8i`m^%^�"�%|iL�B!Fѐ5M�@��9�z���פcT�R ��S�n=2��^�/`�$�B �.��y�W!5����R�N�/ N�2�_���gy��
$ �h$�H�m�8�i6$�V�Xq�G I�p[���)�<~ѐ8B�fV��E�6t����w�I�2&Z}R�E�
_NttS�=E��Z��x��A�yD��'6�A�wF�&~��O����]@��¨��'UDuI�d>��Pq%	! �
��v�G�wObC�I�b��*a/A�"�	5�8nH<�H�@hC��r�6�x��1S�.�uSğ:�-Cȼ�Co��f.1�V�LQ"��ҧ-$!����7�a�!���sI���?���(�Q��Z�3�}4���I>E�įձYH�gL�m�"pA����	�߼U���>Q M1U�c���R.�Q�B���\UR`���>���TVh����=6��|���hH��KN j�2es�jX=�C��q3����,�B�v-Gc�%/�=�c�\j��3&�0�Ӣx�v��SA]!�^q�eN�a��B�I�M���;�MI�r ac0b����Dں׊��Gӷ��)�h^Lē��-�ڔ�$��awnM�
�'�ت3dvOdU!�'3N�I�*O�!ɥ��e�.ec˓$!��Y>KƁ��g�G`Bm��	Dk\AP�� vp� 3b�F�Z��8��E�%���YG�'���QWGO0x� ɳ� t��@@�1L��@E{2���.J��+���@�jS�y� �B0��W�T�U����>)���+6�E��݂zŤO��ܝ�D`�._|�h�,��`�N��%a�J�铘��ǉ�:��� A�{��Dq�ȏx����8b
l�W�O|����'(����K�A0�8��A�U3d�Ol:A��V�b�X�!��(�	<W�0�I��&XP�}����Ú9�'h�<��VwZ�yȱ �"�џh�t��7&�{p��.CZR��e'}Z5h5����O�
yi�k��>Ő��pYꀮ\XT���	u�p�q�'��[��V�Z�
�vgH&.p��{�S��xp ��0J���"���D�Ă-�̤S4r���:����r��_	��$������ �K���!@01���kͿE8�ĉ
|3�z�������'IX$0D���r=	�fY�:��d���t5�=�@a�
er���شaÖ�ip˙*�ٰ �G�{ǜaC�,������;��OJ��AOM��q����i8�h2��'��I�UFH�j�rSß<���zV�M����3i[��]����)f��~�D�3"��p�FOX���e���'�tQ���אÒ��m�9&j��C�~r�+�W�"�0�),Chh$Jo�<I�LRM���Y��Y	L����w냨F�*Հ���"�������x�>�F���O�a�E�X���fa&�`��"O�X&,I�:�^���I,l��)��e��P���?�����q�\w�Q���0�ƐF�b��
Z�E/T���%lOPMk�(�(����!�Fyp`�c��RRg�$P(�a�%��d�1��tp���T��B�Ϋ5�O�ᛣ���%�@dbb�L$f)\�"`+=��.R	bt,����/%��� ���;�yB�[�Ξ�C��E�A�xj�+P=.'����H>!�Hb6��5��W��~
� U�A/'��ա'!x�<��"OP@Ae�A�?�zg�o�D�aVMETX؃m��Tx�����d�����\�cMСY&��On1��B+l�a|r��,bVyk�nX�#�`ŠEm�\�^�@��\���9��V�[���J�*�m�C��!N��kuKM:�Ol�Q7$աhR\�2Ǚ�A�����ق�%���c�Nü?*Pk�"O9P.ΜF�����z4�@�1b����A��x����g�O?���n]���F�cD �7�^b!���h�~�ĄݷhVƘ��W��IwݨEI��A�j`V!��ɼJ)�/ۖ���.i�Hӂ^�l�R"VP8�@��n_ �la��e�,s�V��e_Z���͗l]a{b���q����	�S�T�� BPp$U��L�`�>1��"H6
$%'��-�0K�>�@� g�]�iP#=Q�*NL���}�w��b�~��ak�)�r�Ӊ�`}�c׎Y�Z\1��|����3P>�Ȗ-�~�r��d�[�}�F
�Ҽ��=E��4n���S�`��.�-Ҳ�Q���&�(�ѯ�ayBێoM��{�ܫ ��)E-���d�B�J�ߓ"�%�t�$s�މ�����R�zq��ɑW�n����'f�i㆘���X��C7gT4L�	�'���2��Ȕn�4�;���,��D���Ă&c�"~2t�ȫi���fSy�}�C�[_�<�ᇍi�	P�bƔ_�����Bg�<�5i�	y���CeJ�v�>��%�[�<i��\�.��y%cn����S�<�c,�,Do�eh�'O�uH��A	�N�<1�f�
{�("�%�;��h3@�H�<�B��!T`�p$��#Q��a���F�<��[���q���j�$P1�B�G�<�"�Y�n�^�!C�A�@Ú-!�D�<��X	��G�=[An($d�B�<i��3�l��BI28������g�<�E�n}�d�e%����ScNZ�<�櫐�5y��+�|lp�!D[�<�$�.~�Q:�l������l�<Q5ΐ*=_��� !�,�XZ��Zl�<��ˆwՊ0��nJ���<�#�E�<�C��v]��d�"0L��i�(�[�<�i�+X8�#���mgX��gGT�<�Ń�_�T���V5|��YV�<q�۸��Mjr��]dd%� hDW�<1v'N2%���ChB0Rn͈Gm�I�<	&F�$v����<���i�<����k�Pq�FǺ�5�B�i�<14)A�B���N
�v�yЭMk�<!�GM�>ҵ�1�Ҋ@bL�lRy�<�3��.`BmQ���pB<2��H�<i"�Kv�ޭ��i�#d�%�gF�H�<yk��T�"�P�<|�C2��F�<Y���@��b)<4섻�J��<��*)�u˦�ՠv�~h�fl�x�<A�����l�D�M)�pCeGz�<���b��1�t�3c�����r�<��/
,3EL���)�*��hg�MJ�<a��6��Ti6���\�FH�h�<9Q��=|v 9�H�
4�`ːD�_�<�t��1w���3�ØO��1V�<)a�ǪLET���.��i����%�N�<��*n�Sl�	(��ȧ-Ep�<2�� !>r3C���>Ȭ��Cj�o�<�BF�!��d�5���b�hB��e�<i�l�!%n����O��t�a![\�<Q��$�qd��v��1�ȇE�<�pgT�Q���
��٘^a2���L�C�<y�;.��"�cCE��f��}�<� ��򰉌�
��*Ed�$�*Las"O�����t�ܜQ�A	�qq*�;S"O��Wʄ1�ཀ�o�U���Q"O� Xah�2�܌v��YH��d"O��Q�Ո�t���+]-�t"O��G'	`�Ls��G(�d�J�"O�m!�	�f�-AS���V޴sd"O�8h�C�L| �O�X�y²"OLy`#O9�%�5o>T�b`�t"OhD8V/������:>�J�V"Ox �E����ĭ1M���r�"O�ċ���< _ܰ���T�VQ9�"OT�E(�Z������Ӽ�zV"O<�����y�  U�!hҜ�7"O���.��~��Q��@�5Úp&"O(��� y܆53d��M"l�"O����(�?���M 	~$��!�"Ov�KR�ǚUъ$�wKݥ&/�k4"O��PǓ)�^@2��W 81ʵ0�"O�&�f�X�����KݪL�a"O|KW!�p8L�����(�"Ol���+�$��Z�lW��ۑ"O4��w͙�W���C,T
g�(D�@"O�*���;�\�:6a�0%N��%"OJ�1��25n���.�m����"O�a��[��$Q�tN�ot��"O�D@�\<q�B��E�[�1 �ݺ�"Oh0�O%o�4�� ��9$��DKW"O�1Z�m�`��� f���X���"O�<���;�<�c��?�zI�6"O,�`"��rǠ�`��ފA�쁱�"OR!0���-q鎕1pBƄ|*"O|��I��i�4PKr�H)k����@"O�1P%��7�4�1�/^�i�����"O�h�,�%'��C�ᆏ(�PQ�T"O�Ai��\ +> ��a	�f��AC"O��"�G:c=R�0���P�\�"O�����(���K�o�0a	.��e"O��g� "�\��Q]P��S"Oޙ�q��6pu4��6�<~Cdm2�"Ot������K��qZ���"nM2��"O�h��"K��S ��1,%	�"O$��R#��,�D[�`b�Q"O	��C�Z���C��xw&A(�"O���p�E�?s��K册8t���x�"O~�م�Դr����Eă�l�AU"O��JEA�)0zl�E�H�OQ>qC�"O�Myq%4mQ�t���<����T"O4T#�O��H�dр#��I�h�ء"O�#3f)��"���}��|B"O p`���	=�l4 �#��+[���0"OKٳ�����R.�zhG�U/�y�K
Jhmj0�@� bkw���yR��@RBDA�D�q�!��	��y��A�]1��#i�M�A��oW�yB�7�h�����BA���� �y�s����T�0�
�bDlV7�y�L��L��w�F�7j��R�,�y�+R�5��,[rJ4+x�B�'C�!��+�����7E>v�1�!��G	Z:����Ǜ%d�Ԭ��Mgў���Oq|�D���£Z��ӶEG�A�l|Ѣ
<�y��U"�����i����RR�F4�M�cھ3<9��A0}���i�VQ��	��Q���< �"	��� �,[6�GJ߶t윸Q(Tu�F�O�X��%!`�ʕj��;,O|� K�_e���g ��`�'��$BZ�"P��ǖf%z��SJ��(�
T�҇�6/!�$̄;A�4H�j
;J+bȩB)�7L�Q�t��l͇=M��ʊ{�'An\D1��&>��2�Brn]��3�L]Y�G�-i���uTy��3�j� v
����[��)�矔;s��"2�Y��|�سg�4D�hP`ֺdvE�w�R!��ۄJ����k[����Z�e]fX���5
�g� ���4ӎD���7�O�\��F�Z�h�rp�U>_٦��LU'm-N��aJ@R\C�ɳ.eXXbw)�3��)�A��/�g�<%�"fE�u�H������^8@)֜P��L4*�6��W*Ǉ�yf��Qy2E%-�>x�vC��M[�,�(J�����6}���i�`HhѬ[=)Va�q�Re~����Ͼ݃B!��%*��D^0Z��L	D���*:�2M(f��I�o4
��P��t�*6 �r�]�d���ek�rl�q@�hR���i�b^�!��S>x2�`�
>p�����Բ��O6�rf�����d�D�A��?ia�c
�;�$�a��N7b�1�L�$
=stO&�A��ў`�l�6e�s|������E��y��G�dY���gZ�M��Ȟ"?�&��|�'��С�S&@���#cȒĮ����d�M��K���ħ5��ur�a[�[�u鴆�8�X�[��&R�5ꥀ\�Kl�1�sɕ~�`�$�����Ƶ#��M[���<�W��ݚ��w-)}Zw`<��d�lG� ���Ȫ)��:W�Wq\�!y2�q�(d�R Mo<YDCE�0�������7R�}��;G6�n���/��s�p�h��ڽ0�����
�i�ZYZ�w����̐=d�bQ�t��,c����l�
��B#�+0�R5{&	�(6pt�NӆZ3�j+Աb�ȵ��� \�0}����3�V���1n��ݑ`LL�fv�D�Ă�#�?9'�37���YC�3�	�4!���*�'E�]Ð
�d�L�n��^�I"D�6
�T�c6�'_�t�"�թ	���R��x� ��,O"x
�/�=L��	�X<�{V��+i�q�a�Љv�4�Q�i]�:���k�������i������d�!�d])	��Ƙ>b�I�Q>5���N�"���?U��#�y7�#������t)4#��]��x"Cޟ!��)ǋ�X��ɦ 
LZՂ����s��Y��m�n�4$�"}���X��T��R��ũ5a�F�䜓1���K��* (R9&b1O��������%$�!N8Ց|2dE!	JDzr� (ipݠ 㗷�LD��fK9����G�9)2��$�	1��I�ꖗj2E�F>eEў��.�hpƩ�����8Т%��jъ��k���<�!�� ��X���#]�rM
�@Ѐu��)����d��S�f���{v,�k�p��f�$;�� ���*�CbjZ���#@@}�*��'H��N�6����ɁiO6�B��Հ�(ER"@�v����	y ��9L.���ɏ� ��Xwg!����'�� ��"� ����'Ȝ��a#��䀧>��EF+��O�����9W��<���]�e ȋ�'[���W�c�jD��ĳJ�b��y~��M�Jҧ��4H��f">�N�yI�DiJ�p�<D�8�-K�ΰÂ�)W��؅;?q��R�L)�	ϓ1��d�B&V'���V�^Z���ȓwe�5 T�ϋR�̹Q�@�;W�<A�ȓt<l�33�a����'/�j��ȓW�"�1�D�q.�X9"�>� Q�ȓOTl4ҥ��b<.���"��}j\0�ȓ>�\Xwo0+0@}@�&�SVZ���C�m;4�,=,J�����4`��ȓo��,��C�B���B �Tf5���N��H�ҴP@<��LR�O��ņȓ]�D�qRl���A������ȓ2J:h���ؓN��9��
Ǿ'@��ȓc|�J�� �&�	R�Ղe�
��иqS&�ΛɊAШ��$��ȓ*��)1 ��4@��ar�u�Ȅ�PjEbg�"� !��I4]���T�Y&$U=~�R���Y�$�t���S�? B| ��N�����g������"O��j�c�,���%|�<�D�I�<�����C c��bD�[�4�$y�QmL�?!�Dߺ�����������W�r�Ʉ6kl�8�`�}�)ҧWo������L%����#e4�ȓ/��)�ĀR�,Hش���@�O�Q�Љ��)#8�
�Y�ʄp@�X�o+
ɋt(�r8���C�ta{��ˤL*���&�ޙɰ��T�OF}b���a0`�#��
QMN���O:%{֋�3
����d�ݴL᪏�
��apE<�y��v�f�� I���\��璷�~cGM6��DT��Ӄ\j޵)���Q�����C�	%V1��E@6?���34�ת@���'|
	��O�P�����I4e�M�$m�r..aP�.�183���D΍aـ!+�+������0�N�wk�]�֠�	�'R�=@��5{�!i�et�p�Z��$X�6�05iӧ���O� E� �����ta �����'g��Ƥ�6$NJl�鉅@��0�O�)Q�JM.�O�>9���R�]kHx������aH>D�����?�`�{�� m��!�g�>�� l����<i�E	/���� `*� @�}�<��e�*� $6�̳\m�T��*�t�<!�(��kF }���,f*��F�H�<��G�8)DF�IG '}^���b^K�<1ӮP
 z��Y��P$Ȧ͹�[S�<�2���f�qdS:�VU�4
�H�<�a`�DhB8 1��24K  (NC~�<�AQ�`*� U�ߨl�ʅ�PÍ{�<)�o-v��Z�B�=/���C�*�i�<��O[?\l��BVRv4����}�<���a¼E:�χ!�F�򳄔z�<�q��FK��%Y ��j���S�<��ǈE��ԅ;V$�2��RC�<I��~,����Ϝ}b*!Į�~�<�f(�\�6�sV���P�W `RB��5s��#p`��AZt �i�b�C�I'3' l�Q+؎(�Y������C�	4P����*�-lHI�s"�7n��B䉟*�@�Q�J��w���HGkI���B�	**&<��WhW�<��x	��YψB䉅hۄ4@D� v `t�E�T �B�ɭ9 A!�/�V�:({�ߐ2�lB�ɍty�����ծ	@@�r��!lrtB�͊�%�NxAT�H8B�pB䉇V���̍�
��4�WB�*:l4B�I�1�00�ì��
� ��ԆJ�X��C�	�y�h8��*#�P:�l��%@�B�ɷ[�$�{v�V=���t�խ�ZC�ɍ-�`��
>&�+�l�d6$C�	�x�)(v!�	EF(�#�b����B䉪
�������VD$�>Hu�B�	�aB��0E�1qx�vF����B�k�E�M����B�LB�B������(W��Mې���c�B䉢p�\�ҍ���BÇ��\�^C�IK888�d����_8�:C�ɔ2D*t�Z9t�Ia��C�ɏ�M��,�<]`8��.G����8�d(�$X2|l�Z"I��N�V̅ȓ!Ø� BY+�y��
��6�~���z�.|���ſ A��h���z"|�ȓ,�y���<8���u�XX�ȓ)���d�Ԓl@�30!�͇ȓ(��<[B�S!zS�9��`�/!�Ї�S�? �HǤ�'(H*�+� ���qY'"O���*�Y��(� 䆶q���۶"O\a��ӧ1���)�B�}�$��g"O��{��yŊ�ȶ#R�jD2T"O�)�@]�[B�Ő��l��);e"O�M8G�G$e�<m�D�țP� d@�"O��qv,�
|�ܴp)�s�$!��"O���1��l�<����Νsƅ&"Oj���	�Jl�!��D�[u>��@"O�ti�LO��X򤄗��H�4"O|+
�&�!����k�p�'܊�`pX%���z�K+v���H��d��P<�P$�;\�bu5�����
@�b�����(>Ь��+Jk�!�$
�O6�4e^2%�M��L�_�!�$C#1>4���"H2 �k�!�D׃`�,�1�Ç<t��/2]&!�DI�b:�$��M�)O̠�qE)ؾt�!�$Ƣ}��I�g��C��y�a	S�h!�D�0 ������?p�)�q�N�#�!�$�4|�[ÅR�BW ����^3!����=�� ϶;.T�!6cǶ>!��O�����fNN
��K'�]%`!��F�Ot)kg)�!I�Q�C!�[ |�V!L'|�48�ᡀ�AW!�d `�fm���#�:�p���;\!�D���`��^?Y)5y"ϒ>$I�O�]ڏ��)�T�f�}zs& �8Y(ׄǹ�L� #�u�Is1���~*&J(�D�)p�sD�Q�G�(b�6���i؟�9Wd��%~։����T��� ���&��aif���j�6NU��'��Ȕ����W����1����
>�������P��(O�O|�ɀA>ձŅ��u�
�p��� ;A�����(OQ?�S4��2U�)X�A�g�q�Ǽ�(Ox�}�O��Q�o<�CHL#B��'>���?�a�P�1K��x�x���)	rI��OS�hhFLO�b��Ң�� ��'�"�eo>��I
S��8W�T*T��:d��`��*	><���%��Ʉ��|y&'�b?��nW�
\�eCP�杖9cD�>aG�Z�� �"}r�(��Q�q�$��2HT��PR�<�B�/b�	1Iַ+0��"*D��SF�n���TAS� ��#�d(D�l����qK��qT��^4b��8D�<pu���81���YJ�"A.+D�< Q�S���Ň�P�8@��l'D�������*ό!�"���?��L�%D����S�4%�`��	�l����$D��b�@���h�揱�2&D�\x�ǘK�h���H.0(����$D����� ��L{P�F/(�2m@r!D�t�5�C�Oo�@H�X5��3D�l��eȹ~D0@���V����1D�d����&JJ�8ኤA �d�c<D�L3a�<yFJPQDF�ojI�p�;D��v�B(<B�d���\��&D��P
W�S*��f:@}�8(0�8D��5bW
;N�J���ʨ�x�%7D�l�AS�'C*�Pb�K�h�#	5D�\�O��Y�hdIU/W�k�D�� �-D�l!�nK�6�f�
B䀦}4T�$� D�Tjf��>�R�	�)�#R X�T@>D���u�v��@�L���i{a`<D��*�5i���0ROJ�:� %R+;D�D�!mS2o<P�hLˍf�H���>D��(�\4��]j&�
28�V�I$,<D�X�s�NxT�*����ؠ�'D�����f� r�Ƃ�M�=sV�#D�� ��K0k��ze0 ���^�~툜�q"OvAbS$��o�h8kF�Ԩ~��	�"OT��djP� kBp�E7;�X&"O�uXÍԍA��je��mF
��"Ǫ:�n�*c?�PS�$\GX��"O��0%�ܗHuL���F	g4�LS�"O6l���=�j�Sb�Q��h�"O` �b�C�%�
|#��?m�@���"O����U�3U.���BK-�xZc"O4ᑄ�ϲ^���v�<	�$��"O*��æ�6��-�"V�w�͋"O�k�A&Jb����&Ώ(����b"O�|Z(ޱF�HeI�����18�"O2��B�! �vd�B�<1Z0��"O��AB�ִ$A��2qJ�l(�L��"O0���[���� eB�,�h7"O2�(rFS.8���"�H�J���R"O8I�1$�(�t�G?,��@�p"Oh�K���%�<"��P��L�
�yR-��@��cve���XđV _��y�'
��(�9%�7d$0����yR^�bB~�Y��R�|x~�P&L�y2"��`Sg�>c	<�`l��y���+u�I�e�S-d� ����y",�(`��`��爗G:��p�K�y"Q1w�L�z��M�P8��V�y2'Y>L��iȏ�H���(@�=�yV�4@R�@[�,�4bD��y� \@ٻ5"�"3�		�%ה�y�eG�<�[��Y/�z���lV=�yR�O,����lS��:�3���y�RJ��@8�&)�X�ҥȝ�yr�����aAc�����d��y�̛T�*�qvmO<� {�$�y"H�7I`U�@G-��%���y� L�_bts��R<;x�A��F��y�bB���⁕�3( ��y���C�E�F�*��3�B�yR��]�d�@��޺����"D��y���8>yDB%E�U:���.��y�f�"�F�)WE�O�Ȱ��˾�y�
�`���: "#E�t�����yb�ߍm tp�&M�:o�x��
�y��B�44d�
#$Ř+nZ��/U(�y��JRI��	���vi�xi��ā�y��S�}��u8�f_�m�
�x"�V-�y�(ˣ/�5�p0�M�Qi�y"�"=;�H`@&<�@a�I�y��n  xZ��c�^yQA���y��N�w�ĉ&�ޱ�%F01UZM��c�����"�^+�h��Aݥ
}�`�ȓqxi��'I�������P%��@tA�Ѫ�>N����Ha  �ȓv����R�-U.�
D�uo�y�ȓ2X\�hj<8����	-�.H��:!�y���Q���!�V��}���ȓ)�� 9E�I;vk���6�8�pI��/uTirV�](�;V�ݢn��Ʌȓ٤ՋD�U$@��I7��i&��ȓh�^u�Td�iQ:�DLO4���9���τN^I���:��D�ȓ`�*Ց����~��H�]9u�C�Inp�IQM�q/fD;uq�TC䉓w�̄Ý4Bu���T-~@C�)�  ]+��3w��I���SR��4�A"OF���m��kG�ՈpA�r�p��"O�$�uEݨSʐ�F�d��qXp"O�ɨQ�P"~�a� F�\��<��"O��'��;d�)��Ć��� "O$��W�)���1�BɯG���"O6� �:O�&y�OY95����"O���]�O�m�T�?�-��"Op��dZ�m��#ܥ&��e"O�����O�N��p��Ќ9����"O��:�'v/��[���9�r"O��Y�·2���y���!	���	�"O" **1���S��jT�d"O|�p�LߺVH�q; ��p6u�S"O�)�P�1P�{7��d!te�3"O�|8��M'���q3�#6a��"O*�a�2��ʲ+R�0h�"ON�v�ŏRpHE*�J��XI7"O�Is֦�$Y�j<p�HS�"O���P�(�@�����"_��(i�"O�X�nΰP���J�"D`*R�"O������4#dR��va¤o!&�G"O�ip�Y�4�����	
�NJ��"ON�Y���,ihdEAfHR8*�#�"O�T�!���a��<_p(0"O�͡��G�}���qV����!��"Or}�v
�a̖����U�#���J�"O�)�F��m\`�$�[�p�(9��"O����0n��r�J��r"On��4���v��+�!o�f}��"O�"��ʠ669�EJ#|aJ!
�"O�ip�D҈X`�hX,Y�\�9�"O�qѦ�#x� ��G.?�:�"O�5҅#"����W�φB��!(v"O�(@&K�0�	�#P�~�"�"OB���lH�kvN��r�*�ڭ�"O��)֦�4tyZ����.B�H���"O�$��a�d�J�S`'F)DsF���"O\��"PY"X�v��4�*`�"Oʭ⑍�%mS8��eKԋ�VH�"O�E� L'"�fH`Uh�3k҅�"O�@!�Z�O�N�rt�L#ꪘ!�"O�}�`Q&�ݪ�#� t�|T�"O6��� �([u�IQD��r���Qs"O�P��&�j����ծJKF��"O�!��-��)3����N;x�"Oƹ�S`�v.��0�̽9�6)B&"OH1B�"��kb����A3�"��'"O�d�b,��1ʨ���jY?,�FE	�"Ou��C-b�L�C��	6�� 0v"O(� &oE��hb�Ĉ'E�p<jR"O�S�J4`��ӣ͝sd�QP0"O�U��N�9��A���5��p �"O�A8���7x�zq�	Ӎb�4��"O����E^3o<)`r(�Y�r�9D"O�L[���Di
����Z$�8�KW"O�T��E�|�e����V"O���&��?�x�qb�T��z!Q"O0:��Ņd�Xy bI*�d���"Op��'�؍�傑�I�$Ϟ	�5"OzB3��#j\����u���"O���Ta�60����2��y��y#7"Oh�� S��<Q�n��4�|2�"Oژ[�*�v��e ��{j��S"O� )�t��5����H}jZ�*e"O8���m	)����@��/]p�bb"O�
f%�K�8�En[�U��[�"OJ��U曰	b6�q�� V׶e�"O�b���u����8<�\%�!"O� ���(-<�{��8�B�H�"O��)���*`r1�Q�:Ɔ��E"Of�b ��/$��*$Ǎ~��A�Q"Ot-i�o�(H���W0mP�IQ"O ��/���j��0%��J�xI��"O�P�J�t��4k�C�Yaz��"O0�1�8�J���@M�� �"O�-��ƈ�^�P���g� :�"O\�P�,]�]�Ea��=x�*pJ#"Oԕ��׈#,zaxG�^b��t"OP���@oܘ��'�1![��"O�y2T�Y��!A�õ9Hvp�&"OlԸ'K�'�
=�a�N9��;�"OB��f�9Z�z�=|MI�"O�A���;D
�H`ꑾM[z��A"O
8[aC
�]�F0I0 ��
H�U�"Otq0�aj`�P��P<Z����"O�𖉚0��<���a:Fp�!"Od0h���)i͂��臊$��Y�"O"Ab2]��0�e�����*O� fD�� ����B��	�'��m���nm�͌;��	�'i�@�wb��pI~-Z0�V�I�Z���'��@2c�?gv|�J7�:OQ~�A�'��<���[<�I�J�7T��)�'W��LѨ9��!8�i�=4�p�	�':���WǙR,T����15��h	�'�p�V'�	��ku%��u�xE��'�v�s�kE&[�6Cf(�1<e��1�'֔ �O$Ema5g��0��2�'�V�k�X=A���%D�*���b�'{>Eb �T!�1y0��5�t2�'/��+֧1�$ @P*��N���'j�Њ��=�V=��������'E�p�����p�Jp���� ��'���9
]&��!k��h�'��%�  ��