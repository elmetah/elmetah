MPQ    ��    h�  h                                                                                 |�B=S-ʵ������*�������0�%��Oh��0�4u.����r���@��,6�6��Î�I<�{ۻk"TI���a�x��������0�.+E�������L���Y�O�^�}.p�A��.jU��	=XB�W�t+'+S��V��4ϗs�Z� f�AX�]}/�f(���{^���M�"�͢���UMS�͜�o���\���H��0˰���L7L7e��.Sz�_ȡ��d39�.���A�ɪ\ ��H�~F��``�
r1��98��/�6�]�v8f��6�R5K�衧�"�v9����ݯf�8W��1GV݆Pl)j�j�Z����Ĭ~�,q�๺������`x(�z�]�-%'�*��JEV?�q�΍�f�#$i ŰN<��_���ʶfl�	����+BD�lBP��Z�B�bNŏ�#Dkl�����xqԧPE��R������8	��9�.#Q�-E�������sVW�	&GM�dšU�4D>�bDq������T�����|2`'Vt ��g�C R.�Ϛ�P[�(j�*i^C�u4�yN���#�$����`�:H��$/�ů�Y��<3�Ȕ?��IV}�e<K4􏻢�'ك
�W9L���?��r��j�4f(M}� ���1?J�8.gQlD`�.����vLl8,xo���3}��t'���~lpP��7
5!Z�=���l�ʟ>��=l�$��� ��?�nBw( G����� +���)�7�8�2޶�1.Nz�.~恃'���4����@�&5�D�3BƋT���!��V�Q���ຸ�2��?�9i�뒇,�^�H�ǰm��ع�e������\����&����%[�᝷d<Q���]Ĭ����������[�9o�|>_`z����;���gt<�I
���v��ZS��Rj��M芸�c=�������wD�fk���9�F3Y��t:^�n�:۹�2�/vKΜ������vT3�6R7q�j��d�M�|���{[�xʑ{�d{h`�A�b� t�=ͱ3l�p��>"|��Z���G�Dzg��60�t�=k̃QN�-1���+����,0�*���BY��;�&w���S�H���=`~��8�r:�(@�~C�y�Y�q�y>(9����pj#㪵e?$�s[jLnu?��|h&+��YwR�u��5]�o�3���\1��OD�A+��nzb/8�P�L���3;�q�va�~Cpz`��a.�D�+H��!�_p-t��潖$|=�E��)v1ngMQx�A����#���4/��'�H;���Rf��D��7��� �l9�*H�0dƍ�s^��+ �$�����ʾV
����T����*��	m�1%+ua�V#u��9��A�D5 X��-ۚ*�*��p��	�����uo`{�X ��Y��66�h���'�k�#��+��k1��w
%,� �����s~�S5�s�Ċ~��`��B+�׆�ó~P.i��58���՚�VMz3"���_�Ċ=v��xQ���,~�C�L���n����5����O�J$����W���Ed���b>�gz�1��X��W��j�[ڂK��wg�p��r�]�%�^�N���DNA�.��:��]
�+w3�F9�1�����^�ݑ�{i���<�Ww:��Rr֥�vPڇ0h�c^���Ŵp�/�H���J�_a��cb�����}J&��#�ַ׀h^H�_4)O{�F�[\�|���o�6��i�襅�"Z����2~*=�~l�z�_�Y;Z܋�hp�H) !��"����ʝ�qBzp�W�d��ᇖ�w�X�D#�'����&��4�'�*u�6�9AߕG]�t1�6E�r��D�)'7�k�^b�� m�����j�.�:��cfI�*X��O�<f�n|�Y0�"�1�]��-Ω�}gdð��tM�5���{�D!c�� ��뾤�i�3:n����1�RB��f8��(Nk!V6�0�	8����F[[~E{&���Q�4�u�bԻ<d�p����D <����R�u	5�͑�=w���g �}��z�8+T�����]c�B�룘2*��aB���?�S#�ݯ���~�!�P\*�ivɃ���t�re\��B�̃E[���������ڔ��ع��G/���5��щ����^�}��0�Ƹ	+(C	�J�(Vb='�F��콗�n5;�ʪ.�;'�LzEJ]�qb�W������[s����2]R�$�'XY�WZ>D��Ԍ�/���d�6��,�'����W5\�_��.��lD[�v��F	��y��e�8$�{2"]�:�h�|')�o�V{K�YݚٟmX�F�0uN2�Ö�C?D��JÐT��EѦ&O4h��7�I�7���h~DJ*՜7ʹ��Qp%�m����K�@�d����T�n3GHv#n6r�:�007��v
�����XY��hh�7a��~-��@�H��fd�Z��b��X`�t ����)�2Eѯ�����t�H�ޙ,�`O8��X�J?���৊�]�z� �1Q#�@>����	^V<�Y�*�������$��mSL�#δ  6@�j��=�ꪌ���sfY���`�VӜ[#"��s�[�x�|Hú��ml�;	w��b��;fm.S�T�r_c����	��s ̋��$�f���L٤��\����qς�UG��dl�άrϑO���d>��
��{�YH�E�yE�����/d�G5�n߉?rk�l�H;��4���f�/�Р��@�~�����ͮA:\O�gZ�5�rJB�L6����<E�ғ����Sh>"4j�2Z�I���{�إ�F�ޘ�נn�P*m8o�5=>~��|ߊp�s@�V�����XR���4�x2AJ/�ƌ��p�[����j0hY��@+n�BM�Q���b��0��qL?���ǧxxLL�n�Gi��YK�Tb	�d�o.�v�a!V�}j=���[
<d"bP d`�WT�3��4�IS�@h+ �����gxi~�x�����z���P�sYû�\Q���;�,S]m�	�9�KU��_�%�A�{8�����<���/��0h�<Z0���g���t�>��b�Al�P���ξ��f=�(��ݛ!g�@fB�&7t�Ǆ\^X��K�G�2-F������T��FU��w��F��2�Y��!��^{}�)�b8(lt-���e>��U �t�sm*�8d����慒4g���J��~z�~���_֒�+�*���9��^�@�WO
�pJB�.�Ţ���U8d��_s %�~^�Ӹ���~IK�eN�8Cv�?�<��xB�3=�����A�%lDҾjk�"�}���H��nk��j��� J]�xC`�zl�-���e*����V:(:�)���!Zd#?��@�PNL��V䐞Rfg �;����D	��B�KZ�T���Q�8b[kg̾�b}x,Q�P`�WR$�����sk;���.��ƈ���[�\��r�WP�j&"�d 缱H>�
�q�g|�]� ֽ�3$X2;�t[7�g�+�C�ĉ�*m�P�(��0*����P�Uy�i��v
�Ԟ���`����0`�/h���4�j<nQL���知I��.e�~���f/��
�5�L!��?2cE���jA��(<� ����d���Q��Z`XZ���Pv^��8��c����!��O[��p�l���2tF!x�=��!̇Q9�.��K�$�Y�����:��B`K< cO��v�{e����)���89�t��1�N��9��Bu߯L�r�z�abDD�Ɔ��F�Ce�l=���i�������K|C��(��N����#��S�e�����="
ێ���&T��蒩+[��u�ߢ)��C��-����92�N��|YM�z"�����Ԣp��䍚��m��)6���h�`�3��=����0�E�3�f	AO�ڻq���"3tJT���^�GQ�u�����vF[����Ů��TN�<R�Xj�Ӓ���f��m{VA_��t,��D`��b�ko���n;����>��i��^��gW0	6Dtq&��.N�����p�,Kq�*JF�B4i�v;w.�OS<=�+��`9y�8
�U:��Y�@��R�{9�h� ��p��C����?��
N�BL���wX2&&�YҀ�u:�uP������\l�}O��+���zr�h8[�	g�~���L<#a�p��\ ���e�HJŰ�zw��d���$O��|�����ٞ1�OM)�\}0ڑ���q�>4jz�'��t�R���j���:�Z��G��9X/bH&#�ƈ3�^F�[ �rU�7���F���#��YTA�D�%]	���%�(�q�#�AP(��lp�|�X��ە�*�}����8Ax�
�uJ���< ?겞�ݙ6���Uy�k��KǦo��Fm�Բ��,�Q5��3Y�βT��/⌎1��=��G�}��!��y��wE��Ø��q��*MU�R����_��v�����P��p�CɖG��1n��H�p^�+�x�E����6ձ'd�&Ub���z�3�������e3U�ݨ��2pp*Чr2�%h�`���mЈ�N<�w�j8����Q�*ew~�F��6��ܫ(3^����.$��0�<�M�:���RM��T����cY�ײL��p|�H�b�JRd�������
���s�&����1��#���z �O�2���\��4��6���i����?Q��*��lןd_���;U<y��υH�s� <G2"z��ե2eq}���=��g� �X��\�_��'v߼��=4�b���	1��A:K2]��r�Q���(����DpP7�y3YϙbBø (�Z�����{l����IW�X3@��7�(nג�0�-�Lҵ��>g΄'4��Bd^�����iQ5��Ė�*�~�ŘZ;]'���d��:�������mf������!��g0|�A���F��9.u{A��׍��$��QW<��{��jq��s����D��Ff��~i�x��~�G�x
>Xb���X����!��]>�<�&7��$Q�j��'��C�S>�~�%wO~�d#�������d0��Eo��$Ot8�r�z���0e̾��������=�e�����j�iQB5��a�Ě��%��^{,k����r�+CԪ���V=�q��T+�X>�n0�Q�%d]��L��Jر�b�F4��6��-�s�aAf���XtT�Z��:�na�jk����86���΂��R�P�_m��.��l�u��oF��yt��� ,�$���"؃z:�X|b*o��AK��m�4XaW�01��2��ڂ�AՐ�lb{�9��ߪhp{��d�d7b���+D�++�����[�Q���mRW�f��߈���NT�z�G�ی#ur� �0����_8
q
��yaTYγ�h`6����~��S@R�F��8��kj�=����t�.��í�)*o�E�w���qr��XJ���,&�C�[��S��J�,Q}k ��4H��xȕܜ�1�[7@����<�V�)N<����P]��k����LlŰίC��{���X52��¡f�������Fӗ$"Y���wA�����H�zmG$�	R��Zㄖ6��.��D�-�Qc�*Z�\�����P����$ERl��Fp��#N��	�ݲ'�'����X��	~�,�����t���ѐtt@����E���������n�~�ͳ)�'��;�,"f�yH��U��%mF~����vz�i�`\j�cZO{]r�>G��ƨ�e���7�a��߀�b�&hY2j@��5ww���]�s��F�b���8�)W�EE�oS>Y:�|1k��V�����3��ڝ4�;>2g�J
���~�H�[���ś`h��@F�B�Pm��r���q���:=��">�x3���}�G�Q�4�TTP)q����.��_a|4}%*��wX
��"=GNd�ڐW�6�3�7���?k@��\;33XF�BQi��kx�E����s�Y�"PEv���G��e\�(�,�������9��U�r��@͚�� ~�w�|<1t�/@�c�$Z�c�����7������,A��PVaι7;f���(_G�+<����C������\�D�ޏ���-Lg���5�>zҺ?���y�E����2z�3�Y:1�<ߒʏrh}p�K���({5���n>��y ��-s��ϳf��E��!�s4$�z�@��{NS��&����p�ҿ�t�3�����Rx�
q���+��I���7�U	��N� �*n~Y.�.S�تd�K�ç��v�P�w��U�.C���+���l_Z�j�Q5�X��"�зb����;��o��Ypx^ӵz���-�P�ɠ�}؀V5�1����#Z����N�SȌ�}\�+�&fb�r������.�D$9BF��Z���������kb��v�>x��P{;R�?q<����аI��.����]i���Α�W��E&���d;���L}Z>��#qM/s�<��Ǽ�q�2t�ρgLːC�W���_�P��f(�π*_o�+dwy�[���a�J�`X��K@f/�l%��<��C�uN���AI�Oe��D��1���
�3�L\O1?�C0��/j��(�� ��7'���_�Q�%`����v�h�8�+�Шv�B�*��@�l��f�-��!��=T�̢�/ʕ=���I�$*4�V��50�B�?P �����X���䍹�Q)�8�+���Q�N0���m�]c��*���M@���D�0Ɓ
���c���ä�c(����n����^������ި�éؾ�k�>�#��e�3�6�	��'��z�&�3v�MU�[�V�Z)�x]��"�M ?�݅��xJ��|t[z�us���݌&�1ͣ��j� ����-���!����=g;��k˞�A]f#��5ݭ��/�3�.��#�^��$��B�ho�vAH�W�ig�Ti]�R-��j|�Ь�0e� R�{Q���G���� E`Е#b��Jw䱩�j���>�)��~��*4o?g�x$6曘tF�5̹�(N�)��>hq�+��,f-*��VBll���sw�ػS.����`�|8%uA:����4���ޘ���4P��[�xp�g��a�?�-)��L�=��T4&!�8Y-�u���kߎex��޽\�_�Oz]4+�/�z�4�8zR��~���'�a=s�p��'�W���	�H�C����j���s*�$�$�|s����c1$�M��a�w���*�L��4��'3xf��,R�@������}���"Sl9���H�5�ƃ��^�#� �C�R���������7�T�p�� 8	#E�%�t���ڲ������$�b5����ې�*s]+�q� �S�q�+u%Os�V� �=D���U6P�D��PkVC�!<��!�1���,M®��}�)���,s��Ž�t& ��N?�Ϣ׼�ѳt��AE��'w��v�����M0w��V�����v�j��Т�C� ���@�n�Z��V�ƅY�@��8;V�l�d�{�b4�kze!���ׯ�<��`�*�8&n�혼pE�r��E%Cc����6�#��N7����২<��U�w�/�F�7��q��Fi{^�=b�O�^oV<�c	:���R(���xއf��cT�Ͳ��hp7�H�cJ͈;�]���::��T�Z&��5��������HOq�]b��\?�_��R�6�X�inqx�X�}0̇*��2l�_G��;P��O?H�޲ W	I"���Հ�4q��Ȁ�Z���W�[��X����z]�'�/���6�4�F�`�X,��A� }]ZV�l*�#���D@��70�}T�)b��D ��f��}�$b�����I>�8X��6�2��n2�I0:0��g@6�xp��_���?#d�����B�ħ5d��ı8Y�	ڠ��v�q!|��_#�:$��DHЈ�S�\�B�ޛl!�:�0�î���F��e�{\-���������<�#��B}����v�E���ޚk�C����������G�s�3�d�Ю��-ֳ��G�]D��a�Eh?��y�1��OSY���j�~}Ǩ��bKC�_i��9�P又[tS��r[�o�n>����B��n���=�I�ߨ �a�ڳ΂��5\@���n���Wa^v������+^���@TV勔�3���n+O�=l���L�/2JS�baUv�G���#_�s�f���Ez���LX��Z4�1�(F��`�!~36��,���Qmk �_�P.�v�l���Ĭ��F���y�����$	"S��:\h�|�'o4�K��ښ��X��0L�^2�:����1�SW[��J�vG��܏�h+7M�%�7���fiD�L�m>�۷�Q&��md����&�Zj�_�T���GM��#�Dr>'�0���i�
�6ĽT Y	�h�T]���~���@�x��,jP��Vh���t6����j@)��"EG_s��P��j��i�,a�KnP��N�J���8ޒ���(�S��Y�1ǳ�@t5&���vV�ۂ�X���-��޶�Ә���<L�Ϊ<b��~�[Q�s�a��/&�|y&�To���.Ӓ"�ȋ�ъ���>����[m"�	�I���*�1�.	����:�c�Ŀ��O��%1���$�]
�����Z�����D��Ȃ�>T��l�D�]�������z�"�sX���ђ;~�E�N��ZD��}��nՓ;(h���o;#>'��%fa㯤'�5���/~�����Y��$��\��Z���r�S|��v�� Xd�2{��IꚐ߁ht�j�Vu7��0<����F��b�NB���7z`=�oU>4��|U��ԩ;SV�\4�P���~F+4y2��&J��6�HO�AA�[���� '^h϶�@a�}BC���3&��㠧�A5
�}�x�/��6�G_.��T����{�.��2a��Z}�6���
2>�"^ld��qW�p�3򤅂�K@�w�V�Ӹ�ܙi��xH�A�����_P �����G#s��,��؄�/��9f�UJ s�[2��q)��R��<l�{/�}�^\�Z���K���R<��jr�����A��P�Flδ�~f�@�(u�Fw��6�Q���f��\������t�w�-�������ҕXK
04��J�2խ���W���
��}K����(�������>:~ <�s���.��ϴ��\�H4�����>p�'M6>锽��	qA����aߔ�X�Mb
�����dv���U��.�ծ� [��~T�����ej}K���.��v�r���wH�Ǒ�)iD�B��ݷ�plzjja�3�3��](������,����ڠ�t�xyf�zb�--��������V0����I����#u��6mN���
�ƥ2f]
��^��A`�D?qB�DZ�6����n?�k]PѺ�d�x��vP�X�R�L��Z�䕑.�M�>H������;WF�&�B4dvIF���I>���q������*)�2��tчFg��C�
u��q�P�Y�(��*�'/�,�y����ؤ �ɞ�T7`���f@�/^pB��u<�ͯ�����IgV�emF��a�d
\QL�(9?hD3���j���(~2 袯����(�Qe�`����av'�8]����i�~��#Z/ulAtU�(�}!.�=��̽���m���hQ$e.����0�*BTd x�x�+��q:�����)C�8o�i��.N�);��x�/ߥ�#�(��� Dz;�|������ढ�ۢ��ߺI��:1�a��ܴ�=Y��y,T�Y�Ileg��q�IX�l���&
���!�[K>�����Sӽ�]��ny��� ��5�j�|���zgt�̣;��)��7���-�k6ʰ������*�)�=BT٦��Hp3f�$+����j��3�2P��M^���qt�	=v<�W���'�$_T�L�R��sjW����w��V>{LQ ʢ��i`�o�b`%D8���7�Aq>E��Au���O4NgM�6�mt�7��T��N�Wā�U$��+�,��P*@��B�<��Hwd S���a`��&8@5:�P�M>�*��B`�/����pFq���h?�
}fL����on&�Y�=Mu���PS�G�c\��<O�+܉�z(�{8�>�r��qI��Lax�pK�#�R*(�U�gH�Dۻ���,�N��$��g|l�����1�,M���ܒ�xڇ��'�4��?'�?�\Rw���i�/������"�9Υ�H\hg�~�^�h� B4�m��<�f��r��Tw����	~��%\�C�����7�V���l�C���ɟۋ�*��x�,�!�nݓ� 7�u  �,C  u����M6�[9��|�k2�ǜ(ޖ�D��(�,��w��u��=I��y֊�]/��uU���}�W�og�-^y�f�.��C�~MI�鑍d��H�v��b>��]�jC����_n_�%��nja��;�������'�bd��b��z@IQ�	��(�L�[��ړ�[���]p`pTr((\%6���tо��N2)�� ���xmԠ�wt�Fʵ��������^ױΑ��y�ί<��:w��R�'��k�cO�����p��H儐JH��8I�u�p���f&~�Ⱦ�3��\��tO�1=xV\z+��j��6{-'i����K�Gb�*��lMJ�_�};K\(�y�HDi� r�"p�[�4q�jÀ(����Y��v�XC��˕*I'l�e����4P9_����'A�(]�!��E�ߋ�BD{\�7���O��b��P ���<��h����VIyYXi���-j*n�	�0��l���������:	�.ܷd�������5��̱����O�{�|����
w�Z�O:9%��VУS�׎.��r�!�z0������Fl�w���{w|�׃.���@���<5�Z��:%�U��1�˜!��!Ͳ^����o��v��np��x�i�H���)]� ���zW��e�S�p�St�x�~�~XJ��A�޺S�Z�Dɔ��J�tn�Rr�0�Ilm�4��������
��du�ۤ����Z�_�'57��:c��[�X^q���A�Ը:��+yVƇ�H�V�hv��2���n&	��6[�l5�L���J��b<�����2���^s��+�Cj��U^�X���Z����;��u���:�6�=�8U9�����g_c&U.���l�H�G��F���y*�?���($0� "Τ�:7��|�JxoϮVKګ#��/~X���0gM�2����oP���U�%H�q���7`h��ۚx57��A�6D�����?�3�Q��Im��w��,V��k�:@�T6�G�bb#�r�MG0a��,�J
g��/��YDB2h��_����~>K�@�^���@P�zO���#	')t�a���G)�G�Eg,�P������Dl,�Hh	eF�I)
JP[4�pI����γh��6T1,�@����VM���#g�ܢ �!,��[��}�L�zTΥz]G��D���y���5�W�.
�}�1MӍ�"�����_��鑺>�Hm��7	��&�D�,�z.d!��"c	7W�R;5�q���<(�${�ঙdkٵ ���:D�����L�r�#�Z�b���B?�զ�.-+��,˒�m�Ep-���i�ڎn����<�ȝx;>��"`vf<m'�b���[&�~��O�,Y�ߡ\��SZEfZr����F���/�-F'Ҥ���T!h�I�j6'��ùkȩ�F|n�ީ���8�{U!o�'C>0�|�ݼ�D�V��i��yv�9�<45"�2u�J��F��@��Y}[���{��h���@|�3B��(�m�I�	�Bw'0�����x����~G�*7�T���5j�.�\aa2�a}�c��߉
��O"�zd�FW%��3�1�Zx�@D/�qq�NK�����i/�Ax�Z��6:�n�P�ۢ�\�� 6��!�,Ʉ.A$�&9�r�U�b�v����Q��-��<���/v�YJ�ZA�v��m���������A@P�L�ί��fN�(�a�9��AkƷ��JCR\/���w�X{�-w	�#A@�4��p�NEk��ܼ�̙O20�'����r!�ʅ�&}&u�=A(=�M�{��>�db ��(s�
ϩ�J��C�ܗd48Q���#=�����M���Ғ�[���%��ꈢ�/�ȻH��
'�qȡ�4�h�-$MUɲ��/� ��~Ol��&� �}K#���d�v�a��I���$�������rS�l��j���>2Ę��'>��=��% '�{��x��z��}-t���HضyCV+\<�:;�RN�#�!�v=N�UьK���a�vfX�˙L�����DZ�%B<�nZir��Nk�	ޱkX��,bx]�.P��9R��'�c�$Rذ��.;Eƙ�&��u�0CW�S�&�ԏd���F�>��sq����'<A�l�2�Zzt`?g�j C���;��PG��(�y*U ���y:��P#��8� �`ΝӁ`H/ٓK���<�������znI��e(�e��'��T
7�)L�!�?eN�(jRB<(98N �Oe���QXi�`)�����fvo8_٫K�����Y�>l�j��#r�!���=�ӵ��UUʋ��⩧�$�H��e�+:Bq�x 3B�7�����o{;)~�8
�ȶ��fN�jQꃓ�	� �1�JJ�6DR��w@B�WX_t�A��]W��̺$<��ul ���ת:�u�4���t�����eB���4��ҩ���m&e�c��X[(�.�P���.iSĘ:JV�˞�}��.A��%��|��|z�x����
�S%�ǵ�ڣ�-��l��>�ˈ�2|��5|=����y���af�F#����%)3�VꏈR,^a���&����1v7��1��vJT�[~R#{�j29}�9��V{4{G	���:�PF�`j5b�V\ 1��t9�� M>�v�z#���>Hj%g�i�6���t��P��{�N�����b7���,��\*�`vB��|�'��w��|S'�<n`j�8[�0:|����:�e����0*���W�p�}��?t����LZ���H��&�oY��<ukk���_[��`F�\�ZO���+�pz��U8�#����tq&�ݨ�a���p���Mo���&H{�v��L"`	c�)>�$ �Z|�������1���M=�?ܭ�5��/�4��'i'r�7�R�5Z��*�l��s�?��9	�H���yŹ^W�, �D@�����Ҿ|��ܙT����	�E�%$��¯`��S ʭ#E!Ec�)�ۆZ�*)�f���������{�u�GgO  E����6B���.0kM�5c����c�,��㮢I��߆���A��MW�j�ʢ`�[�.�L����j�����!����w�� �M�:E�̺��0@v�n�����	�C5:��wn:t\�!�t��C�60:��?U��`�d�eb*�z�ؼD`d��qŋV�j��cJcp{�r��^%�(	�:k%�Y۷N-�<�{���lA�DwלּF�S7��s��|JT^�EW�	��L�<1�;:�CR�9�b!���V�cJMn�]�p��FH �SJ�1F�sᙰ����&y���B��T�u��$	Og�$�\�����6v"2i$zK���f$��\�*�N'l�ϊ_}ɹ;F�ԭH�� ��n"�J��6�dq.���i��Mm�aQX�.�˰�'�0���VW4��ˌ���"^AK+3]з�좺kꙺl|g>D��7fb�J�=bS$� YZ�!����J�a{qI�
�Xj~�(V�n�t�0�����|��n3���Ai� d/�M�Ր�z�N5�f��J��yS��VF�R�W���U:�����о���R����i.!B��0M�/��e�F�p�j5{��������N��<�.��Ri�h�u�4m�a��9��)X��Ofo�iSSiɢ�$���c@t���u]�
�װC�Ԟ�����+.S��ѯ��~3��<?y���U;��ﮓ�� t���rQ���$���o�z�P���N<��'���ә����M\5��uw��n�^l����Y��?+�G@�6]@V�1�2R��)�n!�8�6P*�'zkL�ǿJIpBb�ʤ�ភY"Ps��K���.�X�IZ*.�]�?��6�W�6譝Γč����d�_�9.q�Al0Z����$F��=y�)ϕQ}�$K0 "I�:��|�oja�KձH�E�CX�IL0��2�1��j߁��Ð�e%l�[��Ph�s۵�7���@�D6樂�/����Q��lm�Q������P���4Tq_@G�V!#	JCr���0�MG�?
�ﴽ
�'Y�h1����~���@�����t�F2d�΃�D�Itl+���DX);�5E����,o �` ��f�,�՘����D�J�"��#$����I��m3�1=��@�T����V���ma�������E����Y �L=�jΠ�4�����:��uy�x�1�2��E� ����ӈ?�"j9��G��贑���AmؽV	�%+%��'v.����^�c$��ʹF�LW�w��$�#C��|�H��.6႘���M� ܺ)���i������0pָ�!.�Ÿ,�1}=EK,��������n�(�0f�X��;Y:���rf��������~�����x�͚��\�HHZ��rp�v�87̧6'(�(1$��^����h���j���Ṧ��DpBFw$���ZY4���ouc>�ڮ|���߶�V�>��إ�}�4PE2�yJ�R猾QKw��[�Ԫ֝9hE�@��B9e��H������E+"r�3��xd�����GUG��:T?���x.�>�a�I}V�c�þ
(� "��xdLW�C�3��Ƃ�ć@�
�@�����ӿ[ij��x~����j�7Pv>��'K=����),?O�ɐ��U}9�U�ۖ�\W�g���A�<�\/ӲTXZ�kt�����<7�`y��f�|AX�	P'r"Ϊb�f��(���|M��, �ƒ.���i\ʖ������-2��>���:��K��߸jة���2�*B��'ȍrp� p�}y�N�A(�N^�vձ>��& �G|s�F��$E���G����4�"��(��QP �}!��;6��e�����%����лC��
��{�\ux��z���yjU����K�\ ���~J��?������K>�ѧ$�v��a�(�!�̑�E�����-$Ll���jW�������a3�3�t��n �P�6�x��zX.�-O��Qo��Qb�V&XuZ�5+#��f,�9N�^������,�fSxҙ�����#�Du��B��&ZD�8��B̏��)kSTT����x��P�`UR&{�_4J��u.
������G�=���W<�&���d�����>��q^E�IB��~2��{tGXlgj�C��P���OPu�(�n!*���ݼ�yu�W��3��.�[/H`���Ӝ��/T�@���@<Z��Fo���I��e�<�S��a�
��L;?����|�j�B(�v ��>��DQ���`�Hu���v��8�(ޫ!Lxt�xֻj|�m�lw�;�\%!��=�(Z��A��,���$ۂ�'��&�iB�܌ �!��R�0�g���J��)�Q�8�����q;NA�%�ރ�I�ߛ����D�M�nD��y�r�(��/|��
�����������O��������j��Q��%��?��e��&� ߎ�H&�Ԛ�~o[C1'��|�	y�ӫ&�6��)�щlZ�� �|�Ehz����E�Ԏ�L�Pܵ���h�!�^�����ԋ��@=��+���~-�f��w�F����|3���w^<c?�av��9��v2��h�:Ś��T���R���j��t�؟��{B��X3�	`!�:b��=p�Zo�w�7>	k���%ߘJ�=��gC?6wct�}\̊�&N�s�O���\��,�qP*6T�B�4-�btMw�	�S`颗i�`%H�8v�4:� C��H|�����x!r%�?�l�yp��.�1T�?������L�Z����&�eY>z�u&�r���֕�;�\X�LOKQ�+ҝVz�`8G(�ӊd�oŸ�6a��p���HԐ���H6D��ӳ�s%���$;�a|D�����Z15�M����ȅa�}��ݓ�4V��'/��2	R-�qA0�7�r��E��"�9D��H�-��t�q^�S� �u��5�2��W�����T��C��2	4�X%��n���/�-�ʈ��\f���:�ہ��*����+���O����u�!��{� ��H����6aHc�A Fkh�ǒa4����Ԟ��,y��;�:�p���~��A@��,Ң;#R�i6׍�e�d�����~���4��DM�L��w��=v��h-���{�C5����=n1ì\���DM�1�o�I�4՝^�d;�b�J�z�����(�^<�Q���I^W���p���rOM%�;��u�J���N(�v�֙��m��
��wj�hF�a�"����^����`<P���N<Lf:m��R������+�7bucE���]ph��H'_J>����I��q�%��&t���&������pOⰪ���\�?*����6q7�i.���!R�[{=wp*���l�tj_�;A�G�/�,H��G �~"f�����qi�T�^!����<�lkX��]��$�'b�>�m 4Ə��1�X��A�`�]��a콲y��9WҪD��~7�,E�b��� ƣ�<�V��լ�<�I�ۥX�bF�#b�nC c0k�<��J���Ĩ��j��t�d�b���g,�j�5��R����/��1��':J�f�P�.:5���u���6��ͽJ�o�w!}�^0������F"}5%�^{�z�y�{k䉆�<k�����I��O��C�O睚�|�r��d`���u��dV}�+��O<�~� ��]�+D���9O����	z���fS�L�t~�ټw]�f��P�e�Jg���s�t���r�4Պ�'�̪����Qd�����Z��Q",�+��U7�5�*9Ѱ�U��*�^g(�������+�X���DV�л�m�����n�衑�ٽ��L�"J��b�Aݤ�+�����s�U������#X�0�Z��`8U�V ���6�=���S��}��6k_Y1�.Le�lk���}a|F�<�y�㞕�r$f�"�E/:�WR|No4�K��I���iXM�.0�}D2��M劅ށZ��[�Vg����`�h\*���~&7	|���DqpL�>�̋)Q70m>�(��-���W��T��Gj#�rO��0��bD}
]|���dY�P�h�pl��5�~�ME@>�h���T�	�ީJkK^tb��a)���Ex֪�G����"����H,��?�b�?ٷJ
�i�"�.���n��HP�1x|=@EҾ�H�V��(�Q��^�r+�d�~����LدXΛV��2���Ŭ�ua����r��_��gX�Ӄ��"š��������4LGm��	>u��%��"��.(F�ׄc?���HN��' �̲��$�@5��W�k]�.��I�Y��"�(h����Ϙ@m��v��Y���6��d����<E&K��Ӈ�N=gnƒ�9E%��G;t��5�f��F�ت���_|~����ⷖ�U�d\���Z;�rKR<�sG@��>�#<��Z�i�N�,h��j,(��6O��--���Fr�?�_�y��'���o��>ť@|
��z��V��ȉaڹ��I�4k�Z2kA5Jv������[p��1�h [�@�B�V��#6���r�xޚ&Y�����xu���!GЃ���T<�Y�k��.�@�a�\}�[
�t^"�bgd�c�W[�N3�!�1<@��K�/D�Eͮ��i�:hx�T��Fq��|�P1���B�j���,z�E�d 7���9w�|U{��!����㸙<�J/��oO�\Z�X�|#������,��A�wA�iP·qΥ[2f*�(K7��������m��5\eG����8�)-�F]�Y-�*���&ce�s�����2��Ea9Ȩ��{}ܜ��[(s�Ʀq/+>Kw� m�s��
ϟ$V�`�����4n��MK��g�Ô�"�z���q���`�a�eHq�>x�
݈��P࠵�$�#�3U܆�Y ,�p~EZ���ؖ;JKY�f���4v[���cy��U����SX��Pl˺7jҿ����8��B��¿���?���x��,zӄB-*(hɌPd��j�V!t���QS��;7#ƽ���bN^ך��n䗠�fN_�R��r�WD�l3B2�*ZJ���9}�?{�kN ���xӠJP��R�]u����6����.��O�� �:N�W�8+&iXwd'켸��>�24q����Gx]0f��2�4�t�p�g��PC��X��hZP�21(�*KHݗCy��������+����`Dtӷ �/�:"�{�N<�����deά�IxO�e�a��1�h�	
�jLHt�?9�~�dj	�(��r 9�8~�ZCQ��Y`_y��K%v%"	8���<m^�7#֖>o��l�2�f!?2E=@���Nʁ��_� $ݪ��!�CB'Q� �!U�m�3��i#�%�e)��8@�N���N��h�F���+���Q���o���DK!��m������Ϥ�צ�������B��R�0���<N��ت�e���U��>�e��"!�)N��&�Q�9D
[^�'�F����.�=��8����Y��m��|��{z���]ƹ��=l���ȣ� ��|9ɰ�z�����NQ=�*P�W�L���f��'���_����3��V�~.^:Ӝ�(��ԕ�v-�o�ÊD�U�T��RR�7j�j��e'��$�{=�ʳ	����`<��b�1Y�jT�������>.��0Ht��v�C+g�ڊ6R;�t2Q��%рN�����}��0,ҁ,*�gFB{�M��R~w5�S�ʢ��`��l8��@:r��vs��m٘2�  ���}�pw��L:�?�s���L�N	�~�m&~�Y�H\u�~��cQQ�.3\��O�7;+�W�z9Z�8M^�Fbj�$œ�a)�pj��CY�fۤH��{�V�s����$v�||�AN��)�1�cjM�����R����14���'�V^�M R�
,z�RF��i���R�9�eH-��oq^�� s�&�����x_�2�3�#)0TH�o�<�	��z%��ʴ�5���w�c�����_���|2W*ߊ"�]����7��q۪u�R���< F̺�� �6�n����k�:���Q��xl��5�,�Jf��M��	��n_��V��`�E��8䤘��(���`�}>s���n�4�y���)M�~7�Bu�f&�vߞ�s��ЎCCP�y�u6�n�Z��w%2��,�`���T�X|�d:Yb �zр׼�FA��&?�L)ڤ[e��{�p�P$r�(%�n���g�ЏfVN#��1�(�u%Bw� F[��]�ܲ��^�ͼ���+�J��<g�:�4xR�+���IX�ҍ6c@k����p#
�H6��J�Z��ɺ��&7���$�&oh����1��z���iO]��δ\+�U�;�O6ll�i��D��������*_B\l�9^_���;<�A���fHu�� �Q5"�5Y���Tq�{���?���ȖǕXt���Q�'ݱ]�H��4k���$	j�A�i]F�����o���2]�D,��7��W@tBb	v �Q��W��<��WI*�GX:{&��n���0&˚��8��dv���K��p�de���^0A�5P�M����o,��IbA��vb�Kk�:�ݚ�0;������H{�J��!�þ0�C|��_�F}�����{�)����VM��ģ�<v������f<Wb�5�j�ؚWZr�������q煥w�_yc��К7��*U��)t]�c��M���鵆���d'�ࡿoSż<��x�~������kI�K��ɥ?��{W�t�OfrG�ڵ2�����;�{6�����b�F��@J5�cg���J�,�^bw�R���k�+ʉ�,�V�����v�__�n�����h��c|L��J?�3b��ߤ3�S��e�s�:��T�ˀ�-�X�7Z �Pz��u���06��~�I��=��(�_�f.'J�l�:
��F뷂y;���Ǩ}$��"?ƚ:��-|��do�&�K�'����X�u0�Ea2x��e�M�?���� �b�	�H�}hf���1�7�����D���٠��g�Q�i�m�������F0�˒�T�G��G#�w2r��f0�A�}�
�(ֽ�LpY�qhgw���~O�q@��+�=s<�ބ1��gt�����`)�|IE3>p�b]�Ve���i�,MP6�b��:�xJaz$�E�Ig=�?�c�#��1�T�@��о�yV^���<-�-���Jݶ?�k���kLs�Ζ�wX�Ku���ߕ1�n������Mb���~�" *��������Xm�E	yn�aF����.u�V����cZ�����	���Ԟ$L̳�����;\���ڄd�������+�0(%�37���@}��b
�_k���0(�'��E�|�F��鞇n�'�y���W�;�Zm���f����Q�,,�~�]�=��"@\�l)Z���r&�1��w�lṽgRҵS��	v�h���j�X�|v�i��z�Fm�A޺W����~�]3ok:�>��B|AP��"V��򉼺�j5�4��2��JQ^،4�]�c�[z������h���@�bFB/h���v��y���(!�ʶ�[x�v6�[�GK�{�Tw����.�baC��}̩�#�`
"��Ed��~W��.3ޘ��k��@u��>��p͉#^i�x��5���v� 4�P�c1�]�23Y��]�W,�?҄��T�;`9ҹ<U6����]����P�<X�/G�JԐZRf�7�&�<�V N��Aκ<P]�Πtff_bo(Z՛��U�"=�H���T\ +���iE�-�u�t����� ��x�'�/,�F�2A'�� �%��t���}��K��(|��l� >�0P (��s��$��;���Hc'4	&N�钌���"=j�)ꖒ����L��웨�� ũ�9��
8����Jl���/����UZ!���o� �p�~@5��6��Q�Kt�ç�9v6rS��dKR�A���lSݣ%�l��jM�g�����I.�i ʓ�0�6Q��# x��^zN��-nk��Q�؇��V�;�K찃b�#Ứ"[�N9ȇ��z
�24�fIf��]8��-g�D�U&B��zZ����P��y!kI�G�=�'x�ݮP��R���^'��X
�P|:. �ƪKĈ�l��U�W2��&DJdb>��Sd�>��~q�&����x�tՙ2]�t��bgSɌC��L��Px�('y�*�I��r��y���!�"�����`�w��Ҁ�/J���V��<�F�|z+�uI�7xeYUv�L	&��p
��L��!?Ԇ0y�8jc.(jT{ T; �Q��5��Q	6�`����ߪ�v�`�8I4�W��j��q22F,l����=!���=�1O�)z��j��:$�$QWy]Jy���B�� dA�؈Ǿ�]d� �)/<i8��u��ѸN�f��3��-�ߑd�����Æ�D渘�h�)�h�.�����z�|]���9�&������L���v�eoްŵ�57e�i�]��Ļ1����&v5���)[y�0���:���t�I�'T���O�?#!�V�<|���zm1�8g���?ǆC�|ד����ov��
� ��=�vDْo��j�f�l4��c��V�3�)��Q^�0W�����o��v(Ip�wN�~T�H�R�<jþ���B��'��{8��!����d`W=b��Y��h���v��o5>�m֋�I������Zg9â6-3�tmDp��+�N�O��K�����,��*,��BVZބ�P#w�tbS�1��Mz�`�o�8��T:��e�{���wJ��b~dԮ"A�p2}�g@�?�psp��Lc!��&�Y�6�u�8
�T6̞���\λ�O�>+�18z�s#8��	#��/F�n5�ad�p����>���dH��a�BoѨN��$��|zd���a1��iMnS������s��򓽾4�':�����R�I���m�?�����i�J9��H�r=�jwu^h�^ .7���%��(����^)T�ē��	�%H�����#wE�>�.���+5�w��*:�����ڕ�����ul��4Y �d��g�6�����k��Sǈ��ht���,T�������z��)���0�J��{%��P��s����[��K�R�6�O�F��ǚMw���}��[�v�ftΛ;�I�(Ck�����n�
!����c��'�������BdUb�[�z�(O��魯�1@�G�=��xӘ�D�p�0�r��%�������*�N��
����@lw`��F6�d��?��M�N^�������~<��4:c�TRo�$�9�m�/c;*"�nzLp�seHQINJ4�����aè[�&j�S����o��i6Oد���5\f�u�ֺj6g�;i5���� ��)d3s*:�l9f_N�;7؊��H0�_ ޳�"\ۤ��Oq�k����h����"�`X/�����'X�H�#�A4<f
�g�� <A\+�]�1��N�
��Dg��77kz;��bd�� ��`�r�����#Ie�}Xճ��~n�v�0����F��GRΦL��d ����u*�7N5L�8�z��H_�翂�hT(���FM~:��,��V��a��l�%�!��0�V�}�F����\�{��L�o8�1O/���<�Z9��Z����~OL��;���W��ʫq��� � ��Z�zP��Uv���q�r%]`����J�o��������y�\82S�LN�~ĕռ��J���Ffw� 89�6[Wt��'r�Ѫ��c?� ���!S+�vڌ�2��=�ar�Kj5��E�&t���h^]����i�&-+��^��Z1V_�A��o��Ŋn1]�G\ؽX�L7!J�N�b�Ҥn ��*7�s�?�¯;��A]qX_�Z��<��
��(m6ٽ�Τ�K���?�:_O��.O�l��]ĳ�SF�R?y�������$��O"�f�:��Y|�7o;9�Kƃ��V�X�[ 0�-f2��@-�z�ǐ�~�]�Z����h��
�87��/��D��U�t�J�cQ��m��j�e������CKT"d-GT�#�>�r'�0M���v�
S�X���LY0��h����9�~��~@��ҳ#���+�_8s��ct=H���)Ly�E��9�}�W�����f,�=�u���5	�J�8|����d�f⺩�����1�Ly@{�|V�7L��L�H7��vC[����
�ILe�Α���/0������@��÷��[A���A�yzu"{�	�x�͸9���*Ivmiw	�����Жk.Ю��4wcu�2�>჎���(�$�wj�� 3�!:l�y���#�	�(�ޯy�kW)��M)��*J�A�t�����kE��A�'v��  n�ܭ�ͣȉ7�;�1S���f�Ԧ�N���~��$�����ˌ?\/Z1�er�W���ħ�2�����ސ�kHh�=�j"�W��Wč�X+Fh �-[��{:��^o��4>{��||��԰�BV������%A�4�n2a��J,)�oE�H�B[u���翳hvh�@�МB�����ט�5������'Q�Dd�x��6�+��G�\�V�T�tF��dO.���a�??}�V>0�
��"_�d�g$W�p�3٥K��i�@0N��m�:�'�d��iU�xO�����{nP�&��x�����8�6,�璄�?*���9-�<U�d�����3H���<��#/��qEB�Z����
�٬�����v�A	y�P���Λ��f���(�����~���{K�#��6�(\�x������ -c1���6� w��ܴ<1�L;����2���4���%��q�5}�D���;(�B��gC2>
� ���s*��ϕC��?܃M�4�W%���I�b�]���Dq��pE��'M.�֝qߛaz�4��
��Yȍe��p�:�U5���o� bx�~;0�P�;�g'K�Q駕�
v�D��o^��f���	��^V�l+�j�6�zi�ĄD���蓸���Y�g�x &�zɑ7-����s��"��V���$�>�;#�م�<8N�$�7�I���fD�O��>��8�D�^aB(�Zա-�:�[�u��kD�˺�*xI:�P�R�,���H��X��Q.�n�����xT��p�W���&\�d����X�>�"eqo{ލz���+��)28��t� ,g�(�C�i����/P3�(B.�*A���M��y&�I���^��lg2`� ��� �/�a��1��<������^�I.@�ei��g������
��L�F?o'�t8(j�O(%�' o�`	����QD��`�)��)�v۾�8F��r� \�LF����lH�)���!�$$=���DƁ�w:D��$��;�+���kBݙ� ��أ����~���b�)j��8v5�ֱaNRF�V����O�s"�o�U��6�D�p<�c,D����`n�)����z��{�a�6�����¯$�� P���_���e�Ԇ��X_IO�� �&ѕ@���[�zA�<�g�� KĄ�4�	���aњ�t��|Pz��()�?���!���w���2�ް*�8�%W����V=����V�O9�f���WEy��31'd�t0�^�G˜��
�v#��y�X��`T�GR��j����%@��M�{3)��iX��<>`r�:bx�l$���H�HH>�����^�{5���Qg�ˆ6KEt�Wx�[��N��`�D���,�*���B1߄o<wkZ�S�ʁ��2�`V308��p:h�	�V2�Q�O�I�(�Ȯ}$p�_�f;?�Y�K�oLF����&��YOE|uW�fcG�Y̕�\	�OeO+�+3z�}8x��$�`���I�a�P�pRm�9�І�#Hg��7)�Ls���H$�C�|�~)�1Fb�M)ά��+���(�n�|4|�'�+��R>_����舠R�_] �D9�}HcEO�e��^ã/ �ǝ���+�������T~���)	E�>%��.<β�m�{G����Ԗ�r�h*��^�ӿ�����g>�uG0S�) |�F���6rC�r5 k�����p�C�j�ODF,�'I�����K��丏�K�k�VSq������^i?�V�#�����j��w�MRBj鸯�����v�N�)����2C�Z�k�n�'�Ȧh#��"<x�Z�T���dpmb�z���0�n�/\�B<�Z���O-bp�0�r���%e4��&�s��q�NV��r�{�[��w�&�F?�����'^�Ւ�q�­��<���:�G]RJ�@�N�͇Eac6	���8�p���Hl
2J����b��������&e������@���7kOS����E\�Ή�q��6b67i�󅺠K������*��lt$�_黛;2\
�@�:H��! �5�"נ�բ�q|��/J����}J�X�E)�''Ӳ����4w�ǌ
���A�� ]��/�[�h)�ҐD��$7�X�6�7b�e EɅ��Ky�i�͒~I�HXp/�F�nTb0�XC�	u��Z9�΁m�U�,d�M �����M�5�-��S�Y�e�!��د�ób�AO�:F@�����*�i�>�� ��!.H[0�V��x�]F3bSVT9{��8��
M�q��:>�<<_m�}��K��ц��F�Mu���x�9�d`�Ud�����ϔV�~ڢ];3��ý0
-��g���XS��G���>~����(x���ŖA_��[P��~|t�e�r=Ч��1��[ܿ�3�q���kuè�λ�|�o�Ƴ�5~5��aR�bx^Xu�z��f7+ L��"�V:�<�b�L�n�!���'��LRx�J5.�b�N����ؗ�(�s�d��
 ����X1�.Z}�#������ɍ6ԭ���� ����m�_�1�.�s�l���NX�F��y�Ҏ�=T`$��O"5'�:~g�|��o�kQK�	v��JX~L/0�5S2n�3��|��|�,�XM���Q�h�=��!��7zc��D"����	��QH�:mo���#C��<S���T]P�G�dN#�%r`�;0EC�?�
��'�v$�Yk�h������~�k@o�]�>��2P��:_�0�Ttؑ-��xY)��]E�mԘ+��LJ���,�J$���0Q�J���.��[8�5w���fA1)ee@��w!cV�Y���c����[����5�E�{L��3Ό�+�r�/��6��d�Z��1���8���t#M"֚��3�3�T!⺥��mD�s	�������m.+�X�J��c�����E��:��c=7$�CY��_��|X<�4�����t��������ܦ��i���4s��վ��4#�1)Ē��E�g�ἁ���0n���JBc�D7E;�(���d�f��n��z��b%"~|}��5�͆c\'�Z��r�p��$8է�EQ�q�k�y��<hj�b2Vz��?�Ȱ:)Fc<��p"\�FZ�roa��>VƖ|�<��K-[V��:�r�_��lR4��2���J�	����㴰[pt��Brh1=@_B%� ��X�p�U�I�������xP���F-+GA��1*lT�{�<�.��a��}B#zY��
˟":��d8�W,jV3���!6Z@�*����k�?�iV�x�e����V��kPb	EÓ>�)4��E,+���5���39��|U����0��S�^�t�x<Κ/}��@ЍZ�,��R�����L����	ADW@P�H0Ζ�f3^(|A���y;�ڡ��%�q��\6�޻��l-������ 2ҷ��l�;���g2��,�v�J������7}m��:��(D)�b��>\� ��sEw�������ܾWO4?�t��|��!��|Ô_��Ϥ�'y���6�/>
���H��?���U��7�� ��~6K�����,|K��֧ǧv책���PW����d�j���l�.jC���UDĿz�������r����%�"�ixy�zDH�-�Y"�=�dؽD�V�r�����4#�>�N�	r�r�<�h�f?�F�e���*�D��B�/�Z�}�u߈��yk?ܫ��lx�#P8��R���nLZ�K������.�K_�`$��3\a���aW(��&��Kd��F��m`>{��q�"��5�q���f2kbt3y)g��-C��ْ��P�+�(]�*���({&ya�Wxr�.K��d�`u�����/@%O��<FC�����gI�h<eϜ��?��z�j
~� L�ߎ?
�?o4j��(�x �G���k��}�Q^d`07����v6=�8�������`���'z(�j�l�)�
D�!P�c=q���_2Q��)���`$ǫ��-��B8n� ��VؾUm�S�����)��R8���ѱ�N�E����#߇���J�9�DH��^���N�#�D�z�r�d�k[1��t��#z˾X�_y��P������+1Se�_��sQ��d�Ձ�&,x�j��[�}Z��V��u6�Ŀ�a]"Ҟ����Yh�̻j|1>�z����i�z�Ǽ*S�r���\���>�@0L��K=dn��^B��'sf��a��F����3L���w�^�~/�M����BvC�ԯbņͯT&��R��jybF�`]��]�{.���į;��S;`�,�b�i_G�!�F�N��>�6�Ao��6��rg/�66��t����@�N�"���8�H`@,#r1*"b�B P�N��w`�S�W�-`X8�R�:�Z��1�������#�Lٮ�'=p��[㝬�?wc�&��L��m�O�e&�
�Y�s,u�(���'u�yT\DZ]O���+�E�zJ�83{B?;��N��$3Laں�p���4�3�w�H"ý�R0K�]��p�$'�F|�7X�y��1��M�h��4��i 0�Igj4B�0'p�%�^�R�9]��}-���V��90	�H�79�`��^�` �x����{����ԋxT`����	���%���Iｲ���`�H+v�0��mf*�<m莆������Yu"�b�l� a���6͡��-�Fk�u��~Sr�̡Ԋ�d,��>��C�ᦽ����]�fR���J)�����U���rK�Q��O����]Ә�py��,!M-���|��7$"v�V���5п�`C�gF��~
n�d?�H��������4Չ��d�O#b��zb�.�k���ʦʋ=�ڵИ
6\pQr
A%@�9�a�i�`'�N�7�B�i�Y#vZwV��F�H��\܃�^�	���I~�{�><�~�:Y�R%��������c1�$�pT�NH��]J*��Z��e����&`fɾ	�0�����R�O�.�_F\�葴^	6]ˮi�?]�u`��wm)!�*�l�I�_���;-�؊�J�H�I �K"R�@�}Y&qU���?����Ԗ�ԫX���7�x'N���U�4��،��*	��Av]w[��)��� �ý�D�!�7mf�1W�bF  �.���?��/���(jI�`�X�W���n�mF0Wύ�$���J��\��%�d61y�A�5�/��n(����/ڝwf�^g�<q>:����a���E�ҹ�����!i��0Tt�s�F��l�{���e�B�粇�u�<׃9�x���w.�t圻y�Ȳ$��e��P��V�h�P�~0�7��F���y��b�]�M��P��y���Y�u���҉�S�)���Z~z���c[�<��<xyɶ�}��%t!�r�k	̖���W�R�l������=�ހ���A�5Y�ќ�c��X�^S$U�c4���.+�ۇ��NV �YΕ�0�nB���W�αDLm��J�-Hb^=���	�`:s��/�e�	���XLZ�bI��J�B���^F�6Ͻc�Z��n�I(�S_E��.�� lW{���?F���yL_���7$�!"��:YW�|:�Eoq��K�����X9]�0	^(2�ʭ��0<��r�����S��Y�chH�Y�<j7���c]�D]��������qQ�;~m*�<�>A����\�T�\�G��%#�,�r��F0����(D
I�B�Q�uY��$h8���޽&~`�8@*�̳YY?��!��;k:ts����)��Ed5�Գ������f��,�w�����+�dJr��U������dl���1d��@�R�rTrVo<�vX�~A<�l����*�0LD��·�Oih��ڬ0���'��y}�l�[����o� "1�#���o�
� ��m�c	*�2hU��.��I��c�[�4�3����̞�$/��{���ז���V��;��]_��w������E��^���>鸐ɚ�LU.���rE�����4𺃹n��s��"��V�;�?��_�f^HG������Q4~w=8�N��Aª\B�Z''tr�e3�_��=�'���ƲT�:�th1�Ej�~�(���>�K=�F^�p��7�����no�l6>1�|����kV{�X��B���|4���2W�J��z��P~�6[k`���v�h��h@�B�\}������N���,#u��p�x<��aƿG���v�T(レס:.��aT��}��t�
�ҍ"~�ds�KWǃ�3�f�|"@�},[0Z:��Zi��x��i���0�1�Pî�{������,f��������79� �Ug`��v����A�Oظ<	�M/X�;~VZcNh������:ɥ���AUpP.`Α�fp˕(7�ț����X��st���\�IZ޶/z/�-�A��Ņ"���Ғ����q��� 2R��1����.�g��}Hlu�(�/ڦ]ש>� Y_|s`S�ϋ�~��<@����4�<��!9�f2SLv�z�$�fzJ�� ��L������*xZ
I�����!�B�U�H�r�U ���~1���؂K�k���v��O��	؎�R��\���Il7Qj�-��0?����?�:���C��G�r�ݶTx6�%z�]-����x��X�V$8�\�v����#2v��_�N�Zo��_����f:;z�n���^<cD�ЯB�3Z�yᜰV���5�k:�N��x�S4PS%�Rw{�I�[��Ѱ!y�.�H?ƻ�b��4��
�W���&��d���$�x>v�q%ꭍ�Qbɘ��]N2�gTtn[g$H�C�oҒ]rP�i=(x�$*7�=�#�y����^݌��"�`0r�#��/����(�<��U�M{N���I�^e��+��
���	�
Y�uL4��?���j \jt�(��m ��Y�]��&TQ�"�`˂��Їsv��8z�s��1�ۉ���[�9_l~Ҁ��!���=,���z���m9*����$��.O#�X�B�b� �`
��̐��$���{)���8�|��чNe�̱5������%g��t�D�?��Y��y6?�(�_L����F[���o��s�˹����ؖq���	��l�ed
z���r��U&��/�%3�[ʠ{�2��P�����"�Z���e��P%���w|LL[zu�N��	YԵ���W�F�m���R���[�[)N�� �=?�C�<�6�fܲ��h���3g��j�B^�Ճ��1��@��v�Y�/�l�A�TAV]RʑjTd���+���s{)���'���\`��-bngd"^Ʊ�E��~��>�y ֜J����g�<�6���tބ̑�ZN�4�S���,>�*���B�1���w��S�\)�^:`�8���:^9u�n��R�����3K�pc]A�B?�{4�L�_���(&�y�Yu�%,C�=���}�\�sOR�+�=z��8��ZwjV3���iaE�p��*�/��Ҭ�H��q�mW�Bh'�Ky�$bN�|Kt6�t�~1��(M�#<�O����U��$l�4}�'5����R�3z^J�z��U~Y��Q^9k�H�J��[I�^y�� _I��*~#�f���B��B�T�����?f	�G%yjc�dµ������f)����˅��hb�*K��Im�+p��]!�u�UE�8� �Z���\�6(H����0k�%�����'����W,%����Ֆ��F�Z�����LbM��4�a.ה�ϳLR������姘��ޚm�6M���.j��Ҹv�~�߱��z��C��ڟa,,n\�������F���NU�D3�d���b�_z=������eT�8a���^��^�p�@r�`�%z-�������4NH^杣a���.�w�#zFǦ��I+���!^�]ّ'ڭ6�<Ӕ�:���R �����>|lc,'�=pqiH���J�,��5ʃ�4��,�_&[P�d�E��v�m�OI��:p6\#���ߌ6X��iF�ǅ0@�O���*˩�l��_u�;(<C��ɏHa� /��"͋��Xwq��O�e�4��/Q�3�X`[�RF�'�3�����4�>�8o;#AmKX]2�X�DkY�{��ZD�-7��,8buF� ��[��1��N����IҘX���
~%n
�0f|�?1��P|��7�ˡ{d�4*�z���5<Q�ĉ���[^��x�N���p��7�(:�"$�.2�`K��4cu����!�L�0�鶮n�F�̣�{4&���Ŧ�L�XX30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�#ڜ4Pz^�o*И�m�9	�|�I8~�3ݛ�m�}=�el����iJ��z�*��ى�g��ʅ1��je���*��7�]k6=�L?����:��:�W�Si��Y�IrL��m�u�?���D�ݑ[]Z�3��m��C+L�8��O��ީ";�KL������<�f^��h�nAj���I�^�j�:�⇺�:���.F�D�� ��]O�*�x�T�Ew�p6a�`���sMjLք�Qc=_>)��$�F�gy~�y������KE�T��S)D8T6&Id��]D�w�L7��a`�j1U�SjrHطO���dI��-��n�rj` A��d�[��Q@F���4�"�-,�*��~��� ��f��kY��B��=��t��W:rk�Y/��5���_9)�]Y�x٘�a~�� ���AR����6��ۅ���n�������8�R+���9��Q�����T����-{h<����������c��Έb7��̚�gQ�̦�Ek�p��G5�kNTYG��*Y5"M�F=g�T%����a�ع����q�Tq$n �c��C<&�!!���2`e�7�����nL S�]��?M��k�(N�i$p����@%��)-#̰�����֚`�����꩓Z�Ϲ��&"���o�ɕh1Z~�Ig�bEf��go )/��"(�܇/�p4|iJ�hm|�@��p��o��#tN���xO �^�Id�
>C�|"�!+�O�-�I�K�W7��[I�����#��*�#��|$��_���]c��p��w0��ј��#��w�S�ou$�'4���z##>��0~^�UG��U!�@n�k|k�f��ŵ\����b+����ќ�X�r����g���� ;[����5�R��V9�4%U),�h4�?��r�
�?t��?Y4v���U�m�>�C���%��J���v�2)��#�D��T>�#N�Pn�}o�棘���9}Rۋ=q�ݏ���,e`헦O���]7����*�=�2�h�R�;�e�".*��7�86�%�?��]�+�.D�W',w/w����L�pm9��?���D�N��OF&Ч�dݟ��b��L�{~��SFޝ�ֽ�+��d* �.^
~��e�jU� �=!��ޥ������P5�ی�׸�� �B��X���x �.Ek�:�͵��Rs �%P(��Xg�(C�Z�Φ;������Ӓ�_I���;���!���2(<n�Zڬ�(��l�p|�X��̐a�E��gH�Q�M���8��U����B�}���\Y�Q�F��%ngLn{�oF��y�Ƭ�#S�gc�10F[�\�\uN6:�+�~x� ��+?CZh���	�B�[pn�~�'���l�5{�mv��1hl����#����pY���µsѣPG5~�<�G����jM�� %������b0'�5�1�s�U�\6�=�^#�?��-a�歠���g�ɪGK
V+��\�}����fvY��jS���7k.��ʻ ��:~��À��{�v��[��Z��~�=���-�OqʯM�1 /Hm�rB�����C,ަ�Лb���b����eB*Y�Xa�s��b��o���nn&ww��Hƣ*�H��3A<7�-ۄ�]�[奮��w�6j|.g��Ys����QU8��<�=�)��vr��_�޴h?3�Q��˖Am?#�;�:��+���,�M��P���oJ]�þ��k�8���n@�+c�ڰ��+}��k<�v[Vs�F�:�8;�]��ʬp])�Z��lւs� �)���Lv��AfQ����x�J`w���|7A��`��,7C����ʑ�(6߅�&�D�1=�pIy���z�;��0��5��~C��]J�F����k���,�3��N
g�꓃�����F� +�48X��w�_�v�A��Q����y��8�Ф�amkY�����JEšK�26�=�b�p���V�Ѯ9m& �2�a�?9�%>ǂTG����#���_��Ӊ�9:T��Su���Gߋ�L�d���$p�	��!��f�\T\# ���意�ŇT����!�Y�f����ar2���h�.��'�0� JF���������L��D���#-MDŗ4B����Bʞ�-�7�/�����b�.�C2h	Փ�a������;�F)��/(0$�6b��2�2W�t�c�<�����c�?ܯ�����
{T��@:�i���pJQʏ����a[>N6��-fBg\w,���w��hό[�����cF��d�`���J� +�(���G�=�p���c�]��ms��D�t�=���~���p��;��ѫ�5�a���F�֫ͯ=q����ix�i��������[�/��ܬ}{�+$�#bE����f�(��i��x���jRಫ��$;	~ɢ�7�WhGR~�dqߴQ��i��6�I�m�cB�'N�O?��+�~��uc�w&�����g��"��y`e�ˈ��P������t�٥K������BT�6��jrO7�%�2}OC}G���bj���w��Fv��� �x2�:��rD���㐱y��	��ܣO��o���Z�*�y�� Y��v��R<S1�#����rp��OG��LYo��]��+m�<�xD3�$�4�)�1�w�q�m���L9 @
���4�3�dø3_(�l�D=��!LN%P�@���e�=һ��1��?�]�{��|�9� �g�va)޸d��"h��ښ�U^��q!���K�RE���i�����D�9>h�xkD���l��W���ʙ���Ye�8 N	sݯ1����E�����:��j뛲�.��N�3���`dQ�VRӨa�Iy�����Q 2G|��Sˬu��uf��a��'���0:u���JU���@uu��H:�KXG��'F�u�O�U�нh����g�F�C2����\�&�}eV�O.��T�<'����[/�)A'�Z�\�B; ���[`��?@��tn���)�Nn����M�z��4�o϶h�ܛ�!p�1x:��R�)ӿ�-����@��NOUI�?^�I�zɍ�or5�Ǹ����m
j4O.K�� �F^>�%��5/�Q괷�Z(8�<j����,�|"�/�����3�ќ��'�μ!М	���H�%��-Ru���8V�iTzV=�5N'�P7b6~������cf����8k՝.le�
,ٌ�[ 0o��O�ڦx`XXR�kk�b�~����<|67PEAD-�L)�x��Ν�e�
8Esi��Q���_���gET<�
�#�=ƓFb�DѤ��VG��]7c
���zC0,�M�V���h$�ruq�鰌ǝ�]�,��'�,�!��M���ϝ̍>��m���}���w>�lf��#�J�q�����G:�_��kS!~�r�������z��D�X�;}%����*��֨� ����E7rrAF����:�cp:����Wr
�N�R�~�}.�5Y���g:펟m�dL}^��J�ez`��#x�j���ģ���ʹ�a�t�"�fL�W�9MŔ&P�����V�4O9�a�e�i�3�&�ڋ;�U�<�i����c� :�,� 3HCi���;a���a��_�/L����
VAOUH��*m1�xں�Z9|t!�>*&�����$�ڤ��t?�~ܣ�pWB��^�6�\�R��S�M�4!����ﳲk�4f�A/S�}��hc��d-J�Q��������mY�V���Opɿ����U���3׉��㚤��V�";��lh��̇�ܰ��NQ_Z4�b�(�&G�Z$���}Q.�cU���x�Ս��B��c��O
"��E}o�B��aO��]N��Wh�U'�
*��on���T�g^dtm��x7WmR\���� ���f1�K�>�d6�[	���"����3���a�1��v~g��}S�/9[0��:�������������Č����CTt�S*�X+m]Ƽ��)f�6�&��;Ԩ�=Z ��Q�	fYruO\S����r�)-����߶w�T����@�+�reT��τM��#dL^�#���@ƿ�ǹ�q�,P.��3��Z�З��X�q��`^4�@=&��&)�0�ZlްT�k(��
�sT�;t�k�&�[m5*82��W�Q���!��Ds�;�fBš"J�@KM��c��g�#�������:q��8�)�6pM'Н2P���%'[�����r�[�?/��r�I�6)�4Cv�U��B'0��,8g�y�t��.�!A�3�C�4�v�~0Ƶ�����C��Ɩ��wPr�FS��j�Rx��۽��[����s	"�P)�i&���ĉ\�O�uq`�r�-��l�����Q���j���⸨C2�z ���u��Blj7#�-��&�zn^X��R*�0z�|��B,�⧷J8T��x�v��r �*7�9�G�n�<�z� ��xi�c*nϜL��A��k.����h�����Wq��i��;�eU�;w(���C���DbZ�����E3@]�'d�P$UM�V Cȟ6������'T!����~^MX\P�u_Xf⩊�AL�^�d��B����8R/ﰿ��4�M���x�5|��b.��[+IҔs%��������TIޜ�t�ѫ*S���4������6�u�ˠ^�a��9��ъ�o�g�F�""�I��������Q^��C�HFp�Տ�%���xY5���[�028���d!���Å,qƟ󪸱�4���J�u���V#{��g<��@7Js�W8��V���_y����:�j�wk$���M̫lA|��Qas_�d+�c��>����9	R���l�i���������rƶ��'rWw9м�~ڳ=�U����z�V���?ƺ�[����GSr���2 �Z�I���I}� �eo@�$�">�A��.b&� �i�E��j�L�I 'z�O�[X��|C���/:\��TYǀZH|��z�N�� �hEA+���� ɮ�J����̱ ^G=�X����2�b����R��y�z�f�
E��.򲫏n*�����<s5��I_�{�n�|��.ޝ(��4@屑_��=��G�)Η]{�< ?{��z	+�:U�����]�@;�T��F�4yo�D♁�ø�U�8�'���&�N/bQװ������0G9_=��l����<pD]Z��/�(�4����
yo��n�	m8�wlN<�rG�� .��a���o:���^�2�8	�]�Np��T��ZVwa�\�fH���Z���o`�;�W���bs~1C©i�#Yʚ���0U�����[�0���bS����(�twg��*B���]ݣX�8䱴Q�����@�麉MI�J�Ͽ�#C�a��Nƾ-�k�>w���d�E��d�[n*�ڟL�c��d�>�K�����$(,i�Gcp;�E��c'Y���ԵOd6t��x=v>g~ jWpI%p�z+m)��a��f��6��n�=�<,��p�&��ט2}�ʞ�4/{K��<�{>�$I�EPq�r���Ei�èjҬ��E�;b�$� ��2���磛�D��~��D�{���6;?���L�B����
�̻é~N�c!Y�����A�7ز�y�����(P5�=;q��m���3��23ب	��ƛ�j;�ɵo�2��t�~�N�	j&7<wOB�v�`'n�� !f%2Z����)�Dr��� �یx�.�l}����B�Ѻ�k{�XY�K�ό��17�AyZ9�~��d G=UY�s��PR+��b�	+3YPb4b����;w�W��W��`@� :�Đ�3z ��Ì ��K�D͒W� N��*@x�e����K�1,t���Y{�z�B`Ґ�`�C�H��sh���U��;c̬�Ks�r���r�43�����9���x�������@}�i����-�z��e1��N��կ�B��t�:>�l��eĵ�BwD�x��N��~3RtO`�$����I	v��K�� ����a����8u�z)��6a����ͯ6:3i�h�����u9�.:k��G.YF]�OA���Mp!W�gD�a-�Z�5�)\'�/}��1O�e�T�z �Q����
)�T"��Eu\azI�#q��[��I��@~g)Z�sn����Kz1���e�o���j�#������`�U�*뱽�X�-��0<�U��+��ݫ�
��gW5L���.�Ai��j�~�K4���ֱ#��I��Ŧ���SL�R��8�Tj,Fϼhd|���hQ"Ħ�B�a����ٽ��mq	EJeHLg��w�R������i��Vͦ�5�T����Oԑ���֤�c����m�ke�l�r�HBC��0���OK�hx�[�j�k>>��c^�H��|�(�E�g�Zp�	�-�R@�M��%@F��0O*%����>�Wg`C��u�2,�\���}2N�O���T\��n��E�) !����\����n_��n�L��!̰;��)��Sn�����?znˬy_|������1��h�]��Vܱ�hj�����U�`FkL�� h^p��5����K��j�ôK�U�3�4��Uïb2��S�/��8	��jIX��y�?|��e
*�C}A垂y��Mռ.]w	b))H	*đm�R�e�i!ݣV���5[q�������p֡%�c8 �ۦkBwXlr�o��� Z�0\�OH�"x��L�kY������e1�|�2�E.�[��+�x#*��?f
�X�i�A��t�s���EA>
mcj���������-�Ģ7bXx��I���,3��M{*���t$�mq�L?�ٹ��JL����,=����.��1՝�E�H'��;m��ы�>c����rJW?F�{P��ؼv��yk���	�󷢽��4�����/�<�ZX�m�%�O����û���|�+:�wr�>���t:x4�b ����Cr�x�᱅~w±��7�ֈ�:�쟺�gLj�'�풔��Ƶ�奇����-I٘5�La�^�"��i����9�&����9,���Od�aZ�����3'��s��;%�<�L��Y-Ӱ�� '��m��HL��<�;�J�����[�L�1��9V�-}H�^Nm���'�*9�����(ЃB������15f����K���pd\�`���H�?�&S�1s�a���T�� \��A=�A���[��U�������;�5�������m&�V/�g��gɬ�uI�,��3� �_�>�%���V��;1�lh��Ň������Q,�I���(�4A��-�lIb}>���𡽰!W��Z�@B�����
����&}	{,B<9�O �N�?�W�W��b�Y
��o���H���-�d���W�cg\(<L�����L1������dcob	Ӹ�����������$�1��v����ނ��.Ȥ�����Fgԣ!�YбwU�QBz˲��i�AАe��]s��Eݐ�#��&����='�̪j)	&��r"��SSK���,���$ݷ��G�D���@�!�rӶ�c���:�#�8�P��L����$�~ʶ�@VP{+�� ��ZB����#qW؛^�	�=3�&�~L�}��G���=kU�%�h�Ms���tҘ�&:*���28�RWl=!�2!e�	s"�g�s�R�NNx����My�ˎ��H�P��cA4�7q����vk����M8d����i�('�=��S(ڽ@^?|��_����ˢ4pj�UY('�7V,E�yF���{t�.*����k4��K�$�"�����Q�Qf`�e�u=�RF�5��D�RE���*�{�h�����sR�R��+l��g�	�-�)���sj`�ʲ-�O��E��>&���J�!M��zm��ق��B!�#$�ʵ�<Jz�1��Ɨ���dߏ�*����B����T�z���U����Ց��Cڔ{�I�C �(7i�l�*�^H�y�A��n. �&�<{�W�?Ki��ޮ�߬;���meCF�Doc�pH�ے��JL'�PQ[�]5�C5X���z�U^�Tn�t�/^�\2P?o�u,���`�AY7���H+�4����_�œS��2��c��z�jx�uЪd�
��W��s[��s���%��'��O�!:I�|B���ј(ے��Ha"����c�ub�u���^�]��m��w��u��s�^"N���M����o�^��CC��p�m�[[����Y�ëf�l0?l���q�?
�F(�,f9�ޢ�ݸ[�J0�O����Ѝ9�s�l�J ]�We#�Vvd�_|1��\`�we��$p��ڸ�ln����T_	�d8����Tf9�����l���ɸ��F�K݌�@�c�1'��o9��~g����z�NU�k�g\ �cF$�49s�54P 0�,�d�^)�|Me$�$|��.$#.�� �[�E�6@��3V)zS�/[��)�ic���-�\	�Z	��ZsH��z�=��=T��U+m!<�Mu���{m�bpH̾�N�7�X�
m�Ì�b�~�<zy})�f��E�D�.�
*�g�s�r�����sbj��I{0Q|"�{.�R&� �@�E�_��-�Ǌ�)�@�{�� L�=�'���T�U�o�!�X�m:��!���by|z.�F�Ӑ�Wr��XGbR)� ӹ��|/Y؝��oNӒt���i_ f�ICM8
�RJ|��!���G��^�<&�7�J�IX�f�S�쌚}S�#l�$�s��Pe��nl�� E	�0!X��)�=#}U �$b#u�U4*D����>B�0���Uص��>�2!}S��\�;k�q���"���w�m�9΍��ׂ::X�牊�V��x�5��ŭ;�X��n�=.���3���)!eh(�pd8riOM䰳"�Іqv=�hURC�>�ӭ�«p�/���(^݃�IOzR����N��#0>�`#_�YP�u\o��`��V9�;��:����݀�[�9Le�������G���"*��>�3�򯹮ӐL�e�U�*Tk�75�y6BW/?�e��.{�X�W!���!�M�Lwm�b?1F�D\iё@��и���ڳ�LH@�T�8�N���vx��n];��&�^[Z1�"�"j�$������B���&��e�D��	�� ���b���Ѡx�h�E\��K�1���<�r� >�%�^^�aa���arZsǔ;�6��#�>��l�n�f��u"N(�Z���9=�l�
��8޴={{��?�ʱ��"HU��r�8��ȁ��Bn?�O��YI�{F��%?I�_��o#�f��[n��-2S>��jv[X�\Fq_+y󏓓 �+�?�}�hWV�	'~@[!�{�O[뭧�l505��vδh�z��`�����Y`�¦���adS5�g����P4.��j���[�����'¼��b{ns#���f=S�6Ծ5Y��a��j�)�=��ʪ�r+�<���2e���э][}vJ���{���ڮ.y��q��:��1l��LO*v���[���7���HEО��q[�\��&H>m�c;��+|��'(���5���U,bD1}�6.�*J�r�@�̆�bc��o+��n�i�w(к�2*r���<h�%��vZ��w�?�vwM||���J�~
��Q��3Mń�j�)��#����L^ޥ�?D��Q�A��ۄ#At���*+{[,�|��A��Àq���Ǿ��8V �����+���>}�8�<�#�]FJ+	8�Z]6ޓ�]��)}�]�|s�)Z�iʝ'�ײA)�sL��)�`H�o�mc��".���C���;N,�r��6=��A�1.��pZ�͹�UXz=ok�����~�:]�Fq��|,�*3����[��̠
�00�4v����F�EB+�a�X"��w��}�A➓���kor�)���̼�m�|:�m�����2�t2�Α3����q��ݶmW�2H�x?��Q>X�G�Cu��&��_�_�Å���fT��uh*�G��L�������]!�e��x`T���z=��5B�XN���?%�j!�M�f�f��/j�r�� �]=��E��}�1}s��I��VH@)���Y��	�����M5��E���!�?��;%�-�)����Y�
bԅ;CC���ļs�b��% �����|7�0��Sb�y��C�t�~�3мjˬݤ�N�Y�L��I�E�L@K�V���J�	����a��"N�,?-7��X��w=S^�2Tι��[O��ڠk�c�jd�!���B�1d�(�G��p V�`cH��Wo˵���t-ke=��~�6p*�B�{,�J��a��I�7$`�m=��9�b�jqH3�|r�ss���XD/����ݻ�{�$*��EQTl�U"�deix*ب�MS�1����$�xe�3��xp��M�~s$u��"��6��w���7B��� p��̉~���c��ÐJ� ���ؓ��y���9�;Pv~��se܅���|R�����؉T���B�j#�f��ڴ2`&T�����}j�Z6w0��v�x9��> b�2�E��$ZD�+��;�Y�7�m<<K����0���Y�-E�A���18�]����C�����RG�g�Y��螮�+�#C�	t3z�4����"S�˂��7ˁ�1@{ (��l03�|i�m���3�DN��R��Nv��@Y$ke���lÏ1m��Nٔ{`8��o�Q*c�皎�I����{�h�P���ߴ��9I���6K4c���A�K��UB���]9/S�x|���Fc��)��J����&��"*erJ�N��C�&����n�B�MKf�#�c�t��N�3�p`��9���Ҁ�I
��lp� �C��a���n�u�ek�huਘ�Ͱ)f:&��S�0r�$��uڨ�:,!�Gm�F^��Obu�Ў~b���g����7��!�\��}���O��T̓s��3��l~�)Dr��e\B�3�i������]�e ��i�)� �nc���,pFz2J����@��Y�1��rc�b��!,��F��*�U��qhYU��L/V�L]��c�HT:5M:}�O���ȵj%EK����w֢vߐ���r��]G�s@	8ͫ9j����=��|S~)�ćCp�b��شμ�	�qH�z����BRƭ�ĩ�+i��V�d5E\A�GT%�PT��e;^c|���nr�k��l6%�ĲM0�1�O:�xѡ#�8�k_���O�$����|G(Er ��Ixg���Y��
�ϙip�IҸ�S��	�E��g
1W�����-�|��{x����7&=
�H���,w�AM?тBp$��q	����"���U�P�,�lnѩY4�?����1�������Y���>ؐ��;ұJ�aӿ�uԜ,9�P7�kd~ɘMq��fo#�x�g�w.`Ӏt�X�a�%Ż���X�I/��� ��eֵ r��ѦI:���&�b�5�r[2 %��~;�և�ʌ��.:�*�~�tL�@���*Ҕ֬�����K�����܅���a��4"KPܔ�Б9�F�&I�=��GO(aK����=�3kϲ7](;i*
<s�W���}�tu1 kJ&1leH���{�;���\�PߎLȝ�}�V�{"H�d�m�`B�k�T9Ma^�/� �4�+1��O���b-�Gʯp(p��O�
G�`��bAS`�����*H+��dw��PA �1����ə������졂Wz�2n�m�oVsL&��7���*�w�
J:�_���~����sV�;�7�h�\m�kЎ�?Q��'��O(�XC�K�t�0n|}�Zྴ��eu���BU�]�c��
���Vzk}M<B #�Od�PNT��W'�&�
��o�����R��d�+o�t]W+)�����t�(�j1_����D,Ԯ鷶���~��
˞��Y@[���Vv��~_tb�#v�(��(d1�_`��Vɭ��-�>?F�SM䙵Tv�blp��=l.��Y�t���P���i:l��늋�.�b�xR�x_3H�V�ga�j.fk=< �'���xt��&�fl���8v��W��рI��!\Gs��U�*F��12�C�M�Ɍ��`.�g�%�Z9��)q����|�����Mk��خU6��`�}'��f.��Tr?�I�~2��)�4���UP�M't�4,�)�yݏ8��_�����r�4*��B�2��8R��,�������/�r[F"��[��R<���Y#�֖�4�sɔ7�ST�-�p� ?]� ��J��`�� -1�켗8���!�.�`�&��9zD+0�9h�B���#��ɵ3*z2�h��M��Os��t��i*Bp��{b�TLؐ�<�!��.�̃�}t��2a���  c>�i1
*2�X���A���.�5��ǩ���W5��i��Į)vX;�a-��mOC�DD&=��Y7�	���;'(�-Ph���T<OC>bȗ\����T姬��^�PVuu#���,�A�J�S�t���6;{��������w��Q�\xs�����8tFF�Q;�[�y��%����+����IT)�C(��V̑xB�{�S�L�uEB
^/�(��3G��*Y��v��="Eö�$Re���^K�AC�vp^�����
�[=Y��=@0��:��W�}Ņp�=�c4���7�ݯ�,J0��V�g֗�+ ���|&J7r�W|߂Vm�T_S7��~��ɩw�e�$�G�Ml��ō�_���d�C�7���+9M�y�ּ�l��w�j��p�C<���@'6�f9g~�@ʾ�qlT� ������@��ڽ�؋�!�le� G9�������p�e��0$�z���!.&h ۣE������;az��^[}?���Z��쥿s�)�Qr����YH@��zb�ߴ`8���
+�'��dB/����9�H�u#]���XT�4���bQ�xԖ0�yt�|f_��E�U'.62�������� �sy�,�	3{Qj|�μ."!�k��@)Y_������)�ſ{��� *Z;�e��|�UC�X����/�q��py3������|�U.,��'�&��/�?k�N���=2yG�֗��X��Q�<��
]�h/��ۈo�?s�}����K�����-a����jǇ��UN2��xQۥ��pjG�w�NWv���3�l ��2_hX�H�]D� �����ﭑo�����Q�ѿ� c�Y]����@�g*�1\��>���g"p梕JG⦥YD���ҟ=+����-�%3q�4����ơ�˦7���RJ��
@1��Y3?6��([T���Dr�����N�>�@��,e����<1��N����{(KQ'��unXߋc,�m�.�d��h�"��Z���R�\KYKX��������'��9��9�1Mx�@i��zg�%5_��Pq��˓�?l�e�ȶN�f�J�.��R,����V�^��V��sN�f|3��`9���y̨v�1I.eu��M '!��fl����u;�S��-Ѩ<V"��ze:��ڙwI�����HЋu~P1:P�SG���F�9OO2в��&�Ag�;mr�ڳ��\�}� O�HT��C�Vjz���=)�����{i\�l��fJ�c]�4��	�K#Y�)���n���м�zV+ea��d� ���@��ER�#a�EX�>�<����R����U��1S�������s��h�5q㝢�w �J�j��$Kـ��¢����Jm]�뀷rt8�j1ǘ�a
�|�|�M�V�+ 冂w�|J����	J ZH���U��R�i"�M�i	E�V��5Cs��bk����)։�Qc sS⒫7k*DlZ&t�h$�ݩ0D��O0��xu��V�k�{�s��M@a|k�E�����xa��}�)
��+i�{ �\����E)
UQ�R�&��p�_��6HҬ�z7J�������,��Mc�Z�]�$�w�q��r���:�2�l�t�,%���E��������0���#�����]>������J?O�c����φ���k����Xɷ�Kj�㉁����$��X¯�%i�t��o���������ޟ��r����{�:`:J䅭��mr�"��C~_:3���p���:�i����2LRTX��ؔz9ŵ��t���8���Oـ�
)�a�o�"o�j�l��9L�&��-�b��{OL�a�҈�ލ�3pӲ[F�;8v<��E��#ӘP� �hU��H4ѹ�T�;�_�������I�L�\r� �V�� H��^m�'�u�9q�3����*��3��e簌��3�����pL���8kZ4�'΅S�g��I~8l�P����)'�A�2)��_��=|G��`?�#�V���-��o�m?nVG�䆝ɔ�y1�����$�9�&�C����V��;k�h�����\l���Q	�����(�V���R��T��}&Vʾ�w�	���B��B��d��jq
��t�zu}�sB$w�O��Nx��W����J�A
�A�o���m�»vӒd�hÅ��8W� \�[�w~���!�1k���,MdK:	����w`���پ�#����1�K�v������.a�1]���.ί�	�Й8��9 ��M��`�)��M9�][�K-�2��Y&kӜ�b=��Rz�	�r
�HS;_m徽D���Է�L5�,�T��F�@��r�q��K��"�#ٖS�8���4�7���b�f���G�Pc��"�Z����6q?pY^��M=Dw&��5�e��/Ƨ�%�k=4|�P�xs��`t�2�&"�j�+8�aWT���!M��s
���[���6��u�Ma=юmF�8�U�KO�_�q��
�k4VM�8H��G�Q'�rb��%�ڥO	?d�+�G�e��Q�4X��UA�'��Z,-­y..,�c�'��¸��4���3�
�1��eَ9E��MIm%�AFȋw�,+/R-e��1��P�[��1�s:�����ٿ�=�����{s�[T`�<�-����-��&/��pm��G��zU��j��B8#�n���lz�������������&EB�z��/�T�S)��ɜ�GԽ��e��PE�c���1ҥ ���i��i*㼧�a��A�9.�����R�$ʁW�k�i�W\�ڥ�;����yMaC�"aDWݍ�X�t�zG2]|'��}P9��E}�C���ȝ�=}�TV��\Jr^���P'�mud���AA�H���.�!ǻ`⭑p���H��z��b�Ax�'��L���YE�⼶[�-�`%�ai���	,�I����Wр��}f4I��l�z�]G�uv�^���n	9�_��]�3�[�t"6釫56[��Y�^�
AC+�Zp�Fx�C����G�Y�=�Nw0'���h�"���/y�l���e�ݠ{�J;�����_�xX�T�J���WMN+V^�
_d�>���H9�wM�~$X��,lV����._�,d ��������9����Wl�����.MV�tǕ�K�$'���9��~O����4�b�H�
:�Ń�O�'�K��*��B� �u���3��И�=�e#�$�W!�}".�|z ֎�E�Ɵ���^>��z;�[�;�Q$2��o�D��Ba��OWHq�Iz���% �=+*+Ug��5xh����J̦ͦ�x�nYX����wb0c�g��ye�fpD�E��.��/�O7-�Z��� �sJ=����{A\|
��.sY���@���_hRA���A)�؂{`	 4�-����o��U�Լ�	�_�U݃�	�����yd��.���	 U��,��'��!&�Y�/��ʰf)⎭�Gn����pm�WW�<�h�]��/4�Nȁ�H���0	�u���J<������!ͥ��EՖ2$T�g�	�k-N�8��io Z1��x������� {��4��\��"���4��w(�ギ�h��T5�~��W$����V���9�D��v؂z�����J���+��U��r1�7#X���"�[��g����JڻL�&��\X?5���R�D��Ż#��M�����X(���q�Ǟ2G��Fw�I�u6C��D��M��_��q�$���C�&��SK�Q�L�W�	��L<|E��/MI}X.�����Kt�� :��v��\���%��f�{�X�jF}2���UI���e���H:%�߮�1:��ʦ���T;��|������O'%č7�c��tق-�d���v�ڲ�Qv4"����ٳ���f�^�~�"�J��n}�A�f١D��9���3y����*tWh�4lI��Of}��K-�$x2���o���Xa�Rs��	8�w%ҏ��x^b��S��@*�s�'��tR'9��w2O����������u��$�������e�������h9(�Hx����dD�ZQ����.�E��T�eK��N�3�?B��NP*�H�Ƴ� ��G✒�3N���3�m�`�QZ `�K�<I��՛%�� ���{���tu����xh���Ig�:�vO�,'��2�=��uN�:�m�G�D�F���O'�gO{�fg�5���O��\��"}��O�2T�-n������)}i���Z\�-�*B��ŭ���:]�^���:)4A�n��#���bz˫(vK��Rq����ț4@�z��R&�W��g�B�J]�U�,�H�Z݅τ$'�865����q��j} K�}8ݰ�s����B�{Z�,�8�2�j��w�V,p|��;�c-� ���������ռ���	���H�$���9RB�"��i~��V��5�]�:C'`��jD־�c�V��
�k?ql��/��nj0�p~Oe`�xJ��|Yk ��(`N����|`�gE��8���Qx�N���6
���iI�ұ����6E�H=
���'�|p����T���ׇ7?{�£�$�,��M،K���$b��qnV����������,��B������v I��5?�C.�N">1$^˴��J��x�xXf�u�9�Iʝk}pO�����K���鍁�S�9��Xw��%�7��׭@���8�J�o��o�Ir�iB�s:�	�?�ӭ;�rr������~�eF�sw�:��<����L���6�e�OO��$�
��ш�hi��ռ��+a�w"�Pz�A��9w��&�"e���@5	OA:8a��j���3�ٲ�`�;"��<L" ���/Ӎ�$ �u~���H	��� ;�N�5$�I��L�΢F��V�V5Ho�m[vy�$hn9&A��(���n�)��N+P煻� 	� <�p�H��`����S����`�R�&���F2AIA��@���{��S���+��
��1m�C�Vl�+�ٌ��)��fᙛ�4�]���;끤���V �;�h1~]�����W�Q��O���o(d%f�D��IՅ}������1�շ��BH��</
��o�}���BY�	O��N�~W҂E��9�
��o�p������d^�T�c�W�;�\�,�̲t����1  s��|�d ��	0E��~�Ց$Ӿ����1?�8v(�F�^�YI��?IC��У����.`��n:1��.�m�>�ӐfH]�L"����'&�R(�^=�2�g�&	êqr_)}S0�*�So��Ӷ2���O������"@nz�rO?��@����t#���ft� �,�p���PX�X��]DZ3n�̷�q�?^���=�&�ՇZĖ��ƚ�Z��k�1��D�s�\to��&w]�_i8���W����f!�UBs�����ŋn��j<M�ǔ��#6�&��M�1,�q��+�"�r�`e�M��c����2ƥ�'ń�Lz���:�?Y����΋��4-;zU���'�+5,���y����XC��Ԡ����4�h٨�c�,��~�#��:j�B���"F��k�ñR��_�'5��ߎګs/�/�y0�"�Ƽ:�����pz`�%�-����"�D��W���?�̥`m�mzjp��R�BV��#���>��z`����͆Z���\���B����c$Trw�"�͜��X�2���E��W%�`� �E�i(%�*'��6�TA�.�C�C3�y�qW��i���ui;a=^�C��D?&����o�D�^�'*P�A񺒀C2a��}䂕���TK���}^��'P��Du���7A�����q[��\G?�� ��^ڄ�wL�xY8Ȫ����kJ�w^[Ր���%f�����!%I����S���u��.<|��\��ru+�`^�MS�ce����G�0��"�7�JSX��k^���C <*p��7�x���� �Y_��c�0�b���䂼�PU�����Ic���C���J-���<7_E�C���,�J'�W"1JV�)_y����6��~mwB�$���O?l+u��{w�_��d���ݜj��49sҋ��}lu�	&�7�C���) Ơ+5'���9:n~�K'p�֊�)�i� Ƥ�h�@zرg��R2f ��s]_�v��@?eY|�$���D.�� ���E=첶:��z���[�����룲�����������H&t�zp��� �ҷ�+��m�
~��G���_�K�[��1WnX���@ogb7�]�<�?y�V.f�X�E�= .���DOɡ�����sMP�s��{-��|�<z.�K��!�@O�9_��߈�ک)���{�� ��d�dU1u�>x/�*�I�~9���nyZ���W��XUT$��S'��z&SF/���4����.HGchF�'�ٓ�Ԃ<Z��]�t-/)|4R^��N���A	~e7�!r,<t-���8��6�v:����T�\��	 ~N�:�>�PZ����o���i�[��{����\���WvY��g^��3���h���5���Ldݽ&`���j�)�[������2�J�+���1v�l�͏X�F��l��-��-�J/[=��\����١�@��0�#�bÜ�&�'$�(�}�q+U�2|W=��I�ރ6X��Ŗ�����_妚q�����rC�r�����K���L���^L�A53�`/�S�X�v�P�\K��еV.��S�\��%���f��1Xy��}�,����I��i��7w��f%�c�f����

��p!���W�ꔀD���"��c�6�I9*-M�y� ��~yQ�vo��$��H�.�F3����w�� ;}��f.i���ٯ�C����m�*���I�Y�b�f�~K"�7xǪ����
a%�R���8D��'aa�mZ�a�D�u���H]��ccR<���,����d���<��R�
Q_W�8^�ʿgF���d�|��[�,����3�Gt���q�g%$tl�������JA֠s��t�������x�)�l/FlA%l��M�=.]�E�x39hy�wε�rv��$k �&��(BO��i������B�m���,�.���)�6h��(��oM��[��şY����c�4��iD^��.�~*�ƽN�ϱLFP�?���K��#�����3�v���{��W0Ϯ�fԋ\8!b
`u©�<�j+4�ܱ0��n\H�MP(�6�X|���
C4�b�{T�����TG��B:6	�3�iH��fg�W��	r�1���^�G(�-d��N�Y]\�g���e�7'L�,k�"���i�������Tz�]<�"��/�.B6h7�$E����`O]�s�b���(�sDw�eBf7��S<�"U���l^�ARx�E��DW�D���=���^B<�p���f��`YVe�q�kqbNA�U������̮��c匰/��ϋ�\�@
řB�n�pp�Aj=ٙx�f�Ł����V�}9|(��)��/59Rh63U���m���la�)U�6!p�DnJ ���R8�޷E&�dXR˔
�fT3�>��y��H���'�0=��y��:����yQ	n�>�U|��|�}�g��y%Mľ�NFK+P���)S���T\�� !����݄�7��O`�$��S��q�ݚ����d-�=nߓ�`憺������AQf���k�����-�w�������9����6�Ԉ�Lv�#_k���̽ډk�;�r5k~���VO}'Y�Mݘ}���kim���"8䬹=�A�P�@�˔�nwT^�G@1�Z��&�(�Zf�2�8�9�23�n��S����B�����i�׻�aJb@�������p�uH֑u_��y�إZ;'�O"�V?��2���Zuȧg|�ffo��o��"�g�"	n�f�'4����_�g|��/�'r0o4.jt�Q��ϰx .�I)�n
5mL|�!�E��(^�)�֢ؐ7�I�I �h����af��u�#RP�$y�?ֶb��1�臊*��0����O��#cB ��� u{��4P�����;>�.�0U|�U�c�$
!##�­=k����ܘ�����g�γ6��h33Xf���J!�����;RѲ��!�T�O��Zrܫ�)��>hN���V��r��G�����v#�U���>>���N������b�	�>����R��/�>:�#�L�P��o�H�~�d94���K�i#��V�(h�ew��F_��4���)*~����u�� ӶAe���*�A7���6ho�?�����4]�F/WGt�#壴i�L���m��#?��Di�������x��'�Yv'L��A�z+q�4�\�6�j�Ii�a��R�^z눉�j��Ԗ��U�ʦ-P��rJ���^ׯ�� ������[��xw:�E¯�q|���0�I�� ��%U_�G�y�Z�ӎ;�q��Ғ����\Ğ��ŧ[cU(�+
Z1{�_��l�Np��ﴣP����w��x�����9�&8��m���BF����Yo��F�g�%�2�ŵzoI�ف��>ƣzSx�a��x[>��\�;�5��D: �I?:�h�=�	MR�[����7��l)�p5�W\v���hC������w�Y<��㮣���5�I3�>ٔz'�!�0}u$����L9W'�6�H��s� �3`�=y������=�a=$��O���~�u�>4-<���C��m��v�/:ס����M�.�iF����:5v��cm��""vd��[�aɈǻ�4����q�i���cH䆽ɉ4�Q�;�ǧ�ޝ�!�r(��ϓ*b*4C�܍*�o���ݝ���b	��o��!n%n�wY0���C*�F��~+<N�a�{�2�ͥe��w3�|���ɰ�0EbQl�ٛ���J)���	����~w�w=?j��Q�ٶ�8p�#�����&�+a+�,i�0ާ�zæj������u8�O��%��+��ϰB��}��<�ݬm�F�K�8A]\���C��)#ǒ�s�j@	��C�e�}�֙���7`��5����Hyo���$C��3졏�����p"��h1�Ip���ɋ�z�a��k���z~�C�]���F�+�����d�*.���'
+���[�O��F[�\+���X��wy���(4A:����`!�E�Ƥ��m�D���1�!�[�X �2�Q���_Z�F�|_�����4�f�d8ŵZ�0į�&�� �V%�	�+ob)��q���ݞ�~ǃ#����wk�KJP� �/�W/�n�EpO��=�)5�&1P�A|,]a��|���x�W�R(Qf3�8�Ԭ~�p�L��X���H��� {��R��B�.�d�����&D���%ʟ�X:��}�x��0��2y�@`:��p��b�Q�>O���su|�g�Dy����DK뿣ʺ��SO�T6��p���X��;7�,*`��E�9S��؝�R��,od���-׳�n��r`�v�u����qQ&b#�+�e���'-R7M�~��TxB�ZW�hȈ��ݺ���^(|�}Z�k�~(�x5+���"�ՊYL���=��+�V�4Z������e�/�l�5b��xj��/��}ܬf {��$�L�E�@-�� ()i�t>��ق�j;���D$;2�ɢ��Wя����~��ߴ��i�H6�R^�m��B�p>�O���+@~�kmc�@�yA��p��"��y`��ˈ�)P�`��6�t��KyN��%�k�6+7jr���%��2&yCF�����j���w�v`5ވ� ��2ʪ��a�D⩜㐺���2u���#��̄�Me�*4���Y�q�v�/�Re[1�l��'��r���NDG�l�YoyϞ]�+m�]�xX�3ɍ�4ң%�1��q���͉LB9@
�7�4P63��+�3蝅!D=��!��N%Y�@��e���һ�y1�?.�]Y�{��_|��� �r�v��޸����(h�IB������:����<K�[I��Ji,��0D�D��9>�xk���l��`���h����%e��YN	h��s������ceճ���TT��G�N��3k`d:�V[¨a��Iy�i���� 2�������uk�uf ��j��'$�?:u�噂�j*�	�u���:�T9G�*F;�O��н�0��zg���,o����\�O�}e�eO.ET��ݡ��\�[�g)*=�Z��\�ko CU�[���?ɲ�t��b-)�7n����v�z�"��o�w�h�����^�1a��[�)�%�-���Ո��pU�Q�2�z�Kט�5���N����j4�K�[a�FG��%���5X��Q3R���n8��Oj�/n�,�,|"���N�����具'n�!Y)	��H��䑀�XRu�~�8�iT�-V=T�5N��P�6G=����>c����D�k��le>�,���$e0o��O��Ax`�TR
�k�˹�~�뽸�%|6 NEA-�L2rx���ȮZ
8�vi�I��ǣ᳤yET%
�,6=��F�uD:���0�Lx7,z�Յ�zL�,VM���$���q�������]�n��0P,ȁ�'���0ޝ���3��F��䛒>�u���LsJ��R�2���Ў�_a�kS��[���������Q�ϭ�X��J%Ԅi���֑��)��ҏE��rA����k$:�������r
Ա�{�~��w�5�F�e':�?�m�*L}GG���e�=��l��j�s��M���+,�}'a�]�"�o��W��9MP&P�����VZOa���i�f3�O ��#�;��Z<����D�c�� :n6�	zHl���L�;aa����`�_bDL��F���VAX�H��km1%�ں�9|�=�>�Ӄ��V�Uڤ"�盝��~%C��}pW�E�^�*6�x�R�US��4JR���M�4��A/�̀}V��hL�d6u�zG��/��]�m�YV�Kl���ɿ����y��8w3 ԣ�L.��C V84;䗳hǺ�����Q_���b��(����Z͜�M�}Q�c^�����Ս={B�����A
"�K�E��}X�B��pO��MN�g�Wh���U�^
*2`on�^����pfdt�
���eWmuI\�p��F蝺�1�4��>$�d6#~	�:�"�]�熑����*�1��"v~pz����/P�[|��d��oi�Կ����M�����O�C�MԼ,�X��]�e���6x&��'��N=Zi!���	�!ru�5Sd���[ժ)6y��!f�w-���|@Ĵre������M�S#dU<�#(���J��0��q���P.J��3�oZ��n�́uq�^4P�=&+&)�0�!�ZU�ް]�k(:��S�sT��t��`&��5�82�HW�Z΀�o!��ss���f�gš� �@�M���p��#��H\ǁ�q���8���6��M'��;��8��'[���x��?/��ro �62�4C� U��'0��,8�zy���.��Aq��C�Y4�5��~MCƵ#s��nM��o���P[+FS"���9Rx��۽?��[�!��s�j�9��i/h��BD�\���ޟ`���-����P��Q���j�>���AC{vz 
�uBl=#����zng釙{܆0��|O��B,�����T���x� �қ�sg�9K��n��#� �k�i�)*nR�L��A�%�.�@����VkWq��i��ڮe^(;wQ���T�C��Db�E���-�E��]��'d�P$~c��C�{��~ԕ�*T!I����^Ma�PBu_�z��AL=�����i�RD৾�r�7��2�t��O�C�U���5Xj��%O����S���&?�BsO�86r>s��r��:�s���NW�r'�7q��~���23�f��:@:��J߸L��멢n�"�W?E�g��[+%�(���6a(2�"�)�Ώ9��&MɅXǴ��#O�G�a������+3��k�V;�6�<?j��?)��@�S �����H�-��GF�;^���(�;���wL���Y[WV^#KHB�m�+4ڷ�9�{��҄Q<�����X�X96��8s�z�p�)Ȣ���0��XyS,G��R9l�G�њ:AlT�Z]M��.ϊ�h���NFL�~6�m��wV�WI���|�<�=ٹ�VJ�Z���D����VS1;���hD���7��ca�Q�굣_��(WBn�������}΀����ְ�^���B��}�/~�
_j��"�}���B�RO�\N �UWe���܏
g�oK��L��fd1-�@0?Wj�P\��^�W�z1%}�[$*d�&�	cb��ՉՄM:�Z$Z��1R�v�=/f݂���X�<xq���ˣ�.C�A+o��g�[��2�������]ڹ��j��&C��Y=�u����	���r�Y�S����f ��Fjf�w����ܪ����@a�xr�������hS#�V6��L���Eɿ�x���C(Pퟙ��sZ���̊sq���^1EP=ÿ�&f�|�!�׀m���k�8���)xsQ�Stb��&���/8���W��܀�HK!���s����v����^EM	Hǎ��������8�}zq�
@�u���M�kR1=��	f��'X��?A��M�?G���N,�S,4 R�U���'-C�,�_y����8�}!�`�Y4�U���d�Ʋ&��q�ǎ�%���>�͔xFp�����R��ۺ���C/�-:Cs�ܢ���Ŀ�e��<q��,��;�`��1-*/7��蒵�)������H7��z���h.B���#��Qзz�7��VO����y��2�Bi�駔�!T�� �C����Ƚe��6�������z� |��i; �*��a�	��A@�g.��"x�̚RWNQ�i2򣮂�;4l3�!�C���D�`�� ���"U��h'���P�����C�s��pI���T�.5�^j2�P��Ju�-���A�T�Lf��~1oΌ�U��mJ��l��
%xL#���������~[H����!%R{[��\���O�IMlʈ\ʍ�(<�%��Y������uS�^(���v�9~�=���"�R����h�u͋^D�0CӸGp���� ��D0Y�4A��=�0�Y���$���1��	BƼ���n�*�H5tJ���/qW`��Dƛ��@J�"9W��#V�_�|�z��w�4i$ �U�j�l�Í��+_���dȻ �0[��?9�q�/�lH\*YBn�ֳ��	���'O��9M	V~��C�Ǌ
24���\)����\�����̉��99 ��6���9���^e�#�$�m8�G.�� ~��EEp�I��\7z��[5y%�� �:S����+����}V�H��z[]���e���Et+��r��ܣ�z�'���M�N���Xm�١S`�b�Ǚ�4�y�f�%E��N./J�����:�Y�rs���%{���|�."���@b9�_:W��)+J�{�� �8�ͷz���UD����ԁ���筱~�C{2y������Õ7iUg��U+('T��&?�/_�ڰ'28�6�iG��:{h����<-�z]���/�-^4EB�G�j���6	���ʔ@<G�n�17��ޭia�ڴ����	(��N,�	�Z�j%�Y��x/Ζ���{����o���ʡ��^�
�*E�h�Gh53_7����9���S�����r� Ȃ�8��"�J:�+f���DE!��JB�+�Q�G��M �`J�쉯�ٿ\ :��qN��B��c���� ������zXp(><�q>��2�Ԥ��Iƾ�6�d�Or��l�_�h�q�� �n�7C����/�Kc��L�u���C�����^/��X�U4��m�K��Ш��q$\Xi(%��ffk�XLO$}ڕ��w?I�<�����VI%�����Q��r���7���q�݀����=�#�\��5"�cT=��-�.O��u`��gQ}�N�c�[Ÿ�����>����|9�}v=5f��ǐ���(!�����*q?�ܺ�Us�f%UK�V�x�W���'2��?MaX���}��87�FzP�� 4�tށ��	������R��$��5Q���V�ڍOYeRD�_*�^���g�
���;i���;�,��˦#�t��%���g���lȟ��1����y�A�ٮ�s�t�i?��~&�����|E/�Q2A8��Cl���xQ�ƦNl�+��ҳ%_'�7j����|(_�ɜ�WO�v�5pLmE��,Y*���C6�_�([ҔM�z'������cw#�|	a��z�Q����^y�Dc{P�(��� �0����3i����������A���~��!��N`�i�����j�!܄�P�#�bn�$�MC��6�#�ѿ��1��ձb{��DE׃����`6\
��H6ag����S�1Q,@��-q�<�Հ�<��Q]ob_�=T�
,�_
"�|Ɓ\��'�^�{F]SA"id/馬.uX�7V�x������O��u���V�DJP�eu��7;��<��[����e�T/�Ҹv�D��"�w�s��Ա�QCb��Ӏ���sCDV���>-b��D�袸��\՞q���2�B[W��������u���AIp��a=,�`���Ŕ��,�)k�l-��K �"�uR�	3���'�t�#���"͖iU��(� ���R�-���;3dk�`>��9q%�Q�۟���;HA�v00��y1�,:Cˬ��XQ<�o>"�*�n�o?gҭ5y8��J#�K���-�AS"�TTO��S��붼L�y�7Y�o`�=7
R'Sc
=�г֥GTsd��S-*�nR�`�/��q�T'hQY�⺾��x,�-�2*�M�h�g�K���3�Ո��뫺v�TQ������kP�<���5�G�~��B_:Y�mL�0�O�~�%�=�����p���ȩ���Xn�F��m�m�j&-���-�o2J�ػˤɼ%�n�vSǲ��2	�#H���r$i*����K@���Ӗ�̚Ec�/��b�ȸ��ԭ�ZΎ���<�"2CYƫ��PZ�wIgO�>f�هo*4Y�Z�"�X���y4��y��/|h��ZM�o�o�t����"�� �ۂI<~�
��L|�n!��M������m;7���I3����h1��V�#�W5$l���	V*�Gtm�#�^k�0Z��т#�,4��(�u�f�4���۸>'��0(ɝU1KO·��!�O�,k�h������R,Ϧ�|�栍���XY���B��Q�����;���䧴<���׀�{ܞ�)ֵ�hE�i�r�հ�����)��v�tU�-j>�����P�(+��A퍃ܻ���n�v�"�T>��#8�iP��co�W�Q} 9g�8�g�t\���9d��ۿDe�Ღ�o��0���D*�����t�h���i�(e��g*mT7n�6��?=���ǉ���9�W����7��' VLW+�m#�y?���D� V��E�Б��2��ϚL�@ � �ǉ��)����LS��,?^t�[4�j?���gB,�H켦�셋��;�3}�"h� �����F7�H�Kxj��E/P$������I W�U%:`�ڍ��Z,��;�������W_ß�p���Y��(�zZ����lƴ#�!�v���/�C�C�鬻����8�9u���B�1M���Y�g�FI�%؟+�uo�@6���)�)]SKr���L[ѹ�\�PT��	�h�> ��?���h��J	��[����î�`gMl�'p5�IKv.ۼh������;Y�q�_��: �5��0���<M�T��������'�A%�[��s<�|i�=���M3l���a�^���˨���� hI��n�:����4v��T
���.)���:h��ê�.��dv�x�[�쌈0����
M0,�1 ŇP��T�m�����8(]����%���}X�m��r,�4:��V6#,=(�'My˺�� N���L�:c����4'�f*Ǚ���8%;ό�uP	�<�L9��߿{�8�3��k����Pyω�����!�`��.�j�E|��y0�k8n7D M��~60�(��G�e�r���{7����c��g�Ą:�l6��0.�EHM��g\��$�n1�I��ܖ��j�Ș��I�t]�u۞��R�R1ϵ���"��*��G��ob��O�]b. "�W/1t�.��7��c�G���W��OX�����?��b�D��e���7��<��V����g�O��� K�D4"g��C������L����a��v�V �b�5~bɺ��0:��0���g��^����V��F�1�[�G��sE�bp�=tPL�a3L��ŨX���q 1��M��(��j�R#�3P���oa��k��8����{��� �x/R�J�@F�d�4�������y͙㸟�� ����S608�oyy�A:���� "Q�^Z>jUl�lW��gH�y����o�KF���ue�Sj:�T��T�����8%�7���`��R�S����_��Ud���-rMn��`��0�5���Q����.��-�m���������%u��tl��m&�����Bk�S���5���'��Y'��x�m�Ƶ��rS����z�+�{��pn9a�B���7�&u�2�u J2���Z�m{�n>`�S�ՀU�T�k\���iV 4�<��@�FPH��~�wB�L�(� /r�l�Z��G�|"z|��h ���8Z0�Og�xf�_tor���N�"�ća:P4��I|�(C����o��t ���j�� )#I��Z
���|
�>!]�],0�d���=?�7ۃcI[v��Ǟ����5
#-�&$�A�Q�"��6y��.f�ߡ0����ʫ;#>�ܨ�hu�>4K����>o�0p��Uy�����!^�݊]Ulk�]��7��:W���d��.ה�C�X��ʊ�3K���3�;�d��	�Ϥ��ȵ����)o�hI'+��6fr�i5�1�q��v���U3�/>ْ���JU�p*��If�$������j�>�;x#�xP�@oP�˘�*9��F���M���݁u �#��e�d�\o�OS��EI*Y�2����� ӱ�"e�*���7�&�6���?�4�"Q� ۠WB���J�o|ML�0�mk�A?�E�D=aA����k�O��NL�<��#���@�q�Ϧ�ӝ\�`�ϡ^�+���j�Ҏ�I?���0���w���l�M���j<� ���M@�dux�SE]�*l���'�� ��%�.��"%�ڝ�Zt�;��D�B�	���5��]���6J(�Z�Z�/l�Z��lxBN���<F�w1����&���&8�{]�\�B�%O��V_Y�BF�qZ% x`��P   7
  Z  �  r   �(  �1  58  v>  �D  K  �R  ,Y  m_  �e  �k  <r  x  �~  ^�   `� u�	����Zv)C�'ll\�0"Ez+�D:�Dl�&X��;O�{�'�jn�!3� ���ٻ�
��3Y�"`�j:.5Z͐�%F!5�̢�(w��p0��?U`���?MR�*\�!��y��F�]O�y��Z�LA6�ݻX��$����*�@� ,��냊�(���*��ea��)CN�!2EcR�b�L�ps��,���A�'���Ё#[�H�2��n�V����O��d�O���O�"��G��"H�J��UP���b��O�����%`D��By"�'�Hp
��O2�'~<��%kJ^�#�A[�>�q�P�'�2�'��'8�;b�'����O��I�{�
U(#�S /� Ҧ�� f`C�I�|��TO��}�N���(�F��O�I<Utȡ��?Ū��"�|�+�C��NȐ2	�O*�d�O���O���O8�D�|�w4cpd�5�Da[�͔�Z���;�v\��h|�V	oZ��dզ���4˛F+eӮ�ğ�����{E�%
�����UEz�ʅN�>Q�ӂ堰�7�J.�N�
�/�3�*�s@\�}r�<�	D�B�oZ7�Mñ�iA���O9�U�N r�
���,��"7D!���X#&d�3�`ӴA�"%���k[iv6���E��E�,@B��ߦ��ٴ-���.K�p��@i��T�n����p��4@���@��v�l�o�M��ׅ9VR���Ɵ%?0�X d�ե!�)���|V,�a`ɟ�<���9q��"k������2��.s��n��>O�$��$;�6�@!Dͨ
��T��&#V�010��$uǂ1[p�	��M�S�HRĸ:��0J_L=a7�N��?�2f��qt��C�I8$�<8 �*��.�B��O(�D[7*"ilk��<ႃ	D�:��!��d��?)O��$�O���z�8� -C�~���x+�ҟ�J��ޗ��)���P�g�t	[��.O�)�Ȕd��=[�m�	8�7��5R����m��j]T�1��@������M�2���O|�6�r�g,ͦ::=J1�9���	П<��f�S�Oޞ��vM
 a6B����U4}-�p���!�,
x��-�We vxxؖ�Ϛ�?	�����\�ݳ"!l0j�E�>��Pq�
AtTB�	;LNtL���ܹl:L�`F�1B<B�8Ic8�ɕH�F
,[ 6�B�ɮT@�x�ݝSN,��-xR
B�2+񐡀"ݾd�M��B��$)�&�J�A�j��<�R�&{����{��"~� Ò�j��p�3H�;K=���&�yƈ)�a3���@��`Spc��y�� =��k&��C��A)a�P>�y�il���ڨ6��<�U�@�yB��S���ӎ�4��|�T�ŧ�y'd9tL�e,"�8�R׎�2��d�+bO�|��٫|��[fiV��Y:m���`�'ަ�#�d�1L�5�	+Zi��'�$9�����_����D�=B1��'r�ɲ���}�h�S�ٮl	j��'	�hBF�|۞�qTkƚlCX�ϓzXu@�i���'���K7!�+c�PXň��R��]:�'�$޸U���'��)�62(Eb$�e���s��O�����?�p�`PF�<��<s��'�E�ׅ�
J�Y�d�X<�&l_�
�29�4� U>H� �ߧZ���a��dӓM���c��o���s�c�j�^͓!8O���s��ty��'��OQ>ŉ	K'��h��g�Q��f9�IB���㟔XKK>es�d��aV&�\ ���O��O�\�g�6JO1��v�IGa[�f�����Ѭ(Į��2D��c$�ۙ� �)%Hѿ~�^��*D��K�� �B�@��ٷT�E��+=D�ӓ�I��r}����."VI �:D� P�쇰;0��qQ*\T0Q3�:D�xzbb�	�>��֋"\�#T����$�r�f��?����@��ey��C�ve�G#Y���	�g�X�6��Y�*Y�J[\7�ު3������|����$���0CN
;�XR!�%@,��]���$!���&�T"1�zVг�'���y����+�����v
4��i<�>����IC�矬��˟�� ��.袸��*Dt���}x��Ɋ��W?DOb�&8jq9s"�(��dBܦy��4���|��'����B 2���9P\rԳq�F=K������xxn���O2���OJ�;�?!����4�݀ ���R5�ȗqZ��+���8-�ba
�'�(s�DU�.Ȱ-�w�V������x��U0,< ���~o1��]�2�������2?n)m�X,Ew&�{�ŉ��yb��O�����
?IlabB!���@��֔|��\��n7�(?��$�2T0$q��lw��5�Č��l�'y��'��l�y:��#���_���;O� d=r���s��yK8߼4���'}����SxRT�%�ĄU��q���=(%. ��&ŏTӆd`q���)�*T�ŎN�'R�����қ��'Q2�FJ]RRd���p`�Ca��'B��'$2��4��=y�8M+G*AqLhT5�_'TV��
�O5�wm�W���T$��I����'E剈\�j��޴�?����)Cg���Dۺ��0#�������6+���d�O��GE�nV�a�h #<Ɇ�I�(����d�?M:����m�V��S,A�x%�R-?QA�
��qRt��z�ܐ!AK�4����`�Mѕ��b�+@�jf�� H'*�Oȍn�/�H���)��N�.�P���& &�9U�6GfC䉃wQ��:T�ƛ�\�bu�A�D�"�?��S�����e8O��(:�Ȋ���4lZ����'�%Q��a�����OB��<��=2c��c� ��茁��+�?���O`�*���B����$�-@ODx!��þn�H���
�?#�\z�B��/�HJE�Ã`�
̀�����	;:�.���"�8�.\�aCR4H�8���O����6���*�<���E,8��l��i�Ǳ\�k+OD���	k̓Hގ�#�M&"\�� ��@��'���C�~I���?qDd��8�O|�a+��ÞGJ����ʜ:��ݺ0�4oZ�G@��'�"T�4%?I!˕�\��MJ �B�PC����J� ��8�,Vx��L,��.J2���#ХB���F|�^4SQb��zV�ݢG.�+@`��I2%`x��\:�8�+w��0��H5��O��d"���O��?�	:uONy����P�0���I�Q�e��;'`DI1	R�-O�c�B���zX%����O�ʓS�i�!���_"w���Ɗ�� m� �*�?�*Ov���O���	W�fC��J7P�p�1�-�)�M����6C�$�X�XK� �q7�A�T��ȁ���{�m��n��H)U`�'^Pm��O��M)B�8EL9ǔ}�r�	':�V���O�X.��L�/Vs0�0��G�JNU'���	X���; �ǲ?%���c�a^J��8�Or@�I�m.�@	g�.4�L�;�e�&:�&��<��N����):-�<�0h��C"�U�.�D��B%N.����O|	�Q�Y�t<��qf@)_�
`��t�O��z�� z{�×"h��m{�O�x�̊4U�BM�����i&x%B߸O:FP�Α5��tP!_*I�L�Od��4�'�b����<�URwH�j�.��De���ce�w�<� ��XQ*X�E��%�r�'�~�}⒨��iش�31J�q'zɳ�ă���<�&�������?����ّ	^�1��oC�IS%͚/M҄�aA%%����b�~E��� �3�	""� 0���
���4�[<;3*�#�Me��4mZ��|��a�~̧���'���F��a�fm KѮ1���x����V�]C��'�ў���H�I���R��59!�K�<AE�M� � � ��B4}A�,Py"�+�S��U�����5TzR�+P�G:M�CA:��U�I��,��쟤���O9Hxs��I.OD�)Ũ.T<���Z7.@\��Mt��eC%�4<O��R&�I� ���h'	A�j �as��Қw�F�	�N�P��0���r�DU�`�		4!��H��E�Z�v���&L&0U`Isfe�O<��!ړ�O�i�A��m�����|�TMpf"On,r5e�nwBU1*\�0�
��P�|�ţ>a�2F��� �-:d�b��:Y:x59��M�y¬̍�-*d�]�HE�B3�_��y���Nr	�"OE�ĳ [)�yb�_����"� ,	ݓ��T'�y�*��:����o�z="}�e����y�&��Q?���4� G���R0�hO�A��S�?<�GcUW긜��.�)
��C�I�*�� ���J&[��x `�zh�C�	�r���X�X������
��C�Ɏu�DY�#������+�"&�C�%�
EG��_���d��*�hC�I'TE�[���r
X-?Q.����"~R%ߥl��l��&<:,Xō���y��+`�P�z��W�l��ĀF��yr� �6>6܂`(����	��yBⁱx�x��(G'����〴�yR�͇G��	9t�>{�� ���'�y�hE�F�fL[ ���n�FaVD%���'}-�|���%�
����h�0�YF)��y
� "���^$/�(�1V�2��P"O�T�UB�F��p@��A	��P"O�(0�`�9 f�)�� ��!{�"O<� �%[�g�-��n�1c����'i	s�'��Y"&�.P�Yr&`Ӡ>�H�#�',Z
	>��b�v�b���MJ,�yB��<a�('W���hB"���y��U~=�d�2��X*���y���|h��ېe�9�$Q����y����r��Ŋ��{�"(�@dC�hO�P���&y�NX�,E?7~,��m+[�|C� N��Y�a-J 	��#�:=z
B�/[� ف1^�7��}���K�N��B�Ibw�%w��2Yݔ5c�f��[R�B�?_9���T"Q>�T�BtI
�}{PC��8l#V�k�m	-<���3UE�<=�>��
)'�"~Z��Ŗ'��$�� <X�Vha��6�yb��%t�p	�3g�FTaD��yB�X�����K `�����y�m+&���W���ܴ�0�S#�y���5rt�ɢ�ᇱ7���Y�yr��SV�݊i}��Eҵ�L�����:��|��k�~����n���L3�y�%��8�TI!m�6c}p����ɔ�y ��>4\�k��52K���)��y��)w��H�`��%�Z����y"#ۗIl������&��,�1n�,��>AƁBS?��L��v���r��{���a� b�<q�O�7!��� g�-vu��	c�ZF�<���Y�g�� ����`��I��A�<)di�<$H��q"L0̴����B�<����&FV��0��d��WlI�<�"�L'�6䅕F���҈�A�'��]3������В��]s$\c�
�#2�!�d�r�FBeH�8�z�R���7P�!򄎓I4Tp#h�3~&���ņ�nj!�d����H�h�%e�()=E!�d��[�^��%$[�:e�9`�-C�<6!���9
���jJ\a\��l*��N��O?AH�g��c�f����Lh�G��m�<a�9|n8�|'��"oAi�<A��K�4tx͙�9w�D�f��M�<� e�{�j��'K7k��PC�G�<��j߅W#b���o���$&HA�<��困S��" B�-)^9��gyB�W?�p>IdV�U�r8�B�C4��Zr��f�<Y�G�3���lI�VxI����Y�<)Ŀ_�cF�ՃK�ͺ��L�<9�JF�I����l?�i��
D�<��&Ƥ��@j  &ڶ�c�&[x�h�Eɹ��R�#�i��yUe�eW���d�,D� ȑi�1&�#�i��~��{U%D�<�C �*	���#��.T ���ċ/D�@;�p> -���Z @���&�-D���W�ժ&*1E��W (8�%*D��H�m��DU�AA��l�.9Zan"�vЬ�D�T�1<H���.�$i�
�,L��yb#fQx����r������yo���D�C6j�X��zCc���y2C:i�.4�5�JMzr��SY��y
�+� ܪ��1���c�@��'�`���۞\��b fY4-��@+�C�NFx��)O�,���B�*b�
�-�7^w2C�Ƀ$eV�aš� /�
�p��M+Eh,C�)� �����j�C��P�@c&IP�"O�A�`H#���v�pX.�s"O���O]:8�.�%��v�0"O�tIVEĺ	��D�T*T��l)£W�$9�,�O�<b �Ο�]��/X�ʼ�S"Op��O�g0$���+{�P���"O����I�LY��H�N^4=�B�
�"O^�����@&1h��P�C��mBw"O��g��[��K��pt�!�1�'���'���0\e}����V�~6�d#'�4D������	M�%���Ԉ)��1�(D�t�r���@��kT�/�8b�'D���tL��"0#&��5d߮�S��&D� :�朩 �����ԣ&Ԏ��0�0D�h�$;;k��!�R�\�l���!-�K%��E�tiۃtE�$�D0E��u�!/��y��ߏf(�E���p�.M��X�y2-J�<�&�B��J�j�(�q�O��y�愰aל��Ei�%fQ�Yk�I��y¢�x�l��Q�5��L�4���y�n@-]yzq����4�^93h
(�?)bH�X����t]��`^�B�2d��	��D�8���<D����(S��c"=d���:Ac?D��Q�G"3�,L���	� �;�h!D�h���6���Cb��4oi�];b�+D��[w��-#���)G�{t��@�(D�k��z
<���C�2�|�1�g�<��d8���6�R>
�x�����_�nijci?D���bN�a�Ҥ����#4�:RM0D�Lr�%żxH��K�.�JD F�.D�H�E�I�fi�`�ը�0�i��+D���):sizhJ�=\j��*5�+�Oj4���O�m��bXvS>���:B_@H"""O���F�D�g�d����>omĵU"O�4[SB	P�I�Ըk�4�t"O&���oӴ�48��
���i��"O��C&z�|���D����׋�y��Q, \�9j�8ِ5*����hO�U����	T`A�B�>>R�`���i� B�ɑh��qHb�"��ɪg��0<�B�	2��T������x�� I3ZB䉥S�x����<�~��!���C�+!u#�I� �l�8p�[+j^�C�I�E{�Ź�B �ZEs1&��veX���#t��"~&�G�A��(�&ϨT��dQ�ψ%�y�֒!��a �'H��`������y��̆!�کz$I�0DV��B� �y��ֺo��|P�C�r��bJ�yB�
5]	`��Dk?�t)GOY�y�+�Y� �Y��ZY��� �F������|bE��9<
0��������I���yE&.�
-r�ڈi�)�"���y"�K�i�ǣS�^|�4a�̃/�y�Q�RSLPa7�� [8=���A2�y"!Mw�|mӆĽO�ƴj0K����>�ǤOp?y�@��(x �G�ON@%�!)�g�<15��6Vr�:�햂X}8���IPx�<���@!(f��Ek8>����1�Z�<9�`Н^���3aJA�$�`��AMT�<��J��-rB鞴[l0��ff�P�<���H5|�Nɀ U�:@Ш��v�''�ۍ�I:X�v�
É�;�� �0ꑧ�!�$����I�z���j��B7w��1�'�q��92��X�A��n(E���� 
	kC�\.*\^}�����o���br"O�Z�����\!��i���"O| �c��/���I�<XpZ}�B�'Ũ� ���/�5q!�1+x��)�->��L�ȓ=�`�%g2	Rp� �c�e�$�ȓ W.���6_E��#g+�*F�؆ȓH/.�' �T�X�R"�
U����~U=b���\b��J=z�d��ȓ$T�I��$�������7]�F1�'m�I!�V,2mX�K����`w�Դ]��ȓ��ĀV��(���[c��5砐��^�i��.m."|K�fC�>��d��D��u�T(���A��V`%�ȓ4*�@SB��2�����gT��	���I)n��q@�U�&Y�TV��l��C䉹 h��q��M�4�H�*�[��B�	�D��`rW�,�X��!�$ UB�ɲA����fA�1����Ro͆Y��C�ɤGX����|t�h��&JQ�C�	��f�3�A��u�����Ԣ=�t�U�O�d�@@��
�:@��(ɮ"��j
�'ȼJ�K�3q�^i���{>Ա�	�'Ҩm���;R��[��#;����'�BY��"--H�Y�ڳM��	
�'yJ�����9�ޅ1׆�8B` %r�'�����d���g�̬Y��~@mGx��I �V�jm*WiZ�c��p�Μ(*�B��5V;���B���*EcP�-�C��9A��#�J�HI0Pq�LT�|B�� QgPD�0��
��Ha���5r2C�ɐ�P��یy��i�a�P�C��"(!�h�P�ǥy�t����
	����Y��yy���:1(c�,)c��#&��ј���!e�N��%���d�O����Oj����^q+��U�%�d��i>i�2OߨX0=�&OW�?�~���$2�e?Mb��4�t}C2�^��MC���"}��t"I	�xYdEs� �W��������Nc2�'�1�H���F�3:�&��S@� ~�@`W������DQ[�/��B�"��qL��A����NRyBgץxP-Q�ꈓQ�m��cS��D܋_|D�o��ؖ'�����I�W� ���Y�\!�r��U<g���	�' pѳ�2D��Qz%o�;�?E�D*G�X�����'5O��`�Iޮ�y��W�
2R�*�B��D�<I�0�i�����鏴5?A
&��}mdP"����@�$Ф`���'��)��9?yD�aM���`�(PU���j��-C!�޺5�ZX���Ӵ2❋����ў�y�����#����P�B�y���t�����<1 ����?!��?!����ԟx��n�L.D�zF�P=��%�򮋛}�x�Dβ]��m��R���3���}�o�;f
�@��(�2����S,�M��)|w��+�$� ���S��'g��"�]1AU�xKV�
W
���O�D��'���	�<1���qx��Z�Γ6c�Y5��g�<�qEʉpLB1+��D3C�
�P��O�`��4�����<�bɄ���9y�FNi��*�`I���2���?����?�)O1�@(*$��9Qn@���.A��UH�&W,g��A� ͸ ds���\x� �C& �8 ��q
�>*�V��U�qst���@�g��i��¦�"`I!�P�ɳf�� c�R:cJA��ƐC4`���E�'��J�h�0*B��$j|F�ۦI?D�{Yyl�ѡă�'I*����^���d��M�	Ky�k�5j�7�M�P�S�~�����XN���pL�,P\��'M"�'�"�\Ix�1'B�N�����O�)\'}��+�愳g�(MS��\8����J�qwHZ�_#��mZ�p%n��ƃrb��	��8f:�B��RF�'�~p`���?q��Aʖ$x�Ó)�4$�Nt���d/�O�C �`�R���� Ӷ�`#�',H˓%�T�2K�ko�$g�D�D[��'�����,|ӆ�!�a�<�)�X�I�O��h<萍qC��vK�E�O����) �Fij6��g����)��|`��B.i�`�R`[/������@�U	�16� a�T(S2�M3�$�[�O��t���-Lw`�T#���П'�v����?��O�OD�)� ����I�&Av ����D�@T��"O���A�!m
��ŀOuD����ȟ�P����/�(�*�/�5����Ǻawd˓Q�zQX��i��4�'t"[����H0���,A.+�( �fT�/�6|�C"��?)0�̹'	��o�n���	cȐ�	&M�i�
0W��'�X�ye�e�2����UP��-�E:ҡ"4�)r�^��
"p*PҊ��i�N�G�P���� �Ik����T	�)>�������*.fH����yB�8D�xtq��W�JD��g r����HO���O�c�`��_�	\�`Ib��vvԥyk�O�a7�' ����$F������a�����'���	4�ť�h99u�I5i��d��'�t1�BK� P
q4e�a����'�l<��茈1�thk�bD�faFI	�'�HR��4�"���i�\���)����#P��n�����	�|*1ƒ?	{�)W�L?a���G�L�<Y�Șҟ��I�ic�"w���(vE�!a�"����|2�:u�J���N5�J�y�cEs�'�h��� g��iEC��F�X-[�栋�JG,>�:�BG/�8g� #1�I�t���d�O����O��22��X��]�`Y�eA�ĉ�dj���O��"~�/�,ʢI؇KKp���7ƀ��$7�S�ԁ�<�� �-8���A�y�XkЅ�oyR�'��5s��'5�O�r����g:��,:�,�H�`�f&O��=��Zy�p)Pbfە��h��Op��O�U&�T�f�'��Ӡ<��� �, �9�8�c����AZE��4�?�3�'�y�H+�?Y�������y�	��C঩�f���v��� 7i�f�a���i�"�^^��<O$ASҟ�^wИ��s(�����5�� ��.q!�T�'��w���o���Iן ��⟀̓��m�	�fQ����O�b�@ٟ��ɖ^�<��	�<	�%�pnz�r����sc���tu����4/u�B��'3�9���?�R�k?�ޟ(���?��ɘ�.��FZR��e@aj,ƄЩ��Mi����ҟ����ݟ�̓P������]��u�φr{:`�"��	��HW*
�M[�'�T�0���?Q��[���'�R�Oh�q�'���r�q:G�A `E��ߵ	��D�%s���'���]��͓1�<�禍:� �?�1Ԥ\:(�T��de�> �� �4�y"E�ϛ�Cf�| ���?����?�!0�чF�� PV�������Ǖ�M��Ц�y����?!��Z���y��Z��ԨC V:���h�8���򵨖�Iy�6N�\�W� �	�b>�I�Y�Ŧ	'Da9�oָ����ȓ:��0�� [��h*D*#$�l�'q��IyB�'�U�P��&�\�`�nU�-�j�p,�I.%!�4�?Q����D	Q����i�ΐ(!>�>aCj�Lf�i����3�S��&�P֌���@�|st�+�/��y��
2R�Е�ټw �ջ�MǱ�y���7���{��V~�af�;�yr퀿X���J-|�h8��Љ�y��ˈ0ٱF�Ǥv�����H�)�y"��+ �̵ѩ�^���fؘ�y2A��4U��gM���xFL��y��"�yr�_ 
�PxN��y�Вs�jA�f��G�(���j��y2�V(t�A��햀S�z������'=�"=���d"wb��"���w.�A@X�"O@���ӭR�%�Ń�71�Q��D i4!p��J�R-�fLT[����GBKR ��i��8ǆ�BuO�9S���p��@^��+3�[/Z�,ȓ��A��@l���V%�I�'o�&��Mj��H�&�f-�f!��r�x�8����e��y��b
*܋�Րԕ�e�Q�+�v��5��F���OԬ��Կ��)A�S�(k�!�G"O.ab�>=�� h��w�H·"On�($�X�p����fIY\�c�"O��0�hYj�&���ŭ_(�S�"O�,�EBƓ�6�H$��-`�xx�"O�pk�FO�9��1�"�V7+�N,u"O�˄�]~�ؠ�6ff~��E"O����1k��yC�	�%|&��3"O̐R���)w1DM�%�==��R"O�1�NQ�Zp��RFC@���"O�P�C�"��i�4�N/뀍3"O,�K���([��t;T$�V��1
�"OFT�i��]r!FT�z���"O� ΁�� �/Z,���� Jd��"O�Ir�-]1&�����B"O�e��*�a#�K�D�:��8x@"OXt�nX(H.,c3�Њ<����"O��q%h�d5��ygJ�BSFt#q"O��#���aж Q�N�_ti
�"O=�����k�-2MPe "O�� �C�I(��Cg�Jj	J`"OԌ����%>:=�e��&3�A�"O
��U�{���R��нl9`�҆"O4��0ؕge����; .��y3"O<�GM�37�L���,X��;�"O8�Ȕ�����r#�5H���"O" �-N9|���)�a�K�Ndʀ"O^� �i@<�q���@
{� ���"O�̡���+8踴����QЦ��u"O���S"M�q��IS�S�Ga����"O�z�l��bZŐ�c��XO|̙�"O��c2Fjr(E*3	D>'&0��"OЁ�S�9z6�(A��N
 c�"OĤ�uc�7���*Tƙ�^"���v"OL� �`�8��#����Bp�"O2�C�ԕh�	�D	�5.��]�T"O*}�@�*oF�����^޴e��"Od	�W�B_8:uqe�\ G"�0{S"O��֢��n�H1!�"=Q�"O������^��d�ՠNB��Rw"O�ب��65i�Y��M-c�|
4"O<��%L-�l傳�v�h�r%"O�	Pĩ]�?v��R��1(���"O��ӣ 7&y,4�&��?����"O^��"C�&���pc�<h�AP"O��s��7sM.`ׯ߄6/Dy+w"O" ��f߻�8�0Ձ�=t�`X�"O��BE�pP�������o���8V"O(�`��Vg����Ɔ�s��Y�U"O��2}�	r���3��!85"O�P�jHh�hB�6~:��"O:(���(za��H�ɇ	rkdY��"Oƨ3�LO�9�4�`UhG�qp���"O����e��|y;"�^Tuc�"O� [d�+S�V!��H�r�2=�a"O�@�&��&oFa�qg8o��1��"O�Yd��!��4s`��3\d�|�"O�������z��A��I'~|ha"OT��U�/Yqr�Yg�˶_(�3"O�|��ēvN&=*d�[**r�"O]�%G��_Vmj։�" �T��"O�����>t�4$	G�h�r�"O����ijdp��jƒW٠=�D"O�P�>�X��I��i�w"O@��J!rO��nw2�"O|p����`��њ��WaJ]�"OL��dךa&�ȢgK�<F�x)"O.����Ǉ=J4��e׽Qb(�'"O��!U�������$�t)��"OZ�!�J�PD�*e���v�"O���P
� ��p� ��|"s"O�� �cڵ5��T�v٧Y� ��"O6��V�A������-[��X"O������_� `����=�l9�"O�e�F'Ӎ�>%�A��*\�dő�"O4(��\�=X�P�$�B�8�"O>�q3�P
���jV��P���8�"O� ������MS(԰3��0�&�
�"O�,a��8 ���Ł<<��C�"O�e��e�F%0��Kl�|qje.�k�<y�G��P�h��)� ��!��c�<��G:���c�?2��g��_�<Yө�n ��&C�t}��QW�<����{�H2��Z��e��#	W�<���D|.-��Iː�V��)O�<&%��[tBhsDM��"c>��.M�<���y}�E��'������J�<��C	���9�Q�9��H�A�E�<���އa��f�:/D� ��\@�<Y�H�tgX\�Բqa��a�Xv�<��h�"&U�ӷ�4p'�T�J�r�<Q�Gx�1�Ԭǅ.m�tˆr�<��e��/v���l��z��7a^�y" ֞6�z��W�8CZ��bTͫ�yr��$t�9Z���@�SW$��y�J�Q��=�' ��ly�e	7ǖ�y҈�=6y�T�4��j �KL��y")�O�e��Ț�v
L���ϴ�y�'	�TK#�Àr:�U���*�y���4=��9qbk�)�n�i4c^��ybɘ*-k(4˰�׻z��Z���4�y2�ֳmQ&�7>+~�q�R��y�*˿Y���p�Ո0�=���]$�yMe1���5�ۻ,��Ca�ʼ�yR\�xb%.K�VcF���ޝ�y��_(����!($��B�䘳�y���N;��Ȋ"�6y^>���ȓ� �c�%��ҢЫ142�|��D�܀0��ƛ1��;�%B�*��e�ȓo|��T�pe�ȱC/�"#�����|�F�pp�Z,c�)t�R�1��Ѕȓ��۰�W6(,q�ܶ:���ȓz���d�{�rE���ޚ]0ꍅȓ>�L��w�K7>[|h����~2��ȓX�����9>��Q�VF�h���#-na��"'w���#B�[j*Յ�C۪ �G㢉{B'�#�@��"���;�8�9��r��@��Ic,��2̛�N����+�G���ȓ9�`Ö�5z�0�E�-.��ȓ5����C-YJ|��6&�y�`؅ȓea�t�4�`����f�z�\@�ȓC�\�C�!�,���թ�? b�(��~V
��(.���T�ۄ_b�i�� 3:�@��J�k��Q��'�>=lFM��)�遠H�?<��(  ��4;����\{�m���%��!(i.,��x����u+O�9�8	*��&6�\�ȓm*�h�+�h�%'�C�`�ȓF�B�S �>m �S�E�%��d�Tչ���>��@j5NSV�a�ȓ	��@2G#֯A0Zp3E�ȲT񺠅�4j�Л����<HjX;�n�-%$��q�pX�)�r���"łħUY ��ȓ+���$��7KbphKaK%g�襆ʓ&O�ca�\)$�f}1��ޚp8C��"D�i�P�YE���`��C�I�Rpx���G�[:HC�	���d�=r\5�c+�+l�NC��:E!�l���D�0�*�$�X�1�2C��-r>ށ���9��Z!Ζ6"�B�)� �u07dLV��\)qgX�c�����"O4%y� �,f7���5�AC�挙�"O���U�Mbi���ˏ��e��"Oh-�q�]�s�؁!�(`��
�"OX��Q��&k��x���>K�"Q"O�l�6��:n#�E����/)��"O���Ӥ�咀̖7�d�25"O�X36�����	�1iZ���"O*�{��
�F���R<.Pę��"O:��p�.��X��9IDh	�W"O�@�ݱT�D�#"τ0B=ڸ��"O�A8�� Py ���#�=��p"O>��EK�r���dd�:dݣ�"O�
V��#}�&A�A��$"O���p##��X#CO y��02�"OF ���/lɹG"���8��"OV��SǘU�@UÔ�M
!���"Oʴ"����>�ZEnQ��!��"Om���y�� �AS)m�*��"O�@�d� a}����F�}qP�{ "O��z�`��:Z1�1�4jq��R�"O�9��^� ���)�,�z^`S�"O���@o��)��8&�,"t1k"O\	jQb4v���t��)Z����"OtQ��F�Oz`���
/(��XD"O ̠U�ך(� 3���1����"O TaQ)<��@$ͨ��0�"O�|�S��3rL���	��a2@"O�m�'���h8�5p�˞<Urp1�#"O�ei��\?5Lf|�e�/6f�1�"OH�6����|C��dY�M��'�vU)"�1Ҷ� ���{�� ;�'��Ms�#��0����&As�� ��'DL0!��8AF���+�B� ���'�6!��Oƻ�:��f49�b�'��I�蕏!jLcG�S^�):�'����9?8������!g�4�P�'��0�g����A���U�+�''&��n@�_IV�"R��#V-��(�'<*��w�� {3:Y��풛U���C�']@�s�C��(�6�6EU6Na��'(����FFC7���f]!t�hr�'ӌ�8a��J��h��e�@�~=�
�'�$�r��"���SQ�/$��	�'ǜ�� �r�0<q��:l�L��	�'{H6��F^�I����Y0
(��'
B<J ��J�:%n�%O);�'���D�t)��J�p:4c�'�t�HGON���;Q&�2V�\I�'3�jJh$�@��(~Bt��'���P�n[8efPiVn��#ߺ�'\.�hd�"�
3 G��t{	�'D��B� E�r�x�%d���!{	�'8lE0�h��Ś��ɨh�U+	�'Q
D���M�@L��	�d�s�'�����6p�b�8i�C�'���0g� ���HI�w���"�{� �+f�����)k�� �4jO����6E��{�>�q nƦMX>E��\�$��#5D��<�2M�+w�`��X�80B1᜘J~�"�� +)�B���y|.L��D!f����R��C�`�� � L�Si�8/�T�p��QU�؄ȓp���	2Q/:�����BZJ�	�ȓ"
�#6ϊ(����N�t��S�? 4�(��M�{����A��U~���"O�x�BCXt@ x4JLZdH[a"O*�PkV�1鵧�Z娄�"O�{�K�N�r S���<�jU�"O��"pcԪL�`-�E��F��12�"O=(�#��r���%�\�'��!k�"O�ZB���6��< ���4)��<@`"OdHJ�%�!z���Q8;*u�s"O����ʦ;t���/8&�)��"O��9���rjVe��4��p��"O��Ig+�Z�48�րj��ٳ"O�л1�S�v^SGB�'�8�%"O�X"EI
[L�P����|���"O8�ru"A'�4���ړeX�"O�Q9 ɕ6Auz��4	F7�ԃ"O>T��<�<x���Ҵ>0܁+�"O��@�������+�� ��:p"On ���»	�V��D�V�<ة�"O��Afޣ:�B�`�B�"����"O@}�Rƌ�,�l�xD�˰HƩ�"O¥��ȳ0A���E��f�p�"Oj�3����^2���t�J��!�"OF<�B�ۡL:��1A�2��D��"Oz��w��L��\��6�B�Ip"O��,8$T�0�J�8X�����"O��ba�6���ȓ�=Ϯ���"O�HvɆ�*��I���Z-�*���"O�d8��ѯ~��
⁚������"O<�eJ
���)��,����"OMq���A:B�i�+�D4u@�"OX��$4K Y%��8�HA��"O�(���.�4c_�mS\��A"O�Л&LBx����G$]�6�@�Z�"O~� BH�
�tʵ���F
$)�"O�8��$ӯ~ۄ@��0y�5�"O<��c��<w�| �C�� �i��"O�1�.��OA4L�RA�5�*U�"OF��s��)Kv��@^�h���"�"O�հ���"ك�mg^y� "O�<����jn�y7��3I�QR�"O�<ZфA�C�> ��!Ɠ�F�P�"O�u"r�U4��< ��
=�4$�"O�	��G�;���g%����e"Or$�s�%�d�j���!n���Z "O�( $�3Y@�K�b��oĚ)۰"O|A����[��	k��F }&~�HC"O�ن��#"Phy�Go@�BkP"O�� �lY�B	�
"O��2{� �"O���@.J���.�����"O�x�S��� ��y⁤?1!jay�"O4�p@�P�D*,���G�bcq"Ob@ABb�G6Z�rhف<���4"Oޑcw�Jr ���W<�P[�"O��҄�F��Z%�
D!�l1"OX��E��}
��',��S�"OP��+
�b�[ �R���"O(�x6HM�>-��ȥ��~�.��w"O`5���ۘ~x�P��� ���$"O���5f��0��5�p�Њ�*��"O�qCo�1@O��^���6"O4���T�[����� e�HY�"O2Ũ�L��pvl��	�1�(�!� �jx�!�I���!��.S�~�!��6�T	ӣ�K>to���t.A�~!�� Lqv��n���c�k
�5� q#�"O��9Q)�s���X=(� �!�"O�)��oZ�=tzl��$��bY9�"O���͛0(G� �aM
�`���"O:|�6lS$w*���G���{�(y��"O�ܛV���[�ͪ�H����"O ���a\�R�x����5,�H��"OZi���^�t�V������s�\)�""O����&R=QqW�G��Y�"Ox����c480!��U#�8�f"Ot]�gU���{���.�(!�5"O������,=�r���R	^圅Q�"O��Yp,��f8F�#a��Q<��0F"OR��Sb�El ��!Һ_#��b"O�t���̔2k��Ӈ��S����"O"��ꑢZ��EI1AЬm��Y(�"O\��R��ed�$@<Q��xAp"O:�U�;=���uL_���`�"O�h�F/�6*�r���ٸ)�z���"O��Z!�BX�����3<�X5�b"O�ə��G�]@ťO�=��H�E"O������ў1��E�&7lƔs "Oj��Dʏ,^���#E�tFR��"O���Ki��.F��U۲"O��30L<�A9�׬�܅ �"OnA3��ň36���Gc�!�
��`"Od1�)��WݤԂ"���b����"Ol�3�N�4��1;@�K=���j#"O8���>h0�yPQ`@<�$P�"OT��- <]���V��@"O=��.W4�\"6f̖yd�"O��D�Kb���N�28�q��"O� K�`��P�( �s����DA�؟H��I��.#���i^D�:�%ԁ��5��'%��0����{�Z)j%a���(����Y���p�&�26��;e(��Y,�!`A��j�<B�Ɋy+�#�JG�A��� #BN.TR`7m7!$^�
3��?V�D�S��M�w�C�F�|DR��W!0.z,��J\k�<��
N��p]k��H��0Q�	^}��J+�򁒀&��:��x��Q�&��Li���w&]�w��0>�7ႜoI��G�q�RlzA��#�Buۂ&��]]�X�&Ն��?�F�C L�x��!��|[6���I�'���3��� ����KTWx�O����ڴ#g�ԛ��[d��@��'��M�B-uʼh6��O�qђ�Ȥh4��P�ě� �h�p��h��$^�v�}��0M;~=�� 
?!���1P��@�G�)����T??�`��,4�pE�6H��>�L����ϨOv}:$#Շf��Yx6f�6$l�� ��'O�Mӂ��T���p@2!W�{ 5ӄ8����Ln� vA�G��~"˅�iv�C G�W����X���'��x��WΦH�AU \^�p�~���K4�.�*����e�a���w�<�eI
�Jq�B�˟iLܡ���і�r���l������:;�J G�T�O��Z���+LO����3[R�9�1"O|:- �-X7@��_Ũ�j���3Qr!F���5�Y�Q��&��<�`D�#���=~a��K�!	�<���,ut�2 ���@A��)��Y1l�����x�Qb&MY�<��q���h��XXԆ����#���Q��1sq�'��&�������O��<��OX}#�O/��$ѷj��e�'�&^���'�D���W�B��ັ�� �l!�O:��ǭe���hi��~r�LM�AQN�؄XE���y�MO:0��͇�%��mh�	��MY��Xl��.C���'�X=:��VZ�xXF�W6\s��#��=b�`���99S i��)V�'xP��
Ԍba���7�f���"��W�4��V*Ž+#$��'�7�"�~DK�@_()%q��-���5�*QW�B]*z��g"O� �-����yYh ��8P&�OT���R;@h��&��}�ԣ�X��1���($�5Q#�	f�<� �ߒIIDH�l���MA�eC���$��jra؀
;<OX�ha+P"Q���Z��h����'������V�M	f����!�� �Vg6J��B�		H�����"VF��pl�8w��B�	�b�h� ;?�ȥy�eՉv�B�ɴ?h����$*G������9bg�C䉓#�b��c�� @��9��N�x��C�	*S*��3J�,2^�����Up�C䉈x��)�qk�"l��逫�m�C�Ɇ�B;s���OH�Q�E�;"�C��G]�qg��v}��0+�5/�\C�	���d��+ �x �!�͋?�B�	EO|���*.��I�X�C�ɤl��	�����T�X����W%BLnB�I�z}�%sC������g��+�B�ɺ$�hq�W+Fy�L�� R�[tC��6n�&仧E���JՉT���~*�C�I&!�4a"�ǆ4�4Yh�j�8M �C�	�Kk�E�ś6��D+q��l��C��3#����r���|�͍${|B�ɵ^'z�1T��*#?*Q*���HB�	d����'Udiq&cɒ��C��/
l�%���M��*�����9I]�C�	�BK�!SO]�/\29z�A�pG�C�I�U	��c`n��]'i���s[C�	�r@h�F�8!�u�S��^��B�(:"��%`��IR�h�%@��C�ɝA���s�+�kJ@,Aw)�6Hk�C䉡p5̑����R�F�\>�C�I�!���pϑ'\x�-*��	-��B�	:)U�   ��@;���ƈ�q�B�?=����A�R{if�CW�F<rC�	�*�xܢ�D�'N�T��Y0�2C�I�U`8���/M�c����;6"C�I�hZV�q��]�E�bYY��EJ
C�	�+Ը�TjJ�x�p�+C�[�K��B�*l�P����U��XE�
hlB�� \�,��%m��=
���FV`B�	;#�^��4�W�Qy��҈{�&B��3I����Ԕ#W�IP��  �B�	�`n&�㵌J; ��@Bf��B�	Dt��# FӔ�^�Hā(K>xC�	1+�h6�R�5����f�"�B�{DR\����дp"�F�lC��8I`	���J���h #�̩za C�I�W
��XD0�ȰKr@J�lZ�C�	�f���H�cD�L�f̓!�(ZݼC�	�Y��D���3'��j���\B�	�̫B��)`���BB vB�30�#���J�-���h�C��#�`� ��(�|�dʇ4��C�9����V���"�VE�5�jB�	�@):h��ĈA�r���@A2Il�B䉈aB�蠅�s��I�2K�oZ�B�Ir�����gN=}`1�����
�hC�I�h�����
�
@�+J�2C�	pO\���
����T�H�U�B�I*��h!$$�Iqԍ��1D��B�IU$Q��a��!�DB��O��d#��ͷ/�J�� �0-~
U
9�DXyѢ��6�֔7��� kƷ �!�d�&d)��@RI�XZ������!��K�m�|��'%E	M9�SSh �T!�� ��%�$��ղg%� :mpI�"O5��ǼJZ,�֭,]bR�"OX�'�	?��L@0_H��V"O�9Ʀ�7�N��
��%.�ə�"O��X�l�1y�Bx�ŊŁ0���{"O20apM1H�بke�7<����"O�  �"T�Zj� O�!s"O���tO�X�r���� -��E"OMkv���6�15N
�l�0=��"O>�H2�E.?ɦ��1H�>{x���']ޱ��% �p9��V�2C���	�' By�rO����(sɟ�}Ī�R�'�4
���R?�����֒`b���'��������2���Pr&P1M�n���'���{'�\Hڝ� �JJnI��'�H0'�M�%֦���Ɣd�c�'�V5
��8P�c2�H��Ͳ
�'~���G�+?���K�d���Z���'�ȴꅄ���ݡ�h�� ��':��q�X�1;�}� m-_t;�'(`�V�)z⑌U)���'���L�PF�X T�U�Gj���'��R�+]4Yy|��scvf�[�'��:CC��#^`�R�ƍ[��8��'gn�q�(ٿr��K�F҂W��
�'S�(����6d��1[�H"d`�'���j�Z�����v��0(��'�*4��o
ryЇKO�K��a�'k$t0�'�>Ph$�LXv���'�X0��ti�� �˗e޽��'Jl���`��f
�}f���'�l�f�D�P �a���W<r/�5c�'J�}�A���b�T����(p_��c	�'�.Hk�
[�_h,�+��&c�L�'~��ӭ�4Pt麤�^^b���'W�zW�<`mR$z$%.S�Z�'��P��¾jX�	t)O?f��#�'��;�G$ p����X��'�vh*�$ƀ6�����ފ@� C�ɴ�v1:�#�Y�lA�k���
B�ɟ8��������=0��Կ%T�C�	7,xYB�%ڋ'�,p�o!GC��&~Ej��e#S�4u�4*L<W�BC��/�nYj��|��9K�"��
�C������&KȞg۰�1�%�7]|�B䉀Ю<0$��#�x�q�S�B�	�,H�J3e�3�J�i���H��C�ɩU�R��pmC,/l���רB��C��f���)� 3���+��U�w�C�I�+���F�(Δ����G�@B�	8c����������PG	�� �ZC�	e�0Ya��#@ƒA"Q��u�C�
e��%i"�ԃ'F\�Pb� S�DB��3m;��Bd|$QQ�c��G0B�,mENݩ��Q�R�=."�z1"OZG�ѐD�䔳
�1<�yp&"O"���ÕM�-���в`u�tz�"O,���đ	q@��	���1~���"Oz�B!�> W�!je`4����S"O�x�Ѯ��= �4�o�6X�Z1�2"O��ѱfF�R��h�7L��0�"O�ب"�X9�.-��Y�:����B"OZM�cB��&�ȇ��Z���f"O��p�Ӌ���3Ai�)V0t�1"O� �<�h�?c�dٺ��Ƀ	(.��"O�UH��W �Ƅ(e���m&�QCW"O4uQ�H�Gˆ܁���=�Z�"OAB�k*9�2H��Sꔱ#"OXTZ�E�&c���H蒷.�j`�"OH`1��z��L�'�G�%nܕ��"OfĹV�ú5���å�Z&�2�� "O�L���mW��6�� �h���"O��@� }9���!�.+��b"O�,�eoJ3u+�-A�AB�Y�a�"OxԨ���9T¸����l��"O��k�mѡi�0��ŏ!f�%��"ON�[v��\~mU�І�!�"O�I�B�4<dh���k(��)�"O�����N�=�^�+�LN���I�R"O���$+Pr�|�Q�GP���5"O�l8`��ƊBt�����"O�*��B�Zz0�	'HĢ"���"On�B��
�`���iS��.�,-�0"O�I�͎!@j�)��EƸ	TPá"OP�b�Ķoj�xR�\>&��Zf"O\�0A��e��]�F��#��t��"O&�@c�N%l��`p�-�7z8��V"O����zJ<���{~]��"O\  1��% ���3���q� x5"O|���EP:"���RĆ�*x�f��"O��P��B�M�D+�+	�yz�<��"OV���홨e��M���+�x���"O�� /e�^�*Á�vvR��"O q)'��6s4py��ߘDt�J�"O����Ɉ�8�ԘY��?v}����"O�ȴ��UP�K��ǺGrLH�"O�RN�.#�F��ƌξg�8�"Ohd��c��[0�k4�^9J� ��"O�4ȕG0m,]���&j�$�"O
Pg���� 7�>M��"O��pH�ivi���ф_I(X�"OlTs�+ɪ��)Jd�M��(�"O�	 0���}��c��-a*l!�"O��Y��#DtͩDDO�DVm��"O���A"
��Ѣ��8E��"O�c��`���+A%I�P�4"Ol|8��L�£��u�8��a"O��J�":`s��5�>�C5"O�E��%�-fF��pCAY{<q� "O��%���=YG��,��4��"Ob�s�F�b��4�N�Bt%�T"O:i×��"�,)Qubߺh�h�1"Ox�+W��50��\Q��5H�S�"OTݘ�Ǐ�	Z �Z�H��s� U"OXȠ�ƷF�$�J��"�<��"O�U�r��W�ځ�#,�#�<�z3"On#1��IBf]#���!1���Y6"Ol8��)��6*|9��\�T�&|��"O�ij7�G	�-�lJ6���XS"O�=�'��?�ȀJ��kr�l��"O�E����$iМkD� ([������ |O�`g̀�PEl�Z��V ���"Olp�CMG�c���*7���0����f"O���r�Ղlx�5	!��l!03"O�A9%�_�3��U���γ�ͫa"OL�ч$��>�z�S�'̓P��4*$"Or]x$�|vPd:F��3/8Y�"OB�`! �%e�UXӄ�+X�X�3"O� ����_O�1A�O�3�6	c"O�ѡ� ����C���:�"O���jS�*��!+�oD�y�n��"O��0ƅ��n�@��q�P/c��|�@"O�!c��o�F����ʡ`f�y��"O�%b��?| �iw��;���C"O�!p�ň&�8T(Cּl޲5�&"O�I�P[�f�~Ax�%�v�Fi"OVi߽sG2��5�Єi����v"O.�f	(n�]ѷ�%*�଩�"O�9��h�E��.Yj���R$*�y���*Ȃ9@�L� ���ɂ���yS�e���
7.�7D�H���y��5k�pv-Y�X�ܼY���,�y2	P�B�	V�Wu�|6AU�y��Z�dZ$�3���I��ϊ�y�'D�3�&�Z�CM�Ph��
2�y�*ǠL���3T�=4�LI�B_�y�T�1쒌)E �.9rΙ(و�y�
\**zH�i4N�/qh�p�f���y�΂GK�т��Ʉ�Y��y�c���\��_�zGй@���y� �^N0H#�(g�,�4m�"�yRjC�b�����2�:m9�@E��y�� �~�����~�0\�����y2�+ ����&I	�h���D�R:�yb���@� |9 �Ӭ^�����yhH` �ɺ[�&9B欋��yRЪ\C�КL"��5�W<�y�È�8ā�F虽I`�R�U�yR��@�,�¥�D�<8����y��1*��y�`eP�A`�@�5�y�L/YZ��b�@B�=�fH�Gh^��y�g�7BtB�
ؼ�"&�ܫ�y�+@"~���B�[~��8��ٗ�y�`@���`3��q`F����y�fI'{BR屗n��(���y�C�K���7e��� H2����y�B�S���2�#� wl՛A�ɹ�y�) �?5Ҥa�Mޘ<C�9�@@ �y2��(�^�ȑC��.��Xea��y�nB�G��#���t[t���y�Iťg���`�#	UV$`c��yb�K�oE���G��v�1�y�f��Z2���-�)��,i֦�(�y�+"h���ԝ-Z�S����y�"P��8h��,О�
Ub��9�y�R4K����,,(��/�y��#7"b8X*1��jT�ʋ�yRL����a��'їv-J���y�����P�GU�FXR�o֩�yR�� Cx �%�U��Q�����y�헐%�dlq@�P(��g�C3�y�'�
$L�� ��F���F$�y�Ď����S���o_T�RB���yb-��4Θ��`�&d߰�iP�@�y�[$"�Lu��OB\�\��M�y��u���!c��-C���M��y"�%0�������0��i�M�3�y���P\��0�%7�a�&��y���l\��f׊(��� ��ʝ�y�)�6�*dI@�L:%�M��T��yB�g�~p;%,M�"���h����y"H��h�-�mS� q��	qnְ�y
� ������~��Q#@��`z "O F�1L�����ϖP�
��1"O�Q`��ڬe�����X#��E��"O���p�DVS42d��h�l��B"O�ly�C�
x�0��e� �"O,�c�ETa�Tj����OaC2"O�DH1��1�Q�X�S��+�"O���KB�`İapMD;@K��""Ox�â�X�ޙ;r�U�>�P0t"O�}�0�n'\9� בj#�Y�"O��U�ELߐ�J��ɓ;���f"O6(�.]��9b��%P�4�"O<,�M�FX�Js(@/x8n��r"O�PV���Dc�d���87$0" "O"���E/] P���tq;�"O��y��<����ƅ�<#�%cb"O&87�Q4�X��e�@��2!"O�!�e�D���'E���j��"O6��e�Z� �2��F)P��9	�"O��ɣ� `�:���ݠ���P"OD��r�ձ�N�9��W*�(�9�"Oҕ���2��qH���%)���:�"O�Uad���"��$=v�R"O&�;�,Ʃy��̀�"o���q"Od�`2,EN�f��ϐ&pZ�Y��"O	f��˒��Mʕ<��d" "Oj��O�K󦁡um���t�*�"O�UQ4B� E~̌��Z�L�Pm��"OjY8e%��+��T2���V)*%"O���&���rVJa`��Ř8$��S�"O��C�R�aU	�h�
i8p�u"O�؃@���y�:C$CJ-�Q�c"O����r9.�$�-*�4�c"O�-��e�0�`�$�ˮ����"OL������c��9G$\'Y�p�A�"O�R�(O�-{h�0QHI#��0�a"O`��Dؓ1F��W�@u���U"O�}���R�~��M�(��p"O2E�[-vI<I���p,��"O�؁�g�"J�4(wlM7c< ��"Or$�W-W\&4X��
7Qb�8�"O¨��3��]��T�?D�+�"O�r��
x���]��\���"O��`���P�m��lY$|q2�"O��:�GY5��[ье ����"O\����|�z���T�h�\r�"O2��we�>G"���R��AI6P�w"O4,��
U�f��Z�Ș^<X�a"O*@J����,�� �ڸcB��I�"O(գ��6x�� ��|7TiRv"O���4���:��gT=O42-��"O���/^F�2��q��Q=0�Q"O��AʤlE<�I�E��3t �"O�䈥hR�X�J�(sfޒG��i�"O�h�Տ�<`��ۇ-(�d��"OtqXSL����ዑ�ֿ|%��`U"O��3�Q�6E���!H�,2,���"O�`���3  ��J�.p�Xb�"OM�`��pk���H�.T���a�"O�03��"[	�	qg�#r�Lr�"O�x��i۽Kz$I�,2ѺUC"O�8������m�#($�*�"O�D�p
��`^j� o� "m@a"O0���!D�Y���e�H��"O� T��6/�n�*{e���S���"O���@BW�d�.0Xd)�1Pf0��"Oj���`�;.d�S�燲p.�c�"O6e*B�6ea� �%f�0#ZD�"O"e�W����Yҡ�tJ���"O�����/1�X�E���
4Y��"O�LH��(s������?X���r"O��I�e�5���
D�H�=�"O(1��� /�n��F2JK����"O�Yӄg�-�B- �0?�T5"O~�;dd	j�b<���ڃ���J"O걪���<-"=�ց���9d"Ob�ؗ@�k�В B,+a�Њe"O�=	e�ս��btN�,�\���"Oֵ�Ł�*�TH��������"O��ɋ9�謰3��(?~|���"O8���e�%J��=�Į;8��`"O�U�B�	9�x�(�N�z���"O����원Q8=h� Q(��jP"O�=��$B�.��}(�9r���U"O~�Y�ޜ(7�[�M�8ek�APG"O�bW�I(�S�A�~W82C"O��"�5��8��<O!��ٴ"Oȥh���6l�T(k��фb`�"O��(�"��?�����q��IY"O>,�G,�)}��D�띄c��3�"O����H�?M[* "��+� �"O�{���u��噠	ݑڤA)e"O,����
N/���7. 7�$�k�"O셋b�Y�nH�����x�"O�0�B�3�auǄ�x��a�"O�Q(�S�hs��"?�Ja�"O��Fc��72���S����"6"O�4��²&5�u�P�=�p��"O������F�Z��׺
�<P0r"Oʀ9�FCw���X��B>a�(ɑV"O�,��+�C��G;%�2 `�"O�t� (ٌ�����Q�:<z�"O.|h���1F̠XAˑ����"O<|��e)'��$s�H٪�޽��"O�D3�B:����6!��� "O�!���˶G�4�3��)>�XKQ"O�q#rW�=�d�J�i�f/y� "Oh%Q#]�-� ��!.�[�"O�����/#��(��(�PX]P�"OۨCO��]�ӂ7Id����"Or�7nO�B��H �k^�f�!��ɮ*�Vx��mZl�{��Y�!�Zd�
�1Ǟerh���f}!��M�.n����&P�N�"��ޝ<�!��P�h4Q�*ԋ	�T`�C� ��!�bX� {a�r]>d��Ğ�!�D�|�cf� HV�C�-#d�!�Q�!v��"��-\���)�!�Sy_�:�'�BU�mjg�ǺL�!�ͩ,t�<�d�X-,õd�-�!�Dʿ���y��$��0­�s�!�V"�������(dw���V��.!�D�^�ب�`o
 \�5�ŊL�?�!�/O4hm�1��[���ELT�!�dC�����D
�`�x`B�*�!��7p�4J"@.I~< � iV�!�ĝ:n���OT( ��зH��!�D��I���r�)|aB���şW�!��  5��ӹDp�mB�&���lإ"O��	pH�-g���r��O��0"�"O�l+�׸���.���=�!�T,="qG��c:�ܲР�9'_!�$��Zۀ���!�,:~4���#\;!򤚶Y#�h*���0br���B(!��/ �h�k���7p` ��!D�W$!�D^;JX-��] 4����!�L�H�!�Խ3z%� bK"��c���!�T%MTV�Q��c��ԑ��h!�ƣt4�׎�l�b���a��!�dŏQ�b8#�
�8	�L��g���X�!�-7r�U�$Í2�PP4��,�!򤘁T@�5�t��B|���9�!���>
�ӱʓ��J ��F�2F�!�����peį���Q �U J!�F15�P���䙍D?05�BQ�~3!�X�Khl��I�+Dժ�G�'!�DΜZ�h1P'E��n �4KE�C�2�!�DR�a:x�SE9���R��=n�!�D�4MV�����^��3Q
��7�!�D�Fp���s�I�b���P2�!��ӿ�n����ԦI�RP�q&�DZ!���-�Qp�O�&����6���/C!�䟊K�V}�F�ٞU����v�ǴL)!�DB�b�c�eA�����F9!��Nޠ$�D�Q�B׬~[�9��"O�����S��17!Jz)�x��"O$�Ac/�0ZKF�0���^mZE�f"O�͉�јBDr����U����"O���B�?$���R8A��i�"O��Xs�[��-I��Y<�P�s"O�E�C�=HR`+b�9I�.�"�"O$���)O�+ǀ8�E^P��,`�"O�q!FI��S |���H"����"O�qe�<3bM�\�*�����"OFHS-�-7E8;㡘�θA��"O�p�`�l~�=�b���2�X�`�"O�(�q�n��1�.��g�l�"O�C���� :28혶j��R�"OT� �'�72�Q�@�o�rdv"O�	��ʞ��^%��#%�*qs�"O­ ��+ui杺�%@�JA)�"OD�Pc�/H�T�R'�&}*MѴ"O^ar��ُv��TbG�3Sf���"O�8����&K7<u+4%��DO2�c"Oz���Ƌ�Ā�.�JD�!�"On�9V�ڂm:b��C,P�"O<=J���9�6�'Z�%Zv"O����oP.Cy$li��S���Up@"Ox�i�	��  +�=b�"O�p�C�(T< �®� Hnb(��"O�q"���,Pޠ@C��&���"O~K�mU#/
��@��:SG�Lq�"O��ӑ/_�maz��eΥ :���"OvL�g�� ��݀L���C"O��H�Q��Y�"��X�ܒR"O�Zp�[�,A�)�g˼s�(!�s"O�0ⴅS!mW�PP���W�f�)%"O�1Ğ�k�"��'�<e���"O`���	��D�T � �Q7"O��"0�L�s[6L��ʛK�ޙ�e"Oȭ+@E�� ��so�p�f���"O�j� I�4F���H�
�:�ʗ"O� �g��.e��R�nM�B�<hʀ"O<T�%ERT��D�Æ�3 =��g"O Q���Ӓ#mҲc�/&�	�2"O��sNFRfN��@�_�)���"O�L��B�w�|z�B��'�壓�	����Q	*>���I\�#�����ń�^9�t'�4_�qO��DZ�y������	�>tN�ٔm<�tE��O��\#B�nD� E�{ A��dʻ;�8�9b��zRb���%)����'OS�0�S��Ok����͝�vҖ�Ez�L�'�?��gg�OU�vȍ�e&�%��m��_ ��Ӫ���$9�)������ª2"�5��K�\��p��$}r'7�#՛gg�v7�\~�F�a�c�4OPI�P�K����0<僧l�՟d���i*��W"E���ұ!�2R=jt��"@~!�&oG�/ B��J�}�aQY_�ʱ�}����M�&@� d@љ�'�9�pl���s�"��1��3	�Ċ2%T��P��k���(�k̗-;ɠ�7�É9��4��a��t��v��?1�/�V�'�?7�,:2��V�ȱ'K`1En���O��=��}�(�.������^'�@�@&Ό�(O2�lZ6�M�K>��'�u��!�L�FlE7^g�1Q&�!w�����YF�i�ay"O�=d�������3zI �� H$8�� aT�ol�);¤� ���)'%����7��h`l��i&
����۵s ��Q�&��9����:*��2�V?1��D۫K���p��lܖ�{c�W Oe����
6�.��I��M{��~�'q�tY��S��@��5�vg�hy��BF%D�Ъ�T�K��C�*L>G��T��-5v���~�V�O���˓2Kd�딄�57�T����I*N��t0���&�vY����?	��?)5È��?i��?9�eI�dGF�B2[�K��R�A�p�p���e��Т�#��شC��*��,Lqfb���r�S$I��YnB����2��0 ˠq�(�/1�:���@�'�%
���Ms6.��� ��0r�И@@��2g��O��D�O��ʧ$t�3l�.�>MpGB:,�eFy��|����"W����"D{��W�����	�M���i��I�fOU�4�?�O|²l
7�j���п38l�{!e}ܓ�?���Q�e<�8!4�*�E�eіd4�=����ᒅ+�Ѝ V�YT(�#=كjɇf�!�sI�F����,L�#��	S�4	A�A�+�9�B�bɑ�C�O %l�/�MS���	p�X��񈘿Y�8��8���Iry�T�"~�	<E�y�ć��Y��u��]�J2���Ӳ!l��] &D"#،[�n�e���Ѫ����S�۵�Mc��?�/�j�q�E�O���t����� �h(���d�a�b�^�x�ʔ�a�V�^l�LA�*9Q05cFٟ�ʧ�"]c�~UZ�MY��~Hӈq$L�2ߴcD~��Ї8�����ȰP�Y�W�s��ht_�p�m��k�,Ȑٲ4/h���k��']Bι<��y��M#��2'<@*��ީ)��W�I?����>a�EҀF}j��Z+���+QC?H>9�i�.7 ��ֺ�uB֜{!�x���d��b5KցZ�'Va{rήY   ��   �  [  �  �  �)  \5  �@  L  hW  �b  �m  �v  V}  +�  [�  ��  �  8�  {�  ��  1�  {�  ��  (�  q�  ��  [�  ��  C�  ��  ��  ��  A � �  O �$ J- R4 �: �@ �F  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1��2*Q��'/�ܱ�Dnٲ�0�rG-E�ws���ȓC5p�yaL�!	:Xy���J+K��X�ȓY�h����a�$��'AM�D�d �����f�6n�4�B�j�?���� H,�&��+�b@Q'n�%+Z�Ąȓ6}ܤ�2c��p��������\H���'ba~�a[�:$���Ӧ{�2����y���?Rچ�q%�F�	����?�'�`�)Sn���D$à�S�U[�'Cў�'��^p�A򐡋0+߲5.
�ASl��W��F��6SU�<�L�As�A�'y���OL�=�O��xI#,�(�C����k	�	��'tD;Ue�46�8�q'>jæm��'g�0�¡��kI��0p�ј-�|�+�'��pv�F�m;�y �RuK����'�,d��o��۰�B���sh�0J�O�6M'�S�O�B��t��U��f�����'��p�pL�<`�н�D̑",/�m��'j���7K�7nfpd�5�ƟZo��S	�'���A�/�,;Ϧ�0�V�SFxT	�'q����
:8��R�F0}h��[��HO�8���_>bW��:O���"O����
`�=Un�w�\�#"O$�e��"Z��S��u�4�s�"O4��G�|bI�c��.E���w"O���׫U;�X����,��[�"O¬	b�2x�~!�W p5�R"O�}i� �%z�R�03�� a!�$W,zb��Х�Z",���fI!�D*8v�x���%x������!�D�t��un��u�F��7��7�!�D�sp4�b���B�j���b�!���'7	fE����$���r'KI!�J��H���ӓI� ��$p"ONQ�	����B�Ŗ�j���� "O����KƢp몹���)y�>��"O�(%��z�`Z��S3�D-�""O�!b�-,l��1�^#"�(H"O���b&ܛ.�{ �KX��a"OyqsMZ	r�x&K�9I|�b�"O�x��[)*��z�I�R+�ԩ�"Op�W

�M4�X�T�#�q"O���֣̔T@-�S-[�;���"O�-hf��!"��*��=��"Ob@�&�� ����תJ<Y�T� "O�I��3�.՛0̆0Wڤ��'"O,� �nŦ2��\c��׃w,��T"OΠ�D�X*F>j�!���x!�(�"O"i����a#2����]�#t��"Ol sG�P%�LC����~�,��1"O� �i9���;"mލ؀ҏ3k2�`�*O�9{��5G��� ��D32ޠ)	�'&��S��?��X&�Q0�> (	�'V8�r��R�!�$ޚ)oh��'���N� �|@�C��0�12�'A4Z���rQ���G��5�����'�8�����<1�놦@\4 4��'�
�a��V�M�"��wn�f��A!�'�4�s���BaG ���L��'���KQ��x���п}��L��'*48"6�ř4$��j�xHe*�'hf1*'L�U�H��A�lA 5@
�'s0QR�,�1e)2�3��2!�
�'�,�X��_S�>�E1��I8�'I�̹0L�9|�V�{E&�"\����'"�d��[�n^����^�S��ţ�'܁�E#N -��h0��I	MJ�'t�������\ �a�	�GcT�2�'��mB��Y�N�i�Z�v.��'�25JCHA������ŉ�Z�~ �'4"��b�Q�3����r��D�&���'��臆ֆtaX�s �>;He��'t��b�Ņp���ʂ�Ł%� ��'n��E�V�n�	�)g&P�
�'^�� �O�o����AD�7
bf�3	�'���
��E(���K�J����`�'��C�K�!vDF��O�.ych�i�':D<�'38�8�@� ��-`�'!��"Ǫ߳殩��A�r�"�	�'�A�e#�3��,i����f�ꁱ�'H��Е*ڕY� {g+�]�H��
�'�vM)�敁4߆ȋ�ɋ�����'�h�I�T��I��7ts�T��'Al�*��	/x�؁��ш~�z�j��%��cu����I)t����.�b�<yҰ���%��@ɚ��:��B�I#@e�Z�D��YH���N���B�	WH@)��B����F�-RڐB�	�Z��aD딉?������5Q<C�ɕn�Ҝ)�j�	5�`�z@�A�JB��=3����P���!�#aRU\�C䉹x4�<�`g�%o�@�gH��M��C�|Ѿm�4p���A��	�z��C�	�oI���e�Ӣ���ٶD.,,C�ɰԵ�ӎZ8
/J`�� �N��B�	�Ѡ�0�?m<j���ӄ9�C�	0*�[fN�p*Xy2&荞z��C䉵c,����yCV%�!	�p��C�Ɏy�P�B!�ӸO�huh��H�_>C�ɘ�Υ�f$F���|�w+F�c
nC�	,f�:٢���1r���Ӭ�m�TC��	2t��!P�qO�51dݽF��B�I9	�̼s��A�^�������B��2`nTI��ǚ3��A�g�i�B�I���I{T�ր;H�)�ו\�B�	�m��9�����(��k����B��
|L=*6A_D��`��Qx��B�I7䶁k�o�+9*D��&�<:�^B�I�5M
Kp��$i�\B���&@��B�	���8��)v&���a.�FC��y¬I��˄"�Q�FB�'�`C�)r4�Ɂ5,�51x0����g��B�InZ�0cB/�8ao�kw����B��u��@�M �ϰ\���â5c�B�)� I� ���8"S`m[�"O��8S����E�'P�~��=�a"O�$�G��}݊p�v&T�_�z�;"O���v�אg}@8����=�4��f"O8�BG`Ѯ���+�>�6a��'m2�'���'��'�r�'��'c��N�<V�3����~h�'���'�'g2�'@�'���'���P���%\b$�����p��ԉc�'��'���'�'��'���'����@"�7�h�A j�6Ik��';r�'�"�'nB�'���'�2�'zP����ٖĚ��2ƘTc��'RB�'�2�'	r�'�b�'�B�'\��9' رlP.�p�B�=��9���'��'���'i��'F�'�B�'�����p��bro]*[�*}���'.R�'���'j��'��'��'A
5�dBE/\|x%CR"ʑ+�X�V�')R�'"��'�b�'"�'��'m�ʥI�F���Sd�W�P�8��U�'e��'��'r�'A�'���'k�h��c����6�ܠTV"t�c�'0��'�2�'AR�'�R�'\��'>�I�񯝘3h��"1�P�{d�Y�t�'�R�'��'`R�'^R�'n��'��1��� hT℮N�e����0�'���'���'d��'��'���'���/ˈ<H-0!)P?N���(��'���'�"�'��'��p�n�$�O�����X��>U�uA�fBa��WXyB�'�)�3?��i縬Q5����(v Q�Z4`v$N���d��m�?��<9��g0�a��N��E�����ˮX��{��?qgb_(�M��O��S��J?��r`7R6j�����\�l�"`7�՟h�'��>��U���3x�:�$�� f�Y�Nت�M���IO̓��OV7=�n@jJO��P˲�W�~9&y`��O&�dk��ק�Oδ�ڑ�i,��G�wxh�T���/�>���&E��f�\���*�=ͧ�?YsN
�S_BL1c��c�\m!�-��<1-O��O�m��u�b�|�EaϺJ[�h��Ĵf�
��x�?3Q����Ɵ�̓����8~���
wj�p7�P`C��K���џx 5bF"Q��b>y%�'������!�d=J�ˍpEh��� ��5��'��ş"~�V��QƁI�:�Z( ���  &9�L&�V�ڝ���Ʀe�?ͧt��ز!��9o\<�0bśP����?����?��,���M��O��S���c��P�Θڣ����AW���B��O��|���?���?��J�����A�e"��+1�l����-O0al�45�|Y�I�|�	�?9��ty��<8�J̈խ@�vO�0���v*6ꓞ?y��Of�'	��1��?��ɷLҡl�|u�կmԐU��Y�H�◽7%�u��}y�J�<QXx(���_Gd�U�ۀ9��'�r�'��Oq�	�M��)��?!B���	"2�� .D|\2�c��?�P�i��'F�A�>���?ͻI"VњVI�(jfV�Z�.T�+ф��4 ]#�MK�O�D��Ј��ę��w��]�!�<nhHT����3��tɝ'R�'���'�R�'=񟦴�CQ����5[P�`@ڪ�?���?��i�`�R�O���t�r�O�pb�gP�BJ��Qro�$q��{q�d�O��o��x޴��'-z.��0g҄)
��d�bbj��S;�?���)���<y��?A��?!�A+T*f��'E[�s����1����?���dM¦5�����������O�ډ��߫	��z(W#ի�O(�'�b�'iɧ�I�<X�$4 s�:r8�u�eK+.�f̃�*�ZɌ6M�dy�O.�����;�PؐDG`�:984͔*g��8���?A���?��Ş��妩qԂY�B��[T��FXD����8pq�]�'{7%����D�O�Xƣ��p'z=i�`�<P���O�����7�"?Y0-։TN�i9��*��U�LP���"%s&�hĦ��y�]����ԟ������	ӟ�Oj�X�"HiLY���7���@�a�^�S3M�O<�$�O��>��ئ�]�Z�3��O~�dp#"�1�Ƥ��Y�S�'h��x�޴�y�!��"ClQG�~| �����y"�@uH���I ��'N�I�� �I/ ��	��\+�����Q4t��9��۟�	ݟ��'=v6MI�G��D�O
�d��=L�i��)Q� q�n��"�.�k�O����OΒO:�@1ٟat����Ft%�����������~�o\�'B�.�	ǟh�� J�k��aJ�$�z�� �'����I����I�0F���'�5���V�-�T#�#��aZ��'77Jmaf�֛��4���uL�=hd9PDȅsX,I��3Ot���O��č�'�7�)?!r�A����1�p��#��J�����-μqϚ��H>�*O���O��$�O`���OP8�ub�=c���ڒ{4^,�#��<���i�l���'yb�'l�O{R�O���d�%5{����qo� ����?����S�'E�d���O5Z��$�FI8N�L
"�ļ��|�/O<ѻ2)
��?��6���<�vo���ɸ�!�!��A�֊�#�?a���?���?�'��ā��2̑��@�S�D�b��*��,��ؘ�ʊ֟�޴�䓨?AU\�8���L�I��~��!)��Z�\��3l�:~j��.��M�'Fꐨ�E�?aʤ����� F��g�ߞjnNxR��T�O��L��:O����O`�$�Ol���Od�?��T��+Mv�H��@M���� ؟��Iȟ���4o�+Or�o�[�ɕc������r��U��mn|%��	��0$���l^~b嘳}^�ᄨ5�&�ٶ��3�@MQ!�؟(Q#�|2P����H�	˟H E���&T@��\38�h��V�����PyR�v���1��O����O`ʧ�����l�;+�H=sR�!r�P�'B�듑?�����S�� ؂})����^��}�b�ԂH�-�wAC/K�F�<ͧr��k�t�~��a �,ʵ�2'��{��'�B�'b���OM�I��M�Qg˅<Ch�[ƃT$4����L�6^�X���?���ig�O�8�'�R��L����+ �E����K����'(�H�ix�i���j��?-�W_�`C��ՆѲP׍��J�t��v�l�x�'{b�'���'��'v哗��d(��TV��T�OԾ4�ش�q��?����O%j6=�a�tA�<�v]��@��`S�PH�$�O$�d6��ɇ*0�6�x���ť�I҈�cb��5Zy�����}�ȑd�Ⱥ&�2'HN�{y�OR�X�L�"-����3{�n�+������'3b�'5�ɯ�M�%�ѽ�?����?`�)�^=�H ����C���'�t��?����3�b�dFԅ����͆A"l|�'& �R�DT�'�D��dT��ب`�'Zp��$V�R޺ �M�������'^��'���'E�>u�IA0� ��됉H��,wF���	��M3�$Q��?���4���4�^�0�� �J��'+Q&`��Ѻ�4O����O��U�W	f7-+?Q�	� m�������VgZ�i �3'�&+;��$��'+��'���'���'���2�	�W\ �t[5��8��^��شC�J�)��?�����<)������)-,��Q���h�	����{�)�0T�$���Ц8V8�Yţ�	f��(%��:����	� ��O�9�L>�(Oݘ��Q�C�A�2��:��S �?���?q��?�'������F ៜ��N,��UJ����L9���c����4��'m���?q���?��dS�dRPP
��ؚ6rP��nH
�t<��4��$ʻ	a8��'��O���.w����@V�-��jT�݃�y��'^��'F��'�����A>�$Vڄ#Of�3Iΰs�����O��dM��i`��TyyB�b���O�,��+	=2���ڤ�7�\����*���O��4�Խ�IӀ�(�F���j�)(w
@�6��t�4���hڕu���������4�@���OB��� &�a�&�?�x��CK�]F`�D�O�˓���*И���'B2U>ys4���y8~\�&E8kxmU�&?�]����_�S�T���mt��62\`U ��X;�,���h]�`w�xsGQ���t���]W�}��x�#�"!ʽ���+u#�|��ޟ���ӟ��)�SDy#x��	��G?5��]�A�A��<�Ԍ�?t��O*�oR�� ��	���9PD S�4��!�,r|��f�����O�LdoM~"�2$<T�����6����烋;��hC�ܒ[��<��?����?)���?�-�(�	 #�2\�����"DV�qX��X֦�@�m@������@&?�����M�;Bn4�p��S~ ����#�2] ���?)M>�|�c�
�M�'a4m�n}��q� �P��aX�'����F�\?iO>I+O����OL5�T'\>�h<@$�I(= �j*�O��d�O��$�<it�iCp��v�'W��'�*tţ�(ӠԲ��W0_ڠq��d�Z}��'3�On�0$A�C�ђR���qb}�Ò� �E��=H�v��� 8"ǔ�d �'+/��C���A��b��ʟh���������|E���'����cڂ&����\�	Ӕ�'j�7��5uBH���O��m�X�Ӽ�6���YBn��GF�,|����m��<���?��3���4�����Cč��~�C���Y��=��H��4����݊�䓶��O�d�O��D�O6�d�>l�A����/0��ꃋ|&l˓V���U�'�����'��<j"-������οw��`䩯>9��?�M>�|J֧�c�P���UJ�DC�I��+ ��'��D�&p���)���Oʓ�`��!�Y�z�`�m�"]��4���?q���?1��|�(O|�o��WM��I@d|9��Fr��i��-�����5�Mc�2,�>	���?�;Zup9�|�� ���"h}���X��6m.?1�CL<Pw~�I]���ڿ��bV���02���)9t�r�Ӳ�y"�'6��'�"�''2�IӗA���f_>J���qBȝ�>˓�?�A�i�j��OF���b�O���d$��@(�u�1�ɯ=��E:���O�4�ʱ�0������L��͈�c��X �e��,\H�P�� �t�0��OΓOt��?���?��"~��4�,[.��Юdj�e����?-O6Am.S\p|�'�\>��AȞb5萤���8,�h��??qQY����H�S��c��r�\���,�;��m��Γ/v=Ʊ(�c�=W��U��[�擌���}�I$��q�j�6�yz��]�=��	ϟp�'5���\�#޴8u��3��M6��A�_�(�	����?��Hw�v��\}�'FFA(�m�C|РOU�jh<)c�'�rĀ!rٛ���L�@�М4,�t�~� bQ�P:no~M)����b����5O��?���?Y��?a����=����`�<;m6�+�델N\^$m�I���I矌��^���)�����JU��v�HW�:�B�r�Oň�?y����S�'l�Ta"ٴ�y��/fpaPlR�-���d�&��	r,���'�]'�(�����'�"m3 nƂJ���KG95��,�B�'���'��X��KشiEк���?��`u6�aJG8/I���c�� n�0a�R%�>���?�J>IG��)��5E�C!,�C&Cl~�k�$^
p��4�i;B��4��'��@W1Y+�}��ŝ0Q��V�q�d��Iڟ��������R�O
�E\3i0e+J��R$LT��$;RbDt�p�rB
�<YR�iJ�O�nM-~HPd@�Z�	���b@�S��O��d�O�u�R�hӄ�Ӻ�Bѓ�����0u&��;Vb� F�p9!�0~��O�ʓ�?!���?)���?���i.M��8e�<�xToә^�P�+O2�nڂ!�����؟$��p��؟| tk7���ѱ�I�f���H��ӂ��$�O��b>���)%��	�u��>9A������^)R�k�ryRSpiJ��	�!��'j�ɫ;Ӫ} �˸+�||`�o�-�f���ӟ�����i>!�'Yl7��_2Z�$�)D��bհ�L%��&��$要�?�wZ��Iݟ4��7�حb�(Gw.t�-�H3�B��Y���'L �q���?�}Z��7�
<����e7H\�T�_�d��Γ�?1��?����?����O�9RG��?u׆�����7`��'���'��6��=����O�mZs�	�&%,�*��V�1�������=H�H�'�t����S=u6�	o^~��IK=�`�A9w�]�gF��J�D -��������O��$�Ot��!H��xم�L[Ĩ�Q�I�+sv�$�OTʓ0b�6��s]��'YRS>i�b�%&et��c�K6�N�{�&,?��W�8���X&��=AA8�E_oӂ��GP1x����u���p7m���4��s�� z�OtY��H݇[�H	;Rl�:q��ݰ���Of��O<���O1��ʓtl��.	��li���Y!�`,�0m��3��'9�Cmӄ㟨h�O���� G��3��� .�z�4%Q˓
:F�0ٴ��dM=hl41�'uHʓ��u���1D���E+q+��<�-O���O�D�O:�$�O`�'!��5���yȀ�j3ccZ�иi��E�T�'���'F��y"�l��.�?"v4`1iZ;t��hҖ��&5��d�O��O1�\[��a�~�I�Sb`B��ق6�N�X�銍�f�I!T��mx�'���%�|�'~�'�Z�[���H4�B@��(���#�'���'�Z��3�4n�,%���?��)�ͳQM�K\�D�㘔w�����/�>����?�N>����
� "1�K,�9$�Aw~bbց>5~��KB�+��O"z��Ƀ+�b���EnD����:?R�P��^�!b�'�r�'B��П�xb���$�^]@�,���]:�Iϟ��۴w�$��)OJ mZn�Ӽ�A)	)$�t�eG[�L�rT����<����?��R�pi�4��䓩4Ո����a$���&Y�4�ȃGV��]�pB?�Ģ<�'�?��?i���?�co�2d�X�g`�Cv��a�*��Ϧ����ԟ��Iڟ�'?��ɔi� �Z$��%�"� R�LY��O �$�O �O1�(��%#.I�~���ȟ�c�$�D�\�n�
��D�<i�$�y��D�����Œ,����ڞyD�@E��8� ���O���Od�4��˓g�f˔�v*��םkj�ii��&Б1M�>u�R�~�~㟄��O��d�<i�G�y)�T	^z>pB*��|m�!޴��d���9�'aP�����#���KD�p�S�/��|��d�O���Or���Of�D-���WN���dI���#ư;����� �	+�M�� ��|����V�|�#D�)���rt����ą�&Jݣ;�'�"���$�:d`�6���ݿ)�V�@�12"�ٓA&�[��r7.��8#��|"^���	П�����a"E�e�3p ��.��hq�G�̟��hy��~���!��OF�D�O�ʧg�u��M�Pk���r-�>7HT�'��ꓞ?y���S��gA	T��t35K�~��	%��
M}�AE��.ɛfG�<�'k�~��d�	�S�p�k�x���x�$&&��Iğ ��џT�)��Byrie������M>��⥌����;T��]X�ʓ;�F��O}��'��bS#B�z�H��^D����'=��_1�&�����cC9q�(u�WCJ;IiZ�8�H�[lB0�p6O�ʓ�?�7g&�?����?A��?�'6�����%�U�����ͅG����i�@�
��'"�'i���O���'�:7=�H�ˁϒ�	�\�Y�e��sC��C��O,��$�4�~���O~D˔�l�\�I�p��%f��U�Q�h��,z�'�@Y���䟬���|�X���џ�30��j�r�a���B��sO������ٟ���my��}�F�J��Ol���O]�����s�(��&�G�a���0�1�	&����O���&��.Ѫ�ɤ�����;���2R�	0u*���ɦ9�|�D$����	�,�6�B��ȇ�pA»W\�4����8��ԟ���B�O^���r�i�`�F��4�s�I*^��e`� ��h�O��d��}�?ͻ!}����jE�`�����-e�n���?	��?�F���M��O뎄-o�`���O�? rhb�JL�L**t�@��I��ub�.�$�O��$�OR���O����Ot��eP���v�̂4N�x��'hw�ʓ1��/+ �Ƽ@T�'J�O��������]M��p3�S
��P�Nb�	�X�Ily�S>m�I⟤86	�p> � t$"]z�;uI(*��<GC!?yw�8[Ub�ć�����D@ E2l�`oV?H�}x��M?KB���OH�D�O��4�tʓD%�	I�ROS5��ٚ���$�ɢU���2�~�d�ܛ�O����<Qń�}{`�2����L`BA� �(+޴��$@9����\��^���$<M���eO�7��A��H_���O��$�O�D�O.��5�ӏ�uxiS�8�x�I�E
j$��	ǟ��I��M�BȄ��ݦ�$���@Ѩ0��D��U�#]F�0'�{�I�d�i>��F�릝�'�&�P�J�+�2�Fo�=|��E�A�4�f��ɼh��'��i>��	՟���	KB\b��ي �v!b��7I���i�M++ONTmZ�ks@4��ٟ�	^�$R�N�؝31n]:K=��o��y��'����?����S�$#ї ������uQ��V��4B3}mӑ4�&�<�'b���	T��d��1+3Ꙡk_ĉhd!�EK����柄��՟��)�@yBD~�Z@cv&�
 �*aZčC��Ĭ��$WfH���O(oZZ���I�P����)f����r.X0�Pe �ş��	�U��n�H~B���n�����$�)V1�9�3���-�z�(��C���<����?1��?����?Y/��ģ$�G^/�%�B��c����h���y�������џ�%?�	�M�;d��S��2?.���(�;SF�A��?�K>�|b���M��'�@�ڵE]'M�FVN�(�T��n�hQ7K�:s��"��<�'�?�$�9�̠��:y"��c����?i��?Y����K�I�w$�syR�'  ;��Z�T{4[V���s|TYJR�Mk}��'��O���'Έ)�a����R�R ����tBW�KD�5:� Id��JA� 	�����A�5 ����F�x��]�·�L�Iџ������G���'�U@�%J�=� ��G�?ydF�"��'�6��^�˓ћ��4��Hcզ΁Yu���N[�D�6�h2O����O�����f)N6�<?�-�G8���T����J%6��Y�b@2fY�JH>I-O�)�Ol���O,���O:V�ĢO�Ԙ�%�W��R��<���i��u���'���'l�O�2"�B���0!��9�,�57L��?Q��� ��W,*dxUnu��x�="(�������. 
��� �'J�'���'_�Ի��Sq4���	�5y��:��'���'�����^���ݴ8���Lg����cR�{���U�����R8�&�$�O}"�'
�'nthX��E�:�
(G'�l��p��M����xr��V��4�I��R�BTG�|���w���0�½�;Of���OT���O~���O��?�gLȬp9�5�`8�|5�2��ʟ��	��Qڴvp>u�O,6m)��H�mdX�[����X�@ ��K�6���O@�D�O�)�.��7m*?��@d�=2t/�	b�IP���\��̨�X��?� F6���<����?����?����.PJ�	[��W*>,ZЌF��?y��������FW����	ܟ�O2yBRo]	ġ#�a�$'�,c�O��'�"�'�ɧ�)�3_�ܸ��I��x5��m!L����e�PDy����S %�RBEo�ɺ%�h�K��%K2Hp�%M�	x��(�����������)��y�+n��z�`Ĩ�$������Ԇm���J� �<	��i��O���'�h54��Ը4��J��̈��2<���'8����i;�ɺ>.q�4��H��b1�E�=<}lA�Ń$��<���?���?y���?	(������E13�Y@6Ƌ�Z9��%�æy�aCty�'���mz���TAؑD�����M$E�& �W��ޟ�I}�)�S�B((n��<��eT��B���=0��M�dI�<�AX!qZ@�$ݤ����4��ر
�������#��{0�8,����O���O�ʓ��N��^�	��$��aD1t�n��	P)X�@QU,�B�`��I���Ik�I�R6.y���7��N���=n�%I��$<2�|",�O
��}�9��,�
���ݜ_�л���?����?Q��h�d��Z8q8h8G��.x����T-���MϦ	���Ny�|���杲K�-St�Wx�:hs�(��pԌ��ҟ��'2�	)c�iV��6'����ON����R�l�x;cd^�W��I�[�^y��'�"�'cB�'wbR�5�eRtϜ0n<t$��O&o�	)�M�G���?a���?�O~�a��$s�B���H3���j0
���\����ٟD'�b>E ��V,�����b̌&˔�jP�1v��RK)?�ՠ�h������F6�x�Ж's�p�3�A��%�'k�'�B���DR�Գ�4�������Re�ac���ENR=���)W�F��T}�'���'�3$i�$V$k���Bo�xqW�	�tܛ曟�����D�������I3v�E�X�q���T8TjJ S3OZ�D�O����O���O�?�E�o<�� ��B�CI
��X�Iɟ���4LpM!,Ox�mO�d�������7	8T-"�̗	�JA'����ϟ擔;��AnH~Zw��� �,��"�PO807ʖ''��T���M"�?Q��:���<����?Y���?�W�=s���Z�O�I!�L+����?�����ĎѦ��C���0��矘�O�l4�T�M�(���T�_CF
�O�M�'#"�'�ɧ��U�S�p��PIH�c��
��^e8��\3�$6�cy�O��1����ah�3c�]:s52�,D14y���?���?q�Ş���Ԧi���)$����f'�jMD�2���5�"��'=�7�(�I
����O`����*T�4AǆtA���
�O���Y�! �6m9?i�
���>�ہ䊾8ZL��#�	�|D�4
a��'���'��'R�'���&^$��7� V�"8�t��(�@L��4)�~����?y����<����yg�.Z�58U)�*sv��������'�ɧ�O_dH��i��D��E3`��w P�!n�j�ָ|�DF�V&2��3h�O*��|���ebl�kW�H�P�*�ڴnV�V�����?���?�/O�l�#l�vE����L��+88��yҍJaB*�@f�ʥ8�t��?dW���Iԟ�$�4 �?B�����O�{�l�X�%9?�� �^����۴��O�����?1�J��dzΩ���|�x`�H��?q���?Y��?	��	�O�KQ��">�ຶ"�#8H�����O��n��"�T(���T��4���yW��0-J 0B��?�`�!	��y��'�r�'�NtQ�i���-ldtJ��OI��9�@ԜJH (��l^��BN�^�	�i>��I̟�������8>Tqa��@�]���#U��;1�<U�	�Y�����j��<�������8�M���<��SC���3�-�(�����! �lq���P��?A��?"ɨ�r.�����O�ܛ��Ha���!K/j�,gR��$�@�B�<��D�@�l�D؊����dݢ{y��Sc��1��:	�����O��$�O��4���uv��D�����G�6B)Z������I��;�I���D�O��$�Ov�0�P9t�:1��iȋn�
s#�,!O�7-/?!`��Z-
�|���`1b$�f�.v��H`�� .A�Γ�?����?q��?����On*ٸ@���4��)}Eb�H'H�<��r����X���$�'��7�=�$�|� � !�l�Qi5�\P��O����O�)���6�<?���Y.KB�Tـ�O�2\yIf�ވn&��4d�O�"K>�,O���O&���O$9����@����j���O��d�<17�i��Y��'��'���3
�ҋ�c3fP���@ Q����IП@�Iq�)jd�K�rx�d8�kI����;&˕�G�4�VO��?���*O�iٽ�?Y�!�D�o̅�� �;6*����9�j�d�O<���OB��i�<I�i(��҆�c~ޅ÷�4��Q�D��(i��M��b�>����3�MY�${�Y�@���R��?�E�M�O�R�.y��	���X�F�`!���G�f��4+U�J��d�<q���?���?���?Q/��Pq��_H^h��o1c���@��ۦ(#.I˟��I�P%?�I4�Mϻ"N��C��e>��3��<&��9(���?yN>�|f�.�M#�'(d:AgL�Tm���+�h6h�#�'v�dJ���П��v�|�W��͟|�!�A:_$|)�^� 7���S�D�	ܟ���Ty"�i��-@��O����O�H��8Q��Pڕ-'l� ��gM1�	�����O*��8�Dݪ:�ZQQu*B2\���f�"��Ʉd�Y
�� $O�b>G�'E�����j�ҥ��U�s�LU�%�8z)�M�I�P�IПt��n�O�e z�@�[���򑯆�B����G�6_+]=�I�Mk��wH�$m��Ks��W�\�z��\��'�2�'��n�~�֑��"��^�'��I��!F.��x�2�)����F�O0��|���?)���?���^�������8O��՛'���Ʊ�/O�Qoڤ~ ����l�	f�'�ƽ��l��SŎ���?��p�p\���$�b>���E��q��0��Fϒc7�ea$�� {3H\mZ3��#9�(ܻ�'M�'剬4b���NJ�>�d�x���5w<|�I�������(�0l�|�'Q*6��/l����y��t�A�D�h�M]/����Ǧ�$��ɓ��D�O��o�^�`RA�n��	hw#ٷ&!����M�'��'��t���ӓ%��I�?q��3I�b��BHz�NZ?���П���������I^�'L�ޥ ���@�-I/'d���?��G��R�@����M3L>���Ít!ڭ����
�:� Č^̓�?�,O���Hp� �KT���
�:��D%�4<A��Sj�b�S����$�O8�$�O��V>w�0G`I:d� %D��x�����O>ʓ���a;���'��W>�Jb�Y�B��9/æ_�t`A�E.?�X�`�	���$��2�p�j���l���iF)�
O� ! ���C*��ݴ}��i>A��O��O�qi%���j@(	�	ן5%�h#��O�$�O��d�O1�˓Wf�v`
8;�����(=Zjyx�b�#�z�P��ݴ��'Vj듣?�"G "�\:��ŗ�j �t,ҋ�?�J����4��D�??��%A����S�x��YR�PEDM*1hR+�4�Iey"�'U"�'���'�bP>����5;<��J�g��u�F,��d�M����?����?K~ΓO���w¤�(ݡ=!�&��he#"�'�R�|��'�.˛�<O� ��#ƂY�O� ��B����2O�9�O��?qA9��<ͧ�?Q4k�,�� ���H���sĄ�?����?�����H�u����Vq�f�d�,%�X򐮊�5���g/� t��O���O�O,� G�\�
q�]K3��l�N~r��:Vf���6.Y�ؘOp���ɀX"����<H0!��K�0��FGB�'.��'���Пxxtk<���QIx%��[ş,a�4Rn&<*���?Q��iC�O�������b�U�sj|�x(�m��D�Oʓ@=�y�4��䇏�����'��8(��95�fXA�Os򰸒�'���<����?���?���?I�F\�$�a��,��g`6<�3/ٓ��d������ߟ�IџD'?�I8d�`չ�K�"59��3�Y=b�p�{�O����O��O1����H:8>	�S���kC���Gj#Z".�c ��dQ#�T�F�b@�g�	Uy�߹AT�	�% '&I$N?BB�'B�'��Or�ɕ�MKN��?aV���}	�B�	<L呀��?)�i��Ob`�'�"�'��hV�0L�I��K��^�3`�\��i���*{��l��ԟ쓟�Θ�B#x,1�H��1�DK�d]P��O����O��D�O���6�ӏs"�(�
\*3N���Q
��`���˟��I(�M�$�^�|b��^a���|Ҩ�� I�O�o�<0�&���'������\�L��V��0�D�KŤVA�1���!�=biP2�Rp?�K>1*O����O��$�O�L�C!2;<0ơ;<���j���O����<Q��i�^���'O��'z�Ӭ�,�i0.��T�0H2CԤ���I��������Z�)��dR�F�l�ڛ&踄B�$�.1LNur%�O�����J��@+ǔ|�旣+����|m����'�F�J��?���?��Ş���Gᦗ\�حP�I3.�y�L�4�8ж)�O���ަ��?��W���+'���Z��'�T,@��.!�ּ������ئ�'�V @���i�/O4��#E�*)��p�A�=��I��0O˓�?Y��?!��?�����	�:�\<+���vc�)�fbӧM�f�m��j#v��	��@�Iy�S��<�����!�Y�~��)Qb	ϫO{��[�Θ)�?����Şz+l9�4�y�$�"	眼PjКQ~$�� ]��yb�I U�������?�J�e�y�
�?E�@8�	%O~%oZ(u�R�'��$̹y@`��vg�,W+2�2�,F�O���'�r�')�'����v�*hD*��g�J<n�]!�O�T��݁a�a�� 6�I_�?�� �O����&j�M/>��!��ا�y��|�.�#�� ��}��+Y�w��u��ء��O|���Ӧ	�?ͻ��!��ɉ0��5Q(C�rb��?	��?�oS��M��OB�R%^����-�9�r�RlF�C�L4�V�
k��'��Id�'�&$J�b�[d(���e���On�lZ<_2���	�����Y��&�����J=E��l�S��41ҵxR�(�I̟�%�b>�jT&;\E�Y�&AZ�Bߤ�V�{�"n���D��rؓ�'��'=�I�x/"�J��,��0�ᥓ*F�����S��):��^ڟܛf�Y"A�	����#\0�a'�}��4��'�꓇?q���?�bѲ{������1B����� -��4��ܻ[ \�`�'>�&��v�n+<�[W�I��0�VS���,�O�4AC��t�"$^V�F`HE��O^�d�OB]lڰ,˪�I��&�|��P�Jn(9��W��QQi��iy�'�R�����5�&���9ԭ�d�rHX��V{ZX�5AV�cV��I��Op�O�ʓ�?A���?A��5r��s@ P!]��a dE�/$�:��?�/O�lڱ��U�	�� ��T�����2� �PF#^I�� ����yB�'�n꓄?Y���S��n��lc8xe�'���mR�6���FG7 ���<�'2{��ID�ɛKq��I��OY�P)����&���	ɟ��IƟ�)�SUy£u�e��Ӿ7F�H@f�O�J%v��`���I4�d�O��m�L�	ܟȩ�OH�ğ�,E"�B$֊���oXf�����ğ�B�X���u��H�6�$�^Ny���J	:h�jj_vU��Խ�y�P�x����	ʟ���ߟ�O����h�$})�T��h��{��f�ڈ����O����O���������]	����#�.
R-�w��	7���	Ο�&�b>}� BTզΓM�FL3b��53pr4
�v�̴͓#f�@�#㡟�&���'�R�'��a!���L�
���Ǒ%{��h��'AR�'c�Z�H�ٴ:�<�3���?���S;�1����s��Ս�>8�XM>���9�	Ɵ��n�I�	v���/F<5��Pa���<fV�xjp�	2�I��Mџ�T�ٍ.�|�"l�g�r Vcv���m�3p�H�ࢅ�73e��dͯU�����E�?:rH��Sw^���h�(<��gΦY�:uD�+v9��L�x/��bߓd� 5����/2P�=Z�JH!7BR@���&�zQ��L�*�ܤ�b��4�R�*�l��mBIO/#j�����,S��1kEI���aDѕX�&��&I+WE��p��'jL�)��ı>Q�D�g�-+��b�G֛L�vlKS$�2{
d2�E�<,�e��	"(hd�S)��(Mf��V��M;�� �v�&U���'��|Zc��;�&�倽y���6F%��J�O�14	-�d�O����O�˓-t� .UK@�|��!���:�8-�s$�`��Iy��'��'t��'!:�sw�I�D^�YX���t��̘�DK3�'���'|�U��	�A����͜��2����Jc��x�%�M�.O��� �d�O��D�� Hb�InF��{p
������Ɛ-���?���?a)O~��'�@|���'G�-#�d\4	y����Y1���0��yӘ�D+���O���و��p��RC�y��b�4@ӂ8�2�w��D�OTʓd��Q?�������`�J�N��ԣ�Q��E�J<���?��"��?AH>��O1]sw���PB ���K=��K�4���.6HPnZ��H�Iٟ��������u�c�H�6(H��j*p�F��³i}��'��0�5��/�	9�~�ÕH$_�Ta�shΛ��7�
�d���mZ���	�<��'��İ<q��d��p�EȔ�� �eL܏N��`��O��?��I�d}b�� ��1�@�� �;�`��4�?���?���H���qy��'���%���p6h��Q���0UIÉ"��O�F(�d�Ov���O����`�^Ji���F01�1�/����I�0~���O���?�N>��[P|��'J�Gj0�x��rPv��'�Ҝh�'��ß��I��'�hp�T)��m"WGǷM->4�M�N]����$�O��OX��O
Q!5/��(��ʥ)̓��%��\���O����O(�$�<٣˃�F���q�HDTD�0M(	u`]�H�v^����`�����I�B@��8��-��.K9a�%����	ž��'i�'��]������I�O�-2�(ʇ0E�<�����`�f�Y�A��W���D�	-%�r��=��I��u(�I�W�	;nF��s����	��0�'�&��$��~B��?a�'].�t��K�<<Y:1��L\�#Ŗx��'�2�A�1�ON��
0ʨӲ/�B	:����-�6-�<	�ذ\�6�'5��'����>�1pY� ���Y�b�I��On�dm�ڟT��f$��?����F��;n 4�W�&.��HSj�
�M���F�4�F�'��'��h>�4�����?.�Z�:WaޓF"�鄃Rܦ��I��`�	d�)��?i���?��Hc&��"���6�)i�V�'hr�'O��9L-�4��d��@j�JA�.6q�4  �TH�ȩpb���%�$�~��'�'8�J�1E�0�*�"ϭ9��)�@� iK7��OfEs_����4�'ɧuWl� ����7:{T�a��I����?�*O���O��d�<�f�J�1��0A�?/=�-���̷EE`�'�xB�'���|RS��"Y��3b�7a�|��Y�CHX6��Ov˓�?I���?�-Oҁ�a��|�m��X�q��c�V,�j���~}B�';R�|R\�����x�EL��2r|s"��V���1�H�����O��d�O�ʓC����������v�$���7(�q��'*��7��O�OF��|2����Y�r��Gf��&�\���oF�>�6-�OD��?Ae�,����O���k�֙E�
��GCҽro�eb�'�T��E�(�Ӻ�g$��4(uj�:�Ȥ�D�x}��'���XV�'�2�'s2�O4�i�Պu����ݐ"!ǟOI������$�<��H�p��ħOt`q4E�:�ƙp���;��o��ͤ��I꟔�I�����Xyʟv`yp�Iް�Ƅ��2�M}i��O1���D��Y������A� �0Rql�mZ�����B��7���|*���~Bφ$98��b���}��x:���M����?v�s���������$94N%����\� "R3.��\۴�?�4�U�?����'|ɧu�dѝ��x2S�S�
�v�"���ē�?�L>q����$�O�!��\�.�$ Q ͷ/��� ��SX���?I���'hr�OP��V��\�
��C�Z�x��������O��$�Oh˓S��ɀ8�B�xSH�(b���A,�q�vX���ߟ$$������'D
�#��0H^�딍��mY��(�L�>Q���?Q����dڡW�b|&>����J�v��h���ٵ",�ZReͩ�M�������4����2�D��,٠�Ӕ����� ��Z��M����$�O�غg�|����?���3b���\�L)��f7%���Q�is�����'�zi����Ep�k��QtТ��ЗA_��d�i��;*ܼ(�ڴe���͟������_k4��)�l-�|a��c���v]�d����M|�J~nZ�O8�D�Q	�r����LB�7M;d2`,o�֟��	П��6���|�A$H�7���ۦ*��:*�5�� Λ��'���'�ɧ�9OF��k�Ҕ���4��l�g�_
l��ɰܴ�?���?��O�<e���ty��'��$A�v<�2���K��m��똆U`�F�'$2�'1�1������O�$�OXء&�ܵ*�d�B�,�7{�"!R̎ڦ���8F֒%�O�ʓ�?�*O�����'%F�&����: 8�y��U�����v���ԟ(�	ğ���Qy2�N�/��l�#?.�B�HP@Y�?%n��'�>I.O��d�<A��?)�(������ϴ�yv�K���b���<i���?A��?A���$T09Ejϧ^�"-*a睼-��[Q.ɵx\�nZfyr�'Z�	柸�������i�lZt�C�� ���	X���;-G0�M#��?A���?.O"g��l���'E� Nhʠ)%&X�s�JI� {pt�׺ix�U� ��������q���A�ܴ~I��x���1R��д�Ͼ[nNoZٟ�	qy�*܀$�b�'�?����"��� �J1�Łf�L@.? ��	ʟ0����$�2�~�'C�iP#u
U�S@U�Bjm!�m9s���^�0��d��Mk���?���b�]���� ��5��ܒ�EC�9- oZ��0�� 扤��9O��>�94�ՈmE�lx�*]����Xb�v� 궍VЦ��	��\���?1�O�˓]�^��� �_Sl�����玔ã�i�`Қ'��'s����l@��taF,�Ȣ �X�OK�-l�����ПX�f�
��d�<����~r��> ��xg�� Wb�exp�!�M���?1�7���S���'v��'w�؁D	�5���aV�`��UY�NjӒ�$�����'��	����'�Zcuݩuh�j�E0`�A&tL��O������H��ӟH�	ן0�'�"�C��]�T�Дh�2v�:�Zwn�4w������O���?����?�C��L lP
Cĝ0*�\��©C�ZU����O^�D;�)L�u��x�'H��pC�_OД}�U &�T�nYy��'��Iٟ���꟔ 1�~��߉s �@*B��.(J�4�F����П��ϟД'�h�"f�~���3֮�k D	� ��|N��q$
���@yr�'QR�'���'��s�d�2G �edD�
�JQ�f��D�ik��'@�	PL~��������O��Iʜ]ھ�!e������ 0�}I�4�'���'�����y2�'��	]Z�"�>m�ū� =�X�1������'l���r�����O<�����X֧u���K����Bi��=��c#��M����?q7#��<����?	��ʸO,��P��ʅ8��)
�L[0��	�ٴT�,Y�&�i���'��O,�꓈���_� 9z!$ԟK�ȒPb­t#�n��\�D�Z��`�'�?A�(	�C#��q��@tL��p^�:j���'�'z�ͣ�(�>q(O6�ĳ���E��0"Lx}�U�̒��i���j�O�q�2O�ԟh��Ο�#�Lp�nP��Ɵ8'�P�9��J��M��w�������O�OkL�V���%��{t�a"��H�ɦ:/^���Sy��'���'O�I%+��%J6����@Kam�
E�q�H\��'�|��'�fհ�2�d�U�W���j��u��y��'��'�4k�y��O���Q0��%!2�*��#vayO<������?��s�����0
��#��H����R�BO?���c[�P�Iܟ�	^y�j��?�,���â����zs�΂M7R��0!���1�Iw�	ʟ4�	;O�d���J�䂄�+I3�pq�MF��Ɛ:�4�?1����$��-&>q�I�?M@�k�9��8�ׄjꎜ��Ȅ���?1���}������JY,��� �l5�X )K9�M�-O��%¦݃��H���R,�'�>�`�g�Q�*���K��14���4�?�� �>������O���D�5+X|Kf(K0���)�4�̘��i���'jB�OK�O�������1It�=:)�5
g3\��n�v�*����~��_�X�	4&�4P��!n��\���-J��ݴ�?9��?�oI5>��OB����Hf.��@64I$�̎����f�ēO��K�K�M������	�����ߐdp��U$S21�ԁ��J��M��Z�`����O@�Ok,�5W5ش Í* g��@�E/u.�	�'A��IGy��']r�'剛Q|b(��nG/ObR�_ -��YQ�����?������?����� �b�'0ttfF?�D�$!�<Y*O ���Ox�D�<����<�M(x|�4#�ǌ�S�X#ń�tg�I؟(��^�	؟,���k羡�I<>�µ�I�O��hr�Q��fۯO�D�O���<i� OkN�O,����*��:L����~Ӽ�D!�$�O���E�%b��)}BFݓ^\�*r�Ƅ��HO��M����?	+O^lk��@�S�<�ӗ��I��'7R�dqs�԰N�N�rI<���?��"�;�?�L>)�O���j
�*4o�i��kN90)�9kش��3kr"�m������O��)X~BG���
Y !��)��l!�Ц�M����?A��O�<�L>ɏ�D-Q�c���▭&N�i���>�MӐu�ah� ��O��D�V%���Ɉcs
  � �+m()0r,E�ap �ش�(8
���䓄�O�r��l,4��&�}�j �� W�P��6m�O��D�O��� 
Y쓘?��'|�!�K3[3��[1��'w���J�}R�H:��'�R�'���C��`ԄQ2V�n��P(r*7M�O*H`�
 M�����ID�i�������u��.,��\�"A�>�g��<�/O,���O��D�<I��?��#�B���1��D]�v��U;����O,�O����OV,�Uh�(Z\E1�����!�L'���$�<����?����D
7�y�'J��b�!�<H	�����)�6A�'P2�Dy��'wh�PD��=������M�i���>���?�/O��̎y��$�O��䉜7�ޕX�aӀ/�:�z�lI V��o��,&����cy"���ēQ�(�kr�X']��2��^��h o��<��Cy���:_|����$��#�M��8���I.f�B` ���G��ӟ����iJv#<q�O��<�q���$�"�[9�%��4��"y�$�l����I�O��IH~
� ��!��']��:V		41�h	V�i%��'��Y���8�ӄq���U�XC84�8�C��&&b���f�~q���LR�������h�y!�ʋ�A���VJ7D���+�%K�'�m�� 9S#�(^�z �AHR�nn����
�)�]$) �L��'$�qۀ�y�!�"J�*��FE��.����t�Ņw�J��f@,x2JO�E�t��������G��:��T9���D�p
 �rh|0��k�,��<�A�J�
X@�� ����uxb'�ן��Iğ��I��u��'�7��H���Q:�p��c癅8�p5��FT�M'�2q�["B��P��8��"�X�h��ǃ:k��` ��bp��Y�K]�\s|�#&�ل��L0%�ց#���f�G!X�R�K>�V��L-*��\֌����3n����I�(G{����W�mQb؏C���壃0B�!�d�h��ue�an}A�#��hr1O���'b�I;L]�	�4�?�Rnb���b�E�Th��AU�� P���?�S���?�������?�O>��O�<�F�%��*;T ¨KV8��c�:����D��*Yh��p�)��f�V��dS�d\�.5��8^���́�n�d1��NȐlD!�`_��6�Ӄ<����!�W+!�����}��� W��Jυ**\��6H�g�ɾ>LH����|�����	 7:�Ċ�_��D�i£-� )sui�i����O|��._)`�� ��eĺiԲ���|R)�t���\�^9�E
�嘝~�����>	�d���H�4�ȷe�9r��iV��z]��NY(W[j0)��KO�S��T�I�F��':��0��A3T����b�H�
f�s
�'w\L�F�O�^q�&)��P`�	Ó-����3b��AJ��ׇ�*}_�h��	˸�M����?���#� ��`/ҏ�?����?��Ӽ�HI95
X2��9+�ƅ�����'�5�ϓd�
 �������\3A(P�"����=�.FHx��8�B�^���#@c��ۂݲ�/�K�߂��)�3�d� �,�R���SZj M�4
'!��[$4q2慈�ܾ�[��O���ɮ�HO>ݣ��5q�L�d.,C�5��Ś�3� ��`h�䟐�����I��u��'�b9�@���.o݈�Q*\?R�`"G��l-�����U��?nR��IQ�~p�j!,�h<�9.�
�9�L��se���3l�=
T$��	\��(�cj�C��}��o�f�B�2F<D��IaS$���XA�60���i9�%��'�FlBib�F�$�O�t����}���-�v؂���f����Ol�3
�O8��`>ѩ�H�Ob�Ol�0�*áW�9�J͒4�,E���'���8�BG 8v)�@�޸S�=��eJ��p<�����|$��aa�ϑ�4�1�ұ6����Ł;D�`�!��3"e0B�Ҳ!�T�Jѯ8��c�4v��E8uf�BSB� �HX&SgЄ�<a��8R�v�'��]>y��)���1qkоR�%D��
R$&� ҟl�I�s/I�	B�S��O@��֩ضh! Er@͆#:��Q�>��T���OJX�Ӂ��7W�L��p��D��ոO��2qa�O�c��?��$��	!�%�RJ߸z�X���=D��"fT&Z��z��\��af�=O�,E�D���	v���K�5f��Q��/_�Mu���'Ab�'���R��,b�'�"��yW�)R\���_b�0����>s�1O�����'2]X0�_�51d�х-���2�9�{�-A���<�c�"d:`�����H݊!��.��'ڂ!1�S�g�8kv
q�U��"B���A����|�NC�	��¹DcK�Fc�a�� �5r��"|�ԁ3f��`�t�9IE��y��K<��u�q�6�?)��?��gG�.�O��~>�R�	V�v�{�LH�#>t%p���'GvxC�I�a�2XYЧ�lD���ۆcb�P"��/�Dy��vZeǜ _��,��Eǯi%���4�O�1�v:v@`���a%P��"O�<[�ᑸG�$�BU
��FB�*���XW؞�;��߮0*0�]�6�j؉�f=D���ůףmG<�0 )�?Oh�Ɋt�%D�d�vI�)��:E��0z|� �?D�p�P�گHղd"3�,j��JDo<D�hK�FZ�96���� �1>��[DJ9D�h�A�[�Lq��GH��K������6D��Y�`�� b�y�Ȁ�	�:�l5D�� �Q���қ�r!�$�	=H�T,��"O���֥� |n~�BS)�.F��"O�ăt-��"�q����Lx0̉�"O���#�3u}�1&�ĕf|~1�e"OdA�@M�2�|�@fkw�Qx�"O@��Q�U$FLbx��	��~j��Y "O�u����Ag�9�v��1[�!�`"O��O$P���Yp�y�b8#�"O�ԘA
�U���;�DF�Yo�	K�"OD�ӡĔJQzy��l�5)rX��"O:���
DN5&1h!k�@� �ڰ"OZ	�%��_8��J�5$��8��"O����k�X |'�˚vwA�"O��#�O;?�*��"gX\�v"Oj� 7��	�h�i6N!;�H(b�"O.HZ�$Byz�m��B�S���(�"OL�ۂ)�+E��ZG䒉X��p� "O�В��	�a���6cNeްm�a"O�1��H77�v�Tg� l��<`G"O��I�nƬ+��ȁ���%��"OF�z�/��DJ��Î6>�Mi�"OJ�1A���C$�	+��f%��`"O�d��B�ZY���\@CT��3"O�̙�A�p�hIG-T5��W"O.�@C0?�����f�1%{�"O��b�L�gY`��D�6q-~x�!"O�lǧ1�� �5�^"N�c"O",���[3���c��4Ɖ&"O�+��@DD����K6n�k"O��{�e�Vb�P�'cB.$�$� "O%�)0!$`C:���+�"O����mܣ?��h��n�r�؅"O�Ԫ�
IP!��9�B2&��A`7"O8]!ᏎO|�g�]� |� �"O*q�*��tpu�D�>���"O��wT5Ob$�A ���ڱh�"O|��DK�< ��S����8�2"OV���aӇ-� �@��T��P��"O�!C3��0u�1+ʎzv��1�"O�0rӃ�o���iR��:���"O�X�7�T�}����aɖ�,|z5xv"O��1� #'T�@���W	W̤4Z7"O�@Ӥ B�,�4�� ʖg�F�#&"O���H�Y�0�{��6�*�&"O���-L'Wɒ�r��$4eL�"O�	(����9��x���T�R���7"O��ZEF�mv�W��rr���C]�<Q ĝ�+f���/̷R�N���_M�<�� �*�B˧1���Ӣf\a�<�5&�:����#�N� ��D�[�<��Α%`�m@t�Ӻ=0�H�@�k�<�0G�g�F���H$�X�"���o�<�&��Q��؋7j��
�Ta�t��q�<Q6cݣ-DB�k�b��o�b\�㈙A�<�QNA�$�0�HG�R"B�ލ��ORC�<A ��p�Jq����ZQ�a2H
T�<	�-	I�)г�LYL�2��z�<�e%ۏz�`D�֯J8rp����A�<Y��\<B��t�|^1&
�u�����q���P��0	�͙DR��*���I"4�&�O�����ͩIf>�����($[0		�"O�8����An���h�o�@Z��d�4Y��b>q1�E�RE���b$Q��X���<D�4C�&K򞡀�.��pF-KBBF3pt(`� �)?Y���l�S W���䧀 �@%֨F2��e悠���*T"OB��� �69 [�k|@�ɦ'�]��qk���?����D�,�B���� � 9A�6���c܆d�P�x�'Q6���k̦$~P�z��O@	'$�x��Ș�/�phw�00�b�$��]n�I����	1�5�	��T��SjT]>ƭ�J<Iu�Ĉl:|�Y7��_�<��l�����Feڷ�Ќȥ�42
�p����M۳�`).��>�Q"E�)�>P���є"CTq��@)]�R���/}L+6\��j��v�Ӻ��Kx"��#��RNT��# /��ē/�9��6� I��)I) (Q�$8O�L�3���@�p�C�� Q��A �`ǜU��K@:"�>�E&�}d��sf�",OD|'�\>r{ȁ1��إj�p���G g�ެ��,�>!Z٠��v~�X9� ��E�6-��
��ĻU����=Ig��Gܸ)�2����� U�D $�L���/F!jil8b���b��O�Y�6�O<9:����C$/��90���,C�ő��_�n�<E�����5e?x�<P�A�$�}��Ш���������=1���?�H�<vir	�A�@�m>�����f����>"�,��#
!$�4!��'ĪX�wO4�&ekF��[a�U_p|!�oёj�( �6�π]���ςcU^P�m��A;�X���}�!E�U&1��t	� }�='����KA��ay�G�a$ȱ� N"��d�U��-�*E�ح"t��:`pO�YA��5�.��ܓJS�dQ�P� �'m
A��X���!GÁ$�$}�Ю@�P�89����\�4�뉪3�p$� e�-a�lڧA��s�*�:�W�I�&�����=��D%����k�:k(f��C�2Xz`$�1!D�������bI�����	Y2Y���IX� ��ɕ%R2e�"�ѽS���B�ĿT�B}1�f� T$y(���A���o�)j<��e��P���8�n%A�xp�V䟾x�qY2 .�䗮X�qX0$F�shvQP��.���CD�e���ɈЕ8�
s@ �#�"�<8z�#<�O_�Q�4�)uf\f�A�C@Uh~B%�k?*�8c��f�p�ƤLh}���­s�Щd�7�Ju�@-�7+�ў���Wd*ĲwfA�[z`(+R�1�~DB2�R;������b��"?��烲CJq�eN[T���c 3W�	x��%;&4��$6v�2�r�]�I��	j�=�Baa��$�%W=�)�1"\�wQ���MƖ�7eU%Q|�!+CΘ&T���I$���׌��3�,��IQ�qQ%�8�&�xFf�-��>���9�b�=6��uQ�7����gҨ'���`��'��i��(Y�>qr��$9���,��|"r`��S+2|��R-��I�c � ����Ytl͊U�Af���{$����A�ƌ��"�aT�#���I������7g;�8�f��jmlD��!M 
�xq����-N����v�ӧ��u�%E����^�Ԕ�f�v $9'�/[Zl���<r�xݺ���>���B�E�6:��!c�i7��}[��	���E��&|h>��Dϑ��3���FR���+��1����wx�����S9n!�(ص�D|j3�X:���I�2|�DԗV#ģ�E@�!ۄ,� ȕG�=M��ژ�M�R�#^��Ma��
9{�a#ALd����et�XɧO�9 f���;��I%ǜ-L�(��j�,Bƌ=�e/�����Ĉ��l��!b0����1�L:,����0���m����7}�iF[�����O|���
�}Lqrc��� �%O0h��QA���30�V`x�x�D�2^aX�˕mڊ+�:���4��51�Nx�@�>�؁ȓaº���'F)j������D���K�+��ȓ9k��S�Hv�t�B��������y��c#D�D.�`���I�On]�W �H����JK�K6ph#"O�\�k��kԪݓ�ZRB]rw"Ot�1����s)�c@��a&8�"O�Xb5@F�<<F�G��'s�܉"OT�r"�6B?N��d@� ҈E��"O�p�Wg�43��P Q�a<I�7"Om�֤�G�p��B �?3I����"O,e�R͖�7$�ΐ	-�<Z�"O�4��a��C��=���"OB�Ȁ�Z-C��x�鍑Y�M�0"O
@�)(Y)�p�䧈<	�U�%"O��@J��1f���:��D�1"OL�P���P��Y��DT��<b"OP�(!_7����C�c�"Ot)�Ө.2�(�����]2�â�>Q���'�O���� Gy}�ǡH2��QQ"O�8qϏyب2�/L'L� u���r�N�z	Ó"�@E���=gr��Ə1y�t�}��� ةSɑ�ɜ1G\9W۲��b���5�!�ğ'm|�(N�A�PX@c� k�x��U:]g�L��
:�!�	.pE�aɑD,D��Ð׉(�l��������!S��*}r�VS?4�&N<���T�&���S�G<@,���k�"d!�U`�;%f4vTa�$j��[�HŁI<�I�,k���>�O�!�p�C���c��$�
�s7
O \����0��k�S�#���c��CC�K3)�|��0�7hX;m�ĸ���;I�YA�9O��Sc&�G��O�;s����$d��X�P�F"O�`�@eE�*v�i� ��+�FDh7�>�DA˿^L��P�x���H=B�xxr��4N�"EPI�%�y2`C�V݈�Z�`�I��E��M&4&�d�D��6<
q��'�Xt QǄ�
�U����@Fh��'$*��&ɊA��i"��ʏ6��iY5��zi��X4�<�O�@%��d*�P��0�b�J��'+h��`�`���#}�
����:���]���%�d�<�w���U���rΜ�r���t�V��;U���3�q�)�S6}�T(�'J�t�T)L� �C�I9]�Q�6(�(��x�'MIAqֵ�5�8}O��6���}&� 4����B�S���|�P@j;�,Z�@��8�5H�"L�.@:5�ׯr!�!����[�qO�N⟱O��!(P
�$٤jS Rpl�V���p<!d��I	Xc�d�rfO �(��+Q^�P�j�� ���F�s�qO�>ei�M�l11C���;(f�>}T)('f0�=�"��ɪ�$�N+3��h1��x�D��RnP��
�N��UB0-�f��p���Id���=yQ��&6�r�<�%zΑ� MR'+�\e�`NQ4l�m���&$�`��h�]�,iH�.�T�(�4ڰ 4��l��uW˓����E���7�$eC�V>�1"O��&��^Q�!!ŕ�#)���"O����I�M> [�DD>0�-C�"OZ�8�GC'L"�����A!l$�h)"O�|a�B�9�<�{��&t��mS�"O�I�b'_�P��uʤN�% ��8�"O$��*��6�B�h��qz�Y�`"OLc��G��,�d��0s�cp"O�L���*�"�H�]~�إ"O����ޤdr���L��eZp���"O�) T՜%���Q�J�*>�z�"O��R#�X6�" �bJL���(�"Ol��j�#ht���)�,��"O�%��'�@@5�3Ȝ_�lJ"Oѫå�;rc����խ#`8\�"OY:�3FjȚ�eRҸ��"O�E��/�M�rL
���֨8s�"O�l!���*	��3P`׊w�<0"O��م`�L��U�0��%`PFd�`"O���Ů�e��v�&,�,�"O����S���2#�x�Y�"O�()Vd�3af��pG��.t��!�"OR$�E��-*�h��@7�Du�q"OHP�Gŀ�U� �d`Ȉu��@0�"O. 3cA�S����N֕'l(���"On����ݻw�,�#!��O[�bc"O�,��V�!�浂�-3,R���"O���vB\$X�&�W6#���	�"Ojm���$(���c�KZ��ui%"O�%��N�!&{V;���?nN<ۃ"O����"��P�p�\3WLe��"O�=���]��tYU��DU<��4"O�İ0`1������NZ- �"O�83U�I�ɍj,�m1�j�7J@C�ɰuA����]/-���`� D	3��B�)� �q����M;�K/3bf��"Oֵj��_�IhB��`CG�?��]�%"O&H���?,���`���m�4�E"Ox)��~x"�S�BY9��=��"O�`���K2a�aX#�;*��A"O�YA��S>(�: ����;����"Oօ�m��$��hEH�&��0""O�-��ˀ3�:��7�><0{PÞT�<i�@[*P���fҾ1���5D�V�	{d��#��.�&0Hv��.�Py"A�882�0�g^�2w��"��
}�<�Ogt&h�qC�-?��:C��|�<����g���P�N�uf9�F/[w�<��F�9��̣7��$wN�aG
N|�<9��ȷ4�⭀�AZI�Tq�N{�<YG���Q@�M���_���	#DV|�<ɑ�M- ��� �I������u�<�a�w�8�;#�&P�����\�<� �F�gW
�sd�ދ=�����N�<���pp�xp�`M�f�@�	ǢI�<qEƉE�b46�j��lqD�D�<�c�
4/ސEx�M�K������v�<i��	\%ĐYթ�2�����Np�<���ߔ�
qy3��\n�h6fOd�<IA 6�1���q����bH[�<��@��Mx�iQ�#�
E�P��y��
�usDC�!��0���%A"�y"ǈ)s|��u	�:Į�S��E6�y���`�+"	<,��I5��yRL�7mޜ�A-�@E&�Q!h��y"�&[7*@cÊ®D:@\��4�y�D�9hp�е#��Q$����y�B�v��a���ٌm� �ٷHB0�yAӊ��a�C�#j�ڈ9�%�y��[,q�RC$�F�h�� �f%ʚ�y2�Ʈ{�>]"Ǖ�Z�REOC��ym�
}�|�� ˕Z�6  ���y�n̦�dqq�@=ZB��2"oĖ�y2�CR��&d�9N��9!��:�y����kޠر�\ I��Y#r!���y�L�,�z�x���39��l
���?�y��H�<�h w��F������y��L�<�nxkÂ�%VR��匐-�y��& ><�A�i�4�C��yjC�.̉x����։�2��yR"�>�pѴ�*rc�;RQ$�y҆[�}ژ�# ;j�n��KG��yb� �J��f�D�U��d�D� ��yr��\m�A�gG���l�y��_�U�ɛ�7=��\÷h٨�y�LЈ@����V*�3�B�Y'O���yX$#�xš�I�#P��aGb��y���]�~\ڥM�qV&�aN^�yB���H��!�fa�A(1.@�y�
,9w�u��@��_�t;��^*�y�	N�$��dZ@z�ߨ
��B�\(�y$�΂ub��2��4B�>P�H�zT��vl����n��B�	�b�!
�̓-7��텵Z!�T�.]�gG�>̪u�@l�iC!��(#STXa��W��"�@��6O!�D�r4i�Ο�5�
<Z3*�-H!�d��7&��H򢀹p�T���#W�0�!���z�n@����ԄH��.$2!�� &���Qh y�v� 4��"O lS�Gl-rphV9�dɷ"Ol����6��Y�Xn�,9��"O(r��c��E-Y�p��\"O�m Rft���yc,����J�"O��S�"J�:��iQ;"�nXHb"O<�Am�7)�`X�玀��U	"O���dO8*L�S�+]'G�:��"O\\i�-Hs ��!�ʙ�o��$"O��S�2r��6�XrU٫0"OVE*�g�T,��
A��K<n�"O��a�홝#d��'A]�]	^q�Q"O�A*�L���i� �'a��Y�"O�	�!ك\F0�����E�4�D"O P��Q��V��"�O�s}v-��>���|IŐSJ�\�sϔE4���$l*���/F�_� �B�nT�,��ȓ65 c6+1��lg�A�z"x��Apl��,�7>�}KT���ޔ�ȓ|� S���{W*TsA�\)]����ȓ\NR�r�P�o�n|g`C�6��хȓ�F|[�o	>���b׬�ln�����^��(�� ���
�a���_"��AV�c�`�i�+������:�6�a�ѩ)�bɸ2,8X+|9�ȓ �P�£#�[�����M����ȓr_\����ǗJƦ����]e�8Їȓls�s���|����n�_��<��Rq ���G�>~ܠlҧ�N�I{ҥ��J�5�5(��2�a��
 lU��8�2}ڴ"�/�Yu‾MZ�H�ȓ#8}���Ʀe3�%��˴3���~aZ��`J�9VluB3"Z�f$-�ȓ9�t���ס%<��F�.���+Op�� �1�FH{��� v��8��A�V�h��e8�lIq��8�r���N3t�����?����a��%�Z��`�pM)ǉ�H�>�K �#U�`ȇ�Z��qp����a# ����);� �ȓCr�k��CT'�j��_�l�T��A'���G�A?�������V9�ȓG�$��u��?b��co	�b�`�ȓ3��8��T(^X��s`�D%'�F)��~6<# ����T�v`vE��J@|�=ci��KG8=?��ȓ6*�Q,�
ў�z�� #�H0��#���zD,���	�<���ȓ+l��W�-5B��w���#�ȓ�|`�DI��lR�!{�Z݆ȓ:W�L�g�
�k�x�Е��9ְE��V�RP>�d `� �S<8���,�$�����ĆP�Ko@���+8U��!�a������52��Ez"�~�Ȇb���V�ār*��{Pn�Q�<�VJ\<X6����P۬����@G�<y���P/�a�d�2bi�t�M�B�<���Ⱥi��@a�@��Y����/�d�<��m�6��"U�0�4ܣrËg�<A������j�I�����LY�<����'O^�" '�4�|�p��l�<ْh\�[K�)�+��e9�E{fb	p�<�E��6n���ǛzW��*	x�<����Pp"F� #�`iV�IM�<�V	5;�����dB�PHJ�<� 4	� �!�d���N	f�Q"Or�ՃF�h���%d��#e
h�6"Ob8i��۝
}���ce�	NJd��1"O��Y�t ��9�dL�6B0��"O���)�ы")�{�@�b�"O*�`��)i)���a�9���(C"O����%�^4�Taݲ����4"O:Q����3fh�"6��6�Z�0�"O� �>����i �;ͺq��"O�(zRk�}Nfx:"H�7&�ȵ"Oz�&""R-�&�:'Dv�4�yb�(s
�p�@P�@F���1�y"	��r���Z3;J)�g�֐�y�dN�tD�u̍;9>:��GJ�.�yr���@�(c6#C�5�2Ǝ̎�y�j���l����B�2W��p�H��y��C�ȄBäJ�S?�r���y��F�#�<�����!�ȑ+f�Y��yRn�2��1d�H�	�D��M�y�N��.�N�k$V���fώ�y��2���[7��9g���D̉��y"�Cb�z��1/�����T���y�L#^C0���L̢&�r���gֿ�y��$�$|c���/�2���y"J���T=�e,|�v%��H����x�%u���q�!��� 候�*X��'|�#$�-fl@��F_(��:�l�Q�8�M�"���A �L�m�,�#�=D�` S`�7?��|�`a��k҅±0}BF-�S�''G�ؠC�^^�PI¯N�a��ȓJ�T8�)L+F�����jW�}+�0��} �f!X�*��t��BO�4x^��ȓd4�E�Rm�1lg8�����L���ȓl��,�G�?0K�s�ʔ�>h��ȓp� �Y%L���
����ȓ7�H!e%h���S�k��.��ȓN��-['c4,�Uk#1vܐ�ȓ.���C+W�RL��#{� ԇȓ^�.T#iV��e�	֗Wx�-��G3"yq#�۔\��`��)J�6�DԇȓZ�V�#Uo�0��� �גi;D��{ӄ�Z{��b�?h�Zp�"O;D��+z� "�~�����b�B�ɜ8
�Ps�T�2��$�M��B�ɀu���W�u$��E�ϮgބB�I=�����(]0�J�**.�C�	#-Ը�W�3l���zGI�?l�rC�0kB�uKm `��R �B�	�mX0�і'��@�#�MҔk�B�ɔ!6�4���n�N$"�%I�B�ɏ$�.����&a�T��"l�YbB�ɯa��Y�'ύm�||k�@ʲJ� C�I�P��Ix����`P�8�/
�9B�Dn�A��7|r���4�Tc�$C�	n��-ƃ�r�9I ��3nM�B�*0����#~�^��5�\�z�B䉾�pw��<�8��]�rO�B��X�!��E�5������ϯP��B�I�B���j��*Z�E�$`��/��B��+2 �P���X������Ug �B䉾a����T/�3�f�b�lG;m�|B�I�	]J@;c�ˣ\t��!�ls B�	�4�4�H����_.V��$���Y�$C䉚Eb��dȄt`�d`���+j�C�)� �Q��
�/��K�,^x2�8`v"O~�YƉA�v��P1�k�~K��"O�����s�:�K7k1HI�S"O��9��WH����Z6���""O��#�Zx��1��p��ɐ�"O̙� �@�6AN�9T�6�A�"OJ`�eQ;XD�ISu�7	��P"O���5��0[����Jަ+�
0KE"OzT`�lX"q �t�Ei��![@"O�q�X�x�r�r0fX�K�4�:r"O8��H�0��Ɩ*q����"O^�����U%�P��:)&�i"O��5���m� ����'^5!t"O�]yf�;�l���%���QR�"O*���|굓��<�,���"O|Y�%�
�t8�%��6�6�"O�q8È�j��1DDգ^�\�8�"O2	�#	�83�(�	��8N�^�a"O��)$�H�,����Y��,y�"O���S� C~�����j��V"OZ���/y��$�_�|-�1Q!"O��c&	(7�9a Tz+���"OE#gDUX�c�ڒD2ź�"O~��ࠔ� Z::�O��5��=+�"O���Qv���OM��u3�"O�s�¨5 <�C �[�21g"O��af1PG�0�0����{"O$Q� B�r�^D�R�0DE3"O�h�k��H��@C�ELd��"O��3���bcj�S"�1���"OnM���� &4a��S��=�"O =��nߏG��p2��:�8�b�"O��˧A�ed��DT�nr�4�G"Oz��d
%̦��#C�h$m"O���PEK�.�(����݌F�0A@"O�-	��$..Ա���̊Y����A"O�d�2�N!RrD�X�gC�,�*���"O��(r��$���E�~�2MG"O8������:"�)��C�4I{nA��"O���u&??���-N�G�
�!�$KO��	����T�,R�C�+�!��&'`	Qs�G:��E	��K�J�!�$�%@}�C��O���F<�!򄞹�����A��ԍ�d�N�=!�
���>�JM4h�2}9eJ�"O*���l�p�t`h�lB<N*i"O�����^ق8[�dQ�L
t4��"O��ɢ��40�b������"O��qq��3r��Ф
ɛӸ%(t"O�%����9B��v��(M΂Q�v"OrQC"
GJen���ä�h�"O����B�D-J�
��_�n���"OncD��/?��a� "5����"O���2kY�_O�<{0��d����"O�9�G�ŕ*��F!6�� �"O.��T��&"|Q��?�~�#�"OP D&Ǎl薕9 f�����"OF��&�٫g\���`��A�֥�"O$4���(`Aj�#II"#����7"O��i �PS�LБ���>1�^0t"O�X)�
Nx$��� [;eߚ=J�"Oʔ���kJ!
�Ϙ8)� �x�"O���(W�~�Hr��Ȇs����"O�X0U�|��K�(��>tc�"O� �HR��kEVI 4��K"d 
&"Ot��CE�!�t�Q��P��2�"O�l���*3܂�:��^�m�Sf"O2�
�h�� �ţ*�D��e"O�AB�����t!dE�-�3�"O�P�⅕��p�S��ױ]���"O�x8'"ĩ^B�(�!V&_�b�S�"O����˰�x�G��1�0I"Ob��p-_�Э�3��?%�rp"O�Ah��� 7���L�"��"O�i�F���P�� ��O
~��C"O��k3�V;K	`X)1�#!Da��"O�U�F[���u(�O�k���C"O¡д�W4��X�A��b9R�"O uh��K	
D�tHoŎu���c2"O�5�4#@2P�:� �A:��X1!"O&L�i'�����&S�e+a"O�͑f���%��\�1i�����0#"O6tI��	_�PZ�X9C��i!"O<����_G2��!H���MI��*D��t�%T���Mڴ^��LYFJ'D�PUA�gи3@)�82�E�o"D����g��l����0��5r5("D��C5��x.M�j݄>��be?D��7�Q'�Y�h�� 
���>D�h+�__�m�V�W�����Q�:D�,x�IS�Q��Ai�V!B���a:D�<i��լ[p��S*
7�����=D��@Q�@�8�P8I���;MH�`a�M(D� QP� 2Y��P��=���s��$D�\@!�,fFV�k�kF>X�� "g-D�|c��Z#/�|��b+G�%/\$���6D�|1�h@�x|]�����2:<l�Y�y2a�7ex^��6��/$	ڀ�B,�y�#C��r�Q���а��y���H�$��@�Ͼh#z�x�Iû�yRH
�0�QǞ\0k�%��y��K�A���d�G�*��%���y�-A������n5T�0�S%�yү1R�\����[�w^��0ccR�y2��=	|� ôx���Wk�yD�J�b��:b��:�� �yr��]�.TA��5TFx���o�*�y�S�\Q��[��AI���Xq�M3�y��Fb^�tI!̟US�|�7�	%�yb�U�U�ΘX���S�ZQ!�I֚�yr
�M�����(Bs�ER��E$�y�L�?�����A*��=�y�E�a
]x����.���B�K��y�HP8
}�E�s��)'llMU#��y� h�Q����i>�l�$P�y2���MF����Ua^ Є��:�y"�թyԪ�iUϓ�a�\:uh_��y"I�:f�b`�"JE���㵇Y�ybfM�M�1����+�.H9�o��y��Fd%n�T㎀9�d��C�߃�yR��+&�UY/f�%��A��yB�J�Z�2�x��[(]�P�R�T�y"�� �,(� �Å^0M����yr`*�u��PS�X��҆�yR�ݩ��$ �D/x-�+f�H��y��Ɖ�z@�m��DZ^PB�IB��y�f4<}��x)�:=�V�S�)=�yrE�6u����T��I�Q�QhҌ�y
� މ8���3l���fЌ~�B�"OZ!c�a��0�r�Ȅ�	�|�x�@�"O�%RuG7-G�*�#sڲQK""O�ԉT�E�
��b薔ň�s�"O��1bHS�Sl��*�'�;#�XD�u"O^���Jl4D-&��'�B`�!��U	�ms��۰,\�ȹ���4\!�L�*�tհ6�ޮm�^t��hÈ.��"j�LI���O6HU����.M�;%�B�IP22(2t��✋p�	R�2��d�O����;F䁘P��4 4�D�UnV4��5�����fX	O9�L��Mޯp�ԅ��7	0䢓�A�b��`K�K
A�ȓ��5IS��OJ8l��n[0s�Hq�ȓ}0�a.òU)��ЄM�����za!�c��"����/�=6o⼄�Y`�!#�%��Hl�3=z:�D{���<��H�0���Vm
3j��	���G�	B�D!q�O�h�})��(�A�?D���F�p�\�2��d�����7D�ԣ7�D�$�HY�4�\�RC���4D��86��pԐPT�Y3v�	z�3D���#	ƑQs6��"�D�Eo�E�a�O4�=E��H9\�p�-
 %H�0��1S��� �"����v��cȔ�\�@�=�	ÓMq��3ah�9L��tɄ�!}7�]� o���M.M����r��.�IpwKêT�nІȓ׺�I/g��4�^%A/��ȓL�� ;eA�Z|�(�`�*OqZU�?�ӓ?ޔ�!dL��F ⤤��%L&=��vQt����ǽFi�D��' ��%��b6���@Z�DW`�������H�����_�S�ʹKr.K;��(��\I�<���8'�Hb%[8O��\F�<�Ԃ�7$U�h�c��1�r�W@@h<A�K�^�:R�Oc��i����y"�_&u} u(�-Q\�$2B�ć�y�a�Pu�h2���<I� �$�����d:�g?	�ƌ�m �[l�*6���T�Qq�<�B�ȰF�p�J�K�&���� 'o�<�f�9Ib���Ć	z���e�P�<)4�C ;�N}�5	��X0a�`��O�'�ў��Fa��,{Di�3㘅���H#`�I�<yc��7F�2�F
Eڌ���H�C�<��49�Z�2�l��m�6ԑ��yyr�'&�OQ>5���6W9�Q�� ^n�����?D��s�
ɛ7n����xxy���7D��bрF2rZ̒��W�L�6D��X���+@����耩3�D�h��0D�|�b�%"��BB*�8>�jW +D��#VE�������$>�f1F�,D�,!���gO9��
X I�n%D�$ MR�r����S-T�$�"'D��2`��S�VE���� ,��07�$D���%ϒ�>���s#-Y�n�`��&�'D�X',�>��M�t�׍pl�(���&D��Si։f2HP�,TuJ<����)D�dqdGN,8�P���!�4� ̘Q�<���9}b�e/ɢ"@L8�ÌL�<�v��o�&H�A���"��t��M�O�<a�Ͻ[]M;h�G��x�A��a�<1S�R%W(�Y��� ���ce,XH�<9%��&N�{#(��L���V\x��槀  �[f�gh�	���Zh�ȣ"O����A�=o��(: f(1����"O�Iq�h���)d�^��ed"O
�;�,/1�`K���T��+w"O-q�F�\
`��fϛm��좇"O�%��$C�V�6�,��g�<��1"O�$��A^�����+�� �-q�"Oj !2Y� �P�A+\  R�q"O洃G�8mV�YZ����~8p�"O�Թ�놁4���R � 8/Πd��"OpI�v��$�H��X<�$(�"OR)c�d�%|����QE\��d�	�"OƱ��Ҭm@�� ��9Q��mٓ"O`3�'S�q���j$@@�l�.E�W"Oؽj!I\�t��E1aO�T�9�"O�@8�nN	t�P��?#(�)�"O�(4lɚS�jMIa(O7,�	6"O�)�&�������D(P�PQ"O�D�a�K���X�͒Y��h'"O�h�a[�M6��6hP-���a"O�\����jV�y�Aa=14��;W"O�)�ē/?�[1!߿M\��e"Ot8��@�l)�(㠎ɯs��B�"O��0�K�-b�JR��=�x��V����#��#͚�,��l��o�,��B�#b
���c틶-�`KV
B�[�ZB�IR�
d1���"-�TY�$C;O�B�&bs�S�mH�(/ؐ�/�
��C��9
��H�N%_��ZUH��wbC䉻(��+i��V�h�i��^��dw�4�TU�U�b�Ǝē`1�I�5//D�P:�-hԀa��M�*��	J/ D� 5$\5:�X���'r�U��#D�����O�P�J�#`�;D���i�!w��IP�{�ڼcrM4D�,:4B�9�\=:��ml���4D�P��Hi�]b�ӣ+[r�PO'D�0	�9�|��ê�]�\����#�O�扠 �Œ��R�%B�����V�C��;�6(H�l�2y:��Kٽq��C��"j��!��K�����՞N0�B�I���4x�-ԟvx،�7�ѯJ��B䉟d����D
�M�<3d+U /�NC�|���( BO0Y`�U#�&`0zB䉈v�a�źn�⑩�� -\B�ɋ>hV�w�YH@���F��c+�B�	�oH�l�!�@^��D"�7`bB䉀 TK#��?Z��I3�I3T�rC�Ɋ���{�'X5h��x���
F�C��.ưU;��5N�܉��F%j��B�3g˲$ʒ-�c�s$)� "O"��q"��eX��ȯEx�]�"O�ݣ��Ƣm%Px���۫WszQ��"O�8�fU�1¦�q��Q<4p�"Od�$�6+��h�EֆTl� �"O�	���� � rue��7� �1*Ot �Қ-�TkM�:���K�'�Pl�Q�V���2�AC����'�25Rԫ]4!mҠ�Q�װG���j
�'0���M�(�8�a�i�2��y��Q 9r��O��z5�'��y�]?5$(A����<Mr���yr�E���a�7��<�n`�F'���y����4W"�(��C3���ö�y
� lDC"<+Z�Q�eҞ4ْQ�P"O(	I�d�'Qj�]!�����]�"O ��M΃.&$D��ɞ�p� q"Oؘj�̕Pl)r�9�1�3"O� 2�� :5��>lc��"O�AЦE�y��(g��vb��+�"Oz)�a\�מ�Q��#+U6�)V"O��� 4�����&r6U*�"O\񰀨{E���b�_�u��!��"Oʥ�DL�Yg�	AU��,Z4� �"O�q:���<&�{# JK�Vy��"O��Q!��=�D餅�'�R$ٴ"O�(㢉�P;� r��D(�"O���A��4~�@�▏��L��"O��3�^���JO*pv܈w"Oȵ W�ˠp�bX��.Z�EN�`�""O����r��A��π
�0(8�"O�5�6Ǔ$"�~��uF�}��0"O�X�7��x�����"�2u�G"OƁ�p�ɉq�@1�l����"O,�@�_������L~P��g"OT��T"RLl0q�iڡ(V~q��"OR���Ԁg��m�bϝ<:���"O���c�5,��0�DL�)"�"O�Ap�0]�"ȁ�N�,F1
ę�"O<��抚Gq�n��#%�"O
�u�Y0+�-SuN:W)�s�"O@� �����"�x�mM�\��p"OFQ���يF���[��x��"O�u8㘤��M
�j��E�BIc�"O��s�.	<V(B��qI��A�l�Q"O6��dEI�0%P􊐟?~8�ӕ"O�i�� Fߺ���h0M`�y�B"O���֋�#>�%S4���dBtX�7"O$���AӀp�*����]�F9ҙ�"O�i���&|��j�g�6����"Ovh�pM�C�.�P��$�)�"OJM�`&��u���{���4�V�r�"O\��Pw���f�5�P�I"O��w&��&�e�կq�^���"O��� &=�,����`�RD"O����_F�����J�ot2U�R"O�]A�]X`�@V�,VrA�R"O$�A�Q�I)y���A��)S"OR�Kg�:��T�QC�i�����"O��c�TΦ�k!"�'�"���"Of��bΥY�V�b��ȟ���["O��F�D�3��y9�&2"��3"OR��B�.�T@�%����X�"O8ݚ�̿9'�x�p�G"����$"O�Y6j�W�l��d�Eq����"O���u*p��Ru'?n2�xP@"O�����.��1�&8=*d���"O��B�خR���eT.�`��`"O.\zWB�"�����T	���"O���� �(���(t�R��9��"O�	P���7	�Bէș63����"O�IكEU�>FhQJ� ȧa�d��"Oh��q�Bk���HP��$AZ0�"O���Jn�X�".��D?�%y�"O��+R�Ls8�@�MS�B<�"O!���4{*llԉvݲ"O�h�"H%�r+��\t��"OhIrr�[�Ψՙ��(Y���E"O�  z�	�?F�>����=���@"Ol%(�(�
o�Ř2cU��bs"Ox�X�*��:�6�BT@ �h�z"Oj�&�� Q��q&�'H�$i�G"O޴�@�Y!'j�9!a^*3��q�"O����E��5�jH���d=`P�GZ�<��#X?N�~L3��g����,�Y�<A�%;J�� �/ڵMמ�k!�A�<�t�+QQHaQ���S�N@�<i4���N8􀫆D_�~�U���U~�<y� B5r�%q��G��ʑ�|�<	�a�I���`�/فRmHC�%�z���䓝��S���L��%�=+���`"Opj`G�T޸)zq� �CLq�c"Or=��g�.qU�xn�49�Má�'�z�ųY�8�;�$]�Y�"���'D��)��)uu��RśSG��)c"'D�@z��OU|�	z��5I���)8D�$�E�7�B\����JM��� D��)UL��c�y���H��|D��O`�=E�$�]<g�Tu�D	�
&Ma#�-�!�$X�e�-�3� ����;U��y2ቍG��2����ލ�V�Y�"��B��)�1�'Wj9�d�=L�lB��<x� I���\q"V�i�B䉹L�عI��E�*��|���5'�C�	 ����,@-A���3��F4�C�I�jW��q���+p�Lr�B<D�����?�`83q��0d��s��ħ`�l���OD�S��yǕ�V�~XS���}h���Q���y2 S�b_���ЇHg�\��pJW��y����hP[�DZ�d����	�ymJ7Bpv8C#KگQ�ڑ9� 3�y���`���P�U�FY6!���y�Ĉ�!���`���[2U"E��y�)��˞��%f)Tk���ۉ�y�[ ug�t��CĨM ��!g-[��y@��y[ʄ��IҜ?�
��	��yRh��JSD���Q�:v��f)���y2J'u�Z�4,J�f�D����hO���d¸ �~�r�E̎	�45k�LH1F!��}���1"m�d�T��$f!�p���W<rx�8w �Q92=�'i�@�S�F"�:��V���0r
�':.�i7Dǖk]V��Z���	�'�����o-6TAɵ. T�<�	�'>��:U��(q�m��X {'HUp���)��F1s�|K�K"��]�֭��y�*�����,f��q��N�O@!���A���:��3/ƀ�xUH/@!�Ă^��0b�f�=3��5ʧ	�6_�!�"\N<�ğ�����Ϊ�!�D*h�ne��-ߞL4�q[��-D!򤚱�`}�)��#�4���˓2�!���x"��lM~��!jA&W&w!��F�8\[W��	j��=�U��1�!�䁳%h��ؓFT�`��e� C��|V�y"ቪi'�E�4� �!�����B�	�gN0��B��U��<��a���C�i�	�u�V7h���o
a�QY�'���8t@�Bu6(��բo,���'�B|��L�M�̹y�I�����' ����%sF���
�(�`b�'��jª\�2O,� S�y�b<Y��� <��e��M ر�Sf�F"OT�ф�*<F��X�M
	�ĩ�"O�e��!x'�!;�,ӻaF�ZR"O��j�bbJ�TQ�˔uG�L �"O.��U��'$���(�>ȼeJ'�	U>e�c^2>y��ط/�/�ny�� D��A�k^(%�ֵ�f�%R��xt�*D��$ f�����fל6�����"6D��q��%�T�f��:bu�U�dM3D��	�,��ȣc�5N��E�/D�((�,�3g�!��/�6'`��iW�+D�����A�����݄P�IX�)D�t�p�P>5�,��TJ@�n쬘�%n9D��jq�ѳf�,a��+��N>���I,D��c�m�*!05 bd�}��� 5) D�x�E�;u7*b4m��a�̥��F9D�� Wǖ>�Zh�S-��3
�W�4D�p�ҡ�j���2K�e��]��<D���!�|@��#I�����j6D��30�L,_��M�0���"�z�� b5D��,Ԁ��	Q�}B�(��1D�tT+̛g��i;�
�7�h8Yԅ=D����N��VY1��/e���r`<D�$���ɿ c
�!�X:�j��!�:D��K�Q/u����9B��'5D�4��f��g�=5����i2D��#�kI�F��\�ʋ�A�n�rE�3D��K"�Ǎ'<��0�"�wj�QUl&D����ǎ�(>Y:��T�:1x�%D�p;ĢM�'� ���Ɵ���C�B#D�l0�F�(�,���Q/��""�&D���D{O�O�,�,��赪	�'.������/=+���E�-$���	�'Ö�JS�F�S9tY����8$X��'xfq�,��.$Rש?|��l��'T^ �g�;lcR�bF�%_T��'�҉��;�"�v�Z�!�L��'ɬ��b΍,�D�s��6
�p�8�'= ��wE�D�\�����}�d������,�ZI�'��H���p��k�!�䉎pB�Lyg�6T~h!��(J�n�!�G�*�
s��Xcd�hC�m�!���.P ���@�<1�PQ�HI	`F!�d��O�FT�\�w�8��'>B!���J(uzg��c���2A���#!�$[%[��A�t\�8U����!��,ZD����M�sz�(�I�_�!�[���q��U��D#U�ƣCl!���-)�*� . "�rű`��a!�$�S4lҁ�J���9�+��N�!��t P�*G�z�2c�D�W�!򄕝<�V�iu J�
�&yb��t!��L;i*�I�4O�8x�{எ�eu!�dL4j����N�H�K�5�!�A ����Ú2�
Da�I!Q�!�$D{T�۱�?V�hI���ȬA!�$ֈ9�J�󄭄<(p�ͳ�Y�8!�Ĕ�Z�
L�Fo�)cY�w31C!�IQKRh��D=H�(���&S0!�DP�X���sI�C��p���"r!�d	�;�(v
�\�F���(��A�!�D��]BTI��^&&z�#��F!p!�Q1U)��{R���,�	H2h�5n!���"R5��W�
� ȸ�� ^N!�� �TX �F�cb h�3i:-��4a'"OjA!f�8K�rq���IW�~��"O҉s`����\x H/'Ҕ�(�"O�|�ř7��B�z|�"O�1;�J����g�4�x�y�"O	��̍ ���{mH���"O<�xc �c�p�X�Jݢwp���"O��4�M4�pE;4�B!6���B%"O^��k_ XU��(��S��"O��tV#xT��ˣȕ�f0.���"O��	�b��[�����s� ���"O*�A�b�6�̍��D�;2r
}-�y���G�01�\�D��9o4�y��$�V�۵�G�U���p�\��yRH��0z(c_?Z*L��'fR�y��E�1`�Lڃ��!�
L���Z)�y�a0D2�E�$�,s��1�
�6��=�yR�2R�~����2��$8�mX9�yR�jI:��d���_�.$�aiΨ��:�O����EM0�`Lq��L
9@8H8D"O����h�0%� J�s/����"ObE+��nG<��W��qL^�"O��IWfZ�LE�%j۱t�� �"O�(
�
Q�ab6!z�K�(C��m���D�O������R"[�a�p������L{�Y��"O�|:�V�8!e�`�$SB�p�'���k�	�ct�Q���"�¬J�';2�	��MM�@$�x��{�<��
3!�p�!��r��cJ�p�<�i�*9�NA9c�E9Μ�'��e�<i��u��0H@�=J�g�c�<)�A�q
���!�Z��F�w�<Q4+[O�2	�D��?}�j@��X�<�Ӏ[�Xl��@�߹`���׉T�<����@jt��fՀ3�贀g�Q�<yT�LsƬx ɽ{pxp(姑b�<��9�x���)I:k��X�m�b�<���@�-C^q
���:�v��_^y��'�h�@�%H�P���j\�D��Q��'U,�a2E�A�Z�蒋��}�U��x�j�hf�$i�C�"%��d1����y�I�";p`1��\�	$d�@���y�l�"�Q"ADސK
=S�NJ��y2,�r�ʨZ�K�q�Ti@��y򁇭`,`�kq S�n���+��Y�y"�\�H����T�y��A1ևM'��>��O�=�RgF ��f�6	�T�"O��Y�ᖕ*+��i�k�=�h1�C"O�*���=�<�W��U����"O�2�"]8� k��^mF���"O�� �'����R�HUSN��"O���)	�j[��@M!����a�'�ў"~�dA�'��a؆�:
�H�$�ѳ��?��'�p�y�%�U����eG4G���C
�'�.`�#	�u�t3u�3*��	�'M��2@�K�&'%z��U$�H�<1��ɸK�ĵ ��̡�J"q!�A�<��N~ڼ��n����y�`*{�<�2㞥Bn\Y���_��Lbcw�<YìX����5ř� "r&Uu�<�P��sE0�! � 8�� �!�DN�@ܶ)�T^0m:�:�	�$%!� �H�����_�����Ǻ.)ў��	7|��3�ȵ���#ω�&C�)� �ɉ��l�Ȥǃ-<�<�0r"O���JG�)�Q`� ^ώ�h���{�O��0k ��͘���f
�Zz�ȳ�'y"@��O�kF)(un��z���'��t�W�[Ø��E��&F�t@
�'3h-`֍�[ {u��)%h��R	�'��m	���+c��eK�-�Q����'�Ip-����4��_V:���'e �0n�
ij�l�Ā�Rk.��'���!m�p��቏
PF�y��'0J�B䚛8����Ŕ����)O����ՠH�kקV�oD���r3!�DEj$��`���]�5�Ȭu�!�$��8�pI貅��M'hQK��H�*�!��	(��ܪ��6`|�:�
�2$�!�
=��)����.;`XÀIY�q(!�$QuF�)���L3.X�U"	�<!�D�8V�q`��US}3�j��*qў����<�F1U��u�\C�?_ZxB��e0�hP��6` ��;d��,L.C�	#Y��0%�LCR�*E��pC C�	w:B��)Ț<��(��$�B�I--��A!č�1Ԝ�4l��k�\��!ړ�?9���$���A���4wF �׽pq脹�'����b� ��EJu�hH.�ʏ�$/�o� P0'���
�n��f�1#��� �ژ0�g*X�vL�K-Wc�E�ȓ~�8�&&d~��DBG;���S�D�:A��5+��}١�ۉ���ȓb�ƥ9f�K� ����)�/c��ED"P���|:e��@P�2��d�t����<y�c�T챡���L�:y��`���hO�'�8��wb�����h�%�a��$a�+���(D��n'�Ն�b��K��  X ��T�p��s4:H&C�' W|�Yw!�Ah�܇ȓ<�\��'ሖ;@����4^�F2�'4��)B]�j��C(^Fm���	^j!�Q!#pܠ#�j6A�&p�#!���T��&��gܓ(1�|�U�M�5�\Yw�[9��m��C�(�d�'}v�A�&�qm�8��)Ĉ�`�֭m���E�LgЅ��B�p�X%��2Ȇm*��U�w�v����z4ˑ ^)d)�3�E����ȓoq�P[���Y�t(z�J
�H��a��k`��-@�\1:T�Ո42�?���0<!ao��r��Ї�R�f�,�����l�<1-� _<�)ۆ�ޖK�싒.�k�<d��^�<|ȵ�L�F�`�� 'Cn�<��_^�В�	�%s��a��f�<�͋��z��+����_l�IP���O������Ӳ?հ�#�!��l!�/O��d�+f`X���A�Z$X(��C,=�ў܇ችE�T����
�x�D�J�8��C�	�!����E��-n�0#�!�kR�C�I�J��Y꓆tMV�r��z�\C䉩1)L����
� (9���?�JC�ɏhW�h+�ɂ�\���P�[�c|
B��;mb��S5([�"�9"�Û�u��F{J?�(�̆u�,1bmst��b�;D�H�@j��oq�{cBƓXˠ)�d
8D�ls��4g��aq �;�l]��i#D��r��Jly gd�W�F�j"/"D��`Ղ�)�Iz�,U�ݩF�;D�� hPS&K��(�zV��=Y�h��"O�!BH=��1׮�\q*�"O �b� � &��J�`U=Z�2"O=!uk�ł��i~���O@�cޘ_��a ����B-�CC0D���h��b@����[��<�JQ4D�D��'�oC�RD�6Wj]��N<D����gG�/��0�3l�5�@���=4�(q���!0b����++�i���\x��Ex��	�G)�ƤԪw 0�`�F���?	�����RA0	
$C�n�d��
�,�?	���E�v)ZS�I�f9s'GH%9��`��'��e.�<3>J��ϟ7�	�ȓ9V8�@[@NZ���Q�xj�܆�D�i�� �w�>\ӆ�M1���ȓR#�5��A&x
4%s1�=g0���?�ӓ&K�.�L��e�?�Pi˔�=|Ob����j�(��(	v|���>D��I2���i�bP����eV���F�O8B��Y�XA��.gL�p�$�>SDC�>yL��׻q�(��ט�6C�ɝSE�̛Ѧ�%�D(�Qĉ)(kDC�I�n��Y�3
ݭw�ܨ�Ì�K��C䉞L�~h�bO
�2�c`J }<��?���)Ο5��l�c��:�~HPU� .��'��	y>�"�
]�����4 \�3����$":D���&��&jњA�1�Y u %-2D�h#s"ܔ,��<ȗ ي*����a<D�@ &♤2E�u�&󐁘2g:D��1�W�L�����L Mv��Ɗ�O���G{�O�1�B�y���P�cN�^����!�2B�OύAx�)F`Q�T�@��1�p�'��O�hp���W��UPC��0B�4D��HSÓ�,7��ĥs.틠C%D��*�)�[�
���(cr0qpg"D�@��iP
h��s�b�`� ��K 4��K�bU(N��HՁͰ�(�xg�|�'�a��o�>w�9�#Ɇ'��}1����<a�����-�j%I�$�
6(�`f�$!�d��9�����c�s3� 8�E�Na!�>O�̙�`o�g8�UFH�(K!�DØ�x`���@/}	�p3�,t�!�d��.�ޭ����'�,�N�>;�!�۫�p@�tˁ�7����ӌB�m{!�P�_���$��-wh�
u��d�'fў�<��%H���(�p[�5���~�<A«Y�d'N�)���$/"lĻQi{�<�"��7UlP��ܜu����y�<�6�0s�������J$a �v�<�� �\�*H�`�˯z_Z�P�t�<���Йd���#��--)8��Pb�q�<9q�^�}��H2�H�
��TpS��d��hO�',Y���f�:B̉R1�{�M�'�B��SA�Ta ��W:/�D���*�
C�	9-�U��	}�L�"�,�`C䉹x74X
���K���EHϦ5S�B�I�!�Ft:�'�q��H`V��-���#j�Fp�f�8�ea��6fP���#�dх�о>[���r�4%�b��ȓ�ƀ#q/Q�䡨$�,6,��?9���~:���"ސ\3�dךR��`�T�h�<�e`�a�^5��K��&��)�SO�z�<A�K��O�jw�/e��ɂ�@|�<1�<A���k�ό�E20�e.u�<� �$ �o���.��ïX� ���:B"O����b��IX���12{����"O��s@<�a3#�ˈ;�� �"O�X��F��B#du������"O(�{�H�_xl��V�L�S���r6"O���NڠX.�a膀S aQ3"Ol��D�(Z�츓3Q=Y(���"O �6B<�Trࡑ	I�´��"O&���/Z.���A��"���R�'��O8���%��D�T4j�KX/K��}��C��y�o�J4p�l�#L�0�0����y2����؂��={p�[�	���y�& X�*e��ɀ3�p�Ɇ
L�y�.�"N����Wʝ *G� �v�	�yr���S��Ik��� e��&�2��<��䝱�2ܱCm�).в���5)rў���I:!�+'��#Fv����� b0B�I�_hB�`�D/(�@�� 
4C�� L��D��$��8"���>��C��?T�X#��O_~�����Fg�C�	���p�E��Dr�`I�/��C�	d���% Rj�pt��\�rq�B��P$y��-T�Y2(�"kv4C��\�iY�H��w�$r�L�XB�I%i��Ä�լ)�,I��C��RgB�4^Q�	��35���чW!K`NB�ɝ^dZP�J�=�����hT�B�� +r8�D3%a�A*q�C��93��� �������C�~�B�	�h#���@Z�L~lQ���G��B�I���S���1/F	C2K���B�?,nd�yg@�j�<�r���5MA�C��e��԰E&�BTr�h�a~�C�I�-��ug���yB��u��TC�	e��t�A,J��2B� ��B��m<��B��"6�p��X�m.�B�-gqx@�t�9HP��-A�	k�C�	�O>-����-:Op�c�đ6C�I�'�(Uh��[+bh��k���>1OC�I�Sd�*�S�LPbQ���x��B�l�|`��M.r���R,�B�ɇ#qDl���?�
����f��C�	(~w���dB�`@�����)��C���h�#H<9x��%��>`�C�ɝE;��aE��#f�V�H�jΡ�d��T��uʡ�Y�GQ�D!m�-W!�$��D��%�F#<"���ޠL�!���@N�yb'��DHj�Y �Z([�!�d>Q4�)YblɄ��I���!� ?V����\�[���H�JD!�dO�X�HB�Bۄ+���p�-�+-�!���\G���ݧD�x���>0�!���G���K�%��(�*�1A�!�d[V$6�9
��G�t�[�mp!�$ǐ3uJ�S�̒5
㚴��ӢN2!�d׏	��e�T����-����A%!�D�bJ9����\yT�� ��7)"!�d�s�q�&��tb�U�#�0g!���nG.-yF�ڱ3�(�*���|M!�$W ������M��r��Ғ3!�=>-N勁$�x��Ty�o=�!�ͱZY�#�Q8:�0p:ά	!�$�)\�Q*��7O���T�� p�!��G�0����a�ߕd�p�tŵ�!�� ���!��ڪ�Z0�I�3��(�"O���Js���Ĝ)j�t���"O�eT�$B�p)�e#�VBT�!"O~�)� S����aM�f�Z�h�"O��금&��,n��S�ÑK!�)����-W^��9�G�,o�!�Ē�v�N�Z�F��=I����._�!�$"	�t����]�T.L����[$0>!�+N���\�-�,�1�K,�!��+�)S�	2d�Lä�H�Q�!�B�v@�2'�ŦVBa�3��9�!�DB� ��]"���\HN�S���=!�D��r��A�}B��ro\8~Q!�D��xȍ*�LN4N��'O��!�DP!AؐU7�҇\:x�yÃ���!��H3���u��o2��2��ȃG�!��"뎄o��PB* p�	ڞ	��B��	pZx�:���&�$���05R�C�	�m�LY��Z={ۤ�`&!|zC�I�4�02Wo�('hua�
Q���B�	R����Jp�8��OV��B��-b�L�c�x��k��S:B�*c����_M:��ac~�"B�I���	r! e���@ЍV#@��C�ɴUN
x�uG�n9�1�P	V,j��C��5b1�$���ؠ"��� ��.l�B�I�<��MN�X����bC�I���X�E�EW|��W �'x(C�Ia�Z��RB�h�\�QGb� �8C�I/<
6Yz6&��w#@d�T�<O$�C䉓[�ҝ��X\s�����-jy�C䉼q�v���nS	 �Ơ ��	r¦C�ɸW��Lص�B �p�+�/�2)�hC�I�Q��5��MD�&p�S��̌s&XC�	�t��y	�)��q�vd�T�T�mdjB�	6}��I(Z�/h�� �a#;�C䉫q_��A��0%%���s�Do7�B��M�D��$M2HԾa�g�yHXB�	�)2M�WO�}l	S"�~�NB�'rV�	���5RPa��Z@B�I�m�:o�"`�6�;���`KB�Ie|t�K[�-O����H��"��C䉙r<t��R"�1C�-D��I��C�Ic�Ta����r��O�5�C��!�Z�+�q<�jt�٧"6�C�ɱC:���b��6�X`t���C�ɉB��5
Wć7RV]pv�|�q�"O�0� ��X��xe�˱Tp-`�"OȀ�&�I:za�l@�ܣjp���"O�}	��@��4-@�J�Aaʹs�"O�䊷�P�\#.Y"uh��+�lD��"Ov��uOE�u+��g'H-���j�"O�<�Ћ�p��9�抽[Ffi�"O���ď F��7/(=����"O����֙w�f(���N9{��)�e"O����'[&+��mRDĂ
� 0��"O�X�`J"�*�;���&�Y1"OD"�"�76hЉ�G�+�"psQ"O�H3�Žr_(�!7HB1J�Ρ�!"O���#��Q�\���l��3"O
� DƼBWd5�'�1H��Ȓ�"Of�ٷ�G�7�6�^�y�Ç�!����H��<#��d;���A	!�Dۆ";�}+������r���J�!�� z����&g��L��S81��Ӂ"ODI�W�%o�ZW �?i����&"Ormˣ�� ƬX� ԛmX��&"O�-�eÐ&_>:�$bw�X�`"O��S�iĚk:챓�-�"O�eC��2V��VB��U(�H�"O���� Ц/9^Q��1oJ�4cW"OP�Z!a��B���`M_���\�"O���5��y ���(bv\�3�"O<�*�Iߊr*<�z��G�|RXt"�"O� �£�ay��B�G�E�u3R"OByc�Nޒ ��5�pi�`�,4��"O��	�(G�D��h��"l�<��"OpQ@g�A>a] �摣hF5�"O�@��AL�v= �҄D3mT@H�"O.|� ��'7�쒦BOk8���"O�	��J8&��A��)$�HS%"OȀ�4&V0c�)Y` G��p"O��ǂ�9r1a���#C�	�"O��� V$\nn͸���G�\��"OҤ�dU.��a�
�D$Q�"O�l��&�I�}B�%T�x�d8��"OP�N4.�T�v�V2Ըғ"OL�Yt�S�C
�)#�g%)i*"O �uj�:/���)cg�^�$cp"Ol9r�D�"�h��VA@x�f"O�Pڂ��
L��#��l �"O����#�V��x�Pk߈Z�5"�"O�� �:-5�����Whv9p�"O��WJ��J�2�ަ"�F���f�<��ĝ>�P೎O<^*^�i�<YVm�&�b����$��]A�G�d�<!T 6l�h�$Ɏ#C�U���Y�<)A�;,���+ۊw�p,)5�G{�<Y�.7F��y�k��p�+�~�<q�J��1�R�;�Ȏ�b�������p�<�G)��yh ��S�Y+9uJMP�RS�<��)R�53ṡ&2t���B�Q�<y3,UJ�~)
��O�)�����^K�<I���E��U���������bD�<9����"\\�S��#O�=�� E�<�%�-��A�` E�t1s(WH�<ᐈ^*0��Y�lZ@�tyb��@�<�Bܘ8�[0-����-Ik�|�<��+_?/�Le 5h˫iBn�BAq�<aa�
t�z���U�|1�6͗S�<iDEX���AQ�iA"�t�ȖK�<�WK+\���P��������A�<1S/Q%�Ph�.�:L5�!��|�<9���K4X�c�O�V��mX4��y��`����?��t�	1,�=D�8Y N�R(1�d%I�E�8���<D�Tz&�U�JV���;y���&�=D�@!#�B�:~¹Q��0Z���c=D��R�o
�ik��@1�^M?� S��(D��
c+�-��K
M���D(D����BC�K:���gϝ:%�b|:sk%D�i/.J�����&�3�'�W���'r�J̓��ċ/y �b��	}�����`vLhIN2i�n��dC+P⬄ȓ M��*��ף��q�a�=�r���P�[r�Y /��DJ�@���I����V���IJ'L�D��� ��YsZX�����!�$@�p�C�E8B$�afہa��6�id�"~n:� f�A�0�ٹ�/ŕR� �"O�4Z�,H)j�b4{@O�d�ޱP�"Oā�w��?xi�q7 ��xۈm�d"O����k��t��d�=iɦ��`"O�d�GE�Ng.H�'�X�5䤸��"O�h�ͣw�Mq��=F�N�Z3�'z�ͦO:������8����.ň qs"O<�	�BK�.r\�䏽/D!a�"O>���DM�o|8Q� a�[���B�$0|O2��w�]�2`��D�`t"OڜJM�u�X�'ʸҷ"Oܐ;�eץcR }	>Ha �"O�
�j��>�̐ٱʘ������"O�`�!�5@��Չˌ�̹`w"O�)0E,�7-F��!6H�3( t"O �(�(4��HN�\���"O^ABS�\�w�yap
� s�Y��"O�}�f%Wy״�!���:.�Ya"O�m�V$Z��,�7�,&Ѩ�"O�Q����#30��ڢK%Qh��"O^�q�V�p��H&BFh:c"O`��3�P��4��sf��(���"O�RM�"j���;c%вh���{�"O�@�<;�}H!*M6)�VdB�"Oy��Ly:���/�>�68�U*Onԩc흘0[�q� ��3~���'5�p��E�^�6tc�.L�p�x[
�'4�pk�������SY�G� ���<E��@n�Q���K�<-b���*�&)���y�P�*E�M�+���+���#'#h��V�(h�6e�6fX��8���%�2P�'�ў�|�7��@�L�x�5� ����|�<��N�4 �"%�}�����x�<��2�6Lbu�~�n���`Mi�<�&ElN�=���ѣ�\{���I?y��::H軂����
�Q�h�E��	��=�'e����h
]����&ΣE����%?D�Td'��Bِ��$5��U�U�>�Ic��ħ�T<HeNN�E�8��;�.��ȓ��`+C2abʨi��4@*P�G|��!�^�8taS"p��J���rdB�I�:F���B�^st���@����'���\���'SF��4?��u!�� vnV]��4��}�T?��'��(:����DF�v8B��S&[�Eh����p?)�?*^e�� �9o���a%TFX�ܥO�zFfʞ1z� `�ۘk[ڝ�"O0��G(b�f��`!ɸ3HF��v"Ov�� Hݍ.4�J  �j�J�c"OlT�u��dۀ�@_��d��'��IV��hOl�馪�]z�8YM��=����'�1O"���B|P�m�~��@S�d5|O���FZ�2�DB�*����{��	m�O���S�i�,G%C�oZK(1
�'5��p�N��N��܋q�9pF�r�4�����x�"9o�Z�S��D���С��԰?�H�@}�!���l�@B�+%���X�����b����:�`QG�9t�PC�ɝve�傡HQ�I�b)�@-��Q
C�I$[���� AΜ?x�#/ c��j������!Z��H#4b�,*k蠨��yr�
�']���!)�12G�ep����(O���=H��ଛ�0It�+� �`��z����	�j��v �		. ��Ro�>�!���6��5����#(����fN�nca{�]��է� �P9�.�?��`;�
YKǠH`"O��;�`¸�p|�� ߮����&�S�� `����cɎ��"�����()bB�	�~�b�s�+�6ݺ̨�`W3�C�	�K�ބ����&_�옂qI=�^��$�<���W��v�X P� dZ6iCq�'�a���Ϲ�B<#�G %y^�Pi��ԈO��D�4c �d����焻H����@B�>�yBg�'8d�;�Qr�l�������7�S�O{P�q�<_Uh�0V�F�k��1	�'b�8�d�L�BSJ�ҐCCd�r��H>A
�I%��[sko�"�8��D�,��!�ȓ>ot
Aú2�x���',���>�����Ā��(!3��_���<SAEF3�y"'�yJ��j�Sr^@9r�H��y�K�0m�� �U�L����Ղ�y��`��[D��x� �`6�(�yҤ%p��H1f�t �L�y��D�:���v,�-u�gMW��y�혳~�֜i����q[�G3��'��Il�O��1�eH�m+@A��	W�J|8�'
2��G�S�O'��KI�lg24i �XL\���'�$�c�$����;<���+O"��ā<V~,�bǭGY:��VMa�;\OV��'Cع��MZ��M9w%D8�H4y�"O�q�Oo�)����	��a[�O�C�eP�h�p�C���l��uq��n�<!`�ĉEV*T�7�ʇB��Yq`��m~��i$�O֢|J3.�r���{&�މ_t1��T�<�B!Y�v�(�]��e1�'�L��oӺ#<���Cά@C t1���6π����L�<)�1Y���ɉ������ɦ�&�d�	ӓHy*����@��#�3<8�Ɠ.�jر�'V�TQ���#҃z�<�2 �*$�� ��ըG��X��o̪d1��(��2ғ�hO��2rP�c��`� ��\+@B�(@<�\� ��/K�N�ru/�_�B�u�@����:�#S$Y��C�I!44I
�h�78��摠l��C�	�}K4�2�°r&��I�DC�ɬ^����Ʌ2�ĺEd[�R�0]'�Ȅ�I�&���iUK�+Lt�rr�X<6PC�	����N̵4uTKdm[�g<Z��F�,D�x P"��&:� 灘�@���$(+ʓ�y�ٺK�_? ؼ��aP�s ���L~�<�U%�vq�`P��=7��|[�d�{}r�)�'l�tA�a�֙]-��k�/LaU�<�ȓ��T��F�(m��+*�8� �?!�7��ؠNH��@SQd�D�-�Ɠ'�"�� 8Y����g��75B[�'��i9q`�\�6����%Y�F��'��m�:�:!�CJ(_j��
�'��Dӆ��&��ͫ�ؐKڽ�	�'���� �A<=���: �5A�d�Q	�'t0��$N}�$��J#A���� ���A(�`�0�0C � |�� �ȓu$Wɇ2afA�@�C�=�"!�ȓP~������"�Q��]�?�.A��8|L�%Q�d,��D����m�ȓ~�n���]f֑�c�:'�ę��i���H� �<�~��O8f�V8�ȓK5nP�u�S�xN|�f �	#O�X�ȓ�^���� m>Ehq$�uujɇȓr�[�
�71�d�"�*PB���S�? v�;�mі1C��A�oE�Z� �"Of!��"�	r_N$rn�&f�DM(f"Of�0s#�)xH��T
�)66�}��"O�m��&ޛBZ*�Y�(Ys�4	�$"ODm��f�։	�i���)�yR� A*@�Kڤ�HC'���y�cZ�]�!���ˈ	=F���h�=�y2�P�|KL� �X1o��s�!T��y��/>�6 P��R�4%�ِa�%�y��A7�"�*�n~�W�(��H	�'Ab�@��_�l�2���9��h�'?8� V� m�.��6֋:���'`���皶�F+ߣxp|��'0
yx`�H�<)��E:o�@��'��ԘR)O�uX�"�+S2�ȋ�'��i	�����,GB5z�'/��0�LUtz�2�eH�>��'S�l:���9v�<��éb� ��'��$3�J���>��㟆TɖYj�'���`�(��O�\�r F���Y�'���p�L=5R����F�A3��ӓ._R�q�C#��ԁ��v�T\0��̜~�
�J��\�D��u��:���"��h��Ҷ�L��ȓ"^��`!�G�h����&ʭH���ȓp���K;H-�с����s��a��6���k+��3�Ƭ1p	�'��t�ȓ9� 0Z �W/�쌻cg�4}���ȓuR�� �zG�1Yb��/f"�ن�B�t)�dDhDE[�R�D��C>^�S�Gs� 	x�%W�	x��ȓS�^M(`*�;9�<`#�Z�%i<��T!F�2S�ߨ%��k���[紅�ȓ��ɐ(È.�Z1J����P�5�����C��f��y��>*�z��ȓ.\��fם����V�m�h}�ȓW\X�1��5~,���2.����J�֕�A����"���2;�L��w�
Ii�n�E�
�ɑ.Z^V���B��+]>9J�92�)8j���P�r�R)L�M=^Y�B*	�pv��ȓv�P��@iƏW}n0P����L��Y�$�TM� ��KN,8�\�ȓ]��LƇ�B��`��*�3m�T���N�b��ʹY 'K��4H�ȓ~�(̳��(i\�����^�3�6x�ȓ8��I�s�˹J��I�hCռi��cP�=KdB �)F�䐷�Ҥ/�ɇȓL̎� č�g^1�G�	�'q�9�ȓX	�|�!�!�<h��Чk�l��,t��C*W,9`H�Yh��ȓ#�����)�a�R�#8����Og<�SB�W�����^i�t��/�yK�Ē�ٔX��#��#D�h30�\Bzʈ��
O�Y����s!D�����F dc�a���B����L(D�X�Sg4W� 0�/�;g��Jc%D�D��K�<P���@e��'b���a�#D�����ؔ==|�&,�kHTs4�?D�<����<C��r�"1`�[��!D�$5��Y4$(��։w8$�0D�g��'H:��E����)�q�0D�L���5������ƴ�+�.D�Ի��\0����Qo�� 5��:1,+D�X�egNM��,R1#P%\~d�`�m=D�� T-��.�3FT��s�H�ԡ�"O�4�&��K� �Q'cWS���ۢ"O,�1 Pl����BmD
���E"Ox�Z���Yd8@gN��tJ�"Ol-i�B�.
(�>�8U""O����M�5]gą)�D-�Bq@�"O�-��KH�B)(�#�^{<�B"O����*C�l�V�	Y"4�1�"O��·��.l� �yƀ�Ɖz"O.U�7垚fV�� mS
�!e"O���UeQ�N�D��[��
"OpM��F �b�xjqL�?b�>Yc"O��6d�(><����l�p���"O�%�LZ�G��Q��F*N-�6�0D�DkR�ަ9w2����4>���V�*D���㨏 ���z�㜹 F�P�PD?D���+�>M�40�p㖢i�(P��=D�Dh�ͶxӞ��!��k�P�Rh9D��U?X�<�y֣
�>�"�0D��kR�?(��C��T	���q)/D�{�F�Ge��agP�Y�I�ԃ(D�Tʧ��2d�����#Lј��2@)D�s�#[4@�Z!ꑉF�V�2Ŧ'D�� 4 �Is��!���UT���]�!�DɷR� q5���!"�`�|!��\�9�8=⁩�2�ܡ`wlO�Ql!�$�7������A�N��U�-A&-�!��4\�\�sÓ�M���	�,Q	i�!�d��mid�HbJa� K�5�!��W���A��[^�hh8(��w�!���$LPF�d��m�t۴��*#�!�g�Hᓠ��<n���3(�!��LHRt��R
��v��@�j1!�$V1u�(� ��3|�Z����!�Ĕ�mcH��҈�1��Aˣ/M�!��ݣe�2P�Oف%2���O	:)!�D�1�@��L�p�t��"
u!򄁰P�PbsG�M��<
��I�#�!�$٩d�.��)�<��<SC�/T�!�dԇ;:���KU����X=y�!�dG�!�D�
5[���r��,�!�R�<��	�#D�OD`���q!�䂕ed<����մ\B$h�Lњ*,\QV���p?�B-�}C$q�)68n���#BX�L"�D��ms�`Q��j�-Rb��!���X	K?ޔ"��!D�0���10Zv�(�����: >?1Ah1�		4J�<gז�~�*�<X�Q0_������x�<a�n��;���8�	&vQ��Iw	
�4�l9�3h�ȟdr'şv��'?㞘�$�P�Q�&�9��G\��y�d3�O4��d"i��1��\�K���0���J�q��P�����j*�OX���CI(aۚ ��ŧVD�
��	�IJ�l�y&.�rb�������wuX���D��� ��C&�y�h�00�K�N&v塰�����AmX^hr!k��xeP��U�ȴ�h��]�C-4m�r�Q�@<�v���"O��7��A��t���!��0!��~+&�9d�I� h�)�K��g"�'��'��u�&� m�691A���I�|�������{V��wNL�����T���8��\s#��#'$��OS8hx��=��$
�lA*� e��9i%����W�'O��f���WZD��S�� XΠm������a1cU�R��$���Z74�lJ�"O�12�(_�#�H�)B��E�|�0��Opy�Mg_~�KF��q�7ҧm��Y���
	��(t@�~�4���!�*�23'W%=x�RfΚ+{Q��{"�)7tx5H��W�gἑ���}��'������1eM��(�Lu	�"N�47����o�R`2�٘)����@]:AmIj�J��o)���P�	�>ر3��0lO� �����ͦ/��j��.+K�p��I�+��t�p�
(c���2�I�����;P��s���%�x�i��
|�� ��}��k��Tlm���Q�S�͒��'��pC��MN�>� d?Y��F��T�>��Cf��\�90M��y��� ��TrR��N�-Q��16�11p�%&t�%y�ě� QK|�>1��ޯ`3�j��@�GX�`ik�I���(�+��J@�ISF��^�\�ՎڵG_hL���T7c(}y�E�E����"�16��3o��uS!�H�ԈBƌ=3A@�K�e̹��d�G�~��0�/�|�@
'�y��.BFȌY��4�<���Y���W�#`hQ��2!_z�ʍ�ɒ�p��5P!CDyƌ�й=$!�d�:=px��3.&%
�E�i*����#'?A4��%�Z�>�O
�$�� dd=B関<�-�f
OvP"0�0吭X�5�@Q���q[��Q��ً�0?�5 N5�0��H�Ȥ��v8�|�l�A74�
�b�S��ѡu��U���Y!�W`O:V�!�ă�}s�q0d�1@�1ZeE�]_���b�.<D�Kq��l��/s�O���!�ƽwRƱ�@G�/ܸ�
�'����o8K.�H��"�$j,�-L}�H����.,�PJF���g����(�  /R(@����xj���<��LJyh�">����>>�9C����1�i�Z�գ�Á�	�4�_��$@qC�'?l�v��4c8^\q2$�x=�1p4�[D\#���P�<��d�x����W���.׎o����f	5"" �萝Z���x�H�5L� ���, ��h�)�
z���ϒ3���E&3 ��K�H��@�����H�2\��FI%Eƌ����
E��cU� ,�z/(LR��PBD�ؘ/�1�*��DL;�N�U�CD^&	�?t@܄�KT>Z�0�$哓kG�ϸ'����(�t�2����*�,�Y���U�X�m���B�`+�)�0�e�ݴ,��X�FQ��졧fM3`���N�i[z�!��`�36�/O�X�r�Ϫ^1䔀#mS�I��ܗ+ƂԚ����d��j�@	vV�uB���IM�,b>}(s��`"��qn@IN��B%� �r�,sQ�s��ƼS�
6��5��� }���(����@�q�}�rp 􏒴b���j>�G��I t��p A*`>�!p����݁ F)��D���D]�>�,(0�؎��'�-���o�+c�˽|�.�p�\�+�N���c_��TI8�3�$�4���"�] P�19��F����8���PΈ�}4xN|
uA�p�b��'=.X�g-H�B箐7 F	o����
��,?&L��*WsƄ3v��s Πٵ�&Фz-O� #�֥J�tP��d'>fp�"V(p���Zf��n&ax"�˦�F��'$91B��w�ҥ84d@,K��I��
��\j�;��J؟�#7�+o�-��!̬I^:I�2'!�.��!�Ƅ�2�$�&�tG�6kW ��˗R���"O�
Hܣ[L$�io��8E��Y�8��ؾb �4�>E���[69��" _r�N@�'�C��yrK��V�%k�v�RJ�<���'��rT)�ϸ'p~0)ǂ�`�,�+���Y���
��*upI�+f�6u� h�kD�ā���Z�*#�O~��S�п
�\�bc��8��1xe�ɹA�>@B��Kw0�O��uB$%�`6� z$��X�xh�'w��@3��#�:�s���<_���,O���T�P #�pirL��|�V��=�ĸd�^�ܰ�P_�<DNg�۱�Z��N��A�԰@��\5,�P�c�(��g�(o@11a:yy�!���
�E���(mTqƧ3j�A�������D�ey�8��9�T�I��ȍ\R���DE��F]��	#5v5X��$O�\�qPC�T� ��(U�Pq!�$?2���(��֧K������!h�!�+G��d)$
�$)����A�y�!��ʬi(4�xf��*��BU!�䆘��	��K_��T`��`}!��ؽX� [�&ߒpy���G�i!�d@�<�b�*�Jogx�X ��8+o!򤃇�,��#��1�윹�g�?^A!�׻d���tEL�H���ʆ��6!�xD�����w�<C&

�.!�$C�0A��	7e���sIN�'l!�� ��0��I9�H�!����C"O�,�a�ݰ`nr��"�:�l��$"O��6�H2b�мb�N��V�"O@�
2��5�yi�� �G�R��""O�4��AJ$�|�*'�_*A���"O��@�_<P58�1���39��ĸ�"Oޭ�n�f�������	���s�"O�ܳ6�dW�A�1�
�x~)y�"O�r��yb�r�XCr���"Ob�y�m_�B���f-��b�`�T"O��ǯӿ;�7.�4�4��"O��iA쏅e�b�ᶭ�"O���nG�Z���I�F>Gy؄"O��(	��* ��ˎ)���y�"O���)K#5�(���t���Au"O8)�V��Q�lt94���^���s"O ����V�`�`ܰ����9�,�q�"O�T�&�4ZI�a�@٭��a��"OJ��A	�5��D Y8z�ã"O�(1��׉��@���=��a"O���6���l3�URR��k<�(�"O��:�I�!]nHtj5�� BZ�b5"OZ�#���٪�+r�	 #6�CV"O��(�@��ŀɕyԄaG"O��+g��`��9�_<���"O��F�j�z�xD'V#7��ي "O��C�;(Ez�f��
�,)�f"O�|X���A��9�eN����"O-I�Ô�1z��������xPT"O^ �p	+R�yJ1��?�Z���"O���0��	V�@})Х�!�d��E"Od���ư�a�Ä&5b(�"O��I�I
0����&"H0b�����"O4��2l�-��i�cB�'� �e"O
�3���*4���-7�J��"O­h�N]'H1�5��޲��mkc"O.-����khe�Ag��C	1"O:u�� �A���(.2dS%"OJԂ%��zN����B		�(��c"O≐e��:�j��&DY�T'�Ta�"O����NW���D�5>�LQ �"O`�a�/�%n*-�@�u�FA�"Odz3�N�MI7�W91�:�sP"O��p�V`r&e�1b�#R��h3�"On����aᲙ�!�����2�"O6�iQ懞O����/F-���"Oĝ�d+)wP��B�'!���"O��J�͚eR�h�I�5Tv��:�"O<ȸ1���Ran��r�(8@"O�hz � Z�����5<V�2�"O��	w!�b��rp�8���H0"O̍�@ wgD��%'�U91�P"Ob��6�W�`�'Q� %�"O̤�ԦJ4Pa�XIR�_k>\���"O Q9Ǝìs��3�%�`pn�"O�3c��1����m	�F�H�d"O�Q2�m�>Z���QG��o�;�"O���bÑ6<f����K��(��t*O@l���G�wW��5bW�I����'?�(� 	�wD`�;���~�pJ
�'��(Rn@ytpL;u�X�m�FxH
�'�
�i֦���P�)�@t�X���'�(�+s(CJ��x8�b�n�����'��ea��'}�|
%@S�b����� �(�L�j�H$)�
��0�H�X"O"|�CgO1.�}B!������#"OVt���9lj&Q2�bV�$�N��"O$�U�P�"L��da��4���@�"O�p�uM��c{(�Q�� �~< 2"ON�
��������� ��3"O
D���	?h��ײѡ�"O@�U%�l�!��]�_���"Ohl[��\=a�f�(s�	t���ҷ"O� `#�W"Mɶ���J��>̪��@"O����-±�j�cZ�}L� "O~<��Y�-� ��wo[�C<�"O�0�ɓ:y�	藮�CN�"On�@7e"bZ��1	�U�ɰ"O���W�A{�(�fk
Z��sv"O8�����h�6}{)�)):>uX�"Od�#�jN�E���]v��S�"OxT;Q��[��(��A^��x�B"O��hsD̋[�$̨e@G�E��4�v"O�T���'����0-Nm��Y�s"O����%�d�Ԥ��	
&����r"O$y�Ȏ�!\܈ӵ,��.��Y��"O��bu$� 	��V.O���z"O���fg��Hevu�Y�r�a24"O^ 
g�V�Y�H�Ҧ�:[���"O��e��)&L����ƍ�+�4tJr"O��9ѯ�x��1bŖ���ж"O�-��K�q��H�a��g��M�b"O�$œ�?��ؐ�6}�y��"O@�x�a� ����s(ϥw�ą8�"OzM����8�0�cd�Xɪ��"O�9�O���*-y��H��(�ybŞ_�e�ѩ�?T�`�HMS��yK	��^�pd��N���0��Z,�yBhf(<�*&DU�ALxK�ˆ/�y�׾7�x4�t	�<��Q�b-���y�� J���1�Ꝑ+�h��ɻ�y�M��
E�d���P��  D��yB��-t����#o�@��x�A@�ybJ�(�B�r�vj1�'���y2����Y��E)8�L�Gl���y�ĶEY6��j�1/�B�Z���y2��z/Ĕ�!�"!F�8wK ��y�!��<2�X�Lƒ/�T������y�ȏ*0�x�:')J�x�I[��yRC͖tP
�K@FF5H]�p��(\�yR�A�UA�@h$ B-N@t��Ü��y����m����!l�LA��ט�y�lȲK?�0RE@�u0:D�u�ũ�y�m � �ĩ�e�S�mLڄʍ��y�P�SR��;�E׸c��Ysԉ ��y��.ζ��,�	Z�B���9�y����
U�0��	(l� j��M�y��߽(I��b���c�J9��f��y�o^ ��\�U*-e��$w�&�y����uP�ė]�D$:�D�yr*��7#��q�׈X�E	��C��y��I�t(�(��EE���G�y��M�(�8-�$J�a��YsN;�yOL�N|����by�h���Ӫ�y���#Q\����E�Z�^)����)�y��V�����A�P�d�q����y�I$fʅK��9�.()��'�y�(�(A����fc����Z�"H4�y
� �@K��kf��$g�+9�z%+�"O���Ս�,������	;ېa�"O��Y=
�s6���E�����"O��t�V�?s����& &T|^A0�"O�dY��J��z��1�:]�(�"O��R��H?bԖ�˱�X0���t"O�=rv!)�,P7��S�`��"O��.D��tsЦ޾K�`Pb�"OLY�`�]��Q��
{���"O�ĸ`�${E��C�muv���"O�|�Ε�|�����Ē�m��"O��{����"���!x�5�2�'���2ф�a�	s��;���Y;D`�l> }�C�		h6��1�˘)j@Sa���P�OPܠ�b4+9��O��)(���77BxI���&IfαI�"Oh]�cN�*?��Q*�#��sj���A�>��O���"�3��#xHy�#��:s_�	���T���?�E��E�/H��]��X>"�n)�/�Uh��$~�5���,��ڢ�'�΍���$t�$��+J?yN�d+':Oޔ�w�ѴS�@\�0$�4.=�D	S"O��A��X`��A*��j�y#I�h�,�`�.��B�4L<G�T$Nw&�]�AnB9���Q���ybom� ��ըG|���tcPE����V���c5ʑh, �x��0��ĕ/b(�l3��ԤF�JT`�g��(t1OH\p�'%��O���LīfW@H�B鏡k�jBǖ�	{Ҕ:�E�6)��0�O���p<Asj�i�,�cĬ1����1"_�I��@j�K�hO�� ��-gtz����Ӿ"�Ԥ�Z�� b�-z38��X�� ��:rwb#?J�<D\�Va&���)	lAفN��6�0�h���9�剺O-�ܻ��X�}�L�ʅ$��YR�>	�$�!o�h+"��6#@����j�>�Ā[4ߠ91�-7?�I�#`�c>�!�FP/W�ئ��*a��E�H��qa��A�lz(�*6�Y�7����qO�"A�B=( d�f*C+v�� ���<	������9��DJ[�S�QN�c�io�b�=��	�a_�	Ȑ9k�܌d���A�!e����s�,���Ui�Y1I�&i�f}	% �6l\y	u�^���	( �ܨY�
�2���t�S5f����|��_�x��YABM��L�'����ĐZɐ��'2�`���}|,p�߅/DT-B�%��=��	Y�GG��%�+Gl����gо#/��H���\7����j\&?������\w���T�J��DE���;t���z�" �OY�(�*�:g�����?�h���%"P���{�'A���f��g�g�	���qBƫ�o����(_5^����'��`GO�@���B���_�=��IӭO�R�h�)G�Ht�akElF2����'o�z���
>L��A*�_2ǉB6AO�ٹ�S� [f�$�!G���w���E��փ'�(��$(>  J�O,�HgNɑlGL]�ǫ��@����CaU�(�4��Դ��?at��~2�0'	�q�bH
��D�'R�i�#\9'��]&>]���ɅmbN5W�X�%�8�YBc"D��qA�K�;�N��s%פb���A�(�<)�ϗY��M�SF!}��)�hŎ���EѳH~�iA#G!
�!��,�������0��O�	1��H f4*��qO��)��C�
4Z �U�:<�A�'��y�?��LA愛�i��T��M�l��#)JT؟����I	XO\�2�&P����@aa9�& nK�C|r���0�U^"��e<)�f<�"O�ɸ'�/2v�rF��t~m�[��A ʘ�N���ٕ�>E�D
��(D�F�tH��y��Lz�x�Ś�L�`M�'7�z�'? �6!ZLk�ϸ'��<j2�C$+�|��G�DG�	Q�'��,B�i�-K�1ӢdP$�4˅K��$��M���'��`Yg"G&T��mhg�v)Ç&DH8��ؤj��1O�3u�Ĥ;˄t
�G�"�V0"p"O����	��o*xy��c׾��"O0	p(�E��DW�1��G"O�aba�J6�P�����V�}��"O�8�"��K�'_��V2�"O���Θ�6`��U��o<8E3"OHDQ�b �G����&�c� �p�"O� J(4�A�nu����߶6��|�t"O ���&�#b��Sd�MΈT��"O�4�D���@!�,/�4H�"O��!�ڗWq�y��*rĵQ�"O��!�Gh�V�:��<Di;"O�J0���g�d�XDA�Vɶ��"O��+�e� ab4�*J�,]��"O�U�Q�
	V|��j�K��x�4"OR	s�m� $,�D)�
�
yb"O��PDNS�:@����W2ua�LР"O��q5�]7p�,� �ށe�S"OZ�p�)	Qv���P��;S"Oj0у�8�P���\.COba�"O0<b1Nʷ�T�ѐb�I��"O�I�T&�6�@Ţ�3;��D�"Oؠ�@�Q,S�q��2[�p��`"Oj�����	[�b����U�>�C"O��3�ψ�I�D���◡H��仴"O|c&Aā>APHڲ/I�a-DM�"O&tSL�!�ҙ���C1T����S"Oʙ�Di:]*���,y�*)�#"OܘJE!I�DЩ��_���͓�"Or�#4�Z�}|8��*�tT�H$"O
ꖢ��"P���ç�2`����"O.�)��X� ���d���6��y��](&�n@�B�)��\b���&�yB��9,��P���^���KR���y�	�{�b��E/G:@�6��y���{�&a�G�P:xޢ���0=ـ�ܿh��q�l�R������.y,���O��I<Tt���SQ�<ɱ��K�4As�#	�"(��05oM�<�M̃g�Tx�e�ɍK�<	@RE�<���TM�P��V��� dd�B�<a�A�7<�(����L?8Gr�pb�H{�<�퍹����B�=V���&c�<�cI�&.}P�A[�n���Yt�XdyD_D��چ�� ��Z�12�dH��|��H\M���cJ��!�O�Dn:�fʡ�4J��h�AH��[P��'+�M�4������A?E��b@8��	��C��!x���5��b ���� =���Y}
çe�<a�G�?b^��YąQ)�
��A&��V&�+����LIGH&�Xy ��7a���'�w3������|�'1:��6��� ��O�@�3$�)o���ˋ�
8�8�W+D�C��ɗ	r|yǧM�P��Y��Ea־$	�]�%A����,}HԳ�kN�&����4�IP#��1n]���ːY�����O��I�f_�Ȋ�<�}ʶiݦ)r�.@��Q��@�������$�
V'���h�ӧ��<Q�O	w�iz�Bۉ)��I9#�Sj�<�!�X
I9��U9��ؠ.c�<�7oN���0�� a@&�C���]�<��-`��Df	j� �S�+MV�<1F$�CA��9���. uKc/R�<�$$�G� F�̄�<1[�n�P�<Qu#^�t��UP�ɍ�Ŭ �U�Cw�<�`�$
6�j�e�  �
��[s�<�F���Aӄ�QE.�97���s�b]l�<qT	N� `,�yqJF
J~]��D�e�<	��^�^���2�-�!���6Da�<�r�L$�4#�-�b�-��nIg�<��-E�k{�m�m��R7E`�<�"CӴ`������;�٦�R�<�Q�O�9q�R�.3O��S��P�<1��X�Gr�y�B0}�FA��F�t�<� ���kr%�-5�aC�Op�<��b�
]�hH��B^x�ף
W�<�E��*�3������2&T@��S�? Z�cd�Z�PYy��Y�Q��0�"O�@@F�C�?>����Nu��]��"O:�a ��`t��چ�#��pf"O�$��K�Z�p|�&�R��( "O�9٤��n�0P���QV��z�"O
���2MΤ��܀M<�q�$"O�L
�e�
��W��j "G"Ox��7F^�O����fׂo�L! �"OJQ#�.���l-$g�Ĉ�"O�J��Rǆ}2JU��b�"O�|X�G�'|�ɹaˁ1Z[E��"O���l<� ��C��~&�9�"O���g��4��,ճAr��"O�!; )L 4�� �*H�NQ"�"OFBE*K4���sҮ��Y)�%r�"O����
a"TMW:\��\�"O�9U�@">h�7��e�dMR3"O��+r�;	��� �ՅԞtH�"O�Q6��z8�Q�:B�کH�"O��c�G�>'���)۳,�=�"O.�k���k�l5��h�#����@"O�@8`I����EH��w�B�ru"O�9W�ӡ?RL�j�柭px���"O��R��z%�%^�<�C"Oܼ��"�&=����T�H�s"O�(���*��G�j8�eӕ"Of{��-�ܬp"��V4فA"O^��R�;M�z�B�As�^�Y�"O��C�� nN�0��c[�8�P`R"Oh�E��8��Gc�x|�H��"O$-heA:
��i���7~o���"Olc�J8 7x�k��c��p�"O
�@O��ܔj�ΑbTFQ9�"OB �X^E,�j�h�~����d"O�� �̡hR�D��O�Ҥ���"O�̺�)�+42��։��&ʁ,�y�]�PE�$"'k�M't 1
ڭ�y�Ǫt�����II�l(p�c��y�kR�"��A�4Δ�C삥8K�$�yr�,#ܨHG�4�f�yB!�yB� g���"�ӂ.F�`�F���yb��u����f_�y�Rܸ6d��y�A�g�$��f�3q����P�A��y�a6��iÃJ@�drJ{ ȗ;�ybo�t$�Q8���W]��I�k9�y�o�(w�@�� Z�!q��&����y2j�))$�#���8P`"G͛�yb��)�T��rB2w�TR�"�PyRn�*,$h��<z� #��o�<�R#��9�Z�����G�,�2�n�n�<YǠ\q^=�wO 6��,�֤�O�<�ՠ#Fu)u�5d�i5�J�<����FR8�bQm֘��Q�5DD�<e	�7q̉(6L������u�<��N�u渝y�/�#��2#�s�<yA��J�@�Ȣ35V�Z�F�n�<Q'`�!R	�h�S WM���i �i�<�ui]��0��.YZ�¦a�g�<�0R<$>�w>$P����Hd�<��A+<T����t�I!�{�<駮�u�t�r�iPR"�LCw�R�<іHF+��cbaR�IL��t�O�<9� Ձ<������$�Bb�OB�<�$,U�dà��F"��p¡Bh�<� ���@͕o)Ԕ�2��C2�AK "O
|P���[��X���1��C"O� ��腖h�@�X&+�N�H`j�"O� �d-k:��	�d�+P)@13�"Or]�#��LH�4s5���c�8�I"Op ا���	Z��)&C[�P�0I "O��bDA� PV�|+4��3b#�eb"O�ઐ��~DR���dZ��"OB�ۗ�Ӛrp#��"6 2<Ѓ"O6)i�k�'�.+`M��A��E+w"O�P#D��)*��!��28���"O`�35h��A ��惐�I���cd"O*y��L��S�9�������"ON����E�4�tm)�f�/�xB�"O��#�ܭ/�.��Lȳ~����b"O�h��&��.��0xA�\άdI#"OL)���Swֽs�*�3D"�ڳ"Ov��Ģ�O^� � P�G��"O�PST�0A���h��Gz���v"O�Yx�mM +��=)��
.iøɛa"O�D�U��i�Ea�KX h���"O����T�&���C�jK�A͈�X�"O�%��! �1�,�b�IH�<���q�"O܅���ӂ��Y"�'�����"O\aJ���(]��׬��6%�I�"O�؇��iъ�v�ԷM�Ѳ "OHY�aܚT�0��d@�9�va��"O��1�I��,���N�t�$�w"O,g� �1l������;r���s"Oz�b�H�[F�@����y��t�p"Ox�b�˃$��`	�d��KH���"O���q��)B�zSjT>JH `��"O 0*C&�J��i$k-���E"OF]P%�	
_xS�GyXhf"O��9&�֮k&R\"&
]f�,c"O������$ɴY��D��.fFx��"OX,�m^�t>�D��Α<~w�Qr�"O8��3J�S&v ��D+y`6��"O��;b�S�{v.Y�cA#1�V���"O0`�Ҋ �y�Lp�!�N�x���7"O��+&U�#V�1 �Zh���"O��B%��* 1�lXtN�>n��"O\�(ѨQ�0*1��J�ew�U��"O�Y�6&�)Ax@bK8k�p�q"OHѡ���q�h�Dʆ�\[�T�T"Ol<8S̄
���C��7I�I��"O��*��N8%��H��'=E�l�`"O��K�����1�"��0���F"O��O�+Y�}� `39�z�I�"O�x�'%T{(�DOÿLR��"O��0�A0�6@)���sD��["O���0kނ� p�L�E>P,�"OJ8���=j�U#��EvA�iH5"Oȸ���%c��Z`/�--L��"O��a���6	������#'	f�kB"O�\:k��;�v���P�T&��P�"O�Q{��Շ_�.a9%gD��Y�&"O"��w�� &�H��FB.��T�G"O:��M�n ����r���+�"O|�Q4�$vaH��f�%,��"OJ�b`�2~�v�Q���wL\��"O���q���d��1 F�)U�" "O��Iv�D-m�,��oq $��a"O�t�'��pϰu �G;�	j2"O� q���ǽr����V�3�İ�G"Oz-�ˎ=�,�%`ߐ�bq�"O@��1����k�_r�\�T"O�q� �_� �`�Ĥ][$�K�"O�D�%�
-X<[!^|F����"O��3p`@�I$�p����	8:�`"O>���AQ^N,�#�N�m��UAs"O �P �*[���1�N�!F�E��"O��(�˅�6�	�Y���ht"OV )�ZN �%睳w/����"OڬơN�noX�g�
�2��"O����F��@ ۽-\���"O�jѬ٦I�B�"K1o�Qr�"O�Zw&�f9��KD��h���"O�`�֠�M�d����Ĝ�"O
����
/�d"�H̞J�&�J�"Oƕ�V�P��9��`/Z$2s"O�x���ߦ�v`�0��"��"Or�� ��I)zPQ��0upt�"O��Y�Ι�~!�Ȉ�$�q��"O^���A�B��dX��"Op9x�L@�c����"�>\�Y�V"O�y�5�^�d��#�GXԩz�"O�!I�+�B}s�ыxD�$�G"O�@�dO<X�,��źᠥA�"O�D(� S�B��Y��6$���&"OJ�[��1U�+F�r�{�l���yb��)��3��E5;��0�R$�:�yR�K�;���`�N6���8E�Z�y�C�SZ�+�*��^���ځ���y�%E�7و � J��'��i)1H��y��ٿB���1�I�$�:��c�!�y"oA���w���L�C���y���M��t�4�47�n�!C����y�a�6� �%D�3{�D����-�yR� P����C�5�SO��yb�ےh�V}aMTG`b�!� &�y�E�DDS7FM8��@��΍�y2������`A��nY���%��'����³<����"���y62��'�V��oݳ.��(��º �|!�
�'$�2Ə��-�.��p恸�FAh
�'WNEy��+T��e�g���q���	�'5P��R���E�+hB��	�'��Q���!rj��R%ӵ[TʹA	�'TV���EݔX��-�� ҺTÊ�b�'"@
�蓯6�&x��U�Ju�m��'4Թ����*KC,4{gd�K���'T�35MҾB�Z��ϗ�-
~A��'��XKH"[l���!@-\B,�'���Qө��SN��V�R94�:%��'�����J@� c&��`�'���'�,���"��=�������q�<�q�'����Ȇ��-�%��uj���m�$�T�ѽv��=1��]:��M�ȓ�8UIn�PRr��hS2&�,��r��)����.-�٨tgT*	=:Ć�~,����O��P����E�xd��
��   @�?�   �  ]  �    G*  �5  �@  QL  zW  'c  on  !z  G�  V�  <�  ˜  ��   �  h�  ֻ  �  ]�  ��  �  ��  ]�  ��  �  e�  ��  � : { � � �" ) 2 3; uA WI wR �Y �_ =f dj  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�OL ��-ѲS`x�F	�P}�$�ר9D�4���rN ��������$?)��?�S�Or�prI�;�؀7��3�H\��'�����U�7��	SP�fY��?!t�'�6U���ۤ;�t	��1�n,(
�'���f�B�|�+'��+X�U��I�$oB�	2I��u*�	V���#�mI&O�C��:�Dbe���A�p���xǶB�� 
2(C ,_�pN��E��$4N��%�S�O�(�ZG��1���p�-�	���'UV����I�';�9pT�8Ǫ\ZM����I-od⼒�@�O�L����A��B�IަّS"�=�-����#���&�-D��K�U�<��њqI��C~$�B&,D���fB�)-y$�Z%�#�r�re 5D���e��t�����Oɰ�3D��IV�!�XM��I�'���!� 3D��:CD�9CF��"O�&7����.D�p3P����h;��vJb�ꂢ7D��"��.�ɥFK�Z�d䂑�3D�����p����Ȕ>W�����'($��1 ���r��zZm�	�'�>ܪ�`1F q`Q-K,wtҔ�'&.M����w܎4��C��uE��[�'����0�[�^��)��Κx��QQ
�'8��@ ���J��E�dqlm��'�\T3��L�9Cf���X3k��	��� �񰇢�����pl̊^�|Y�"O��Rmń>�ܣ����i�421"Ot]
�n�%�Сf`C�'��Yb"O�lY�H
��6�XQ/��%R���%"O<m�$!�6]h5@qm��zHLL�""O"	�tjDZ��*+\�"O�qQ��D+x���O3#�0"Oxq��BUo�Q"rN�&/!H�w"O@q�%��+���#BJ|�v"OL���#N����՗`�L���"O�`$DHA5�Ţ�΀S���1"Oy1V�K�:�Z���M˷BQ`!Ʌ���HO?�F�@Tř ���e��E!f�!��J+slp�{ҁF�,.L��e�͜vg@L8�8O"�p?���
$�Hh��-7���k7�c�<�4��#8SL$3ĭ'H�ē��_y��'�J��M�n�L}I'֣^*�L�K>q�O��?5�O�D���#H�a��hA��P}ڱR�'���	��^��Ҽ�@CU7z�H@3�'����Ȕua6�{�O�?j�n-q�'�VPa�̃�&l��r.N�ZYF`�
�'�p ��2`�����(�����	�'o*r�凔�<%+�$D>�{	�'vt�C��7*�Prt �1B�ѹ	���?K8H�6���m �
@m�O����ȓ)�� E�����h�6J=Y�$�ȓ/ͪ�yE�/;ԙ���6�-��P��6��1�ISSjױG��A��~�4�+C�G�[ r���c�[a�,�ȓ�Q�lP�L]��	V���ȓa�\h���Ͷ.p�A,�RC�0��1�.b#��A��\��Hڊj����gm	a�D0KM���M	@d���-R&����*t��X�ĒlQ@D��oLؽO�Sߖ����pzt �ȓ
9��ײk������-�$Ԇȓ#����KI�=�p豇/&�P���HR!�K�B���qcM$"��@��;�\L��R�*hea$B�)r=NQ��N�J,cH�M}^pzQ��&j����ȓ{���`Q�gpٛ��,t˦Q�ȓ` <�Ĉ8�4�s��*p�-��Z�&uP��G7�ܜ�G`ƿI(Ј��D� 1�㇣��L�D͕9/����ȓtF���CH�MkH��nR7N!p܆ȓCUf�Am�,�r�#QA~��d�5D�@9�ƖY���`@Z+���0(D�x��@U{7llc��C�n,� �q
&D���Ç�5�\Af��Kӌt1g&#D�ĢS���PДI��m ]���� D��Iq�¥y��)���+@��$a,D�,���25 ��Ӊ^)Cl�	��+D����[gE$����dZ��6D����$��F82��P�+��4D���G+�o����+��g��pQ�7D�8�Z7��<B5�A&	x�V�9D�<���J�O'�1�Ği�NȐ@�+D�L���] ~�V1����t	`�C��(D�@S�C2q���S���c�V0��%D���$�E�r̈�i�%O�F�GH/D�0����,s�*Qh�d�1��0Zq�-D�� �}��1�Q�I�+ ֘`"�+D�\ɱi�4r��DJ�'g�l	�m*D�,ĥѣw����!A>�躄�"D�� Hui�`̎L�`@��/�B�jq"O�G��6��BC��NF���0"O���P.1x,$��� Y��#r"O��!e�3�J���l�#6��1%"Oȕفk�:qVD�1L97
�P�'�r�'���'���'lR�' ��'�z3C�&�l��	S�[4����',R�'��'�b�'���'>R�'"�q�SfVL�k3n�-������'Z�'���'���'zR�'�b�'���(��12�"�1D�U�n��Q���'�R�'oB�'��'�"�'�2�'�V���%.5��L�5C�ɒ�'s"�' �'���'y��'���'}p�����"�Pآ�#P��$�G�'��'�b�'�2�'�r�'���'ؠt�Նm^�X�'$P�Z��H�w�'R2�'yR�'3"�'hB�'���'E�����t���EL�.�<�B��'R�'���'�"�'�b�'���'8�t�_����LU�j1`!3�'��'���'i��'���'r�'��%��� !s�\�цD&4ݒ�Y�M+��?���?���?I���?����?Y�e��[����%)�f������?����?I��?����?q��?���?�᠄����Z�$���b��9����ɟX��ܟ�	ퟌ�I���	ҟ��	
_~�����D7����]>:�J��	����I����Iʟ����ڴ�?y�!��ГH��$���]�n@H������D�OZ�S�g~Bd|�fa!�g߫zgB� �� t�.��b��Dx�	9�M����y��'�)0fLG�p�E��0�ҹ��'���[��֙���'{!�4�~Z�g�#-�и�fw��0)6��B̓�?!.O��}�w���Qب �"G�!�q� �;[�vf]���'��(dlzމ
�+��!V%30CF#
,�� t������	�<��O1��m��n���I+17�-��G-sP{�*J������<� �'���D{�O�R��>`/���7�ӑ
Ŗ�ZqF��y�R�'��۴-$�Q�<9Qi�c�B8�t��Z�Pi�)���'7��?���y�X�@���'o[H�(�Kx	2&�E��	ϟ����V�b>�
��'�D��v��8�B�[*6�� ��佔'I�ߟ"~ΓY�Jh1'��2>�8���I�
#� tϓP`�F�J���$Q��?ͧJ�|94  |����EΓ�?���?y�,�:�M�OF��j�E���"(� �Ҳa�~X
q�H�F�O|��|*��?Q��?���`��F�V^������N4.ű/O�1n�:w�m�I��\�	n�s�t�#��O �X'�ʚ!�V�*$,ǩ�������ڴ[����$�O��陇%"�}�bD�wQ�,�>�4��A�X?h��J !ZH1�Ӊ�r���K�	��$�^-zĈк.;yr3 ��*
�d�OH���O��4�˓p���?�B�D;[0̢���;��= ���yb�c����h�O�o��M�u�i{�+gA��+���'Z�s` ɰ @�:fG��:O�@un	$]> �H�����zI����֝=��[B��2u�0�y�&P�<���?���?I���?���Tşpؚ��J����H@��&Q��'�*jӞ�֤�<���i��'��L����vބm���B�A��)ӁO.���O�7=�X��G�q���|p.�
�D�iCT��ȝ�'��V,�K.��Byr�x�0��?i���?���MӀHK�P�U���@`D�m��	+���?�-O:�nZ�v馽���L��w��jH:)
t�R��gNh����_���DAy��'B�� 7��O��$nI WYLaB�!�W��tG�hՖs�`��kM�6E�<����"���'�����Q���9����H�c���ej�ݟ$��ɟ|��ߟb>�'�7��W��m��ӄI �d8҆�ie��9Я�<���i��O�d�'��6͛��6u��N��<4�p�`l�=P��nZ��Må`W�M��O6}��nJ���U�(�����;4,��5��a� ��T��3�M�*O��D�O���O��d�O�˧&�U�F�!&V��� ��#c<tX��i��2�T��	Q�ƟȈ���[P�	1")0�3���m� �2HʬeԛFe��&�b>��V����=�{��2%��2=���%l�$R`ΓP�`,�����'�7m�<a���?�b��5+˄�b�
蜈[U� .�?����?	���F����mE����	ПD����tN
��a&�U�&��	��MD�i,Obq�焳B���u��,���*���d�G�VU��n�������;�
�����-*���P�7��ԫ �,��@������	�����j�O�$� l�ȉ���7&v�	ؔ��5L��z�:���D�<�3�i��O�P�l�*�XAȝ1$D��5	�]^�ͦ�9޴B.���ӛ撟r�oR�0��	!-��������b>^X�@�@�R�,��R���I���I��I�L�'Z?>�l(g�Ё}���$�@Sy�z�N�#��O��$�O��󤕊�
���Ȯo��l��ɲ.��'�t7���5IN<�|��8:�^d�r��O�x I"gI�y7�`ٴ2剓9⤣�O�ʓ%r��^����@��U�D��E � �D���'Wb�'��O��	��M�%�X��?I��L�R C�/!��QE��<q%�iB�O(�'�6�զ�bڴb4~x��G�A&0���؍o��h2'jͬ�MC�'����
M�n�����d���3�{�? H	{v�71f��s`R %Q����8OH�d�On�d�O ���O.�?]���N�@���0�bYD��Dy2�'�6M��~���O�Em@�	!�<I���%�|��B�Fl�J<a���?�'$� �k�4��D��M�[Qc@���{T�K�)32��uj���~�|�^�<��П��	��h5�ڲbP�q	������ϟX��dy*`ӀXs=O(�D�O��'��`BT�7g��2��6���'U���?q����S���_;rɆЛP�B����S0BЍR�o�u/�uq޴��4���8�'��'���(t����� ,.
�����	�?����?����?�|2*O��ͧD���i�&�������	ٷw-^��A����۴��'����?9�EW�u�����a��>��@gC��?�::0+�4��d�/w>}h���l�w[���������Z����y�U����ן���П ������O�$�1
� _djPs����-�1d��͓�;O����O������睍R���SfmԇA@Z�Qs��'�f��IϟP$�b>= �Ŧ=�p̤��f���@	"tBw�CDS��͓nV��0�࢟$&�����$�'���b%��:(�a�CMÕO��A9�'p��'�RZ��x�4x��)��?���"��m��,N���;�i�#~��b,�<I���M{��xRȝ�1�(��g��ECr-��H����$Ϫ:������(�q�DM���o���|��K�e�<�t��UN��i�R�'B��'�R��h��n͎cD�)���N62�L]�S�՟�eӴ #ug�<Ӵi}�O�N�x�h��T)��Y�����D��Φ9ݴkW�v,��~E���L��bψ��T��.#Qz��K=� ��no���&�����$�'�b�'B�'y�|��ٱ�M�P�m����S�\ߴz�h����?������<��W�	u���$鉄�x�J&OԋL*�	�MKĻi��O1�֙h�/����}�� Ɨ$�$łRKM�e �|����X�ŮV�R�s�	]y�e͘b
�`�oՍpE��ɁL�N��'�"�'*�O�	��M�����?Y�FZ�I%>��Q���*�D<g#O�<)u�i2�O˱>�#�i�h6��ۦ�[��� �<��v�V"���cEj�<��m�x~������kܧ��cA�&"r��s��x��י=��ϓ�?i��?���?1���O�0��T��U1�@�UK�	}���)��'���'��6mSm��)�O�m�|�H��׍� �D!P�n^��A�L<A��?�'}�8��4��B$*If�:S�L�'�TЁ4"��&q�mH#��+�~2�|�R����͟��	ǟT�↖���� ��Y��P�� ������[y"ei���V;O��$�O"ʧ��K�.�:���E�3��d�'O���?����S��fO�f)
�y�@1rė)Rhv)�
�:{�搟擣P�D8���1&�cE�6.e�d��]����O��$�O���<�E�ib���`�5�ڹ�H¨n?��T@��/�M��BH�>)��i�x��v���w�"Э�;�%���wӆUm
�ll�b~r���w�4��[�I��;Rl�3�B��H����k�<�
��H�Q"�<z�J)���L�q�< S�i"����'��'!�Qoz������I����v��Y`���`�	��S�' �J�+ش�y2���B��Wd�=����#���y�)T�~_0�������D�O� 08_�h˖/��\�$�s�H���O���O�ʓ�V��L��	ʟҤ)ߦY���Hҳa����E�c�e���֟��I3�ēEp�
2JH�`6-Z0L�&_���'�|[�*�V+��m8�I��~��'p2�)�G��ΆXX�1��'���'e2�'>�>y��1"��a'��2H%������"e!(���M[�Q��զ��?ͻ`1xI2��9>���t �����?��J�֭ƞi��斟X2P�K�	�	rܬĳ�	^.r��X"$�)�r�O���?)���lZƟ�����H��O�9]��r͖+jn�)��ly2�{�,�f��Ob�D�O~���$Ӵ[�^(V�1C��	�Cف,F�'��'�O1����%���G�Q���7'�֍�!�Ah6m�sy�n��������]�V�QKD�^�T
���݊|�$�O����O��4�D˓H��Ƃ( �2��3O:���7
!Nr:��6&	�y j�T��8�O��d�O��m�e�8Q�'ۭ �*�H�
w�49��Y����'(4�HSYb�O~z��[��`��[<R�U�gAt]��Γ�?����?���?�����ON����܆(d��7�4Х�'��'�7mBR��	�O�Em��H�'��)����Bg��rJ�q�6yAe�9���OX�D��h�zĬa�H�	�|b��V�#�,0&D�5@�H%�'��=@ f\�a�O<�O(˓�?���?	��.�
$��*K-V�%:��I0^�����?1)O�Uo�=x���Iȟ��	l�ĤOj�:�#�-o�X$�F�ܬ���X}B�'�ҏ#�?�In�^]��J���9X�RE@�E�d�&��a@���p-O�)���~r�|2�T�k����T4� K@0����?���?y�Ş��ߦˇ�]�X���L��u�28)fo�!�.�N������z}��'�L�I6%�I(.�3hW/�$���'X���?�&��l	�n�K=q�� l%���ɍ�A��@9?�l�z�=O�ʓ�?����?��?i����5n�������9cPJ�rU�B$��o�����Iȟl�Is�s�������dݐ?�.�H1�@����s(W�?���򉧘O4�)��i����b���`��"*��;8��!40= �'��'��IꟘ�		ISt-zpʍ?]ɞ�F�V�" �	��h�	���'�z6MQ�<N��O�ğ�@U���_���[�ƈ�����A�O����O�O ��� 5����O7T��`��� 	R�Y�`�l�q̧.���	ß��aJ��X���
C[5B��AS�	�����������F�t�'�aq�m�+~I�g�'cg��h��'��7�U1y�Ɏ�M��w�L9k�J��=���l-�+�'/2�'�"ƞ�:����������)�`�h�˳~�}�����X? �O���|J���?���?���i�\�D)\m��8�cO����/O8Io�B�0���h�	v�s��#��P.�r�!5�/P�(MRч�6��$�O��3���I�/���PWb�/y:�ԫ!���>B9ib�gӲ�JB6�9�d���%��'.Bљ#�ې{
� J�%0�]BZ�M[��?q��?ͧ���Ҧ�,	˟��U�ɶ
�����#E�D���f��;ش��'�*�g��6@w���n�1/v�2Al�C�x�5E�8��D����'�����K�?A�}��*Mh��`G� N�P�SA�Y*o3*�̓�?q���?a��?i����Oj¤��-�,�bAӉT{�x ��'I�'YP7m�!!�ʓ��|�-CZ�ٔ�ļ�&I�A:w�0O�Hn���Mc��'���ܴ�y��'�24��� '0Ͷ��ajE�
�$qF`H!zP�I���'�i>���Ο,��6	2�E;�MK#4���c�"նI����	�Ԗ'�B7-S*A��D�O��D�|�Zmm�!:!h	+.��(D�Q���I����Ob�$:��?�����4p��m�	5��=�`(�|�d:��������@j?1I>�@�B7=H�t��4a����?Y���?a���?�|�)O�n�@w�rT,�',7J��k0�6�Р�X`y�MbӐ㟐�O`l��{+�HSc�9�V�Rr���(�ߴ h��ŝ$ܛ��@�hY�9��4�~jc�� ��3�����9���<(O ���O����O����O�'4�Tȑ�J�"�.���'7���s�i� MR�Q���	X���P1����$lY./<iǀҶZ{,Z`����?���w���O�(���i*���<�ys��>R��!Js%$.��7����'��'��I쟠�	�R��a���P���9���1! $�I۟���ݟ��'+<6m�`�����O
�ēH,m���/\H木C��.w�:��@�Olho=�M�c�x�A�&��H��	��QS�"��.L�ps�e�?N�1��t3�D�0����t!~��%$}�D��ፅ �"���O����O���%�'�?ɵ
A�ܮ�!�]5�uH�ʊ��?��i
\	�[��ݴ���y'��N��t‎�*	}��0����~B�'���k���T�v���>X
MhS�⟀tjU+*/�ە�	�3�@�)���������D̛��s4���i��-0��'��6�Meg���?���?���gيm�!&"�Pb�{F��?�*Q���OQn�9`
�I��jƃ�_`�Q(̬pΛ�F�<�"�ÎLbl��v�	gy���'*���-�����34c����'�b�'�O6�	��M�a	�?���1B��Y�d"��:l�p I�<���i��Ou�'�6�R��Ya�4h�<��u�L�g�>�˓Lؗ]/�Z$D�Mk�O~�؁�Y8����4�w�椹U$G:[l�7�"^��@1�'D��'��'��'w�QrEm�7��S�(��R��t�wn�<���el�g\���'A�7�8����P?�dJ�%V�!!�J�nZzt,-&����̟擱��,oZw~bIQ��4�p�-�`2Q�^[��M�s@R?QL>!(O��O��$�O� ��Jۣc���(� ߂���Q��O��<���i��]y��'aR�'u�� ��ŢK���i�W��!��	蟌�����|"�pY��ID��*=��HX0�$dwn�x�%W�Ӝ	�4wC�I�?q���O�Op���"��0[�=��虇�Dyr���O6���O���O1���қ��&C���EB�A�.�c��!����On�L��Z��I��0�T�
f�i1Lή<S0L������( �oy~B�9IX�}�4����p�ې�ܚPDp���W�<I)O`���Ot���Ot���OdʧfAh��c�ػe�FXI�@،6�X4�i���q�'�B�'���yrEc��.F��,���֑L���3h�}����O~�O���O���f��6-|�x���j<0p�D�7w{� �t�o��@����H�$ ��<�'�?�rl\�y�h�#Ak!2��C��?y��?Q����$�ɦIjE���ߟ��5IF�jl������r�(2s��k�Xt�I>�M+ǽil�O��E	ʩq������3���%��S�,�9g��p��'�S�o�ˇٟ@��"�,af�I(v׶��!hF�������(��ʟ�F�d�'F�Ey#�6Ԓ���=7a�����'�X7��s����O��ou�Ӽ�
�K�Lܰ"BޱP[�) %��<��i�@6-U֦pe��Ϧ��'���Q�+Z�?i�� �P��=�lY��0=�\��g/�d�<ͧ�?����?9���?���/2x\�`��V.E�$���D	��uC����۟�k���'ln�3�(*�b0�G�Rm�٠d��>Yt�i�~6�L{�i>y�S�?��c�_��	p����M��s�C�177$1�+'?1��mm`�dW������8p�8��#�6�h���p���d�O0���O��4���53�v�/ED�d^-娅�f��)�Z��Ö�y2�xӺ㟤��O�lZ,�M�#�i�8�۰,TW=ڠ�����G�f�Ap�@J�&����A�N��T����~	Kp�\,z�=���G5Eh��R?O����OX�d�OZ�D�O��?!�ABه��3WoTy�Ԡ!0��l�I�P �4t�\%B,O��o�D�ɟe^�d!��;�*ѐ�iJ��QN<�6�i�6=���ȷ�m���=��U�'��-��8���%1E@�WIQr���č����4�����O�����4kO��y%~d�WХ5�h���O��c��F�E%�y"�'6RX>i��)]Bk\\�E.gd0!�0?i�Z�������%��ǟ<VeճC��ѡD�7^��u
�?`3V���"��y�'���`SJ?	H>�PĄ497:�� 	��>��r��?���?���?�|")O��m�ts���'�E?`B�Q�.��x��Г2-?���i;�O�(�'T�oӢm�>�s�B�
�d������}"�'pN�R�i��D�O�}:��؅��s�(���u�M�ӇU�V���@�L�'-��'g"�'>��'�哜 *2�i�dО#���d,�l>�ИٴT��	����?q����'�?����y�,M�&�8��b�w��k�˓iR�',$O1�"q���iӂ�I�H���"ECE�)��
2|� 扟.4� �O�O���?���x��pѧӋAF�4���A?4�0 ���?���?�+O�<m��~ј�Iߟ��	R
��RPfВl�D�BJ^�X���?94Z�X��ʟ�&�'j�' �ADI�H��RqG%?A�H�<5���z�4�OO����?U(�1֤��c����\�j5�]��?���?)��?���i�O����]�@�9	#C�(����O�o�nw��v��f�4�4���ޱ\l�KāE2!�r\(:O����ON�d˅X�:6M<?!���%��Ә��`q���A^y V���%�p�����'���'"�'�XЊ���e�i%N��LSP��#[� ��4i��a����?!�����?�f
�`�*<�2!T*B�Ă�$�|y�	��	���S�'|S��#�jҀ
q4%部LP�l}��3�8��'�ܱ�䦑ʟL�G�|�V�0�a
�B���Z�o(g	�4I�@�ğd������ڟ��Ny��ӤɈ2��OЀ	TAvC~1d-�=~��1�4�t��4��'�`��?��46a����}�d�Q�	��Ö	[�9yL"�i��I'l��;��Odq���n��Q�u�5$G.��\a�A��P[���O,�$�Oz���O���#��z��P∣g���SP�\)=����	џ��,�M��}�D�{�l�O�y��53��2�� )�B�h ��g�����lz>����ݦ=�'�<9��%�Wt�`m@��@VN�^N��ɒ��'L�i>����T��D�4���Bۋ1e"-[Ӆ�C|��Iߟ�'h7
q���D�O���|j��W`��7��tѱ�~�-�>����?9�xʟ:akS�g�(и��K6K4�[���Ё��	|T�i>��'��p%��+c��r���HJƬx��n��� ��ğ���џb>��'��6m]�s�n! ��Гmc�ؐW&�)�6��ժ�<�B�i��O���'۫�լ���L�&;xݨB�&o2��5�{���mڠ
�0o�r~�/L�&%z���c��R�!�ؼ�@̊�Q>�a�����P���<�ߓ@�Ԑ
����&��"��a뾀:��i�"x��'X��'����oz�S�*C00��QZ����*�#�gP؟���%��Ş9Hb�:ٴ�y�A\� 66�8,�1$[���vݤ�yBcӟS�$�������O\�d��_��"�@�c0⭯?9τ���?���?�*OH�m�g�b�'x�&�# tE�`BĖ
���*i�O 	�'�p7�Ȧ9�K<r%$;<DL���M�%	>����
u~b�ǴDwlXs����OlL��C"IɨD��� NO
:��E��ڐ
���'�2�'�R�s��C@,O�K{b��B�4���;vȟ��p*�4��!+O�il�f�Ӽ���G��A�#k�m�<��p���<y��i�f7�������Ӧa�'۴��U��?)!��ɼT�Rd�U�!%<�-�-�!>X�'9�i>����<��������o�݋�C)d�d��`RN���'��7M�+�&���O��$4�9Otd����>/B��〣��d��p �r}r ��9m����S�'w�d���"G�|iᐣ0��8��OZ�#}���'d�s�`������|�P��y��٫�BI���Ă#evt�G :�O��mZ-f����	���XY`�X�%��P�������	��M���e�>���?!�iڬ�(��b����&�0/~����L������E'̰*8��+�	��ba�5B�8baҷDI mCN}8�5O��d�O����O0�$�O0�?��%�$i�Ɖ�!_�����!
Zy��'�7m�:P�)�O0�lp�I4(���˚L��Q��@e�I<!��?�'-�FEAݴ��D�9� .m�p��4��%��BI� �P��?9�j!�d�<�'�?���?I���u����h��[i�9�@�Y(�?!����D�ɦ��a��<�	�T�O�#�GV�?�a�LZ�Z���8�O*u�'��ir`�O�zS�9s�mR=Y(�ا��g��Ԡ������%B#?�'8%f����LF�x7���o�|�2�kИl,�x���?����?i�S�'���ߦq�V��0���mU�fT��0I-"X�i�'��7�'�I�����Ѧ�1��ԗ(c��@֭��u8@��wK!�M��i�r��d�i���(�ΈHV�O,�'a3�T�Ħ��B���S�+5H�Γ��d�O����Oz�D�O^���|���ܩf�|D؁��2|~ ���,N���ֆ�9�I��l�:��y���	V������d��A�ċx�6�����M<�|�Qω�M�'+�����n��,R���UW\|{�'(��������Ze�|�[��ßd!�n )�Y �,נZ`͈���ߟ��I̟��	Ey2l�"�����<���vu��(�|N՚��/E���+�˳>���i��6�Z`�I̺�Qc�ڽQ:e������y�HuR�]+v ��|���O����+K��AS+{V����Ь vސ���?���?���h������inp2eb�� YΡ��I�R���}�"������M���w��(K����	`B�G�N�"љ�'<7����1��4S�f�ڴ��$�q��I��'`IU�cK�g�"xSr��f�59�0���<�'�?����?9���?i�b��2I�U��Lq�D��4�˜�?�d��a!�3w�����?���0��6^>�	����!K�T��q�E\�4����O�nZ�Mk��x�O�T�O'�Haq��>��¦�I��f0Y�
6�����Or̀�FC�?ѧ4��<���b�m��H#~9-,Z���?���?9��|�)O�Elڗp�����N\�5&�d6�z`gۧD���I(�MӋ�I�>��i?7�禹�!�O�@�j� KD$�)��ځ�l�oZR~�̗=k�`���~�'տÐm®}|�D�u�ODA�!b����<����?���?i��?A���`�waL$��ڃ&d���BߋYB�'��bg��)�#;������$�x�)۠^�zQ`�k��~�;�L�%�ēu#���h��IC�]�7�8?٤gA6o����u�+e�(M�Be����	6�R*Hb��Hy�O�2�'1��U4wڌx�I���`�#�g��B R�'��Ɏ�M�w�щ�?����?�+���U3�����)V�G�y�e���i�OBqmڤ�McE�xʟl�y�#�7f��h*���4�$AZNƞi8T0FϞ�d�i>�h��'�T'�`�� �)p����ʈ�"�����V៌�	�l�	�b>��'ފ7-�
M T���Ȝ4^v�4mծ��i��d�O��D�覉�?�[�4��4�`��Mʋ�4\���	\(�<�g�i��7-E�{{6M;?��-��:�I1����8� |��&Nu�`�i�2�yb^���I�������4�	ڟ��O�L��-{1�:QB�q�4(ԉb��(wO�OF���O���D����]W� 9�+�LvyS�|1C (_ɦ�3�4f����Or,p��i~�� �H��!�9\��}
�g�!H�$đTx����u|T�Op��|"�d��m�g%�{F�XnG������?a��?�/O~�o%\�]������	��r��"ʉ,6J�M�Ɲ�0^��?!0W�8��4	n���3��N"&"�,;���<pɛa�9���D��$c�Ȍ:}r�=�|��(�O�=��*#��24B�9����U��1q��1���?��?����h����	�IY��I1�s��kF포���DЦq���RXyR�i�B��]�K��8Z0	��Ju}`D�5O�\��MB�i�6��I[�6m1?�4@�d����ޝ'�2��s�۽�Dp��#
��t�rJ>�)O1�1O�)J�Έ�k��@�s�U,!�r�A����۴c�֝���?Q���O��\;D��l���逥YQ�����>���?i��x��M�=Y0�ez�hʤrP5�W�Z�t��ӿiS�˓C��Т����$&�\�'O�X	�J��	��v�X�XW��J�P���ØdK��`J$�h|�HEh�m��Bd�b�L��O����O��oڅ,� �� N�9Ú�@�l�-@ PuzRJ�˦9�'� A�@�arM~��;��:u��5v�⌻u�I�����?��?����?I����O�&E�(�r���vjH�)4��'���'��6-��@��i�OP4oZx�I�G�����E�5��FŅ	hx5sL>���MϧcW���4���أH�&$D��eWx��r�̘`=�$Q�����?!v�7��<�'�?Y���?I��F�%�l�b"�I<=(E,Ŏ�?)���d����$��Ay��'��S&�y�%&�L�F��[�v�=^��ll����S����;,�12�E�"���3/)V��ȸ��59PZ���O�I��?I��!�dF7.�u��R4w�T|rd̘"4J4��O|�D�O���	�<��i�����2L�6)��F�\���a�R�y�2�'Z�6�4�	����O��qu1P������e�$p9��O�o�+,:��lP~�显|X`��q�I8&���5'89�]�vX�j�<����?Y��?A��?�.�~�c��ݗJ&���#]�$i�aC _��5Y�ܟ��	���&?���2�M�;u�3,Ї
@��� D���A�iC�7�CP�)�S'h/f�l��<� 8�QD���a��L"c0袰<Ob�ib����?�1&#�D�<�'�?��i'�n)ժ
�,ix��G��#�?a��?����D���P.y����埼��a�P��1#��#,��
k��/��	蟐�II�X��
A-^P)ؖˎ����5��!I� l�ŢuB�����sѡEH�����b��.��1�c]���	ß<�I֟�F�$�'`�%�6���J��`��͕.�0\���'G�6�F0#����M+��wZ�i�b��ज़`(ǻ%�T%��'�2�'��C�V����8ʑhɹU��Iw�\��K0�B$B��2�ƓOJ��|:���?a���?Y�^�Bp��_CZ�YV���0n@�.O��mڗj&f������Im�S��t 僕�;x13b�Kf`�a�)�	����ɦ�ܴ7N���Oz���Fʔ�G��0�'��չ�'��=L���O��sw㌎�?1u�(�d�<�%BWȌ雂V�hY61�C�R�?��?����?�'��D�ڦ��g����/;�\�� ӣ ����X�� �4��'��'C�&�s�Z�mZ�&�x����.UiI�cΓ+L1�`D䦩ϓ�?9se�)ZN����E~"�O��f�Ou.�KQeW?�@��B˖��yB�'jr�'���'Kb�	Ǌ-�©ATC?���S�5�v���O"��F妵��v>��	(�M�I>�ǂ���4az������+f���$�Hش7���O_ji���i>�	<�>�������=g�|1�2/G8r�yڱ�'(�'�h���4�'�R�'sbQ����}�$�%ͳ���Xw�'$�X���ڴ@.�8���?������;�~��&���5�9�DcH=,���%��d����ٴ[*���iTҡ[���H��w���q����Aʴ`�a������h��AII�Ɋt/����M3l����vC�	��T��ӟ���ٟ��)��Qy�f{�6L�B������Gl׶Fc.`��ܘ5����O%oZG�X��ɑ�M#5��!)bF(�L��5VL����l�F��w�q�b�/`p���矐�Oǖ��
<f���J�A&�.U3�'��	��P�I埄�	��Iw�䍌�MI(����A��=y��C5��6-ˌqs�ʓ�?�N~�����w�0�1���P,�ْ��{�t<�r�'��=��� ���6mu�����v�h�F%�`.H�§i��j7���iQ�d#�$�<����?�m|��� k���P/�?���?Q����ɦ墒o���	џd�B#�2F�����t׾�y2��w��!]���	�ē�Ne8�ٝ`{���U����'����A鈍����/����~B�'�<�[eɔ�:���e�T� ��'�R�'���'��>��I%+��(;s� �u~����s�6e�	��M#F����?��WD���4�NPQ�n`p\p�H�H�z��08O���O��n1(�!lZK~BT�T��H��.?�XpM��!1��Ɓf` )�H>�-O*���O ���O����O(��p'V)T F�G!��}\8� �<)��i��I��'���'*�O���ߺuʤ���	��^�z^���>���?�"�x��$�#5���.��j������I�p�\��'"��!�)
K?aO>�,Orl5k��3�r�xQ�8Z�:	`�'ɠ7�ޏU�z���}���b�eN�E-T�r�d���dM���?�2[��	̟��ڴe�T�:ƷdY5��(�D��LB��]l�w~2%V#=���'��'促o\9+� �x��Vm�(I���<�
�2#�Q�OǶy�\D���L?{�H ��?��~���T���)Y���'����Y�Zg�axC	ߕa,���oC��ē�?��|
����M#�O��{�lI�I�t�ڵ��Ptd��Ąޢ���'��'R�	`��B��X�=�|qQ����q�<iGxR�pӦ�Qs��O����O��'5uPu�F�-W� ��:rd�'����?Q�z`������s�����#��n�8��M��L��*��zF�7�Uy�O������"<�H��'D*~��|x�d@�(���j��?����?��Ş��D�æe���B7i��P������s��H�2�(|�'�F6=�	���$�٦%�T���.�<��ƪ��9�0b4E:�M�Ƶi��-���id��4.W<��F�O��'"Då��#1�ԌZdc�A�Μ���D�OZ���O �d�OH�D�|
�gD�i�����?I�}���F�J���	>��D�O��?�r���c�g;� �@	�I��F��?�����Şƈ�ش�y�fG`�� �߷�9�$@կ�y2�B��e������4���$I�TM:4��Cq���Y�����OJ���O@�D�<�i�~��'dB�'���8$���P�`�3���8:�h�G�dF}"�'jB�|R!��dh���}�t��䚊��ė5�Dd#df��c>�&�O(�d��^��0h��n��hw��<�(�d�O���Of��&��#7!�����B�l�@1H��c��?�Ӹi`�R�O�l�\�Ӽ��IW5th��IB�P�#{.��%��<A���?a�=�LKݴ���ɞx82��O*�"U�R,踑��P���|�T���<�	֟��I\�㋆�mn��'%�T:��v�My�y�(���)�Oj�D�OR��h��Ђ{O���G�M��\�0�{�xe�'���'/>O1������ R�l�6���z�y�H��7	]0\=�ɲ��Ո��'�zH$���'�� �"�)s�H��e �qr�D�#�'p��'7���4V���޴`͘ԉ��Il&&'ؘ:(����,��̓z`���\}ls��Ulڥ�M34��Pܞe���%8��<S�a�y5,�	۴��ĕ�0�����O�'�F�v�Z�*� �z���6���y��'.��'f��'�2���'����Mʢ4?���soHBKZ�D�O���ঝ�rMi>-�	��MSL>I�B�D�z�%߆3���Z2*�@(�'Gl7mM��	�ho�y~�HE��r����/z�<��������J���آ��|�Z��ßd���<�$$�(Z*����k���֦��p�	ry�g}Ӭ�� ��O����Ohʧ��F�]��,�`^�1��'�:�!���Ӑ�%��' �T�iLuծ���E��,`��( *րK�t�R�@~�O���� Z�'A4x13BK�T�bȱ'�Qjѹ@�'��'`b���OW���M����}��QC��K:J,���*B�L����?)հi��O>}�'�7��c�b}z�햧�rYfo
�)��nZ��M$CD��MS�Oxu���U'�
N?��E9�bQ��%׀,��< �	q���'��'�R�'8R�'#�+4 �a�'Թ?\X$f�1�@!۴ט���?	����<���yG�)�l9�Ć&��ų�R�|"�'gɧ�O~8���i��D�Q�,�a� ٰ$_`:p�X��RU
�	{�'��'��i>��1#(aqW�Eh���LB�d�����ޟx��ǟ��'=�7�S�j:�d�Oj��ק/���a�cc���f��%�|�p�O��l���Mkb�x�N�5x���هjX�#���� ���հG�˗�
21�8Ћ� 2����1�\���)�.e��0gM�$&\�D�O �D�O��d1ڧ�?4���_�P=��B�IB=��X�?�w�i�t$AY��
޴���yWl�l��8�ߚ0�8�"�+�y�F���o�M��R�M#�O`@��Y�r�����օ��fˮb�"|ö!P*^51b"
ӄ@hTC�H�2f:���&,�h�h%@8N��܃7#U JvѢ���$���K� �+�~��G�-c�|��Q�.8	�so�qe���V���@��3�=!�. ��E�ʁJ� ��i[��ũ@KCW�$X(� ۂ頁�"�(���P�̀�,�]�Џ�m
� 3��K�t�h3ވ��ax6���S�^Y(�*ʘs4�AK#O[�W (�Fl��t�z<�"�:۵�����9�/��g���M^�K'p�Y�Ƈ!8HP��;���Q���+}� �$O[�\�����M����?A���"������
�M�,u���˙L��I�ez�T˓}�(Gx���6�� Z~P�-k����Mc�8�>7m�O��d�O��	g�Iҟ��WNC�T0tx&�U7(�*谵Cʁ�MK2X���D�DW*4&VX8P�^}݌�ks��6z��<oZǟ��	џ���+�ē�?9���~��P�$�8�(��2o�D���S���'�{�y��'�2�'�p+&� ̚ܐ���@d��u�����US��&��	ϟ %����,�&�F�*Q*�R��׻3	��3J ��<)���?I����K�}��Q�Un�!X����7ʃ�q�f�;Í�u�Ɵ��	A��Fyb��"�I9� Lw� �Ζ� ��yb�'0B�'�ӆ0 �e�'Q>�Q�m�����6b�1��'����P�Ly����\�"ü����m�<xc*G0f��IП���՟4�'_Z-�6�"���0x�9C��u	.� C��,\؈�nZߟ���eyRT�����%�'ͬ��0�������ŉOc�)�4�?�����E׮e$>����?}��W�:�,r��&:k̥�G��ē��/�}���	�CĆ��� Ú]q��Ӧ��w��fX�l�f(��M��X?Y���?1S�O�A� 
\��*gڻ&��8Rf�i��� X{P#<�~B�وe�K�~Ɲ1��ej%[�Mk��?�������$; P>t��GYo��(�����F�oڹ} D"<E��'*��R�KϬO�J�`YK~���,�'�Ms���?��f�8A��x��'Lr�O�tc�P;�
}ؓ��&B���5�$�P1O����O���:c�x�m�PV����<���m�џl�Q�����?��������C[�f�Z�;l�B���.Z}���$̘'H��'��'�r���⭐EM�o�1HP��9�_�p������I{�����I�H���إi�����Ԫ��#��mc"D�0"e��?i��?����?�r�����ȼAB�a��>���KT�܋�M����?I�����?A��B7P̓���A�!�݇&�
!���BA��Q��>)��?����?�M���B.�t�$;d���a��J��c��U]J,l�8%���Ijy�/����$N"��F��:�d�F昭��oџH�Iҟ�	�kw�L�OL2�'8�@ն~eYE�M�9y)�2���GM�O��D�<q�U��u^+A���	Ѯ>��z��D��Mc-O�14��q�	Ꟙ���?�z�OkL�$d�X�k���
{��8sᔻ~����'�r�Q�;d�O�>=��f��|>PUau��,��ER��p�t(ȁO����I������?iA�O�˓-3J +8$uq�g��1�hQ�i��L�a�d$���܁�)��m�`�R�>$��}��$��M[��?���_(��W���'>2�O�Dƀ� .���ś#ׄ�0f���e1��O
���O�DC�? bHғOR�q�St��.2NB0���i{�	�tB�����O�ʓ�?�� ��4��U�q�m��O �;HD��'ϖ�Ӳ�|��'�R�'�I�tɖBmL�ರ([�9~&y���K%����<�����?���F�\ʓ��$#N9��`�vjB,a��1���?���?A*OM�DY�|����</��h���$������'�ҝ|B�'����	���(_2�hU�͕} ���E�6G~�I�D�I�<�'����ϯ~Z��_d��­R�Ftb���8Cڜ[��i�b�|��'��'�7u-qOJpc%Ɨg�D��1�Id�5Y��i�"�'>��6f�	��t�$�Ov����,hh��q�����c�T8VW L$���	韔i6"Hl����t���1�.�c0%��v���ǋ���M�.O�P+�F	��m��������?	��Ok)!��$Ⲏ�+d������4ԛ6�']Ҩ[oI��|����r8�D���~HxW\Y˛�e�aHn6��O��d�Ot�	M}�^���o[9cuD��#Y�O�ظ:����M�W�ƪ��'����$�1C#$ۃH�L�u��}>��nן��I���Y��
��d�<����~�(�>$���"]d����#2��'�����|��'���'K��R���P���	�5�,z����F^��9�'���h'��X&?���`��1C4`P
��4���l�D�I>q��?!������P�~�BfB�#�\QXgԩ�$���m}�Z�L�	U�I�H�I���-A�M�W �9RG����b�X���`�I̟��'�:؆�>�wAƔ!�0	���fa�G�p�$��?�L>A���?�%jF��~�K�/�d�FC��q�iA5�����O|�$�O�ʓp]
������˛|���)T��6X���P�fȨQ�7m�OL�O���|����S�w��8>�����-z �4�?)���D"��E'>����?��/�"�� C�C|U�U%C�cN�O��G��L���䧦�)^�n�,q�CҋO��@������O��O��d�O���r�Ӻ����
8�d(��E$X��a�ަ=��ڟ��M�4?�c�b?!�f�Qh��`A��%��X �hi�x`m�ݦi���8�	�?M�K<�'"��az@�S��۷!9S�%�f�i<$����'�rS�0$?���q���}�ԕ!7�X�����i��'����"�)JO�xz4[H ��uA�-�ŨE��'#�q4G:�Sǟ�h�L��4F�V��I��#�y�5oZ��3�uy2��~ڍrj�FnL���`]).Ъ�L؟	n��. 9�o�r~��'B�'�剥V��T3$EW�6Z|9P�.�^��)�dK��ē�?������䖄&l��� J�4�Տ,q�\H��f�O��O����<A�n�n�{�O�9���O<T�B��k��H���4�?	����'�b�'����a�H��M��?V��g\�|,�* ��n}��'���'O�I<��,�H|b�O
hN����K�S���ԧ�.9��'��'s�	����IR�i�5R�(Y!ʸ-
-�QfW\[�V�'<bS��&) �ħ�?�����Gְ~д��U��E�<AB�S�IybD�.���ӟ<W"��3\�����2,M�+�Y�����k+���Iן��I۟H��YyZw�N����%R�������cܴ�?���S��̻ŌGA�S����	a��,C���)&�V�_�:5o���N��4�?���?�'����\c�.x�b�W�Z�Y�-�D�*�Yݴ"���b���?����?��'��I�|"��X�Ni�%IX�i�>Izv
=-���'���'ײ�˱W��'��n��}�u��`�`�� ɞjJ��y�$S�b?��I~?A�@�[�P���O&;R�yQ�����	bN���'��맸�'*��E�P����m�8P�Hd{���>���4�8|�<i���$�O�ps咿bV�S�ΐ&CPX8uj��V,��?����'2�'-�EP�M���T��[6�}bq휛T���+�yR�'��	ٟ�!���u
� 
�&|�ш�6�����-��ǟ��?���?����\3<�oZg��}�G���HtKf[!�>��?����?�,O�ԋg �I�/r�@�!ҝ1m�58��]�;Ċ�ٴ�?�K>).O|Pa+�OL�O+��B$�n��� 	��	��}�޴�?)����;$��`�O�r�'��4j�\��IAT_$aj�DYf��hF���?Y���?!�H�<+��?٫e��v�:!ڦ	JH�����vӢʓj�D�Ӿi���'�2�O���Ӻ��퀝/%4�nJ3޼�㵁���Ɵ�K�N1?!(O��>�p�#Un��� ����Q�2�c�y{�
��!�I�H���?a!�Ob˓��	�`��<����f�$���i��(h�'���'�����O2(@�o� W�zh��5l�Ԩ�LCŦ��I͟x��(Hݖ���Ozʓ�?��'G28��@���U��oJ�Zaش�?�.OT
G<O��˟<���<ؖM��6H�Qo�p�݊�ɧ�M������S�P�'@�\�TZ�wI���L��%�wɂ6-�1m���ɗH|�x������֟���Gy@�P��0�&�kV�y��GCDhUƫ>+OD�Į<��?��
���0���9�td��� Y��<���?��?q���D(6I���g�? 6u�������7]Ntv)��iV�I�<�'W��'��/�.�yB��4�P0��
�=�L��lHv��6M�O.���O��ĸ<i�J�
<��S�֘�
m���Tn�6!��	����7��O0��?Q���?�#���<�,��v� �E:���i	�Y|�m��e���M����?	-O�t�F�b���'r�O�p@e�$��4� "Kj<���>9��?Y��X�.d���	�Oz��!l����抟��	���A�v�7ͺ<!�,�g���'���'��d��>��*ll���3)�5y2A�}U*�m���I'Wx���e�	w�'�0I�ER�d�y"�Y y>dm�&;��ٴ�?1��?���_0��sy"�I<k���Q�#�M����{k�6��y���O�ʓ��OR2	�w��r�E�	��͂���6��O��Ob+�AP}rX�@��G?i�K��F$:d��e��a���j�"�㦁'�̺��o��'�?���?��[&&�ղ#JO��	��U�m���'���`ƴ>�.O����<���sw�	�93�D�֨�t��zC���!���h��(�Iݟ��ǟ(�'�,��%EN5I��)��H0����@Ȃ�\��꓄��Or��?���?I��(;<(0�#@&S�8 aC֊0��0Γ�?!��?a���?q,O�)��"�|�BAҊW��|����y�⨸���i�'|"V�l�Iԟ����E�	���� R�ޛb8�Th�`,xQ��ܴ�?���?����ؿ-Q�9�O�"Hz�v�2�J�tc̴����B6M�Ot˓�?Q���?����<�I�x��L]:j���y��x��a��n�,�D�O�˓Nz�2�^?��	�L��7u�41��g�[���*D��%�X�r�O��O��dW���|Γ��4�ŞCL�1�L<�z����M�+O@	��kB�Y��ܟ��	�?��O뮕#�����Ş:`\@eJ�✘3;�v�'��Y��y�V����pܧz�
%�C�kO�q$>钽lڗ}r�dX�4�?���?���pH�	ly�+Y�%�N�7�E�UaDP)`��>�@6M�����O����O�r픢y���ʗE9fi�
A6�O����O̽y� B}�U���j?9��G�}�:�s�޿mp@�d#�����Gy����yʟ����Ox�Ӡ'[:T
��@�ԡQ�L �7M�OШi HCz}bP�$�IByr�5V�K�n杸�m�EP������Үh+�d�O���Ot�D�O$ʓ$'���A)b����
F�^B<4���ԍa��	ry��'��I�������X"��!-�J$*��G	KjFi�a�#i���?���?Y���D�zn�D�'eEX0��
Ϸa"j�J�l�`��}mIyB�'��Iɟ��I՟p���x��؄*tv<�ĈP���(:��O��6��Od��O��$�<�˚	3w�S���q�:���Q$ȝh�H���(��M�Ȧ��'j��'T���y>y��4+��@k�e�,7�Z���KDϦ��	͟��'�,��o�~J��?��'К$��ܶR��!�Gz`�tQ����ϟ��I6����D�?�Ib�ِb���V��B �8( N`ӎ��@2ַi���'���O>��Ӻ3�i��D���c&n�\��]����	��d2�h������(��ZM>�X���S�4@��쑵fX�7�[�.
��n�� �I֟P��!���<��)C�_�D YFL��
�����&y]��n\��y2�|��i�OΩ�j��cp,(cFC1ö$��RѦ���ǟL�ɤ9�b�1�O,��?��'49�㫍�=��L��i��,���4�?�-O��a%?O��ڟd���<�3d�$�� �0��v;8|�b	[�M�@*�u��^���'�RX���i����W�l�)��
޶�~P���>馅��<���?���?!���䉣:��S�[-}3��`�X�6w�$�s��`}BT�T��gyR�'�B�'��3n�E����ڂ0>���C��y��'�B�'d��'�剷m��p��O	0X� Y�U�`�bA��5�ZT޴��$�O��?���?	�)��<�T���Oz��zCĝ�xu��O����'UB�'��Y�<��n7����Okl�;����#L�d����`�ۇ��v�'��	ş���ş|�t�X�O`MX�+B3q��0�C��!Z[<p���i���'z�I�Y�$ȭ�����O��i�..6��`��G����5��0	r9�'6��'��CH��yB�'��n�!'%��Y�P,��-aW�W릡�'ؐ� me����O���P�ԧug]::H5x�5����0���MC��?��.��<i����?�S�G<޼�u��?��8���N':7-�'�2�l�D��ɟd�S���'8ހ��Z�P̪Š����U�=c��~��0 ��O��O��?��	�k��}[b"КK5"��v�\>`��	�4�?Q���?)�h�?D'vB�'��$�,fᥫ̷ ��)3�ǤK��O����2���Ot��O�,��h�G8郄��M�������		�r<zJ<���?�L>��+�	�C�R�H�b��#'����'I��:��'�������ٟ(�'R�q0�$%<��+�5�B8��ϛ�dc�0�	h��4��	�(�ܷ6,6�! ��?����3���t�'kb�'��]��zDnj�OܩQjG5�h4���N;=;B�AK<a����?i��K����#�m� AQ?֦�+Ю�(e�6U����ן ��uyb��u���*H���9+/���"�3X���@���1�IQ�I�4�	=|YT��	\��\	����n]�p�� �Y��!�ݴ�?����
J$�I&>��I�?!�� ��c�T"E�&�Q���-vp���x��'���>{|؟0E����.aC��  N�Gop0�i��I6	�a�4/�������䁇pG�$"P�I&�"��sE�7d��'Ç��y��|��H���X'fK$�q�EV�\T��͍�+ �6��Oj��O��	�X������W�<ʂ5���DwP���i��I���d(����a���n�0q�/Lv�H�C�:�M����?��O���x��'S"�O��M�/^<y1ah�I�)�P�i�'`��&�8�	�OX�$�Oh�r ^�v����Ii���kZ���IY�8	�J<���?�L>�1C���g��K��%Ya�Y�<c���'�F|[��'����I�8�'LjY��͔=Qq@5�f�ǐ<��4��?&Jc�H��M�I�L��J�r=`�n˷0=
ܲ��.`U(��sC�ßl�'�2�'X�]��£������j;�,a0L�=j�U�����?AI>Q���?�a͜	�~����s�<)��g�� Z�ii!c������O@�d�O��%RvH�'���i�X뷉���L�W.M�mo��o�؟&�p��؟��dy���O�$S��!�ڀ�� :rĘ-X��i4"�'>�	�/���O|�����J v
�k��]+/\ycQ��9p��'��'7�T���'i�'��)�,�z��I*�6����U�TQ�L��M� [?9�I�?M�O��X���`�����!g��55�i*�'H�l��'��'|�Sh?��D�=삙�'�Kz:T���U�S����M����?�����g�x�'��e�#L�/C6��ԉݕ)�HYc���Q$�O<�Of�?��	0���S�^#c H�Q̋�9.myߴ�?a��?��뉥Y쉧�4�>с�:�:�e�ܱ*�������=�?A��4�'\2�'����@FK�~l�SQ ��~��(a���Ĝ]+�-%���i�'u�p�Wʱz��8ȡO��FQ�UyN<�����D�O��O�"6�W��anP�ɑɔ�iC�R�R���'� �	u�'��DI�G��#��01�^p:��R�g����'���|����L�'.��u�v>��ȁ8m��m��Y 6�h+ct�˓�?�/O���OX���*v�=/��0c�4�\y�Aڀe��Pn���4������ISy�A]eF�ꧢ?w� �.�N� ��S�-G"���¬<����'��I����Iϟ�YVn&�s�>�ctj��,n����"ض��зi���'剶'���!��0���O����)B�l��P'j�bB�4I�P�'lB�'��)D4�yBV����jңI�M��}Pɓ($��I��@�m�'0�x�%z�z�d�O�����FIקu'�� <d�h�NӺwH���ߵ�M����?a1)��<��X?�	zܧGp�s�*Z<,�Y+��G)k@��mZ�h�T���4�?����?	�'H���Oyh� NZ4u�P�U(ZҞ��7����6MԜ(��O�ʓ��O��D-b��)��DV1X����Peդ0��6m�O����O�,b��OT�$�|���~b���/>������$UL+���W�f#<Y����'���'7��:�A��]ZĜ2P&
/�x��es�0�D�P:�%����8�Iu�ɂB����3��!�7�\�Q��	�2��b���ן�������I�@R�gޮXϐ [�"FO�P��f�YyB�'[R�'v�'ZB�O����m�1� �cԩ5��<�3�i�NP��OV�d�O��$"?�S����ם�cP��y��@�=�ȃ�^�d�O��d"���O���֓���3'�L��㤏% ݲ�2�O(t���?Y���?��O��PC+�	�	�T��醺5<hYf���H�l�ҟ�$����ҟ��6�.���>�x��-�_J Zo�N�P���)b�>�P�J�m�X�'n��OA�N�M�������d���.���y�̆*��W�,��a��4��x���z����/Z2#����c菀'��	��T$�����l ������!V*���U��;`Ԓ��*lŁ�7�UC�e
����,�#�-t�	�u�[�6�01��I��$� �^5K��l�C.��tYg��zȒ�2�� ����C؅Kk��ao�(8$>�����t�����2_w�u�R�ԹB`�j�,��vv�M�G(W
��*�皭l�����V�o�1�Ru�OT�QR�ҽ 2|�y�^/zVj�pE��5�e!�Ç�2�7D�RԘ! �a�Ծ�qyZ�]�G���3��}��Eە��E��M~�KW��?�'�hO�d��H&�h4D-B/8�ȑ"O��Q�!�Im����N����6�����?��' ��6�� X@��-�b]�Y��H�@~~Q[��'��'�b�qݝ�	���ͧ
��iSc�)^��Q����03�����O<��%Z15i�XS.�6#`�w��P<�����4k�QU�ɤO	�=0*�hӴ�!$�I��`�	q�I��T�	w�_�v,�Dg�.`�"�!T��(E�-�ȓWȘ�:��ѵ��5@���X5�<��_�X�'��kᅯ>q� ~�1�L�;ר�17I�/y*����?�6m��?����aA_���TO��CK����i�r1�F.ؽI���K'V.��X
ǓH�ƀ WH���-)E�/�M�1kB3C�i�NAR��4�@�y8��D��O,�D�<!�n®R	ZA���B�~��㥨u���=� �P9�A��T �YK�/�h��COr�n�$h>�3��#Z��!�oU�<���I|y����w����?Y.����O�O�uâY�`��$��`�+Dh!��-�OZ��L�}$37B��j��pPd���ʧ��i�/�	A���`0գ�$�#��F(�ӤM�	fDy��L��H����u�_�|*ݢ��O�0ޕ���>�u��ןt�IR�Ox�B@�=�`�qG-������y2bV�(�� )u�Z�$�-B��;�0<�2�	�7J� ���>2j��	Q!B2|>, R�4�?���?i��w����ɟ��Işt�iޕ���ތ~�!�l�XŸE�'y�{�`Շ�ɖD����!]?.P,D��̈́P7��؋�D!<Ox�`F@�/&�8�L�YCp��1�%扩[Cx���|�㘻*Qp]��ȫgyH�����y��'Trz ؑD�a6�9)������Vq���𜙷E߶T �䑕A\�;�,A!�O�m���O`���O��ğֺ���?1�ON�@�)�%�`�b^�@���:��[�x�͙>b�F�@SEػ0�`{B+D�kɋh<�v�Dl���� i��`�-i��t��	|�����ML�g	@�	u ��c�H�1��"D�<B�獼������%-�f��CB5�	���'3(Ćd�����OB�ҵ-�5&J�J .I+(���7��Ob�W�����O��&��d(��ǃ|PTbǔ �2CZ�&��x2�]���'��("�)��$ �荱|��u��3pXL�Id�	��Bt�L5L��R�l�6_(C�	KЄ8�-�W���YRd�v��C�ɹ�Mc�S�L��+@M]�U�=�S�G|̓f�v�C�i'"�'*�ӣj���	�0ߐ4��J>����Ӭ�p� ��I����3�Wҟ��<�����Z\rd��ߺt��1xS�ɀ��V���Fx��D����ѫCJ�Z'6L;è�'��I�^�F��3�)��X���O��V��1{���:�TC�	)2�}iG��}܆�8"ΘG����D�'��L rb�2]�0��­iO��ْ�>A���?����J������?	���?�;;���a7��6	kz�ӵ�J�N������\�F�\�8z����]�g�	W�N)z��T,E��y�!.D"t��l@&Mݺ k�	�FU��$��|��.  q�@��0o���Z�E�����$�O� ړzPbP(13�� &; *1��C	���J�`-r�*��'2�
a�'>�#=�O+���ݸE�R�6�Fْq���Y�(��
ׂ�,��I��L�I��̰Yw�R�'��D0f����U�ތX�� ��F�>�n(�M*"M���Y&ޔ�P*�Y�'@��s�>_� ��I�.
u���BfĨ �a���4�\i�!Ł����@;l� �Q$���aE�&p�v�e�'LB�Y�8��̀�q|����� 8�ȓA5r�1��V�1�uhƵH����<1��i��\�������M���?�Eևb��dj1I�
A��fY��?���j#:�H���?Y�O�hԋ���Ab��F���ґ�!&&)�px���8	S��T�T"MR����.V�q�pȩQ�5O:Yɲ�'[�'H��/��lH�i �R�B�4��'2��H�a�7���'
�-�4a�
�'�j7��6)��d���Ku��=+Մ�z]1O A������	ß��O���'��C�F�2�����D��V$1��'�"�C��"�T>�o��9HfE�j}���Al6j��Ot�j1�)���}O*�Q�/��]\V(����V��'���p�����O�8<I�O�#��CR)E#LE��'�a$/Q)dM�b	6E���Óv������-kZ�3# �S2��D���Ms���?���f
��B��	��?	��?��Ӽ��DNbZm{ÇԆ=��Ϝ���'z�$��d؜!�o�"gæ *I�Z�n=�=9g�Wtx����G��M�._.rB� W�H̓qF��)�3��د9*p�$/As�1�U��Q�!򤓯"K,��q���F8� ���$M�ɜ�HO>E�!#
X� I���9]��[s�ѣ^� 
������I�|�	��u��'�R=�����2Jm|�#�cR�w%�I���B�!�$)|��Xq��*9w,w�s���P�O�Hq/\�`c�9R�Q�X��U�y�r�'�za�0Τ%	d�fѦA	�U�	��� (l�0m�C4�m�K',y�dw�d�X� �B}:5�i^��'pkU�E�6��uI6�
:���;g�'uB獪d���'6�)�� ��|�яF��dp�-�-SR9#fL�p<!`G�n�~�v$�ŭ�F8�}�#Ƌ�W�����ɶpF��/�D��i�HC�ٖ&1f��P�+>�!򄁩BX�;��U#OD\��'��B�!�d^֦��u�Y�q}
������%T��!�5�I:=o���ݴ�?����I�z����
rꎕ2�`�9��QfV�[5���OF��j�Odc��g~�揭:p�@� ��#���ɩ=d�#<�B���>P��#�q�X��l�dG9�����̊RT"� ��j ��C�\�v�!������PzAK
'�sN�u�r�'��"=��ѶE�pe� &��}�X��×3^���'C��'���ٟm���'�2��yG/әQ*N�I3�s�H\��.�
b�1O�ਲ�'�����T=o��2�ˤc׮<�{�ߪ��<�cm��Թ��0`��-peL�?��'��-P�S�g�	�u�X��!!�lp�fR�R4�C�ɧ.Ŝ<�׭M�W�<A����(E��GP��"|�fCI4�Z)�l~�&��1N4��3FH���?���?��4�N�OT��`>�;ĊאA
�򆪁4�HtQ�d�*Q�C�	)-��0�$ɕ<�j���+I8f��gD3������/&�T�!�͔R8P��Z�?�
��V�r|r`���x��a�`M˶|*�e�ȓ'��wG;]��Y�p��L|���<y��d��Hl��l��T�I<��e�s�ՑZ�ƉA��Q1=^%�I�* `\ڟl�I�|�d����%�b�b�'$��H��T�j��`(�e5O�,9��d��z%Y�$߾3���Å�MJ��x����?J>�wAѻG�P�)� L� �1�b\c�<)�D����CWg��4��� ��u<�0�i�n=k���V�麳�H����(�yON>4��6��O���|a�[��?�A,JM@�� �,� BaM��?��O8�hr�iA1O�3?�A\7;��B�qV\@�L�Y��
��z��?�{�b�$�^U1�B��+����+}Rl���?)��䧛�'�1[��X*L�Gk�mӸL�<�����<�w+�w��b�@<EJ���D	R�Dh��DO4�rIp��qW�h�C��-eB��l���ן(�M�0	����I�������6&�X�(_���H�$`�rh�<�N�}x���j�.6z��P�АqA�81+�	(V��Y7hx�y���)J� T��)�OF���&?���S��>���O��d�=ukRp"$ ��.@��)G6:^B�	�-���3��Y8U��(�CE\�-*"�U����DC�U
����	!+ml-"���O�!�
/t��YFJXDP,����fy!��d�Ƽ넊F;��1e�P�Py�h�#��Q)&�
p0Y�ҽ�yR��-(9�]� b|�ax�@T�y��K=w
��d�Iz�X�b��y�m�9 49�)A4I���B�y���=Ev�	i%�|��6� ��y2e�0ODq�dI
a4iC�ʵ�yB�
N�v���lCM���@��Ű�y��S2��pb�B�8�"ԩ.�yFE"I��l�<�H�!��Pyr%�"&�dh�1�^�hD���V#L�<9��?ݨ�H%(�a"��H�n�E�<�@���G�БQLΤ!�dY���PV�<���7D6�9 D�ɩH�3ǮR�<�7z���w��"%R���y�<�0lL�C&d�2M�Q2 �r�u�<i�)H(]�N�ê���4�J'�s�<!D�Jc��yZ҂͋D�ȡ�/Iq�<��T��L� 7�Ɇ}B�urXH�ȓo\�48d`��*�� X�c$X^u�ȓ)�� �P@֢m4�}a'H�l� ��S�? z��a�PB$�H��×=�pI�1"Od@*����/�P8��Ƃ�t�+"O�P+��ߩ.��Q�S@=t��x%"O0���fY�+�@B@��1�m��"O���w�\?B��c#M�8E��`"O����Ȑ93�Ā����*ӞU� "ObnsS�k0�H���c"OvD��<�T)Cĥ�e���`7"O�꣪�9!>�$��d �dV4<*U"O x���J�t˞Qr�G�8�|���"Of(�t+��VZp��smʣ'���"OBH��b��h�ԫ)�*�i�"O��Q�]]�@�뛎��m0"OZI�7.�!Cht%��.� 9�"O�p�w"9���* ���a"Oxr�B
b�M����n�ʕ"OP��a��1��tha�O'2NT�"O�Qr��EX&�q[��Ŗ	DTYQ�"Of�[���^��m���G?1H��"OޠQ��M6� d2���>V�:�"OJ�
U��|MvM�4@&SzU�"O��� C]�=�F�)�X�~0�#�"O��`�
�)���'��� �>�)�"O�q��/���*`�`�ժM�]!��'~��_���z2�ݲL@��P�'��@i��Y+�>\Q���RlP9�'c�$�&�ӑIP���J�T�"�'�}i!F�0{E�S�ɍm�p݈�'<�9YE�_]T �
  �<�4̓�'R><!�a�8B<0���=j���'�6�d�*�B�����wNU�
�'.ޝࡉ�WC�)`UGI�P��*	�'`J=i�IK*cff����P�y
�'�@��`+Y�}��j����F��	�'� ���\|�U�U�D =�����'�lX8ԁ�J|�)GL3���'� a��@/J���zWjݬ-�z��'���۔b�;����F��O&��!�'*�,
i
��`xѣI�3V� �'y���
���H��F�D�6�`�' �bě�xIL�cӍ
	DZj���'!�PJ�ě�/&�x�⡑
8��q��'/��s%, ��<��.�7�\+�'q�k�+�!;�8���l��6?Z@�	�'.��T�	H���3V�29��	�'W��s���Z��1��:VŊ�	�'�̅ˠ�S?��13ԛ{Q���'���5$NT#���-"�4�	�'�\m�f���;��/ �H	�'u�����x��e�������'b��r-�t��d+���&F�Tp��'� ��i����#�-r�2P��'q
 �W-е{��x��؉eT��r�'D.���j�#]I�@K�(߱��\0�'�h�ـ(B)Q�V(+Q���$	�'���
���|�!�q�а~�Π��'���#�ށH��I��U5s%����'6@�Eb��>�J�a�L����'��K���B�I�B^h���'�I0c�Վy���A#H�A�x�x�',dtQU@H�dP�hى1��m����Q�IXH�"�9�'N�B��D*ݵ2"�T�t�h����Id�D��T�wNp�9v�X �E�Ɂ>ަPx���"}h�!s���ԥOx�a[w�p�)���'�v��Ь�*+ʢ�q�[�k�8t9�y��Z�o�(Ty�n�IMZ���$j�4�0_>� ��b�AW�\8l@�����&�'��1�̇7����#x��EM?+>��JU/C��_�U\�����H.T�0@!�8 ��O�d0%Z?ט�R)�ѵj�9�(ɹ6�^�F@�B��	��U��G�U<�� ��P�v����D�o���Ac�,`����i�~��i�(�~��g4 {��kF.�����r<0�6K̨�0=�W�
��}ۥf�#P��Y��c�w�&�cG��mf0��`׀}��a9a`�
dLC�j3I�ay���i2Q*�+7m@䵪�l�*��'H���l�(ј\�B(�2:�q� HF�:6����7��裔dԒXY��9!��4U�P�80A�\(<��P�CN����Ԍ��9��zd䁨N���
�I՘:B����H�#�������|�%���ۂ�͚HV��
,V.��p����!�*NH�1�J;��)���O��Qf�M+�0�������1��(FX�q7K9Xs�(�ř�$Ɔ�<`�ѐ1��z���`�%LOx��EN�v�dpR*�v�|#FN�C��؃qc?=ۘ]���$@9�x����5��'�ax�̇-����z��p�L}�<)��q�+��Z�6���)��h4�t��&f>D+�iڬC�(���d��L�m�QZl�����x�A@��%'Һr�� z����9
�BpgO�4� �)���W�ji:�Y; ?�$J�ø������yW�V�l#�4��g�j��X���yB'ݯO5�m���dȲ0�W�a<Bݻַ��٣���]:<��o �07.�j2-��x��%�2?y� 
4�:d�p��u�(I���z��D�Q�ǚ$�y�
ͻF���N]�M ������.�a�CZ!:l���*��1�:����6e�ӭ@R�)�冞W4T�&��+�햾�T��`�F:� ->�Ӭw��,��Տk����K���VC�I�6�� (U2Q���'�gF�bTa�N R$��p�8bun4�|��U�J��6�HWkX��$��!�R��x%j�YҠ�!o��(�2��G<)�i�!�<QrF��6&3O��1/;&� hHq�C�~P�y�'l����)ՙO��@��A 6�j͑4Ã���?:�Ԉ5d8	�<C�I ?֊��K�.V���ː�[}�O�9RC�{7�Y	��J3`pH���:�)U7n��c�]�4Ti�OmV�C�ɗ!5*<�f"��+y.A� �]t|V��-��踖���M�v��n���$ '/i �C&��Er�L�A���7<!�DY6"�����瓴P�P���kԠ:)�d!��~���AJ/�RȆ�	���K I��FYnD�&�~���N�l�"yK��+�(�� GI�
��L0aC�<K;�!�N�fO�4�Tb�d�S��?1sǌ0�2�#�&O�IB��z��T̓	���x��4s��	�u"3ʧ{�(�DN\8,Hv�91D�- u� dĄ��l7�O�p���
8�\Y��[��,�s/=a��7ƅ��~�mɼ��O-����g?Q��<x���y��sJL�F�E�<Q��ԀpC��q��� { �-R8P��Ġ0���s���@� �Q ��?��'#�<%���G�?*DjE��A�%��	._y~���	[�D{��I���C�>/�tJ��ñ&��%�i�H�����_��y�D�X�@m�Cjգ3�|Sc�?���Ċ���(�:?�|����M���d!F +j>0I`��~ݪɘ�D��y���4�֨��Ƀ^Ɲ;�fڠC�A��E
�eD=��m̙�H4L�O���UN$�g?Q�ڍHΪ�"�`�� 'D��#�N<Q��-P���#��ch�(�GD�ި����O�"�:��2<�D����?���ޟ�d��χ��QpҠ�`�n�[��'�Dt�����F�X�r�Κ5�2�۳@ǅo�r�k .ʮF)�D��F��?�b%�[}R.Z/P���[��2�|��Y�b:i�l@7CN����$��$Ƞ.��) �	J�8�Q�Pm�J?�	�dv�KeN��44�3-3AYzQ�EnW�f4ȉE�'2�A4�����K9�&�� (C;��>��w-���2�ę��!q���Z �DJ�^pY�j\�����gL�h����r��$.�hq��#��O�`ֆڥj�I����"O���!
9o�:��"Ł
���1A'=0.�⟄���92^�tx�M�!Y�(LAg�>}�I�T���f��)#o�t�ai�<��D��w'��;�E��s�`PG*�dEQ��b`�˄8@�`���X@�F��M��A�U�6Š�5��Q�&0ZM<Q���W� �fcG&;0�ѷ#O�~�[��|�FX;_t��Vχ=6��T�3k�s섒O�t��k'�ėv!����eOA�]^�h�T6O��(��#أm��z���e���
�`� E�~U���؋[s�ѣq��)A��fI�9_B�'���b�O^ݘg����Mo�̦);�CؑW
t뵡��/���"�f��;����{���=KFXMS��H�M�]�ѧ��)< ��)Κ=~8(y�'ٶG�X��'����썿$[�`qN�D�2t���$N�s�|�I�F�,\���%�
=f�9s�G�T������*�b��ף	�tR�oоQ�vU�"J+/�p<ؕ�[}�	�S�? <)�#�:C�PАN�i1 ��#�OxyVė��ZP#�&w�h�W��o����v�����M�eZ�x�募k�"�h%�!m�������]5�kǦ�,��O���b��vv��s��"2�Ƀa@�
80ZpAŝH�6�RV;0Z�����U��86�%YV+n���1�ϦJ�'�Bلd<�!�)�^�d��.O�x�0� �$Tz�NK'���R2��?(h20� m�����$@S��$�	ڦ!s��˩m̨I 0m�h�"��e�O��<�C'
%vG��2�b�5Y"!�f ���Q`sl_��">��k@& ��I(d�I�um�vMl���Ú=�JŃFN�W6�k���O:�ۗ��?O��OI�T�ʡL�((�C�]�z�\4x�d��GP<F�t@J�b��Ib�hخU�%s�CNt��T����v���SMO��C��_u8�\�C
�
Dﴙk�
.��\�i÷<�p��>��O���b�H˺�qv)\�IW⑀���t���p6&�0 XD��!R~,�0�`��B��F��R�Ӄ/J�h̓*l�)�ɝ�jU><��̛�pu`��Ʈ��>��$��r`> k��U�Ml�Y(p�;D�$A����Zs�Y:b4����LD2T��*�授uך�!F�	JD�>%�̩�,�]�^���m�����/D��:� 3�ٹD��.o�	{�
,D��0�O1%\��`q#�-�l�P�E6D���#)�6$,�9��O��1Dpd�2�7D�L��o�l8"�ȃDܙ
d��3a5D� k�Ǝ7X�)�	ۚ=W*4��&D����a5�f��䋗SU<S�7D�@Y&"�`mJ1;ǉ�#4>T�8D�ԋ��� ��{�ʗ�^� ��m4D�����!m��Y�I�j����?D���À�#F4s���;�����->D��+"&	J3<�EӬof���B0D�<�O�x�LI� *�g:��Y�.D���#ĿS 4!�ņ�/]�ij�+D�X�u�G��%�UA� A͆e�)D����H֒>�d���V(Pup�i;D��HCB�R���	A�
��"-*E�-D�tz1�>g|�92�I�j��|;�j+D��a�j
w��zq���u��16
*D��	�D�_�8��U�p@zHg�=D�H�0����K��"Z�Vx��c0D��1��,z��a��@ ������/D� ����i�*`�� <��T�-D���gd��x�t��bŖ�.�t�P�+=D�H�j�ph6(B&�T�;>`�ᇇ;D�p��D�s�j�J��� �"���H:D�pb�jA(zrV4�a�لA��BP4D�<P��Y�`�8�c]�]3��@�<D�`��&S�S��k��(K�~X��5D�(�b#0j�jq(c ݪi�1���4D��C�d�@1��Z8
{Nq�tD=D��{b �$ݕ&�bX��8 l��yBaE"x�b��:&���yҍ�m*�USD��4��Q�N��y�C�'-�qj%�[�0�^�uo��y�D� w�����{*�d1�ȃ�y�a�9h2e��C�^ڨ�餥@��y⊜�]K&���#��jslXX*Y�y���"�:����	.4sdPʰ,���yR�ɥH�jD�Ꙕ:�l����Y��yBȽQ6�1�&$���xG˃�yR��+*AjA����&�<i�&��(�y�߯I��<#f#a{6nH.�y�e��/Y<��,]�����@P��yb 1_�ŀ�$M�$��!9/	��y��V��� ���]�|���+��y̓�~ ��iǗ��Q���y2�D
r|p�R��qC6$�aͷ�y�L.%��S��)us��c�_��y
� `p��"��m`8�bTMZ�"��|Zu"O$e/�qy�]��������"O���C3_ ��O�7U3x0�"O��YG�˼o5ZT�a�|1Ptӳ"O�sA�V��ru�!C�)b�"O-qB4���h��
��"Ol�Z'l�7c�8�H�KI"��� "O��������Pụ�L�$��;�"O�����9*���)�/��u.����"O�!��$_u�H����	.L��s"O�<R��5��`&�F+���aw"OB}z��՚&�r9Г��z���+�"OV�"�V+n�{����l��a�Q"O� �C&���yb,מJ�X9��"O����ű\�HqZ���Wˎ�h�"O1����nk������� `���"O汪6�Ɵ(B����%:�f�k2"O���֋�!��l1%E����@�"Of��QQ)?~�Z�d_/c��d�1"O�	�EHQX �����I��|i�"O��i�D�����r焸<f6!�0"O�`[儉���� T�S_�E��"O�e�JJ��D40�ٯ`E��ʦ"O. �B	��qt��T��87|$�7"O�5�A�Pd����;��&"OT���a�^ז��N���P�"�"O��H�V�T#.������X��DK�"O�X1�EB�vľ�a�kկJ�:h�"O�(q&ąUK�!Ã%\�]A�"O�Q�蟨1h����ML�EN�E�R"O�� �v%���M��(�$Bt"O����ϝj���Ѐ"։zq*���"O�����b���C2�Ţϲ���"O"e��ܦ5UxD�A�
�~��"O�y�A�F�<�f�QR���q��Ę�"OJ,�6�$g�@��0�^O�N%��"OZ��G�7Ű [0C��T`{�"O֭@i�d����O�z�-�!��Ϲz�)�u�]"9�5�&I�H�!�$̎B�v�à'�Zbx�;�Q� �!�;
(]��.�5.+�p���o~!��U	T ����7)��Z6`W!�D� �d��!�&N��d����
=!��	�D0�A!Z-^ނPp�B��d!�י$%5Kr,K8˂�ѐ���7!�P�~H,���9%�f�چ`	J!������#ݒ.ĶUJC!ǳ|�!�Dۋb#�ix��$K���q�٠C�!��%*wxh�qg	�G҄q�"�&tA!��e�C�Ӥ:��AB%J;!��P�r�2�e��a L�q���8=V!�D��, �j��:( ��2��G�G!򄍨AA���&t�$�	��		!���;>���C	 �{}���N�n�!��6nCj���i�'{ iC�MF;(�!�$V�uk��8$ N���(��Y�$��I\����$H��
>
P�@;�B.{f�@AC"Oځ��$�*�Ruk�'@fXA�"OX� ��I2K��)�) �T�>H��"OT�HN�T�,0"�R�iղ%Z6"OX�y��Ѝр�ґ�׺n� <�"Oƌ;��?>XE��A��c�""O�`Q\8��"�
b�PxD�,Km!�d6s�x��A֮�����ǐ�!�� �I�CS@�IK�yZ)��I���vl(�'#.ؘ�) i�PS�`۾^u�Q�ȓe~� ��Gԡ�^9CRH��Wkv�ҵ�i 0�O>y���O�����L� ��ef�=9�^�kw"On�Cs"S;z1�!"Gř�5�:`!��'P2u���p>�g����܋�;-� Ep��w�<��M�SvP0��D�]�.��/Zo�<�F�ΰ_
ԥ6�N�F}�a��E�<Q���1We6l���	��P���A�<ѡbJ6\�wE^
�X̓���U�<W�GG�]��?q0���'Jv�<�6������kQ��8@7��R�r�<��R�B��ej²�d�u��i�<�%	$n}�AS
Y0|�l�ǆ�]�<�f��m@A�I/��E���V�<A"+]0#ڠXq�a�ɺ���O�<����EzFxѳk��`���Y���J���0=�l��fڜMqMLM,�P@��$T����T�o�
y��� �q�'�Fh< ��'`�6�:sH�n;p҅Q{�<��oÐE�M)�N	xHA�c�x�<�ҧڜo7�x��i���X�i���p�<�&�ԦJsH�0si�-���i�qH<q�)2v�6��ec�"�J�q%K��yQ!�V�B�r��c�)XR� 8�i��F!�#�ݺuN��3"��h
;0&!�T[��q�G4�@��FǾ,y!򤚛#`l�D�S/'�Θ"d`Q�H{!��%cFah��M'*�x���{!��.iWZ��iҶ>�^�[�.��q!�D_?j@n�ZpǑ��&	ao�:v!�d�y}:�S�?P��)ca-�#q!��ʟ)���+��{��E�EM��!�D]�7��Y�k�$f~��X��j�!��ɡ-�T��2bZ�ZڼѰ��f�!�d^7�hcl_�3ʹ���X�!�	
���s�5�H8ۃ�S�}�qOf�=%?��+E�!���ꋁd�L��UN+D��X�CL�1(N�(�bH�G�ҸB�K-D�l@�A�"f���a���}���k,D��a lC?}�H@�A�M�9BPv�(D�@ �Eƴ,ǲ�1��dh���<D����l*a��U1ǊZD�z�"=D����K �:�ʱ&�� D=�[0&<D�P��T-��`
�� ���bv��y�
��wir�Qs��Pn��!달�yB�A-eH���C�����`Y�ye֋=��y`�
	�$�n�i�.� �y"�!<v��M�M{�4��/��y�X/i��7GO�K5H�(6IK��y�H�ĥq��I���elٶ�y�˓(��0�$X� Ⱥa�Ƶ�yA��@�@���cC�P� )����yҀ�+u�ba韢@+1�7�N��yr�^�a��R���5=��m��� 7�y�k>+� �CBN�Κ"����y�c���U� )�{��預�9�yϋ �N��C��|l���K��y"�H>+ǂ��,Jr��S�%-�yB��wh�u�g�/F#���S�p=��}�A"���ҩ'=a�5%aZ��y�	���^m�ej_j�,�Ȅ����y��~T&�J�!�'3���C���yRI�7��EV��1@�\�K$Jׯ�y
� �q��N\�H^戁GU�oD�P&"OTEPd퐡_��*�뚇�d`'"Ox�ZAf�'0Mkfd Y���"OH5����9Z/�T�MJ�=��#"O�f`X�+x:�x֫_�d�lp%"Ox	�U�L|$z9GꙄ�(ؑ"O�u����o9�@��ܷ%+re�"OP5Q��N,P�:���r܀u"O*):�I��Uȱc&$h���"O	��Fגl�꽃#C�%���U"OryC�O������hU���"O.�!�O� .ʥ�w(X(~Kz��"O,��1!B��a(�(H,�U"O�ĳ� ��X���p%^�%p|�"O��x�e׉�� "��Z%��"Ot��ʆ	[ыTA�y��G"O�8�OA��([�MR.A��u�"O^ e��6\!��M��v�V���"O@�8f �|�Xx��B�ya܍J"O���fN��~� ��f��PDb`"O1��\�^�;����/�4��"O���P�Ԙ[V��ԉZ�D��a1�"O"�['b��rbXI�g��4�"O�	OB�K���6��8A<D�b"O�4a5'Y-LҬq��7�6D0�"O�cO$�p���!XӘ���"OB�cT��+ J��[7����y(�"O<mh�����&��ǘl��`)2"O� �ҎN��r�ВJ�4A��\�c"Oly�#�2K��@�/�?�x`:�"O��"�@�1�TY�qER%%��8�"O�TX�!П�Č;Rg�d��!�"O@d�FJ<�H}�P���:�t���"Ot��%ʚ`�|`t�ȳ�����"OF(�ł����� &�D�R�"O(}��"4%�q9��_�0pؕy "O��0!��%��%I�P?}]r�p�"OX�j򆈊|HH����.��!"Of�����,-be��&��(��"O�2׈4����U�%f��Y��"O������ ��AEKۗ{!"h*q"O� ��ᛜ2�p��5�� ��Z�"O��cV!"�ƽ�&O�W��|�"O��  �**�R"�2�L=z�"O��+C��X��&�A���"O^$;�;Rxx������C�>8 "O�R��SB�|`�"�T��5Ӧ"O��P�EI�) ��%�U���T"O~�C��M;rr�=�BMćq	�pГ"OJ �*A�;lx@��>�=��9��x$L�Ð�S.0��j@�de�مȓU��!q��X���  8`*H��{r��W��-�.���d�r%��΀İ����Z�2K�Uj��ȓE�PX�V��SxuҶ���w���ȓX���R`G\�z�l��毞/}��1��kVp�Ո�ₔ����]u�=��S�^]����<�� `�(��8�N��ȓ)��;� <p�ݣ��ȇF�hm��+t��9��P�w�)!'a\�)����ȓ
��xh�J�d|� %���>"��� ���6O��q����I�ȓNJ�m��U%�B40�JJ=\����ȓ=��MS��[�T���:m�`��S�? �t	�e�+o��S�eO�2�ш#"O:x{ԥ��]a,�ؖ��z���"O���Q!ӗv�hT��.�B�f��"Op��Dŷ�\(Q��FI��,��"O� �OE$?��@s�ڶ6��Q�"O|l���b$6�H�k�
{B8�t"Ox����R6Y� �����<*_|u�W"O�Yq¨�"LVm��K^0���`"O�5vi� A��<1�
K����	�"Od1��
bY� ���8 ��"O�[QI�*�%it�[�VGfȸ�"O�c��'�H 3��#.�q9�"O�̓2�-g�!b�K<0 ��F"O�	��F;hx�s��l~�J�"O�Љ�o��"��I[�Ꮯ ��r�"O�t3�j�`���Q/+���P�"O@�ӈ��G�� 
u.#W��1�"Oܵ�$ �P�	(� g�L`ؠ"O���΃!%��i#A�Q}<�d"O��b��A�6?��kV5Jp�0X�"O��S�	�Y-���d�bp]�s"O�d8�@[ 5�,Tˣ�P)TB�s"O楐�k��cd��P,��
1�HS�"O*����ˆQ(@(P,ƀnV,�r"On�+$0p:l����H��$�"O��5�M'�px�D(��0"O��C`L�2�zG[)����"O�%9�)綸�Ak��v����"Oe�!�YD��I/q��;�"O�E[ c:; ���Ѳ0���"O`�����Q��2�Gʌj��"O\�H!͋���@Hǈ�6��9"O�1 �߶rN�٠��)�i1"O|�F_���`b��)uZ��"O���Cl�/ /L�4�<[�"t;F"O482& 0|�f$�戝5|9\�(S"Om���}�����H9i5DyRv"Od�R@�@�Nq�X�g�0d#�5"O�Х���%��CW��$.�,��"O�q6��N����F�1nR��3"O��'#N�7O8�!ģ�T�$Y�f"Ozʆ�CK��=BU����"O~�#/["��كQ�P� ���b"O`$%�O,��(�&C�@�p%�b"OY+Q��B�:���[�	��E!�"O&�J�!)"��ц���U����"O�x)�C��8�z�+ʖp^fu��"Orؑ��D�)�
����ƞoP����"O���`ҝ{^��3#L^*/�l]c�"O��Be6V|���"
;�Z=��"Ot��"0����)�j�Lx�"O���WD����Pibʛ�yU,)�"O�Yj7D�#Jb]1�盭+�F8�"O�-Z�ȫn�z��6k��e�P"Op530��*CM���R�,S+u�"O�e;!�Y�i1t�i�'�
P����0"O�uztO�<Q���;|}�"O�=� V�Z�88�&ްu�^�
"O���l^%����FÈ�*�"O0m;/�OV��aW��)&N�C""O:���h�2�x�{b��-PR�3�"O@e���D�Q��u�� �B @�R�"O4c�ّI:,��o�=�u!1"O�YKp$c>v�Tָ<����"O� ,��'��}�� �L����"O(��fĝ� S� �M�)�QD"O��p@��0!r�� KA�n�Е[�"O�i�4FL�����ۏw��T��"Oj� �4�\�Q+Mm@T!�4"O�\0��ݹ�r�s�̘_#�xYU"Of���ٛS�����̈́;
d�"O���0�V�x�U��O�n��#"O�2�e�8N߲�s�W����'�ek��~* �*Da�:�[�'�vUq҈�Yz�;�j�(���'�\U!$�;�@Z�l_13׀$�'��)�c�6)����ݹ(�荐�'9��MM�1% �3�C��%?�u�
�'�h=Z�U�Q���#���z���	�'��+�Ɔ%$5���B	�}�	�'�{bf�8��pYԊ0L�@Y	�'�4q�(��Y��S�X�<~��	�'��5�@�(�&8� 若3d��'����%�bG���L�%3f<��':�R��١/v�B�� 3fr�'{�@�ǡ�:o, �B�Է����'���� @ <M��#�s��`�'|X��(?\�x�#t��u(q��'�h�tl�O^"D �
;k���
�'od�r"!NwH�S��z�ȸ�'�)�P@��	KaG#l�C�'�ȭ�A��'��|��CkVd ��'�0t��CN/Bv�	���iF:q��'$ȩ��
�"c�e���]�BT��',���IS6D��A�'�V*�eS�'��@5���C{zt#WȘ�a�x���'P\\0�R^�ȈsƊα�P�' ��C�F2t�������*��'}���JZ6���Qŏ�	�x	��'�L��5���j�T	���	Hx<
�'��)�C�I��M��a�<T�rU�	�'7�Dxbד3f�1 ����@�2	�'�����\DT�0�J]�
,��'˶��#�:6�L )c��V!�j�'w����O�1V�A���P&*��'�Q:A�(?�P����@�,�'A�lB�F���� �7�&xH>Q,O��?a�I�<�`�I�4�Bs��A8�i� ��z�<-�8��-�-��#�#�t�C剱uP��趤H;J*l� eÒ8?
ԣ=�q�4��*��p�x���̝p�"���2��Y�rHN6�d@�R��T����R��0SC��_��d*��G����#n��ce�V
�HR5�ǌO�م�	A~�剐@���I
-;͘䢣)�	�y��bW~����p8e�"�J(�y�-[!��zr`A�w�x�9r�Ұ�yҋ#ur\� �F�q�e�$(�2�y�ԅ&�. �IЄ|U�������y�jE?_9 -tB�7 ��\aT*C��y�j!$8�q�@H�q�px��(�7�y��Z.[��21�So3Jti4�	.��d*�O�Ūe�1N6n؃�
�B����"O��F�ϕ$��U�s ��l.��A0"O��GO�	\�	�	�<5F�pU"O��R��Ш^�%qPB�*��Aye"O��؇�.y8�l$�*�J���"O~����+jO<�
d�S6����2�'��)� �T0���7In*�h$.�P�&X�S�h���\�?�}��J�<�ڢh�h��%;T�K�<�����B��1A�vsg�I�<A��ԏN�¼�1A]5^ �r��o�<1��ޱNT6��!Η�42��TG�U�<�1�U���@['S�71�5!DQ�<�ф�K�C+��;����c+Bwx��'axM"��L���{�Ӳ1ahl��'���6�L*?h�Y����-:��+	��'�2�z&��)T��H.@{0�	�'���&�f%��ڤ��ʍ��'�2H�W�ٷ_�d��TC��cB��	�'�.$C�n��`1՞WĂ���'�ԩ����apuB��ǝ{'�e��'~.u� �� �L3�,�X��g�<I�.Ƹ:�}���1ԅ/���?9
ӓD2�[CN�.mTl@�ՠj�ņ�Q�z	b2i[:�уn���ȓz�vЛ�(x�H��It���ȓ5,���E�p���
H���9��̲�'�11�cCav��"���C�6F�0��I5�X���V��B@��OL&���*mQ�ȓz/F�jӢ�<�%$\0@�}�ȓ<�<�ه�uX� ����|��}�ȓJG�P�&�
�yb]�w�֎"�*��|��j�&��0j Hs��S��]��_��n�n�$���k�;�x�ȓ(���X�b�$8��cv��D@хȓE���W�F�<8�YV!����Ņ�z֮٢W��#6�����9L�r$�'�a~�IIa�Ԝ�R��w��E K��yB	==�%P�� �n(x1c�A#�y�� ����m�c��xw�^�y�W 2���"/7]�j���/��$,�S�O��1Jp�!>&dZ�lW�Zex͢�'*���Χ;���tꕵ)����'�.�i�P���F�:3�0ljT�|2�'��\;���v�J�BV/K0o�t�"�'������>P� 	�E*48�d�i
�'��X8NU�H�>Y�R�;45�j�'�D)���+[.e��@ͼ/�0�R�'M�@�Zi��)��#P�0���'D �J<)��@��[�(1��'F�}��c� z
9�FA�y��j�'8 K�,�!o�U�0�@%b
���'D��׮
�@΂��$h�[@�a��'�bi0Aǎ(|��z��^]�&a��'���qىy��j���OA9�'A����Sk� D˺t}z��'��·o��i�f�K�K6hYʸh�'�t��Ud��3Q�Q��hG�W��|h
�'�0�����oL~(K���J44 y�'F��E-N]G4�I�I� ��q�'�Ft���]s9�<�t�Y9\�b�'�>�q��U 8�첓 S������'��]�R��7f��0�V� �����'z�h�J�|�0J�e�X��"O�\�c�B8U�t�%�8f"����"Ob}Fx���Ý<H�apb�A(!�D��^T���؈	�ő�cS�W"!�O����!WW��eTÉ I!�Deh��j�C�j�8���I%H��	yyB�|ʟ�+�` 8q�G�-�0j�nV��x��S�? �i@�T>�̠�%m�� ���5"O��w�ʲAj=ë��재�5"O�U��%����B�&M�����"O않�*����%C�Ԇ&+����"O$�	�y�fD䈡r"O4����C0�z�Z�
��<�l(V�'���hy���{RfQ"�����M:MQqɠk>�y)��hV�Q���E�:D�&
�y©̦1^�� ��4��4w���y��ʠd�J(�s��)'r�K7�J��y��:��r�����$1�T�y� ԎU����VĀ��<*u��2�y�F]� ��֌���	Z/ȕ�?a���<�|�O$�rf��(K�@1����q�
�S�"O���#�Ҵ[2qC��;R�!�vO*�����( �ժ^�t(��t�9D���D���9S9�1�&cӀ�[�#D�|�'i�&�ʙ���Yj��yR�-;D��q�O��S^�xPDX���5B�L=D��ŏ��3��Ń�ռL@����Ox�8G��'���c%��!
mstOR0K���"�'�⡐�j?Q��i��NI'F�t�`
��y��
�7}� z��ϯc"`�3d'A4�y⦖"7LZ�ral]��A�C�Ѥ�y�[�,T�|s���M̬�*FNŻ�y�d�z;L]{E�H,=�6P�f��9�y�e� ��8b���duܘ��"����/�S�OD=��e�t�\�e g ��
L>A���)Մ8�(ݪs&�*7�<�؁Y	F|ўT���1�r�!��ı��@jA"��˓�0?��|E�����a�M����]�<	��˭n��t�b��"T�� �c�VY�<�b�(=�,�C�ƙ�i����V�lx���IP�:�n�����d3�]I����|�ȓ`bB���HW�T�y�5g�s|�'��G{��ԥV�QE��ľ_&C#�ң�yr�ʎGc&1�1�����ò+̲�kM>��C�Y!So�B��ʡ IXX,��8t�1�J+"��
�"q&��IN�pKb ��^��l:DB�����?9���䟑2�xI#��T�3�)`h�?:!�$\�p���Y��|_
�6M	$����ݎ=�avH�ms��z��88Ȣ=ɉ��?����H�vhCt��9%�D" ',�	G��p9��)4n���<\̭��"8D�h��MׂJ6��S��E�f�RE8D��H�2p
5q�!������6������Ɉ�7%XD�l���+!��W�>�luZqf�B
���I�j��r�'�xLqt��0)�ֹ�06V9���'�!�D� N���c&�V�Y���%žr��'��'��đ)�����	�w�j��D�˕l B�(�<��I��fa6xHEɲO��B�	L��(���P��a�CG�,	v��#�nq�їo{���+P�"� \�Ɠ<3ލ�����{k���o�	9����'�x��&m�)/Wh��ѤK�>�5��'�B�x��^���U�@hF�7#b�s��d!��倄
X->�6иŪ��V�4-��"O��!Ҿ0�@Ʉ���5z�-��F!�DP�ND�`�Aݷ3Ӻ�	uBC
S!����=�#M�)-�,@��慰|"�O>����.�������m�1!��K���S��(�Ȝ���U�)B����,C�lp�5	Q"O� РrG��DbL�r0��KHb��"O�A#�v���@@G@jUf]� "O  ��D�L��<B����p�$"ON���9 ��P�	���F�7�'��DN�X��$��(J3�f���R ���d=�g?1�)�*�d�Yɞ�]�8!��GAy��'��OQ>Q�0�ҒRL�+��?W\4}b�O=D��uƕ�f:@*RʍXL(�b"K>D�P胎�uP̥Q!'�ҴAy�<D����ƍF]6`b�X�k6|���9D�\��5Ī�����Y�>�Z��<ɋ��S�!��`�c�y~��;"�Q��(C�	 �n���"���Aǋ� �
C�7�~Ԉ�
�)q�T#���5j��B�I�hA&��g+�6�&���ԑB��B�I7�`�Ə�3���b��S�A�JC䉇a�xlꅏY�t��X�Qo��2�C�I�|~�� h��2�Hȡ���M;�ʓ�?����#RM2���AH�T�s��߬B�	�^���0�OطvB�l	�)���C��#MFZ4x ͌$*��E��"L./'x���;�"]�
4��4<z��Z�~�C�I�\54-��E�%v� �Tf�-w!4B䉹/�,���\���)tN�9>@C�4�JX��CUF���棐d@4�O8���<��x���%n:�Y�p%V%{!��O.M���S�7S,�#Z�e^!�Dڛ!�V�	FCE:`�yS㕾UT�}R�����Ȗ2;|�a�'�F��)D��ڃd��t9� .�7s0�B�&D�TA�]����q��E�g�����l!D���T��*s�H+���.x�hi��!D�0R#�B�b@H���A>E�f��S�>D�\�S��+{������|�>���ǽ<����ӄ�m�g�Ѣa�8W
���C�I� }���#Om����=*���d?�S�Oۨͨt*�@���hA��'S�H�C"Oui���+��;#L=�~�2t"OT��AA�:�X �lжbʨ��*O�u�E�K	L�\��@ׁ"Ԛ��L>9���	��Y7�B�T�Al�ǉ�+"�!�D�{�y�A�S>t�`��d(R1v!�dH&򁻢C�#�u�(�?o��)�'�Ԥ �o;����ǘ�t9C
�'�t�sL�A4�u��8 `
�'�rӰ&���S��<tٜ�++O>��2�O(��C���*����n�;�"Ov���� 6x\�`��5-z�"Of	��`!y�D�4f(���"O�p'j����P���ƫ)@���'�ў"~�%��6�^7*��i�0��y"O�*I΅���3�����dɱ�y�b��n��Bq�ö*W4�qnؠ��'�az�)�
3��ZF�݇:���pЭ���yR��0 f½����8kI���yrb}qj]� � �>����A$ܞ�y�o��ky|��D�=�N�#.ѭ�y�S6cqf�J��،3���	�c��y�
~�}@�"�\ل�eO΁�y�n�<>��[�j��fԹ
�.���0>��߮0�蔺�fɩ-�h�c�K\Y�<IZ*c���1�[�>�*��U�<�'�D	7A���vI�!g�~A�c��Q�<q6��   -�5�HxeM�d�'a��  9#Aפu�D�!�X�>��"O�zPG		�T�,�b����"OҤQ�'RQ������w�N�I�"O�];�� s�gQ�u�
%��"O��`lܧD�&x3$�!;�
�R�"Ob��"W='���&D��0��"OV���
͒����;��cf"Oƽ�'ǡ"� �ٷG_΀(U"O����ɝ#��A�DmM���I	�"Oh�z�ǫ-�֘�G�����"OA#R��%y0 '�U�<���'"O�9�B =窕��$L1G�r���"OV�[B���)�*Զ
�`�YT"ORdᶧR������i�b��X"O�bs� DP�����
f^�8 �"O��#�ׄ��:r�P�lJ6���"O�mIC�J<aˮec�+�-/z�0�"OԱ�p%Q�1.�q��U2H&�'V�	�v�i�QAF������=V/~B�I�mm�E!2-�ʬq�D�fFB�I*O������3oy���R�][��B�	4+4��`���M�����
�k�B�ɕ,��UK��Y�<���Q�����B��J����5GU���4ˁ��lB�ɻ\[Fuۂ�<df���o���*��$"�ɯl�Z����MMn�H�m_�%C䉬Q��d�  X6jV�x� H�^�&C��T�9j�ʈ<
���!	��`��B�	��R�YT��U#�e��'�NEtC�I�s�|Rp�Ov� .]�g�,B�	�E0�p��H�j��Ԙ��*��B�I�?��q"!G�3<������0�C�"Vhye��:Z%tD�E�O�,��=AÓ{O�$A�':aط���W��H��[� ����Q�,�-�t��I��a��Te�Uې�H?z1hD3Q���4�2\�ȓQDN|�o�j�\�f�@�JT��)�n���"ء5���FP$|�8��� 0�	��sn��0�',�����Ҷ�I���Eb��6@ӟOԸ���q;�I(�Mk�́U6��ȓ�`�����kI���Fb��i�\�ȓf�\��iڿ$v`k�j�<~=$��ȓ&�<�3��L��8�7�S5L����ȓ'g�f��D�b�h��ٳ6�Y�ȓY�$���E�T�f1�#A�2z��P�ȓ@_M1��ӄJ�P�v�_�!Ͷ���$���)��^*���H@�_JNP��M��@�$��d��ꃏ�7!���\��{w�L+���a�
�5�Y��$�t-��bK.7#��P��VB\8��T.q���V�{�؃F%J�@kjQ�ȓ���Bd�;0�1 ��	53��X�	}����
9�@ɰZb>V��'T���J��y2��!K�['�R�X�j���yb�2���r���u��-(�n��yrۏJ8��4�'qwl0���&�yfU?��Tж[�L��&�P��y��
2z����X	��u �)?�y��$Sv4Y`g/麥K�L]��?1���S�BkS&f!ۦ"I�^���c�D�<��I��[ffr�Y�#�<!��׃�Z�b�?\8ijf��y�<Y7,�>"Ĵ��3�^�L*"�d��x�<� b��!ʎC�akV`	W�C1"O�[�c4>g���/
07Dpz�"O|-B��9�vn��!72�k�Y��F{��韢7#2���HN�&� `��O�|�!��Ɯ����`�G�^%Ȑ���!��]s6xl�����
�f�a��޿e!򤅚t�N��`��q��Hxr%�	#�!�dlo��U��?�^�锣K�E_!��4C"�����Y��Z�|!�d�VAd�T�ˉ,���jd�!�DZWq��`�%A�pA�N�"m!���rg�D*׭��vKF�1t�[ mM!�d['�i9�g�W/ �l�?G7!�d�.9�"�$O�Z*2�"��ث3!�$���z�[2�99,��:��ƥ�!�d�X�8@S��W "�\�b�H>!���?QH������,S�D�6�!�	)����$� O�"c��(Tl!�$�"k�X�-�b~p��cLF�x�!��)��aǓ>��I��F9KH!�D�%��Zo\�]�VXs��
*cM!��P�E/^lX�����5���(@!�	�H�qT��y��|�� �+xt!���)���I6f[+۔!����3{�!�di�R�Q�m�\U���&�ʤ�'"O��B׍w���CG\>g�TԺd"On�ń֬Q7�)H�刃r�z�"Ozy`�W7J~�|��D_g�P� �"O�h%.���~��C��kfLˇ"O2$��'T8�����hc~-q"O�%+H<�̡CV��v��"O��t��N��R����!P�"O.�S�X�Ȉ��
�7�H���"O-zSLؠ<��i�D�/44@p�"O�W�J9Ұ���N�8Y�"O4x�Q��(gWtd�#ȁ��ʕ�'"O<�SWoKi�v�酇��^�ف�'��>O��e�Ǭ$x�LRf�`�
�Q""O��D�6{(h�%�/=��ˑ"O��9�d�'L&M�@�C�em���"O,� ��ĜKe�`�Jq�Є �"O:]�"Õ�u�rb�f��	�B"O��R�i��掹��Uq��s"O2R�V����1`I2B���B�'jR:O�K��)e��5P�H�c$(<3"O%��矄fZ�H�@;F�ͫ�"O`,b3�U3K�
����c�:�"OH�Z%kE�<'N��4@Ҝ����"OP��dQ�� ��-t�8��@"OƐa4HQ*sט,*� �@���*�"O�� *��C}��yjDJ59�"O��y0"�gA<��jʯ}O
�3���e>��Cݱ''*I���D9f�� �.D��Z39_�l��e�ݥ /����-D�,���Ăs��J7���$����+D����ܲH�j�`Wƞ� �v�b
(D�S�D�%�
��ԍ�(�\���9D�P�e��#y�����c���@@D6D��eI*��e��e��UyX��)��O����3�$h8�$�q�T)�.N'4!�DY'H�Y��.I����̝J�!�Rt���Y⮘,CX�Ѐ��S�!�䅦:!� �U,X�!A*=�ө�g�!�������.�,F"(01�瀑N>!�� DyBd�P�f}QW&\�Z�"};��|2�)��Z����X�t�؁P����u��C�I�-�(��I�aa��piB�	LԐ�;��^��#E�X�B䉧@�zt�q,�0�P�r��Ճv�C�	�F��q���PL��KX~��C䉗0��$2���)Xcz�[Q�V�BvC�	.\����_	` |xA�g3<�C�I:g��i�EG���P8�Q���|��C�M�D;PKA�Y&6@��㍸?��B�	�f��`��+<s��@2�I�TB�I116*���D?]���eȧ{�B�Ihk��QA&��E��J��7�vB�	�����D�^�� Ä�x�C�ɟD�^<�4DN��9���|��C�I7^�f��&���,u�	��CSQ��C�	����0!
��3�3Đ�u�nC�I %1�U8#�K/�$%���*:lC�?8b|��!�?�4H2��M=.B�I"jz�7-K�m,��e���B�I�Y�|u���*�(�`�*�]vB䉝	�L� 6�*�����P��B�I�4T@�r�îy�J��cJ�M�B����,0b��
Lt�H�
B�B�I3S�8s�=,J���-�n�zB�	L����׶87(�q���H�B�I�8�
1J�nU�*�1U��$2��C�	�o�,i��G�?2�ū�D���C�>
���	t��v[@�����2c��B�I&1��Ap���@��A�0�	�O9�C䉆J���D�3%	�{�K�>��C�	)q�FVT�dP��f�>j^f�x�'^��)C'H'A� `��K�c�J�c�'.,�h���������Ҍ07l-�'(�Q���J����w�Ǣ)�1�	�'�f�K�_���2ئ�����hO?	c�e�5_��9Q�%.6(�H0FXB�<�4H��7B����n�C���S�~�<��È�5���)�%�	K�Yr��`�<��	�%�����L�=�,m���]�<�de�,��!(�m�8��@D XB�<�֏Y;�����_9f�@t�R|�<yS	�0 ����`���Cօ��$EC�<����l���ID~=�頤fGA�<� �V�p�ta���K�B1�'�{�<!0�_�d31�u��2���Qp�z�<��엧b�̩#" !)��9!��t�<�����)_�p ���$�AV�Bj�<aSKӗ!�R��KBN>b��4��A�<�A����9u/�b�P�W�~y2�)�'G���r�@ڳ<U�ؑ3�"z�i@�'��s�6i���	amH��k�'�DkS�O���$�B��fFz��
�'#nq��/ѕgL6���&@�(C�	"T�U��C�+��G-Y�Rk�B�ɕt_4���o �� 2e�`[�B��=y:�ҥ� %#��X@A�,i����k����פ))��j�^�4�@<D�\PC� <��k&��R+hh$�8D�
�D�Q5�#�V#J�U	:D��7!٣H ]Q�G��FNh����$D��s�G�(]t��ĥ1�@̃�o!D��z�,"&.hV�X��yu�9D���g�F�k�Z��ejӕH���x�c*D�� `���/D]�\Xx�E(�X,��"O����oQ���yZ`�^'-�|A�"O��вf�2m����E���r��"O�3��T�?e6�ɣE��w�h`{b"O����MP,���h�Ѯs��-SG"O<a('*L��:�>�ĕQ"OĴ`Ǡ�?yfTJ�hڌ<�<`�"O^�j1�,��� �č�(��]:p"Ol%��.!j�j�8��Y$(�dY�"O>�D�	�Ot�kܥ��pڡ�ȓ/%�@���	2T
Ԝ���ɴs�����.���GL�Jc��
G鐳	xن����'!H�Q�#7���
���p�<yΕ*yK|M�1��4Nư:3�j�<	���#m����(��걁b��f�<�V������q���bM!��Yc�<1 熓I*��r!�Ů�Zt�_�<�h�1�|eAՋ��t��e3A��s�<y��R����F�@�`V�Kr�<quMS5M�0��)˲z"��@�c�<���!~��7 \,Ql{���[�<���[�y/Jt �)Tz�$�p�X�<a5�X�l�h��	R?��r�`�W�<���O5$�ȧ�P�y`���A�S�<���˨v�cAF�>��J���t�<���F�W��yS��^�E`�]p�<9���6@���30,q�Y��.l�<T��7$Ә9p!R���%3��f�<Qt��R�>����۪�j���2D�l��.�.��y�􌛱L�6#P	/D���w�  s�]!$%�A^Liku,"D��0BN	�AJ�giұ
��Ȃ�+D��u��A�(^�C��(2�?D�(�r�:[N�0��ݘ���(�)D���O$hu:);�+G�|(��'D��s�F�f��T��目<ߘ����%D��৤�$G 
D;Tn"y��ZA�"D� y"ő�a��s��#B[|���;D��Z���<d��X�l1�;D���R+���)�U���q�8D�P�#�ąA����M:�����7D��CQ%
�q[�^�Bz`5ʡ4D�L��ÿQt�9�qȔ9�(��E�0D����.X�3��!�4S��!�EN0D��𐨉*�����O�Kg��� a(D�����תu���[e掸	|t���a+D����U5b53�.̭{�0Xu�'D�@��NC&Ը鶇K��phʥ'*D�p�C�Ğ~㴙�w�݂8RDJ!N(<Op#<9�皒h�Vh��O1YZ<0u��P�<�AΏ�@9��z�/72����#�K�<��\�{���	�&�n5���\J�<��8&�����N���l�'��m�<�ǅ�Z&���2)	�y��j�<�c�PHU���Ɗ<�&-���A�<9- {������4>0-��Dx�t�	l��l$*�
��i�Ժ$�޻V��ȓ �^Y�T�ƾ)�Q���� �X�ȓ7.$K �$p�u�,��;B�I��pa5�����G��BN�C�I��cW��V!E(%ˈ9:��C䉌.f��T�[�e@��aĉ�HښC�Ɉ#y"��0	\z#�fƺP�^C�ɛj{" ��hn�]X �<Up8C�)� DÆ�������3t���{#"O�Zn�;��aS�
N�<n�"Oz�cB��+՜"c�ͧ4+���T"O�	
����<	Y�GC ]!���&"O������r�@T�F�K��1�"O�6�߼5�֘�`��80e���P"O�p	a���VN�a0e�	/�PZ�"O���#��@��p�Â�)��̉�"Opt���'"��
�+�9�%B"O$�)�=`":�@t+\!+��B�"O$h+�K�BM�Yа`Ә��"O(��⭀7��=����}�Z��"O��r�t.�aӄɎ3�� "Ox !��:W�\�V*ܰ�d\٢"O�4y��]2l���"�"�
d�`�e"O2<�qj_�"v�c��G�)[��v"Oz��c�6�m:#�<qP��C�"O��yR��I��7a�,"m�є"OV1q� ^�n���%�K�8y2���"O�h+�bӄyH���l��m�(�"O\�j϶laP�tIݧ} � ��"O�4�!��'�00�T)�a �qC"O]y��Y"x f�� ��"�"O���d'؁}60L�ժ�8'�`�"O�q��W(2~��;cd��� �"OT��/���P	$��'�l��"OE��C�n)�d"r��<@>`�20�|��)�ӣG�~�(�#� p�4���=3YC�ɼ;V.AC��B}�2�X DS%^CC�ɴh�А�7,O4����
�!�B�	�32�h��C&����A��o�B�I��8]q���l\��f"�|RDB�	7���Y��H�.@k�@#%�|B�	�bs�y�¤�G8C�	�"=�p�3)N��2���/g�B�"nz�;�bQ W�V5s �ыo4ZB䉔2d��U�Dnl#eGK�/*8B�\��]����>��AK5`�Vj,B�I�b���ƹ5I��#��8�<C�I4p����e�k�	����x(C�I%'��;�������-`QNC�Icݚ51.K�f�`���
��
B�[́*���;/�̩��ۻ~��C�	�CMؖ΅���D!#nL89'�C�I"{�|�7�
&$U���3�J2�B�ɲ����H�:q��)�W&*�zB�Id?�M��/
����1A�B�$��IQ��1��	�C���
�BD!X��2r� `5�C�I�8�Z�$h�/4g��{��Y��C��6�B�
��]>ɼ Y#���cZ^B䉆;�DI�T/P�=���d&
q�B�	*�B��rJԲb̦�04�@|�C䉦r�����jK �@��1�]Y��B�	�P�B���"g�-�Oƴ�B䉰o�T��dē"�$��6����C��7J�� �V�C���F��(?|B�	�N�H�X��
)��@��@:8&�C�ɛ	�")���1v���j��f'~B� ��@y�@�Mg��"��Q-Y�VB��!,��A�ч��ԑzf���/@RB�	,N��eb5*C���䃀��#%Z�C�	z���a7��d���R4*��C�I+:)�����M�qXtЀ���g��B�)� @�ҐH2L�\(T�ʃi�5�c"O�9p-���(�4�ׄP��"�"O�Y+u�ʒ`���fR�~U�t��"OQ�u+�H��1���r+8|�"O���c)�#K.�Btk��M�����"O������O��(B�]���"O
���T�,��T.w��a�u"Om����'Đ21�
�2��k�"O𱂑�Ȧ��,�w�?T��ћ�"Op} ����|�I"��n����"O��@�2w���՝e�A"OpD�@o�plX���dɕp>�QV"O�*��. ����B�!Z9��c"O�R�g��Z�zUK���,V��"O��!��ҷ:8`�zBOސ�&��E"O��c�M��14|��q�� �H! �"O>��i\R~��Y��H6�� "O�:�ˈ$*}vX�)�9��"O�ę�`�,H90�h�'C�g��ܰ"OR�:Ej���caċ�l�4 q"O"�����1D�l<�@AF�F�B�u"O������*^���Ê�Q�v��p"O�i`�Ȋ������k�.���9�"O(��T醜1��$Z4h�(+����"Oy�O
8����2n�
=���"O��aU�R�e`�ȣLӶ\��څ"Of�:vO�����+�:EڍpA"O�4(*ՈTb��k��"l�8İt*Or�)t�*a�9���Z�lz�'�Ȱj�:�x\Gd_&�}��'N����Ն��M��-�A���`�'h�8�l�b������3�Z�S�'�\TC�.�����yr��2t4,j�'�l,b%۲�T�9Q�Z,2^L�
�'~bݛU���Y��0/r�	�'P�H�A�� �F`	���8,Y���'���c4+��>{PL�`�M�q�Y 	�'E�P8��@�ц�3$�c�<h�'��`�&�z��Mֆ�')�(��'��	s�3.�J���'̝p�'~�M�ⅈ}�rM�1oJ7#,���'�<� 䔞|�x�!���N�Q�'b��	#�n��q@!��N���!�'&
��I��z@.�A��4L�-��'�x�1`G# �,�i2$��y��(�	�'j��U!��6��`(���aް��'�vy���*� �#"��^k }�'�8l2�3�~u��S�g"�P�'�@=A!��<u<x�sf�_!X$¹��':�M�d+\�+�L�i�o
;ߚ��'�� �ѧ�+`~x0�u���6�L��'�n�R�
>`��˅���&�R%�'��x�@h�u�R��,,!e�c�'>�,��B�J[�$ъ�D��Q��'�H�`�?���h����>�A�'횩s�A o�����˞ o$YX�'D0\��-�Nq���ƧG� �����'?\)F��dD�4/.Ά���'yp���N�z�m
�r$���'��E�#ρ���C��Y�W� �'z&(h@���'��Y��.��P��l��'Б+�g�1q����"P� �	�'�E��f_	q�҉�iʓ�ܩ�'��s����a�'��I0����� d�+��E�Y��|+�ق2�eC�"OH���'y=�UӡaȃB��a�1"O�H`^_��с���lǂ���"Op�c D� ʢ��"$�M�f��4"O:œU1h azU,B?�V�Z�"O�@6O�#�*t��Jd��K�"O��ö*L/'����3$�Y��"O@%��\�\�"�(�����q�"O���G�8� $�j]�]����D"O�e��&L._��Mc4�H;8r��E"Oʈr����ޙ��������"O�1['U�bq�c����&��(�"O>!��A�c��m�dC�u.�0#�"Ol��a�L�Q"� H&m�9A���{G"O���2 K�U1�ِ�⌑���zB"O
��_>�ܨ+u⛴vfAp"O�M3 ��re~���F�7UA��³"O^�# C�PچQs��3m&~1�"O��[E�[�0�2�I����0����"O�(�Cիz�2x���}I�"OR8㍝x�$�C̀�RL�A�e"O�e�� _�'Vb�a��y;���"OfI�e��:��<��M�tR"O&���.ą3s��ƞd`TT��;D��*�8pj��H�7u����4D��9��Ҏ5��a�oO+=�y{�B3D����$Q�l0�[�"�!���12F>D�TI�+��@ޔ�CO��I�ܸHB�<D�\��~\^AX%Ce|���e.D����	(,uh����¡^�M�V-.D� õjG8�����J�u�h�pS�>D�d9V��5؄Y���	�/�J��/D��yf(��1&��!䊇�(ZA`��,D�`��D�2� ����h�:�6/%D�Cr��(yz�=��ݦ*��t #D���C4�BDa٘*��k$"D�,�3�XR^����v`����<D���6iM'_�)C4M%sKb��կ:D�x�w��P����m�T��d�7D�p�
H4.E=Q�J+7�<9�A5T�I�A  8��×��J��D{�"Oe�A�J'mg�B�I�rb�x��*O���#K�:l]�dD�<��ͫ�'���Q晈X$���d
}!�9�'��8���
�w>�9d�E8q ~�K�'��Yq��:��|����
b��}C�'J���
�=���e��D0�'�ܩ*tf��|����(�-rbe��'���0΅�jl����\q}�Y�'$�1Ц�s�@93�@˱z����	�'{Z`���	���7Ȋ�zI4�K�'�� ��	�&������݊C� ��'�N��TkX>C�@g�P�5Q~���' ��� �����ET�(8� K�'%r制���Ԝ���	��1	�'�$]Ӄ�A�,YtADr�T��'L�@`n�Lqɢ��	?����'�����,m��2.�>EXr�'&n�p#�Q;'�B9�m3'�Z���'�6`�v+L�-<j�K k�P,�L�'"�"�ڃ:�� �G�U�T0���'���& �24�M!��V�>��
�'M
s`�A�q�����%�쀉
�'�@{'�i����ث'�\[	��� �8!#��VD�J��cj���b"OH�R� B�57���	Du�"E1�"O&<i��تr�4]Rv��8Gy�s"O��
�Z)_���
��ǻ>F `��"O�t9Sou&l�Q�A���9f"O��R��]�^h��������0"O((D�� ��i�իX�t�-��"O2��6�;<p�9S�F�
LX "O����K9 k���@�F't}���"ORT����*M����P	��]P�g"O�	�Rj��qil�#GH��+F�e�"O�P灋#w
���C-��k8�pd"O@�:"l\�,����CFBDiڵ"O����B�a����f�?(@$��"Ox���LX�t5����̚PD*��0"O�4���K�`)`d³��O`4d�$"O�"�� <b�6��ZP�۵&!D��B��Y�p���*ՌN�juصI !D�h��ꖁj���cč"U�ʽi�?D��0��3h��ɑ��#���9tm*D��"�3CF|$����[u �S2�(D��@un����AFd��2�$dxw%;D�<���<x\�U��@�l���+&D���S��1������+�B(r׏%D�xz$"V�4�̽��I�w.���`$D��q���q�e;� ��=�bL�%E"D����re�B.�b��� 
 D���J���
����A�C)\�ZWl?D���#a�Lz쐫Kޙ�8���7D�<�`�č)閈S7�H'I�\��3D�ԩ�⃤0�F]��'
NPNŨ��O�=E��aI7�Xl��@їAU��z5���!򄞘V�,�ӀS��Rf�M�!�Ď�H�@Y�mPXFT};��P�!���&_�T`@��=8�p�S$� �!�d?|��E?5޼@��?o!�D�JQ>p��F�y,d�)��-rP!�I%�^���N��&yZ�J�.E!�V�1Ӯ5�Hݟ#���H#@5!�X*����F���] ����A�0!��ǊNj�Ă�R�` �Ee� ya��O������[�8����^= M:�"O���瓔Y�pY��"�D���"OĽXG�3)�ЭƱ$��I�"O�r�Ԉ53 Ĩ�
R�{oP��"O��	 ���E�C	]�`$�#E�'�Q��3@�����3����q��8!�<?e�'�~�<s�����T�b��Q�w�Is���OK��	���;Ɍ�۲���$��'N<p�!d�����H�B��q~���Ob��D{��/L��A$ץY�В�Ǿ��Ԇ��f^��\�f ����q�n�����39���	@�S��yR�9t8[�Ϸ@&����߆�y�"҃Y�0���	�5�F �!ƅ�y��'s��c�>@�����!Æ�F���'L�IV�$j��"'d�4� ���'Wr4B�A�:;,�}`g�O�3�ƌR��D!���Qpl�n@Dj��=a�P���'}qO�`�����O��ժ�e\�P��"Of�\�0k��-;"�D8�X�2�O��=%>��/V,)�`��+�i���+ �;D�x�C-_"!#�-���J8D��PBLȤh��u�r� �fU~!���7D�H�w�&)ZF���+݊s�&�,a��G{��� 䵡��C4Oмس��?)����1O����2��0��E��M1 ��L���!���S?���" G#j|�-�vK�!�!�DW,*J,���L�8*U��	$h!�ĝ2�AӪΚ1^�b�\+*��}r���`�ϸ<6�PƆL��&�i5D��@��ݞg�ʵc���U�����2D��{��ß>��X�m�
��l0D�|��HF�2O�ݳ�(��S�>,��j���{B�)�'�\t+�b�K3<Xi�փe.x�ȓ� �����8=hا�Z&�ܦO�К	�0ƕ����;S���A�DI�.�����<��ς:Ɉ]s7)��>����kM�<1��C�ww�h ��-{�(t� � F~�'YL(R蜉(��r�Ŝ^Y�l�ȓq���ܙ.tV<��	/rv�ȓIԠICp-�r`>BT �J�I�ȓ	Ȭ�8p�_�B�^�a'g3uK�х�Iy~b���ɂ����&����UOح�y��)�Sg}R�]�N�|��+�,�5KJ��y�b�4pt-�g�	#�A��yr�74qp��}0�������p<��D�zB!� 'M!\��,�wC�/>���ȓHB�k�mZ�}]�%j$���.�"��O<�c���i�',���0jS~�eY�i+s!�^�_ P1��i��p��f	(���՗xRW��>O��KGmx�cei]vR�)�"O8=zJN$�Z��P��-Xb����O���d�%I��@�F��;B%�V��{��`~2'W�f��$O�8�>�r�-�:7*�C�2�h���/K0{w�aVdȩs����M1a��"� P�&�A#��@��I�`�Φ2�B�(g�� [�_΀�fk_7-��D�D$O 	P�Oh��~҅�:�pӀA�$۞��g����>�U���#&���ԼQ�F�L%�i�pϱ��5"�<)��tGe�+ ��?��Je&(�HO�c� ��t�D�D�l�,Q5P+rd�a���u�v����/�2]e���R"I*q�T�%NL*�hO�O������:m�=h�Z��Z.rnJ8C�U(�x��\��L�%�8˂�b�&���D(�O��Ci��g5H]qe��;>�:e��
O�堔�]'UF%�1eI!Za
8��HO����á,H��n����1$�:V��x��	��� �!�z�3+�l,B�ɗ>GNd��ꌹXLV 8���0���'��I}�)�S�G��\�����RB�H�X#�"O�y�E��QQ�԰'�X/E ����J����2KI8�P;�i�<n��ݸ���y�з3��j��j;HY�>�yBd�3:��,�u�=�=AD����x�	I�1��HS�1<x[V��nI`B䉔^K��@�E����:!ɍ�&�C�	
sqn� M[
�����g�5L�B�I:c�̋Wj�p���=x��B�Iΰ5B!��q�JyÐG8�tB�I�k;J�*�����-{�Mc#�C�	G�6�p��oʍ�d�ZbRfC�	j����df�̲�l��"-VC�I�2�� ��ψ�rr������pB�I�]��d�g�n0i4F%	��B�	#Y����F2[��sa�ޑY�2B�I�~���Y��R�.Х[OR�KG,B�ɺD��㤌E�Q��Ez�*��{��C�	�UB%��-4y��4�N;&�XB�)� 
�xB�P�Q�,����?<^�!)�"O��/\�J�j�ë?3d���"O�8a������Fȇ�bL��'��	�_�4�+��@�̨�F$�G����ĸ<�@KM!H6�if��a����0��O��~��^$��q �. @x������+D�����F�����ʚA��QJš6OlQ���'?�>�g���~튐�FNpa[uAE�<�Ё�(G�k���,�h��Y}�d�)��'w>Q���d�M�0)�1e�P���<D�l��FDy� 
�%{�|���*<��j�t7m0�D�?馟~�h���k+�q�W$�Y�!ɳ"O�����5+�1�sADw=ޔ���|r"U���Oq��1��<�
��k�;dd��}r�)�I53���W�I{J�Y��C�.�!��\��l�q��/l�I:s�ay��ɣ5B�)9C���X��eRĉ�/�"C�ɰ�J�p��!J��9 ���9a�&�	6�HO��=ɳF����Ip�C6{�@d2�K
F8��&�4�$e�D	"�Ǐ\�ٺ�˒�kӈM������$Bc� �4�7�E"� A��">�����y\��ȕb77�J��f@G�bT�ɴG�}2L�9G�X!B˓.So�u��F��HOĢ=�O� Ir4��i���x�H:��(q�|�$��	�3@�5I��G9����� :��b�IV̓�McL|B�)6�h�'�[��xh���d�'���FyʟX� �5��PѤ��-��"O�U��#�0W|�0'dE�~�
���'�1OH	�&�Ѫ|���h�E(E�E�b9D�@Q���*D��`�F0~�~Aq@nv���b%H�'�����V� z�1 �(| -pl:D��Q7IW��is���3�%�U:D� +���)xJ��6�L�;�,0q��9D��*+(f���H�*�(�3��+�O��(.F.�pp����<�6����'������.!��XA��Ȍs��+D�H�k��X��B�%��j�!�9CR����N��D�hg.�+;�!�ā&P�ܵr$K6;$:�x%n�|�!���4Ǣ�6B
-@&��NԴr�!��f����燏�Q&�ݨ׋A� �!�$�<�ܕys�ɤ}�:9U@��!�DF2aȒ���eJ�v��*��X�|�!�$.����#u��kt�j !�u�ԫ4��E��	����,p<!��
}��D�-�B,ڰ�Նl�!��9ix����B�v�$�Y�!��=R:�%"%�ў-���N,M�!�D�6�h�x.ށ#����T��g�!�J���y#ÉN�[�^�j
�5�!�D�+P�0���훌6�d�T�!�$���ܼzf�,2$9c���t�!�DҐ�\���*мt�d�ib	z�!�DB�+	N8S$fQ�&y�Y`Aʚ�:p!�T�c�T���
�S��y�(˙c!����i�L���©u@��gU`!�&x��B�yN�(#����F!�N�{Rd@�qm�6~:*-(B��|E!�^�V��5��6I%���W�&!��+!)d�j��fI��K\�\`0��'��x��V�c�V�)p�ŀ~m�'��SF��T�D�`)��Z��'y��P��1V��`u�T%8&�d��'��A
�q}J��4m� *����� 
icҁIw�h��B�P�O�R�Sa"O���R--�Ub�˔�*3���s"O��$c�?0���J�Ș=,�Y3�"O`��ԦJ�x��e�1�=]*&ЛV"O`�ІOɺ�����h��m<�J�"O�I��!�A��+�	@�{P�R"O܁o�	
�(Lp��V1c���C�"O�(�%���:$�$�\>��XC�"O��2S'N�_�.����6S}R$�"O �R�	ԘU�b(ŀZK^�X�"O�� ��ذ*�iw�W<K���"O�Eo~3r0akɏRfh �s"3D������3$l)P�
5x�="��7D��`�j�`�8y�]4'{���di3D�<��%ְ?�`=�R)��i)��&/D������@�@��ƧO�s�x��*D��""\�L��������N<2-(��+D�Pp�L� /�L����5\��M*D� ��(��<�x]2���q44�Q+D�l0���z\�A9 �	��a���=D�x��"9�깁�={��0&�,D���4�N�hF=�E$A�>-���*D�0lĭ�|@
��Z�ղ�#�*D���`Lůgz8��bj�;@��A%"D���YmN�Mq�mDj�Q� >D��� �;����	B�0g�\;�).D�|kPD@*J��a���LJIaP�,D�@!G�!��j]�%�Tի� -D��#�B$����G��Z���>D�hc�%:�V�{ֈ�4O����@l?D����ND	��D�������` �=D��iQ��bδ�`肘=9�l�� :D�\���� )��i���aVLxC	8D��eNz;�"�2H�j�9D�$��M� [7B�+�kܼMȥ��`5D����"]��)�b'�][
1ڗ�5D��)�8_����-��I��3D�$ӓ��a0� �w�� �J�2D��K��_�*o�]
�f�2l�i�=D�8 G�۹"_mH����a^���@ 9D��:��a�p�a��R8l��W@%D�<��Q�.qkGl��`�{�%D���l�	`�~���Ɍ�8�Di�wH%D�l2�,�rD���	O�akD  D��R0�F���`稅7�#8D�hzT)�E�*=`����|���7D��`��V�4�B�	�1k�P���7D�,R�%G�3�d�����8�(���2D�D�4>��"�j�E��	)�h4D��P�7td�FL�(nX�e�)$D���h"/\���JQ�q�r�1D��z��F�<�2� ��0(麝��#;D�wI  d��PG��#��%�4D�TC�o�1c�9]Iȉ���5D�L����i��̈wmz1b�iC�yR+�.L|C����z�����)P�yr�,r�<=�"�[�M�P����?�L��?��>���V2Z=r��P�Lx^<D� B�<`�T�b���$)N�C��X�o�F�i��t��(�<<Q�T���!Şm�U�=\OB<�r,�0�����9p�Jslʸ
*|�+�3A�!��Y%B^���t@� )�R�t���{R��+u1PІ�>�1���V Ȓ"ԗ>\JC��6�V�A�ƻ[��9D���B>�4Y���� �ħZ�� )L�� ^�:�dX�e��}ȀHU�&n��"O��h���#�D+�`�	K�����I�����OH�`ĭ����9hp��ժ��uj�Y���ͦ��ɲJ۶��OZ����8�8��j�UN���x�qO�hY��Y�<!�a��i��ICQ����q�%9D����'
B��2���ܤY3�Y��@�P�;�O��4@J�.P ��
 ](
pe�'ö���J~�j�y6��	��+vvZ�i�,��yW�l�
�@$
�5'Y�\Eŕ���'g$�����O>�pH^6JD�LR�oS)�`MJ�/'D���#s��!�䂸�Afd�o;�O� E��O4̫����Z�G�DE�.�9�"O<�Q�ʞ�Sς�5B���4�Q �'���3��iX�$��b�P�Lq�	��uR�6ʓ�n-�B��<q�dL	@�<!`E;��Mu�-"$�ه�Վ�*�h�"OZq��A��aJ1i�'>�D��a���*���@){�$I����U8��"����yw@	
%®�!�f��[A4R�\��y"O��;,��p��풥�oi��nٜ�z(Q�($hř���?�qQ-G�t�`��@�N�x���I@�$4�(�,0|OYrc� ��I�2hb`��ؤt��
�l�"QH=�v�V�-H�Uzό!Q��zʐkm`5�s�ߝ-�J�QR�۲��'H`a��ui��斂9��Ⴌ�!��5D��k�MQ�	��4Y���!�D��r�'�n}K��J�O���g�9��	�V���$m�uJ1Г�X�$�~a{�`���䧡yw�T�2@�fL�ߚyQSa�-�yr޺22Ȍ�̂>'�y�2�Wv���c�CM�J�>������)ipe(��37Ƥ�dL�-�'�x���M:���Z�gJ3#�F�Bߓx�c�+E�w�D�	�&1Ψ�R�N�y#>�����j��MBS/��`�WBn��y��Q���`T�.���5d���'>v��%�mJ�CP*/T_��[$��P���v!T�R,Z��rf�.E�`�5�^�%����R�
Q�"*�<Y����&�A`��
P�.����Ū��`V�{�@�>T�q��4x��S�Z��N�..����DXG=,����%�!���%���(�+n�p�R���D� z�H���h�,9D�����?/���'hT�l�d�O~	#F锑sq�4yw(�:=��B��'I�1�nF0�����l&)a"���5'	,TBF@�;Zr\���H�i+2�C'g|<��[�N,9�o�|J��BV�[�BG^��=��홣&(F�
&�I3z�`�k�$��В=rr�,c$��z�MY.d+ �l�n��S�nh<�g�òs�P��M�52Fh���Jy!2$;7�::�qcD��_済��bC3q�V����Mq�w�<����	4ݠe��>A����'ԈY���2Mtи�I�;2'b���r�8�'M
H��C���uGe"��N͊Ș'׸�E��U�<҃��7��� 
��x5�t��ך� Pk���#��0���aSx����cSl�%&
���ɒqB�Xs��T�|D�e�X�	�>)A��3�Bq�nǥXц� ���pB���@�V� ����C@�̚��=D�4��BԑL�L�۶��8��u(��l��_�(.�1���/A�ep�f�O�NX@�CF	t���"�/`�f��y�T m�jh`E&LH��AH	�F�F Vv)I "D�"���L?�Xj�$�6g%��2���P܊(3�*�O�]��d	�:����拰=O�!�5AÖ_ڴ����j����'�Q�է
}UƅS@���T��I���dן+�]���ň>���ܕU;��XE-ԟ�y�e�S��I�cM BM2������y�nʱ-?bIRj;2�<��R�
��y��ƽA�l�[ �U��p�����y�A�.T��=t�Q�`�n���g��y�+w=V 4��g" u��H�yr%Rbh�8���ǤeH��p4	��y�V*N��0!���,/��� cO���y�bٕ�����"&���3/�y����3gM�`,�A�͢n����'V̕�����K�fi�)ڸ
�( �
��MWb˲T\h��aj��K�',�����MX<�t��/,���	�'�L��Q�լf�|J�MP�>����'
f�Z0&Q�@}�%&2J��`�'�^�R��P�� 2!��]�
B*��UfN�kT����'r^M��e�	E����*o=��a�N55)�=���;�Pxr*7��@Xq���"�$����� l��Ş-�'7��s�ı2V�O�'v²-k�	0I���p��)wl���	�6H�]:%n�)3$H�'���K�J��.�T�a���)��� �N�a��H�b�(}��\J��҆q��a��J5V��B��<1��ߍC1&�`QK���" B�<4�,���=�@�*���k.�g�����'d�;��W����c�=<����ٲP�z��Y��i�1/�B̧[��Y��oO�0ƛfN�	s�����Y� ��JU�ϋ��?�7��$T�G�@�3�����.VxY0��ÇzX� ������S���?�뢐>���R#F"1�Ͷ4y�<�����N�(�Ō1�����T?}���{�J��&
�`���vmۖk�T���iԹ��Iv��~¡�$.�,1�Ð�9�倢�X�򄈏@��h�6��1eRd����H,=��a3�
�v�r�dC�2 b�[7�̈1Gk؞(SV-}����F���?@��"H0`}\���'���Ab-��D�O���a2�ՒF�����7�pר�~�����5�򡀖0T����G�KpR�X���VG�)0򠅮h�p�TgIy��H�����=�O@1۱�A� `+�u3�uN��@�z�Tq,O�%R �L:\+6��1��QX��c0"Ot�*��"h���@��X.��`
�(��䞰]�a�d��F���%�=d(65!`jϏ�p=!aO��LO�ҫOD`Q�B��=m&y���40���'o  a1�Z �0ʓ2�͘`�ŦY
�����"^��<��m��\�	
c�:�'&p!����/3���3��:"�ACB�Y�8�	<�vԈs���7!p�S�'0ݾL`E!M�*WĄՂ�k�,Y9�U֐�'�͂U?�9E�2�^��O�qaK�6&=n<IS� ;1�)0��ѝ��a�'a �h)�3}B�H�Nᢁ�ϓ�n���/[/M��,��n��5�,E�v��!)�����>��M4�)�6�8�� ,�P�M<D��1��:�
 �I.�D1�ՃL?A��͓w?��*/]L���OG�5��89���h�䟏+cT�!���� `%E;�jt!�Z�|��(J�X���I,sD���%0��	�p\��Q�Q��|���(���wē�qG& B��P7���-ܒB87���G"D0����V �)�SH��u��/��-n|����n9�����;���GǴ� �Os��t%L�*�*0�'G��Y���|���㷯�bK��@ dZGx�'ǜ,1����$z1N�-����AG9	��X"�S������pv��@-�&g�:-�O��2��4��L�n%�F�NNX�t�Y8)�:��Tn��hO��Y� _Q>�J6nj�$�ӆ�*���2���.%�t�MS9i,�'_B����d�g�
I^�!̎:�P�*��qtc��:����sq�Ё�S�%*���DV+-�6��i��6P���#^:/Ih���'�J�p��x�0�`�'p��!e�V�"�O�)	������D�":�'��a��9|Z��B3s�>A��'��p��ݒmQ��a�aօ0%��YM>i�!V�1'���>	���G�<Q�T��wx�h���$D��"��� $�<%���vJ��ej D������\���c��?(J}��<D�<Y��8O�t���8J�H�ѷ'8D�d	͔%<�6�iԉ�/
�|���3D��0�c���@��Q��>�����1D��+"�2['���� GK^�Y��-D�ܹ�O�o#Virf�G1p ���&�*D�H�g�XV�o���i9dM&D�P��I�/h�$ٖ��9��RTh0D�Ƞ�Mk>)0���V{ʸ���/D�Y���G���guBY;'�!D��1��	$<J�I��L{F9��>D��u.�#���3�tI���N8D�Z���g��A�틷A{����9D�؊#�G,^��uA�o�9�|�вB3D�@�s��.����Ac2#V�m�t;D�V�C�{����@�*F���"�6D�|�ԓk<�!�Q�G�a �]i$�8D��8!��,<;pe ��«s���7D���Q���&Ӹl(`+Ļy���;'7D��&-H�L�ꇁC�X�PV�;D����3:r~����Ě}C���dD8D�� ������9Iml�h��S*'E��D"OJ�xȧ#貔a�
k�0��"Ozh�M��w}+��N�R����"O��bp���{���C�&L��0�K0"O^%2� ���d�
";E9ɵ"O�}c�)bU��k�^�T���"O�M�&W#>Y�8r�%@��:P�"O�@:/L?l�0Ջ@�6�2��p"O��[3ʑ>W*�h�e��>@��}�"O��0��-OZvdI�"V�'�D-r"O:����ɃEm��d#;���Q"O�q[�c	a�p�%,M�@T"OH����8%#ZԲ)ʂcN���"Ol`;�hV~��B�	-��C�"O��Z�F�"�TYd�M*R(4�g"O�(�璘q���"S�Z�x�� R�"O���W	�� ��1i���%�NDR�"O�h���ܥ����C��`��IQ�"OJ����H=X�4�EC��|@i!"O��br#h�&�j��A�����"Or4z��Ju�,�*3�Η,�@���"OX���'��i����$�I�Z�(��0"Oz�JE.�5��nA��*���"O�=�3��?I�X�÷ظZH��Ig"O��c�)�&j�R[�1��`�"O0	c��D8A�z�hEMT?�����"O���B?�� ӅF�Va0s`"O���0���9�6I���0Z�x"O�x��"�/r��dP�K�u���"�"Oδ��㖩'�:i��G2 x��U"O8�ۀ�R.L����XWV���"Om2�
Q�-������O�&8X�sU"O
����\�v��41���<1�H��e"O@�U��Q�D)hu�߾['P��"O̼s��X?�����U�:}�"OtؕK p��	30Y�p�*}�"O�� "�_�P��$r7�#=�¥��"O`�v����#'nW�-�>=4#.D�ȡ��V ��3y�0�@�-D� c��1<pRE�!�	~�*�!,*D�08s�(��ȫ�@�-T"h�*O��ˁ��*���u�$ɲ"O��9'�3m�=&�,c�ԡа"OIq���6�������ڕQ"Of�)"P�9�ΐU��8 C4a��"O�c�&��~Q�b႕	�Z�"O�haB	bྤJKN�h=��"O,0 �HmʁQ�(@n�i��"O2��J*6@Y����u�e��"ONi�"ڞ=�l�Vݺ~z����"O�	/}I�9ⵌɥ����"O�oS,Jr�V$�?(�My7"O������0��ɂ���(s�$�$"O�-3���n&�(���@�nU4��"O�y3�[{�t�b�ę&OP]�"O�]	�o���(�혘?.�irD"O�ӣ�T�K:�%{�b�8@z�9�"O�)A�������1���8��� r"O�L)�'&��	!J�=��h��"O��)+�v�-�F�AE�$ �"O�D*�
̚Vd9cgC�D/�s7"O(�9Q��E]8�Z0e��m(SF"O~��'�03�l��t� �3n��"OV�zƖ�0��}XG"�6��|"5"O� :�y�a�2GoZt��O"Dh��"O�9S��J5:���t�� T�|�"Oh��UK�&�=��E^�	����@"O��K"��1y�}�6�S�fy��"O\����7��5�ת�e��J�"OZ��2�p����l8�d��*O���J�LjX��".n�s	�'�lA'�$S�(�;�MO������'�t�gDW">ʠSף<*�(�'�����*a��qlR�/a�S
�'|V�d�)p\h�V臷"c\�`
�'���II�ֈ�bÀO�f���xuZ(p �V6)~<)HFڜ"2����d�F�����;N��BB�����2���ӍH��{s.�+\�Ġ��xh��@�LF�U�Nɫ�`�ȓZ���wL�!:bء���,W����D)>�8����=�lU�� às\�Ey"��E+:�D�4��z���*Q���;-�	C���!�y��ѓ.ً��e���x���-�b@��I�ɧ���D��`͞��2Û(i��Щ!F�}�!�D��kL�� �Q+F���k�D��d�!)�" ���%��	r۔ْ�-_+
d���Ѱebf���@�
%���pޞ���C�3Q �,(:�%T[9���E�>R~I�G`A�jk�L��&�80��Oܐ+���Jw�䪴o@F��b>]U��<;��� +�-'�PA�+3D�L ��C�&Ǫ��A
K�vIf�⒠��s�&��L����Z�$�ON�}�N�@�� �TU"u����"ap��ȓ�\�8n۞@�^���\��)��q��i���}W��AQ(R��2#S�(cx|���۬F��LZ�&2|O��Z�ML�`f,�R�:/~��eF�D �c�)�*a���7�X�S+��J��d�7��|'�,
���D�F��ՙeE&{O��3"/
�JD�O����ʔ���qFҶ 9 �'� ���oO�/���S$@R�:�TɑJ�)M����҈<@
(�Z�#��F��wo�p���Ə}I؀��ʝ	$�q�')\��gH�.!X������f�z�"�m���2��)"�bI����.��$��W�'4���͍.t�+g��v����
�s����G�"�=p��Օ@��k @3d�~Z����L}9D	!�O���Ed�+m�-v(Ϸ((>��0�	�^C���b��L�B�B�!�I��@�x���i��y�@��A�5M�!�0��ؐ	�;>������l��ćO�٩��&��\Kt�X����h��'��kW(V����[�"O�ј���<`�-�=j�0����o%|�+&�[�3�D��fH�K�g�*�
A� (�(>��u��R�F���I87�|Rĥ_|1� � `G�o��Ѱ��/X=�I�wc��
f\ڶ�'2�
���+>�PP�#���-�zЈ���)e�����E$<�D��rW�����T٦��G��(�x�1��;�y�L
�7��H�&L�&��~rĚ1k��PP�H7[�J�R�"�'{�Z�����+���*C;�l��!�T��
�r$���a���A �E��R���}����kZD��$!c�Q��eȈ���kE&Գa��A�@ð�1�G�=M4%��)��)��z�b{��Bd�|=
�f�F C��0<iūр)�Bb?��G��B�|Y�7/4�.�O>D��	%�\-W�T����dS<�r@=D��@��K0�����CF^Q腠;D�`��*NX�`V�� ��5D���'�22����ֈ.�09��.D��:� ˆ$:��tf�:p7J=	b-D���5�P	��k� /(�X�Q +D����h�J���I��ղ0�4D�$���H$>�D9�@���"��)[�5D�`��NL�yN��������H%@��2D�����#wf����iæx��BǢ-D�� �2���ofV���bF;kH� 
s"O�09�J�_P	���24Kc"O���j��	��`�6"�k\�J"On4 l��q�`�V��K�$Ub'�O��c&#�4�0>�kͪA<���ҋR�`�^�0�O\y� [�J�}�Ή�I�f�-Y�Xf�#�E�u�C�	3�&dxv�ZK�B!����;
�C�/f��͡�Z�,x��	?��&�>��4���gŰ2O^�c���w��-���'*��Q�
�4���v_��jb�K޼��⢏�,H�X`TΎ�%n(�d�.��	]��~2�*!���R�k:�S�o���dQ/:�t+P��>z�����)��@IJX>�i�G�4Sjn�8��'K:4�De�#~�@��I�|6\H�G�#n� ����_��̛��Ä�~"���PzЂ%�)Y�Usd��U����1�r���%Ө-
0�@6C�x	Ŭ-�O�$��� O�t;�D�#C���K��F�iP�J�UDz-"�'h�����OP���O�y�"S�d`�|��BJ$5D(�,]��i2MO	$["I�O��u9f�;�<x�U�¦��8�([�f.!��#}R�܊�ۏ]��4#2���o�:(!0ͯ<1�lH*D��`A�<��#��CF�^Ė5b&�V�,����D�ߟp����eE`�"�'�
��� x@4�o^<e�Q�d|�	0~���@)Z��~������?1�_&v�Hd�V�� >���d�R��,!��'�<�p	݀Y.��7|`TC
C�t����Q��qM�(<qO�5&�,#s!5Cj�dR&W!h^��D��	�rS���0�˓m���G'+���Db_��d��D���ToW7ri����"Y��O 4��AD�|9�'���q�ߩ1,�Qf�S�9����Is��t'N}�<7�ey"�Q&R�U����<iO�&S	�E #Q���2�L7`�[aMđz7��7扑{3�0B W*r?�g)��*��V	��Ds�	$p��`��8O�D�0	�Eٔ\*g��b?y���OgzH�'�±4�B��C�_I���X��<u�� ��iK�.L��?}BB��V�. �VSˮe�TVX# �;��"?�0�ɮ!����W��H�u�<�:�$�0�� �	�6]���C�I�OT^m03ʏ����& ��O�z�I`���j��Dh��W8=��с,���󆎏��(O�Lp`FV;;����lu���0���Щ�����>�j�e�7<�'(�e�u
Jj���*�>e8Qn�,���ʅa�b=3 ��x�-ȓ�7��'�1�S�״��@06�Sc�:x�@��E��){��+<�:�킴���s�i�z�1Ub�]ͶI��O��fQ��Cj�D��ѫ��C�P)���3�}�Z��k�lJd��*=7b %�<?wO75�qi��ũSB�+
$r�Ze#I<qW薕����ě:|{�! ���Fv yҴ [r�p��7�� 7r�It�%K��gL7}�H�ḑZ�(��gۂi�z,B`�D2IO��%�Hy�%D{� ڿ��ጒ�E��D�hD�5.x���0�=��10��>���.p|�>�Ol��A߱Z(2���fќ
����DQ�����JF��H�����\$����{�H�h�̜0W8ĩy�l@��0?Q珹vͤݫ���#a���2T�!ts��{ǜ|B��a�4�^�d�Ŕ>!�B/	|��:�6�A� T�<)ߞ6��\�vN�y�.L)$�|�	�x�*D94��I^�FE��#W m��!�.W!��#wr�R6� oqs"ùQ!�R	�l0�HFVܲ��gs!��;�:e��B��e2�q���NJ!�$���F��u샷|5$)��ȂY!�S�0�\��6�5�ڸ *�h
!򤖢db��� �vg�5���/
!�D�9Y��W�!5&z�j���) !�<r��s�H8y��xbc�!��Iz<���˒	+��2C]=Q!� ?�x�kW(̅i[�T��b�=!��,�r�h���A����I(�!���3cp������i14I�d`�T!��58��8�7	�8适K e!�ę�9�j�I�)<����/dX!򤐨"���3A��\��'`23�!�Ď	�Q�d�������e� %F$!��^9�4UJ�C^ȫ�k�(�!�$����X�d�*)3࠻6i�7X�!�� �ɨ�MȦxI�XHc��_�l��"O�Q94��fR Q�c�ĉpB"O��S@cۉ�6� �HW3N�C5"O��*���p��E!v�m��"O6� �Á"s�%�6M�4m@���"O�Q���.���S-
�)�"OZY��#	�) �:��X BJQs"O΅�W�9J�IX��ï["�"O��95G֊z]��Iq��*���"( !�DF�j\����[P>���>�!���'H���V�+rOLɠ��p!��>dod4��1P�A"�Gmq!�d�0;)��p$���_H� �a1Qn!�Q�wn8 ��&*6�b����8S!�3 �%ѥ�����*O��pK������µxJ6<2�'.�pƇ ���d����"	�'��C � X�>h����^p�'XR�	���6u��
m��
�'�^�B���>�*(15H;�d�
�'����'G�/܄-z4��e �aP�'�0�n�������	G�� �'U \�W�FJ����Fȫ.p<�ۓ{B1O�]"!��*%����A-�<@��@�'��s^�Z�	\���S�O���2@A'6\&%�W%-B�9��vuj�E�<��8�\�S����6�Ld܊t�,)[��տ5jH�'*��L	V>5 тM�T��`+��F�5�6�C&	��Mc����l�ݠ���w��%E�Ԇ�[CZ=y�MW��u'DB,m�U���VN�y��y�� �'ԉ���?��m��!�tS%�B��Ջ�$L�A�$�*O���G���M�����\� �㰯�	G�I(ge��,~B�*F2��a۰ҧ�O���q�K»i��#`L�`��i1J<V�ض�j�r�8�g͇'�����ψ	_CD�a1�>ٖ'��~GN��Iq"|�'���B�?L�J��a��yO�9Iߴ?S�D��t>�ӧȟ$�	��M�85.P��aW��hum�P�� �C�"}��:&��:�����.)�p� �8�Ⅰî�|�ɩp5p�	ç Wp�p,(2�\|zTHS&e(t$�����&M�T� �Ӈ;|�u�&
6 `bL�2��H2x��Q�	C�ԟ@���O��2f�G++����,S~  ���cgz��"��<�%� ���(�!�R ��(O�G�T5"O��р��-:����
�}@t���"O`�ȵ���,-��;_�b"O��� $"��F�c8,��'"OV���iX*M3��֞DH[�"O�y���̠5��B��Z��
Q"O��d��"T����p.$8�n�R�"O�,��!��Ds��!.Ȩu�h,B"O�����)""�(�gQ�T�p�P�"O���ѤU�s�{��b%�EX�"O����"R�b��d�
�V�S"O���W��3Y��Q$P�N�έ��"O��K5��.v6��7�L�Z!��!J��������Y�AKk!�_U�2`�c�K7JR�2V��4_�!��ӢG,R܉Ҏ�3u'�9�3̄a�!� (�E��6$=D�ɷv !�$��Y���#�@^� %��C@�)K(!��?l�D@����P*�hwƙ,G!�Vu쉸�Jܲw4(�䦂
h�!�R� �ȃǺ"r\lrb�F��!���otq�´���+ m�-P!�DY�5V8����1��ab	5k/!���(�����pe����:�!��"����G&H&�\@uG!�!�$�d1��j�)۶}yh�
c��n�!�� ��C`�2�\�p�Cg	B�"O�1b�G�s\̰��.59J
=H�"OlYK�,��"�OĬx-��r7"O�ũ�Q��Q@T��;B+�M��"OR35��-vV�XЗ$�'FA0 "Of��!l˰E�J9
vc�<�p�T"O����Y�2�a(v�5T�,(4"Oj��׮9μ�p`�*&�<�+ "O�\SkX4N[X� �N_~4̴�!"Oba	aܥ�v�Yao��_
.�&"O l�B��4p��\�p �o�!��	�=�a �b�RM�e�!�D Os��X�a<+���%�Q1.k!�D�3_6ΘY�̌�{�0�IŦ�@�!��
5Gw����END���E])C�!�� $����KI���	P��#Ei!򄅻|̄��N˼���{�T�[�!���;p p���׌��؄��y�!�$��o̶	y�L�&"��$Z��H�a�!�D�� &J,gx�*�N�X�!��J�KE ���/�-"H�e�!�d�#
wf�C1Jg��seZ'j!�d@�c8ȡ�&�"Wej�@f
�*!�d��eW8�sSiR�BG(E�I^��!�\�=�`)I��Á=����Z!
!�G����K��u!Xm��䘱]!��g��͠w���H%���x*!��Vݬq���ؔ��I`�[�
!�dJ�*�H�*g�Br).-��A�5 !�{&�(�)L�H)l8p[M�!��_���AP�sD�{t`�6�!�:_�x�%K�o�����F�!�dW�p\�Dz�ːb��dp�M�m!򄉾s	Jh%���'��e1D�^�d!�$�)55zL���~f��C����. !�$��n�(��%E�O�8z�%�"�!�#J��6A�vB�my�N�%�!�D�X,x3���(�T�Em\3+�!��E3��X�K]�nh��a�зe�!��_��ŹQ�A&mX�dۛ&�!�dX4s����mճ
�0� B�#�!򤂂A�>�3�أm�^�B ,�8�!�dM5?pXYrS�e�D`2����C�!�2f�^<���P�:c��y�ʆ!�d΅@�&����G	�Z����[�!���?@�0t�Ìy�A�JDO=!��d�@�s���3��I�1�M�Y3!�D�����Qc�˒�T4S���P!�$Ƌ$�X(��"q��e&C1�!��/��݂�
W�cRdh�e�պ9!��C�L�4�'V�ಘyӮ�3^�!��]�ade��O�8J�&�fD9x�!��)Y��a�1f�-P漌�`D�-;-!��03x��`�S<� ��cʑ+.!��:D�(��.�<*Cv��bJ!�D�� '@}4��s��T鴮K:YM!�),��Iw��"9W�e��
�!��� _X�
G��PKX����%0�!�J5l&���`�� 1�[�!�D�'(b�hDJXz��s��(<�!�$=W��1RǊkvx��3�!�Ė=�@�ˉ"\��M�s�!�D�A�1"���$Y������!��R+b�$Sa�3��}ˣ�Ē_t!�� ��8���}5Ȁ	\,(�b�"O����*٫ �����H��m��3�"O�Y�"���[u��-�	0�"Of�[b��L�
L9bg�.C�@�1A"O`akN�)M���1Kx�4�"OB�A�_a�u�σ�p
4�k!"O
�qF�����,rAԌ'���B�"O�P��¼?��� 
�!�J�� "O�<aCD�m���:c �Ps�"O~�a�M��!�\�.W�Q��z�"OHxѓ�ܵ_-X(+V/�
3pz��"O���'�D�K���W���s"O`�3�V0lpnic#�7�)�"Oΰk�"�Otسl&1܍ҳ"O��å���`�!��+jLQ�&"Oa ��}d:}tD :6|�1"O�d�T��;��(����U�e"O����Q�n
�3dO3q���R"O�0�� �a��,3���C��4"O� ��H�#�����߿]�މ��"O�� IL�6,�H3�%��BI�F"O&}ٱ��?k��@3BK�d��$�7"OP����x��H�w�2g����"O�щ@�L�yy�	Q��C�k�l��"O�
1� �Xz}aã�8LԐy"ON�V��oj\�R��-�PqI@"Ot���L�'>-2���%N{��R�"O�Q��O���EK�o_�4dh�"ȎCb`J�^��2o��(i��#"O�"�h�'LV�� ���@6t���"O	XW#Bc@��3��' 4+�"Od,�a�
�Y�$9yR�A,}ܵ�C"O��%շ:��-�rFʦ;`�E�U"O���G��:]�� �ߡhJ��"O�t8(�-:����mg8 ��"O"UB�,S��	���0(��X�"O�4�,�[�"���J��rĥ	6"O �#��Z�D&��s���9���+G"O�`��hOt�ht	�V(��b"O����攐�k�$w%!
�"OD��+�/WjԹ�gW�
`��U"O��ܒ�p �$&E	�X��"OPh1!� t�$�Y��T�⁺�"Ov��фN�f����AJ]N��%�q"O�h�&D
`-9T��W3�)� "O�J.Ǭ2
hp�c���7��}( "O\�XA�#�t��S��T�YW"O��A���0p�h��":�����"O�$�7c�Zv��S��U���a"O
9	��MP�Tk8w- A"O��p��U2�����Ň�Z̰�"O��Y��)z�8�����r9D}P�"O�E��X��(�d$F�y8*-��"OHۧ�� .2���E�7ƽ+""O�)�#�&dl�{�C�<4�8Zf"O���3	>5�H@�ĳ<h��"O<X��$�w����9R�ƭ�"O�X�cމJUVe#w�?>�&��"O�� �Z�a��� ���"OL���ǝ8�zP�7��:�P��"O��wEʟp�r����;�H�"O\���l��8E� �oE�yB͠"O5�AЄrNh�1�#��bU �"O��#QaB�h�X�ya)��65�"O� ҉���\%�	k�H_�z��I�S"O�4r�����X�Q�й<���Â"O�h�@��H�|�,�4sL�h�"O|��#��H|B�|a�k""Ot�3TK�oJ�|����r�� �"O8�`��P�ln�x�֍�/[�j�"Or4B�Z1�@�#�F~0��@"OҤ�D��b\8S�G�/i\���"O�AC��6��4���
<i@�;�"O�aa�I�H:��Ä�WC�c"OH@�&��*EI8�ś�f,�$�"OXX�JJ
#��x���\�w)���"O~��&��C�Pivb}&u��"O0�S`�цu�(QCF�t�@�*T"O���f$��hDPY�a�:K��#g"Oڨ���Z:iJ��Y6N�<@h�C"O���,�o�ʠhw'��@��)�"O�U O�#Q���RH�Z����"OJhJ������q'4m��1�"O�DKe�X�)�����>�t��B"O��b���uJ0�+b��I�R)9"O���(Ե[���ȳB���ȥ3�"O4E���6w�6�X��G�DZH�"OF�9aB��xN�!�K�a9L�p�"O��/F�Y.�=�`P�;-�)g"Ox|A�H��r�s�
�:�!Q�"O�	�%"�9�(�`��ʊ9�E@"O��ɇ�L� Zt�*� �"O.���l�B�P�'¥h���J�"Op�@���3z��Ҵ�'��)#�"O(x1f�O�a˾q�$Lƥ *]�s"O�x�rƈ!"�$!1
��!�"O�i���-s�T���	X |�Ep4"O��I����Ċ%�I� )o����"O�E·IB}B�� )�3�`�1"O��Wg�E�\���C�z-rL�7"O�e �H������A'�(Ԓ�"O�0�̇XP�D���ֈ��PXD"O���)�%6jd�� ��M{.�R�"O�`IB��#�t�&#�&Cb�d:�"O�:�a�b��|��J�p$c�"O������,�(�æ� -� "O�9�p   �D���A	&�����4(���B�?D��Ce!һd�"�G�U�_��Q(w�0D�d���#���Hս^:`)a�H2D���f��q�(#5�-�,����$D�H)Pa4��@�'�~�A;֊"D�����U5uE�E�e�Q8���B,T�,ٔ� �j�b�R�h_�(��A�"O@����/��%p�肖N�p��"O���w�fR��8dM6`��%P�"O
ͫ�AЃ?���<�"軰"OPZ�b����0Ɏ
b�P��"O���    ��'���{s�R",� �D�8,�f,�'k�T铤�r��*uI��
�'���R�������H7\K<ň	�'sv�1���
6� ���.JBF�@�'94�9�MҫE��jD�ݬU�|�
�'� �J�#΄GU���D#Ve�us	�'�N�;ׅ
��� 0��]��y�'��s�>K��9�g�+W:"*�'o,m���*"x5bp	��T�
%��'���q��ã��:���=K&&��	�'��`�&G�L�1�� ^�F��	�'i��k �w����%b��2 �5�	�'�|����F>n~����䘦D,���'.�T��*=���EÌ�=&�٣�'�@T9�h�s��U�R0��S�'��0`�ʻ )`9��e�5$��'�nT��n�o4��f)܍w�]��'�hu�7� ��hx[F+�5Wz84a
��� �����α�v�˯^����"O��) ��u� �I�M��F�� "OVô�ѽ},��K�Z�x�"O<� 񂔪i����"A�\�H�k�"O*ᲀA��R�>�Y��õ����"O�)8��ƥZ�"TPO%{�nqq5"Oxy�G��8E�p:�o3�����"OȬ����,�~�ӫ�:�Q�Q"O�-�ୌ� �q2�P�O�(X:�"O����H]�p'�YͮD�C"O�����y�|�K�a�����"O9k���ZS�)��@�[��t�F"O��1S��-�|L!ƀ�v�88��"OL-��J$ߜ=�N��/{����"O�0jt*Xz�Hmw,��5
r1�"Ox%:V^Y����5�j)��"O.`�6�Fqp0��"�T���@"O0��ץ��6��RBaC%#}dH��"O��;��̵hZm�f��-ZT"O��鲌̝TfQk���0�8C"O���EM4�`q���ht�w"O����#M�A�� ^&>�0��"OX-��+.6ql���%�5��H[�"O���ƪW�Ҥ�w���p�F�Bd"OB�9V�ݷu=�"0�Ogp��ɠ"O}ӐO��^�dIЀ�>Ki"�04"ObP����"G4�����WH�*�h��*,�=y���OPx��o�@;��]�3^� [w"O� �/X�
�E���:>��Q��i��c���)�|B L�`������#})�p�$�p=q���7tXk$�l��j'�	g�0��G�, �͒;=!�].�����]�-₨R��O- �qOP9�r痂��`1���D�p�b�(��.����
i��qj4�	�A2vx X�9ɦ�� &I2XA�J�ㆴ�}�O�8�M|��%�faDK�O�P�gԁi�P�"�BO�|��"O�Q���O�%M�Ӳn��R����&o��[<�"���/���:5o�l��I�����~���$]�g�D�p��2a�1WC�?�p=!�XG|�����a��9���8=h2�p���
K"��I�.�!.`��ӦS�&�N��X���?�'Clhi��� ' ���'H�uX�e��{2$A;(�&|[��[�Ol�%�r�]h������R;�3"j_#(�F)8�e�����C0<O�84��qJ@ps� .�tx��I�B��\
��>���~�d�ev�-�aB��$ d�֖ũЪD�;���9�[(`�T$��y����%��$v�9�k3\%po�w�PY�$ �;�~�Z��f���ѧ
��u��)�H���A��c�bmxG@�Q�{"lV�v ��'�<�@'P�'9(��d�9x9�C����RӞNs���ǃ0��OD�'9�s )��m~��c�ªrM�h��'�)��ʵz��x��o�1\�k�5r�x�_'�����V�E�4��I�/Iސ*dE�W�qZ��t����gP�Bt�P%m�=��k�4I��b�m�si\�.�$vm����D9$�8����'��#�a��1�U1G�5?9g�C_i�5�N�( �Nh�QD7q&���,��&݊3"ZĨ��ɟ&�\C%"OVt�	��J�ڼ:�ML�=��d�SD�I��9�d)̨f�ʨ�JL%=y�O���$����%Ƅ{#��f���RPB�e��G�);0��ɊD�Ҹ2�f�q�L#	���P�2%�|���I�ayr+]�v<1� �k����VD���On�yPD� Nض2�F�T��*�E�3x��Q��5,��a��9�,��'c�H��d�c�N��i�;��.O���N�'�<4�Z�.Z0��X���O���	Ն��ب40�Z��ܽ��'a���d�@<"���d۫h�p\�d��>H�X�S���H��ꆉF��'	J�ODQ�$֚
$�!ĬS!��T�'�Ld ^"��x���P��ؗG��/�B)�EB�D9�)9u�X�{���DV�%"�1�p��	1.� Ŏ�h��`>T
!�<�/�0�@�� �؅*s�\sWKM���49��G�V�"�+S�4)���n,$���#*#�����_L��y̂oy���:|i>b�0��h!�	�x�:�M��QE�b�� ��A�G�!+&��'��P�)[B�'��q�燿,*�����	'$�q�ǽ t���B�(O��@r!�VLt�  G�//���OD�'�6x��H�<k
��]��0���#f�`�y�5��'	���pn��%r�1���3k}T���1q�a�tVZ!���'��A����P��.�К�0(OZ���θz9T{f� ���O�)����$�D
�a�"=a��ԦT�D
(�Q���dH<�"
z���3�K>�ٻ�+��(��D��h���#L�>�v}�B
���#�>�w�����Ȉ �J�[Q� u�B�y��f���ɦp>����
e�^�{�)�1;ǡ�?YI�@pf�5}b��|��D����d�V�Ƭ���R�U�pq�#c�	�џ�:�N��O_F9�eM�q�.�Χ*?�H��JH�`|l��+�,lڄ�'6���"�W1X��yÙz�4���+�3��0��;��/1¬*P,C2t�t�� �>�S9v4�h(CO�,n�S�`N�|=�q���=!��2:�%2��.=>й�Ċǳ$<ۓᛳ"��$O�r(�0��͑"����Ο�h+���'@6()����kf��a)G�Ch$��Ü�2'hQA�M��j�X$�B/�0>Y�k��DZ�yz#�@5.�*�h�fBF��@0���5ʸ��1O����N������E�A"Ob��`�,�~Mz�&�<p_bأ��D�8-7���q���~"�A�I��y�O��d;AN@�1�LBR��$5�}��'�*<�#�PD�Ī1�O�(��<o��v����ӆ
'$�mG�A~�y ����j��`^�~�4hTj>D���᨝>\�.��BA�&��P
Q�H.�����Қ�~R��qC���n�'xh�r��主lH�X1��',֡�ch�!q�@hhD#=|q��睻?��1R��FX�L��%Ķ]�4�#�F#)A*���-<O� ��iG /K$��O.�*�1z�Bed]�ʰB!"O�1�"W�"T.�#ǡ��r�t���|�K�w�j�Q���c�O���I`f܀p5:	9��e9��	�'�>MQe�P��� 8 ��&\O� �hR�V�
�'��PQ���>qCR�0�`s�p֤�Nh<�#(�"�*9�R��#*���O����p�등-a����֠78�	��ID^>A�U.�&2�y�	|Y0]�nZ[}��I�)�F��D&��~���B��y2���[\DB@$[5P�d�"V*�'Q�t�r�V+f�?���.Y8g�-����6.��)V�8D�,+���.R���*Wm�;IF���X�yJ�xpP�<1G-��!2$�L-uLJ�藨Xn�<�A��F�1	�U�p{�ΐk�<�A�̂#_�r����
��5�g�<)�)�"6�^)�E��*E� +���d�<9�߫@�p�*R� �n'�	{�`e�<�4��_�j4�H"ya�Hj�Yb�<�Q���)ؒ�1 �
V��� l�Y�<�'���qP�D�T���=@�P|�<Y��W0�Ћg,��2�8E�ǈ�q�<��ƈ4R{��I��пRߎ�3a�`�<�`M��=�hP���7G>��(u�Xa�<I�+M�WZ�"痱yS*2R�_�<	�#�9e3�`/d|B!z6AQ�<����)�n����
�:)M�čCT�<��蛧N���{���l
]1�f]�<1�I"o��k"%�:\~�QHL@�<��2nv�q��lU�M�z�P@�f�<!f���+>�8c$�t*����d�<��Ç�/*��#s�Zj��Dc�<�7GB ?��03^�R/tM�f�Q_�<�ISy�ј�eƱv�E�"IAA�<�"]�,%(ոE�ȬdO.�@��Hk�<q���~��m{5k�6�d�HA�	`�<Aϔ�UVh��@�=H���D&�a�<�U�_3T���Ap�,�����aMb�<y6��::�=S`$ۨL�L��4Ze�<���#�갺��O�\Ԫ�᥍y�<� �������=
>��pH<zmx�"3"O>�x�"��VJ���ND�Z5����"O~�eۂl�I��� 2t�r"O�i�bf��{kL��풥l�В�"OT`#���X5�`����<�"ON�	�^k� ���=V����U"O(�	�%"y�Xm�_�p�A"O4�ɱN@��L0��͛[�<IB�"OL�a���0� �wƌ>ab9�"O��1�^�8�r4b�L��W�e�"Oh�2�/Hg��ɝ�^��P�P"O2���ӧ�8=s�Ͱ8.lT�"O4�����0�̊�b�Q�d�d"O��ˁ���(��Tz@M���3�"OV ��� �" �)��� ��P"O<術/�=g7^IR�K�Dװ��p"Ot��]�:�8��-9<�*�"O��m>6b�yR���9����e"O~x��#��"�8�B��r�z�Q'"O���E�7�x�fM8g��)U"O�X҆��'؁�D����.XZB"OF)H�=Z���U��~Cj���"OFPk���n���u��pD�Ug;D�꧃ʯvj��I5c,N_b� @4D�t���)6�X�b�,�,��0D��󵤛�1��ӵĈ#R�&��a/1D��h�dC�8����8Iol@�02D�P4�(M�a�Udƣo�R��0�0D�`�V-��N�}�K�$x��=D�0s��!t)���ȵ�(��K:D��zak��>O��@a��= ���E*D����se�qB�F�>g�-�@+D��c����).�dX�$Ům
c(D��#J�	6pɷN��jXd�c�%D�@S�׭]�,�+	�>`W@q#�>D���W/( a �?�N	�&D�l���ѷd�TX�aW��� �A*'D�lA�DʷQNh��U�m���"%D���`�Yr��s�P�}�|�(5D��p��Re�јªU�]�l��3D��0͚�y=�ČR��\dp(<D�Ps@o�99��d��K�TK>T���6D����
�&Δ;���Y���ȱb4D��1�:nv��p�A�;><�H9D�*�K��d�@�:���Y�^�A0D�0:� $:P|�D�\.��a�#D�<j�x3��HC״����Ư>D�4a��*C�Ұ�0W�	�ҹq�K?D����g$�(�cb�=j�5(�?D���E��e{������:���rT@1D��c���z���@��qA�	,D���Vd@�Zŉ׌fJ��379D��P��;���"�eJ��v�8�/7D�Т5�*iй���y\�53D�\�πg����c���>3�3D��{Gi�z��K��<}Fɋ�:D�\� d���GC�P49�Ǝ8D�P�@�X�qIZ	kJ��A�7D��Q�%������R`�JD>1%�5D�@�bjߩzv�p�dC�i9
����/D�@���۴fW`=��"
�Z���&D�,��,Z,6�h��@ަ72�$�8D�l�A胴eP�㱋�z( e@��;D�C���
J�,HBÅ�+e�X�A�O#D�� F��듽v�0��Ȕ&`d"OnMaԨ�0Z@j�PA��0�x�e"OHaP��13w|�
�J�&�p4��"O�bQ��V�c���8h��`"O��0e��0��m]&vl�"OX,�A/��)�y �jC.Yg�8��"O�)�/��Ң�Ӈ!Lt`z�"O\}:«̪"��)�$Ö��>�Ї"O�`��A�?�M��eL�h3��3"O����YmL�01G�-�cv"O�H�M'�f���w���җ"O$d���P8#�t�Ă
�Q8 "O&��.�
=ߨ%S�N=�p0A�"O�q�Ƭ9�*DC#l�p�&���"O�M�� �R���eғ4�t[�"O��J�G��t#�	ஓ< ��(E"OԐ�s��{��YómĈ1�N���"O��K��s�����@�O�&�Q�"OR�Sse�R}|]�P��N�"���"O@��G��>.�>�h�̆�� Tz�"O���o�e�pջ��(>댬Q "O����B�'� +S�+Ɉ�J�"O�����p��3���f�d%�'"O(m`�����*�&թM}���"OR����rP�!�H�
y�ݒ�"O�]rd(D�%�� @�\��X�"O>��ol���qò�pqB$"O�@!���"�2GH9��,y@"O� k�@�&��uMR%0��e�"O���"ט��8s��miʴB�"O(�A�IL�7FXI �F,�p����e��`�=ي��O*E	���/_�@x��8Z�HX��"O�`�`T*v��4͕!����i��b�NA���|���+X���a`m�k���㵋�p=&@Z;u�v�
��s���s/S��n`��G%lӺ�ӢI/D���䟜- 8`S�B]1F�*��

��0���L�"�?=�A�9B���U���4�1�(D���aᖐ:�t)A̓a"E�H*v!��7}��Q����		G�LRF�;Y2=b�ǘmJ!��9�ܲ��?D��aT��$R#��{�����k�'�,�C曩y�dwa�:Z�Z	�1��uxt��R�ɿ(�D����{�U(�R6\>�I�����S���_���9�T�pډ�$��05�\��h�P��%�"t�:`X�����ط�N���.Թ������<��6��t ��[�8�v	��:NTP�mG�$���OBFʒ.���W�;��R��b@�v��mH<QB��&J���rd
�_a�u$Ŧ1�� Z�H�'�!"I�#.F�>�';�J��5�˸>�R@�'��8�X��I%|p��_�$��K�]r�� R���q�x��ò�����$?�
׫�o�4�?�'�d�{�B��|�!@ɆL��+�'�����>*����@�*�i�ߙ"։���B�#�,`$I��<yF��U:T�`�A�(M(�1SEx8��@�BI�Rp� ��g���)5c�7h8�١�N�-i:���&ԭ8��q�ēh7��PtfW�j� �Y�A�:5�'	d�8�ʌ�!��ezR-�������@6�-\M
��4jK�$6Tp7��;V�C䉄��(�
��
|�q��m��`��i�	Q��`��c�Dɸ)*�I��ēe��XE��G)��%� AS45��ɓg��p�����`�*U�DoG�@?��)g��$_6h[�ҕO�bDs4cp�ayR-�?lb�5 �o��HMzM��ԓ��O���v ���:�e%�PEjd+U"��:�	�,fx�D���-9
�'��U�ȉ4@*���#I�^`8�B-O���(��"n��tK�x�"�͐���O�����$ڻ!�J|��$\�F���'Y��я
�Q�Ӳ�[�\�����Y8��� aN�.���`���',��O}�� J,!���1�^���i���'>e�� 0���#¨v�a�fbS)D�]�%C�,<*�B`�&n#<�aD><O�u&ͮA�9@#�PH����>y�T#/���3k|��(��S���JbG\.�R�C�ַ ~�!hF�UR
m����q�lC��;r��QR0�Ny P���ǘi߄��'4��hՂ@g�m�N�(a� ��~ݡ�G�٦���4*�;�N�P���
#��b�ҁA�R�$�j�и*x��3'ֶR�t@ӵ�R���" �:tha;�	�4\j�G�x���x�?MI�m9�jЕ(T�4���	���O05�7���D_�@K|�P��4fs���ui�^�<=b�@y��l�dţ�(�`X�\B6b�S~�r�(�V��P��<��*١jdB�RC��O���>�!T�_�M�R��%b�K�\�ViQgti����] !�B����82G�.{��9�gC���  ����yB�]�}:��	`.°���xR�Kn��|�1�ލVc ���P�Cs$�&�'�O~$:�)�=GҰ����A�
�9�_:gf��s���.���,@��U2P��aHA�t��E7F�/9ᠨa䇝CDХE2�\}����f�|	a�6��(�Z-6$�����f4�p��L�E�2�l���!5��@�J����1�M�=q�˓Up@0�/G-5����ר���Oz��+�f��f���µ
�]6uA����<�ȓd�S��Q�}5�	�gO�*i6���&L3p���􌸺6�J@�g̓��`��
C����գ���!�Rv�@8�n	�gJ�XsO�<'�bQ�'˃�R�(� E	6����$,pڍ��H30���DE��z�$q�y�!��<!ucLV�6U�rj��@`�M���G�<�ǅN�	�.݃�A!��!��Aܓ`B��#��,v��8R�r�?u�b"�g��x�N�_��	�$%%D�tAB�U)����3`�ܱ���B�&�V�r�O�	��.�<��|BQ1���+�*�~�4���BV�� mH�"O��)
�mM22S��&y���/>m����d�`?� d����4�(�D�0P!n�ky耂��4��+��ܚ2'O%E�%�B�шu0��k��ȯ,y�tbT <�O�y��`׆t~���q�ї^fL����'|�퉱DД[aF��'SP}�d�/�TI�(~mK�'B֙�A�L�B͊�oV����3J>���ֳ���r$=�����eN��ۈ�b0�(%<C䉳g"x��!�u��m	TO<�	�b����	�z9��OI��\�"̸-��L�E��9�OK����<�r%�t��yӄR�G�0�b�3ɜ��� �sԁ	�"ɟ��ą�I�r؝1�≞��	��$�fL�!	�E�&��#��C�"6�@Q!q��<'N���GKI��Fb����	�B,F���ɍr��97j��5������5�y"��5L	�6�Y�'V
y!��3[��Uˌ{�m���ګ�E{r ݣ7)�9@$)ʫ�!��V_��'D�%X��+@�!�D��0�	X�-]"&f&�;ЀW�6�!�D ?o�A	p"���ʠc�K&_�!�P�(�81��ؿdM�ӱ�T���ȓRƄH�	�x��(8�eN�;T,ԅ�a=���C�a��#r�]
�Jy�ȓr��V��L��k�S��� �ȓVRΨ��Κ�`
�8�	��G��U�ȓn���e��8r��@��3����H0�X�r�+F>��i	0O����1��+�n-L���df��j�b,��hp��6�xx�Y	ԟn�� ��Ak �a�,S?�< '&J�c^���%�~u�"N�()&��J �D�&�ȓ,�h�Y=e:���m�0b+.a�ȓ�&�cϓ�3PI�],g��l��l��uK!�
l�^��i�+�b��m��
��Q�3%zM@#�Q8A^لȓd� y�e$/f�d���`N�H�$��ȓH>ʼ��ˬ.@B��եLHDF���!�|���G�6U�lO�8M��8�D|��#�V�x��>3"|ه�S�? ���2��LA!7A�6f��"O��S�
�5����p��	�����"O�-�g�:z���6�$a�d[q"OK��.eT�#G��=}��3EC"�y�+��j�P@M^9Z�9�bƐ�y�ע�y���Y�_���PbNR.�yr�V&���a�C�T��0��(���y(�
�&�����V�8m��GP��yR+[<�L�E�I2xtB" T��yr�Ȯn-�����S�MO�8P�#'�y�+O�s�xA��%�T#���!��yR%E&�x]�rcA�@�Xt;�D��0?1�!�!-&,�P�L�3�<1��+(�d��Ù^�<���^V�����ѱ~�����Z�<�b��G/]�cJ�(X3�I]X�<��Y�6�J"@O#o�-�f���<�Q�]�Y�$�ul��3���<��ȮO��D��ǻ#W0S���~�<yF��=�8���-��4{��o�<)���(�N���e�Y�<5���@�<�c�ІGL��4/�/.DMP5��f�<)g��=Y�@���P�V<s�Ag�<�#.�97�+��ǳ>ː�$y�<aUM&n��)BE��x0�M�7�|�<���!ef��Z���_v~�%`��%�M#V+
���	��uw�7����-0�CҨ��8c2e��B��~��^F�~��	Kw�퓓<�� ��F�~A")|38�c�H2.N8i��7}���_*2��7gR����Tm�?%������
zr���0|2T$܊XB굱&�K�c��h`�J��CD���O(���Պ�&����iS�@�ZE�҂�94DZ��'�\�O�%���qfLM����&H���*OF|�B�F���a' � V8X�X�'b�}*�K4u\�����F��� 	�'�jm !��,��@�Ԉ?�R��'��P��	j���8�� &t� �'&�8+�Xl�԰��5i��(�'�:��wc�<GB�����.��Q�'w�!iQ�˂*�D�B� �~Ġ
�'��pBǙ\,(z�������N��{����%������.3��ȓ�f}��ӳ!w��õ�"ݺ܄ȓB����^&L�<!U�ު��1��_vl����=A�Fl�*_�� ��x�F�2���%j���u <Y�h�ȓ �4�n�6+�`h�S��/ͅ�"z��$@Yd�Bt ��3:����9�2XʂʭP���j��D�x�����~X%'E!A�Vb!���:�q�ȓPCH���X�2d t#ė,"���ȓb>���NԪ_{�0p`��r7�4�ȓ]���r��B&r��}J�/¸;='\��D�/����ȌZ�f	8�	PQ!򄗄3jd��֪H~�Iȇ���!�÷d��e𦭞#wx���AZ�!�D4����&XU�ĊQ�Қ7Y!�d�X�ۥ�B�W��pq�ƘCO!��X�"�H�z� +�͚p�!��*Z���a���,�9�r#�15�!�$�1jQ���I� G@��`	��y�!�$�����'d�c�H��	=�!��'@��Y���ɯl�x�Wg8`�!�$dJ34K��}�^�'�bi!��`-��M�7Akؙq�ȍ�_T!�d=��ъ7���9�r�^�]8!�� ȐY��6IJ�(G�ÿ*�����"O�����$w�qA���2�D�"Od<B���}�Za��ƥ1r|$��"OL((J4������Uʰڰ"O���Ke40�٠d��Z���j�"O��$D�4>���dD`Ty�"O�h�U��)P��4{с?���3�"O�tUfJ�kM��Y���23."O�|9D�;8Q�b߆e#��"O"ٴ�3�4j`L�"�$"OR�V�Cұ�*���pKd"O}{ (ZV-��c7iE�)�D��"OP�K�EUPt\Ec��[��q"OxŃ�M=gV�,{�eM�5�L�[�"O��I��)6Nm��eЁ>�)(0"O�a�X& E\�`�ق0xk�"O<&��_m:|���ԋJ���"O@�v��.`"��TM���
��b"O�i��c9�6 Y�Р�!��(_�l�3��1Ҩ�cΚ��!�:*l����M�N��r,��YO!��I��~,���LD���H��͝HL!�dCq2`z��#v0�j��!�$S�~*�5j���jZ��t��\�!�Ĉ8ܐ4��G�&cE�i6)Q!��Q�~8T	�e��k^�Z���9I!���p� dq#�D� �E�Bq�'�8��ف�d2�lǄ7h�x�'��y�eC9#�d#��@�,�+�'p���ÿg��1�G�ƾ8 ��'���6C�v!�`�N�\*X8r�'�r�3�'��h٫��ٳO|�l�'��P���hm�\(�$^�NG�}c�',���3OA��{q@MR*�b�'e,�U��@�	�
B�.�{	�'J~Ha�a�c��Ɋ�
>$��B�'B�;��*	�E�R��%D�Lk�'� �[�$^.qD}�¬��B����'tV��+E&;��1ڡ�WLH�0x�'�f)r6�^��`kV6���
�'xB���B�d�xu�2'ߌ�����'���:��Y���%$�p�S�'�ʵ����^)���v�V/)�9�'�`�b�O��4�u�Ɯ���H�'3*��[�<��t����A��'�V�a�`�)T�K1"
<�'�`�BA�5{�~��B��t�q�'	�m;��A>@y�у��m$�b�'��(%��9���&�/lg0�
�'F@�U��l%섢7���v�p)�'����u,*��A?��p �'��b�PJ:0�YQ�S�<+��
�'l�p�x{��S���7�B���''d�
�C�Z��K�`|��''��8p)A�Nv�+`㞣+��|P
�'�.y��.("n�I�g5(��H�	�'��]��ț-�\��S�#���K	�'V2�0�%��	��Z�F=!�8�#�'I�,ر烣}ښ��с����\��'p*RlY2F�������L�2`��'vj�r�V	!Ϭ�yUA�*=Ƭ��
�'ZݱR闑*B�h����<e�`�'{6�R�r�X����!H�|�	�''Jly���hzT�4 M�BY�	��� LMc(Z�X���s Ịk�� "O�-��4;���S꘳j��P��"OĜ�ƃ������:���i�"O�h��)�IrHM��Ň<�$�"O�`����0� Qz&D�-�n�F"Ot���n�4U�w�$(n����"O��;gɤj�x#geA=YE&��"O<��b��6x�L2�C��Ө���"OR�i�H��(LXc�(/l�`$��"O*��b��k.�Ag��J3:|S�"O^�` J?�	��+��%�$"Oh���Dr5����V�x�#B"O"E��	v�j$��c�h$��"O���
#�XC���O��d�"O\x���,m˲ ��y��"O0䂂�T�Т��/
HH�0"O$,R�h��8~<�*fk��<Q�hW"O�!!`MR0~rF��%���"@(�"O ���bئjwv�������b"O.IѷoZ���3��,7�ft�7"O$�Y�d�/$9։:���f��1U"O��`�Z��������(�"O
,x�y�x�j��23�"OY[���=<S>��Bq��}�"OtL���^�r�H���/uZ��'"O�$���KJl9P�_b��`"O��a�C8ː�3��S8#PN}C"OZ$ �I3@�ڕq�N��cW���"O$9����1�`�@$	7F԰�"O6Q�rfs�ְj�S#Id%�"O5�.('��a0���Bp9�"ONU2⡍�V
t+'!;��9�"OA@F�ψ:��ҕ�ӘTtI�"O|+���$T���1�#w���T"O�)��Y�P>x#Ў]�I �P"O"����R��Y(BR"�m!�"OX	�1N�:N��($[Ppw"O��yd�@��t�"C�i��ЁQ"OP���;|�>i���0y�ШT"OB����!Wj��Q�܀L�ꜙ�*O��ď9~�T�{'V�fI@T��'#�e	B��$X�� !/� EK�'\�����#������)�Ȝ��'�
�[�i?I'HUz��N�|����'�&���K
7l��@�ǇM{�� h�'h^��Ӣ0�^S�GǶy�@��'/R=�%+
_<��sF���b�p�'���#@�s<��Y����E��	�'G�\{vdI 180�բ�@�H1C�'Q����X�YyF �4�� �'b���-�5m�6c�eܩ	r�i�'u�I�ص	+^�Q7�^�g����'\�x��g� J��X���]��,S�'Y�@CfѶMK&�	|�92�'����\�|�t�4lU���'0\�Ǧ����14���,���'r����D@�u:Cɛ�?!�h�'tlɒhU[�z\�R�̜O\F���'��R����Tg'{�&���"D�$ia��P�rA���I��ܑ��2D�����T����9Wn,�f	�Y�C�In.�=�磑��h L��C�	.G�:�u�e�F0˗I�3�JB��#��B��A5`I2�#sC�+L�C�)� Z�hTbO�vY�)��ˉ=��r"O´�G�R�6|С��_X���"O�\�"�	NP���N�C縕)E"O�T�S��;L5�Z�-9(/���"O8�� �W�rMSS��1yZh�"O�\ف�$B���􄐠w��b"O$�ᇆ�s��� ��x-�A�"O:��w�v��ЄB��P�"O�����|9(���G�0�	�"O�*2���������5.�y"�"O �a��G2И�M
�,lh�"O�P+�!�Cɀ5�M5|��D"O���Qi�����rz��"Oz�9�EÂU�V�K�!̐d��"O����
��hK4!H���2"O���f���q���+��)J��h"�"O(�ɔg��/��Xw�ҡm%h5��"O&)����%k�J��!BԺ!�!0"O�|S��I�u�T���7�z%��"O�+!\�M�iPLҦ:��i�"OR"Ƌ�;.N�P�J5GRXH�"O\UǏT!�	��� I����"O~|�G͍Aƒ0	�'�2C��"O@��^�y/��peW�h;���"O	*tÒ
�$=�p�Hz0z�"O�p��ؠDx�"C"/*�H�"O�\�!��;A��A�K�2L"OD1d�P);�tiP��T�%��IA`"OJl��&�	R�*	*�]+�V< �"OD�p4n�'R�Jq�P�r�ЙJ�"O�������܊ mR%I}��9�"O�<���<H�����ܸfy\$( "O&�S&V%e@��9���!` U��"O�I�����V�B�@CF���"O�0y�&Ogj��#�\$���e"O����-L#`=�{�A&\��"ObHH�� n�i����;�L,��"O���$��sk|ᩖ�ƫ?^�9JD"O`PtO��|'4;�� =cAiu"O��qT'/no��:��(@B� �"O�{#��:��-@��tXf�r'"OA(�   ��   �  >  �  �  8*  �5  $A  �L  X  �c  
o  z  s�  �  8�  #�  l�  ĥ  
�  J�  ��  �  ��  ��  F�  ��  J�  ��  ��  �  `�  ��  � - � � �# q* C3 �: �A �G N R  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#����!LO� ��!צ[�n�V��G!��~�҄�b"O�%��$Vݞ�x�` 7${l�"O������$|(�bE� ���`�"O�4;A��c���A1�R9�\+�"O��:�E�M�&���B��C�"O&��T�Z	/ �x O"g�<!z �'3&8lZ"i�L�V�У#��)!%`'VB�I�`$���(E%D���(H0�?�t��E_襲ү� �bEx7�ͣ �B䉙s��u�"ᖵ?�z�P�(c�h�'[ў�?�v�g���ԯ�J��xhsL8D���D�,{�TͣE���&�(��6D�����SƸ�6�f�8H*f2D�l:�ЧZeN9�2@�PpT@0D�n�X�\0*nJ��{�/4�4KbIߤ*�pQ�͔�-K��)�r�<%�1��E�o�%V��n��+�-��&��C��L���5�	-0.24D���%
.�����AG�R���-}A/�S�'}Ѡ(�qk��j�����R	al��d��)��  �d�jDeN�mFM�=��'���i�<�*E��#{N�Q�	�'� �,�x4��`(���^Đ�"OJ-��-��h,ч&�9`�n�¤�'-�O�y�JW�����w�b}PEM�+�y"挤$(��B���p�L1���^��y҆��!}���B�x����mÙ�y���l�f��wpu@�.A��ybD��~`h�� � �څ�F��y�X�\�j��#C�?�ج�Q�R �y�V\QR.�( B�TB.���y�aǟJ��R��#'ABX{��=�yr�L�o�8dpe�;!=�8�3�y�hө&�$�R���zt�����y��J�aA��b�<	u�Lh��H�y�+�9�4��D�X-��\Y6 ��y�)�mv�pr$q�M�U�^�y2d?��̨�G Р�)����y�Ǚ�hV,XLY�Pu2%��/�y�ʊ7S���c���޼)P@���y2��=`di�'MUy�V�ǥY��y�fT<a���Q��� �v���.=�y�J֜'�D�;e�� l�x�����]�<�#�:c���ۓnծI��M���i�<I`!�CC�="� 	4騜���o�<����7)"^�c����8Eok�<It��/NQ;Gi G�Z�k�P�<�hX9
Դ��P.Ż. Yy�#�J�<!�ŋ3��s-Az0�+�^`�<RMڤC|��'Δ ]沬iQI�_�<Y�e\�6�B5�w&�$W�$h����p�<ydiO5�d`VN֕$X��aF�T�<!C��K�fec�A
���AS�Ke�<���@�>���y�b՟P�|��F�F�<����	��������.m�3��w�<���	14��$C�k�2�b�cl�<Q#l,� �P#K�,eV�i�Kd�<v�!}	PV)�Y&�Ih�_�<�KU�3F��9�ޜv`���KL^�<�F�C���ڔ�.]Ʈh��nGZ�<����]��	3�Jۓsq��� �m�<�5 ��7�Nx�&Ï4&��b�Ǖm�<�`":._Zt�"!Ս0cV����o�<�Ɔ�*o'��z�*\/��1׉Ai�<� �	�����iR�JM�1��І"O��8&�?s7�����I��Lx0"O�rt�S Y*P�a��$M�Ms�"OPɘ6���^;d)ې��*Jp\`�"O�e�牂��^5;�I ���)�'��'���'vr�'��'���'�*��@
X�a}�(��MJ��j�Y��'��'�"�')��'k��'�B�'�@i��
�-���Kd�@~�@l�6�'���'���'�2�'��'���'�\��Ǟ3tK��ШV��i��'!��'�"�'k��']��'�b�'a��K2G�3e$���+�d� �c�';��'���'��'R��'��':�x�l`�.=��W�L�p���'�R�';b�'mb�'�b�'��'�R��tOF
z	��
���i��'�B�'U��'���'?��'�B�'�H����ܠ4V�}���
t�>�RW�'���'���'M��'b�'���'��Z��Q bVb���Ȍ�qn�[��'h�'uB�'y��'���'{B�'f��ZE�[�m��12Uf�g`A���'+��'~R�'o��'�2�'j"�'%S��?c�\RtIץp��q
2�'��'�R�'t�'��'���'
��:c�Rє��ɖ1F8aY��'.��'C2�'���'���'L2�' $X����7M�8�cûΜ�0�' �'K"�'�R�'��HcӮ�D�O���!j��EGV$�b�*T!���,F~y��'��)�3?��i��$
�.66�ҍJ��/w#8M��e:����䦉�?��<��:��Q�G 5/����9#�^�����?����M��O�����K?Aj�N"a�PYp����P3��K��1��埬�'��>IS5�>/� ���<3�<)�'%�M�`̓��O!�6=�tip��.�1����t��装M�Oh��~��֧�O�q�d�i��Q�?���z����H:�D�{��Dk��3��J�=ͧ�?�v�Z�8����k�4��q��)U�<�+Oz�Ol�oZ	,�c��r�eW�4�r0�3��[,6��q�Pm�:�I֟0���<��O�p�T/�0Wa�l�%�*|��t����x�I�D�4�`�.�S���'7��	��4(�udV�y2_WZ(�@_�4�'[��9O��õ�N�b��9��4;H8��c0O`�nZv��0���4��բD��!s�	��ъ	^J�%0O��d�O0��OG�73?��O�@��9E�n=BG	����@i(i.�hYL>����?ͧ�?)���?����?�2)
�S7�+�`R��"�Z�i�%���.6BP��k�h���O��oz>��>6��p���_�M`D��3xTx�	�����I4�Mk��i7m� y 4�'�B��yϺ|P�SWp�5k��I�L���,J�K�T%A��S;�p�to_ 9ʺ�\wI^O ��'�:�3D�.	�:��o �����'g2�'�����U�@��4]�D��V��9����V����� �;�0h�@��dE~y��'��j�LL�"n@�v�e��N=%��]��Q�;�>6M!?�w:P�������'��{�F��Vqɤ�ϸ��YQ5��<���?����?����?��T&��=���0⮟�]��L0�f�7Yg��'��eӄ��4;������%'�PB4o����c��U�j
!�n�%�ēԛ��g��IA�3�7:?��(͖R����"��Y���K�i�`��|ɕ��O��O>�-O����O����O��q�摿����7�Hz� E#{"�'��ɒ�M5O��D�O�'B3SB��LI94C6X��'�b�R7�&�o�Ȝ$��
���9T�/FS 13��_�P��`ɚ2i:$�4E ��4�����4ΒO)Ū�6]�`2�#ίd���sB��OP�D�O���O1��ʓe����8�=��e�b;X� �(�&?��ɀ��']��t���`-O�7��$$���8t�>͂Ԫ���l��M�e�^*�M��O(�C��Ը����<y�=4����bJ�)
�����S�<Q+O*��O"�d�O����O�ʧ(/�,A�n
�a�T�.G�o�Pt��i`�|��'�2�'R�O�Bgu��ȉ|��a�̇]}���
�lڨ�M��x����^.%u�v?O�p�Uf�>	�4� 昘5��$=O>�C�ΐ��?q�O"���<���?���1�hzR(ϊ2xZ�kݲ�?����?�������ߦ5�PCELy��'����hReSn�CC�;O��`Rv�|��'��v��6�f�p`$��{a�۝x<��wk��"�0��+?酯�o=������'a>��d��?Q�A��+W����p6���Ȃ��?���?	��?Q����Od)��ۭ^��ȃ�M<1֌B��O8�oZ�P5���џd�4���yG���B���m�*{;ZA����yb�x��inZ��M[��M��Oz�R&����_w���{�R:�M�6O���y��=�Ļ<a��?!���?����?Yf@ႁ�T���R����U� <Y/O�Qo�hk>��'����'.P�¤�.�
Dp0�N,Lg�����>9���?)K>�|j���ki6#�Z�
4�Ӧ!G�ZN��&����1�F1���M|ƒOB˓|h��b%�Y8���E��
趥����?i��?Q��|�+O��n�$>�P��I�k=�"��ҡLY0qb8��ǀ�O<9nZR�����*�M��iV�7M��:�S�
�g��`Z�c����E�k�x�s�
�K��� �H~
�{�? �=`sl�z�v��  �n<�dЃ4Ot���Or���O����O�?�҄��3���C�ޘ%N�)���0�����(�4�O\�7�$��ԡ2��)	�����˧~J�Ot���O�I�U��6-2?��ĩ��BΙtM�h���3��1f�:�?��!�ľ<q��Ϡv��L�kςAW�@�4�O��l/(��	�	�h��A�$Hϯ �2̠�E�26F��fBL1����I}b�'��|ʟ�i1t͉9_w4=ZF N���!�m�n��e�F�ã`xr��|Z���O��K>Yt�U&3N�� �/A%� ��n<i��i�.p�r�D���cq�X=XR��ǲ/S�'��7m'������O�� `G 6�V�i`-Ʉx+��Or���Ԋ�ش����l��F�|$S(O���$�C�)��'-ڋmݺ)09O<���=ie��h���� �WA,x��ԝuț��q��'Q����Φ�9C�xD�4)�.;��5'�L��:ܴX��F�+��)t!�6mb�H�P��Gt�A3!I+њKE�l�@y䎝��B��b�sy��'ar��g��h��O�9 eJ}���̂B���'�b�'k�	��M��lY�?y��?q��*T���ُmހ"�L��'o��j�&K�O�O� QaR	���siU<O� \
s��(�s�%'����fE�ӣ%�fAן�r��ǐ#7,�Krd�l�I������	��IɟPF�D�'�L���[�0ؑU�X	{��
��'6|6�#���$�Opl�O�Ӽ#�DY�n��	Jv+�d(^�/x}ϓ~����vӖ�lZj�oZk~�LEw!D��ӳh9�b��K�V�2S@ҼmT��7�|P��Iޟ��ǟ\�Iן|lD�u�UZ�� )���wy2�d�d�.�O����O �?���_��]�!ږX��yr�����O6��JP�)�Ӽ,&Y�KG)}w<0فc/�HAj��K���?^ԑ
�
�Ot!M>!,Op鹦J��7X!��
#�����O��O��D�O�<�!�'������8B>�R��C��0էܹF9�Q̓VE���ĀS}�'-�ghӀ�X�VA�.,��σ�D���@.PN87m=?G`	9*!���1�S��)��Í2
��PRjX"/��R��w�,��⟬��柠�	����j���|S�U��)n�XmC�	4�?���?�t�'��Dk/O��o�f�y���23.��bd��A�[��y�O<��i�6=��	�rcaӜ�
�}qq��#!]�����R��<����eb��ѥ����4���D�O��d�.V�p�ڗ@�~ĺ-�!��������O��mě6cҾnh�	��|�O���!֢���$L�|�0�@�'&"��>����?!I>�O�ְ�o̚n�!u Kr��*�j�-^���9ׄPlO�i>����'G�$��A�/(>��7�X�)�cER�����ş�����b>��'��6M>�<,��7�.l���Ԫ��i���<��i��O6l�'��6!�
J7�r�I�W��Ӧ��t�6�Gæ�]̦��'<�s��?����I A�%G�1P���,��P4O���?A���?)��?�����I�,X[,���-�$Nz)䋓�/.X���2T�����O ��=�9On�lz�=��M�H䅀m��z\Xu�����@�I���Ş�8�k�4�y��	Gs\3sL�A�N�S�f��y�U'3�0��	>Uj�'��i>�IEJ��R
�<���!N��6P�	ܟ�����'6:�d��<�"�'X��˃v0�����U74�X�Bj�$.�O`�'���'�O��Y�
 A?$٠7����)V��D��j�I�i�,+�S	NR,�ݟxrq떥A5����KYz����I�p��� ����PG��w�İ	s�A�Nq�2��'l�̝c�'��6-�)HQ��i��4���)��>�v��`]�X9�;O����O��d C��7M,?��M]�P��gP��rG$m;���P�3W���*<��<���?���?����?9��hz����@.�4�#�D��Ă��9 ���ޟ��IΟl%?牺w���{��;(�,�W�Gr�!�O�d�OޒO1�f �@�����cSA�q�d�[��)8>�'̣<�q.�~���䟰����d�g=zYbC��#�,��d#�"˸�d�O2�$�O��4��˓(�e�-ەOg�2V'�x�$�zqj�2�y��⟬�O�Ml�!�M���i��\��R�8"���W-<�<Y@�k�*��֐���	",��$�)��֕󆊨v*��رN�:Oy��r3O��$�O��$�OV���Or�?%R��\� �J5LޡbթE�����I� �۴&־�'�?1��i��'�v,F�Ю;l��);*D���M'�$�OF7=�f�tDg�X�i;��2n�;F�ඁ�Kh���F�"�h�Ā�����4���D�O �D�?h�le�!J��3�ư_����O��8��V�Ӣ{��'�2S>�3�b[X�R���#�)h{$9�bC??	�Y���	ӟ�M<�O��Ā0��h�bAX�k�?��Z����l�/և��4������z�ON0�����p˂�+�ʈk|!�ƃ�O��D�O����O1��ʓ0��蛯D@L��ʂ�7HD8��֦�x�C�Q��Kٴ��'DDꓔ?�4c��":1��Y3x����E��?i��ix� +�i=���ǘ%J��O��g�? �a!O�A�����{�@�&>O�ʓ�?a��?���?����:�P0eC�0�B�YS[��T�n!R��|�	ȟT��Y�s�������BO�FtF'�9�d�15�޲�?i����S�';�.=�ܴ�y2�з�<A���m�X�C �yR�M��d��
1M�'�	ӟ`���`����Ƅ8��J8/NB���ʟ���'l���(1R�'k"�^/�xTZV�$�TW�	�:��?�Q���Iş�&����Q���ȓx����1?�IH�53���i<��'>1��$��?�m�0�Z��҃�^
�� c;�?)���?���?)��9煮� * ���,ۧ�ݕx"V[��O�hmZ�q����'�X7�(�i�I�S�T,#����b��#Ev<�3n����џ ��)!`�l�v~Zwvl�C�O�N�ᄥG<�Zl��A�P��n�L�Ry2�'���'s�'
�FҴ;>���V3P$ ����!eH�"�M#E���?i���?qN~b�]�B��f��\T2 ��p���X���4C ��A3���rުH8��K�"��q�c�.�a����*�	l�Y�Fd�ON �J>�.O��b���P�@��X�N��.�O�$�O���O�<!��i�*Q
G�'s�)�7Ƀ4^2�j6õYr��&�'4*6�*��'��$�O�7�������l��x��X�(��ʲ�Z�	��1m�K~+K�k�z��%)�O��F�(!����`G�e��$A3 T	�y��'-2�'%B�'����jب<�/�5ky���%n�n��O��$�� �r>E����MsN>13ER0?�v�!���%j�c�F 2Q�'$r���t��&����� X�d�x���JC�+��`6F-9e��J�h��my2�'w��'�	�`]�Q�DfV3ۮ���)K���'_�ɷ�M;��$�'�RY>�6���I��g5k>(��/1?��Q����ԟH$��&��A��:D�����9�IyB�l@�UPB��'��4��	��.�:�Od��ψ�o	z}s`��  �q�C�O����O ���O1�`�zO����eR��x3Q�F��`�g��J�(-Q�'�B�h�4�<j�O��~�X�ń�)Aڨ bt�^�i@��ͦ�YA��ڦm�'�h�c�T�?���q5�ח/.)i��CSɒغ"5Ox˓�?Y���?����?�������5{J`��D/�,S*�r �£�dnA�����d�	F��_���w:�<#7�)e�=����&HP`���'�r�|��jfD��6OL]S��N(d@ L��`NM�|գ�0O섒�@�?��>���<���?��%��qT!�4�\�4r�����$�?���?�����Ʀ�:��]ܟ\��Οt� �!���%�<O#�-�Og�P���П�n�<��Tڽ���_.ͬ��$$�3%`��'X�1�!³o8�z"��@��z��'�,x0lκ.��}� �b�X{�'���'*��'��>!�	�t6�U�ٳ;T%�5��r�б�I��M�@�ʪ�?���E6�V�4�6����R�r�j�Ҳ��.J�E�E=O�oZ��M����E'��M��O��R�Ę�����M&$5��M�gh�تa�ɷ."h�O�ʓ�?A��?���?y�!Ƣ`霓><�e�qMӏvGX�:+Ov�mڣ!�|���؟���^�؟̛���r`������*�6�z�����Ʀ�ڴW-���O��)�c�"v� ��%��2\*�w)�O��5.���C%\����D�X�O˓s�ℙ�돸��1k�N����L���?��?!��|�+O�n�H$����]����2�@?xϠ\wbʔ,�����M��ϫ>����?���a�0�BU(�4^*r(�Alڍ^����P��?�Ms�O~m���ګ�!�>�	��~$j_
t�
�ٰB�r@�0�;O����O��O�$�Or�?Up�i1�^���Ĵ
���5Zğ�Iߟ`��4�H�s�l�ߴ�������V4�8��sdP�q\ڠ*H>����?�'j60i�4����t���<wW>8�b@�Y3 M�a�ٟ)-$���������OD���O��$
�ϊQV��5�����7V����O,˓$����gWB�'q�P>�S�g�?w�J�M�X�����@.?� ^���4a��f/#�?�Bw��FzM��
ʳ8���D�/t��X��Rm�X��|����OX�pN>�Gn͇�ȱt�T�'"�=�F���?���?����?�|2+Ov�nڀk�ɱB>rO���Q�֯Ae|��%Kџ����M�R�>Y2�i���N�5Bl��`N(a�T���`�z�mZ�L�R(m�o~��ί5Dp�)a��	�Zd�$k&m�u��A�G`�z�	syb�'G"�'���'m"T>�Ed[5F��X�C�T��������M+��Ȝ�?����?q��D�v���tL�eyWBͬЈ��ҿ5k��$�O��&�b>�r�e���]��H�@ȃ
{����	bb`�;0<�G�OƐ(N>	(O�	�O�%c�/��qo�1� ٬<>���m�O��O��<i��i8>Q��'�r�'R|#�+�6+�d�����������zy�'��ƃ>��V E����/ɍ<�P @� ��#��I��(�h���B��'?�p��'G���I�]���d�M.����܌a��Ο�����It��y�Lx6`�a�-c�PɈ��ȻO����b!�w��O���L���?ͻ�$���]�b�D�C�
�ވ�~��VJc�$Yo���L�nZ]~b��t������� ~��s�?tFV!��2U�� �>���<����?q��?����?��H	�u`����?[/`2��P��d�����5$qyr�'R�O��S2��wЀA�6]:�M�yj��3��vLsӾ%�b>Z�k����+A	W!"�0�C	L�H�e��lyrg�0�$u�I�[��'��IJ3~�b�����T����$3$x������ß��i>A�'Ib6�Q�?�$��2p�6� L-ņ
����SҦ1�?�!T�(��ʦ)��4|�Ԑ�åͨ`u]!�����Z #H����;?)!�-v���I,�S��E ���15�$dyC.�< &��-i���ܟD�	ڟ��I�������J2z�t�j�!b^ĚQ`Ƨ�?	��?I�i�Π�dQ�dR�4������S���Aק,}hTi�x��oӴ�mz>Ya����=�'+>�(�}�2WY�t�Pa���)��<�7�'g<�&�(�����'�2�'�`�7���ڶ���ІvdxT0s�'*�_�����iZ��������Y�D-�N��uc�L�x�V�C�nȔ��LX}��'tB�8�?!x���F>��u�$n6��j�	˂*�����_���|�A��O.	�L>��% ��1�Q��D�������?����?i���?�|�-O4�mڐz`ȩ���&aE����sAn�!"Fܟd����M�ҍ�>��7���u5vf��EHX�;Fs�X6��+����̲���:��Ԝ~J&�=P�<���/Hv0���<)-O���O���O���Oʧ)&�<�)��d��@�GZK�����i��I���'���'T��y�`��nֶuy&�ذ�	�hLhb4���9�&io�,�M+��x���c�T���>O`� Ǥբt�ziiS�(��8O\-�ŏ�?���.�$�<�'�?�a�$4�â��S������?����?�����֦%�U �柌�	��am��[�n�ʂ�<��lr���o���˟t�������XB��8����n��%\H`�'sE�͇n�� ���EƟ� ��'�.��1�F��@S��T��M��'��'�b�'��>睷+Jp��sj�܄�$+vi�Omm�
g=�|�	��ڴ���y�K��RI
<FH_�Ș#�@��y��'��'Uv�Ѿi��i��"T��?*�e�e����G���8Zy
4L�0=�':��ğL���(�I����Ii�29��̕&u�HE�&j�޼�'�H7͑dl4���O��3���Q���(d+ݞA�v�N$xǰTC�O�n��M�$�x��Dl��@v�L��#F,��x)��^�� �4Z�t�C�L4zB�z��ty��M�q�E; %�{�����@��R�'n��'u�O/�	�M�7���?��j�0}V��: �K�]�s�&��?�ҵi�O�Y�'�x7��ۦecݴ7��`iB�� `ջ�O0)Ȫ)2�큐�M��O� {�(*����*�����9���/��, A[*`�|�JG=O����O���O��$�O��?i(G��t_TS��<cjSkƟ �I�����4{��iͧ�?��i��'�ޤ�KD)T�41�F��;gy<9B�-�\ݦe���|r���M�O�9;��!P"Pn�(�̈�w�́�B�
�?)�&�D�<����?���?�@��z��ܐ��1i��ʷ-ε�?������W�Dė���������O��`c6&�D>DȦ��R_`�S�O�Q�'�b�ia&�O��U�����^'7DF�u�R�?��X�݋/n-s�[by�O3X��	�o��'XJ�ʗjGl����&�ďRj͠b�'�b�'���O�則�M�`-�
wp�v��t�~�����vBz�`��?q�i�Oʕ�'��6��#�|��D"��1��Vz�lZ��MS�b��M;�O�tՄ͢����<��I�( ��*Y��,Ԉ�K �<1)O�D�O����O���O�˧F>$8���ڍL�L(��݇` Y�i���'�b�'��O�km��nD�:=~*�N�B�c��ÁSd����O�O1�
9��h�0�I�%��+�n�04�J@:b�X��扸r��US3�'���$�X�'<r�'_���`��$Q�0�i� N*5z��'\�'�R�hhڴ Y�`.O�����)���g���{��� ��W���O���p}B�'�ҕ|Ҭ�1P�4Y�ЍB�o�&�B�ρ����9ߘ�;r���?
������?���Ȓ1�R;ab�}���#FJ�!�$���f9KpG�9{��� �ڜ3�Z�d�	�����P����M���w-aL����" J=u8`���'c�i�@6m�7�+?!:3x�ɑ2ˆd��ָ%}�e��;h| zI>�*O\�?��l�G�D�5&T\8h�q��G~��e�0��WN�Of�d�Op�?�d��&V?�uY�$]�zz����#�6��D�O�7MD|�)�)��D�[��\�z�����T²a�a��07M|�|�f�	�O�4�O>9.O0K�b�e�8թc��0N���Q��Od�d�Oz�D�O�<��ih�u�'� �3��
inN`$�%F�P���'X�6�-�ɼ��DH����M�C��DԌ`a"�R���]�5���4���_�2e����$�ғ���ným���5�D4ݨ�Ss�-N�$�O4�D�O����O��d"�S4|��$Ѵ���!���;�U��ӟL��=�M����|r��Y#��|([L��U��f�Nb�y؀/M�-��O��o6�?���F(X�lx~B([4̀ � B�H�w�JP�	�3rJ�TgJ��?��-��<i���?��?�H�&�b���_i�p�(���?�����U���ߟ��I����OI"и��<�fy0d�� s�$+�O���'C"�'"ɧ�i�1!U�Փ�T���5�����SV��X��H���<�'/
�� ��\���{��L�x�28��S�F)hx#���?i��?Y�S�'�������l�>	l2p3��Hq��Il�+Z���'�67m,������O L��� G��c��,�h�Cd�O�$�l�7�=?�;G��[�')��˓
r��`�l:iV�3)�yx̓����O����O����O&�$�|R��dy6) @$��AQʝsr��*F��+
� ��П$'?!��4�M�;���t�rL�!�oP< |����?�I>�|��"�+�Mk�'�^��caW�b�
T83.�?�:xȝ'v�*��ğ@�|�\���I����i" ���C�M�Q��
B�ӟt�	ß��	gy��a�X�C�F�<�?�rtb�&�D����ҧ�#>�p�K>��p��	��MC0�iP�O:쩖�ҤV1�Y!�D1(N y��ZK��tW�|�6e�U��4uPbeǟ,���	�6|z����'j��X�g����d��ϟ������F��w���U�ڸ~Y6�Bq��!E�q8��'�27-Ŭv)f���O��m�d�i>睔�@b��ߟy�H\� �[q<�	ԟ��I՟T2�����A�u��Zv��͇Z�����j�6Ǆ /oFX%��'W��'R�'�2�'��;���V^�Cu������F]�`�ٴ3�di����?1���'�?���n.��p#Z�0Z��F-�t�	�MQ�iЬO1�-��ǛLA��XWJƅ�xE��� _2����â<��Vr�$S�������j�p]��j	�/�p��IH&B{��d�O����O��4� ˓ *�&C*=rb�?!�d3s���V�|���#�y�#g���L��ONem��?1ܴ^��})���y�<� ��B|Ш����M3�O �����:��/���﨡S�'L���	�(��� �c�=O2�$�O���O:���O^�?��qE�uXE���;FYR�s�����T�I矸�4"=���O:67M5��P'V՜`@�a�O�h�@b�}&�T�޴C��O����i3�I�N6�=�thS2]�����T��̐��^�M�b��O�Idy��'#��'����"";��)��Q
SB"����ܫo���'�I��M��T��?1���?A*��Ha@	�;*bpi��95�[��h��O~	o�?�K<�O>��#U�/������F�%��Xʥ��R��H��K�&��i>%K��'"��&��*��
i���³'��//��z�dV��L�����I�b>��'�6M86�P}pG\u,JI��iʼ7PT �!��O��d@��I�?A%]�(��(�0T�C�S)/8�i�f�%1~��ş�BҦ¦��u�S,~(�f�wyB
�z���υs����(�0�y�P���	�8�	ğ�	ٟЖO�vm�A­,�{1dD<@x�P)c�~Ӹ�a���O����OD���dZߦ�]���Ap`��V�s��N!!�`������H<�|b����Mc�'~�@r��R,�VM��`_�}[�xZ�'�.���(��hۧ�|�X���ٟt0�/�!g]�hTh�)��	�E ɟ|�Iϟ�	~y�p�ʼ�& �O���O(�:U��hJm�'��*C���" 2�	�����O���v�	Ez��4+�� ��5� e�����v�["�]%<e�|�.�O"e���.�Ee^�d��˗f�s��)@��?���?����h�`��Cs��(����+�Pi����
$�D�� ���jyR�f�H���?>Gz��v�E�Q�T��阜m��	#�M� �iݨ6]�*7-(?�F�13��	I�I0��kFi�#7v��ǅW�]����L>)/O���O����O6��ON������P����6"� ;�
!�b�<�iri��'���'��O����1 �5�@�8s&q0�7U˓�?�����S�S�]l���3/ͺ��i�� ?�9Q�L�?�*��'|�z7��̫��|rU����#��9���Śt � ��S��I���ǟ�Oyr�t�|:���O�',=���iv>cn.P����O��lZ]�u ����M�q�'F�挞�k�(Ak���6T~Ei��ڍf�(�'�iQ���k��]���O�Z�$?1���v��|ڗ)�7��#��Ү;H�����I��t������C�'AꚈib&��+̘�Ia��"B�P��?���2�F`����'��7�-�dȧ"6,�!��-RI�aS%A�{��t&�d�I���S '��lZM~r��7��联C�$B*^Ay��74M��kJߟX"�|�[����ퟀ�I�d ���,�E�$�(8<�w&�ßX�	Qy� w�\��e��O����O��'oJ����9_ڌ��n��;c���'����?���zA����I�h,�E�v�[<CX��(/��tYĂE�
fչ��S�e���B�#�t�A�
��W|fT�B�7��Q�	۟��	�4�)�cy�i��PpW"H^�0r!�.0澕r��ۖ(�v�;������n}��'2���V#ǻM�����4�$�'�'=p6-̄$�6�"?�֦����*���F:LB���PɁ�Ts1���5�yT���I۟��I؟��ԟ|�OcD(z�'�H�c(�>^�VjW�m�F�
��O ���Oޒ��D��݌NwMq�5�I�&N�<v�������x%�b>ᣀ.��u�S�? n��p�Ⱦ��i�#�A$�d��<O��+e(6�?�g$�d�<��?)��p�~��6��|R�y���?���?A�����^𦑹B`��8�I��p��O��li1AܝO�"�Ұ
�L��	��M���iu:Oʕ�fD�ژ-:��ѽ, <Ԋ��� [�-�40��E��k��57����ɜ,8��5`�� 7���4jRҟ0�	Ο����E���'���HE!1S,���F97?��j��'��6mXh�����Ov�m�s�Ӽ�T)�Y�u����4$�H�JuG�<���?r�iW��i\���2��W����&7>	��.�70�	O� (T1O>�,O��O���O����O���� ӊ`����a;D�"EZ$G�<��iS�}�T�'aB�'��O`�	-�i�t�
h�e*�T' 4V듣?A����S�'m��\W/�,\���`��T��`RWꍾH�v9�/O
HRh�)�?��,7�Ŀ<qF�)Ox�[��9h� ��&O�?9���?q��?�'�����a�3�A�`؇F1Mr�����D��0IvD�Ɵ��ٴ��'�p��?a�	����= p��D��i�DK&�X"��C�i��I�vT8zw�O q�<��B���%��8�B:ъ�$�OJ���O����O���#�ӹc� K��֌+�c��PP&��Iޟ��ɠ�M����D�Te��O�p�ï�-0ڄ]��(�:{�ؠtb�W�I��M[D��i��M��O�p��/ڈu?L��씜CVX�U�
i�� ���ܓO�˓�?9���?a��X#�iWIO8&�$ԋ�	��-W�a���?�*O:dl�t�4��ԟ��	T�����	zv��lѾ���"�����c}�fq�84�	x�)B��\pXI�d�Y�"t��gAR&	�$U�H�vf�%k(O�)��?q��(�$
0����$�Xf�<"�ϛ(0*�d�O��$�O���ɦ<�`�iR��z�ʎ$fd�)z2&�� �V���Y9�R�'��63�ɛ��D��(d�9{i���n�9<��P��M3G�iU�}��i���8z��r�O��-�'i��`�]"\'�չUʠmߒ���'��	şL��ҟ�	��`�	�����P��g�RyrX�5"ՙg�6��:{����O^�d(���O�nz�Y�֖^�*�ЌQ3m�$i�����M�ûi�O1�v���Jl�@牭{x���A�$EU@ KԈQb^�I��=J��'�D�%�4�'ir�'�Lx9B��q�L	ӓB��xaJD��'%�'"U����4 2�����?���	��V(��d�Q�b�1�d����>�B�i�7]K�I�t�(�آn$���P�g��'C�
H�����I�%O���K~"�m�O�����s��Al�#�P�&��NX,����?���?q���h�����7o��<�aE��/tt���%S�@�G�)���Οx�Ɂ�M���wsXZ@ν���A�%ֹf��'��6��զq�ݴ6��Jش��ˬ>��!��I��r$�C!f<�rD�<����"$��<��?Q���?����?y% V�VLؘ5h'rXS�\��^�93G�؟\�Iǟ�&?Y�Id)�U2����œ�A]��˩OҕmZ��M�x����½;�Ѡ��0�*h("�X�J^���Zd�剥c�*	�s�'4�m&� �'G
� ���?\�x����$@SyRR�'|��'�"����T���4m�-)��#�r ��#n�6����w�h!1��#{����\}��kӞAn�M+S�
�z�B��'��
GS���A�PR"�Iܴ��� `����'9d������v4�i��K�^���F�8���O:���O�D�O���3�S8n�E��I]t��	�c�$#Ѝ�'!�i�hh{�>�����˦�$����C/(@`��&[|���\.�䓈?���|z�M���MS�O~���!I1j�b��O�^u� c(؝"֪���)��O���?���?!�k��jvaЫp�Ȩ�F*�?D,a;��?�.Op(l�F�b��I��\�	_��(�#�z C�DP.*��뒍ΰ��$\b}��n���lZ���S���V.��У��p�����\�ڹc�O�� �-@RT��ӹ e� �C�	#F���%$�7K���1�\�Mh�D�I��I� �)�~y�Lx�f��	��R�"�nɂu�|;�fH�j�H���O�lV�#����(g�+
�ȐѰ��W���A"��쟸�I�>��mZg~Zw������O���'�B�2S'��UZ(��&�'m$�B�'v�Iڟ��	�����ğ���X���ĞhC�0�`�Hf>[fG�D��6mD�m��D�O���7�9O��lz�q�C��uڞ�2($ S���uo�ɟ(��n�)��-S��n��<�c�<�:��V�J~hBQ�]�<!��Hd'��d5����$�On�$@���E�/� h�-�M�����O����OʓTn� ��?	���?a��ʕf�������:��܈����'t듖?���>��'�!�1�=j-p��IE�#����O\��%��)SPK��i��?1�,�O�XD+�6*,��ʾ[윍!"O��ū��U�C}��2�b��'��i�"l�r��OP�D���?�;��9@��y���@#I91L�$0��o�.�lZ�
�Pn�\~2�ƴr|�<�4�Z�K���22,n��#)�jl�m���|Y�(G���1�0�#��4�q�f% �����黎Ra՟<�	ğ���b�A�%�^�b�oQ�سԨټ~��	��M'�i�O1�ء	'� b�Ҡ��;Z80�5��9��Mƨv�˓5���L�O4�!L>/Oxu1 ��ӄ٘C�ؑ��HD�'�6��o�p�$�.]����ũ��:�Ҩx��,¤�$��-�?�Z���	ҟ@�	�`�i8�$ՏQ`��Y�_�Sf�p�c��U�'�>$��f��?	Iu����W�U���sad��uM��c6�֌5�`�ȷ	:Rn�&3p������b��p3�g��iu�`���ӆ!�0�6,5�@��ƪ�&��X��b'��!"$Jӥt�V���ʉ# �E3�9�V�0Qj�C47|@��fl��D J"a؎?34Ӄ��{�����:.�Xr F>+D0 �o��5�
�c݄k�T1�؎S2��� �!'|0�n5o���e��ج�#C��N�c��݄O
�x��@0����f�c#Гw�܅�LM{�7��'#�|�۴�?����?��#ܯ$~�On�$�����7m���������b��/�I�M��c�4�	���&�E��@�4ɘ&��^d��A�-��Y���$�f 	N<���?AK>�1')��X�nH�\� }��ђ�:��':��=����?�����ۓX��CՎ�`wl�!O83�]��M��Iڟ��x�	Zy��ƞe�Т��
uT���v~�p��y�'I��'��ɗ%Y:X��O�h ѦI��&5 D�@D�2+�(�O&�$�O֓O$�Eb�'(F�t.��U��,; �]�v���s�O���O2�D??�����ħ��!�bH����Y��.Q؜iKB�i�R�|�T��$�=�I�(zڐ��H�+5��!bU�YI57��O����<��bIn�O���OZ� µ�[� �ґU�7�T}���*��<)���f���)_�R��sV�C$�� �����P��iUGP��M[UZ?1���?��OHMu��"ň!J�W�Ƽ� �i��I	����?�g�%im���O-"���0V6MȒ�Ddo�ן���ş���:�ē�?�CN�A�(2t�ʶ	{�(qc1�v���O>	�	� �K�i�I�`�	㊏�@�$��ߴ�?)���?Q���{��'v��'�����	�v��!�(�&LJ%��ʱO���C�$�O����O$�à��k("��!;���ɦ��	�&��\+�}��'�ɧ5�#S	�����*f܎�h3jE�����(z
1O���O����<���\�ml�nM�g�Bu���� b��񘰐xb�'D2�|r[�ȊF�O\����-B�ĭI�f��&�c� �I��	]y2F�a�����BǗc����eT=G=ɗ#�>���?9K>�(O���\���"���a��"N,̤���>����?��?���t4p���?���@�V�ڤ�	�~�Ƥ�pƙ�Yt:!8`�i�Ҟ|b�'�b��7^�0�N<	�a�,����j='Ęp�զ�	̟�Iӟ��$C����џ<���?BSNG������Xpb�L��h�����?���01�L�I�S�T͞�M��؆�E�>�����ז�M[���?q mڑ�?Y��?	���)Ok�Z +eL����_�u�P�Z;f3�v�'��	8u)$"<%>��p$�:ྡ�'�	b<�0Յe��Q�P��O��$�O���J˓��)B�{�P��\�+6��:����Q�|��*9�S�'�?�0DJ�cTdR��F-}�M!��# ���'��'��I��h�>Y/OZ�������Ă �RU*��A��X��+b�ΓO����VD���<�	�4:a�
�|)FJ�	I�ZE�U�MS��;���qY�Д'�Ҝ|Zc�~@Rvb�0+b�b�V���H�O�msQ�6��O���O������AS*L�R46ϴnh������H��qy��'��'��'D�C��ƺK��A�5	NGw�\a�jv3�^���ៈ��{y��L�FEP擾!�� V�76��%����6M�<9�����?1�y�(�'�Ȉ[��$�����@����O`���O���<A�C͑j���[��6��A4��&`�h9f���M����䓴?��b��쀋{�)Z�t�ܸ���$�˵�
	�M����?Y)Ox���z���'�B�Omҥѳbޙ"�J��p���.����&n�>q��?���90��q)��Ix:�-�#'�0����5U�"���ߦa�'}��ӧ�x�����O����$ק5���8XE�$:�`S�[ބQ��͂�M��?��I���'�q�Ɣ���5Ng�i��) �m�D�R�ig4D���l�@���O����F��'�剳V�@�	(�:�����L��P �4��X�"���OnAx�!E(|~ �e�V�$뮴a��Ʀy�	����3���ڨO"��?��'T$ e)�*r! x�cMUs�a�}J��'�2�'�" �S5X����[obY�	NV�6��O�P[�͛l}2U���I�i�Y�ց��mZH��W�2�`�3�>!F
��䓖?A���?�/Oj����xB�)`b��3ކ��Y�����'��IҟX'��	ҟ���� �u�XQh��2���"ƚi?>@��Ny��'\r�':剤Ob`��O��qBeMG�4 ��K8C^\޴����O��O����O�7F��� �(�_�<Z�#U/�2�>���?Q����PTJ��&>!���{̻���>�6�&K.�M������$��L���D=�Ĩˇ��xk�U�D���
�^�Mk���?!(O@�[����@�s���D!�t�0A"��<d�)(e3�d�<���5�?I~��π <�Sr.�3we) � �4���ٶ�iK�ɝm �޴{��ٟ����d�Z`�`�LA+X�0}��Y9�V[� 3�aPğ|�K|�M~n�t)n=s2��l�h�i�A£1��6-�AO��$�O
�d�O��i�<�O(n���Ә]�v��&�P� 
���0�b���p���.1O?��Ԃ��,o:�Q&�/1�K��ݾ�MS��?9�ꬹ�/O�S^�D��2���ЭII]�A9�k�(4����<�@S�K����䵟0���X�q���-��5(@�\_�&�'�vѸ�U��Z��N�ૣ�Q��k�$��3~F�"�������_1A`
��D�Ob��?�5 vb�Dp���ft��Ic�B�lB��i/O��D�O0㟬�I�أlҾ:b����7cx��JC"z�P�I"?���?����䘄1����'m�]0��ڒ<�����Ε1�~L�'���'u�'��I�0�M�ɸ0@䡝�~�
 �D
[�(?�Eq�O ���O���<c�p��O� ���3dX�G�π!0�z��s� �$#�d�<)� ,�?�H?	IA��X�����o>x���u���$�<��q���.�n���OT��Ɗ)fLO
T+RɈ�V43�6��s�x�'g�K��:r��y���	�$��Y�$�C�j�*���#��i剆j�Bp��4S��S쟨����䕵h�<�kC�~�`���B- ��]�L17�����L|�O~nZJҾ`��!6�25'�]R7�ŗ�]��ԟ@�	�?YIN<�'h_��q2�n�+�N
�7#���i�j h��'h�V�4%?�9Ӹ��L�CA:�H���;*K��Y�i ��'��	&4*�)�N��Ҡ�U<�p-�'��-5D�i�n���':�}�3�.�I�O ��O��JԮ�3d�.*����x��G#�y��)"�U�H<�'�?�����3��YK� �,���(��97�o����IR��p$���	ןt�'�Z�⠥�y��Q	7 ��Y��B���\O.���O`��<����?�f�A�wN�y���$�𑁵�U6�����ON�D�O�˓0�䑁�П�h!@H�,�6�`��ȕl�����4���O�ʓ�?)��?q��<�B�߼}����Ή�1Y���ˀ⛖�'92�'��S�@;��"��)�O�r�ᇦ&2hHd���9���Ȧy��Iy��'���'$��y�}��OJ*�YYP���텂$ZՒ��4�?����D�~"]�O^2�'�����=F�f�����-h�}��Ƒ�skN��?I���?1��h~�V����G"� ���[��ق ���R�lZXyb���P-�7M�O����O,��v}Zw"h@"G�/]��1���j���ش�?���~�t�Fx��)޾-ڸ�'!��$�x�mT�, �f���"6-�O���O���D}"V�h�H�V|��Z6��ծ1��@߬�M����<Q�����*���DhƊ�x�VL�7C�"pyЃ�M;���?��v$�4"4_�L�'�r�OX�C�R/zutA�B+� )ZF�jýig�'�"@����I�OB���O��C�
.J�%�JT,S pJGO�-��Q�@i��O4˓�?I*O6����(���(m0u1s���* ę�X���'l����̟��������IyR!B�[H��4/� MĈ�g�]�V����>)*O�d�<!���?I��T�è�x��|�炏�v��XH�EX�<�/O����OF�D�<��"ǅ`\��8L4��u�4n��9��O�@C�6Y���	uy"�'���'AĐ��'�h��X�<
��ҡ#T�H�m�p.f�<�d�O����O��mm��&Z?��i��˖�P�T�*=��Q
�y��aӐ���<9��?I�u�ϓ�?�����q�(��tѓF670i9��i���'{剃 ��q������O|��W�~tp|�Շ`��Y�M=.���'���'�B*���y�'��TҦ,F�f�̩B�A�h��@��d�ۦ��'��<�obӠ��O����@ԧuw�
�x� �� %�:I�V�ђf��OP��
U���Yy��Ɇ�[.<J������l���7�ˎ$��o�ߟ|�	��������<y��B��L8�lL4I�Ʃk3�W!ϛ���y�Y���a���?	&�V�>:��E���7u��9R�HcR���'���'��a��#�>�-O,����L��_n:L�*�J�� �<���d����<�#L��<�O�B�'	��_�-w��ڇa��v���ä�3.�6��OPA Ů	p}bR�$��Wyr�5F�LL!��ſUn�$qEɇ��$W�4��O<�$�O��d�|�N��vKp�����Cj~D�#����Ny"�'6��Ο�������H;YhS��ү0�&�S�mǢ������������8�'B��1Ff>�S��r��i��"�6KF��'!�]����ퟀ��e}0�I�R�P�aP1��;a��9҂��4�?���?����8bl\��O�Zc����K�%��,�1�ŷ@��]�ٴ�?1-O����O���W&ft�;}�A� Nu�<ɖ��VXc�#G�Mc��?Y)O��(2k�g�4�'�B�O�8�1�M�[��}CW�R������>Q���?���.�j̓�?�)O��?V��CƊѽlV`]�AB��6�<��)A8_!���'��'�dD�>��i���P�˗.hfH���	n�ҟx��0?Z�I��$��˟��}��M6��h���":ܸ�d��;B�>�M��?�����R���'�\@�D���Lk��O�p�)��{�^da�3OڒO��?a�I�� �E��K@��v&�Oʴ1yU�i��'��"�&W������O��ɜR�%
��A?���"�!}K�7��O����OJQk@=O�s9oZ��h�I�dq��d��r7:Л'�]<b&|��4�?�%'��'=��'ɧ5�7
v�
7�G�i}H��������!:�<����?������ΠG��a�"��q[���'�,R8~Xa�W^��?iM>	���?I��I�u���?��tc��n�T����$�O0�d ����9jXΧV�)`��l�(*�
�sC>&�8�It�	�<��c��	#ѐ��giK32�̀d�ܽP����O���OJ�d�<)3U�m��O��)	vf��
�Z��`��� �����Oj��3�$�O��}_�0}�	>V�č ���QVt��.�M���?�(O*�9��k��۟t�:V!(�Ҕ�*Oy��)�P)�U�M<����?�B����?qM>��O�"|1a@�x%����@��YH�m��4��D�#۔�nZ���)�O�I�l~bGL�:�V�j�쇩z�;��6�Mc��?a��N��?�N>9��$�Ȏ"0R��ǜ x�P-��M�$�*w���'�b�'^���.�d�O~q���2 J�<T	�����`7-O'l3�D!��'���|Z��!4��AǄD�f�4�C"��M���?i��x=C��x��'S��O&�9t��Dr�:u*K�s� с�� 5;c1OD���O����h+��!cɷf�(a�\�'��Yn��B2n���'�җ|Zc8	C�K�#�ؘ��Ь/���O8�f��O`��?���?�-Od��2�!�J�0�/ǲM��	頹2�\�H<1��?1H>9���?)�d�-x��Be�5�t���\,y�v-Γ����Ol���O�ʓpi��p<��u��gf���E���D� 8c�Z�,����`&�(����<i�q��:�
�Vh�ы�¼
J����	���D�O��d�OZ�b��E�`��T�1Y4��f!�])�(X�ȋ%:�7�O�O�$�O���!%�I3,�����gX�3��p�3�K�b��6�O��$�<�4�Tu�OgR�O�����%G�6ͻE���p��s�)��O���F'2�$1�Ķ?URj�*CDV�SB� *�p89�f�H˓	_�T���ihj�'�?��E8�I)R~��阂U�4=�ѧ�?jV6m�O>��-T���-��|Z�'KrB�-�(�������;��y�4�AJS�i
��'c"�O�lb�BW�%���1�)��cB���5����M�N�<�N>a��D�'Ӗ�ї.Y�? �9�X��p��}�B���O$��0U�r�'��q�d�|Q�1Rdk��=�@�"�N)ZЛ��dt�Sӟl������0�Q��Cz*��$GL��M���޸�T�x�OuQ��0�m�$Y�\����M�4��i?���O�ʓ�?a���d�OP	A��Z'Jo���#	��9y��P��¼$���D�O&���O���:���O����.�T�趫�3��r��6MDj"��ҟ�����'gz���o>�B�h�:"�4����&�@����.��O��Or�$5�	�V����)�W��C���F����?���?)-O�����p�)vj����'c4�I�i��}lz�4�?aL>����?Y�%�k��@E��CJH�"x�C�E�"1oZ����	DyB/�cH�������`Ey�� 7�����
�,9c�l�	՟\��#:w4#<��Opj�cCHթ�N ���D�ag0��V (}�o�<��Қ��{�\��� �{L�\b��y��>- ř!!�?F}F���CQ$����!�f�Ô旎5!<�1�X6HQ�P�5RU9�RAV*��5@lӘ,_n�k�KЖ�P�b�+��]h�bˣp�,=ٱ!25��j؎ ��6N՜'��`�7���� aH���媃#��$�dJŢn7ء����a����D���{^Tl�Iݟ<��ɟ,�Xw�R�'�IR�"	�@�0�91-��4���ȆG�<C�D���΄�n�!������7ʓPTD�c�M�8�z���-��RT���RCE	��T�Po��_�"| �c�x�7�I��Y#��j��Ɇ�L8D��	�0<����O��=*OJ���� �~ဗ�e[�
C"OR�8�(w86�����/�X����v���I�<	�H\������kKV,+��.O�L�V��n��'r��'��J��'"1�r�2E-���ԍ�	q�v0˶�/u�8�Ӑ��+H���+<O�|rM0X�؜y�bL�6�[�ʕlG��G�nI���?<O̘���'{"��E�n���h��i�JU��JLm&ў�D�C W'�ɛ���gN�] ΂&�yR
�5R��%�^n��l�/�y�j�>i(O���T��B}��'���Z Z��F�B9a�d�
�%Fc��Jb��۟�����DE;��E��Q���2�S�tC[�7vI����)k1蝄�(O~���ֻ'm�ɱ��.���@���Ǘ 4h,9���/ ��2剚 � ���O�?��&�}|�9ʣ �b@��ne����I�1@�Iw@����ūn�*����R�.Y�D�8'i��&�
t�RL��7����*�h�O��d=��@ӟ�����pH��߾Q�����8V,���|�IbVO�1Bk�jd��?�O�1�
� �y�*��G�8�Q�H��8記�� � d7l^u�^=�HG  �&���hE�q�q����4�bH��
�
O����6!��K��'Cҗ�����O�Q��	�"+{�,��f�w���a"OHy��d�� ��S!���n�<���I8�HO�S*@��YbG��hx|�)D�R>P����Iן`3�1v�.��I�4�	�)Xw��'"�է;WܦL2Ԭ�<�8� �'}i�ţ�)Qۤ��$G+O�qۖ�ѻ�LI�&ɞb-�;��O~	����,Y�(�c
�A8��3.ގcO�쫢�N�L�#�ĵ� c���O&�$>ړ��d�*ȶ����\��e�Ƥ֮>�!�݈aD��Q�'�b� ��*.pGzʟ*˓)à�`%�i�^�Uh�PM�	͍���s��'�"�'�"��w���'r��+B�'��H��hA;1n@��T�<��uI�w�<dj�#٭��d��˖�Yz,�r�	/���0�O�D���'��J9�X5��Ȍ.i��z���:m�6��O˓�?i���S�t�jӶ}"�d��,Y�	!W��'�yҥ�mx"	�v�	�R*��A��:�y��mӦ5may䉍~>�7M�O���|:��^�=����#��>`�j|xJU�?*T����?�/����iv�'_哖-6����IX�i��)ha,�:D�<�"e�A��4§)b�k�����C�(�df@Dyr&ā�?���iT�7m�O�˧"$epd�|���ED�-Tn=h�������Ğ�_�@Q�/UJ�.��d�������A{ش�?�a��-O��ed��:�JL�����<����\G
���?+�t}�c�OZ���OdL	�ސ
�i8�k�=��H�H�t�ݨ�Q[�|����Cz.A3A��H�i�!�A!uL�9���/*�|���|���'?�Kq��OH���i��6��l#���r�'���';?�$�4��e�CKP6�ڼ@VD_����O8���s@���x6 	�M��c��J���?�bA�F64Z2����|d|I�S�ݟ4��r���J7������I�h�I�u��'3"��I��X�@L*{F�j�.\�G\t��G.:���F�H&P��y��hO+B�X?,"2d������2����O\�.�� K��p���xh��%�ZID��#|����n�"��c؞d��	E�W�L��::��xs�a$D�,��P>R~��� ��2Q���� �HO�	?���Hh��m�>WjI  cN�c��x`b�H�[`���Iɟ��ß�0u�
������|Z�Eן���2rCx�
��,}��b�aS�[����dQ�{U�I�MB�M�f�[$T������`�������'��t�Ϗ)�$��f���X��'�� �(_֔ �qmǋ�J�I�'r6)rR��7G��pr�Y$�rHk�'�v6�(�S�O}Z$��O�1�T4@��2 
� ��'|<	��`XV��V�H'MF����'%4�)���X�M��ǝ.<ET�i�'gr�AlD&02(K�#�D+P��'J]��
F�&-�T�ٓe� A��'RyY`D4�rs40^ɼl�ʓQ�1���,yT�l� �[0xJ�y��]��@��
���P@�*(|l�ȓtzF�DD��PA�&1��ȓ�  "L�*i��d�4)Pqq�(��;�����0p�n� �	��4o��`r.�KX(����İEN>������@� �	0ѡ��)ȁ��X�t��ch�*�G��}Ot��ȓL��\I� Es�*�á�4d�`U�ȓ"�}�	$��̲B!�<�|��ȓ3��ŌF�\ z����ԅQ�8�ȓ�
H9Pe��)A��� N�>�r1�ȓ&���i�I5d@��.H:l=�p�ȓWb�yӥ#,a�R�Y ���A�e�<a�95��lp
_E���:��N�<�I�:F� Eŉ6��8�Aďn�<)�m��x�dȃCΞ�2ҁ�F�<���H>2����眡� �ab�Y�<a�O�l��N�?�(��oFT�<� �`��X��.���,+lD���"O2���H�7*P)�� xX��"O�d��!֏N�ȁ�Ԋ�| �i*2"Oj�9'"ϣ7�n}rah�$;H*dʁ"O���I�p -��� ,�%��y��)rv�KR	B$5ֲy���	�y��='�V�:�eP.;��7����y���sX�AC�� �腒�M
�y2K�5h�v(�� �E+�B^3�y�䏰r��T�g� +_>�J�և�yҪ�,#�0��@�
6A2�Z����y2ԇ(u�Ū�`b(9��# ;�y��Bk�@�HP	$:��X�M���y�g%��ˠ��|@e����yR�N�B��e�v�,R��\��yD�#��(pdF��PtrW ��y�N� gdQ��`����	��y򧔫v������/K�x�XqN�F�<�NC�DJ� ".�bX`, �Aj�<�'��f�$!�3�ْt���
�Q�<��&-���A��
g��DHp��P�<A��6f\���#b%\{��kgRq�<���F�?�6h���}�ze�j�<񂩀{4T�!i�~%��a��X�<�b�K?�� ␁=f���`D�y�<1 �Z���ʃ� ���qS�_n�<�&
�jf�]vKD�
����D�b�<	��Z�DZ uYi՛Z�V�XQG_`�<�L�,Ω��I�%d�<Y�j�F�<a2�ϾD�)8jM Lj��E�<96H�/_`���GM�6�����l�I�2����9Oba)  �1K_�zT�ͣ4�"��' rAi�`T:S��mc�)O#%:&��X�V�s�O^i��c��v��E����D�	�5�n`��
V̧]�IzqC_�	H\����=(�8�ȓ;L���O�ќYڃ#�4�*4�'�F������|������tw��/ ^,��A	�Y�!��03YD�{�#�'<�@E�7'J-Q��'�Pe�'K/U�ax���N��P�� c����?����l�H�!�z��j��a#p4S�nɄ�x2l�T�3�Ҵ'4,��Ti<�0<��F�e���<y��G�AK����C�h�A�ZU�<Ѫx��}i������UWfS�<�b�#o�R}�� ��t��iC�L�<��@;^�-��n�E��p1�	E�<YG�f�X�Z�� �L`��C\�<񵮞�)�.�Z&;�d�B�P�<ٰ�F�t�	�ufѧ��0`VFPJ�<����$!p��2��!ظ"OI[�<��o�s�`Ճ��[$�BP�Kn�<q�d��]�̈��PI
 BA�<i4		���|�����,�V��x�!�
�d�����+O�'�u��-M!��?!�rt��F�0殽��*-@!�d�Z�D�s�I��9s�IEC4!���|<u٥DF��Z�;��U�2!�d��s�����O�r�8� �ND�!�A ���T���x���*� ~H!���<���f���ju,��D���7!򄊯HZA��(�gfz�y�H�$�!�D�%,� ʅ�ӖlaxTE�5�!��@DV�e`v,Hq1�k�DҧC�!�_�~�D������Q��>p�!�d�#@����!��=:(9�ւ��Qm!�� �}����~�dUD�m0Z4Y�"Od	��8Gv`�͉� �~�`t"O�Y�e^�@E9��M�=�n���"Ox�������$eY�+��*y �K7"OTy�g�10�R��f�B-i9���"O
�pIݴ(�(c'�ʎOD@�ñ"O$���MR.r���0Θ'
���"O�Ic��ՑPZ�P[����!�� Q�b	��Dλ/|I����!�D�eq�PkQ�#j2���DӒ'B!�D�:{Wr��hF�*���-ւn>!�9o7�8�6����y��m��9!���^�~,���	AM�� 3����!�d�?��x��P�F���#�!��G?G�*<�Q�Z>���BG'�!��ȩ
6�T�>�H�1щM�q�!�d��(�0�c��X�x��?�!�d�V_����ϕq�q��F�k�!�D�ѫ3P�l�DQ! �Va!�U1 �1�`E�O�9R�F�+�!��72<x=0�nG��53J�d�!�ŧj"���"�6>�p-�N��P�ĥn2�g"0�9�g?�d ߯K���a�ѹk_�)��p�<�QML�'�rI��!�<�rdZg�ğ�;�)�6hB�p�'o���4��T����m^/L>Y��x��Ղ����yg�6J/68tÐ<�q��M�%�!�Z�'�����}�c�(c��O�Z�W�HG��{��	��P�"�# D�*5���"���	�!�$*���e�dU\l���7��:�HO>�h��Y��b�Ffʼ7�t�ID�rG�5�a�'�=ːN����"��g�1�}���'��Bk�(y6�8*��  ư	�FIS~�$k5I��<�a�G�i���0u팣��`P�]#^&�'��@��LA�O
��i�'�-�e�=0��4N�80��I�'���g.�_�TD����N�1dfA	��DU���Q[�Gn��c&�M����FUt�1�K
Dj� A�`9"ayb��T�EC��>�%`�4SMR	+fJD�BM��)F����f�Y
!EL�jR@Ёi12Ć�Ih��$)���8V�d���� v��1,��
�Al"����L<�N̦Q�\���̎F�ts1m��|��m	�'����b�M:�ܠ0�V)�����}�֌��q6BI'�h�Eﶟz4�~�)�1L��#�L�f�K�zQL �O)�5DQ;_}�2!��;Zt�$y!mֈ �(�O�%{%�O����π)��РO?版"�J5���X誠"�=N�?��"żn�0�a���� V���T"L ���F�g'L>���L����'�� ��'焱��ߨO�>�ya�Q�5��,��'�ꭺ��B�S���C�*g������� �:����5 �(A5OA�R7��{�9%�S
Op�;G�%��
D!T���@��S��R��0�@4����\p�]��S6��4XP����N��Ι&+`xY+�!��鶸�@�фF�a~RhC�h�$yA��=H&�Ȓ��06��!&�%s<���O0L�%O]�����ɐ��p�&դO4ݠcE�z���P�.�e�
�A��������䚦�K�"�(H����-���c��K\���)N�W�P`���Y?�za��mڝ�%{��'Ѣ��o.E�.\�Q��iW�5�'�����Ӈ�<�rMM#Q��c!8�]�W��#����+a*�x��XZ�Vm���	37o�!��2��yC�_ �����G0�p�@�l^�w�������@a9 �v�PG�]T+:�H +�7�DD��O�kz<����}r��Y��'��9�*�? YAS�E����yA!�?f�2�x�&��$�*|1���܃h���&B�&7����'}�+H�]9��;s�Єo�ɻW���Oh%�3#�1=�0ؔ�ڒU �q|�ړm�'s�^��#J�A��Dj3N$f|1��M+}"�1`�\�vc�@��	2�*�I.�)+tn�&H��牪ā����o�l�0`�)BƲ�)�E*Nr�((rb�>1��ӜO����t��&|��Z/D�8���'a:q��OF�<�Ĺe��]������hxd��%MQ�N
��g���$\>I���pTĐ^C`�λ]��%㕧S�a��Ҕ�'�DI�5#S�x��!��H����Q,D�g
H]�2��#��N�0E(#sAӈ�E� *
j��W�>��$X��d��ҒH��b�'W�$K��g5$AdJJ2A��[��Q��� ����� r��\Sbj�>b�h{�f���"�c�e&�|�'.���p<Y7�| jx��
�{K��;�`�͟�������Csg�0g-��fu8�����%�I�W.VݸS	�1u�%��Λ�k�^�z	�'�
��熔��t��� ��(Q�����(9�H��!LF��M3-� �3�6 �Z�Z�p�*�fE(�����I*���o�a� �̾|#����xu$)�N�! ��@����W8�0���(Jgd���P�~���W�'��,���Yn�3��+��T�'%�*<��	M�h��� L@�2@��V�B��&��x�N@A0��!H����ɘn� �	4D��0�VB"~Z���>Ә)������Vc��y���@��!��2,�)[����Hhq	c
r�DQK�>���Q��Wvp���I�G;v��ȓS�I��Ƅ"� �z���%s�D�n�i5ܙrE$�O��xce�<#]�q� C���8Z"O���@�4:,BCG�
I4x��"Oҩ���Z!H���A�l2��
�"O�h*$J�$�ء(�.əC�F�g"OX�b��/9zP;���;z�2���"OJa�'��Rv2�S��V�|�)V"O�-9 ��2��8E+�A�܀�5"O��&��;�8�P`�o���2V"O.(�q�C< �H`a�#H������"O���jM�G�ݐ �ЋT!�ӗ"ON�!@��rT����(; ��б"O������DCBd��΀8W���"O(��)L��� KA]Ӫ	�4"O u�Ƅ�sz^�0@jN#5kz��$"O����-Nf�ɩW�@�!�|�C�"O�����6n�~5#�f��Hp�c�"O>U�`o��p�VEЫd��1"O� �ă�,�#㮒�U�u�s"O�t���E�N�[��4!�@��"O������V4<ȅN38��0qa"Op�k6M�-J� ��B��s�X��7"O��u�@'Gh��r���C�ZMx�"Ory�e��1��5r`]�b�ԡ�"O��b���M�00��$f��p�"O>dK�dNt8���oU.H�<-��"OJ�b)��[�$8� )�PW8�bA"O`ă����
Z�eYg'@�^%�q"O�e����^�������;:
(*�"O��yD��|j���MZ�tZ8��"O�7�٦'2˒,Y�0:�"O�pI�NB,
v �`"��a~rA�"O*VH��������)S!Yk�<q�g�%��%�'X&��{��M�<iD��8I�H�#��D��!�&�M�<��F#(4�ӓ�[vh�K�<I�g�x��t�B �Y<�D��
I�<��T�Ew>\Q'�gDLU�Rl|�<!򧍴A� ��AH�%�&KJ�<��O�T��T�q/�؅���}�<�gN�j�h0���ϸ}��Ia�y�<yu��0(>@Q��>Iծ�aciFu�<�FEQ�Z`�T��g�%I���J�m�<�r,š:��h��CL-j"k�<�F�ܮC�@�����`��{�a�<a��S3�����i5p9[q��_�<��KI�nݦM0e��-6Ūdg�`�<�:p�0uwT� %��Z�<����|�)A���E�`t
��5D����Wh����}��=1�7D���̍;q�����_)���c8D�L:��I��(��#�3�V���*D�� ���L�9\*d��'��(�� ��"O |��Yk�a�`�:^2`�u"O~p���cI,{�oQ=Zt��"O����+G$�P��Ζ�<�,s�"O~$Pd��?���q%MZ�u�� �"O�"gg]b��Qc�MZ��!"Ox5Y��0���Yf�7Qj5{�"O`���=0G0RUi�#U�I��"O��P�H-U�����ǭHA���2"O@��d����H9�nˆd=L�)3"O �y#J��
��ૣ�.k3�(�"O���Dɛ�~�h�GB"w#�]�"O(;c7?��e�w�= �"O,@�B�Qc�H�F���@ɓ�"Op�2lˣU^�� �K�d�2�:S"O�Ȓ֠ۍ{���Be����p��"O@]P劍*p��)ꡪ
�?ڙˠ"Oޱ ��T��Q@Pd�$�"�"O��Ӧ��6s�(ѡ��H���ȅ"O�����N��*����Cy�!�V"O��2̏z�T���Aöwup}�G"OT����:\�%���>id�<��"Of�bA.I��m���H�Mm�\�"O4 ��!��MΨ�U�:iX��у�Op��D G^f\��'�,�c�:z�!�DX(7ᾬKa$�i޼�I��*>!�$�����ϐb�"�G�4!�$�L0�
 ۔4n���P��!�*;'�y�f���0���S��֌%�!�I#9<*�Ҵ�уN�����.�1�!���9�x@��ƻm����tc!�D�� D��Ib鞒���ۑ��(~�!���:>��$�;��ȓ��..�!�D�6��PA	�b�zTi�(jp!�^�\y�Ybs)���>�G_&nY!�$O?�AqRS7f��q�&@�.Y!�AQ"`��`dӳz��9Hp:!��Z��1H��<X�F�A�:!�ˬBx2DX���-`�E���")�!�D��f%���Q
46����]#�!��n���S$w)���S�Ip�!�$Z�:�P%bJM���5à�C�<�!��I(:F�p��P'*�]b��T�
�!�$�)��Q�6f�D9$Cٷ�!��?I�B�qB�|ڲu�)I!�D�;$j(m����<�(i�$"�bN!�D+e%:�#��	�h���bg/!�D�]��\�E�E�q,���&	L!��]=����Q��S&b<Ð���*!�w?��[ ��?h��������G !�Dd)�Uq�c�4� �)�kG�U!�d=��eȨ8�$Z3j�:V!�"�*� ыߩE>EQU(�6_!�Z�_�0�1Nkz�y����r�!���><�ASd�CD6���Ɖ+F!����5�pa��J�<UH$��	@!�dg;����I� �P��QdR/L�!��[��� ��y��h���-.���mݱ��R�OCő!)�9�y��
� z4ږ���TJ-Ʌ��1�yb-��cg���D��*$h��ir���yb���|K����j�$+���K�����y�oؕ`����
,-1F0#�3�y�m��	�\ xâ�2�ݘRb��p=ɏ}
� |�'�ؐ��l#�ٱ
G�!�"O�A8�n��o~$�9&�ɪg��4x�"O�Գ���s�\X��Lt�ł�"Ob�Jd��.2�<9���}g��A�"OZ�u�-�6T��ՀxVyA"O���ǋ
%a�mA���?-�Q��"O�IhY�����L�K��`x"O���e ��K_��R��*P�x9�"O��Q�ԧ�T$�aE9P~6<2F"O�qS4lZ$�~-� fz8\��"O@�I�1�9�v���m>���"O�U(C	)Gńqb����QU�!`S"O���a����A#����ճ�"O��R�hs*8�!i��*���u"O���@��Q���r�ū*bQ��"OFԛ���\�i�dLN�PASE"O.�gNƀfX��F�ϬM���"O$��DbF�=����'ϳ+  ��"O��bG\O�q�D�J�ze��"O@�a-�rvIYb�)����"O��	b�~k X#G��
'ѲY��"O�`�/��T.��8chU�%ꀔ��"O$
թS��>)h�!�,ָi�7���OIJ�*1e�/M�p��;^�Z z�'U���C������P�ң_���:�'N괸D,��q��%˗i�_�~(R��!�S��?�U�I�S�:}j��Y�=1#�	n?��]t��m�$dN�5�ʎ�za��	,�t:r��=�f\�vݳ�^H��CI�E�V�E4�#c����	�'�Ѕ3���MCj8"�X���k	�'�"�`�O},�+�)Z�OU���'��2&LA][L��Ƌ:Ju��:�'�l�p�	�^��;0�̖?�Ý'��R��lR���0��}(�b�1�y� A �t8��AIq���c"��,�y�$��ms�`�㋂o��HQ�`�3�y� �l>�jw Fj�vQ�&]��y��\�][�j¢�a(Ґ�m[�y"թ(p�ģT��-��DY��yb��f�p� ���*���ұ�y��ǇCH$0Q�ϊ3��H�E���y�#�?&k� е�3u�z��菀�y�Q�i�#r�'l �F��y"ԻK���p�b�4t�4QF Η�y��S0?攈ǎ�< ��1cdnF��y2Bc��UK��Y2#�ق��yb N*��y�3.a��#��S�P,�C�ɭ'B��S��C\@<<��oP�i�ZC�I�#h����ȝ����A�6�tC�	"xΥ�G�Jh8y��,�J.B�+]4ReP�b�9�ʀf�Q;"B�	1WvM�5�4��L�Td#J>���r؟�k6j�	C�̠���X�{Hl�$!,D�(H���#�8Q˕�>p�3`�)D��T��e���79��)�1�'D�<�0�����B�"E}��l
0� D�x�q,V�(pI�JĊ+u��95�>��MdJ����R�T�~�y`Gߑΰ��MpЌ���\�����0(ߎ����r�|���C�G+�	*�C_�v�1��dR�r��;%'�e1�X:\}�ȓv ��.�:1�$qQ�
L�\��K�'��I �c^��l���b2S��� (a��f�*k���&$ڱ%�(A"O�s��.$��#�=
:���"O�tX����(���ߗ9���<Oj�=E�dB�g��`	�AD��ٲ�͔�y2φ/]<�0��-1�\e˕����y"`�+B8pH#�0{�$h�@��y�./v%��k���36��#!@��yr�!6ߔ����Y#>���ה�y�o�e�>�z�b�� ��0���y2B]�4{�!��k	�:��a�Z��y��T�L�&<�������fė��y҉�4d����ª�lڤ��@6�y�b3OABd�RB�1j/f5A5���y��Q,ah$�bpa3,Ř		U��y�C�s� 1Y�./f*5�t�H�y¤ƊgGCBg�<+I���JM%�y�lR�S��B����8�!�X��y"N���z8��(L�,��I��y�.O��� �ޚ	Y�������yR`U f&�����*.bi j��y���r
<*TF�Ud����y2��y�L�W�Z�HV �L[�y�-�I�|�
��qDX� b
Ɂ�y�E۬7ꖑ� G��y���ש�y���3(��Y[�BR�4)�J�"�yblw3v�:􉒇>�0��$@��y�A�8s��DTNQ�2���� �>�y��W%=r ��ߛ+68�ŉ��yB���C���(����)�9�y��Cy ��� ��$
�@�T@�&�y��-Wn��C��VlF�� ^!�y�,�1X�@Hc�K
2=�P� ��y҅����u�	�"���*$�� �ybϞ�x�6}��l�>���f[��yRH�%��P���onu9aJ���yR�V~`�&�� /��}X�O]2�y�o��Q^��R�Eֲ:K�\�G��-�y�)	/�����*+�Td��T	�y��A���MSD��)���˰��y��T@��8�'#s�4�:E�]��y⢌�,��.�z��0I�E!�D�����b#�5�$�(��H�!��G#Ĉ��_!�*,��ҩ#�!���t�8]B���j��4+��]|�!���,!u�\r	̍P��b�b��!�Ė�I��i!h:z-N�����!�DW�iO� x��;"?��Y�Y�4!�d�WI6�S�d��J6�(
2���;'!�$�nB�y�1㔼`-D��sb�/!�D�_��)y��v����&˛�?@!��[%�r`��`�8}���	��Ղ9-!���1Z.�5a�!9��i5�ϵW!�Ij�E���3�Rx��CT�!��J$�0y&�G�`}�`���F2�!򤈝"����,L���u$
�d !��Gp#���u��:� �ţ�?�!��i!�Hif�{� �k�]�!��H5���'+��S�0�C��K�!��.�Pk1��.u%8y�_��!�$�?Ä����?����uωT�!�$^�3�V�qI*ц���Qq��,TA� �ʵCx8)PB�zJ���ȓ]r�L��˛A6�!��\ B*.���c�F�`�)�yR؆�ے4Hh��S�? .�5
�t�v���;� ���"On����Ն�ӱ��,��"OTh3c�Q���sV�(s��88a"OnD3����>���U��:D�YJ"O$la!cE�X����Bl�X�b"O�-���6!�d��.�m���"O:�DƗ`x��lJ,h�yq�"OB����[�p����E��=���"O҈��e^ޘ��Þ3���"O�s�KK�{����chP.m�J�`�"Oд��@Vh���sP�;&~��۳"O���g�8����&xc�H��"O^ʧ
�*WJa�Tb�#w-��څ"O�3C�ކu9P""�&exfh�`"On��A�G�q4T�x5a^���"O�<�q�î!�D�B� �Z�(�H�"OM���<�U��Ҁj��)�"O���W�7�E�"�i&����"O��j� �s�H��a�$20�W"Oj�@P
@�)��@W /hi"OX馤G$|D�����V��� "Ol���ò]׈�����
�@4"O{v�_�ML�1�'V�b<�"O�=� �%��P�C����"O>821(U01$��X�����ͺ�"Oh���G��:ULܯ]�>�y "OzɃe�F�?z��P��@/#\>���"O6���NA
;��Eqd�5ϖ�y���s�e�j��B�>��w�V�y��� �"�Ư�:#X8�+�yx~���^ܤ���H��yB�ݍ���Y0��Xd�ћ�N��y"��42z	yVFQ���1f�I��y�lX�&PD����,A��JҀ��y"e�8R�`qf]!K1��H�����y2(;r�ЁH&���I����l�.�y����J�~1��	=�~�����y")���@���H8 _�R���y"�V$s*��df^�r���[��A�y(�P2D�#� T"|@j��P�yfE=_�@���o�+8�B3L�y�A��D�,���ͼ��c���yBk[*t��u ����h21���yr��R����^�t���;�y��X��3�	����h�T0�yRɉ=���7M�t�$�{G���y��'��5��L�m���Hף	��y�����
ͤ\��qh�D;�y�l�;���!�_�<<Փum�y�
��.Q�҂~����3��:�y� �$*~e3�]5j����M��yr΅�,�����;h>�A[����Py�,N4h�:�P� �d,I(&�o�<YW&�v$4	��!YvP��&΍i�<1a憺N��) �N�E�$��Fd�m�<i�'��a� �1��*��N�<YA��F��	q��%��Q%"O���7�Z�hp���Ø0�@ya�"O�M2�a��k�2 z��@$,�@�"O�m+��AmAI�c��q術`"OtY��_��<q"��&u���W"OhQ	�K�XBt�6� p��1"O6X�$�}��5�f�ީ;XD��"O���6@J��HM���$>�ܠ"O� �D��f �-����Ũ\0V P|(2"O8Qs,���&�W�	�� "OB����ݾN(��Ɵ 5S�i��"O"���ŋ�Bv���C�͒4i�h��"O�4�'D�v���`��(0J|�"O,�X��F�,��yh��Zg5�"O�I:��J.�d):6l+o�i�"OvIY:a���
�@�Q��@1�"O���vA�	�4��
*M'�ݲv"O�4�����k8�,�@	T	D�u�V"OB0�kݞZ���:��]S�"�V"O�L�dB�,s�x"��`��Ѥ"O��A�̞�A6���R�ʵGʬ�ӡ"O(��deN�;B	�Q��1Z"�t1�"Or�8���|������P5i�� �"O�`q3�
��`��+d8u"O�|C1ǉ1FC�r��ՉU+�Th�"Ob�"�K� ���Q�,`�����"O�b��]�WĄ�@�R L���{�"O(��+ם[�X)X�Y��)�*O�m� ��|���2ю�,z b�'�H��½1NLȧ���F��'�,��.�!�r��v�)1�X�!�'���%��I0�Ц�ֶZT80
�'��6b�8�Z1v��a>�8	�'� W�0�
��5AF�Qn��'d��	 b#4҆ a��ǘGS����'��xcr�H<.w�L�L�(=� ��'�Lm*���[�BA�bd�$�(щ�'o\uY1i�mmRB'n!s	���y�IL��d@l��j`�2᫝��y�U��am���9�� 0�y2��!|lH���P%Cx!�1!���yb����P����4R��!�1Aϙ�y���rj�c��7��hj�!C��y���������*r�,S�l^��y���.���x��s�F��tbˉ�yRBY�AɃ�Kh�FM0�
���y�b�#���w)%vQ�	5#D/�yBfկ}��,�v��� ����y�h�L�R(a��X��Z��yB�DjT�"�*EF:0�+I��yRg7y���kQ�I4;���p��ybcȓ,d���,/g�3 �_��y��0�&��`7,:���%V
�y�J�C%TQ�3i�/(�(0��mÖ�y"H�<�Q	dˊ6'����9��O�"~
eOǸ�L���CM�8���]q�<y���^��y�ċ�	(��(y�^o�<ɣG�-N���[E	ˊaH��#�t�<aC䒡x^�M��CNRL`ԋ�H�<��?f�"�2�k�sr��%i�<1p�֨S�Dxۘ�(��EE	�y���!�"	idBhI	����y�
Ì)SP5��z�ʬ�d�ژ�y��[4�T��,�jx���)��yB��@�2��S-rs�i��M��y�,PW���4�X'YV`�{�։�y"A�#D���3cڗSO�]�g�G;�ya�e�,�"�i�>A��l&Ģ�yB#޵g������P�7�D #�!0�yn/(Ҩ��D70z�������?�
�',f�!T�Fhޥ%�E<okX�	�'��*��݆%��-JdO�k>��"��� .��Ő4Tr �����16Xc�"Ol�A$a)$�WF!ޥ��"O��R�E�RH�-"� -i��L"O�����B+/}\MÕ�$u�"O�al>gn8�1,��V�h�Ks"O�Py�&	0)�� 0��45j�q"O�ف+І6����Y��4"O���C��'?B00�jE&�8���"O�%�v���qi�g.n�h#"O�*��r�� k�^'�U�"O��!��́L�z���.4G��k�"OP}�smL4qɂp#���28��Z�"O��ӏ�7]� �]�8&��!"O4�p�A���)S�晭Y�����"Ob��N���Ɓ�!,�/9t�"O���rC�w��e��n_L�bB"O��j���V�v=c��Kf)�3"O�y�q�P%V��b��~��Dj�A ��ϟl��	2Fe0����ґE�tyԢQ�hJnB�	�Id�a8"�C�,�3bMZ/A�BB�	�'� &K%e��苲���@�6B�I2���!��=��x���<B@2B䉮0�"���b �=�T�!ˀ�"0B�I�%`�:cA�w� sf �Rb�C�	�O�A�HӞ=�D���h�*��C�	7?ި���ސe(s4㙚NRC�ɼK�����5��ɳ��@2:C�I�)p$3'�ÜX*�9���DQ�rB�	)����'��$�h��V�dB�I;*��r���`�"\*D�;{��B�ɝ0i�Dh�(C��SQ��"(�^B䉘h���PrƐ�����r�+rG`C䉵f��Bf�ͮ[.��d�J��XC�	�;dr033#_�~�d	�%�
~��C�ɦ<@z�R�S*�tiVjJ3��C�I� �@�B$�w�Y�S�M/v[�B������dL�g����熥��B�ɷ	~���Jǩov��Uh�(\AnB�	�K��������V�� ֲ;��C�I%V	h]ؐ�0#���q.�9�\C�+(e2�Jŋa�q��&��e C�2Dl�uE�
��E�"��:(�DB�! ��]�6A�<@�48��b-vB�I<2sBi���x�nh9��Y��B�	�^1�}��o^>&��3��+��B��7p�,�f�H2,��! Q��B�ɂL����2+Ƒ'{�=HW΍oi�B�ɒ<#�E��ļ-��8�.�;]��C�I�y�x�����3���b��)��B��	=���H�ɛ4Z�1�숟.�ZB�	%>K>��f��68ĥ�dAE;C\B�ɨC�XP��H�blv��@��C䉘B����C۲�T$"U[���� �d�]��YBʗS�N ��Ƹ-+bC�ɡ{�����ZH���6�Y-RC!��;����a���?��k%D!�$�n
�X%��&u��pe���!��8s�dL���N�C�U"�_�r!�$�$b[�Hc,c�	���y5!��L�P�f�acÉ<M��@�V� ��:OΥ�@�I� />����Mu�H8R'��F���(@�3�0�sAEn��A��"D��ʤ�ϲ�l�� ߟC�x�V�#D��:qh�<��أ!k]�E�)��3D�� &��C��_܂x�!n�,kS��Xd"O���$EU�F��U�@ tJi�"Ora�Q Y,��Z,ƂuG����'�ў"~��O<ZHDZu$�+Q� ��6����'�az2�H��Fl��G�JT�]s5���y����Ek��%�O�w殜�4hJ��y2��)^����c�{Q�I�åS��y����b9�#��,B\|Ȫ�"͸�y©ZD"�Е��1g�����y�Z�x�v�H*j6�P�F��y�JC�J��Q�Z5��Į�hOB����5�*y�m���A���#a!�{���2��6K��������!�d�>lR�*�h�0X��ƤC�!�$әo��A6[��ڰ�!�dF8#~���DR^���sh�0z�!�DJ2g��⁉V�d��psHFx�ў̆�	-������q���õ'�m�D�d;�S�O�����
�a���(�S�xj�m�"O���Z�r����ˁwX�t���Y�'y�$O�Bo:��DE�����ƣ��-��O셙A��`����+9�d"O2��H��	�
����?40b3"O�	[Mq)���)�� n����D�OJ���Q=A��`�7��E�T٩�۩�!�X�iu�0�!�a �C]�!�@�/g�p`��x\"��wC�,t��7O��@C�:~��8� �I'k3�MS�"O�8�2��r<����,S��۰"Ob-�h�4�i�CKL�"�8���"O���`d����
"�Yc��IJ>#q�)^g$���+��A`��`f	$D�0 ���+�|�T,\�" !F D����G�DJ���r��(\�T���=�O,�d	%,�����֔@��r%X����$#�����[GnUIB�	��p=;w$=D��z�3,�L90 ǻ_j|](w�9D��I�H[�-��!�ɝ�j��t�#D�<14��3w�6}�ר,	�ӂ0ړ�0<��噀V��E�r	�+C^� ��KQ�<A�O�ư���5�TPs(Jy��)�'/Vq� �$�Ḇ�E-��ɇ���ط�~�����i�Lm��&A��j� �,Uw�%@p�H��z�ȓp� 4)�B�#��#�F�_�4Ԇ��^,����Ȣ���Q+ Q(�	ڟ��'���>Q�+:<0�TϘ� J�_�<D���t/\ɩ��2A��w(^y2�)�'7� �q��:�@]Y4�=�Դ��o��I�4&T�p|�\�1I
:���ȓ*�|d��Ձf�>���)�h_Dԅ���q�2��6fV��P���/R@�ȓQ�$;G�_4�:PC%b�:p��'ў�|��
�<m� �!W�u2t1��,�n���0=�D���<n�h�V�ޔ~�:E�1@�l�<�ga�@C,�(s�F�Tٞ���Ng�<�a+ϱ?k"��(݄N�ʅ�c��c�<�7�/K���%oԿ]�ĐS&,H_�<�0���8%�B�&�(�a�FYyr�)ʧ>h�آ-�WҼ����!���$���I�Sܧzk�I�T�-~bLQ�G������4�5a��+.K@i��]�5p�T��^7�1�`j�.u<%� � .��$�ȓs\���.n��ӇU�V��!��S�? �����z�H����7/�xK"O�]q�M�x���5�h��g"O`���6#v%Ӄ���:�0�["Op]BԨҎYk�б6�FB&69�3"O$��bfT�t�x���<�D�IZ�87�&F�oX�vZ���#�R�<��� ==ڸ���`�<t�j�i�<1� \�R�`q���2r����F�^�<��Ƙ�1�z���M�g�ti���YD�<1�lާ5S*�"��#tIҵ;�P~�<Y��7HP䨥��enb�S�B�<��	@E X�q`�M�a���q��d�<A-�
�nEQ�(�V�<����Yl�<i�����0�����w�Q�<�$��,��Bڹc7�	`��N�<���_%B��c֦��	HAb��H�<a�$α8��V
�| \)I�aV�]�ID��t�����Œ���$(;�A��?D��Ղƛ.�l��ʖ/��E��<D�X�V�g�AX��z��A�Q�-D����66-X�K�Bӯf��e��6D� C����y��"5.�!/�!򤉚b�f�J��0m�&Zo0n_�O\�=��:)p�,�/*t���ΒiO��+��'�!�Dh� �d��&u�<�Q�CR�Q!򤂄 �Y�u%�2�r�U�zU!�$��L����)ިXkT���l�7!�$�2(�H(��M!]d���ю�Y2!�˨Qz���Z)K��1�-B��Py"��5[��m!�.�	M ��X��©�y�O9-V� �!M=l��Bϔ �y��Κ\�R1��iK��f\H,�;��'Uaz��	�Z�تtJQ�^-����y�f�F��@�y�pḱ	C��y"K�]�рMѱx�`��e-���y�BM�e��(=T�I6퀗�yb Q��:�a���V��a)v!��y�c�(a�@!�eN;B���O���y��Kg�h��Q�+�zEå�E�y�K�jxE:v�&#� ��3�ԍ�y�C�*O�����֋F����y���H�#��ΏU��qoQ��y�b_D�T����8..$�w�K��y�W�'�vYp���}�(�Rwh���y�b��S�d�u�&t��@��	Z��y��:jؖ��$�Ѻ	xݺ�)���y"�^(a~}�#Ě7a^P�JFC��yB��j�9��C�RInM�RE��yR�Wd�p��k�B��Ep��Ϙ�y�Ѵf�.����A!|1f�\��yrU4�}R���"N��L�@��y� �s�R�ˍ�fY���yb'J9���k� �4XE�[��y"��j�2- �)�>~قс7. ��y��B�t�ԃ@���w�>��՚�y���J�z�����h�F]c����y�$D!��=�#�1HZr�y��b?D��b��ŤX7Rىqi�1/�`�*6 #D�\KI^�,�8]E(0N�BV!>D�D��N���b�Q��LC��dB(D���@�<d
:����3b���j�c�<a���Qh��U�P;^Ul8�Tl�
B�	�U�A����$y>��ȩ)(�C��(�"4�d,]�y����T�4H�C�)� 6媣�ȅ��]�2oZx"�7"O��H�i��Z���M�\���"O�� A�$���J��ؔN�<љQ"O�D(1L�$R4�Ҁ]�"���"O�S��ƕ[&M�L�/�@��"O����ʲH��4K��/�D��"O���A+�?@`�c��A�S��r"Oh���Jʪ)��Ι:+9t$�v"O�Pp��5(q!�MޯyE�$�u�'�Ғ�����2U�����mNqc|$h��-D�$�k���q"���h�P�c-D�`�@�L*Y/& Iec�=8\����+D���a@
�g,�[�Ox���)D�p� $��Z|�[�C��]�Y�L2D�81�]�*�����iq4�.D����b�1+Hl�Ɗ�E༥�j+�Or�q����fj� @�BԢ��7>��%��R,H$P���8zb�J"*��g괄�:̬�5�ч�I:��Y�}�ȓa)@�{d�V)Y���*�{}����Tq���>)���g�!w��l��Qj�Թ7���-��I��*�
!Bh�ȓB�Mp��6N���N]�f���#�>|Rc�	W�Τ:e,�{o¥�ȓ]/Dy$aݩG(Fˤ�R�R�JćȓK��Q0D6g������|����+q<��"�̡v�&|��JQy�d��1�B�c����$UV/��`�2���Z�X�a�ϓwjHb�#ӊy9(M��D��Pp�/~���1y�&��'-D����H�rb��E�'7� ��b)ړ�0|
E�̋M��� ��΀+�2��`bGo�'�axR��@?�0j��7w֜� G�Ö�y"���+Ң`�A��)u|�������y҇�/��AO��y�D�)�y��1/��g�NG�,�u&K��y�ʊ�vQ�NÙ9�U��$��yҬ�!���"�I>@��X��@��yҊ<2�^QsMO�6��������0>a$/D�7䕢����N��$l�T�<�F�	Hd!`#ʜ�Y�|E2��Q�<i�Ȏ�$ $e�u�@�kA�=��C�N�<Y�(^�y@��i��r<��y���Py��' �1qwO3l�a�('8� � �'�8���#H�ŚH�Bh�Uk��D%�N��R/Cn��]�#�/J��L��"O�r�/�3L��aT��z�T�3�"Orػ5H�!0��x0B�U�x �5"O\ի���f�@����E��)q�"O Q�Aa����q"_��c"O�I
�I˄5,��uK�I�K��'O��!3��#Q�f�OV��@Y�+;��Y���� �!j��F�5�3 �v}�C�	�(���C�*B9E�e���=X��C�	<@j!�mWN]N��_>A �C�	�=<� ���2���^�L�rC�ɜF?:ȹ��U�P>q��.�0w�B�I����aVGu��m�4��7a����$0�ɏo�����W0D��Ё�g�
J��B�ɓA�9���RP��#M�
�pB�	|�`YK!D�_�N|�>7pB�I�>C���W6C_:L�e�ШH#�B��-	�tC ,��V�5��/TPC�I4��@���=RS+FM~˓�?q��?YO>I�y
� <�Ia�V�2i��x��E�'��(3-�b*�!��$��1�5�d�Oz��>Q �'�&��d�7�?U{"���OrB�ɢ=�5j���F���4�M<C��69���S�LQp���AaK�?8C�I'�(�P��BK����N	�36��d-?3%�|�ѡ������oJt���?���On������ �I�6���q��3�S�i�	oPl��!皢y����eo�m�O��=��P�!��2��	�Ճ��p�z*r��F�Or�`yv��>�8��!c�7Q��dx	�'�
=���s��)a,X�Yv�1X�'N�dI@ 'U:��� #B:Z`�9��OH�:�
����cfR�k�
!�t�'��[�)�'U~�u�C�=`^Ժ�>�V̑�' )qdN���VȠym����'8 Dyw�zd>�9���p���'�.(����!u���	b�I�'H��x���$pTܐ���2f����'��"�#�5;dx ��	�W ��n���$J����e
 &l����!�5�_�R{as��ܾ'�v��ȓ(�p��߀n38�
�X?�l���/�J���`��	*�;I���$����ɐ|��p��ˇ=��'���H��C�	+�xih����G�U�C�ɀ6�����q�T��JB 5�dC�I�h����c�%ZնxJ2�@���hOQ>�8 �\�[��x�d�J�wI�5�,�OP�	(�<��C(,e�7�Q*��B�p�lm	�'Sɶ`)��B�/p���0?i�N�<$p@����U����?-M.-��4���Ŋ�NR9B�4b�xń�	��m��-�/4~���Aq�.��F|
A����$?�t\)���U��m���+!I<�r�RįW%#�(G{B�'��>��#�W 0��@���V�b��k�<Q���N�𑹳a�㐸���i�<�2䊸N~�bU��TxV�13�\�<�v�U��Lx(�h��^h�p��V�<���Eô ��#[T� 7�V�<��(N=| `\��*qQLu�ALR����<IW\"���B�_\�@f��'Nў�OrDl��
P���G`�5sMs	�'N��M	�s0�xF&:�$ta��D,�'rPșv�	1 �.x�c�t���:�d�!A�&$q��ҴDS�p[f���^���8�kȤZ�|`؃�S�
@�E��A�d��T�����+Q	m�zԄ�	F�'��,Ti˛xf�(y��� ��'��B6�M�{�4�A����~�f X	�'���*̌�բ��d�|Z||��D�O�"|т�rCJi Pg� @
h��Ӭ�B�<�
�=�p���/ʮ�5�_c�<P*�5���Qg�����i*���Y�<���� yL}� � d����/�l�<aV��� ����W%�zn|x@F]h�<��!�"q�B�Z���Q*t�a�<��Q3%I�=���1��1"��D�'a���ܭq^���Hˡ��P��A��yfR�HQlD�M6d�!�D��y�����n�Y���.54D��L��y���9��l�v��5.�2��e���y�_$+���rc��[쐰C�Ȕ��y
� r!� dKm���Іi� ��ٰ�"O�����4"��E;�ιOR4 I`"OPu�� y	�I���)g�D�"O�H8S ۇ%� �C�%Ҙ<W`��"O4ij!��kJ���K�!i���T"OTe�!��:+$�Mz���n��r��k>1�2�F�{'܈��nW�/(v��7D��CG.�}�Li��O�PJ�Y��(D�$�+�+�@�r��L: �j�+ړ�0<q��Wowd[�
��<�y��L�O�<1,߿�P��@��.bN h�m�e�<����	e�U���A�f����Y^�<�K\�fð�% ���&��G_T�''?}�%�xw4y��P+8�� Z�	*D���� A*N�������nu��'D�)2g�-#����$n��tJ�J2�7�SܧM�����2a����2��a�\}��_t����ӛ(tސJ�cXQ̰���ޤru��<LQ�	��[u��Co�����X�<��Rl��s32�&�$G{�����M��aV(E��i��1��x2�3S�KØz�
K4HP�2�J��'�>�!���u9A1A�T�%+�1�)O(�=E�t�	?(�Jq��N�j��`�ݖ�y��j��s�Ƒ��ڳ���y�`�:Jk�tt������y�ȏDJ������?�^��cÕ���'ў�O��T� 
�R��GY�0/D8�����M:�����B�mM�4��\yG!��6��1�)���6DZ� &'5!��/bq��bȃ0w��ը$n�0_D!�d��@�j�����x�Q���y/!��Z?J��KC�h�:p�6E�$!��Ok��eʖj�$QJ�a��af!�D
qjJ(р��LS@0��Һc��'Ja|��O�U�9�'�F��n�n
+�!�D�O�X�pT	�%��ǭY�!򄝖���2Dk�\$(Cc\&}�!��	'���RC)Ս⹨�Gʴ�Py��ۅ~h�A���9RĀ�4/���yB`H:~8,��#=����d�Ȗ�yr�����C×aͺTa��_*�y�C�-$ܠ��o��%�&`��ybj��&�[FȔ;d.�X�H�+�y�$���T�?]xL��UmG��yRğ0Rf�%��E�br ��.@-�y�/��D���(b��*�����y'�;i�N%�C�@7��-d���hO����F7SBdt��gI�z�e�a Ց,!�:|�xcF�^�0Az��J�;m!�ƽ>�����#[REB�O�Df!�Y�'U|������AI���)A�$+!�A�s��@#�BO"|V� ]I!�䇔	H�Ӄ�\MbYk�f�$!�
 D* R��G">$��p���S�2�)�`~�17-*�UHa��"�����'!��j7��42����^F6�
�'mȥZ��
a��:�l�	����'�`�W��n�����*��~�C�'5�г�Eֻv�!zS��r����'c
0�$C�'���'��>�0|�
�'���`�7D����v"��5�d�	�'8�L�梟� ��"��'��e��',�0��"��~���0��#i%�y���� �ѱ�o�)aZ���G%q�v��q"O>3�"œb��-�΀��B��"O�� �Ƚv�$�r�]9L�v�Z "O�y�f�B�4��6�ֻl�>��"O���ƅ�u4�D�ƋwI80����?����CO�9�C�5�b�B5*ȿX�|��ȓ}��ԫ�� �4�x��AO�Z���ȓ3p~Lz�j�->�4�+W�S5J����8��]��c1N���!#�٭!nV)�ȓa�a��%8���2���fp�d��'� ��3b�t��q�U #jh��.�n�S�cH�m���KQ� $��&2�}��ՃDN� ���@ ����|"�1�%{ܽ�'텔h�2,�ȓY'���U�4���Al�R�\)�ȓ �lX�th�)i�È.�­��n��4RK�5�FH3t>�:�ȓ>� �d�
�����QF�lh�ȓa�Α��+B���FC�����'��=+��Z�s�l�H�	Z�}dŢ
�'݂MH6��3-���G�%r�,�h	�'��|����Nnx�r0����	�'�L�wnW3r6�B���T��'A�LCv�;�.݃�c�	O,��'�qp�l �~�ā�& �Q��5�
�'�4�s��N/)L��D�#A��a)
�'p ��*3j͸�%"3t�p	�'�Z�9���4rA�H��mG92)��'Y8 6�I#/_j��s�)��Hcj��x��i�����g*q`\h�˟�yR+%�h�'!�U��ia�M���yBI�T� m*�B����;S�ۡ�y���Tb0)�qOז�¹벌L��y2�W'$�l�j�Oؑ�PU��b��y����OM���G�=	(Z�ࣀ��y"O�S���i�!��^����U���!�O�x@S��I�p��3@�x�0e�"O���p���U�	9�-]�8�Je"Ofx	Pl�rZ��a, ����"O�|Ѣ��'��驅@�̊��"Od��e�J�T����Qo�>q����"O��x@�U�*�����.�&b���"O9���Шc^P�9D8����"O&m0D�G�"��
 ���IQp"Oܰ83nVNЅ�Y.[�n��2"O"삠l����L� Jг�"Orda�+[�'�{���"�x�"O)Q����'���#7��""O�����9R%�0R�~|��"O�(�9{<z��&C"�$�"OԘ{WF_�gy(�P���i��!R"O��R�@�#�Ҁ��d=�d�x4"O�ݑ�l+-����P�m=�ʠ"O:a`  D�0|r� ӏh*@�Г"Or4
�BI� O��['��=wdi�"O�9�����U,�y* �Y�Vt��k#"O����N�� B���sJ��"O�1A��J�o~�ƄR
6�̌��"O��{1+� lQj��s�D�\��ܻ�"O��0 �!B�x�XE�  ���°"O��0�lK�z6��8�G�<xR�: "O���-H�|k��dg�n��i�"Ox	0���?M� �����m��13%"O�9r�G�X�B-z匂�'���"O� !�C�3t��1�O�H�]:�"O0ɛb�U2�j��W�,I<8��"O���ލe�~�:ulv%�d�"OFݘd+�4(i��$�	�Z ��C�"O��p H��n�+��v�	�ǋ9�y���<�<���nޜtW�9�/;�y"FWtYn(�A�:6ذ�Q%Y7�y��T�H����n��4ȮA�э��yçL[r����
y�nU	Do�<�y�iI�aD�i��
�o�49� �J��y�E(kPy�!�7�2%s�c�3�y���6@DuU��j��c���y��L9}�}�ԆG�W<ܫ����yBg��H\���9JF�����yb�Sw�h�Fb�<��`�g��y� G�?9�֎H�5sh���P�y�[?" ��XY�zT���<�y"�
�9Ă����U?O�M��!��y�c)�U�] ��� ���C{^d��+P�bB���u��	�6)��g}��ȓ���"�/a��adm�V30%��3�>�����>1�<���1�q�ȓVd�����[=�,��wo�0�ȓ��]��0J^diks�u����ȓb��4�����%�D�I��ߢɮl�ȓgH����J ��#�j�a� ���3t2�,D!"V$8k ��}t"���<��,SD����0� D4�ȓ=�l�O��2�&��ƒ7i���ȓ8:���q�F @y!�w-�+d���	4��pA���p��H	&B&|���ȓBry�k�y\��(E��
p���u��ٙwg��'"d0���+��h�ȓC#VYj��
�~Q��rCM��K� @�ȓ!=��˴��G��Ы��?1�ņ�ʆ���J���.�%��4��4�ȓ����,�c���!������ ���fJ��4�U(.��\��M}b���+Kp����$%d1���iqe�ǆrT�Y��[�ӆ���*>��޴]�q�	�e�( ��z�B<���	sv�	�0a�g=!��j�>��C�(7rą#ю�:3Q�ȓY�Ȅɰ���uh��Cu�*TSz���M����&�3��#!))����r3��v��u�` �BU&/D�y��A��y:�GH82~,�
�) �e��44��ѧg"Q��իK�!�ȓ\c�A��MZ�>��1ra��Q��l�ȓB���ac$]�	���IFN��=V$�ȓ+Z����H��t���\����8�d�2��Y��ma�Br�0s"O�T�3*S�5�ã^QLĤH"O�9w̕�\ȅSB	� m( *O(ݢ�d�(A����Մ17�,+�'c���$�E7�R`[�!�'�&A��'�8q�oɆh���ТZ%U����'H��Q��"Ӳ�#H�($ �9 �'�آ�аN��x"O^��n��
�'P��)Z�BiI��C����b	�'BTT҃��<`&!B�EC`$p�'K�1��Y��b�P�-w��|��'B�}(�,	�9�Yh!��?���'h����T�N�vPrņ�5y
��� �u�0D� M�� BQ�[�8[l��""Oh���ȓ�,( ���3|Hb�"O���3� �	�3�' "pek�"O����Oէ/ x�G'A2&�("O�m�E�X���D&H����T"O!�E��Q�xu[��)�I�5"O�p� A�8B��`&ܜC�){�"O�`" ��
堡e��S��"�"O�3�ڎb'�i�$�[���(@"O�U97oĜ,�U��˓&B5c"Ob�05�;�ΰ�񃓽d�&]�5"O
�9�E�Ma�%#!$U��p�d"O�4+!(��f�{�#K��2V"O�=R�oD���飔I�P�d=�!"O�%@��'4RɊ2"��	���s"O]ҡf��~���$D���T�!c"O�����E���7M
?�}�"Ovu�T���s3L0~���x�"OP��VRv� �jA�k��Qy0"Ol�D�K1WJ*�H��+4�6-��"O��Kת"S�"FJ��v�ΠA�"O^)��B���~mp�� ɘm�a"O�l����s�m�V��,-Y"O��{�O�/H�s�P�~ق`�"O�3CJ�Yx��5 [:7�Ω��"Ob��0�
�}�vx��(ѕ��ݢ�"O�ղ�e� &�h��!���?�8��q"O���t,�6VKV�S�왊��}Q%"O���D �h{�j���j��P8�"Otty��BE�Dk�J&��b�"O�����b@�����?�H0�"OX�vO�.2*u���״pIz��"O�d C�_ bpV��L&eQ� ��"OD�k��5����.R*�"O��+��T�s�f���)êDG���"OXȳCᒤ#��Ӷ������*�"O0-����0pp��*W��"b⸁�"O4xI�ǘB�U�,F��zs"Oހx�ܪ�(�'�C�o.���"O�H�2�#1�$1���*iR�G�<	'
N-i��@��	'
 �q�n�<� O��#��@�*VrgD`ic��g�<I# X�d��@����K3@����Y�<pCL$:�M���N0�9+��W�<Q@�Ƙ>Y*@�+Ȃd,d C�DQ�<a�W�<�0���$��C��zDA�I�<�t��2=���녷wR���lOD�<���'�2�b@�F-p5��bsf�}�<��N�|�2񋲋�?���"��Fv�<I�+��@5`�:u W	}B���J�<��A�"UИ�0�8pVM
��D�<9�ѫB0��b,�28j �+��~�<��
��h���.hL�SQ�`�<���
�/C���sJԨ(�j��B�<)0kN�HO (A��%����AS�<��ٺc��ᢑ+�#S���(��HO�<�B��]�E��$&c��a�hf�<q#��}�,f�7�~M@f��W�<�LQ�D6=*�m
�@\X�vny�<�:h2�T������9��<i�!��I�i�8����ߐt�p�3ԣ�x�!��L9h��3\�\�r�Y��n�!�S�d��u/۝j�r���Q�i�!�$a�a��,tX0`�~�!�� ��Q J<��2��	�l�B"O��v���mG~m���0M��!Ya"O҄���	�,�)�F�=�~���"O���*�"b��<8�۝h8��"OEAͲ���+Q��4Y�Ey""O�@�Q�GXh��c�.1x�1�"OԠӤk�x�-ђo�	@b 9"Ox�B�^�L�:D#��T�/ű"O.�����(Ya��M��q��"O�yJ�+Θ~ >�rӎR�{�hg"O�ࣷ��+0����˓�s�a�'{��C$�ǺP����M8zߐ��'��TX��ًDQ֔�s
��&V����'a�ebѦ]�d�ִys��"��i�'\�iy�O3�B�	ѓj�H��'���hE��*E���3Č�a�"��
�'����S�ɣ1%2�:'�Wzΐ�
�'�(�fi 3h$C��I����'�Bu�Эژ� ��d�LSBn%��',h���O+
�$�z��,u�q�	�'���Qg �'%����F+m��L��'�J��)��F��a���s�`A�'�p<p��H̒��#Z$��]��'���SQ�Y�DV��r�m5��'�  )��եC�.y`����&�ݺ�'80�# �@��dG���=��'��YPb  ��|у��	�yC�'~������(F*�'��-�X�r�'�L�ӔɄ���1#�Ś(�X-k
�'z� �dŹ}|���1��4��'�zmA��3[���(��$��I�
�'��]��ŝ*]b��d-���I�	�'Pi�+�w5��pdc
5�t��'�L�����j��qz�69��!��'b�!�Qȟ�1u�C�+×)L�� �'φ,���"��y�(y!(h��'�D��fdj��U�s4�̣�'��x�MM$���pUȔ�:��!
�'��䂢iN�q�hq�Sl��㮤��'��c�i�7���#A����'!�[�U�8p����(�:dh��
�'��8��H6}n���� B�0/$�(
�'��=�f��L@@���=-�V�q
�'Xb�p`AG0r�(j��U/"�z�B�'a@�B��P�$�����/*�b
�'g�,�*Z�g����LH�#�j1��' �0��^>y7N��	����@�'`���/���9CW�Fq*	A�'if ҠO�=e��9��g�=<�&�;�'ޔl�@��?�pH�5��
9C��`�'a IA��L��@D+u�<���
�'�0���Q&u:w倲9��s
�'~f1"�Tk�ea�gȲAݬ�0�'��@�1�S(^�A!R&�3��Y3
�'� -B��!vQ&̐B�%"�X
�'�x�'�7<୻����Ot��
�'7`��$ ͗R�.����ŽF����	�'c��aM�66@����G�/8�!:	�'���H�&6=��:�Jȅ7���H�'�9�Q��4aN&�Q��_8*�����'�ĕ���#g>��$h["`�4�'�V���X�L�5���&ȥ8�'�p�B�DJ�ȹ�\<�݃`��{�<�F�W�w�A"�o�*� h���n�<� ��A�\�/#����ƀ#t�V(x6"O������-P�-Y0U�gT긠�"O�i�&�ϕ]�Dm"��M1^?Pٰ"OR�y�	�@f�� S+g*���"O �1ʊ,~ƾ�Xtأ3��!�"Oji҃�+2j���qbϐ1�H��"O��BbZ�����߮���"Of�2��E	�F@dǂa%"O��2eK�}ޱ���Q��V��"O6�:"l�&0���qG��n�dAB"ON�#�Ⱥl�~}s��#Ti|бr"O츑�@_�F IX�K=d�����"O�)c�!h<|]�w)\�L��a�f"O�}��L�<�<��GۍQ�
0a�"OhɲC��}h��H�ѯ%��S "O@r6靻zZ�I���I�x��"O����a�&��Z�)�����"O���BY�{
�4��.D#j��A��"OtA1��9:����G��Ez���7"Od�ir��"@Ȃ��Xit%d"O�1��ڿ.��<i��	%]@��"OT���Hm�2�RQ��
yR	J�"OtԻ�$���hq��.�6ɴ�6"O��q�fL�H�8Ej�o_�Ld!R%"OB��ѰR���Bn�T�At"O��D�(O+4b�MD^��	�"O���A�lW~y�3�
D��9��"O LC�`Ҡkt}kpl��\�z���"O�q0��ßH���*F̏��<c�"O
uk#�p�΍ZAl��o�DX3�"O����l��X2-BCk�o|p"O�"��H�3�xؖ�ߣOr�('"O:��a�] f���*�N���	�"O �#�0u���N�#�`��"O<��Š�
*r0R��M>L�\2"OVt��씅A�l=ZS`ʦ�޽Sw"O��ä�NNq�TQ��I�����"O`HO��U�S�6� ��"OD P��2��풤M�"��=X4��\��I9:�X}ƮۀnmD<�@�P�{�nC�!< �X�4K^�����Ȑ�1�6C�R�� ��$bk�E��2P���D7�0�&�$V���N�(tΨ��2D���Xa����ѮG�CnD���H-D�ds�J�A2X�K0e����/.D��c Ǆpgxu���d�
ٚGH�O�B�I�{��(!a[q頩2B	'i��C�1:1��&K�)Ȧ���m�/J6tC�6J�I�kA7>@|�Bu��(K 0���>�-[&N��р�,�F��CvfDF�<qVł6���*��L	Z�xg(�f�<I�o��m�A�3*�l��Rl�d��hO1���x��@ B܃��=� 8�i+#=E��4I����5t��ز! 	f��'����)�|BD��d?Ry�6)F���d*�<Q�)�O�����
JP�x"c�=�:a�N�M�ax��I4)�T��BN*G\�n�$5�NB�	��m���{ax8S�U�[p>"?�4L�Q>��jЋ:��A�ą�:M��Qg� T�`s ����@�qCa˦37��""Od˄#�%�� B*�@D�Q��"O$aM��eԚ�q4*O�=6t�s��D&lOJ�35,�*�.�Bj�G�|i���������S�
�;!FP�/�X��2-Y&oL���D~�� v��e��'��\)Kݴq&60He"O���c��0PJ���w���-��5���	g�OY�ܠreL�6Y�:�տo�24��'��|І��"g>ZL�#i�!l�T�	�'-<h$N¸��U
��\�Mo`�	�'A؜3��L�4U#!��OF� �Ǔ�HOvQ�kb���2�`[,��DR��'��	�2��|Ze��UfD�j!��6��C�	�Wr�y��h51ҸQ�.�B��#>A���$d����Ƃ2.~�$��.�I��C�I �h��#eQb��$���k_��IJ��h�9�.�?�ɓw�F@DƁ�""Otp��c�CِE�d�;4;��1#�>�	�0�h����aKD,LSm��ȓu,0����K�qy�D˔*��q΄��ȓ.�� {&Eϸ��e�DF]{k� �ȓi��Dۂ银Ft�[�lυ-�v���'3���"+S3��� ����+��<X�' ��r���;fKXU�&'H&&�Vai�'9&A�vL�:Z�.x6�S4 H!��'�ў"~��2�2]����?�$Hٗ`�j�<�1`ϋziD�0#蛰j��!a�+�]�<y�f�(����/��A��	V�'�Q?	�t�K�58���Q!6��#Wn&D��Ҡ�C�E���;��>�H���i�O7�<�S�O��U��Ty�Ić��*�R#c"O������N ����	�]6��7\�����8t�}�sd�
�	��'Ľ: ��$d�d�3Y@�*���䎊^��d�>D��H�kڽ{�`Ԁ�],��qa.<�D��d/>�N3"˼V�� E�A8�!�<OM����D׺d�jq����9��xR�K�'�"d9���9��Ic&㇫y����'	Z�a7�֝2%���Es��z�'L�'��)�!�-ؠ���1����<�����W�DS�dq��� �L�x���?���CA����K-	��\�BD��a��KF�7����$Uv�ڡ*�7�K�.M�>ݺǪ>�S��y⮝�4�����.cY�tB$�
��y“.���H֢]{�8 T���x��'/�S��)5�{��A���*�'�(@���^lDb�d��~of�a�'��qz����K��i�T ͖E��e!��)��<9��H��H�OW�3���١�	a�'�ўʧP̱sS���&�ؙ ����4͓��'�ay�Ē�^e� (���61��U!ӎ��yR��-fi~�Z� O%ㄘ��K�y�F:;��l(�KT�8�Hr��F����hO���d�E�Po��P" h�m��r"O,����N��e*", ϞI"O~�c���6U�&��ɅR���[��Io�OH@�{�ėEW��p�ɑ�D�<�Q��d:Or9Bo��rT��A-�^��`k�"O�Hr �2��8cpΘz��8 �"O��H�.�A�������y2`�UP�p�vOǋF7�`�����y�`F;�v�`��"�RH��yR��24��9DM��Bw�$c��T��yrg�#BZ�(��ӭ�@�@A�8�yBd�<G�p$&��
�J�;Ӯ���y'Z%V��2���|���,¡�yB�	����VM4&�����^��hO����W��P9�c@�2rES!DG�	�!�āi�h���	�*jZ���N�{�!�� >� c!Z-A[,��#f�8۔ȺR"O� P2f�&��A�E�"����q"O��K����3C��PZ7%�\5SОx��)�Qj��S �F�*ĺ��%RN�C�	�|�c�IH�a�$@�����x�B�I
N���i����'��%	�`�.lY�B�	\��m�7e�p��J�k_�l1`B�++�+��B{���� +_6B�I�w
�2�G ά�"��8.���s"O��m�t�@����R�O��Ec�'	���k����7X(]��FQ8�H�C	5}24O���D˝�Z���Q		�d�ZrK��N��	"FS�I1�H��7�`��)peC7�P�b�O^�\S"On���B�}�%�1�G�5��m���'D�ꓑM� ����'�t4�gI:|pN�)�!]�>}��T��f�6�FԣcH�0v�Dp�@G��'!��Iz�`C�Nӝw�:��"hj��rq�6O0�Iu?��'&Lu#��ݠ-��@�U��iM2�Xw�P*r�!�L3x��S��e-J�9�BƸ6��|���?�J��S/U�c>�$Y�3�����:+��A�c�Om!�D���N��n�,3Jy�@�ء	X���,E{��D���
��Α����{ŧ���y�:$�x`�r���4�D�	�򄬟����-G:��#Q�]�,czy�Ơ͸w�>��d�����q��i�mȶ#b����1D�䲤"ԅ&_A��i\�
��%`��/D� h�O��3)�0id@���U�V%-D�A%��/	j� ��	�7�E��.D�XN�.��Y��H*lٺ�A D�@cӣ"CQJ�{�`\<#����Q�<��s� fBR���9�s(��?OR���Ig~b �%FM�)p��٢_�.�!i�4�y�HS�u��P�%)�>Q����fn�1�yBJ��D)2@��I�f50Ƭ�y��B=z)["LӲCr@�B�T��y��
�j��@#3U�p�@� ��y���)�qul�;{��3��X�y�㖢��-`RbɌ�H[6�K��y�,و Z�y�U�ժ.N�Ҵd��yR��?QnxI$D�)�p(�M�=�yb�R����#�hO���ge�,�y�-�?���brEˋ0,�G�Y�ȓn��h�
5	��qPgߍ[J���ȓd�X�[ Q1]~�PCB�<y���
b��T �'X)s�
�!e��e�<YT� �VL��Ȩ,I�E��v�<�bM�%w� ��!��.��YF@�p�<��(>,x ��Ҝ1k�k�<YѰԑa�At�B[$VX�LC�I#e��Qk���8f�*��3@�/�B�Iu�!0�
�s�l�Ā
=�B�ɤ	��xsSdM7C����7K�B�	8hľY�U�ߨ������΁W�B�	��d���{J�`X�lX;��C�	"AF�����$⨤��M̹<�B��TYd	�)ޮ<��L�F�I���C�!C�8���h �)\���� B�IcԽI�ă��N�S����k2
B�	(:�)1UeأZ�jM��=2��C�	�~8q�E�"@	0��eB�L̶C䉗t���J@�F0 �����b�C䉐M�,��E�d'��I��͔v�C�ɏ�J�����8��,��lׯ��C�I�K
f��7M~�f�0�I6W]PC�)� �� �V�,���JS-A_�M� "O<����l�0A!����(�H���"Or\`�E�.��j��	�"�*F�#�Ԣ�␛T�^�	�A��Q�6�ɑ;���'$_	b��`���+2YC�Iq&��$1z1�% QK2�B�ɦ6F��@v��q��\��K/�dB��%�h|��̛{��!��]��C�I�4��M���ȣi8�),Цs �C��BbL�@�M"Ǯ�p���<l�C䉢%���q,HG��9�bT%K�PC�I/0��Pz��Z��N�i�N'8�C�	�}�$Q&�t��f�ѕv��B�>Uq��i��i�^���j�;.~�C�	�l�t�gk]2l�\D S�]�4a�B�ɴn�L�HgA��<`��D =:rB�IR'�m�lB�	�(�.Ao�|B��+*ɨ]�� Z��������5�C�	.)�у�.%��y�gi� Iq�B�	�j�R4��f��t�d!7��i)�B�Oe"�i��	?b���Q�צ,��C�	>�Z� ��B?#����3s��C��C�A�Ƒ��̂#MFj�@C��;z��	����OK�ݡ��ĸ��C�.c�y�HU�Ybb�[�kC�Z�C�()XX(@B�%�z�s��́l��C��5��a��}�"]c��ͻX��B����9`#H|�y�J�;FB��0g�z���#J-B�lk�cȵ8B�ɏ/�p�&k:̠�IՈF�#(B�ɐn���k�M�x��'9�B�	!^�c�/_�a2������ �B�g��11�KJ8|��L۱�ܧd^�B�ɛP"����I6=g���E(�x��B�	�Y�x���F��h�Q��k�C�	�f]���%!�� SbG7B�9Nx�i1E�B�s	΄�	Q(2�C��6: 4e0΄�S �$�!�N���C��F���J /Y�^=r��+B�" �洲���p�(�+���O( B�I�8(��f��12�H�dϑc��B�I'`�*4+uj�|��H�7L؟H�B� 	�FeH���AR�8ХH!@~B�ɋZ).��ō31Y�}�B��`�>B䉪cBQ&��!�`I[!n�u�C䉩r�����%A#Fy�7G�m0B�	8y�v,��L�8����;
�C��.	<(��@b�	�R����L9��C�I�̡B�F� qV�Q *�3Jc�B�I2LOZ<(D+]�Y�A�4n��L>�B�ɘ	�\՛7⁶p�M��ʺZ��C�	&~O��"#�-g)�	����IR�C��W.�*�ʰ*،�SFMD^4�C�	�8��!��f���~�P�D�?����D�;sɓ�%;��4�F$�zT-������x�F��7~=����n��8�����OV�J!C��
�b?5C�n\.-`�����	����&/D�T�d��! wx9�"�zW��� �n� �@ *���g�>E� JcB0X�pD4�d�����(�yB�܇1Jh"N�&�8����/��DD�YE�Y����p<a�G,�Z�x�䙓�.%y�AW��4�P��M1v��K]��6E��DJ45���H��D[�QL��ui�X���Ss'J�Z>�`�F���:Q� �IK$3�B,�R`�?;־0D�1%!�d^�^J�}I�D�>��S����0)�D�@h�c��9��)�g�? ��C�a�`2P��DW�+���9q"OB}ғ@ֻ��a��:~��xʔ�����p�X	Ѵ�'�p���K��|:�E�
��DB�tu(9p�+L&9��ء�GC$98lq�j��{(Ļ�-��*w'F!>�ҁz �4�n��H*�ruj ʃ��(��O�8��SmIl�ՑpD6N�]8�'6V��`��'zVI���ڡ���ҮO<٣��渧H�>�8�i_&!�٘5"ي\��
"O�!�4����[�,�y�%Y Y�!�d�:	���c.M5i<��q���!���1���w�U.�dQ��ȓ'VJ!�B��a�䕡h�*��R��;�qOR`�S�U��0<���dG����%'O��#��h<�	X�[���q3B8&*R�qe�(Z�A��j^���?ɕ�X�\��-r�Thv@-�/�g�'�&pڵ��]��1(+iw�O�~���ش m(Q�b� )�(�i	�'�@�wd�#H�j �bD��2:��OD�sB,)��m2*L0Y��s�?�I���pAb%c��(�S�K�v�<B�	?:��m)peݤk2���p�U�28䳣�Y Q�Q�F�J��@�K#C�Q� ��$��It��iɡO�L����<|O�ʄ�U���5�� �k li[�eى9�rիЍ){J�ئ"ַİ?�t�ƐU�vd�T��qت���LQM��Ӓ�1i"�*Ũ)G;����9Q#@ 
�2[Āܗon���"OV�X�+�H�B�1PĆD���C�� �|�D��TD$I�0F�>�I2e��q�Uc ɺ�0>rH��"OH��-�|U��zQ���R`z���4kވ���%ٯb`����ŧd������yAh�9+n�5@�,O�T��{���eB�	��9s�dK�6�L0�6�X�v��M����2%K����Q�,u�0{@J@��lH�JU�O��O\��	�"_��i����)�@Iɰ�5R�&óa��5K��V�.qp]"�ȓ��!��+`X�š���lW�Q�OY�,�ָ
��
:F��&e�%�h��.�H[ػ���6OE�)��]�'!��25�
���
�G&��q5A�f�=c�@�<'��I4��W �Zv�O��FzBR�"�Ő0l��D������=i�����AR���l� ��	J��-��jih�g�$�Pt��'�����	�-�t���&T��t4��"V�c����ѭ�Y&��S)L�,b��O���V�#]3���M�q�h��'��	���Q��d�h���0 (���x�� �F�I��j�J���|��wQ���!�ڃ͂�ˀ(����'" }�@�C�<����Z"^����Q�^ N Q�N�9�u1�%���U�$�B��:��P5��`�a��=�����@[2@����H�<az�H�-چ��@�M�|�����V�V�a}BE�<Q��⑆J�9��H*���'�D��2mJ�z� E1�cM�U|8i�J~�N�l�\�1�Ɔl+�A:��ڢ�y�`X?d�.L!E��szzPA��^�Q��k�M�S�����F�%��s�AIo�p,FY��ɘ�$�:� &�!D�D;U̎T���@��@�MJ*�`�дR��xI���%�|��D��$<�3ړ[�*�R��؋7�ԕ2'�R7y�����&z~���/��`���ֈ��Q2�G�Ig�PЂOp�Ѡ���A��pR�;"��`�I��y�ʦ'�1�&�YC!��*r�e	��TΑ�7"OT0�q�Q��䈣��z+��ID�O4��Ħ�[x�KI��}Z�*\�u3�<�u�������	R�<������X(��'�8x�p�+�OVO���r�JѺ�H߭�0<�1$HG��pI^;Bi�&*o������F�%o6��� �!xֺ�
T/�J��<ʇi��:!��1GH�h��
N����8�Q�c�@
e��P���]���b)�z'�a�a= {!��!� ٙS�X�\ܥ[�+��.����{���n�B~�-�9��~�ug��x*j1�B��^�Zfai�<��i±+��<#�AQ�<�~�Z�&Ue?����	��m�k�~B�Q����H�@k|��A��d��,*����!�,Y��+�-L%#�\m�$i�1$����m`.��'Kw�-�,�Q���v�Q%D�B�x�dP�,d%��=�O�R��H:|�d)� ��)f�[R� ��%(W����wZ�`U�m(��?�D��ƯH*�d�0@.�0��Ez��͞K'v`�'��Y7X8�~�d@K+0	>T���̀A�-9p'�Q�<��kV-&���@�U�&!h�P���6(�b�Br랪�L�(bB�\mG���{W��q���c	��<�vL��}9����d�=1��BL�F���#ω+��i ڑwQ:<�$��OF{"�V(��j�9w��-
�����=y7�"r]P �����-)�����pi&��z��<`0�,9g���1�'>�d�!��/�<�c��/'����}��("��p�F=_�(���ؿj���BB�"~�Q,@�E�D �$�� �\�!+Q~h<�GK�=\��'A� =�.�CGV�y����u'��x�8���#?phՑ�4y��1��|�n����C�KN��������i.D���`$_ H���@�P�b��h2�JF���O8
�9Aƫ��&��� �_"M�����Q���S&��ȷ�� Q����&��$��Gz�ڄ�#4BT��&B�d�Y�`G�m��d;l��kдq�F���O�^ ��ɋHl�qQ$ϓS�x
S�ҝrD>㞌��O�%�Jd*c쉈$v��
� ��Ms��	Og�}k!j�|b6f�
H�1v�6��x��T 2��C*د'kִ�e˷#�V5Bs��=���"FL9M_�d+���"7�٩j�|ʢhށYt� �8T`�X�Ȇ+v�:�K��<D�4��5sv��� ��(��=0e[���_"<PRH�0[��5�S@7v|�����BC�I�w����	�$n�2���l��.-f���[ :n #C�
Z�.�)򭗽:F0���lI�Qq
�@r̜98�t��#dS
Lΐ�%' �0=�&`�I���b%i�8�� w�Kw�+ �Iӂ��(�#�K%G�X�J?�rSŏ�@CDy�EM[$��Ѳe6D�T�A˚�	>��HҸ.��td(ȅ�u�G�1�d 4���O*�a������h*n�5��"O| �pj�(�v�����ow��f�G@?Q�#�n�Xm��$G0���ɒ(�2����Kߘ�C"B�;Fz����AH���ONl��p�@��U�l@��B�2��l��'���P�ۅ7���a��=ר�����o�ܢ����L�kM�Q�d�(St���Oϭ�y�� 1�d�:�k��I.��J����yr�խa�v�����>G}�dY�(��y�O�%.��]�4~z	 '�'�yR"��v�ҁC�Ñg)�h(@Ł��yr"A�M��������]&�8rg�4�yr`�
8���I�8!TC�b���y�\��}�VF�'0~��$5�y2���t,X�!Y�.&��� D��yB�/:�8 r�NRB8��pd;�y�\V t5[����<z�@�y�7<��@�5���d�x/D�����ǚ9��b�"UZ@ ��5D��s��& =�}�`��4!�ir�2D���S��s2����OV�'�<��PE0D�|����%���Do�v�H�7 D�h���Y�t*���D�T9ZL��"��3D���ꘃf
Lg�ZSi˷�;D�H��d�<D8�􀒥�t�̰�H9D����d+�@��C!P $�q�7D�8S'LS)C7��Y�g&�H�j��?D������7v�\��)Hc
��Ȅ;D�$1�B$�hxQ`�0Y�X�'9�C䉵u�L�P#��>a��S�D�4Q^B�I(m��)s�M�섈�
�Y�B�	�fɰ��3U���M6b�C�ɵ �mc%.��B:\Ȁ M�B��C�	��~`;B�ͻ|e�EA2+��L�C�	�E�>p�R�Y�I$���0"o�B�	�i�&�EiZ2,���� '�B䉶c��k0��*~.D��N��6�0B�	�*�-��@F(�8�u+W8�@C�	�P��DV�sn�a��ۖ-�rB�I�P�:$�&<�A:@?8�BB�)� �1@��#!�6a�ǈɜv�B��`"O~���y�������PZ(�(�"Od�&C�mo��S$nl�\�"Ob%rv�˵OU 'hR�[�,4yg"O�T`�A�3v\���R)c��@�"OD����?E�Vc�����t�@"O��	 �����H*%�W�C��qa�"O̽�q��4~L�	�眷m|� b"O8��F�Ly�I�+��?bz)$"O�����s�(�*�i��LP���"O��P����>�S�fƐ&x��PF"O�r�̥7$2���e#b� �@"Ox`cG���k]���DZ�EaFY@�"OzL����:k@<9S�E�Tl�"Oưz�#�0T��$b�CN�EK��J`"OTl	��
~=�wC[=3 v�c�"Oܪq&ʒ]Q�xi���#a 1"O�|��Q�~��X���:G)���"Op܈`OQ}ZB|s�`�;+����"O(�aB�Ӳ[���3w.�,�t��"ONГ���:{h���Q	e�@��`"O�<0��;�A��-�)X��"O����@_�h�L��I�`g )(�"O�!{�b�o�z���j@J�9�"O�|q��,����c��,�F�S5"O��˃�� �(�h���)�Z��$"O�������d��!̀lҡ��"O^9(�� X��0FT?UB���"O�E���<���s�S�p�i(2"O��;��ŉF�����O
���7"Ox=�$mݞ�*���P�;�z�xW"O��HW��tQuAႁ	�
�"ONyh��
<.%��Q�k��"Xa�"OnQH藩{�U�+Wm�r�X�"O�<pD'��]��}BI�)H���&"O����I�R�0��˗}NxI"S"O@����*͸WnH)|V�D*�"OX�䈐9Qy��Rt-g��)"O,͊3J�:��xږ-��Di<q�"O���o��A�f��T��FtA�"OmՄɠ!��=8�]�l�49�f"O�$���Ӳu�ĭ�2�R�|$��"O ��mN�$���%ظ}�"O��1�� +.��@��:~$Ո$"O���d��LD�U�*6��0"OVcW×?�Б��Cʙ?"�{'"O�e��'@@�+����(�:�yB��za�@Eѽ6�xD0d=�y�bD�?��ڣ!��6��,j`��yBo��{�4��D��r�z`d�,�y��y؁pb58���3w'� �y-�!�8��#L<��3��N��y�ܢ^�V�p	N�F'��&��y/�w�����M�RY�.ɠ�y��"֤�;����O��
`&�:�y�+��h���ꉲC���H��"�yb��$uE������(���m��?)��H�N�qώd1p�.� 9JB�$4�Ѓ�9*�@˦D�����-5�X㨌{1 ���Om�Tz �� J*�}3�-Xj�H��'r�`��a��2�B�ˌ#_eXyq�'2����*7��<�O?�����"7�U��/1B��*w�/D��	���C.�`ˡfW[��؁�J-?�փͬ-��сCe5O(�(�B-lz��hFd��\f(ك�'�����D�� *q�6d�P�V�Ge9p�&���DR�Px(�@�J-����:*�cë
��O�Z���c>��B����R	(�S��2�<S7��y2"�
Ʈ��0�Ͼ"N4]Y�C��yBLJ��{��SU���/K(d2�B�	SRX��l�'P��B�	���S�BVؐ��K�Xb�2��q�!���*����W��-Ȑ#�,FW��t�MT�a~��H+m�2�*�+̒F�6��%�#p
�hS���i��(��@��	����Pt���E}Db�$Y�`�ɗ29��ġQ�L'Z,�d�\F!�䑅3��h
�f�P R�]���GQ4=;��铿q`l0�Lׄ)����,��c�B䉝*���{��s��aq�ܤQͶB�	2j�<,C�E�Dh�հ��G�QvnB�	��$P7�H�+p�
����Z�C�I0a'(�T!�<!�L����8>n��Tڧ�6�axo�*.�.!�G�Gz��=g���x/«,�d�z��-����ǂ�E���2��fx����7T�L�u��+2ޝ���;�(O<���C$7V�T�#�3)0��T��ʙ �@��٬dڨ� g"Oh���+�$��BS�ht�p�y�PX�"�#:' ́p�Ǧ#~Γ~ �=���42�P0@����a:إ��8�������Qr�����ԩSj
_=fya嗿ml� �0���?�>Y�k�,H��8�
��&Ҷ#'Y���HBm3z��q�+�/}�6ِ�`��?l ��E��_�.���)R�Ka�(�`��L��)����A�`�
��'��P=s�����R(h�'>uk����x{��:6��+�u��ݯ�yb��$��z5I��}����M�p��e 2��/T����'iY�2�t���O�9B� �*���1�RG���*"O^(��m�FC~<�#'P�r���;Q��2I��1�dƐ=u��+H�0����Q�q�μ���\3V�BԡJ��y=�{���>���ڷѠs�l(h�a��34a!���U���(�aƃ����Z�)c��!Ƅ�T>Q͘>�O�[���4GU�l9�	N�t:$�:J4���+�,)q.�d�XQ���U�<�r�׺'�����@k꤈���*r�Sr_;�?	�&j�bա��9�65)��ڸ=�X�T���d�p"OR����&�^��E.	k��X	S�E8zY��Z�U�X���f�̔3R��ENl�'� h�`j
��Tpwm�*E���H�vӺ��+ˉw�h��偖_�JKT��{j��Bs�	5]H�%�U�G�<����!`YІAY1A ��Yp�,��O���|IԢ�M�3a�{ H����5j{>Y@�F�J��e�R�	s�!�$�<�&ذ���U�|,7`�+uh4�s��� !Q�n�t���R�Ow�ڿ"H��۰"�E}���V�ho!���4��T��V�]�i��#~��`�	H�v���qR0 ���O��HDz򈑎~�f� ��T�1�t��#Ԗ��=	���91VMɰȑ�P���㜏:��=�"㈗Y��B%�m7�٘�I?�O%XXkN\W2�����fV�O��i�,
!g��J8:�>xJ�˛���IH�a�D�a��/-`Re8'�SGX!�o� ��ǈ�D,�z�"JzqРFOnx�\pD�EE�5�T�7��;��(���V�'Q4����X�<�
-(��I`�E��@uVD�WOH~��Ԃ��Z��9$������g�'G�e�m� >'�="�jC�"Z]���6�	�	�P�! �	X���Ș.;�|vԐ !���.�(��f��Li�nX�5Q��b�"��Wq4�H6�	.#n��xЋN'Q�N�8t
¤*�!��P1'1���dۢAd8�ʕ�B�}���M�&�1BcI���)�'"}�q���^~��"DCL�n���=`�0����x*T1���U92l��OP�Zt'ƨtj��^E^ �ӷu9|��F�/q�=��Iu�h=)�L�9{�� n��vUv���JZ1{W䅓wO�`�O��</�9��$�5e3����I g�����ߒ,N1��\���j>��!qb�N�!��"OhTKA!�e�T�� ��i�R��Ў�$ ) $�"}�W�T,"a�)�WO��3��Z�O�!�� hx�2�Чc���F)� ߘ�ڰ�|RiTݜ����Z���4�� �gI	�fz����'$ҀxC�<�n�o���@�')��@�DH�&��X橗)t�<E��'F,���%��U�L�v��'�FUZ j�"[�p��D�i�\Y�'{N�2�!"j6h�ᓞm�X�(�'�,�y&��1+����C��gm^\i�'zr�{k�$H��mX���Q����'�� �P�m7T٩#bM�M#����'�Li�d-U"Mt�	c��410&��=C�
402$����S�I��&ƭ!'&�q^�1�ȓ.�m+%"�!�Xy�"ٗ!�-�>A֥	vβx����ED	���!�\9X� ""�*9Mn	�.V�a��%��'���P*M�pęa�[	J9fq2S��
����L��n��] t�U's:����y�hʡj�,�-	�.����!D�x���F�kd��xTŗ-J��:�ς�[�n,�FF��AZlź�O����M����&>7M�������9}���k!/�\{�zB�_65�B�ѣW�<�1��7 '����.~�HJ@�V}"Ԛr�]��&����<Q�A�\�%}(�`�D#L�@�]���k>��6퇳!�� �J�G=�RQ��"�$�*׭R(�B�O<��!1�(����fN�/{zq�����']���B�5>/ҝ;����ѝw\���� #/C쨛�f e�h�#�',`�b �L�G� � *��['~<�B+��P�.!��'
p��V��F�O

4�o�g\�����|�|a2�'��i�7ß.\��͓z4-�G�N
%�r��ek�+J��-�'H�� K&�0=	ԩӠ�)J�@�P��x-M�*��U���'Ψ�dʂJ�M0νK�@\ Su�DyD"O~@��,�?=<V=K.�u~Y�Ө��(����=a���Oƕ� Y�"`
�ps�W{PI�"O�ya��GR���A"Q�=���"O|���vx$4��ᘹg�(��"O��U��D PU;���;!�@AC�"OZ���X�|��%�3�ʇe�D�"O�B#-�%�\����=nE�4��"O@)��쎉=h�(�&��3��S�"OpP���J�0��`�%�%=0��Е"O`y˧O�?���Ō�֨ɢ"O�y:��M�A�����2,�y"O��K*wv4ؑIR>A�1"O4��c��5bP�$a�#C
8���"O\E���'n�H��OA�^�܉%"O>��拍	 &}*�����* @"OZP��Ċ�
^ݱC�	�y��Q�S"O(0[$L��nd�A��3Ӹ�X0"O���W��6���D�l�&�Q"O�9�a����y�E�Z�jC"O��pMF����C��/|��r0"Oj,��Ό�=��2�*֡u0�S"Ot}a�,���C�
�2S��m�"O�̳1#�Hɰ%��k��b"O4h����U
�|��Ķ<��D"OH����P�OڰYxwϴYm�@�f"O*�Z���p�h�R�R;f�ܤ��"O�):��O�I�Xer�� �=�f�	"Od���fɔ�t�1�ᄑz��m#�"Oc�®-�\J� K�>y,!sV"Ob���ė�@<�֊�@|�TC�"O�D��%E�A(��jI��	Q��h�"OD9J�5�Y���]?�,��"O�d ���(I�Y��ˏ6q~�j�"O�����N�j.�b�_=n���"O���!a�j<����,c>�d"O������@��R�۠A��H��"O� ���$-�+[���;e�M��`J�"O� ��柨@�a�j�i1����"O�`ֈ���pZ�^��I�d"O�] �B��˖��3�7.�	�"O��3wi_	H�j�)s�٥iX(]k�"Ob�B�Ղe�:a��� X�M�T"Oz���e�2j^�LWH��&ѷP�!�$�qH6��Fc�$98�42WE��!��"E��TpD-A<yS�*��!�ӵ�\�!k��d!jx��*�	;�!򤟋aN 8��j�Q- i��FF�[����,ȇ �D���Jģ*���P�+|�tɳe;��=BB��fxTTA�=D�����J7w�����>UV��=D�l������l��%L�B��s@<D�P�ъR�k�
�����cX�m8D��A�â���y�+�]�PX��7D��ZΌ"9��z�bDv�����*4D���C_1-:V��ՃޯwZ�TY"N2D�؃�+��5��Ж�ɱ(�� i@5D�؉u;l�1��Ҿ6'<���"3D�a0�Z >~���or�q��K$D�$���X�t��!�KK�r[�l+��/D�$�` �
x�v�zv懪B>���!h#D��P�.' =�2G�:nr��"�?D�8�!%�8>���k�G��2����:D��ٳ�Х1B���G�O�؄��K.D��S䝏l�l@�Mð|��x3��-D�z'��8�@sG�.����׭�ON��1���M���:?�O�����n<�uJ�*}��x�Ӂ=[�����T�1�6�ڷ͇>
ջ].�����0|Z��"x�kf!ϡd[�}Ð�� u	N%��	1f�J�E����	Z�������n�V]R!B$>4��2v�W�?�-i�U2!E �K# �c�z!����o>Y��M֢H��R֬��yX`agL�[�f)����ę���%��vǶ��	C�T��j�+�� O�l;Rj�`g2PB��/f����$�6#�xf�~����c�8eR5XE�st��cC �-;�CUUuX��!g��87��
�'Vp �#q�ņ)i�� Vk_qQ�����\h�����.MFD{'���P�%�?�x��tdD1��������2���o�1WN����Ц%�!�D@�&�V2U��9���f���!��or"ٲ�o�4W�M���H�&�!��ĵh�t81�	ȧ
@,x�$��V!��O�"�b%���N8l%�Yp�LN�-&!�ϭvt��3B=jY07��4Q~!��hb�����!O��pp��l�!��|}����Ŏ9���SB�.0!�dU�n�^%�7ᑃ��1B
�I !����Z�뤄Ł ��M��gG�m!��;s"��5l�!�q`$Ǟ�4!��*�jmZ֌��X�U�c��R�!�d�>&�2QF��&��zGhVF�!�DՆ�VZ�Z�B,��
��`r%�ȓw|t0��	��͊��!^i���ȓ]L�E�v�Z:_b��,�$!��^Y��h� ��,���K�ImRE�ȓ7�D��
��
��uK���Q%(8�ȓxb�E_�D�E�
A�豅�"�p�˂�^�YCj��bcQ$z H�ȓe��PCV$���҇G_+m�����g���#��!k�<��
��n>N��ȓ$�{��Q�TQ`��֬��t�vU��Z�:����0�"�ʅjG�/�Y��s5�L�3�ay���t���pz��ȓ�@)2�G�RD��)�!��Fʨ�ȓkȤ���#ܿ,7v-a���mT0��ȓ�<���*'���V�	-ɴ���S�? rڦ���Q1H��GGNp1�"O�i05���X��$��G��Z���"O��BG,X��9ڦ&
�/3VI�"O`�;`�(>�\<`e��,=+����"O����e'�3��f��U!�"O&E��W�%���IC	�Xu�Ż�"Of���UHp䈢#��HB 5"O茻��+*8��y��$
��V"O� !D ��0�j�cs�9t!faڦ"ODa�� �'��-bQM��Z�Hv"Oh���ʐ9Z| qgLy|���"O���VH��� ���Y�R�͈@"Od<br���Td��n�s�(�d"Oa	��ɲH��1b��9--�\b�"O����-��p/P���Y<`��"O&�kҏT�I���+�J�u�"Oj���L��E�8�vˀ� Q0ub�"O�r���#Y�Qp��3#6�H�"O
P7nb��Y��j�*���""O����#�d}6y�2��2��)�g"O�D
a�60;�T°��T�@} "O�0�A��#T�j��%�+���;�"O�Ż��[n�xa�dӫZP�D"O���X� ˄�2 !��V%~y!�"ON��u)��7MH�Hp��03��yp"O`�s�gH>�8TS�C\��5�"Ox%+���#*pN d"ŵx�H	 "O΄ ��i��E#"@ڧcf�"O��a��H�p������I2��"O�\b��R
����& �5�����"O�������������WYN��g"OJM���Ɛ{=��s�iM�g@x���"O��Y�	�
pFҵ���ʹ��hrT"O: ����z��8v/H� ��,��"O�-B���9Jt<x0L�	Q��K�"O�P�����b��$����	<<q)C"O�5"�ψՀ��S�ƌg6��W"O���Öz��a�v$U;��HA�"O�33 �x�P"3Q�hl�!"O���6 c����?Ј�z�^%�yr���0�`<�'�	�2��8RT�.�y"�ʛY�`�C�))N����)�yBe�(*�m��jB"1�9R�O�y�Z��U��L�*f��X�KK*�y�D�5~k�e�3�\� ���
L]�y+S�Q�2��c�
�"��J�L�'�y�aD,O�@ъ�lJ){�gɯ�yrB2^��]��ݨ9P68�5k_�y�cZ�K� ʒA�1�����P�y��&�fXˁ���<[Ih�
�/�y�잙��Aǈ��8�%PAC��yrf��s�tek�iޚg��	k�'��y�K�f9ʅ��'.-]�	���7�yb)�#6-Pp0���"�����y!Q`�0xq�.���h�K�$�y�b�����ab��'��8����y"�Y� 7H�:ׇH�zt2�re��y���7�����tn^x ���:�y�B
�T�j�#"�o��p�BɁ�y⇊8f�yz���:�Q���B�y�k�v#��x��+B6 ���K�yrL��*��D	 �&e�azt����y�J��>�*s`�+�������y)��'F,`cT�?y�h�r ��2�y
� �U�a��2&��4�K!�yR�"O0](�g�d�AX�����"O"
a���q��X@��	3Y�0s"Ot����Z$X�Ġ`0bH�J�yI�"O�)�P�۳'�f���t���"O��΁�\�f��u
�A�R�2F"OF,He��!Z�p)�H_5hؘH�"On`��%$$���RrjX�<���i"O>(c���.�� �镐g���s�"O�ir���~�������U3�"Oƥ���>F+I"o�A��H��"O�����ܨJ�MF�߻ �ThP"O�]���" d4�r�զ��E"O�1p�J�\��1�R���'�j���"O^ͺS��.��]� oT�]����"Ov���팗w4�c���	��t��"O�)���E�J���D��,��"OV�1C�6�<�p�̭"�0�0 "OLq�ċA�ܐ4���0��C "O�4I�N��H&�8q$�_(l:�"O �%� p�dhdN/�8��B"O��1k��_�`��AD��qb"O|�G��"@���S�+7�x%kb"O|���߻<�ƌ֙2��p�"O�Di[=��}�0F��fܨ,2�"O }	��׃p�2���]*=�|j6"O�%����[B�1!ՉE�bD��"O�A��JW`DD��?���"O�T�� �l9��+,D��A2"ORm��	ػAr����M9@�]��"O�p� d�8�4qƦG-.\U�"O^m	D�K�iW�0KFE^d����"O�xH�Β̱4&״vm�1P"OH��J��N��Ukae���8�F"O���Ē*�X�C� g;,���"O���K�["(��#6P貗"O�4��E��`�V�s6��+� �d"Ob���3s�����ƊD���u"O�d(C�F& <�#��1;@ܩ�"O�Ie㐽L��	���B�P7��"O��j� �-����d�`���"O4Da/	59�bb]�'����"O.����ߝ@�:�Z�k��]���e"O�X�K� ��ԃa�)[�a�"O�+7��
!c �y�g��n/����"O���
��E0�@r1��)S�\�"O���BH�_��#�l�&��"O-�%ٻ=u`� !|��H�"O�u�t���p^�$H�%����U"O��l��Z)N��K� &����A"O<���#� <�4k�iI?A`E�"Oⴁ�j����)�����@Q"O���d��4��`Rh�P�"���"O�1���h���!F���!F"O����m�A�
`ْ�0�*5)�"O��
�B݊\�EZ�$M-9�<�:�"O.�R�gVc�D��"��z�ڱ�"O�h� 6Ҍ�t"���$��"O����,B�@�~��@�P"O�X�3BWs$�$\(H�4�p�"OH��䃲⤡�r��Z���˦"O�=�
=D4e"��0[��]A�"O �KQҩu�V�e�q��!�"O�l��Ů��I�'�Lu��{6"O� �-��`V��Z��Qߎ|c�1�t"ON}
wM�i��B#[#D<$0�"O2=婅���c'��Oj���"O��)Â��Y�Rt���ـ"KHI{B"O(I�5��#x�	�c�
20�#"Oڬ��,Ba�Z�C�� f���"Oޅr@�B?����`C)) �i��"O:$4͓1Y��T�w��(
hl��"Oy��E&��X�����L��"O�dA���`;���6q�^��"O�}	s'�'68�Z1�%��mT"O���q$�' nb��%
�v��К"O�����B�S
�r��*d�F%�0"O�(�l�h7+
�=��$��gO�<�G��lr��G̙)��	d,Ge�<Ѱ��?`�Kg%]R۴�@!��]�<!��_�\���25k��9Y�IQ��_�<��`��F�0�`%TDY%˓X�<a��#X��\��&M08r�P���W�<5aٖxʜ�i��M�.�U`pI�V�<9��%I�}��؄ZJH�K�� H�<q��/p��v	�*���@B�h�<�c�ѣ)�ٺFQ%x��?H<C�I���{���`������^�.C�I�IϾ@��LK#�-��L
8^ C�ɚ �x�f�d,h��a����B�	�xx�RLۦu*]r�`���B��!V�bp��`�T�^�y�)�dB�I:��tB�]���B%�^�kSXB�	64���ĵg�x��A&%nC��}��;v�ª-�"�y�,�YExC�ɾ_�ltb�"��DE�����U�SQ"B�	:�j�*���7��
T�@�HRC�l�x��ݧej洡��S�A_C�I=P:��tca���wM�)t��C�ɑ����V�6�l�e@C��B�Ɇ���������ʧ�ոfuzB�I l2�%��_�,�{5,ո*3~B�Ƀ*�@7���=�4=��l]#K9�C�	(n(�&��$��Ө�n`�C�I:;� @  �P   b
  t    �   �(  �2  �8  	?  LE  �K  �Q  X  Z^  �d  �j  &q  nw  �}  9�   `� u�	����Zv)C�'ll\�0"Ez+�D��4��M;�(��<1�Y̟H��Y����4gï���b�愙2A��11��A�"�Sb��{mX���c�u���2��t��?U���C�}����B&PVD�S��(*��P�\��h�'�#4�Ibr�λV��݊Wh���ğ��5�^��@[���m&��P���Z�[/�?���F1���۶��j���Ӕ:o�'��'����ʘd�Z��ܼJ���$��'�Rh0w�mӾʓ�?aŮ�����?i$�^cᔽɇG�8m
.2��?!��?����?��C�%�?�p�G~��O���SQ��=J=��w�Ҧh2L`�"O g��3]B���!"�	8�U��S��Fxr�Oh����H����� 
��=�BZ�vz��MU::�';2�'���'��'3�Sμ��H�w?"A��=�"�A��@�ߴr0�v)|��	�'1�7�IҦ�Bߴ���'6�\�č<���ӤI�&	�=���I�-��>m�#T�&�����"4u�!��L�H���k�]��C'Wv�|lm�+�M[�i3��>�ƙid���X�"�5��9M��)R�܈cP���'S�a�ĨKUf�]ñ���JI
��5O˄M��Y�g���nZ,�M�B��6
ظ@mF�EI�Q���É�jU�2��t(F���ix�7�P�2��>&P�� �
,]N|��JH��la#  &Y��aa�e�a����q ��A���M�Ҳi�86mʱ0e@D�� r8p��eU�LL���e�M�4�3���%v��(bcR̦�aT��&<�pE{0�	#`|K��ݟ��?Î�"Y����eڎY�<<`afO�?)���'�R��,�r7m%��������-H�"�W����\�'�r�'�rD	4�\9��,b$�1m�O6��AĐ�e�X:}�F)�7�ù�0<!� �7�TmR7J&yq���4}w��{�5鰑��Ҵ}�؄(r��cԧ�?����N8'M��i�"ϵZҨ�c�
#q��'<b��S�D���bG��T�v-��,ܦR
>����H�A�	h�x!������,�6,�O���k�l)�'�y�*�Č8��ˬ}VM1��W��yB�V4C=,�X� �A��+���y"�YE��E��<_�Ț��y���FY��{�o�'��2@� �y"�µG_����Z�&�����Z=�y�oU�|
|Q �$��L��H��I��?1P��#<E����"R`�����)y�1i���1{�!���uΈ@�N�[L!2�T)!�!��G�L�uȌ�0�2����!�I*a����i�c�fl�a��*x�!��=<�(�ƚ&z��9`���o�!��ɶL6��3U�C!P�(7Ð�=J��=��|��	�&�^ir�K�����O�I��C��� ����(�����t��C�ɹ+Jс��C*a��0PL�%O_fC��lgȀ��b�Ysf��9n`C�Iv0�z���/c"���l�����dI�a.�m`~�^H�Ȍ�`�/t�f��s�ڙ�?	,O��d�Of�$R���	��Һ8�\�堋������*nXl��"��Jb��S�#O���!Ę�*��]k B�Av�6̀�>�T�	�ش(dɋ�gɢ:�I ��p`F�����UP�4�?ya��.���a�%dbI�Zbd�'�哑}���ʳ��{�Du�4	֨V6���\�t"	�M,�AEҴ	�j�����OV�OB���c�8_m1��|ޕ`ea���Z��I�&���q�<�������YW(��<��Y��s�<�@K�
��)���ݟ���Yv�l�<A�@�0��0�vKA���1fO�j�<9#g�8T�P�ye�[��hC/Fi�<��ȍ�0`��I�q�n\I#� ��M�H>��A������?�����dщe���T�i��i��9�Xo�:��3�iu��+�F_)����'p�Q�j��f�b�1c�[�R��5�Y��R-R� 3�����-�O�^!8�+Aq?�U�\�~����!*z����pC��MSt_��W��O�c>�D�O��D���LB(yN~0��J�Vu`��Di�6�X�z3��	:n����P].H�'��6-զ)%����?ɕ'��H� ��'�<�R'� 76�`�0���	��7��O����O����'9��9uHQ���EZ&愥7����ŧ\0�T�Yҫ=U��C�Y�����=x���p'.�:<Δ�2��@�X;�@�fM�A�0��
�+S��(!�e%�c[V�3DH
�<	*F�Y�5x�Xb��џ���4����O����O4���O$�	��٣�0b�V���ٺm^H����͢,�����

���j"C�	5�M����)Lv���OR���OD�	���Ȑ`����Ëc�B�'���
��'T�>������S��=d"��Q��� `��dI�G8�Ps�HW^����B�' ��a�k
�#��)��~r��׌���=�/�4��@�k�$#?!�Q�P�4%	��@��w�Y8XQ��1f�Ԉ�̒O��7LOp �1�cu� ���2�$%���'����P�2]NI��Y%	Q�8�ꁇ�S�lx����MkO~��O���'\������I��g	��Xl.]@&�'�o�@��Y��֗V�xa�;O>�u�F�'�~u��iO�}Ʋ0��+?q��_�{�R�`��U�DI�گ��q ��6�ԏQ`\y�Pc�6qrd]���䆮mcR�hӼ��O&����I����c oE#m���L7a~��O�d�O��$(�b�Ф�%K��	�"��58џ�q��)̊dК�R�H�C��H�dB�<	�ꓑ��� Y�m����I��8�'Ѯ���D$x�����S����Y�����g*.Ip�O{�i�n;����CGϷo	��{�MU��,l��, ,��^(,��c>-�u�>���"UH�Û7�v� ��ϟd��ş�q�m�ݟ��|�'�B�Y�fmLْ�M�qm����	�V�:">a�y��o�� 3��?7�~ة� R���\P}�[j��'�������鈶Sa����\�DP�HK��[�p��a��惡��؟��	]y2��D�)@p�ٲQ��*��		0��-���~�t���V۴E�@'�6 �ɦfͧM����S ѽ"̤"3�ǁ|<���iP3>q�>	��<D���h'� ��F�Y`�d�	˟L&�h��J��<a��ЧU�v][ŋ�7o��(���y�L�,�����	{�Q�ǂ����	gy⇘50��$}9�oܹ!��S0I�&����C�'�����	џ��E���T�#%��$���g�io��#ɽ>�X(Ԍ��(���	�1*
Y�"���U����7�^���Y���t�(���74����F�5?��>q��Rџ��Ia~�P�_q��s���`���A�!��Oj��d� =7L,��ɓ.*M��R�J,�2��OJ�Ӣ$͑|2H����-tRs@�'�	�r�N�A�O�K���'K~� ���G�Rt�+L� H���'��L�?r��
q�~L�E��h�ʦ#|��V%t#�uaV�]+!���0�h�q~��'a.���f�Q���H�=�]�}z�o�Bl�F�T�p�7��p~2���?����h�����G� ��`�	�O���3w̖`�0C�I �P��T+7J����Po�(0�?��퓌��İ����7�t����Mo@��']�	8c���֟p�I��4�'H�����T�$�H�g>�MD�P�
���F��O�M�u�R?P�1�1OX�EB�0v]+cƆ�W� ʰGI�D4�tAЇ{�>�	��Gs9(b>��P�>��� �h�,@�e_�l���
g����'�B]1��?����ڥ'� 9�@&u��lQ�Jܐf%�C�I�V���y�'t�|eI�P
>|�˓\c������9�t��G�C*dB�)r�<O�"2m�O��O8���<�|jm�)i	�#��-֨ڴ�.`8�+`Ƃ�u�@5 3D��z|�yb#�,A?��Ҁ�!=(]#��P�  
P.������S�]SǴixг���
�r� �H�"�&��s��!e2	hP�'�B�h�'@��I�%O ���`%X49k��R�'p�H
�.�%,a�����RHm:\XJ>W�H�?y#Iz���B#Vm�(8�I�U1���	VR�<��Ài���G��X+�=T�B�	�H;���'�/�`P�%�~B�ɰ��12����xȑ-P^NB�I�:ԌIѽ*��d�)K�W8<B�I�oaB)�ЁK�bѲ���>�Ң=��
�g�O�u����E�"�����s
�'<�D�q`��*Y����싺i�4x	�'����K[9U^�Bƭ�*j2�#	�'���"��%On�j%e_ 	٪<;�'^|� �e�[�b��$dI�Ѡ���'q}����<q7�0Tj�>q|���7�F0Dx��)�p�(lZf���Ur�Բ&��?�(C�	' �D�f��/I��gk�*�
�':�-�p��kv�e�ɣd?jEs�'��(Z��r�~@$.a��л
�'h6j���-t�:�cK]�G��
�'��T��*��h��� f�$C���2)O\0�'�,��BG'5`��gƮ7���3��� L�9bJ.��=� IXW��0�"O8�V���r�
4Q4o��Hʬ��"O\Q�mH<�Ak�'��.1"�"O* Y�D�=�D����P�Pm�Ha�'�n���'� ���޹��<���${�&��'�X�k�MUh�K�L�w��ͪ�'�����0�*�$�Z�v�B���'Hz�/�LTԁA$D6�ٳ�'4IÆʌ*54�$�3 ��D+P���''`h��E�!bY� �7-^����d�g�Q?=që�:A����K#pA�@���(D��J3��r��@K���#V�؜لh'D��P���c�|�B���C*�x0�1D�`9���s����"�2#Q��31e$D��! ����JWo�,t��K�� D��oZR��]��Vԕ����OX(�R�)�iv0��Ø�ef��1H�<p��l8�'*|��c�>������ �n�|�
�'f�!�g��e|�����kEv�Q
�'��8R�mʏ|XPj�0f�Q	�'!b`�¬�1/���Y^�X-)
�'��-J`��)o~P�0�Z'�\1c(OZA��'���Gn��ǂK�&�����'{��ʵ�C�h����e��%�Z1��'">�1�U(r�>t�@�d�R5��'NL�Q��w3d�����X�z��'����a)?ky�	i��;i�ma�D�8���56y+1]�H4�劗��/�~�ȓE���h
8c`ѢD9A74��l�F��f������0o�
qi�Շ�b+��V�U�A���� �!�����>=���FOXA$��bB�pn1��%&��cC䈸K�ڍ�᭎��P�F{2�V����X�I� 0~U��	3E���PC"O:��`΀�+�����#�0����"Ol��� �0��Mi��M>G� QU"O�t�2l?"_�0�jQ0`�Pب�"O���f��M��B��Ψ�2A��"O�-��S*�N̸7g��vm����'B�X���S�i+�DXr�E�x[� "[�-#,��ȓ,|��2$RJ(�9��_�5��$�ȓ^M�l"㥆�'/
8��#	_H��ȓhT�M���Ā#� e��EűWt䰆���]Y H8����F�-������������>?�Y�WP�	���'�{	�[L��Q�;�*uztlB$)4ZՄȓf �ٶiʮh{�����ģV�N��d�p�S.�9"���2-47t��ȓb(HP�'��:�����%M-lTT�ȓ�����)��X������,i�pd��	���	9 *�AЦ��tԺ���OI�d�*B�I�)���b��m�Xh�Q�>jB䉓f*�K �@0�Dp�%�3�B�	\�RL3@��w,0���c��C䉖H�6���oT�={@Q36�]�eƔB�I	Kg���n���k�F��:���=��-f�O�%:�����X�ac��*yp�'!�l�#�ƎP��I���.�p��'���7&r	��$���m�P$a�'Ǻ���:7��
%mȋ2�\���'�4)�ձ�h��쒴9�x�1�'��*�(��^�!.�	}�^4a�]t\Ex����Q�,"�-�0r|;2�R�C��9O�Ȥ�nѬ{�`���ێZ6B�)� >��1 ��L�ZU�$K�11}����"OT�;6��q���y|��9�"O*�j>I��JϿ6��v"O`l���O�H(�ۆم�����Y��Z�$�OJ��pƑ��q�p�%5�|�"O�E���L�	K�c�R# ��%"�"OP(@kX�+7�%��1b�L��!"OL��$�_�x,�<��-�~��"O�K ��-@���cD�E6 ���'���:�'��Ac"��nl\��,G�m��;�'~<e6�֥g�Bic�-T;L�'&�����C#����!�Z'K����ȓO2]��!�~9PD����>�� ��VXԹ����+vT�@��9BK4T�ȓ@ʼmBPO	2M�ջԡY�w �pD{2�O�����t#��	ֶ��胦f�\�I�"Oĸ{GAҚP�mj�	�JOv8�"O��O�J���f�i1��2d"O��h�/D(V��`1��ɵR�ܤ��"OHp��C^�4���uA�!]�b$ V"O�Y�d��?MF��9D@^/Pr�tB��'9V(���
���KAh��A�0���&���%(�R��z�VA #���<���ȓ\��9�凚%`FPP�dP�aZ���qFx]�qN�s�I�Q�0s,���[����-�1? ��!K�,��H����8еO��	z�T��eH�s��u�'i�R�tL�!�цF�`!�`ҥ e�ȓ@�6���% MonP��٬2�0��_��3�h��
+R��ֽG���ȓc^�(q%�Äl\�[ģ�Ec4��ȓ��`�E�	!ۊ��$_�2��Ʌ��*M?T�ɐqu�a�f��<��иg�E�C�$bZ�A !�*�<8�I�$�lC䉵
Yb@�Z�I܍�⫔3*�B�I]a���BW�2e�)���6Z�B�ɱw�f�D�!�ę�f@
���C�I�2Z�)�#(�%/Ӝ�"�h��idz�=�FSi�O��a� ��d�S�M��?���9�'�>�H A?2^\������a�x���'k^q���"����w��'��i�'B$1����%��N�TD�3�'�d���a�*�$Qc'`T�F��pI�'��A�@36���Y�Y�
��=K��K���Dx��	������F� ?�հ��?^�C��*g�@�j���O�u�ר݂_ٮC䉍9�l,K��xD���.]|�8C��kd��A�ԿNuz��r�\$tC��R圝���Շ*�l�-�=#�
C�	����J�o�zq)����ʓW@H��	8k+�̚�E^
K��T�b���;JB�	!�� �	�\�d�#f�Y�-�bC�IE�a�m��~1�d�Y;~�$C�IG}l�����P���R'ͧf�B�	':{��#Vj��*H���IV����Ȼ6����v,�=a��];b����e�i�<9E	;~���b��NeΌ��Nb�<��k�l�����*�x��KY]�<��n�=L��wA��b�W��O�<�3撨�v-s�W!D���0j�L�<a�I$%���K3�V�@�Ry`f��S�'������I�~��Y�l�1	x��R!݂A!�$� H�P@�bƯNzx���.[�i=!�D<g�ȩ��Y%rt�Kկ�q9!�� ����[8nhQzWL�+�h�"O$�+V�R�m�d��&$p��"OJPv�����Ct��'T�֘���'��4S���әf��m��F����x0끕sG��ȓǴ�Y7-_&W,��:w�U�k<���&%��fNu�C�W�@�ȓq[�<�1��xx��
��k�2�ȓ������J��0y���0>�5����H�-�zӦ19�.Q�/E��'��`	���5Qʉ��N�,�c�&%D�`�֫��RJ��B�8��HƧ'D�����D�R4���� �8D���rFAj�r�t��TF���T�6D�,@pM	�3ۂ�cT�T��	��5�O4� ��O��q���(l˳*��A��0ӗ"Oj(p� ]�O8�k'hQ��\�3"O�\8�kA�=S�H*�M(j$���"OTq���E�2ے���K�yK�$S�"O�ဎ�edP���	$�&dh�"O�q�燞,F4��Ek�����I�8�~���ѳ	[D3�"�9
��iv�u�<Y1j���Y�E��#��|�&�n�<���� C��h�"̮?�JpQ ,�h�<9pjA3x����*�;܊��� d�<�g�ܕ
��MC�$�'c���� ]�<���W �ʡyk��<r)P\֟(��E#�S�Oux�HDHԷ��e���H�"O�И���&n�]�CCE�XX��"O��҆J+��i���q�>y��"O��NY�3�E� Q=�*���"O��Bd\�@�a�3�p�CO���.�'  9��ٳL�e�4m�O>�'f$�'�5����� _"U)�$B�#�(��
Ů?��I֟ �	��2�Έ;�ظ��A�:T�z��|��Ft��tj�7[#4���?K��L8���k��u���ȾA�l�m�!�����E�0�DqȤ�T,���`�}�'�ȸ��?���癨?Y����η{���բH:��D*�O�q:�T�7���X4�T
-�NEYA�'[�ʓ
��F�X��У�*R���'e��S�b�R���<a*�r���O2��?�}xp��+�p��!��O��r)�0��$�1��/렌�)�l�<Y�͍�E!ni�t(��r���̓	�4l#��R=x�Rm!d�r|7�͐VQ>ay�`ٌq��Ų��Dsp�{ �h�� �*�O��D!?%?��'{p��4&C,e(R ��A��|:ؐy
�'�>M�����&`��o�b�ۉ��N�O�q�/�5;��}Z�.�X����'�剳2�Q��ן��I��|����k�&O2Z(s3dK�Vy�(��Ё�~ȃW�'h�#fဪh�L=!ʟ����J��4�T(Ǉ#8jp*�vC��l���A���}��4�O���=P#�#.�Q��և_(�I�n�s~���?���hO��	I�!	��<�`(1�����(B�I<:D.1x�ox�!�H�;0�˳�'h�#=�'�?�,OND)@"dm���Җp:���X:B���O*�D�O��Şc�����T�SÒ��d��7�*%�B��^o2P*�~'�D	 �'?��{�쐃I�K�Ńy������.R�ȍiG)�+f:�\�d�iE�l��$ܹ1��oЀT�܅��&�P)�=9qS�|���If�'�65�4�1%�#t(�$8O�X�'<E/�� �J�,Q�M���,O��l�T�'ցp��$��(Gudh"KW-Rm�u�� ����'m��'��Ǜ=pDp�$���e������O�B7<F�q�1��a��,S���@�D��@�b] �]m��
�, �Û�H�
��JG#wnܑz��DN�'C~x����?���4�'����慐 :M��3�Ȇ��:�O����CO������Yf��	s��'0.ʓ)�T���(���-��#_�&\ؖ'�&t���nӠ�d�<+���D�O���!Y�#��5�J
a���i���O�uC1��%f#v<��ׅPa"	�)�6����e�J�E٘Y����7��u�B� w�]�. Ls ��M��KK�O��aaH�*��{�'��YA�a؟'�b�8���?	�O�O��)� 5"�k�`�rM�c��px ��"O�s&d�Yz`y��(��$�퉇�ȟ�4 �k��aeoƖZ��Yh���~=�˓�p�2v�i����'>P��I6 ��Ź5�է1 h�	%e�hv8 ���?�1�H�f>��e�Ji����<P�&1zB��Hr��7�r}JV�~����Y_`0d�b�4b*�ɓZX�T�S`U�x�)�$�ʨ�*�e�D��ٟ���R����$`�61�j 2q�A�/�lq�"���y�b�9{
r�Y�$�����G��?IP�i>U��G���W��`�Q���H�.��5���Dՙr{6`�m�/�j�D(E�n�!�$ʔ[�8H[��M/)D`S�G
�m�!�����*�─����,�!����9�f�W
K��Q�-Ѓ2�!��� ����(�_�"�A ,X�C�џsci� ����O���1��̓#vM�eIC,�|�����D�(���OR��;���9G��B,J�` *�'K��jXw۔$Kt�۠�ܤ2���T!v�+��$S	S���*� �d��I@�hOq����%(��r��x>4�Z�̻#�H�D|����?�5�iVГ�nH�햟fO���'J��*3t��3S�\�	o�𰃫��uqt�;��.w����Rj(�Of�'x��J�x�M*S��>O�Z5S)O`�צE��Q�'���O��h�b�(7�����эssj�#0�'jўq �
�����Y�(�@�)��eO�c>��I�?3���(�+M�$PJ≇9�M��X]�y�'@>�����?����?��'L4�zb�B�+�Hő��W"�)"�l�)x�F�'���Jg�'E�B�6����u��#�1g
l,�T��|�8!�v��.~4�}P�@�O���"m&��Iĺ+��?����?y�'DD0 R�õE��KG���S����D��?��S���+���yrf�5�����S�_?a�"Gs���q#	?�$�����Oxx9��'��HR��~�'�?q�����y8@�y J�1T�H�he��
I�lL���'�d���?�ɇ��?q�'�Z����M��T����Qf���'�ܷ`��I:�!�"��&:O����'�bĔ ��I�O6�$�B�鶄̟{�*����&S#���\"k���	�h}N���O^%���?��'�T�x��M+�gǞKtD�cF��j����*ޑ �n�d�i��$֖9-�7�	��]��;r����f�^6�`
�+|��ic��3c3����9`�DO8;oR�'U�$�'W�$�g���ƮO0ɺ��X�W��ciƅU�L6@�^�����<����?�|�' .�'�,~%h���)e���ئ"O̭	g�V�^��u.��Yny��V�0�'��'�'�2�
�G*n�T�ϳ2k�u/�(2�"=��T?�Y%ˇ�1�4d���[ !��,��+D��`�#�=x�����J��2����)D�|�rH�h��pՅI6"b���)D����	%E:8G%e�A)t�"D��r��Y"L�j5h ��2 ʢ p��?D�ȃc�Q~56�`qAS�m1��ɐ&!D���~1\��u@��%`��Ă�U�!��ϯz9�e[ y�2}��/qy!��X�z�<�!O�Q�谫�B �ip!�$�<�3%�&(��SU�RR!�dֲ�V(r�ΰ;}��d#ð2���E{ʟ�)�L�6t� ��� A��"O`�[S�C*X�u���ŌG���c��D�,/�Py�n+
�x��&	' 6�Rҏ�U����b+�5~�Qc�ʍ*C  ��ō�:��S�2H����D���h�P�.�/+X�"̂4x�)+F���
�j1Ȁ�o p��0���B8X�/Q� �$�ZF�D- ��ہdi���s�̴^J�0Ӄ�ԡ")��z�ݳ9֛��?�$%��m�?2�i 5�Y��D�O�Ո�E�O|c��gy©$�U��V��4h�e�R�hO�)��)�S*a^ő$+���Z`��aVOD����'�1O����W�n�ze�F�ɮ��B"O	�@��|g6f�!�V�c��'u�<�"�/y�$D���*O�f*��?�<7��O��$�O0��E�"�����Oj��O����������Q H�������>N�%Kb�"^
^����
��l���;�����N�*���P��a�v@W7~�l�Y�2QtlǮ�H���F�)Z~��ER��J�I�<$�Zؐǃ	�S�0amZ���$F<�O�����R�J�r������d�Jgゝc�!�䘧*�Ҽ�b�B]Rd�&�շ��c{����Od�!;|��N�8 ł�"v�� L�X���*-�z�bH&Д�"�6f?�܆�S�? �e�֮��`p���� ƈ@ʒ4)�"O>�ҩY�Q�੃����W���"O�C%e	�^/�z@�Ǚ^�(aP"OVXB�&�0	U x �=�� ��"O`Q��JA�r]S�n	2}���a"O�`*���@���Ц-�/���"Oڔ�tK�7�"�����.]��"O��#�S!V��5��Ô1�P��`"O�iXŎ�P֪��(^o���ж"Op���g�<��1 a�0Y8�A0�"OJ��K܃(j�YE/ ,�	�"O6�q�$��gM�d)5d�2}L����"Ol���d
���)%S$��}�G"Oj�3q������bmP9:�аr1"OBԨ�D:���S�$X�|W�R�<�N��W�~<@p�2{@ EHO�<9dmH���(	Yl���tE�<1r��
����P��/�t�Ps�E�<����]zLA����+g1�u�2�W�<��ђn���1U�lSv�r�%�z�<������a�$�$@����#N\�<�'	��S�P`��#�M}�)1�N�[�<��e\�8M�ѡGLP/D Je#�/�Y�<�p��b�gX()����E�q�<���>jE�ԯT2��L8T�n�<鑡F6)���#���/B�1�en�c�<)���9G�P�����S���K�CV�<�S�(\�	��牗,P����BY�<ن@D�PWj����Mva����I�<��.P�_��iyp)ѓRlh�$��A�<�V�'R�Z]��߹]WjLڳ��e�<��h�6�Ass�G�K�n�2�k�<�t��+4����F�M�x\� ͝j�<a�MN�@��@1R�u!~�P@�/T���v�X@|��h%���,�����?D������9nM����4X�:�yK:D��* ��J�(�cb��7;C�9�j2D�@�1��6EህB�i�%���L-D����:0_�����_KՓ��)D��d˜���@0,�"}2��j�'D��8��U�V��b�D�5l[���)/D���!�U�V#�-;�� Y0>���0D�����E�xh!.#1� �:�/1D���񏏓$P�D0�*��RGָ�6*0D��կV��q��,�����p�� D�\JFi׋]� ��%��w�\,�I2D��z.ӆ2�͚�#�:@YQH/D�8���X�`7|���h
*s�����*D��s�.�	T�$���F�\6��ƈ)D��rG�r�t�)�C�6�ڼ� ,(D��� ℐ.�@yɴ�S�\t�X��%D��x�
��"x��!��=�U��c$D��i�!J ?����pʓ�N><�� D�`�"�4jc��a�)~ul�d+>D�Xrrd�4/\r��*�	���tk)D�Ti�'�^Xp@G*��Q� ��ӄ<D�<)���R.<A��! �d:��9D���פ�k��M����ll��^<!�$X<W<μӶ�$sP�4�<!�$�9 A������}bh�8�ʚ�|!�D@��$����3dN-�SZi�!���!ܬ�x��^�XN�<��*�3Y!�䆀[�؍A�h��ND�Y��	FR!� A�b��� M�FP�3G�	
3!�� ���s(Glr*��Bh~��B4"OZ��'҉��i2*�2cz�db"ON���5&c��s�Sc�a��"OT����ג��rH�)q�Iۆ"O�	���^az�Ȓ��I��"O�`�C��+F&-��̐'
L�"O&���,Ӊ.�fi��K�]v]3�"Od��G�N
$ ����"�����T"OPT#��^�IbO�H69"�"O.QJ�.��a=-����R6���"O,�J��@*Plz�m�?*��6"O���0��F�����%O:xQa$"Ol�����"Yb��RC�N
�$X2s"O�a2�F\�SF,J-8�"O����Bˆ5I�9ӗ��<Td�"Oΐx�IW�j`Y�#ś3$�� "O}[���0��倝�Y^4y:t"O^5����U� ɹ�&�=N���"O��X�bW,� �����9�x�"OĹ��(݆-T�a��ak.T��"Oj�M�*�t:�$��k9�i�"O�!ԍ�ql�K��I*/�@Ct"O�h�gS� P�H���zl�$"O�	b�ݱ+$�y �;p��"Ot9�b�s4���)��"���Y�"OЙ0�$�{@D�7OA�tNu��"O��cg�ަ$P�ݪ��i�z���"OJg�2Qt< ���%B�����"OZ8H�	��z�(��=p�� �U"O0)x��-ԂMC��,(��"O���4,�V�1�BնJ�>���"O�1[��ߊ-лu�Y�Y�"a(D�\��j�p�hy���ԲX|�d�WK,D� ���
�v3.�ÄU:-�xT���+D�p8`���9)��2% 3W���c'�%D��!��̒S9�uۓ��*=���a�%D���M�Ov���gn�{!L'D�8#�P�ZI�����A�j��8D����fX�w����kF�<�`��F�6D�X�p��7D�ܼ�ED�Wv��C�3D��ч�P�kv(�g� 6XS�/4D�B�Η�w��Uc��(�'"3D�3���D1~��סU�+�� D1D�l�S�� eB$3�B�?��ɱ&*D���	F�.p�q �`>N�%X�'D��آN΁3@�L�i\e��#D�ĺ��6s�������ra0))e�"D�x�K߄bѺ��u��F5�#.D���`#^,;R���E�V�4�B1�ǋ(D��qu�J�~��<��ϳ{f*m��G4D��!R�&��)pLM�/��k��4D�hhU�8�z 	�Oހ˜æ�$D���葩(�4dqBA].�$U#D�1DKݣj�0y��R�dt��� D�d����Z��Zf�Ց�"D����[�oք}�A��.!
mX�&D�P�29�0
��x����'!$D�(���5z�̩O���Y���!D�� `4��|���	�Uc׀+D�,��
�5N~Z���� K *D��J��Z�(Vu@�ʎ�9���*W�'D���$(�M.���
ɿJ:�I�N'D��s�B7S�T�w�0pp�R��(D�x����JBDH��N�QK�98��'D�� �04�T�L���u�+�xY:�"O��1�
��!���3.	s�yc�"O⼉�擛.��i2�_H\TA��"OZt�4j[7b,�٥��D�Ȅ	�"O�,x�.E	�Xh!�N�s�$�r"ObѸsB_>N�䊲L$�`;c"OJtw\n�PY�Ė�f�*La'"Od}p� ��J)@��Z�N��U"OĀ�� iB=��JO��ܙP�"ODJW�o��M9fI�#b�h8�"O@<zc�l��� �� F[� +B"Od�B W�5���"@�]Y�ع�*O�M��ē[��@z���R�(	��'�^��!���tu#@�0F\��y	�';z�����<8+���嗔S��y��'y"��WO�}I���7�v��'J�����E̑��� /PD]8�'�8	KR�Ϸ4�J��!��4#@�x��'�$ufϘ�a3R@��%��iJ i�'5����d]7��I�` �o�Ă�'�N4���"2��Q��x���'3R��9�1���:s,!�'�fa��9a��D�V���6�Q�	�'�<l��^�2wй:�N��b>�	�'}��珝gyΤh���":HS�'$���棝�c8�P�jǪl�d�
�'������}�r(kC�I/8���
�'�0�`B8CT\��V�,Ǩ4	�'�ج��HP�,0��٥ye���'o�䫑J4^� �'$_-c�\��'��qZq/y������W���@�'e�|�m$E�PC��O����'s,��v�	0�F� Ǝ�1�d��',$�2&T"8\j�ce��/@W�� �'�p��%�b�Z`j��2�>0��'q�PC��YL����遵X�ݩ
�'���x+��}i�����Uo���'z <��H،2�Jd�1��H��'뢡�'Y(~����$Q!z�'R�æ���q�lY́� �,D��'ƶH0n� #����A�!t_l9i�'���k�싲}
������re��3�'���(2*J,�f�p�k	5jI9�y�U.�RBfѨm`�
7č��ybi	�%0���	_����F���y��$_��jT�;Z$�T��ŋ�y��JU��+�I-Y���H�y�΃�ƚ�J�M$;p�2MV��y"�Ǌ����օ�(s��13T
��y�l�;K�a����.���	.�y�nΡ` �Q��%e���cJ ��y�&��P�Q�˓�Z�\���(��y"�E�|�9r�nR|��������y4Tu��b�eFM��P�ٖ�y�iWKU�HV�שBH�|j�
P�y�ʎe�QB����= 0$k�ҹ�y2(�<5yfɍ�`.�Q�f��yb \%0������\h���e�0�yRd�,�0��3h�Z�	#����yFJ�S�@�uHQ��Ɋ��yb-�"7c��!��}� ��4�y�8}�(q��O	�U������y�eFsw�e�}�&@���3�y��H�e�B@����r�̜��L�y
� 4�D�$35p�QM
8Z�h�c"O*1�bT	)��pL��7��=�t"O�M��͈K�:���kWG�~�B�"OtS(`Rr<���Z<Nh�`Z�"O�e�$�MM �S.�=.��'�54��*r��a�V��F�
���M,D��ÅKL�FSq�ŉ�!��)�B8D���c�O�F�T�֢4�r!�a%D�<����~���B֊L�2�F�0D�ȺT�ݑi�񋇡W��,`n+D�����[�?,����XT�X���*D�8i4�E;�e�#��!�7D��T��r�Ri)h����Z��8D�+�Ϟ�bL�=��ᎉ(>�*��&D���T��9e}h��聪�]�6N9D���+�1���3����J��� �&D���f�Z BJ�bD��C
�U� /D��P���"�����bL�b�X<P�J*D�� t�FA�� PF�ưT�̃�j)D�pkU!Q����B�%����"D�h�5aR�U��,�V�љ&� R�<D����B`��Y�P�p��@�%D�H[�eK%��p/�޲��R�&D�L�ÎY�,1�L�p�]�X����$D�t2�'I�z.0�q��}	+�%D�tTF�88j��En6�����$D�8a�&i�5Y�F�f����#D�x9��)��SԄ�.✁ J/D�89��D�[�(��"K����U�0D�0��@�'��kf�����*wI1D�(���-��$@Ư@��J���a;D��K����2������=#W��B�3D��z(O,`ZN|����'%A1�	4D�����8Q���3fAE/H�DQ�`�7D�  g��~��l�֮�31Z��1$b;D���5�آ`ࠤ�S�A�J�6�'D� �d�۬,wЍkP�ҋ!�fqJCj1D��0WE�?�<л� �@&��W�>D�Xi@E��n���$
P����w�9T���4Ù�I�Q�c-M�90�[�"O~5I��Ϊ%��)(DK��\�н84"O���l	Q��)����YA3"OH�,���h�A�j��JP	ק�!��ƙ�:�CQ�=���*�a	5*�!��Ġqx�%����x��Ak7 
.m!�d��
�CC�ŉN5�8��H�z6!��G*%2�	��șW�d��I�:R!��� y[����@�0�4�ZsE�)E@!�DGIGd�*ah�n�ɖ��:�!�$V�y��I2��6>r�8ȱ	R0k�!�D��%t�p�Z6:��+��Ŧu�!���=c�ny��Ŝ��=Ywa F!��h���� ��&Jf9CCaƓ:�!�D޴Q1FLIEHEH�0��D95�!�F%��iX�?��	Hv�ܯ|^!�$�
i�X�X�%҇f�����_1|!�ݷkIB��Ҩ���nlcbƚh!�d̟z�x��p�
�v����o�"8h!�D�9Il��D�ԛ*�dxan%:!�	w�B&-��$X��g�qg!���]�0��G�C|�|�dHK$C{!�E
�`m�&J�h��!U�!�Z ,��'��~~��8�
I�!�Ę�T'�-��d�JSN ����$>Q!�� �k�">�r����!��S�"O
��4͂=y�@�0)� sĜ��"O ɢ0�TR]X���nQ�x��Ӧ"Op`�v
V'�@�����g&	 "O	pU(q�,{vM͂��`F"O�Ɋ�"�.Q�1JS�� �m	3"O��S��+7B���H�	�"Oʡ�u���^��v��0q.�k�"O��(�%~�h�[�"\�2m�4"O���O'KS���!�1c���"OR����9rb�JG S2��"O�M)p�Ӻ,�=Z��Y7~,>�z�"Oʜ�t����H��&>��IY"O�!K�@TkiBY�'*�+'��uS�"O�E1�(�C?bdPfhUr�ƨ	W"O���D��RA�0(\#MժĂ�"O~)k�!�	RN�jǯ�;88��C"O�ɲ�a1�d�so�#<H@"O��zDj�[�(8�gK�y�2<�"O�:._s�:��F���t��-C�"O�@p�&�SI����狵{ÚH1�"ONIq�+Y�iN�!j3'��%���1"O|�����4��t���	)�� 6"O ��A�Q�U�LQjd�^/�0"O�x���5VUX5@Wl�-' �ڇ"O,8i��OgTx6�[���j� 5D�l�7	��k�xD�/ET���'5D�����d

sÚ2T�25SĦ D� ��݇~�@�Z�M'�:Q!9D��(" �ag��D����!�#D��X��Ӊ2��f�1q���㒈'D���@��=-��	�P��\q"�&"D��� O�0i"<���۪,e4�Q��/D��Rce\>LD�C� ��bK�\k�D/D�X����1K�&г㏇��� $�,D�`���>S�Ĵ�SG�Fjh+Ɖ*D��`Pl�!R"(�P׏R�5�\9r�<D�p ��3,\J N_�=�\P�:D�d�E�_7��]B�#߂A,yP�#D���'�L@�ʤ2DK� 3g%���!D�0�@l�4���7���2m2D�L� ț5D5R�Cd/c]�Bd�>D��h#��uWH�`��żSjd,çJ=D�p��B��XYfd�$C�}���a5D��'MA�D�xp��Ǡ�o/D�$��˘�T�2-��M�fUx�:��9D�zV��_�|i�d_A�F��Sn#D�\ڃ���p0����W�5�h� 5D�0z�&�d,���!�H�~=� �Ņ D���+���Vk"n��Hb��,D����F�#8Z���L�����P@�,D���S�|s�Ȩ�n
��q�� 
o�<1֌�,
�N("vHӠ_�J�v�a�<�_L(*��]z�εI�/H\��B䉻s�0�C�ڣ;��H,lY�e�)D�d�.&���J��4�V){u�<D����.����P���-��"�9D��:4'�?�J���ָD�@��d�%D��2bg-�(��mp�r�"D������A��p��E�R`�G�%D�H��EA*Y�<iҭV�k��'*/D�̸���bƐ���iDm�׮9D�@ˣD�V���QA�L��T8�#&D���Bf�=mev�����2R:B�*#D��  �G;/x�|�a�� <��"O�y#%�,!GT���-L ��"O�<�G���WG|��v�B%(*ك1"O`��џ_Gء�a�(lr""O���s��y��KV*&��##"OTt0M
�:s������Lf��g"O*��E��r�4�hRI+�([�"O����]�9�T�t���-t�Lk�"O�I��/?F����)}.9Ȃ"OŐ��L��t��hZ�mv��Z�"O��C�#0ؐ�j�e^�L^tp��"O�ez�O&Px�����N�(U�9�"O��1�<<��Aô��Hg"O���BK��Fd�yq���b��c"OF��!M	����!q�SX�6�@"O(\;@�^%(
������LAV"O�`h�j��8Qp<p�-� ���(�"OpI��g�t"J�[�٘}�Ԙ��"Oz�zU�B�A���3W����@�(�"O����T�x�,�ؤmQ�/�&��v"O�!P���h� r#kM!(/�A�""O���`Y���
���b&���"O@!	lڗ&��9����X���"O�${�䅭/!:��d��? \C�"O���Fa�$[�Z��Z6� �#"O@(��iL8�qi����*x@I02"O<@xA摋,�V 8#��.v��X�"O��K3a
"c�|̱W��0���b"OnY����%��B�fŻK���"O\񋇏��I�4���E�i~^��A"O.����AM�����W�Ka �@"O����%փ'd����Ǯ_F2H�'"O y��S1I<�9y��غS܌�y"O���Ɓ�P*���ǡS�:ݡu"O
 r7�����Z�#8`&�Q�"O0I�
�>�\�v	Y(d�I�"Od����?��aq'��p$@��P"O������!��Hl���z�"O|x�.�!D�t�2䏘.I�DX�"O6�PC�g�԰F샾L�6��"Ot�9Ä	�:��As�M)��J�"O�u �ڵ=�F�Q##S*>A��Y�"O~Q�H���:��,T����Z"O��s뎴�����%)��S�"O�ˁ�#�p�z��[�TjZ8��"OX1��T5���eƘ.U�@�"O�}1W�-_�<��$V6yAlH��"O�ڦ������J�8���"O�S�Uq�Ր��ÏO��"O�4k�ϔ%]"l�7�V/3K�K�"O��a0�� �����¿oPL�e"O\,�E�Q�8#¼I��j�r�"O
 ��	��QV.�6Y�&"OE�7M���ّ�L�I
܁��"O�e���%�fp�0zʑ,�!���e�lX�n��)
�H�c��9%!�W�n�j��E�@"uW�Y�F�*S�!�N1lPD8�CM"]Kz)�ag��I�!�$��'R��R��I���$ �!?!�d��DT�딝v����Ə�i!!��׺.�B�KVe
�(�()˰�@�?!�ė]�1�ҩ��}u�f�� f1!�7w
.��F۳0��Aj��A�!!�R�xn��""B��,d�
�.u!�� lȀF`��fU;��Z�/�T�t"OƼ�Њ��j���\�=�>�c�"O��x��O�r����a��G�N)2�"Ob\[�@�g8��Jv��.A(��"O,Ѡ�iO/��D��"_pԤ �"O��fߡM�f1I��ϳf�)�U"Oj�	D9�~Yb�Q�NJ ���"O�q[ŝ�R�ұѶ�� jEbYj�"OD9��EΉ <.���@ā>	X�p�@<4���+�0$K�%�/YB<|;��$D�d�gJ�Z�>!�q�R�&��%M=D���I�f�a��' o`��¥<D��	P��igR`-�&�D���<D�t0%ビV�2�їhХH�&��CD>D��CG��B
69�L��2��r0�=D�l2�k� 0ä�G��r��8D�t��U�#�0�1�@�$(�$ʲb8D��j�Ǆ2WO��P���x��Q�"D�� �>q��� �_+�N�A!.D���6�H�5�c�R'e�4`:��7D�D��\>l�t� !��
�F�D�8D��K狑�IrԠ�)�!����4D���D��A��8��*q� �Zwo4D�:3�?�&� cD�<�� �c�3D�$j�O�k�H�Bw�uA���U�4D��y�o^	bZ����	�vkG�1D�L��=a�X B-�3�^! #D��*a��BcA��$	�b�;5�=D�h�5j�2$�Zi
���t�x4�C�.D�4����n��噲�M�9CRԛ�d.D�8��nS6.���1k�@2t�A�9D����S(rr
�a�fţ.�*�F2D�P�b�i󠈃e�@ ��%ô�<D���g�]7h9h*"&�Y3��;D�����!Z^d�D� m? A��8D��0#;92r�qfk� ��a��4D��S�*�/!��y�B�f���S�'����+붌�.��]��AJ�'\9�h��1��-�0�,'~�b�'6�P�7-��e�8��u�K :ʝ!�'��BC�z=��+�*OJ0{�'w�H��H�w���`���A��'dQ��j޽�B��!J�\`}��'�^��fC�9*b����OU�})�'���8�\�OxX����S~���'5�t�t�C�	H�u��-��N�ɱ�'����%VW�A�K>`M�'�<)҆�HN�}��*X�K�'�&�QPl�b�(4��/Iu-��'����цۀ?�^�Z���~���'�\��gN�xP�hg��;u�*�'��0IVH�6o�F4��M��}=>,I�'��ق�b���$��>>�K�'��v�L1�����0(�\��	�'k��� �6IѢ9�陰%����'����y >p�dEA����'(��i�@P�6�>������
����'��I�։�2qk�9B*�|s:x�'�,���eГ[ ���-Ӳu���'����U�'���8�L_2uf�@�'B-)�'�I �ؖn/C�V��
�'�F����5ph�c��X0��-k�'���"DŢi��r�O�
H���'\B��f�*��ő���#��
��� ���dH�^��H�dS5�2L "Ot@�Q#ʆq����)l<��Y�"O�I�d��{RR���I�qK�97"Of��N.8�y;�(�MHF�K�"O|q����hI+"��5\�逤"OT���D�_�-�e_�&���P"O�I���w-�L���\�l���"OLX���!J�b!�Vm�><T�p"Od=���U��Zhy2�ƀ@:��u"O��!e0����D&:�P�A"O�M�2BV�m$dp�Ȍ#Ar%"OD$�s��>t^�r��^�j�""OΕQ���Q4� ��8�R�7"OH0)4`O�77`���.�>�P�"O��tCϿHی�A�����Y�"O���cfȫN�6��%*X<	z4�R"O ��1M�7xґ87��^]Ԑ�"OԽ9dB�q!���A�AI� т"O2����J �c5�Tr�4�("Ob�!��	�~��<�E�E��p�'"Ot�f%K<�̰��!�>M�z�ۄ"O~0��$��'<\ �� ��aÎ�z�"OP����ìY,�2���'�jTy&"O)1eg�=�N)��ށ,����"O\�"�@=  B��Mۭ_����"O�)�P"�+v�xy�����j�"O�%���<d=x�kǊP}.�"�"O�2G#�� ��*�� �th�"O�s/
.9r-�_(�%�P�l�!�D��p�$��i@�Qrq���%!�dU(�
=Q�{�Ni¢�> �!�Ė(z<��5����1���U!�)[�Xْ#!=����`��?�!�$�=_��p2J^#Fth\��N�)-6!�7k2]
�ɋ#6�-�pmɣw%!��i.�)�.w"�˳ʖ��!�ש�\a�`+��w-�����x�!�D՝#Hݠ4�J$v,��q�G6-a!�dV�c/PiHБg*:�Rg.�!�45�&�jGϺ[���@,�1�!��2xe�"�L}�AqIM�z�!�E8�v��ɭGo�����62�!��i@��u�W2N	J�{�b���!��X@�&��ԏ�T�x�j�U�>�!�dI�vy�,�)�;&���QfAʱ_�!�$�5i��Y�wO�Y������ƕKO!�$��Q�b�SFE��!%�\8��E4?!�D�'H� �PU�ל�$X/	!!��ЀrABI�E�q��t��nH`�!�$N����
<�v8ӭ	�+!�D�%i��M��۰vʹ4YwG�C�!�$L.!ߠ@H��޺%-	�P�H�!�DԾذ���������'�!�D��9D���lQ�I�� i�?<�!�U/^4�G��Z҅�[X�!��8'�,��R:ޜ����j�!�DO8t͠��s(�$>sg��n!�D/.c�|���W��{bF�Q!��,����g�]8�B���$,H!��(.�;���~�����'-!�ۀ? ��@�/t��YBA��,&!��6m�
�UϚ���IS$��y�!�$A$N5��0h����`��(=�!�D��]��̈@$F%��](�K�
;�!�� ��& [EB|�#V�E���S"Oj3�LM�2?�X��%L�8�L'Oh�D�|T^�QfJ	�b��ZD�T��Py��,b�|�+kEt3�5QԦ���y$]
K��'ʻf��q�F!���yRn�&KjQ�PA����	Pb��y��/�ĉF�ԅ[W���p��8�y�?~��r��M+t>���M��y�M��%	�P�W�?:X��MY��y�aZ�b� �hq��1���0E��y�!�/, Z9�F�^�)�$1[Ѕ	�y���T	1
Y�x�!'�;�y2�I�.�>M3�)θF����fb��y��>=�p�IP�t�
F���y���Yp
8���IK�P�v)^�y�	�.�~��׊oU��z����yr)��E�\�h��C1c�Z��O,�y���8< �Aӓ�l��S`
�y2��0�0��� Xq��Q���y���%T��#����
Ӥ���y�B5��=��
P:M>xmP����y�˛���� S�BY$�(���y��	�ȵ�v�9<  `cL�*�yB�b��9�b�C�/u�jw�ԫ�y��G�}������#=Z"e��A-�y"ߵ$f���׼3��遥���y"a$GZ��͊$~N9��	̈�y�k_�N�"Sc�����7���y"�[�d�|ŚЎ�7t�f�ؖ̒��y�%�+/H"� E�v�\Y�a���yb��`�D�:/ղiZ�] ��ё�yb�8��Pw���L�)X��y��N"9�&�q���' Mb Ѝ�y�ŌBv0��$K �����ɽ�y".њJ~�zDK(b8>z��ܧ�y�)�ti$82�ǻ'Vqs7뎻�y�.��qu.I�UQ�UyL��#��yC��h-h�ٱ$��<!�ջ�y/��t�R@ucÛ�� ��&��ybKA��`D��
j�	�S ��y��N�X�
9�fB�4�Z�2��y��^�o`*��d�۽2�F����yR�I�}Si���,g�]�-Ƃ�y"(��.���z%NϢw� i���ʔ�yªJ�|~�<��Λ{�n��G۹�y2$�!�>4B�%�g�tAZFN��yBɟ�o�v�PѬF�T5�yzf�^%�yrg�r\���덊U�,r���>�yr�L$R��d>��*v�A$�yB��+��� �`&��4�~!�'�ژ�vE��(���>2ҞH�'�z5�u��t��)t
E
#��`"
�'Ў���ώb�l�(�B@*p�صz	�'��U���R ��hU!��hcd���'A\���.n��FW6Z]�}:�'w��˷�	�R� Tn��<d���';��C�`9���aVE2K�J�#�'X���@��8]�(�F������'{�8	� �(��DɁ
i28�8�'��-kV��L�䙢�g�s�'`�A��lǷ8��3��2Z�u�'���E�̩�lH����:��Ĳ
�'����HXC�H�rr��3gt�C�'�f�`��K�wwb�;�@�MR��	��� @���e��a/R�� ��!X~��u"O�,��ݝi.<0�'�/�B���"OJ������B�(���Y ��5"O.�x�N�J��(QD]����"O�mr�Ό�,��q�B��R���T"Ozܢ4��R�H�d������P"O�0��*��S@�a���G}�b2"O��Xi��F6 �B�(?ZE�]�&"O �A�A�<Uh&�E�
�8:lL�"O�i�G]�L�ܕ���B9(�9�"O�#S�$g�	�SxP�:�"O��	��C`!10���q��Ja"O&�[��ƣ)�+)\!D��"
L~�<do�"{����U"?��!�FB�<A�d�M��A{��_��%�fJ@�<I�'�R�,�b�����@�2SNS�<I$�e��d �a��ž��r�Dd�<iB׃w|��3�F?ff�Az�[�<A����YX���l��:�d]�<�@��*0p�2���xA�pB�,Xo�<����_~L�A ԣ1]�)�D��g�<92�Z�<3:��QDݟ?�ڴ��H^`�<Q��S�	�^�C��=�2����\T�<���{ 8
!	�4�RD�r��v�<��;,}���Gµ=����u�<��jA �`*4
�]�"��E�V�<�t����I��̣W��@3eM�<���� �-y��!1��u g��R�<y7�)Ad�R���xL}�CaO�<���7J�XR��@�x���ǒI�<�Gf�{l69hd��N�qr��D�<��W����R�Ĭ��)3Q�h�<I��B��{���+B���"Fd|�<1�&QH�%�@�n{��"��x�<1UCZ&�,Y�O<�:��2��z�<�)Ǣ|��Xq�G�Ctf�j�AK�<a5�G�kC���!��S��1�.r�<)�e\���yy�l�-l���U�h�<a�$�=�|�Rf�փK�bq���d�<��mJ����G�n��JeLA]�<	�L�|��� Q)h��L!���g�8���y���܂9T^�ȓC*�g
��.��J®�[�FH��uXV�I3AѣW�����?D�j!�ȓ$,��`�N~��Z֤��H
���!i\����aJ�A��ش��L�ȓz������4P0�$9�ȳ48L<�ȓCJmj���gcjpH5C^����ȓ4�b�\�#��4�)���ȓc��y�BI����0h�+�f�^���[l8Ӧ�X0Y�x���B&Eb���?��,8��
�2�4�qV�5ܢY�ȓ{,\�@C��@���i��
�Ej��ȓYe 眠38-yA%ܑO-RM��@Rf9@�oO�l��(Z]���ȓy� �BaI��O1~�+��쥄ȓ��`�@^#�PcSK�?(�t��ȓ�3�$_(g�\}�d��mc>��[$$�7J,�ܑ��H8Pp��JR�E�r������`�+!����j0	g�Z�ij<Hv�J*,|����B�~5)��.g���g�){,�	�ȓD���&(2��ѐtjΡ!��(�ȓP�ޔ�2�W8T�6�xa��! �ц�S�? �͖�l>&BP�#>��B"O�e�᥆�b�f}�%��'���"O�	�u��)-�yb���<Դi�"O��(��ж|bR�dB�G�
��"O�As֣�el~���J7m���)@"O��1�(S'L� ��$���+��!�"O���D��H�,�QU��n>�5"O�4c䩀%^z�A��0^̼�W"O��Q$OG,��!B��ZE�Tbr"O��!����T� S3E;_Л"Ob�P�1u{��Y�ڿd����A"O��C�Y�1�M�<� �!�"OD��#e^�fw(�职S%��Z&"O�5�D�
���#��1#"O�hN�:�������X(�"O(P�ݍ �a�� �2�"�@d"O��2�k�:R�ع�<j�LѶ"O�����
;z�"���i\'V�hؓe"O�u�-~��lw:�"O�}qQD2�Ν�!�\Ќ��"O�yvcW�ORp��I�^Q>%�a"O SsJ�����iD��'��E�"O>�Y�a	�"�n}p�(�0�Ձ�"O0آ$��5��Y��D2
�����"O���w�َf� ��L�t�Ɲ�b"OT@%N �}0=��	�l� m`��I�Έ�>m
��߳���3,�*Y� "Odp �,Vc�\�K�4$���"OdU)q"��s���3�Ǻ7z�Q"O�$C�^�h-�T뀁.��"O�ɂBN�u�@$1���T�@c"Oh|#6�
@�)X�(	0�J�H1"Oֹ�@��7g(��#�g�H���9%"O�l[%�+~L>Tk�- |�a(f"O�9r�ㄝ -|��҅�=ʉ� "O�A��l�8?�*�`�$�=Y tt��"O���j5XJ�9�-�z!�"O�=�"_yd]���X%�Ũ0"O��Kb�SQPM"���`��0:�"O��2�f� *D��
�*"���"O�ً���
i�ڜ�D���33����"O��k��vN�x��ȃ�R'q��"O��?G>,�7(�*O���%"O6��B��a �PWg�V��P�a"O��hb��0��7L�Ax��"O�=�1HK=30 ��Mdq��"Oޱx�k�3Y������9Q�`��"OZL� ��H
Z(�r ��;h�A"OF	��b�!�v�sD �+ V�d�"O���1e�Xq�\�%oǫ"b}��"O�iHG��(]l�S,߃J��X+�"ObD�D��Q����<�L�x�"OD!06(ٗ7�p�Z�
�L,�"O�� *�Q�$�;0,T;4Q䍰B"O��Q� ��kE�0	A Qd��3"O"a���#f��#����LiU"O�Br��
a{V�5��@Ր�`"O����"Yz��B���fo��""O �ɂ�(O��g�� S� �:S"O-��#�t�˷OV�9���(f"OhY@�ҧ
9��h#/�-�tX�v"O��R-�<�u�% �6D�!"O�0k� ^�D4�S���_�%Zd"OLh̇�w��}�#DʮK�Zչ"O� \�(�)a�GÖ�7���a�"OPy���
N��2�� =�ƥ��"Od�! Kߵj�½�r�
��i��"O
Az�
X2n1��N���`Z�"OT�i�iD�ȅ˱�RG�����"O ����_�4�mT�7��IR�"O�	K�)�"�v��ĭ]�;��P��"O�C�ς�m��{cMM�\� U�3"OT|k�a���P��k�.~�J49c"O��!��o�0���WJ�i�"O��3u6]��HN2lȊ�;r"O���s��?;vx�v��k��A�"Ol��`�$t�@�υ*�ͯ[�<Qu�ۭJ��p@��X"%�݉��x�<Q�˪!�J r��$j��@ �/s�<9�I�?h�T���E#K��S�T�<��I)(><xZ�$Y��h�E�FO�<9C�ߎg^�e���)QҬ�8"ώd�<�A���������D��AHTdEe�<��v�t����D'i�E�PU�<Q���$d�D(�
��hN�u�EP�<YS���P��)�Dټ)��	���RN�<1�`�"tA���!S<Z�u��F�<���bL�p$�� �� ����@�<q�-S�C�*�#��O�!5�F�<�-ͯ7X@�Y��*g���V��\�ȓ!c�X�`�'�2@�����rYN��ȓl3�0��P�P}:}�D��@I�ć����ȶ���8�����.mWҥ����$��M]�c�NUʆ�L� >9�ȓsh�*��V�?fl��$��] Ȇ�Jv&���R ԘY�pˇ�M����ȓfD�)b���N��1��Y�`4���1�\�r#'��}�D0�w��v��ȓG���!��h��a�/�x�h0�ȓC�6${rOƠ���qaO˖�����0�:p$�ՋD��؆�"pd���ܔUNL��`̳��ȓ��t�d�	#��A� +\$�8��褭���=o����"O&�2���p+ �3&��j1�DY�e���ȓp�q�R*C79��ea�� n̈́ȓ,;�l)D��3�Ae�W��]��D�	��d�/U�Ɉd ���,��%�9�G'�9w����s�U��<��qd�+æ��?���X�P\�,�ȓI!�q0C��&�:�gҺ#�ȓG/�Ya�A�NP�7m�8M���ȓ�6�{k�<����/��H��Z�*L8�A[HK����Ó?H�(�ȓL���c�Η9K���*G�&�8܅��z���HſK'� 2���V�ڤ��c20�ƙ٤`i�
�/!4�ц����̜Tt���a?:-�ȓ/e`� A2���H�,������ȓzq�P�`��r�0[(��I_�(�ȓ[|���Y'WX&���� �h��CS��@��44�4��W�?Xt�Q�ȓ{�$�:w�B1�hYU�o�*��ȓyZ�&FJ=Un@��'Q�(�� � 9&�аW��C�<#<��Vt��Q��$o*H�/��8lx��ȓ	� Yi�/)Y��%e�;��ȓD������ٸj��X���͐��d��S�? ɧ�(�f�ZS�ɖ&;���"O��"�(��		0õ'��!�I�"O����+�|���ږ`��!�"O�� b-Q��$�z�����0"O~Q�Q#\%�y���{���"OH�yR��.��ӕn���n���yBk;+\Dx ��p��Q�reB��y�Ɛ�|Yc�I�d��%X�`	�y��<%��Y0%dJ
�*)��$X8�ybMZ� ����W�|�� ��_9�y2�]'4���eS�w���G�'�y2�N�6�ژB���Y�<�	?�y��7�"�f�R2��l�7�I�y�w((��� ��\dK��y�w�y@"!�3}9�Ix�՟�y���8l�4��q�
�e�Y9�yRLK�u2DY`3K ����jtJ��yB�'�a�6�惡��	6C�\PROE�1�^�p�`��v�8AЂ��J1�,X�i6 aÁ��Z�k)�sj��U��\vn��0�� d8;��i���A�m¥Cs&��@"���I�A�'��d����U1Tx0Wn���4H�O��Q#�O��lZ�c���<�������N�Ókŵ�e2�oߩ	�!��˱�欳b��#��v`ѫp���شT��|r�O��_���%F������?(���!��5J�@�:�ƎJx����5l��5;�#@u:��qB?`��p3�DM�C�.M�jڧ$R�`r5.E�T&��P3�/ܡD��1�IF�I����*��4d��QF+ÀK����,��m؈�d�2Z%��\<����0�ٵwְ{�cOKNrQdm�����<�im�O���'z@��C�΁9Z�\�TK�;y�ȓQc�4�E�=x�~�1E�G����Z����ѳi)剉y-,�j^w7�����~	^,� Oi�~P��ʀ��'>rH'K>��K�MPo�R�Eߨw?�|Χ-��P��"�MՎ�EiZ"<�Dz�a`hhX�<Xg�	�g
5�擮c,)(SKF�#�˞�v#J������|���O�'>�l�%z`�!�"�5Y�bǥ۶\���������:��F$�>z���rD����I���O `lڹ�M�ش;���!c���p 醷$3> a�O�!&"���m�	Nyʟ�O��&Ĕ{�8�sgMT��V��=I2��4�J�
��ׇK"^T`xr�����7`[�s[ū
�2	�P�@�.�M��źh��!�����u���Ug�-�~�|�1+	�d�GJ@"hv޴��,v��o�,�����O:ym���<D��4t�n�A�
H�Qs|,ۢf��p<�}���?	���,��,M�����6l����=}��<)��i��6-4�����(��"ڪ��)�D��C�ax,O|�pȂЦ���&I���T�>~���d�бr�����2u�L� ��s#Uf֦�d�$g�M#�L��jTBRQ5yV^�b���m��VQ4�!4]N�4"3h�[efۜD�F#vk�$�Ji8��'l��I��'!67m�.��Y����h}��_�O#
�@�o�jFƘ1q�V��y�N
+4J��O����,WK�|l���M�K>ͧ�
(O��l.dT
�-}^PEx���D���&<OR��!!�Ea��˼q6Q�*#-�>�S/�DpC3֨��!����OPp�s1�����KB�>f1�S+ V8��A\��P�P� ܜ�G~����?���R/IIX�z1�G�a^��9B/!+߆�"D�i+�\���	iyB���/-�@�NL�H�����,�!�8��`I�A������U8?[�����i0�4�䓌?���ēL��H� @�?   X   Ĵ���	��Z��wI
)ʜ�cd�<��k٥���qe�H�4��6X8$<gT��"�ᔩ^�"u�ǣ)z�4�L��M��i�Z7-�Vx�,a�K�[����݉a8�-q��D�Q_��b�iq��a��	�"��6��Xb>:5H8:�UC��Ǯ���Q�Mx�ݴ��	+hf�(r@[�剟R1Qq�#2�HY���:K�De�R�RT�6�[�;����mbm�cΉ>�l�y�t<�FH6���Z�(8C��<k�H��<������l�����U�l�Hu�O�	I���^���Öo���AB�Oꅡ��N6xP1O��t��	��'�^4��-ԒM��1��Z���'"B�Fxb@�W�'r���O�W�Y��@�+g5�&->�9�Z"<�#G�>Q��d�>x�ÎL�^�q v�FM�d�OM،{���P��rg(Eg��W A�M+v�(aŰ#<3L6��
c%���\�Q��Z��Ȝ�>A>�y(��;J�*#e�}���)t��|��'���Ex��A�����l����kR@J�-�,|�!&�P��#<I��O�x�r��g8�̪P��9L����D���Ot��H<q�C�f�H�"�0��,x��^@?)1�8r%�O,�&B�U�M��4y��	�-J���
��IgˎL9@�$OHi�DQ�O�l���(��S��LB���(t,L�/O��9#F30b�'Vp5�� �ēB,�����u���xS�A;+]$�+��/��$GyB%�M�'�����	�`��xH�&�k��X�'R��:@ ������iC�	9�x��ٴ:z�Sϟ������KfJXYcC�ZO�qy )a˛��'j�R��|B[>	��RL�Y+���<�����o"qG�pn��U��m��4�?��?1��qV�'er��v�"��-�@zX��¥��".7���X��d/��|�'
"-�9HI�@�cD�w�DT��/�W#�6-�O��D�O�Q �j�^��埌��r?!����ۮ�8t�ǀp�A�rm�צ�&�prGN�(�ħ�?���?����6*͚���/Fa��/��
B�V�'��L�v�(�I��&�֘�Sv���N n;�L#4C�'*:N�xP]������O��$�OjʓF��a1h	8� �ŀ��j�.�ZHTj��OT��8���OV�%&{��b � �|>P���OT�rN�g3Oʓ�?���?(O��r���|J�D	    �    �  �  $"  d(  �*   Ĵ���	����Zv)Ú'll\�0R�P����=9pn\�Ёba�#������{�<I�d� �t�Z5$��vT�aN�!@ i®�,]Q�����E���I�A���0�2rTƌ�&���L�/xP�A�^�M� maf�E�m�];g�0'h{G��PZ��xv�Ӳ]m^X�S�a���N�y�D�{�e�>;P`���H�F���_<k��ac5���0$���72>���)�-#��d�O����O�e�;�?����$+H1p��Ւ;o|�ԫ[�gS�	`'&��d���A�4L��HR4rP�шw5�	�6����0'("ݑ�<J"��V.�> �ɕ��<\O����(��@*@9����3|r:�"O���$��A}�@85A�.� ���ie�"=�'��+�B(�4��f�D ��,����4R����%+���?���?�������O6���*!���S�F�j�/[�`��p��l�QЊ�0c��_�Zz���[?Q�4�U&�xUXv�վjxƁ�3�:J��X�t�M�W��Q��`�S�'��QJ��gl6�˰iE�|�2���lB�vT��t�i�07�<�I<�H���LH0Yx�P^� �C��y�&��*8�����ɠ��Ƅ����JM}2P�H��G�6��|`���L8�"nӪ(�6�\�g��t����)w�^�"�"O(���ou�J\(^�12"OJ��g�"L�x�&���{pj���"O`s��]�hZǡ�=
TZ���"O08���̹)�y(�B9M����"O~�����q>� �eI��vr4�"O0]��,�a��ə�\2X���"OX�r��4W��Ҧ��;>H��B"OB���#�m���Ah+ [�"O�H��ݎh��8�t�(�(�"O��*d���l�J�qAhU<3�b�Xv"O^ݣp���[�
�ɣ��S�"OZ��N�e���5�va�Ivl!�dV5��@��� 6�bA���<!�dK�XmD�� ��[N�,ru�ߟ !��G.u��ʷ���a�p�ˎ�*!�$Q�8�ZK�d�h���F��1"O��XD@ l�:��P0���)E"OX�Br�]�f�^���@�~ H(��"Od��o��(��smN�s"O�=2RB_�pʾ̈RΏ"QFڨ��"O(���Ǧ^T.���c��_樘`"O�\S��[�+k�D�0�B�PSt��#"O:L(Ҥ�K^d�z�g�\z��s"O@�tH�V_
�qD���9WؕpA"O�}sr���f�B�\PҍZ�"O<-��X8�$��G�8�.���"O�)#7�ғ|+Ar�%J�Y�p�"Oּ"���-��jZ�u���"O�@��eT�l���Q�)�#�=!�"OH!�d,����I�M�cp5��"O&@�Ť����9��3G�F=@�"O^���`�n`��{6 Ʒ<xn��"O���r.�/5ĩ�&6�� �S"O��4��dP w�� n����3"OD}�ag�[U��ҷ.]�(���ir"O��	3�@�0&$쓒��X7"4�"O� I��ء.��q	vlThB�1�"O����_/��#(:�i2"OB��q
ɢf��D����}nb�Pc"O�(ڇ�#e��}`Ҡؼ4Zڵ:�"O&���k.4^���PO�u{Q"OX��.s�a�T����		C�AK�<Ŋ�;����_\:�5�d�K�<�7��n��)ǊR�H�(�B��Q�<�M� bfŹu�Q�Cm�Ty���s�<�&	+!P��d�@b81��ər�<��LH�0i��js�˘4m�YjW�C�<� :�s-rXEa5e�?�f���"O `0ǆ D�����qH앰�"O  
��9����0��\JJ�J"OΠ�&i��`\�9���$i��l"P"O^�
�$� h���7�"O2��aȭ[�`Q��^/#�~�x�"O���7�3,]�̃��t�P�`�"O������8���ԯj�����"OJŚ�bL7������(@ʕ��"OLY�qf�/-���U�!8MH!32"OL�뢏ɲKg���!$S�;����V"Oz`P���'�U�7�y���"O�H�dFEm�b\�g�� k�p�"O�`` ���m��9Y4��[���11"OV�iQԒ{��`s����D8�"O$��k�v����E����q"O4035��T�r�Q�D�5HF�y�"O0���V<oE��(�˝���"O�(�s���^��Մ�=�ht(�"O�|�qm�!.��E�檐�b��t��"O��Bc[�&A�D�1�#?���"O��´m�1e*�A�'[8w�NU8p"O�]�"@D�hP^p�f��P�,E�F"O�$�֫.�2��֏-���r�"O�a������X󮆩^�.���"O:��m�w�9в�Q=+�|!C7"Ob�r$e��f�Q-�N�r�Q"O�-R�̭t-sFX�d��u
#"O4 ӣ�τC��8BP�P���"O����M�)9�Dd{>Qr"O�`� �3���fĕ2q+��@"O�%*q6�1����0�"O�Q���Km�ő��D�	0���"O�0��
ӐU�4qG.7vd��"O\��nI,2�����?�^�Ia"OL��6�ڨh��摜-�=�S"O�6��?�$��EN�	r$Ð"OxH�Ʈ��z\�kT"�4}�ܔ#�"O����a�H�ٶc�F�90"O�L ��J�h�q���?����!"O�(Yq�1Cю(r�$��h)b"Ovi�Ə˕G!f��j	��d�a�"O���I3���G�@��A�"O:bC�+/z�#F��9_��M�S"O 8:$#����QР��woB�@"O"I���իt9�,�N	&4z죒"OV�sB-E-oF�@��B'j$��37"O�Ib���c�l�3�E��w!,��"OZl����Z��	
"Κ�X�� �6"O�q�BL�~1����/H���@"O�4���H��=s0͖�d�J�0"O����	^Ď�s����.���"O(��j�I)��&�._�،s�"O�$X%�ީ:MNm���%j�~Ő�"O��V`�'XY���b�ΨH𠃃"O�ȇ�&*�XmS$�5,��"O ��P P'\Y�\�$��Xll��'� t���'SN��F�J�i��t0Љ�
��qד�u�eO�"����y���Cf�Vbb]�P�>[!�D�>GҐub�kM�(bN�3�E�_��'�N�1�M�7#��q �r@�����>�x�2���C�	8L�0������%	p��,��n�����{�
˓��D9��L��2��->�����bU9V��t!��0���d�� �z\����t���%��1�	�4��O!��I�I	~؞� ���&G�vXtqr��<\��2�'}�Hb���=@o�q�G��'b����n�zESѩ�c�X��eM6�y�A^L��iu�l5�)�K%���lXj�Q ��.
� jăٳ�(�N��݉��T�#� ,�¤�4"Of�p��̶'��8��w_���n�(G��my�F�#yP�x�]�l1�1OVMS��![1��:R曨؎$���'�VLQ��cǢ�`�
��10�C���0(�l2r$
)6/��)�T�az���&/4�3䞮Vfʉ�A�	��O,�JԈް;:Z�+#f�|���R>{ CF���9ˊh�E�Ĭqu�B�	�&�x�y�E(ҬA��!)���- TI�E
P�q@ê^��dӊ��F G8`b��J�v`F�P���!��21���;U��E"c.�.-�M#�=a,�QkOrfr�PԚ��d	 z��	:��'&���$�w�rh :v�(��M��>��	�Eݎ�@I�"|��ejd��8  �q[��'h$��e^<�AK��$�>M�Óls�آ�J�E^�!K�aC��Y[�)�.\ )�M�o����#�M�<)G�R�}��1ah >b.�y3C�M~bZ�x1G�
�2�.$�$!�'^���(vI�7� ����W�̵�ȓN��a��I�-9�J����C�Wg�H���ݐ��>����O�u��aB�=Ȍe�e�i!�`B"O$��`�1)�"� e�ҷE1hd�Ʒi�:"�F$U �P�
�9�$"r��6Y\A͜�&t̬��+a蠘�Ԍ���yrHG�k�d�����W�F]�U����y��g�ȥ{E�=قT�f�.��'�D���C�F�"~�"�=��M��	n��@�3n�B�<��KmR�a�҃@V��#�W�<Q�U�Ԟ|�GX����R4q���pÓ%�z5�3i��XT!��AՐ Vǒ�ܡ�oL)}�RY!"�a~R�@�����[�6���f�ݩ�yB�]�S�~�H��$\x&l4�y��ɡ�ʈ˰I,X|$���y���U�b����i,��q����y�,�?l�nL ����6T�@�ޠ�yPs^0�(��U ,���y��'A�I���H<B���P�ώ��y�A�X"�`�cY	z{�g�
<�y�G�"Wg\Dx��7t�"���/��y"!�4z��$�n4��9�(F�y� �h ��4 ̄l�
e�R�߻�yRϙ3��j�'ϻi�rJ��y��?3<|FiҮn>�U�P��1�y¥�4�"��6m$9�
������yr��?&��QIŢ]6crrt���T��y�&ʼzĚ<F��"��=�Pb�4�y2j�1sԱ�׺P�կ�4)
�'�@]�v��1��-��Eϖ)4����'S���hX0�L��fK-c$�:�'�l�@��f"��D�%N$ ��'p̉�O�?RLT9�U 2��yA�'�+cN (�`�t�F;0��p�
�'�v�X��=j��hC��R.5�����'J��Qю��dE2�z�L^�;��M)�'o�	��L�=rt���I�$�^(Z�'��!j�Ϸ^*(�� ,H)VE�'�VH��ݮ����q��y:����'��Q򋞷[�m2�fB�r�.3�'c(,Q��Q���;��� �n%��'�F�����f��Qz��Lʶ�k�' &Ы��8�2ё6蒣qߎI�'!�-+u,K5��Щ��Y`��0�'Pt�)���e�4���9N Ti��',&pY5��/���W@��@[r���'���'Y��6�P�l���'�I��-�"N�x�!!F����
��� j�Gܠr|���F�	1lP�Ц"O^RD	�d�UY���u
����"O��P�Ë�#JZ���ɻ-���6"O�ӳ@�\(e��"$�A�q"O�ؒ��Ƨ>_���������Q"O*�S�Z�V�P��@�1`rF��2"O��k����󬑙hvը'�;i!��	���-G�{���W��8~!�� �pP� A.�:~��8��-9`!�D'?'�$11�?q�*pk�J]�nI!�D�.hBJ��r�M0�T=;��W��!��%6���&�V�C*dbQm�3�!�E64K:u��c�8=`��#�Ȟ�!�D�=t=���6U i�N��2����.2��y��R�f|�6�O�y���dU���kX��ָ(�n�=�y� ���O�4[m&��PG�5�yF�4A*Νٕ͈�(&�� ,�y9���I�*�#O�j;�hÇ�y¦�1��a�AHԌ�Уϛ��O�Y7Kb�欙���]��HbѾi5M��m�E1�
�3
͊�X�'�Ԩ��;�)s�Ӆ*oL��'���c�Ͳ,�� ��-}(���'�z��'F�_�*<�2��%�A��'��|ZW��Z��偱CC�[pE��'o���Qň9�x�� '��'�<�
��)tz� P��ˆab	�'Rr��Ǆ�,'�+6-��J�B=��' ����.uE��8v�<<�!Q
�'�R��PkɕU+d��5K�-�~�
�'�l����R�|��e�C3J8S�'!*�c��<�B �-k�j8"	�'Z�Q��
J��VBB;n��x��'������y��d��L=O��x�'�v�q��
 GF�zv�B@P�1@�'h��s��J��N|9�������'v4�PC�n����~A�!��'?��6��u�RQ����}��Q��'�J��tj�Q���o�&���'5�xaF�5b�\(��W���X �'�xu�!��U�B9+c��!<�	�'�~�p鋑{�\$�A킎���ʓ�~� �˃2jՀ0&KR���ȓp�	��6,����E�� ��G�L��� �!i������ȓ{���.L{a#�o�P`�ȓ!G�ja	!xNk�O6j��@� �b��B�`�ڄ������=(��u��)��z'��v����)4:�0��ϑqS����=�ȓj�(uy�c�%�Tm��='P��9�f4�#�U�n>@)��\��vY�ȓoOڴҤ�<ȴ�P�
2R��ȓ$W���	�3]洼(G��]*l�ȓP�X�J�AJ��`Ո�DYFA��}�lȣ�B��j�8��Q�8����ȓ8�p{�N�>0��˕ PA�`���R�\I�%M_�/�jh;�,���}�ȓe���b��OB��mb�mSbOb`�ȓU*T�uȅ�g�Ș�2�kA\�ȓ	6� w*�$H�V�����s��8�ȓV;F��P�hRtax�Ǔ*��5�ȓ�Ve��)�M�E�P�4	�����Z���hǷB�5#ײz�<��S�? v��3�B�ɁA'�d�q"O�@�3
A)/��"!S;JI���r"O�iȆ���/R �aMΤ7���$"O:��,�(p�* F=b��H!�"OP�
pB�جx2%�T�h�.��#"O��؃�F4y^��I����&n(��b"O:��4'��*/�J'��.zp�`�"O�8������#ł+ .d�5"O|����N��i����2�Q0�"O��AN�.r�>x���>���"O�(����|�E�'�q�"O:|�b��Bu�H�1΁%�ޥ�U"O�%�#Y~z\jvL�>ڶ�JV"O"��e� W�~�T+E�@��f"OF]�VJi�U*��	,$����"O�}w���IE
���T��`t"O����<�$!I�,�q��"OD��Γ)O�tq�E�^0�i�"O�5��$��4[��:�Ē�F��PS�"O�A
�fA7�R�1wn��t�� A"O܈d�&�%�DQ�ģ�"O��:�)��L?��q` W�2E0�u"O������h)�Yp�N/l%Ta�"OjBF��+
V Bb�je�b"O2M2�ۼG�<����^0�5�"O0M���35��1�É3zp�h"O�����."0�胠Ə2@|a"O��p��߂xH�e���WRX'"O��h��D&r����u�ǯN�B4"O�d��Gɜ\��1��Kn�6�3"O0�@Dm�(r5^�*2�Rz]�%�A"O]z�N	�8�t�g�kW:pQ"OT4��Ǐ=�f ����	J���"O�= � �n��l#�b��V�t�7��h��D_����`E@!6rAb��@)ny!�䊷9�	i�C�
	�Qc#Z��!�$�5c�AZ���k����Q� i�!��5�u�"�W67�.h	ԋ�%�!�Dʪ\q�13�ᕮ��=
�
D4xG!�כY��ɉ��L���� ��;tW!�$�JP�hA�DG�~�i�R�� 0!��1cm6�"7��u}JY8M8Nr!�d�g&a"�*CRRYH�@�)�!��-��JWc��\;�)jvJ�")�!�$�)�|gI��A�y����!�$]Xn�0��_
4�vfo!�䗯,bZ�j6,�?a�F��^�T�!��V3��5�R�A����s���4D�!�C�mf( �@;���X���1OB!�ڞ`u����II6��ń�94!��ݯ�vC�⓺C1>�@�m̤1!�DE�^�J8��!��J/`u	�m�(b�!�0` *���Ė <Y(�͏�A�!��* p����P.4�,*��[z!�
�"L,hڴ��N�4"����.G!���!�� �Y4	^�IEJ��P>!�Ȫqm�:��7B��B�oݣrN!�	-� )�����]����o;!��N��x��T'*�Hp 0�K_;!���5M;n��k��ȸ��KƯ
	!�$�<��}H��&r�B��k�)\!��Š��FA�T`���e�!�^��\A� $6�蜣��O�>�!�U�.��do�7ڀA���V�DF!�� \Y� #�:d����q�N��e"Oڡ3d�æu)*�G7�
T)�"Oxp+�.�<�`�6���>��=r"O���@ Й`��]��@9]{|i�"O���۟��ժ�V-m&�!�"O�XȢ����Dr��( fܰ�&"OH��vc��C����bMF�y�E�"O�y� ���i;�=p\�{J�a�"Or� �cڣ"X������?:<c'"O����{�l�s,�F2�x�b"OV� /	� :��!���&>��L�f"Oܭ���%�u�ː:h�@e�c"Oڥ��`�1�a�#�ؘ/�H�"O���,q��y����%ea���"O.4�#UrK|� �J ����%"O���3h��VP��h��V�n���!�"O|)1�\���|�ӫD�?���"O�`�b�q���f�V�:E �""O�]��E�(Q�Tj���%`h�"O����!y�`�+|�r"O�dCq ц?K:�J�$>��lQ�"O�R�-ƖK\����t�,)$*O<h1��\�j�:DE��ex"�{	�'�{�lO"	� �#�a���'��٩�G!6ot��A2�5��'�r]� O�A�x�1�9 �'���Kһ*Jhad�Y�\>X�*�'��b`��L��=Hs%]�%�V4��'��x"�]�%�
ăR�%r*�-;�'�p#��2W��� RLg.���
�'��gN	"~|1a�׭Yr.(��'�􌩥 ў4���(S'T6���'10X`�C�	��񪶤֜S�B�K�'jڴIF��
WE����AB!%�X��'���$ڂ��Y�H�z1��'��}���M  rf]r'�JE�^-��' N�� �4lL��0&*/-,���'���L�]qDh;�͐�\��'�T��,�<rЗ��-*�����'zH  !t86����&K�!��'��qЅ4$���I7E4�i�'^��i�bK�&H J�Ϙ	Qh,�'+�I˅m��1O��
r��; 2n�P�'�ҽsTf����ؒٹI�� S
�'���`E�!�l��/ےB+
�'��F���a Pc�4w2��	�'Ӥ��@������GO��].���'	,�:�`CH�� � 
��0dq�'؍ʡ+�6"�&�PCn�,q�EQ�'[�-20�\�6C~A�E
l���q�'6,���@2�AQʖ2�|���'���#/��f�R'�b���+�'��zbIˇ2�f��E�D�]�ԋ�'<��Y�A��C%��$7lT��'�����\�j[�U�TB�2@��'��)(���2�����E�}�0} �'�P�����'�0Q1ġ�.L�C
�'}.�����#���S�öP����	�'���+djL�s(9���������'L*ܙs�_s�b��e��2!��' � �1�@O�!qAOJ�
���'8�=�0"џ_���"b@�O�JB�M@�Q�F-�>͠gC�t� B�I�S�8)Z��5�]��,csZC�)� ~�8gM�1ڂ+�Ɗ�7��PCD"O���e��UFQ`��Md�2"O\hg	O�>�(=p�f��	��Yt"ON�cB��[sl���D��9��)K�"O�2��S!|��
D%�����"Or��bE.V�(s��ʿ�eX�"O�āRD�	"� ���t\^!�"OD�[���'$���E�;=����"OB a�R�� d�<���_�yB�B3F�x�Y3�\�&O�u ��y2�M���U���53���*��y"BD�6����Zﲥ)�ʪ�y'�)H��2���L�F%�y�`ܹn6�dqr��G�H�����:�y"�!�AzS �II���5Ɉ�y����F�h�@"m�E:�)��yIΉ�Fy�`a�-�� �C���yb$�7d���)-{P����Ђ�y�o
�u����$�A�i;��`�cy��Ec����bۊ ~ ۶m]'J���ȓ(�r$U�^- T��Ц&U���ȓj&���b"V�|��H J��d��q�ȓYEqЅ��=4�{�B�ì@���DC��޽|x(i���\j@	��[��X� @�?   X   Ĵ���	��Z��wI�*ʜ�cd�<��k٥���qe�H�4m��_;:<u�i��6���K��=�3g��2�R�9AfN/>��m���M���i�����P�O̚�+������ch�i �o	��M����O���4]�B|S&j��.zU�VnR�q_0��'&Z�Q�����݁-O�p6*�p�6h .O�)�e�Α�Zm���
9HfE��$$�4��4M��!���OZ��E�&�s��i��L�6䨰*�3�R4��GT�+��1�nC�
��ɯAhl��j�th�'�����)�~�f3{��T�u�0Pd����k��~�O�PC��J�yb���GBxx�<ID��%��l¤ �P`���<�%� '��"<���E���˖�f��-�!�U�{P�LɅ�I�)F�ɊE�:�q02�*��En@: ш�'���Gx2j�Hܓs�A��&�.+��{v��4B܁oZ��0���8F�޽�(�(W�б��	+2��%�	�L���f���cq��-Y(ȑz���5��d"q"�<�@
*k�⟬
SB�#y���ї-vhV5�6�0��ܠ��	���k�7<a��n��#�|<K��ܘ'|�Dx��Cp��:-"I�����y�j�'�Hm�f��"u���YT�xB"��P��g))��9�'��L�Y'�O�h�'�NxD�̜P��'���fDM����ݾ_Y2���&ͨJU��3c�$��ę:R �Q��D��j`ԭ�M<�����8�L�q��:�p����J}bh�s�'��Ex��a���0�zpH�Wo���y�@4. d  ��D���<��С�'��(=+��:D�X��F!��,��(ə�DJ*7D�İ�����²BSw�LЇ#D�쓱C���^'!WCF��$� D��P DP9�=�ԅm���s��?D�0�4�,m��S�Nl�~���;D����\,Z��:�=(v����:D�,q嫏	m�� aMF!�r��-D�0�R#�cv u�b��8rԂ���)'D�p�J��e� %*�-�5C�D����%lO���AmB� �T��[�6�ˢ�-D�t�d� D@6��D�e�8EO D�x�@D6r��!�i�<P�Q��#�O������$�&��3����ik�	�ȓ(T�{�jB����tj�-�^��H���B��l0� 0Ɓ�+��u��S�? ����NQ�:q�=�&"C�J��Aq��'����    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �P   b
  V  �  p   �(  �1  �7   >  zD  �J  �P  YW  �]  �c  'j  jp  �v  �|  ƃ   `� u�	����Zv)C�'ll\�0"Ez+⟈mڛX<�	%6��D������&�:)�����B�<5�eO�N`���.��-f�A!)ߓzY��;0ʈS�'"�Ÿ�'x�zikR�1툘��&L�`=�̘c�7<򬃂*�a^4j!��cx������������3R!�0��D�꼑�n��
,�BO�4�����%R7�S��
�ٴFw�(����?���?1�jT6�ZHU1y�*����rn��?��E.-;�Z���ɰL�d�S�P���%��@��K�i�x�مώ�$���Iٟ��	ޟ��Iݟ���k���n��͓thhY�b�1�!��0O�D%����<D"�l�b �T�l\�ڷ
S}��ID?AU�[�K��Bov	��
/+�u��#�&]j�H��ן��	�,�������O��N�4c�F��5�.'�p0����>"�u�f�o�8�M�Ӳie҇u��m��M��iyA��Ol�@#7F�:x�=�G͋�c��"=ɤ炧�����C`قM������H���{#@W�=���T�L�|xh��!~Ӵ�n��M�'�R�&�-'<�"���u2h�(PA"�l!��n�j-8��Q��卂�HQ��KF�H
 ݴ-��fr�(�ّ@��{��8R�C�;�D%��T8����`�lZ�M�c�i
�����ć\x��y"�%*���@ Jém�f	����r�qa枽a(���ǢY�Dq@�wӜ�oZ��M��ᒬ &�<@���B�=(g�׶ �,����
BA��d�A�>a�6�i��d����h����"��LE�d��'�OXօE�_�MqC�4�����b�OX㟜�	�d�D�M�ΟTA0(V�Du�9j�N�2i.��I��'�__�� ���;.69"S���c��
�@Q�s � �U���'<�C����7�!2rGV6!��1r�7=��]I0�Ӵ-�U�@ME �|4Z��0�����P���E>����'�˓p�	O�5T��u
S
A� V}�	ݟ�Ib�Ş�y�剚vzj�&�>z숐�ƈ���?�c�i��i��D�R��q��xBLapw��D�$Pj�D�����oAD�*�j_�n�0 �cڱ�yRKɉe�n�
!�D�h	`a�	��y��έA�PY{����g�La[u!�(�y�,�d�h"�L�ZT`xQr���y"lE�5eJՓ�$MX�ey�)_�y�#�}��(v��H�4p���?!��w������c�H\9I�r!�'oxF��4a;D���`N���aT�
����9D�(�A�-l�|u�6D��l�����8D��i@lӭƅT�r���bV��nRC�IE��HQ��<������`��"O�]�'Ƃ8��!�p�X�pX�Z�]�,Aqc<�O��T��:i���Y�F�6 zq`�"O���nT8|���IF�;X0����"O$�*P�H>9��% 6�0&5�XPa"O�8�`[�[<^���!��p7"ON��QbɲS��DH��	0��S�'��i��dy�>�J�9�H�h�[��G�0 ����UyR�'��'G�#F��F���S�	0�7mDw���$��#�B��ь�?[����DG;�rԸ'Qs�i#f�h�f}0ԋ��/n*P���ϒ���w��y�Q���f�OD(m�+�M3��$�x��	�h����3ǖ�q&l��,O��+�)�'E�ha�P�M����J�>�"q��ɘ�?Y��*�h�%�^���s��⟼%��s�j�b>���[��ƭq�`h�nα`�;�H�w�<��aȊ�6y*��רT��C�a�|�<��I�/s�(�a	��DMz7�t�<A���#?t���R�\�f�!��n�<���&sJju4K�*��Y93�d�<���W"�:*�p��ͫR��Lm�Y�	lM��ܟH�	ßT�'`��
f��"x�b�ѳ�Y8�L\��4Vy.)�T�j��	�!�9'�ʧ�R�yR�G?S��0cV'׶G-��s ��Oe�T֪F�U ��z�ğ='����Ćҥ0Rh��P�ѤMNUk���t�;Z:P�ش	��	�Z���?��O��d�O��X2��S��!VB�%;�t��*<O���?�!A�%q��<҇	�4D����Iy�|Ӟ�mZh�i>��Sfy�MB�/��b	Y���%8th �Lt��Bl�"�$�O��D�<�L~RW'�$����4H�C ����-'OL���)�}��0�$̱�0=yV�U�.mzt3��X�^V�����µp�0���D�.3PD����Uf���`"��<�(Y"p��Q<�aאh�$���͖'�R�'7��'��?�I@Ç�)��蹕��'F}jْc>D�lI�O�{XHK�f^�;��x�K=�����9�	^y�/�7��O^�d�"G�v	���ϬF��9��)̚A���d�O�sM�O��dp>�H�O�c�� $t)p�.I�vOA.+�D���'��0*���
c82)Z''��r�0���Vax��Ѻ�?A�|�bQI/D�k&�J�ufF���B��y��ߥ{����kiy�y2���?��'��%nA�a�Y����8��r�6�Đ.X1(�o��\��x�D`��#��F�;$��@ ̯=n��qA����'D@�P`��@�b/�%��T>��O=�x���Jm���]��q��O����!B$����-�;/�t�}�@�A>^����Q���a��a�A~2��?��i�$"}��'}�Jd��*"p�A�n�0�Xk�'	8ۅ�^����a8BV�����E�O��ܡWM��H�0)R憼q��Ƀ�i���'`�Ϣ(I�M���'�R�'9#��
D�$�
�G���"!�ˎ=�ĩ�V�0�ɐX$�Z�	�G�� PV̝`��ăZ�� �!O�DH$ݐ�O�K�	 %1�1O�D�˝=X��	����0���'��7��O����O(b>˓�?i��.X����-�yT%K&��<��'�O�����G{��n��6����0�� lZ��M�M>as�O'�2.O��c���U�*Lp�C]%-<�x5d�6%�m�r�O��D�O���ʺ����?�O�J���->Wk(�jk�(@sDϋ-O�\xrt�L�Պ��%�'���+��H��2�3t��<jG��!D��XV��^ w�i��'_P�(#g�IK(9�1���Xˠ؉���?Q�i��6M6��!��OHa��K��:H!�M�;�M�
�'{,�mG-_ͺ�Ѳ�6��YSO>)[��'@��0
t����p��!Ĥq�|�T�+�"���}y��'Y�'��͡��ѱ~������!|/�6M��v_Xh�ڲeffK??M��𤈹5�N�0!��0=8I �i�����V����8�.�a����Q�H%�Q��h���Op�D)?A� ̜/Sب{Z�������oN�,�	ܟ���M�S�O��\c���z��E逎�t���'	�&#2:%�م��,30!���?�)OT��d��Ħ1&?��O�� ܱ!���P̍�E�qPr��;��'�z$ȷ�5��,�A�P������4\���"A㛑��hB���Y��
|�G�/|���e	g]h�2�1�+� Mz��X!,?��
c��1���A[~X�	���D��'��MK��O$JR�
�b�L�z�"OV����F�Q��H6I�l�Z��S�	��h�܍�#��)m�y��j�˄����>�)O��� ��d���O��d�<��0I��s�[�L�r��.\ `	�,�Gʓ# h��Θ5'�=
�����Z�>\*`��(� L
Aթv�-����>6x�6-D,�K��1�~U�=�<��"��`6�`�#U�Nh`��	F~Z�
���?I��D#Қ�b���^F0ԁ���=ThC�I���p2nC 0j%�"ď���r�����D��1�#H1w��|�E��;�
=�#��O��d�O8���<�|"􁃥r� ��o� ͫ� �
�jP�g�*g-&���˟�Jf�72O��E��9�~0Õ��1��F	c�0�ĔBY�����3���&�O��"J��be �D�xa0Yb!�D/52�'{ў�Ex"�^HPApf$E"!�Ba�G���yB-�EfT�E�7�2�pMS��H{�IU��~(�H�'�  %��1W`	�([�[I|x��V!~��p‴r�����.
 $�ȓmg���u :d�])�j�N�X�ȓG�R��F�<	$<	��#@���|��䨰��@l�(�f�T�;�U�ȓD�"�󔣎�tJ��>?
�F{��N���.d[cޣ���f"Y#���G"O��SÆ3T!R� ���J�0��"O����ze< {�[A�ݡ"O������B��7g�&
@E��"O `C��0-��%M���Y�"O�8�F M�O������6��A�1�'�,�����e�j`I���*������7x�A��)��9���!36���0Eg� �ȓR$��S�ױGM�8Xf�ݗ!鴀��w�r$e�
���*[��#�1D�x3�.٢M�N�����~�Xp�f/*D�(�c��43��X��ܣ>���Ǧ<၌u8�|ٲʂE��Л�jZ�=MXe�Э$D�� vQ 'D�!	�SE�!T�6uH@"O`��D,�m����æf�̕�$"O����%l@~͛�'�%+��I�s"OY1��H�dT�iܴC
���2�'�Li�'C  �fZ)ޮ})4�!{Jޔ@�'aJ(���߾r�B=�C�YRl��'Z�E���� �T4���4@x<��'[�]�d�ɚY����d��7����'����	� $�W�/�49)�'�,)�n~���u��4$�x�B���
�R�Q?
c����\Seь`,��+pD3D�hB���8y�h�*r��v�^���/2D�0��&��\=L��JK>p2j ���,D�K���*^�-`�`��e�P��6D�c1΂z�j�j����O��ᓓ�5D�$C@�e\�x!g ���xC��O��1�)�{P�H	�j)�j����֡c�M�'�t�a�`�1)�d�p��'�ڹD��\g�L@Pf����{�'� �R��|ļS���=`���
�'��y��$S�5��%�qi�=̼��	�'���cr�E��H�aѶE�Ze)O�i��'���X�����-�pd@�'����.������P3 �&]��'|=�(R����7#��{����
�'ʲH(�Ėf���󠙆x���'q�L��K5R�	�c�w9�� ��z� Vi ��wtRUQ�ؠUo���f{�;�؍A���Ҥta� �ȓkΚL���Z+&�2)�v�C7p�D�ȓ8���ٷ��1_J9�h�G�Ԩ��;�&ԩ�b5K�X�Ȗ��5P����5�\�ߤ��b�^�/7D	G{ң҃��� ģ��+l�Z�$[�t���"O|Db�L�i�:�0V��
s�M	�"O�e����
�J��F�*�( �"OXX���ʘ%���T��� ���"O����( ^���c�aN �f�;"O0\#�cܨ� ���@� m���i��'�8p1����x䶜3��]a~a�Ȑ�7�H��;5�Q�G����yvE�. �ȓY2�Q0���/��8�W9LE�� ���q�+
�MiC)W����ȓ6�����!�N��@�hh(�ȓq$d��ؿI�]��M�_Q$�' ؀��G�I��#1�,,�Kȉ��ȓB(8�C �"X��Ò�
�,b�͆�(�z�RBē$b�C�
�o�m��	���xr��>f�h ��!["iK��ȓ}�Xi!���xvH�e5 ��%��Ɋ_r�I6D��
�ki�̲&f]+V VB�I6Dj������gۘ��Ӊ
A�BB��?p�i9�!Ю/V�Yq�P'&phB�	�5��j��X6����&B[0B�	62)6�I�K��"i�ͅ'P^�C䉬t|~"��޾y,�0� Ǆ{��=����`�O�PPjǋ�_�����/��
� ��'=�P�eڰB�w�]�~�^���'xR�LX�zME ����z\�(9�'���Y� �-S>@Y⯖�ue�И�'}�a��m;j,MY�Nހi��<j�'d�i���pn�y�k��r�Ѫ�9��Fx���ъRX�uh��\8��a�i�{s�B�I�9r��+p�
!�����(W��*B�)� x����B�e%l4��R����"O"Ā�e�k�j�X$.޹($"O�x3TAX?A�*V\$������W�<釮�0 �>zuD�7'S�����Oy�
��p>q�"�Nu\D�����ܭ�b�N�<���  �c �k����F%�J�<�%��>b��×�@=}�:��'�M�<�� YgK"y33�ӯV�n��1jOs�<ك`�R�԰gj�*z�`�'RCx��i�ୟ���ן[��u��j��&���V/!D�����Y�
�:$�6�W�A9��!E�<D�4����7W�.����z�V�b6D��@�it����ӪAuL�@�5D���I[�}�`���V���c��1D��(�bޚn��)(�ᐲZ��ut $�o��UG�t	y��!�q�ҿF`��C ��7�y�B"[����肱C���
�V��yK�C���m�4-䘠$E"�y�.�zg�Y���0#Ą�d��*�y2.�$]�`h�A��y�FӀ�y�	�7 ���ĕ������?���PF���� 0�t!��@���b�5�z2g�,D�l�A@��"�܀��m\;~j���-D�X�D�_��]�t�Ͽxx�E)D��ZTCQ:ITz,Z@ɏL0����*D��D�m�Ҝ�-&	�(��E4D�@`�(N>s]P�b�ˆ�la��<��e�K8�̉�f�,P�Jݛ���{�IA�'D� ���Q/{fH�S�τ�$�T5IӠ$D��	T�q�l�R��U�R9�Vn!D���G��MA`�m���ب)�i:D��!��'e�PqaE�P:Oi����6�O�V�O�	&�� ��P�C�H�<o����"O1VBD*:;���#�C�5��Ȑ"O>5�ƏZ�2Wd����^	~-�x:"OJ���h�:���B�Nŵh�90�"O���#g�~���#mݧI�K�"OF b��Q�*���ˀ�d�x����8n&�~"$([&�H��@\�*X�!��F�< �4���r����\��{�<Y�
0c�@��	�4����2ɐN�<�p�V#3��I�l�iT��AcXK�<a�H�_H�� 2BV�fJ�s&�V|�<�t��H�*�h2�ED$u�š��|sE-�S�O �9�7c��z�&�T�J1��U2�"O~�D�ؽZ����Ui���"�"OL�B���L�|��tJ�a{0��"O�l���4Du�o��hb~�h�"O�k&�ST��йRd��1�*�	�"O�4��$D�( &(�WEѵu>ư�]�|cW�!�O�9����3����	
s2͑�"O�\��K�~��qvC>/�P!+e"O�L��'NBw�� +o���"O^hy!@P)9�i3�F+7/�xw"O�;�!�]&��r�^�"��A�c�'x �9�'H�� �Ų8�"��wL��40\�"
�'bT�)��&�#���3̈!�	�'�V)Qt"B�����M��Y�(��'�L�f�LW^-�C�M@�J�'{�t"IܺA1V|�&�}�}�'�f9�'!�78�PC��v��ē����&1Q?ݠ���4�q��`I�%�d�4#D���7�޳$��(����-"13`F;D��Ё��!L�Z�ɉ�~�=�;D�� �$��tm������-t�m��"O����&T0^�d	�FC��n�	�"O*%�F+X��H�ao�U��	pT�'��Iy�����ȳ� �Q�-���=Q�h��ȓK��!� ��>"5:l�6X2�)��[��Y[�^�G��й��]�م�L�� i˸gJ\)5�ִb�r��ȓu0��F�}HP�Q�ߧY�bi�ȓjW��ҵ�hc�K�)�"?�:d�'�^p��'�,ax�CW*`� Вp��!M8Q��n���0v�D*�}�D��n�D�ȓ:��`C�Eѐ ܅�5a�Kl���ȓ�ze�Gџ2��� ��3_bX�ȓ#�ؕ �Mw�FEA!��y��q��IGv�	�x��i�jÜX�R�Z��P�"�B�I�z_�9i��L�
-���o�:d�B䉮z���x5�� _�����JS�B�	�3�` j�$Oڶ��D�ř@T�C�	A[�l���xr�Ax�m�O'�C䉞h#h�a2	�s�đ�O'|.��=�Q�w�O�������V������0^�N�C�'�ReڕjI�8@7��W�^ur�' �����I�.���d��?~n�P�'����c��84���I�c�>0-t�c�'�h�ل�J�9גu��dV�"bA	�'H�m� �kL��#%��� �S��pGx��)K->��,���ޕIE�� �W�C䉅��t�pj�H42k�63~C�	9�6�� N_�b�4L��C�7	�B�'���" (@�_��"��[�y�B�	�s"fM`���(�-���ڋuTxB�I�{F�
��:=5��rScձ{����_�DUyrOF�c��]�/]N�(c�C��Fe�<%�˓�?q���?i�F
'BX�"���UY~�h@�i��i�.\px�e�`c���Ꚃz���h���57On43�� �J��n��=Jp���Jk��8������g�CV�'��P����?�����6k��x��U!-�:�ӦCԉ��$.�O(�Q�I*���sE�h4��k��'�@ʓ{�F�;�����_�`�Nh�'�0	���x�D�<y/�X�d�O aYOS�$b=I�+ڒ) �Z#��Ou2a���|�h���k�l��O�E�79"D`�%Q����'dp��c�O�Q?R���&�2i�F�ƈ�(�صQ�e Dx��MJ�'��A�E6O\�@�'�Ҝ�����|�:��M�'}�l�SF@>.��ȓ,L�m��.X)���b�� ^<�PG{��4�'M,	x�e�	x4�$Gܔ5y\�Z���D��,��d�O��d�OV�S2s�%�����
���
6hʹ\�hٴH�(L�F�;b�F��͟���s�їm/��@F
2Zx�yA��$	���lZ�9���8�Gϔ�e�Os�U�=G��8�� ��E`n��%�g~bK�'�?����hOX�I=c��`W!]�V`k5��3=�BC�əR�"aʵ�F�"�d��S����'n�"=ͧ�?�*O��V��m<�[�����bܢ�ʜX����O��$�O��Şs2��3$L�8/x����(6���� ^������*\�-��iJaxZ�`h2!o�5<��S��H*D�:�MX&����Á��E�\{�4�^�F}�����?��M\�u6���L=$v�u@E�A��?���d#�m1~�t$W�3vv��iZ w>�E��&����b��5A�1�ɉ�}O<e�'�*7��O�|��)WY?��I�|Z���!(f�s�㊙bPȠ�4^���;�m����	⟔�bAA&�&)B���R<����|�%#o�q0n��`D�L�'���"@�9@�M�х�	{��-�������	����"X^">�������^�'��S���3}��ik�$�)r�L�'�a~2jЖ��	ĩ��]�i�5�_���>I�^�`�j�b����J���\�*Cb:?1dL]����x�OL8c��'��(@�:b�y�uB�+�8u�dLZ<Q�"GV,gNJp�3L_�i�fuZ���O�k�'.�p�B�~y�� BlB1~& �E�Ēt�䶀:#A����UasjZ4�0,(�� �'�z-y4O�IӁ�'����`�S�? >�CĆ.}�$Ղ"��0�"O"�
7��W������m�N�����ȟl��ǁ���5R�:��bG�
��t��~�����p���OD���O��)�O,H���M�[)����ƈ�D`F��٬���I�-^�8�	@P�g�'
�e�K6#�TMk��8:�h`�f�����)����匔���I&6un
��?D�d���M�^���}��I�	�G{�?O"��%��{��Պ�J@8r�!1�"O6L 6�;:���T��p�\M���'l$"=ͧ�?�-OF���R��ظ��TyT8�`o�N��� ��T2$�����O����n�d�O瓕y�x��,��H�h���?:�(�I�M�jƐ�P��k�Fe��ɉ!,�S"��aY�Y;�-G�DL��(	�in��GA.ݮ����hn��Ч#���j�f
$$b�ݚ�%�%J:��.ړ��O��kzn��"C��)�(0c�"OH��B�èk���Ӂ�L�0d�0b�S��Xش�?�+O���t��B��'�鏹��1i�
�:BF���45��F���'�R�G"9�`m[���q#�XAFi�O�)Φ��e�#�"Q:|���Kz��̠���2{�"tWlN�88�O�2(��&Ǜ]��%�����n�����d��R�s��)$?M�lD�'��Z���V����RK�<���0>Icn�o�^|j��ƻr�����Z@x�\(,OT��g��9�hD���"J��A�uX��	��Mc���O{����TM^�o�̤`Wc��X�����d-O�=���%���I�`� ��*]���?��4��>;�c>�)�Z9YP)��g�,BUQ�a;?Y4�OPQY2�>��y�-M�ն5ȷ�@�S���C7@&�>�����(�K����� }��!�)P&$d&�"�uڌ�2��E�
a�M���'�>��K����7S3�R�d�2Ǒ�I�~�'y��'��I8K�\a��r#W��v�� U�I���Bg�'�IO�4���0��
Kd�!q*�>���Cs囉��8����`�OR��OZ�j�>�i.��Z�E�	;���^/���/OT��B�>!��S/{�J\��%��1�|��$�-�~�����|�+KL��'$��Ґ+����C*\8.NĹX���	Y��)v�t���`�D铀spz\��)N,+��1g�ځ{i���G��~���9���?�	6����|"iq�nֱyp*TE"*l���R���?i�*K�R#���R膆\),�9WO�N�<�t��a!�l� ��*T*��-	Ǧ͕'_r�'Hb���'OZc��db�$i�̸�8: ��O6��O����O���<%>)C�Bܰp����xR|���!�d/�S�'x~�x�Wሶ!��ڧ� Cp�e�ȓj��̓���$��oDjcd�ȓ3dHq���M��DH�KT 1�<H�ȓxr,	����)���!��[2:M�ȓ[FZ�Tkܿ�y�E�GKO���xf�����'�V���Ъ|����ȓI�����.� N�\��Ɋ*�t���������CȦ鸲��'R4�M�ȓJ�i(�n�K����#��%\����/	tejFヮ{S�x�JͪI���'J��ccP~Rs�U�w�����n��16i��j��������Er@�?ٖhB�*ڊ9��Ӊ�~��jY�g��Hb,��2��U2�]Rʄ�4hY/���B^ I{��$O=@��U�M���sw�PK:db�oV����S:}���Q�L�5L(�@��h>��<�f���l)#D����Q�n�?T�lLX�*��~Nx��"�|�D��}^��C���p�D%���Ԕ�y2�X%(*�9��׵j,P���ǳ�yҢ��S�4(@T&r�@��ta�8�yb�'?S#��d�"t��kO��y�E��p�)a��`�L��ʐ�y�*?NN�B�F�-`��,�d��)�yR+_�AXY��G�%Eמ���� ��y"��!0����D��ʑhL��yr��?���e��7���K!!�:�y�Q�]�|q�_�2>.]JdH���y�n�>/{��òdٛ$}D��Ӌ� �yr$A�i���!cIKR,Q�􀖴�y��I4c$ti�_�C��S턯�y
� �ف�]+L��2ԦEÜ���"Oڐj��YK�)���7;���A"O�՛��cZh$KŃ�o���P#"O��x����;D�����& �>�ء"O̍ف�A��`Y�ǰQ��T"OZ$d`05fT�A)h֔dc�"O�����lq^10��ԓkHQ��"O�,��A�e�e{��2[OшU"O���E%�(@��ߜ`aPa�"O�Q$��<l��1@�A��a	D"Omc��Բ/��a0È)2Th"O�h 	�^ X��#��K��Q�"O��:�l�2Y���]��I�c"O�8���E��V�A�|�H�(p"O(T�P��26 ���!Wr�>d��"O��3�	
}�� �'�Z�
~��6"O��`GJf���X�IN�~��J�"O����E�IG~%�b�<|ňUj�"OjD��E�
6��[0%y��H)u"O^�p�B %b݂���$X0f4ڶ"O��fi��s$��x����رu"OCa-�b��Eͅ7����U"Of9)��[��
`�P���W��x�"Oj�r���8ceF��'@y���#`"O���W"�J�|��d�S�D�KF"Ov�0�'�n� %C�07�`��"Or����W.���ⅱt>�"Oh��R��?uf�l�P��$<���F"O橊e޾�&-sq�
����"O��x0��N��H����K�yD"O�U�e���T����&;��,�a"OF��j�$]D����Ι-�&��`"O�യ��a�
�r�]!_���#"Oj�
W�:6��,��l<u�4ibw"O�2�*Q�K��{zq�c"O�xZCN�O��%�'���#~B5;�"O�"BM�}��D��f�2Jv�!"O ��޻Aj P�rF�&	n ��t"O݈�0��Qk�+�&tk�I��"O�!
E�O��,R7wDA�"O�}3�b]�(�����Ý�}E*ѹ�"O��H���g
��b �6l\K1"O��:�f�clY�$
^�k���'"O���c-_�Z�� �h
����"O|�Gg�<SFuZ��%o46���"O�xiA�@-@5C��],V�j�"O@d�)O�A@2� Չ9&)�"O��f�V���Xc��7)�$�*t"O\����_9VV�Ԏ_�3��"O���	���P� �g��:�"O$Y �A�a�T�p��$����"OB�����#L�G��2~j�p��"O>	j�����i�ë٘f��av"O���v�%?���jv��</d|�+�"O\�iU�5B���"#��xJ�"O�l���1HMջR� l,�}"O���4-�2��V Z;q��;�"O���"���}#0��;G��ّ"OȰ`ਏ&SV�I4n���x�!�"O��bF��1�D��3�)j�P@ R"ON�v��9*r:q�$��,l��P@"O֕:�JEr�����	]�x��Q۳"O�A��9S��q�I�<�^�z�"O�\����)m������S�.���f"O� ��ĭʩ
F�x��HF�Z�:!p�"O&��Ț|'TP0fB��nb����"Oj|1ai����sϕ�@Y���"O���B#���b'(۸f�)�B"O�TІd�B"@�е`'H�<�"O��@`U�O�D�f���U��# "O<e��/���
b-ƿ|���"O���H	b��yRk��y҂�9"Oh]@�ʟ�6���iF�A�a'j	��"OphДm�el,�P&o�}N5��"O����.�*dU	���7���"OV�J�fԽ2[4=��iU'o�����"OX��-D���Ũ8Q���c"O����Ɯ&l���` (�q*�"OX�[4�˷2	E匪
�0݂�"Od��wR�y)�;��5'^t J�"Onܻ�.�&#��ũgEX�GFX���"O�)B7I�Y��%Ǒi;\��w"OZ%q���<�1QD�>����Q"O.�e�Нm'Ɯ-Ԁ<YQ�7�!��;)x��eǝ(c-�����ŉ�!�d�8�����;^%�A�e)I�!��]�-����EMV0[dŻU0�!��>'�f}`��@/S	��ub�@�!��4ۢ�q�&ґj֖M�B�J�!��3�
i�s��(�ze��Īd�!�d��\:��3�έ@�ꙩ7K�i�!�Ě�@z��a ᐥ\d�DÆ�˝f�!�D�\z���59g���@"^�h�!�����
�k@,��1�Z�	�!�dFB�ʤ ���'��;so!��a`1�#$Dbji��@�`�!��
<�y+�5�~ԋSb� �!�d@QX��*0.[�v�)�׍~�!�?x�����W� y�å�~�!�!�ly�J�7�H0�iFK!�$ҧaj���f��:��h!��~<!��hֶ �! ��7�=�-T1!��¹sۤ0%'�?.l��MI9Tz!�$@�>�ܠ����/qX &��l!�$F1|wZ8�6m5q:�aR���jV!��.���b4�G�$d<����+!��[<,��0@
�e�:����2!�D��"�B�it �O�Hr��4}!�ǧbv֡"D��$W~И�,� i!�a�2��a�6A���X+I+^2!�'d�BĚqQ�8NѰg�ʓ�!���C�@I�b��)&J�C0H|�!�dE((�c�����BT�%s]!�DȒŮ�@�G�n�� Rm��&�!�D���I�1G^*]�8L�`f!�$�?8�0qחָ��W6kM!�D��h�2Y���Y�0�0u����;�!�$.|�� aM+�A!n	�_'!�$H;#���E/$���"mF1m�!�DG3,u`6Ì .�����հF!��L1�b���V����dŇ$i�!�$�,1��Q����v�pm�T%Q9�!��lLM�� �T�v�I�!򤝢$�A: �Oݬ%�2C��R�!���#� �*P)Μ
ٖ$H�B��W�!�B2
��i�E4(�b�E��!�DσF�
��EO\ 0� �YFC!�K�U������>u��ãA$8�!�� X\"�^�2�ص�@�*�y�"O*`I4(�8~@q��N�XC"Ol}c�/Z�!��٣b�{�	��"O�1ҵ�I����6-��*�T��d"O��3\�Ja����k�)�  �4"O��Pb2E#0e�\$O��в6"Ot5ò�� u�h��O�|tf�;�"Oh��Ю�&����%[t�C"O���XQ
l�� /�*X��a!D�x��$��M� +A��c� k!D�h���/H�Тæ�*&����@=D��x�H�"5��Ԩ�F	��h����:D�`�W��6r�t��wE�-e*�de:D��*ѩs�T�5ƅA����<D�Tks��b����N��e�F�8D����\�KK����CO#k��@x2�7D�8�5J�83R���h���܄��(D�x�āX�?9�1��ܑ]�vհ`l#D��`ңK!�%���Z�9}�� D��@�>]�>u2��q��$$�!�H/5$r�$(	9Nbi���S�=�!���G?���$�	@(Dy*c%U�A�!�ͼ~�������ȢB"�!�dL�6஬���F���+!�Ă��@2��$m��( Q&!�D�,|��� �Î+�y�.A-W!�طZh�I�$	6(�x`�p#!��9/XI����(A.��r�!��H\�ʗ�ʿ}��eO�3�!��<3��Q��� �Ν�bl0�!�D\f��T2�dY-L����ȇ8�!�٬�����<V���v��)C�!�D_�1����lFoT�5���I�s!�DI�&���J$��Mf:Q�$���^g!�D�E�.�pA�ϋ5��*�EE�G�!�DI�=����-�Z�����A�7N�!�dM*r���V�
'o]"5Q�� �zQ!��д\>"�5A;]�[D�ߊlO!�..T�y.V�`"P�W�5GK!�$��8!�U�J�J��$9�/��;�!�$T�"lBĪ�d�"�Ι��.��!��R�H(b�E��L	��E&hX!�ĝ�MO��I��1
�`i��0hH!��a�t`S �,���J��ըZ6!��:��u����S��<"V��%_}!�dU5}8<�cc�Z����M!��ޘ t&[�n��k�F��!�D�2A4�����1�S'-��B�!��K���R M��<�0� m�6g�!��/�.sG	�3�6\ل��>A�!��**r�-�p/�Ǧ�ba�� �!�D���j(IW�A!5P�=�����!�M�A���)��2d4���&�}p!���t�f �W%ύ[|8����2x_!�dX,SZh��!J�!Ǽ�pdD�f!�RF@���K:y�GcN� �!��]&}Gp��ؚ�,U�a��Z�;�qO0��)�k���:��F�A�\d��|�-Ce�z�L2Ų�)$  �y ��1^�5S���#.�t�b�N(�y��-(6=����78��4*U/�$�y�� � ���J4�0�JN�y�H��X� ��,V�T���!��y"J�(���0�ć�F=��A��9�yr�<ER��雱.�EjĎ�y
� ���#&Ih�0@30����"O�$:@�ڀ���PQ

/�(���"O�U���� � �`�H�=O�,T�t"O�as#a�)��wh��N�N���"O2���M՞mL$���0�~|��"Or�BEa��L���I�O���M{7"OX�A�gq���3O?�jA��"On񣴢� Af>9��,/.�<c�"OT�;�Ս�P嫒nӟ}���5"O��*A�Ӈid �'ȑ<܂Uy�"Oƈ�r	G�/#<<�U�=7�e��"O�Y ��Q�\�JdI9J�.�9�"O�����ަpjz$;�+^o�~�"7"Or X��<GY�9`ba��Vq4"OJp�Hأ"�8��v� |ծ�XV"OH�;���"-=ȨX5GE�s�iiS"O�U�#KφRKF�e����"O �@��ة^�� R*�;�ڨ�"OⵀëT(L�+ 7}�L�itEJ��y�E�FZ* �#�\6n��0�I���y�ʞ#��2���i��f��y�'��ƚ���,D�N��l��LR �yrL a,&t�����W� �G��yүP�v#��"��â�2�sW��=�y2(	?nҴ��Kµ�j(���#�yR�	9�M��!�?vp�+�A��yBb�lǤ�z��S�B8BF��yB�� ?��*3������@ժW3�yB�6sn���B��6�1�c4�yR�A8^�h�d]3w�$���`�y��Pi��˗Ě%>�N��%�K��yR��:e_�m���֕e�Eq�ET-�y�,U�%�8�!�C%վ�fl���y"�R$g?.i���N�7v�@�B�H=�yrM��S��`���9a��x�����Py��R�zt����ˋ
8Z `���S�<�a̅Q)b�	���Y�I���f�<iq�2I0�{�a�;�XX�C�[�<��ݑl侨[�g!S����)D�DZ�.�?J���C���33�Ĉ��k+D�Ě6�S�l��iٶE�;J�^-�v�*D���Y�%6��EH�^���9P�7D���dU"�Ejp R5'|�e)D�X[p��lH1��'
��š4D�����҃��� ��
�X��+2D�(C�	ތ	�����+�x�$K;D�8��\�b���¡B�'.�(T�%�=D�0s֎�<�nP�v!ں%��S��;D��['ɦ&@�$A].Q#�k�/%D���v`�&!���$&�;l�h kg@?D���t��NLh=�a��b���(��;D�z��V�@а��G�\���q��6D�\p�" T��D��o�h7x��f3D����5v��	ö�	�J�x��<D����	[(	�H�SD5�yCG7D�tc�K�a��Q�C$������)D�(����:w���k�
�6I֩�G6D��i���w�tAe+�uX��-5D�8C��H�:%T)�I�|�Z��7D����Ül�Yp�Gִf�r�
�;D�<ԆF�.� ��!&҈djE>D���V.�d ��X2 ۦIh��td;D�|���Ǎ=�0����,��<��'D�H���H�vxJ ���[�D�H1��%D�� �ءUm�e� #���m����V"O�cuoʸ��]�s䞴T����"O�H�J��䐂t+Bd��J4"O�i��#��<In��P*?a��H@"O޽���	#��Q[	� O+p��"Oj��äH�7*Xs6{�!��"O@0��M�wl$D��'�{\�UC2"O���C��q��=�����Gc�e` "O6��'�J ���F�Y+I�\*�"O����c^=�L �N  q�m	�"O���σ���t U�F;g�@��"O�ei3C� ��HH�BLr���p�"O T���A���I��H�#""O }�g+�'���f�(����"O���Șh12u�8Wގ���"O|m�E.1#P��'�ze�*�"O�h�1�ΰf$1��
'c2�;�"O`=�@=9�¸@㛟)DV��"Ox��g��_�@�p#қ>�� "O8���V
 IB�)�!�}�T���"OHH ���	�*��� C/g���q"OTs�D¯>.��7�! �Y�.D� 2�o_��Z��3/�'�j��a+D��;7����Z�O9q�2P�)%D� �'@��I�b��c'�*T�p#�!D�x�&#�=i@:-(B� $��Hӥ$.D�lѭ��M�4�	4�yK�O*D����mN�BUM������Y�Uo=D����H�sd��a'.�4OS��Ve:D��06���YRQc1�;����#D��"� ]:��C�s�l:��#D�����J�&�,t:� �X��-D��i�j��tD(����z8�\�aA*D���w-^7h�T2����OEB5�.D�<xq�P1k�AJd*X�;&�A�B*D�h3��A�I:7�~Q`�H+D�T����xĹS�ȿ~�@�''$D�����a�4b���2j�@)b.D� �"�i��@�m�,:z>[��8D��٣W�b,	�PB�훵��B�(}�񹰧çW8�a!�c��O�B��5���M�h:x��� c�pC�	VQ�=�4K�u���@
�i�ZC�	��&5D�Y	�d(�J�7�.C�6n���x��GV�*�b���bZC�	�_��0�¢B���4I��T(�C��#xN����N����7d��@/�C�	?)*8\�e�Q�;�NH(f�(l��C��J����ʐ<+�v�i�֦Y�ZC�)�����Ļu�F���`к��B�	!H�*�2��G�W�`a�јC�ɡ1�$8�V���^�-!��\'"YbB�I�<��`�*z#�M�,:�B�98�h؂�Ԯn* �*��2h��C��|� �AO��u�1
��#R5RB��	���Qe�!G�
��uO�>d;�C�ɿE�HB �̜�@�)#ɟ�z��C�I��2�bC�6�U���3��C��6m�V���'@x��ãGE�3g�C�	fK^�
��E4w�8p��D�*�pC�:�N��&b"fٮ@�5�MpC�I!rX��S��R�xH���p�C�	�[�*h��̭�T�p��ՙ\�C�I	D(
C^6s���i��e��C�)� n�	 ȃhEY#�MD(Xz�Ц"O��""�#ⱡ/���'"O�8R�'��Yx2�8y���"OR��(�l�zةVO�.V��J"O�ز�ݽwod0�s��"}d���"O������$�X�$�;F����"Odc��X$%�+w�>�X\�"O�x`�a?^��Ę��A���i�q"Op���!H!R�J)F"����iy�"O���g֘#v|��b^�@)��"O<���V�M!"@ч���d$402s"O�ph�,~N��rN&��a�"O��Jǘ#KlA����سG"O�� c�A�u�B1�g��{���"O��ڂ�C�;.	�0͖�7�rE8E"O�aɣ�ٗ`���jҌ�Dp�q��"O`��NO'b�� �L��Rб�"O�X�d�� XJ��%�Y=�|<Y�"ONك�5@��(��C�$��|��"O��¤-\�m�d�yWe��@� p�"O
�J� O�W�t�C�䎽af\��"OT}S�m�d�ұ�Ƈd�
hSQ"O���"ӾYB�"�ڇu���C"O�Xja*�D�ȅ���;��Y�"O@��#�>.4Y�.S,/��i�"Ob�q�$�4TW�P���T�A"O�a�,�"aPz��T89�a"O
T��!>9�X����P�E(D"OPQk�ť�6�Ԧ��m�dt�B"OT����X��ك@J���e"O*,
3C�1ک;��cJ���"O�P�@�ֿ#�M�w(^�e��Ń""O����p����� >�����"OX03ì1�`Y+�Y
N�H�V"O,*��վ���A�f�c��S2"Or\��.��{t�  kΖ~�<=&"OV�tn���Й"jD8`��KS"Oj��5��:ZO��sR�>T��:@"O�e�J�#W�0)3��=Y��D"OI���M��d��R�]#�"O�a�#A�n�rl����`AJ��"Of�d)�z3�\sI����U"O�z��Ld>��r 	�ʀ�S"O�a��c\�B�P��a�i� �e"OxXDǅ�P�j�Q��֯7��i�"O��P���
�t�֠�-z���"O�6J�8dX��R�F0xf�c&"O�U���9yu�0���]2�B4�"O�����>'����ַ��֋�yr���Y��!�$�z��#P�y��Op��$#�X8���,��y�C 5H^ @EA���\�C ��yb�E�O��p��
��#fI��y��� "�L!dNJ�8��S�*X3�y��	>R�$�a�f�?i�0�U����yҀIv��3(�:��I0�yr��� Z-��O���%�ȓ�y�� �K+x���
�Ȍ�j��a����Q����1��ժP�ȓ,�:�� P�@}�BK�[�
}�ȓE]�݉��� jA-D6E����=�&�2v<�,��F$%^`�2X[�U�Z"�*I"�B����O���B�	%W $�rD |"�%J�B�Ic|q�a�;YVMX���Z�*B�)� $%��	���zWgF�F��i[�"O�$��A�b�28pFF� 1��W"OH��f� <(����H�)�"O��$OS`tD��ؕK��!�"O�l��]rΕɶ��Y����"O�9s�C	@�J�z��y�l��u"O*Ї���5�x�vg]3g����W"O�uB�� l�������(�"O��S��3��KՂ5@�Ypf"O&@H�D�A|Fd�� �8�V��"O\K���Cu`�o�>0f��"O8�*����v���!��
�"O���'��6U��wn�1P	H4�w"O�q�be�����I�F��
��"O����GE� �����p�"O�ȓ��3��`#S$N�l�h:�"O��h���N���tH��?&f��"OX�k�61w�!"ƔZkVXSe"O��(҈ֻ&�v=r"fQ���'"Ob�QW՛P�|�wŕ$!lf�"O����L�^�QD�19��H�"Ol8���:P:p�J�%�=;!����"O|4�,�<e�ݘF*Am���U"O8L�[&3�Z�4��->X܄��"OL��&eZ�0�ԡV"��t�aa#"O�aپV�s%��{��(!"O��j��Ta�m�s�J ��h�"O��	lR�j�Ƒ2c�MQz�F"Od�׃?1?�`b�Ǟ�J�\�u"Oe��e�%z.���U�,��"�"Oژ9Ă_  !&�C�B�x�b)2W"OHq��,�x�#B�?9�V��c"OP]���vn�a&�22f�+�"O�d�� N=i�ȉ�`d f��W"O1!�@�
'Ȧ�Zv��F����"OT����;6����@>\�m��"O\��F�r���ԮA.�6���"O���j��k��|[$ϗ�K�>�2 "Oxa�M���0���`ǌS�`�0D"OT�#$�=�4#�K)�d�(�"O8U!�L��'!����m�o���"O0S�9<�Z�-�ɒ��"OizA�A��~ux�"�(,�V%Ac"O>�87��h,���r��D��"O�H��IЀYg�:%o�� �hY�"OP���oئE�x���Kְp*4���"O��"*��΀��i�6$�ʅ"O` CB�A��`�����	{h� "O�T!�a[�R���d�][΍Q"O�:3L'���P�h~�d�G"O���GC=Jj���ț@��p�"O:�H�@E�wpl�B�Ө92]A�"O1i��@0_YSlS (Rm�"On�1g�_�	&^c��5���"O�(��T�� �;f�]�&q�9!�"O��!��-#���*�Kg��0B"O�d"u���n zC��X^*%t"O.Q�vB�8}*Ę��$]&��H��"O�aCb��<J�J�3����	�v"Ol a펒2��;���:a�|1xe"O09-A<2�l�$/��ʌ0"O2�3�G�	%8�u�7���m��k�"OV\#g&�0Dtջ���?|���q"OP��'*�΄ѢbL-�<ȓ"O� t�����&)�|��"��a�&���"O��K�݊�b�F`G-���""Of�0�(����LE�.-��"Ob��[1�ڽ� �gf5��"Oz��3.X� ��W�M�6`h3�"O^4a��IV��T�V�WP���e"O�8���]w!��H�:?�{T"Of=)%��=7���H(A���!"O�S3 �2o
�Q�`V"���4"Ol���@_Qj��F>ǴA�U"OZ@Qr��1�r��g��4S��2$"OXՃa�.l����j�5%v���"O`i���Ҋa6�#עjo�h(�"OFś���8j�:�!iPeC�"O
�+���q�X2�ye��8!���0������a��a����%[!򤁴Z0J��VcM��xS刐�of!��V6?�`r��.oC�QX�I�,9H!�D ��o��WXxa���DA!�$�<�<)C��˴j��p�'ճ2*!���p#��+�oJ3?��,P5\!�S63�t�r�i>��I��2I`!�J';KT�� �Dؐ7�ތb4!���eCm (@+(��9%�+�!�Ĝ�g��(�hL5����ǆq!���ȁ�M�PAKqלn!��r~�Q/A0��:��"0z!�d��DP+�M�ˈ}xQ�Z�ps!�'w��U �OɖeR�*Eb�6B!�k�mK�j�9�L���^>!�Ҧ1����c�W#
�P����H�!��S�2~\u0E/ o{T���e��!��i��x�B	��3_�ɸV��e!�D��l]�@��ė�g0ZI)ƧL}T!��Ccl���lB�Gz��A%T�)�!��ΌO�H��N�F\BM���
2�!�d�J�[��M lJG����!򤃌f	�U{�75�B#�>Sg!�� s4�@� E�3M��J �'�!�dW�1�,��b�8&��	�쉨C�!�SuR���*Y�h(�I���!�%T#2p��8@�ıX�NYl�!���_�~-cF��_�"9���]�b�!������P���L�`%��#N?(�!�dGev�Crʕ���! �44!��@}���)���_Bа2���=!��?$>H9p���,t��cĐ{�!��s����3�,�����Ud!��3�@�vo
C���&ʆ4bc!�$S�މG��8eKn� ����mb!��Lcnm���,J\�R��o}!�D�
j&͈s�5�	 E��_�!��")n�Q�%#��9C�P�C"p�ax"�	�S�[��<'.eZG&'_5TC�		 *�p�$V�Y�"u1���b}�C�I�Uv(Psuˌ��J5{�HG�E�LC�?��miFJ���C���'� C�I�9�j��*��^J��[�K��I��B��2% �b"F&��҂҅GB�	�U���O�8�*�@+־�6B�Ik�x�
�Qi,��C�5<�LB�2Z��9�A�؟7�������DZRC��F����sKT�Lbt�v�W�n`\B�	�e�2��@*�:�H ��k�0�VB�)� �C��W�N�pL����Xh���"O��b�"\�z|qe'׆i`�I�"O6��Uˢ1�L� ��!z���"O�1�Ʉ6J�@�0��:��9Q"Ob� �?L}ʔ�s*��hԋ�"O��9�b_%XH��k��~۾]�c"O��Bʓ$=]dEWHбo�j���"O���`G�R�br6�S�B����'"O�l�d"�slp�UJA���If"Ozq ������ϟ
j�~��"O���B��K-�,��/�m�,4��"OL$:��)�0T�lP�	���`"O~E�f�;����3���C�-:�"O�P!��G�^��i6��/ 2�s�"O� ��H�oSx]S5�2��9��"O�h��ȭ��
1��"O��JD�PH(�%��"�q)�"O���ċl;�}�wl֜,����F"OF��HV=97�5����9�1��"O�ph#��=qޑ�����:�"O}s�� |V�P0���RAi%"O��@�gP�\> ����$6���"O�t�ch�G��ڒ�/3����"O����/;�V�"b��w��V"O�䪷n	�$�I�Ъ�%(a�DJ�"O�|����4U�ج`U��5BX���"O�ձ�'J�p��=��(s-pp��"ObM���j�N	X��
b:L9�"O0�Y�-B��@*�I	2&���w"OX��GOR�Fn�)��N�t�t�x"Oh�:ԇ�,-:hq�R$[t^�"O
��OɁqe�ݺw�!�-� "O���5-O�j鎈�L�4�Tp"O,�cP �5(�P�R���=Q���s"O6����{2�N�&�|paG/�+�!�CI�:@���ӎ}~����8sf!�*yѮUcWaG8%�p��,��
D!�đ-6���$������,�=9/!�+y�qس�A8f��r��S$!�Ě��}@Wɢ=�6�,�!�D�@$���e��G���jR*w!�C�0	��{�D̓}]j��(Y�
!��=(����L��Mp�T����G�!��w�
��'�E� |͐D
�+�!��J�����˖Fg�I ��]�k�!򤟵~Yh�*K+B���%==P!�䔧]��B˕(8�8��I%{>!�䜗Bx9��c� ��Mʶn6!�䏂zM��A��-,�&e��Ͼ`7!�dݓ0��r����pQ2��1�!�$IE� P�3
�����ǝ�&�!��S�y����E�E�J��H�,`2!�������$2B���jȕG!��GZX@<�E����Ht���&0!�$� (W�)�%@�4�T�ȁ�ƫX�!򄅆x��1S�.���8���֥v�!��;b��a���P��h�^h!���<�����~�`Ţ�L؊= !�$E�/��Lv  O��I �19�!�8l$��@�DE�J8j���*�!��:�
]�g�ڨ[yZ��e%Տ!�!����Me�	��I�;`��0�m�M�!�dC�_X��#
�Zh���șf�!���"~��-Q�N�#�|�� �$D�� ��:�$��1���P)ԇ]���q"O�-h4կz-Z��"T�1���R"O�b�H�P�2#��N��u"OH���J�����L�]C�Ȣ�"O�؂3N׼`6ށIf�[ 89@h+�"O��Y��G�@6}�F��6�A�"O�1��eA<�����ں�p��E"O ��& O�E�4�јw���E"Or8@e�A Ȩ�	�/n}hZD"O�h���ָa��iIs��8�R�� "OP���[IG��hS �D���B�"O��GB�
,�:��R�=jm���p"O0K���|0������ d�K"Od�C����
����N^O�|xf"O`\s�N����ۥ�L�M*�AB�"O��!N�6;� �7�:A����"O�-� B�C���ǡ�H�l�#"Oz=���Q���Pp��.TXٕ"O�a�Kl��HA���*��0`q"O2�.]��}�dJ�fz|�b�Z��y�劎7�vi�"k�_�$�R���;�y��S2 �Jd�"$	,+\��)��N��y2��"o�~�(���>*#d�!׏�#�y�PL:�c���3#�\V���y��6'��X�a�ǘ{�V����P�y2삣z���3�@$zm(T�����y"��-��q핪Gz���X+�y2H�"4�ȋӎ��+�N1�5��;�y��C�s��|@@(7�Xi`J�0�yeT�������07�>LS'Lŏ�y"
F=S���s���$1A��
�A�)�y�˂\�ni
Qj5!�~���E���yf��	�*}d	�;T1H�:�y��J
��3����|ȒT��y2oHG*��Jt��
ꡨ�,[��y	HE2��/H�	pi�ǡB8�y�N��\�ʼ� �-6ɴ����'�yC)$ q��k�2~���t�P�y�L;��4@��T)�:�"c��8�y2�ْZ�ۆ�����1B����yr�V/��z�ɚ�L�����N��y�oS�\s�e_�C���Io���y"$�
1�W�2���H�hW�y�X�V�' �t�r�� N��y��_,�8��ѣ�$<�� �R�Y'�y2�[�;��|��H�iNE�����yRn�Z68��DO�}����y�-P�+<u�%�HF]FI�`��$�ybJS]|.	�P .�� �uƑ��y" ��1[��Q��� !�� �$A�5�yB"x����)媰�I�y�h\+=�8%$߸y��YC����y����6��;C��-���2���y�M�jD`#aL1Ht����y"K	o�j�32�%R��=ۑ ��yRiΊ����� �^�L��\:�y����t4.���dM�\��|8�;�y����rLS�t� ���S��B�	�5��t��|*���jƜj��C�=��jVEP/@�ȝڂECU7B�I�g|ƍ0��Ɩ���f�C��60��<�r��/;k(0���:^��C�ɫX ,ċ6�x��K�Y]B�I�Y���"Ȍ�>ߚx҅�X_��C�)� @�����"3�����Ǖ8�쌊�"O�Y�`!C�PߖTȂ�N�R�TI�g"O	�Vm�5d�M8A �pw�Q��"O�*FO�?d��I:!��"9S$TѦ"O�ei�	�M��4{&�3O�L�P"O�������(`�fF�~<�P�"OJ�(���Ua�H�Gd�@2�\k�"O�pP�N��i�0	6(*9�"O�T�c)C��B�n���"O�l�v��O�����_���q�"O��ʦ�K�wy� S@���!�N��"O�$�GMI�mG|��UM k�`ɘ�"O�Ijvb�+X��܂T���� a�*O T�vǛ�o�Sg-�0ɞ���'sV��%χ?)I��c3}���(�'D`�u�Bq�}��F��͠�'Y�0I"nM�eö�#�_�9�@���'���ifd��U�t�!@��;{֘��'"�����E�+�
H�ᆐ	4��k�'��Yh�͈U�z�01 ܘ0���
�'�`[0JV�NT.d@e-Z�#v��	�'$��ޙ$�� J�@N�#�dh	�'�*�� N�(tu��(ۜ�:Hh	�'�L0��ޥN���c�

.�0���'�D��)R�C�� 0.|س�'�� ���-6�y�ţņ#<|J�'jPLآnȈ&(j�H�Y�aܤ;�'��	p7����x��e�7�X��'���gZ��ՍO���"�'�:��Ƙ6bTX���ۘ�h9�'t�9)�ɳg�,�0 ꛞzb${�'�F$����3����M�����'��╠-?)����CG~>��'g�1��	m���Z��ǯ{Sb�#�'#r�K�ݜC'� + �+h�ްH
�'�j��p�]�<h� �'�/d`u��A����	�l�\�De�.8�N�ȓJ�4�F�(n�
�!I.l�@�ȓA�4���/U_N+MQ�WV؄j�"O�h��,G!ҽ�a��bQF��"O��:�G_�W'�4)���Dx��"O�m���c;�-`�ǅ�$=`U��"ODLr��D�9��ѩ��[E|�m<D���C�ț��I�A�4IV\�C��/D�X�S��9=�f�o�� D8�).D�t ��B-GN��j��1�� ��n-D���U��*��ᓶ���iB�8�
,D�ȳ�H�x�U�R��'X���W�'D�Dj4+ȇe&��#`GJ�g��%�v@'D�0�Nu�H���MH�!�\:Q�/D�����&4��t�6Aٺ:�<8�2�"D��9�d�E��H*w�T.}�$���?D��CW�0�>�f�҅e�"�C�<D���Q!OG@z�F}堣rG��y�M�5u�8p]"?8ά��iY�yRlU�%-���ʂ=7Q��`���yR�[���,8b$Bc6`}�kY��y"Laa�D~��]pV��(%
ޅ�'v�����GGJ�Ds�$Y=���'g�U�Q�ąa3ʱ��ZB�I�;���s�� �F�:��$��uG~B�%j��t�#%�>c�&�J�*%.shB��s<d��!Ѻ2_I�tG?_�`B�	!`P%KNU+2�� �S�հONB�)� �taHϠu�(��`U�a��D�Q"O�!��;CF6����3il�0ˑ"Orm��H�]7$x�`�N��Z�"O�S�IK0Z���UI7��@"O�E��2[C��:� �"OV1X��6j�8��A.>�^�f"O* ��!�A8���l�h,A�"OF�IĢ���.8�������"O�M����3b�`i���.��r"O�P��O�5y�Q��/3���ڷ"O\81��8��R�Jh���w"O���`j�*\��0IJn�`��"O�L��	_8/	L=��)H��X��$"O�x���m���"_��Uap"Ox�@Ĕ7�uRP�I��h�q"O�<�֎��5�Z`���@�`2"O�m:р>��48�U=$<��"O�@��q��$�	!tƤX�"O�:�nD20%V�)��x���˧"O֩p$��h	��r7lA�gMHr�"O��B��P�<��⑋�c.�d�"Ox�y��	�A9�|A��'b�B�"O4����au&�@7���m�"O�EA
Щd�@P��m�zh�@"O�@%c�6L�1Qgɟ8���р"ONu N�\��U�ą��谓P"O6A)U��6dF����D�=�L0w"Otxs n^6
�� �vBʉB
�,;�"O�2窈�W������T���&"O�᥄�~6[ړ`��YJv-��"O]�փ�	j+RAʰ,��h���F"O��񤄼������-;Ѕ�0"O�)�4�E>����E'O
\Uމ�7"O�"�H=w�<A*���@��`"O�)����w���t	L@-�s�"O�-�C��/9ˤ!HW�Ѻ^�|mY�"O� �B�I�V�C>��t"O�yI'��$/K ��BY��a�"O�e��L�N�xRq͑�]����t"O �r�&*W�Qb�l!U�<p�"O���sG��c�2�"���?����"O4�3���:�P� j�q�R��"O��{�f�I|N�c�
C	a^i#�"O����ݡG�ƀr#�)Y{X��C"O��P��S��x���K2=b=�"Ox�U@;c�D-y�0D�r(�"O��
&q<qʠ#9Wܞ
�"Or�y��U(Q�ʜ���k��b"OF� ���&R�z$)`%�=�T�u"O����m�,O�� ��2�\q��"O`��l�)m���F-������"O
L�"��9o�X�Em�����"O�j98�*�Z1�������"O��a7�G� �� �`xX�"O�=[5�
��h��d�ئ!�lqK�"O����K>l�l�����Xp��"O8X��ʇ	�}Rg_�T��]�"O�����_���J4䌋�^���*O�)��40��Kr*�:ߞ��'����ׯ�
>��]1GlP�[����'/�U�g):5D|1�N8��
�'�pLK��Ks���U˛/0���9	�'X �Y� �U�`X5j�� ����'���؁䑃{�8C�&B�0��� ��B1�Ξ�����A�k�@�h�"Oh�!��]3*k0r�gu���T"Ob@�eDC�B}����<E�x�"O��"I?%A�� ���)d�KW"O�X��lH�L���)�$SH ����I��T��]�����U4b����7pt�s'�53�\%3����<�I�+q��e�~h�F�*Em��4HY���i�����à�'�������q��(1�&�\=  �8`�z芝Z��e�==��C�#�v{�Xp���",Q�0�Sb�,Q����mڴ�?٪�����O�r�PLSnG�|EL��$G]ƟD�?E���i��*���� �tCӸ3<���)�2�M��ߟ8ѪU�7��9�$E8�ڕÄ�O\��UOM榉�	dy�Om�<!�ɀ�;�V������ �:����H)������	%X��I`��2z�B��S/^�'��]�{6X{aÉ�j��H9�g�b�`7�ʝ[B���S�_��P�V��0^��ȹ��
����A'�|��>�,	��/�\Q��ѻYRk�iJ�����FjsӬ�d�|���ܴ*N(���F�|��+��.< ���?�	��ay���uD(t��$�!Ӏ�p!�D�Ϧ�ܴ���J\w?V Qc��eo�4���T����<1��ݧ~2���'PS`�ƅ0.��K�s�j`�4��,b���f�ᦕ`��<�4(��*���Ձ�
 �i�%�7*U��1j=��	3�S�zp``�7���)�0����:�t�'�>qP���(#K.�)��\��+1��O��:���O�qn�`%��<ǻi%��8)�����AD�`�0,�D��%V��v��h�n	zV�Ak4��c���h���CW�"�M�v�i��y���dӳ@�	�|�cK�4E�JH:��}��ly���DUj�q��$��<q��D�����N0E1��C�\H��1�<��p�������� ���#?�סΝ>P
���.NR�<�r�Q�L|�	ؤc��30P�x�㇚��WA|_� ��	��|]Ƥ�����a)ڶ@@�̱���`"�H�)��'#B�'K�O�Ӽv�ܹ��[�'8����цw�t�<˓3�ha�C��N�tAEI�)�����{�F�iӼ�\�97�i�b���*�:&-:� Rj��)����E����'��`�c^�9�f�v�v��Tȋc��ͧR,Ԡ��㏌lJ.�a�$��P�Ez�F�4Q�!H+%�����ID8���k�ܠ9�OW"{��H7�չC8�`�%@*��':���O\��㦁�I`���(ܑ���<Y�����#�V��$�)��r�	>�0�JQ�ٷ�If+ͅf�f�����ժ޴�M�uW%*��`d�1 ��(�'��E?awG��z��H���4���oZy≬M��[��ɺ'���Ƞ7=������'Fz��O_>+Ԫ�A�1;"b�>����P�q�[0?�n���kWT8tۢ�i�0�2�]e�y�0���\[p� 
�W��`�7%��s�MR�M�a]�� �cG$Y���{� hӴ%P��'�r6MNcyJ~Z͟����-�4�ᥟ)�BA �L���	}���O�Fm`���'D�	�K�h��<r���榭�ش��O��.Hi�2$��O̶Bpd`#�U�=M��'�����7`� p   �   a   Ĵ���	��Z��wIJ(ʜ�cd�<��k٥���qe�H�4m��_;:<��iF�6��/F]�1hA���>ᜭp'*��,.�n�*�MSַiiD�E���$�j�2��['v���Bf�f���Hy�%{��[�'���nZ�^�=AS�M .�B���i�a����xQ�D}��1�'�6��6�J�X�Ŕ'�h��pE�N�pYⲋO� ���3��=[$�qشHE2���'АQ�_y�5�fT�E
g4�52э׽	b6����(-h��E#'���Uv�� �H���d�3X,D�S�q>i�"�̫2��	�/J� ���������$�
b���EFߤa.1Ol���,(|��)t��(ZflhtOe���2ቾP��ѷ��[FvXҢ�j���p���O�=x��$�3��$���Y�����Ĥ㶁I�\�@"<	Q�=�I�.?$���-(6�(i���}�(6X�OD���D������d��`�pqꖣ�#O�j��$L�O��q�OxE��i'g|�	BD��M��qY_�
��I�A�O�92�×:+���ٰlu �#R퇣�OT����d�
�?�e���+N`���n8[@�s�n��#<)��*�D��fz������U��PȤ,�;����'�OhUK<م�Oth�V9$���Ң.GR��h��'V�ʓn�Iv�_��D�1���|2���<��y ���>T\4`���~y"���R�H>�u�Q8&�bq%��� C<9 ъ�e�*�Դ��d{Ӿ��[�'��EFx��]���af�G5��EbF��y�C�y d  ��%CI��b�0!�Z;[y�a+���:m��8Q���!����x$i+`a<��E�!b�!�'=��iAQ,n
T�wEExA!���!:p1���#[d mJQO"!�d�@����`�
*\�\s��	�Py"j��F�)b��*`HLs ��yB�s�v�Tj2(�p��� S�y"��.fD0�u.����&�D-�y�.G�d��������}~PXG��,�ybI
~3�x��+8��	B����y�'�+�p%��)2n<�/�y2����2�A/lz!��]��y��q)\HS�")�R�nB��y��E�0��❂	<��*C��	�y�-�+#Č��@�2 �써B˜��y"��q����Bu��Qr�:�y��S��t+rhW�P   �	  �  #  �  �'  �/  �5  "<  {B  �H  O  ^U  �[  �a  -h  qn  �t  �z  ��   `� u�	����Zv)C�'ll\�0"Ez+⟈m=�R��/{|@�D R�ؖ�_�}�X�stM�/q�L��J�0����` �{L6J�G��,�;�`y��H���{�')`d�5F�y�x�s��8'2aBLR=�>��"o��7&��Ha��U�ѽ�����:�D��6
���0�AGbTI�ֆG:l}�2���δ��*[����S,	�RLd<��4iq:���?Y���?��w���p�Ν^����1�!~/������?ɏ��'I��S��Ip��L	�.D��Hg���@|�	3���'�R惓B7��^�?)�'��4c�[3�0�5�&F�����-I'�R2O�Բ2KRK���ˠ��
G�V�*Q�xFx"�O�e�G*ɺ���[/��%�D&�1a?��
�JC$)���'y��'���'���'���'��cq�Q 'Ț~�nBb���LY�4z��&%}�NDm@�4SE�VB}��o�Y��ٸ�p���99t�A3�F��x2��.xm��@��=��� �B�0$�키�/x�� �N?��je�Бn�?M�;Y:��i&W�����^�0O�[�.	:wJ�Iݴ���k#k���!�l	)}�9����'+v�pJز���V�ѿ$����''B�'�b����x���T(�2Vsx��D�O ��3�S;-e��y�(@8[41�&�W�0�`ʓ�hO>��	�:v�X��L#-���j2$_ğ D{�'�����Hj�z�'D�$���� ||��K@$A.+�>8�	vy�'��>������P��	��/;��6�9�F���	̓ ��`!���6Oxhjĉ��փC���dCp��Tj��˗Es^0��(�+�ax��R��?Q� �Ij)L�C��p���Q�(�;p��D�O��.�)��<qG�W4F�X��IŰ����'|��<�ߴH�d��T�mk��RBcD�?��1BǾi��O,Lh�3�I�?y���@�r�h�"I{���#�Mk�<�Vm���lU#]��a���\�<����C��x��2G����gRN�<���_�ؓ3S�5��Q�l�J�<�C U�`|�� �+N O�iч@SC�<���X�B��=Qdh�"�^!Ae�ş��'�S�OQ��5NJ�7����%o8t��""O%	Ƌ�~!�`�aeW/r��c"O^���K[;8���mE~� ��"O��	IĈZ����꘿0�@��"OX�⁢�+���o��P�"O�FJ�(9������q
J��S�T���-�O�1��f�����"�#u��� "On�������O��P�"OT�Bb��r�t�;!D�;R��u�W"O�
GoD�6Q�"�ڥv_heI�"O�
[jԡl�_R�=
��'gҌ�r�fӢ� ��A�%זT���UO[���I@y��'52�'"�����58�,ݪ#�֦�N�$G�K��ʒd��@����'-axJލ^�|�E�7�*����'UƩ�%g�r�:tX4�}��d��8jv�I5�M#��ib�<����C�-l~�!sOBy$�	ߟ�?E��F�G���qD�?+��!w@�,��?�G�'����G�P�g���p��DeJ�ő����oJ��a�%�U��<��w�	`�CU��ta� iF�|�	�'~L��L]�1�*��GδJ�P���''b���P'�޸�#�ك?5��9�'�N�{w�]-@��`HâW�0��\9�'�A��^ʔ� 2N��[��<��'����� pu�u��N,G�D� �iw�'��)�1�Oa�'Wr[���2/V4��鍌{$�x��,Q���b�G���M��+�9����,��X�?a�N�B�Q�u�Ѡ(u�<蕆[���!��c���F�](���|�p` �gIf�ɭb�Qc
O	A[������_(�nZ)��<v����'���'�@�,ӪkyZ���̖��aI4�'�R⟔�p�җD�P@L�
:����p��<���i�X6�=�4�v��<�F�U�@����a��P�6��7`2�4�i'2�'�P��$?E��N�94���)�"޳{*�`���N���s�딃a(��4�i��tafͅ|�D;t�ܥ!����@�� g.n�e��gb�S�H�?��"�Z�l�Q���F(��R�q�J��ᾭY�O�TR��A٦��'���'
"�'��?�i6����L�7n��]�C��#�y�C�!��	���K�a�cF����4�f�'��I������4��)�8-r�آ�ѭ6�~��N�kYax���O� ��T��=6Q伹SH׮/b,, &�'�0���DD��q*Bǂ���X@D�UaxbS��?aE�|��
k!$���>a�:��Q�͚�yR���H�N�r��Q�\{&��5��?	��'<�,�r�,]��%���[V�hL>�Ì�_W�&�|2Z>=��y��b�BL(J>8R��%3d�����Ĳ�N9�<�Rѧ� Cf�Z�S�O0�HG�ǌ4���h&�<���+�O%�b.�=uY��ԎH�=��}z�O�u��a�Z�='��1�
�`~R����?Iּi;#}��'K҈C���qJI�'�/[��}��'��£�Ϲ,��o�*u�Ƀ���PA�O��<0����A�����5H�,��i�T�l����M[���?�������L�p*J�YV�[4�G<.2���B�ٓ?�|HlZ=J�A��bJL��.�I)?�l�c�(�,z��ũ�dI�K��0��K&O��T���@*\D�i#�3�	�@�\���b�>.p~�8�K�w[F�D�ۦ��	��Q��Z�gy��'2z��1�B������t�b`p_�����5�X�b'��U�P��qʐ/u�|�M#��i��'r��'��D_��)y�n$D��wP+��1A��Ҧ���ȟ��	Fy��� D�}�v��[-�4I�%$�wvaoӫ0"q��k,|��$0<[���#Ď��t��$ b`�Q3!�bt,�R��_�����ܵ:Px�S�3�Ґ�B��\l� F�'�&7m�ئ]�?�!�	�%%H���)�{�<���$^?d�!�t�
�K'�=C��Se��mu�'�����t]l�T�t���?���@��L�& �1dG=�?q+O(�$�O����33��A�ް	/�ܨ�	�����N̾��5 ��x2�C�+O�T�5�' Qdųg��1����|�fC�I��@��S��
!axr���?�����D�4Rhª� y��5��.�l���'�b��S�n�@@��Ā��SG�ZL����D�ٟ$� O�AW<)�E�٪a�,P��L�O��M�|�PU��'����O���	Ǫ�Lb�غ`�Q���O����'<Vjub��l�X|��.F3�MG��l
�Bb4�r��
-��u(7G����ص,5VUꡨnS^�@�R�O��=CRG�Z�A����=����O�M��'�Sȟ4q�@@	5P@\�@fJqg2q�tBP�<a��Y>��|q�kA��̈�UFAr�'��}:e%MD͘���L�d�{֋#��d�<i�����J��?����$����!jMj#
��c�Ԑw9$``q��(�
��I����/�3�/i]�@�f��Zh��DU�+=(`�W�� �P�I�4���a/�3�ɸf���yт���L �L�8x���<?�0l�ğ���u�'Ԅ�㔁_�g[p�S��O�eV��c"O��u�P�[�J\	��Y�`��fV�TЎ��?y�'����I�]Y Yu�U�yɂ8ʄ�V����'���'9�)�S
s��Ыa�AQ��R2$�/8� 9"�n	
-�ZX!���5"�A�����0���{zd���5wE�e�pT�4VȜ���0���J�7U� ʇJ �X�CAk�e�hmx����H�Iw�'��p)D�W!+ـU[B���[u�y	��7D�,j��#����ܽ6ЂY���7�B}r��G
5r�)٭㔅c􋀊v�~=3����!��*/�	� ��k	<��ř,i}!���-�84�0Ia�ᘒo?����P�M��b�>sY�ܠ��ԌL�z܆��L܈c�8�h��B$f\����g�BE��F�
w����m�*At��F{�%	���x\�3n��%�Q�^���9g"ON����,z8�CfU=�S�"OBLk���
O�@d��@�P���J�"O��Q��yހP� 3$�6Ay%"ONN�J��E`-S�_���`�"OX�S��E�"� J���?�=U�'Ԥ	Ӎ���
Ms:1��.�)ow��
��߀r�RԇȓeT(�f��:�n-3D �:Z�q�ȓ:�.�!�"�Bn��{�L�9f����P�@!�Ū�2(Ű�bTZ(ʰ�����gM�bLܸ�Ua�(
؆ȓ� ��g��p�l�p�P�Fp�t�'<�H�x�1TΝ
y�4*���.��I��S�?  �O
�(,��N}O��`b"O.$XF���2�:�m�Y9��y�"O�F��Y���!�U�-:�e�w"Op��PlE`"����-08~(�#�'ǀ�	�'e���W�R�V4m
A�`�'�z|����4�����F��:���'y
��KA!����fS�4�"�8�'����KA�ؼ���Ɖb&r�'�8 �C+[��5 �@�����K�'���Hǫb�0�H��9�R�(��D� �Q?�K�ǌxhl]Y)�p�C5�+D��iDІd��)�:�*�R�*D�8 �I�;�0���B[<kv�q(��=D�(8��ڐZ��p%�6F�\i�5D���)�:S�|�I@=LĐ�r@b1D��Z d��j �2�ܩ@Z���O�OH�P��)�禙{B���zt����V0X�R"Op���'�$��	VD�}yG"O��0�!�nP|L���H8!C�"Oؘ�r�E�ql4���C[����"O��w��M>dSu$�|Zұ�""O,�6��!/��
#�1$Y�T���3�O耲���Y�`��N�*��"O�JŎ�@��t��Ńy�t��"O��Č�)��(; \�P|�] `"O84��a�73��aI��dvT;'"OX8��/J�?Q�Q�;ezz�h��'��Q��'�d���V[Y9�	ȡ<�& ��'��Q��wi�;�S�I���'�T�%�|� �)�G�z�x	�'���زCP�[�(��tƔ6z�:���'�b��UDϽm�IN�'��#�'�j� 6H6n���3e_7!�
T����e�Q?[U�Q(%�T���(�0E>-U�;D�\ȰP)U��A1�34�;b�8D��2��O�/��mXb�\!#q�(��6D������_*�<
`4����"3D���S��1
�p��զ��(\�|��D1D�\��1j �P@�&�;6pr$j=O.�X��)�'4hP��o��^Х{+�R@|x�'���6�`����
�EuBj
�'��P��>�4�Eiկ=K>X
�'�`�� d^K>���1#ȭ�	�'��M�+6JlxnB�@�i��')r��R
[�A��Ih����y*/O����'ab�y2"C�~��$�D�Ko����'���j��D$-�Q�TI,��1�'���Q4B�
YE�����\�S	�'��=�S�/1�xd*T!4Zp$a�'Xd����:
���c�X/�"x��s@܅�5ݼ�k�j�Ju*��Q�����"��(�Ձ]M�2W(�p.�E��P��5Q�ΟUN��d�wT�5�����Ѫ�$z���VL�u�͇�טy�v���W$x�5�:s���ȓc�����C�rg�ѷ�B

�ʌG{�G�Ѩ��1��'V1ha�խl��j�"OE�B��}f|P������#"O��pSJIH�RM��ĺ1l�G"O�dx��� ��"WN�@��0�$"Ob�zj^-d�	A��[�!Br��T"OTA��李OvU!�A�b�I93�'� s����N���^�.�:�Ir�ZGe�-�ȓ[��P��	�F�@`ͤ;<��j��� �ʁ�ؿ?�����j�pˆ"O����ʜ�u�Ȩ�'/uM0�Xq"O�Htg	y��X[6���G�a
"O>�0�Ƃ�fp�]�g�$FN �2�\�<r�� �O +D�S*_^H�g��0�| Yr"O�@`CA]6���cp��<t1����"O(�@�6��J����)|���"O>�{"+��|]h�&;R+u�p"OF �sA��j*L �fͪ|��us��'r���'	
�c4�L�g����R�;AѺ�@�'� AA&Ϲr�R����Z�:u����'��lїǱ? %3a��2���'r&�Ƃ�7>��0�1/��9q����'XlQ�ɘ$W��S��@1
F��'}fQ��AH���m;��)��`��d� &+Q?��튷0�,�ɶF+
p2�IU�-D����Z7D���[�Zc0
�'1D�8a��A>I�	ū�!b�X#%K/D�ȹf	�(WK��𱪖�K;�c2�8D����]y�J�����#>�(Is�n8D�����S!JJX��shZ�[%D��i�O��YS�)�OHL���2>�B �F�0����'r�ݫv���	)P�Z֯�,u�\���'����5́�B���&a�$pӈ�:�',��B-7���C� X��2�'���`䅕��je�#N�j���x�'��)�#A�)l�z}�&L�2�U�+ONt�'"6�B�/I�5�p�"e��A��  �'v�L�����XįI�b����'�X�r��$[�`��hͥ�����'ώ�6�O�+�G�?U�88�'�1��ɎBlPȑ��)<����Cf��g����%B4�ZV��/!4��U�6m�2�^�Dd�����=?�Lp�ȓG�8hH%d��!��	
��'��u�ȓF��ÇaQ�3cr���.�"Їȓ*�Lx��eH�	(�kg��T�\]��~JH$R�o�; Ԙ���%"�.G{�c@��^|�� �8]=��b�$/��c�"O֩Jѣ��Ќ=�2�3�m2"O�`��CѪFU� ��J6~ 8Ի�"OR��$$ݍ;ՠaj��L�	h�c�"Ozd�a�صf���$��T���"O$�2^�<<N8�r�(bI�lQ�'82���Ӽ6&(��W�XW
�jt�3KYȄ���B�c�#{$��Y�lc2�ĄȓjDn<���!&F$�)+��2�,��ȓ|�ȝbeV$����hV�8�X���^%�C�%���x� 
p��p�ȓS�l��n�5P�	^�Fd�E�'��E	�@��
7�K�US�(���>48���dfxIa��׀/�TA&Ø�Iz���=��!��^e`��yE�E�ȓ<��꠪�D:�ϋ=-�T��Kj��C���2�z�ڣ�@�O|-���0����Nۆ}���x)t�p��բMgjC��+D�����ǏL�tUB"�$m5(C�uo�mq�')ng8�Q�G7� C��8%�жG�V���1�ӧA�C�	oS�P�0�B�S�L(�v	g��B�ɇJ4�5�Ce��4�k��Խ1�Ģ=�N�r�O��,§a�7a!���U-S�(X�'��Epb)D1=�a�F�%K���8�'����ϋ�]'�M�"f�.��EY��� �-�ҫ	�R{��*s��K��H'"O 0p.�	9��}з�/\>@�"O����lǀ}Êu�u�@� Y��'0��#����3�:hp��0
�Ղ�̳%����ȓQ�����#Cb��p�U䖕��ȓLX�u���U�(\�0$�(�`�ȓ�Ru`с�A��[e�_	<t�$���\�0DE�Fx�z�O6 ��ȓAJ����	��xz�?R�@��'��]H�
a� ���ɐ v�dZ�&<k,�ȓ����^� �����^	���ȓ�>Q��H�7��0��
1:�����M��)���|Xn$xD��"g��Ʌ�<h%m�;ej��f� ��ɬ|���I�5�$���@f~�1�9+T�B�2lyJ�Z�ɄT�ld�'h)Cp�C�I)r��cE�tN����y�C�	�9��J�Lk�]d��
��C䉘0������|�v��RJ-�VC�	�`��i$�XVѪ���4�=)���|�OM($�@�fu�����ݷ{5$б�'Ϛ0������*�cwA�,dv�[	�'���U��+Z���s7����'�����y�YaF�6�����'� �j0hR�wJ����\�.˄z	�'mN������e�w��9%��1��^���Fx��I�	Ӑ��эޓ[r�I"���
@�XB䉧Uc�-a�#�3x���#���B�ɮX`q҄� v�\�B��ie�B�	�|j�c��Y'j�^(� g�5T��C��6T&\pU���p
�	y�C�I
����P��0U� lZ%�N!p����b��Mbyr��r`�c����#v�xD3���"j��J�	�����O>�$�O$���4)��q6Lς���i>��SjHL�����B6X��H�`f*����a��Aߌ��ōَ��L�#OJ4�4���;,��F�ͫ'��Qq��O��D$�ӌo ���R�>/,�)'̀�F��˓�0?9t
\��ab�I��8�`
zx���+O~��g㉖b4�3��^<{���]�pX��Z&�M���|����?�R�I�:���h ��4)���.�-�?)co�2M��9�dĺO��}�!���� �����3�D�huy��+�3Ox���Y�F8<��e)!vW΢"�h�-�!!�G����d��<������R~J~��O���i�(��| fb��_ՙ�"O�0�-ڡF8q� 4V3zhZ��I��ȟ���!��?]�X�����?B^H����O$�}�x�p���?���?Y/O�iW?x�) ���rl[��D"e�Eʴ�O�`@B�J�U�d�?#<9uL�ybp�e�&!�����J�c��I���v4��k��Ij�T���O&\�l��8d�Ɵ��T�򶟟��)�O��D9ړ�y�@=`��1�����.1[P)�6�y���,e4��(�U�Q�'�?���i>}�	Hy2��-i�<Ps2�	1g5�e�䆵"�0;p�'�B�')2^�b>͋0j��8�ܰz�h��7�^]�dO�z@�VB�4�Ƭq��X���<��KƆ�4�^"YK����Ń��dt#�G[�~x��vb���<�G[Ɵx��!�'E��R��3`�y�����F{���2sXM-5G��!t� 4OTY��"O4��s+y� $J+oev0	�_���ݴ�?�+O�� %��m�'[7L�AE�:%���բ �#*O��D�O���ʙd5�!RI���1��F�ޟ��	2`a`h�PB����o�p">���H�mLq� H/�*Y�,��0 ��$@^dl#���K..=��������O$b>�I%��&���8F�DtQ���<��gǦy���O�.��$ ��e����I����/��pR�jD>���KԊ�W���3^r���OB˓���O@��-�\���k��R�F���	���'>�|I�&Rf ة𲯑���S'y�!3��~��l� ��	ܨ�Ʉ�r��ĉD�
��SK�~�OMzD*U*�m��H�1��,C6��'�4�����?Y�O�OZ�)� @�� 㚃S��4�r�
�:U(��"Ot��W�T96:L0�a�	<
�#�I��ȟ�Ț�D8��9����)�<:E�J&��⟨�3�`�.I�
�A�԰$��!(C�I��(!�&)v��H�)$\0C��/>圬 ���i�D�LC�	�,������3����i� �>C�.U��[�*��Gv�9�� P:dB�	6n�����]�$Z���]�9*�d7F��~�
�8�8p#���%zl-���$�y� ��"(B�:��E#d�,��T�J?�y�∃^X���C��쉺��S��yr;Q�䃕��#sN�͙�����y2�Мq;�h� Hѵh��@�dS��y���V��M롬��m@� ����y��ψ2d�Z���9`f�MBG*O3�y
��A�R�q�N^Oێ`s6BХ�y�)]�
� ��YE4����y��E>%�2rL�{s��b��/�yB"���=rEɆ�:�)�N����O�d*���P��$,�<0a�JZ��B�ɣ)#HZ�����	 &Ļ)�⟐x'�>�D-�.-����A���g傻EA��!���;E��S��'�t=�'(�4S�h�3����I$a ��'1���)��I3Ӳ�'��>�M�<;	����đm'̘��eS��I�~r�s�x�&J�nU I�	�!Z>@��d��l���'�N�'q�Q�K�X�����3��JJApUG�i��a��'n~(XK�H{ӎ'�'5�Jm�k˨V��Cs;vV=�����p�O�OP�>ᔴiRH�.���`ӀF�fL"q`)O.\��>���S;
n�3�;O��@j�L�)6�vx��'��}RJ���<�Es~b��|h��lަc�l��+�d�ͤO@�"A����5�޺�m�<J.�U�W,6H����~	Ψ���?�,_n�	#!�8����K$hM\-a��Go*�$S���?��l"N��۔'>�%B$�\C�<	��4$�:H1���0���	2����Q�'��'����'�Zc�Aq�Ƣ>�̠���O�6KH��O���O���O���<%>�A$N	-�����a��`�Q�(��,�S�'q@��֋܁7h$�wI��{�T��~P�ɡcX�h�pD[����f�d�ȓ8�v|�sa��L�s�B� ,���ȓ(�80+w�T��0��#TG����p�"AH&d�0v��jG"Q�n����Cm(��$iα&IF�BQ�P���ȓFJ����̚�= �@��� ��ȓF)X�ӳE�"-��aUfFS�$�ȓ7��eP�:�������@L��g?ظ�j� f����R �����	�l���W�JP`� \�
B���ȓ9s�H�J;.n~H� ��Y����?��4Zu��٢�pR¼��c��F=C�͚'9�4q�$˒) ��X����qU!I-_�\yB�8e��թbImaz�01"ƈ`�02�W� �,a0�'D*0�f��l��ԪІ:���+g��;`���@�8F������ Jt�l�Ek�$ v�x�w�|2��hw�Yص(�+&Hi���y�� X�A��o΋d�8�Î�yr�\.p�*ͫ�E��a��=�c��y� �@})��!#��|�h�ya^X ��gc@"!P<iC ��yR&Ҥ[��ܨ��,$à�{�Ë�y�/\f��§I��f�@A͌��y����l80h�A�)~��Y!�
9�yRn������ӂG�԰p�O���y��*���Q�	2K`07�݆�y��Y0P)�ꧠ���$��yҥ�w�#����褰m���yRA�1� �c�͇{�t��J��y
� ~� �d�D�$��v,�8I*��"O\�$��"�KUj.]�*�+"Ob*U�&	 IkT�[�C�,"�"O
u�0�W,N&|c��v�%ѳ"O�T���+b����Y���8�"On��j�MDH�/Ȳ"O� ( GY.I�f탠��*�*8"�"OF�z�̓0ഒVL@0*���"OICjZ�vjn�XA�z���"Ob�c@!@Dz�)'k��$�h!p�"O�E#� nr� 
�n�5+�"O��r�ku_L YpH�$`^�9�"O(uP��
jy��+u�ԤB��qq"O�p�R`�-pD�0�T��b9	�"O��6D���`TӇ���V�(+�"OVHb4��:k.�@S�\r���"O��ZW��.����a�� �깋 "O�(��c��tTn�BתZ�A��;�"O��7/MR��̀�OX�f��\�"O���4`'B�x+`��P��Ⱥ�"O|�W� 1�%p��%;: c"O6!1q��V���P��-/��V"O����!ɔ�8��XdH&���"O�}�L�W�i����&�JLxu"O֔ڕ��25j�-��N��?���0�"O�5�B��wy$�x�nI�L?
$!P"O$H��d� +�l��MA�-,��"O��h!n���E��8`&n��"O<�*���'�Z�4J�-��[�"Oy�&�W�B$Zb��-k�Ɂ�"O\�����o��d�b�3NQz�"O�}q� ;=h�I�OB3�g"O~��)��H��$Kv��*(�ٸ"O  K�A�`�貇	ֽT(=�"OЙq2�(Z�}���K�,�Qw"O��b����M�ᏘmҴ��e"O�%Yǩ�"�*M� n	T1vՃ�"Ov(�B�O� �f�&�ܽ ��]�G"O��%;x����TZ�0��"O���v�N`����'9T_$�3�"O� A�LW6Ĳ�qG�H�P$���"OJ	9�F =6T�P�&�)��Q؇"O���al����i��T���ٕ"O���7c�%sn-K��<��v"O��)��4|��z!�Y�v�@)"OP�A0`�p�v�P�F�5Q	Le�Q"O��h��Xvt��GΏc  Ɂ�"O�e[���I�R�R5�ȑ��x�"O荙���1+u`q�cK�o��Ĳ�"O�)Ң�W�R(���S���6"OP�Y���Z��e(�D-2�&���"Ot�PB�X<}�����h��v6R,B�"O����gȪ$~1���H�+��r�"O\t�q���.��n�?�J�C"O`��	rd�%D���d���"OΠi�� �`t*�䏮,mF�b"O�-����I�LP��_z8J-hA"O`G�F����@�*�|`"O�ٰAhE1H:2��D@X(*	�8yg"O �3cIG
-�r�Y�Q�(\��"O0����H�S����!�BДx�2"O�( �C-�����.'8��"O�T���Y aXx7M�F�d+'"O.	+T��>@�P����A���"O� 2 �Ŏ�]ט�:�m�'_�J�	�"O�	��0
�pE��z���1"O@9��b,O)�T��D�R�Ъ�"O�e	r�̦ k�0a��R��V"O�X�G��FX��'5BX4"OD�i��p�%�&�D^O` qV"O�	�RD�LҎ�!�l��O8b��6"O`�cr��"&����,	0"!�4!�"OL�!�ފP�:��1k�!U2`���"Of�(��1qkR��$@�62xi�"O�e1��D �3�M�!?-�	�f"O���qB00�M����X����"O������Pp3�+Ԡ#d�$Y�"O=q��7<��{�l��SV3�"O�%�A9)(ʂ�F|u��"Ol]3�k֜����� @�6���
 "OzTCR�6j�-YfO� �1�"O����o��'�|��r���
�ڽq"O�a���N'cOX��d�&NՂ���"OF4���(����ɀ,Έ���"OT�	`��� �-;whV��D�"OX1���a��]��������� "O �+f� ]�4���I�+���"Or����5rm��pR�Ûl2���c"O��� !Ԕ�{��J��R"O�غ7��>����.�'qHЁ��"O���@ ��0�7��Vf���"Ov�H�닩mq<}vm��~���"O@Ō1Qtt�R�a�;U�d��G"O4����=_Ք@�EG����̙s"Op|�C�N/2j��'�2�xL� "O�)����QEt-Q�L�{���*q"O����'(3�4�چ�ѵ-��u��"Ox����"��D*pDѤ~��ۓ"O`�ӗ�Y�2u����4w�#�"O��i�K�g?"XAh�9}�Ȁ"O��%"��nf��DGroJ�U"Oi�}<�p��Ƅ|b��F"O�������#� |R��:B]��a�"O�]�F�!��͂�/;<Y��@A"Of��f���h!rp�0C/
�3a"O ��7�$3��U��6s6Q*3"OZ�5HZ�Zw"9�jɏ1��0�d"Ot �CmT P��`��A#
��	��"O �{g��&o�T%�d �o�]�"O(�� [�ٙ&#
 ���"Or�0K��"��Y GB�,�X@��"O�lZ��Xl��1k�q$x���"Oj�
�i[-k�"���KW �,��"OV�֠V�E�.�AӍ[,{$͓�"O����*˪+�NiK�̀���i��"O(D)�ҋL�$t�3,�
��i2�"Oڱ�e�����3FE���c"O��pF遤X�P�tdK,
)$��"O���Sj�?T�������|8F"O���F�?"4�B+��Q�!X�"O�1�ʁ�b�8ax��
�@�|���"O����kZ:9p��8v�&\�J@��"O����ն_G�ũB�K�$P"�"OН�э�!2LS�o�:_�8�7"O�L�C�*{`XC��������"O���ӣ��Ȑ��Oܬ_�@�ٔ"O��S��X345���	�u����"O�l�iձm��b��˦Fb���"O� �YAF
@�i��,ɼ!d�%Zu"O��iPɕ� q�L`���)w1�=sc"O⨣1��7�a�,�
8,t)3"O���J���n(1*��`!�(Hq"Orl��G e���0���9	�@X�"O�Ao��,�d�'P�e�(0"O�"�LL�w��Ȉc���Z�p"OB� ��i��ܫc5��$1"O��ꡀ��y�b�����z).�k�"Oz�``��{���(V��%�PRU"O֙���E#c�bъ�`gT,�2"O*�3eF:0�֌�G(�J7e$D�tvÉ8m�6���Jڧ
�܁��%D��S��C'.���r�C� 2�ٰ�9D�ĊQW��b���@ܘ%4��1�"D��Y���	^:�{���# 1t)1� D�� Lȟ_���)�ՠ���� =D���'�����;��)@�e.D��x6�": �s"AS.r��%��'"D�X2a��h��vL�']Ѭ�BP�!D�8�"��_j�,qvi�bB� � �,D��Ȑ�#0��,cD�� 5~���c+D����W6s ]�1,�1	��*D���CE^UҘ�e�;M���&D���P�*Nw�mI�&�<ה����8D�\"D�M�~�ZT�Ԫ��=�k!�,D��d�ͯ5���`�!uQg(,D����TVب4�'�~���ঠ(D��	3+�L&�)b`?p8�Iz��&D��#F��<�� 5�
u<x���6D�(�!�0�l0g�ْn�Z�36A3D�����1/:D ��W�8T1�J<D�DrjX Mݒ�0���;dp0�7D��y�KGs�X�pl\�t6JțC�9D�x� ,�&U�����"=��0*D�d�B��4�� ӑWv�Ur��:D��4X����&%A$��o#D��邷5�D,��I��ģt�?D���䮃sv�$A�鍐�ڜ1RO(D� �wO��a���u�;cᔩ�D�$D�,s��#H�I����ǅ6�9�ȓ%����Z���D��'��)x�':"�	6��"+]rA�̓�	<�i��',TmQV�#9+̨�u�f��	�'�lYsA��=n}�ɠƌتg�p�+�'��	���3;&�X낟]�N)��' l�s�-y(
iPw@�[�
���'q���-*`邸�mM>Z��1z�'L�X��ÄL��yaB�c_�0�'���2®�E3�@�T�����') ���O�/�����y6\@�'c0I�DH
��5�^k2�s�'L��o�9eKT�2��,[��@�<���.6L<3B��8\?欪`�A{�<�7��j}�4뀫���20E(�p�<ѓ��^��ꑥٯ.��K�!�p�<�t酐i�r՚��ڬ.�B�BU�.���C��koLb���$\��m%��B@���(4"9��X���=D�hj���_��IQO� lQ�l�d<D����B��-R���D�cc �b�C<D����2C�&��,^-�r�n;D���&�/a�(�*�n�T���h0�5D� S���!|������\"!#�5D��	�-Ze �`!�����b�	4D�� ���ɂ�i�H�8ҍ�vZ�l�"O�b&�2~TBH�į$gR��y�"O
�{�%�'���Ir�6P���3"O��[7���X	l ��?n)�+�"O�T+��2\�@8P�W� (�T"O2y�偢,\0��щ�!bi�"O�*�L4
��Zg+ɳU
)E"O$�%T%����i��<�I"O4P�փ L~��Oճ �<a�P"O��X�ɑ�n檬O_ ��B�"O�D����R��b��U��ȫ�"O���Ua�U���G�}�D�(F"O"hPiE�5�(@ ����l`�"O��f��1wF��:��F�Ǡ�JT"O`�J�fD�"�&Ap�LY*�X{0"O�=�U��:I�d�;"�G�~�0�"O���eJS<u%B!�����
�a�"O^U;6c���D�� 6�Yg"O0d�Z�đ!Ĉ\����Ď��!��-zS�H�Zh�!��G�!�ě!v$ٱ��=C b�����)�!�$�#3�����.ر�ʘH�!�dܓY6v�0�.Q�lx ��	�Fw!��&5b�(� F�;���j�敇�!�E	t6�)2 ɀn�רY�*>!���#r�0�+�Cҫ8m"�P��cW!�Ć1l8�����*!z��8�D�w�!�$K�|\�d�BFb����ɫ+�!�W�v'a���]�7i];�ʡZ
!�$D�bY����R:!c0��v���((!����@��]fl��e�R<!� �<���jV���q��TP��J�Pe!��X^0���BQXQF�Y��/QO!�$�	���R3���'��ɩ)�-!�dٳJ�Ơ��x�h�Fjʁw�!�d�(��@�biR�.�.z�/�^�!�ՉJZ����a	�z��/�=!��J5���p�M�%�M��G�%!�d�<&ݖ�)��c��K�
Q!���r��f�F�o�Z�T�S� n!���2x�(P+�͟.(�����Q�!���)pc���s�,�~�QD[�\}!�ĐQ�v�鲍�;*㢙X��Q�1o!�$^7j��1`��2F���aW��V!��Oj�X�筙�h9dmz�g��!�Ցu,�#QB�"EѦLC��\�R!�$U�FE�� Y#w��q�Ĥ$N�!���B~I1d�=3�]H�*	B!�䉓O�$� e"�e�%���_�0�!�ě0�j�SDP5hz<���eJ�!���3!v{ť� Q�,uK�(X�!�$5&] B

&cQ̨ؤ"�L�!�$"-T2բ` ��v�)r�H�T!��~���4��a!n�
��O�	!�D��Wd��K�"m����_��!�	�p�@pkl��j �Ua(m^!�D�	���@��b0Hc�gG)Z!�d��i��
��ñVy�1#�غaQ!�$��f�p���Їt�����S6h!��H���	� t��5A��N#P!�G�~��0K�?t�pȠ���)�!���o�<UЧ��
,�6�e�B�u�!��u-�E���W&x��}���ӕ	�!�dL��i1�b�xО阷��e�!�� ��HC"z�Ld�F�7ow��P"O����+\+B������W�~X��)�"O������A����"�/p@�1+�"O���䝘=XM���W���혅"O�Ջ4A۟R�}Qf\�\ʪĊA"O23��B�44�9��s�z9��"O� ���ا@��鳆��.8��"Ove�cn�VG��v5�:tc�"O� �a�G�4�i��K� ��]s�"O�I��b��P��P�U倸˄yy"O�}ԦlSbE@%�8$�<���"OV�xөF��rdG�{�Ơq�"O�	;�M�Q-���C�ǩ~�~���"O�@*P�U�� �HS� }PE"O�i� .��HNH� ��T��D��"O�ra�E�Rb��X�mT�VH�X�"O�B� ��+���Gb�#7�V�@"Oh��G��6��y;5R�-�<�"O�����
%]�tJ����j��R$"O�G���d1P!@�,A�X��"O,�p@d͢oLL��d $o��t A"OJqG��v����F�
���1"O�8�		5�l�#�U�.�����"Or�q�29�i0EhK6=�"O��+��M�-�>���/�x�@�t"O�iW햙F�y��Y���"Oj,��#����s��5��U�c"O.����7k(�L�>-,X�"O�,j�� $�l�tI;M7
�q�"O���ªB�+i@��T�I�1�de"OzU�F�ؓk2�id�P� �ms�"O0A��Ʌ�JTnX�@ȏQ�\��"O���ポ-�Z��V'�$gn�`8@"O| �2Ն��mʄ��>�Q�"O��qXX!p0*
2H8����"O��(V�ڗ΀|���&m7>,�r"O�)�c*τv��u�@�L��Q"T"O�Cs�^�5Tj`���ӽ|���4"OȠ�L��L���	>Ez��"O�h9&H�uä8+)O
��I�"Od]:��ے:5�,	��^�W! "O0H����KG�����+a��"O���uF!L��f�J0�l҄"O�Y���OF����FB^Ȯh*T"O�ʴ"D�H�8ABt��a3v�s�"O�%��*e_u��_�g���"O�����	%A)�)kp��%l��q2!"O��""��6��m���*3Z �"O��[pD�*/v�Yժ	��^��V"OL�c�%�+�v��4'�*L�ʈ�"O6]�n���E�%��,m0�r"O�Q�F�K�IG�؉���#=U�R�"ONA�J'\ݚ��C� '�z��u"O�T�� ǿZ@<�����<=��B�"O^aHT*6�l��ߊ,���*�"O��
$�ȷL�&��V���@�v�1�"O�H
��4��If.0O���"O��4�Щav~�Ҡ�M0!��Er6"O>�����Z����)8s�f,S�"OfњD�rB��j��l,�"O��r�!~]�@�#Ã�$�b"O�P�M��wh �R�~�>�:1"O(q��l`bd����eB�p"O8s����V֌_arC5"O� �IS�FۤU�X=�EN��'T4á"O�d� �+z�X#�GSO��=�`"OF���	��*(��¢�M�l�δQ�"O>�k��3O��ً%�2}�X��c"OԄʤ��n'���b+����U)�"O�)�� N�6)�
�5E����"O"� !�����)��2-�X�6"O�ð���lY�	+	��k��d"O�1�elF0ۨDHA�gx��J�"ONY�
wOfP0��K6v*Ł!"OhD !k�/�,�V��<lb8�q"O>��vKO#qu 4U�eQ�T��"OT��F �'=�pu�f͐=�l�T"Op����d.��	�F#��;0"O�AvD�D��H��FHH "O��֎U�3̊�*��WR�9��"O:<q7��UI��
ݿ���؃"O&A��
G�LM�]�#i*�*xq6"O�e�C�ќZ��1�-�9�����"OrK�,;P,��#P1#�����"O��!�@�~������L���"OR�����MUz���R�l�B`S&"O�X��͇
uj>�Cv
ΐL�( ��"O�D)�'W?2!�(B�(U�Z���T"O�A��n�0|��}kd� 5DuQ�"O����$�Q?x��	C=E��3"O�}�e���%����,�f"OX�iV�k*0}����X�~R�"O��k�-�
bC��QA2�fUaf"O8��7��;hw����P��iJF"Ob��μ��%e�D����"O��&g�	سM��b���:f"O^8E��2>R�b�q�X���"OέاBC<>"�bJۼ�n��"O�[��5I*Q�A$k8��;3"OL���&Y������D�1�.�J"O�)��e���A��<(zQ)t"OBI�C�ȭͺ���A9]|�� "Ot�#4��fÔ���.�,y�JhHs"O �Q�X�iB0�󣆇A����""O�%�E	5Ԛ$�tDה@��2"O��XӉ	�J��jpi	C���P�"O�c �Љ,��Q�7.ٗ-��� D"O�$i��%>�b�O�%����"Ot�b�5!���� ��)�F�c!"Oz�#� ��Y���;��T�:<,)S�"OQ� ��G�Τ
g�gS&���"OҬ��$��FzЗ�J��J"ORd�g)�M}�����(c��ܓ�"Oi�u��Ir��6�W:	��݊�"O�9�amZ5\��!�5��Z "O\(��.�eg@A�c.�"wP���"O�I:6�ŏv�
d�[�Z ����"O8��=S
��N�`^�<��"O���K>R��Q� /�3D���D"O�́2�;к�Y�`��8�"ON8�S"MLh�q�`�3<�P�"O�	� HǦ,���"�]"5�T2�"O��@\I:�q;j��KF(�{q"O�UWd��ΘB�	��Pa*ᨁ"O����'u���G\+�yQ��$��5�<(���8��B����'��� �>SW@�zA��YfLj�'T �P UM<����_pT��'�<�p4�Ό!'dy��!"i#��I��� �<
�ؽKܼ��b�ډ�N-�"OX��w"W$Բ�2���c��x��"O~P)u,@�9P�T��̛�"O�ɩՃ��Ql�9RbLLk����"O���V��Q&� �U�ΊIL��!"O4  ͨG�\�Z��89j��q"O܈�b券Tv�RU��?�	:6"O�b6M��S6�� ��]/I�P���"O�ġ�EM�C@���&ܭ�,9�r"O}��-M�2ON�SÊG��S"OT9+эҡά���#x��]�7"O$��@(� U��X28K�Fк�"OH�s��	�h��
^�W����"O@]PR�
�,R
�cu��r�P���H�<�f�];+~|$�(E�0�h�2�i�<�/�:0f�ѐ����+�n�i�<�Ǔ+4"�$X��ۘB�(�5%�b�<q�L͌yT8�2�C�F��X���^�<ɧ�ˬ��̻���(:\e��Q�<��ܓy f$P1��;�V0X�ONP�<�ef�l(���8f�.���I�<�wi?(]:���ڱ!I����H�<�7f�?�4�o_-0U��dT|�<Y�/�p*��k�d�,*�,%�7��s�<�m� wg�C ��%��5�\i�<q1eG�i���P��'9vl�Y'CK�<��d�6�z7F�P���E�<I��@�H�8�"@�'�����{�<QfW�>��̛�/�&U/���'� N�<9��*c��)��9^&� �@E�<�V���7�,Ủ�I5��8(�]i�<�5k�9̎y��҆mQ�)R�P�<�U�9$�
����F��\���JN�<�bGǢj�Nyp��J�i�����d�<�p�Y.^n�-�sb	�Z���fC_�<�N�J�T�����?���נ�`�<	" "�:ŋ��
�oK�zSF�Z�<ф)��T�Ƽ���@�M��C�N�<��*Թ1�����H��	���L�<1�BŜ7X%�����,k  _~�<Q�ٛ$_� 	�\����q%Qe�<)�Ƈ�W�̃��
�hQ8�(�X�<�c��V�@;ҏ�>j��a#��W�<�2͓!�(�g��7@Vd��KW�<�Tm�4#�z#A�54<�S�ʑV�<�2	^8\Q�fAJ�Tk�#���T�<!��	�o-ܼsb��q�8��p�UE�<rL�]��(0`�;S3���A��@�<9�JL;��e��7Kk��� �u�<�D�3e���p��	�\:{�� G�<1�FËOW~%S i�2 Bh���m�<�"��'�LR�@��s]�Y�%aMc�<q'�_�y�t���H�.Wu�����c�<�����~ �%����3O
������b�<Yw��=C)5j�i_3[V� 胣�[�<I$-�#lF�!�R��a�TR��SL�<���=|�hyG#��W����XJ�<a��H�Zzh������*D�l � �I�<�抙)`L [& �#=0y`%J�|�<9�(�
�d��	�����sv�<a�צW&DR(�D����Gu�<IKب���5휍���Z�<9��#t�T�ꦡU1"D&��
�o�<AR���{z<��H����(��m�<� ��UOƄi
���C*��#6T��"O�h��֓c�Pq����7,�t�G"OnEg�D9/��"%��9&���"O���A�W}����q�;�"OPV�8L�ƬBu�X+kj9b7"OHx���[�6���@�ߣa���"O����p�(yq3
м=��px�"OV����<&��),�_��\��"O2�)F�^K:ys�ɷgǊiR�"O��Q�H��4�,1a�j��M�L�`"O	�!!5�@���@�[���Z�"Ohx�T��Ap�Qz���B�"Ox0hJ�~��$I�	B�<]���B"O�P��H� &��3���l�=iB"O\10��ٮl|��q&eͳo���j�"O ���.�	�����cF�`�lqP"O������Z����`SA,"O<� �;r�S�d%(|���"O���P�\�����޷��Z`"O�j$E�6�b�IƵT�l!%"O(ECu�S�݊���c��I�"ON0�FK�Z��x��j��E��d�"O꘰&-ګu�6���$��?��`S"O2-�T���$�>�7�ڱS��)�"ON�q���_4d�A m�Ny$)!"O�a�Z��)��M�YLx9���y�-��҉���ā~#���bJX��y�嚺{H���7��#-�¤ꐩ&�y"	
���I���_0�!�a���y��
�&�����!x�)#��H4�y�KӆL�$`C�\3&&2ҥ�y� 2�@:��=�����ņ��y�eM:jiz��[$�VD��@N�y�bGt�\5�C˃NT�����/�y��m%l����½>��9�0%���y� ��P�ڌ�U�0�0:�Ċ7�y��7�� ���ʆ*&N��m��y��_���qR 6�[��ʉ�yb�.W吙�� �E&����yR�;hB�Qm�1�"-��F��yr+�i��i�Q�Q�7/���؅�y������?\jl�$�(�y-ʃ0��IWGD>U'z���#J��yrm�*A-��(�!��;�H
s�+�yB ��n��i�k�8(�Hr)�	�yB�(?O�J�IO�_Eڐi���y"�^?$��,:��*G'�сv� �y/ �D���J��F�u륁@
�y��oU��%J�>S�(���%�y�+�*`�<H�eȰ=�"��3#	�y"������)� � �����y"ËJ	H��[�i�5ц����y�k�	V���Y�4��Kľ�0<����آ�C��>}QՋ��q�!�D��f>��R!�WGj����|�!�[7%��z�/N*[Nٕ�ƺ>�!���,?(U���	�q�� Q�_;�!�DDtNЫ �&�H D�؂9 !�̏Fjp���*�6@@Vl�h!��
�Y*��i�B��	j�X�"�!�D� `D@
"��)@���ԫD~P!��A0>��Qh�i[�S�>��i9E�!�D�&r��):� �}��M	���!@V!��&���s�=diҌ`Ņխ|B!�� .�
�͊�e�2H[���*M�,��"O���U*�!2H����?�0"O>u�t�ܵq��1	:��"O��!�B�V V�Ybf�D�,�c"O"������53�$�q���R"O�l{B�B�mx������
&��y�"O<}���.'|@�"�	5f�"p"OZ]�&O^2F�,�B� .Fߌ�x�"OV9�UHK:b"D0��S���KU"OR�x�oRT8<�Ul�T���i�"O��Z�ʍ�%�=B੗�cM�d�"OpՉ���Z���J*=��"O<9�ǅ�`P�1��ԅ�d��"O"t�'�ZAX�і(X��9��"O\�#�� %P5wh 51%�4qp"OD�i!�O(:H��3Ǜ3?�0�T"OTy����� �T��eޙ0�`�J`"O���0!��k�u���t�6)��"O�����x����OЇ�5ٳ"Of����Z�#��E�dOXT1"O��r/��fЀ�ѶI 5��y
"OV��l�"=�Xe��43��#3"Od ��Ψ�6 �3�""����"Oh�%(^�n2Δ�QG�3~�L��"O��Qf��F�D�%��#]��)7"OXai҃U�V��  �F�H��� Q"O����lI+m.<34��Z�@`�"O����ȃy��R'`_d��9"O�%1�n��1��=;& ߥP�e��"ObM���ߚ���N�-dBN�a�"O���w��jҍ��%��{V"O�����;T ����6OvZ��"OP����>?�Q���fL~@JC"O�qx���Lɘ
^�$�A	"Ov���d]�4K>�0�	�,H�q"O��Z@G�l%a�ۄ:lQp"O,�↩�6�x�aJ�	s6dl "O����	_�A���s�K�/�`�"O��Rfc�W7�|id@�8e5{�"O��{p˚!i>�2��9)ލ�!"OB�rpd��]}za��P$i(��8�"OƄ[cOU����;R��"6� �"OE�r���[��2�G4K��"�"O�亥-Ȇy��+��Y���"O~a��<|
��3�B�z��M�"OT�����N�� R�	�V�p���"O�y���� v�Kc(�
�&	 �"O^�I�--NHS�F~�0=1"O"�	���8=����(�H�K4"O�a`��Ø�F�I0$q�0�e"O*���"'2%�����!�.�*�"O�}�v�(E ��.�8EQ�"O8�"B�9p%�8F�	6��lj�"O�A� bY0vH�T:rdҎzzz,��"Of�Ce��^x�:6��KQ찘v"Oh��ƆG-Mό<$��-C�m��"O$�c#ÜGa��"#T�R��"O�y�d�P�x�4<q"���p���y�"O6�g솧~,X35�;y�ԕz�"O�Q��E�T�!4�@bv�D#q"O~��å��g(|$1蔾�4��"O(hq Cl1nH�� : �Rxk�"O�CT�@9V�|}��4(}Q"O<����Z�ugB�hVL#l��@E"O� `���Nåko�QW�$i�`D(�"O���#8�R݃d������1"O����)�$̪���%Z���f"Ov��%�=*Qv=�ΦN�^40�"Ou����
j�$�dIY�|�b"O�l���(��w珡gE���"O�-�V%^�0�H=@��
5X<�d"OX��W�I ~eB@�#T2A�,��D"O($v̜�{�N�a�a�:sڸq�"O���H^)-f�[C@A�?T����"O�A�czoj��JS�Q(��&"OU��[X�|�f�V3ҝ�4"O��)�Q�<�5��"m#�D{�"O\<�#+ɲ4#8���!=�A�"OP�֥��lz���⥚ gƌl6D�,"5B�	�z�0�fM�p�D�`
)D�Pv���u���"��;���GE#D�<�a��5DlT1c��� -��Ie5D�`[���fPX���BZ�t��3�-D�D�7`��?�p�A4��)
�T�c0D�0idKؠ+F\��.Qp����/D�`z�hZ#- �T��;
,�A@%;D�����
x@P�iX�oW�X	�9D�lHw"�>����W$�x��I8D��� �F�,q6�@��Q�/z�\ۓ'!D�H�hD����a�Ŝ(ٶ � � D�0��*V��� ���#K}|�"�8D�����Z�1Q-�:5Tl�D$D�����u&���I��|i3�=D�<@����q����̓z!�=p�,=D������m`^�8�i�|��a�!:D���`EB"C�{��P�Dgxt��9D��R�DH*�(U��α
�f���!D�tx�)/Kʀk�$�52�dH�"=D�0v�/[5̵ku�ĥU�B���,9D���o��m��1�#)B,60�g�4D��a��,����6�\�C�(D���ҶW���*���>���Qb)D�P�ǂ�AK6	�c
�y�l��h(D�8EH[�d���F�tDTr@'D�ܠ1�K�`l�ł�/8Ay`ef1D�\�q�>(@QoB�����3D��5��%�����:"`1��	2D�t;�)��)��#B� +扫�#D�p��^����Rn͓@�t-�6�5D�8`�F �7[����M�XjM��4D�l;GK��z&�'M_QH�� n1D�(�jY�~i�hx") B�I�$*D� ������&���{V3D�43@��l�r��V�RR�x��1D�@0��{�8H��ґe��
�"D���3�C�B]2�2ЅP�]a$�+�%D����Xe�~5R�INh��1�/D���DG���e�f��6(��8+��/D�ș`e��4hȅ�2M��*�*���-D����H�$,N4���6PE�آ�-D���Ǉ%�l�b�? 1ц�,D���-��h����"ɕ,Lx���f�(D���֌�lZI���++�܅��*D��Qŏ��7A��0�_,Q� ���&D�l���D��)�7��Y{���?D�d�����)��[[���@��0D��q���D�)0L�!9�,�*-D��@��F���턞{ۄ(k�)D�� ,�aag�$y�`�Re`��]=bܛ"OtT�2���p��mؐ8"�"a"OJ	b�.�	i_�(�j�9b ����"OR��7�А]pX$J#�&b�ڜ��"O��C`�Ȃ
����Y�6��"O$d{����ac7dP�{]�8�"O2�#�\�h"�����~\:�QS"O���b!Нe�n5#D�&C�`�Y�"O����g	R� �5C��,�d�"O��g��A\��k�C�}��19�"O���s!ӳP����v#	B��R�"OҐ ���-	�
 0� X>rh�"O ɨł�[o�Mi�쌝 /�@"O�ْT�T�MN֔�O'
h�jd"O�y[A�Z6kp�1�Q*Dj*`��"O>Aj�!nu�b�'�>Vw�A)�"O��P�\�},ܛ��?����u"O.%P�
�/U`)����|n�z�"O��!��M�tzTD- IƵcc"O4x )D�4�i{D$�)G=�"Ot@Q�� Ȟ�bW��"1[@�Q"O:���P�N*zQY�V" ?e�"O&��#�>$��Hr� �\�j�z�"O���SD
4!��� �>TQv"O(��Dc��ow�A:�I#��)JA"O,� �fI�]�Q�7j��"�氻 "O<�0��g@�YkG��	��UC�"OZ�iC���NP
CG(\�\u�"O^̨���)w��@�!�@����"O�����)C�ʟ��0��"O�41�o]>`�TU����$ a�x0�"ON�X��C?�pU�!)��!Dz]�"Op�z%lE<�!�Y+�$q""O�qhւ
Gh0�'
ړ)��B"O�: �o�"`(Ol
�iR�"O<P���/�4QVbǴ	�Y#"O�͋� ��<�n�y���lր��p"O��	f���i2��*:4$�I"O����	ܵK,�S&Hh�"O�@!�T�^��� �
E#X%���2"OP����U<m�H��I�� Raa"OT]�V+�o��sd�H�is�u��"O�ܙUoC�!�)�b	ѩseB���"O���T�]�<@\lz�Ú6*��;b"O��{pl�0]ހy2,J4,̰ "O8A���7x�ȱ�D�{�~2a"O�L�Vd��E�� "U�%���q"O�5�bA�#�y� �V�H��f"Oސ��̛'D�.ajr/ے�l�s"O|��g��5}���N>����`"O���Cˤ7o�����؊U���"O&I�%�����q!ֺV�.qE"O����ρ��Uc�b�}��DC�"OF�bE�ԡ ;@A�%.`JI#�"OD��Њ�<��L@"�Q�A�,[�"O}��}��H��)VV�h��e"Of
p�M�3��Iq�j����"O�m���{��������b�"O�hSg
�h�e�jEz]�Y�p"OF<e����%@G���@U�pA0"O��ڻQԈ�㧅�y�.���"O�d�%�On�@Ĩ���7��=��"O8$"aO��j��cnܣK�*Q�c"O����H=��T)G�.er�j�"O� <}I ��A�j@ �MCfZpq{"OR��k�V�C��3Ei Т"O�|�c甐A5d�fJ]�BX�'"O��0�cD�v;��Ɔ�����hW"O�as Ȯr<|b�O�{u�,��"Ol�SG��5�D!ӄW�_��|YP"O���$��.
\،���_��)�"O���㖾beR�S"�H��0��"O��1hH�y�����AQ�)�:���"O\(�H��c�9�w!��w��Y9�"O~�.�R�r��rA��`�Vݒ"OB�*fg5P[J����Ͽ#�T���"O�@X��cm��r��.@�
���"O��z抝+�=0҄�i{T��"O�̱1ꕝ)�H&�;*yB�e"Ol�aJ˕B�Au�ٚ�6d�!"O@�
t(I&0��`��်u��{�"O*�)E�Sh�*颇��(%_ր!"O.�Z��O?f+(�jI�M����"OX�� ��&��-S��U
���"O�|���(?�J�{ J���"OhВ�͟�b�B���IA�v�4��"OjPA���`t��h�1W�-(&"O6�z��-cS0 ��j˧9:�J�"O�ĳc��+p��"��n|���g"O�"`o�ﾴ�"/V�z���"O
	��k�1��K&l��`n:m��"OpLЄ	�M���5- 6a.  x�"O@i�#G[5X���p��z��"O�p��M���O�-v�,�+d"O����+�(ȩW,ѧ"��L�""O����Q>s�n��R�۵X�*D�$"O* �@�?V��Չ��E�\����"O�:!��+�b`���$(�.���"O�+e�	�
y�lᒎ͏}���"O�y�B(E�T�n��OgR��"O
y��^�(i��!!V�u�E"O�xqĦ�kX�%���ڑZL.��"O�qX���8t�=!��P%s'eJV"O��h-�GW ��T�*�R�"O���V����I\ 6 �E�"ON�*��+7������$���4"O, 
���J�J-0 �Y}bjd"Oeq6��s��tI�C�fz� ��"O6�2"
��I�� �qÂ�~c.���"O���
i��I�a��/xG�`څ"O�}���O�!����D���Ȗ*O��VH��"V	�L� 6�T��'�v�J��Y?P>(@�ߦ�2"O�� �Λp#�I; �6"�Q"OQ�Ug�ݶ�0�O�(�@B�"O�ȅ�U.�� �V4+�*-��"O�`z�oɀiY�+j�9@�U:�"O$��Pk�+�ڱ)��E'0��Aa!"O��s���6N��C���%s���g"O���P̏�����ox
a��"O�ph���al�h���4_k�8�d"O�%B��I1N���M^h�x�"O,�z2���R�ްf��,>`l���"O����ĄC���`��;"�`x�"O
}ɒ��%�@S�M�"�"Ot�R�f�24��cg���@�A�"O<�B-2r��Hi�׫R?`a��"O�i1�O�����!1#,��"O� �`qd�E�|�.��r�Ǣn��22"O�1a-F�>�&��l��=�j��V"O
 ���2^��Q�%e��	#%"O2�J͈R�2ݣ@*W�I�^*'"O�����(b�����5�ai��	�$��/�R̛��	�U�ze U���u��L���(f�Y�ѦWX���l�0 �*��(wF�L�`Xs�����P�sԈ��M.3N�L��F��W���*��ۚ)f��[@���)z�y�j�7������J��#FF.&#(X�'؟,�4��h�m�	�-�:����Y�M|�ܴX�4$�i� �p
u�	�$���'��O�i2ғf��l�B����8�Xr!�)�$���	:�M�U�i�����.#5�Y8���q%/��~�'C%?��6-�O���|�6��>�?����MÀ*��$��5Q�%֙Y�䠢c��2�Z;Qރb/bM��NN7�F�b�qܧ��]cU y$`Q�06�z���H����4N��R�;f�^�ȅN^� tX֝;�́�Z u;B������)F`u�¥�"&�=j�.�¦u2���OL��L�����R��M��>l<��[��'V*���OX���O�ʓ�?q�����v��{姗�@�rlIs(��(Om���MsJ>��Ϯ�uw��ȩ[��(�*A)2�*]g�ʓd�q*��$�?��?���NX�N�~bvÜ(M���%		6���"K�	]S!QbȚV:�(Y�����Haf�OLXDx��NF�L�BQ8!���	�o��'W&��'���sN�J�͒��0�3��\%r�.Xo�����@��'� ��C�D�p��>�6��ןx;ڴ.���'�i�����}Ԕ�� ��5-H��Cܓ�=�q��P��$��=~���q��7MUܦ�'����?��'(\t����
FҔxf!�����i	�A�@�'��'���O;
D���x:�Lͪ�`P�̽w�I�SB�  +F�H�b=)�z��	D��yQ�	:)���E"ޡ
�ޠ�FHA�G��)�"e���+��]�d��B��� ��� ְ	H>������k@��q����!�ʩH��[,V�,S�4�?9)O2�d<�i>oZ5`L���ƀ�88@�BT.U' �C�	�gCjI0���&ts�@ߛ���ɩ�M�'�i��I	D�jش�?iO|�w�s��x r��f$-��FϮ{O62�'�R�'ynP+B޺@�Z�)Q�T�]!ҩ�B�|��)oLԸ�A׵��� a\/�HO�U�R����|ˣIZ�l �Z7-dJD��=�H��~�����
,|o����*��J,|P�j�Ȕn����O�ŉ�c��B���d�N�� ��Of��SG�'*�dQa%F��i��P-Si6@�=����`Ӕ6�E/=
N� �[�g����ÝTv���c�Ro�Ο̗���#�<w)2�'ݛK�6�"M���
#�8��H��1��� �ެX�F0³΍��,�PlЅ��O�����8H1f�v~hTS��vb`��!�i�(8H�]�I0�, `,�a��ڦi�1��#8>���u��T)J�@̍�SB��2�̦�Y���Ov����I�IT��M���0M���*�ԭv$��"���A?a���,,OH��jNx�ҴgJ�]P*TZD�	ݦy��4��F��!�Xw��y��m����*�A#.��&�/�<lO:���  �   `   Ĵ���	��Z�ZvIJ(ʜ�cd�<������qe�H�4m��_;:<��iF�6�T�T�2Ts�V�Z *��4e/s:l���M&�i����W���DS8Jİ�B)���z��5'S~�As�̦N�Dl��{�i�X�'�4�m�,H�4X�*�"����!	>!;f�?Ǹ J��r��L�'�\\J��$j�l�'pHbVO�y�8sm
9%����C�æg�$�۴~�Eh�',��1O�_yB7�ĥ;�]>/�vq���VI�fhV�łw�v�P�W���dF�	RҹZ�DE;��D�3Wqd���ci>%���5�̴��I����@ໟ�3�hO�nPhb��	&�
8�1O� @C�X�)4�;����<OJA���dY��O�-K MD���I6� "��b���h�'���Fx�eRm}%�:h1�D�蝛���6��	6>w���6��1L�D���?�t�#$�!N��vTw�'9�|Ex.�/j|(�9J@���K��fR$Yَ}�Yk�'UB��'��3'�P??hF�[����df`"-O���D@���'ѠA:�e+P�Tcs.�������[�'m\�Dx¡M��<�g␗s�����oS
��� 2��&����T�xb�/Q��+^*������~���y�'��%����']\�1.X?0L�r��G�dH��c�I5B�R���GQ��5W��X�1%n>��K~%������+s���fn�<�f�".��%��1dF�:6�Onj��](��Q�h�(�$�ǻi�r��"ʓ.��#<��������cV��oX�4�4FLq�<Y 
 2  �s�����xӺ�$�O� Ĥ�Ks����'�����8�Ġ�A�Iz�#Ʈ�z��O����O�EQU�~�A=
��p,����rOЦe�'ъ���K`Ӏ�O���OE�4�����a������(i�<nZ�����#<���Ď�� ۼ����.R;y�R�Џ�M�!��7x�&�'���'��o/�ɷ �i;�'˥^�v3F�+�9�ߴP�րDx����O� s�ϐw�}�g�==lY�K����I������"�tɨO<����?�'��=�e���+����%r�}��6Θ'�b�'��xa����5��Y9p�Ķ-f�7��O��B�f�<a�^?��	j�	��T���ؐ0����%ɉu"��O��ؘ'K��'��V�4�TIW V�P$+S�
P   �	  �  (  �  �'  �/  �5  !<  }B  �H  O  \U  �[  �a  )h  jn  �t  �z  ��   `� u�	����Zv)C�'ll\�0"Ez+⟈m=�R��/{|@�D R�Д㍓QJXAA#fN�3�fIk�A(�n@�(�b�iukѬ6&�;6n.�z��4��p��$�$�Ǿg$��ȗ�*�H�:#%*H1�L�
�I���3H��V� �4�Ic)��E+GWذF`F�U� �)� �٘����~&d4��Nbܝ��B2u�%��49T������?���?���>N]1�-y݈13R͂>i��s��?�bǌ+��*O���F����O��dPN-��e�7T��pK!��wx�dݦ����O��Ę�1� ���+2<Or���7Cn]��A\�d0�`Q�	+iCn���f�S���sP,��4bi�JyXF�>������\�L,\��S!����_�I�0 EL�D}���?���?I���?����?�)�>��f'��ˤ������$
E6_������AJش<���Hy�`����	��4���"o�X��D�:y,��P`��
�a�WZ����ƓQ�Ͱ7d8Z�����[8e�V�"#�є$`���:o5�� �43k���g���I�|{��G����p��7R���B?<����#�q`�b
*I���s�g�R�bD���ş �?� f�9=3:$J/X&�X����?�?���0?�f,��@��8Y���;C��h���i�'���'�1��/<��vÈ}���H1�Ӣ��d6�S�Ot �F�ɐb2��#��3W&�䁕�'�ў���*H��{ڴ���
0X�	A����
1!�@�y�T���Iß�ϧh� b�k�`��<>��lZ>~~q�3� S-,T3�
 Ak~t��IIhF%[b�U " ����,!�N�d��B�H�XA�iR�;O�-���'�B��<��O�i/�T̈)!�j���OY�D�I���?�|j�'�X����_=a��P%��r�&\K����+T�4��\q��
4��y,�T�N7-7�	,F,!�?��'DN�@DlٓUoX,@�hH+pH���'��#gQ��1��-f頶�'aL!��Od����0R���
�'�>,x�V^�lC��K@=��'h�\ѷ�Ud����+P S�'��ir�9H�f�Т �(#�t Z��XBlDx���Ik~]��H�<u���8�ʒ�C�C䉂&�
{ӆNkp�@��4�B�	�'Lq�䏝�n͐��T$��B䉺 NlhH K^��l���B��xj@�ᥬ�L�T����`R�B�	�n)Q��86���COG�t\�0&-��I�z�)Qj\���-C��/*OB�	9��"���Y����Ϗ�B��C�Ɍf7�a	X�)����s��*��C�	�K@:���l��hرq�d��C�ɶW�.TC�
�	�F̻6��<j�����l�J�oZe~Qb\���R'����������?�.OZ���Oh���S�X@�C�)Q���B�ʟ�붎L���0#*Y�g �ː 3Oءg#�C�
4�s/�6���L�B	�ё$�X<y��@��+aax¬�$�?)��i�B6m�O���	˩���k���U�s��<������(��,�Ɍ%�^0�6��r�]��'�N��#H@�E:�	&qB��@ 	�^��|!ɰ��y���'_��z�`#vA�L�5�1<U!�$+"�>��!�
K�Ƅ��ɏ-�!�$�f�`-9A͏���X����8V:!�d ;�`5�7�X�@�&kǈ,�!�d�g�ޥ�D��8B��m�b�RNY��dU�[�>�NÀ^G��0GრP��|�l�=F��t�'���'��ɭT�%�5Z )چ)U/�,5zd���V&�|��|�2���C�?t�L�'��O��S��	0��l
qJ�,#.��+�!�<8	`*��)���Rb�~���4؊ �����s_�(��G*y4��:�%.>�<T0�49/�	1/	f�$'��O~�D�OD��A��"E������?�d��%o&<O"��?�B�x�*5���N�B�h�}y�Dw��ln�M�i>��Cyb!�&S�b��C,CEqz3�x�Q��*D0�6�'p��'��s��:Oڒ�"o��&����R�ԅ3�5�8� �^�H��|���S�>��7nP(Tm(�נA,2���ӫǺ]��� ��Kc��*�/��ܴ�;�(O8mc�(=MO��K���U����o�09y�no�ʓ�?���?9���?�ϟ2�X@AJ<x�.�z�i��R�~A�"O؜)b�8	L���G�O�rH��{P�|�rӒ��<AAj��<��6�?Ugƾh�Z��N�?H� $:Ox9!P�)� |HP(�]��Q�eO�\���'�X+���8]j�HŲI��!;�m���ax"G��?a��|^�	�l8QmM)=,�a'OG5�yR.Q�q�T����>���Z�j�!��?��'X"�2����0�@�Ƞg�Ƶ�O>�`Ϡc�v�|�V>��əa=��S`�D�6�"�Ѐ-5�j����y!�ObDQ2AH��[Sf�k�S�O��b@'�p��(��Z#\���O��('Á�u��w%3T�h�XԳ�M{m5Ɠn�0 ����f~B
��?�7�i"N"}�'l�|5�VEʘ4ф �����H����'��й�_A�(s�N\\)X���w�O������pz��E�$����t�i!�V��B�5�Mk���?y����.lxm�ɲzyc���V���%�ګ'�@�nZ�F/�Aۑ�L��d9�I�>��SfE5.h������5(Vؠ���A!\v����&N��S�!�3�I�N,ى�&մ#���q�C��D�ߦ��ɗ!=N\��H�gy2�'��d�R˰pP��uM�t�d^�l���4(!2���P_|�S̛b͜��M��ie�'�Ҥ�'���I�I�rA�dOÉϴ�ذ̏Lgb�@u/V�]��֟ �	hy����1L�z�ڦ%�Ri$8zd�\&A&,�ó^zz��8sH���(i��0a�2=}�a2�C%>�5��� 搅�PA��GT���D ���sjA�uB�v.�?v}�A�' 6��ʦ��?i���ɹ-�$�����Y��tV嗢D�!��>��q˰�
�%�D��E��8:�'�듫�B�)do�T��'�c�A��Y$B�2�Z�M
�?�.O�D�O$��P%$4b'��L�Dp2 �Ɵ�X��H�@���Y��M�&	�m9p�-O̩���b4q#�E ���3e��X�1nĨJ]�(Po_Sax����?!�����92ђ)��ߕP8�f-I="�'����� e��$��\������&������X`�O��-�J��Ĭרl�=�t*�O��t�H�k�T��'���O�yP
J�Vz4�{�U�\��3���O`�D�/6��e�VI� S@��b-�.�MG�ǮxI��RSk֓���������V�Y�F	�4�Yy��EM�O���2��v����V�o4N�B�O2`+f�'���Sןr��E���r�L�c��q�r+�P�<�'�N�'0���ꆫT(p����3��Dz�>��g���2��6E��;00�3�o�O}\��0�E��?y�I�(�	Hy� F�A��T!Y�)I�����T�]�YFg�y{\�䒁A'���4��=t�x����qjEK�g�7c��Y宋�I� ����>��27��$S�s 2��lM���C"��0�Rm�OH�d$���t96 ��7�i�', 5c��i��'-�P�7)�8z˖�+JX��(O�Gzʟ�ʓ7U&��̱T�����0r} ���?���?!�����)�	���1��ǋHt��j�8��iر��(�$����3!����ɖ#\v`D �0*�c���6����oQq$��rL�&|�%�牚p$��x���@W`�!���:���O��$'ړ�O>`�U+ �Qx�Ȉ�ʖW�p
D"Or��d�P�`��u�A�ř}��٠Ô|�j�>���%A�����5U�8<A�%T�Cm~lN<�y�f��*���Wo�.
�j��"P=�y�/��Md<Dx�B m�J�������y��� N�ֈۗ/�,y�p$� &�,�PyR�X� t��aQɸN�6��HT�<�+�5D�r1XE�ׯT�������Q�'��1��I�tt9rt(A���Ʉ�GZ!�o�*�����=z��Q����=!��I�O%p�IRjN�k�0���NۻP)!�$C�pa��JS�6!�F�R6!��`!Ĕ�*�,�"Uiu���!�d1	���򠮟��֝� �
���D��O?��	�W��
���lK*�ɥf�t�<1�Ֆ��YQp�F#��,�`Ii�<!��A4\wr<2b#�t�ڑ�]�<)u#���L�8F�R�\0l���U]�<�5�U�9�8��gV��m3��`�<ٶ��dN���BRE�ހ����[y��Բ�p>�d��5p�����͟Y�6|)�g�V�<� v5�E%�2S&��FU�N���"O>�RB
U�8���+%dQ�Zy+"OX5!ƌ�<$Ժd�Oh��P"O�5��(TZ��8R��4X����'�&�`�'�5Jg�B%O8Gȁ�/#,yS�'��3t �4�<�[�P:8�}��'}�� ��8�LY��k\?��Y��'tzб�&A�u���uG  �x|:�'��`��Ж+,\��X'w��Q��'ּ9C��8,�Mk��x� �8��G�1Q?a��A���z	�FO�>W�U`G�1D�@b5���Z&�b��c����0D�X3�h�*H�e0��\�Bf ����2D��j�`���u����&=����+0D��Xa�U,q+T �墙�L�y�0�"D������$��5q��8+��d��O⡳��)�'H.0:���*�Wc��0s���f D��K�j}���#�	7P%��k;D�lp�� p� �Ϧ`���;D��p��Ri�0�j@ M�A�y�8D�t2Ӧ�1�R5S�H�_e�]���7D�dqFF�R���#%'L�a���@[�Ʉ	pj����f0�9�E�e����N�s�!���~x@�hJ�v�S���
�!�ĝ�s�Мa�K��x&�ؾ�!�$5�AW@+_�$�aD��vP!��-��}80�[�'��Y ��Eh�}���~Rץ:�����P�-`��+��yr��K,�	����B��J��y� �1{v��W�e�dX�%���yr%��E� !A�.�%M�l{��Y��y�*V&�,9x���dd QO��yB�N�Vm�����0zG�Π�hO�|k���/��h��!E31���J���
�C�ɐ<��'
T�<R��Uh�-��B�=`K�M��D	3�ȃ�jDTC�	�FM~Uö"	�D�C3hد
�"C��+UT*�P�'ۙw��Y�P.W�d�C�O��a���A�f�F�#w����i��"~zp�t�Li����Gց��H�/�y��z)J���T��9��V",���9O��(� ������k=��G�dq�̗��J0��R/{�r\�ȓ�0�`��3-Z�ݩ'�[-I���ȓkq>+fe1��<Kclq�6��';���yXhQ�! L�u	惚0R�⩇�!�@\R4m_�/ Ɲz$�ҫ3�FQ�ȓm���PT�4:@�e�H����ȓk�� �@{���Fm�9Ex���h6ĉ*�N�Xv�pn9@���Ɇ?� �	�{f6�q��0"����#���@nB�I��9r�I]�v��Q&蓯%N�C�Io���� �j�,�K���z�rC�		
Ov�Q ���1��
��B�%�NC䉋B����sDR-Y��uD �+�B�I�N�!�A���!x&K�B@�.��=��A�x�Oʂ�BG�R�3<)[�Ȍ9}r H��'8��K�C+RQsŨӷ|�p�	�'�>�K�S��$jt�p���
�'S��� ي�P���K0`+6aB
�'��Uɑ'�5=p�Sv�ʠh�H
�'��dS��l� L�4�­��N���Fx��I̗�vu�wJ� "$@lP��y��C�I���e�kH�h��l��P�$C�)� \*WI�/\	����BRԎH��"O��3.�B��@���֙d1����"O6�P�*� %�|I K�\�4! "O��VmP"x���JǮ(W��|ڤU��q�"�Oƀ�f��U���ę88��$PU"O���u��'d�( Q&C� =f�s7"O�u��-���z�Z$��*���A5"Of�0!9N�xPB���="��h��"O@( 0��/4�"0C��\��R�'%�(��'�}k��p�ep��X0}2$��'��5�c��%�`����9C��9�'n�<(�b���$ܡ��/#�8��'{���&�N�H��!)M�v��9�'�9��ܖ nL�0Fy�^�!�'<���t�L%x������s.fP���$ɰ�Q?1��C�hj��b�Sx��M3D���Uʘ�i�F����H#[��r�B0D���m�V����P�PI���+�-D��wn���D|���M<����0�?D�0�,�!h`�����JW�y� ��m�L��d�	&���@sf��?�&ik����^��g`V�Kq&�:CF 3�:��;D���B���FX�C�1[�� :�o=D�H��)K!0�������H�=D�3*��F���2�9�Lq��6D���kI�����0;P�N2g�4D������82F���@�8>���N�<�%}8��� ѳL� h�c�J�Qw<�Ɂ=D�(��V&"i�YB�J0�$���9D������(���^10����j9D���#	1�>ѻg���<���xS,4D� �nS��\���E�I��d{t�%�OF����ON��%
 !0�q����WD@{�"Op�$dΝL.Y[DeB�(2E�"O| S�9g{��� ��H��t"O��f@�m=�A1Ď�0A�6��"O��횆4l��lH�Ut�S"O*9� �8��]p3	L�Y]�,!��<u�p�~�\��p1���ФWB:Xy�]X�<q�τH���sV�J��(\J M�Q�<�#��
h.�`��_� >@�C�k�V�<YB�V�U���J3I�2��hc��R�<Q�L�/  f�q₃h�b����J�<	DGA�x-P���aL�E*hP���Ɵ�r �:�S�OItы��1�"l���D:Q$n%�"O<ذ�H�D�(w�ǳpri�"O�$�$lǏd�QZ6lM���Y�"On���D�)�т�1C��@"O&`���:(��u��H�G���"O>)Q�k@륎H92�*���m����ć�]�|�&	�9��E!�
z��4�1L��y��1�Bp��B$0<�9AF���yB��H��{��]�t`� �@�I�<y'J�_���o��^�ȥ1�F@~�<I�HT'�9�A�Ƈ	��,��{x��*�
��$�%딼:�E�7Ȃ�7*.��7D��%��W6� i�g�&'@���5D� ��H�<"$���)eP:����3D�0�`��O���AgJY�Ur��=D�̉��J�4��LA� C�tb֨=D�t�F�	�kؠe;c.,7-,�׏:ړ"D�D�TR/�luD$R y2Zh�"c܆�y�M���D��� U_�miҁB8�y��v��YT�U�F�~B����y
� j��%�E�%����ǨYM�=P�"O���BI�_'<�I6!��!c��21"Ob81�X^8�:@Gh���'LAz����,3��Qh#�� @*��� C 	��%�q�� xX5�h*�����4�T��(+��}U�Ӝq���ȓ=��J��ҁv2���]0 �"-��[�H�2#��WS
8P��^1EL�ȓ]��T���)Fla[u�f)��'�Z�J
�/��bFM�.E��DK1^�l���_;��AؒO�� Y��V+f�*хȓ1L}i�#B={�
=�A�VǄͅ�T�萛����<`�$���уY�-�ȓ3"PU(@�~Sz�K�nG�s(����*t������ �xF� b���R�
0~�~C�	'!���`�!ԿJ!�q�pB��\ZC�h��@�6�\1)�hhq�Y��>C�	?K��� ��48#L�Ls�B��6�,<j�̵_hhyޤE��$�ȓẅI��5K�F9�r�R���G{����˒�ȒY\p�g�m&2P�"O(U�(�b?fY	�`�(L.�*�"O>��F�+4��H�1&��
D`e"O���a���Z`�rV�0�`B`"O���	RH{e(�(G�txI��"O�U�+�.Y����X�YPLѨ6�'O�i����9*���@5~�����7�-��L�#�nX�kJ ����6
^Ć�eL =@���1?v`dʡ�\�>S�-��w4��[d`Y�g�,���)ݣf��	�ȓ/��y�Fd� X�J��44������xq��/�˲X��,<[-����􉑇�ě�Si��>��]�(��FߋQ��0�A�4����'?R�'�Bg�"0�09�eHG Ƽ;���O��
�3���S�I*AR�ur�%Rj�x4��CԥH��ƣxgbؗO��R�߁;k�� R�� ������1qR�'r1��lr'�ʽC�F��ٴ@�B(dT�����u�~�Q�!B3q���/Ԫ�R�&�OT<�'��Y��F�h��e`�f��)O��Iq�������Hy]>���ȟ,Z�B�^��Q�_(wY\A��+AßPi���/��9C��\?���a�S�O��d"`�f���%ǝ�k�Be�'�" (E�Cn���H��?% F�C�x�#V�i�����}�<)�k�O�$??%?!�'Z@i�ƠP�O3,8�T��S� �'` ����R�b�HT T9Q�f������g�O���!�яzĶx�`�h��!7�'��I(�^5�����	�������$!� y"F٣}7�)C^��ca�'2J퓄�F�r��Ο�h2��##P6��#��$<*`F�>U2���ɻHN0��ìO�.N�g�'qlE`����O�Y�E�/:٢=i�O<ܳ��'F����<A�ɻL�b�����Z�耤f}�<9�����M�M5�@*�HKϟ\q��4����<	wh�#W��ժq  �2�X�#���?�r�����?!��?q+O1��4�$
�O���@EO��u=�5jL�:q���9`A�z6�P��y�K��T.�q�M'n���Y�CN�rv5�@�PI�T��Oׄ2^�y�m@��?Y4HT�GW���r�\<���Sb@��?���7�J��|�"EB<sޮ���^���ȓS��0�)C�L�"|�H7[�樗'��6��O��#�n��e�I��3�ؒ⏖�`<�A�jV5����?���?�v��xx[�'�Sq�����T��(������щ`T�)���O
�!�_�Ԓ�z�>���'+4r�pè�[8�u�i4*��F|�F.�?	����O�}��,@&X�m�Ů�XxjA�,O*���������NZ�RF�M"L�Q	�2�剕!��Qh(E��(WÕ�1��&I
����T�'����P�	�{�d���b�\u�fh$�
���w^�%P�ȑ[�&�;���?E�4Ek�Pmh#m�p�LlT�_�y2���:y���r�$!�D���>�ȭ۶��+R�1�&%SD�.�	;l�����OV�S�f~
� �a˄� �:#�+�+a���r"O�� b%V��N�RCDȘS�=i��I��ȟ��r�˞�p�u����[�8I{#d�8C���3���t�׊Ľ@�����`X�H�0م�����?(;&0X-\B�Y�ȓ,~&͚�H�	E�f�� %d]����7��QZS�O���H�H�>F��C�I�p�X����)�|�9`Ώ�*�B�Ɋ=�]Kfo_40����+t��d
	�~B�T/)�45�`�D�A�`��C�B�yb.�:�}Q��e��J��,�yR������$\�ʁ��Ӟ�y�g;�T}��+���Ҷ%���y�'��yC�5Bd��#&Zi��9�y�/H�KMb=���ӭ�V=�F���y�F^�>�0�0��ӽ *�����$�y��	�l!�|hW�ܪu��2Rk(�y��3s�ęw��0szh8P&�V��yBoM�u$@;G惶f �-xBmǗ�y��&[b���ܻ-X�09�+М���O���*��өp�>��W '�v,���h�B��:vȘ�If��Ǫ%�c�F=~������O �D*���!d����S�^ `��oS�9��V=�D9��S��'rp	�$L3T�hy�����o�M��I-��<ͮ�'
d�RJ��8@dȡ�(H	�lB� ��I�~��s��8���?+�͋'������㓆�an��'8�'�x��I�豪���R3A�7����%�6l�^�jd�'�P�L����$��	���e�����+�-����Rn�!�OBͦO�ĝ>�i4,���	)�N��eK�� ��+O :E�>���D^�e��UnR�0�ҢB�LJ��1�'��tkM���<q(
K~��Y�Y���P�fI�I���W���O���6������S����yu�>7Pt�a�=^o|���~������?�I�}����c�x��	O�b4��
*�f�$I���?��ϨS�Dɹp�	/X[�(�v�#D��:���;C��x�"k�>�� �`Ӟ˓�?����?QN~��?���LЛ��D�_�z�aa� X���'.2�'��'*�R���m��FU�YnVuPt�\SR`��x��)���l�
9*����w���a�#	<3�B�II/�)`h�m��IHB��\��B�I>e�v� ���)(�)ª8)RB䉝h�r��Я֙;�r)�'lZ�t��B�I� {��CM�7�>y�-%��B䉁H3"���)a�d$�0�F�o�C��
}>mC�&'mX{����h��C��4Nst��6���9gfϼ\W�C��?+�D�Q"KI,r)�M��΍h,B䉭V��U��A��c�\4�� @B䉹?�d8�m�0
0|1���1�C�	�= =(�ƋA��4��!p�����N9	|$*���,�<`x��HwT��s �B�v�T� �+P�y[��`X1	��W,$����៲� �a��Zʄ5S��1dj&�����\h��He�Z6j@Ƀ�&פK' y+$Iq�
�1a��9rJ=Z����8*J@aĪ *5�M�����x@��zH>IA�U4C�ر#0��P�*ј�l	z�<Y�����Pд�Šj��<���a�<Ie���=���V	�v�y3,R[�<�M^,��%�(�\!���a�<Y%	F����B;�4��`�C�<��	PN�.1�b+���p!7CJ~�<�3����L�0��V	V��(#�G�<�D ��/�T��f��=S��1AUu�<A���"�69�1.P�t)���3�Rn�<i� M�[��C������oA��yBI�+�J-Z�X�m	��t�D4�yr'�"or i�*�id�ad�Ʈ�y�O�&u~u���'�p��S&�y
� v���-_��$���Q�.(�"O�$+��&QXN���.Óg�V���"O���DL��zd�M�{�����"Oz��*I�	���bef�lR�"OH�r���<J$�t�!IsX�}k�"Oƨ#�͕�I�|��Ʀ�oO���"O�Mk��O�H�X��/� Q,1��"Oj�)�Ç�sG�B�	�c�����"O����9sӾi�ՇU�F��"O"�0��@V�=B �1,�XEqC"O김���r.�����1�"O6d���Z�O�e�0#&��"�"O�5j�&�|�'��s�� "Oư[�b�"���W�Z�$�#�"OB(�K�,��(�9�hi��"O��l�%}�J��'SȞL@�"O^-{��Su�va�%i1q�����"O��WD��XS�AeG�����Rp"OLE�����Y�n��,֏)��HR�"O���n��h���$�	�=�"M��"O���1�� T�u�,I�/'�(c%"O�!�W�\����.4��0�@K�!�D�9K�]Q��Ŝ/�hp��?�!�D�E"H��vJG�D��!�P�[�!�P!��`P�� @�����M<�!��0h��Xw�=�fr��W�!��G;o������M� �.�`�S�!򄖳l	Hd;1b�y���4GC�*�!�Q5(h��'ǒ,�B% ��O9!�F49[���+I3���!��(�!�d܄O��x���)0�yxŊ�5#�!�X1GB�����R�%,~A`7�F�!��р#���p6I��R��!���T�(EZg�2b�U�����!���/��yN̎{���%��
�!�� (�3`�E�2ۢl��]�!�Ӈ�6��'�V�T1�V��T�!���	�p#���xٸE��;b�!�dP�ߎ%� ��r���FF�!�$��>䦭��"Q4`�n�p�O$h�!�D�'N��и �ѴKg�D�Q咞?�!�U( �҉S�΂�B�A�L�|�!��i��jtF��ȡ9RA��!�3D��Q�0I��C�p��v�Y+L4!�䇑J-�Ec�.\+W�����9k�!��"��r��Q�8�������!�� *[�q���3�*�ô�'�!�$��y��ѐ$ԩ2��%�ccS�!�/RJ��)Ґh�(`s6O��!�D� "$ ��&G�J�����E;K�!�[�j������W�� �䘐y!��V6�L!�f�<�(�(fd5Ov!��T�y���^�n�3FbM�;!�dA�a'�bV=j��!1m!��G���H#�S%X�� 2�C$<�!��F�F[��pa�(p�p [�l��!���t����OQ_�C$l&(!� �G.���X�=R��i�#M!��e���	�j,q�	H��8pb!�dÕ
��}�e��-T�")NW!��c�x �A1(82���ϴz-!򄈬��!�%
9��f�\�r1!�d�j0���B���J̝m�L��'%n�c��,`�2=��ϰa�:����� �8���7��EIUMG�~X�X�s"Od�Y��Z)ȴUa�E�;0p�b"O\��)��F%���-�:JX"�"O�%{��<\0�qի�1�F�ړ"O:'U�f��0r��<?��@��"OI��GD���P�A�s�i�A"O����H���v��I�	}�~�h�"O��y�����5i��d|��30"O��%�>9}���� Uj<܁$"O��8&�~I���¯ԐQcn�4"O��ڃ)��d��A��$J(��!E"O~�j�g�L�6 c�N�@�D#"O4�9�o�]ɪ��IB�t�"O��.�o��x:�ǲ�<��"O��d�i7��Dkoj�`F"O`@
���~U�L	�ܗd@:�qW"OB�`R�dF��C����e�n�"OTYy���p�F�z'b���"O��DN�=,D��Â
)��i�"O$��mU1gtn�����8!�$���"O�3�g��c��a�b�>T�ȵʃ"O�EȢ
W9g �y��,�6���2�"OL$�A��;����e_�W�T��"O����j�0��I�e�Ü8kB"O��Ä�$PR`�#���-���y�"O�@b�bԛp�J0إ�V�Z�\�2�"O�0�fHN�����H,��is"O���J5f_.5�׉ں=����"O҄A@ ��@��.K�`u�"OXqj�	D�O���ekC�C�ܕq%"O68����S�p��S띌Xφ��"Oz��p ��e��aK�)J�#Y܈("O"X)Ǌ��?6��h��}?(�C�"O�8XAD �������F^��ȓM��X��٠ v��%���OxŇȓ'�,�i�MN6�SI֢.��@�ȓB��]�wJ�1G��\�3��JPr �����㰬P�6�9P�)���Ն�G]��P�B	^���c�j�
H����7;��+4�CP�t�S�d�%��Ї�4��2UM����;)׃0N�ȇȓ2�p �Š��[�J�r#��?n8���3�:)g��{оajw�5e��z�� U�sD��p���2Y��ȓo�2MX��@,\�����9��
�'�.E[��K1T�za��ܹ5�!	�'n�A��OH��Z"�Lzn�q�'Y,Qa�G�^���i��ѱx��X�'�
�x�o�����뷀�G�V�
�'�00p,�]�� �ń�2�����'�����N�������X6��1	�'�0X²D��I��$j4,C������'�#��I!^du��/�GLvb�'x�1[�/0�*�;V >=d��I�'�T�;���,x�ǝ�!����'���	�%ч;
)(u"7,tE�
�'UȜ�A)�.,��x��͗�EF��
�'[�PO�� |�Q��±R�9�'{�I:V��5>��� 5�	��'Ҥر����fz�k�k�L��'5���$�&_��Fhd��'T����'ɭax��8ňV8TU��'��u�t-ë�ȥ���*
�@P`�'���G�R���A "�*d����� �\����]�$�wA�?��S"Oԕ��fր\���ATfɫ:ᮩ�"OF䁳`L=)czei!� = �
9��"O�8��D�:Y$Vm@�
B�y�%Q�"O��(���8yn0�3I��v���"Ory��*��������D��&"Oh�ȂDΛ	���Ie�C1���"O %:BA�"�đ L��@��Ub "OP,s��lL���̪|{�)!�"O����{�(�
�NE0]�@��"O|���lO�j�d�
Ug�3��L�v"O�y*3��	��Ɔǰ0v@���"OM�҉ k%
]�"�ʜ68l�ش"O�
���$e� a� ��z+f�b"O@Z�-�hv0�d���{�"O@p�rF	�$x(zW%=$N|�"Ol(z�Ŝ !�t�%�\���j�"O~�s�ND�U2�ҧ�.��5��"Ox9�ց�;l2���ؖKʹ�Cf"O�e�o|��zRKX�HUK&"O��V$M����� 3\;e"OL4Bv�[�v��P�fB�xJ:�P�"O��J�m�. ;v���)<�� "O�,�B�ĝpi�Q�te�#g&:�P�"O�9�S��/W��MZ�$H9Ф��"O�#ʘ}�<u���%F��M��"OZ�!� 4t�B)�����9�qA�"O�� ���MP�p@b�M�v}NlR5"O*��& �/�29�BJ�h�h��"O�td��<�Q2h��y��\b6"O2 ���K�fh=�q��5|����"O�y�v�H�SX�(Q-U#&�ݻ�"O��Ck�3h]T�5��,2�CQ"O�i"DE�b�I�f����իs"O`��'@.z\3/���@�"O&����Ґ�����А�N\�w"O&�#�Ob�؀���f�Y�"O�����/]�j���zH�y��"O"y;7�Ф4�@L�&�۷\D���"O�D�v��u>YX7��1�P�*�"O�����?C,-��R�8�:U��"Oa�w�>61�i�qh4$�(lS5"OJ]p�.�:8~>L���R9a�Ԝ�"O��r���nv<�0�-?wX�#"O��X�	A�����4MܔL u��"O��ye���� M��l^4
<���"Ov}��.=�(�rq
C�]� ��"ObI��CK�4�۶�\;w}B�"O�8Cԁ�9�"a !���5>�h�"O@[2D$D'����fvK�e��"O,	�&îO�
,P�c �q2B���"OV�*�e�8
��p�s�ۇ6Q(�8�"OF�@��IJ~h�"�8]�PP1�"O� Є��_^�=Ab��0tM�U"O>�"b�ݢ@u�m`� �cj,4"O�0`ūE~��� fȠ��u"O��� T ��=ʓcԷc������ӡ]��Er�A'�z �Y�<��'KJ!�^+mҘ����
	�Y	�':��/�#���E�O��VUI�'�h-8��P��`tdF�j	 ,P�'�$���(N�X|�����c���	�'�����5)'j�q6����I	�'��x��՗\�6���	C�	��a)�'>����U)d^�7f�1,����� �Z��X���do��.�Ҭ��"O��(b������1�~���"O���p'�p�L�8� Ý�����"Op� q�ۼנ�#��ΆH�0���"O��6
�[��8 �*Fv�z�"O��WlZ�ՐTi �Rp�)�c"O���WlL�~��UْTB�e�%"OT�㕤�tC���(�t�K"O���V�WB�ĖO^͛�f �yҪ�9=�&�Җa�K����)Ӥ�y�gA_���/��X�0�e?�y2�Z3�}����|�����	�y��1��ڑeۚ&�����^��yr$8	��|wj��%�jMC�-��y��-�{p�2t����£\%�y�k�!/H�p"R�Z��UW��yR׎����` HP&��y�J�T ��N�3�x���Z.�yh��1�"͎�5o�퐅���yr��:����	�0c�Yڵ��>�yR�^8�>���K���e��gE�y�	��F�F�3�,�>85��C6	ג�y%��*z� r��$>S%�!���y�7jqM;�.�2�ୁ`���y��	���T�;<�i+Qf
��y�Ό:|4[C�
.<X�=� L��y�'��:ZJ|�`�69U�:C΃��yb�˯D>]a��*,d�z���y��Oؐ��$N�!A��Q�CR'�y�d�5B�T�!���<G+�\z����yb�I�3b�cB 	�wF`�C�����y� ��X��|�SKňnK�8�d���y�Hg>ND2W���6��a���y��ҴY��{�b&�i�3��
�y�g˸J�Lm���V`= `s���y�E��`��s&�C�9�a�܋�y���<������P�zu{P��y�%��B��� Xp��S�[��y2�2t�:�򣓞i������yb���S�M,U�]�-��y�V%U�n�!�*BGJ�ⷉG��y2��{�����h.y��=;7���y!�.[\l5��d��!'*���yb�ǹ���+ґ�"��+ĳ�yJMW��p$�֊<����0�1�yB����|����1@i�`g��y���5/�J �5bՙ9<"�k0��+�y���RU�b�1�V`ϐ�y��ϦW�1 )��*����@��yr�:�օZr��0�"<*#뛅�y��5o@�	
 ��0�Rh ��H��y���oj��'぀'�����dȻ�y�� 2+1c�K��:��^�yb�܏Q�xxB��-
Č���l��ybիI\�yJ�Y�Q�dA�J�y���б9����F���-��y�צCp��k�L�6�&�.�J�'y�I��^�lJ�H͖\��'� 5�A#�a����rO�[�DXY�'yT��qM���Ѡ�̂�'��mc�'��>*?�Mrb'_�X�2p��'�Ї#�+�n�;!B��W=6��
�'Bn�)G@�ep0oɁIq( 	�'�0,p"�ܳw�� ��kME$������ b�B��8~w�1��	�=� �˦"Oz�{���,"�j�d��;f���"O2�1�Ʉ=�� ��Z4|�n=h4"O2�k@�*w���hw�͝u=�X��"O���C��(Z{�X��ȟxZP��"O��ҵw�	:`Ņ.�*�)s-�B�<qs @ y��`�0�ݗ-�����V]�<�W$�n��ܙ�O�Q� !x�V�<a�$�7�Ѡ1 ��uX��fU�<	���h�L�5�X�>�PY���OP�<1��	�lA��o�
`��Y���Y>�y�mV�{�6sQ���d�5
�����y� ��n����W���Y@���<�y��--44̡un��x@�4�yB���i@�i����݈D�n
��y���i<Ce�ʙB�a�mH?�y2ʌ��Z�Պ6G6��A	��y��K�r���֧\� |��a��*�yrK�U�6hs�ǡm�]p���y��B���;!.����D� �F��yBkA#m_f�C ����0bʭ�y����=vؒ�C.�$���+�yb-N0���$e'&����v����y�*R�cz���D��/(��a�F@��y"e̲��@Z R1\в!→�y"ޟp���w�A-3����T�ʄ�y���?j�|Miӫ7'����f��+�y���c�=#��F vE��@��y�R�&ъy3��Y�2�����+��y�h��D�岖/�:;���zvd���yү��B�BH�1Ð/,N�yF`5�y�)�o��š�E�P��KQ�	��yb+ -������)X8śƟ��y��^)_����@MO�_��H�����yR��=Y�~����8)�|��e[��yRF�)fu����AÀkb�9Q�Փ�yb�D0��"j+�`0�pB�$�y� ɀpɒa������A�?�yr ɊA�ޔ�M���ajd
���y�(�=�R�;3n��6F�@Ï^9�y"K����J���d6�|�2CJ��y%��#�vѡ%_�ew8�E���y�L0q8����e���J��W��y2$�10h褙T�I�ap�<����y2#�<RXn���	-aN<�qWJ���y��5j-�C��v	 tO�/�y�Ї+��L��$�4(C�!�:�y�(��<�*D�@̀�U�,9	"l��y��v��s��,S*�D`y��a�@����͂��q*@�e�I@�'\q�T��6;�N"$'��K�xj
�'��(g�Nf�`�7�_������'׼�3�jT��l O����-"�'�|��쐙dn�h�!A�3�<��'�5�2�!��H#�ɇ�w�f�{	�'\\��,P�h`��PE���"�k
�'<;�Y)���[%�۱픠#	�'�ڵ�E �*v.�gH� H���'I�m�X�[��U�����9|b%�'����D�=�v�KR+�>p���'.��ɴnQ�`�f�Hr���q�F�)�'��0����rN"tRb��zO��'��$x$'C9y3*=1R�Α&��XK�'���#�^Gni�����Q��a:��� ��9��e'6�4��Q��|�Q"O��Q�ȷh:A��#5�L��"O*�e@���0��f�6�(�x�"O>ԩ�Oi,����R9:���P"O�-RƦ�q�\��_��,݁5"O�X�,�8���#��.q6�� "O�|��'�<r\b�h���?�3"Oz�"���$�>t8�N�"6A1�"Op���M�����:�m�(*���k�"O�$�r��)�	3 ��Y3��"Oxd7���&Z�(�X�#i�b"O��hc]�)`��t
�vg*��"O��(�)�-8-�T`���5d�	P"OPI�e�C<��6)K�.N���"O,l�a�	%:�(`� .�;]HJ%��"O&����:e�|(�+P�y�����"O�i�@��@�
mH0�^&c�D�p'"Of�цM� @��+I�Sa&ٓ3"Oּp�a�:c<d�6�ޗAdT�5"O:��v���_lN�"��+���B�"ON9��*��/��sb@E�~d"�"O�P85NU�E���s"�!<�!"�"O�%0A�H@¥z�@l�D��"O��R	�0S_DHڳ'�/�غ`"OB��_8P0�q����LC l!��=N����AF9��E&�g!򤏸Na�pI �0$E������d^!�=�OR�V����� 7!��*XԀ"�/L;�n���� �!�$͉�΁Hꃫ�n�z�I�'G�!򄏠g�`Q��/�Y��@1H� H�!�$K�6<���E��%�V�ܩh'!�8J�>`��K��Y�6yy�"��q!�d��"�h2�ߕC�P5@�
DK!��"���K��(@��2r	�7H!��qݸ`C� �йS��U3N�!�8����BD%~��,aNXk?!�D_�=���i6#J�'�������!��P�l,��fۭp�0]�����!�x8L��#�zM	��V+�!�d���L� �	L�F���)O�!�dգv'$q��A�=R�������+b!�ȻJV�	&�S��0�� A�c:!�F�#mT�SF�M�;�=0���<�!� !�)�p�q�j��EP?04!���CH$�Cf���S�ͰQ!�Ĉ�K,0�H�Q꾅��CM�^�!�DߛC������.��0�G�ȻD!�$5*����j@Z�b�Jd�!�D�&�Pnʰ#X�y�aD@��B�	�Nd|�&cRrLed��%�C�I/S��x:a�+{&��r�9-�C�I�w(��9V)�	F �$v�B䉀x�^��;jF���}x�B�IK ��b��0�:�RDG�3��B䉘Y��5�
L��F4��e�7w��B�2`�:�rGb��X�8���I�lC䉸�ԡ��/�*:��|�6� 48�fC�	�ZҢ3a&�;7�}�R��J�~C��4)�4�x�\�l��5�bO�\C�	�EA���[=vi�!�X�$���c(S�sC�-���6v�"��O;�D#K������ؘ@�T�9&��&J$!�,rI���OșZ��qqb�#{!�M��c6IU�G�!��[4`�!�� |5�U��#z0fl��M�2t����"OdM*��/6x�y�= ��"O�9@�+R07�Vm�g�� �$��"O渫��G)�}�k�:m����"O��XS�>p����-��QyE"OH���IG�8�}┎6��9r"O�E:�W�]��ec�r�ҹ�"O@ �R##gc"`�WBZ���"O�@D�5c� �D���m�,4"O��#�a� >�$a� �B�A"O�5�4�H�K�vd�S���\"5"O|�[�mS���`k0���Ur*) B"O*�a�sȔd�w��4^I��J�"Om����Qs��4�]�\Y��"One�WOw�*h����!�$� "O�0I���������K_�Az& �R"OqG�D��n��Pk
gZ,�"O�}j���N����Ą�JH�Yw"O�$q4+�,5�|�6���	��<�0"OD��������`4�R�8�0�"O�}�Ɲ=oV�@� ��b֬��'"O�,P�Ayȹ�sb�*H�^@ru"OF�p�D�1 ���h"�x�%�$"OT|�v,\
S��H#a�/���"OH�0����(�k�ŵM�d��"O���SϞ�W�R�$� @���"OB����T0)�@K��� �bl�"O蝪�hŀqQD��-�?_�@���"Op)���9�UB%�@/p�!3�"ON)�+'�4�C�+� ��p:0"O�� �Ѡ4����^&{-�l�"OX|�!E�$>��i�"הQ#�!��"O|�L�[��w4�#"O�Y�3�=����c
9{ <�R�"O�`�7*�Q�ҸH�W&W��)��"O��E F9p��  �,=�4	�"O��Jg�؈Q�"��7!T(&>�U�'"O�0�b��s& (���Y�lDH-h�"O��`�ޛSA�9���!3���)C"ON��O�3D�����J�wm
|��"O�pEb
�ro8�jV�P*^O�I�r"OZE�#��[ezUæ��$Z"��"O�YvOܕ�\AA gݤR���"O�}����\<PA� �/A�V8R"OD��0�cK�0�rF�5z�i;�"O��/G-��h$h�M�&�{q"Oȴ��B��n��ѻH��%�t]�"O�*��y��)[E��j�,��"Of`9eL.w|�A�y&��p1"OPAW�����}��Z�18�ipw"O������#�z�@5@��L�s'"O�p���t�rݰiu.��&�!D��`^B�v�Y��9@pd]Z�=D��į�*2������:v�S�?D���T��b4j��h�/X`qp$ D�l� �!c��R��O0:��t)a�=D��cև���� :�c��/D����mr�y@wD�98*q���'D���" 
L���L<��ؓ/1D��Q�j�\�T��q�Y���N#D��ۤ�؀U���z (� 8�|�6D���h�I�@�VHo��ec$`2D�s��$]�x�+2G��W9(1
�-/D��أ!���9Q��
Vu��d-D�� X�q2([�-E����6i� �Q"O���g%؝3:� fo�>5]�8k�"O@{�HD#X���/�e����p"OFhX��O;M�%E�
�� c�"O�8�l�'Ҙ�����%���"O6�E��4>���C��Dy�C"O2���S ����S ��=Ϥ�W"O8��Ʃܪ_�Y���ˋ@����c"O�ك����8�f��_�0��1"Ob�СV0#�CN�T����"O�5iUAS?iOm��M�5��|Bp"O��,b\�m�%��8K�8|�q"O@鐡��L�|P�"�$�g"Ov8�1`ͽ<����(n���R�"O�u冎 Z|-S��q�
)["Oyp ���mo,y�W	]�bD��(0"O�@ �X9'X��]7
�Q"O$�RO\-,Ր�yQ�I*w,N[�"O�EpUG��u_�ܳã\+�<��"O$d�Q<$��iN䍣�"O�ĳ!+��"I��X�x�("O���W���R��Q��1��͘b"O�tGZ�X�8=���N�Z#J!A"O�ȓS���g�����U�P@�)��"Ol$y��		-����wN�n!�2r"O�X�˕e���$J�Jx��d"OV�J�#�+c~��B�С:�p�C�"OB��!��09�tX:BO	r�(@�g"O�$CDW�S�P�'��S�̉H"O��K�sb.�)���1��i�f"O��+�)
�L��bXk�d�@v"O�4���A�,:B����ۇ"O���BB�>�@밯O~�<��5"O��Q�_�df���,ًl�*��2"O|$01���hx��G��qz$"Ov�z�_�n4��Xtn �^�P	��"O��`�=.�x!���))|l�R"O0<H`	�=�L� Ս�" D�V"O�Ku�Z T��ۣ�I#WB�	`"OF�Ce�خ:���(�+�� �|b�"O��1�l��}�AB2놢�4�b�"Oh��Ѧ1TL,(#dD X��Y��"O��[%L1J�����1(��1�"O��	!�@	`�]����r}�ۀ"O0|3wkģy�ՈEȼ*�B�kU"OnE��I:?�l�z�B J���"O�(9&��Qf��� N�H�)�1"O��d�đltay� 9<��	�"OB*ؔ歈p Ή�r���"O�|��'��`@�L��J �c"O6l�K�v����V:J��B�"O4\b�d�+M�9CE�!�Ҥ��"Oe2"��:Mb�1G|�p!�"O��"Ro�Y�"e�`.h�Iѡ"O���dތHd��z�R�3@]�y�OϏP]D��J^�%bQ�1�\�y�ɉ'�p���+���ʒ����'��{���Vq��Ga�$�Cb�ǹ�y���O���V����`<�r�
�ya��[6@j4��KJ�Rr�M1�y2�=J���ʱ�D>E+ur�HP �y�
<��ȕ
ę<q�eם�y��,����ȍa��3�E	�yB��k��\�a��]��t��H �y
� .�;�fü-4:ݳ`R4TᚌR'"O�$��G�4����� U�Dp��"OZ��U#X�A�TX�f�CUx҂"Oڥ����$b:��PBE@�@�i��"O�2�i�||���%ŝ�I+�!T"ObE�a�P�a�h������u��Y�"O��O(d'Н���5R�h�H�"O�t0�g@�'�z���>,��iQ"O���&�N��H�'АP\<=B�"O�B��Y^���@L�9H���"O�|�⋘�&�l�rƎ�=,L�3�"O��H҃A&�f��5d�9t��`�"O�u�G�\�T��D�ےr��"OP�20�Z"h�p4�!-:I�
�)q"Onً�S6Z���B6��c��ᐑ"Of�HS%\��l���lI�[�*ܢ�"Ov���L8b\|���d	���e�f"Ot�J���<M�%�!dP�5��Ai "O�)1AJ�e�aw��3�Li�5"Op5ð���T @90D�'[�n�"O�`W�ҫv���9b�F�awY��"ODQ�tl�Az<���aB�:�|�"O�E�ҺLp2�9��N�4hQ"On��e�ٹ.mD�{�@b�ȗ����y�",�P�!ibz��6�2�yҍ[�H���2�Ib%<t�ӄ�y���3���s��Z{&p����+�y����n�!�ك>�Ա	�FF�y2�<E��*E���>�:4 $.Ҷ�y��ɟAŴHb�A�$˂%s��*�y�̑�@�B�!v��(��$�FƆ�y2+A�$IR�#'S	%���5h
�yb��t�������qPjĨ�y�&��T�pl_�-�T|y'a���y"gؒ��uȐ��%#�<|"B�D	�y�B�Vr!��.e�n����T��y�%�A%2�
Hd>t��v�^��y�M['!��[��N�l�td2v)ؕ�yg�$+���k��gڤ0��%Z�yR��y#��2�˚[�,ћ�D�?�y�杙!=Bh�T��W\0X`��yr�߸�$�q�n��T���V����yч�H-M�Q@9�U�Ұ�y�`�-b\h@!�	Me��b�� �yG�6��t����FJp�S��y��\؞P"�«D8�$1�-F�y�W �����*;:�pl�W!�]�<����-��� #kSx�sq��!�ļ�d5R��Y99jcf��0e�!�DEu�y��Ϟ0<,e��-��$�!� ��YS[5bt�V��Z�!��\�k��lP$N�B�ѽ<'!��!Dd@�%'��l�&� �<�!�$ɨ~���	d �KҸ��AKzG!�D�4rP�H� �r��c����o6!�	ZtpKWIS�^A8���5c�!�5Y���v�G�W/zU�`�|�!�d
J�vDHd�N,���r��
�!򤘻a,���눟n����'�F�!�@#�L����|�2u��@�:o�!��$+.�xE���t����X�!�0��ě��
 jB+��T�!�d>��Y��F^����:�!��f�q�R畦80"A��"��!�� D����؇A�{�V% %�V"OL���KU��\e���ğG	��#�"O�h[c�S0s�q`���+��xI$"O��'!}h,$�����j\�"Oh1�A0��e��Λ.(��J�"O��PB"�;��X�&T:$Lˆ"O�-c�eD�E�%R��@�K�x�"O�,��N�]�d���ޭ1��J�"O����g
(���ț#��̑G"O�]�')D1%<~�"��@!JP�"O�4�`,�)!&�c�G@����"OPܡ��C,$'@1a쑷~��m �"O �B1�`�,�iL\!Dښ��2"O��:�I�8Z�ƈk�� L����"O$��f��,$�
IpCʄ�I�� �"OJ�D$�x�f��hǂl2��"O.A��b��3�.u��H�-�t��"O��  �Թr�c9<nx�:s"Otdq�j���&�X���"O��QT��OAޅ*��1;,�c7"O$����	T�,s0�߅#P�ӓ"O�|a� �3}�ܑy�K6g

�;1"OР�@cZ���pc��I(.�Re�@"O<�� Mt�5U,
�m�D��"OƁ R��@a�1�d "s#��C"O��A �;Om����r�L���"O^��\�9虈$
pZ��C"Op	���t� �d�ER��ab"O��"����2��HAd�H�!�ΚT%��v	F�����c�(p!�$�p%^!�RNU�c�v��3&<!��
C;VZ6�'K�Eb���!�d�m�c��6iSlu�v�0M�!�DF�RZ�qi7�<� A�4T,5U!�D�?n�I�,�?��p/J�C&!򄔿�<M[�/ڳ${r��u�	�!�dJ==p@Pa"O.Lk����Քu�!�d\L�^���O?Y�5��:�!�DȬ;��������\/���!+D�!��J<�+p�W*�� �M�91t!�d��L��7�H8\�\��#���s!��!/rD�@*=F�&�@ �'S!�DîL� �䩓�d���	�&�!�$�r�T��'��~����p�!��5Q�J8�������%憟	!��fb�]0M��s�Paj�%W?.8!��.��@Nv��$�D%�i!�P_�ԁK�A��0M����D4D�`�GoG^�� ���&���
�)4D���M[6� )�a�<9��@6D�,j#�[�Y��\�4�דf4i�4#3D�@��^+5�ysw�ϛ�Q��0D����B\.]�=���	�-��)��;D�j��M�=,¨󄕖|��\��.D���Y%�`�pk��NނC�G.D� i"�.����T�*Lx���-D��ZQdW�y��	(��U��(l8� -D��ե��`�c�c��j�=D��!�K_,6|ʔ��p��I��$<D��H�AR*_�P{BϢx$I
b/:D�`:O�n��@�/�&+�<���k$T��ȴ��RJ�%@�ߦ^�$!�"O]3FD\9j�Y6�F�$���b�"O��X�eJ T���m�?��z"O� r�ru*�~p��[�y���S"O�,�w����`E{�k�^"���S"Oε�U�K1�@
Fm��6e�1X"OH��%L-P%��Cw���Y%��۱"O�󷬊�9@T)
���{r"On-�7�_�1N~�Ȧ�2x��w"Ob�C�M�a�H�4��\�%B"O$����P[t0�d�H�0q�P"O
��HU#:ư�vc�7�2��c"O&�r%T�]@�b5# �q�"��"O����'T"F����$�
���$"O
�3G�^� �����zu��"O���uA�r�����o��ы�"O��$�F<`�\�����a��v"O
%9e�P���4�E]L��)T"O�Q�D�Zy��A��\��U�%"O�`��V�ט\R�.@Q���(v"O�@���yJ�� n�5�ʔh�"O�칅���L+^8��\6m�Re��"O�9�^"wb-8�薠�&�"�"O�@z�*����� ܬh@x�Zq"O.�{�M��6���"X�V�	$"O2�$��@䚄1T��	��dҥ"O�A�����lvQ�4B�s�N%X0"O���7��X�:�Ӗ�+b�^�1"O]��@�!k�X���­z��"O��H �M��);�L�tDjD�F"ObuY�؄]��H���9J���
�"O�]�u��B|�@DM-$����"O~�B
T�-W��'L��r!�}BG"O�l�2K���X@��G�o taq"O��#	]*DM�k�(ʉx�^�X�"ON�:�b&q<�K��p� y3"O��V�����ר>��=�"O&$�E�N��b%{bD�.�Ԙy%"ONH��K0.�6���F'T}���"O����&�-�V��b��PY��"O�<��o`�-X8�䴻�"OȀ�gH�P{`�03HO>}�8őf"O���DŒ8b�t�K��2vh��3"O|�;Bj�"�=9��\tX��"OhY�T����R��T79�� "O�����Z3:Œ��� ��k��q��"Of<�Q�B�RQ%��
�2B�>aCb"O"���&� ����r(�>V�x��"O���,�Q�v�Ac��&�֩A�"O�tH
�S8�h�h��.��C"O8�Z �
2-ȝCq�V����U"Ox�3q*�t~�	��@4�	u"O�‪	.'>Jy٦Y�xE�"OJ�{F�Z�@\\�Dݨu���"OF��h� NQ���s@��c�6���"O�q�gC0-��H��%��u��"O�1*5�Ч3��e�"�͑��9�A"O��@M�Mˢ\���Rժ�b6"O�pc2��W��k�Iǁ ^�J "O�0�Ũŗc@ �q+�"9�8�"O<h{KM�a��4S�o��^b��`�"O���/ύ(�pX�-X���"Ox��@��r���G��=;TM!%"OLęG���.~8�b�[1M@tp�"OJ���䙄Bv��9�H̋8M��"Od�f΄�G6��bjX�4/�	@"OD�b�I;N�zi�Q �5e��[�"O� ��Kpɚ�U��|�)��@$M�"O�D���N�r�a��(T�>��J6"O~�j��ӻ5�|ɂ�JZ�Eb���"Of����:6�%	F�� o��`�"O� �)��x�aB�	%f2,
�"O|)##�B�x�P��g��tW��r*O�ݘe�s�¡���:"1ʅ�
�'��Dc�On�����+L&�
�'!�yh�GÂ.�"���sV���	�'gjq���X�+eB��&G��6��x	�'�" ��W�K�\����'��$	�'����$�	R��@�R��� ��	�'�� A׿J��4��N��)�	�'e<%C�W#~h,(2 �2#ݬ�b�'�2�jJ�,���9Q��	0����'4�`Y�th<SpH��xf���'��9��T��p��!rZ$ �'��9ń��.����%g��B�'���`�س	��}��O�'��S�'F�s�J�{E2�U}z ��'��-�����D3 @ri�j���'�*��N�M�PB��&]E2Q��'W�}crkۄ��4���MNX��'�&����<��1 aD�F���'y�H�v�Y���"���?\��	�'�d����"<$��C$�b�B���'~�=" j
$A86x3�"O[�Lĉ�'O�	�Ac#+�#��Z�dl;�'���qv�R!�c�S+M����'~$�#īB�HwF��v�SG��lK�'C�1x�.��&'�-c�O�'j<d��'����"�>��آ� Y�5!�'{h0���Z9|��UI��Fcxt�
�'`N9��C�5&�Ԁ��	>0�p	�	�'R�˕dRL-:�3i�* �a�'�Ή;���gѐ<i�H�%�X��'o���ӈ>n�.�;@(ʓ�2��' !P����>=�M�5���'o`ɛ�.Ә���kU�w�U;	�'�xY!��Y/|����)�;F��@Q�'A6�9sۙ{Q���cBѱH�8�'��,����J���=�����'?p�F)S��P��g)�<e��H�'w��P$*I"GW/�< ��'�ʥ����}(�!go/�`0�'LZ��1�ږM�Pm�'<�b+�'e�PJA�Τ :�Lbg��m6�	��'x��#W��|V\��ʛ�~���'���VL�I0���I�P�
���'�!�螖*؅#+�S����'�$9*��gz�%�g��FI���'`�l8�#�"^�<I�jڕ�� �'�.��Dɋ!}�r5�X�Bx�`
�'{����,�
~~���G���Z$
�'���@m��z���!�#�h�� 	
�'�\0@m�Ku��{!әW�$���'��y��S/�5�F�S1M�RJ�'����ǍA�
����!�J�d��'zx�r�<��ꆬ� ��'��u���_�Xtx�G��/C�hK�'�8���!n��(�Anͪ9/~��'�[!�T�u�n� ��e�$��
�'�q���9pf9�b�?^��̀
�'ܲy*FN�0n�
P�Q4��	��� (�� ��Uݐ}# ݃�D��s"O`Kr+D�S�v��¹$d��"O�Y��l�; !�����	�k���'"O����ލ"�5#Sc�E�0i�"O��[E�@.o�0���[V0,c��ǟ�`��%T���	_+>YԠ��5o���JO'!��RGJ��	ƟP@$S0A�0`����*V6�a���O�I�k�T��$m�?���c�*ϺKe��X����aE�2�%�c�!I��-K�Wn�8���`ԇ
Nu`�U�چ+�*\��NR�	�*�$��@Ҧ!I|�ش�]L��o�X�jո�.Q6>R���	E��|���߼/e�,XD���Qq��K��IQ�|��o��Tn���9@iB>^�D��ɮ¦��M��X�2!��M�����4�6=����O.��lӞ��m݃~��G�B���EA��.�
���ڴ{ ��K��WS�vHka�	�v�؇C�f����.BB� ��ٽ�7-�#��I�Oň3�ԺW�U8�u�<v�v���B���Ɛ��L����N�mO�a�#�i��p���?�R�i��sӐl��I�5l\R�(P�#�!@"�O��D�O\�D�<����O�ESQ	J7zkdP(�j��4��(��ʦ��޴��u3�y{\w�ؠ�F�=��� s&�1MH�yu �<!V�ސ4X�5���?��?���P��x %dG�_X�9�@�ޖi��x�N�h*��C�=�L���a���\T��h�CU?;����͞�����ޔ$?�q��&M:�tx��� '�>�4��I�C�F���'b�=R�a��D(��l(���O�lw�'�x6�z�'��I:1��ę��ɤ9
��B��W���➼�퉂�J�XѤ�$~N�2@f՞`��(�&�iS�6�?�4�T�i�<�Y��J���ض<V&]�3��\8���s�)�?I��?I��2A���+����P���SN�*b���gΒ\˸YSU�H���ѨK������V.��O�˥jUP���VfRfjd�GMU�Z|0!D�	B{��c��K��7M��$(S�~�	��8���9�Lx{mݮk�8m�Gߑ	�L��a����	cy��'��O��v����oʺ"a�%��"z챃�"O~0�#��$Y�
L˦�_
y��:��O�n� �M�*O�Mp�����J�r��GGR�zh���F�ri���?����?��
I<]�v�	c琰���z���S�.�paU��?"j�[ejR�OvH#=�Q��h�|
Vύ�'\ =3�����F�Ǎ	4)c�	�J�p�*���(G���2� ���G��$�ɉ�MӀ�i�bR?9�gc߳t�zX��N�=7��xBE��?	��OȰ�G.eј�qs/U�W���`�1�O��n��M�ڴo�`E�T-J�_�"x�*z�,y��ES�	���i�U�擡Cc@�IПoڳ��7��'1�,}{u��d�<cpeQź��� q��˧ �����Q����Ok>rVt�Ҥ\��"��E�F+��:ڤR�D^� �����K/|8�lZ�r#���|�1@�<�+0a�Q�V�A�(JX�l't����O��o�ǟ�F��4ED`(0�F�aL���"D�V���?y+O���D\K
�r���gJj}�!
�l����lZ�ML>y�m�8�u��ۏR�H��*ް �x��N�T(��O����1S 8  �   _   Ĵ���	��Z�ZvI�*ʜ�cd�<������qe�H�4m��_;:<��iF�6�T.T ����A���v�@����:S>�n���M�տid�	]����D��}:�f��U�i�5#��K�x�
D��Dh����{��]�'�r\n�e�8!R��G�&y�lQ�$d��X�d���g����'��`V˄G�d��'tX�c`�\ :���	a�[�V^L��W���0�488Ht��'��tC#by�?��,5PR�8��@ǟ\���8R���:f�I������$W�@+���������й��w>=8��$gA�=cG.B�бǎ��Pq�#÷r	�b�8KS�7�1O�I��c�!oB%��. ���[q4OxH��$��O��҅:'����GA�e�М8@��s�'�h�Ex��R}�N��F�"qa[�O�fU˗m�"��	�`��#a��E�4�|Qc�;Q�+�쒹K��fiXp�'^,�Dx�KB{��U15�L� g�۳�>���}��Y�'!`��'�Z��$CCǦ]rF� B6!,O�c���V��'$�S�n��Z�PF�D"�భG�'�)Dx2mɟ���\ �P�2�'ը^8��6�	�^��X�"�xi�,R���qm��Q
��"ł��~�C�r�'�~t%���'_D%q���C�! �jE�y���+��h��I*Ҫ�	���Q��*�k�y>��H=0�P#���=��K]�	"I��18�$��NM� )���x���>(�p g��~ތ���	�.�M{�͚qQ�P��I�3B�u����6p���2�E QªB�	7XW� �  ���yr
�KO��@��ML
zx�T Q�y�'	�Q��#TA]�[QV�q�α�y���?А$�
Ü~����Ad��y2 ��*�q����}K,es��A��y"��=?�*��DV�z��$�E��#�yr@�����#A�P�;"�H��yb���7��(#�ް-@��f���yl�%u�~$�5�)v�(����*�ynDҒLAe�H$ ��y��+���yb�X
t����;tĀ���Q�y"��?
� ��@�yJ���M7�yϔf!,q���7VH��Z��y�a����6�SN�P�p����y�"͞#�`"֏8:��b���y���>[^T�9�d +0k�x�S�y"ˁ������H5`��ˢ*��yR�y�=����XW&q������yB+�    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  ��   �  P  �  �  *  �5  A  �K  JW  xb  �l  Ns  )}  d�  ��   �  D�  ��  ʣ  �  ��  "�  ��  ��  T�  ��  �  D�  ��  ��  ��  �  Z�  � ' j ; R$ �* u1 �7 �= e?  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C�'g$˓T����[x��3��&1���ȓ|� xKB	IX� ��nĩThEz��OT�}2�I�*�x[����I�'(�L�<����)�� F�D*2��	+�J�<�FOɲV3Ĉr�f�o�D44��G�<��هyF����#$f 	���A�<1f`�I�&�	WdJeE;�,GU�<QW�@�R���[��A�Ca���T�T�<�#�[�VXx�*��B�j:"��7��N�<��e��jZ����g��EK�J�m�CX��\�����$a*8���A��S�#D�чm�:-4���Çr&���D�#D���iӢo(� �ᛉ�� QH D���$�A5J�| �rMڀv�X�<�S؞4��/�3H0�J�D�[��A�6D��P
X{�>yzd��+����f(D��SFfJ�3r���:Yd�Y���%D��U��	jO~|
s�@�-����6D�����!=�ԝbŲ�ܫC��"�!���!�jaQ���L�~��CEϟj�!�D >`�P����*�.DR��θ6�!�$Ҧp�&��b��E.<HЧ" Q�!�d��S�F}��'�=s��	���+~!�6����Ğ�U	lRR@Cn!�d[�:��yi��]�LAY6a��]�F{���'�!��/�	T����'j�H��'�PM��iMkh�U��&�#�Ș�'�,šg)҄��ݹ�^fn�8���=�JHɇL�7KJ��"V<z���}�V�s���5b]B�.�>J��$��qA����m�{Ա��D�-kD��)��\��L]�l����ʞ{�p��rC 5����o?��"6�RF.�Ȅȓ9����(��'c�0��F�A�cM�e�0�5 5�^�ȓ#�\9�$�9j�LsW�E�Y��Ԅ�<S��ye�/$�lH���7H!M�ȓE�V�.ʦ�`Q�0nջy�����<��� �h`�W�Z�E4L	�J�l�<��JҤ�c��ۼ�6cFf�j�<��*�yK%4�F61� S���d�<� N<���03�<iv瘽_��hS�"O�tc�L����$�&t�D�z�"OH�9Q��S�tɖ� dBd���"OBp��&'E	�dC�#��x#��XF"O��妜�'� ��5�
D"z`�"OJ�*e�Nm��g��R �Q��"O\Y��W�r���+�)�2`t�S"O`\s��D<,��Z�(F9 +�"O������$������"3j#e"Oƌ",Ҩ+���#`�.��"O������a�%�<
$��"O��2��0X����'��e"O���3�|����������s"ON���Db%H�3Iؕ&f\@u"O� ��N��,���D�>"DK"ON�r��ܴ,R�hx1ϐ&�ˁ"O������5�v	�1���]�iK�"O��A���t������@0h�ȹ`3"O�!VD���q�G�A%Bt�W[�<-��mB��R�e'24�Q�P5���ȓ~Wb�]�?�D��O�.Zyn��7�\��o�&%�Ĉ���f��U�������D�c� ��a�(O��H��vO��ґ�Y�>,�0�k��mba��S&ڸ(n
�H����$�˼ "x��-�LKc��R@Ap�뛏$ڎ�ȓ�Hij��O�6�S�g��-����ȓk��L��c6 ����c�PB���X��1���O"t��US?�����D���ALM�k,����5렱�ȓ!�d�q�ܸYZp��� $����ȓq|D0i�%W�t�JY�,Y�Pm�ȓ�H%�gh�$�ty�CX !�D��C!��$�Y�$rd���)X�Pa@͆�ka�l����H��W
�4�ȓ=����dL�7;Ѝr0TKB���%���sL�
pB�B2!��DU���ȓE���[E��JwΉ�⫕��Ĕ��[Z�����3)܌9q�I�\��a��5����FL�DtFY����d�Z`�ȓ4/b���o[� ��9�o�qQ¹�ȓQ�b���(в{��s5�<֐��4\3�^�n��RB;a��t��gήT���' Ra�@�W!�)��H�`]���5)jL�bگ3
�m�ȓ?� �ҧf����S��4����u���K46�� ��&Sq��ȓE��9�c@�
\P,��C�^��ȓl3lQ�'L��둨,�����yG*Xp����ء+������X�ȓy0��	㡃�bոX��/B8e���]2p}äM�<{*��S$��W�����G洭A�ǡy{`�(w�>,����T�⁁�g]�s�4���	��"B�)�ȓ9�����$bx`F�-D��h�2��%�FL��(�f ��i���ڽ���J�EɎ���%CX<��n ��jD(Զ%��}�MH[�:L��<���'�7Hf�����\m贅�<��ȩ��!L�0��'iZ(o7��ȓt)±z0�ݻy�R�+#�F}�ȓ�`(S6`TK䂉z��#!�|Y��PrAN��-���Ԡ�k����ւ}XT�7H"3E	.*���S�? ��cN(���hTe�
��T�W"OAUE�8��؉p��;�nXh"O�d�3b�#�+h�5��"O����,Pb�jƓ%h±Z "O֠�E�L�]��H�� P 'Q��c#�'��'1B�'%��'���'[��'�1�W >nm�∛�a�����'��'���'��'n��'�R�'hH!���<� ��1�l�(�'{�'�r�'��'
��'���'u��y�Ĵ���rd	>Gr�$�C�'���'\r�'���'��'x��'����0�ƐPnYP�QqR�9C�'l��'nB�'5��'e2�'{��'b6�5�\7����ɂ-킸b�'�'v��'��';��'���'�1ZD�ŎS� ��ab����Kr�'��'B�'{�'��'��'5�!��ր`��S͚�R���'�r�'�r�'�B�'�2�'"�'����f������Q�p$a��'���'�'<R�'F��'��'��12���}!�YүG=��-�`�'���'�b�'�'7��'���'���`Ə4���e�z�fB՟d�I���	��H�	ן(����<��ן\� m�N�E+rK	?A�^�П��	���������������ҟ��0"� P�48��>Z18��@ߟ���̟�IΟ��Iޟ��ɑ�M����?�#�&,����		�����!�\1��ʟP�������Ǧap�өe ��&d��6Ph!h�v�:�Xg�V�4���O��FF�y��1C��_?�h�D��O���X��7/?�O�R��/�����ƥ�G�a}ZE��ʂ,��'|�Z��G��Ǡ(�N��daF�Q_Lap�� pL6M7�1O�?i�����&cj&���jL�a�pz����?1���y�^�b>a���R���Γo���sm��'�@�d�ѫ �͓�y�-�O���4���ɛr���3䭚k���Q��(5��<AN>�i5�ڈy�KN�_
�݋��1��+DoO�|��O���'J��'��d�>�r+���M��"A�Ft�J��k~��'�V�Jd,_>�O�T��	>dP� �(/L�B%؂�:�Q�c[>Q
�IUy�󧈟�$�1 Or�R�&T�z�$�QT�7��N��Af/?YѼiu�O��}Cd�)&֘T+�E�
�$�O��$�O*D�ҥa�H��4����v�ĈP�P�6-O9AȦy0R�ނ����4����O^�d�O����h"�Kw�Z�YA��Ă�}�J�L�F,��xb�'����Ă<!��U蔻u��:� �l�\�'g��'�ɧ�O���E_&HT)�p�ۛh����@�L<d`�XP�S�3��`ER�	Ly�畧}_��mɜ4Z]����!Zk2�'���'1�OK�ɔ�M+BmV-�?AD�͍3h�Y���,�<i��I��?#�i �OԠ�'���'��n�h��[� =^p�`?+0 9G�iL����<�˱�O�V%?���9ӀI	dƐ�(p����ʋt��ԟ���ş���ݟ,�	|����2c�N���e%�_[�		���?��zh��-ש!�I��M�O>��#��A���C;^y�0������?1��|��i��MS�O����HG):�$���a�r��(��?{�V���X��O\��|2��?q��yP��x����U�4S���?Q/O��l��sZ��I�����B�t
رfp������)9��,�c���D�k}�'gB�|ʟ^�ZP*�5�P�ba��_�J�J�Ů-��sð-q�i>a��'Q��$�tB D�5�&l�F�m?%��'����	��(�	ɟ��d�^�D�ٴW�r���d,�i�r
�IP��;��Ѫ��d�O(�ON��<9���v�!r,�
��%����0�������?�-�Mc�'E�i�
�������DC&\��Q��	Z���"��d�<!��?���?!���?I)�b��1kJ7�]��ʕ�Tj@�ԭ�����g�����IΟ�&?���M�;0�&H*�+�<ِ��t��'����?�K>�|J����M˞'3.�a��Q�=����m�Hp�'<j�0q����Ƒ|RT��S��d�f��a���x��VI��A��������ğ��Uy҆��Ѓe��O���O4��0%؛ n8�e�аɊ��3���O�˓�?����Mkh��I��lF^�`2&�I�Ԥ��?Ig$��t@�t!�4�������'�O�5]��"�A�w�$22��
�b�'&R�'"�S��4��%&�(�Ca)�v�z���d�4�D��)O��mu�Ӽ��U�sY����!_�u���<9���?	�SB$�R�4����(U	�D5���>&80 ��@��n�Ӗ�G�䓑�d�O4�$�O��d�OJ��^�J=�p���J �ĭ�8S\��IZ��o��n�B�'�B��d�'����̀�n�(�IB���f�&�;�)�>��?�N>�|JD��U�j�{��K�hs�\j�n�."NŐ�4���A���<!�'��'K�	9i	��2��D�R�B��E��2"l��	��\�I����i>��'�7M =����ԍP#��a�1&F4�$�q��ܦ��?y�W���I䟘�I:�Dd��O��( ����!3���`��]�'Ć��ӏF�?ɀ������� �!A'�5p~$��%%��%	>���;OP���O$��O����O�?!k$#�,-@A%FI�<쩳�,�D��ҟ��4���OMD7�7��)��p�mֹ=F�<�"(ZD�O��$�O�	�C�7-$?�;/�P(ಅV���ś�Í�v�A����?�!�3���<���?Q��?��̊?�b���c�

v���1�?!����D�����џ���ǟp�O��w�� �Z��ƾf��O�)�'&r�'Oɧ��
 ������#\�hB#�s)� " ��!ň7�/?ͧ4W��	@�9z��9��U�.�*%W���<��	ʟ��I����)��vy�Jy���Edֱ&��Ç����#��uE`˓0���dB}��'��@aF�
�H�����H�N�،1�'\�)�����t�"-&~,q�ԩB��|�%���H,E���=O��?��?����?����)ӈ6��K��� ט̚7틻 ŪulڠTEtd��ҟL��d�ҟT!���S��Sz�d�B���1��'�#�?����Ş�¥��4�y"�5.����BL7jђA��CL�y�B��=?�d��䓝��O �DC���9W�F�4(���pOĸ���O^�$�O~ʓ4x�v�J���'�n]�P��x٦��18ع36��<
��O�}�'!��'
�'ԩ�FBܴ�<}��g��@$�ԙ�OXy*��J�o�6��C!+����?�C�O�m+�$�"g�� �2��*0��@���O2���O.���O��}���pb����,G*^L�������=��j��������:�Mˉ�w���jGV%-���3�_�1�&�x�'���'7�!2��������o�+	"�t�1��U�W�����B�m��'������'U��'��'&�1�ٱ4���儨9Gd1S�T��Q޴>������?�����<���OR���l�k@k\�o����?�|z��	�!θ{ +Ψ�l��F�8M���BL����z�l<���3��O`ʓo�r�2�K��x�x ���+��,a���?���?���?�-O�Eoڴ{b�p�ɚA,@`Q-ڼ|�Rm��Bԗhc���	ҟ�'��Gy��'2�'?zQ�f���-�݂�@��:�����lt��3O&��U')`���'[���?���
e���Y��4:����R��4{����ܟ����I��	|�'e����70y����� !��	I���?a��46�&S���I�ܦ�%���5aF2!�^M�eH�X��4pv�Pz�	؟��i>��g�����'�b���)uچ��)4y�LL7�r�����'��i>���⟨�I�bL��:�+&=��1@a׫Yk�'�^��k�4� x��?����Y�&����4scМ�ţ�'&D������O��D>��?a��־>��9! &�d��v�FPl9�A������.O�)��~��|��@�\I �!��S4)���8$�Q�?���'�B�'���4\����4j�r�r��2�zP����,�$���1�?9�c��GZ}��' ����o� ce�2F��X�pP���'�n`�jL�?�!�T��U�͘�n�2p$M4p�\���j���'4B�'
R�'�r�'�哵U����W�ٶV*��+P�f���MS��p�Y����	ԟD'?牕�MϻU�$t!�� �+��Ի��Z�Z�q[��?�J>�|ff^��M۝'���HN�!&�@���v��Q��'��BC�t���ig�'BzT�'2Zwv�I��0u�t͌�bH�8vk�Lq1����4(�U�qk�O0�$�OB��źK䐭�?����?�%�D0���L��P'���?�(O|�k��F/I�t���O6����OFk̀�<���/Ѥ(~*ؚe6O����`�$`�B��\���?m�@�'���	�{J@HP���0� ��Ҋ�
L����џ�	����I@�OR���K��p��իxKB���"_��Ҵզś�OZ��R�)�?�;I��=�	�f��I;Ԩ=B�~���?a���?�B�I�MC�O5�Ao������5Lt�-�*P{�K̆k�"02�<�d�<ͧ�?A��?a�����կ]���d�[)�P��0 ����$֦AKE��ş����X&?��I�{&�y�@��o8���p�!#
��O����O�O1��	� �3wd� ��6hJ@�
vh�z 7�~yBV�C*��Of�O^ʓ+�a�6�C���b�g�+�(�����?)���?��|�,O	m� f�T�I�e	v�!� ��˰!�3��5̓?�v��A}��'���'�f!I��Y cK|Pp��P�J���V�����d+� 9YM������֜���PNpt�[K���3>O"�$�O��Or���O��?ݫ�O�0?Z��1��	�l�a2T����I۟,8�4(زQ�'�?Yöi�'I��a�-"`�f$X`;,!��|b�'{�O<�9��i��	�lJF��w/I*z��	R�L�A�zEZN̊{�"��`�IKy�O��'l_;���C��������:���':��5�MK'*ڿ�?����?�,��T��#�)�E��E�6@����s�O��D�Ob�O�ӲMY�Zĥրfe��@$8N�(��Ɵ�N�=i��=?ͧ�����;��}��,1 h�%��8a���:]h���?����?a�Ş��������I�u�~�A�L��z�e(%A�h��ܟ|�ߴ��'��듔?���*�4r1�_7v҂����ܿ�?�r��4��$�
3�B���� ���J�Q���p$��4O�ʓ�?	��?���?1�����Zu|t�Z�y�nqۡ&Ю�r�m�5@�pM���4��\�s�,����ˤ���DKaVi�%��GJ��?I���S�'%�4mjݴ�y��M�^z20���f.)�֠��y�'�8�l	�	�l�'��i>��	�H�Ě�S#O�B��X�����B�O �d�O��<aֶi���'���'vDH����f���b��A�aT�-�А|��'?�۟��I�	slt�"�A(U���e�/I��I��X"Q��	�p�0$ ?��')��_wz���
w�,�D�\�R;��D���Z�hT���O@�D�O����O���1-�;2�D�O��)�>A_�(�P#F�X�́��`�Oxo�<wxh�I���	m�ݟ���͒�n�uh�x�nY`7�ʈ-<�Q��ޟ��ן�4��ĦA��?����Z~����2�r�O�kj�,t/��3y��3I>,O�i�O����O��$a�;!gC��mc�(j�k��<�T�i�pX3�'er�'���y¡�:]ٲ�0���H>� �EA#^��?�����S�'�P��!ȮO�����L8}��}qE��M�v]�����.(��3�D�<�㣃�j%��S��8\�P��#:�?���?��1ǜ]�'��ئM�'ޟ�C@�P'v��f�5�킅A�����	~�	���'V��'��`1�F��!��^��<�3(����Br�i\�d�Ob���"�*���[���S��]+b�٢P����?{���ĥf�(����H��ԟ��	�,�²Gߔ(rYZ�n��^:tYw��	�?���?���i�J@9�U��ߴ��!���
7�L�a��I� g	=NK��J>���?ͧ!�=�ܴ�����
D����ǭ	�4�ղ�:rN���䓺�$�O��d�O��dӾ&d
<1e&J� �i#�Q	�|�d�O˓a[��&T�2.��'�rX>�8U�5V�fE�bc�n��릢1?�U�l�IПT'��'VP|��a��t�-Ѧ�n��iŏ�;VM��4Vh�i>����OB�ON��U�BSD���	ܤ�T�O����O���O1�Jʓuʛ�"� h��TbEaC�?�y�&j-r&�}�&Y�@޴��'���?Q�ǉ�F���&-��R���F���?)��,�.}�ߴ����48�MS����&=!����b�@�-���yrR�@���l��۟,�	֟��O�du�D/F�:�H�L#z���U�q�H�����O<���OV��:�Ҧ�S"6AB𡖧.j}E�I�>��	��p&�b>A��֦��|["a�o�=��p�1$��_=<�͓��Mi3����'���'�B�'2�[��ϭ�� �`�j�&���'���'2X��ڴ&�����?9���vLI�V� �d����Y.�ܬ(�B#�>I����'V((�ԯ�*>�j����n]0 �O�ո3(ސc��a"0�#��_�?	0��OF��dKG9h\,�S!��m� �$�O���O��d�O&�}��GP�䑆oߥ��A�eXK���Jƛ��K�"��I!�M��w��ĉQ��):�#B�M�)@�	'���'P2MQ�!͛f��HiSn
�u���'F�>~���խ��" .U�pA1a�X0'�L���t�'���'�B�'?���%�5�8�1�Ȟ�k�`8aR�(�4[�$Ys���?�����<i`�6���@LP�8�YQɮ
��՟���H�)�S�N�M`�J�9O40t�5Ƥl�F����k8�I���OV53O>�.O�p�������m��4���g�O|�d�O&�$�O�I�<�F�i9F���'�H�+ᨓ��I�%�	�{*�ɛ'�.7-4�I���D�O�$�O��C #��~��t
7�߂\�H�ؠfM&+of6�??)ţ��q��|J��y�����E֜8��|���=d���?��?���?1���OB~�����)X����w��,���x�'m��'Xb6�H�/���NЛ��|�n�7�~�`CL5n$Z�
S�3Q��'�R���g�/4T���������/W����3h�84���b�lȇ2��zU�'�V�'������'r�'1�8���E�� �E�˨"��*��'g2_���۴{¾!���?����ID�T�4�	�\)Y��[PC)tj�����D�OD�D"��?�:w\����C���P�Z0q2f�si������覍��tNRr?�I>'΂�!��c�$�s xX��H�?��?���?ͧ�?a`�������!h0�_�[f�ׂ̇��p$	�w����͟<�IM�i>M�'��ךN���cX�&�b��bᄉ!b�'��y�#�i=��O2)�@i�0�����������>��� w�� [��`���'�"�'���'d2�'���fb�3� �w������4E��Q�ߴB�~����?������?���y�c��"�(��be\�p���%�#*�"�'Tɧ�O\ʄT�i3󄔎�-�6��YR������8��B3����y���dK1g�d�<1���*�k��Zj�0@� j�ЛU��>�?����?�����զU�R�Gɟ�Iߟ�d�?d�Z|#�D�:g���� �^���'��_����矼'����� *�.qX2 H��qMe��ɊU�0L�����5�'*���~?��ZxȱT/�-0梸Cv
F�jI����?���?y���h�d���=]�,1W/��65XF���VB��GݦE�q ��X��)�M���w����č�6YrDB6Đl�Xy0�'���'A��������l�\e�S�� �1
�?1�> )u��P��%8�"1���<A��?a���?����?����a��'-�����D�ѦYs7���	ʟ�%?�I":��c���*aUxm;���'���p�O��d�O:�O1�V�[��Wh&Y���@=ɪ=��mϫ6� �`�<��D��4���D��䓷�؉R�6�87��h��5���t�*�d�Of���O��4��ʓh�&/5x��L�~��E޶M����U���r�fӬ�t��OZ���O���M�:Ǫ�R��1g�@p�ŗK��f�f�4�_&,(�>��]@� y�K�(b��s �օ)u(�	џh����d��͟(��}��3o��i�-8g�\S"j[�Xf��#���?������e�>��4�'z�6� �d�|�V��F��0|��hQW)ϵٖ�O��$�O�i_&��6�4?r�Y=�D<+���5z��hY��鮑����O�]�O>�)O�)�O�$�O������ ��@��9q8%+�e�O
��<�v�i+f4z�'�2�'��S�M��[�m�){Hh�ehP�p��V��Iȟt�I}�)� g:#D�yR@`WE�-�Ai��r"����>7b.O�	��?�e`1��ާ7(�	��'�y�� 	J���d�OT�D�O��	�<��iO~��t�߀O�-��a��4(%�HJ���'�6m$�������O@�C�"]�M��r�MQZ:| �f�<ɐB��M��O��iUnH����î<a�B��Np��Q� DҴ�5���<�)O���3 t���O0���O��4�F�zH�!�Pmy�P��P���	��a[�x�	����O������ܤa�1J_�	�DhQ�*����	֟d&������I�W�plZ�<����V>�	2D� 2�6�H&mA�<i�!��%B��	r�Sy�O�r�M�<�D�I��h�)��HH���'��'���(�M��'J��?Y���?��-[�g8�p�Ù�y�MP$(S���'�듷?q����"3&o�(�eF�7=L)H�aPm~rˌ*\(qx�HC"�O*e�����'jD|K����z��,��kݺT���i��'�R�'���''�>���>r?�M���*-��ԓq����	�M�L� �?i�x���4�v�bG�
Kp��V�Y>p��a�1Ol���O���V&1�6m8?9��)yY����=�䙩��ڪ:it.I�����`<�ĳ<�'�?���?���?�h��|�=��aO�51D��`c�#���ȦI�5�Mş\����t���?E�I՟T`qOU�E��iPp���1���ia-]���D�O$������!;�}
�!�}�k@�X�5��I��PN��'|j�IG��,9�|rX��Z�\ X�p��i�k���[�����p���� ����\y�}�ܕZS�O�Q ��U  4��P��\☐0��OZ-n�[��S��I񟰗'�(bcmB*�� [�-Y:�t98��W�"��6��\Ӆ�T���D��r�S���Ҩ��t���!!g�2b��ɀ)t����џ���ԟ��	џt%?A�	33� ݂��;T��C ��(�:=�	�`�I-�M�E�|����?�M>Q6��=�.����׏B��i/up�'���Ɵ��	�#`��m�<Q��eD���D�}�U�A�O�T|��ǀ�ZN��$Q�����4���D�O��DZ%1y��!u/�#%YV�����O0�R6����<���'��^>!��$�y<հGd�`���3?��_���	��%��QR�c�
��#I(��f9Dn
�`ξ7�f�Y�ă���4�����
N<�O <�sať(�܀��F�κ)9���O��O����O1���&q�� �%[`��L'Uf|�nJ%0|!S��'�2%g���d��O��ԍWE��#V�y�X���'���$�O�x01*hӖ�@������O.�#W�YF��B�I#��'>�I���Iҟ���ş��IU��ȗ���XgH�(��9s��
�c� 7C$����O��D1���O�qmz��xqa_7(�@Y꒎�-@���R�����t�?�|3���M��'�@�ZgK�Z���QQ�^��T��'�����/��u�|�_��	柔�����w���9�H�v΂���џ��I՟(��iyB*z����5ϡ<Y��A�R�)�j�
70�2K�+��!�"��>)��?J>a歐OQʬ �+�)�*�@~b׮S�`b�$�.2��O�|�	,2��J���{�득����$	@�*���'���'��������Y�Z4T@����4(6�P���͟H[�42b����?��i��O�N��-�.ՃѮ���9���32�N��͟��	ӟj������uG��63��q])%��X!���R
'@�%�4�'x"�'��'��'+�p��AUH�e��$G�� ��P�p�4��=:��?9�����<i��J��]�G�>�I�I�s�����0�Ik�)�S8�����0H^0	����S��8[W͆D��OT�*U��?�M8�D�<��*�[��I�`�}�U�1�ن�?Y���?q���?�'��D�Φ���O�ğx���ʴF�bЩ%�
;4�bbw�P;ܴ��'�듥?)��?)�@�W9F!�wj���=����&*�`��޴���Jv�� ���T�x������!����6*�2[FԲP	ٌ���O����O:�$�O@��1��A,1�g	9����!�+
7<��	ҟ��		�M��d��|J�x��|���v�ܫ&%%xt�g�S�AZ�'lb�����wߛ֒�d�$�=� ���F#�B�e�$A��Č�&����~��|�V����Ɵ|�IߟT��W?�u�'���x�n��a������YyR�`� lq���O����O|ʧO5fp�0�&I�"�"ܥ�l�'�b��?��ʟHD��\"rgL҃n�P��AţD�k��$DJ�?����|j2�O�<�M>�!O�6|LmX�
�S�C�
N��?	��?A���?�|�,O�0oU$�[a.J8k�\�W������a���H�I��M;��)�>!�i��q!�#�"m����,[������?����M��O����Y���_��􊆸t%(��uK��
u��Jl���'"�'���'
��'��S�[�t��"�A �e&��X���I�4/��58*O���'�S�Mϻy����-��'���bU�"O����?YJ>�|z��?�M�'������fuT��iK�=7�PY�'z��`fU��,�c�|V��S���B�ԴH����֮ӿpO*�s�EV���	ܟ���my��uӰ
�i�Oj�$�O�0�e�[<A����Ci�g�ڥ�1,�ɹ����O��$-��ى@�* ���qi��*�I�>F�I.��T��L\��1L~"r	��<�	'؅b��u�������,�����	����o�O��/S$)�b��2�D7fx~%Q�@[3�b�q�v{�L�<�7�i��O��.3%�h����V��W�~]��O���O�TX��uӄ�VpJ��s%��ؔ�WHmV�������hɔ�zC�����4����O��$�O���].\e�O)1_����S	5n�˓��楄:`���'��W>��	������&�0 %J�8#	�F��xy"�'���|�O�r�'��@���#T�R���˝���J7���������w)��T���5���<!s	���1P���i"BacB�R��?A��?���?ͧ��Ǧa���ٟHBS�&���!,�3`���@(�$�Ѧ�?Y�T�`���h�ɥʶD��<��l����1_8p`�F���i�'����	Er�O�WM
��0���*��@8���y��'���'0��'�R���(R�� ��Y38�$ ףѩ` ��D�O��$�ͦ�12+ QyB�x��O$P9��S?{xD�PC� 8`qe�"�D�Ox�4�<��cvӤ��Rs��Cg��h�K�	F�T��� �j�hE9$�'���$�L�����'Bb�'��Dz�@.t��תp��d�$�'�Q���4#�9K��?�����)|���!�#S'�Lz@�9iW�ɤ����O���.��?��"N)/�̀���*`t-AV���L!�-�Ӧ%����v?�H>���k#��`�O��|k��#�0�?!��?����?�|r-O�Umږ{�`�X�CҢ$H�K�*֍EW,MJ�.�ʟ$�	��M��/�>���gN��(�)#<�����
+Z�<�{���?�צS��M[�Oi������M?˅�X�p	 �Ꞑ{����bv��'C��'���'F��'���>����,�$���F1u�(]ڴC-|!���?y����'�?q��y㋢!����%Ϥ8#V`¶�K�>���)��07Mc�(#��жf&�2��_R��ACT'l�h�e�)R�RiZf�	hy��'�"�[��r!K��N����UK�sB�'���'�	��?����`�I��h	$�V�RAhG�U�1/6Q�w��W�/��I����Ia�]C���K	j��֣�%Veb��z�0���&t��X�|B�-�O�X;��T5*��pB�y<�`VAļh����?q���?i��h���!/'B,���-5�A��H @���DM��k�����I�Mk��w��(Ai�21b}2�x�Ṛ'"�'s�G��1=�F���u ��}|��Q� ��1���ϛ[��"c+�F<��O����O�X�+�3C�fXB��M��H�P���A�48G�A�*Ok�i8��l:���F�� ѐ̓�B�)��D�'��'�ɧ�O����%H�-K`�d+_��a2�I�	��<	��eI��IX��ry�A�}
^e�a`}���[0קZa|�Cy�p��@�O��ɆI�$�r�铭W6O%�1Odn�l���Iϟ$�����[%J�7h��@�r�H�l��S�ʼl�t~r_��TP������+G��C�����.\>��1l�<9��o{���j����a���f��.O���ɦ%z�&�i��'��%z��ܒr:]��'[R�KR�|��'��O��(�iq��9~�^HA$T8͈�_ ���i@�D/��<ً���?0Ĝ���m�n���Ə͖�O`Im�?�� �	�����~��+=)����9u@���+���D k}��'�2�|ʟޜq�D� w��q��JF��%k��Jv�P���Rl>��|r��O\��J>��J�r��%ʓ6��1�d��A<ag�i��}�E�¼}�rt��&�°1�b�$^Q�	��MK�b&�>q��S�Lܻ�AQ;s�N}xçS���A8���?y�L�M��O�dP�N���U�JF�4?Jf�b�#B+]IT{�Hj�D�'��{h5�ź�!T|�4@y���o�Z7͐�~<��?Y���`��Ι� ���Z� گ9��!��HF*b\���O��O1� ���v�
�)� Ν�!&�3a�)�lX�L���F>OP�1���~R�|R]�P���@�󬌦p�����
B�%���T��|���d�	Jy2�{�d�sE�O\���O�t�#�U�
*�d��CȪq��5	ǂ.�������O��D)�D(fS.�z��� e8�B���<��	1�p4�AJΦ��|㴟���!cBp�b�� 4�B�������ȟP��h�O���R�Cs�eP�'̜94����!�? ��Cz���s!��O2��R���?ͻ|G���!�X^\��k��/�&U��?����?�΀�M{�OtŪ$�.�����2T���͊'�����0x��'�i>��	�����	R�p&f��AF̹�$ټf���'�z7M_�7���d�OP�D?�)�O&I` �ܧGW|%.��dI.<[T"F}��'�|����7q"�] ��]:#z���-+Q�y��ic��H��p��O��O��sA�@����E����ak�e�̝C��?q���?y��|�.Oz nڎ�̕���5貸
׮�$�vTH��F���ɫ�MC�R*�>����?Q��Lq����^��}X ��H��x�ω��M�O MR5Ò�(�6�
��`��G� (#��W��$�O��$�O����O���5�S>A�xxH�?V���B��8NH���ǟ��	��M�VkB�|��u��|��Q(�@4��]�T����	��'������ϼ	Û���kt
�Pe���`o�S� p��o�%Xl�A��0��Հ���;�V!Q�e|8�3�Yb��#��0�7C@(U�Ӄb��c]����X�������(e.�kD�8�Oб�#�ŗæ�B
��I	�c�!�;9VdQ�LK�1�Z�����x�O�7�����@�X�j�j؂9��i�A( .s��\Bg��RQ� R6�ѫ=��P�t��8*~�V" ?S��{�/0G�V��a��~	Z@���ڽ)���ӥ��+���pp��K��]���>gb�=BiyG�qa�k���M[��?i��D�%��E��.`�H�����d�'���'������?�Q���19�J7L׳E�(ܡ�#�צ�'��[%�nӮ���O��D�T�է5F�Ac�`�١W�V"������M���?�s���'�q�h���ų�n��>>�
��i^�\q��p� ��O���蟦�'}�ɱ75>�����4���bDׂ���ME+��?�O>����'���
@C�,vn^Ÿ4�q���`�el�6�D�O��$�,-.��'o�	П��g��w��?^���QDF	���Ԃ�/Qc�I՟��	���oE�XD�A�5��qc0U��M��Y��LڗV���'2��|Zc{l�rf�(Ģ����%�0�O��@5K-�d�O��D�O�˓Ad���DKTp6�!���G��HV�xM�IHy��'��'���'�2=��f
2�t�P�I �=��(`�	�sbrX�x��ПH��aybc
�v���<	dz(`��UB�p'c��<'<7-�<�����?��(3�,�'� Y�#GƔS�d)!���O~�d�O����<���ײ��Sȟ$Yq�/4�X�R���:%vm�d���M����䓯?���Hwؑ�����I��%C��P��#��+��ӳ�i���'c�4E�8	������O��I�0'��=� �@�H��59�
�,Ҫ�&���I֟܂�*�p���do�&(�]K@���BJ�+C�O�M�,O\�Aj�٦���X���?�+�Ok,�##�$1�@Or1�Q����i��v�''b�	9]�O��>���dT8�HĘB��;W)j��BEl��I���ɦ��I˟T���?"�OP�=���P���YM��`���iT�{�iCꘓ!�D#�Sß�(�$�+����3�J�5{VD)E�9�M����?���leNDxБx�O���O�p'��`���k��#B\v qհi,�|��~Γ�?��?p�1NP&�Zu���UlLL����T���'#�894�-�4���(����Ա��jU�
��$B�A
�'����Ey��'���'�趝��EX����a�K�	+]l�¶Iۃ���?���䓒��DX�P5�Xy#ǆ>]:@���i��Q������	Gy"G��(��S�(�DU��H��] �eÙT����?������4���(y������;Ѿ:Q�t!b��'%�'�[���E ڭ�ħl�~��ޭv<&�`h�D�:��i��|bR��🔦��V`�1�ĸg!�=P�����i�"U���	�y�
t�O��	�?��	LH~��
�LQ���F�qq<O��ĭ<�D�q��uׄ�"��";V-�p(����Oh�S��O����O�������ӺS,��	%*yp��T�FTTy�傋Ǧ!�	eyR%\��O�Of�"ƙ�L}v`9D�^���4�v<���?���?�'��?��!i�ja��N1Y�X�&����䜳/��"|R&��Hy��G]<Z(�2�
�Hc��'���'ގ1�Y�����D�J�H�J�x4�K(P�����o��?��'
Z�bD:.7���t��Qܴ�?�C�M���b���u6l[g�Ɍ/s����q^,�%���aL(?���?1����d�^���	Pa��6%���u�6��eyv�@]�	���	A�IiyZw�B���τ4���B��!_��a��4�?�)O�d�O���<q�'U��OJ�;�F0S�KŌ(��<��� H}2�'��|"\��ʟD;� �D2�"B-nVy�a,?��	Jt�x2�'8��� %�@�4�'�Zt�w�̀���*1��D��`�,����ey��]6��nY��BP�p$n�32ޙF��o�⟌��my2�V,,/��'�?������N,�ce!��~a��b���7>l�듋?��?I�
@�<�����?�g��:ADU
g��H��c �t�N˓?�FD��i���'��O��Ӻ�tc4&fI�J��YA��2�F�����㟰#�e���	ޟ`�IJܧ ���0d�/����PeW*O|�Hn�/9r�X��4�?���?q�'w���ny��.������/'��U�E"�(�&7MH3��OJ���O�O79��ʄE(\|x��M��7�O����O��e�O`}�U�l��[?���8<L� d�'j�J�+�@��I�	Gy�@Ł�yʟ"��O��Ċ�d����D�-!�� ����Ѭn����3�)����<������Ok,�Cy�h	�A2q����P�He��$oV�I�@���L���Ж'WV��hYH1O��'dAKP'��tPv�I�U��'��S��	$�I	Wv�qtb@�#Đ���۵"��"� �����	ҟ��'.��F!h>�B��X�U�cK.!7�T�Ay��ʓ�?!)O��$�O���4;(���*�^d� k˝*׌���[?�|�oZ˟��I՟t��oy2�Dk���'�?a��7�����)jbI�2O^�)ћv�'�IԟH��ٟ��5�f�H��Mf$M�,!��`�;�Ġ;�M��q�I��'�б:Ȫ~R���?��<U<,��Dk�"h�Eg�uϾ�ӥ\�\�����
�.��t�In4�.�|�R!��F]�ʁ�K���'8X��rw�����O~��^�֧u�O�	lDk0eB� vµ��M���?T��<������6��` �P�V��#�]���a7-]�|޶1lZ㟠�	؟d�ӈ���<�1&���!)0�Ԫa�ơ�ll37��6bf�D�<����Oq��U�D�i���C=ZPI�݆n��6��OD�d�O���M�Z}�R���IB?����64��%Apf½okN�S����ݕ'J�AC��yʟ,���O����6E�����hΡ$"����&�.��oҟ���b��ē�?������ f��"�6�;��R�!�`#1
�n}�+�S���	��'?M�`E�
<c$����	���x�+��M3Hۋ}r�'��')b�'�����D;�4m� �Z|�xq�O7�y�^�X��ן���zy�o؎'����<~HFi���fy����ږ3׈O0�+���O2����J���ɨ)َ``��`d��`O�Q�8�'���'��U�<�T���ħ!^q 鑢 �-8qt.��pD�io�|��'n�b���'?(@h#ln���Y����۴�?����D@0-��$>����?M(��"V����5�b�l$H�	�ē�?A��I1b�J���䓒�4M�{Z���`�@�*�^�Mc,O���"������N�$��r��'� 
�*N�a���[u)�JD��8۴�?a�m��������򩧟@i�̀
m�ʵivK�H�����k�@�-����I�@���?�+�}�� " >zL��,ā�BA@���6��\����3��'��ğ��!L�	fu<�q�"LU}��	����M+��?!��a�jU@c�D�O��	"���X�J���Jѳ#��'?�b���D�Fr�I��	��D��K.6- �a�" �7�p2���M���g��  Ėx��'��|Zc�p�+�c��l��ϝ�G�y˯O�Ai"@�OPʓ�?����?I)Oh�����$��6r1b˶NJ,�>�����?���[9������g�xq�D�Q͞XBmS��?a.OH��O����<Y�G�%���e��m�v��6k\7qY��ǟ0�	t�ǟ4�ɭt{܍�U��
UT�/����aBP�~�:��'�2�'��Y� ��J�
��',�,ي��A�DՄH�mB�Pw�4�`�iўD�'��>9�lώ� � ��E�g�����̦���͟���ޟT���Y^���'y��OkvT��D92uFȹ�+����7%��O
��4lFxZw�8�1��	��M� ��8�ٴ����)��lZޟ���ڟ��S����b�R�ȉ>7��⑇G��p�R��x��'ў�O�Yr(�7��d�p� �xyPQ�i�ؠ)��''R�')r�O-b�'員@��`I��\"|5:Ӯ�^��9�OR��)��ӟ Ic�a�ъ��<'��2����M����?���<�4T�*Oj�'�?a�'�b���B�-���Q�_�T1Xq�9yԉO��'�B��7_ܽ�r��c�
�F
fM�7m�O^Miq�]�i>=�	����O��i���D���A'hȘ<�!�\���U�(�	��������Iɟԓ�뀄NtEˇmL1���bբ/d� �'Y��'��|��'���I�j��kUi��I|,�yvIE-0����J�����O����OX�h!��O/n�ٔ�:ب��8tHh�K<���䓲?��s�*��'o��+Po67J�|�1� ,U���˪O0�$�O���<?�w'�=��'|�C�i.^~���K�a�~���iI|2�'H"̠��'Zz�SI�-$�
����!>����p"�%X��(���,�g?��R+�H1��֥���sĈYU�<� 0у-��4gV���aW#�Zd�p��?�Y�Ԫ/hu�"���4P#L�0:yh��S�1�����+�� 4oU�<�Nt t�
�	~��V�{��e+�hKx�D �#�b� �P�iX�������%&Q�׋o�
�:3�fc@@sd�F��$e�l�����U��{���)�ޔH��O����O��D�����M�2l8ԘՌݗ!Ѹ!�Z��� �n�حP��5��	��h6}"��%z�:�۰&�2� ��
N��(��k=��5l* z`B![���$W�����wމA����I�q�#S�}��Dԟ��'�"\���|J���A/�����	��!]�i�3��/�!�dK�w�>�؀
�>T���p��-4����HO�SyZ���G� (�.��V'��{��Q�HK�*�6  ��?Q��?�G�����O��Ӷ�����K��=���V(>Xȹ�C�	�`l{���}@���I0>���c� 9"=��W�ȸ�.F�ft����;7��ه�&f��gb�(ko��r���V�����O��-ړ��'�D�����-�P�ā�p:2�:
�'��Y:gM֝"�(<��ʦ5�@P��yb�>i/O�sr�J}��'ڊI��CT%���o�))�����'-�g@7>���'��I�> ���B��!�@q��Ht� ��	=��H�,$F#<����'��\���	:{�X��sH17��&�� %"��h�l�;/bt%B�����p<1s����@�	Ry�h�C7����J�+�x�#B#ϫ��'��{�c�EI�P�S-Y#!*�h���0�x�q���s�@�[Aĩ)���W��Չ0O<ʓ%a�\�E�i��'��ӣ%���_���I��N�"H�t`P>5�����������Oyn�Y&���O��	�Mش9)B[�m����HІ4��'�6��ҥU�>I�
�n�,"�����nɨ\/ �Wl�+ 8�e����W
|�D�Ot4m�ʟ4�ZCi�4�8��A�%gg�R0pc�8�	Nx��R$�X�rPT%�`��m�}�#/��?ýia86�;�I�J��M#V	ҕ8��Q�H*5�<�nZ��I��pEI%>m�������	�p���U������}�����F�
]��Y�kƇV���	�'R�����g�G�<�ē�Č��H�3��d��#6J4(��+�FtC`̏&^´j��2�,�F�0����y�CG{xx �Q�<��T?
66mCͦ���9N����i>�������I̟���a���Áp"D-���2	@9D�'(ғg�x��mڈiYb`�+0J�p�'�L7�ʦ�%�L����/�^<��L��l���`��Z-gʆ��lE�Z�����?A���?�������O��">?��Y4�<( �Bա�p	j &3�� �-^�$�����V�L #�̱PD*C��	�bQ"3*�
�֬1A�Z�i��a#���O���d��`U*E8cEI�r�]��J q!�D	�|wx�
%L!iV��E��1_1O�i�>a��L�{�f�'Ң��Ԇ�"�ˣ#�z�Ys��$jB�':��9��'��0�����'��'����+���B$V ��{	�+o���?�gj��)1���$�� d�T|bk�B8����O��O���q����<
��%J����"O
<z�L?1R���ůn�`��O��mZ?> !��k� �I��U�o�c�Й&���M����?!+�½��m�O�y��/P2���_����8���O��d��0�<�|�'�4hsP%O�j_�i:W�+V�ر�M�P��(0�S���d���#c��['-'^��9�O����'�1O����aY�q ��8�N�s�$@"O~UӓH�.H�h��-T�zn�����'�#=��OP�%@ h@'Ú"Tf���Q�~���'�2�'$��U���FR�'%�yGc�  �Y"�I�3.-�A�����5�',L�{��'ܬ +lƐh��R*��L/�����G+����'JV�S�G�g�	�:�;�`V:NV�B��048��O~�F/�?�}�I��	&A`��JO
 t|r�,T0���6S���	�X���X�%��'t:�r��kQ �lQ���'qɧ���<��j�k�6MHvn/Q���s`�2\*,�i���?����?A��j�n�O��$e>�ɳ��0 )���c��<+XΠ�V��nP�C�	�7EP)�F�C*,oR��"��&U���2�9�4�F�\�B�}s`E&9 	"J R���D;�O�Iʑ��1v���C]�I��"O\ )wF-%�9�cA;����r�D�nK�1�7�i���'�@$xOJo;n� �[�c�I��'�2��,��'��Y���|A/rv���N0\�5&i���p<�W _C��8�$���▱e2����B�~��\��	�Yƞ��>��Ǚ�,�K�i��q�xCQg*-U!�� ࡛��T>o |ږ�K)G˂!k$O\l�9;��[�-	k|��囲,MZb��3�d2�Mk��?y)�d��Ղ�O�1D��.dsD��i��n�J�`���O��D�;�>��4�|�'�İ��`�F�vT�
�O{n�9J����9�S��n�E:#�,^�`���?Y�vy�O�\�d�'�1O�F(x0'�U�~$�G]ʂT/T!�d���,���@T�
��6L
9bNax��:�_�|8[�!bg���-G4���i �'Z2ņ�)F�$s�'���'C�w�>E��"��ڹ���9d�ԝ8b��Q"R��y�i��U���%/�
w�½ g�K��'��0�ϓ0ʴ)I"�^�V(��΋�2���j�y�N���?�}&�XqƇȐKȆpj�LϿ21��03K5D��� ���u�8�E-N�a�ƈi)7?�W�)�'}��e��N�	jm�E�Э�;���ȓ{iv�p0A��\�:�CSc�/^Ό��
��y9�������I��%l�ȓf��Hr�O	#���

%��хȓ|R�}3����pe�(��m�('��A�ȓ0��� S�[�҅�5��4��4��[��Q�"[��I�͇?���S
�H`�>����R�@Ƅu�ȓd�� ։^ D��'��$$����m�h�cWiI��l=1%#M�F�bL�ȓ1)Vy:�I�+{�V�AFq�ȓK6(�JóS���H5 B�"L���ȓha����C,�Z�	Vh�	ot��ȓ~����r���J.8�f!5�8��GHh�(���=J<#�M�=�� ��B!h���C�;�J��W���FWTQ��!��+o�5���1Լ��ȓ~J�(f�B_�$�PQG�bCd��ȓtD�9����.���'è1����H��(S��H�B,|��#hh1�&E7)�t�S�U|��9Z���A[	:��a�/&.��ȓ�8��D8{¶Ts�Ѿk�깄�x��)��a��!�
�p��
��踄ȓ{��`Rn��6#���+��i���Z��6�B�/8��1f۟��ȓz⎍F*(l�� 1H�I�B	�ȓt���D�N8	8$�]�u�D	�ȓg�Ƭ0Fb��j}�vn��ci Ʉ�qqec�	\#hUT��Tt�Vl_�Z?�i�P�5�]���>L!��C=px�G^�J݇ȓ0vDbrOބL��/Eg�mK��=D����Hغ\Ⅳд~�:��b�9D�40��"!������Z�\8�&�+D��ZBkē`��գ��E-(P� ��5D���Vχ)hv�+rK�	2}&�� �1D��:��act����_�&�8�H�4D���Ej�6yCgF\ �p嚇+4D����B,�$!���bZH�!P)7D�ȳU��6r��C���"qـ�1D�\G��8�f#�DN�JY�-	�y�G�"BU2���@��oA<�y�O�A�N�jF��
�@��䓈�y�B�,��F'���z1i�.���y�1U��p��I�v{�Ң���y��F=A�D�e��&8�.y�ȅ�LLy������4� 0�.�ȓ)�}K&(F�l(r��C��}�ȓ�j����XT�P�`�^0�F��40�l"A)��=�`��r-N��ч�S�? ���'Bo���&m"ZXt��A"O�鑥�-��	R�k�'z�0�b�"O~�
E��ܔ�g+՛d��Y;�"Op����>	�^tR���qe�a�"O�؂���/l�d�� XK2���G"O�Qv�D+j�^i�G�Q�BQ�T"O��CO�5L*��0�[㈥pE"OQ%�1E�P�& ���ơx"O�,���  �Aׯ��.A��"O"�C^=^��S��5i����"O�U�5GSJ�,XE�ǜ]���f"OԜZ�oʇ_��`a�U0��m��"OZ��7���Y�|�D��T�" "O�ٓvmO�4S���d�ժ'�.5:6"O���Y�wK�1k���9B|�!G�'�љh�o��Ӗ�@N���M�Th%jw$�)iqԡԮ0�O��*�B��'X�H�*\9U�ɗW���jBß�S4'Y�L�����%6eݛ;�<�d�NrdB�	�ud���T�J5H �FOz�Aǆ�H�t�t l���7 ;�����4'z��g�ízX��H4�9D�43r �a6,HB`�+x���"'mL1'`X�Ã& �̐
�/v���3ړMN]A"/M$&Ji	�#ɯl@�>I��$حdB��5�D�Xd �H��q�oZ�B]$x�'�����Rix��a��m�I�Kƌ+��'�����YD��@� �H0`%����Lџ�U�Os�4����]�
 ��,K kq���O�BiIv�S�O֐�����Cۀ7̍�g��$
�O`�l�!�=q!\��<I�
2X���(Х:�|՛��ȯl8��P�&������4O��ȂhX��S3(�R��}0����!=	R�E�u��3�I�$��O�q��U��!g6t����X)=�,8��@ji��%GS��A�h �#� ɼ@��M�s�	�/i�˓ds�@���|ל���nI�(���⑇�����#v�C�@����1�;x�ca�"p���,�a�
l��,�0�N`rC�0y�(Dx"�I"E�� �I.������9���\�|��c ђ?Ld��BD�HN����;�!X�o��l6P�*�ٙ��O��6@��-�+A�
��� �L��)�-(�
͐R�a�t��0Oax��� �H� ��ئ��Ȗ�(�r�zh �O�8�8%p���e�ǵ:D�)P�h��S��zr�1+��9̻7\f�qw~�I�����%!�8��ɭF�,���;n��P�-��ƌ��B�-c
�J��;���|	�(K�I�ƌэ��F6�'�������3��!��V	3��J���Q0�t����
�zxG@��R��I�[4�Q%j��OD8�\��D�Ak�9"��x�,P�3��4�%C$O��1���0sh$�E�A��)t=C�q5�V~�$����wax�o�&	����AJ��*�T���Cu}�i�8�qR��fV��Ҡa�$z�~(�� !LOph�4a�5���C��r$bԭ����]�ƣ?�-O����`��ۅ"�������\J�p�Ê�����t)�3,�^���[8��㢏%}҅�5yȰq�c׃| ��x�l��������Rr�L�E��uc�j]>r��$(!��$�'gl�� �ԈZ�μs�"�,��r�F�N2L����w�� �&��p8�l���%����	 M.�0%cڤ��\д�Y1|���CW:�mډ���/E�Hy8�+@��:�@5�[;I���P���kCM�9w�遅A(�j<Q�E�������8O�ũ�L	&T��p��oߎ-���ق ��/[Ԑb��	z "?i���6D�]�&��t�Lѹh����#/�=h�z�t �i����t�2�\�#NN�;P��
1�P SB<�'��0oĶ@&���� rk���'��6	���戧�|��+O\t@f]X}"�@({�D�����'�@�{��MB��sD��h�
�r& ��gX�p�(O�Mj��8�	MĠ�1�� ���M+:k�(��>D��3�� �v�L)>c�z���6�p��A�U�l xR1〵8jJ�j�Q�DC��H�S�t�K>1�@�	�䗻BPc2�����ʞ=w��|M�;v�t	��SR0|�VƝ�)=�Q:e@�8tT]�?�����M�pmS��I>~"�����3*�x���� =�^���K�MM��=��^��6H_�W:8�����6���LXv��Gc${��1�� �jk�oڜ_��L�f��>������v��Ck;�0���<�Qm�'I+�y)F��m(69Kת�ԟx��ʈ�"4X(҂j��4-���Xk�`y"�W�)"�����hb(����B�S��-�OX`�"��)�ex��I�>"����	�T�Qv� _c �;�j�>dn!�D�Oc�l�4��Y~¥�{�Q�� |�3`�(/ ��+��2p��3e�OQ�F���'��1d��-��a�4��8V$}����'V��I�i�ĳ&Q���`��U��L��$�%)�����<�msC��G�Lmi���2'+���rH�hO�0cD�5WS�M�����	�V�p`I8L�Ԕʖ͆�k{����e8gV4���CU��M���)K�~��L�5���ڗ&έi�ܩeR��?-h乚&ϯm�ҧ���x�#U%r�ݻuo<:� 0BÎ�����H֌wnl�Ak4&����O*�x�q{0)��)��Y1P���T�ʌ�'Ҷ����A�j�B5&�l3�Ǜ�v��iRjLj(8���^�	�R���=�j��E�زD %�Si2\Ot�c6�L�P��f금����n�X���N�Y�'H0Z�b���=��l�L|��(D~����?E��E�áC�'��aC��3&c?Y)�M��S���Q0�Y
����g�z��9ã�.e��t�Z_y����4Q��5�s��;R�	R�$J��yr+W�4�6�"��9$԰�iކ��?�9�g�ÜM�ax�J��^a2�1ta�K��X"�OR�y���,\\��K�dR�Dъ�:Q��5�y�"�6 Mv��w#ڟ/��źp�A�y�
@z�U�s�]�v�="����yr�
��n%2.��W���V�F��y�`Afu��hSd�Q8�U�&���y2���S ��o�;\��ٖ斛�y2E���*p:�ル5��C��R��y������zcܮ'�~��dh˒�y�/�0]��Y��m!��������y�/[#e�9Y�
O���
�M�y2��*�\{�A�t���`V�y"NJ"��5`r��{l5�֯��y�E�(�t���w�*�[A���y2�\J�Z�튉j%zlJ���y���1~�c��\/>y��DB�yB�Z���p��X�jḹ�$Ĕ�y��L��z���(��i�~���ɥ�ybhKvn��(Xf���3�ę�y����-CT��J �̛��ñ�y"(ɱ��l����qc�T��"�!�䆥�T����U������оN`!�$�2�l�93\<���	� !�dL�4�̙�K�1�C)H�!��ɣOnV|�F+V����A	��T�!�D�0t)�	'ꁘb&��(�!�$V�Y���H��^�C�<��%���!�$�� E<� L_
;�e�A�K�f!�D��7������؉\�X�D�=�!��\��(<�c�Mt�I�D�C,
!�D��A���;4�As�����U�
�!��B�v6�Ty'�׋q�[$�՘!��]�h��%�㬘�Y2 ���G&!�d{��1�t	X.q�)*-M#�!�D�$��sM6�� TjϨz~!����3@�� =���{W�إL!��i� Ã�V��,ypN�!��'�`�W$ܷ]�3�mA��!�䏃�<���5WpC�:Y9!�d�f�x�f��8i�z�ò��4n8!��G"<� ��
�6����!�d�(;�rըQ�Ý]��ѓ��(�!�DM�K�.1��ˉy��������!�dҁ!�81@(l\��sQDN�t�!�Sͺ�AT�?Pm�peT	L�!�dZ(�̤��H =¨��fB$^�!�d߾!��:���a� D:�VV�!�d�(p$1�d�X�(bE�<EH!�	L�P�GdD�d���т�^0a!��āeRi�"!�=V��b"�X!�]�Pf� &B�e��������w�!�� H\��DI�\������Y9:���*O���3@#5x�0��R�^����'wz�H$�&_�&����<x0��
�'9�)��ꆐ(=��[��N~K���'�΀kD�_�
_d!�Q��t�JX�'��9���ڋO�4�3��M�Z��P
�'�������(k�}(bM�R,$���'�t|�W!֩U���FaW�J���I�'n�к�%���y���2����'%��F%�O�Ȭ���,+�����'w�P2�>����p�������'3 Dk: ��F�=Ԏ�q�'*�,�%Nž�,�Y��9��'ܼ�b�M�4��TJ���YHPز�'`�y%�ȽHHD��	2S6��[�'������X�(�Z���JI�K�<I�'rjV�H�n��1࣪��4(�u��'NfY�䞼�����&� �'H��� �ףd7��7��;��	�'LΥ"���4Q��(�F��
ͶL��'�p���O�3 ����q�b�i�'L�D����n�H9�J��^}``q�'S���3�
-�t$����U�����'� �i�]1P,��"J�D4~��
�'o���GnhZPP��:���B
�'
4���L���ǭ�3�����'=��S�	6$����8/`�(��'�����@�wRA�g�5��8�'3�e��mǕ���k�L��*#rY�')�M�a��5uQ��i�%�(n��@	�'�~q�W�D8Nh(�J�b�`U��'[�\1V-�o�V�ᐁ0F���x�'�IaP��j��-"/҃7cl!:�'~�T:0-Ԫ�$T[��>*�j���'�T������@(zisd'� N�n�@�'�LAS� 0a��h��,�4D��'��}�D�L	���V`��FJ�z�'i��y��{��%�V!��f�+�'H4�S�G�O�zՑ��is�K�'����B�5�f�;��	�2��a��'��I��׍D��D!g�;zW"A�'�ZE����$��pc�@�8T�:���TyHS��^m��1�bP�<0�`�����X��2c���Q�˸i����ȓ=L��m�H�Z���f��Ї���!A�ؐ�p�BW�ɅrG��ȓ,rLi�ЌЍ^��Չ�~�$Є�c���u�D��tc�o�Uw�P�� q�q!���v�ꭀ�$�vE�݇ȓ#Q���$�ݞ'�:, +�N���ȓi9�@�f�$i�����U_$���n�\�cEI�4AX-#"L�m<Ȇ�S���q"�M�6劷��{��ȓ����� w驤+��N��p������0:�����͐^���@
z�	e���')J�IѬw2t�ȓ60U�� ��ܹ;��
&1�!�$G���Ph`D��Hc<��`n���!�$���쨊a�ݠL2��A�ϻY !���#1dT$����	 �h\�Ӣ�&!�DAo4PP��<V����¡̰0��ğ)Z�6|H$�o�P�#�_��y��r~j�&ѷUxXkP�B�y��C�a�7oN�RԨ̻w���y
� ��QPF��l�V��G
Ȫ�$-"�"OJ�4���o9bt��bC�T�2"O
�)��^�^^ �س뎀;�����"O�}�L̹jP��eY�����"O�ɨ�,M�0+�<u�  �'"O2Y"�b�#D2�iF�F�v�8�!�"O8��bMɬB��l�ѫ�$?��<p""O�#��= ���4E
>��v"Of�:�
�<l�]�U0c  �"O� ����X`f����}ʜ "O���C��
T4#���
I�d"O��⊃8tHʙ�fO��n{$h�u"OZ�7�Q��&y�P�[� `�B�!�Ϭ>�����m�"E�lIq�%�23W!�䑀�j�Q`i_z���Μ�X#!򤖋W�dWo��g��9��E!򄍶<s�0�(�9>T� 	�K���еY �:P�R#(��׎�ygJ�m^�	�C��0�~@;6����y��@) �iF�QUE��Y2��y��'�~y����}��PS��������M[�j�C�%<�8�O�+ y�@Џ|BC�	'"���IO�؄���7�8��hyr��y��w�2Eʦ�Z�W���*�nμct&C�	 p�D�br��Zwͺs�tG2D�D@DK�%���F7Z���bb%D��*������I�� ~#�8Bw�!D��q'��=�𕡦�
y�p؅B3D�d��>S��,B$�=�08�l6D���q"SwT�+ �R0^��y4,1D�j��OR�� p2`�1��D��=D����-F�t6�\�A��%8[<��(;D������W�T�ʆD�${A��&��O�B��;5�Th����T  t�4>�C�	�#�0ٹd��6QI�A���	` �C䉽%pT��rW��p������V��C�	�gN���AA����ƅњr͊C�I�R�T��R�d*������l�nC�	{��qi�,V�tP��D�_�P�fC�o�>����\�_F	weZ�8�RC�I�E��qڗD��?��h����)FzB�I=j|�@E�#��@��wnJB�I,�B]{ �����Þ\���p�"O��{����&��P�Wo*i��"O  �ǭ��1�o��(b�$��"O"�cU()����DRB�s�"O.����*(j�HR���L�J�"O��eȄ>|����CG�.H�u�"Ox �R�E`�Px�E��MC�d"O�yP􍇵tB��JU�Gy��ԃ�"O:�I7������Xun��"Og:��3-3�Vt�u�ʔ,�6C䉗Y�9�6cF�\���K�e��N�C�ɸ:&dUq�,�Uvɛ�k�1$��B剞 f"`a�֮�b�y�H��h!�$ÜV3��E�M�0\��GƧ|Y!�d@yq�D �oA�S��iQB�SY!��O����;�E	�+��2<��"O�@���ҀM<\�t �y�>L��"O���yގ�iw+��lƩc (0D��
��O�L@��L�\}�;�%.��$�S�'b�f!�B�P2[.�x1s���E�e��i4��p�#�6 �r�]9A.Ԇȓ@�0tဣ	�+�^Mav*�1~ه�S�? Xᕩ5����ME;?�4�Hf"O0��OR>x�����T|Jq)�"Od�G��\u����HL��"O�	�UFZ��R��P/]Z
5�t"OZ9��4;>�e�f`�(x�e��"O�������8xb!߲o��<h�"O�ТBĞ/&H�1���`�ZE�"O��)�o�8S�9J)E�x)��"O�T�N�r쌸��cDjԆH�"O �;C�-4!J-�U�]p� �b"ON|{d���3�h���*�8AǸ�Q"O��Hu:��G
�2�����"O��֦"{��x�ȕ�Y��t*�"O��q%�$�V|� *�ɲ�hb"O��zb"����p���
0��"O�ƋSItt�6�f9 u@"O�ƨ ;��;��R�_6,�"OL��r$(@��`ׅ��{O<�ؐ"O�JB	��4ȡ1QĜ-�8�p�"O�]6])m���bDڍ���3�"O�0x�D΃+��8�R,6�*���"O��k�P�n�ҔQS��.�:=�"O=��mJ�d�%�c EBO��"OD9@�38@�K�ƎX߼��"OR��'Y�2@.�2�ш
��+�"O��:��Tx�`cNWp��d��"O��k���(�f`#�-B�,,�(6"Oj�8��'6<�X�Q�0�Z��"OQ��:$Z��@M�+*]�`�&"O��)e�\�[���B�k�9|6su"O�x��@d��XxODu�TP�"Ot�1�	�4���ŀݱdV�x�"O���7J�<=�hM+g�ދr�����"O*���j �a��Kq�	\<�`��"OdT�0�j�X%�f폲�F��y���#^�Q���7_�L��Pi�(�y�n�!��Yd�U�k�6�j�1�ybV#�Z�a'j���1i��y�̖=p�<b��]�v���S1l��y2o��l]`9�bBT�i=���c놸�y��n�>x��M��TB�p�f���y��^:��!2�u�����(�y"���Q�N܋U��@|���e���y�T>L3 <!Vォ%��(s�Ś��y�@�\����G��acN��y"�+�bI��7'��I`5���y��Ȏ �u{���>#��<�4n��yR�  g@�L��U�A(D`sф�yr���.,�@���T��`�&V��yҡ؏d-�Q�b
BN�j<�B7�yr��P*����Q+rή��3��=�yB�?-C�0Ԧ;8zH�!$��y�ȋ�h��d�HB�X���2�d���y��֤�� �eĜ �줢$A��y�Ā�BL�x�d��xz!������y�̘1�ر@�e�3��h��)J��y"��;=��0��?0�C���y��X� 2�i��J�*ǈ,BGň�y��؃4 L]a��>#�`��B��y2$ 8LZ��O��&�Z�����y��M!A��1��~��&k��y���O��9��'�`��:��[%�y�ùmx��N�հTJƉ-�yR��8W�Լ���َ B��PE��y
� ����՟j:�]Rb��`��@��"OPX��&G	K��E	`
��-�ԱT"O9��W��Xڃ�]��M:U"O��@1F�/`�"h̙�2L"S"O2|����)@f`	 GQY���B�"OP�R�%�	B4��ee �l�`�p"OT�+ER���Ԡ$��c"O��"C Q$l!`��^�u5"O�0���1�uȀoW!-!��0"O`E w��r��R���@p���"Op|��JՖ?��B6NS,}H��f"O�
3��h�H��eC>pŢ�"O�i�7�Z�{cLh���ź83�(Å"OpMR��9voؔ��}�<9�"Oj�{n��q���[7!V-e���B$"O��2�O5=����	�����"Ov��0��=M!��yP�6?/�$�c"OD�su�3{��	���� L)�%�&"OP�p��0x�Ѷ̍  � 9%"O���B]ϼ���E2B�7"O��r,̣E��Pԏ�%S�����"O�=�E�AN���tLÑZ�0A{�"Ot��#Aȟ'S�T�f�M#1/����"O�I�b$U/�-Y#��1�f�r*ON$Xc�݀6���&��RlB=(�'yx��!��(6����d)H.V���'N(��%�U��9䢆-AMv���'�� �5�ݿ`��+���b�$	�'�=jăZ�\3��Q���}�(�@�'�nA�鄾)�J�ʵ�X�}��ģ�'ôԹQ͒�4pt0�ǅ�{�J=�'����'*J����+N�@b�

�'����G�I�hR�^�Le��'>���(5\An��O�5�Q�'���	#@M|3�b Y1nC�Ek�'�̜�Q���^Z�y�� �;��2�'�D�*�
�8g�~��CT?&��`��'���2�[a�[�.�
y3�'&�PB蔤0����0��"J�@�'>v�y���CZX���!���2�'L��F�Y$����.�9�����'����-�:Z���`��3�H�	�''���!���=X^��fN���'���q��'2a�ucJ6s� �'��cq�F�$��dH�}����'N�}���ȥ$#���/
{H.���'��r�,�CK���"+�)=۬���'�D����1;͐� Q��0ǐ���'��t��W;�L�xe��,�8�'��V3;�0��0�ְX����,:D�`
�C��E���A�-R"�9@#�8D�����$p����De�G��M;֋2D��p��ڕL����cB	DJ@�Ae@6D���	L���1���9��H3�!D��K�%<.�� �8�ҠP�K>D�<KqO�8FJP�C��0pzX=��l'D��Z֛>���۳BPe�j�ˣ�*D��kင� B�{�mO>YbB|��L(D�HӢ/?f�*���O"4t03�'D� fF_�p�l}�4�*[baك�7D�\�vE�49�V\"eo��Z{~a��*#D�lS�@�S���&�Y�)�*呦A5D���C �$F�p���%��f�2D��[�)��M�|d�deV+O���R#�$D�� <H����<^���*�:�p�"OR)#�F�H8���8/��su"O��t ��X=�Jf�K��$}�s"O�!:#ē�J�n�Z�@Gy�l�
�"O+��Sf`��0�Ԧu
D��{�<bl�7z��*R�4C���΂C�<i�I�uS e3�B�7|��"�K�<A�
̮�t3D���
8J�I__�<a�aBK�^x�1c�{�1zd��Y�<�/%-�P��U�W1 ����S�<���w�����A�.8kŁwL�d�<���*Mf�,"��4C�!4�I�<�-O���u�G��lHq��Ei�<1v��*_m�����"=&J���f_a�<�	۲�V�ˀ�X:����W�<�#���p����W�<��ٔi�V�<!�l,lݚmb�̊&iv�"`��I�<��ͺxT$�b�ʣv�Z�+e��}�<i���^nF0�Sy)@,��J�{�<��l�!Cn��3�L� +�Dn�<�Q�V�О�+"G�!�����f��<�DT�m��b �|��viXx�<a��ĵ%���i�#�D�Z��C�ɛ�p��ޫ>�m�#'#!*�C�I�B����(H�)iy����*pNC��)H���g�|1�Fs]FC���(�0���2{���Q�e�1,l�C�
>pb�6��$O��Є_�0��C�.J���䋀=[��p�]D�C��P��+C��� �	xģ�"MA�B�	� M�հ��5z4F�V�w��B�	�<Q��Ԃ� �8��0(B䉺V���#h�>y.���:8B�I7q�B���+�4Yc���^C�ɝJH��gXt�y�O�sn@C䉪kq�]r )puP��Ä��o
C䉱^�n�4�YF8&處�B�A��B�I�J�$m��c�<� L��*��Vw�B�	EN:�$Ϟ�^��@�A�!V�B�ɨ7������Z>VS�ٻ�����B�ɟXs��i� �N��SBXC�	f�1p�ݨ?�jA��'!f�B�&���u�C�N��qө�/�C�	�j5T����u��X���W�tD�C�.xO�5%F�vO��(A藈;ǚC�ɔ)�
FB�j`M۷�H/Y�~C�	:'Ѭ��i¹KZ���hY/D$<B�	�1 ����*D ����W�/12B䉦���x�E۩<y����oH�w��C�I�1�h-1jT�T�a*���U��C�0�����ʖ���n�bX�C�	#�V@��)uY���"8�tC�ɍB(DQ����
d�n���$�==�jC�I@mص�l��#y��Oo*2C�	-V6u�)�����d@X��C�Dh�Eh8�x!c��C7A"B�	�����PL�� !��rB䉜R�ʁ�@��6$?��h4&D�J�C�I�`��YD�X�(�Ji�FI��.�C�	�7
$���!#k�D9ʳ��(I�C�ɣ}����ⅥA� �CH�0��C�	"t�̢6C��<X��0��?E�B�	�K���q�d�[.�|rF��;��C䉾'���;%��7H��2��L�s��C�)� `8��oѥK�e�ˢcV��cd"O�܃Q'��ap�Aʀt�B�@�"OJ��wmǟ,�ʀ!��� 1"Ovr��AQ�բE��c��t��"O�l��kX).Z2()�.� 'zyA"OF	#�O2��q�]���I�"OrM9�K��a\�q8����]I�h�"Or�CG'J���a!wLҀ-�4��"OL9�';"+�<;7l�N�钡"ON!��Q�r����j��t���"O�T�)�.[�u����1Y�DyF"O�����]a�Z��Շ1���"Ofi3��(K���A�,ɐ��W"O.���NC�l P�׬J�%�B��t"O�M����b�t1��\2�@���"Oޱ��*��E\`�����s�,�#"O��$��r�HFָ[�f3&"O��jvDU8U�:�cT����%"O��A�����4�x"��9=����"O��3���(f>�aP!Q/f\n���"O��KsVP��M0wZ�4� "Oѫ' �3^L�LA�n�} �l
R"O����ȵuH��L,v�B�"O���B ��S>��CL�/~a�DC�"O �� @#�xMku�1��u9"Oĕ�bnӒ(w��P�Ah���"O��)G�@#1���+� �!���S�"O������
zw�$�t/�:@�A0"O����,�<+Ct=���^ڼ0�i>]�"C�+b�ӄP�9I�ɕb2D����B�$�\r���%kb�1���/D������Sm^uHk�)�|��U�8D��0�ȣ%G��ÄmT5�r�c�K3D�8S�aٞgM���T*u]N��D�1D�lj�	T�lq���+{�P�",5D��B��ͻW���O	(�x�S��4D��� A�x4�÷-�2O8�K��/D���%J<6�(�"Gꈸ~>}*�8D�H�A�.C�I˛�>)B����5D���p"�!DN�*���-���2D�X����:$�����3LON��GA2D�<jf-�6^RDv!��GT:��1D�@3%.��X�x���iӒVS����0D��y&HK ;�hpy��\���d)�O�=E��%@b}l��󢞓b�J���!�!�$Ǌ9=	j�B��ld昂� b!�d�.IeL�S�/�Z\Cu'�:w\!��P�)R�9��c�4�\�W��kC!��I�@��ѩť߾]�\}@C#
9m&!��>�.�D+]*%��H£�W��2OP��3K@�}^u�3�Z�:>p"O�h����qTj@��֭p�0��T"OX���O;o�n�VJ�3-� 9��"OI�u�гrO�5�4*�P���"O����ǋ.|��M0~aՐ�"O�)1EÂ*$�����D��K�"O�
���w|��bCdߗ�)!��$LO�)h�cV,x��S��#�f�b�'��D�\क`�e	Y�� �%/&(3!��4� �&��qQ�X;��v!��C(!�|�S�Ho�0d�Uj!�ĕ5O� �'�ޏW�&$�2�\��!�$�%��VKQ�ݮ$� j��!�F������-.טX�)�)!�� �HڵX9P �q����0u"O倴�G�4�¹��A�=BT���d.LO��zD��v�i ���d�!�"O���/M�m ˌ ��"f"O�u��=5��)I���.1��w"O��U��(Y��AZ�N����"OT)���u�T��`Ƙf۞4�"O��Ћ�[���υ*��\1��|r�s̓�0�o�q[��.X���˟`���]��-�7��*`����1��}6B�I�"�1O	t��� 3(��C�I�H�d��%x��A��h�%�C�I~$Z3ąϹ]��9 U��K,�C�	����a�Fϋ$�v+�a�;�nC䉇y���d.&��DP�bX
��=��c���51�x#�n��5�6=�S�/D��b�� �x�����O?�Z� ,D��3���$m#ޱ�1���B����Tj4D���#�,	ɖ�s�b=f갑4K7D�3�������s
$+4�6D�ؐ��3/<���l��$-���4D�\��FR�7�ܐ�mJ�] q8d(&��+�SܧdJt�#��J|�=q��C D�,q�ȓ���
�Ԫ>è1�BN�!G�'�X��'K\h��љ6��t�L&��C�	E.�!@�I�on�,�VG��6{�C�I&y
4Ȣ�JR���i���!tl�C䉈F�ΐڰ.J+0�� �UKܵdU\C�I��,]����?��\ �3K�@C�ɤ
��2��4�(�)#�EC�	~�юO����'fѢ}�@B��2 #HE�B��^{�M`�JO9�|C�I�i{��Aw�׻`�F"�L�`C䉟
k��c6���A�p)*pF�:��C�I�'�|����گ]�f=�N�)���=��':ߖ�B*ҍ�`��π�"��`��ʟ0�<�gA?Y�@e���ҥ�L1�Zy��'2��Qf�D�sm�!��]�'�l	�3MB�hspQ/��Q
�'Q(��ef��UA�q�V/V�~�{	�'� ���ώ�v�P���!Ȝ1�	�'����i4xz�7#;�!1��d%��rsJR9�$I�D�>!����"O���*��eL0*��B��'y�t�bF\ P��!d��a���!'D�Z�V�@�|�jb��p���b1D��[���c8\)`���M�	Z�;D��,�@֭��Bn�Y0Vf�.jB�	�Q ����[�̡s#��-K
B�	!{���4� �J#t�j���h��C�I�I����^�
��2ҮA�:V�C�7w���02O	n��؃,߮!ɂC�I	��`� ��UҰd�	�fC�	&G���4
��t�8�pć�)6�C�I=x�H�iGi��+8��:7�ȬK��C�	��Tp�㜩m]��G�� (tDC�	�B2q#&���|3��� n�&(��D4�S�O���2ġ��/�<p��bS�p��'�'ў"~��@Q�8�
,��0}�ho�!|~�'a|�#�k����C
����CeNC�<�々�R���#���t��!3� �X�<)!j�%7��$a�bP_�83��	M�<���!��E�$��|�a1SN�E�<��Eɰ Ra��Z�~���Y����S�? �s�d��jt�i�?i��m�4O ��\/!�� `ᐣ<[NU�g�OF�=E�dN�7���j#��0l�a��hQ�'R!�ѥJ�9�v)U�JOL��mC!�N/�,������j�����=!򤀲S��y����v���päT+!�䙲R>bu�f�Y2k�5qG͇�E�{"�'��I�w����&�R�X�'̦8M��,E{�O���ɮ?!�r�u�\҂�-K���)�W�U��D��}!��܎N����'I$�Ï��`	��ъt쨝@�'�,Hg�_�{U�`@��W�sʐ�0�'ΰH
���~Y ;������	�'2���cΛ>��!�B�;��DA	�'zP 0G
�A�l��OQ�QZ�<�	��yB�H>A�L��dD�}֊=�'阬���hOq�<��eO<fF�� L�0�b)P�"O�Hk�`ۄ4ĸ�ۧ��`%J�i�"O�iH�B�<`Dq����
8Ty�W"O����,b�vHɑ�	�T)�و�"O��{�� '��`��v��{�"O�Q�#(A[+���/�%g�X}k�"O��f�"!<zU;d��.m��"O�(K�#��Q�͜�sK5�a"O��R�@�zD1h2��2t`$���"O����ׂ�~����&OT�r"O� Zpgʹ`������Al:��'��à$��qaT�m|����|p!�Lg�p����6��
	vi��'\�O1�����O�U���n��D�4
��ܸ��O�=E��&�,%21��*~ж�*w	'
�!�$^+AJ��1%1�~�`f��n�!��F�I�@�z���(8�D�k�i��i��In��(�~8q�D�C#8I�䨕
#�Ԃ�"O�43'&W��DyF�"$��e�V"Ofy�'T*EH��Q[�.���"O,��!OP�,�\eyc�*)S��3�"Ol�8���Yl�ɦd�EP)P�"Oԩ�T�3|�)Y��Х0�|�:""O:�[�N�?/����>8:0p\�4F{��G�Z��}0qȊ�.t:��e!>Y!�D�)t `� f�9ota4�єRh!�@[#��*m��z	E�^�6R�"3O����aA ~���c�]�М A"O��!R3�D�y���5\}`6"O��8D(Y-j������N-af�q`�"O�zF�d%���G�X	\[<mRp"OR���,\�$Kt���k%lRZ��"O���2A���*�fC4!�7"O`�J�WM���ZUI�>U�,V"O>��@@P�"�0�	��a{ "O� ���ܡn������;A�x�"O4$
�Aԇp�*\���"���"O���ES���hX&�Hr��-���IR��v���W���AU�׶�� ;D���E�&Z-��1+P�"`u�H7D�H����qp2Ua���x�,��r�3D��iTo��vQVX�K2#���s�%=D��:
���6j�Y���BsK6D�y�_`v�q�Ꝯ���bg4D�`0�Ȥ�8m�@D�(t�x�RY�yr O
Hl|1�A��)}bj�*�0�yb�ُX��"7���_Uv�:����yB$O5\�����8a�Hr@�*�y
� B�Za�E�B|�I�B����W"O�U��$����PШ´ttd
G"O�8rҏT�k��� '�E��"OtL��Ŕ,	�s��t�.=*��|��)�S�7�������<g$��ғiרb pB�ɱs�a�*|��Q"Rœ�V�<B�	*KLd����6�Xh)DN�d/2B�	�'����O^�@9��O>6�6C�ɏ1d�(3���,Ni���/�B�ɧj4����Y2E�E%�5{��B�4
Q�	�F��ZA"�`EH�_gxB�	�W�k�D��oX��S����HB�I�lx�t��#S�G#��ac��@6B�	1{x��w)�0s8������W3&B�I97H�D�A��+��Z�MС�PB��#,'0E�W�C'7W�x*3kY�<?B� r1��)VB�^v�r́J�B䉓OLR��T�CQ̸
���fB�	�ln�S@���l�lP���,\��C�	�q�\yd@P�ą��J��F(���?Y���*"ޝ�� �_,�9k���L�!�$Q09�$�v��|��$��%Y~!���E�)iB�+���/ZG�\J�'���Ь�2��L�ɟ� f<�
�'e���s���("D�ʻ!Q �*O4�=E��ʘ<p|��U�+>;@���yR�J?vƈk����J#���cߎ�y�BN	+@!j�=2�2E肯�y�h۽I;&I�-V45�pJ�k*��'�az��A���i9��0�P�JD#��y��/�up��R�6$J��͟�y�cD=1&�x���3�>)�����y�LBS4�k�*�+_	���%L��yN� ���@e!Q����Ö'�y��U�)V��D�?Nk��"�U��y"��/y����5I5ȵ�Q�]���hOq��a[�b��5�Lm�H�$J�1`"O���-������V�Y"ZG(�Ag"O��� ˑtf`��B��<21�jǐ|��'U"�`A�0䨡�q�a	��
�'SH|x �Y%��3�A��T�v��	�'�����V#0&�"$
ڍG�V��	�'��q'�U�8,�BC��p�RaZ	�'`z�ʄ�U�W�Ȩ���6\����'~(P�Ԃ�'��T��ƈ#'�'�eJ0�ėNCt��iF����'��I�'Uݒ�H�KM08��'`T�g�"o��BC�r����'u^�b"G��qJ2�I2-�;n��8�'�h��ʽ�:�"|{�XI,Op�=E�DǛ�L틖KA$4��4�Y�yR�{��pk���B�@ذ���y"KE|�H#uf��R�<
sC ?�y�ƞ�rq��!'�J�R�<s����yr�Z{l�	��y
�0*`�] ��d6�S�O��貋U	�ɛ��C	�.��'&��O�*^h�g��.Y��
�'T����F'j���H(M~���'�J�[�hܳV�	=�x��'�,���AӄP��@��ā�'� �C�#+&R�!�&��_4�1L>����)_s}�4���X[��[Vɍ�%s��s��t���
g�"����Ն3��LCk0D�h�Q@A�Qb<��J�4��Bd�,D�� ��j���H�*r�-t��p!�"OL(��<.�f�0�
\Y��˔"O܍��Lۚ?��� fH�G��܃%"O*��&�t�dy%�K�����"O@t�D�S7{z֑��ק[ R&�!LO�
���>g�H�p�ǎ]�"O�H��RDPR�B�NL%G=.1y�"OXT��Q�c� ��ΩM4B�r'"O8���`�7A�{�lM>z!��'"O"=�c�#����ʗ. 8ڨ�q"O.��v�?On��*@.R�d�O���h�*Y4IA�.��e3n8+D�9D�h9�Ŕ	w���e�	R���E�7D��a�ԾQc��:!'Z�2�x�+��O:C���5�*$�5"V��v%��b.|(C��!HM&�r%�B��X�� �%/�B�	&P��X���&,��h�\�VB�	�m��i꣥[�J��R%�	@�2���&���|>Vy��l=�� ��C!`��0?�P ��)������/.�p @*�_�<AR�%qɮ(���.Rlj<���X�<��?\��)+��]���u�S�Ij�<a�m[HOp�1"��	X!�E��g�[�<ٷ� #D��t��oK�0]�H�A�<��LX#4��yi�JIC��<q�M�z�<yC�p�8s��J8@q��3�`�<���_3?g4����3x{���B�]h<yUD
/���郧�]���	�,N!�y��.w��l[&��h4bq���L0�y�B�)�>��Ţҷ[�>�#�"Y�yR�X�t�~��KI�Wh�D�е��5�O�=C��y��l�j�ȭ
�"O�}"�F�Mzԁ�)�i��`'"O��C�Y�p���4�P1&m���"O`!& ,�"��-�>
=(��'A!�)��݀�G�T��l�$O��G�!�A�.i�Z�ϐ���@E݅s:!�DǸ �%�p�O�h���5,����P��٨t�*9LV1�W�R�܄�'�Y(�*
2+ F��Q-f=p�7"O8�o��!���D�_�G�`��<O�!��'_1O?a��B��v�9al�1.& ��Dh7��#�O�	�![o�l`*�AB�`鮬*S"O�Y	��V##^���`X%EȤ�	w"O:�S  ,�HhY�/�^�p��p"OHX9F�K:J�lT�䣏�9-\�C"O���u���-YK��� "O�E B�:u��hӄ�ͻ?�~YU"O�3�O�^��с��=���c"O�%����W? pP#OR/9�����"O����)��XҢD�tB���!"O����
��ZPxa�q�	[-�t��"O��;W�&-���!�^�4y"O��Y�$?[��5Q�ly|)�""O*%a5E׬
&�ГA�0Z��C�"O�+'L"\֜��w���)΂�	"ON��i��|*	c���q�pkT"On���77<�}P0+
�b���U"Op���/;H`.)N.��g����y�	�2�D����xͨX���D��y��G/YѸ��W���uz05@�K��yB�Y/r��-X�}g�r/D3�y����@&�0}Fr���Û�yk��*���hժ� |`�,{���y
� P��e%
�>�d��=+���@�"Ov	kA\� �����.vp��|2�'�D����xs ��V�B��X��'y��w�s�fe#�޿ �X 
�'��sEa-C>�(�,^�q��0�O�i��)§�*7�g���F�3D��D��L����
���J��둡�LZ��rT.:D�����0ZuB�$*;��!ó $D�D��$΀a�%OtKޤð�>D�T+�9E>�܉#JK
e��\�xB�	-m�t�E*Жr>d��g-߅�xB�	�
�6��M8j�T� �Bg�|�O��=�}�b��w�ԅRV�ѝ|V�E�b@IS�<	D�%|垭PP"ٙJ�z��"�Z�<	��* :8�䝞7�5Hč�<�k]�E�x�Qw�߱7��GC�<YP(0M��Mbv-D.���!Ԡ{�<I&D6_���P�idW4��Zt�<9�)^6'Ĵ�w�Ўm��dS��r�<!�b6ˑ�]�)(F�{�jZw�<�ecA�U�<,I�̑�\�9�#n�<ѳC�0� 1�3�H&p���-�_�<�3�A<h>B�KCa�<ܲk�&�f�<�T�Ǉ+���� Q�rV$�.\L�<�!���_�ܘ�Y.����#�C�<9	Ϩ����O��F�
[S�B�<��!8w:Fك�蝱x-�uh�'y�<�3(��r�t8�&%B�p8�P�<����=�P�P�$�+`�j�CQMX~�<ɡ�
! ��TJ)eB��� �D�<p� (RL��!ˍ�C�����h�<� �� m�|��'�A,\��	{���}�<)e�R YS��9����� �|�<i�!������,�'� ��K�b�<9-�Y�t(��@�e�iR�K�b�<q��99�:���6Dt�{���f�<!��̑Tw|�Ԯj|��eWb�<I�#�[������޿1a�81l�f�<9C���qczAB�N�rL���l�<y�cP/d�zT��@X�i��4�DVC�<9¤��-�4%{b%S鞸2���}�<�i�5@lk�H�	)R8�$ �m�<9P�¸,��i�Is���7#F^�<�b�ľ(%�ͣ�o�q:�0�	C����<I��J!\�X��҈i%j�@�<9�$�����N���Rqy#��R�<)��Ǽ�RLKqg�5a�N�<�vbR�'��%����m��B��K�<��+HQ�(4��̕5"���ʣ��H�<	���s�ڑ��IW�(�J �D�<��l�zB� V
É bur �D�'v�?�٣�ܠM��TcpH�B9DB0�VC�<��mL0�*���6N�q��f�<���E-�؁7"]��F��a��m�<� �A ��5���=�^ɐYa�<��) À͉�Ǻ+t$ÓY�<yң�����A4e��Pc��VU�<�#�*J@��4,y�D����I�'?Ai�n �t���*�T<�3�i.D�0�Uω,^�R`t�W27�*:D����J��A9!�8i�I+��8D��k"��y��s���
�ʨ�G7D��I5�9Ltt�c���)꾈��6D�\9Ae�~0�Td'�N� )��3D�� D�2����h�$�x@Z��v"Ol�Aę�GS�#����d����"O�Uɲ��,� �nz24y�H4D��+��׻<@ �$B�1���k/D��BdaʟO$>����t,� ��,D�h8$A�&\`같�o�<���� D��ʧ����bh��!-����� D��B��Z�
�H�.��{� �a$M?D����b�u�ތ��m�$�\Ի7�=D�R�M� ��衫6Ӏ���g?D��ȶ�E�vZm����","GN?D����H�  �Cu�>H<����*D�d�͋2L�൚2�0t��˔l5D�8�!�B?e��}b �G6ws@U�D.D�`�W�	~$����3�Ay�.-D�����C D0��c�ߧ	J��d.D�ܒ���f5�ܡ��ݦw
kA�*D��#��	��8���r���s%(D� ���cT�0✇
�3�$D�t�W	�G��%3�n�2��@�!b!D��)'ȓ�c"�鷏�-�� r�M*D�ęB �My�%[k/O�\@��c2D�ܩ&���4���9#����+D���ׄNz4pa�R(�M��$6D��@A@W;���Y��D�Gڜ��3D��d$ �����C:xlFq蠨,�In��L#E�LIv��K�U�<]�s *D��c�U26TY��A�G	�]�r�=D�`��%) RY;���
0�(0��;D��(��١��PY����w�����8D��8�CN�|1��b�Ҩ��cb7D���T ����F?t�4D�px���g�d��h�� ���L'����x���(A:���:]T�8��"Ojq�1)�3GH��RnZ5OQz\X4"Oɪ�Á=b_ ��,Q�^���"O��CԧרiJ�l9L�<<@���"O2��`.\��\%za�˦w$��`a"Oaj  E�Bo~m!�E���h%"OYiB,�)&��\�PB�!��Y�&�'�ў"~"�OQ;<'x��)[�	c���#%V��yRA�&U�X	���@��2�*`k�yRK��j��u�r���,���׭�yr$��~�D	����8��H��֑�y�hD	}�!Sp�X�}��M8���y�� � yQRD�	GR|�bb��y�C �7�8�=D;��AqL��y�AFAЌ�t	):�9���y2Ci���b&Â�X���y2�ڝz�XA�%WBxu!��yR��%Pf�,!#I]�{d�s!Ǯ�y"���b�ydN��x�5i4g��yrAԑG.���&B�-x��i����y��4hj֑Rp*Lƴ���J�?a���0?��TK{t�V���p���XW�<QsE�&m��0��3��j�*�Q�<�fGH ;��r_/=���c+�w�<���$ψ�j��p;0(��Ds�<	C(ڵ-�B\��֐r��#�hr�<�C�9�<p�F����}C�"p�<�'�
;�^�H�3$�F)��Q��hO�'GK`��kO.V-2T��Z�ń�Ty� �"�	d\З` 9L�I��'� D"�j��VCļ�%��8O:�|��S�? �-u%[7>U�"^$&��KB"O (�A._U��`��l�3�|5�F"O���%A�L�FXƉ@�}�:`*!"Ob��9&B8���h�_�0��',!�d�����&f0T�\��AJ�"�!򄖈]/��i��D�mvE��
K��!�U�1id�h�"۹`zT���ٛX�!��O���+4	��\Lv�[���N�!�D�R��I@�(J9vP��)_�!�$����Ij4+��/C\&�#,]!�$�?��t�p��QH`�� X!�d]�L��h�K�L^8!qb%�wt!򄝍�����!C�.��i���� V!��P�t����Lْ��I8qF#BV!�$S[S����D�<a�-ԅخt;!�/jc:@�`gџL��}�T�$!�D��euVib`��f�*|INS!!�ĉ^�`�{ o��j��!P@�X#b!���:1����J���RH�G�v�!��Ģ594D�S��q:녦(>!�$�&M���9�fGObvt����9!�Ę�+�3a[:B_�Q�H
sE!���	omp�*F�VD�P.��!򤎈�6���D�T&
E�W-�.�!�����䚱��p��E\��ITy��|��	K=%!����*��>��hY��^9!�ʵSJ�����L�.�p�A�]�!�*\�>H��X3]P� �/�-~!�dRK��%b�<9��s�.�'q!���1J��1�%��l�rtzQ�Q�pl!�\2�Hz�*^�;�ѯ�!o�ў���ӫ1�Z$��ȋJ+��dN[1'ȓO���5fl�X�蝴0箑3�,=�!��G&�2�a���*M��x�$.[�t!�D�r�:�@A�VS�t)�'£�!�d��DM� $���'f�`�!�F��y	��OL��1E�:�!��,U ؒpkVEd'es!�i2ya%͌ke*\��(�*Vj!��)���lִN;���s�R�qY!�Xf%(���dAR?����@V&G�!��в_���[Q3t�脡6B�l-�ȓ6=�\�)-Y��#F��`9$��ȓ.�:|�v��. �[�/	�E�B$�ȓQ���gßee ��$�φ_0��ȓQ�E�mV5L�8�R	�n|Da�?A�Q�.�X��)�H���ʽt؄ȓl9�$f �5�:=�5��6y�Єȓ?���ϒ1�2P��/`e�E��z]��IR�;`S<�d-{�t@��EJ04���;z��������6�ل��z��5�ģDh�M�q#ĉ1֜Y��0����Iإ-�e���O�ą�'�YGN�&���ˠ�L��ȓi����j5+vDK��7e&��ȓw�D�bpnD�*{����e�Je�!��<.U摂���\���j�/g�!�߻e$ p��D>=��t���D�!��,x�qp��'C�\$Շ�?g9!�-:��,�!�<al�єgX%6!!�dO�G���-)r`�!9c���2&!���T�
���&ю,�H����_!�Y�L�s�C�02��1�U�[�!�T	�u�5%�'V�4lUӝ`!�� ��J�-��ad��Ғgԙv�8��4"O8 s�I�R�ZM��/"����d"O��A��G�r~|���ג;���k�"O�y�펳Bd���E�
)�4ٲ�"OҰ��j�%Ed���mPAp"qH�"O�2��D~taa�l�#g����"O2�Q�iWb�j��À�-dȭ��"O(H�e�C�v������ǽk[te��"O>Y�5j�J��� �Π1U^<	`"O^�x��+���S�ߚ��IS"O^X)6$^�t0z�H��,�"U�7"O<-0g�4�����:�`�5"O�QP�a�9 �1R��&�TM�g"O$)��KʞC�J��V��=s�(Aq"O�E��L�%��<8Ci��MU�b�"O`�Y$��	H،��%^�IE�U"OQX �7���˴�եr?�	8�"O*=��ɵ7�VĘ�͌�t�=Z�"O��"���8�`q` /��[|��"O���IW�.#V���Y�LvJ��S"O0��l�T�.�JSA�&V�����"O�P��n���ڕOF�g����"ObP�u*[��0�]
bBp�j�"Oh� 4D�<\�>9�Rd����0"O`�i�bJ�iS�}Pv%ߜK��M�!"O��;EQ�����pj_%!Ö()4"O��P�C�y�@!��h�-�E`�"O�	L�tXەf�?7� Q�"OV�/4XT����l<�8���#�!�	-R��	�&�'<el�3�P~�!�Y
����ʈSZ��Ik�5!!�D��@�B
U=p:�% U�_!�d��2�򌃀� ]Д��N�w!��ԫ)�N��e�#&�"\�ğ*!�D�-�<��'��A���a`���!�6�J�P$�qÂ �\!,!�d_Ql������7%O@��F�z�!�U�|5@�קǎj�@P�K�!��3*+�� ')�	��q`�@��*�!��=��b$�U�L�&�`vn(q�!��
��ʞ�rzR�[�a�!��+	��\�����JHF��l��n'!��m�L8��~م� �\�!��#���M��tK�`\=2!��$@^A�ڊ0�d��N�!�D�0Wp`���j۝6�H�q���#[$!�G8'v�`�@��A�b��g�Q7�!�ĝ!O1N�R&2wֱؗ��`!��{}�pX���߀Kn>�� =D��h���/3�ر�S�L�3V�E?D�蚗�S8/rF�aPJo߬1S�m8D���l9w�I"ċf�vk"�4D��iF��	�٣F�?$��%�u�.D�Ԙ����۞�*�ͷ��y��)D��JRȄ�f4ӥ�
� 
�:�5D��Y��^�+����Q��y�ޝbӮ1D�0
s�}4�L�&S;��usT0D����B#P)�QcT��$&�M('�/D�d��)҄B�ZLp叔-�n	rƋ.D�X6�]Ɣ,c���MzNq� 'D�,0 ��(�@���h�i,Ꙣ�"D�\��0B�&d�#�2���RS�3D�DzB"��!bƊ�U�h3�&2D�H���zabkȦ5t��N$D�� j��5�_�G 5��F�:ʄ��7"Op���MG�M(v=	D��
e�3�"Ol!�� \�A�`2���*I]�9�"O���ȃ7?ܰIS�ϦzCl`� "O �Q�bB�@�Q��+����"O<}������]h���~�C5"O�	qP�8�� ��n�M>U�4"O!seP0zƘEC���kH���"Ov���P�p��0ȥ��%"a;3"O�	C��+s42�{�$�{R�*"O�G�E�.�X⭇�)��R�"O� �M	vG>�8�D�g^z0)1"O2�q�A��c~PHa$� JT"�"O���'��DsF��E���db��ѷ"Ol�!�'�1b�ܕQ����Z�`���"OX�!�e�,��� q���P�a��"OP����H��L���[�D��T"O����+X��@��"(E���"OlXR��(�^D���VB%��"Ojp�(n�bh!a��-Old�x�"O6`�ET�ܠB�
�`�"l�F"O��0u��L��Ys�,�=b�%ڶ"O��DH)K'"��D�H�Qr�"O�h{"b��xe�m�&?հE��"O��W��3_{2�d�9VR���"Oz8꧌R�gp`�4-��=���k�"O=j�V�1u昺3bD6z�	�"OF����Q�\��(Da!uo�`Rt"OV�â��^����E�:QV���"Oް!.�40��=r���S�Y��"Oh}Kdȋ	z5��� �%R:�#A"O�숐�3Ua����J�V,�ػ"O��`��gL {4!'` "�"O�@x�!�!J^B\�7IĤ2v��S"O����ai�KA�Rx�1�2"OX����"s�|H`gGC�zl�� �"O�9z��΁Y
���.+��XR"O*�S����;�� �)�F�F"OH4p��ܪ!��<��b�*��E"Ovh��C\� πi�5��6��`��"O�P�`�|ݾ𺀅R"g��q�"O��1���
���K�$UG�hXX�"O�=v,�85�t ���D�����"O�,k���<Q��� u`���"O�9VbY�09�	��V�`dڵ�ȓJ4а�ݤ/fr����C�>&ԅ�t+8e��C�2�H����n�(�ȓx �P⥢',TRa�NX2Dt��ȓ:!�����{�x�7�0-_��� 7ƕ�#��[�0��E0Aᜠ���б�b��2�l��#�
T�ȓS �PH�#$�@Xr䘎J��e��~T�M��Fa�0���B�@��ȓ:�8��O�-"2a��ff���%]�����,:�Bd��� 6>����YQ<;�܍jZp�W�Ѿxw�)��\yr��/H"� )JDJƳh�̆ȓ$��a�娖#p+����Ͱ8���ȓ,�H�[��T*~���`֯`01�ȓpp	��D�n>�)a��J, }���ȓ9���X�'Xfb���[' ��:A��盀l4^���M�j��5�ȓ/�R��A��(�
�j��k0X��7�(1b�JԧwdT��S���\�2���S�? ����E%7V�����;,�U�"O��x�"�#{9mD+��r}4\ f"O�IR<CZ5���X>g`j�z�"Oح1�(A�Lqc%PX'�[q"OD�s�Z�%n��I��D5��͑�"OrĠV�^�y���I���Q� "O���-�&�,,)C��^�p""O���1��i����wH�+	�`"Oh�z���3�
+��A���]H�"OF%�Q&S�(��I��,D� d��"O����Ηr�m:A�F�+Ә���"O�y`/��v�Ȱ	@BX0��<�"O�-:1C�2���D�L��`�!"Ox��V�ٺ7��P�H���{�"OT�a�n�;E$p�JŨ3���"O
���>:���ȧ�6.?�(c�"O�Y�7'�/�t( ���1�1�"O4t�����!��������u�"O���ωR�~I8Vj
�fy>D��"O����M5'Z��bC	!X[����"O�T�!E�,�����+2E�)�"O��;��B����6�T�U0���"O&D��Eʞt��(tJ �"O�y���֬Ys�-����Y9�X�T"O�����.=y�hK�J9,l�'"O���&��	4{���K�  "�%s$"O�*�ܔ��``W�+���B�"OFp`D��y��()�� �_�!�D��yb��A�*eߐi92���"O��A3!���В�C3���v"O"Uq�n��=E���bKS�.�bt"Oh��a�L#^��j�d�vy�s"Ox�a�@�F}Y���&��L�4"O$P*��R���@��2���"OX�j0.]�p٢�k��)`6.2D��ϓ-p��di��{���"D�l��=>�<��!��8*@T� A+D�P�ŉ�!hZ$�b��M>j��",D�8�0�+2��0��b�E�x��w�+D�0X��	/�z-�� ǱY<��&�+D��9�ӎR�)����6���%D�X���S�7AR�2�G|��(�ǋ5D�(8�n��Tk��17O�j%����B)D��4
_�o9�]YGMg��u#cG!D���E딊/��z���L�Z��5n D���͆�>,&1���=~�v4�J!D���o(?N\��I��vO6�a�2D�ܑS"�@�D�"	�g�F���1D�������R��"K�n�$�!dI0D� �C"�\X�9j�	�y��T++D��cC��$S'��3�I96t�w�=D�@"��[Zi�G�',	��{�A;D�@ɤF�*G��M��L֘XR-PW�:D����hR�Y>r 8`h�k�j���&D���F�,n��bP��(bF��#k7D�X%F�5��8[Ѩ˗*��Փ�m5D�����.}81"�+*ru0�'9D��c�ݘb�6�#���!u8�a�8D��@G��#g��z�)�2]��-*D�`r��E�Z1�MK��
&_NC�	!U�T���b��%v��C1m\�� C�I�a1�Ԩ,G_0��� �چ-�VB�	�K-��Յg}hJ��P�B��@r��S"H�"����C�)� 6�Q�!L"1���)U�ú|��	��"O�`{�NE�ȵv��W���a "O:��¥�m��0�.�jE�g"O��ٕ�]�W�H��-�� �B�J�"O�� �-�}|ıC��O*T)�0��"O`x�I3K��X��"O ��t��C�0� ˑI�m.�y	�h��}�1IC�M�n��OI��y���v8RDt@K�j����
�yr���J�킅,�)A'�x����y�Ha{r8���2xD	J2ߩ�p<i��D]�Q]$E�r��&NԜ���/�!�Dּ%�ɀ)�7l�Y !O�}!�d�?�@���8{�
���N\!|q!��u��<�s%�._�V �퀧4p!�� �(�(�Z0@P�e���j�I����xr�ɴj����)�1L_t	 V.�x/�B�ɡmu� b�HV!r��Z����op���$ ʓH�T� Cī#��-��
^�-�ȓOVv`�!&	IZ��TY*sL��$�hG{����{YR��@�Z�����!I�y�,�	V(�0�u��}E�a��L��y��D* ��$ZЄ�%Q�*��O�yA�\|
�е��9q�8I�M��yRB?z8ň� Y�
9���y�ᆴ��橆3#��R	���yR�i4����|��*2��6�y�`C�p��I�jK�?���y�E�;�Hz��՞FPT���O�y��)�'v���#6�����E�k��Ѕ�}��8�HݱD�	ů�r5�ȅ�E���P�!=HxP����޵m�A�ȓ.s�P E��1$�TY��	�&��ȓ N�q�@���_�(���_�pmZd��%}���i��Ę���C��ic1(̮w��c	�'NnhA1e��r
Afͧ�h�'� 7��>��yR�dA���<���˦6~,�A@D��|b�x��X5���H�F�P1s��c�h�IGy��O�#?�wI�l�$ة'Ɣ�}�J4�b�v?��\�y0�d'!V�%����
����񉯍ē	�$"RdE�H���*U�:�ȓ[��	QC-���2uD[�*�B\Gy��|*%E�3��\�X* (�сB��t�<A��� .�h�� ��l���c���hO?��?g��l� ����t�E�G�c���4��I/WG�A���C�*A� �ڐM	�C�I�aH� �vm��0��Rh����<Yڴ+�	
I4fT-�B� ���0���|��r�S$Yl���6�%@����g�'���b��7n]̠{��M�>�b�	
�'��@��hX{Y<P 4�=+�B	�'آY"փڎK��s嚍2�<�	�'�bŸ3&^)[d̹��B(U�y���2U8��5L6)z%�N>��?��'�Ą�eA��=A&Ɲ=o��'�V��֛+���u�q ���$Ϊ�~��	YT�t�2�8H�R��"��@!򤌲0�J���M�r�'I��d�<L>�O���O��xuAJ��h��c[Z���1�h}�^��8C�'�$���J�PAp8j��%B\nؑL<���D=}�W�\ט�Xt�_.3]��HT*���y2�L�fcx���G�0Lei�g-�O&��d_�}��#&m�--X�h�f��a�!���|$� �-��%r.��l!!�� ���2Ί'��YY$&A��`�"O.1G�\�hB�d�ܜ̺0"OL@C4j�T�j��܉�$ �t"O	Y����J�ȀCV �- ��'��D�"���2l�#e�c��ؼ@q�{��I!C�*a�Z���t��eK�SK!�d�x�q����1���aqOѳV/��b?��B,�ŞSoЩ�A���&4-*���=�	�� �"0�G%S$[^2�k��0jt��{1��C�/�����p�Q���μZ��|���3BH�B0ެ��f��1�gN<N}��z�D�X(i��
DN(���A'[��AB �3n�xE�����L
��*Z���.}��ȅ�B�q���0�!E��9���	}yB�X�� d��9�-y�.�1�yB
ʄz�b:�d�<4�;sϗ+��'F��;��|�v뙍O��wL`��p�WtH<�eCͰltJYؖ�.F*=��W&��'�ўb?s��<eƂ��D�Ű\&�I�!�&��e�>q���e�/7g$���(>�I�T@���'d�zR!� ���O�y�襚�
ۛ�yB��?'���P��^;oi8 ;�E[�y�� &H{ �p�H��1X��:Ua
��?��'�l���mBL��b�I��a1��y"�Y�lx`����i�?��=Y�y�,��Y=,a�J�@DBP.��O�i���޿ �Ό�ef�a�X�ƀ��8j!�ߤD)�#�+��9�T�Ei��( xQ�"|�e�M>b���ƇD�$�ZL1��� �hO?�ɼ�
ѳ�B�72��`̾{;C�ɜ,T]��4.� K��5N��Ij����ԍ��d���2�MO$����(LO�㟈�l�7L�I�� h�^e��!D�\{R�N(%�~���ݲi�8m
R#D�0���
�M�X�c��q�\!aV<D���N[U&���G�f��`>D�A�&�;�\��tJ�j�n��"%=D�$ ��N�A�����Tj	{�L6D���Gn�e���q(Ϛ��q�c6D���E�٦�id�Km���4D��J�7�`QS��U/Np�<��'2D�X*G� H�ʔ(���h�:%crd-D�@���A� 5�-� d�'T2��1!*D���"�R�&���@M
�a�Xc�'D���#��-4��
��m9�ıQ�!D�3�+�3����%���"8�h*D�<+cg\F�F+���y�T�Fb(D�$z���T�ֽ�� �?N��3��#D�H���֫E�Ly��"E+S���1��6D�|��A8qޒ�b�%C�s����5D��g��F�� j���� P���3�O���p��P����R�o��Y)t�ȓo�2� �� :EZ��AX�~"���^�IAg	��ZTk�":M|T����-ipJ�T��)�A�)nn�لȓIYX�pO�<���*N�}���7b(
砙����{�n�u���b��)��pz���pЀU���,&8C$1D��iG�Kwb�+&��=���`�$D�4���n��0�qD�8���8D��� a��a����` ؤ��aN#D��ȳ����P��ƭ�#z�V��F D�(�w�I��>�Qb
�,0����Ǌ?D�� �Q���7���H!JTd@��"O�i��,�,���rD��=�p��U"O�4 w�ͳM���Xd^�z(�"O�BV��i��Xi!�^�`̀��w"O\���#ܹB1C ̐)�r�9V"O�`b�m[8���r�.B)��Ö"O����������Ǹ���"O�8���'j���ĦH��(��"O�ub#^�U���wlU=�<x"O�帖��J�}��HW;5�yr�"Oly"�#�6�T�;R- A�&���"O���@��xj.�`k�V�> ("O����(C�E�!�/�h�y�$"O~��w��jW<�f�@;}Œp��"On9;B`[�\�HY��Oթ
�H}�""O�<��0@�2	�G�Ȩ?���0$"O�\��P��Y���E[#"O�p�c�΢K��j�n��_ȌK�"O�H��չQD���#MR��v"OF�a�A�`Jx��\1z?���1"O��a�b�J�Å�d��Ё"Od�`E�S��0�D�]�Ѩ�"O� ��%Ԯ,v���M�"�`"O׋]�}��¡��_���"O�81��̜p����BU� 3L=
�"O��JwD�+�(;tK�	0P*$"O����,F$J|iI+��Z��s"OP[����<&��G�=��B"O�PA3�^1Yp�h�E.|�D�q�"O�L�����9x���<V���{"O<I�A_8a�
�yA$G�`�T�"O�P0ЋM^�PEB܅"��}� "O��0p��7
jFQK4�W���0�"O�yi�LF�!��y� B0f�Dk�"O^=�C��8Ȩ 2 �F[^h�G"O$ R��gS�-b��>X�p� "O� 9�� �ͱ�F�P]���"O"����)>�,�b Br��yR�	>< ��1��+-�P=@a�A��y�c��j覕Y#�ڮ,i¤�Sb��y��
i����d�Y/Y@J��R��yb`N�X��K��_�΅����y���n���k���4-k�a��yb M;8O`򥣂�[F�#�ր�yr�X�)۷�C�Y(B��rD8�yb��� h ѫV�J�i�Nҹ�y�H37*�;�*@�Jt�t)���&�y��VAD��T烃C���Ǆ�y��+;�B�	�a�",c�t8���y���{-0�A�	�	1�Nd�7` �y2i]�!l�릈
���S�냱�yr:���7�
g&D(1�D#�y����]�U�CD�6"����I��y��Z9��PV�F��Y"b���y���D����V��p�D����y��p�x���ۙC�$�����ybjL�U]��B�N0>���+�y�j��c��1�0p��(��Φ�y2ʂ!ZH��
R�`_�T�'h#�yrώU�&xA�
=^��P�&��/�yr�M<O�,����8P��2�)���yZ���؀$F�C�|��KG��f�ȓ��19�/b󲅹c�G�����ȓN�fz&��S2�I��<v��<��S�?  �0&Wa��H��E`��p"O.`0�IU�^R̔᧊��NƢ��G"O�@�6��m��\	�i0P�|Y�"OȩX�AI�xI3T�Ձ2;FU2�"O�*4Z 7\���`��"��D"O��صF��&:�|��a��mÕ"O�)����?c��-H�aBS����6"O@R��"�x�reU��vA �"OT�0�(q����E��.��I��"O�Q�E3"V�Q;AK�<�:v"O~��ӈ�#}t�yX��P�K�24�"O�X�c6l`����^4R"O"A�f�A< �:]/����h9!�W��	"D�� �ݚa�Z�4!�䁄D��'� ��=bшGF�!�)\T�z$�8)���1���F�!�d �`Xꖮ\�[sj)���r�!�Dٸ	W�(�b��;yz�2��1!��O��<�s�J!B��m��8!��Ƌ3ȸD:�I�m���VBЊ@�!��X�ĉ��I�d�b0���B7�!�C��,q �!F�g�<X�" �WW!��Kr00@#ީ��DK#�֞�!���'��)�g�t�Ȣ�	�H!�䛠j�8	"2�ܨ��ȧ-O�-E!�3�ҙAg�1)��"TL�K�!򤅈{  EV�c�r�ӆ�z�!�^�^ .����\:���W�W�!�dB"%7l�ˡ3lDj����M�k�!�$F�F�UŬ�(�v�cBD�T�!�d�1[ Fek0�*(��pA˻v�!���J8>�'��E�V��O�w�!�Z�t|~�I��D�?Y�Q�RĆ1%#!���Y$�q��('@
����?P<!��.��i����?�����.?!���%;r�1��&�]���0�CE	f !��2s��M�q%K�d��Z�(IE+!�ĕ60_z���H�d8�����Z!����M��E�0��Ѣ$Q�:!�'4���#�JO�j��5ʥ��!�M�a[<0X���5�d��'f!�$Nh��X�"L�p߆ a�e�4b
!�ċ:]6��prB��I�z�Dv.!�D�f>��Ġ�dBȉ��<L!��
B���C#M��b�Ӊ(9!��==g���%ǋ�))�����ԓ%�!�$`R�&mU�f|�T��ܡ�!��� ����)V,/�P��&�-v�!�$E���AP
����@0b&�!?�!���Y��،����U�?�!�Ϧn�l���`M�b�]��ń�Q�!��g��#�D��ʄ�,*�!��]==]Ԥ�U�Tz	�]Z�ݑE�!�Dո1>��d2`��QC�ѼJ�T�C��+BbIN4fɧO�DS&��ē7�|��5�͠e�ŉ��E>D4�鉲K������_#��y���QsLh���Zi���ǅ�<�ʐ	%W��3�^�@�Ld��]���X��O
D��Ђ�BՓ ���'�`ͱU�E+$�����>,��y�\���^��H��!i(��9�ts��f��B���~�����'eC��#�'@1Z���׮���Y���>@z �5̞��ɨa��%fG��3䇠���S�&@���#5�z"o>[����!���ѥ����4��
�@�>Q(��#��V���h��Od��� "Z�<`��Ov���"Γ`Qdxڗ�Vh��|����:I�m�A)^�\=��2�N�����F,0��<�4��Y�0��B�l����(Xh�5`/�����t�٢r��3>����5Ҏd�I���TZ6&�;N7
��C�=n��찀,�fʡ`L���� �x���"{pգ��īf�t!�fI6I�!�$�(I�a:��Q�y�����ۼk���2䛤g]�ǚ���{&*O�Ijv�Іy��� �O�A?bl� 5�8)�~��AL��?���=dV�DJ��Q4i"D�Ao̶z�����&*U�& ���d����~��Z5�ؐG���Mv�I5"L�Zr�J$Rц��e,�--��?!���3.�\e+�j�0Z�*�-��z���ab�"7l�+ע��Qk�t	�G��~��ݹP��b�D�?_��D|�`� ."�ito��P��̲k	���Q='@L�3SkҬ$",H��<A�S�O��v B�6�h�W(0Ј��S�#)�B�|�6��AC-�O���B�IHF�� ��Z|ֈ���)��KXyܘ���.���Ф��$������͹
��K�d`5*D�D���A���x�����2��сr��\Ux�{"��%s���
��\)3���e�!D`R����a��ى��9O��Ґ� "��P@(w�P�I�"O���Á >L&k���(���:�)̯;
�s��B�%6 ��N�E���ɮ����@Օd��+��\�&��D8#�r���mì� ՚A��<t���EvF�:�$��̱��=�O��
��C�<�7hX=d���;5�D�s��0م�^�
@��P1x�"�'���_='lp Ja&�$9RЅȓq�X)pፁ!�y�`j��$����H��4@�aܥ��Mj�!\^�O���Y�h�a�)�����i,�!�$K���dPaē�8�D�xl���Wxc80à��B4���F�u��%#p� �O������7�Ў����ڜP�9�aC�&G^��"`��5�[��Ԝ���6�B+
��aC=,Ox�v-�'T6m�8�mx��U�>e��q�%�"��O�miE�4��L3Ta�SI�ن�9�DlR,;K28�s��*/�R�s����O6�R&�%Zs�lx��ɝ,���3�y!��p��O%qPԭ��ꋌ=>�bʎ48�X7��x?$���}��q�,D).�=8q�D@�$��&c�F��'L�>��+W p<jdk"c� �K�LK�gc� v,Bk[ f��+
�ce��]H�'����+��=0��#ǙE�Ź��-�~��#@I7~��}� et4Q��6l��{��2z�:��'b��TqB>D��-��'=4�U'��&�=zG��Xu覭'x-܉ҌM l�O��iSD͏,.
��@M�0M�R�O|j��Y<����<[�4̲��N��Xs�5�!��!>�l���/`h0]�SA���`(R8a%>�"��>����O���&�F�P��%�?{z��j4�����tY� E?W:��g'�)E���h��DߚD��Xc"�9�fȐUa��m�oh8p��V�$�$I2�l>#>)�e��f�*)���G�I"r�Ze�N؟�HV�0�j|�D��m�'�L���j�2@��Ñ�I=%�\P@��d6�)Reɚ&U��k2�(O���9B�0a�d
�~L������(6�j�!�,��WJ����=����G)3�t�q֌G� �h�z���`q�A�1����#<)2!޶7H���$'�'\�|��Ū��=ֹ�3�^�:�q���\��E�#��>���3��O?�� l�3)v�бF)�=n�^��v!Ğ�25�B��j�ɧ���Ǐm�I��eq���WnГ35|�	�A�#�޻DG����'-�ɸ"i��YI�1{�{�ʱ�
�+/�р��
�+�.�o�R�ҍ��ʰ&:���r�2�Of��M8OR�9�2ӬwV|@�'�i��m��x��'���R�Ƈ|By�7)ߘqD`�'�ZA��Z�!h}s��K-֜`�J������;[qO��(�լW��i���ջl��ň"O�}��`�(.��y�e��.'n��"O,����,h���ڴ< f%3"O� a�nT�)m��Ą�<���9�"Oα! Ֆ)z����c�8�<�1�"O>�K0�_ i(p/^�Zxx�#"OF�!5��%%F��"mߏ ��$"O����{�@�ǎ�GU\a[�"ON�1o��Q�@ C��$1���1"O�M��!�l�lt �F�k7�<�q"Ofd!�%H�-�B\He��*
���"O&�*�#��"e�d�J8���"O��mS�*�xs����>۰0[e"O�9���[��x����1s�|�3�"O�cs�ӷ(��a�J�F�tL�w"O怊q��/�����$�uع��"O��X��T�6�	��BŘUi�܊�"O��I �=d�n���>}�i�"O�  �X��F�c�H�� ��L	�1j�"O���2B��Z#�2�M�W�����"Oh��5��HH�h�E����8�"O��b���7kz�L��j���"O"q
T��X���aR��G�8�3f"OҠ���@�d���XÙ�U���"O�st#����iN�j�jt@�"O��Vh�.d������0A�A"O°���	PI��I�ʠ|
�"O�B�	�]v�Sh�z���[�"OfA�D�Rn�^|��G��BL�4JF"O����e�sxl��"���s:<���"OR,3��%V�8"֥R3�	�0"O4} �(����QD�g��}��"O��R�ƿ[K*1�tD��
G��� "Ob��у��`S� *��ͽ�T�0D"O�5�%S�12�H�#�0,h�"G"O�Zw�?:������0Ѐr�"O�=ɆI#aI��%�;�p��Q"O�1-J��d�r}]�goA:�y�l�"��Mɡ��1���@�H��yb�_!�Pi��ʡ2M��@���y�.�W��
�5/H؈�HY�y�AB="�q�[�7��PI�F���y�g ��h���ӼT�z���.�y��A���G�Rez$�%���yR��B���Zt�^������E\��y���DCe����
�(��r 9�y`�4!д2���+v��Lpb�B�y2�N:(Ӛe���n:L��#�*�yb	&7�<P��K�n?P(�rl]��y��H6
;��#T�*��=Rk�1�y�j��-�H�*��P�-����T���y�圴H1�r��#j@��j��yb	��-�9p��7&��,�ҁO�y�CK� "H�ʠ�eC�둄�'�ybdI�lO2h���G($�z�;ѤF;�y�#��2�$��c��N�������?�y��U�$x۔$$Bp���F��y��Y!T�ex&ȂC�X����y�>Rpe��EX�{�Z�y2�4��@�ɢOV�ȰV̞��y�J����8%�OL�=�����y�R�h��z��CP�j C�yR�3G�z%���]18�&@��ݓ�y�B��yC������h��! �yb��9$�$����U:��![�cJ��y�����eXM������Lsg����' �@�)�b���#`
s����'�y��y��B6IE�ocDx�6A֨�yB�D�DGSj�ӆBR��y�ȅl`rEC2����!11��3�yr/I�B�V�c,�f�c�bN�y��ݱoHV�qǈ���mK򦀖�yr� �leBCND�}D-����%�yf@��,9�Wz�<\ĭ��y"��g�؇��6s>�qk�MC4�y�&�5|:!p%(W�ib8����y��f�P��#�kp8�1�E��y�N�-j8��D�dW��bm��y��=J���&U��`Ep"�J��yE�6#���hD&ÊՌ�p����yR�@/`鰸��MƘ�R�#����y�T�Z)��ѣ�٨Ќ�O�y
� ")C�A�r(��͝H�l��E"O�m�E�J}�(@��X�M����"O�i �: � �2k�@�\uY"O������l*\k�	�]-��"O��P��4{K�͂�hPV�qs"O 	��D�=�~\� �� 3�x"O���%.�	��`$�M��"O �I�C ����eY"���k�"OZ�j j	�A��iZ�d��d휡� "O0�䐛l��0`�C64"Px��"O�1q��n&Bq�ϝx�lj�"O�!'�T�B2nT�S ݱnj�`"O�m����B��1�ÀByN��"O������`B$��0�*
nD�	2"O$�5`G�+BD��lU9Yn��"O����/L��0��߄iKlAx#"O�i!U��E�����dY�"OĨ��"O ����Y �d!`C�3QM�"O>�ƣ�y�V9��p^���B"O�+�[�&�p�j����-$Ԩ[t"O� ��T�(��9K,��$Lm+�"O���R(��+WB`HAi��^ؤ��"O� �tg��%P֐��	��GZ���"OT�a"�S���sE[�0�:E"OL5yԮ��nN0�4S'�A�Ǝu�<����Z�Z�BGb�Q�IcOX�<�ӌ\�Yl`ũ��jƒL1�IW�<���5#�Z���*X^>hQ@�RQ�<y׃�u_
��m�EI6M��CQ�<I��Ӄ
���*I�G����Q�<�v�	ۮ	C@O5c$��X�+\I�<)�+ܳ1&0�ď�`��)��|�<�" �,"FX� 
���ad��W�<a.�w�druU;W�	����Q�<Y`c� �ƚ7>���ç��I�<�� "Lxr��'�E3,FZM��n�<�eCR�6�@�׍\*h�4E��i�<���E>:�>��4�[2+�x��~�<)Ҭ�4����sl^�
=p��r�Vz�<�v	�c� �$��w�<�aHNw�<��,[-L�@$qF*��1Ւ�,Rh�<1wC�3]Ǽx�u���v����C䉙ܤH�!��1'�ܺ#A��! �B�I(�*�	����d���l�HB�	�� ����2f�i2P(�0��B�ɱ!���Κl���@;3N�C�ɻY.�a5��P F�ڸ|C�	*�X+mئS�Y2��3g�B䉙,;,�{AH��{2|��cJT�RB��9@��t���N[�$�����,XB�	�7� b��n�8��Gߐ:B�I. �P=*AG�bEH�+����"OR\8�.ǐT^�yä�,E�8��"O�%�OZ���D�T�"�r��A"O�U��|�� @��j�:�A�"O�S0��vu��
Rj%�FUBe"O��;Gl0���`���d�8Q�"O��i��;�H��T����b�˝'ؔ�P��'-J	��( O�$�(0^�H<YM�6L$��ZG�ȅ!��1GW���3D�GΌ���j���Qc��Qwji�� �|��P!�	4��	�M�;E,PL��	t��,�1�G�4�9���=(�'�daH#�M�U|LX���f6����H�F�S ��w��is�°^R,��c��U��p�I 4U.B���e�1�ӱ���f��"0a	��Pv�2=@�bFƔXX(HIn�v�*=k��aB����;A�@<tN��b�^�gz��2�'r� 1� jm�E���F��4(UM�/{��9�F\(B�$�H�Q���/\�;c�DޡJN���h�����Fߜ�C!��'h��BG��$oUџtSF*b��KTJ�t��I��dдM���:u,׵��̊E%�2m�  ��m�n?V��.,��A�UA(O`�"@�V(@�I�4� {�z-IS�V��"���udD����J�fU0���$,l�h� W��H��οA���-4Z�it/� �B�	����Z0�2]C@�r._1��x� /ʫ F��E�+��)C�m����
��0^G@��Ү���.�c��HP̈�!ƥk� �|��
f�x�`J.`�-��
��e	����1��!&ۢ��AJ���:NH���3�Ahe�3��u�Ǆ�7�˝$\l"5�D-UG�K^+}�0�)��Df�xt���#��e+t��� L�!��C2�\��7C��I�	��ZTö:��DۖfP���U,����W��I<�W�x�B�;- �����U:�5p�~��K1�VYеk
�5I������"��H��.X���I�l�T`Ҥ�
�K�G^`�z��v�	�FZj�Rӆ�4Qrİ�8P��<�����p	�o����,����Px��ފ B�!aC��*	��q�ra0"�� Zҟ�� O)h0s�@�ly��6D)fL"@��?j�J���!�"&iz���}U� �_�X�<J�V�4@$�7yz-'?�TI�#�,p�z�����n�-K��-�O�Dyc�A��S���!F���뉥y2��AD��>V�����=k��q�p�542x[�5~�џ؊���sP����-K��])>'��Ae	Ø���E��y"k�^7"y`�ѝ&Ru��C1��䎣9 F���E���)§;N�K��hb4�!v��x�`��[�@��)�.f"�aǔ���|r���}&�Xi��֘_SnɈ�l^#
�<��c*D��l��=�$�B��!dH����2�O�)gCIA�7m��+T(pqfջ\��i������!�DؕO�
PS��J(I�P�GC�����#��1)�����S�<�m�u���3�T�kDlk�C�2f�j͈���4hɜ�7�B5+�!KFM;oRT���<a���O ���٤c��Z�a�y��r�"O�P	��
��Պ���x�~�
��'���0�ܯ}�(�g�'UF�kTb�9.l�T�[�>�$�k��υG'"%���1<�0�Q-ΆB (-�'@ `�x��m�9G�p�i�}��CfK�m���%� �\V��U�ETW|��դ9�	�\��{����E����
 �LY�c�5��-�̃/��D3h���hְ��)ʧ^'�%`O��׸E������h�Y �,�K -�Ty���͔����Ƈ�<渐������{$�Yq��J`�3��){��UR�(�#9?f����J�!�X��Z$F�6�S#G][��?q!*�+m����"bp�����=��أ����r"$O �K�D2�0$�b��p�P��`��7<��I�g.I43��?Q���D���*wi>�I��[�4����U�>�=��۞)��t�s%�+��yl�3>�ޜڇ��,#l���7`�D���w����7"_*{ӧ(����� Վt��k3�LY���m�
N
V�XG��}�)��8BDሜr�(�N~��)0�"��	2<�(	�`Op�3�ɗl~H�J�+�\�y8�!�1����$KnxF�t-�6J :���-Q	JE\�%$��B�8`��y��������!���aчiF��I�f�LK�ɲXz�[V���,,��I�ޙkA B�	-�耀`�˙ z�����j�R�' �`c�GQ�S�'s� ��0C�X���9R�W�}��!�ȓ�f��c�n�|�iwcBn�܇ȓg.���t���	�e)`��L�ȓd$��w�cߡR2���IJ�^�!�Q��29)r���� )�i�W�!�dֳm���a�\9k6U���ɷ�Py��<������g�ޝJ�ៗ�yr��'Y���҆�\p��#aJ$�y2	��b����\W��q��GA�y�Ƈ3l$6�b+�L*FQ�q'ȕ�yr�,=c���7.�*:)x�J��y¥ʹuOd����4 �B�G�2�y��[� ֲ��6@�2�����
ƒ�y��B�5�\��ӧƌY��Q"ӠC�y
� \���KS	��z�m["W�hC'"ORE�®E9v�X�il�� [�*""O�x���R�x��ͪiNTC�"Oxq����R�1����Z(���6"O���X�.jmڒC+���d"Ozj�.\�Rz8�b�B�M�"O~�hUn� � ��u���:i�"O�����T�y���!>��A�"O:%3��5t�۳���{? G"O
�z� �w>t��1)PE�"O� r�dէzXT(�ۨ^�*�cu"OR����8J�|���]�e�$"O�hC
�>_m3ԿD��1�"O�Yڱ,I wb��t�Q�J��a3"OB͂F�@�e�$��PS9v^�
D"O,��#z��tb e �H<f<��"ON�[� ɣ=Q���q�r.^`��"OZ���,��5ڲ�].a2��""Oސ�"-�3X�j���
�;r��J"Oh���� �@8js� ?����"O�Ěpj�5s���B$��A�t�B"O"|��2D(�B��\��<5�"O�e!ԧ� #4yPƯ�j��5�"O����n[*ʐr�2�X��u"Ot��dOG,a�����s��"O�9�'T�9�( 谌����Ҕ"O,hS2F�9~t��fN�J���"O"��GO�rT�5D�7Y��u"r"O����n�-j2��򢘈% �}�"Ov%�V$L7 ��"��&35��i�"O��8b�
ẉ�@)�' �Y��"O�-��\�B��y��& vd�ѓ"OZ��ϗ}
T8����!� D�"O��� �v�zW  ��T;�"O�u8��
>N����W�4v�T�C"O�Iƀ2?b�1��]�#otlR�"O h��E;�B�Ӯ�F�N�8u"Op�p�X'~�zm�7L"�%$"O��׃�25����`�%k����"O|�;�M�#����Ϛ9�r0�"O ȹ���e!�P+DP-��lI�"ORy
3.͹��(YC#_Rc��7"Oh,� ��s =3���Nmbm�%"O��`eJ�&�TC�fP�\4#�'"�Ii'�@
T���"M��R
�'R�zU�S����=���@��e�<�ÍR�h.ź&)�Q��ٹ6G�]�<	Pk}Ƚ�bܘ���T�<��)�'g�z�lF�Mt��ira�{�<�p�8���Е���o� ��u�<�E�=��);��IJ�R ��:D�T�$G�;�x�J�	h��R�B�	 g讴�#��'^�x H�-<�B�ɒj� ��sAI
�R�� �C�I_��q�c,Ȱ4��a��B.[�!�5o��A�� ��b�إɡ��_I����9�����J��X
��=��	�4FNĳrh� ���#w�Ef�`Rp��+��� ��߸�yr�i�O��O8�� �("N8��V(@��JL����>	S�&�H�çrb�Q�u1:<������	�ܔ!7�$�	�ސ��S�&� ��iך��lX5�é}�O@ѠJ�Ӹ��O�rt`��\JϮ|�T/IPV���O�Trf��'����8�7(���-1��ݬ1������V	q��\(�M�������w�>N~�8$�	fJ����(�j(���C�1Oh,D���|� �L�e�=\%
�!ciT�w��u�"��4�����De��.XF�$�U�k0Υ꣌ۨ>N�Dps���G�^��*>˺��+O���Ͼ
��\�ㅅt��Qp&\0i�裀i�����8`1��?�?գm�!�D6@��\�L����x�dܳ#���QΎSt�!�ߛ��'	�z�Wn��xV�Q� &E"��yBh�,����$�Ђ/^��a ����y�)�M���	�:$R��Y��Y.�y�*O =`y�3��)"8�A�!�9�y�%�� �8�����):�����y��F?d��"�� :+R���aD��y�+�	��t��/E��&d����3�yr-�09S���:s x�/��y�^l��Pd�ӄ	���F%��y�J�8������՘�PNѩ�yr���^�D=���I�I�<@�7oI5�yR��@�b�zt,��H��q����yR�~1�����99bekP!���y��4��HAF`@�a�m�G���y�.����1���RI�0�g�)�y�iW
T�ƅ�� 7<)�!��K�2�y"��=�,�ɔLVB�U�5oC;�y�����}
D��:c����H���y��Ц}9�H#��Yv�L:,=�yr�ͥT��Ro�1I#��8���yRc0_�`�!�RI��Qa��W�y�$�r�MϠK��� ����y�-ԝM)f��2��D"l[QE�%�yR�. 'ęY&��l	�,8�JQ��y��6�D�@��)h�mȡKJ5�y"�7�ݺr"B6Z����Ĉ��y�IV)�21Yv�U�Mw|���`h�ȓH�$H+��ݽ5W�8�`B�1��P����!�Ds��Tu<��ȓT��[�L�Kd�U�s��C\T��ȓV��Ai���*��R2J�y�����x�I�+U�h�XB�Q*{a���ȓ;w<��5�Y�~5�@{��ȓW���k���^����!�[����ȓq��Hi&FF�?���C�5y��P��U���r�(���g�/9���Uڐ�2v�ЃC����G�,]�fA��%pɓ�+6P�踋��Ʀ���ȓ]N)��%�6$\�6�D�%\0��1]T�CE�@�m�p0�b�Z2� ��� �z�V>j��1W��RM�ȓyR���,�F��a�ԺF�Մ� �� Fm_:dp�C�.W:X�ȓ^�Z��Q�b�ܬ��8\��\�ȓ�������U�!�F�&�����Y�x}"5��$r�$�P�Dɀ<q�Ї�o�e��	,Z��r����t�X��9J�C#	Ѣ	����nK0r#���ȓOE����=���*S8ņ�f-�5��� �{w6����]�ȓa���!�ߣ{�T�a�u�t���]B}�!MBl�|Hr��/ꝇȓu��;V�ϲ@|8��ļkX�ȓ#d��f�		VH��Fƴ1�����zSp)C�썟d6J�	���
�\ԅȓeR<%�VB�6f�ѓD��~�\<��P!��7O5fq��L����ȓ **Wi��N�sP�h�@�ȓ��p�d���d��n���:=��S�? �e��Kl�9�-��[NU""OjZd��x���",N�:E�|��"O�5Z����qă*;C�s4"OJQ���e����t�!.rP�"O4��T������Yc�Y<N5�)"u"O.,��m����e���O"�}�7"O���̘�N�;v�1){� 1�"OF��F+�(Qp�̀d�.T��"O�f��m����a+�K�Q��"O�]k3�^�E�����
ߐT�*��$"O��Y�F�fzZ��i�M���J�"Od��e�D�\`.4Ph1Ƨ��(�!�O 7 �T��C̄g���V�(ie!�غ۶9��F� Å�;yt�4"Ot�@J��q�-ˮ} m;�"O:���LR�_KD	ZE-��1� ��"O����f˜<��l�*���"O9qcE](�T�P�ЂIݜh0�"O�-�Ҋ�0l[2��׭_���ա�"O �7,/�80gȬwrt�S"O*a����b���Ӭe�$A�"O�	3���h'�=î�m�n��!"Ob@n�!yu����40�����"OB)�4��v�u8���=!���w"O�qR��͚4I�5ٖ%�!@���3"OrY�s
�D�ؒ�J��~��a�"O��Cb��Z�ll���8v���E"O�%P�B
G����F�@,e�}�"O���&J�6/0#6�S2�\��"O��rBU�a'n�
&��#zvP��"O��PbÎ6p��単'm�-�e"ON�A��Y���bLK4/k�-J�"Oʈ���	V���rhM0h�C"O�U�㩀�о�2*ީK�0s�"O(pŁN��m�'ę�0H��Su"O���G�R�xcx�B� �%<>p` "O�t���N�T�9Dʞ :3���0"Oryjp��W,V��0*S(,�k�"O���ʛC6*��i�1v�٠"O^��3!F���#�'�|�F��"ONx� �H�R�B����	�_'b�8�"O�e��@[70V�yq&W6]H1 "O�E�a���?�0uZ%�6����"O�rb��N���9t���20h�"O�Q{�b�3�����9v��2`"O�)wn�N6ެ�4G;_^��7"Oz�q&�l P���Ҥ}]����"O�u�+
*/��<䀔*]*��c"O�I�!X�2gj�A3�цvU���"O���Ô!{S��	��M\	�F"O<m�eŐ&32�ܩWi[��[�"Oڵ�E�V�p������
���6"O�}��'�/lH�Lz�f�0R"��"O�q�!$Ę> �E��Fܗm�@E"O4�)��k��%���UkHp�c"O� �욄~��B�=U>`"OH�آ0�4$qv�є(8LL�R"O��Jh�uY��n 5�=�"O�����Ұ J
�С����q"O&���$a�d�Ӱ�Qm*���"Ol�r-�d��Xj�E� /�91w"O�(�[���A"�?,Y�T"O൚u�4Z��Y3�ƭ8 R�"O���p�\/���gc:�����"O� &yY��Z��y۔�U�\����"O� ���,�9 0�E� �.uD"OT��卐	8(`٤3M`"O�=���\5�ބ�n	7%�"1"O&���D�4:�:���^@{�"O*5�g��3O<`1�N?;�ˡ"O\4 f�>��0 ��W-R�G"O8�!"R�f� l��sl�!"O��)���0 ���#H�&�HV"O>�p�� ) �E��W���0�"O���d�@�q�|��4��'��:�"O��"B��6|L���d�zH�(�"Od�9��S+g:@�i���]��̘�"O���D��[�J1Ţ_9{�h��"O�y�蕋 �<x�@@םt���qB"O�X`g�(�n`��[�>r���U*O�h�����9��0qe��^�p�'��L���>\P�X�`�+o�<4�'�:$��
�k�ޡ�w6��iq�'{0�(2�֞=g�a��8A�pHa	�'\��D�h������8	���j�']f�³�[�c=����Y#5���'��I��;sF�Q	��K	Z� �P�'����˘�x��*QIжU�4��'ʲ$�Հ1n���0/�� H�ݩ�'���s�X� *�����!)�h���'� ��(����@�pd��s�'�؜���ɻ5̺0@b�ƭe�HM8	�'$���	\0�p6 �2\��Y
	�'`@��%�&�@z��X�j���'@1��˅|��m�WjK�NG���']�ʚ)T�9���Fv����'�(P� Z�L�i c��(��"�'�,PLYq�$E�獉/s���{
�'�lJ�h�<A�����q�,�
�'�D`��A34���h���>~�>m�	�'�.ᘄf�܎�7��td:��	�'�40���%n�h�������y���_T�=óOX߼h�v�U��y�	�6�ᢷ�� \�*ţ��y� ��_4`���@7,ep�K��y2!R�0�)��L�/J�PL�2���yb&$�
d�T��/p����G[��yC
�*;��A��W�#���8�����y�(֥��骱͘3XJ��M�y�N߇%�n�2��B! J@�� ���y�h�v������*f�Ax��O��y�օLJ��03�����e.ό�y�BSp��d���X>�F�	b�M��y��H�>y
�̃3u�,!�)�'�y�aI$�pݱC�!V:B�k6N��y2K�>����N;S0{�l�
�y��P%��%�b�`�n�Y"�T��y��R	V�Tl:�錑+H�����y������AV�%�j�y�C�y�!�Fw`5��3� �)��!�y2�.��j�� %�p�a���yb��d����/ǀE�������y"��%f�B�	W�_��P%0�a���y���" 	J)�w'�%jA(��ӕ�y2掉x�dC�$U
�Dp��c��y��u��]����{gΤ/Y�:��ȓ5���b�&~���ட�C���ȓM8z����i�|��Q&N	D�N8��S�? nl2V���"��!"�范H��]1E"O� �P!=I&���l�17��"O~]K#��/H�@�X��X�G��9�"OܹاAʳ	6�8����P,�z�"O��@nY�9"�B�Rx!�ɋr"O�\3)߶T@E*f�� Q}����"O�U"�Fʘ��2ta�'Zv�ű"O֬he���v�ȱ��O�7���Q0"O�]I��2f�M��Έ�9��S"Ob ��� C�\�nH'k��ɑ"OT��� Ao}�u,]������"O6�Z&L�/�reꗬߒwrZ�"O�F0�@sEVc4`]�"O\�I�q�P87�ǿR��� "O�!Ȗ   �P   t
  V  �  m   �(  �1  �7  ,>  �D  �J  Q  KW  �]  �c  'j  ip  �v  �|  T�   `� u�	����Zv)C�'ll\�0"Ez+�'N�Dl�l|!9O���A�'j�e�>=<%
�ǁ �pp	�JQ0K%:����V�E���r5掐9��"���H�A��?m30O��?���B�[,L�7nI6r�diq��6j��L�I	th�� 4�"���O7�u ߆d����'4$UJ��´l��̱&GI9�b� Q��v6=I��Ofi���C�oڦ�×��Ӧec����� �IƟ������b��Ld�`@2��4]3l�#&lڟl��Z|�a�ݴ����OV�Y�a�J���O:92�*E�h�M�5�2 @Ѝ��F�O��$�O"�$�O��#��O:�Z��'A��Ə{�6!���=��!�s�6�Oh牺E�x����17z(!@ F�U�,��Oz�	=��90�?1�LL' �z��[ N�H!	�O���O����O��D�O��d�|��w�^��`@��5��)�e��,��<��?���v� �o��M���W���kӐ�o%�M���-`1�(��q@�re�� ,�͂��I���G��^-Hؘ���%r��)����'X�����Kd2H'O�",ڛ�Dk� �o��?��"#�>9)���?��R�I�8:IZ#�O�,$l���4x����W�X#	X,�ɢڍ&LX�C�g͸YB�1ґ�iA�6�DӦѣc�8SQ���"�ʳ[yp�"�+�W Th��
�SR���ݴ��/uӤ9 rټ+W^��#�5_p�+�B���IxA�ַ,X0���ԂB�$h�*'�E���٦!h�4E[���
�0��K�.�|YBe	�PA汘D�űb�TC�'�=V�"t��H~���BFL�6m)jX���!	:�!	�Od�Ё��� 3���^�k2):�I6"�D�O�����:Dn�}��h��@��1c���'o�5�f R�?�,O����O�ӶS�� ���Ǉ{d��B������Ǣ1ˮLX(<=d�B�(�v��Pubs9}��2{P���$6�t1xh߈J�M2�H�R�L��A�@��'Φ�r[rIc�	_i�D�3�^,4�����D�Ix�S�'�y�*Q�ZUd�'�@�o#�Lr@����?�&�i��˷�-�͂�M���v�0&�nӲ��S�� Z���B�K�	��$�2���zC��$%��y�kD�WFܘ�F�n��ʓ��=�y�g��ei���#l��Ysȗ��y��|� �'Ȇ�f�08�W�yB�ݛ��L�4`�s�  "�N�y��޿*�Х��'�$�ĚD�[��?Q��U�����<�t������ވ&Z��:D�(�&��KB��y��$0 ����#D�؉����Ř2�G/I�@i�ք"D�Ę7�T&m0��[ �b��5D�Hd�"$���UĞ>u.U�� D�ܳ"+V8k�� ��A]��B)�<�t�x8����C1d �ܘ�hU� �<D�ĸ&j�=5��#tN�☉�4�<D�D���M!z.~�z��3V6(��;D��,�:B���xEh�[�r��D9D��3ufG�x�����H�e�T�۷�7<O�eA��I⦥�I�XH5��q�� K�^�x�����؟��I#"G����Ο�əW�0�#S�^��y�P�CgC<�cn�[&.s���>��@�O�����Kf\ <w�|�2�]�Q��1���6�JtSn͍� !1�͇[&�B�+I72�0�?�V��ߟ��	��M���'� ݐ��	nh�G-rJh8,Ob�D$�)ʧvf!q,��z�%�5�_<��E{��I!�M�T
߼b�P�+��G��$t�Z�9����|�C��j��``�D�HC�ӯU�irSI�tAV���1D���`�f R�X�I
ILc�/D����LN� ���T!]�V-3#D�8�����3V�aK�Z�-��02��"D�`�B�Rd�y�b؟&}&�xF�-D��ӳ0+.���l�"����6����Y$�p9���?�Iٟl�ISya��Ap8p���֘u�"���@��bô�s��'_$�7�V�j����rk�|RR�d���Ny:���a���b�8Ɇ8���=�����i�>&^c��iQ�y����'o�-����/ɰ8K�Ɵr�����i$ʓ4�Լ��e�矌�I��I��.���¬��H]L��AT}x�����P�~��S ��[nE��I]������e��4���|��'���ߺc��4�	�U�@k%'�61Ξ,�Eg�O��$�O��ī<�|r�! 1n"��2!�n>�@��KX<@�(,{�u�����E�\��y�*℠�r�ـ1(��g��:2���cԈ�A�-1��A�N�y�����c�%���"#L��({�TR��?ы�$/.�ZB/N����pD�Q�l��ȓb[��`/�HHP�CE��6�%�`�޴�?�+O��(Ƀ��e��ȟ�U�:�j��3�X�|o0Y2��ԟ��	"g��)�	���'���s���OO��SS�O�0_��� �8hTE�0z,�b��P��	��'�P0���D��H�SצC�( �����pgZa����nr-K�Q��0<�
�ğLcK>����'v��C%��29��m���E�<	$m);�A�	#15V�B,HC������
oԚ��#��xP��޷9x�'��p��7�M�O>�(�����)Q�0x�!�I!@�HbV*T�c���O�T{g(L?Q��m;�.�1g�,��)�'y��;C�}�
�Ӱ�*\�'��šT��bl^�33�N �>E��/��"�h��Q�7D`�5A2?)������	h�O��D�"�X��ƭ��҆H�\�!���J�pZb� J�!N f������V�O(���F�ݦ�!�ݶ�U�ij�W��k��?���ߟ�IiyL	K�2%3�F"j��EJ�1< �����(d����m�(��`��D֫d��8� B�Z�����T4$�c�(��;E�$:��N�
ݚ9�%���:�p�8�'��L
�e���ę�7b�u����i@��'�B��p�'V�dU�l�	�D�	�1���;�+�8&��Ѓ@e��i��ȓE���@DIƵ$�N@P��S�jҽ�'(l#=���i�S������``��A�W9��4#��DU���	ҟ���񟬗��O�����֐r�IZ�.������7v�����A����x�6<O	yBG�I>���`�:Cz�tm�_G��&��hkDzG!-<O��D��_1�P�e�-�x��~'2�'aў�Ex��l^�yA�o�j"�CU�м�y��X��P�ra�$v0�ȴh� ��[����'��7���B����d��y�,+B@�l�J��3FP4�����O�T
�(�O�$s>Q2a�D�&����"܅����I�"$r&C��C6��E�.	����D[+ ���C�  �ݡ�H�OT5s�	��V2T@@�(K	}o<���'������?Y�O���Q�o�R��@)�"[u8�)!�|"�'aaz�ʾq�pI����@ޢ�Q7m@���?!��'"jIRq矟R6dl]r^�����d�<yk�1�'cRY>Q7�ޟ�`��;<<�i�S��q��	����8����Zx�;sژ�R����?�O��ӌ4�z�RT�q�|!� Z�PNN��\���ů+�$�ߴ�h��8(£�g�T�C&ӊc�8Yb���:Ч�O��D>�'�?AJ>�!��L &29ٵ-C=�y��L�.������L��������OD5E����~0as�ƝQ^���NV�L��	Ly�Ö�h�2�'1��'-�Ɍkʌ�H���#.��=���6�lĈ�΁tWX����C����ɂW�g�hkJ���/��\�B�Cb��w�వ�]0�����i�$��U�g̓FF�X;��L�z�E�c�D��f(�O��$Ŭ	��ҟTG{bM�����3q.D !���W��(-!��s#V��#�FYxެ�d�8��I��HO�)�O�ʓ\�S@�>R� ��� $��`q�����?����?�������
5�)����RN��X!�É6n�&��A�BE�@�S-�[x��/=��H���� 
�,��!��>I�t��O�oQ�����v|��Ưov9���S�<�9�P1T>�IaA�'���	�'OpU0�Ɉ�\ޝ���^�@�m��'&� W�ݳr�����M>	�V���?�AWd*�AD�3�ԙ0�(R;Z��]�W��m�<r��.0��|�%.�6~��F@i�<�f+n�Š������i�y�<ѧŊ�O�$��W��/Y. ��u�<уhHI�$�6�N�~`�{�s�<)&������b�K���8�(l�'Ott���D�J�rL����)MV8E{�bN�u�!�Ĝ�L����i� [)�����#�!�D��FlJ�z�!�o>���c�R�!��Ә<�Z����>\�ȻҢ�Z!�D׎�	���\�]KN�{&#�!FE!� ��+ei�}I
T�U�����͓ �O?� ���>,��A�f٧c\x�k_s�<�P���JX�ka�ި�k��[s�<1e
��')�لgU�|(��Ts�<�u݂YE�R,D_��@�b�d�<�B�hi�d�rT�x@�bb(B�	�Z��蓦[l9��0���9�H��N��I�5����Su���@�^�9	"���S�? �eJ�$H.(�
�K�3��tئ"O�d[�딚h���@0���f| 0:a"O�h�9Kh��RlNEt�J�"OR��ĭ�?7\d�PG�ާ�\����'�0�'8����ID>k��Ku�NA7��1
�'�����CG��氺�9����	�'}���W'�(�AY�1��c�'o):fG�[[b�[g��,8�	�'�̈i���,�^��K�5$@d��'}�P�6O��y�w��`nV0��D��WkQ?	�i�?|!ئ`��*��񲕀>D��z&O<�<�x`�	/�6l�g8D�8Z�L��?��g��\P����4D�<���d���S-]H{��$E-D��hg%��!��!�'f����+0D��J��M�v/����M��~|�� �-�O$� �)��m�`�Y�/���nML<��"O�ѹ�@�g���5/��|F���"O�J4��a�5��F�xZDD)�"O&8sGl�6Er�ԦE,7y�j�"O�`q��N ;&�I�!�I-" �Q�"O���F���p�hhg&M�w@��RT�<bTN"�OH�y���!�`*�d�1/�YAr"O&}A'&E0$�h�+E���A����"OzXYS�G)w�l%;�S0k�.!��"O���C)�����U�+3����$"O"m�� �|�pQX��/	�X}�'^����'��=�c*��Lۇ$E�Y||ez
�'�(qLԄN�ޕ�FG��M(&	p	�'�:(�e��5��%Z��Y�E����'Wr2�C��6�5��[+9����	�'�@�B��Q^P ���ϯ2u��c	�'�z���/	q�"ݰ ���%yh�1��$O aQ?YI�O@�Ɋ�k�d�R� �2�0D�p�6�[VX@���8 �Y'G0D����%=\<�1�^�B�@ "-D�pYp "#vu1'�Тc�̀��8D�\W�b���O�
��a@��$D�Au�EU)2��jL�,� ڵ#�O�ɪb�)��r��rC�	�@Y��M�"i�ȍ��'p���d�Z�����u+Œs7:�Q	�'�f��SD����K%-$g�޵��'.�������1V%�6� 4��'ID���m�)l�|HD�?)�2�"
�'eN�:0%ņ8�zYQ��^+����,O���'��Y�����EP퀕���r�'|$�iw�W�c���� �[<ā+	�'9LA䈹$
���B\���H�'v�i`g#�1f4 ��c���	�'�C)������D�P�N�6�	�1-��_R������&��\�%ʄ�<�T��B<hR�ۆ�� �d�T<���ȓ|a�l�CڍOWJ�Y҂�H�N���Ct��IA��%x+�@7D�t9��"OFq�c�=|���B��-;�|$	"Orx�g���9�����ᑭ �$�F��.c� �~�% ȄX�ЂI�}�A(�M�<��X�H� e��a����LS�+^I�<If.�Z��1�3(��=�6�(�BI�<�H[?A�{ACB@��C��^�<Y���'g*�S6�J4m�IY]�<�CF*t F���(`4ɩ��؟�[��#�S�O�݊�H���I�	#=_��k`"OPհ��ͧLfTE3�m�>d���at"O� ��:�F�M1�����_H��R�"O~�+��#|�����	l1nxÕ"O� ���Ǯn�f<��  }��"O�����GF}\���3��ܡ\����#�O�����1��5o\�H4�i�-6D��25��$�9�p��'f��u�3D���cV�;�(5�F��T����.D�Dj���/Q�ը�ɀ�/�i%�+D��AC29�|���(�/e��؛t
+�O%`��O���&`�t�ȫ�F�lo�i�"O,)�Q�ڳd�A��#_Z��:�"O0�"EI���(@ZE��cT0A[�"OB}zq��^���i�$��2tEQ�"O|=+4��_��3&e��#|��`"O��K��*pTRa��*6n��@�퉍l�~�� Ck6-Ƀ�ԫU�œ�	�p�<@F��u�xҕO-`S��hk�<y�DZ,p��I�� �S��p�	l�<�2���7�4)�Ϛ&.�5d��j�<�4`�0<����3FC\�
����k�<f��=c� (V"�c��-�D�埀*ĉ3�S�O_�h��T��<�`D2`��-��"O@!�Bʉ�U�����	����0"O���eG+n��UC���r�R�x6"O~���	a�d���c�`ݎ}��"O����� �����!];v�ޜ�"O$��Qj'WFUj��u`|���S��㢆7�Op�q`˾�a���B"��"O���Y�o�x}Q���4�Ty�r"O`�8S�áxꥠp�
-���+C"ON���c�%�-z�/x��T"Oʸ��˟#w+����L��@ڥ��>)1�Z?��gٳL:^�o�V�TӓaUO�<�E��Q�����6Q9����h�B�<ђ�	(պm��e]���!�L�Y�<9E���s$���2��#/�����a�<!�� �bi��o�*���Md�<�b W�s��8��R����t�'/T�;�����A��l3-T2��e�E��W�!�D
@���H�ɞ�;}����;Y�!���x
6���&��j�h�b�-H�!�$G(XfHè�-lyN�y%!˾D!���#�A�E�8�a�'!�dK�9��P�6�B�i��@	���d�:�O?�
��_a��1��4��}Â�z�<1G�^�|dICg�-���r��r�<��%_����4�H2�0l��� r�<)���܈\�l� 9���(VD�<�uDQ��h�+�=
�����f�<��W�z<���3�Yb�2QPt��cy��p>���M�H|l躢�߂/�pA��G�<���P#����񤚁U<�	I���E�<�叕q���
�N�<�H�H5[�</ʆmML9�ƻZ� D8�.�S�<�L[�.ܴs���^�D=�a��Qx��3�f����Ā�k�$��T��+=-Ll'@(D����@�~����g����$&D�@§���iBd�BJZ�k[u���8D��ˤ��6l�dT�%��$�`��0D�\K�I�������tY�X*A<D��K�� #"�0J���!-V�cm>���G��R!k���r-�<rDB7�y"B� |�D��0`< �c��y2��h�!�v��U�d��Wc���y
� ����J�o� �)3d"�ְ#W"O` ���ѓS;z�C�B�6Rt��a"O|�3RO6@�Z�W˃2lL����'z�����S!Q�>�H�N«z!l�Qw���1�ȓ3,t\K!�āw:p��r���g�JІ�#�Z�#�y��邖IЁ1#"���JӾ	s����l���H��ˀ
F@e�ȓCV���F�*ZU@��Q��\8��u��3u�0:a��A!g@3F;���'?y��r��1�C@�~FVXS%����@�ȓ}�}*�A��D#�����Q�ȓD�άG&Ӕ�\ ��!Νp��)�ȓ?�؁h��S�t��ꖪ!���ȓu�����(ÜD����-����I.r�`�ɹz��,{�jղi�2@���H�
�B䉥A��D���%0PZ1'f�RC䉿Wa�P����:^,r4A�B�	�|���ʥ� <�1�`B��^�|B��;T�X|�D�P
0iw�v����2D�h`f��8]�줱�#��PK0b1�:�fdF�tK���& ���IYC�|�Q�S�y��R��f��5�A�Swl�Qa�*�yb�
!.t퐤b�J�����P��y͕�YRqe�Z�k1�:�Py�T9&Dk����~�X�-UH�<As� 
)�(:��_�~�I �`ǟ\k�N0�S�O(���F(�Fa�"lԆZ-G"O�����=h�� �O"VI�P"O.p��k� N)��+ǯ���(�#�"O��@���>b)����;����"O�%Qch�C���'$ )�#QO!#��x�"]�C�ė�D��'�O��'���'`>E�r�O�����?m;�)�#d��ZC�
s���ɷ�oy�'��'�n�ke��`�P�@�9Yc<�4�8$["��,}�X��1�\�X�.�"c�	S?�͒�&s
��\�4�
y5\���i:���a
�ԈOh}@!�'��P9<��	rV*��x�h}ڷ�K�kl�i���	V-�2�0Ę��S\��a�1�'�Ox��'8��#�P�2� �1T�*`V�9�)O�Ag���H�#�JyBV>E��ʟp�Ȏ�\c�)B�f� E���"�!PߟhH� ָC��cg	Q�"r�M��S�O��0Mu� ��/�:B�m�'��ʝ�&���
��,	��?9sԇ�J�()�P��$7���u%n�Ĺd��On�$6?%?�'��0� �E#B$B� H)6�r%��'V�P�����T���� Y7�E�]p�'>R#�@�,0 4ez��ؒak�,S\ے=i)O��ʇk�O����O��$�<9���E!3%R�*hu�Ć>|mJ��4��]�i.�h����-���I@i���0N�-�A�N25���`����@�E�)�j�RR�#Fx�&Ae��<K�ߑ_��ur2*�?��d߾#���'�ў��Z��}��"�< <
��dP21��	�Y�mK�)~f����d.���.�HO��Opʓ��bfM7��p�"�υs�,�����?& ֨�?9���d�O��� �JP�/a�9ↁwT���!$@)[��U �غ^t��@�s�b�YV�K���1��m�k��'x(�܋�쐆./���ϓ{+�\�	
'F�� % �6a"�j4k՞O�@�Ib�'��D�v�X�~Rx�B���q��� ` D��:p��mbl�pr���\E �R�̼<IB�i�Y��I5Gҟ�+eD7�q�E�(5�M�
� ������O6�D�O�\K�b�1}���2Ə�7�(��i>M�ӄ�!Z���*⟢1��Bք*�r�K��Ӌh�hZ�@����IG�z��B������@/^L<��PV��O���9擭!��zA�A5o�q���-��C��0��K�6�R��w�׊L6�=��!�OD��'�v�U�_�����+Z��A�O���'Jv�1_���O���'��<8s)o-�1L�����'���QE��~��F-#5�R��7;�(,�я�}\\�pG��|��/�U�ħM�?�i�CZn�O/^�8�k����.D�E�\�`�'�БH���?��O�O��)� ~��6�a��� �޺h�s�"O���"[�?Հ���(s�Y����ȟT��R�Ĕ�48�EU5W��H
Ѧ@�Q��d�O�Aj��̅lm����O��$�O�L���?�+��������0�AՂUԊ��ӌ�_N��(���&R5�Ο���Q��!fuʰ��iHc��-T�*���E���T�@U�`���g�'�q����D����p4<��Of����?i��Dy��Ӕ���jP9$��8Wht��DJ4D�4"%L?AL
}S�,�e�	r�C�O:Dz�O���$RB��8�4a�0t��ڳ��:���P�p?�ז9HHi�'$^{��; ��]�<�4��<;t�"n��p$�u�d
R�<�q!A�<�v��1��%FP�7��Q�<�gBR�/�fy��Lν\�&�:���S�<�%FA�D�L�3#��� EW�'#�1mwӊ�O�KP�*D1���V�m����<����?a��{���I��YL�Q�M֜�y�O�$D6ܪJ�^Q���T%�Tȏ�$�X�* #6/Թ�b<�Тڒ;���U��e�v�1%Hz�E����M�6�ȍ�$�\��'���'��ڃ1klxS1.^t}ڨ�/Y�Y��'���'��W>�GxB$�`� �A����0�� c� ���>�_���4.�,5�8�T!+9���I �<I��3��&�'%�Od"�� ��2h쵢�.'Q�H�r@.O��=�b��P��D�R��.=�s�U�Ep��&�ܣD�'��S�H���ԧ�q% 4*@ʏA�|�hc��ΌAs�S��':�D
�(LS���
�IH�F�%f�q�'@B�'�p�J���H|� o�>;>��a@��/����Q�X�'[���B��yBo�&s���f˙ft��C�l�m�,lJO��O��Y �(}��~�� v���`�	�g6����� Xl0}�IV*���c D�^��-p���Y�(�2e�O�x�5�>ƛ>Y'�Iu�d��U�����WI�i�W��Z�xb��<E�^���[�O��tr�'q�}���N�l|IA�趟�s�,}*���(:��ɋ|Ⱥ�E�$�m��Ae��<�'� ly�m�<��'��eF�t��F���Yv�V�z`���ǯ�?yh���+k=?��y�B�~%����Ts�hÝDm��̙�?Q0m,�O$�r�P05\�8�&�	9k��B�"O��C�͙<)LP���&: ���%�i��Oj˓���Oh��Y�<���s�E�$�U��ѹ4,��m֟��	y"L�~I>��%����>X�$a�̷���RpN)�D�<!O>�~����?{@�h;SfQ=hx�� bN�<9���a��M�Rc�#�Ԑ��SI�<�f!�,�@���(�lM���H�<���QX���`N�(�i3��B�<!!�ķ+���*a�H���	��~�<	�iϮ6�����F	4��T1@�N}�<'�J� �����E�YlU���x�<	g�T����%)� �%�~�<�Ղ��29[� ϳa'�}8#�r�<��ȗ	e*���˹���xLAj�<	0@��os�p�@·5B��USh�<�3듇=�Լ�r��9��,����f��ll��i�K�3#.�B�l�c�Iģw�Π4@�#V�^�:&�āy�����+] 4���%k�m�pl87iM�
�
��F�5bΎ{��ɛE�4p,R> w|(���W�d�x[�JQ'm��s�aL=_$�y'��+�,r֍ӥ ��@q�\�-Nz��.Y��i���H��ml��9|Ze�T-�
nְe�^���x���?afă jcy�R
F�|���$���	�~��lGF0xT�$���5�YY�	�&q��	@�Q��pӋ�U�OFT$K����=��0�g���eZ��J<q�� �|��4:țv�'D��r�P�b¤t'�a/�14M�عv���O����،4���)�'@� I�#!y�x��3�h.��Ån��M�%�f���r`����Z3\���'s���P�eߤ��E�W}���Y�'��e�@�]gN8t$�>F��'V2�*���	Gdށ�#���;)h�'|���"��{Lr1��jɒ.���i
�'׺MzF(��y%���[�$O.�	�'&�@�*�G$� pM��T�4�*	�'�j5��CI�A��L�wY|�A���� �����$U�h\KDmыV��9��"OV$[��
)�����iՠi���"�"OJ$�w�@F�}"�.̯R~����"OP<�PG����TC�mIU[�a�"O4�i����`ܰG�]�<"�u��"OL�{C�Q�1/>4Xc�_`�
�y�"O�i���ܒ��GA6��y�4"O�����Jnb�8���7Q���aw"O��'15�K/,�4!�-�y���g��	Q�ϯoM��:��W��y��حms>�z���� � "�Q�'��)��� G�i�@!W�JX�y�'���{"�j��Ȍ�vX��'Sb��%���Ľ��ィ(��B�ɢ[~@qr�[!p_�4� �֯
�jC�	��V��*͆~j
Tɓ�#�dC�I	����Q�%����Ug	�/<�B�ɟD
��0*X!$�Z�,E5X��B�O�:�a�ܴ?YR��&l��B�"&m��+�V�O2��6n��a��B�I�s���#��8IL��Ї!ϴ �2C�ɺp�X��(B�v��({Z/cF1��G_*%8 ��
1֥�\s6|�ȓ6��YAƢq�F�pU��;���ȓ&kXMa�LP,*����!O¹\�݄ȓuPS��ӂiv�Y[�n�+����8�yw�7g����g�-�v����h��nW0I�ɢ�V#;G��ȓ l�c�ߨK�l	+�G�m��]�ȓ&�h��j߶��WMC'R)dȆȓ��q�o�2T�
`� X�p��ȓU�hh
V�%w���Zjh	�ȓJg�	2G
Q�Kc��0�2/� ��Iu�=H�e�1��1�Sj٬X>��},���ɜF��0�UR��VT�ȓx�*�R��S�!�d����om���dx��a`�� T���B�R
X�� _�5
Tk2�:P�"�d�ȓ*��t���TxX|��KN�*V�ȓY���w㍢	��H�d�&�n��ȓ8���0�C�(<`a���7ę��k�l����/M�g`Qz��Y��6�<�ga@�K|Tpqv��E'@��ȓf��s��
]�i��b�):"lM�ȓo�rh֣Z�X{�� C��&p4���ȓw��yg�ۅ:����WB9�n��ȓ>Zp9�6cK�0�� @)
D�ȓ	���G�
�ib����%n��ȓ(O�Ygąx���V\:Y2a��gv �����i�6YB��4̄�|b�I�1ס'α ��N%�����Y�Z�W*̈́�V0 &D�m�d�ȓ�A#4�3<8ܳb]9"�b�ȓY��	8B�U�.���`	4W�d���8������ד���(`���j}�ȓFH�aäB�o*����ł��昄��j���n���H!����NC�H��U%�m`3l	�ab��4蚣?�$��R,l-��1|�ܝ��Z:]�e�ȓ���S$� ��ȣ3d�(�=��8��
@�L9u�����Q#z� ����u��A�m�x�R+߇4�؅ȓ�H"lU�t�Y�ĉfd�a�ȓ\��`�6�S+8�l	n�'�y��S�? ���R�'R�)��	�0T�"O!�*,�|S�D�&=nF���"O��`h/�D�h5�']T�%K�"O�:��$&)pq)��,s����"O*�ʕ'�>-�.V2I[��8�"O����քY�Z�v��s���y"c׀]����3�X� E��1Sa���ybya6�O�RKtl�$D�.8�9k�'IB SW��/8��]����:80���'rDyi!
�C��u��OIbE�<`�'L����O�=0S
	�B�CU�9�	�'34�BÃ*
���aB@ 	�Ł�'��AL�=F�Y鰢\.v�,}�'0�H���9�,1eL�,l`�M��'R��G�f;����V�g$vX��'�����φ��]��.���'�	2� AvUY�(�w���'MlP��K�&!��D*�����'Ix}� �8(�8i��> ��K�'ςX�6	սc*��$��F^�̊�'���tC.>����TN�!i^fܑ�'AVEr�C��U�p��Df�P���'W,8k9�z����S0
�c�'lآd-�z�.F9JlȨ
�'�jXhaE��d(}���أDe.�	�'6L���F9Z:X1E�/<{n�Y�'�R�r�j�,S�^U���'4�-�'���[�
�r�c��#6O��'���@I,G���:/3�4��'��E᫔��-r�� ����'��4��JzD*�����Y
�'p��V�}����s�%��+�'-�|��(D_Wpqj #��q ��	�'�"!"2HU'=���y���M�IR	�'����e�]qD\�2×:��=��'���0ॊ|��ݸ�m,kJ�Eh�'A�IщɆ#�Ș�!N�\��50
�'�`ҁf̬9��h�R�E ��}p�'�i+@A͂��(�5c���'��� ����:��� :� 
�'ƨY# ^P.�5"�.�Ш
�'�LP`6Bֵy/)H�K�y���h�'jj)�WK�<��u v�M�^�X��
�'� `�!�S61��`r���;C�P3�'��=y�HE�L=���?e� ͨ
�'���B���XZ��g%����'���ٳ�F�����0Δ�k�l\k�' f���k��!^���qN)�'����5���Y�j�C#���jXiJ	�'~
qJw�S�}�0�rH@�
�2��'�D�g�D(K�"�x��\��"�'U���E���(V6Qy�c X���'�jܢ���W,0|;�Cځu3��3�'���(�&T")�Z�íR���'g��KO?%Z�}�tb��Cr��9�'�q�3�ɂ(�Nu�C��%q]tp�'s��a�F��	T@���P%U0���'0��"C1N
��p5Z6��V�<��F�6[�����t�RR�<QRoX�`Ӻ��"�Q�C��O�<��ɔwu�PӨʆ]�t��ae�M�<Y��my$���cq��0����G�<q�m��_{H-��O?'����G��|�<�%�,��r��J?H��qj%TP�<� B����p1(�i EK>{�@,�C"O� ����"V�)z���8w����"Ot�s�G_0�8D��^�Y�=�C"O����nJ6��1�����]���jC"O��1��)x���av��d�DI��"O$�8c� 	k��|q0IH(c`6���"O*��,�-��;��6>:Lb�"OĴ[6
Fo�E �,�craY�"O�\ 
W�6��Ì[�v�6���"Oj��t�M*pQ�9��M-
sp�#"O�����@%_^,�T ֎)S���"O�!�o����e+�l�q*`�cW"O�Ē�Ǖ /�1��k4�F"O�L!�/�=Sen�k )BT��"O�H��GK�K�4p�GW�y��T#"O
tB��N
=�b,��� ���쓠"Ol�&`�5[�Ջ �]+�K!"O���p$��-pF��n�_l���1"O~�凡k�����:]�eK�"O�,RD�C�R��0�q�;2�Ⱥ�"O�����X����[��"O�aV�jTb!;u�_�RZyq"ORuA�.�9�� C얆=�1"Oxy�4d���`E��Ri��"O�� ǋ�Q��|"�R�֤�d"O��%g\0��}� ���WS����"O.�
���+9��Yٓ���)h*M�"O��+�e��,p�j�[��F.]h�<�w�P%d�!�@��^���i$��b�<�aʕ�/@�i�H� ,��h_g�<��G5X�<�їHR�L�������N�<��-ݎԊ=2��ݑ\b���iK�<������*���-@��4� @O�<��vkN}�hH^D�z�R�<��Ī/��Ъ��8t�J��ZP�<au(uq�XR��Xc�<:�F�D�<Y�N�;P���J%]�l�WnLF�<���T4H,:�c4!��&<�yRE�<!VaV�|�Je��LM�rrq�"nN@�<�'�K#D�T�(cS*�@k�A	d�<��)"E�U�4���~6F(b���k�<�������%�Z�iV5�VHP`�<��ނ�4 � �<Ar�[Cm�]�<a1G��:Ԫ�Ǌ��j8��̘c�<�aZ�2�<��!#=�ji��b]�<Y�� �V�t�D'B5\0P���]Z�<!cf�*�r�hG��{�h�7��|�<I�ċ*.3���5��Aj�RD�_�<i��H�>�t0#� ����Ge�<A���?�����N�Cf���� �a�<��g������*i���K]a�<�fX�-��(�s�UI+jD�u,�^�<a7F[GM�L"Q��f�̀���QX�<�#��%? ���(��Kl����l�<aD��j�`�����LP����]m�<��	71s�EQ&�-�djck�o�<�.�*b�b�+\�C��k�<�H*m{����틜���p�h�<ᅋY+qP�s�!ؘ~��;���`�<Y�ո3���g�jE�q[��AC�<A���4"����Bޔb�r��a�{�<馋ʳ=ebg��4^��&�P{�<�S��u����JD%DX�b��*n�YŤ�*x��TcB�M?��<�����E���)"��"FC���g�<� �<Y�V4�H��aBKI��K%"O(��e�H
<,}����N�8��r"O���2��"��$ᕶ	��Y��1D�[u �4F�D�x�/M9P 3l?D�<)�-�	"� �`L7d)&|���=D�캁Mǰw��
7@�k�+0l=D�@!��O$s��A�b�C	k�P��:T�L
2K� ���:#�Я8'�=��"O���B�=��i!OO�nx��"Ot�z�ڿDa�P�G.tr��"O� 條�Uߊ��&�!5z8Ӑ"O�E+&�T��CE&Ĥr��I�S"O{��0`Ý�@�K�k�"O(��1�
��5;vZ4��"O0��7��o_>��Ǝ]82���d"Op�Zg�U$�����Zf��:6"O���U�_�<yR1��$}���"O�@���]�0�B��jx��"O��4��9/����]3"O��r@"O��bFւSvh!A��L(yL�Ě "OX��"ၹP���DN�$��09�"Ol��4L7�qJ�ʚ�n��K�"On$  �
k��d�'H�P��u"O:���,,KZ�Jr׻"�|ّ�"O�m�FÒ "��������P"O��0C�؍���c�E/Q]P���"O�噇����(�M���
M�'"O(�U!��|�'�͜w5�3�"OZmyv��nmH����>{,$�x�"O,8��;]H�ۖ�ސPXш�"O��r�� ,~�Q���^����"O�T�B�+������ǟ9��i�"O򀺖`Bn.)q��<����"Oj}p�)	�Vq�$�I��h��"O�Yx3G�%t�(0�A�L�H��"Ona�$�«���#�2tԱ��"O�ɫ0�И'{֙s"��4,���Q"O�m��T!%�d��d�,�8 ��"O�{C�@6a�歙u˖7:�F��"O�����/ӆ<1���kd���`"O��A�*�S��IZ���e����"O`��&F����;$`M�x5"Ol������hd��*�LR+��TH�"ONU�d�(\���a��L�	? �s"O����"b�Pѡ���R!���s"O��#S�ik��������[r&��t"O���6��"l�H��ը�R%��"Ob$�A��.�r��t��A��ԘA"O����IN�E�|\!�$�x�l,D�`[f,O�)%��'�:Vq�m���*D�ZQkM,�Ѝ@�"2y>QHT�7D���E�^�2��P��R�zU�&F4D�lJǅ�2,�B��0C���L����%D�4"���&k�P����M0ڀ(�#D�9tEX�H��@ p(H%fU�H�t(<D�,�`
\=P��#© q��@#7D��
�W�5�5:v�A�xp`��ǯ!D�p#4�I.i��Y�E�%�.D�D���=F����i��"E�.D��� L��?�иՆ�|h��#+D����x�<�Q�C�*�J|0�º�y�+�Dp2�ǐ'Ac�I��y�h�=V�z@ۡ!_7o����2B
%�y�̞�?`�� �DIe\��L��y
� dz�G�!]�42�m�%�^q��"O���O�c|
h��Aـ�D���"O63$�Į3��Lc`���n�u@v"Ov\��϶ތ<X���xv��"O�4��H�$F]�g&�6 (�x�"Op��MU.X�D�3Х��xoX���"O&LKs䃄?\-�q��-lm��"O� �0�V�Pr S�-�"\b���"OF���#Ft��@'Z��%�"O^���k
e�3���B��7"O��q��a�X`m!e��h�"O������`r� �d�
���ss"OA��E�C��`J碊),���9"O~Q:�ƒQJb�C���O�~��"O�j�KM <;�)��@Q�^��e��"OV�J`�����@g�T�����5"O
�*��9�h��u��u�ȉ�"Ol�a!n�`?L%8s�َI�pbD"O�(	�ֹar2\����/���*�"O��hU�4��E⡤U�?���a"O8��J��i�
���y�ܵ��"O&1"ծF>�p�$F-(�L��"O��8vNI�oHt[�ŝc`���"O(E�� �.d��:�*K,:���R"O�a��"�J����J�?�F0��"O�I��PrR8���I����"O�MX���9r��)�!�ƃl�xĒ"O��b�G��Pt<���Ĉ�z��aV"O�}X�I��7�|JU�����@"O1��j�<K��Mqqȗ`,hA��"O*m["�Sv5z�(��O9�n4h!"O�Q�"Κ< �j��{�%�&"O�YB�կN�ڑAg���j˞1µ"O&����
:����m��k�d�x�"O�T����P4%�!�ε\�Q�"O>�� ̀ݾpu�	xpt�h�"O�C� &O��@�dȽiu�}j"O��J2�\�_��4@S�N!<_�,�"O �c�l>� �r���t5�u[�"O��I@�1�l(�t-�	*5k�"O9���C�� ��!�I"���"O$A�KN+R�ڼ�$�
�jP<�5"O^��H/}ώQBR�u�d��4"O��#Aդ,9�ТU��դ8��"Ot�S��R,
��T#c��h$1�"O�A�//PҼ-����aex��B"O��%�-�|У����)����T"OL�i$�O'��)iՠ�v��Y#B"O�ͣ1��[��ҳ�	*p�C"O �0��\4I��h����2Jf�K�"OJyPT6Lw�$	�Ɵ�O��ل"OT,`CJE(}"�p�M�}[��X�"OrL!��ҏ/��Z�E`�a�a"O$�7��w����aA� R>�|�$"Op2�O�Dtp��P�z��)�"O�����+�F�  *),�P:�"O��צ�}Z|X�5��#?< ���"O�\˒�ę&{���)@u�"O)ڥ㚼-���t̜�CN�X�"O��9���:4�R�J9Xn�܀r"O��;��:��%	��"!��M�"Ol�
w/Ι�t! ��/ ��+v"O�(����D2x���W�L�P}��"OV���kP /u���v�<�����"O�  �8A�ڨtk^x� �
��$k"O�D�S�G� �c�ƚ.Mg�X��"O���A�[�tnb���W�
�"O!�
ەO��#$�.~�L\��"O���EJ��%�^�h3N�J5��"O.��9w9N�j�
"	4���c"ODT*C��(rl��#�R� ��r�"OD��B�/��8���L��Zu"O ��&��AŐ��@�ʏ[�Z<�4"O�Ic�AS�[P�
E�_�|��8Z�"O��p6N�)���aP�%~��xP"OxqꥭY�F�<� )F+_4�l�5"O�⠈N �BY(u����$"O(U�T*��=|ZT���=.�9�"O��W�4��$��c+!.�ԻP"Ojр�CL���s5��l�,X@E"O,%0�fڸ�D [
Z̨"O��˃��]|P�X��\�ޮ0�U"O��Å���Q�$İ��4"O���e�*=�5��+!9ر��"O½!ra�E%j4#P$��)4��3r"O�؈�AH�#H�1�ѺA&�A��"O<��! ��Z�.y�!Y�u�y��"O\yxSJ��U{
�����uH����"O�) �T
f��A�%J\J�"O�A�����%3�	!�mʓsd �"O�p!�I�4���#�,�'5c~=P"O�D�`��0(�ޱ��������E"O�!j���`�B� EI�<Y�L�#r"O�Ӗ��]�B�hO2u��"O�]�0�E�U	0OɞzoL]C�"O�0�D��U���"OX-Q&�����Xx�+��"O.�0��Z���U�hY�X�%"OL�a��K܄@閦�v�Ly��"O Ű�잒?��Rs�L�7;l`r�"O�l`@ Uv��c˞q@�X$"O��n�7#n���g"�Z�
�:d"O���ʅkl�Q��@�+u�=bd"Oܡ�����p*`J�~u�)3�"OPmXU΅(DLJ���,e�4�&"O�-&��;:��@�SM���"O������n�8j�!U�Q.}Z�"O�)4�l��D��Cv���"O(=�T䀙o�Y�'�]�� !�"O(3'D�,�|�1���'#V�ɡ7"O�j����Y�)#�t (4��"O�!����+D�l-��8q�"O�)�5lG�Ρ{Dĭ�����"O�X(���2)N���%D�$����"O����s@��$�:=ִ� C"O\p)��+gf �zbk��Jθ�"O�E(C �;@!���Q��!Qk��c�"O�M��!S�
(��NP,w���X�"OL��B�V��x� �V�p��1"O^���G�`���G���m�""O�K���gM(����1W,4S7"O,!�ń�|�8Y@�'Q_����"O�%3QC�?;G�\QC�.MK@��"O~�p3) �lwT|cv ɛT�ڥ�w"O@�TNZ�
��ī��[�D$J@"O� .Qm��Bu���h�8�KQ"O0��OW
�$� թC�F@�2"Ob˳O_	��A��7����"O� �Ի����l0�'A�07oʽ�V"O؈��&# t��9q��"OmI��Q�^���nE FT����؆d�������$b@=<O�l#�%o�l9vg]��d�6"OF���)h� r Sj�hHc"O�V�4g�64Y H��k�r-�C"O�����$���4H�$�jjS"O��@Be�"n
��F<,0��I4"O�E2DۘrtiyU(��5+d"p"O> ��?����2�V�}7TUJ"O�!�BS�%���@�z�1�'"O�Q�I�"�D�$dÀg"p�@"O
mS���94��;UBiEZ�"O��gF%XZ�zFl��Ld�"O�Ҡ�����J���+n�q��"O�x��$̰*4��:R
�ir���"OF�y��מNWոj��9� �a�"O��Z��N �>����̆t��\��"O��ɓ-V�<sV�J@�
��¤�d"O"����-�����M�q�̼0�"O8�*1ꌍ|r�q7L@�cȈ�1"O�a��9>҉����-��xv"O"$XPFZ48�0 ���E$���"O��P��:&�����<Z���BD"O6�p�E�lм�Kw$R�*��(��"OvI(ס�r_�J��В�:�f"O~��-] Z=�:!�[��BL�7"O�)�@��[Q��h@�"~'8�8�"O~s�Y�c%��q�\&*
��F"O~]sb@�#���d�v����2"O�x�t�9@Tx��˭9����"Ojja!���`���\"R"O�� ƀ׃u�t�#+�/��d"Or̀@�Â!ӐH�'	��=�q!2"O�B%�w�j��1AF�euD��B"Oa��^sZ �)r/@Fٹ�"O�Y��$��u@ �k��L'-.zD��"O��Z֍�5m�xaI0&(z(�t�6"O��D-� 5p"���W"Oh�) ˈ�2�!I�&#?ܒ�c�"Oh(��V�yL�*��҉sf��*"O��󫊹��|z�q���[��yB"�	 �p*�"Ϭual%�6�L5�yb���0
P��Y�m����&��7�yb���v����Lh��l+F����y2��K���)�H�2wɠ��
.�y�� �z!���]	Z��@&KN��yb�����p`�E��VF��5� :�y$����X�؋�E �Ѽ�y�Q20�xKt�ó�8��DC�yBi�85\����
�u���Xf	�yb�Q������R>k7P(㰂ݨ�y�C@��eB�6c�-i`�S�yC�lH��%�W׮����y�f�T',��'ăU�&�Y��
��yi�
��9B�]���$Ή�k�!�DL�
~=�&�I�|�)#_�R�!�:-�>��CMޯ_v�2�5C�!�D�%G1k,ӣ����U��'��Ep!Dg�2�KE�"zƀ�'�����Ŀ4�P|h��^����
�'<�u����q�e ���	.�|��'� l���0ឤ;64���'�8i�KFU�XD���)���h��� �L��=v�H�s�=���d"Ol9���)$=�E��f���H�"O���4GKs����c�� B�H��"OL�[q��?���ӡE �|��ɩ�"Of���,@�Z�����P�5ã"O@h�cJ	���X�J-g�8��7"Oֹ�%�t�:����`�r�"O�p,��)On����$~�0<�5"Op\��/a�u��Eçr�.iZ$"O�\0��M&4b�h�u%�~�|-��"Oȅ�5�tkbB�Ē}��"O��2�,��u���c���T�d��"Olh�
�`(�� �K�U�j��"OZ]h7K�
h=�pujҕ���c"O�����ԇ,Z,���+�f5�	�W"O�L`t ���D���E-*�Z�"Op*�;*�4����VfIr�"O��!�ӷa���X$�]2Hd���"O(��ԊB� 7 M9���3�]�y�'�,!c�=c$D��*ӡ�y�#�/Y��cE���7�p��S��y2�ù?�P��-�&:�r�3#)�3�y�mTA,��K� F|�{�L2�y"�C�8�E�D�W�|��|�lۛ�yң@9�<�r�B�9!q,-���@��y���5�R���JW*�rx�����y�/�!) ��ʒ\�P`p�0�y���*u�,s����BO2Ya�h��'O�i:q%�:Y�jU��+N2Te,�:�'7T��BP���<�퓄Wv�8�'�����B�΢|�E�Ҟpd!S�'�.����}�d��*L
r�p�
�'^Θz$�2��a��G���r��
�'�C��;((��J��b�2�'��,�ܲ0��9K$b�J�а�'Z�<�gDC9��Y*$�
D[40��'ᘩ2�A0U#��T��3D��ݨ�'��|�����ɨî�@��P�	�'�Z(�Q#:5hXaC��	#��X
�'�Z���F�'e�$ܣ��0����	�'9* e�I!���!�:���'����˒w�t���XG|0�'1.\B�E�hÎq�&	���'�^R���(���f÷~�fb�'�"@��h����[V!C�&I6z�'�x�B" -G�&�c
��'Hf�P]����&s�T�!�b�<�2�V<PZ��iW)B�T�UFEX�<���E�"�� #�|Z��i�W�<YU�1:[R�d��4 B��x�<�P�ޗ��wL�2>~�+��A|�<if%�(q��i�$�.��u0�{�<�A#D�b��.G*m��e���a�<���Վ@hl;��J=R�H�cPh�Z�<!G.R�F]��-�q�,T[K�J�<�Gh�F�����\���IG�G�<I$V8Z�#u��G[�`�M�D�<	aL�]�j��qF�8�lt�3A�v�<�&�E�K@kw�W���عрAs�<��.�<U���*5�,|��y��Zr�<y���}!�uʓ��1Q��ckHm�<Q'�Hp���� =�9�a�n<Y��v����7,�(9�H��,L��ȓI7P�c ƓX(M`���C�)� dm���*�����E�0!h�3%"O�A�EU�	>�=c���/41��"O���!Ê�*	Z��ŀ,�Tj�"OTț���1	�n3C��!y����"O�� �>oo���v��91&I5"O�M2R
6��@��ŀ ]	�"O4�C�JJt}{a�[�LZ�HP"Oj�¢�W'"�����Z�I�"OX0�Am�;~F�s����BŹ�"O�D	!f��Q��-����"O�Ix��S)�2E�♎�����"ODi3�+�k�D�c���!�"O\�Cd�ahA�⍚$2�R��"O ��E*R���9hEl�(0��p"O2�K֋N#q�Yp`ȊQ0�$J"O��K��q� ˆg�6(P̡d"O�RU�R�$�����GS�9�T"O����D��)ӧe	:jeS"Oza��әW�A1���5�J��A"O�(�0�`(V3u�U%�j�Jp"O��QK�i��\�%��pn5i�"Oh���9>n8�0���\j��kD"OB2�Q !�Z�Z��ƞW�Y0"Oj����L��6)h��ՓR,U��"O^���>:y�`vB�D8S"OzHZЇR/DY�v`D�z=�ua"Ox|`�O��p_!���I� >��r6"O��f�0�Ι���̸p�2lpa"O�I�̲6D �@��2��u�"OD��R�ʳA�N��%��A��=�2"Ov�
��.����љv�I�7"O��� ��|��0R�V�6�$�rb"O����h�ly��/����ɴ"O�Uې狠{����T�T��f"O�h���,��,*�n+S�,�h�"O$�9�O\�iT�a!�7�ؽ�"O\=q媚�>v|�X�Bμqp`��"O �ɲo�v����5�;kn$:�"O�bwQ�M���(�cX.~dܭP"O���2�דV{�$ ��K#gh�SA"O6�ɳHB�	S� �Ƅʃ9QUr�"O|��0��8��T��[�@�X�"O(��G�+2]��Dώxx�	`"OQ�a+H2=�P�˩t�@EA@"OTm#��:����C=f�(�X�"O�1���(14��c�YN�W"Of ��I�VL�J�aC�uB�	%"O(@ق��#��%sr *E�e��"OQ[3��8'Dp#!38TX�#"O~�%��!j~,Ђ�R�u(B�T"O����9l�d:գF-|��"O��� �&+*4�7�<���2T"O�1�5-��z���*$bJ�d�H!�R"O��{�I�"��Xp��9���Rf"OX�a#&Y.'D�jsς��(Ӡ"O���6'��J8Bea$�Z����"Ob��#��xEV���^*{�l]��"O$٩�Mں(غ����G��9��'P���X=W���6�M3.[����'"�"U�]����&�*��l��'���^�X���B� a��H�<�lM��x�;��	M�X3��i�<qED֩y�攙 !�O":��f�q�<A��T�L���ρ_�hA�c^p�<� �$�����~��$2���,a2�0�"OBU�Vٸ>SP0`OA$GY "O��gK�txT��d�w)dg"O�PTl� O%D���U�\x�"OԸh�<��%b�59bR���"OXk��Ì1 ]pA'P�p��ɧ"O���+Y;/�N��	? 2y��"O���́D�j�95�[�M`�"Ovx*q�G9Q���
�C tX��"OjIc�BU�wb`���\�kp�`��"ODV7+5p��(�.�!�&M}�<qѧ\27R�z� �R4��Q�Dx�<�"�y�
�I��E5���)UZv�<���\�\a�ኃ+.|P�U�\M�<Ɇ�k�HAk3��*��8���L�<�U�P�&�r|��2=Th�@�O�I�<I�o�0I[���cOE����sh]G�<Y`� ٬��� ��� mNo�<�gH��RsA>=������n�<iD��KE䐙# 	�{����O�a�<����h�� F��12���G\�<q��-DF�Ҕ�Շn����p�WA�<�'�9��b��ȟn�Jt��|�<y`�V_���ɶ���0}��Em�<Y5h�5]��7lLs�6�+�&J`�<��� |�����@�b, ��G�_�<����i|�A:`!�u�(y�eL@�<��h	qޠrr�T.)�̉��-MW�<�M
(dtY�
B�V�,r2H_i�<�E���  �Z�m����e�<��f\)2L"���	1Z���`�<�R�̶.��qӅaY�_$0h���T�<Q�MIq$ryCg�G#m��5�v�<2F���Y���V�����Rq�<y��GuˎH&�^�H*�<�R�<B䉚�Nt�E'T�7Z̸���һPC�I�_@d@�gՏ:\�Vd�4Z\B�/;�(ً 
G�oF]�Ąê*�|C䉭��!(%��
�vɠ��.]�C�I�g�rK�>wN
|;'�$7o8B�
8�dpMK��p�B��T�FB�I"0�����^(s�P�a�=�<B�ɾ<���䒳 �!Zn��"O��q�T�f'��6��.�@��T"O�9���'|M>$���Ys��˓"Ofp"3��$�tq)�ˋQ�$��"OzD���˸D6~��	�8૕"Oּ��΋u=��FgL"=�,ё�"O�	��Xa&*��`���4Y�`
�"O�e�u�^�F�<T�S%��8H0��"OfH����#Y0��s� *6lG"O��Ѥ)!�N��"]f1��`#"O2��(� {6.DqU��5,��"O ��Ď���HЗ�9�"O��R�b\F�fm���x���p"O��+��\LRK�j�C��\3�"O�,��4Y��h �#��~��X3"O���C�W�8�n��#D�"�`5�R"O���G��K*�hWa��#�<pB�"OJE�I�(*�(H"Nˣ�����"O��Ɂ��zYt�X���/�J`@E"O�2���Q��-C�b͑ �Q�@"O���P�,D�(qwa�O��g"O�\җ �
5���� Lt�F"O� ����MQR�jTɶ(��m��"OJ��#`_�e+`00bY�A�}�3"O�)��� �\��&��f���"O�t�k�H�00�C\�<4l�X�"O�Xڕ�m4��0D��WKVY�"O�]B��F*���8�a;|Gld�"Oz`xϊ<���0�a�� Iٸ�"O�1k ��u��b�5�>���"O.}�d#%�m�2a+ְA�p"Oȹ��h6���RQ�N����2�"O:13���k����NH�k���j�"On�h�� �4+�ٲ�!D�j!��"O�-��g�����̎�-nl��"O����U�|�hT�d��
X�� !�"O"	y4��P�����IZ�d�R�""O��i5�ԝ�8�h��Ȥ�R�S�"O��8B��t����'T����ړ"OB���m@�B��A�%U�;<���Q"O.U8aI�n��i��E��)��hB"O�Ӈ�+e$����8_ =�`"O�$!�n��aZ:��1�^.m. �)�"O�ຖ�G
%�24t��@&\=:�"O"�C���PX��a��F�/�|	"O�U��H��6l3aƳ7����$"O:��
64rdT�`,v���W"ON��S�d�0��T	C	L�J�"O<y#a�E�X�aj�>&�*��q"O�͠�Xs�%�I��@ߞP	"OR)�5C=�$�y#��*4��0"O��!�)Hs�D :��R7QI�!�"O��E�wH���g����p"OHy�FE+R�*@k�f�|���1"O��sB)��ELҘ�ӅQ�i"���"O<튒��&)`���G%.Y��,x!�$��<�#J<
�.!�t�
��!�J�V+����(�Űj�(~�!�D�D��x��� 3j�u2b�i!�D�?.0�I�3�g�T80'Vx!�$��k���y2A�'kl>�	�Ɨ!�D��@Ѽ��J� z7<X;�,[6!��,��zTOڱO)x��*��W!�$��u�60�����ZS	�%(X!�!h:��Ё�M<	���4hX��Py����nE�5	í_�}Wt�������y�"N�5��q('`@������yG�:~`��'�Q�:��a��7�yBM��Tx�*rmߥ\*��q*K��y�,ǦB�Xڗ�ɮ%ܮ���`E��y2 �	iU��ڶ�R�L}h�0�
E��yb�Z�nM|��=MS�u��Ӑ�yҪJ'Ebeq��Gu®�i�A��y����T7NM���ʲzW>IY��ۇ�yb	-:Th�[��a)�P���y"$ԈP�*�AJS�XE�xצ��y U-`�\�j�ٖ|��-)V�V�y��${�����`�"���e]��y2�����!�ĲY�D=���ɽ�yBL�lC ՘�CD�Kj�,����2š�$�<c�tx��AEw*�paEO�co!��'1rq�櫗8([֭h�D��_!�d<����.T^���e��	\!��:C�ZT��∨so�SFĂYP!�$E�y�ZԌtm���!$БV�!�DE�8O����ԫLVF\��	�9\!�� ��f	?���@2 �ic�"O���'�^�Zen��J��I��"O���W���jE�Խ6,`�"O4���dC;}o��Ӄ�x��4"Ol�A& �k'�1�T����5�t"O�h±�T�1��F��s�jAB�"OZ��t��;c�!�Ty|�`"OtuiT�ؽ8���J�GN�{��"O�|᥄T3P�(�@FMχ�@)��"O����	<��P�GmЫA�@�4"O� �ыћB9�A� ��LiH��"O��rŉ��8���L� Wؑ�"O �cSa�=c+�>���V'�9�yb�N���r��B5`p^���iI��yRA=�<��A��</�H\���:�yb�Ps�&m('��sO�\Y㠏��yJ%W;H� �S�\�J�	�۾�y"�~]N
򋜓P�}�#)���y���(gb��-�^fX<{V���y��Αl���7�J�e;����\�y�a��8�4+G�E#Z��)CR��y2�O�
��YC��'g�p+�mМ�yҊ��vB�40��z:0`x�N��y���]Вx�)��]a���S��y�ݲ@�x�Cv	)Q(��"��y�� CT���܉T�����)�y��_%T�8w�>x��2��� �y��I�%�T%�*ţg'@�g��=�y�D��U^Dc���m����&�T�y��L�A$��v�X>�y��6
����%�O�s|:��E���y�́X;.�飂�y�l����yRf��e��L�1ɖwn�8u�0�y��q|R����
�ەc[��yR��w�p�*g� "I(D;����y2��WڔE����_�Ԁ��9�y�GE63��D�V�	.-~�GM�,�y�`�0?6H�pa����8�*�y2b��6$��`c�V�-&n����Y��y�/|�N�j�k�`�i`���yB;l���O@>\7�u[a�-�ybB[i�*��^#}��qk�-B2�yR��� � `��z��c���!�y2���e���/IA��
C̗*�y����D�H�.�%��Y����y2�X�+�IxtH�a Q?�y��W�l�6=au`�0E!R	�V����l����27d0�Q.݊�ȓ:f.˷�� Y����f"m\��ȓs��H������elL�o�ȓw���`ƠT��4�I�3���ȓO4��dh _��`w�؝N�RɅȓ;q�L��O+��y�R�M�%�i��?�����8�%(u��U��x��P'F4r�Ø�N���`�J'E��y�ȓ{z~t�����41�a���9f���ȓy��� e��	~���KG�Ha�ȓ'� �q䂓�wI>	-�<�G$R�<���!�����|Y���L�<��X��ё�EK���Ї@	M�<	 eX�=��M> }�H��OD��y��X9+����&��.an�j��y��V5�4��b�,��ؘ�'A,�y�b�S�� ��<�،h�D<�y
� ����N6���@Ǔ�-�H��#"O҄(���#E!F)J� �+)��u[�"OF�I�,�)B�@��S�^s���"Oj�q/�:T���׋� ;��t�"O0������S�1��4���K�<٠(�dO���� 'z�N���*�K�<Y`��?/ĢijW�U"l��GʕI�<Y�g�3>�=� �S�V+j7n�D�<e]�=p�U@ѥ�[��	c�L�<	"H���[���Z�м�0��I�<��#(f@�{�ͮ;
�}qC�C��?)��"#�6�>E��'�(�鐊U#79�� � /� �he�R�2�X�㐣�6��đ1��V��]����Ͽ���
Y���6O	o?�p�c
�㦙�rm�������G��.�z`!PJ�s��5��	N��]��A�8�D�t��49��'`6�Ҧe��k��M[a&A˴��mH�Ig�9�mf?Y���:�S���]!���!�v0�`)��(O�lZ��M{J>��'�u�ޜ{��Yj��VQ�6y��M��D��mbde�d�i�ay�
��U.)XF>r�lأH�?�.�Z��_h��u�D�ǎ���*��,	��d��3���:�&�@T����E̼P<���i1wq��K&��9'1LcVU?9��HR(�(��O��@P��$a�!P�.���m�Q��̟X&.�۟(Sٴ_"J�gy"�'��	�f����^>�u��)�T3,�(.Ol�����	��-)��è.i���݃l���ikL7�Od�oßț`k��?��O�R�K�nC�}����Ca��u�q��7��l�G�'�b����
�KmL$���JF�\�|����d��� �'}��j�,ZP�'�2F�4��2�)2'\�l�[�&�{f��?|�� ��8�^h�6��"^��OD�Y��'��D�k\q�ށ�F�ɄC�9r�nO v�7M�OPʓ�?�*OLb?= �iE����{@�^�c��{�̣������T$��KѸ$��)c�)T�>�(�R��A��#{Ӹ��G說HEmZ��M������w���#�jͣ*�*�`�kV�q��@��Ⱦ)�����O��d��4�@x��n��*��=E���q�1�OV ��F;@r
1��&u�q�����͉���x  ��}�f̲W/N�0ul��Y��K>J+jA���1�ɭh;f�$Eަ�޴�?٩�X�{ѬH(A��Z6�[�*����$��d�)���d!Ύ
Oh]�7��^��c@�6�O|�o��M�ܴ9��]����'w�*�1Dd��8ŌH��y	���ֹiF�[��S�?%��ؗ%�:u�ac�RL�X�!�ʆ}<j��ѝ
�l��%�l�d�#�S�?���:I/l �c/A�*��Iz�W!�Ht �x C_)I5�4� d�e�|-@0�1`��\c||�K� 7�q㯗h����4(ތ�	�LZ�4�?����i�|eH�ޙX��D��o<J�����'��T��E{*�N}�ab�]mZ�,�*0�.���ɶ�M��i��'=8�9���,�Ձ֍k5r��t�Ucu椛$�՟h�	�X�.)R&h���\��՟���
�u��'G��.ɂ
��E�U��('�#"G�A�L���̑�\'�x�c& ":�D{���u�����qJem�Qא�h3��u����b([�C���h���:*AY�_?�se�J�X��O�$a�e�|Kd�ӏn�u��ӟ @�aIԟD��4��gy��'���k�*�fȮh\��$gL�k���<�˓K 0[���q�Z��0"����b�`�nZd��?��S{�̦�;s   �   K   Ĵ���	��Z��tI�*ʜ�cd�<��k٥���qe�H�4��_?8<�q�i��6m�i�����X�p�Ո&�J2m#0�mZ�M�@�i�~��v쓞�䜀A�]����u����흐Pd�ZF�v�	��{r�D�'�N|m����$��AA��h���:5��M���6�ÑtI�˓}��J�pd��"b �ҔJG��Ȱ����:Q0�8~�t��b�0#���/O��8�Ba��Ɔ3�G� ������M。Bk?��O�x`�'���c-xB��	�]�
a�����(�8�kF]���	����`'扴7��8�DU
�E�K: *,��B
��$ߞ�O��#����8x���Kv	�
_w ���k��F�Gxb�w�'����'nn� ��xD����L+�4y�M����ɮ8qOf���/WWN�7䆍MA�P�t�i��Ex�I�'L�#!�Ʋ�B=ە+Ӈ��tq����'��|GxBJTd~��.'�Iᢋ"~ �h����2���OZp���F�`Ɔ8����~�T|Ps ��!���Gx��RK�'mx��	����5�<�p��]3_7�L�F9�_��D��xrL�
�5ZG�\�Z��AK��~��E�'�v�%�8��'��������f����I�LD�5X�q���OC�����	�OF���Ӻ�,�Mu�)��M!�FQ���K�θ'\��Fx��j��In�B���x	�a%��,��ɭ :�����I�,v��T��x��ˢ%�B䉹Q�t �  ����f�0 ш_����'_��z���I�O#G�S.&��&��;�d�$��.�y��'|��'b�'�2�i�?4�,�J�(	�ʹ(�M�<q�\��O@������qUkp>I�	�M�N>�r[iM(6��5%����!����?���|se ��M3�O�\��A/uX�١�/,rqѳk�Cs����'��'��I���	���I�t�M:S�9)E|�Q�T�U��������'�j6�^3)θ�d�O��D�|�7j�v�PG�*+b
4�Ip~"g�>	��?H>�O�VL�#v44:u��S��M�Gb���Q�醊S���|:���O�5�H>Q#��{�|���"{*$[�._&�?����?���?�|2.O2d�Ӆf< �xW!�4p���+Z�!h�1`҃�<��i��O���'�2�WV���@$-�}td]�qگ`�P   �	  y    �  1&  �-  4  W:  �@  �F  9M  �S  �Y  `  ]f  �l  �r  &y  1�   `� u�	����Zv)C�'ll\�0"Ez+⟈m�f�`�	.[	��D��v�P�o����#e��5r)���(�>^��9���:U�$�S�fa�|�;,t�����F�&����a�d�h���& �P��ڶ$�J b$��+ym��:E�ұgl8�HޜҜ[`��운ៜ�dG�	Q$�S��
=_������R����k�`��T�	��f@��煟QC�- �45�@����?����?	�.�����bB�cL�;#�&{be����?���'{^�:F�'��'��0�Cܦg�~��T�F3�<h3��'�:��A\����,�r|��ϲ��'1�韶Ђ@��#� p����w�ͨ��)�O��ɹ/*�-�Wa�{~�b��97��꓎O��	�l�=���?�[�4nd I�h�Ĺ�A�O����O����Ov��O8�Ŀ|��wg~�1��2;�q���NC2��w�fMq�4�o�9�M+��z�V*lӄ�o���M[��eO�Aq%aʌô=�e�Ѝ^;�J�Od�F��/-",�Tio�[/9Vnc���	�lr��	�47���j��(o��?��S.#�z�2!a�RU^$K7	Y'F�0�!�M��!ݴ}�%�m�r��<�� T1p������'��s�Ȟ,"�#d��80
����'	"�'c*��ճL͊�o/�<�XbP�'�2�'\1�ZՁ0���81���2¢v�5�uQ�DE{���Z�V��cA/6 8�R��hC�D!��?����˛�?�#�؇R�0h�T�Dlq �O�˓�?������ę3:vrb��+-��3��i��Yb�B����d/YlD����'!�ݩGfK/F�԰"�&�-1�B�>Y�x���[�*GN�ԏR��0<����0�ɇ��Έ^V�I�ŵfе� G8��'M"��	f���@�/Q��U0$*I 6��#�%�O�}o�.�P�
�c��%z��O�AJ��ٴ��'ߞ�f��1�ՠ� ��j3"�0_A`e�t�<D���BKI [*�ȡJC�6���+?D��(�J�k�^�Z�HO?:Ī�i1D�+���v��HQڵE���K�#.D�dysgD)o�Y��ْ���-D�8uČZf$�H� D��-9���O�1S��)�'!��  �o�!j!I �d�qC
�'��q�� 4XU���E*J�S�8I2
�'� �`�)��9}��ꃰG�@e		�'^��B'׳�<Mp�j�
Ba����'�,a�1�Č6�0!� �'�BY��'���#�F���ʧ@��8 )O��s��'_hA�t�Уj^M��kϥgq��(�'Sr�h�Äm%0��\����'4�0���L� ��C�ՓL����'��1)�C��Ix\X�xv,]9�'��@��G��ł�������ϓ��H� �i�I<� ����Y�k�� �l�(s`��$�<���?�'|̠�P)������<6��f�BX�!ǝ�@Ԣ�J�ꄬ�ax2&W)� ��#)cI��'�*a���W$`�٘3��I>��ZÓa�"��I�d��4�?�+ɖ_%�0 ���g,�\�p�^0����O�㟢|��
*I�|��E�Ĵ; £=!��d����#7%D7�25�H�"Q�D�d$ŷ�M�J>A�	K�Xy���O�j�3�L�ҥ�eh	XM��80"O� #%���f���b�ƍ�s.�-�'"O����DQ,n~��f��S��4��"O��C��eq�݂�R�5�\\#�"O����	�̑�`-B�Xs�ȋ�"O x[�@� x�����>}~�	�c��O��R���2�$�O~��<I@J�0
�0)���b��@ڲ����:��i
�6���^��%�|"��DT.L�d!@"M�s��X�*@&2k5��Ȍ2C8�d���C�`���s���Z�'Y����+�>��cCB3Mf8��i��ʓ����{�矬�	��)L�^�����H��L���yx����cY�7'H�C� [�HT���+Q���Ŧ���4���|��'��d�w�`�HR�S��B�j��J��t��O�$�O���<�|��#ެ6�D���	�]�93
2��8`�Y�O�pa3£����ybkT?{��͛@c�H�V(���2$��s�X(>R樨���||��B�H�9�HMGyR��4.�DY�b��\�@!&f�������?A��d1v�8�S@^�
Zxۖ�R�l�ꈅ�(0�M����1�^PBaM� =8�%����4�?�+O�5[d������O$^��t�,��8RCg+衹	�0h�1Ex
� �;A�Ғ:�����M�B#��!��'�Hdx����8�֭s@�"5a>LY�o=3�ax���?�ԑ|bl y�\j!�D?�
� t��$�yB/�P_�=rrQ@�(RI����?��'ƺ�sp�9c�p�a��%ՠ4J>!�
�ԛ6�|�V>M���l�Ť�Q/ЬA���0���������#��쁃�,�^T��S�O��B��Ҡ`�*1"ScS9 �Q�O����@K�2k��X�J�n�ޢ}2F�����l��E�y��� �_m~bC��?����h�l��>`*֜�2��+KĘ@�G|��B�7/������8Oϊ���QG���?���Sp�|��׌�CTh�G����mZ͟D�'�P@��O2�'J_�����­}�j�je�օ��x"��X5�X�Ti[�<�Rk�"v�|�<�')��5�@� �=x�50�,Jl�<H�%��<A���@�|\�|�<qW�G a�XeX�/��Q[^� fɵ�M���?�Jˋ�?��'��$�O����O0��V \_Z����G�F�Z2H+D��j�D�H�Ƞ`�;?��L�'�<ن�		�M�����̃it����ɱl���� ��\�X�C��O����O ���<�|jb�FF��a�R�?��h��+S�lD��YQ�)�l�Р(ì��yRB���Yb�Ouc�Q��ʄ�R^�U�� ��y$�W�8��y�f��T���ޏ|e�r!�D�(,����?q���!��0T�O���L!â
�i�ڵ��u���{ՆP7dH���!���%�0�ڴ�?I+O0i��W�S�
���0	H�\1	��2&�$�<���?���|d��{QƉ2f*���j�����_g�nIC3F՘K�.5{���0<�FԁƆ�v�P-�<p �����bA[�rd����kĽ8�n-��I�
�`���O&�8M�<�$EQ�+�b����
���'����O��x�hQ5c.���M�O�F<��*)�Ol��I)+:r� ��� �g%A�p@���<	��)��O����'80�����R�6i�q-҆f�&�+6�'��Y%���i��N5F�	9g(�O>��G�� ��Q!iβsl���$.?A��S���q����m�,LA�����o�V�F<EBք� W8;�	y���D�O��}j��=�f9�WA�<@b��@ɞ$GyF�*	�' �Er�.�.y�.�;-�G)�i��$�E�O嘝k�'V�{|С��kY�c\R�qf_���'�
��'}��':"Y��y&�T�/b�]Ȅ`�|b���D쁰T����`W�?A���{�^��|�<��!4Ju��I���0HP�tMUZ;Ԫ��R�?�q�~���|�<Y����T�Q`a�Y
p�a��ʟ��'�2���?	��D {`�I���F�aX2E��:(@B��!;� �C�#V;�Z K�P�$�.�'���'��Dg��)�d��!l,ƃ'D� �B�Of���O���<�|:��ٖ�Q��#�C�P��AX2n+8(���|Y�i8g-Y�
{�ymH?���(+����C�]V=&��EB��+ܝd�@L
ϓ+2Y��� �Ȍ#��Z#�}
�K������u�'��$�5�	]�@ �Õ�m� �+9D�@�1��<Kq�+�;��B�7��g}r�D�~���7
H�Ѧ��8�X�	f����!���. ��ਃ�4Qr�1`�4�!�14����1�#E����D)0!�D[�.�9�c���:Y�e��,!�$�� X�mȡo�HӠ�H!�A�h�dP��܀b���˒	Tq ў����%�|T��w.�}\�M���Dz� D�並�̀!�Di��^7�(Q*�?D���`		�"�S�D�+~�c�B;D��7c�"/5ِŘ;,�h��U9D���w�432��J�<Dy�,9D��wE��4�*�yg��5C�����O��$�)�'z���2���}դ�ʗ΀^�b�R	�'Q\]�T�C;܁�g�	��2	�'1`��#A�0�d�pb%zzb�x�'�<ѣ��A�-���2%�X�w�X܃�'yH�PA�Y��(kT�Si㖕��':,� �Ξ/(}�=s��\�
5I+O^	j �'�rU���D�
ԙp�K�V�I
��� �l9RO�**䠡��o��*w\l�0"OH�`_,��:�q�\d��"O��u- 1؀`r�(E��1Y$"O@�����DW�I �.O�^f��F�'��D8�'Z��4%�"W�4�H�:Z��z�'��z�oG8A^���n �X�"�'J�H �
�0���!L#�,Xi�'�r���)��-j��)(N��0�'o0����R�Uޔ���+��.�C�'���J� ѧ w�d����v���ZQ?%rb�7!��p�c�(7�bl(�(7D���2C9d�E��� �LB��4D�|���֘yF���!I���(��@3D�,Q�GC�8+��\5,F,��n0D�����q�z�#3O7>D2�I-D���3C��~V\͚W-�6r�&|Q�J�Oڵ��)�'	��*P�	�g̼���G�m~��	�'��'�+���#e&�Y��'���x�(.@2��R�&*=�Y��'�<����!�@=!b	XxV�8�'��}���tt��#�XAR�I��'iz�f�K�JK 壠�\�4P��)O���c�'>�y@%�*&4[p�&c��'���!Q��kޢ�"3��5z�`��'LZ�J�뒭i���qB��<W��%��'���aE@��Hبec�bZ�N`H��'��A5�ݦ�N�h ΖB���c�=kXM��T�l�FK� �xē�"�De�x��vANy�Qcׇ�(��D�dy�܆�ERTqS�\�(��;P�Җe(�ȓC��y��V:;g�EKr���<Q���0g��+% <M1�Jq���|��l�ȓ���"Ȣmg��ZP$e�^F{�ǘ�����j�J޴~�j���?�q�"O���§��%t�`�Gy>| "OQ �+O�2�t�%(��g�Qx@"OT��F�ѡkJU锄�:�LY�"O��3�ŕ?<仗�AM��Y[�"O� ��<Mr�,�,B{2�C6�'.v�Z���S4%���Ao���8���� g.i�ȓy��T��8�(�"��ɰ�*(��yuTE	��ڙoN���`B7>� �ȓ3����0ʁ6'��H��5 Pl�ȓD�ҹ�cK�Kt��fЭ*#2Ԅ�%_.�Zɟ0:�t
�%�)"V&`�'�>C�(Il)��$�p�n\jV V.}�⥆���qx���}��'C�+g㴅��s��Ñ��8܊���l�'r��	��7Cv ���:�z�Ph˯L|���ȓ|g�Y�S��?HLѷ!,O����ɓ0R��	7�ʰ��۹P�x�PDGU&%'�B�I1UJ�� ��^D@�P�V�C�I%�|����>4p��[��, � C�i�� ��b�b� ��#I:V�B��W*��6C�b�$��L47�C�	�v5h�dL8}�)��	4���=Q�@�r�O~ep�OHgZ�@�������	�'+J,�d�K?=9$���#.]�~���'-\��A�W�C�&�g����'��m���ȕXڨ��č�l����'5�I�s�[��%8��9c�VD��'܀Ի�+�/p*��`1M"`�h��DD� Ex����l�L�H��۩0�2 ��0�C��*bB���Eԯ��5�v�U���C�)� XT+���&q.0��䘂B�Ɲ��"OHᨐ?�6Tr��̶�ƌA7"ODi!S �(�$!cabGpuxJ"O����]�$4,�3�vwDIqZ�,K��0�O\)#sB]!x����AC�jA �"O�Ma�f?��<�ċ�<��<y5"OB��� F��q�t-k �W"O`TL�(��� b|V���"O\ J�)�]�T���&8Tr����'��Qx�'�"iP$��%W�	0ē��z�S�'��q6��V+�]���<i��Q"�'Őy���̼T�t=�*��Pb",��'Č�1����ּj�L9��'*Jt�SF�p�q:��"G�9��'�lq0x���QW(��Ap*�����_�Q?�E&�IR���f��t�d+D�8M��W̶���e�W��L%D�(!��D[����E!
#�p Qg�!D��ׁQA�i�E�SѠĉ7� D���îA:Zz.��V�1Ȃ<Y��:D��{3�
��~@qAAl�H�	���OV����)�'*��� ��#q�z����>�
�'��<�E��L��h'`�ؼ��
�'&�l�o�5`�С��ܯ��$
�'w$XJ3�O�
�5�U�B�'\��#�'v�𱄁�>i�VtB�T1���B
�'k"�s�JV�u�S�D��ya)O���#�'�$IHaȋ&vR�a`4�B�?Xܽa�'J^u�RfN%�v���m (b7��
�'$��3`�$�
q�BB΄cT!Q
�'zVL��OCp�b�ֻV�m�	�'�-JU��0h6Xi�Q�O�G9���	�8�FD�z��͂� ��L�Lݟᜑ��~������\&3�.YX�$0�Ԙ�ȓ�6�����,`���́:k �Q��Nu��Q�N��	�D/�6	�L)�ȓt�V����u�N͋� ʆ9��I��U 8A��VOb���Η�ZM��F{�J����ݒ�"� 	����C����:+�"O��
Am�8��
F=,���J�"O�DZ1�M4!6
����_l{r4�"OȨ�qD&Gt Q��S��	��"O
�Zƅ]P/:�1��S�"�r"O��&��EYF$�#��>w��%�6�'�������[b��sʞ�/%���')ҩ7�U���~\�`!��i0 t�`��WL�������Ԏ�+9�f%�2͋=TP���ȓ7pp[���=ڶ<� OE��V��ȓN� �c"�4-�$��	W6��)���<�S��_8*��9KP�2#���'V�	�J���i0�����3�11I.��ȓ�؀y��18��9`'ߩ,꜇�Hnt�)��+�,�����$puFx�ȓFW��A��B!Z ���bMM'i���ȓR�8��$�UZ#���B,D�,����;�t�I�q�p�0�ĵt���#��yB䉻:n,��g/�DkpmS`�Q�&/�C��>s40�9���b��*4�C�	 #��BE\jk��z`��xzC�E��Ӊ�E�P����F�[�B��#]�l�"��P2$& t3�mF�"�=���K�O{pB��,�(��"�\�H�'
�	��f�u�)!e�K�^`��'b���I��-#�x)<��+��� r4Xe�RJj������*\Dp�&"O^L��iȻ|X�q��[���E"O�Թ�BC�,������%m���Z�'�ʩ2���S�U�P����%2���U5�,�����q����5���m�$���t�j"	R u �ы��Pm����V�d���O/_��y�bK�i��B�3(����Տ̍��h�'�o:�B�=7P��Ȑ�#a��!����ʓCqz���
�,l����)v�p� �C�c�B�^��%#�66���N11XB�I����T�`��TQ&_�SZ�B�Ʌ2�~��X?h)�i�p ]5H�B��8zpm␀��p��	3"�~���ތ]r�D�<Xv��Q�B�H��uB��':!��]�S�\Q��ҹGf���o�3 !��Ƭb�@���Z�,
����E!��^9gc(P��!Y�c��u�!�DQ�?U�(2Lp	F��,!��ΌP�:8�1AX-}*�z��X
"�ў�I��+�'o�����*�!y�	ǥ3P1��^a�\-��d��%�yHLRӮ�`�<�'�*o����g�y$
��C��B�<��H-��� IS��E�<���ыFO`�4�V	2��%d�D�<���TD�c ��U�\X�l�ǟ4��.�S�O�V��k��0��,�d�Úa'Ԕ�7"On��ud��l_t!���Q�˲"Of�� (���)cmM�-����T"Oj�@�=;z����S�`�f9qV"O����&؛s�N#�܊OU�d���E�饆X�uyh���O��'	�'�8�';��˟���D�Y*.="Li4�?���3l;D��sJM�Z�41RС��;ąHP�9D�ʄ��	 �]`f�V�{���S+3D��x�o(tX��t���Kw�yP��0D����,�*�0Sr�
�T�v��2m)D��	e��"&� p(
�T3V�i��"�	�Nr�"<��~,�b�Ƿft�`Rr�B�M��L��"O�Ҁ��70Bq8�H�N[�e�5"O�P��j^$	��HCҢ0Ue�'"OL����تS�1'ӆ,���"O�Z�ő�V�xd#Ւ<]�"O�̀��W�Y�L��֠�u��
����OL�}����}��?� v�؝8j���ȓ0����fސ$ �$Q%MŅȓ'�RT��n�r�8���}"�p��(�	����;	yF��j�V�����@N�jcƑs�r�j�m��L4HՄȓ�܀��˅'����؄-���ɷ7�N��d��MH ��@	=�z�4��!n !�d	 g���BL[;���*��B!��4�X�����YC��0|�!�D�
����3i�%L���BE3I�!�dC(o�	4�X�LƑRC�@2,��{2�Ö��ɣj�|� A�]3�$
3�!X�FC�	�|�� �	]=R���!�Y�]�C�	�V�&`JE���0ɀ����3��B�	�%x�J� �*)�l��G��~�vB��A���pmm��Q0sB^h�fB䉸R���83ɗ$)|m����P���Ĉ�e �S�)I�>7*�!3�����p�S���!��D�І#��-�,p��+<!�#��)�e��T�f�{V���Py
� ȱ��Jyz�h1T�Y6`j~��5"O���!��-R����q��0%�ʩ��"Op�9GÆ8Ҍ=E�@=c��W�H%�O4�}�ke���A%�e-h��Wi��ȓ5	�1�ʀ+]�D#��=|v��v�b��#`�3b�:����4�~B�	�H�`AEQm{ܼ�wES/��B��8?6��q�<YD��'C�B�o�X�I�
�T�R<�a��;��dJ$;W�~�خ-�"M 2@�9^G�-�ЯL�ybN��DX�
2�$I����_��y��5�ĹHP��-f~U�b�,�y"�R��Y� �d�!!�)��{�'��e��B�k���P'�5Y�`��'��Tzg�@�Έ
���>3R(B�'�P�C&��U y�F/:���(�'<"xS�F9�Zu��%�V�-+�',� \��fq�N�JaT�p�'Q��+����P5�ըF2CP|i�'���C��ܬC�����^2�@�+O���O�O�6��A�4��N��bU���v+�B�	���� q��9b�(@4�S7_�lnh�ɭi1�rm��UoxT���O�-R���)㖟� �'�¥�L���<Q�kÃ5����T�L)v]z�Br픇{i�@��O���O�tz��>�6���ʖ!�5zU���#c�t�f�J�ծ��OΠ���h��>8���2v��0U82%b�-�����>aT�>���Z�Y�4�T�P�jiD�ۢ>�t�1��?)��Vy�����?����#Mf@ ���d}`}�c(�� �t�;}2g-}Ҭڷ���MsG�?I�*�k��=T٨��c��my�����	9�ȟ�){Q�)b�6mz�NF9M�@�I?�iT�T>�I;�6�����TG��{2�"׈Q�>]"�̟�����Zg��$<%�>����qEE��*X�p�^őS��OڅH�'�~���O�s���3����u�Ш ��6̄�b�F��O������pYU��3;,��eo�t�B9�ȓ[������.m����?|S�o�x�����<)��?)DՇiJ�EJ@AՎ!���E#ݛf�'rT�|讟
�O�iQ��Z�o&�e�w%/*8���M<�*O��O��:�"S�ԩm����?D�dI'"Op���	R�G��5�FJш!�2"O��t�S���Zn��/�<q�"O�`B�J;,k(yc'�8�,+"ON�ꑨmVe�U�!h���˵"O&͂Ƣ�|��	T�՜4=�"O�+�.J�
�8�p��x�̈e"O��wLΥ`&)��*����0"O�:E���C�F<�g׍g�v+D"O�4SԆ�:Y/�Ty���.D�@h'"O���0n\	m&�\��ًw 0��@"O�I���@�<�����<<(<E���f���y,ġ�RA�c�5pl���ߛ9�j�3��ѣvȄq��ͣz_�|K$�1�0mʷ OIN�l
7cŬr&���3�ܹB$0'�½F'~����+1����+Μf8|���h��Am���ʜ�FB,�@���̀3�4�BW\�(+���r�I�X��}YW�8�йZ#�>+�C�I7\��*��<6�!עI0�hC�	�SEb�����	%����(qGBC�	�2�� t��l<��˂B�&Y�C�	%I��%@��8����ᎂd��B䉒 ����k˲G����,X�C�B�
|A4��t��uC�Q��B�	� ��:��G��+�fڀr)�B�6B>���c���e�&�!]�dB䉊l@A)"Ę�A�GX�#�B��{����c���dh�	��B�I5h|B@�眤5�n�+�枣0%@C�In�LA�� �j�G[�)m�C�)� XMh��R�>`��"' <�H�"O2���#�
9ȑ�2*̍4j�K�"O pz��L�
�h$���\mi�E"O��y�(@�l�8x���;�ظ�"O�pf$^'4���H�iЃZC�qC"Ou�4�B�n�����;4:��I�"O��M	'���4K'��P�"O����Փ%BXIC�J�(t�YX4"Oћ�L��/b:���eZ�X(��"O�d0s�Ԭ��cMz��\�t"O���w:Y�5��H�~0��'=����E��Z���Ev�a��'r�ȋ��S}�<�a*ݘ?��43�'�\�X�)��,3¤��s59�'�8�C@R�>���`�12� !�'��ؐ��]��IJѥ�:/��P�'C �z# ����A��,! M
�':|�cA�Ōi��3�iHq�:���'|�0Y�^*sIʱ�ũ�b��A
�'e-(�c���
�g������	�'Ӹ�Z��N�Cv�)4e�)>�X���'!.��V)� L؂鈤*���'��T��+º7�0Qq�f�U��Y
�'0��!4Η�y%F�����ܼP
�'b��Ι�L��KgS8%O� ��'����OZ����x6k$�*�:�'n�yb�O+7�R��r�x�'�ʸ㓨��]�\%Y��^_ȉ��'�"(��_
��ɺ�Z�98D��'&<@�C.�1�v͊��)���c�'x*��׏��P��Z$M۟C��p�'C�Ӷ�·8�L�V曦A/D1�'w�,B��O�0T�QGW�4�ʨ��'S|lZ�L�Y"-�p+L�/P�d��'��$n���H�iQ)~�p�'j(r�ɧG2-���w%zE��'nPa�N�ؑ;4C�kj����'��܊���|���;kb��0�'�r=����t�5��2^�,P+�'�J�aw	7WV"���+�=R|6��'B����� =�8m�R���U~�{�']6��g!^V�!�"f�M�"|��'�(d��Jőn��uF�!D'���'M��'�R�D^^��tK�=j���'5Mq�� *q|b��4��$-���'j��0�%�
���蒹*fx�
�']$L���X�Z ;�
V
1���
�'��� ��v�TbҊ9(��hK�'ǚH�C�_!r� �!a쑀0dX�'M�x[bՅ`D��( �_�l�H�
�'Ax!Y�L��>��-�T�tb���'�F���B�:�EpÌ�)i�H
�'�`���M�T>MKc�"7��a��'[��%����dpRh8!�5q�'�^0k���U�`+"P�f���'�� qao��|���u�פ^}�	��'��c�Mˬ[ ��i��\�����'H�9��'�/J��P�4aZ2SƮ��
�'tJ� bUG�����%J�R��
�'�j�iRǛ�E�ܔ;�cU�F��Qh
�'al]xU ȉ9��C"/ڡDq��
�'���#��ٚcŞ-!��O�E�����'�.)ġ�7��P��'U�z8(�'=
4�@��*y�,�O�4Me���� �I�
��tK �*� ɅpZ|��"O���B��g��M)g [��P�P"OF,;c�D�!Q"Q�v���j'"OЕ f���yπZ�B�W�F	T"O�t�Ӈ�xrU��'�){H��C"O -�4f E60H��)A.��"Op��4T�/��0�@��,�(A�d"O����N��Z` �ӳ"O!�W�J���g��P͙�"OFY�T�}�d\�%�%u`y�5"O����`\�#Ԥ.az���"O������:��X�%,7��mj�"O
��7G̸G>�� VO����"O:��V�����E�1�P���"Of�%	�Cn"<�W��pb���"O��e��OJ0��$LN��yv"Od���^?���P �b8�l�`"O��A3�#W�X�r�U�8��#"O�ef�M)(DQ��*		sE"O�i�$OCg��-(%��[��"O޸��S� ���O��J��4[�"OXE���,�
��@N
g*}*S"O��R�$[(L�T0�f�ڝ9F�c"OxD0§��n`�A:$��|�`"O�m K�g'P�e��2�|d�"OB���NQ�(��ǅ�Jg���4"O����f�%�l���G&bSp�T"O.��JE=�P��ʕ�\7�"O�!��A+N�$ ���*1b�"O@Q�ªQ/@=�!��h�.��+�"O�Po/X�@zV
H	��,�"OVq�)Eޜ�P@�ϊ"&�q��"O0\�D�	\JIش�\���q"Ot �b�%  ��GǞ0�F��"O�Ibc��g�X=釨�%i����"OƠqgc�(7�и�G�L�����"O���`D����A�/��(�.� �"O��1.V7��j���;f�≺&"OܩRL�|�D�X���/兖I�!��Ƨ}H����ϾX�F�K�k�5w�!��Z�C��]P��D*=�J�! ꊗX�!�=O�Q�AT�o ,��K��!򤈯I܊��娕�|z#U,t�!�M�%�(-�r��)lYy�mY�=�!��
3^��+���B���fĆ,�!�$J�w~�4�T�<*t�rb㜺w9!�� �1�Fi��g��,�!��y�@X�d�޻�̰���� ]�!�ğ�x���-�-0@ ����!��Q�%g`4���	�{����.ԗJ!���J�L!6�Wh.ġSKN	T9!�u�,3M��@ �ݓ��ް�!��W�X;�52v(��pD�9O�F�!�U1���3 �X��]���2h!��.i�b9X#I�b��ЫG�`!�$��w��t��b�Ttr �$4E!�Ē�9Wn	���@��e	��Pc!���`��3���� ��P�qO!���x�Fuа���-0�%�� �d'!�$VjJ�d�⚖#vb�� �[�!�$��	���%ͅRub����!�!��  �i�Ξ%]x��-Y�A!�d ?�bxÏ��gH�	;�F�%iC!� H"�r�'"i�\,�ĦЀp�!�� �)�W�ơt�Z� CB�'��	�5"O��p�}�z����{B"E�"Od隄%K�	gZ��P�+>0
�"OD��e���=ZE�ِ~�P�*�"O�z!�I,^y�%���ޥ|C:��"O�Pp橗&x_l,s#b�x<���S"O
��]9����7!�z:���"O4QcSȔΨ�;�	�"Ap�"O��SG�:�����S	p�͡6"O@��Ν�<*\9q��b��i3"O�d�w�N��ͻЩ���`�j�"O�u�2�W D��c$i�R0�! "OD����̬�4Ej1	Е`���6"OZ]�R)ֶBL@�U�\
zA$i9�"O�	ёѶ>�&E
��01y��"O�|	&AW;1rQ��蛪9���B"O\��͍�2)��:��"U�b9 �"Ox�`�!�	Y����j�6�J�A�"O9뤩�IP�\���[7J��1k�"Oz	j6<0Q�I�3l�	�0"O�)AI`��M��C�+����"O4m8���'��0����0x�j!"O�� �K�yH�a�(�.0P"O�|qHRrr�č��[�*tk"OZA+��phYz���(���"OP� OA�2�����iN"Zr a�"Op��S�Љm�$�����2�b"O�|�s�Yj�l���!�'ذxQ"Oi�2#�WP�x�B��t�\C�"Ol� b�̼[$d�a�Y�n�X�1�"O� ��f�Rl8�8_�|���"OP�	�1C&�0�l�u�^4{R"O�9)gl�"!���r�y�H�b�"Oԁ����4��i���K�Ql)�r"O�l������b�]`r�e0%"O���Wo�!r�Lٹ�P�yc���W"O��:g+U=\1�͓q��75�`�R"OX��3<听��T��0�q"O��K3�l��D��[�<,H�#�"O��ٴF�4n%�� �o%M����"O�H��+�6�䜈���"b����g"O<�+r�.9u����g�����"OL�P�`������˞x��%"Ou��H�)o���G*S6*y�,��"O���m�3T��+B�R	�0x�"OLe�ׅ�>}A��_�H��"O`sD��?"�q� ���V��\�&"OB�KQ��>�~d�t�K�eV�ezg"Ob��Uѻj��{�#�^Fʸ�"O�� ƭl Z�B�?B���"O4�a�-M�]*��T�3R!8���"O�T9S�=I&N|��@؂g���"OJ��Q&�<�q
èW\0��"O�ݠq�1�Y���_G���t"O�2�E�;ֆ�à��$[��"Od��g�e��B�h�'?l$���"O}��<e�P]��'Y�n �䛼e����7�%�`)b��-%�'kfy��N�;:8�Ҡ*Kmw�0��'�2�"R"��_U�������<Q+�'iА��*�N�15��&���'��a���N�&FY�e?X�Vx�'%Ri��fp�c�A�P�z��'}2�#fa��vx�0b3���B>l �'�����U�"
ȱ�c^���J��� P�H�*݌W��$�ْ/����e"O m�s�Y_uDЪ`ކ�4���"O�z��ەm�<�8�M�Z���"O��"�X#��W$7D	� "Of ;3o�6v4X'%�aQ��"OPTQw.I G]�2�$/nW�<�4"O�Ec�(x��}ң;Ul&H��"O2s��%)��d��Q�c4p8@"O� ��P�<���D�C�A�"O�ݰR�%���$� �lz��Q"O���rR���,֝+;��#�"Ob�@7���+K6�;6fz+@0�#"O�Dp����増1\'�� "O�� �iT�i�
����F�-s�"O��JC���`!>�'@#_��"O��hw�ʟ'B-+�6]t��"OЭS��B�z�y e"O+5�: ��"O>EQ&�U!R&��T��,����"O�1R���61I���Ơ�t���P"O`уQ��+���FM�U�|���"O`	��/61P����_WpU�V"O��{c�%&C�=#́?{Rdx�"O:��O����$S�%�*�Ѵ"Od������H�̟-n�B�p�"O�q�"�Zkh��bC�*X����"O�����sE2M��۬?�6��"O.�)��қO?�0��Ñ1�֐@�"ObQ@�6y6M��l_:�d�H"O�{�m�%Z	��؅�s/.�h�"O�)%�hm�����%#X� �"O�-�2h[�nb�ȥBR�a
��+a"O>��@.��z�n}3�!ФgR�
�"O�}(�M���ATq���t"O��9`�0 ^��QS�K�C��\
#"Oh=i�D
 �jH�4N�:6��t�S"Ol���bV'<�L���#G�*$�"Oz����(E�,���I+7�Fp��"OT�q��_2PNi�㬎�J��l��"O�YY2�/H���k0)��y�l�c"O��)�N�*<����J�<a��iS"O�������<�0�X�5*����"Ol��f������Ve�-Z5�"Of̃��@:01^��5%7R�� �"O��3�Şd,���g!ԝx}���"O����B�$CnH��I�!c���"Oj�Z� �1F�xų���7 I�!�"OV#Vo� ��ܹ��ŲHL�`y�"O2e�_�F��0sL_�O���u"OJ9��*%|̸�24�N�\����t"O��T%���i�S�S�1����"O>���M�D �*���GZZU"O�iHυ�q�Ѕ��L���"OشZÁ���RԎ�:��|qr"O�� ա7B4����_�
�ʴ"OD�j��G
j�=*V�q
t��)D�ةgOT}^��3��;o&�pQK7D�@z�)�=�Ff��n/F���"3D����P'8���("�0G-X`(��;D����� �i)�З�N��IP�+-D���C�{"��X�
N�06����&D��	w�[)<TM!@G?f�����j!D�tc�HD?;B8X��虽F��F!D�HS�L/B���C���q�.D�l�#�8d�l���R�{�LC�i,D�� N�{L�;@�°�Y�XAs"OT�j��R,������.�I٢"O�l�A�D-
5��2�NΒ"6��Y�"O��+�ƙ|�@=�t͋�
��?�yb�����x�,48� ̛����y�D�v��s���g�J�;��4�yB�Ƚ#8�a� L�`�ĕ���L!�$�"G"~D�ԩ��S4���«_�!��m�e;��S5��4�ӭܮd#!�deB�гP�ߋ	����U��6&�!��]��,=:�f��[�~]��mT�t!�dC=2݋�N�'�e"rbׇ|�!�����s�*07�d��Xu�!��_6:\��3Ҫ�7".�t	CDܐ5^!�DZaj�BVU#�4h�U�X�4m!�D�(>}.|[Ӡ��id�#�N?!��.+hQ+p	��
e#5��!K7!�䖛l��Y�b,Ź��I��ϗ�9�!�d�G٬�cބ9�
�ۀ)��!�$� F���B�k���`�5<�!��:)�`�P�:ZXa��9u*!�P#0z���xrX�Ju�X�,!�Dλq~�V�{�4��O�/!�J�EݞM �c���0!�oʱ�!�D)E�d�%dB�l�T8RANJ�h�!��I����;�8��7���n�!�d!%Z��e�����>Ct!�d�)�"�+�>,&�'�^%.!��U�7
	� ��t���7⎷a!�$J�`����T&��Z�f�iE��!�S.K�����gǾq�c�ʎRT!��>6�R��-;za!�E֧�!�dڑMP�	��<>�����4_!��ӍC12@j�^�J��u�'�<A!���9k,�!�R�4*�iD�"DN!���,X�Y��Y&< ��2��;�!�JF��d*����Y\#s�Ͼ�!�D�n> ��I)Mx����)�$f*!��[�P�!���m0	��!�dӈBӢ5��� /�Lв1/�K�!�d�+�l<ђ�����z%��!M
!�$ˌ�X�� L�<�"ܢ�$[:U!���U�ti3f[�<"��� Pa!�֮K�F�Ȁ��l��D�'d-N]!�$��!:vq�6(|�X�1�++#E!�$��j����Ĝeגܚ��Q��!��1v(壴��}�
�uN�C�!���qc��k䇅�**$����4�!�d4S
�<*"ۀ:b!��j]+U�!��_@R��,\��Z3T�q[!�=Od��2/UCg�Qg'Ũs�!�"qr] &#ѦNU�<xd�e!�䁗\�>Pj���0F��ݺ���]!�d��q~�j�.��-��}��/��v!�D?�8%)p� I�H�ˢ(T�s�!�D�9k���C�нW
D	�'퐁"�!�$�2L|2����;�B��V�$�!�ʃ^3�Mi7H��8鈱�_1~�!�$�
eZщ`F�B��%����3@!�\$;ڒ�Ѵ(א���P�ۍ"�!�D��gi��b�c	�4�p��1����!�ӝ~T�4��*W�D��"ؐ!!�6gp�q85"�/���G:MV!򄍧\/�탑B��X��P�D�!�� �����k}�P7�[��T�"O�%����8�:�1�	ק_�>�)�"O������%i"�̪pC/d���"Ov�J�e�.	�(�BIBL*�0"OȤ�Q��*N�"��§�_Hb�"O�ܢ��H"Tlfd�%��q�zQʒ"Ol��d�(`^�����;�"O� ����+�
 �"%X@2��"Oi��ڬ=��p�eM)7w$m�"O��	��=s0�T��ݘ]�}�"O(���D�F��)�L="YȠ�"O�b���Z2Ç'�1d�F���"O�� FƟ(1�����ߩ+��|�3"OP���G�?(�>l����\".k�"O0p�D�>b�(�K�<n,�!�"O�����
<Z@�Ʉ�/X9""O!��h��/d��aGh݃�J|��"O6��A��
�й��/�h|6H�G"O�aA�G3��q�r�Ģ]��[�"O, ;��E�|���B�
�VAڔ�6"OB�!2��,��Qf�-��R� D��9+�	"�.	�	�b�"(13.D��׫X1.��,S� �e%\�Ê+D����Ձ]��R���V*� ��-D�l��΁���-I�`�/V(���-D���B� 6p!;��'WUB<#3g9D�|)��@����� ���
��bG4D�t�䒺q�$���6Zu�`�� D���EZ�M}��3�/ˀA����S$0D�T`Bc\�/��d2n�3Rr�@׉<D���6#�D���d\S^Q�O<D�d����,�i�@L��5�ѩ:D��K�K>��e��E� @$<3�C3D��뙑W+P8�'%"�p���<D�h�G! k�<A�fV�X���d:D�:�D��H������ms��;D����'kv��0k��H��9� -D���w�S�B���f��!� 5�P�.D��!q,Z�H>ܻ7ϧh�\Y
TK,D�y`�  r�s]Jf�S5D](IH!�2�<,��@ßM��]Q��T!�<�J��郉I41����X!�:K�4U�6g���'"���!�$O�5;�@�3�.�:VΞ�z7!�Ĝ�9����ꁮ�F "��H� +!��;.j��@ օvҠHs@��5!�DU;��͖@�Z�rv�.M,!��@0j�(92��650�5�'L��N$!�DD���}�c��0, t���_!���qN8��D�+�����^�!��!zqkP,I
�<;��+?�!��[\��
é �c��dˀ�0\�!��[�)�֑�b��r���3Á9�!��S�,d��O�w|t��� d�!�d����BڄZ]�m�W͏*!�d�-R��r�˃=�T���L	�<"!�č$il6��g�G�	�����67
!�dݲ.�QS����A�F�I�0!�D�4h����B�W
dT&u��fٝ�!�$��n���'��T���\-!�$�P
|qg�Y_B�`#BqO0 cʆ�.�l�S�(�����|��U����f���hѩA�y�o�,�
ȉ���^�P���C��y�fH�L$N-� h�.&"�X��Ǎ�y
� (p��V�(Op`06?dI�"OZܘ���?yBP{e��5B3���"O�@�c���v�-*���F���"�"O��BBmªa3ʩ(��̸N	�đ�"O�p��h϶:b��1�]���`"O(Ihu�^�z�� �.@;6����"OЭ!V G�=��D0�BY�M�FL�4"O�,��[�q������3�nh�"Ov�p䪐�WF����n���8�"O�\�U��*���DT3��	B"OjM��BH=� �a2�G�_���ɱ"O�!_&O%�7�ؿK�B��7D��'W�au6�3��W(r�4I��;D���q0􄺃D:Ehҹ��6D��)�ش!�\4Z����<�d�z�	3D�\25Jɴv�xJ��:wf���)<D�ܡ�C¤�d�aŠ0�l�SE8D�X�A�L��eɕ��,�i��*D�y�Ζ2���B��"`<+��(D�<7�]&=&l"E �rM�D%$D���
çc��*���=g�V��
8D����ᕫq�2��ѣ��
�J?z�!�dI�v����M
B���3R�ܸ�!�M��AC�"I>Ա pgP�~!�B�H��p0�٭��եT,!y!�dԡXv�ث���E�p8����=!��J�,l:q�����
���j�!�M�#B����e�D�rAҀ���!��Ė��={7Ή?j�LQt�8:p!���<�̕x�'(~���!��&iP!�dZ�=���Be�H��J���@G!�ڭD����ǤB�7�H Jd+!��Z�:�r c������ƨ�+a!�F�)��Cʓ|���&� !򤒏 ��Lb7,e���"��#!�I�P]�� �X7C�B<xG�1!�!�Ν>���'>y1���Q�U�,�!��T���Eѧ%)NB��E� �!�S�-��� ӈ�_"\i���.����3*��`G�	0e��o�+Xv���gM��HD:�E�4��(Sz�ȓ84|u��>� ,"G���Tȑ�ȓ���	#��2V̱��T:
4�\����E�ю_(p�TX�d��;~+BU��Cj�q���{�fYa�8C.�Ʉ�=���оB��
�f^�y@�������o]Vl4�'���-+�x�ȓs�LE��%Hd  �NBK��0�ȓW��CQ偋lej@�<߼�ȓVN@�L���@u��F��P�ȓ^
F1
�B�4;.b݂��x�t���m30�`\!��sƮ�ug:�a�<D�0q��U�,����1�H³	9D���d�g��A�%(� l��5D�0I"�E"��5�OS6}��y{�B>D�pBM��z�(����F�*~q�)>D���a:|k��KI�F�h���;D�Hrq�J�-���1`�X$R���*:D��;�L�
f�f���G>H	!h,D���TC�0a�1,�9ٰ}��/D��uCI	;��q�c��~�p� �:D��P旙�l��lK1o���Xrg6D��*TbB�p�a/
�D.R�*Q�2D� ����0]��
$�H=s4y:�i0D��  �X �Ӡ��C6&���d�P"O���!N��UBV�ڎ}X���Q"O�CӪ�'=u>��M@+��LІ"O�x�WnΖ.A�u
����C.��"O��h��E�xwj�q��̒i�$[�"O�(�A��.�*�b̪"R��4"O�I[q`�$pw�)0��N�k8�X6"Om�V�?UH���M���JC"Oxa��@�E8w�&5Y
@15"O���h��1ƀ�ҁ��uH^Y/�!�DM �M��ʉ^X��B�9WL!�ą�i�, �t��<��-���T!1�!�dL=Jì��`
M?���c���!�$�N)��#���.E#ph	�R�!�S�@j���d�ܣq<G	U�!�ǜr���q���f�5���6p�!��P?���q��^�Ɲb`�M!�DQ7M%DԠ�\�L�6#A�!��1N� �q(��j�6U���Q&X8!�ؚ[6u���G�I����0��RK!�d� Ov�80AP�V��cv'ف:$!��O�G�VP�3�á`0��� Y�!��<͜�!��?,T�� � _�!�dܛ3��d�AW�(Ʋ�)E�h3!��A��ّ�F��X���A51!�d;WjL0�W� �E��]�c'�*e!�D0��Z��/S��(�wF¥%�!�,��bo�znt���F.Z�!���Z�pՃ�o�2ET����S!Dq!�D(M|U� 瓡G�|)��/Y!��p��'/��A�(�H�<cp(q
�'�*��$��3P24�Fi��h!ԕ��'0�v�Q��= �%	,(��4@�"O�
�C�ji\t���`�d��"O��y���<b�@�q���3�<�5"O�	#�ćr5J��㜠l|�8`"O�mr�A�
^�̘�qLP�|���%"ON�2��9|���C%Ѹ����"OЫD���6ohA���Y� p��"O^�ڔ̛#����O��a"O�+�n���U�Q�}�f8�"OD ����B5�5y�ם=����"O�|�QOZ@��Y{�j�7Ƹp��"OHL�V��
$��I��&��"OFUaU(5��|�U�9v��9�"O&1�W
'��q�6���"O�t�e T�-�Z`�+�~x#"O�YB���nRNѨ�D�<4�`@��"O`���K�l�V%�EH(,��Xp"O��)��R?
_��I��\$Y*"O��x�%��ƹ�I;h��"OR�jǨY�3�$�SC-�-\���d"OX��"F�.4�n��-
3(�Rh���'�ў,B`�O�h<X�����5���rN4D��jB. ��
x��.s�i��K4D�p@R���'pL�@�aİKx��Z�4D�D0�X�X�22#��aq��QO0D�P�DD�0E�5��fԾz�,���(D�	�-\r�8��Z
��*BE
�M!�dW>���K���[�.)@Q��-FA!򤟷�"��dM��Y�xT���I8�!��Ux�X`Cq����4�̔8�!��Ty\6Ar̀5I� �}�!�䎬���p��&��ئ�>�!�� ʕ�4�o�^=��nU�1wb��F"O�}{�A^(d���Í�it�b"O���E�}xN@	�ne:�
�"OD�d��w�h< 2kF�nX����"O��jB�Po"^��d��IC����"O
�)b�[�"�R��QbU.K2<	Q�"O0�J�I2 ���a �<*f�`"O"q����\���ؕ�
*��8�"O�8��-����;@��.o��!��"O�h��CX���� Z_�HD���
e�<���ѯuO�y��D��|�a ��F�<��I#���k�'��:�z����|�<���x����1��bQȬ(��y�<�'o�&X��Xc.ĚD�P��(�p�<1ѫ��8	0�r 埛�f�P��a�<��lS)`��i!V'��$`��H�<�d�/f�)�#@�.R}+���F�<�Q��ED�u���-0�:}CF�HY�<���7H�D�A2�yg)�k�<	�dJ�r�x�1!E@�T�H�2FW]�<	�
֖o�xQi �C�5����<�#�ּ7���Bn�fL�$�~�<�)����k��	D(1BR[}�<	�,=0;Z�P%����e���H}�<�b�]��H�ɓ�W?��aK�d�<9��@C 8������6���i�<A�F�hǾݨ�$Q4R9J�F�h�<�G��5n:6���h���ご�y"-(NH��ab�	`&����Ƣ�y�5��Y�M�VS4��〙��y2i��-�����B�@�1ևV�yҬ�/�J�0E�8b�Q�l���yJh%��2�W�*��L�0J�i��B�Ij�@;"I��M�<A�/��>B��(����0�2Q���c o_�B�>� 4z�HL#=0h}�r�S'#��B�ɛ|���A�@$�w�,b�B�]?�H򳋁�j�X����[�z �B�	/q��r�*Шz�0���c٣'|B��C�^ �%��)��E�,��B�	,.�ތ��d(~QS�@� \�LB��!*���bWI.x�B���/+0>B�	���|y�C1u�P�Sl��I[�C�I1Q ����MT�������z�|B�B�r�h`CJd2䣋�VnB�ɼʶI�`ɂA��	b�S�[�RB��0B������83R�J!���VB�	{��aHD5O#��ȅ��2G?*B�	s~H����ni���SF�1P�C�I3�ޭ� /��NI�5� ��tTB�I	d6J��A�)\-\� 2n�g�^C�	�\_�M�UF�}*B�B�,�>r�,C�ɢm�]P�����f�
8*C�	�4���FF�
-6Mr�N�=bC�	�9�((��Y!6dAr��PC� k����	�8q����Q�C'�C�	�S��u��`�5��Y��\�&2C�̾�P�Fn�UYr�Z1	/TC�I6K:)y�˶N<���,\	N&C�	R��a���H1]ɦ�K��'F��B�	�1�����i� :���y!.X�7��B�I�Y�pA@0��+lThxkvK��4��B�ɈE��T;�/Z�9M,�,�%h:rB�ɧf88�Ʈ�9g{��:Gn�>9&C�)� �`�VAP:��������A�W"O�{�+ITT�[�c
EHY�@"Oz�q��60l��&�z(�l�c"OZ�@�����m�����=(l�"Or4����������څ'��m�P"Oڔ�%��y���j���	N���R�"Od��2�-	��ȷn8g���"T"O���P�N!E���LA�r�T���"O���F��$�|H"iL%ޒ�R"O�EH���0_����W�x���"O8��⋆�����Œ�%��U"O<$i��x5�4%S}��p9�"O��hF����j�b�1y���i"OF0�r���`�в��T�e���U"O\�� �ŷ�2��j��A�٨�"O  �T�Q=@}zĩ�H��>DY�"O��1��G�3`$ߦ�dH[B"Oz��GiM*@�#��8���"O��n>�~��P@]�|� 43�"O0ĒQ�Ы� 3�M���r"Oȍ���Օu^��Ռ-܆� �"O�P��n��J"�9P�]�qk3"O~��5(��P�ZI;!*�.^��l*q"O`Xbc���D�9�	S�b�8��"O
l�&L��:���%*�EP "O������G��S�a�RB�� "O�$[Ch�9_��(b��)�L��"OF
wi��F���d�P�8�ʠ�"O)rT��{�����v��z@"O�̒R�.8:ȥAT&��z�r�"Oh�8������Ő��P��9y"OH �"*�t�F�#UB�!C��aC"OH���]�A��Q��a��P��0�"O�Ap��<=1I������2"O���7�ؐ$_(�S�b�N����4"O^��v�؟�<rq"�)w�X���"Op	jt�ς;��	*S�Af�"Ś�"O��X���?=x�a�H_�ώ���"Od=Z��0�|��gS5��)CD"O��3�ߡwҴ-���@�=���zS"OԹA EׄU�J1K�dƀ���Ò"O����h)���lB� ���"O�X�̚�;`��:t��C���5"O�ihE�HRƤ��"V��e�3"O���6싊&1V𣂍emf�"O4`c�k�����gk��ځ"OZ�bea;6����$#P$��"ON�u�םiO�9zՆ�,ML���"OP����'vbMإ��7���"O
��ac��]�H=k�D[u�B�"O��*sE~��#�c>�1S�Zc�<Y�a���x�83��	)�"�u�s�<р�Իd3��h�BIH(�xva�G�<D쒅%���� ̅:o�ːO�k�<I#
6o���C]�u:��d�<��L��@��D�ٿ?�@�3�`�<)��C�a|�ey2i]�q�`)��AZ�<I�ęs���m����p%_�<�P%Ɲ-��%'�bq�uGZ�<��k�?sF>鰥%� C]���ADR�<��E4G|�����8hk���T�<i��_���剌1���� @[�<�����&�@�^�L?Tس��*T�������0\V���o<U���	*D�� � A�~^�L�^1j���"OԽ+�ؠB � ���Ww�ŀq"O��"@ޭ$��3ģ@�wy�e[u"Ol��#�a�Ҡ��i�3[��Rt"O΍�r�]�6�H5x��_-@H��Q"OF�p�YP�Z�ʘ��YA"O��i��3Q(y�Х��U �X�"O�0c� ���h��J�����Rq"O����Pu�܀����ZyJtR�"O����j�.*@I�Ӂ((��Z"O�q;@�
�9C�]J�BN8,2��"OZ�!t�<�^!i$Ir��zf"O� ��'�MN��	j&��1ʇ"On@P�I�5��*.R8F�6�V"O� $�ўx">HT�� &�)"O"%���N�M����K�6u��"OI�½��ջ�k�/Y�܉�`"O�!/M��Xr2�̥#XN��"O�ݲ�e���X�	U�@�K\Y�"O��!㉝P�lʐ�T�7B �r"O��R&�9P<�d	rh��"OJ��2� �aM(�V���D�U��"O��;L5ȁ���1@Q��H"Ox���kƷX��eag��{3����"O�h�F��^o4��M7qNLr�"OLZ�E4X�Flh�E�hPq�@"OD�+�L�lNf-IF��K��"O��#�ބN5�TȲ���X�;�"O
! saM|��i�7��|W"O�$;W��(?�H����Z�V�hb&"O���&���M��<�t
�y�dl+S"O���ѥ��?Ğ1�ܝ���F"ObD����-W$Y��GO�H��TkR"O>�����:Qx4L��M�"����E"O�h��H�'B��<�I�/���P"Oʰ`1͈��M�h,�⸈D"O�4iF)�'��T��'M�}�ĵ��"O8�8ĉX4A	��V��*
m"�Qc"O8R2�\8}�\�!�	"|���"O.���-��2!'�@AP%3�"O�Kt�D�Fq�]H2h�V�,$��"O���ǣV�b�b} �)��It"Oڹ�b@G/�h|���8j|X�Hs"O���2��R-� q���;He��8"OyC�X
32~ع��<.V��	�"O�@��]�\����F,��I&���"ORt�B�Z�:w���U��)z4�"OpT���.t]���mO�0� ��'�p"�,��Of.�6L�Ri�K�'�V�a�A�K@P(�eד_�j��'������{���*���I
�Q��'����o��q:DH��A۰;E֘k
�'��J����peS��W!8�|���'��% ��ݷ�����ˉ7��
	�'����? �0Kci��-0��Z�'��(��J.0�J�`\pn�uX�'%I���Vs:��k��աbN�!�'_�I�
��E�X�0���'Z$�x;�'yR���ב~ʴ����G�}mN�k�'�jm)�_�S� {�j��M�P��	�'�"�I�ΰ0!��>(�#�'L����F%Pq\��Q�B�`-����'��i)�&���Q"D�X�4�p�'��*cB���8�"�1W�t���� |)�r�[5~2 ��tB�3�Ly�"OpciW+�����Qpת�{�"Ot�˵/
�/� t�&��71�Υ�0"O��㎐�M�p�{v�Ƽz�E8�"O�m�aF�-���@��F+}��u�r"O���p�X�nX���*G��ٵ"O|��AT r�,��өd��2�"Oj���8`�~	��iZ�X2#C"O��  1�h���h.Zwn4K�"O>(!��-1���!���>�D��"O~|x�l�6��$��ˉN���"O��GD9pqVp��e��R�RG"ObH ��(,Zy:�Pt�5P�"O
	3��z� �ɖ��*_Pa�"O��ijQ	V�AzsGF6�$�b�"O� �P���c0xYP �58�h{#"OVIh�o:[�f�qT����؃"OVj&Pu�^e��&D�b�^�Zp"O�5�ah�D�����
" X` "O�yu�I~�=(�MW�+zLĉ�"OVmap'�0�<�Q�]ecf�Pe"O�����\.c���
]294�CP"O�<�r�9
׾}�G�L�^Wr�9�"Oв���_����F�C�1��"Od=B��c�P�w�K+O��`��"O����#pn�AS�	��5�"OLl�Ԏ�����X|+�/��y���:fZ`�p'������5���y�șop����@ߕ62��H�����y"(
	[�H���M�6�#d��	�'"�����R�G}�H12EGH\ld�	�'�aP�ώ2|�Lq�B�ר:R$Y	�'J0��2o̒R�%� �Aփ�j�<��GS�<��H�H�[Hvܺ�'Rj�<!��S�:O2e@��DF�I�w%�c�<��㈥[�4���S�F��p(K^�<S�Ĭ���Y�J�(4}T%9k�\�<��\ �&�B%�\'!� �h��
~�<	�Ό jX�E3Ū�=')nuh�g�w�<QE�A�YjL��<OC
�W��o�<�Go�� J��Խ!��P:��Q�<�'d�rI��B�j#��U���UM�<�B�#��PK݉iή�X&��K�<���\P���ɤ���B��؂��H�<�R
4-h�8�'b��QiKN�<Y�NG��Ǫ��fJ���bEFG�<��L&�.t�Ql�Q��pP��E�<��#ܮZ&���g';7V����<��'E�k{�d�0/��I�4XZ��}�<��d �E�� �L�Rj� �a�<�B�E�`MVM9�lF�N��F��a�<�� ePP%@f�ϞV���xR`�W�<�4*Z��Ɣ���\�5���"��l�<�"��2]���'	��2ސ�+�H�C�<y�6Q�\��q�z6�����W�<yF�ʎq�jDʓ�> ��W�<��	�&-�2�{��t@n9Q��j�<�HC;Ģ�1��I�J�(1QQ�<9v��e�pRDC�9�b�
īP�<AuퟱH�R@�5���K�z���Q�<���7�&�#�͘4ǎ5���F�<)V�QJ�A*u>Ƽ$��]�<	c�F- ��
�g� ��u:S�W�<��II�)hL"��ε�Y���I�<� ��#��WR~����/(s�5W"O�{��Գ-`ô�V�E���"O���'��i��e�V&(d"O��%!��=}N̻�d� /FX��a"O>l���@9RY��15$�uB  w�ßXx�fP�v����'K��T?�{�%R�$L��BF3.�IS�ֿ��� ��?i�<��5�dN ���r�`ί~ʽ��+{>9p��
k���5���D� ͓�O/ғ]�E&��%0�`{�G�h��ᤥO�\(֩�6�� 
HF��>[��"��0ʓU�	>�M#���d�icą0�/%ް��CV37��7F�O`���'ATm0�+K0Tf�	��-
��ɨ�����f�R7��{,�!��iX�;G�]!:���(�l���4�?�����i�0�����Ox7���3Pd(����c�69AeH��e%Z�������Jj\����V�H�k|��A�t�O�kF�9?�I��0� �ɱFK	T�F�ʃl�5{E�\���Mf�TD�\c�4�C��F�D�8� �>���ߴuJR���՟X+O�4�s�Vu�sa�9\�pl��[���P��O��d0ړ��'�NhX-Y����$�=�	9���^轢2�4��O&�n'��Dto�"��#�g��g����	ğ��ԁ��;�fE�	ҟ��	��c_w�R�iTЋ&�ݔ<$�ZN��,�4�$&X��ӄ1��M��şLT��� �O>�����1��4I�b872.Ta���%jJ����ɖ-�rb�f(�SY'Db�Pz���*w,���R�p8c�h�>y�L�ܟ��	���?������r�8�/e��A�r �7Gt|��'�"�'�ʟ�O&� Tf^����!�;s����l±�McR�i�ɧ���O��	#E8��`TF�	vb�X#(
\	��
 lѽ<�ĵ�	ğ$�IꟜ�A\ȟt�	ڟ�J*�0aQ��` L�R�iS
�,z����b�H�z����o� i�d�Ij(��
�Bذc�n@�Rs�8�Q�קV�6<"D`3��   	*	A��k$H�xeb��{$��O�53Ц��S]���So�9|�&�����im`%�x��˟`�?�O{�h8e��R�Nx�G���pE��'4�"=E��_p&��k6��y4��&��9�~b~���lZIy��2(,�7��OL��~R�M?mv�rR�:LK6��RM U�)Ц�'���'�B��瓊L���I�'wN�8����|
�BٴYt�h�r�.2��b�UX�'� �(���1*7��8v�V������@�$�l������p���Q!|l��(N3c�4����On���j��)�TFݾ�8%���� ��<h�D�2�?9I>��S��?�"L΄���ҢP�8����,K�`�'��6-�o�)w�ڝh��ªP�T�dd�K> �*@�iA�DC���>���?A��x~�U����?)�4{�|���� _�������w�y�G�ϰX�V��V	+ڸ���/A���'�����ט0h[hxe�S�s@��1mP�tAt6�C�?ǔ��S�ND\�;����S�ll���s���磖�l�%p� �wS]KAcc�~���'646��ߦ���~��M�Æ	�O�H񪙽��у�m?����?���$�Ob��4�IRm�F���+�?]�L1�u�Vb�Q���޴؛V7OB7��O��%�g݁1$��lmdMPqL�/f �Y6D����=��$   �   J   Ĵ���	��Z�ZvIJ(ʜ�cd�<������qe�H�4��_?8<�q�i��6m�M�X\�W�]�Cqj`�Jʦ�Btm)�M���i��F쓄�ؒ+��I��+X�
)�G��چ/��3 �"�{b@f�'4mZ6��h��b]BzP�{����1���#�-��#�@�� ���(6�ٱJ�\�E����A�eLIY�ĸR�BXC���l��&�ğ�� )O�i�8_��	P@��V��я��s�H��,�M�'c?��L�Rɺq$���튚R��ɋjt(����Lve(SMJ-VX�Ih�@i"* �ɿL�D�E� �	B%��[�J�ℛv󤇠�O����kG<��ga�8 �$Ւ;�EFx��\�'���'�~]�0��H�`�QDR8Q���cI�<S�ɚ'�qOz�� M�'��,�GE��"�\;D�i�5Ex2%�K�'B�xx�o]�,K�HbLD�-].�D����'::�Fx�N�X~2@�����! �'���q���� �O�BL�7e�� 9S��#G8���Ό;ĀDxBlGg�'̈�ɇ�T�ҰP�;.�m@W�	�@b����IR��'&2�cJJ�r�̓��[�6 ��'�*iDx���Z��9�~$�! 2-��E.1��p0�̀��?�լ�>A����e��s�T�O���;^n�5B ��1Y�}s�4��@A�{
�}�'@��O��)�!�:b��G�>�.IµT�l���I�m��8�f�A6����5�؅Č9;fe2D��h�   �$ J](P�y�~�i�,/D��R#ř"}l����B$~it�"�.D��XvhN*,.��Á��f�F�r�!0D��"���;���s�Ɋ � I���3D�`r�� =���cv)H6V����d0D���q�O�H`��DoS� ���/D��ZU.�1@�|� �Ȣ]y�\sq.(D�h[�F��Yҵj�h�S%�'D��y�e�C��\�g�T=�=�v�!D�D���ߜW9b�j�#�8 �Yڔ	?D�ԣS͔T�J	��ϑ�r����c=D�p(���'TVl�����20�t-pө?D�\vF�FxMa��E!R�45K*?D�lcc���lqR�PB'���[�D;D��a��M�_��H��_*I��|#&�:D��z`O�}f�"̟6���ˢo7D��ʅ��YF|�����	`��5D�1��Ȕx(�ڟ�΄q�i4D��(Q�\�j���e�{�0ʅ/'D���#��`��`��Gx�q�1�#D�� �uѷgA:R�8%��lБ8��(@�"O��z���|N�!�e��24XR�"O��C�dǗd��F�Z�_b�a�"Ohp��L�PȰ� L�G�
�S$"OZ1�hE.?X����"���P�"O4��e-�8�0k�&(�N�KU"O�QIs��g��5��K�~�@��P"Oh�aЎ�{�|�˓�%,f�� "O\HJa�T���I��*A[��(B"O�9y�� /�l�|P��o���y2o��!u�;��ܨO 0�O��y�U�Fݖ���@��Ze�fS3�y2�G�{Z�eˌ.i�1�D��y�!��fp�h�3��2r�Z7���y�k!Oπ�
�E0V�\顶C��y�����i�/
#8����u�ǎ�y��;m��5K���z�����y�iR#|j���`��%z�� S�$�y���/q�0�+��,�ubҭT��y2�^��pk��"���5K^8�yb��;8px�4�O��43c׀�yB���"��G�8}�"�:"٠�y"M�"	1�1 �n��ph�G�2�yr H�H�xi���5��)����&�y�e�v
zD�� ���D���y�-2P�(јg�����A�6�y2�1N�Q+�(�v�T���'�y"��K��1��l��|�%���yr�G7��Y��H�]��C��,V��PJ3mHai��x5�N�d&�C�I&-��is�ѯ1��$����#��C��1p��ZDo\�S�X����֩3}�C�ɡ"��8aK^P�|��٢�zC�I"s�ԓ��U�ED�u����V_bC�I�8�|��`�Ǆ%z��,<`C�	�(���P�!K�T�jS�ˡ�PC�Ia���"â<j�x4g�7"x�C�Ɋ�`RD�^(`	�
թhٲC䉘*הȰ�-J3���h�'S�ke|C�ID��!��A�	c��p�,F7�@C�	�,�(l�,F���s�D�"C�6&��$L>/)fA�񇆬2�B�	�cƬ���.��3�Fd�"B䉝z���9�*�)*W���CD�%��C��+/ڼ@ҋP�q��;�FC�FnB��<#r�쉐�ز���Ia��}�TB�	'R�8pf�'~�A���g vC��/�����%.�#U�x�r�:D���bƜ"���[3��kS���7D�0AF�E8<��d"��<QڱzF-4D���'�R�M��;�`�Y�Ɓs�e.D�T���+s�R��P�65�i�f�&D�DٶA��5x��BckɷZ�d����"D��S%�yj,ݫ�
�4ْL"D� �)�}��-0�'���{� ?D���D��7�,XZeН:���3��2D�d;D���s���ƍ�8)��r��1D�<��),��{��N�Ovx"�0D�Tb�Nǰ|4�	����ewxx��/D�� �1-�QE�ަ^�(�3��;D�#熋S���;�-ЮyC� �i$D����Rvȹ�PmX�l��UF"T�D*3B�9n�2)#���;��1�&"O�)k����zG�j )�F�vkG"O� 6��Յ�,c���$գ3�=
�"O� rS�>?� ��7�2�\$��"OF����ܕ70��#�C!�%["O�����(
��9b��$VD|�a"O|�#s`@$F4TVB��r]�}�"O�<�� ��b6��cZ�D>F�P�"O��sHK	uz)q����[��0�"O�$�&mY-�>��Kͅb5�tH"O�ٓҦ�(ڂ��J�L�|%�s"O�,[AOߘXr�3	�
^���"Oj��d��;�X��Jey��"OF�z���7��8*����԰d�0"O�]9���g^�0�%_�#� �1"O��Q0"X�2%<Ј�M�=��D"O�z��NM	�܀'-JX�i�"Ol1���,�=��"4Oe��9�b���XF�PeB[�.�,�ȓ%��`6� .%c���?+��h��?9�T�K�c��`�f������ȓ �p�e؝3����`�7�%��L��Urg���Z9��*�6���k��cE��:p�������e*D��ɐ4]���tO<P=����-&D��thͬn�d�+]&+��sTG"ړ���*§ �����ԓ�=ے���_Ghh�ȓ�*��RB�;�n����;5L��Z-��Y�Ā����с��8��+I0ȹ`%}��$��86<�ȓv�\���?+����q�˄p����P�
��ƅA���!��S?!����M]0�%���Vg
8���K�y���ȓ5��9{�.ԏa��|Jc&�h���ȓȑX-@�%�d���C4{��ՇȓFPu�U+^�o��@h�-\R�!�ȓ�r`1�K��d�v�ѯڥQl��ȓ5=��@�F^�L��Pd�7h���K�� ��E�X͈��)�4o r܅�(�z�Y�4o���aB<;3xa�?��N"L�f���[\�tA�g�by�ȓF��a1!��V���[ E�T����u�f���NUij�At��$a�怇ȓO�TE���?W$�t�&C:�>�ȓ'��i׈J�R�b��x��T��۠��cʘm��$/X�,Y|��)O���d����m��
_�+�Ԁa`�ڼk)!�P�e+Bu�r-^�� �H0�>�!��M&b�bAڂ@�>X}��z�I�!/�!�D
�A1��s�eۇ�L���^-'�!��@�`�����j�;S���(����6R!�_�v͑ӅG����#xȆʓ)ciSf�^
�Ű��&lB�	D���h����vp��i��`0���0?ٗ�u��M��m�3�*�����o�<Y�Ȕ:U�&43CksJd���`�<قѤc����A>^�`I�r�<�%�H(���K�$ж���5#@m�< m5rZ6�PU�6��Dذ�q�<Y7�5o��[���K���aJo�<a��؈`ZPp�`0\��r���i�<qd�g�c�k�^}�h�o�[�<��W�sT�SB�\����	D!�Z�<��<��8���j$,=%d�Z�<��!P)DV+0�P|P�C���!��@%"p���%��	|.9eݶ!�� ���Ԋ.�<|��8gly*�"OPi��$T�[���O��~��_�����=p� �zC�N���s�f_8�"B�	AF\���Y<�(�%�-D��C�	�OO<	���՛F�F�rq�,�C�	!8e1!˓�D�I�˕�+n�B�I�.!�$bB�N�T�9w/�,e�|B�I��p5¦JY�Ax%���J:C:B��\X��#bL?t��	��=3Q�C��%H�zɒ�_$l�<xe#P	-վB�ɁUi�H@S���#V渠d,#[XB��<|�n�(��|G�hIs% 0FPB�>�΀��� ?�n��ïC`�C䉜C�����"���w�3nC�IG�	�F��R��T҅���K��B�I�E�R�V�}_DY2h4:�C��9?h�4�2�
(���H�nC��:e��i�J��&N�����R1�~B䉟,���QKF)I>�
��2�C�I	#u�kteV�K�Tu ��k�B��!G�5�r�Ĥ6�f��-��PA��� B��sd��%I.����C=_�!�N�s�&�.Y`��e�!T��O���dB1�ְr1Æ64ڴ ��V��!�d$Qbf�2��
s� �R"	˪%G!���7�j�/%(��0�&�o��q�'{�$ë�>E������Y�z�v`	�'��9X�c�*(@Iʤ��"ۮ���'�HH���J)(���S���|YxO>1�r�I>L�<	�Ǆ��zeX@%�iςB��V�D�pE���y�n���n�XB�	r-P��ب�V�U��C30B�I54�çX��2���W"�C��P9�ؒ	Ɂ7p��g�A&�C�	3v0�K����Z�8"c�Ӆ%��B��
|'fD���+~��7 ��+�B�38 ���ݺ�>��c&"��B�ɨ=��\�0��6 �2\���Ԟ
�B�I3iV�Q���8tt�
�ֺHB�I�GI6�3����"��;�DB�	�'�v��S�Ηq(�Ape�b86B�I�y�0�!�H�j��rL�wJ����h�x
䣞�M��=0�� w��败<�	X�'m�Ɉ)�����Y�Y��EI��C�	�^�&X0���^��X��aA��tC�	 ��QBg�t����b%�V��C�	<tvi�E�\�{��ؒ@e]
��C�I7�8��R�$fa���E���[�FC�&d��@u	�/uL)���8C��8����(��4�pB
�Q'C�IK��kvA��Gd�pR�����B�]u�M�� �7:-)���!�C�I>l����-�X�$\6q�C�I5E�R<9��%	�m:����c_�B�I1�8���/ƞ)-�!!�̋��B�|�|t���O��)H�	�Zl�B�ɖ<�n)�a��t�D���]��ʓ�hO>a�)��Bi�Hڄ����R�v���I�θ P�!W!��Ee�<K^���#�f4xV� +(j8�V�B�qֱ��/ ���_4]3H,cZH���t��ɑ���z�d�+d��>	�J=��h�J�[�˟�i;�*$K�fЅ�e����dվd�4�	g勗qc�E+��� "��7AP2|�.e��
�yB�z�U��G{��C�-[��I���:^�ΨU䁘q�!�Ē/��}Q��S�;��B�!O��!��ĉ!Fu�ҦO:_����dOX��!�䁀}��Ӡ/i��m�L��l�!�Z#ưH��U1T=2�3�j>?�!�dI8�`Iʡ��q'j���)DA�!���*.�Fƈ�9K&t ����u��'��O?�"f�!^��B��CK�*���E^U�<�v��PP�A�Rlހ�n��G�H�<�m�2R0��c��X�H.J��QF�A�<Y���F��Xr����}w�r����<QV�_7@`����%���i��}�<���߀G�Rа���af���z�<�R"X1kc���$�
s��9Q�+\�<G'#�^�;� Z�$ �����p�<��ObA�&S4}֬�j�<q����? �tCNƌy�@3�d����<	�W�&��d���Bz�h��[k�<���׵/D�=q�eJ�HƖ	x��D^�<e(�|��1�$�n�\��Y�<�v�X�H��Mi���	k����%�J�<��'��P����ՠ,wc\D[�a�<9��Td�����\���_�<��&
Q��a���M:�����[��8�I��،�c���xy��%��@����t��CQ^L	�u��0����ȓ_�9#L��:�@q�5ǂ��Z���<X�+@�F��PJ���ȓ#z�Y` ��s��ճCL8 �ȓN��-�ҩ�7�8 ź�G�z�<)q�X�6�*| `������)Ym�E���O����́*[Z9q��?�r�'�T��)J�=����>�0�'���HG2/���ρ5ogL����O0uy�jۖ$���hui��f�>�� �'���|\>c�擪lM�@�G^�|bOG%�6��k�P�Y��Ě@A�!"��j=�ȓb����,=Z֘����	->���ȓIz�1Z� D�Z4B�z�E�C.�u����=��苽UbH�V(�(h���ȓR� ���;+�8Hـ��gO�I�ȓ_�(�hU*�7�‐�E,!?�Gb�'w>	�f��!�EH4e��zhI�� !D� �7$�ř�EL�t�bI�* D�,y0�dD�U U��v�PQBe=4��!4oܩr�@A�g�g[Hx
��x��?!����ɢf�$9��[�n�'"Of(��UjX+��ւ$
�m{B"OԜif��E��tP�	!Q"O��7�	Vp�BbG�{�b`�"O�P+GFB(�vՃ�Il�~ ��"O��3B�T!S$}�#��l�֌�r"O>�ʧc�!��U1�
�F����"Oʉy'�:@�1� GՓr�l���"O�E0��V��r�eШ
�@qb�'w��xbOG�t:sB׳>P�����(D�x:C�2���C� ��%�,�E	%D���w����}�eӯi6J�P�=D�4S�E]s�pA 5j�>gB���E&D�����]�0�
��c�z�ڱRǥ<I��哾,P��#��	$�.��D\P~B�	�
�|�sB�^]40c#NJ�FodB�	I�,K���.9wLa �K� �C�)� ִ�QŔ�m�ĵ9A�ǡ!/�y("O�*�@�n6xKb'Q�}v|�u"O���J6O%`��.G��""O<�P@��
u� h�K���p��P�|��)Z�'GD�K�Γ��v��㬚7N��Ax�'�ґ��G4!���nY�K�J}��'nΑ��O�'ؔ����=�a�'��Y�B��ɖ�]>�3	�'�b�IĂ�l�,���2Z�E��'V��s�䍽_��Y�+Y�3�` ��'�z�*
��1j��~����'ebX�6��z߬�Bb	�~`�"Oʀ��7u����F��sϤ��P"OB��cE��jR�7�@q� "O�)�%k���F �Q��o΀�#�"O�����=
Vv��ǡT�Y��i"O��S�&L�r�B!BL���"O	�� ބ{�]�PAI�-%�!�"O6��4��F^��¡��(-��"O�iK��H>y�BJ�ϑ"$t�"O�X�잠jǆ�A�^�}{�"O4l�~a���8>ձ�oǎF!򄎍g�|:�˓I mRb 
3	;!�dD,12�Y�.E%&� X���U(5!�d%�m�K�6��5�7�̓	!�I�W�|�ݴA�R�Z��_�7R!�Q'Q�̡a��ZXP��u��/S:!��E�I,��R(�c~к��^�>�!��>\&I&�N�敱���j�!�D΄ea6y�I׾R��C��5�!�$O!L�9:0j�kM��`#[�y��y���%U~0Z���N�bp���2�B�I�A��`����SJ=QR >
3PB�I)xt�g�_X*� !�P�'�JB�ɜM��H��WUu��2�-H-/!�S�0���#����bQ-�t�!�d	�9�X����D��!�w�� fA!�d�>�Y��GH�d��IԌ	L,!�D�	x� �Ǒ)P�a����E��h�D�.r�<�w�];"�*l�pc2D��ZF�A�,:���"<�����2D���SB"���l�Ct���#�:D��(׀8g�B�p��V7F�V�
:D� q`⊩Q�zU����@%��6D�d�g�ņ1H�8�0
.249�cA"<O"<�C�֌C3~��֩�z��`#�GV�	o���O=lqaСՄ'a�@�@�]�"��	�'Ͱq*f�ʐ'b�si��]�� (�'jr ��萧~�"�C��]ݖu��'O������â�S�'�8�r�'O��z��)>��s�
�h�I�'dwm�����"�b�c�'�$)�GI_�}�� $`��bd��'�%��,���PS��8�8�'��q��+f�ЃglO=kL���O�Z �'¢�ZGG�0��4�@��uפ�r�'��bG������Lܑ`p�uc
�'����.��R�U���Z�\���'���;c�1=�8�k���YkRE
	�''ĭ�'��:p�p���1"���"O¹�� �����(�h��"O>a� (� usr11�08���1���8LO�܉�B�'q��׭O��j�"O��@D��w��Q����"�z�"O� "�S�I�mQ��	���RR�"O�����z���h��Ǚ&z��R"O�`k��ٿX��}�V-ϡʨ�0"O6l��#t�Q��m�8����"O�"��B�r���R18�����"O�-��	R6eZ�ʓ�ˆD.d�C"O��C,ܷ6,��c�ԴN>��#�"O�$k�M9Vtۦ*�\��"O��0Έ�r�;�� k��A�"O�9�tJ�g`�q�#�L����	}>��1��lt������>�Ќ��$9D�@[��ԆO!EŐ��A8?ɶF�j���ҝ!�:��չVL䁓�4D�\��Y$s����P�S'��q��%D�|ۢ���A���y��Ԍ(�r}{t�7D�� G(��2z�SӠ5'� �ӆ1D��`�b�,�FPq`D�m+DqS��0D��(�I�f���sl� %nF�3��"D���Ѧ�> 4ٺ��X3��%� �+��=�Ol(h��0��h��Q�	
��s7"O����^&�L��M�.�ة�w"O��ÃB�<I�IhUGȣB�*%��"O����!ȼ��,��.����"Of���"-yt����"Fj�_� ��ɂ`\}����}�Hy���D@��C�I�p���ؖ �B���f,�:H��C�	Z2���G+Kh�� R��A�Im�C�	#��b��=e����-�FC��&CR�"����6�@���	�d�NB�	Zh�0t��K�9�N�| RB�	�WKh4��̀��<|�%�ЁW:�B�I�b���aM �E����o����C�ɹU$~p��g�-;�}䚟"��C�ɋ5�a�b:"�5��Z�KO�C�	�H\���%U'P,HKZ�G)6B䉪AM�$�"n֥
��p��Y[�nB�	�J~�H�狚<�\z�B��fN&��'�I�@q�����M�@������z�C�	8<K4��&��(���^�W� C䉋<���%�{�B�1�NڍzOC�ɕGpL�
@�*C�\�JP�ׂ^�C�	�Js�u	t�D*
L�!3G��LݤC�	T�@�[������JʜS$�C�	J�H]sqk	�oz��v(G�Vr,C�G#.=����0 �R)��+�(c�&C�ɭr
̩�靂!e$��gC$�C�I.�`��0�82LO�Ae�B�ɛ(I:pDC?y;�M��LG.kw�B䉈w4v�Yա]�3MN�84��<��C�I�@���� �'J�6([ց�3
�xB�	3�Cԍ\'%����B�P�i�(��$+�ɜb�̸�g��F���P�͇sf���%�ɷ$2���ר_,���yKʉ�XB�Ih�0cw͑�y��u��ʮP;rC�I)5��� ̗�<H4Y����Y�HC�	�?��(�CKI�Vp�X��-aXtB�2��lV��n!� �g� �BB�I�MQ��x� Ěd�-ȡ���B�I;�t��r��*T�e@#��YBB�#Z#��� ��MMR0�VJWz7��ȓzB���A\6���IZ>��(�ȓF$��۱���h)e*������i��e d!�
mT�)��t$�y��{���y����K
��͛�Rժ��S�? lHˢD�,�� W&�}T"O�(�g��?**�ԁA��	�Z���"O�M�O��P.<a�$��@�P@��"O"��S�1t�hg.RU�q�"O&=1vHD3il���#�j��i��"O$(���E3�
0���/j�hH��"O��B#@�P�0�����b24j�"ObYqE "Z(t��T+&��("O�1p1�����TA�W(a�CW�HG{�򉄟e�~u+TmY�04���N7I!�E�D���E�P��2a.�}�!��>+��ٓ��E&p�T�A��^�N�!��(�6�0�@	ӘM:��֫(!�D�Ҙy�S��*ULT!��(N�!�E�r >�)n��d�D6�M(�!�D�<&����nɶL���b�"x��O����;��ʭB�� KaM��>�|D��}��K1�Ý<����gD�|�ȓ<2�`Cv�:��)F"�1r� t�ȓ��ihs��B#8��!%��e�p���d,B��3e�� "���)F����ȓ
}���$�A�HQ�U��LRS�>���zR���

�B�����Ćȓ|\� 0V˃�ĉ���'
z���	Y�? nY�+ҁ�:�y��E�I�ҕ�ȓlR(�Q"�2H�z$�"�ܝH��܄�qۺ�S B�2��5��N�:0��ȓYź�ce@��9� �G�D�wq ��ȓ.MkP��<"%��t�� F#���ȓ+��3�!�)<���B��K�����H~��K�5Ia�At�h)a�3�y��	���gG�e2"dȖO�����d2����
�lS4�b�H,Ò�C�"O����S8g��*�ቪsH�D��"O�T f�	}�^��5�G@�`"O$�i�C��t��d��9GA����"OJ�:U�D�>��z�,�H4�S	�'XD�`�E4;�҈Y�C�zQ�QQ	�'�$:&bБ~���s�H'm.��	�'��@�@V�P]9Uܨk�X��	�'Ȍ���Kâp��0�ԯ��Y:���'���S�D�_�: �� (�����'
��c�vr���Îٝ$(M��'c4h!F��]`bec���ND���'�,݂G�Y[~�M��F߾;�>H��'w^h�aC�qĜ��퇾<����'\�t��t�Rh"0'�"e�����'���ɲmҬ]7R����Ö��y��'LpD9���G`^� ��!����'���!�!+����O�}2���'������@�Vx�	Ѡ��sh@���'�	)ad�	��]C!�ޤr%Ƥ�'�����1[����CM��byT�0
�'���@O�l4b��ܞ%H���'q�i(Q ��ݞ��b��.� ��'�:e�%G):����ХF"�F���'��(�RL�"JB����Q���'(62�"��0�JiC���4`,
�B�)��,Y(`XfmQ�g�]� �B���<���ߟr^�[��Ѽ ��ˢ���!�Ĕ,,� �i
&]��j�� M�!�D%��P�MB��5���K�=!�,\���)Ą@/����f[~b!��/8o\��w�x3�)��GE	#U�O���-�D!�3� 6�yG�A'cR�{��Z�cvYS�'��' ў�OW�I�$��=5��e��B�1����O~���
$���Y�`O�n!��F�IL>�S�͉�6YRP��5���3Q�+D���V�J'FpP�)P�s=�8��3D��0rC�W���S0���|@JgE2D�,�P��I�m�@���\��#�2D�pw��B���"�s�p²C�O�C�I0����dD�aZ���D��:;ɂC�ɚ*��bj�.��̲�X�s��?���ɆK#�P����:��u��A�	�!�C,UA�(�+��5Y�,R�@�"~m!��H�eծ���z+�;��!�DIT��陁#nyԐ ��8�ў4��S�'���
B@3���޻V��C�I8Ơ�$��>�fD T'�.f�xC䉚����1�ɭ{MX�����1}�<�=a�'p�`��ρ@�Z�x��	g���w�Z�C���J[��A��J�
�Ї�<��}���W�D�l�@�N@(<������6&pK� ����PB
��'��U�?����~Z�h�#&�V#1�*i�R�*�[�'aax�Ăx�j��B�NY������y�΀:����eͦ\�20Z���y�HUlp� ��]+S<nt�fnH��y��N�3x`�k]!}�����B��y2�ȫtM��"M�!0��S�2�y��*�"��4��Ƣl(�M��yb��.3�`�q��
^>d�mC+�y�
�HoVq�a�� ��IAU�՝�y��G.YiBQ�r'A'w�������y�j�&���8Ďִk��![W��2�y`�M9X�!�ߕd`�;we��yR�/dŋpm�Ms��Cq'	�yr�K^����c�(2��}Cv����?��'&�{u�0Z���ZBHݰ&�.Y)���'U�8E�E5*����ъJ0���@�'s����>�HH�T�
o ���'8���2�K�5�L�� RA^�k�'�bD`�� �ẶK��B<
���'�Z�x�G?�T�����2��!9�'=�hXg�³c~��6A�4U�\]J�'ޙZEo�6ir�� wg�z�2m��'v��[��2Q���qF#P1~�.}��'���1ׂ_�/	���l�y��b��;����� �S�803jϩ(z9��"O�樑,v��,ie(�9Ng��� "O��a@%��f����ć[d0i�"O>
nŨ	w�%�CH�-��U�V"O|��sEz*P�'�(��"OjI�6*J�o�${f�H�y��"O�=�b�@=�-+���-8�py�"OҰ*HȮ$t�C(F@���J�]� ����Ic�h'�[6~��d�a*�j��C䉝Q��I���G�&L�]���H�M��C䉬2 y�|i�i��Ѳ �C�I*2�ĥI��J.�Vb+�)e���?i���S�OHTj�.B�	*��`��A]�UR�'?f�g�,eD Q�E(1!(�'iĜ�҂F+���1W��.)�-�	�'76������sY�H7�
*�J�'d�9h�3�� &��1AIb�'^9�*�<��;��N$��9��'K�	V���1<,c�IXSZ�a+O�=E�� 46��E�E�L;=���kfV��G{��	�:$���aU�/�����)M�'�ў$�<i㫕/]b�`��I��Ȣ�C�<�W���\�*T��?Jǜ-q%(Ue�<Q&M��� +"��FϚQ�Q	�_�<�`��.	��U��5�b\���R�<-M��S&�¾oq�5;�ԜR��ʓ�?����S�O���AJ�)H��{�*�c��y�
�'����'�x��-zd
a��E��'�\R�],O-^P�#ϜiJ�#
�'Hdp!�hˉaJ6%#��G�.���'\r (F�ƨ.���P�D�����!�'!8pS�HA�Ex4�w��x����'6��A�NM�Xþ)�GҿoL���'_����-g��֦�� ���'Bx��u���2�"
��"�I[�O�H�[׭B1u�L`�%���[�"O�y�$���L�RT)S"���b�e"OR�rΘ;<��̐�o
(��p��"O�\*��K�>b ZNʈ>�\!�2"O�#�ꊕ��mA&�Ѧmˌ��"O^�z�21���4Y,m�D$Y&"OR=H#J��^��䡆�ʎ`I�̀v"O>l��Ǝ6N=��Ҷ�
�g��"O��	3���<�N�P�D;�����"Or4���׬`���b��7K�h�x�"O����ͬ$�J 1�d��UX��"O�p3���;=�(}���9_�=�"O�T���ʆ)l��{q�B+�g�!��u�*@�e��k,�xAm�>c!�Z�b�c�
4I\���e�Ǭ_v!�Ā�_��h�D�8�V9sD��<t!��^ oDlYT�j�.�z	�?7�!���-�h�ѥީ/��|!DH�S�!���O��mIb��6E��H�֍�E֡�$�	f���ԫT52��XAV"���d6�O:9huEiGT��WD�&R�|�OrdS0�[:cD����g��G6�`�H�<�ST���T�'.��a�й=�"!��hP^�`�gI�U���6��17H�ل�G8�m�U�@W�����e���j ��:XL�IE��D�1qbˋ+qތp�ȓq�,�q���l�Z��-�^��ȓ�"�{�Ù�a �8tJ(_�dȄȓ6Ϻ4h�kP��Srj��\Q�̄�f����(3;���F�
>�-��C.�"7�Z� F@%)Q&��a:b���4��b�:a�fͨ7F�z5R���<H�@�!2�T�i&-;����=�9�LC*^V(	֥F�5�����LP�5���zN��< �QA��=D��G'	��@@� ��E}9qƌ=D�����T�`�fL�:�9Y��=D�,�+�n�����4r���a'D��
��P�0Od��*y��a��%D��	��'�~5���H��	���6D�TkW�֖KѪeI�I��n��A�0$(�d8�S�'Gn���V*y� ���(@.P��i�ȓN�B@K2��'>�����Im����<�<%�E�q����"�[!�ȓ9���6d�p0BE Z�h֡�ȓnv�+��g�6��B�0�D�ȓhg�$�쒲~���D36�$x�ȓ$���"Ʋ9nZl���/-�����S�? �Eh�ˍ	�L�9%�nQ�$"OL9���V�+a�%cC�E�h�Ly�"O�x�B�9|��� �o��R刬�A"O��pA�����JD�9R��̣U"O�@)�ヂ*�v<pb�v��Dk%"O|���J��0G����M�2�leH�"O>�+FdS�U_(Ȉq��O�t9�e"OB�ɥ�݌)3r���\<3�d1�B"Odu����1is�d����P�����"O��֭��	;ڹ�ŁR,ib��'"Oh�˗͙�K���'�QdT�@�w"O*PT�dw�\��5TL5h�"O�ؘ�� �zNp|a��õG=,L�!"O����.��Cnm� �9pTv�y�X�LD{�򩃼J��!;NŨ%�����cHD�!�ְ%�\��  ))�"5�#��]�!�S ��ͻ���1v�$��ᆮ}�!�'� 	���J=`e&@HѠZ�!�+o. ��0d[�,�u)"J�!�	j�4�c�.A] ϒ'�!��5f��H8���d��+�HBv�'2ў�>`P"�1m �M ���r���d�,D�d�'�"3ΐ���-�2H`�8D���F
,e�	9�Ϻ��õa7D���r-żM*=h�*�-`��=��B4D��Y�#�y#���2�!��Q��4D��RG�G�P���b
�a$)��2D��������kb��ZА4S�0D��a@�V��6�c!��$=Lȼ*6'9D���
�>f���k3*J���&<D�HYtY�1>0��CC�8h{pn=D�t�0L��90�M���P�>�7�<D�81"�%�%hק�15�xPcFM;D����I�k��8�2AѴe2쪁F8D��Y�ט;�]�,9��&BmM!�d:S?���U�N�]��S Eǀ@!�D��/t����|>���.c4!� vp�(�K�P682CN<I�!�DZ�2.�)�O�o28��׍�!]|!���'�0���I�/��Yy!�gئ�R&B~i:u�I�
r!��ڬ�`t���/�R����O$`!�O�X�Ve��c�`���fh�gw!�D�P�t���+T��Qe�66d!�ď:p��) �޹2�D�wbÞM>!�$[+ ^���'�0���Ѧ"\8i#!�$?�n�WE�i���8bY�0!��LlG͉4aޓ?�]����/~�!��M�Y7�֏U�=�*���'w�!�D��E;�Y� MؼF��u�
c!��Z�Qώ	⥈V��D�B��#�!�r��K���]�m��n 0�!�D${�41���v��͇N�!�Y��1�DM�R�����:!�D\G�
�����g4��i��ă
!�Dշ!n��cr��w9�<��N�Y !�$�& @�B#I"' QY"U�!�$T��(��%M�Q����Q-:e�!򤟸p
���䒊<G�P�J�!�B�"�ڱA �d9ʵK�Ol!�d��2Q��A�Ň,9���`'�3AW!�D�4u(#-^4$D�E�ԀOYJ��� g�,dy�& IJ�� k�yR�ϐ':����J�r��J5�	�y
� ̝H�+�?j:ĝ�FAQ"B���ɰ"OH|�chU0V��W-���%�"O�t�v.Z�-�*Q��K4���`!"OZ�y��L�0֌��$�
�����"O�d�Һ'>�C� V�c���!"Ot
��P� �Be9�F�L��!"O�=�u\)
��B����(�"O�
ՈW;v(i��/=��H�"O�eR�7�H�GN 0��,�&"O�MA�Jx)6p2�˳_�A�"O�t�'fq�Z����P�4Д"O���%P�jU���%$ۋ&���"Ojh��Rh���i�bE�YFlH�"O��{��I/�uh� �2::�ԛ�"O���6L��qגLQ��4����1"O��k%��>~qd�РOQX́#"O�M0�	��r�mr� �/݄�¶"O�Qk&��	vըw �;B�Z���"O��'U
����WO��k��(W"O��z��	a����$ǿ�jY{�"Oġ;�����p&��v��8�"O8�
6Er�r�2BS�*:�Q�"O@)!E�8`� �	��ܑ3(����"Or`z�	�*��%P7�`(V��"O�Q�tW�9s2�(2�θT�phd"OD�q��K
:Ȱ�H�<q�.U�7"OT}@� �pn� {�&��)�֐��"OL�sRm1m��K#�̰c">誠"OD���N��|2ŏ�1�Ru�"O�<R����I0v�@��2-�'"Oj���$z����"Q=�6)�"O&�����/K5��V�3muh'"O$�EҊ	��4hF�O��rT"Oȭ�E�M'@�X��\�MH��"O�Y��ъ#d���!� i�����"O�5Fi�(:z�Af��iW*���"O�\9�F�:��t�O�4>thc"O�uK��Z�('�S9D�""O��!Hv�2P9�L٤:j���"O��⧨�);xpK�i���t"Oڅ�E���E�6� �»d���ð"O6��$�� ����QJ����"O�u2�@U*Ĝ�)@+��R#"O
�2a�ƀ|2�5?,x��"O�x8@a8Z�:�`a�]�?v��x�"Or����W�]!�L1d2Ax!"O`�RӃ¶#��suE�8o�����"O���EF0Y}*-2��Ֆu��1��"Oй!S��}Y�#�A�o}�	Z�"O�����\2xYs�+�>lh�-�$"Obi0�L�p�RP�����(ZlST"O:�2���"#�|EI� żY��a{3"O-�¬�h�`a1D�E�ԁ D"OD��MͰ9�4�S�ܺ%��b�"O���+բ&i�@d�7S�p"Of�;뎚&T��`'��]��v"Oh���X�gF����ʕg�*0��"O����Ѐќ����Q�7�<Z�"O��d��qg� Y�� �Wp�3"O�s�N��Y�l���Y�&ؐ�kv"O���c$գ0����@eGR�ެ�a"Ot<2��Ϧ	�4e�D��"O��(��=BuX��ȌS��ĚQ"O�@�r
�/<Fd5h�V��f�hS"O� `��aĚ��`�ڷ�'d�H��"O�A��qS�8Уe϶/QRa"Oh���.�<���`d�[���p��"O|P@	�*-�&���K��(��"O�՛�%�2��e���rtP"O,�C��؅V�P��Œ22�b�"O�Q��j��T.�i�!$Ac����"O�tR�G.w\��
#��i(0l2G"O�a���E<0z t��$O&G&�E��"O谪a�ΝL�D�10dԡd���"O@�rpG�L�CԿ"�qe"O�ՠtd�Sx$"�������g"O<�ڱ$�4J�r�3�%�8#��x��"O~݀�\6*� ��*���M*�"O\�p�
ZW ��(!���@/�Ã"O�Ea�c�S[h!�
�(�`�"O�!�R�3��I�W�K�-�4"O�|r���+����h[�	�=X "O�))�K�� Y!#.U.�`�"O@�'I�+U�x!���ʨU�T��"O�]�&d"_�Г엇1�2̈@"O-�2䋦GN��)ë��I"OX�R��F�z�d�	2� �0�x�"O�s�A^90Xl��J��g0�eA"O2	�fI�?^�zY�r��&z�c4"O^5�3Myc2@��ş@(�0��"O�@��6����<�t]�D"ONda���Μ$�$AEo&�b1"OD��o�7p��t��o�<b���"O8T���"o�ɢ�m��,��g"O 5���%'6�)CoK�?��P�"O`RaN���Z��^�T� x�"OBPku+�W������2oݾ,��"O��y(I���[��T'̺ݫ�"O�����(WR��p���v��X)�"O���ԥ\q�t`��H�r�v�r�"OJ=��%L=Z�@#�!�W�T���"O2���GIq����E�O�^�ṥ"O6��lѱQ�1�͟Yݲ�j�"Ov$��-��<��eB��f!V"O
hRƚw�`�q�[�yG
("O���ʁ�N_|��1�T4��U��"O�p3Ej՝fB���7�*��r"O�����)�� ����"O�T#qeۉr�2D󲢇.��#�"OB�J��� :�.Y � �=I��	�"O��� � �dW�|�S����t�yG"OR�QaNJ{.����N4��b�"O<x�#�
;�Hi��l$�
�"O �z��z .0���P�?��з"O$8h!�CE*�@ڷ ]�]!�G"Ojly��՚r�0�C�U�k�}Y�"OJ)Ip�U���ӡ��?u����'"O"��#�3Ad:CӦ�IO�,�a"Oh�+��]��2ȣү��-9���q"O���5��!�*8b��P�w2
��`�O~���K�S �X������&���!��P�\a���K�V�����A�!�+d(���AO�f�����~�!�d:,�6t�W(�3M��P�BO���!��з9Yt�� *m�L��/�**�!�$�1x�f�5��h�!w�3y�!�a;�)2�J���تV�C�t�!�Ę�Y�t�P�0{�2�bSBS 3g�|�x
� ̙s�O�B���Hw{�[c"O�4 ���F�R����9^�MC���N�O��mJ�=��S��Z,on��
�'r ����R+� ��c�(,M�9��'�qO��}��-x�c;|� ="��@+XK�|�ȓ~���AMS&�$�q����O$����f-b1�UW�e����2c�cWa~�]�|��F�+,�RŠ�o?02<dSbn;D��藃�*���{V�+4�X�[�O9D��@��/B}��+�>���+6D�H�D�K�DD����V-_7�c�j5D�@�C��'��D8��J>ʹt+��3D��ɕ/�?f�5:5(
�:;��ؑ�2D�����א>����V ��Mr<Z�
0D���B���� Ө|zH0(�/D��#` J(	���E��x9Ь� J+D�x`�mޞg&%���ªl� 0I+D���+�=SN�W��,�v��$D��3ҭ�M�-ď?f���xC�!�O�ʓ:x�=b���(6H�J�MS�R�hD��
�R!q`D@8\{(��TM��BN(��ȓ$���L�#l�BZrH_�<��ȓ"����� hd�m�1��YX(�ȓ}�&a[�K^�)���D.�qZ�ȅȓ:%`��.�#'�0�c���r�;�']4��w�^"���*G�*7V��p�O.��<Q�4|��e�PW�Y�Ir� �1����\��O2N6�H�F
"�ĸyQ%�)4]!��p,L8H���<P/R��N�78�!�B�U^�� ��>�-
����ў�ቯ8��0AU� �;�x�	��"kx��"�ɓ�H��I�v��Xu�4!��h�&�&$�(mS�'%џ {�؊A�G�	�+��2"5|O�b��`v�T�Wf�s�F$%�h�"/�O��ɩfbU�b��5&�6 �w�\)��B�I�O{$�0��D�mHI%��3=�̣=�U�8�ddH��b������٨	�`��IW}R��ӌ�IB�<F�~ �P�m+�w�H�Ity�ȯ>%>-Kɟ�ref�/������;8�@̓s"O@1B� oei��@��p���*���'�bn�M�'��9O�4��LLfh�Ja��?��AK�O�0S��Qo�f��ʶ�&���$_UD�Dy��I�����@��+��)TU�\����*�k�n��w��{��M`�ݩ7�z��e̖�H`�֩�R��M�'��`���iR�����O>�����~B�Ϊ(`N�b�>8k��#���8���/�O�	#�,�>��qLŲ.m|���]��G{��)��1��,	bE�e��5�#OX�n�!�D��mv)[�]�K� t�"$ʁ_��	����'4�x��0A	�tÂh��O�]�c��y�ڼiDb�k��ڈK���x�����M3�W�a~rl���
ds��D�B�N�sw����>�5�����ׁk#���
��"�Y8E"D��S��X��𬂯C��!
p�!������
ç^��z�N�$?���`A�0RӔ��� m ����CHڱ��*X e�	�HO?i�L��M{�|`Ƌ�9L|���#D^�<��!���l�i��EbKZ}"�'Ӭ����9}�Ȍk�eY
����	v��1X⩜�e��+���.H!��hʚ��f�_z$��ʅ�F�(�S�O� Tc���m�b�X���c����'����T���D��TmŶR���r�'�4t��o�rӦ��T,6I|������ (H���V�F�T��CW�i�jЦ��4��I [��(�6%G Q�X� B7f�B�	\��֯�I-Vp#$`:I��B�I�dpj8T��!XF���9ijB�I�-�
}�
��� H9��{�8B���-�
��7� ��0�����Ms2�!D�� "�2��=!��)!7>H�� O��=��-��n�@(ӗ�@�b�zQ�g��<y2+|Q��Ɍ�e�Qp 
=T��F���_���#9F"�/:D�D��K�A!�ʔp��c�M8D������/RуM��&�2�x�E"D�4���>O���3r���"]�-�ҡ~� 6�#�O��b�֙~�D��f*?���2�'Չ'���B�j=zO���W+��{�J�
�'�Ԭ+��[
n�YWmY&'~���d�M���cf�6% ���Y=N�!��S��� �rN�\�e��ўd��I';�$�Dj��Q)�hN1'�HC䉰�|��Ɠ[��sW!�)KFC�	%5<���j+��!��0�B��t�8 ��6@X	#�eɿ%�vB�	S� ��F˶ �hZ9R�ԅ! "O.�q��P�;=� �ѧT1���a"O�\�	����
����Ќ:��'剜	|�@y�!Ӱl��|��̳d�C�$?Ґ��0�T�XLh�"�	IT|7�=�S��M�ԃ��Q�bJPIɽb��*�T�<q�,\�O`���7:R`Q˒&�ş��'��|��G�@��ш�E܂.H�t!C���=!�y�
L {	b�a���'Z X�����y�Җ~t�8�� &="�BFB��'^qO��|:񏂚5D5c�+�k���8ሞz�<�t���#�9j����x�'ўb?��ьϲu�:�x�@F�����:4����*U�"q:���=f�tU�s�qy�)�'&cn��`��c��s3��S�T�?���O�~�������,Q�w��5���Te�D��:5BY�Q[�m֏)���!!2OZb��Γ~�� r��dި8I'N�Ն���O9����#�~!g�r������<ى��S�;��L�a눉{4� ٢�ז�dB�1qN�Y�������I�E�E�VB�I0����#���+:X%q�߻O�6��d8��9K�rQ��Â�$�BIF��Y\O����kx\Pѥ!���0`��1O�=�|�U)��CD�!3��<�|���c�<�ᎸJG��@�/�H^r�+��K^~�L/�S�'D� ���Bˤm��B�̍2*�N �ȓt�d$�pĚ�jnPp�ڢj�1���d#lO��G#�L����G`&���D"O(
 L�%p|zǬ�01��"O�ih/�'r�Ƒ0sfԄ��P˖�$�Şqa��Q1@͜h��Iy�@_����ȓ��dhP���hό<�MGx�'�J$cĜ1dL�	��Y��'?�d��2��a�1`f~d�'�"d�@""���(A��n��t`�'��X��V�Ed\qb� �'f7>(�'�%�c)�<O��8ه��U�����'Z&U	����t\.���&��Lp8��
�'����a[;$^�GB��8��B�	^a~����KP�k��ހsضC�
>$t�ŉ[Mp���� ��C�)� L�Rf+�5���0�,��"O�P�D#�nxh-��$#���+0"OjP0$�%j���w$��	�H1!"O��A#��{�)���W�9K�D"Opu���ľ��P▃\=�L"OP9�!����@�V шL\�x�"OfY��IE1{�%���L.P]Z7"O�Y�D�1 ���)e��H��"On@S���9Y���s�ıS��T�#"O�$Ѐ#�Հs�a�Y[�ъ6"O�d��J�:�I1�E�$fИ w"O�)�9R�� pХ�\�հ�"OHu{�̓Dm�1h�d
<q�z�{�"OLx��Eƾ( ��uW���qȒ"O�8�"��V�9�2k� 3�ڑ�D"O��xs�Պ ��0Ѣ��/�u!w"O�D������� E�5F6x�'"O�1��/V�F8��Q3E	 "���S"O�li6�z0n� �_�N�P}�"O�QP��s��k����	�4�y#"O���c��0=v"�'�+���X�"O��ۦi6��yXtf��l�h�(�"O0�AE�(X2�9�c�D�.����"O
�X��Z�h�xQ�)*�����"O�}rd`S�tC19F�5uk���	�'<6�c���#�XI�@]	E�| [�'��Ĩ�� >1��bc�+,lII��}�65���1)���
���x�D�1�x���K�Q��(��|iL���E�'%��a����$p!�}��{�Z�@�J�8GR`����#����ȓ^ځ@��<����R	�Z��ȓ2�J�x�d�[m 0�M��M���v�����L@�+�b�{�Hs�⑄�N]�99��K|���g�ѱc�*���AfLZ���4�*Y���Js�@�ȓV�b|9���>3��c��+�D�ȓ8{�I�D���:
��` ����nC�O]�H��jR*�>G�B8��[ݬ��JB�8!���Jӌ��L����ٕ~�lHI�g��gl�%�ȓ	�^���)"�>P��I�TI�T��*�4{���1���iE-SL�&��ȓnf��jWdǠ<��v���ڝ��y���v@�H�̩��f�yҲ���^�5��.�!����з=����Dr��bR�Y������0��ȓL~zP�g� ����Q�܅3�>e�ȓ&"���oH�w�L�R�SC6Y�ȓS-$�K�ʈ�x�P<�3 \ �"���f�`T(�� tX����"�h=����k��EAd)E�m#"퍟D8���!̪d��<Ԯ�btGA�Mآ�ȓ!���Pe&���f/¬	�"h�ȓz��iҡI[���Y�͒#e�Դ���R��ī=;VX��oWH�@l�ȓ.�|i�2o��R���a�&97�хȓq��з	7_�u9;Et���'���wnƕ����V1B@�ȓc�8Eǘ�<N�� �$ձ\�~8��L)�I��)�f4�ɐ��*|l��ȓf<�mԤH
da�p�j�t�&)��� S�LEB��'�8�L �-�
4���� %J��X�'�\��¦�v�:ɬ�'q�Hs�.�4���[e"��H�(���� ,�� y*zX �"O� \m2�-�5��\�Aˍp��Ȼ �U��,�a3*H���)��<��*�?`�����W �6��l�E�<!�͊6 �t�� ��.��)�����<yC�M�Dy�­=\O�����9�
�`vm�y��	��'�����O;3�ra�E YjN��'�K�f�^0��y�"@�lQXt���T���`�!�4�O8��f℃\Ӭ����)�3d��c
�w��Hq! ҠZ!��77L��r�8k3�I� �*X <@�C՚*�`��N�"~Γ^
T�
�W/7:��yqJ�i�Q��9������Ϙ ThY�p t��I�y|��i�'B��$��F����
�J��ez���a|��
#Ḑ�e�ӣD�d��k�d�5	�F2p�a��'׮���AQ�W��-��������䟁?��u������(�8PI�Z7 �h g�]�>m(q9"O2h*B�\�^��m0F��7o�@Г& �Ĺ�uH^���)��<�Q O/OK���8*����\p�<�B�Sx}� ��]l��t����l?�3`E�-��h�e���G�EU��� Wb����	��"1��'��r��>FP"��'��P�<��'�l���%�	N��Cw�I*���'��mV�B8'����JJ?���S	�'�d�"J�"h���8V癈Bh��'�~(�����<�P�됞w+bɲ���^;�>9(��W����S��0d�]�oK�!�$��P_x�T]�d��!�n2p�]��A'O���hQF�S�R('��O����6Kv��(.�~��7"OD�8�P��%��x H���@@��9�s��Y[JT�'�T/{��I�^�Ԉ��;M�� "pD�8l�
��d��E��9�m (���Q�F��"O��`c��)c�Ԥ�sB�`���'�ea��JSB���AMGG�ȓ�}��2 ���K�e��( D���79�O��b3�_��$�k��D�2Vz͙	�'�L�
�͂0Jz�p��@�(^��ao�+�<(�$癀�A�����7
�,�I.�\�șw��К���P+Rh�Ј5q�X	�']�L��;�7��i�����!ʗK3N�p§<D'�u��-L�T�d��'~2�k$�ݗ��	=l���Sႆ$"�KfD��4�4��d��9s2���}��!�L�$S� �i��%����T�\�1Кt ��H��B�J�K�I��q
�'�M��`\��� .� |���B�y2N��~�����7h�4��h�-��wȏ)7�e��[�I�a�$O��CBڇ#�Y��'/���P!�z�b���J*�0R��Έ�T�'O~�ҙ�AB�#-�����|�l���j�(� z�w����5F�h}� �G�ۡ�i	�'����Ռɍc��X"w�Y~��e����Q�0��H&t��e��j�_x��H�,�a��pz�
�y��M��O$��%HBaJ��׌Ϝp�D�	�v�<1��]�\;rAS�B���%C�+'H1I£�.C���b�ه^4�͂"�$>��bĬ�+S֔u��	�;�6|b�˔1n"ɚ�����RjȘل+וO
�eKpi��L�r���J�nu������� �ѱH�y[c���N��AcJ�sH��'�� c�؏wZ"�&#���s��06Z�� w�D�@mօA"�9��(+EtP:�Ɲ% �䑛wo�U�A�'X-(���V0$�~�K��5j�}���C; ��q�РxP`1R�M�^�$�c�A�@�1��E�"6����O�r�(Ѿ,��'��)��Y*6�����[�:��э��d��2s�O�iC�hj�DV+pB |{
V�t��4��2;�:æ��6v�b˓>���`,;,O��[��LUߊ=9!�E,����V�t���W��+�nK�#��1��ն`LL�>i��'�M^�0���i��(D���Ñ\��	1��t�M;�-�H7�������s'N5 �l����c7�>���I�F*B+�? ��K�*P<�3$]�|���H!� "ZM ��UJ�<T����w�^	W 4�����X���۰<�D(�2zz���g��n#s!�J8����j��x�2h�L�A)8���@-?���`5B��7�е� �"O�5�6
Ͻr��m �B��$� �Ap��S�I��h n��Py�#}�k `t ��������
B�<	D �8i��xK�i��;��ġíѡE���v+w��b�����H���G3�Y$F;Yy!��H���j ��n'���f�F�W��	���,���Vb)|Oi�DꄖVy�\��3a[�j�'n�2�ٕ �V)��i����NS�R�~dpG�(�6��	��� "�zv!���Ԉ"�O�rU41����)�Tҷ�Ա�h"}���0@|��70x�y�@Q�<A�jTXP@�`��3$g�`ƬZ7�RE��EU�dC�I�k4Q>˓��8;��8�����[�&����ȓS0R|����l�F�rQ�R� K^�l��u�rm[�T+n����O�]C�:�d��qmH�y�{r�֝۞T��g��������TO �ք�`l��+D���
W>Z�^-qg7p&��@�+�I$V�Y��蔯~��>E�	��}��KH8RP@d"�L)D�����P�����K�_&n Q4-�;}_�"����	N��~Bi�)H�M�1�[�nɚ�dņ�y�k��(JDO�Y�X�"P%ƍ�ybI�#F�=���'eĂ��-
�� Ϗq��x�?L�9��q�$��P7Qф0�W-�7=� 9��-D��p3̝���,��/[� ̼s'�&D�$����r��8�X?�)��"D��:�,�
1�����?zٔ@
C�>D��Hǝ3^μa�`�fN�ɛd�>D��h4(W�s�� �Q�Jt����+D����$f|��f!M:L�6'D�l� �$kVӃ��.��ܙ���� I��eta|Riؕx30q	AK D<�u.�0>)�`�.A�xa��L\�{��4S)����ۢR�\Ʉȓ=�B��� zg^9�4���`�|������	�g�O6�#i�|�ӌ�i�:���k���y ���G$!B]B�nSL��3+-i��5��Q�FĮ8Ѷ���=�Ъ�ZL��~�� �u�+@�؊��U�U��K$U�.�H�㉒V�R�3s,�Uܶ�sPJ�<�h̀6m3~`p�A�V�W��X�!�'��`#��`���I�$�N1�
�+���@�+���W$��W ��V.��+0^�' \i��8|�B=K�N۔Q~�H��^= �7��!��]G0-��&R�}��ɂP�ڠ(ƴt�DҁXa6��G��-@����X@:%��O�"�+���M7g�q�r�U(:� �  �J�5�az�j�A�X̓^j��h�DηE/���d�Q�0�~iI�״SC�|;��N
�`�ח�?)uϵF+����!����'���t�է,��"�h�Z���L>)��CX������@RU�2'ت�2ԐթK���	�'��<��Q���l� j��G6�?��l��$4q�FI�G��y2�9��xV��j�Yv�J�T&%Ё�ì�1U�L�1�H��b�'2b���<���iÌ  �tR�R�z�rP��	\�2K��j6$C�ɽT�.� �GD�wdA:\XK��ζi~<����dB������r��d�V!��? Pp��z?1Ǉ��=�9X$�O�(�x2�݆Y�=�`"$,O^�0��S��<kܴ
i��T\- 	� �0��K����^}��ѳx	,e��Oqy��W
A����Lr�I�0a*W������5�8Od=ڥK��`e8�4E���˷��G�b��� M 'X�]�I�(��H��1��dQ��K�:�Gr���
�FY����آ;� |�b�A�\Y��E�Ơ���K�O����N�R3d$���S�|�Hَ\N@ �vb����?�Px���o�2�90��4��"�+1hn��iқ���.�,��f�n�>�) �n�D��|�n�7\�
��Q�R0[�4XE%FjX� �c�$c�
�y�Z���
Z*:���.�-��)��Dl�^Q{�4q�ص�M�"~nڮ/,� {Ce	,���@�
x�O��!���z���	Wed #�UNJ��#KY'��I�l��lj��\X��y���K��ģ���en�(X�ě6k-���=a�u�'UN�u���?K�`c�Θ	9�<���9D\�%��'�MԋόO�����,L��C����h�~����]�tY�� E�%n��!�CA"�!��ŗd�`T!wj�( �sR�A$D�!����`�pP�
�����NS!�#�ڝ��I�O�
�����%!� w�y�$�.Oٔ"t�)P!�dӃZZBa*QkRC����c X�m	!���+z1�(I&r��d�q�@�K!�$�φ�H$h�03�� ��34�!���~�0��6.ǁj��\��n�>}�!��
Y�XXcCY�f���@�^�!��O5��e��H��S�Ʌ�e�!��Q�Pd�O� t�,�!�� �P�c�P4"i�Տ�mX	�"O�%8�mR�#���0D�٣[�T�4"O����BOS$�q@!4��"Ot���B�*�3R��K�Q��"O<�����H?��� ��Z"O���K�#b��S`�C�p�L*"O,}ᔯ�N"&���Y0X�hٵ"O6���(��:�c7cP�P�XP�"O` r�F�M��2�m��~��4"O�i�ӌY4̖�a6>�%lO��y��ا[�����Je��f�A��y҉&0���0�(�NW�����'�yBL�=�f��̩~e���b$*�yr'S�I�v�C ��8`�ĝ��y҇G-"B�D�E� v��yF����y��{��er��}b���(:�y�Cԛ3ʘ����t�i;�H�y�䞁,<���˜�\�*�:!�R"�yB	�t���Q�"��U�>i�`���y�%�u	<k�њ������D��y2�/'N�,rC Ս�&��Rh ��y��I6O��2���3}�e:3���y���7ܮ%���
5��(٢ �:�yҀ�j^��CP� ����=�y��`��aϾ�����&5D�p���70��d�68��-3@l5D�hj�藇:�%�Y�^��c7E<D�p�bF��\v���f�U3��L=D�L{b,ښ,h�
�'F}�)ju�=D�8f�66t�k� �[�4�91F;D���2��y�ұ� �U>4��#6D�Ъv]�K��Spd_�jt�27D�D�2�Ջ@(�1�?�ѐV�3D�x�1)�h�EJ�C�	��a�#:D�����6W��+"ݍi����%<D��3�IǢK1�\8�iO/� ��(9D���ᄝ�nM�A� �>�ꠘB�4D�ԋ�^W�����	Z����S�2D�3�N
h�N��`�K?v����2E3D�8��4�>���"ǖ{r-
�#1D��(��&Tg��9��ѿ7��(��.D����dE�xAK��6�zܠa*D��!!��DX�X3���8�T�r��5D�8sB�'A�$T�C�^�^sD3D�����ɣP��l�q��.���Z��1D�أ�hK�WX.3��D=D�� 	T�"D���a�v���y��^?Q��QBn5D��	�Kфej����Oe����$D���M�\�x`�R�(�j)�c#D�h����nn���e�!^��1Po2D�Tf�alHU{��+*.=��3D��I��3s(�ّ�E;7P	��.D���𤘋+	Rܱ�dB�y4F����.D�$1��Þ*��ذ��/�:��d�1D��{w@�C���� 1T�e!�5D��qnO�e��&� �Xc�'D���N�9Ʊ�P�S�<^�`���0D��١�.�R���]�~zu�WC*D�8����&OC�i�O۪|i@�o+D��x6��	"Q<�i���6�HA��c&D��&$%=T��Y����0��Q�3D���A�G�7k���*
2����!2D�`�І�F��XЂi_+���ڤ�'D��h��߅>����%�ڷ-{�)׏(D�� �I�F�"�S�]�xK�0��'��)@ �$*CI�&g�H�@��������rd"D�h[5鍽{�ޔ1f��<Fl�\���"�K� |sei=�H�(���n1(��q���$�ʅ��"O��� 6��Irp��H����oذ}g|Y����)��<�qN�xd-��/� w;��T�Mx�<��%A0��k5\6����U�<q���)���a�%3\O����#ˬE����F<�)�C�'�,���X/�L����fA�A�*W ~e 		�	� �y����:ij�l�6l4� ��OM�@����&�(��Ă$	B
d�^�13��0A��S�"OY��� ��!�f��()��Z�Qf��`�H_#��)��<� ��1��E�$�~5"(��G�<iW�^�x�<��w���e�����`��<�g,CzXr�`&J=\Op�z���i�C�?	X��q��' �U�r���!�� �C��"�����m0Bԓq-��y"BʒY�H
�k��b}�q����Oꤢ�� /����$Xk�@iU�4#2p�R �Y�!�X	�����L$T���ψ1(����Ѐ��*ږ��L�"~�|�����U P�j,$�@�ye�]�ȓ_Q��X3�ʀH��L˲(H2f�h�ITP7��Ű=�`���&����!ȝd���
ҥFX���5��	B�E&,���L1hQ��,�$�y��؟z3�]����3�����ą�y��,ݔ���'Q9#,��C��y"fɨQb�:ƂAA���p�dѥ�y�Nʊ��6�M6.P�@�K� �yԀ)��MΫ_�`�Wƌ�y�EM��J�ΑLHμ���A���'Iʴ���R�S�'9
�*�̜<?6�H�HD~�Є�"�R�ʔjR.��cA����FQ�o�m�ɱ�LE��Oq)�%ά0���Ɖp�IjdO�t�&B�ry�s�,�6d�!�#�Jg,���_���>�0@'6Z����i�NR��rA��wX����RM����R�h�Ԣ�=E 49�a�0u�i%�-D���ǤK
��[�	ξW!�PL*�S~!� "�Aؕ�M��B4�c?����t|�9Q�B�#x0X(��+D��dM>Q����F���~�᥎I���+۾Bjn諁H�[�vb?%�Odhk�a�0c��x�5
'd�HO^tЖ�&]�򙛣LA0m�SÁ�n�tQ���߸8�P q��<0l��I�� �ʀ�ߒW�(|`j�"F!��D�>&�lm�� ��D�J$1c��$/�=��"�Pn���Ԑ� |��\s<�󌅠>�f�34��k�(T	�%8�\ ��-����Y�L��:U�ܴ��D���%8t�	���%	��n_�T�t��-�S�r��B��!�D߄V��;�lK�(ؽȥ��/��!y�� �θ��`�	YTX���o��% � e^@U9�NE/,�^p��O�������y�<H�E�-�H��I[wZ�)��]�r�hR�̣i&t��Ռ�iq2��$�'3r��C��^����v��	aO�eb�'�;1)���2/����:�i��Ǻ:R��.8L��M���h��ǉ``�(��ďi߈i��.�|�h�o^��ZQ��N�-e�bL�a`֩
�ꥨ�'St: ����UA���d����V������^eo��za�W{Sv@�O=��]Y�F��|���w�N�x@Ư~a&މ|"�=���h�@�@$F�d�b}	�'�Y�]�և��QKz�+��gv��eˑE�I�fr���%�1��S�~����e
/���[q��*=�џ(��"�/��aҖ/�2|�������@cœj�>�����$�h5���|��]$�l1��I3+������<r:0�E囚g�\˓C��`L�j`��#u��j�|#}�K�P��u`�"^-vl41y�<q�H^4{H�r�)R=Fp�	��E���yy�G�)6�"�sTg_�)Xȭ'?�ԛb��)zc$���lڨ�`c�)7�Ћ")�kh�IW�#3��U��ʝ��=��!Vv� $S�e��P97#Q�F���	Y@��ݰ�O.OA���fw�3cF��y2�g>�3ǓQ�F���A	��y/�q�^u$_*1Ķ�X7-Y8��'�n��6l|�G��됇@��8�Ԧ�4,�Y)6��5�y���-b���y�m�.[�`�V+H�+B�B6l�����:PQ>�S�? 4i���2u�Y���S(~��M��"OHI넀�) <)��,P8.�>4�4L|�R	� ��ă�|��qArخ��r�z�"ܷ.q�C��c�X]�� ւA4���	��y�ꝌG�P���/?k@�ywa���'"����N�P�t$��Ӿɪ񙗨�f`�8P �I�C�I-+�.���O+Q�paF�5N��͊m�X����*O:�K��Y�TA5b¨]�s�Eܹ[� ��!/D�Ќ׀TZ]A���1�lӘ�2��@(,$��J!�'���5S!`Z@ڥ�9$���
ߓ\_T�S��^-(�
6�M�cOZl+f�4t	���� X�Be!�d�t[�����P�S��[ i�O�m; aL(�R����0�`�F�uY�2��2o!�ċ�ٰ��jVH��C뙉'�̋��J�b��OL�}��9�xd��M�હ���,�� ��$B�䓼r��K�F�MB��ϓ|B6����>��=�B�CJ��yI���N%fmb���C8����Ʌ�F�d]��Z���n�=Є�G��,2�!��=w�A��@��!Su�ǅj�!����ad�@�G�T��b���!�Ę�}`^��ŝ�D�{G�~�!��L�cU8a��O㪬�T@D��!�""�I2bo�7٪L�m��\�!�F!L|ꅩJT�i�aPSU#|�!�DN�!].@V������Y�K�>X����VP�0��\��@Ӗ]3�0�$stم�0o�*����̟��gJl��%냯K�l���Ǐ,D�P��/����$q�M���4��O q)`�ϒ�~�eϡR����G��A�O�B�QG�j�)�)��n<Q��"OHi�dI�0�$0�%gG�e0��7�O�@i@sJ�Yw~�Q�'Q��Pb��h��Sq�{�+
�TXђ�,ON�����`�*z��05	�`�E�5,�M
pj�aB�$	 �&�?I�Y��N�)v�/lO~ęU�(d�#��	/s��a[��r@��\�����ȍ=���0�����)�Ŏ^3j���[wb����s�,"�
4v(h�'۸��@k��`pC��P6z\6AX��
�.���F�U]}��eaנ��+C�|J��y[8Yp�w?ęz�^!6F)ф�v�p�(ӓ��`R�*f���A�U1~�~m�b�Q;��QwkI(�q��ו)n��î�p�����'{�nu�Bf�
>���<a�c��98������i���Aov�h���/Q��P���N;O�!�֌@
�Q3���*Bl]���J27زP�s�^+-`M���x��8K���$?��]�
�8�hy5�?ZA�b%��pf�8�S��M��ȂX�<Q N�Gx��r�����
R��h�g/>k��,<�y��E��CL^�1�
O�%��HD�RV� J��J:�L� o�m�T�J��ȠO��{A��#���ʖ�ĬQT���z?�o��A(~K��M��8:�F8��l��F.,O��IԨ��v6��48�]�ʲ�����[��0�$k�K�S!�K�I��= Q�Mcy2�E�+�8�� �a�~����V03�@���oFwVO���e	�<����4k��=�e,��R�:�q��t��}q��n��
���S5Z�j�@��S�\��e���I$�'^:h*��A� \t��#�Kuh�� �B'`i��@�z=�ԉ4�W��h�0�ӼYa�ѻjP�6��m��_��ć1�A�fAV5���u�B-v�ب�E�$b4Pc|��b@g�z[I+���V4��'���S�*�t�@SN��*]3u.�9@Z���:-I�Jܶ��V=9l �$�Kc���!!M1Λf�G�	��� Hg�ӧ������o#�#d�����R�@������z����0|J��ǺC�l����}�̭+���^}r���7����4.Qx����S�}��9"�)��;�M0��P�{�qO$�p��@	���S���\J�@�{� %��i�`�B�	't�`	T���qKʘbC����">)��N-�ȣ|T�<(��S&/��?hpP�,RP�<����7 ���)��w������E�<�e1)�2�+�$S�R�١�%�}�<�a��F��KvC�K2�a2��}�<��JC����j��MG�%��a�b�<���Y�FE6��dɚP�P�
Z�<��k�$��$C�ޛ0��@e�P�<��8y��@�<��UX�+Q�<� �10W�'%jl����ш,Z�`�"O�"�S2�|�2�S�6� �i�"Oޠ���n0��a�T/��Aiu"O�����ОMU�-�BgM �X	�C"O���nV�>�y�#HA�,��"OpP��İ*:�X��S�1�65!!"O�#AF�1vq��"�����"O��J�DL�ð��ʆ��I��"O�\Ba���B`Bn �?�luӴ*Od�Kg�[��=���27�8�	�'��]�df�/;Y �*F�%�"��	�'�EG�D�i����/,l��@�'Ǟ)Q�(���L��ō"e�f�#
�'mx /�fz.��@�>^�0�p�'�
�p/4
��p�G\!y>�8	�'��i��W�� ��g���49ڽ��'0f�	.$r)L��e>Y����'�(���fϨ��i�Dȣ;���'��ar@Z�,� ���5ː`��'�t�����]�T(�A�.[w�Mp	�'��,	��R-Zwba1�W_����'�j%0�ƈ�3R@� O�W����'à����/�8�d�E)�)��'u�x��"ε��*P
M�:"��'m$�Z�Yuj�R��F�2�6���'����cH�,���fX2%$ٺ�'�6T37Jͦi4"Թ��(:f�'�~-���$(�F��$C U�&���':a[�$��n���\ �����'�~i�e�֓M���1허)����'��k��>E|�a�`���_�4��'@ �*�͂c��tBӥ֟C]��a�'����`��7���z��;�8I�'�L�鷈:w�ā��$֪S���
�'4���V�^<�%� �I3��˲#)i:��Ë�1-����|Oȝҁ@�Up,M����<u?�]��e'
�y�헰+�����������L���fɊ�ohy��,�D5��ȓ<�p0C7HY�{@�T�Hr@�ȓP��%��^� ���F�e����M�����G3V%�-�"NQ��b|�ȓ*T�ƭP���ӧ�	����<�ÇGI���O���J�)V�@Er�Dd��
&��'�`7��؍�'���B^w� �3?�')�d�$�4J�f<���V\���kFA��E�,OrE���O=L��W%]�,(�hT�g�B1B��T�|T�	U���(1��	�fǓ0��	�M�d�8 ���@}rh�6i@!�֡@���	Ll�OE�Ub�H��%v�u��h^B�HSd�V���Rr�7��%���O�?�yPƋ4%�А�œN�	�1Ad�L[�@I�A\8�'���	ׂl}@��"l�,xԜY�)�ZQr)��'�,Ô���Mx^Ԃ
ç)�R��G��jѨw,S�R�x��Ż�~B�=c�P����+����O� J��p��cyp%%�����8=|E�X^M%�����۞r��d9�����d��K�UD��!7(�<a�kFy��IZ�a�J����w
L����تΦ����,��	�'�8<'?-8I~�6#�20eb� �q�$�6"
�h2И�0#�V�m�;a"��}n:�+	�{Q��B���=�4��/O�V������������|xX���S�{��@�b�*wU�  BF� @�h���OV��'@�2S�W�?����j�|_�<еJ�xg(%�@K}"��.U[��3S	I%���Z �\ �+ZGjX 5l�	C�D�$�����x�f�E�~�>q(7���>sPF]JY�@��`��S�p�^3�ݠ��Tb�ѩ��\:�!�$-]��J�O 7.5ry@p��
%�!��/1�X��AӑL��(c�'�;e�!� 
g"�9��L�S�Z���O�i�!�d�>.(*yJR(�8φ(K#��2!�� ��S0��?iT���J��p��E��"O�)pE�ڸ��q
���7����"O��!���o�T�ZB���8k"O>�`%o��%���($���mrX��"O�I��ŨN�@"q��M���ɐ"O�h��K��P���	��=A���"O�;��Έ@r�� ���0/2F"O�%�`����	�b�:"W�c�!�ٳBl⸒7/��>i�	�v�ͧN�!�_�S��`��-4hf��nE	2�!��4d!�Հ�m���P�L�!�FY�<=�;U6����"�!���I#���'��I�pxQ�B�[�!�P�R��A{U@V�H�P�����&&�!�dUz�>�o"Z�&H� ��!�DX%=��b��&Z܈c�.Sk�!��-_$*w[�byI��"!�=~�,���@e>NEZ$��'p!�^�@�Z�0��L����-z!��2�`�"�F�SH�!#g�<r!��3WO��j���a>��B#&�:gp!��w`�t%R=r{7JB-S!�*W�|{���-�T���F!�%)�����_�m{�@�fA�$)!���{���;rT$d ����>Yj!򤌆@�T�3b����E���]K!��[�R��!S o�w���(r��y�!��-?���J>|���T%�?F�!�d�.���g#R�tx�U	��aK!�D��_a(��ԁ̏P�ĹQ)B�#F!�כ[� �k��(��	1����m�!�D����4#P ��0Z� T�A"[�!�W�y��q����O�@�	㉈�!�L:o�.Q�q��6�D9� ND �!��0-PZ���ʅ
����Т�!�ĕ�GjLfB�Ut��qɅ�!�$=xޑ�a�: �r��6)���!�d�&@E��
Ԣ�F*h��P탄b�!�D�>|�t��$�Ux��<�!�d�F������'���ǂ���!�$)3��c��-Y4Re)G�N�/�!�]%o����ʰ*w6h`�R�y�!�$�?����ӛjZl}��`	J�!��͒Lŋ�̃{���@" ��8.!��LJV�P�b*��e��rr�̇%!�DÁZBJݲ�	�r���3��|�!�o���`$Z�t�0#� �!��4E@0�#���4#�aD�!�
'��4��([c`��+VN�a!򄛙R�&�3&�8nC�11�lS6rP!��VG;Pp��M�P*Z}��J1%�!��Ǟx	�B�3��*�jѵF�!�D[>Y��ģ���0FըQ��O�!�dNcs�HA`��� ���*�!�d %-���1&a  �0�RW��*U�!�Z�4�& ��LSX���g�<q�!�d:9<�5q��4v��y��Z?\�!�č��b{�M��	�R��фW%�!���}P� �`߇�4M(���G!򄀃=F$`%FP�d�8����ZIV!�A��� Ʈw�y �\%SS!�$������-�-a��7L����R�5�r�!mڹ�lI��y��֬P��D�!��}ɦ�9&ڗ�y
� �D�g�ʁgF` ���!j.�#�"O����Z�<M��$�UW��Y�"O�a����"'K� �C�<o6pI��"Of8{�C�>�j&�<`%pE�7"Oj��b�Ēx{�HE�]�5�Ekc"O�)���\&0�@8����2�`"Oz���ߋ�2��v��	� �r"O:����
)��|Z�#	Q�ؘU"O��q��#ҭ��E%Җh�2"O,���/�`����#�+)$ʬ�C"O���D� �TK���d`p�"O�)sW)��Z��#\K�l�"Oʴ�P�&�>�I��k�`���"OΉ+��ԇX���X�^]�~@BW"O��D�ϯU�����KW3v�� ¡"O����n7����٢#��	b&"Or`z _�
�xE�s��r��a"O���&-L���A��_1R%09"Ob<�'gq�0&j�1��I��"O5�$�B�E]�e*ѹK�}��"O&�xD
N�0i5d�xS��i�"Op�P"i_�1��0��P�'<L�5"OJ��t�V�H�� �%[��§"O�|ђi�"rHhׇ��pҐX�"Oа��C�$���ǔ$��u�0"O<���gÈP����2&�-�x�W"O����
�HO�Ar��W
)��iB"O*���ܧ|X��{��Ü)�X��"O��R%́�#��cg-��#�V�iD"O��qv��B�Ѻ�픛"�d�S"O
d�d&�6��X�M�d.�qW"O5rc�7>l5!���Ѵ(�"OH Z� ˕)��`+2%��[�t�"O��`��8��ph�a�z�Q
d"O������(���OR����"O*��uAH8^�~9��d	�\�R�"ON�"(�;��	t)�._�,5�"Oެ���3�j��'y�.�C3"O|��n�r~���`��;m`Z�@�"OB�+pD�>ڌh9�k^�r�z�""OD�[�N�7'��y��a�t�"O��*���k���U�/b	I6"OȰ!�f�,J�COQ_���V"ONI�S�ޟSs ����g��%"O8���K�{�������|�� �"O0TZ��H�sm����K����"O�%���()���F� 9�(d	P"Or(���f��]��Z�7�P�q"ON`��c�d�YC�k���*V"O]���H$"#j$��l�E�z"O8���ӎ{���I!0�d�a1"O�l�kȗcGb����kYr�qC"O֥�U"���Ait�X?�ũ�"O��{��ѯ2�@,	��̵P�0�"O�;���a�U�� ԛ=A� A@"O$XV�v�� 7�1|���	�"O�`�ǟvg�t�U �V��e1�"O������4C�,��(Ȱ	5�u��"O���#�X�{�����@�&y�D��"Oy#畑 ���'�D� \{ "O.Q�C�Q3
�� �wE�]1֕��"O�9 D_�"����]5x����"On\�g���p�L��N
��"O�FI
�phQ���
Ҥ��4"O� l!pa��	�d ����/��9�"O>�"�[:J�0�"��s��A�"Ox 4
�:|��1uDFb"O8�1�˞I���&��d�)�"O�n�*��Dh3I�����OժD�!��Ƞ@:ݙ�l�j���0��!��Je4���J55�Bu��D�!�ć�?Qr,�g��*�	`d�!�D��V�@кA��"*�j��D�!�dD���1,�!�F��UÁ�_�!�{G��6AN�/^Xj�!�H�!����@�Bd"\�f)`���4�!��V�j��M��-��`p�E/�!�$�L�Pq��C���=;�D�F�!�d��Y� ���
-'��I���P'Oޡ�d�$5�
�p��:}J�`Z�A��y��� i��S��O�]k��i Lӊ�y�Cݽ|#�K�,C�H�ɛ��V0�y(C�nhct䔤R�tH!d��)�y��]1�̀a�ڟ���
����y�%����9�ԥu����D �yb��r�ŋ�'o(D�5��-�y"'S���p�sJ|H���d7�yB�NFP��e�)<m��(�	�yRlZ�r�B6E���!�ϵ��4��'���@eD�1=�A+&Ɛ+lX���'�4��̗�xO޸be'�	r���'�^�J�V�9�rk�/�+�:Uq�'���QmѢG] �td�3
z��'�*B�@"�@�3JC%����'w���fȀP2<�B�+U��(�r�'t�����W�������Y��)q
�'^u;fE�9}�0�K"A�����'��	�n�?w����B��<C,�J�'����a�Т�F�5����'3���@�1��`"6��,&e4p��'��ԁ�Ɍh U��X3�Xx1�'ǾMA&���S�X!*����h
�'֌����+U8Ȑ�tO(u \0
�'�����.Km�D0�	^<t�X�	�'Bh%7��w�pT��9 �D��'p"����X&���#]&Q�;	�':�`E��q�<P6��C�
�
�'Ѹu`Qfխ	e�l��4�\�	�'a�})΄1l��A���W���\�	�'ox9��j�T|ma�\�_���'�x,���	
 W���b�� Pm��'J���e杹��,bả�f��i�'$�����6^����C&'���R�'{�E�biB�{�0��#���P�
�'�B\��c�%#� ujG�H4���@
�'�Ι*�@Z+L%�D!��-#�JiB	�'�xe����b�~l��-ƍ!�P��'"����L�e�h��2l�
eI�':Z��aش"*���e��j	�'l�idA�O���A�0$�i��'��4�P�	��+�F�#@*�@�'�D���Kj�^�"��Dh5��a�'JhH����L�Re[W⑴p����'Lb�"�	qF�]����#��Gy�<aw�'\��UrU'\-p���AFPt�<� ]�L��@��E���m�<�4��0�6i��[0ޘ��#�	f�<�2�����dE��)Nq��hM�<�+w�   �   �  ,  �  �  ,*  u1  	8  "?  eE  �K  �Q  /X  r^  �d  k  _q  �w  ~  W�  ��  ې  �  c�  ��  �  '�  ��  /�  ��  [�  �  J�  ��  A�  ��  ��  ��   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C�>����鞿6�!d��x�^��I��~�!��
�l����v���:�9a��:uZ!�L�,Ƞ�#g��UԀ�e��t�!��v.qc�ʁA�P{U�C-h�!�DD�x>B��cG;c�lK�,��"�ayR�	� Q2���F��u�t��� �/��C�I�Ld֘8����D��T�U�#�fO��=�~bh(e������M?��m���Tg�<� �������T�����R�g��dR"O���ѣi�A	�͖<|l��"O�ȁ�N��SO��µ'�#{u�L�"Oҕ�sGY�>u�0@�'B>]ԕ�b�'I�O 5j����)ɲV�л�"O"}��J]�P#JLa�׊R�Q�֓|��S���O��Ḡ/��l"�88�n�:!�D�	�'X���P��u�҅� D�l7�<��'{���6f-虡4��	.�<�R�'L�Q8�C d� ��욯zA��'a�l�3�F!C����4},0|ϓ�O�4 6g�'���z�h�!�P�R�"O�$Kue��Vrl��MΈӲX�S"O�!X$�ZD��z%��B����C"O:0���b�V�a@���VĪH��I8�\��׆pT����Y)i3	=D�$�&���;�#!a��9��H7D�|��BP���x� 脖~g�T�#5D�H��
�Kh��Fo�Z�s#�'D��)F�^��$H�/ǐ'��(#D�8�\�.V>���bYO�9�4m%D��3"�Pq�f�2P.p���(B��$K
~%x�b1Fb�la�CN�.��C䉮T��[#A�$I����(��AC�C��H�XtN)qH�!!��A��C�IHh,����s�6C K�R�jB�	����#塕��Z����}�B�ɥ~�� 2
?<�[�"��nZ�B�I)&�ĝ[uj	�%��a��;�hC�	�f�-� ���=��d�E۸a� B��;}�܉�e�1(��1��ġ=JB�I�!�\3�oԾ�p��C2h�C�	FxXz�g��dp�Հ	c�C䉇>�6���a9yVa�W�vdlC�	�!2,ҧ�?U�*�����5�0C� XwZp''�q�1c̀�ThfB�I(wM��+����k�I�@�ӽ	LB䉆���F^�=*Q�@GB�	�4�ܵ�!�� (Yv	`s��7�B�	?s�r��d����hj��I(8�C�	�g��d,�(M>�h�h��q��C�	�TTx�5��<�� ��&��C䉿[.� �� �a�P��/ԌV�tC�	3F�!wFY�b �'NV��C�	>=F�m�FǵxZ8U�ց�	tLC�ɦ:�p�n[�u�ҴY�!ӣd�BC�+;���U&�<b��T�@�����C�	<+A����Ǜ �R�I�.ݻs�C䉂Ԫc��T/T.nL���ܴS�B�	->�N�9�N��T]@xËZ�a��B�I�E�Ĭ1� ̮j��� A��'�B�I8[�2�r ͫ���TP�]`tB�$�0C$�!O�偷ƛpuNB��]EdP�o�4'��m
D�ُ9.2B�4$�t(*d�8X�}cRd�+DB䉷L�T���k�2n�i�CE�[SB�ISQji��6��{@��/'�C�	�sϴ�;u
�?�X�:b
��~/�C�I�F!*t��N�:�0�h�-	NzB��<�C��3}"%���CW@B��&`H�ܸ�Ζ)��p��+� .fC�	'�n�x�$t���2�I8�^C䉟2�F�@�╧Nt��q�ŪXtB�I15D�"� 0h},�H���yA�B�)� ��aF�H=�`z�aN�'b��v*O��xc���2�~�0����}��'���� 0����
Wl��*
�'��ԁH>pxcG�o�����'\za�2mF�3��H��ˀ%o�����?)��?����?���?���?Q�=�q���-xpB�ѧ�B�j��9��?i���?���?9��?a���?i�vD�U����;�Pĥ��?P����?A���?���?���?���?q��S�x�+��� &�h	���#OVlI���?���?���?���?���?��j�$X�գ���l�o�d����?a���?���?����?A���?��(b���[tu��+�B�h�J�2��?���?����?���?����?a�I$>�K�m�����Bl����?��?	��?���?i��?��,�lyGm�1��x����n��,���?��?���?���?����?��g�x˷EǂP�C���'�
�C��?����?I���?���?���?�7ⴹW)>��
A�������?	��?����?i��?����?��s��A�N &)*�n_�a ��0��?��?1���?I���?����?a����*��)[�|��� ��r�J��?Y��?���?���?y���?Q�z�(��P��
^CB�ve��A�Z)[��?	���?1��?)��?�c�iC��'�:�i�ƩQ+x��r-dԙt��<A�����0�4)�f����s�P�p��&�:�S�C{~��nӘ��s����9��S�Z�A�u�_�ƚ-��՟�R�(����'Z�	P�?�����uc2&MD+0�ѯs�du�����Of��h�d�Uk�19�A�v�R�q�2�a�����#1!#��L�'Ad��w1���G�[	7��%�ECN��xM9�'$�?O��S�')����4�yR���B�@T@��)T����pM��y�9O�����ў�ş�%�dȌ��#QV5���%`�L�'�'67��-�1O�0�vg��k��Lץ
�ؑ��/�����d�O���u���'|��Gw��Ȃu B�}{�O4�DK�1
>	���I.�?��H�O\�p�n߲iM�:Q�F�Bc�m ��<Y(O���s���$ޑ6��$ѳMyE��uOv�`�ٴX�t-�'f�7-+�i>�ꖉ Q2�8��Q�'�a���o� ��ß@�	�ED�n�q~�=�,��&c�<hJ��~KL,�&ş)���#�|V����p��џ�	џ�Rp�N
W,
��IV�LH*3��oy�u�mIB��Ot���O̓��d^��%D�8Gr��i���Hb�Ʃ<����M��'L�>���O�;5($s �� �h��MM�Kx�S� �>��@jhy`�ьO�ؖ'c(`�C� ��,��D�	H��'/��'�����S��ݴ`� 	�@F��	�/􁻂�D3`.d	�Z�����g}r�i� 	l��tK#�^�p� �G7Y~���D�Uo��m�^~�닥�ܠ��w�'ojk�3=� !e��!'2<)�+�T���O����O���O��$9��b�.Iy�$:?F ���>/�(���՟���9�M�$)Y���dNߦ�'����M��d�di6�ώBb�(CUFN:�ēM���Fu��	]YD�6�7?!g����(� 
����s���?�Jx�$��E�F�$������4���$�OX�$R)�e�5ᛧaU�l�FnUd�$�O�˓Z>��.M�\��'erZ>�05#�+$�����LDA�=�l)?�_���4 ��v
&�?]SGKE!F�:�tB��@¸��4u T0h�I3���|��`�ONd9L>9����IF��Q.2�Ψg�ކ�?a���?����?�|"*O�$o��Zm�U��h�r����L_!h��I�������I��Mc��B�<�4w���E픧��=9� S{$��sǿi��7mC0H+�7�??Ae힧����3��[�j�x���,Ү��qe\
�y�P�L��ܟ���˟(����ܕOΰ5���m��eg��$��XXmq�(x��-�O��d�O����dD٦睈B]�a���q#~-�
ӈh%ډ�	��
O<�|z��0�Ms�'�ص 7���NcHLp���A#��؟'��)�4Ǆş�$�|rW��S��k���FTn��"��6%�Rw�\�������	hy2�{�T�*�OF���O��.���P�C��Ii�r�Э8�����D�O�7��]�'e�:D�P�1R���i�d�	ǟ$#����2U#B|~��O2P��	�x���0'��(e�(ј	h4&ז�"�' �'E�����"�!�3����^�qo6`x3�C���4.G~�S.OBl�l�Ӽ#����Is�y	V�A<e�L��E�]�<���?��i0�a�ia�$�O���WJ���!*�v'z���n�4���2#�F�RUp�O���|����?����?����>4��D�5����LN2,.� )O�o��+�m��ȟ���X�Sȟ��G/�-?�н�d��Y�b�*�(C����I妹��4Sg�����O���H�3U8�UY�� Q�YggI*Ly EY��d�*\�n����*h��Of�(2��2�K�4�X�d��蚘���?	���?���|�+OzUm�
INL�ɺ/?� IRa�8:x(�cC+��H��	6�M#�2$�>��?׵i�\��R�*1ՎQ�G�N��Q3#7��:O`�d>Bf�Z��Vb�	�?��=� vmS��A%1TCV:l5t0s�4O���O6�D�O$���OZ�?ᘡ�.n�Ȉ�ɇ8�Z�#"��Ny��'_F6��+5�)�Or nW�	&P(vă����j�*@M<	���?�'hҰaش��d(<	��E�ϢiR�|
��G{J�#�C*�?�&�,�d�<ͧ�?a��?�U�O�"ߘ8{V�5i���Y�	�?!����������ٟ��I�� �Oh�I���.�J�*��6�&��Oܘ�'R�i��O�S'Y��YA`�<1B,�!!���t�Dy�eo�()ں�s�:?ͧZP��DH���bd��q!�M��1��ɮ�	���?i��?y�Ş��d�ͦ5q���$u��j���v_����+^5A�X��'��7�>�	���pӄ�b��;L��6ʍ[=���EOH��P�4*;r�4��$��X;~���'��5��]�5ɂC�5{��W"���Iuy��'�R�'���'��[>uP�Ɠ�e���QBOϫ�j���gۀ�M�Q�?a���?�H~j�v}��w�"𠱩�
,��(�EC�g�ԵSv�b�v�l��<ɪO1�0�1�}��ɡv�j����W�Jq�偄�qUd�	�js~q��'6H�&�����')n���J�X�����V.TEK��'��'m�Q��"�4h`Bs��?���'�N BT�O9z�*q��@V���i�B&�>Au�i��7�WC�ɤi��9:R�II!b��2
F���*�#ϟ�t�D�|�c��O�D��0��#�d@(5�pBvI�(]�
�c��?1��?���h���$Λ<�f��S�[�8s�Ao҉H���Ϧ�P�B��D��:�Mk��w�t�d��3[˸p�WlI��`�'F�6m�צ5�4}��`�ܴ��Y L�6 ��z�v-c���m��!�@�~���cB7�Ľ<ͧ�?a���?9��?���1]lM)eeA�S3���r�U���dW��M"q�ןX�	ڟ�&?�I2de<��4�E_@�y���إ
��IY.O~�Dr�>]$���[�Ş_4�ځ��o�(M�wӄ#��!���\����B��f�	cy�
�nH����K$t��Y@��f���'zR�'��OL�ɪ�?AE����@g�ż'�� Y��'g�@H  ϟ�a�4��'����?���fk�QθZ�K[vhrYyA-V�2�h��iH��e�X����O�q�d�N�& S�b�ײ�0�����Z>��O&�d�O����OP�d1��R�L0B��7�^	���->t2��'$�ix������?�j�4��7����N�.6�6�`F���\0�x��'��O �Ҥ�i��I	T�{��&L&�`��ǌo�� �p�ؿvn2"Lf�	y�Ob�'�Ɍ�J�4�A()8[P�ԗ���')�ɮ�M{����?A��?9-���(��Ģ|.��S�D�	���8ѐ���/Ot�$g�\$&�ʧ�"�c�X�n-�HA��:G�2�#��D�$�N���"}~�OT��I#z(�'���3V��VT�[r�ϊsjV��V�'sR�'�����O��	��M�1%KmȾ� #Z/��
�!��zF���.OT�l�`��/�Iݟ�w��	[��ٛ!ǆ�}�\E
\🸠�43�pڴ����H��Ÿ����+Z>�$��2�r�U�1�D�	my2�'���'���'��X>�WDF3Ӕ$��,%s@]A����MK����?���?�K~�F!��w�h9c�[	T�V��W!�_wZ����'�2)%��)��+��6k�� ���M�p�!�'аC��б�$r�����#|B�H]�\y�O��Dؼ�p���f��سQ�Y�4��'���'3剸�M���I��?���?�sd��l<dK�C��L�2`C�����'��ꓬ?I��H��'V�Hq*��Z�,ʳ��)+:(	(�O4�ٖ��(J P:`�IN��?`��OF)x$$�3���Ԥ�<�l�`&��O����O*�D�O6�}:��4&Te*��4k�t��0FS!{GR�(��K��f�ɸB�'�J6m3�i޵����u;����$þ���i�j��������;ش�R1޴����(oȤ�'|�8��6?��H���9$i��*v�7���<ͧ�?���?���?���=|&�u�aE�L��%9uFY����Ӧ�1
	�,�	���'?牝T�d-��!V1b(�3���>�P�S�O:�mZ1�M��x��t���k�$	׆��l?�0Y%ˀ��T�aH����Q0�����!"ؒO��.Ɋpk�@��#J�����|���H���?����?��|�/O�oq@v|�I�E
j�!�J�� �VA��ɺ�M3���>����?���i'H����?U�zh!π�(�S2aWd������lA�S!������ld�Beǡ�썣+��H�B4Ot���Op���O�d�O��?���E�`�8����U�3
d��b�Gϟl�I�d�ٴfy ��'�?��i[�'&黳��-������
�i2O�W웦�q��\|6�+?q�ȆD�ШB���3#7�#�윀r���H�O�9;J>�-O��O��d�OĽ `�����)��� ��E�g��OJ�ĩ<�'�i���<��柠�Oz��(�	�H�Ĥ� d�zX��O���'k|6MS��i�S��du�|B�I�Z��"�F6Q��	V'uSB�RS_!��4�P����ָ'?2�h��M�8�h�A�.x��	�'�^Dt�/ƺڂ� ?tI�	�S�~�-Дh"q�A��Q=�P
�e��5<��@�쟃�С��B�ncn���@NR�iX@���HvgĐd<��6错;� Q3�O�R�\� ��e��oP�yh�͹pT<"�̟E�V�Q�'��0��̛���4/���H�B ��A!"��*��Ap�,�8���f��[���,o��kf"O��g�F8�(0_XeX��S���pT&I�c��'v��f�7��ݫd�L�y �E8F�F��q�Ȳ ��k�� ��D�F�[�|��`�`�����N"r��4���Ŭ<a>�F��e�A�!��F|-�FDN&aI?:<z8H!E�bXlaH���-H(5*��.$���%"�K$�� �c�O\uP��� >�6q"D�K�9C6�9Å�O��d�O�,�@:Jy�nW���y[�IG��������X��#E�k���Jg��)�(O�<s��*�� �	�Y�"+$�r���T<E ���9P��a�'Ot�'r�D����?�O~����t�z�c^���´c�:��$K�����?E��'��	�-��`8��`��,�>`����'�'�����
Roâ:�&����O���D��P䊦o�m�R Y`+'4!��թ	<��!�1Bz<�ꡨǽ4!�C&��A��;W Q�pHߋz�!�$�2��|�Df��| ��J�AH�Z�!�d9�Z=K���bg��%��br!�$g��e��m�� L�9�4BƃXh!�$Y�f�T-�5���B�XZt�@�y�!��i���`1�Q�T��
C���,y!�T�{V��%/���P]PP��H!�D�7Ul�@���h����Lև!!�䕘6��B��Q�چс�AJ�r�!��4 Vl�$J(P�x;6�)=�!�ě�a�H�8P�%�9��$�x?!�d�/&�b�F���l��S7@�!��+ێ�(�NA�+"*Q�� �2r�!�d�Q��"U#H�a:(PoZ:9!�$D6~=�UJE�N% Q��՟;!�6NS*���	� �'�n�!�$T�r�p�ra@A���u�<&!�DQ�.o
��'�Z#'���׉�2�!��� �@��A
B9��-Q��|�!�$D<��y	d"F�b�^1"�m՘x�!򤃪q54����YXX��l��r!�ĝ�[�6��GBY��{�K b!�DZ%�X��_�8�x@�%��uK!���*N����(����cӶ28!�"z��Lyˎ��jd��O�_L!��?-h�D� [5G���V!�䃠��(z�SN
}S�f)R!�ď�{��S�'߳7J���Q�T M!�&>�$����
n*�U��O[d!��s�<�)��?t�l�ir��RL!�){z���n�;u�>��Z~�!�$M�17[Q��E��yұ�л�!��g�A��{��I�V�z 衇ȓL��air�O�E���Ƃ�4`�괆ȓJ=�!�*w�x)�JB�d��"O��bR!JZ��݁B%��g}t�KT"Ov����&��)���)���z�"Oh�wM�0�p!��u���(r"OL!	R@>R��a��f١��R�"OvL�7K�e0�����ߘXՊ�s�"O��%� =hV��U�nӪ�2�"O�}x���ј�cW�W�N�V��$"OR�ă��3`ٰ��W�N]�a"O�Ps��ϻT
�#
6`��m�V"O:ԃ0-� &���cJ���[�"Obm��a������#��BGJ�k4!�D��N;��h���)eF��b�>!�d�#"^ �B�B�B �͠���EG!�l���k��W�H̢I�'d�>?!�D��Ji`��Q\�,�QB�?.�!��C7'�8.)v`m�7IM6 ������ i!C$µu�p�n�30���"O��A�a[�F,,l�-C&�nyx"OB�0d��2HL�x3���eې�"O&M f�G0
8���.I�bl�q"O�xcGE�X$A��+�|�"O�ѣ�FG����Q�N-SC�q�"O�B"��@=�H!W#�+vEp"O~���X61���g_�"l��T"O�8I2�й_Z ���'˥����"O��Zu�h�挠��� LN-J"O:��чѧD�9�4i�#7�t��g"O>��C	}_26'Y�<%R�94"O��B��������ܪR��A�"OL���"�=p',ac�Ϗw.c�"O��!��8M�H��/#����"OR,ٗ�qIr��:E~0U��"O�+��"���bg�'5{�LJ�"O����n�S��qq�JE�MD��T"O��
'� 
�Xx)C%'�UI�"O�p���*3`�9Վ��.�Pl��"OD8���܇pI�`9�&��T��*�"O��Y�,���N��e/�g"O�yg"�/v�$�H�#]�*,d��"O|��p�Z�1!i�R��A>�y�"O(	榓�]3&�+rb82�"O��sVk� j�M��K^�K�j��u"O��!��r'��:3Ii����"O���Ǘz�A��s�^(�"O����o"*469 G�HXŪ��C"Oĭj�DI+!����'+�=�S"O���0��zڂ�Y��Y`�y"O�!���>^��)UD�_\]P�"Ob]��HV�+�\y�RC�]�։)"O
�fE$ }B�Ŧe���"�"O���5�V�?�,����Xئ�	 "O��2��������#��9��"O$)ht+�0Vs!���'=���A"OVy@oϦb$ ����A���"O�E�N�`� BfݿK�zE �"OP�A�'8Z�����	�$;PLB�"Oބ2��ԌPW�p8������"O��� �]�%�X�* (V!�@��D"OLb׹�V�ز@��*_�P��t�<A%���}{�ms����"i�4�]G�<9�/�2q���K_=b)x �fQo�<1�4a����ڒ!|�4��Q�<�LT�P,h�!bU�P�:�[��q�<	�	.XP�S��ňb�y�"��q�<a��ݒr�&)X��
�d��f�[l�<�I�7 :fa�k�8���ʑA�<���6N��Q�g��V}�`�+�{}�Rx��	���)a��FF�_�����%8�O������<�N�LѤ0�&mj+1�o�<qS�D�;	�-�DI�D@h(0�KZC�'�rHi�0�k�uc2�1*=
��� �2���O�����G��d$}�ek�.����N�i��O?�ɝDB%�� I(�:X�R�2"�JC�r�($K����
�2#/�0J�$��I�D;�@��$��#��lx��b�ߣRt�Ň�&v<�p���A	��$�\4 ���O���b�(@)*�!�92A�Ѹ'�J�D>�Hr�'IH��'��Ip�/Y!*��E��Oƃ��<ȶC �@=��D\��yr˔;1l`5��D�zH���jS�W7L��&�ņR/>�ZmE#)�M-F��é��9�����S�? ���Q��
/3j80�(�7 rg�i�JX�mV-ǰ>���(�$ً��:O���x�@K؞�Q�aǵR/p ��$��z����Dd~)b����w/v���S����c
�(�b��iH8EDx�	׃H&�����T�9�lyU �4;Sn�b��E�T!�䄑(�� ���L�H��+�l�N��b�/ �' �>���8�pv��~��(�c��*Z�zB�ɜ+~J���Ϩ]�]�Q��(BP6�_�`zZ��R�lCP`\2H�8���I@��%q�$?lO"1K ��d���~h}�1��0��q����7�^��ȓ�$�s��JzX)� -2B���?�AN�Z��H��I֜4�ԑ7'Z�M��L!�Cě�!�d�%/ND�,�$�l��C������թH��b�"~nZ��ҴB6��a�
	+�n�vC�	��`��=%^� ��j�L�@��+��'��xb��U6W�B�`��IM��u1�D\�d0OD���64����*5���r"O�-��/�;l�����!4�)��	�dm���):>@\�a�܄0��IBᏑOb!���u�<�&��?A���z��׬]�����p�=E��4�p�C�\H�I:��N:;�&��s/�x�ph	�K�E�G@]�#�U�'��[D!��=�0�ӗ:=zr�- ;���c�JX������u��6m�p�\��E.k~X��K��^�!��,&I<tXf뚾H��@�d�Iq��H�Ee�D��>���!��Rq�TKc��D�e�*D�<�U�76���ӵ�!.l�`a��tӪ���
LK�S��MKCE�4cBᲖ�l��)Q�Cg�<��Ы-�E #�^�^	�`�g�WN}r$(a6���d��U2QТM�8X@=z���)~4a}��3<��I.���e�Q� ����G;6B�<3ꜰ0&EG	:�i{�Oq�"=�!L�)�?�"�D�.@1C[�t֒��<D��I��J�5�<��Z�G�8T�C�d�4\����w�S��Ms�F	����B�_.Q�Xm���[�<I���-Sr��{ �. ��f�Uy2��p>yA�\�V<��KթH'9bA`D�PN�<iDh�c���#��L0lJ�UN�<A�nX�����*	(�}���J�<yG���'Lx�D�E|�lp@�_E�<�5bz����!b��{�����[�<����m�V)*hj(�S��S�<�Qn��6����'ԦN��Kf��L�<y�Ē�7��r�*�96�飰��l�<�`�ƨ!��I�愜��A�Ġi�<Ap���/�:���J\��xp��l�<�ҦȂ[F����	-[<�ي1̇e�<��f�l͚l8c���j¦?�B�	�nw���#�Y4U�2aCj�i��B�I3&�I$,
�-P���_�`&�C��8c2R��E��x���T!�C��0,-��ȿ4i�ZV�Y0`zC�Aih�@�G��BU���=@C�ɑ*`(�j>>Lr��?��B�I� p���+9�d�x�N�a�B�I��h�;��E<� ��&L��Y�6C�ɷ������( �I�C�	*n͸���e�	^&3C䉁?�b�r�o<!���� 7)לC�	�Yޚy�FK3e�l�h��`��B�I�i8��W�5=���;��B�I�U��Y�v�?A���HԤ��L�\B��`���JgIka4�Ǒ_!X"/$D��� �ϠVbR�gL@%Yܼ���/D��  ��nR5W$V�b��b.Љ��"O���a17U4 �0́�S%�	��"OPi��jY�W�<�d,�?~ZI�Q"O�`�-Ϟ �R��g+�5�@��"Ob4z�,I�U��4
�)Z�3@"OXM�1��X%Z��6� K�l�s�"O��ƒ3>�
���a��I�:��'"Ov$ ��2j���f(s���R�"O��Y�,ʙ�
,1�%�YkX�F"O ��'/̀���CϩR~i�#"O�Yڄ�ޘ\&�\Ygτ' ��sP"O&ܰ�
5Y]\��c"0�&@J*O�S������sV�1�`S�'��񩠄�3�1U���K��XJ�'A��0�*W<@� ���ِ@ 4�
�'ۆ�RO�1`����OH;᎘r
�'BYʴ���V������I,8�ƝS�'�^գr�[�k��Ea��ڢ&@��'�ڙ�D�2<���ϳ~2�!��'����F֟N�,�AY���K�'�R�!B��YD�k�i8~�V�C�'5�y���΂2��ᓢ�Vs1z���'[zDZ*��z49��4l��@P�'چ��g�#+VX�q�[�d����'m
�A�#�~Y�P��,1��`�'W���OA�J|h"��<�x��'͒�R�f 6'Yb��`Ç ���'%��IEOQ������V&��'Ȣ��g �4b8�	�	��}Q<���'8�����'�� J� ��@��X�'#�]s���|��Q�eEm�X=k�'�h̹!a�ڎ�C$�� TT�':���ʃ��,z�i�)i&���'�8��w	�>lܴ�C���̴��'�P\�e-JBg&�h�]:!����
�'�z%�S-S�H����s�ܸ
�'�2�Fn��'�&9�v� .�ab�'-�)S�N�Q�;A��-l�έ��'-´Ҷ�N.@�q`#�ؘ\��\3�'�q+���S�9+��T"?3\���'+n��iNb����8��(C�')�xpi_H�\�h�JP�/a ec�'
,� gV3A{&����(�$�Q�'5���˖8�vDQe�-ml��Y�'�8���"L�``Q�
�����'��2&�Y�2��{B�]�;p��'o���@�6!iQ����*���y	�'���b�# ,M�I0�����I	�'4Zy�AOP*L!z�C��N+9æ��'<�:6�TE u�&��
i�	�':�(g�B! ���R)�]!Ԣ	�'�"I����첢k�,�F���'ў��f�46A�[�&���j
�'A�8*gC�Vݦu
�ψ4#�<z
�',)��	(%)�(���t�9�	�'��XC��O�>	zU�O�X�`S�'$��23H�x��q�����v�����'�xY �#�+�"itO�$�@	��'V�]3�EE���������'���{��& �������"�A:�'�v�9r�
c`�0K����;�' p�AAǌM$��06G�=Z�'����`�pE��b�ŋ�'���	�'$e˓�S�i��%*�iZ���}���� I�F��&v�"�R�P#
�[�"Oj��nC��X�Q-D,u6Mp�"O��V�&���;����"O��R�l�b� ���#h����P"OԚTm�)=�@��bQ������"OP\��&�	]������L�$�D"OV="u��BRx��qC� �����"O ���aֵ���K!�Y�?��Ԛ�"O�@� �ʍRQ��yCAʎ�ĸ�"O�5Xp��_���Q͕�K��ՙ2"O�8��&ڋ��	P���cܤ`��"OJ���gUHD��p��Ы}��X��"O\���])X��-��c�F*a$"O����7
NLm* �_�/�(p1�"O:�!�'vH���l�(V,�4"O,���ۈ	5�pr�˅Mv,��B"O6�K�ʚ20[�l�-ɚG^�l:"O
@1�LD
J��h�U�R�ոd"O�9B��O��KӬ�&8Jص"O�=���L6D�B�"�N5����"Oܘ�@ ��P�N�"F�S"O�l�0N�"��9����I�1��"O$�s�@9jEBT�@�r!^���"OD�r%(T!Cv`u��hs����"O���H�r���P&�V1'�fi�&"O�a�Q��!zZLD��ǈ�A߾��"O|$��K8=�d���۔a���"O�	�#F�h׋�iqL��G"O���piX�R2�I�kÂ>il�0�"O$)Iq���!�/�CGt�JV"O�%#ծM�mBdXc��Qb����"OFk��N�WP� I`�/O�̊�"O��;p'�r�0(ʣ�
 ?@�p�"O��@L�"Q2�[�14��p"O�;3L��(�����:@�y�!"O(x�b��!%��l��0�y�r"O@�5圐i�<���L�;:VFA�P"O"��Sn��`((m	;<h, �"O���af�g�Эj��J�Y"l�"�"O�hT�\10Ą�ɂ��+#"O�l��0W$I�E��P2�"O��t��@�R�3���(��J"O���jLo-������74�,C�"OF(�UGaJX�!Ƣ�C�]r"O��YR�F6�
�i��B(�fd��"OB���cT4(��e9��9æ�w"O�Y.�1%��b"%D�N�Ľv"O���Ǝe�����CM'��H;P"O�i@��Ff��$BɳC�����"ON��ો�V��a2���T�Bh@�"Ot؄��W�yC������"OB�[�d�0 ;�92 �D�g�%��"O�2ri�I��i���oؔ�""O�i
�_��+��@� �|�jW"O
�{&�P1����V��
�0��"O�M	6#�*�N`0��2;�,�!"OtQ�Z/�6����
�Ŗ� �"O&�`1"��.i�gh6�fe) "ON��e�F'U�.�7�¨B��P�6"O������X͊5
C*Řw�40xP"Om9��+�Ui0�_�R�8��s"Of9SV(���-�!� |�"O��*d���P����qm�r��s"O�����4Pz,�r�oΌ��"O� �H���[�^��R�ΎF�!3W"O��Ѧ�;&�
�ٳ�(�����"O�́���P�����b�$�i4"OZd  ���&�9�����F"O��Z5t� ��۵62���"O~���'�uN�� Ê2M0�)�t�'��D��(��h�$ �O�r�=�ȓ;�$	aTd�V�4�PR�6��	��y�Z!�ܬ#R��R��?4"�}�ȓA�ָ-9 a���]�H����aJ4D��u%;\E:��CA]��-c�*O A�T���X�n���n�{���D"O��#6A�JNԥ�$`	�Iѐ��r"O��@���1��(q"�;V'��ا"Oj�:" �>e"͐�A�u
� ��"O�l�r#ʴ<�L1b�<_�	�"Oh	�I:6<f-i㠎�;��u�"O�-�T�Oo�i�f�Y����S"O|ܢ�ˌ5�~��u�ژf�e""O
pA���T�p ���6"O�����K�AA���dR�0g"O�����.���#�N]��r0�W"OFU���&�~�K�B�~Э��"O`T� �B�q �C�CK�"O�T+3)��|�U"M8[��-Y�"ON����.EcDq�
B��d��"O�0儋�R�TÁe�p�ޭS�"O� ;���f�$� ���c���X�"O$H�C��A��U�BM��/N�T�"OJ91$ܤ	��X�ۿD8�x�"O4P9'k�G�������MJN�`"O�IiFg�;D��d�`G�}��"O��@��Ne�%"ǡU
M�*D�Q"O����B����a�����w"O��" = L�Kp/E20��"OVԓ�I�|P�=�)_�Q��"O����Ίd�� TB
:fni�"Oֵ����@�^̸g�@��h"O���CBT�M� �����"O�!�MX-P�fPr�^]�k�"O���D-2rc�V��T��"O��k\/���
�k �5Kd"O��a$��>ܡ���%T��"O�q��b�b�nm�w�[B�4��"ODmQ
������� Q
�I�"Oڬ��@V.`���
T�9�I�@"O��9��\[&@��R�T�D"O^�y�]�+@��A�;Y�0�B"O($�#շqæt���܇��y��"O2aԩ9� 8��BÑ �~���"O���a��Da:�h�n~���D"OxB2��!@������"nl,y�"O� ��n'A|&�BP��P_\�rS"O��>y�bG_>S"��"O*@q"I�l3���#��?I�#"O���R���`��	�m�F��"O��	��̑�nА�핳M5*$�"O����ڦR@m��˕Y n��"O8��`I/M����*��jT@$"O�1�E��d	�
4�J,W�H�+3"Op�P�ˬ�ܘh&��&>�(��"OP�Zq	�Sb;�抣e6&�U"On��g�K�j�BE�P��7��J"O&��螂(�J@/���p���"O� �s���v�F��4�i�<�cD"O�I�$�!0��Q�#G݄}�&�#"OQP#֑��y;�^��:�h"O��[���d}Ԕ��>,$��5"OB):_2L�!��_!:>�0i�]��yr�4͈U����(�l�w�Z?�y��@ld��0拷�쩓VjP�y`����Ҽo��정��$3��	�ȓ"B���R�%"�H���L���ȓ,{r`�3����t`X��_8��ȓ��@cA� �X�w��;�l��ȓdx]p%�C�uH 8�I�b�х� ߆0;AGQ�t�:t҂*R�B����5Z'AV�&d����K7Ji�ȓ˰!�IW��l�Qj7�^Ɇ�b�D�l�!((�֤\
��ȓc��U@�G�t����T�$���m�(!��$C �L��%��(�9�ȓ.�T������`)������ȓ��S�gU9��H�&��[�x�ȓ6̨�cង���Q7-�k}4���POZW�6)F ���F)xp"O���D)BtH��aID�� �q�"O����k�Z	��u)�#j稬82"OR�y�F%S����t� ���"O��p�=c1���ǈ�^����"O޼��-*�� ҡ���\���"OZ���ָU�^�� �ȟ(��͊�"O䰊$j@.K� �ׅ�$�|��"OD�Dm��U��d�#�0�w"O\�`'L��{H�Y�գ�?�Q�"On�Q��؂Y$<�h���;:mA�"Oq�3����}��- �"O~�	@����Lb G�*e~l��3"O���rd�D �{@�P�� P"O*A��OȥoX:�"Q3���C�"O�J�r�X�2�O�����"O$$c��_9>T@��:��4��"O�=��qk������ 8/L�Z"OF��Q�.~�6�!WԌ9(ܼ:a"O&%!����|M"lJD�ۦ$P�T"OjĩE$.A���ظL��|�@"OT|��9MR�b"c��E=L�+�"O�H�񮓯6��H��E;̹B"O�@1�ޚ(��9@,�S'N5��"O���e�9F�ܤS�JX"^�ٻa*O�Y1T	�Kba
���}��y)	�'w�Tѣ�D?8]ڭ�S��<�ޑ��'f"�Ig/њtb-1$E�np\m�
�'&��s ��#w(�f�S�_���	�'d���cԋA��j60T7	C	�'.�C֕B٢������FrB		�'����.�2�r�dK.>���Q�'����6Nͮw�x���S%v��2�'b �����)A��a�NIG�)��'ly�%�ͅs줼S�n�	b�8�'����*)����+�$K	z@��'���H�+�.��8 TI��B6!q�'��@�+<7\��-%A(,E{�'���q�œ?BG����8����'���#��ݵ{�H=+p�X�B���x�'���@�u)���@΃DJ�q�'�j�!C�yG�a[�셞B�ȩ��'���@�ɢL�QcQ\B���S��� �E�$D�yj`�Bc��(xx��{T"OX��a��=3>�)��R!No(��"O@�x��2������MW�@��"O��[�Cѡ}@Uk�$n>T�"O�l@�O��P�����vak "OH��V�c,�c��h��y�"O�CP��c��4�;#���`�"OD���R9"nB��w떈Y|:8�&"O�b�������Z` x�e"O�a2���Y�T�CҨ�!ET��3"O����\����-h1��b�"O�d��	�.�dd�m�
�*p"O�`����tۤ-&�C
�����"O�}���8<pAx ��F�D�6"O440��]3C� GD��3�|�5"O�����DIP��`��d"O��YW��l�a�T�.�xYې"O�����T	�e�3��&\Tlp¥"O4��ꃪn��@�B�F����"O�-�r�W�4������K	1^��z�"O|(�fm��V�6AW�0%4�%"O�R3������!ǰxӈE�c"O������
�z�ՠ�&�F�#"Oj�bs� U�x��o�~��x��"O,�"���>@�$����� ~~e+"O�9�^:(�b�Va3zY��#�"Ob 3eτ�	� a�t�<K$(qQ"O���p K7Z��H�5C��2DT"O��� �E�_R���X6{���X4"OP�+�j]3X*
�`��3��4��"Oh�i]�M���WFP�q�d��"O��B*�)�\�H�l�hH�"O��fhϮ*>,p� <am�5p�"OʱӅ�V'i��J�O�_V�T �"O����2Z|�K � �[�@ �""O2�SƬ�I��`��O�O����7"OfL�UB�%Q�:@1�b@�+����s"O�	*�MVj�q��׋j�޴�@"O�=�e� b��1���_����"O�=��,�%�
�C͂�_��1c"Ot�@`�H���Dk�
�Y""O!12��{����I�y�8��"Or�b�F'uK��qۓh s4��ȓk�����7x���9dN�r
&$�ȓ@)��pm�;���%�г.;~��ȓjhm9�HU�D��Ap�/T��8��ȓr<���ä��F��Y�`e�zهȓ/0��sa�Ia�Qn;ꅇ�&4��(7&M@�	qe�M2*$ҽ��|��}�G��&�z)���O�*��ȓ����9-�)�RŖ=E�r�ȓi�J����o�й�A� �g$��ȓ<$��b��3?`ģ���2#EDՄȓN�B�[��+"��}SU�׬��ȓCe�[G�:]]6�9�_�c\|����BcO�>etT9j���!UVh��#3UA�#�63^<4�H��ȓj��<��@7/8��i��Zk�����a����1LB�m�#$��-f�`������2���`k�9����Ĥ��z"���.а*u���AB������W�L�z�MĆ\ڂ))�-P<Gt��ȓ�����Ȝ�7D�u���� ��@rL3�O	�)�,����Z�D����S�? �4�El^%��1�5�K�
���e"Ojt�7A�3W�<��!�;z�Ѳ"OJ��'B\��i11*�2K��"&"O6�k(^��lC�iY�wH��y��E�D���K�V�"�1D�·�y2N_�B�L(�í[G�,ȓ�'�yR�0�p���DU.	|d&A���yR���P�z�z&�S"}�r�b堆�y".�v��Hۧ�ֺa�]sD@G]�<�al2�ꈚ���.)�]ҥ�}�<�h̰/A��/��p׊��W��a�<���U��h�G�	�t���5��t�<�j�=~J\,�A�Ğ�j4�Wlp�<�d瞽"��#R�v`���p�<�Uf�.>0�B�6^܉�NS�<)`L���z`�Γ[(L�+�Q�<a��	��lɷ%�n0���`NO�<y3�M�i��h塌����eEO�<!�Ay��8���?M�;a!s�<!S!eȆ3���2u�EH�<q#�'LCT�PSU�|�l9��N@�<�VO��ZTȄc�~8Șb��u�<�E�j�����z��0t��t�<᳉S�W��D���]�B=���m�<PB�']Vii�eƉ)�d��c�<Q%1Z����^�t�����A	E�<�w� )�x�	���`*�H�d��e�<�&S2��8ɐkK��4hRi^�<��@��N�t�Cϖ�f4(A�$S�<yeK�Jn6e�o��a�N5��*�t�<�sg�=c�`�'��c�=a�o�<�%�3y�*-�Dτ�6����#��l�<��-C�>Q�JX�n��]�3 �s�<�ӌ�#�P� ��I�tlj�kHU�<a�Ӽp�ذ+��@�1�萫Ӂ�M�<A���O���DD^�v���e�o�<��i%~.�`�ǋ�4{bPk���g�<�v�G8ze:�b���h_^�(�_I�<I���8Z!�ѤX�`+n8xdF�<�P�Q��2����M/��1��-VI�<�nƌ&����큈G� @�Z}�<�7���`9��ˡfQ0+ʰS%B�{�<�1o�D�U�s���P9�9{�k�v�<A�I��8hZh�$��X̮���)WX�<1RK��l���Z2�K�̈���Q�<�⋕{����U��c�:9���U�<y҄�=th�!j�fW��F�`4D�O�<�W�P$b$ք^����aV�^I�<�7�G�*�<0a)�)pnY�BO�D�<��I�6j8t��3J�2�����@�<�3�Bj�zͲ����*M��Dh�~�<)6�" �V��"-ON�!�À|�<YSN�>�V��	ؐ`5>�q�kSz�<��(X�Kyl��ve�"�F�+��vx���'LD+1B���a2U��i��d%O���u�~R�"�ܞ����"O ���A[>��X`�DK�{�La��"O�A7C��}�D���D	U�� ��"Ol��� o|����B�R�|T@�"OВ���3ZJ�h���7x�x��"O&��m��c&Nb�� �"O� 8��� (j�|Ç䒽pC�d(�"O�P)�l\��J��7ߠf���8S"O�,���!���a��3 �LI�"O� ��*w`з,�Ā:�D}�
���"O����Nɼl�������E��S0"O��b OԿ4���a��܆&��9��"O��p� �w[�`��fҼS��=��"O����I��$	h%�랖D~���%"O|�X� ΰZ�� �C
jN؂7"O�9�
S=k����d*�Ch�|P�"On�y���3B�P�Hu��}(��"O~���)œx�.q[�	E�m�"OY8��	,J��PfߋX�e��"O�u��H�(��a�ܳ��("O(�!�&�6�3$�0i�؀��"O����$\���t���;�"O8�ã�+|�L�*���g�2�
�"O@a�vHc|�dC3��|�h�S "O���6![�g삡�$�&���"O���'D_� �WD0A!��z�"OD8�1�Q�!,�TB�$<�L��"O,��^�K��L8�&O�B�09"O~i0D�"�ZX�ͬ%��$�w"Oj�R�k_�
]y��X�U��0�"O��R��9x�t���mI!I���U"ONA[%iEo��t����F�0e�t"O��4��uD��	8*�Ќ+�"O8xp�G�^��uږ�\#�*�J�"O�<kQ�ǒ&����A.^����"O��@4�Z41F��p@R P ]� "O�0J�$��f*T�ϓ.Cab�S"Oz�P��� wΪ��mΝ����"O����ʰ;2�ē��I�߼�1�"O
0��D�5��������c0`��"O���g�dNԴ	0��F'D|�"O��C'��su"�B�Ȑ>E�}���D(LO�YQ#@�	R`���OL�~��pI2"O����\3$I�yXh�f"O>�86��L��xKfΔ�_Z ��"O��p��||<���9iC~�S�"O4��I��"$��l�>O*��� "O21�P(8�rt�LҰ5z�A"O��A"�Y�T��@ ��-qX@Qw"O����홻%�Α)�(�̄$#"O�	� � �BZ�g��d%
�"O�Y�
�8b`XR�o����!��"Oꉺ���BC:IN���uH��|�!�$���`u����={B�h:���!��ğ��q�.T".�=��'_vz�y��'�1O��p�� /�U�5�?pQ���"O,�**��l# �85�I�(J�k'"O�d�D�m7p�����O=D�)g"ODLi��ЗA��UJ�8_�ԡ �"O􈈆!�@�V�����y��"O�LS��J]b���f�lp��I�"O�Jq	�.i�r�`��n=�I矰�	çrwR�Z�!�i[���G"Ht�ȓ]T���\�"�T%#�E]�^h��*�~%��H1DD�q�Ӌ���ȓ?���TJ(
�.�Ag��+�ʐ�ȓI&���C+|���x�$ɉ�p��ȓC@`R��}�"�
 �̯J`��ȓIW��7�LY-��{SL�@�0��NNl�j��2G��	q!I �t��Wԍ���?ٴ4`�%��!��ȓt��k�cUv���OU0�z���}oj�"�拍��S��Lc/Ć�S�? l��5�\?�!J`HYgܽ�"O>% �b|���  IN��"O.���п7҄�SL[8 />�q&"Ox%A�#κ'e�]��N.X&�m�"O0GD�.�t}hւ,X�+�"O< �s�W)�جw��k`b��'"Ou2�o[�\�D)�gU
\U�� "O�Hx�ϋ!V�N�B2G^�{��v"O� R�c��{��P��&U4��"OƝ٠"U,I@ �PB1n+���s"O�����	/6�;�B	_"|��"O��U��,�	إ��9�T�0"O`�S �Bs8���DJA(�"O�e���B�m��|��@�y�n��w"O:�����
.����!J�ē5"O�TA���$�|�*BׄAН�"O��ub�R0�};�@C'�b��"Ov`"�,C�h���@���Je��T"O�<If���%0$X,W�`�)�"O�y{�/�Nr��A<y��t��"OTH���=�l�ʦ8���z`"O�����%�Z� >9ҒU�g"O>�Z�Ǝ�W��@���:�B�2B"O�q�5�[
~�l�o��a�i�"O�P�ii�J��-�t��I��"O2�b��]t��X���M�W"O�6�P�k���z� � h�~���"O�d(	??aDٳ�P>Y�>a��"O��X���(�lh��،s����"O&�vI`; ���"ĥy>�m�"O\����[��<��!ޮN/0��%"Ot�4�/}t�z�� W�HI�4"Ota�s@͔=R�	Ǭ˨#�$�j�"O:�q�횋P�E�ԋO�S5V���"O�t�����Q8�%`*O b���"O��kM��0���2S��0la�|��"O�9J	޷T�
���ac�i��"O
��e��G�ةq���2va\T�"O�Lx�N%t�D0#�֚"�(�"O�,�C�0����b�,I���"O<�āU�A'0�:Adçy�`��p"O2�aɂ�^��[f۷NYf�i�"OȰ��$O�<ĔAS���-��u�g"O�,�B�)�2R#�.��hiw"O�������)�7�U5-��Å\�T�IK�S�O��\@� dB��qgX@+.%`�'���`��оRi�8Х,�=�2uK�'6�=b Nؒh�E��O@��;�'C��bBN�T����\i�'����,�Z����#M��6ܢ�'5����A�.7ɰycE h�|8�'�RAGӏނ	�2�ŚtQ��Z/O@��)�)ʧ�B���ΧYT�\���]1�\��`�L�¢
*(�)��#!�\����Ar&K>C�f0Ɂ��8a��ȓ2�(9w�D3mvI�]�UxL��ȓ7��X�e�.����3O�J�d��ȓ 醨��))}�� b�#4�ȓ|d
2�ġ:L\d�t#�$t��a�����1Vz�@ �I�g;�|�� ���j����Z�.�#���)���0��I�5C�T�S���i�l���.�X@�򇉅n�N��e��%je"T��\����:�� ��"byj%��S�? �y0��]�N���Y��3jq����"O��p��p��pJTA)k@����"Oa�	[�L����t�� \949`'"O%�C21Ը�Ue�8s���"O昀� �i�`h���!H
�"O��i6!)ekL�F�Ն)��
�"O$}�512��C�X�x�"O0	g�<~n���`������'o^��Rl	�<�݈��Z�ER$�'Ђ�Z2�� %��T���U';Ҭ|�
�'�t�ä���P@^�9�
��g�2�:�'�6�P��W������oM�S���'5j\: '�6[\��q@�$��Q
�'8��*EC�#��ps�,��t�U0
�'d�esv#�R*
�1/��a����	�'� 0�	�<Q��a�0h:	{
�'Gb��U����|%i�	ۦg�e�	�'X��+X�jy)��C�k���G��`�<�q&��|�d��̄/ar��w�`�<��0��@��,EK�q��I�Y�<&B��6EtM:3��#u�X}�֭�O�<ɗ��8V��BL��}*ZQ �g�<I4˕�>�`� V�V9�eA�^�<�e-td�(�7��^R~$��+b�<!�9�J���R/k����/�u�<q�gȣg��Z��7��{�TG�<!$M� )J��7�LZ8�q�Jh�<Y��m���郞��u��m�< dY
.���՛v��"���`�<���T�k��xVd�C=h�z���[�<Q5�
6-~B�&����dB5�DP�<	�L���p���_@��r'&
u�<Y"O��'�p��ǖ@�䙥��i�<q���VQ��C!7�v�Y�UJ�<��U�j��J���b�(؋#@I�<���P]�ڔ*��ܲEQh\e�Nx��'?,�(A0�P����L�t��	�'�:(!�*1�^]���L�3 ^H*�'d��j�%�	-�d��p �~���'� ����\�ntc��_6�L�
�'�@�!�d��	�4�i'�F8.�F���'t��%�A!~�J�f*�= >��	�'{���,Y�?�P��2m����t�	���'q�}��-U�{�Z� �jQ��:	�'e<	����%>��������'���R�ѺH�r٣R���߂���'$�+���"K���pO�#un`��'��쁣��
K�2Q����!V����'p�y��B�3d�-��%�* "�xi�'�%Y'h�(@���kR����бr����F&L���qf˚M@l�b	�I�!�d�>w/.�㔦J�tD6�"�d�L�!�@e�Y���8�1��
�g�!�d�Q �%������g�&_[!�$[�9t���_8i�V	��b� 1!�qt�4:TW�U}^�
�AG,# !�<, Q%@�@l�����F�]k!�A!��	�a��wX�m$ �`!�d�SH��3�o�)BFpcc�݌Q!�d0g�QX��@�E�Y��o�?H�!�$�#"�2�ISbB�u�,8�h�%T�!�W�A/�=��مg�j��:&�!�i�jYZ�D�� ����B5�!��Օwa6��2�C�V�z䇔�5�!�� �᳗b��5ߒ0!��	�HQb�"O�-�C��;J^Y��	�6uԴ��|��'`az2݋v,�(j`L#S)p��"`��yr�Q�:���H���`�1�F���ybg�L��Q`��]��0�@�yB�."q�[��A-���k�i��y�ᗃz�%D��y��Q�:�y�ʂ8621��J�=qo�)������OT"~b2���K���"e�,v7LP8RC�K���0=�di�:Pڈ	�"פO�HX�g�G�<q���^4�� ��"���P�B�<�!I�P�8���5x����z�<����r�`�u�H�H�@Tq�<�M˕R1�9C�냒QK��v�R�<q�,:(l�h� �3��0p��IJ��?�	�'6��ɰ��B 56\�^�VA�u�ȓ��h)�EX�k���k��H:l����Q��ab&g�HR<�9@@�l{PU��z�P��J�W�8��c�<@�z���J%`������(����|���ȓA2ĉQ�>&�pR��2�:9��a̓2�B��n��^`�Y�Bl��s���G"�S

��4�֛�Nu��!0ԨC��4A��bG<k?}S��Ò;��C�Ʉ����hU�`�1�6�O��JB��<U���Zf#��)JDK E��
�FB�I�zx�} ��(5v�hn	�c�0B�ɸP�$i���@4A@�j3�\W�ȣ?q��)Zݶ5`��� xr��v&�"�ў\��	�h��@��"��e��Y��H�C�I �ιc�E�K&�� �K7 TLC�I/�␙EH 7L��U�E,N91 C�I8g�ʀ�+n8�%JᏜ�C��2A����w+��G<��iwꎲL$C�I <>�� ��ɿ]R��gE�����d*�)wHh #(��#�8}�"���4B��H !&�����4#�@'��F{���G��U�
e�DBG�������yr��L%��j�W�y�t`���ybAA�.���9C,6�x���OX7�y"�@0\$4������&FB�Q��y�&@j������JG�$B��S��yRf]�l��j��F�@# 9䎏��y�)F-(E�Wh�9d�RC˝0�y2��m`�i��s��1�@ŜpI!����Х2��P�V�����I1!�Ğ0L���A��޼>��qR��#00!��&:b�Kdș�l�8,r�&ײ*!���]U�u���� 
u2L���; q!򤟦j�F)�4k	�+c��g#I�:�!��P�pi�a!�*U^�ab�*�!�DǑP��(qb��o:������~x!�$ԭA�R�z���@1��ի�rh!�D
�\�D�!��*�Ä�
]!�d��aͨ9�����F�I�Ĥ�(p!�d�=�vթ��d' ���eD!�D��=���#���rg�}�g�!�$�'s�ࠃ-H8v�%���!�
*&�4��k��a�@�;!�$#p��0hС,w\���b�5�!�$؈��D[R)��|S��^!�D�^FҥJ�Ê*"T��.� .�!�$X�t�L���iǷR"dU��ݖ{!��DRm �h��jb�\R�� t�!�� F��eG�]��+r�P�BߺQ1�|r�)��;9C|eb����}Ė1B�N�=Pq�B䉡;L~�Kw�Ʌ$����&U�b�rC䉍>�4ɑ�b�h�A�D�h8>C�.6ta@�8W(��2.TD�JB䉳OW0a��O۩b�I��b��H}�C䉬,�%���_ݞ��Ev�C�	�
�n��%#%W��sD����B�	�>�~ɓT���,����H*B�	;��4��1QɢȰaKD�2�bC�	�@|d8b���M�dI� ��B�I���Ű��@�i�((�%!��_HC��> ��`c`�v�(|��e�?@�dC�Ɉ>2|�A���-W�8S��G,Z C�	�1W�0$퍫]]D�d�<;hC�I�_��8UK'Z9\!�w쑝Q��B䉒,M:����O�Y-D�d�B��� ɝ���E(�p�!�"O ܓ2��,Nɮ�	�f���Ca"O������6�L�#��o�ʵ�T"O�:� L�s���9Ab��v�"O`���e(Ǣ ���Y�#%���"O*�����p<x Y���!��`"O��CM�R�.mbBBW~826"O�Up�(��
1 ų�(zYj�٧"O��!��q������qQ��'"O�#��J(lb�j�)?=x@"Oj��GhO����J�wN�Y�"O�d ���+��ݪ���vM��h3"O�%hf���5�6D��M_�>���Kf"O�YKV�-4�Z|a@ύ(%���`#"O�Z�Æ5�pq �����L��y�N�&n��hs�Y�5@00���!�yR%o�U����.��h�Ȕ��yb F���P�X/Q�*�RC���yR�O�ѣߵ7m���n	�?��ȓj�l�۶�?z��}k&ÒGP��ȓ�|��$��5V�I��N�P-�܅ȓ7�*��(�i��튑˓3+¸��ȓsن8��׆G����E΃-�<5�ȓ�|�)�#�R�"!д�]�f�4��ȓ4��3�-�B�}1�ȜHVDH���t���A],�$=c�ѠS�Ņȓ#��Y���I�NRTc����fQN-�ȓ^�b�	�lQ%<�"��p��E�d�ȓE ��
��XP'V�q2� 9x5�����l_&=a�t�ӱn�0ͅȓn{����C��$C�
!���ȓ�T{�瑒2�l��.60\�ȓjt|�gP5
�����pS�p�ȓ)��P����]3�@nRY�ȓ��@���;J�0;#��/hB��ȓ4ƜeK����/�4��Ƣڭf}!�d�20:�k�F�[����E��/!�B�kq"5*����(�@yZ�KM�!򄈱�$�JP�ݯhu�al�	!�d�9mԖ;oO��eHG*	16�!���.-�m�L�$& ��)_�*�!���=,qn�����{|��G�ڟi!�$ܫ,u8�:b�Ѿ���P"�,-!�ǌ�
I�7��<|�4��Вtm!�,:�*qm٧/�|��ʞc!�ɇ;�ҕ+"� B�8Hҩ�<a!��(V�BŨS��X��C��!�� �Ũ�kɚ+b���6�Ӡ8M<MYW"O@-�Eh��GKv9�rG�2נ���"O��i�A�~H�po�����U"O�	���U�� [�+��<��#"OJ���B�x���j�
v�,a3"O�@�D@؎h��p��RchP�@�"O��w�Eb�xDk�K��;^raH�"O9�S��TՖus�HB�~'�u;s"O��kpH�(<8�ၰ�]�I!�I�&"O8-�嬅d_&I"�e��8���Q"O�,[%	� �!�V���H�x�"ON�c�	�vt�aI�0F�p�4"Or�#v�ӸVa�h��4-��P"O��ÀFO7j�qJa��C"`��6"O�\��I�5�~�� H#C�d �"OD5)�(C#a�J�Z�'��{IV1a"O(Y�Ƣ�5b"�e(� `���"OZ�SKX�Z�L�a��Wۖ"O��Վ��!.�"v��=~��Y#"O���G���X*w�3n7\��T"O��B���72h�]��)��J��k"O��ӲSt�&	��(
�cb"O �Y����L�"I�3�^�S�d�QQ"OBM�Ph���)r�ֳ%-|�P$"O���Q��r0Ec��� �|@"O��p�o�!F��Q��["d��"O��sda��%5~�`U,iV��z�"O:	�Ɗ�8�dI�#f����("O
�	���PW
�2a�2��$"OH�J��
3����hI7O����"O�m��LtP�Q�Ι�Ol,�&"O*@� *��@��y��5�"O&�#���u��Y��?�:��"OސZ�I�8=�ԐR1S�c��I�"OJ-r�䇓HV��S�(����[�"OL9�J	�<���sG�$�0x�"OV�@�d��4p�#���hն��D"OPq֬B�G
��T��I-�	Y�"OF�"� �5r�b���fܬӷ"OĴ+$F�f�*B�T�M��z�"OzyX�遛b��+u�����"O�T{�O� ����G1Wt0�"OzH(`�'xl)��_�n>��#"Od��!�3�0�� g��u*��[S"OhI"� #D�p91���h�1ZW"On���V�r�d��hȝ(�vT�"O�]�4��X�,���fٝ~�Dܘ�"O��y��ٿ#.t|ʧˊ;*T:�:"OL�C��,�LT�mְgO��"O��4d���M��,Ǻ2O\Y��"O����W ,D��
C�s���+�"O� ��,DE\d���JT����"O���dE� p ��V��3r5��'U����H�\"8�W焊G.�"�'��;զ� qu.��Z�j�6a��']�E�#�I�h�<qc�� ?\M��'�v�wr��[�a�-B��e��'�V�)�咇�L�iT8<*�Ը�'$f�A򨃤y׬EA��1-��L��'H*�k�j�2Cl8�ʐl��+����'����P N!�00�*Y�[	�'!��8��
/`��2�� :M���'匕�. ����-"R.��"O¨r�'8b@�y��Ǒ
o)�e"O�  �8���a��m�fm��&Er���"O����e�z���8>jZR"O�P��k��t��cf׉G�x��"O$ �g,E5/N���E� ax�"O�Ay"�B�gߞ�sd��RE�@A"O����J��<�h�JtC0JC�Hk "O�T�`E�S�4�b��S>H3a"O�}�� T�D��騐����M���"D��C�`2K������`���3D��ƏZ��H���G�����*3D��4AŏJ�"P�H��K
�Qx4�2D�����/�
Q������B��/D�|����P��e�Z-@g��h �/D��e.ڵh��LcF�� G�4i�f�-D�(y�OZ8<�zq�U#�$��1D���� 12�\�k�`Q(���e,D�$���8z���a�S
����(D���l�|3fK��l[�Hj��!D�����R^¶���%> �����#D���qkA�ل�C�(M1�$����7D�@�#�8q��,
7��:M�����/9D� �5���]���pǆah��9�j7D������%"�̹7�Q]xHqAIb�<�C��4KO����	ژh��嘥�IX�<�dK��d,��tǜQT�MТ�K�<��"Q�l��8fbN�{ɂ��cŖI�<Ag��������ܾ!O�aA1dC�<��fJ9����*��I� !@�A�<���3�xx���]��]� ��t�<��KM�=n	(��X4�셁D��m�<���A?p���8�������`�FA�<��)N�V�nY( ��;H�`Q	�A|�<��סFDv��@!�Y�||q�)t�<���#$WH�PԎZ7w"�9�t��m�<�1d��[z��33��3 ��1��Z_�<i"�Ȗx�bݢ�hX�'>� ��^�<	4N�n.���[�0�3��Z�<y�[58�p0��_�:��SG�Z�<釉*k��ɓH��8\AYcG�X�<1�@~,ze{�Q�Dw �j5�X�<���ԪNS�0� ��&,��i*p�RQ�<���9Ąl��`	";2���b�<���-�*ɂ��8�(��Da�<���V:v�N"���\���`�r�<Q��U�=@!�R/�G1T<��cIo�<�SfX1_�t��$�!��aE-Hl�<yA��2"�h]�Sh���ܙз�A�<A($E�JT�6���9>�Ҩ�t�<9�!�0Ĭ���}%�蔌Ae�<p$�(taPo�WR�YHԯ�c�<q�j��?]d�!@��8�#��Ut�<QuCM/xn�:����B׸ZrBنȓ4A�¯T�$E��Gɝ���ц�=�����m����F�%*��݇�i��A��HE����b�j}��S�������HT�֖�<�ȓ�X}ÄK�.��V�ۑ ����ȓa�B���i	�z��ro��\&���ȓ��\@�ΐK��岷�P����ȓ@�~-��%P��Ja�R%�"���J+ � �\�6��cI 3x ń�L����L�#�&� ֹb�&�ȓm���Q(�7y��<�Ңa!2kKG�<!���ް���ܸa�rQ
��<� L�3��\�N�6�0���
@�*���"O�\	��T!'wv=�6�S�-甬��"O���T<B���$I;ֲ��"O�qQ����.�4 �Ï�K�=C"O��S a]�`}�QJ������"O�}�qg��H��t�#m^5k�F�Q"Oh�86C+%B��*BϳYE<0��"O`hHa�F+M��G��� >rX"O��y�,rI�.�'6,�B�"OPu��G&��{�C����"O�8R��< ���C /��&�T�`""O��JtL�QJ���sC�i�B��"O���F!DV��1)�!A3i��
�"O\�`5䔉S��d�b��A�t�Z"O`D�s�  �<�#Qg*��"O�}���C�OϞ���AF
\T�aP�"O�:iƲi��˳.[�L��\Z�"O,����
U_�di D,�άZ0"O41{7��=h��\�v��+M�����"O����'ބX*:l�R@7nLMB�"O���P�#"�pCD.O�@�az�"Ok�*�T ���,�(`� �"O�0S�쀑*���l�)!��3F"O@}:�����(�j�"�X��"OZ�{n
'?�D��3�:���z"On��T�X�M��<�2�H*�ZA� "O\T(&��OA��îP�sr��8""O��	P�Ln"J\���> ~�L�!"O��j�WfT4 �/�Cw���"O��	h�d�d��\q@��"Ov�{�l��б��o´e"O���)X�G,d��&�ΟCC�i	�"O� :RO�@_,q�Ǌ)d#*�Ї"Ojh��Ę��M�G�;��ӕ"O��r��l6��@O,�� �"O
LP��e�<D@��O�I:6�"O45Ѕ,g�	�1@\! ��� "O�@yU&
=�H�6	C%-�ŉ�"O�P�M�8 (�k��L�G����yB 	�{��k&n�>i�ⳇ���yL:Q�V�X�M)`�@����8�y��\+%�\���]A�q9Gj΍�y�/���>4`#.�V�����n�'�y�aĘx�����B�K^b}���y�MG<l��ٺ����7 ���ì�yB.S�"`~m�2�A�'^h(B��y�c�Jp �V�ܣ@�)�w`Q�y�˓X�|�`*i囶D\�y2+����`kC�HfB(�	?�y�cͷSF���$B�\�������y"hZs��86G�4Qh�$(6��y���2%1ܵYV��Q��p���y�D�PY��1q�F:r0���ǋ ��yr��pv�`�G�ΘcH�j���y�n�+����_�	�V�CF�Ȱ�y��4y\!��/�t 􀸶�ِ�y��V!+,���M(�j�UHO��yR�2�ޙ����M��0(O��yr�ɥn0�2 �ģ%6 �CJ�y�I��P�yO��V�@�P��y�ؖ6�je����V�V�IQ��?�yr�S%{�x���Fz̈��C��8�y"F'F<�d��	ۛx��+�Ɛ��yBoW��ָj ��s��Њ��[��y
� �9A���lm(�"R�75�V"O���b�
\�e!���/2���"O P�2��3������y0 ��D"O�J��U>/N���2,T��c"OB0"|P�8�I�$�����"O.�#%L9y쑢�a�x�� p�"O"u�"	�W��qb�5f���""O �Y)P</�\���}`U�B"OT�p$Ӯ$T���Hp]�I�7"OB�2U(�/3	t�1g(��L�j"OĄp�GN%���7�˟i�(�"O�dQ�\�D�P$8���&DX�0"ON`���ȈR�l%���q��� "Oੁ���%'���jg-��z~�s"O�{Ť�.+bR���KN	�\�
�"O���`�ܠ���{Ɗ��z�|�;g"O��C��;a���ĩT��8�"O��ZNV�IE�u�%�{{4�@"O����!��K���7@Y�0��"Ot��gM���9cK�J����"Or�#��V$��8;q�V�}��0�"O��&�Ӫ}5��@C����"O�qɢ+��f��t��*x�Q�"O:ɚ��W*o&�!8!�Nr^� "O&��1���&�����4�>��"Ot�A���BA"�3�6A�P�"O�嫓A�[�������s�T�a!"O�$v`P�Fm�`.������"ONi��j˧y�Vŉ0(�Q��p�"OҔ�1?hd��'H�&v�>��"Oր�F��Z�z�S�蝰0���C�"O�)���eu��*��|�bT"O^��1�[>Z�X���*P���Ec`"O�`���JL�� 8n��L a"O�<�F���F���j�3�(�!"O���AG^�Wc�ˡIǊ6�h	�2"O&AP��
.mP�9 k^�t�5��"O�%�����[;~490����z-�g"O��cqA�p$�8'`�=,����P"O��`�T�=~~�#�nWC�DP�"Ox"�Ƴ&�RkI� ��U�7"O|H��	�	:�t�8SJ<~|yb�"O�p��4,Y(,@�	���is�"O^��6�I-�b��k�}��	� "ObyQ-S2�$M�$
S,���0"OD����u�Р 	� Y����"O�@Q�NݮQ�ҡ��D�B��<�"O$��ڸ|}�Y	Ą�	c�p
�"Ovc�Z�l~�	w�E�Z��"O��fa׺n\��P� 
4O�a��"Ob!K�����\4�y$y��"O>��W�(6P-0�ȊA#x�f"O��z5O��[�����Q�D+S"O��b��w�y1�/� �@���"OH� э~��Y�Go�?^@���"O�!Aō�O↼��]�r��"O"{��&�`���];(7�՘�"O�A�@��s�j� �_A�yj�"O���򥗦#��Q�DH�[2�]+�"OΨ`A��!%��1BÒ�*x��5"O�!���#J�	�C�
����"OV)FL�0��8CU���V^�:�"O8�Yp-߰� ���r��P�"O�-�T�:���m��b����5"O� �HqQ(�9k0�qZ��	:�i�"O0���MW�t>�JCM�c��MXV"O�T�b��(7>�k1�,	�h���"Oҵ��ӅFO�(
�㕋\�} "OjD�r���h7��եL�"�@u�a"O"i�'(�6ڪ��n[3qў���"OV}sv��;Nn�ڱ��:�0�{ "O�,�iب%\�x �g�?,���"OD��iG�$`kw��W�PH�E"O�9�B�^�&!A�A�n�Ka"O�� �@C�$���o�RO��"O�i����0Ce����hs�h�+2"O2��(R�~�Aᐭ�7ۜ`h�"O�A�� �Q��{b���(��"OT:�ё'���b�k�;y�0��"OP	D�Gˎ�h7J��pLu��"Oz��fI�B�L����Q �}��"O�I���c�� �bIV�:�Y�"O>\[Q��`�~1�*G�V��tڤ"O���҉DN��3�*K`aZ	��"O4ub��ǡH&�E�C�ܿ(�
y�"O.��5/ ,:��S�³T�|�zU"O�ɲ �T�]��K3Q��"O,� ���BG�:UdM��㛝M�!��Q�e�)��2<r����!����,bqgI�V"�9�UA@�)�!�@�z�����."�<�QV�\�fF!�"sr0	WE�e��A���&,!򤜎T�,$k��#LlZM�$D�h!�DTi�ɻҨ-u0t@�c	�o!�d���F%�G�!~�(p-�u�!�:��I㋚�$��ݘ
�!��A6x4,�td��tm����2U�!�DK(\1���1�����	J�!�ė*U 	��ᕗ^Ķ8���e�!�D�&�2- '�C�0f%��i��=�!�$��UL!Pc�{�|��)���PyR(�2hX�Ls���oVZt[b��y�K�-Ҥ8���� ^����� ��yҌ�/KW��Ӂ�#Y1Q�R���yBۭ�jԙ1#���^yyb����y�o�(x�F�TjW0��bsB�y	�=P���&��7b�R�U>�y�BϏ3�>Գ��.�@�����3�y��G�^�����J�z1�ᐅ�y�N0
0ir�Q�t�0�
�����y¥A-G_�e�Ǔ�@jU"����yR���Mn]�蕊����m�y�	�n�nDj��T�xϪt�&����y�D,K n0��_��iㅅ���C�ɳ;6+o]J"����=М��'����,��;Q(pk0���a<�-��'~�y���[= ( R�l�V9�
�'V�=J�a���5c�
QǬ8��'��i���0�����J�n{�'�:��@4I�5�ț1�3
�'�̜ia ʔa�j�3%A>�L83	�'�� �/3����`K?Nꈫ�'�j�b�ǚ�a"� ���=X���
�'X��j�>��P)�$��|h����'� �çh(}�|���ʿ��9�'��X�Gc�"<� �@Ջ,%@��6�\,0��
v{R�{WFMx�t���A�S.Ze������
9Tԅ�S�? ��� P03�V�Y�ʥ~ȢD"O�]Y�>Cf�="ֆ�,��9q"O�U�d�'4Z����W��aI�"O~�fiH�A�����?4V$�aG"O|qiT��~l�Y�D��)@v�&"O�(�F�2*��lY���
GL
��*O�Е��h�\�2!�����
�' t�Ϙ�Bb�R�G���{�'�F5���TG+���Wn�D��EH�'@h�ȝ2�}�PKM�oԎu��'�㍐�j���V���a�L@�'t��S���0�^/X�ੇ�=�z܉A��_�� 9�)̓\8���ȓe�ĳ��ݑl�<J7�&k}� ��H��} Ǭ�?+�.4HS��1$���JO�(ɥE�a���a! �B�)��{�kƎ��@��F(��v� �ȓ:7I�D)?Ρ�lV�3���N���9�+� +�6\ G�
ݜ���7}���O	�AA,�Ud!��@$��H��|�ׯ�*���`�ް�B�É�h-@�={��ȓz�� ��2N��ȓ4�K�7,�i�ȓ'>�X��&�.��P�7�(I�ȓ/�,�:6ףg���#w,ӈD��H��#;�8�V�ɲA�sá�WFE�ȓ$���FB��>~l�ȓ%�RE�wk��t����@&ي4 F�ȓ#\ �#/T�� ��ʚ�=�޸��M��Sv�- #���Eك&�0��ȓ2�b����]�Hf@�k�ޣ:'t-��TT��2���@�"mN�ϪلȓdN��'e�6)D��B`��n�<�ȓV�Py2�@%њ��Z�&X�ȓV���H䀅'��⡦Bv�&��ȓ@&��e�
�E��D�ԅ�i�b̈́ȓ���[��U�vפy+D��a��M��wܱ����	x�����	�lhD-�ȓ6��zRh�i&P�
)���ȓ����ȉ�>�d�'AZ�!��l�ȓq������7�PAx�aF �q�ȓo���qM�4i`�mȥU�VT�ȓs�FH�ŬC�[��҃�|�p��PU�U����%�ԉ�K�(�ȓ{EN��Bo�%����b�ԅ<�@�ȓ?��p��/�aB
09!� �:����z^e���pNl�(G�P�V��ȓq�0 #Տע4�����]�@���$����
�$�3�mQ�6�����7,.�P gC�:� � �f	�Wo���:Z�x;�� "
�@1@��ދJ��I��t��a%�{�8 `�/e���ȓK��1����>�\ccL�S����,�Ry����9j\�����[X�L��x����#��<1ؔ�#B�ftZy��g6��glD�&�����iiL��ȓL��-��I$;�2��ӧ�1H�8<�ȓ8��,�&m]9Y��{7鋖Tr�<�ȓ�|#��=R~�!��̝'��)��&x��&kϛ�n	i���7��ņ�jb(W�q��_`���ȓD�\�����	KO��	�J��XXY�ȓ|A�X�&
(	r�
DK�+TH��g���c��d���"�)NC�)� H�Cdin���ʇ@ƚa"���"OxM�E&Z���ŠL y�]�"O�|�7��.z�`�`�C���"O�4� \�s��Rn���"O�M���źdp*����>/YĒ"O(L@�o%r*TYc��.K��j"O���w)w� �	��ݕvWʬS�"O��	��6z�Ljn,(3Rp��"O��4�_0}yJ�X�M�]�"Op��ԨV�7�6 ��
���K�"Oxx���ʤ��"C�<d��d�v"O�XS� /;r��t�RHan�b�"O��0�zD@����8b�����"Oha�7ʀr��Q��c�5�Ї"O��3p)�	>��V��	v6�2A"O�y豍ƓEk"���HT�kKr<k"O
��玨~Z2&� K,�%�"O:\ZB��	={$��"&�D� "O̫�Gk1P���n�"1l��'"Ov� Í�}2���  y�^��"O
E�I\�p�|�R�"�2p��"O�0�@D���u�P�z|B�"Od�����#���`�\�
���1"O������%ML���-�f�D�0"O�����\�f`C�e
�Ph}3v"O��a�!�5[�$5�%���d�K"O���E�B�\8:�8�ҮO�!��� �zQT�V�mN�ř��%$�!��6i�5`%ɔ*Lڑ�"��M!�dC-!6h`�2�*���nĊP�!�$Y�5�x���VϜ|㴇��^$!���(<"���`�8
�E��G�T!�H*o�j� Ì^�;��<��Ǖ�b!�7O�h��bV��zi�A�p"!�D��]�p!�H����$�s!�d�#=��;EF��U�8�p��K8	!��?%J�ɷ&��tg���虄n�!򤁯7-��!c�X���>�!�D�hC��#���4 �y/Z�(�!�$�	��k���s�t�I�!򄍧.0�Ei�A�cj�� ��^�!�$�2]��C�MV2HR��s�σ1�!�� �aN"��$GW?�퓐CE��!�dI�H��!��ܣqB�I�#�g�!򤅧\��тӮ0W��%¡��+8�!�dMH&�2'�
�Z2U� L�n~!��֋	xt�b�C�ww��(p�$2w!�dC����PWIi�X� �H�,w!�$I�"�z�x�	 R�X-�al!���Ȥl��#����'[H!�䝬=��q�m72�P�0�O��x-!�$��j3���B�� B��j�<��N��k�ŉ�f�:��.���ȓu�������r1��+~�*�ȓ%[.C��(�D�"� *-�`���th8�J�˘�f:�*��@?9C���A��=+�F�9ڎ���7T�B5��@�R�����Vd$�+pV����dUf0���9�0L����N�ܥ��-�d�t�ӇWv��ۤ@X��2-�� �@@�gI�L�J�I*�LV��ȓ ~J��R7U^�9䞼����a�L1�`�-���r�ݠe�\��
��j �øG���j�"^��Ȇ�S�? �=���� w��\��:��(�"Ol� ��;gj��#Oэ�&�P�"O�"UA���r�C��|���"OPD���� 6)2���U�4�A2�"OD��@/]"<�"��6�ˏ1 �ʴ"OH�yA�L�$��f#��B2 !�"Ol96(}�2���#M�� 
�"OZqɠeF�9��[�,ܪ#�jK�"O��d����h7&^9!U�
�"O��"���ifB������K`�rS"O2�$K^'1����}B^��"O���G&@=����±)b !�"Oz�
r��x<��q��f	l`��"O�bk@�^�na����,*��9�#"O��ؑ��d)�B����t��f"Of��5�Y��`���#*yXa���?D�h�@A�$*�h�3i�.-� K*D�\���5�p'ҝ)�6��'�&D��R��EN=���c�ì�(��!D� �Ѕ�g���BGhB5����!�>D��:gA�OLT�DdV�U���
P�;D� ��	�&gP�C�O<B�\M���9D��Z�/�ѸT;� �<�~�h@�8D�:��ߣP�^�q"��*v�p��G<D� ��IC�s��$("����<���$D��+�AE� t��(ǥh��z�f8D��s���S���s�:Fx�p�#<D����L�S5AH�o��&����9D�<2'$�D��D�����b%D��i2�H^%���G� �ɤ���7D�H3R����V ��L� px]�0�4D�ء�ر�6m�#I�>f9�w�0D�P��G k 0�	F������;D�����y]�ah�1V���$.D���Ȃ�Nd:|��aA>�d[!� D���C�� k�@q�dA�ckhQ$T��r@�Ymmh�9�-Q��8�a�"O�]��m�C�*�@&�E<�0���"O�<�o�&L�B�KS%˹8c,��'�(]"�b�-V��a#�P'iL �����!����-�4>htER�H !�!�D�3/�DC��|G0A26#�1�!��V�^&Д[�͟mMLu �i�){!�G�����z$vx�&�H�!�1 ɡbә�4��!�DK0~9N��A�ث6-��A����!�D��
,+wl�,SPa����9�!���k�"urF�	�L	�d��6*!��XlN�SQ!c�h(i��W!��6庵�d!F�p�^�z��Y,d�!�dS
��[rW<���H�H�+�!�䚥N�z�'$?G|$�A�Q�!�D�?C��C�,Ɲ!�����a��!�d�-#:����-(ʮd��C�:+�!��$An�ȃ [1{�����Q/Za!��W�/B00n m����!nİv�!����=D*�"��7(�����!���z��9yu���������5�!�$FzN�M2q�I.W4%y�ϑ�
L!�ė-'�.)����AD!��	�'�����ԬM"�p�"a��R �3�'�����"v��e�"k�U5����'pԁG:=���AG�ZM$�ϓ<��ag�V��D&y���$	�e'��Q
�qs!�d�?0�����=s�ء�j_�1��'x�\���?	`��� ¤��.�b��tp�f�{�2�Yr"Oڸ�j�((4�
��t��SPbͺ)�B�,�(�9�`$�3��ۗ{2QU�?MH��A��T�E�!���y��2�PR�x�yeÉ�A|Z�:˚� �5�XX��(")�4�HX��G!F��ط�(�l�ttᥓ�A]�)��jb7Ÿ;��@�0�2. }x�!p�<9Dh4`h`����`�sy�ᙇwPh�#'���i\
���(���sM�x��9�!��8yg�`X�kA801�EC��(u� ���
���3#޵Wq
�:�Y>�<�Q���ű@��+��Lkc�UHX����F�0F�ɓ	�6�]%
֣�x�Z�I[���0[@y9E�Vc8�:F��� �n{��!��Q�$�q`P�3|4��Q`D*it�=�Q ����ƅ�m�}��K�+�aҴ�y�X��z5:Ƨ�
���!3���I�"`{T�	1	Q=Lxu r�l��ygA�h�(y��צ�~Ma�.�yb�Fo���*�e�}����BX+�|���kX*AP��W��2$��Z��o���Fy�D_P��\k K�pǾM9ҀS���=GL�'.�7$��U�:A����v2Z��Р�bt���]ݮMr ��a8�	�g��ed���tn�uK�����;�I�Rq�U{�F�����3	�j��0;5G�?�°"�m�:I��ƑP�qҮ<D�4J ��p���I�MK!>�ٳAi\����bg�C֪(��iѾ��-j ������@ߙHY䵰"�=4$Q�4�w�<!�.Ҫ�q�#j׉(���g�֮$�6����P>�h�����-{�r�"�Nҫ|��<YքR-xh y&��z�Z�*���i��L�QC�������M�P|+��c@��'�Q�]�p���4U�"\s���:�p>��	7�8�RM��-:2�ã�b�ũaϐ�H��6	U�o�"X�a��I�qQV0I���6y�W���!�$�1\���C�e�,�p�E�H��<�%�^�SU|��2�M�qU�U��0��O�*��;�Z�����8����ɞ:
8D�ȓ|���Y��Cf�\�RaB:q�,1�7)I��* �)�.0�K��ӡ|���aP�"ʓj� qK��ͥYIH�yb��9b+�!���j�|��.��c���JTMA0m~�����<C�(h��
f� �vN�-ւ!��"\X���6nA:�I����	�=�h��K�<�r�F�v�m3� N���謟FAY�R$���@g�6#���D"Opzt�})�!�0+O8�a��v�|  �'��)��D�0@�P�J'§�V��MXa�c�#d�n�(p���6L^C��-�h=�#$��$�nM��4��l�R��=E�s�5-�֘`n�ٺ���N�.:V����#'	P��ӟ��{� ��wj2�9�M�,9��D.� !=�A��@��.A��c��,A�	
�� l ���(��Aѩǒ8Kh	Ex2�-#�hɑ"����Xgh�����ah��oOЄ�B"OH��&j�>���Q��V�{OF�T��)m�2��͍���S��?tR�5�Y[G�\�VM���Kv�<�R��98�N� �EXr��f�p�<9�*ÈJ��X��A��\1AM�q�<3�ސ[�����QQ�t�E�n�<��k=\��)�i�?�`��RC�o�<IM]���yqh���e�A%�d�<��+7~��W&�*8���Dz�<y�	;m��*%a��e�E��`�v�<i����j��+V�!xvB�P��]l�<��Y$n�: a2M�"X��U�� �D�<1ǌ�'ǘ��T	�=��9�	_A�<A�L��:�F�R��W��ܼ�F�B�<S�ױt!��0r ��4�L��M�{�<�Ģ��d�!�Αei>�C7/JL�<�CG�*F1��޽r�4"� O�<q���6eFua����%˕@�l�<��\5?���WI���T[���T�<9�+��d�0�`ې'��H����<9@�ǈg�(�b�ě�88E  ��m�<ѵ$��t�)�:F��DX#��j�<	3���Nu���7�B0MZ ��De�<	�f��$���� �,.�n��i�D�<� �LsE��L����_$~E�T�"O�(Bp�ߡ}��;uF�"x>��HT"O�,)����r�`[�f;7��@��"OS�%�7임 �ޯ*����"O�ڲ�!H�<٧ٕ(�� !�"O.�f�A`�
A��#�R��Pq"Ol�b��9:�c����SV��"OB���N�3�hX�!\�.F����"O�Yє�P�_r�Y:�[�i� �"O�EZeH�3~� U²�4@G��92"O�@��·W���B��A����"Op�ۢ͑(`�,U��ѓ\���"O4|�r��$?,�1׫�3d����"Od�I2j��c�RA�F�D���U�G"OT$��
k皔 @�PZ�0Y��"OLU��ɉ1�$�YBW.(`ڒ"O2�[G�܁`�H�(�s���e"Onњ���b�CF�ߠ��D�U"O�U�����ؚE�<1����"O�$3�ț����yb�5�mk@"O�P�ԯ�'���!�G��d4�@� "O2,���8�}k�� �"��"O�Rab�,C"���1�
��F"OX��Ī$:>D��d�=gPI��"O|l�w���Lu�����ˉqH��;�"O���M�:5�Z�{� Y8O�ܰR"O������>Yu����τ�s4d��"O��yc�A�[(1*M��f?��T"OԠ��9K����퐮z� "O�<��"]3\�j�P5LK.�IY�"ORLr�Z��Y��k�#1^`���"Oh���"3hȹ�)!p>zź "O,Mkp��.%�V��F9Ctp��"OJ�R� �v�����G�ok��3"Oƅ�.7DQ���Z=�0xg"O ����?10�V�J�L"�["O�t ���[�$���&חV���"O�TYюW2*h6YJL[��"O~���Ht����#*�=	�:��F��'w٪�ڍ�	�Kd�)c	;D��1�HٲJ!�d�=j�����˵ l*p��ԁ24@ѻ��I?��gl�|�'�$!Ă�V�`˅EA]3���'@tB�eV�X_��4�I:W���b2j�E\n5��刡LA����	�`���!�9yYDT�%�խZ���d�*r񺜀D� *Y��ۖ L�.�![��P�4���0�l��*���!��ېI$
���F��f�'�$�G��	<"ђG��3t4�F��)Pu��h�+��nO<�Ò��1�yBh�X�vq�F*��t��1�&�U�x��8�厗�n�t�CG���i6P����L>��n�Mc��i�%�v5D"�(<i��n�|P��B�p�9g���Sa���&��pҘ�`T·�q%���G1�������!,�!��Φ/�axR�ߦ<� �(�mX�z~$])��a� �`�T��h���� �̵!�Orh6Ι	\͜-JT眄wU¬�Ɲ�<C�N8澨9��H��!���s���xAAaKG�]0��IH�~x`݆ȓu�HCu@Ŋ-�b�&�Qq�A:7K�7R@�ಯ֟[k��(�G�f�'��.Gf���EW$B\F5y���KV��.Dn���*݌?�n1�`�S�6���X�����C� =(5QC	��<���(D�`��ƥC�u`tp�Bs�$�F�6*��kC#��w*��ʳ'��w�u�%�]�
�ڡ��-��\�Ɠi�0�#f�\��%���R4cS���'���cDMZ�m;D!�m^]dΜ ���L�`��� ������	4�!�$�T���x��`�
t��(q�dG�Q��!��0LƠXLC1�ĒO�`��iP�l(��u�$=�0
O4]�$"��v��9�J'�%��^�8
�c�N���0=� �PB0��=`��ls ��6��@���'���
�A9��T�sF-����4�Aa!�;{V\[�H�I�<��g��&�h�Rp�7
-$��M�ɃoR\v%[�}����$^m�Ojd�d攈c���6L:f�����'�(9�Ĩ	��`��Mv�6*ҒEJ�b������ � ���ē� ��슰(�@�"^sBh�Ɠ�*y��	��.u���ՐEi�y���R�yԒ0
щ��
�Z��䒠pL��/�I%z3v�zr�z�#�	�Y����<�g+R�X��<AR� ~HiR!��Z�<� 
:>��T ���,��g@J��@�c!�v��d�!(�B\8��^�y��.�>�I�)Cy�~5`��ѻ_y���ȓw�@��"{���×0*k\ ��_��c�"�$h�"��%l��<�ȓR5B�+�)n�+-"n�`�Q�"O��rA�I&��óLs˜u:&"O�ѡ��՗r�`Q豮[�w����"O����D�?C�Z�;6�]<��m�T"O(��q�Uk8�R%�
2����"O�)�'f��lF��&*B�*�,1�d"O2p� �(�X��P���w�1�P"O��%�47�`1C�,B
M
2,��"O�tt�2T����A��q�	
v"O �Y&k�<������&h�Q"O�)3a�)Q6`	aC/�zeb=��"O4%����302�{�,�#zEΉ�q"OdS�l�s$r)c녂G���kG"O�p�����*zpu�j�8st��[ "O�}Y7Q��R��d�Ot֥�W"O�̓���o0~e�`�!P�D���"Or�C�ʁ)M��l�� ��p�Cp"O�q1�
�z᎜c�H� dy�xr"O��8hB�о����/fb��"O�a��SC�F�pǫۏXfN<��"Oΰ��a�;%���bQD���� ��"O����C�h�:T+vĞ�[�z%�V"O��r�N�0��X�	Q�a��8�F"O,��r`�#k����ȗ~���f"O�u�VC�;pF���7a^}��"O 9���t�Q��V	)g�ċ�"O2|�2%�Z�8k�)��at����"O�EPT�D�MZ�И�'6P�{�"O*�s#�V�O�u��ѯd����"O�,Z�M�:\�,p�Z8iT^Lq "Oԉ�c�����r�.��N_Z4��"OvuZq� wƴ�'��%ʐF"O��!ਛ/n6\X��ſP �q�"O�]�Q �4	N�� �M�[���4"O|�
GEU�lf�8�ϳy |T"O���I�W���J�&ů\QFy
A"Oh���zҥ�g�[=*�b�"OP)CD�B�iu�\�a/y*�$��"O�cg���>���J�oT
P��"O���P�Φ0��уM�7
�4��"O JN҉�6�Q��D��.�"O^�8�V�Z( @8t��ag���g"Of�7`�*�`�)���W���4*O6����ܱv���
�V�s��1�'e���C�	���cϝ	�f�S�'E��1A`ʐy;Z��1fye����'�Lِ�cwJ��PPѱ$���z�'�81j��p��m G�A;���'��cƊ	#JR�0:'@";�$�H�'|~�DI*%R2��fG?�h4I	��� R�Jt*R�|.DT0&�,)c!y7"O�)�k��v=5��C�?ri�t��'<=��׿��	%I�.IC1�O	6xձ��� C�I=7 ��R_"�8M42[�O@�ib��jg�t��Ef*�0�g��p�y�o��g?�B䉺�Tͩ�)�?H<|9� iU�(}��Cq.U\~�a�+W�T�}&��W(��'���"�1g�h`��+����Ø+}N�H4�>H�Z��a&y�h����GE���K��Eʂ]$t�վ��b�&�w�@Ah"�Ō��]�J�q
g��V���o�J�E���W�<Av��8sD�!�w��*��d�Jgy����dL���"�>,�����	�;|:%q�Ƃ+H4�`�C�f�!�����[d���o=�с��D�I�t=apAڸD��p����{�Z��]>�<aa-��u��Y��)V�8;�Xh�KsX�H��D�5d(�y���G@�F!�g̍.k��s#,-X�`xxU�|��`��	� F���+�e���p�.֊YJ�<١%T�&J�ۥ�c���(T�����O��	�@�&�����6VX���'���w��9\���-�8ĩ(��x�ց[���1%vd�q�I��E��w�rd[G�hW����Z[(�B�'��lĄP��* ��/��u�h�BI��A �#I��R˟4���o�'�Fi��#Z@���j\�t_TX��n��Y
W%D�n�PE�+�!l����@a��q��i��d��%j��^�I���P����&�]�Ipu�fb�f���D�l3�v�c���8^�:܂��51�l�SSY�@�C�^�(�V�%\}�PC�I$	��`��b�K�耺t�F !<U�`om�"A�F&S{^a¢���.Y���4�sޅb0�U�Z�b����u�j�#'=D��hB�+�G�4���$LV�a[^�8ⴍ�t#�/�J�z�cF&G���0��J8 �Kt�X%�@����5���d�9,Wfܢ���6 H6��t���c��y��̒�{�Թ�L7nH��Cv��5Y�$!��I"c�(��F�Q��q�%W�DB㞰����'�-���j?L�j�L�)���0�O*��R�Y�8Ć��k�?T��yC�'�8�"4��mA�XId�<P�zlƩҪDL ��$�B��kE���a�0��~��x���T��sƞ��vg��F�D�b �,D���-̸v�]����(0��A%i�t���;'�i��\Ӳ��Q�����9r�Q���'�~<�
f�XC��b�7\O�	A�%r�����D�thVH� g�iؤ�8��^)d�,�AFĦy��-�K8���q�_�jQr!���U�Sjmke�#�	(����`�f��}�����dȨ�k�t�]�E����ȋ���@a�
�yҬǙZ��BF��Fw.`['*5p�t���.��`͸5P'��v�:M;���k���-�!��
$qiJ��nD�M�!��G�E-D��3�%Ji�A#A+E�3�v�S���<�@L����5�Z����D|�EA�JZ�#%AC�Q���rPEX���=	U͟/S�����AKx�Y�͔.J�x�t���WZ���	�N��	a@v@;��Qfѣ�I�+id�#<i�;.ƈ��F�Sy�O��Q��{�>4��f�!FX�];�'��!q҄٩dH"���Y'7�F��qO]&O��Z�Rz�)�矼
��%�����_�q��\��$D��+��<,��9GK�h�
ݛQ�"D�P!���s�v��@�eF�89�� D����&Ǽ_v@��n"tMR)� ?D�\#�FݏB,�u�p�q$}�cd?D���E��:�\-�fC�S���ڷI1D�xB�ٰJ�=�[��40��L�!�$�PMz�Q�Lϔg�MjA����!�dJ�Oc�)(e�ǝ	�����x�!�dӪ}G
8�D�=*Y>ݐ���*De!򄏛[ǆ�p����x@���&�#?a!�$2�	����7DT��(�84U!򄜫YP�@! 6�������:G!�ĝ3��Q�m��<����-�I!�$<vpƱ�5J�7)R}�흽P�!�YGB�뵁9?�@�\%�!�H�Bx�A��� f���oB��!�^X�u
�@�N�>՛�?V�!�� H�8#�Ϩ.�������H��"O<�YS���@6`�2��<���"OHU�A��_`��,*	�}S!"O��#L*RL����!��n���[u"O�YA.��U���ˁ,전�"Ovyc��ppSS�I49��"O�x�/�t:�h��%/�Y��"O�AbU��eD��
Ts��,e"O�)�V��/)�(b�j�3��J'"O�aCP�2�2H1		��!S"O��0�ǻ�P(r�h3�a�R"O�3 (D�/,
9�ѧ�M��@JB"Ore���L�D0 -8�������"O0DR�����|�*�G��w����"O�����$��xYW&A�T����"O&)�e��x���%�����"O���ូ�Q�O��g�d�q"O�<�P.�DX��J!a����"O4��B��}*8y-ȈD�����"O��FYp���B�M�)
@}Y�"O�i3��$+,PP�6&�p�\}��"O�u�b�ށBl��)��J�
��!�"Oz(c�_�}P�Z�gU�_StJ�"OĘ8@��T$��D��@���*W"O>�s�cI�1R��PD�rQ�X�"O��P*8&�,��Gʞ		@�qA4"O����ZTX��2G*���"O�T8ң��/�QF���]�D"O�,)��		~Z�$SV�F��rA��"Oĉ�J��^��c��X�A�p�&"OR��R�!Z���Ыk� �I�"O��"�ŽT�^�:dM�/r�6(ʒ"O�	bu�R��J�.N_UR�h5"O���Vc#����l��s312"O\m#�L�6m|<(ؔs#f r��>D���,�w�	j�&Gu� ��"�:D�X �/���Ƭ8��?
y��ɶ�?D�8� ��#~[1�2>K���(D�䛃�[�^(��y�R�F�����) D�9d*��/,���BM/~HD��s�;D� �a�Z�H��5���)L�f�2�9D�xa`��b��[@\5B|<i��:D��ۖ�nz�8	d�� i.H؋b?D��I�eĜi� [��W!FdLB�N/D��b�ؽL�V��'l�lE*D����.F��Za!�d��F�z��&D�hI� I�6�J�k�*L�
�����$D�x�����T���3rf̂,D��3EߏN����K�B���� D�$�A��2-��zW���8��<D�xs1 鶴�5&ݝD�
����6D�4ĂT�-�-�]��0��8B�	�z��L�k:@�J e۶)FB�I���p�W�eB� x�W�$:B�s��$q&���8�p@��9SB�	�H�vE�C �Q`�����Q&C�I�� I�bذ�d�b`f��C�	1ne�zs�é�����`�=�B�I�q�D�1l�96eHAk��A�O܀C䉩��L3S͜L�N5�C��m�~C��f��LD��~���&�6QMjC�zZT
�3M%���o��bgvC䉟s��3�-^3k�U�@�	/~W�C�/?L�H�c:&�X�с�8�<C�)� ���T´C�uC�m̊��l�C"Op��3�;v�;Cl�{��љ�"O��Bu�ҏ_o� �,�p���S�"O�]��MތH/tS�!n�x"O�����,
�Y;7l�a/�ę1"O��hW��(F��Cu���[!"O\���C.v�I�'*<���"O��#�P����"�$6.�2�"OI'$D�z�x�x5!D�h����"O8k�@<DZ�$����<k�"Oz�J��;|C��r��{G�!"O~)	��F9k��|���SJՋ�"O<)��G���6a����aZJ	Y�"O��B2�;1�A�a��"���
�"O��{`@�)�\��/iwԜ��"OVؚ�+�b# %P� ���2"O :D�4K�tض���9kBi��"O��jo�������4m\2�ڇ"O,ܰ`Ʌ��89�����9ؔ�"O!���?^�ҁr�(�Z��<3"O`@�C��6}�l��B"5���@"OF���2 ���K"�A�!���j�"O��ѱ*�+g(8��oB��� �P"O�}��͈���bcy�"O�0ʷ�3�:�b,	#(_\�HA"O@-y!O	a�)4="D�[�"O4X���}�RHt��'�]ʢ"O������Lɘ��ۋ�I��"O��Y�A�|�*�8D�� #��Mb�"O�\:U��+��m��'�(�� 4"O�]����`�ҥt�ɉ�X��4"O^�Kd`�,��m!0e�F�V���"O��"񥆉|��,P��FPt�xA"O��' �:�Zm��E%29���"O��A!IQ�����4]-r90"O��V��'�\����w0�{"OVɋb�-���c*�j�$*�"Oh9�Ř>*�����
�z�����"O�ZÐS����rE~�\��"OL�y��Q
��ue ]�`�D"O��4͵EO��aD
 0��k�"O&�$R1=t.��֗S5��� "O$Y�a��6xA���1<�
�"O�E9���$(�9�nO$_>.<h�"O��8g���M����a*ļGJ���"O�E���Lrb�8��U;D� Y��"O�x6�ҜX��a㗢��� �2O2���ٵy&$��1���$�1 ��ɫ*ϒ����,@�X�$�V�f0B�I�.�BMjs�_&?�����('3ZB�o�n�x��=*}�����L�h�C�	��� o\��Z-)��Ȗ����(?q��U�~}�5��M��`�<1ԌˊX��-q��UQ�H�1U�
w�<�a�¢��@` "�k���S&)�l�<�*j.g�=�.Ԫ��_e�<ɶ疼KpxH2'UM�ܐ��J\�<�rُNHcƝ=S$pZ�bRX�<�g,֢?%v���G WE�	��nJj�<���7h�� ��DP��	d��b�<rDث��E�2�r�,^j���E{�G(�����"	�2��x����u��<q�����'v���yU�C�2LP<����&WQ��9�V�4I��ا(��$A�أx�}z��Z��76O�9�'
1��?y�>0nԐK: ���E��E�f^��D	�����?� ���Ԉ;?.�Ivcէm���Z���H�'
v��i�'`��p�A�&��Ua�.��Oڹ��i>��\�`y��S�/ت�����!pz��%�P{7��o�S�.PX�g�ݺ>��S���'�%�'���a���ӟcԘ����! �x|S`�ٿZ�>����(O?1�WDϺd�	�	��ł�"ac�<��?3mZ��kMe�2]
4*^�<Ys�  ���'eV
K��,jEq�<�%[�M̆���d��#u�� ��v�<Q�O q���A(��(�6��G�u�<��d��*��=�t�zA�^p�<U�K�N�0��q�5JӁ�v�<���%(�p�ڇ�w�p�³#�r�<A�čA�Mh/	s$��+��s�<�0�\�P�2��@�߂��!BIW�<�� Й-�0�c��,+5�CQ�<�AI b��e�,j�x��&h�<�r�S��Hf
�*�T�#ĬNb�<�p�O��t���n�"t�ƽ����C�<!4�TPj�!]:�����=T��J�M׊GP�[��(1`��,D�$��h�4���CF�0_?��;�+D����n�?U��P�a��t)�	��(D�v�i�ê���j,�+^Rܘ��'c�0�����8�ʹ匊+j��x��'�\	/Cd'���Tˉ8_(rt��'[D��@�1~t��3����2��'��Ĳ7�ù^�003��%Py�i��'z`a�� ����oV�xXҁ"O�Q��R��m2���e{�"O~���
Ւg|��f�OV�8m��"O��{�jP%H���S�|x�0`b"O��"��t[r:�o#O�\"OT��c�޼G�D����G��};"O<� "Q�Ԁb�G�K��9��"OF,KՇU>�\tq��2\{�"O�Dį��@�y�i�6)�NܢT"O�3�Z�i�D�V��D�aW"Oz��S�L� �q�����p<�"O*Ⱥg�?}�x�Zu%VT�\y�"Ox�Z �I3"\���� ,:̪w"O�$U*.�:�c�@�#m���@Ot�<���4\ܦ�S��R �e �iF�<�0�<QLxPc��X���t�C�<i���q4�rD�O�S$BY��|�<���W|�qhEF�	(�\��NJp�<��-�8vA\�����f3�4��YV�<IuaN��{&b�*�n!s��\h�<���:H
fLЙ�4���Ίm�<��@'NO�E�D
H<�!�:�	���S?�b��v�C�!�d�;�Ԑ˄HG�a�Tat(��=�!�d�)U:,hF���p����>�!���f�p}�$+̀{�d�<D�!��;�p��C�� n��i�cܓn!�1y�J�" ��J�����4x!���+�ΐˑiBS����T�'
!�B�=^�yжK��+�>i	��I�X!���(}���#T�2]*6�1a͌!�σ.2 ��ߒy���cj<'!���x5f�s�)^�+׊ZD�C�{�!�$�|O
͡P#�M�E���	>�!���
�3qO��e���1%�ՐF�!�� �,��l�0���!"�M�!�� �4�se˥H�N�s�)��aQ*��"O�ɘg�ωS��E�O�{1Δ�@"O<4BfIE!g��0���DЀ#�"ObT8��Mӄ�x��>�@��"O~��@��Jy����(��+�"O�ܱP�GC�0��0[ɪ1�"O.��"i�&E��ð�>�.�k�"O@з��&/6��j��LĲ�"OX�C�jB
8��i�>��9;@"O�ҥ�%HcV�۰g��i�DQ "O��`Q��6Yd��(��[�B�Q�"O�lySǅ\��j����\���p7"O&��`�M:����83��ɉr"O¬�0�)[�X��W �F"F1��"O̙��A�"_ܲ��ɪ��/E�yrN)
Ll�����	�~�� ��yG�L<b��d�BVI�`������y�
ڀe�$Qum+c�<ēE%Ԍ�y�X"�YG�C-^Ȇ�B%O*�y«��l���b%l�;f���8 +@�ybM�2<�LAbq�-
^�,��
�y�i�d���r�9|�´3G`�?�yr�7|���8�h�KB�K:�4�ȓ_nq�1�ѷ	N$萦�+O���ȓh0�"�����['Z�9[�̈́�~s��b��!�r,a$EB�2�:Ʉ�,,x2V
����i����%�0نȓ �%8�mX*���V�R�5����!!g	7~u�����ޒ
��-��{��T�&̂��ʔ�We�)-�l���$�.y�p�֨Czm�f)�r�L��t�RI !��+;�4�F��ni�݆�7V�m�"��Q�F��e�%���|g�� 瞹+�A�SI��j �i�ȓ?�*	A%r�lx�Ğ�_v�����s�K�����E���i�`���-��1 !��R��72)h͇ȓP�Ј��ŕpf�u�i�	hE���(yy�B��WQ�|�'���8�ȓj�"�Y��XZ�P�(�*n깄�~�*����	�y���TBD<XSd�ȓ*q^��m��h!<0�&��k���ȓ���1���{��)��ί>M(X�ȓf��" Z�h�b�[�wX���G����׋E�7���$Ҽ~�怇ȓx\t�h`-��7P$�s6"\"h��@�.��b��	=�|�U&�5��}�ȓ7b� �I��T}��	WKP�r�J�����QCːx8�6�3A��9��b�� ϞY�at���捅ȓyŎX�s�R�q�X�x��A�5����^�bd�d�@ ��bBi��<�F���elv��S,�gꌨ*��� �Ą�a7�$
���T�,l�րB�4���qr|˂̀[w��!����y�ȓ	>ژ:�I�es���.�(Y���ȓ_nD���M�8�%�P�ը�2�����cGGD�J�, �Rl�ka*M�ȓNX�z��߁	_$��jӔR�\���0���g�TE�4��c%��sC��ȓ_=4�RDwfe��KW+E���ȓVs�T[��?/����R/T��0��G�r�J�
aĐe��@�7rp��;��Y!	�01�A���S4de��S�? ���O�>+�TMc��	3LY"O~��#cP�Qy�tP�h�
N4Y2�"OJY���N� ��8�i@�dhm�"O�e#�AYN	��&ޮh슑�#"O0�a�k4m�~�c(ҳ
s�}��"O,2��D1,a3L�:;�Q� "O�u�L�� D��e�"Qƭ��"Oޭ[��/�>�D��RW
̊A"OX| f��&q�8r�M|<\�P�"Ol%�r�-%�uʢ�!4-"�z"O��pʍ1m��M�D�A � C"Oބ�IJ�,a��Cm޲|z��"O>�+�(Ē_d���'LJFRF49g"O�8�FJ�{A���*�<1�=�u*O<e�#���KO�M���f���
�'=�Q��#�o���D�r�ؕK�'*|H���M�5vјU!�>�&P��'��%� �!z$t�����G��k�'��G��%�����a��P_�eq�'�����	Ю6u�� ���I�H�0�'���Bl�=���1� ҕx^��z�'njQ�#�!=�TE�F(H�;�xd�	�'�0�ڲ R�,\�+#��?3���A�'��[�l�;ޔt钣%1�XZ�'}d=q�OT(+l.������(Bd���'H60���̅
�;�!V7%:&���'�jh�C���&<0Hpd��(��k�'&F�;�Ζ�5������$���#�'8
0��j�c�m��5p����'�,	#���d
d}8��ye�a��'�ӄA �"G>���mϚ{��IB�' �����C��V8��d	@�G[@�<�&�t����7P��A��x�<�b������(�i��8��ae/F~�<a�fG�`Ɇʧ��
7�N��ZA�<ԅ:S�6}��A�npj���g�s�<A�o1p�u�0
8�l$au�Pl�<��N1Rm켁`!�%V�p��	B�<Yq�D�06U�a)N�q�v�#*ST�<�E
�
A�]hP�L+"pP���P�<��ŋW���	��I�x���+�g�q�<7b�'Z���he H��b��Øm�<9ԅ��K�\T�F�ucd�`��!�yI.~�8�I�G_
���
��y"�,7Cz���^?B� tH�hܒ�y��7C�\����F�"ȑ�V��y�%SA.���J2Bi� � �D��y��b�)��CR�:����ǆ2�y��D+v�^���AL;�ptYrb��y���	�@ب��S�d��ac�B�y"	��j�Bd�T�^�`J�J񫑈�yRf�.j�1F�G�j2 ��֪�y"Ɏ�=�e���K%��M�u���y�fD=���S�H*O˒���I��y��$����hKS��� �0�y���[����$Ets�ّ����yR/�=��Ҥ�O.W2�4�_��yRf�D�n}��K�op �	��y�j�)5�n��FJa8��K�AR��y�Ȁ/I<�0eŔ�{�`��P�y����f1� ��M�k�hI��ˋ�y�oA'!>������dq��T�
��yR��zGJ�B��n��1����yb�?%�R �7.������y
� ���ЂE�'�X�+�.;��2"O0z'�T�[��U�K���6�"�"O�dxV��	�^A��*ɡe��I�"O�A�VgV�m��u��	�$DB$� "O�=��E�#���
--�\ �T"O���biQ4j��-�t� V�z�1�"Oaa�bU*�RP;6�� ��٦"O��X��ǆe=@
�k�=� P��"O�I��6l� A�0�
, �JQ�"O
a�� �Z����g�'g� AI�"OĀ�f:M�T-3�
�[�\�"O�����Ǫ?��^�D���4"O��x�
   ��   �  g  �    �*  q6  /B  �M  zY   e  p  �{  *�  x�  ��  w�  b�  ��  �  @�  ��  ��  �  ��  �  w�  ��  C�  ��  d�  � 
 G � � $ �+ R5 '< kB K &R Y \_ �e �g  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE��DG{�𩊺9hl(&���洠�H[HGQ� D��݃nĪQ��E;^ҡh�;���0>����t�L���:$�0z�N�A?������Fa��d���<�rf0v
���A��
B�I72���H�A8|�J�8z�'A1O^�=�;c�`гNO���7bێ
ޠ�ȓa�m�'�R�:�,6Ή�aLR|��ē���)	,b�ga\v�P�	E���C��%+�ؠ�U�.���0�ūYLC䉕q�(���#�/�m"2+׵��B�ɝ#��&M^�p<�رo�4�C�o�����-(��qW�R�Qn�C�ɱN�<A�0�ߔJ�H��"қy��B䉈~������Dub�ֶB�	�CcΡ�����	般�
�;o��B�I5�݉B�I�-/��{l�"{L>B�<NQx%��,:Hd@���(r��C�I&yp�	u�E�RI0����Z05�C�IlC$,�'��^b0z��r�~C�,���Ѱˊ�-�Nhir �&e�B��+v�qӁ��2n`�� ����C�ɐY�0Q���@�<�A�#��Q��C�I/'=�d��J�>+�"��9�C�I`|�y�O"H2ΡA5�S3��C�	]}�ѹ��b������10�C��8eJHjfE�p�^���֒h$ C䉌+����3�7J\6`3�Ԧ��C�Ɉ Ta�˜)��ۖH�!h,zC�#7�h����&���^:>C�I BDBuA"��>u%l4��>/0C�ɏs����� 
�>t:-�O��B�I
I�6!�ό�Q��-� Eη��C�I}�������9]��"��ޢG1�C䉩G~�z� ��w( ��pG��C�	OF�)��J�x^H	�H�[|B��E*ޘ��C	[S�UB6��lq�B䉶sE�H�,@$˳G�z,bB�)� 0��F�I$K1�i���?7>$j�"O4�����.:����EB<6�ڗ"O��f�?��X�����^)����"Ot��������� �J,��k�"O�lw���7�� 
��@�P�:��"O�XG�ۅ ��P5i3"�p$ش"Ov�i��ĝ�`"TE�"�isb"OPE��zhr�����rG&hJ�"O 0��-� L4���= 5��P�"O88�G�Oo���QF��v"&�C"O@MB"%b�m	�j�7}f�}��"OE�ƚ0rH�����y�pғ"ODp��܁;�P�ѩĦe�&"Of�9e��,���*	�4,J|�"O¼i"A�|���S��%*q����"O�+���GJX����W�БB�"O�iR�������x7�bD,���"O�e�4']QByS� �"�i��"O@ĐP�!ifl+PZ;!V0,��"Oj��J]1R�*�P��Q!7�y#"O�ݹSF ;�zh�oԶ B`�9t"O<�32L郳��)$ى"OT@;c���g�p���.[q�$ S"OT���&v���A̕�)jDM�f"O���a⑌�Lay4��&}� �E"ON����ȚT�PR��@$G�FŁ�"Oƅ����U�4��c�:m�$d�D"O�����b��8�TɃ�x�4tZ "O�<� �'����ɕ6���@�"O�q��O6�:$�Q6m�vP*�"O��b�-gA*����ԫb�^��E"O����yp44�R擄h�\M:�"O>�2��J�>�N-���_S;V	��"O�tp���vB�͡�
?=�)��"O]�aiW�lsN�#�*�:]lE�"O
����@�9�T�;�cC9G D�"O~1�"�(1�lS(ŗ���X�"O�ᇀ.K}<ݐ��4�ذ��"O@hp�(^�{�r�1�ײf�~��"O�D[f퍛^��C��Ո�40��*O<�7T����z�(O'�ei	�'?,�CVś�>�uHuK�3�x���'L�@��+���ű�1*tm�'-�؛�m��M���
BoŀM�
�'M~��s�Î.��L8�C(��%J�'H)�%��|<�@*Uk��]��'V��z�H��9YT��>u��m{�'����ıYa�u��Dʤf�r���'/|��bO""r"u�HQ)T��	�
�'cn{���$��ts��<t<�
�'x�dqM6��]r��ˣW: �	�'��0�qLB�Tc �y͓�w{�c
�'�(�$�Q�w��4a��k��`�	�'� �;� T�~�,�F��j�ޙp�'�`Z	�ұ��Z0#$�b�'1xR�B��C$�H	-N�/�n�!�'VHI�B�y�F�{"�P)�yҎ�,u�����E�:X��H�hנ�y�@���h�h���R��`21�7�y�ꓼGN��!� W�9�`͒3�yb�M�UZ0z����*\��"��y�a�H�v�B3����(V4�y��0a4t#1�W4��ax��Y�y���7B��x���/8��l��y
� �8���,�B�!$����"O(�h�톤&�jE��Hތ-.J]�C"O�9�se�������*\�"O��S1*��.����˘�|��x�"O8�:&U
RI �e��V�Tm)��'���'��'���'��'��'�<�k� D�s�jm�$jұ�ZE$�'�'���'e�'�B�'���'(4�7�Z��,SҦU�m�����'�'���'���'
B�'Q2�'�@�'
H� 0���P�\, X�P�g�'��'k��'��'&2�'R��'����"��'!�E�/�S�va1��'���'���'���'W��'R�'P 9:�fE� ה�kH�!| ����'���'�R�'�2�'�r�'*��'��D��
Wì�#��ư���'3��'�r�'hb�'���'R�'=t���ˉ�S�t�J<���q�'���'���' "�'�r�'6��'�x���Ӎ^���� �o�&��'2�'�2�'�B�'���'���'�x� �N8-�����P�G2F���'���'Zr�'O��'�r�'���'B�!#D	�1��Cwא#:����'MR�'h��'wr�'(2�'���'EQ�B�8U���b%��Ͳc�'�R�'7"�'��'��'���'�N�C!�B�]��@�1��x���g�'��'���'���'I�'`ӫ�iG�˒:���D8	��Bt�P&W6�ʓ�?Y*O1�����M����Ox�e�X�|�� 0�˞{�
H�'S�7�0�i>��ퟐ��GE4$U��7\�ZqF����	�C�an�P~�2�@���@��ʈ-��%Q!� Luc�L�!�1ON���<�����)Wܠ��&�v���f�g>)n�J�b�P��^g��<�z�ϛ	r�6�[�N�Ŏ���O��y}���ʛ�U8��0O�aD�d�6Tr�cT/o�\�Y�:O��	��?���%��|���]H��؏�*� �/��{d����(�D���CA&�I��
I�p�E&V�T���+	B�6��?�X�H�I���ϓ���q���+tB��sF��rUd�'���lj�j��1�c>mb��'0ޕ�	�Wn����.]� 0���.?����'-��"~�Vd6���3!n� ��L$�P-����j�����@ڦ��?ͧw^4ı��Ԩhz��[�M��?����?A�Ɨ�M��O6�S����W10C���Uz+�|���L~�O���|2��?Y���?�ifm�2 :U��h��|%$�<w�iUR�#P�x��k����SE��L�f1kP��5@V�$J!B�����Q��YB�4A+�����O��Ĉ�8e uR�
S���!A�Ui�І�$��hH� q$�"k�N~�A���$4"�@��e�+��@� 4��O��O��4�:���!����dR�
֎� ��RZrx�G�ϥ�yGyӸ�h;�O4�l��M�i�rY�7b�<9�b੤J��|[D�S1 D�ao��;O&m�R*`�����4�OpF�C!�w�@}�&�Z�Y9�u�t�N:}��ъ�'cR�'d��'���'j�RM��"��!76s�Z5f��x�B�O���O:�oZG�P����b�4��4��1!&�M�p�*���ܷd�"!�x2$}�oz>AI��립�'k8�b���')����3�Ġ�o�8$ˊa�	�A��?�Mk.O�i�OX���O��HcƆ,o��8�&@���F��%e�O�$�<I�i��;��'3��'&�	}�`��-ģG�Q�Fg�#9��������M5�iӰO��韈|RG�J��򁪕��c���K�D�'X�8lcq�(]��I�u� �ʟԊg[��� N"�Pq�CD뮑 ���:�f��Iܟ���ӟ��)�SFy�Ld�|A��+��mI��pdlH8A� ���B�&�dʓr웶��Ix}b}��!�T튬G\ JR,<>�H��cE�q��40����4����jt(:������Z :"��.�����N�8HR�4��D�O��D�O~���Ov���|�p�Z��<�Ǯõ3���A��(���@J>G��	��x�´�yw�I�Q�C��*RNN���R�6�W��)�J<�|���H��Mk�'P6��Pg޽k�$L��fЌ%f3�'r䵺f���X�Q�ؙ�4��4�����3?�,���Ֆ90v�x7c�;���D�O��D�O����Hܸ���'��K��/(�\b"!ן��%PPlϝX��O���'�6M�-�O<Y���M��x!aK��Z(Y⋟Y~�BB�z�z�p���<��d�ĺ����O��R�e^�͐�!/n�j�{��Y�b�l���?)���?���h���$]�� ��B��e��P���I"��d�Ҧi��ݟ����Mӊ�w��@�M	{�8:��5l70ݣ�'H��iad6�Ĩm��7�2?#�����铗v�^L���+lNLp@����"�c/O�=m�cy�O���'���'��H\:�v��ɜ9 l���4$��(��I4�M���%�?���?�L~���E�!�N�[�}'��\�p�شE��$��)����WR�\�ƌ#�֯7y�8Z�ʺ��-_5�a��'�:D�'�~7��<qT��t�@���.!=��*�/��?����?I���?ͧ��d��{Q�����Jܫb^Fyb2F>H,Q��q�8@޴��'��������Ox7�ΧN���PP@ƔWa����!J��m�odӚ�	z�2��Ce�K���yq��ߟ���:(��=� u0GG�V�QY�D֝d�~��:Ov�D�O����O���O��?��������ƫ
�@�%,����������ٴqt��/O�4lZy�)A �e҂	]98� ��K�#�v�
L<b�i$���O����i��	)A:���oǽ�z5iA+�'P��D�P�
���Ay�$sӚ˓�?a��?��5S�l���g���pC��%��)��?,O o�2@E4 �I�L��P����q�-@�ìF�Z��%	����XD}"Mk��5��z�)���V���
Â�/V�bD^A+>P[$Έ�,Lر+O���B�������4�p�a��5l'�9P�ݞL�*�(#�O`���O��D�O1�r˓��ᓭi�$�[fɀRV�ԪN���Ȓ�_�ܳ�4��']��\N�ƭ1MZi���ʇJ�.�2V@�B���u�Ʊ��+s���@�D��Lk,O<ت&�,4Ψr	\<%d��bg���'���'[�'�"�'���"1"1%e��kK� 3gD	�b�ڈI۴/u�(X/O�D$��+�M�;�X��T��8 �� P1�iB�T���'���|J~bdD��M�'��9PECJ`I�<��/ך��ə';�LvDHџ�iAZ�ؐڴ���O��D������Ȓ)U8x4��Vl�p�D�O����O��4O�ƥ��j��'�"S	7ö�Q���\��MQ �/+�OԴ�'�7�B���'�H�PA�$i�8��U�.aN�Bc.?Љ*N�D'��.��纃��Oh����� g\;R#� ��ƛk���
���?���?9���h�"����bBP�p%��	F�(c��͚�<�]Ǧe����_y�cy�����n%��R��D�y�t("��ˬ@��>�M��'Ǜ)�I�ƚ� :V�K.A��LH3��0Ɓ/qb�R(	�E�q�'�J6ͷ<����?����?!��?�A*��}�%ɚAM�8'���9�(������ן�&?���|M�X����7�֌�AlD	<�Ѫ�Ov�m��?�I<�|�D��4bl��'
S�@��	UEN2L�ɓ!�G���$�<����PU��V� �0� �hy�����W� ��4��l���������Suybbp�D���ORu�s&��_�.�6���\�l�"6Op�m�G�	v�I�M���'^��Ԣ$�,lJsF�>� yI���*�"�2�i���$,��1�O�Ҽ�'�
�}�5f��������?t���BM8�y��'�R�'r�'���	Υ�]C"�O>^�J�#t&b#��$�O��$��	FId>��	5�M{O>�E�&Z�ur���08L}��'C>S�'�6��ަ瓿���n�B~��0MV�d[���51<�ST�&sz�7�
��tX×|RW�����X��ڟ(�!��j�#��B�6!�q� _�r�'�I;�M{�j_�?����?y-�F�"�AL>TٌE��f
%(��6����.O��Dv���'�����<�Y�/Y -t4z��D�m��:�ɘ�V0 ��L# ����?�p0�'��$���Qͅ�B4��b�X�ӐbE��	�������b>M�'�"6-4�6�I1�-����g��x�(����O��DK���?�Z��Bܴ"�~�Į�HĊIB�3HP
��i��7�ĝL��7�`����!w�F���Oo�i�'���F�����fa�4�گ�yR^����͟L�I�����L�O��I��`Ga~����H�(��{���ӣ�Ov�D�O�?Ux������$}d��k�āBI.i�mEa����l�L$����?��k�EoZ�<	�(LoLH�`J%K�btoք�y��ͫI7D!���n��'6�	�P�	�n*A��M��8S`���*j��I����柨�'�:6�0Xu>���O��$�'_�l��f X;
taz7�D���<b�O��m��Må�x�etU ���Y&�L%s$��7��O�2��a�n�m�H~�B!�O�m���snڹc�J�`�V��A�&Fu�����?����?����h�����c����C��y�4˴�F[�������9C��џ����M���w^@��L5
L(��	�}ډ:�'x�6�ɦa۴�.��ش��ēq�f�C��o5��z�M�po
i�e��/R���Be'�ĵ<���?���?���?I
"���$U�T#�D��������٦��J����Ο�&?��1h��m#V���~����#�(=Ĳ��.O��Dd�@�%����)����w�� �uTf�RG�I�^[]	W�<��jL-6n��]����D8dhP���=<A�����,CJ���OD��OZ�4�X���V�!�R�5zk�m�$AC>�`��	dd�,y�&⟜!�O�Pm��M3�i����'I5�@a�ѽV����@�ɟ;���Hw/�(z���L�����f���5(�F�œy�
� �~���	ԟ���ǟH��Ɵ���E�8!���L�0���"��/�?���?yñi����OwB�y�ԒOZl�P�Ϥ��HP���@�܁���v�	��Ms���T�7M`�֕��ئ���q�D�i\�Xp��g�I�h���`ι�?�%,�$�<���?����?�` �$a�d��#�ve��CBe>�?����D ަ���J�����	���O�8�`Ӡ�&S?�4;r�P�:� ś�O*�'"7mEǦ=pI<�O~�	g'T^��pG��6��(��Gpp�9�Cʹ��i>EI$�'�VT&�(q��T��a����7�ϟh�	����I��b>A�'H6��o`(�4���kK~D���-Z<^E��f�<�Ĺi��OfD�'o 7���)��I�`��C8c��&*�n��MK���M��O�EB� ����<� R �rN�L�D9�`��;=>��f?O���?��?9��?)����T+`�"3B˚a���-�3?��o�4Dd�I��4�	S�������ˑOM+L�fX��*$e�2�㣭��\����~Ӯ�&�b>M�#���͓ubp�@�8Қx�i���Γ> ]�b��OH	BK>�*O���O\��7���N̺�f˲B
6ɹr��O����O���<y��i,TK3�'���'P�cq.�:N��՚ba���������}}r�@��{�( %�Xw�;9+��B�G/q{����+?�n^�(S���K���'8W��J%�?�sh���J,�7�ܨ3��z���?Y���?����h���䔧$O� ��&NŒ);J fiV�$ ٦	Ō���I��M��wM^̑ԭ�>\a���Uբ�n��<���i�^7�릕����ɦi�'(Xu�����?�Ĩź+�F��Wm�;G�V�{�#��'��	��I�����ܟp��?�����J,Q�(ɢ7	&	��'�+���6âm�����	n�s�����~VTµ
��8�Y�������4*����OY�!ႏ�%���B�NG�'��1�n�W��4Z�l�G(X�Kk�l�{��sy��;�>iJ`���VL��#���Lb�'�r�'��O��I�M���L&�?)�(]�T�>���,�B琥���%�?y�i9�OJ��'e�7�
��YܴpsT�;�b�2��AsvGN�p4�u�X��MC�OT��H؝�"&%����
(��O�v�*�Q��H�p�c7O����O����Or��OR�?1#�O�2
gT�Z�h]�g�R�#�$�I���4^9v��O 6m'���A�4�Ы��,n�\�v�@ �M�N>����l��?)��Ħ���?!D-<6ib��c����K�D�99�ʍ�f�Or�	J>1+O��D�O����O�X2Wk�O��4bĪ�{sm�O0���<�Ľiۊ����'\��'��S23� ���(BD�aʔ+��{]��̟��	M�|
�F�\�M�+���ܑJ��H�am�<�TC����9*O�ɓ�?	��!�$�
J����-�7P�� �D���d�OD�$�O:��)�<�f�iTP�ƥ�(�D48A`Eo���a��jXb�'�L6m4�Ƀ���ަ����<s���3��R���Q�W��?9ߴN&� Zش��޹qz���',��ʓK<p$₉/�~��cJ+bR�8����O<���O����O��Ŀ|r4+�+�P��%m�,X�æ�%b���D�r���'t���Zئ�]70J%aѨ�&��s���*`4y۴-Ҕx���甲䛆?OzxH���m�b�,Z2�&� 0O� m��-�?q3J+�d�<���?�r/�mL�i���O5'p�SD�	=�?	���?����dئM��K͟���ڟt�ud�1)��C�N�)<�$}(�,�W��Z���ԟ$�I^�ɲ���B�ɐ��B��N�A�
�`	`�҆� �t��5L~����O�5S���h@6��u�œ��<��X؟��ןD�	Ο E�$�'�&�9�E�V� X3A.��$hPm�v�'�6m�M'��0��4�4�L�"��yd�	�F��t��6O�!n���Mk"�i��K��i ��Y�}���O9���� �:zfLx1�H7��� ��l�Py"�'���'tb�'�nO-vG�)�FD�'^�����J����
�Ms��_��?���?aK~�����C�Ѷh� 0!WG��^�%T��I��M#s�i��O�)���).c�}�uN=�� X�[9��Ǌߧ_/��c�|�F,�O`��H>.ORݲRL��S�h+��X6�8�c��OJ�$�O�d�O�<)ƽi���8��'#*I�t� �Pd��*Ɂ�*��'P6m9��>����ҦY�ܴ���*�";�ν��)��xE˟ndM��ij�$�Oh�ǍQ��'j�<��ԿSr�`Jx%P��&s��*�T�<m�iy��'v2�'�2�IN�}�๡I�R��I[v��=����?���Y��v��Qr�	��M�M>��"_�$Τh�� �=�x̹�gɤi-�'�r���$(�	؛ƞ�`c1*�![V���e�W�D�����W�,�6Y��'ixA&�L���D�'c��'�D٨�JcЉ���2HG.��'D�U�4��4I�9*O��Ĩ|��#E1>��QbSfɸZ��Lb3$�]~b�>a���?��x�O����4��pi^!�t��N͵/��ؐM���2�O��i��?)d�0�V2_��kb)��z��i�IG##D���O(�D�O���<�W�iX�%ìKn�:P�C��D[�'-Za��'��6-5�I���OH��2c��`:��Q` �2v]���O��m���lZu~��o	������Ovz���%.���,�#r�܁�'��	���ȟ��Iҟ���t����##�n�C#@ ���Z�cT�
��7m��Hi ���Oj�D?�9O&�nz�aq�G+1���#��?�p�2�������}�i>����-����L@ЫK�^�C����7����
��N�O�rK>,O�)�OƀC�C��	PiB�W�,�T��O��$�OD�$�<� �iѶA��'@��'ǂ	ԣ^�@�Q��IH�L��@�D�j}ҍ~Ӏ,nZ�ē2�tp�.m�푦'�L��'ܜ9�C�[�+a�h[���TA�T[@�'t��اh�!��X�&BP6*��PhV�'�r�'
��'\�>����P,.�c�/��c�����ò(lz	�	(�Ms�ŕ3�?Q�R��F�4�\�u@ƾ �rыaKϜ25� :Od�oZ�M��io>(ҵ�i���8m:�J �O�� PiQ���<9t�Y��| k��<��<!���?���?����?1���`��(Q��A*m�d�DM�����I�#K��4�I�%?1�	:t��Y�Q��xN.屔���p)�O�oZ�M�g�x���ɜ�G�TX�6*E�T�0K�o8�J X�@E&�剾i�
��'�,�&���'�Q &i�"-NJ� t,��~n@��'��'�R��D]�(kڴFS��#�mqȨQ��4x�a��<D��ϓI��&�$Gm}��'��'n��n�`�J�*�a��r�(�&b����� ���3 �$�����yp4�͵ ��xs"�G� ˄��0=O��D�O���O��d�O��?ŋ4��5u�nI��Gx���A�|y��'6�\-;��S;�M�H>�`�0,���{�D["Pw��v�ۖ���?��|�4H�>�M�O> �3��~U�9eDB�GS��uK]�1������TF&�O���|����?9��)sbź���~-L�0%'������?�.O��n6u�`=�������E��c���,�����EB�P����@B}҄`ӛ��*�?��&���W\�[v'I� ��B#��*lz�x��Ɨ�ex%����+�ٟ�	D�|n��	������0�d��jZ���'���'���DS��:ٴ�<��1NՄH�Ĝb���-���"�A��?��%p��\_y2�iD�5:�f��
:��qd�)��! 2�zӐo'�f�l��<!�3��Tp�蟘H�'ʸ`�	݁F��]���\�5R����'��	Ɵ�������������Q��G��p'恹#���l�(�@7�	#.�����O��D:�9O�Xoz�i���ҁV�kQ������DA�ޟ���p�)擂y�t�n��<q�N>f�� h��#完2s�\�<q�*�{f��˨�䓌�4�4���^`�3�[�`�P��W��''����O(���O��W��F C�r��'ibn�#JQ�����C� !����>��O��'���')�O^q�G��E��5"��*|�LPz���,k��=*g���&$�9+`�&��� ��36�^�sN4�Șq��G۟�	ޟh��̟�E���'T���r>�AY�7*	���'��7͞`����OP�l�v�Ӽ#��ç�.$�7K֚=9b%AN�<9��?���i�,��a�iW�	�pW�O>Fhݦ$c����:_����$��A�	{y�O���'�2�'Sr��&\l���E�)��}��f�$"��	=�M�����?���?�M~Γ�	�� �aK���aB](f�޽h%P�������L<�'�?��'~�l �F
�<mIU��a�������#m�`�'��ih��H���|"^���� ��hp^AiQ�8�x� 	������ğ��I���Ly�kӚ!��O�1���j���Pǂ�GQ�y�6O�TlZ@��}��%�MC$�i��6-�,Kad� ��q |����pN�Ԣ��v�.�hD�=v��|!K~:��8`�i�qc�(	$XY¢�3M$���?A���?����?9���?a�M�����8�!Eb�'PH���%�	5�������?�ʵrb7:�I�WۄU��`y�͸E#.L�k�,I�� ,�>�6M:_��$�O����h��T�g� �ȟ4h�kQ"�� U��s��@����)F��1B+@�J!2�'���A�'iZw��	��F�$�O0 �B�,<���E2Zx�Z"�O�D��E�<�7�'q����'�?���)O�{��c&���&pgB_�7J��ӟ��'��6-ܦɯO,ʧ�b���+1X�j��يy�"E�k�<H��ݹ%����'z��J���8'�|��֞-�d]����c���# 풔q1��'���'���Y� �ܴ4�ڹ��W5^�h�栁(qZ��á׫�?���9���$�C}��c�ڡ¥��)D�z��2�GH�����I�U#�4U����޴��d)@�<����O�v�hj�PeJL�nX���	$_,@�����O��d�O��D�O�d�|b�&ޢ>�Ьh�hQ%BFVȩsK +3E��� >r�'yr��d�'�t7=��1SAʍXvΠJ�jŗK���ab*�ߦɱٴ7�����O\��]t��6Of�qK��%Z��#Wwt�C�:O"��-���n��~y�Op2K��U�a��3A�B[SK�'K�b�'7R�'��	��M;��� �?���?�*��&Zr(��D�m�^q���̡��';���?�ٴl��'W�E�w���s����"�5���#�O6(7)�F1�xs�f#�	�?	���O�(7/4>����r&��(�8��/�O>���O����Oʢ}b��r�X}qǒ{{Xm9���K�]��$?-$��'O87� �iޅ[s����(��j[�]Op�2��}��شBu��w���i�im���,���0$$��P��Ak�5 ��CQǓ3 �zD�l��䓢�d�O.�D�O��$�O��d�6�^�y��ø�HEEɒ,>�5J��ES�*I��'$�����'�E��'E%-11*��&f�Q�v'�>���?q�x��tAˊD:ƀQ"Q�X�@��Dل�v\JkL������!/p��0�H�O|�M���3
+�ċ�C��5���?���?	��|�)O��lZ�9l�e�ɍE�@�ZT'ÖL7���m��*�D��� �M��j�>���?�i؄l0-��K��R�-�@�zs)��6_��<O\�D(ro�����i�֝���C̖�S��J3A����4�y���	�����ܟ���쟈�:��؉2�铈��p��,�?���?��i���Ocr�p���O�m1N҇!vj���'�13��jǊ�V�I������?�B����Γ�?y��Sx�? :�W�Ԗ9ؘH7;5��Y�鑿�?᳠-�$�<�'�?Y���?A�(f`���C{��zCfJ&�?!���Ҧ�1�(���������O��tQs���\�1�V.؊�i�O�4�'x��'_O�)�OT�@�@"- P쨠솝'Od���̰&D<�����I�?1(��'�$�����щB��ea�ޖUn��0h͟���ן@��ӟb>e�'9�6�C*ڸ�щ�� ��-��� L@�e��O���M�?�X��	�s�l��*�L�Jf�� �ɴ�M����M�O�u�����zK?-���'ut)(AS)�v�襪`�h�'���'�"�'A��'y�@��Hy�j��F0�f���a�K>���	����@�s�h �����:e��)�E_�s���F���0!ҿi�*�O�O����Ǵi�dN��=����<t�Q���Ri6�$߃7*��{��M~.�O���|z��qaf?&�B�C�� 2� ��?1��?a(O��l�B#X�����I�eX��%� 6X���Zb/I/|  �?�P_� �	ޟ�JJ<����o��P�-ŔcB����A�d~�+Z�)l�xpD�5��O~���4-�BAT�vU� Ȟ����acoѺS&��'���'���ş|����t��U!ѧ~)hm"R��ğ *�46
!�,Ojqo�b�Ӽ���8(2�@���]��Ě�<�3�i�86����ApD�ʦ��';�bukH�?%7%�)�F�i��ʤ��9D@G�hR�'��i>e��ן���П��	9(�hy��-�*0b�-A7	O�}�|���9g#<q���� (�(��蟨�I��MS*�D����ܑ7�O*_�\,�A��~��	�'���'��O�i�O���²f�r�"���5*�ɻ5��+�Rq�L����ɻ/���v�'�='���'�������9���	栚UH�E���'_��'3���$W����4yȪ��%�Zͺ�ǣ�8�4Aı�JIS��x�&�d@}�/bӦPn�M��ёyH0y��#�<�DA�i��ȁ�4������2��LF�����_�@&�V��L�w�M�IQ�D�O8���OD���O.�"�S�T˰��vB��5�f�kÊ�6E�μ�I۟��	��M��n����٦�&������a3 ݨVm@�#I����x�I����i>!��!��-�'� =zd@	X\�����d�щ��S�#��I�OX�'�i>����t��N!��Ņ�[d0+�/K#�J���ҟė'�d6m_�&ے���O��d�|�u_�4.ز��0�,�DH�N~�>����?iK>�OX�A��	�m L���.��}y� `����g�D���4��ͫ��7�ғO�p4NB��jue��!x����O��d�O����O1�L��6�O�4��*؍~����%	{�t���^��(ڴ��'��ꓥ?)�d��O'�KՏ�r�2�z�G���?���[zhP��4��$�	.�z�������i�ě�F-P��QF�$pRD�|y��'��'�R�'d2]>��v�w�|���'�&4Cݲ��M#�hگ�?����?�K~Γ;��w	Yy��BG:������o�����'��|��4�
�F��1O|���ቦaæ��!FǺa�f1x�6O���X��'�B�&������'����v�0,�D�gj��P<Y��'R�'�bR�0�شP�*����?��z�|a���e��*�⃥?L��R�>��i�|��%�dPyj�Ȑ��_~@\�5�UO9�ɿ���&i���-'?�ˆ�'��	�I3�\��4��Y�I L�B����	�����͟���f�O���L���!�8[��Y��4Y&��dӂ��OP�Pڦ��?�;n��XQ#�?�h8���Pע<ϓ4�fey�2�m96m��<���jo�ѫU���X��Č;ph�c�G�,t�Yۖ!N�����4���D�O����O��dF�| 2��X��hK�� �T���F���@LuR�'2r���'K�3��g6�؛wOV�dk��in�>����?ӗx�O���O��%����'#�V�����,$��)f�҃ApJDr�O2,�Q�X%�?��;�D�<é�t٫gk�kx�Jr�� �?���?����?ͧ��$Ϧ5zwG؟� ����r���5��Tq$�q�ʟ�A�4��'����?������b*��mד?����AG9�P��d�i��OJ�X"����'D����?m���}Q d΅����ɉ�0>��ן<��⟈�Iǟ��J�'C�H�Aw��|y�-Y(+�f���?���fmߟ���禕$�Q���@?�M�g%�.�&EJ�R��=_�Km��I�"�6-5?)��\���XQ�`3#���&�c��TK��O8�iI>A(OX���O����O�X��H8�a5�i����O��Ĥ<q��i8]�E�'"��'��S�TM
�+ �]�nT�f qb~���	5�M�T�i�O�ӫ!�b���OE<) ,��j[��6���(YGμ��Y@y�O�l5��dJ�'���pڦ	ތ����"|�p�'��'�2�O���>�MSЬ�B��Ћv.T%7�f䒆J,y�����?I��i��O��'2,7�:|,r���.(_����G��oڮ�M�3d��M��Oz���/����<�7�a6���:?�A8f@T�<.O��$�Oj���O��$�O�']9��i���3�\�ÀJ��\��W�iݢ7`�O>��O~��8��QԦ�]&����#>��ف��	0�v��4-`���/��ɐ�W}87mn�� Z!+��͑������b\�"�8O��AN�?Q �<�d�<!��?)c])y����A�-+ӾAQD�N��?9���?����������џ �	ʟD��JUh¬V	cސq"Nf�gC�I��M��i O|9H����`��i����2���#���Ӥ+�?X��d�%G}�7Z��G���h�QZ��k"��G��`�`jП��	�8�	ΟE�$�'�i�+�������n򘙪��'��6͊�0X���Ot�m�|�Ӽ3 ��81$�$��L�<������<q#�i�b6m���Ԯ馭�'�L]2s�W�?	�,�F�T)Pǩ.�+s"��
��'����<����	������c�^��C�v��Q�a��(�@�'	�7�5]��$�O���)�9O�<:B;��hqL˖P����`�`}�`�tem���S�'g5� ���-@�D���JF#\X�j!��	x@�Q.O|u(���?y�'0�Ľ<�1O�#������+)<���E�?���?A���?�'��D@��ݨ L͟��R��,c"dݘ��	A���K6 �ϟTX޴��'������My�x\mZ�n�h���N�Μx�M�3����R ��Γ�?�v�N٪���������h;&5ٗ�D'EJ84��	D�D�O�D�O���Od�$ �S4Z����U��Ye�l`��%&DU����D�I�M;�F��|j�;���|�TQ$������"\�p��Ŧx�JO�mZ��M�'G��ߴ����)l��ciѸ7Dh0�
x����M�;�?�q#-��<A��?q���?A�`!}����,�
�+m�g�j���O�˓0s�֊֘B���'R>)��H�0H㴐
����	zO%?q�X����ڟ(�L<�OV����ؘ Ϻ�����`dfYV%�1P����	��4�� "����O�A��)�3������C�D���*�O���O�D�O1���S<�V�Ih����Q�
�J�8�cIm:u��_���ش��'�8��?�'
�39p*8aǙ62(���sB��y�i����5�i=�	�8���C�Ov�є'�t5#� ��~�̐+�G��u�f�'�Iߟ��	������<�	e��凹}���	$GN&��H(�NְM&6-�%�����O��d+���O��nzޙx�o� 	�Y
�*��-:�9j�	�?�4J�ɧ�'z�e3�4�yr������Q�D/���Pv���y�Kڼ�H��		e<�'��Iϟ����
�\�
�<x ��0�C�mE���	���	��'�7-�8�$�Or�W��b� ��9�Zx��ˆ#a�t�p�O�o��M{��x���:y�������=a�E�5ǁ3���N�z8T�K��`�`��|DA�g���Ē��F���B(l{`�9���-�J���ON���O��$:�'�?)�!�!R>����r!����*�?��i��H��'4�b����];>s�(R$�`*�i�(5h,0bf�o�(C�4/��
m�LSC�h�P�Sh�]x�������T�������������C�����D�OR���O�$�O��$����`"LB"x����`˓x���c�5p�2�'�����'�B`sTg]�aB�i�&�	h@F󱃥>��?!J>�|����3HN�p�ƥ�Ւ�m��0��H���~~��&w0t��)}�'u�	,n�n�tC�;$��Da�H��	����	ԟ��i>��'&6-�v%f�D_?` T`wGs'x���_5d���Ʀ��?�PQ��9۴^כ����8E�J�m.	�"�Ń	
�8�U�*C4�7�|�@�	G��1Q��O�\�'J���w�$D�d!�9T�@0��Qª�9�'��'�r�'�"�'u�Ԙ�B�� |�ڜ��-�q��,�O��$�OxmZ���'�T6m'�DI/g� �x`��_d̠�5��ِ�&��S۴m�f�O��C�i����O��2f�?z�tթ"��l�D���_b_���-rƒO��?����?����
�;�f�Ni �k�e�<Z�f�����?�.O�mo�=#U�A�	�����o��l�8��cV�P7j��ږ�߾���b}���܈oZ����|��'%������ Y@���<U퀭�S��UD⅁b�7������@�ғO��M6n[҄P6� �?�΀�2A�O����O8�D�O1��ʓ��&ܖs�$:�$�68(��2��� ��,0W�'N�Hz�⟐��O.�mZ������þ0����&k�vl���ٴ^���B9ߛ6���`��2���kyy�ň�v'��y`�6 q���5�yRR����͟X��ܟ0��ݟ��O�xe�F�P�P��dITB#[�8�+ rӈy���O��d�O`�����HĦ�%��p˖ʗ&B�-��h0e��i[�4؛��0��	)��6�g�T����	h�s$P�x钕�j�� !A/<Nb.J�Iny��'C�� s$�u��7I�|��Eѷ.6��'���'q��MSr�����Op�y�b��ɠӀַ4F�h*��7�����dMæ����ē:��MR ��-gQ��k���V4�'̢���Y 8 (ғ�te�ܟ(B�'a�[i��^vJh��+��'(�Qp�'��'��'O�>���/#�zu3V!�@Ɯa��B�Z���	%�M#QE�3�?���
K�v�4�Ҩ���¼c�� ��B�Pfh�31Oj�o��?�ش4	�-��4���Prd��'҅Z@���F��|�!�R�LJ� �4�D�<	���?����?A��?�֡�$a�C���0�F���F�-��D���!qj�֟��I̟<'?��	u�����!�%*q��"O�
$R�:�O���{�$%���ٟ��V��� x�J�-ȂK�l��oGr�0����ʓ5�5��$�OP J>�+OJ4yaO��.����C��	�ֵ�BH�O����O����O�ɵ<��i��(t�'��+����u�D��XxR�AQ�'�P7-�O\�Ol��'"�'��Y'�4L��)J�6��ds�7]��i���Of�bܴdX���"?������"cĿv�$�Ц*��:��p�Ԯ��<a���?q���?!���?	���&òq���C&�RG�rec�"n��'�`o�L�p3���W��5$�<��K�-�N����Z�%[�kґ�ē�?I��|"�����M��O�H�	��.���2�i�!P6����J1v�!���T�$�O���|B���?y�<�(=���W�>n�����$�my��?i*O,oڽ����ҟ4��R����{�q�LCɐd�Q<��d�E}b�qӴ�nڇ��S�d�8P��mâǧv\� jt&��బi��6�z@*Q��S�;��DW�	!%Q�]�"g]G�\�+�+{�0|�I�����Οd�)��Cy��lӬ��V�̤BT*UE֎Xi��;����@T��
6�����NyB�iG.Y0@f�%r��
!c��3��Pp�r�� nr<n�k~��r���S�3M�	6s$�%;��Y�"�D� ��8���ry�'j��'�r�'
bT>�椕(k���;��C�6�A�qd�<�M��Dۿ�?���?����cf���/7g�8���$`��y��&�,U��nڳ�M�2�x����G4ٛ�9O<��D�]��$��퉍O�TH�2O�ɐ�H#�?�� ��<!��?I��D>.lµ 7�@64�89�׆� �?9���?�����Ц�SE\y�'�2�C�?��EfC�%� �H���Fc}B�i��o���?�d
_D�xaX�X& �o8?���G�F@^�P6����'TDL�$ނ�?��a�	J�͸M.E�P���<�?Q���?���?a����O��1DHD�YUH�
�N?L\��Վ�O�Dl5Q`ٕ'��6-�i�mk1J�,ɘXC&J֕D�8��z����͟|�ٴ ˰�
�4���%"V��'V4�Xd�ԑ��$�L�V@�]X�k3���<ͧ�?)���?����?�aᒮ?���;�a�w���h�T���Uͦ}z��˟���ܟ�'?�ɠ*. ����E�2�[��B !X��*O�Dq�%���^�I��ؔ�����Q���ERsW�M��LaP��l�㞪�2�HX�	kyB� :UW���(�>���17掖w���'���'~�Ow��<�?q������x��Ũ9�PЙ��M>b�E�ȟ�۴��'��ꓜ?����6o�7s��Ũ磐*$��!���}FP(�i=�I�W	�K��O>q���T�}F������|���
��Y�o��D�O���O����O�<�8	aP��ʘ~Ru��O�R�ލ��ٟ����?�p�}>��I2�M�H>96�֏`n<�R��i��I�V�^�gB�'�7٦�ӵW�]lW~Bl����-�RB�����+�F=����0Qa�|�X�������8���ʐ5� A;�i��q;��ӧ�����	sy�Dj��bRe�<����򩈤��H�ć�F���m.*������d�O
��d�)"T,Z.���H�j2?��E�cV�C�EP��{������͟,�|B��5R)���#��3slɪd�Y*�R�'��'Z��R���ܴJ7&=C�I��[,E+GK� &�L-I4�3��H��?qG[��o�;G���C�NG�z4-C��B`�r�{���M��@)�M��O�%��c�=�d��<��i4icА;��P�B��=<L%���$�Op�D�O*��O����|r�`��Px��h�d�y:U���,"!�V��5i��'RB����'� 6=��eCRÉ}��ZA��h���*��a1���S�'5���۴�yb��,r@�+���-ԑ�pa��y�bE����^�'A��ן��ɉty�d����*d���aE�Z�������Iɟ�'�87mˆ@HB�d�Oh��q��0�Pϛ�)C`��P��x��O4m���?�N<9W�^gYz����HR��� �����
2#&��ϋ;^��:��;���%M����v-��%"*�� \� ����Of���OF��7ڧ�?�@� S�Bhk��:%W��3�$�$�?)��i�>QS��'$2+o���杞~��R׌70�T���Aܻ,b�特�M��'P��IU�e��V����rB\9-h��K^>�Bb��L0$�D��/i]��$�0�'-��'�2�'�"0O&��Q�dr:c�ڟ�R-��T����4+o�q���?����䧥?���R:y(�� fs5N��m��l��矘�����S�'S���7O$���K�p�,M�D�%��p�'����ß�ᔔ|�^�(5I�	�
�I��E:���p��'K��'�R���DQ�h:ݴ"ﶼ��qv>̓��XPP
Pˌ�;�z!�jf�F���Z}�'�r�'�r(�dF�=	� Q�cBWzp4%A@Ñ�X���=O��D����x��~�	�?����l��v�[.-����㙂"R��I�� ��Ο��	ğ0�Iy�'w�����$)$Þ=��b����I��l�	џH+شE���s/O�9oZv�I:o--��C�+�.�+#NV1rT��'����ϟ\��>_Ԛ�m��<)��u��8r �L7�T���"%2-9�D����Ծ����4�$�D�O@��H�Tl�h8�,ʚ|��|���B�2��Oʓ2t��P�6Z��'r2R>𐫀c��4�Q;'����5?	�Y���I��%���ϟ� �Y�v���f�ZY;6�T6�,E@���B� S�j��f����?�	��'�V�&�X�ᩆ�T�q��H:K�&D���L�	ޟ4���b>Y�'� 6�!%���`r
1O�lhs��0R���3�J�<���i��Ot�'�B�L?,��e�g�I�m�D-��"t2�'�~@�i��I�r��IrB�O�!<�����7�|R�d�����d�OT�d�O��d�O����|J�jͣ'Ep����	,Y�@y#'�a���	�7B�'c����'��6=�d{���./"`�SJ d4�!c�+�O�� ��	I�946�n�\s�D�J�@<9s%��J2(a��u�|���3R��RF��Vy�O�2!�B��$g��'�)Ӎ	}4��'q��'��ɸ�M���
�?����?�D΁18�T��o��" �C�d	7��'���(��ӎX$��zN]�P!6Oͱ	���#M ?�BL�C�"�����'S��D�2�?Q+Z�ځ
"`~�a��?9��?i���?9��i�O>��1�T�)�^PX�	9m����k�O�En�%8��(�'��7�=�i�997��B�� �4k�<4�|�cLc���	�����!CC�n{~b&�4���Sܔ\ɤ�@,b,�,P)֣ ��(rѝ|bY��џ��	����p��֗5�Z9*B�A�<�%�v�eyB,m�Jp��m�O �d�O��󤍮AZ����P? �Nd@�K�P[���'�r�'�ɧ�O�x�#Ù�,5N���̈&J` ��A�%����O���t� �?��&���<!�*��p�v�06_	O	U���I��?��?����?�'��d_ɦ�i1��� ƶ:�NQ�@NC�`�X봬r���۴��'����?���?9��̘����dȎ<�7��%)j�%�޴��$ހW�f�@�'��O����n�zV�Y�Q�(*�@۔�y"�'���';B�'����P��B�(4_�E��ǋ�bc��
a��O����O>Xm:mM��'a87�"�d�CZ�d(�σi^و���w�|��'��O.f���i��I ^״HJC�.4l~E*K�=�~�0D�	 4ab�D�ay�O�r�'��cXu�m�G�",u��8����)��'S�I�MK��պ��$�O�ʧT�޵��X�?�4X�U�Hi[Tn!?�V_�h�Iڟ|�O<�O�4 r�F�v�b�#�:9���WH�4GZ�	�a�*��4���+��RD|�O����E��F�>�h�L]"l�H�OR��O��D�O1��ʓ����,Z!��
:�X�����=����W���4��'�X듄?Q��_
J��iF+ە�:M��.��?��h]2��޴��D�+TE�������=$���Z� �xd��n�L���iy��'���'���' 2[>)PӈG	։��`Q3b�� ��$�Mf)���?q��?H~z�u���w@�Y�c�
��8�#��(x��xY�'�B�,��)��,��6mp��q�d�&�1[�͌$��b�t`Bd��D�r-i�	vy�OBr
Q'�*�K���b�!0��֕�b�'Sr�'��	��M[��J1�?���?!Q�������P33O�� EFC+Z��)�h}�`wӎ=o����x�C/L�	��A�B��͓�?�`@ې?����+��$�����C�6�$י��(B��r@ǯ+i�!�ēL���S�)6:�y���Kx$���Ҧ���gyB�c�l�杇�2����G�D���{�����	��M���i�7�_�
�7-z���I;FQ2,{A�O�2x)"B��3�r�3!�!T�����D�ay"�	8`t�b�'MA�X�tG�Uަ�k��fN��B���|�R���5�>���R�	@�bb�&0�����M˳�iPJO1����f��\Q��Ն��::�0��G<}�M��ɲ<�� ��-4��W��䓬��R�z���1�敧`�Ab6�Iefa|b�w��0�t��Oڌ* Ή�5�x�б��8P.�;S6OНn�O�!��I��M[%�io@7MF�8x�!	�n'8�08sӨ�O/,1@6fe�B�Ax.����\�{I~���v��c�پ4���� �M+z����?����E�J�H��
s\H ��/�����O^�m��2!��Qכƚ|�I�|�$4C��(�1��i�>��OЄo��M�'z�ιK۴������P#����B��E����Pڑ�؏�?Q�=���<i�ZE	:���⇙Cc(�Š܆|(�"<�R�i�*e�$R�,�	F�d��=`��<��C�8d0��8��D�Dy��'����)�T>�Z���EEڔOs.�tS�#F�E�����`ۑM�D����������і|��8i���S�);6�R�ccB�:�x�
aӰ@勍l���U�W�@Q�,� 'U����O6�l�U��X-�Ʀs�MO=
� ��D1
KfĲҠ�0�M�g�i/�)!�i��I<�� 0�ODf�'���S�1ng2`S`�ϣ&�� c�'��Q��:��K.|D�򠝥yL0����_��M�S����$�O�?]�����A7�M�%�G�	h��c��%Q��"~�h�%�b>�k��զ��%k�F��,�:s!�PN�J�ɁŠً��'*��%�ܗ'p�	�=�u���<|m�""AH�nBZ�����	B��,�IퟄZ�� z���ȏ�N�vĊP�Si���	��M#a�i<>O� ^�#P1I� ��E�0>͚U���A��K�p�F�ūQY��r�2��˟�ò*�({�t������@�zB�.D������2{�Ƒ�acU�#v�IQ�����4
�̨)Odl`�Ӽ��f��3�|�j�dɜ�,�z��C�<9�iM�6������'L��	�'+�yXŦW�?�Q��S$.�ʄ&�*k����C���'h����Iҟ��ǟ��I�Lj<�c*O�x6����s��'�7�&[�4���O��4�9OjE�B�ʅ��@�t��7��Ȓq�g}��'2�|��� �)�\�K���VWЀ�&��P~�%a1����B+���c�uA8�O�ʓހH��u�1䥃�}��1@��?����?���|*(O��mZ�L���Id,(p�#;T��u3B�k��	��MS�b��>����?I�\�(Q͐�3�j,����9@��H
XRpXo�c~"�[
I��E�cܧݿ��@	63#�4:M,5�8{���<9��?I��?���?!����T|��AB�2N2��0c�4i^�'8Bgz����5��<��ix�'U�p�vL�s��0�l�_Hf��|��'(�O�(�{�in��0�*����1���$)MT�J����W%"�/ZX��ey�O��'�r��9@@=���W3*���;� U���'o剖�M���V �?A��?�(����r�N��^t�bm��h`:�����O(hnZ��M���xʟ�	SoĞ3�t%���-o>���@�4���i�L"k4���|�C��O��pH>Yы�,rR�C
^�<v��¬�?���?����?�|�+O�Dn�+�ƸY#Ϛ�q҈ز�O	�8�xHL[ya{ӆ��.O�7��1�f�yC�˿'8li�Q�`�mZ��M#k̛�M;�On�9S��>��<#bV�P�D���=H�i��C��<-O"�$�O����O����O�˧M+$�z��l����FK�Ĉv�i���p_� ��g�'F��w��X���J�:C� +v�@�x�(oZ"��ŞdGĩX�4�yb˜�*� `��)әKhંA��yR 4��MX7a��#(�0T�҇����r�ށ�H�q�I�p�H��2���Y��	�i�,!����BM5���SE�_����@c�'$xDb�j��j8��+����TY�跅H6����(1�sPU��[W� M��t@�@�RW�Q`��J�� P0�+ON�"�I��@O0��p�B��,}b��4%�
m�a��٬
H��(��t'�����L���J@��� � 	  M�W�&B�Z�Ȓ�(�R��Km��8���)�Ρi(L6^aJ����C)�1��ie��'��Iz��+L��X��E[�5h�%�!j�<�d0�d�O>��Q�ݱOf����H$VѸ�,�9j�<%���i���'V�I]��aட����OR�	ڷ_ؚp���C�ɺ�됦\9^�'����៸b"�S�����͊C�I�C��D_��� �MS)O�����ݦ��˟L���?Ѡ�Ok�ÀD-|�C��&({lL��J�?؛��'I��^��O��>�fUE�ҵ�+��v��$�6G{�`t�(����������	�?K�O�˓,�Ƀt�޻#x1��c_����S�i3�l�f�d2��֟�: bЪؾ�uդ	�Fh:�DU��M{���?��9q�*\��'�b�O&4����+��X�` H.��C���F/1��O\��O^�DD{ޠ:'��*��u%��^��4mZ�����AZ��d�<!�����2嚾f\@�`!;���(��f}hÕ��'�b�'�2_��bЦ�P��:�o1|�����@ ��O���?YN>���?v�E?B��P��R�B�@1��m��U.���?���?Y-O���K�|��Q�����t"U�`�9@Ŧ5�'2�|"�'b��).�b چ�����B<V�hl��cJ!S���?	���?�,O�P�ժ�M���'���r�ߡIF�1k5"77̬ @�c�L��,���ON�D�&q�J�|�p�J�`�l��� ���d�#����d�O�}�hxUU?%�I�H��+��5��)�3Ve�i����oz��O<����?i�O�?��'��i��GN��҉�r�H�d�<E��S���b
��M[��?���"eS������㜔+@����H�:8�7-�Ox��G�S�
��/�d(�ip
�o��B^�"�.)��6M�d�oZΟ��	���������|�S���=a��j�d�.�f��)H�GR���s��'��	^��U�4�I�0Bn��#�[(|��#O��-��4�?	���?i@	��P�����' ��@**Z���Yj�,�b@���O���'R�	:b��x�����O��d�O�dPT!�,
�8�Je���f�w`�˦m�		l���L<�'�?AI>�6k��r�Y�Z}��*4N'c�֥`�Or-����Ob��?���?�-O�(����<&�H Q'Ńai�9���J-^�'�4���$�0��u��bANP�3@=7j<������M������?a*O����4��Ӡ+ot	���ͰXl��q�藕!�6��<i���',�7R|P7-K�_3<���k*6�28�"��6'�	���	ڟ4�'�,XHE�5��wp:(q���8r�w���?6��oZןt%�x�'N.���'��'X����lƄ$֨�fV ;K��o�����Zy�eH5t$d�b��k�%n<��oߢr6�d�4.�,�'��=����	F�V
s�������
 K|��������'EZ��C�t�H��OpR�O�H�=Ѿ�H1.�utԸ+sh��|���o���@���*lq����I�O��I�|n:� ��u�n{���B�3]�F� !�iM�Y���'n�'7��O��)�u���~ߜ˧��1yU�rANJ(D���)��E����y��iطGɚ�",+�ђdcоP[�<o�ޟL�����vJ�]yʟ��'�a2g��k��E �C�W_"�jGO"�I/ׂL�H|����?!��L沄(������\u�X7z���ire�kHhO���O����<!�@ލg�Ȩ����J8,IC���=���'�� ��'��'��'���7,Z�1p.�fc��)q�� ��a��ՠ�ē�?���?*O$�D�O���(L�'0�1�c�Hg$�s�L�D����9���O��Ĺ<�e�2)�)�2S���Yn�PAj�+̌\��������S��zy����҈�<s��|:���2o8$R�o�y���?����?)-O���B��G�S�?`�y���Z���!g�?u��t�۴�?�M>�,O��
���O��O�`�6ʑ.U�h�� �q�!ڴ�?���J�Q1�q'>)�	�?��{kr�
b(��X&Ol�H�0��<aW�¿�?YM~��OI.�w�X��h���1<%\��ش��dI�=�mZ�����O6��^~¤�NI�!�̔�MW<dق�́�M�+O�K$��OX�'>E%?7-�fr6�R�aٞPe�MhT�9P���?X�>6��O�D�O��G�i>=��i�97�����,�"Y|Љ�I��M��@��?9����<���PsO�;8K�u��g	���������M���?���&�|�)O�C�dԀH*p�Y�d��D������1����<�بm\��������2u�%u���BY.D��	|���d�r@ʓB���T�{��yb#5G_���Ť9;^��\��r�ϐY6b�x�IDy�'� xp�lķY�����Œu�^D2p�
�W��	џ ��]���?��'dnL"p��S��/���k�46�P$�'z��'5bU���������\��+�Q�R�t%���d�OJ��(�D�<1�C�?Q@�ӑ#��3��.'h%y�͋=��IП��ɟ�' ڬRC��~��#��`���B� ��6��K��E��iw�P�\��ȟ��I*s2��矄��>U'z�!�ޡ[�\�r�_��u�ܴ�?i���_;9����OR�'���J��_����f�Y&H><��3��A��ꓓ?���?�c�X�<y���?����4KE1n�J��H8D�6|!�����M�(O �äa��]�	Ɵ��	�?M �O�n�/P���w`ݢ`kd#2h[dq���'�b@��y�|"���&_f�M+C�ذEq��86(^;K]���.i֮7m�O����O���u}r\�2�nB�ڽ�$=�(��d���0�>����R�):�<1'B�,% �"�d�N U�i?B�'�/�� [L����O��	�-�rD3G��N�P<;�IP�$6�O�ʓl�:��S���'��ޟ�����ܢN��!�e"�>k��izR
U�$KJꓒ��O���?�1-
й���yѢ8 P�٫r�l��<�Át�����D��ҟ<��qyB�X��0u#S&�!`��&[�����>�(OF��<����?��t�$�1&љlx��Q*}0��P��<����?����?)����D�D �Y�'X����U�ͤ42H��3��\�n�]yR�'���ݟ��	�`c�>���M�J(��ʏa�2�ڑ��馵�	͟��	ПT�'Uh�
⋧~��6�de�כGzP��o�j�����i��Y�P�	֟��=	x��It�Ă�?1�xb�������h�q���'�Q��4��%��I�O��D����X�c�-8\�=X�@=  B�qELJ}r�'�'��q��'�bP���'O8)�D�RS��S֬+gb�lZGy�+�'f��6-�O*�$�O
��
S}Zwy CRI���,����Ȧ�ٴ�?Y�<� ��4�����}���[�C��D�6IКɐ6��˦�Z"mX�M���?y��ʖZ�4�'�j��c�.��Pj����m���i��P��3O��Ļ<�����'{!�oN�J�v`��!&&��ݱ��f�j���O6�$��w��$�x�	����ȼEG�iaw��U�����d�&�O�xI7O��ȟ��I؟\�LY+Q|�p�C3$�x�bK�/�MK����y���x��'RB�|Zc�(U֛z�P�� )&&�A�Od!�?OB˓�?����?-OD�Y���-3㠔�E0��ԥʺ�&����0%���� q`!�o�e�v��-Z��,��G�=GXR�	gy��'���'��ɦ~5�yh�O���Sfk��d 
cІ� ����O~���O��O|���O�M�O�)�g�}�XQ*kۀ6�4�u��g}��'��'�	)�b� H|��a��Z2���]�i���	�"[�f�'S�'�r�'��}�!�'@�H1�����4�Bc[=�| kme� ���Ojʓ���P��D�'��$��*wV��q�`�c<X`*��GEBOz���O`�Q5��O�O���+�n�1R��2�R���m 46�<a�KI����B�~
��z������ß���(b���
_)3�{Ӕ���O
@�0O��O��>��_8?�%��
�CY0�Ġ|�T�A�'�����	֟ ���?��N<i��u�b��raǺu'P��0�Qf�,|K��i�Ҧ���|�(O��D�7+V ɶ �K^�A�	��0)�\n�ğ��	��`"� E,�ē�?���~� }�T�i ��)pq2��̸�M+L>q�+^�p��O��'�H?� �� P�Sv��9��iǢe�ҹi�f2>Vb�<��C�i�����z�
 �0)�8�v����>1DOV��?	-O����O��<�T��;W��b���$��RV��$C)Ҹ�G�x��'�ў��%PuT����"�C�>`e�� D���H�Iߟ<����ty"�T�*��S�B��Y�P��J��҅m��u����?ъ�d�O�0��k�OZ��3�_ ajDx�)H�_�$�y���S}��'k2�'V�I�7�0�2�����_e�5�
�a�"`���Q�>em���L�'���'����yB�>ɗ'��x�XT�r�t���V٦��I矄�'�l�����~R���y��h4�����=��P�`B0.��"QV�����t�I#���	^��''�	�"-�ΰz_qV`p3��,6�*�n�VyEԴHab7��O����O��)�l}Zw�b< ��"S��l���E��
�4�?I�@Fx���֟>&kd̅���(C
�=���a��cO�7��O��d�OH��q}RV�)��?:@HS���& 1b����F�MK�I��<������?��؟H�C�"�*�k���oƞ!�E��0�M��?i�'�U�1V���'���O����l�' �@�X�L�d9�!��i9�IƟ,2� |��'�?���?��LQ�<K��+)C ,�q�*�3���'��1��>!)O8�d�<)��3�^�g�,�Sg�`i�=�4K�B}bK��y��'@��'���'��	%ez�Q���`�ذ�i�4<�&*��G�����<����O��d�O\���B�p���C��o�RMiQK�,p��$�O��d�O���O ʓ�-��;�R<��kI�t�J�R�>9e;�i������'��'���y��W�5� +�O
6y�؈�)��lʶ��?����?Y.O:�2��[��'�8�U�O3�$�Kw+~���Q�z�(�Ĺ<���?��SK���>YĪ��6�XU�@�y���;����E�I�ė'�JykU��~���?I��6��,B�Ծ.V�ʱ�C
]�(��\�0�	Ο����q�8�'���?1�"M3T�栁��ȦF�eB
wӦ�8*0bQ�i���'���OԌ�Ӻ�`Hɹ�,l;�/ԁ岥� ��-��ş�xw�{���IRy"��ެq̞,sF��-J=)��ܵD����S0en7��O�q���m}RX�`c�bA7p`\(�pCF�y5F��d�,�M+&��<A-O@��;�S��'��qMy�1LG�x��ȸ�Σ�M���?��'dnĹc\�x�'SB�OMh�ғX���Q��=���Q\�̖'&��O�	�O4��O���o�.l�p�Z�2y�f�\�R,^7��O�I E�f��������\��5I<% �b#� �E�k��I7��DqX1Od�D�O��D�<	qeǕ$����sh=�p�޻]��X�w�x��'��'���Ɵl�I#L��]�	ŶES�Ěr��8zxa�1�I��p�I��h�'r���a�}>5XU�{
D����/yD�+��>y���?������O���6����Z[J�[iԚs�\�B��xD��?���?!(O���a�NK�S��b�PVe9bȒ�Þ=�ʥyߴ�?������O���ޙr��>�R�
:p@V ��o��p�LJË�����GyR�'W( e�'*��'Mr�OD�1S5�+G��-(�ؤO�0��,���O �$Y�)�X$��T?m��n�.�)Ĥ��'.�#�cl��˓D�F8	'�i	��'�?���q�	�?P �Q�JK�Y@��!.˿2��7-�OP�$MG�b?92
�4~��E	�f�%C�x	 !�O����	\�|��O ; O �@ÆM[�%O2�yr)�2+�"���$R�iԼt�&x��^'L��L���G+3�.��8?5��bU��T�#jѶ`�v�SC�N%	%��nƟF˜���(	S��2�?.�N���M<�z@���K/X-C3l��Z��`i���G���r���:9�z���=n>�x��f)&��Ȣ3$G��R�'r�'�z���T���|����+,�J�V�Q徽+��V�T���S��7�q��V q���1��		�B�2̓�k�Ɋ�,�C�H��3͔�6�.�B���<9t	ɥ��UC/�{DRM'�H[/=dri)we�5\���H_��B�d�O$�=��!؃#��5X���K܈��`fh	��m����W#H*��Ezd�
�" ��<��U��'K�q�%kӌ���OVI��ի4�Q�S�1h��!�O~�D��`%$�D�O2���:xp�w��m�	:@G D�d�	(ywD���N~P��[�:E���X�8���2���UnB�G�0T�P`ڵ--�C��'(<B���?酷i���h��SO�,��)����;$������?E����[F�T��\	 �V`A���K�ў"~P�i�vت���ZG�xar�́*>��G�'副C�
� �O8�Ģ|2aO�8�?a$+��y?��%�Rq�!��P�?���Y2��X�Oi@�����~X*�z˧��`%�T�0'��q�� �O�邆�;��)��$>��"}"u�!.*�J�O�M� (��u��^�4�r�'��>���0�(4!�,�?=4���L_�4H�C�I5��Ջ^�]�@��3�G(o�.��ĂW�'\���+� `��P���&x���>	���?q
!~��t@��?q��?�;0v��p/�cي����SJq gC�=���@��'0d�p�gə����S�? ؼ���)4����`��^���h@K�T�х��x���y�q��'ǚ��D�s�"�BPeZ{(�E�W�'�	57��4���=	����Un�/d���#�G�!�E�U�T$(4m��� :�K%UI�	��HO�Py���={�����C6窭Z�nC Lf0�b�d%-�"�'�b�'���������|B�S�c�r��0j��*���W�%~�B�/�:��͢QK���<���1aP��u���	��ڸj�T�i�0]P#����<QՃ��[V��ԧH�*�vER�ˊJ��X�	���E{��D�y�`�z'F'N��`��@�jO!�&09ba�!�����3�d�471Oj��'��I�M�D���4�?��h��x f
�z�nM�VG�
��+���?i�
Ȥ�?�����$�G�tϛf�$T�B���7�ߢ?��r� *�p<E�9L� �Y�I�4����
cO�(h��B�%p��!�%~��x���?)��i�*7��OUpֳT��g�0]3�p� A
���۟��?E�4��F������;*-feI��7�x�aj�`a饌F�uJH �%��,�h��2O��p�`\r!D��?!����J�~,z�$øP�|�SN�#P��՚��+K(���O�,��� ��!�5%̣f"�裐hE���dY>Y�A�5	�F�
4F�*L@�Q�3�!}RL@)f�d۳aH�1X��t��l��>�'j�*2 B����U�W&e��2}ra�+�?)���?Y����O���4,�l AD�2{��Ĺ�\̓�?9
ϓ 0�%`W�ug�SG�Y#�A��I��HOf��UeL�_xt��&��f(O��D�O�����u�j�`���h�~����?�!�d�0&��84	�1�d�(I�V�!�d��1��1��I]�=�;GO�|�!��߶9��,l�B����	l�!�dH5O�0їOلy2 )��bE�p�!��o���b�J�e?~i�'�"�!��
z��0 ��
(Ă]k�a��t�!��B*0�東��	�5�M��ޡ(�!��7H1���h[�7����3�)=C!�dԼoPp�"p%��=�0�C煛<�!��߸^��ۧ��}�Z�"S�5Sc!�dF%S��["!T���
Ef�kP!�D�b����dN�:������F'<!�d�Lb���,�:}�J�C5!��"|�4�t��8i�2�ʷ��+!��5��y���)�~���!��m�!���v��y{�o�@#"�y�!��� f���.N�f L�k�,o!��Jz��e���04�����/�1W�!�6����!΍�P�����N�!��"�ft�Xh�z�m�*J�Xy*�"O���o�1,jU��B;/l-�"O����	�`|�E���!g�YHg"O*؉�@�zʀe�dG 7fx��"O*uu�TKf<��ĉT:��"O�E������*5o�?8�Ait"O<d� �Р�xa�N�&T�UK�"OR�
�7�'��"��=���ȓO7�YWN�_��Y�/�_Nq��C�R �tI�5`UPn;C�V���UqWϓ�5yj�a��=Qi����Dݲ�C#2��ٷ+� ax�ȓi��h񉅱!,(5�GNP�BO������1S&Ӻn��	�lC�a#rЄ�7@��P�ђc��J� �ޤ�ȓF �z1�f�	c�D]\ค�	�(������ր��^���ȓ&U<XxE�хQ�2�lS�[O��X�|��ԫJ=wn��ي&�����?86����5���0��_�@�m�ȓjr@��D� 	_x�V�lβ��a2��R@�$b��Q"i�mT�|��S�? �t�@�x��I��f�f�ة��"O����^�!(��Z��=a�"OTL�r,�-�H�Dm�"t�Z��w"O��u��:��ĸs�
�f�x2"O2�褨���9��˜�k��ͨe"O�ݸw�ШV���!ԫ�&�|m[�"O�,#��`����,9���"O %��e�"��M*C
ՀR$Np�G"O�1��
�ih�]HƂ81�	�"OV�[%�	%3>�-�֠��L�HS"O2�b��>�`�� Aԝ���B"O^P`So˪f����'��=V���"O;P	/�f=A�y>���"O\���X�,�V�4\��"O��
�ƕ?_n�P�6&��`��"O&�#I�em�ӁC�Boڡ���8�l��)��������#?1�RuV��!��VI��"	ftZ��'\�D*D�>0�>E�$L>h[���u']+2���Y���(�yR�V���� h<"�r`JO����|Lx�h
דj��!��|���� &�= �A��	pX�УnW<��h�H��K|nE����4-!�D�eƺe�B�ܢj���a@�p�Q�L�Z���'�����;JP�x���2Y[���$�I,1��ㄅ.�O�m�4쏮g�r�1��R��to���:&,��'���$&���,k� /ah�U��S�j�Ѷ"O�c���������K�X��^�t2�O��M��]�5��H?��cʁ[z�X�!����D���4�O�XsE��-C�5zC�	�����×<���(�$:}��+q���њ��{R*	AM�H�Bϗ!{��r-�
�0<)�E�j�	�VA (
1�N�$U�yR�����SEĪ��$	��'0QAJ�P������!H�\9��D+R�
�k��M���+��f��,tnz�BƏQ�c��Є#S@�<��˽uF��jN,5�LЗ+@y��^�=��`R�A^�ِw��x�OC�h�C��*�lQ�w� 2R�k�'�4�s���
UI�`��5��r��)s�� ��M#"��fD�c�nU*�1�6��	�'��M��ώ� q�1���5����?���GȜ�%Ϯ RE��!|&h2������8���s�	��9���J��}��=s�e� ��<��Mw#�X℈_�<o��s�cK~��r������0V����fT6�?��&�-"��ɫZ��K*��p�$܃{�L�x�Ol����K$8�@1bK�5kc�m����E�gh4c6���T�����SX�v�I��?Ac5��$�`�Ʌj�*E3 �`[�u;#O�%���JjY�R!N{�6s����YX�33��%	UbT��l�G�xX��S�jX�V)^%;6�O����J�(��Y��ͭtpް2u�'J D#�-�(0�n6�ל7���9��űIՄi(B�z��Q�E��(�G�'Q�L��.\�WZ����-`̍��zm�I�BeH==�����(�McF�m޸-릯��~��O�iP']� ���Ļm��ʣI*H��!�7N�=lB�#��T"���!�޼�D�Ҽ�8�E'Z%F�x9" ��O.�i%㱟0��!�?!�yעٵ�b 9sW��X��p=��OL�@�ċE�&WF�cND! e�!�f� 8�:Q;�e$}"�>f�Q���H�)��!�@�w?Y`A�3-Fʉ��#�@ેe�M��4d���A�d=�f��� �t�H!D>zYXdIדw����F$��}�v-�<�	�(�T�CF��/g@���*ߣ7j��>AƥNhN2�� ��U�
��U ����b,�L2�a[�A� �N�A­^?(�2�<�4���[w�0�dt����g`����8�q�'e�h��M+e9uj'���he�UF��2 ʔ�Pe�@#�rb�!�٫\i�m5A�/J�>���L����$�����	(9O^̐��ϥ�$�����DW�l�'2ړ�$��w��Ic` 35��[@��[�P(�竞�*)D�k$,�!F��L�<i�$��m� ��>>�Ȩ�JD�B�`��	P)�g�� �(���C��6m���æy���t�a��
Ɔ-"1{�(�c:����h @y��8^��q"kP/:�M�
��!����g��#����0�ř�l؇6�P�Y4���_�\!�II�iH����V>�5��Vy6�td�!DhԢ�G@#�@ b��'�@�X���'E<�i����~m`��B^7#�nDAfEذ�x�0>�
�+!M��P�e��m۶���@���D�	>��l�6�O� ��;���� �L2��ُa�bT �cƤm;Fݺ��'O~!�	^�&l�5�ƥ_�&��ED�vA�Ӯ�Q��y�F%
��t���6�����#\O P��d�9Zf�h􁔡w�x3���H��	o��bL$*���9C��O�Y�,�f'��'݊�x�L]�i(�0HA�<�dʝ�/���	b��a�v0�'#&�H��H�`fH0�4F��a�O���n?ͻU������8'fd:�^ h�2X�j@PH "��p	��r�@ߧP<4���d≞!xi#����H��qOPh�a�%u8dr�d�|Ҙ#p�'�J�Kg��1T�t�+V,X8-w*0/�괄�d�Z�"E��	�9�p����&F�P5
�I��Z+0� �N��t�Do(� C<��-O-�M�͜�W2�*����'�B�ɖ1�������>OX`�ƞ�a\�ɟʈq�}��I��p]��3�Bɠ\"��*�K�:
�!��4#�P�C$H�n?�Ȁ�U�i[�']~E�ۓk�JX�tQ�"�b��" ]�?�T���\�4��%d�����SZ8�ȓ2��l�5C]4%�����-�Q�|X�ȓS����WOJ�l�Xa"����7��ȓ�R��Ƃ�i�.t2�؋C z<�ȓw�rYct�E���)��K>G�p���pr�=�@DP�sd1Y���:Xԕ�ȓs�#2�ˡS�D�xᅔ6/�@��	]�QH��s��<��(SN{��������6��N��q�#wd��ȓ~��=���|D��&]�l�=���^��7��3 ^ցӱ���kvrA��WD��K �)?������Y����ȓ,D�eK�,�0�UA�"킼�ȓ�d Fd==(��¢ ���2�E��m�
��t�IV冼��77�Qk�@��D �� �4 BD�ȓ|�|:���<c{��kLk0^ �ȓ'f�$WL�u"͠��#oy�ȓ$@��J󬝊*��7鑤]�����*��bb��'��	��^�m�y�ȓk0�8E�C�<h�%X�EV8�`���f��	����e(�I^�s������\4���]�(�k��Ŝ!�X��%Zm���8� q���t6p��ȓK�ʠ�Z9:����7/�.jj5�ȓ7�Y�dǓ�?x<��DA�ІȓM�B��1�H�|�I�� ����MC�LidBɬY����t��9aD��ȓm|h�U�
~��Y+�ݹ[� ��s�p!����lk�Ặ�ŲI��e��|8�����S-ظ"��+PZ��E6( �Ƃ��>-��� �8�J}�ȓX^Qs!�*�\�a��ρ.�|�ȓ*t��	���Iy@E��r��ȓ+䘀l��]��9��Խ3�̠�ȓJ������R74$I���0����7�y#���m�6�	�wР���R6N(�R�W�r����-Z�^X&]��lC������D��@��OP�hF4��3Y��&�'H7�H3�����ȓ!��Y��<젷��*N!���k#�\��L2NE��͟{���ȓ
�z�B釓?\�hi�����a�ȓ(T���`B�|��Y&aC*
X�ȓw��q��-ϒV;P��@b��;𚕆ȓOG]��پ����gD�'!�����𐨧�O~�!x�h׎
���ȓa�E+��  <d	�E|��Մ�xȘ�갋9C݆e9d&�4,X�y��S�? �5Q�.O�ر3��AF궽H�"O�U���e$^9���=P�p�w"O���� �8y@�"T4��4a�"O�ap��-sF�zR�_?<Ă�"O�M��-D J���H�A��^�F�ʂ"O����&R��z�h0�J���"OM�P`@z"�(I5OU�b$�G"OB��V.�\�F����
�-�@"O�Ĺ��.+����n6_f���"O ��Ĭ�8_���U�fMx�kR"O|��A��}tb�@V�B�@�u+�"O�X'���н9��<t^��t"OrX���V�/~��� �ư]el���"OR3#H����e*SH䅰"O	 �FL#.��a���l�ТD"O6ǂ �	��| ƬP�"O(A��NY`@�i;_�P�{u"O|��I�p�HdP!V�H��"O@�����+��(A�"PRA@`�<I�)׻R����raפ{ | �p��\�<�����b���-R�*e|XQ��V�<�D
�I�81ٓ��)�@�2�
�{�<��(�'~|ز,T"<@"çGt�<����k�\MPӠ��T��
FY�<�F��X��=P��-y�x!��R�<9a��x� �2
A* p��R#�b�<�"���3�\��bݩkY$�3�Pj�<	W�D,h���{�jZ�=�`��φf�<!g(±C�vɣCeU$(Zd�WDh�<ɡ ��U����� ^�8PI!�g�<����9���Cb�DE�bY�6)�K�<Q�f�+R�z��fl�m�0@x��K�<�ć3D�.Õ�̝r*�X��/�]�<�cEJ�S��[���j���t�<��E7bfP�2��
M=���&�{�<�a��,+X4 w�z��4r�%m�<�W�B�x
Y�F�}G6d���X@�<� È@x��*��C�vְ�ҍWw�<��Z�q�"��x�mr���u�<Ƀ�ޒ2r�90"jȭ
����#I�W�<$���&���M�{(*�)T��T�<G�F(C\�`I�f�~�Li;��^F�<����.X1C�Uy5@ ��B�<�%��YG�	��
�(��T�áEz�<���Zt����#iU6�ġ]`�<��(��"����-^6�� -Y�<!��U�wB�!�9{(�k��`�<���N'U�I�(��2+l4�SC�<�@��-���y�
	h�0tf�~�<�b�4u hA���;NqL\��"`�<�IȮKN8��sa�[#�ث��-D����f	��8���g	|d��++D��2�m!h%=�5�ۃoth:��)D�<��7md)*��ÑP�j�I�N)D�,Җ@�6>��7a�S}.(��(D�Ԑ�S�i����T��9a���0e%D����L>�L�j�#� �ʕA��"D�l�ë�*z�H����V;|�fX�!?D���C4�2@u� /��p*N D���0en$i�e���	��J�*D����� ��b7�O�U](I�)�O���N44QB��$ p�$�F��(~m*B�	�W`�:�3|ʰhZG
��8�RB�ɹO,�hC��" ݔ|kf�Q�x�RB�)� DP��� �R� � _/wX�x�"O\���k�PZR�HS��&��XjF"O6�1���,kq���kn���"O.`Z ����+��ӛnf +�"O�Bɚ�Y:)P*7��$(7"O���� �dM��7q�%S"O�D��S�_]n��d�4�d A"Oh,�b��J&v���_u�Q�"Oz�Ae�p�kĎ;0GNh�"O�ݻ���"�R���i=�V"O��B���xh���F��#w �k�"O��8U�
L�ʉ�`\�s��)��"O�	��m8x���eW�R��"O�)�7䔾+����e�$nq:#e"O��mɕzg�X �WHn%��"O|�9���]H�c֥Etk�"Oy��2)bB�B�A	$rCL)��"OB�Ra�����"C�A�iB8(�A"O��I�ԁ(BW��,F9l�"O���$��mN*����G�΅�d"O~�G"��pIF=��L@(yfl���"O��8J]�}c.��t�â%W�D"O����i���(ѱG]=KK�DXu"Ol�A��ې
�^d���9.u3"O��UeĂl������ lH!"O�	�J2u�I��Z�%��y�"O>/�
K�)��&ԓ �,�"O�]��K�>�� �"k_�v8��0"O�lق�F�}�ۗ
�\`]�"O�(2C�
��m��۩i[8̳V"O,83Ae�+���ѦBPߪX7"O��$��9��QKuC6��}( "O���G"�%ULA�ł��*�Y�"O
)�p%�:b�B5"ą֬��"O\�Z���:�*�북��T3�pj�"O���g��!$7�	�%�7\0�yȡ"OX�y���x�樉vF��A-Vy�"O�h��yT+N@-z�Wy�!�d_`0��Db�o�lR� ��!�dʧ�\Q93��1i����@��G�!�$�.T�U *�Xc�nV�\w!��&pD���G�r��)8ጉ�g!�d]d?��W�8�!"B蒩 ���ȓ=#l5��皪y~ʕ���G�tP����1çfR�W�Bi�1n�+8l28�ȓR�p� Tf��A?0�˶�U3R�<чȓ
��L�W��8z��o	��t�ȓ^������g8pЭ�����ȓK��411������>M��ȓ'fP��ahM
T�:0��6�F��MS@L2O�<�V"�
�v9�b�Ph�<a-�j6��bn�]��凊O�<5+8��9B��!~7�1I%��d�<9�-����LQ�e�`N45���_�<q���'���Y��O�!��pR��`�'��?M�6��GJ�,٢B
�{3�Б� D��񧫍'P�p HSM�  �d�D��p����<Np�X��)M�~fLn���8���EN(w��6�͒E�ȓX��E���E��MA��A*	mJz	�'q�����k� �I�7|ژ��'8̝�P�6вY��c�=m.��k�'��@jt�C�u�
+�-�.nY$b�'���UaN5<��S�L Ĕ����� `�'��I)j�ye`ңP�����"O���eƵON<��f��<S�"O�hp!�ԀD&���Ϟ3����"O��ELNЕ(�6DyR�p"O� �@^.�`�!��+i\<��"O���/�[����$��6���"O��J������3.��v�@�P"O`y��'�,i��-��I�Y��"O�`:A.��_�ⅹ�k����=�"O��(s�7��m��/=���)�"O�̑2MH%RxP���]�#�0{�"OP4��L�g�FMK��=a���:�"O��(�jL�zp��d<IF ��"O������o��j�:J״u��"O�U"���b��;�b�m�J �3"ONu�ӢZ�BDkƣ�=}l�Ze"O���ܓj+��DH�s2H�"O
Y�R$݄�C�-�)s��)"O~���ĉ�eU���bl�i���V"O����烺#�1�� %�`�x�"O`E�#N�`=�L&�ۛ#��Ȼd"O���G�1��%���<�"%"O��`���2D4䁅�|��"b"O�:׊Oo��P;$�Оr���iC"O�I����E:4� f�/}|I�"O�PEI�\[�
����W"O��Ǉ8��<��B��.�}Q�"O(0��BܓW�P�xrg�R���"OƵ2gJ�L
���ЀA�� �"O��FM�z�:�F�V�6"O	��� ��|� ���44����W"O.Փ��+Oc�UP@$��.�����"O�Pp�B�H�Ќrb�O�_ctf"O؁�F�z!�T�fL��s��x��"Obu���zPZ���A�8a����e"O��o��ct8�0���?�ܘi�"O�415�I$�~�n>S����t"O���Ǫ��̠ g�{�ԩ�"Of�Sᔆ(�v�4,@�~��b3"O�����Ն4�P�YfO$_j�=;Щ�D�������+Xk����i,��A�I��yC��
�*�Bg�Rwx����ȅ�lu��ք�q�r�q��i��Y�ȓCa0��d9v�Y��Ƃ�Z���!fF!:"or+�u3dO�:��чȓ�	 b&έjh���H�h��ȓ�Cw���T����G�6]���'?ў�|bn?` ���J�HG�P4�NY�<iԉVq(Y�VÑ9� ��b��U�<���Ô}��R�2��x�/�S�<�q��/B�XhA@:Zb�kS��V�<�c���)@��k��u���hR�<���Ͼ������]�b�����#�G�<����,�Z�
e�χ5s�J�m�h�<��(C�N��Ա���Fy �z��I�<���C!� 劕�Y^t�p�nKA�<1�D/M��@��d�*���b��u�<�I��ODF\1�H߆�����F�r�<��JÔ[��P��x�l�4Ho�<A�b�,7`�y׃ �{Y6i+4˖j�<��Ĳj*��0�X�}�T+ �h�<� A,T��ȷ � #k�9��E	h�<����i���Ї�;(��8 �	g�<)p:\��i�1K�`���p�m�]�<� :A�h��8<���C@�q��LP�"O�%��e�2s`d�s��V��`���"Ob���dߞctFI�wF�!|�F	�"O�A��jO3eQ-�BK�x�8�B"Op A��:
�8D�  �,�S�"O$8�U��l�H��W7��Eɇ"Op�B�H_6,ڐ��WF&ŪP"O�Z���+ �h���8�0�"O���e�ц`����םCF�"Ox-���23�DM{��M2���"O�!Ss������u�PX��A0"O<9�E�Q�{��3e����0"OnM1�*��-��4��@ tp�"O��K�"�	>
8:�d+f��b�"O�uh��*�;0��0Ud,�"Ot��u �T\� 1&b�����"Ob)B��0 kz�q�K���	j�"O����:J��Q+�PVt)�"O�YBѯ^�2�����>jG�z�"O~d�&�9l
̴x LǤk4�	�"O�`b�P�^�Fɘ��D�B�
;o#!�D�#50L�E�E��yR�X
!�dZ��5��R���;� ^�{!����	�Ѡ�c�_}�*��>=�!�܇F 9#��YτY��i	�	�!�?
 n����6\!^�q�G�J�!��B>bL8!�� ��v��1�!�-5����d��-S�&�
��O�S�!�ė��]�mB�*�J��"N$<t!��_4
Y��U�ŵB ��P� �!򤛷)B�����*\��6Q0%�!�$\�>j��WFPbD|�b�'���!��#>z�!���'4ly{�L$Z�!򤜛2P�Q��+/��gϵ7	!�Ğ�)/��q�T�N�8���f���!�$�����J�!�'b�0�uH�;m!���:or\3��2���&��02�!�$O6�L��*�=+��E��f�!�;}�V(��`�ML�$S"��0!����bXh%��5R48t�T� 8!�䍹_p��*SF'���Ҭ1R!��4V�؍�M�=m����4��5:3!�]�^��iՃ:u�(BE�.?I!�D�0�Р���Xp2��s�@!�$C �=�!d�+%J +!霂E)!�d��#��0yR�%MI*�ôE��	!�D�X�^m����"�8R��(8�!��~���PjP(B(�g�!�dߨ	�\P����?�{Ĭ��i�!�D�\�X���i�\Yc+^�Dp!�AZ#� U.qߎ%�G+��FP!�D�)l��#J4ܦ�3�(M!�Xd[ziZ�e��rɌ���X-?=!�$]% P���cI��� j��-]%!���BI^ SӇͫv�Aœ~�!���)@Q�wױ��L@s�G^!�]D�&m�Sn�p�
�!%%�5A!�$mǮ19�H�,����7aY�R.!�ē2�Tx�ʓ�e���p��DG�!�D�>(�)8 �_�<����P\�!�Đ25B̙S��(s��y��I�S|!򤒂:ڂ��S�-TF���\�Ni!�ĉ�\���h���TOr�ˁ�<U{!򤇺!q�]��!��LL�X�&�*Z�!�� �"Fg�%/���0�b���,�p�"OJ$�Q!�n���P4�k��!�"O��J���9O��c1a@�j�A�D"O91���sI^��󯖮\p-
�"O �@���:N$$ٴdGxn�Cc"Oڌp�ό'd�|rg�:g���4"O>�XO�-�:�s�j�`1~�	2"OV	�7�ڇt�N]ȥ�!W$�Y�"OvTE�\�/0L�QSe�br��D"O`|�#�޷0�
��ccY�*�� y�"OT1Sb��%P]*t���Q}W�"�"O��B�ȕ#V� �������"OZ�H�"iʬ���3Iv���"OZj��M�-����`�]5p�("O$�5F;S~ܽ��&Wm��@bs"O��1����`r��re��!��Mp�"ORI���u�\4�s�� �P1��"OFh�&!߉6�PZ�/R�ݰ0"O
I�LU�B�!A@� ɲ�8!�DN'+��(юS�x"�y�`
�S!򤁧I&.�+��Ld涸9v��? !��%Tp2�k�� ٺ�xwe ^�!�Ā��zu+t"�- r�jG$�=Q�!�D�S�>T�@OH[x�3@ꊟD�!�$�r�@�3�8Y����(ʕ>l!�DT���H�mX+c�~9C2-��Y!��?V
��hdaJ<~��˵�I7P!�$��~F���A�V�3^���q��8?>!�d�{��E�D#T��I�b�!�ލ��QYg#޻*�&�3��+!�Ѯ7�D�z�H
� �zL;pGF!!
!��9�h�ɟ1�^��l��8�!�D�`(Àk�9d�,٠���!��ʒ$hT���ͧ3����u��m�!��N�Lu�q�F눂y���0��|q!���	m���KuA�fT(Æ�OjY!��ʕ?ϴu�&Z�&-������V�!�D���lL1�K}9����Z�!�D�.0%�Y+�g�+e��q�wn��Yy!��5�8=��B�Mɦ�	҇�,k!��)W̹����x���`&э~c!�d�*��kՀ�,>8��cFZ!�$O�8lJ�� M\��M�É�+{c!�DSO�J9AF�4Ր��r��6gG!��$z%�XP��$%�x\��Θa6!�dY����[�I i����E�$k4!���
M�.8�A�/"5*t�⎝�K�!��U�fA{ϡU�L8���T�+�!����bY�eFp��djs!��_�$�,e��^=O�H��cc�+B[!�$��A��� �cȗm̤���@��!�Dh�P!�fB$�e���Z�M!��H���`�u���2Ei��=e!�$A�5{��ʅ�Ȱ_	�i*6��aP!�D�,+,���FC_-9c�� r'!����d��Ek�%�t5���Si1!�$� ��}�#C�!߾�φ0!�P�1⤼äʞ��,���� c"!�URN�|���-�аM�7!�dF�3�$K�Ǿxn��4͏D!�$M�f�B�τ{kb8�f�X�!�D$]��$jBd�s0ɐ�-��C!��#U�@���h�d�CD̔�o�!�DG�yB��$nʝ�~�h�k�	�!�� "�J�G���Jv���|��L�'"O"���Y�a`6�f
WC��"Ol�·n�+ �:H����8�2�q`"O�hi�
��[f`�c�'Q	9�ri#e"O���F%�,n��U��Į;�nȳ�"Ox�%��*����!��v��q"O��W���T$
�V]eD��0"O�L�WB��4 ��)���"O(�@D숷ͼ����I�
��ur"OJ�ᰬ��L�\®�A�0ؐ"OH4���V@2x=�!�H$>��Y�"O�9`J�$����B+խs��aؑ"O0tc� �4 ʕ9!E��x�rS"O��P�$o�a@��7D�4Y"O�%�S��*'�~y��"M�R �"OT1ye��(L(�E�T�V��"O�tq$[2F��e��Wo��9�"O����=mT�2c��	Z4tЇ"ODe���&W튅�l]2<���2U"Oڔ�dGS�}�0M�Ş�Z���"O^B�#_�.>j,�g��1+�\Y�U"O�X"�G77�LS����]�Đ�A"Ob�qd)ɿJ���JF�-6���yR-$�l���� q&a;r*T�yb�5���s4�
�dt�|��G	�yҁX&�j��2�
���5:t��?�y���CTQ�e�m@
A�6�@��yB��k�I�/�k}�)��k
�y�E]�d{fEe�~�fc�+�y���-���e�aɸ�r�IW#�y��\fl��t�X�T����j��y�.�R/���P�=�j�R�H_��y�X5P��zr��6
�
]��y�
�S�)�E��%��;V���y","{I,\ѦcQB��)S���y��^HT(g������G�y"�LDa�@ a,���9�yb�EX��� ��1e��5���y2�X�"�x�(�&$��U���5�y��@�y6�
L�D��!�yB��#j)���O w��I�!��y�l�7���a突���Y����y�JL9L��\2�	�(H�B����y�i��g&���˨q�JԊ#�>�y���6�Ih ��*!�B��"F�"�y��Z�D_LYr�nѕw� ����y�\�{�xpX���$(��-B��y�/޾/�ơ����m�b�Ig
���yR�i�J  `H�b�J��	K+�yrP�US"�i�^\���w��y-ܪaY��� �)��,P�Z��y��ˤ4:�@�#.���2�ֲ��'J��?):�o���X �Ħf�j(@cJ'D��Д,�*���C��(YĎ�s��#D�H!�釯W>�ڵ�Е$�x���a#D����E\�4�0���B�Z��#�y�,�ak�셏~v@�J�T;�yRm1=߾蓤�nz�%j����yB� h��J�DS�m��q+�<�y�ň�RNFœt͏�3Q���DgY�y�o��.|C��
��L�)�%�ym_'�:Y�qӸ�8�)�� �y�f�
V���ڥ<�h�S��y�;p�`���E�5�xH0����y
� d$QƞP�j !!&̿E�ȉ�"O��S���O�bx[��C;	���p"O�q�R��oWj��ޜwP���|2�IN̓
��|��LD�'W�iP�eԤf섅ȓ�*Ly��8S���)�ͬ{XH�ȓ]��ᨔ� W���"�٨F�8@�ȓ
&z�y"*Շm�>�q%��� T����}�DJQnh��4��($�Ňȓ�༁"��ng���0�Če�f���/�2�IC�m���WƈD��	�'ў�|�e��'m�����m��}��d�Ḡf�<�č�� X� ���pl'��\�<9��	�N��A��$"�R@�CK�\�<)1O]�%Nv����$p�\|87l�U�<Y ��>B��9iB��K$�Ɖm�<1����h���
��)��_�<項X0#� Pr�6"�|����H�	j�S�O��=��cٵ_>>m�1�vY� �"OTQR�'��;���+2��YIn���"O<����=v�Z(!�Iƅ�!��	\�Re*Q�B�/��:)�@�!�dy�R��቞Z���Œh�O������m�z�A��bK�<�a&�#@=!򤄴��qr��
$f9���&��!��0yD�*�$1���!��P�FOj� ���0J"��⫝�F�!�$~3z��T2aPT��CK�%~!򄏤P ��7Iے$N�0j�KE�j�y�ት	����U��!Ԭ�SB�U�K��B�ɲ�R����ðq����FcU*k�zB�I90n�g䑭@CjM�e�T��^B䉁"?�������#x��b&��s��C�Ir�t�����?h���bZ++��C䉄}�i'B�$��!�S��B��&�jF��F��V+Сm�C�ɊX�N$�g��|X|�N�`�O�=�}�a
MO
�����ܘ|=|�i�e���ϓ!��!k�0rCVX`Ƙ���݄U�虥c2L�2�B��@���ȓ�|����Z23잁zw&I�f�����V812�ş�>���z0��2����U�|��&�U�V�tEBq&ݫ�Lц�&�ޙ0F�,.��d"1��'cBDP%���	z�S�'GdZ��40R����u�B#AԈ��yc�QkMX.m�ސbuB�`�詄ȓ�L*r�@1��(��	~U�H��- ���i�}lF�P��X�,��ȓLTm��)�,'p����[/g5r��ȓrn���E��I1��t�	���D��I<���f��Z|:� +<�V�&���	v�Sܧ 7�Qr�/4Vr��bN�.zB8��d�'9DQ�Y1� �kw�����YTC'D�|K��˜n/Ȭ���]�o����M%D� 8��(TŢ)���N23�؁��"D�D�S�&���[��N�K��2("D����n�g�H)�d�� �J�`�O=D�<��^w9�U�@  �.!я0D���n�$>A�m��펏G����+�����p�N\� �Db�n%�śq"O>�+Q��~hR�(S(����"O����"��@؄�tHG�y	N���"O�9#�⅃8��J�I"	�\M�"OH��h�>V>Ap��Ġ(��K�"O�A�s&3+�R��E��)B��"O� �,���S�Md,9#��A`�@�'J�����C����P�Cu㰝HD�?D��3��B
(Բ�ӗ� �'�����=D���Ċ"^�i�*[��L�f�<D���G'݊Y� �x)��a�F:D� K1�W,#��L9/\��R�6D�0�&��:fr�jU�e��Q�,4�O��C?���GKNg}< +u
>z JՖ'6ў�|�VK�t�H@e���&�+�#�q�<�!�H�	s,� ��u n��lk�<I�炒8�^E��GB�X�h���h�<3��f�-�%k�:w�x�PM�I�<#d^�=(�-!�A����@P�<�PA�">��i��	Z�9v�rx�P�'J�܊3(7 �
))��Lq$��	�'x��A���q& �V�ùN���'��ة�h�).V@�,.#<l�A�'}|����ڹ&͠m�5b���*���'K�%0�w&y:��4�ȓ)ބ�G&N�}���R��U�F܆ȓh)����ߦ\ �lG���K$�<�ȓy�lM��G��C���h�5�J-�'�a~r��9@h�e�R�'>��6�֘�y��H04�(gボa�@I� \�y�m��0���/L��i��y�+U{���W"�
G2��X�L��yBcB'ܬ	����34"�� ���y"dܽ0h1����/)�"�	�G=�y���"LyLmE@ͻm��D3�K��y"JQ'~��E�R�҅dD0���A�y2I��z�'���bu"����0�y���!=�B#�	]_(�#�^�y��X'.��MBW��h�������y���	��D9�'Ϩf��xER��y"C�R�D��7,��uz��pc����'az���U� Hx�+L�?u`�@���ybχ���k���G��]�.���6�S�O���-WyG�u tcѭm1���'v�@���J�@ �d�h�U��'N����R F�s ̏�=���y�'�bPJ3���C��0y��Q2�ةH�'(��R�k�*a�4��&�T,Y�����$0O�Y�!�ʓ �q�S�%�h���"OD�Iॊ�o�j|�5�Ơ!T��|��)��E6D11��52�e�vm��mr>C�2A���"� $F&M��d�B�	M��I'`�}�M�s*
�F�C�INX�qY���+_�Bɲ$��>y��B�IC� �i��o0�u�v�����+�d�O��?�'����7}��榋/ n�
����يBQ�a��愵e]v�K������'\ў�<�4�֡Kך�3�k&Z� ��k�<	�l�H��P��^���P���d�<YcDO'oC��H @C�:�= Di�`�<�ǨW�k��3�,�!/r�U!CK_�<Y�(K.ߢh����8@Y��Q^�<	��q�)�n@.k,̚&Ɂsh<��b�.sg�P�cLL?�lYA����?���?�L>1�����bC��V��@�T�q%�r�!���I���9�	�,Pu!���!�d?!d�!�.���5"���PU!�$�L�*})D����Y��$8!�$��q��u��������)��!��D�R)��[��P��8�נO�!�� ��BuC�&hֹ��I��pPҒ�'�!�$��:�PrFN� K�BQ�����0!��J�d#h�c�
�Vu<,�K�!�?S�LV��ZH��pcC�$w|��ȓr����+)��1:�D�
A���@�(�G���p�@5ie����܇�a��1:�ϝ-I:����̂'ˤ��ȓ_�*�m�-�`���=,A���	iy�|ʟqO��z���5A3+K70H0�`�}�<�e�/Z�əƊ� 2=�4�!e�t�<3���V�@�^& �)DIV�<	�AՏ\΢̨�H˗dD�Q�H�Y�<Q��E�^+n$����I�#J�q�<q3�I%(�K��n2�89QN�ph<F%��A��Bĕ24y������'7az¯�K��{K\9t�\�A�(=D�`@���;K�PXs��)9��8i8D�tQ%��E�^��'�9AeVI�SB5D��y�ޏ��1��=0ڱ�F�.D��C�a�5WӀE)��.]J`�P�(*D�� %H9K�ȓ�@� ����=D���q�� +>�%��-�(-pE�:D��zEK@�Z��Ԋ����9gTeb6�:D�89��*%��h���6��H��*D����L]�=�X��L�G��p� $(D��2Q%��v=�� ���) u��"v�&D�d��ĳWs�h�� �:= ԕz��$D��p�B�(R��C*�: ���: �!D�M@]vٻc�]	�܀ d!D�"�I	^���ICƟ2�T���"��?���	�N�!�5F�,7.� ��2~�!�D�I���rQÞ���<Ŝ=�!�d�	� q�e�C8;���;G㇈&y!�ǪQ����.�a���Bh�	!�d�+X�x|���O�ux�I"�� �W!��{��)xS��J����\�i�ȓL��ݰ�CJ�f��y�Ǡ�^�D���l>=@�G �E-Rو���M���� D��Pp�YS]��G�� j��|�j?D��e,��N�B����&�Nd�נ(D�̓TC_!"��y����R,����9D�|���sbh��m�V� �Z$o8D��(@�D�:�x�e�%��aH6D���v(�c*�=�tm�4�ݒ#��x�"<E��'���{��
�ٚ@ɝ�q�2"�'��Dc�k۶�'#��Y��l��'��	�Ũ!l����^�J6R���'�m��Ϥ
X>m�pK.APı�'�:Edaڔ)�δ,T佹����yR�ѓy
�Hf!J+^����w`E<�y��['����_:E�X1�5�?�K>����蟜�1g"�4"���"Ӧ�^d�w�0D�@�mX�/Ӽ�
')�(�l��׈.D�\�AB4:ON�
�`� Y2 +D��H��":�btس�ů�6q�g�4D�,d!�z�z�@��G�i�X����1D�l���L3K����d�"�*�3D��kbj�x���	��T?����2�Iş4��Ӝ$��	�Am�����K�h^$G
C�	 R(��[�Ȕ�B��BS�Z�L�C�	�h�*�tH�|���D`�"i�RB�	:?EI�-�GjԤӷ��E�B�	v3�HEi؊R
�arGAPFC䉹-���q�4z)�ⴭ��qW�C�)� ����G�
e�p9��D'������8�S��djV8!%`W�.�@���͇�/�!�Ď6ӠLk�̇�y�y
���,�!�^Y��Ȉ�7B�z��UG�=&!�@--J(�!A���Db��E=p�!�āXY��0�c��u�|[bݓ(�!��]�T�P�S� x̍�!�3>f!�D �����ĉT�d�ptJ񃉹@F!��6\	J��A׎e��ĐP#P�^�!�A�Cw���Ck<?�����BOD�!�$Wt��"�	ȸX����N
	�!�D�)XPt�f\�>����F)�Vr!��6u�<�Ӓ3�\�	��� :g!�/K5���n�<a�gû�!�ە694���d��Lc"< �d�?!�0[�4��r�R�P�~� C:G�!�DӐ*9�Q�0 �┰�=o�!��Y'hpt�@f��DP !�;'���d�<w�������=���`(��z=HC�I�0 D��a����MJ/��fC�	�@��r��><��q�R�0Y��C�I�R��K�M&$�`��.b��I�"O�-�A	Ћl�v�R�-Q !b(�d"O~�i"��A�H��΅L*@qI�"O�taC��s�̑s���:'� �S�'�R@˩,�i��� �~y�t ��!�DҨ^<��Rō&	̵!A)�0�!��yB)�k�&u��<1@f1P]!�$�a�d�c�GӰx�d(��]�9�!�DP������N,�ƍ3�,�4C�!���Bo&��Ǥ��s�T@#l�� !�ď�%2�(��Ϻ9�2�]����DH��4�f���)��9#�<�C䉆@�����-԰(<U�G-� n|C�ɯ
���Q̓�ĉ��LZ�6�zC䉜1E^�RÄ4��da�L�K�TC�	�:�|��D��J�����*�	9��B�I�E4R aڇNyv�� &�&k�C�!�,��f�]�J�txj$,6�(C�ɓ`�4IG���@���g���B�ɴ�v��&M#)f¬�C�^԰B�	���LA"(�)T�1�_)XӂB�	�q��e��$��p�ٞ���=�	�����ƣR��*)P7�D�4�m�ȓe0�2�DE�~����ȝ9NtU��Sm��7��/h�%�dK�6g:|,��dP���Տ]3%���1��S��\��E@Tu�8��;�ՉV����z����2fI#���(G�$4�����Ը8��,f��e�t�G;�J�Ɠ0䩵7��L�D�?MΕq�'��Xg����24B�0A:&��'��,����]x��	G�"����'Hx��Clc�b��*�\�3	�'�~X8�L�0z��1�R+&]J|��'�����N�P��4�բ:����'���a��Ѻe[@�G��/P�I���?!&�A $���̴f&&�bF��y��&�hh']
a�	r���y���-:���EM�R���������xrE�.(^�HQ�	ښx��ĉ�%G#b��Io���9F��!nv��G��T�t on�<���0�@$I��L
L���O�<���)�l�J�Z��"��՟�G{���1� H\鲅��>� �r�Ȣk���"O�����I&�$��c���Z�"Om��fV!&7�iA��J@rN�sO�xY�D�C�������
4?�j���O
B�	�#v&�E̓i/���DH���C�ɿ%���)�/jؘ]Q��T�v��C�� dj���ŢC�P�ybO��B�$m�6=�3`�!.v�@aV�irȄȓ6����S�zth�6<�9�ȓ�p`���ުDC�EP�%�1�5��Q�w	��&����1�![n#�P��AK��+ϐ
^���Ňу[uF��ȓh��)�GC�71�p+��݀r1�e��	z�'�d��a�_�*p�JR�}� ��'�D���p� ��l�rK�5	�'<t��ٗ��L��Ӆ6��L�'��=as`Z6#z�4�I&&����O氛2fA3*�f\ #�:���)�"O؀���`�p�#o�<9�"O��a$gͨ�ց�#V$=�@U�$�'���:�D@R�|Jt��%�([�4|O|b�,��IR	Wi~M�"���>h�� 4D�@��k�9�Q���]]�8�Q0k3D�D��E6�&�q  �C�6�+�o,�����Jd��I]>)
�� �$�Ի�"O�1��4 bu�� �|��H	"O�M[u�;�r�ه8�X=b"O��c̎&��3�
]>�r���"O����P#��v
�(-�D �"O�"e�x<ssdD!���I""Od���L)1d4�Ӏ�P�YQ.Y��I��@F�� �	'7<��aئm�6�Q3���y��
#/���أ�0zچ5@�I�yҦ�iM�8`�;t���AN]�y���N����C�%m��d1��Q7��'�az��,c�4m #W>X� �%�Ķ�yb`8f���KK}��(�UA���y!ؕ:eb�����u	&���y���X8��B��D&l����	�y�'�"O�h)����6G��IcC���yr%��/��}8V��%#80�ks�@�y���@�.��c����Q����D�O,��-LO ؑ�4K�B�I�ޛ*�PP"O�3 ���1 XA��!P(i
��p�"O,Pñn���A+q�T�@%�8�"Op�JՂU���b oM�1�Ĕ�"Ov���터z,,I�s/�6-�(H{e"ORB�KE)1^U����>P���"O|��#qn䑹���7�
��'"OR�@��Mж�P1��4F�H�a"O���"�PB;��Y�Y���"OF��M�f#@ ,�F��g"Oj5r�A�;.Ad/rQZ����'%!�d6`^��A_�wۨ	P3�@$+�!��'Fn��ĸt��"Q-�.S�!���\v���4�TA8��	�;!��(G��:G�|��LA��d�!���1��Uz�ë^|��8%���5!���+v�"�y��Y�w<����!��D;~���qB`B�S3qB�N��!��FR2|�F�G'ft%�Ҍ�9�!��RS�*qF�Xb*MDZ�!�C+�.8��`�. f�����!�d\8{KxHZ���
��I���s�!�� �1v㇞�x�ʴ�M�fH���"Ov��7�^\��<�h�8GJ�1kG"O=P,�/y�z$1�e^[������'����kC7^�T�&NȜ7�`����<щ���&������IRP�!v E�I��B䉭g՛���!0�;���m}�B�	*�����)O)~T�I�5NB��B�	�]�HP�Bf_yi����@���B�	k*BY�a��"I �%8R�"O�d�mթB��DaP��+i
�7O$M3�C�lp��BEZrX��2�$)�Sܧh�:E��q�8#l�zl�ȓ&浺㏘r��5HQ�ǝtzTtG{��O�h݃W��9B�	ڲ�ބbG�4j�'�P���U��J��2)Z�R`h�'�Ze��A̒|Y@�C��#	���'����?oV��"3Qb���'��E�r��yظ��u�ԑG T�K>����i:z��hZg��u��������_|!�đS�(�C�(#�t� ۿqU�IA��(�x�@��K�G�܄��jF�@���"O��$ڣ#�09*$�V$h�T�g"O�4��j�4,ČsaǱ-�>(9b"O��a앝s���*W	�m�mb�"Oxف�IȉT�u�@�Ї"v��RG"OPx5�[3(Vd�j&�W>J.p@"ORlB'���E"� q)?b:5��'��'�ɧ����R�eQCͨ$YB*G��P�.7D�4H���2�ʌ�Aߠo��`C��7D�P�W"%.H���=)~�!�L(D�l�`�!�$�!Th�)@p�� �:D������9$F��1)�	A��Xօ=��*�S�'P[BPz	_�u<N���f��LA9��~B��i���5:�^�SԈ�"hΔ��۟ ��y�)�=�x��'cASӤ��c�C.�Q	�'�0U�p��$��}@���%�J�'$֜��T�<�j"�B�.R�		�'@6� F�� ܐ�{�f�~uzA��'ڮTjEe�j��2v��{�]�'^���C.8���ɴ&�%��x��xR���_H-�c�ЙnP��T՘��d�O����O����O�[�Pa#�DM<MβU���!��P�0k��BF��)�� V�QP!���v%.�����/)78!�GX�pp��:A$���F�T�s�!�D�j�� QĆ	Ԣ�f>��{2�^��1 2�	�e&I��{��T�j,x��'[.�Hs� ��Oآ=��
ɻE&��<��dŁ�~��:�"OHh7(�*D��1���+���k"O��)F"Y�N^m�R'X� c�"O��bᙼ)�X5��?]�H��"OBA�rIIHu 1��n��&;D��ћ|��'�az򃒝(и���D_��� ����<����'jxr1 �Z⭚d�>�	�b�'�a�t����ЬݽE��A�W!�y�휆<�6�[���;6@��K�M�=�y���g�F`��>x*�m��c��y��@�R v��R���ZLdPe�+�y⯄2E뒅�GcR�U���B���$/��$O�1q��++d�ܚC��x��p1��'"�󐤋=(8E�
��=	��>�	�|��M�O!��j���K.`+�͑h v��
�'�R�(��<�vqz0AƺM�:dr��� l!�a�<a��4re�E�t�y�"OP��Q��:ʤ2F�����ӳ"O�!�U#T�2h�8�$N��>\���"OHxQG��\.����B� ���J��'m1O�k��	$C��qɶ"�lY��"O���R(�N��%*� �{l��"Oh�)��Ūq*$����>V{)�3"OX=C�����S���yc�� ""O�M{Bǚmz�dc	�Ue*%"O���C���H�8<���I-_'�)W"O�ًW��t��3b��(�i��X�����k��hȤə�b� u4I��'�@)!���6��ݙt� ���'� eKC�V&ǖ���΋�}���
���d�2#[z����M�L��5Y#++D� hG�>jV,b���0�� K��'D�8+��[�w/t�z$AIj: �	%�	X�'j�I�m��[��I�g��(&�
�>B�I*n��[��P8 *�y�JBE��C�	3"��$g��-st�B<i�C�	$K~<���ƌ.崕pE�މd�C��<@R飠�2	@�	�cH��>�dC䉢(2�F��7k�ӳ��}�jC� 	�J��@�Q"�
@ U�2U����d�O��mS�T�f��C��ag޻"v�C䉉6��J����o�a�!��ӒB��, &�rc�� '�]����2	0@B�w�DqA*������2"$B��	�(Q�v!�@�¼���P;��C�	7�>e���_+��Z�%����C�9pB�[���/���A$��"���d�O��$�&�N�r�ǜjFB��r,��f2��D$��S�m�<�Ȍ9��\��  :D�<Pe�1,�b��N��h��C8D�
/�>U*СZ�`G6��'5D��`QK��"M:D!Ǩ^�FҰ� 3�4D�����9�$\�����?��m�'�0D�( ��P!�F�acA����j�b-4�2Dn�R���N���<#���ן<���4+68��Z.6��+�*��z�p�����)X�~U&)ɋJ�P ��<D��P�l����p�G	x�L�!/D�0�7������JY�`UM@C�?D� rQlx'���"���x��)D��*e�M>�R@qD(U+9@�;A'�<����/u�vT���y��d
��ݠ��ȓ!�\���lB�c�H�`���)���IaTU�,ۘr�6	�2�$;����d^��/Q<~�f)r5C(��ȓl��t�EG 'pxy:�BͲj����ȓWdi���,����Ĕ9Q�݆ȓh���P#_d:�aen�7DyF��'^ў�Dx"D9-�B�H�J�
�1R֧Y2�yB�.�0YqB@T�v#M�yM��*�P%C0�C�8l,�QC �,�y�������0�����-�y�Q2�����)�hx!��4�y���7FU|YHu���*$ I�7I��y2# )�ܩj��6dw��8�?	���?J>���$9��XB`ϒ�0���Y	�'�x��Ō9v� Pq�M|�l��	�'l���Ҏ�]�Ɲ�EY�pk��'�n0��g��+i��ar�Bb�pв�'��	��`�%Ad�9j���S\H�@��� ��;��[�<��Y�O]96��4pW"O"5�r�M�[X��nC&m_�` �"Od詠R�+�x\P$�=vl�ը�"On�TD@��FC�*;^`�d"O�ұ
�8���h�,^����"O���`��u�u&�N �Au"OQ���$��ô
Q�J.�y�
��:�����!Gf"���
��yBJ�HM�%���j����V����y��	q����b̓e��œ5��yRK��]�yz1*�p�r��H�7�y�Nޢ.��-c��Y5mp���D+�y� �;��q���Ӧ8m���� \��y���Nah�;@dK�|,e��i͈�y�`�/T��؄K,��y$l��y�F��S� �Cd���
B�Ac�M�yR��E��@	cX�1[�	�C̈́�yro̔�2<��n�%r�(��Q��y"l�0w���`.,n�������y2鏦H�6U[Vi=a4���KS��yb�9�T�إ�X]�A�����y�"S� `��;��G���-5Z܅ȓ=\�X
��L�m<Z��Ú+�贅��L0EN��	��c>5J^|��Bs���L4������2iLq�ȓCo��C/�e^!3Ш�F"�ȓ`�"u�Gk�)<&^M+���H��<�`�acF�.hk�;�� �Tj�P�ȓ9葐�  nK�@X��C<����IJ�`>����JĶMsV5P�,֜KɌ<�?�ӓ�b��G��7�q�eM�3���� ���i�K!��24�X�����N��q�х�� \�p�n��9�X���,(��S?f;�أ�&b�x��f��H�3NB�}�:p��fU�x�Xu�ȓM�~���W�r�r}���S!GʼX����${�QW(�Q�Kl�><��P���O�0O�ejUL��$Ėa��g̾)a<8��"O$ �Ҍ:�*�7��#uT�Q�"Oph�E(Z�W�4Lc��6+7� �"O*�@�h��� �&J>�B�"O��a2���+fb} �G�B<��"O��P/�}LrHA��m�]��"O�B�ݞ�0�Ā�*H�lm���'r��'x�dI�vD�A�iɿ}�|�����'�a| ��08$GBA�4�H�vaɡ�y����$-J8@�M@�5h� ՠ(�y�ڳr�h(��"������y��W��}H̓2V�)�iÅ�y�H �pt�**TtJa�W*�y�A�vn�A�C��P������y���:�$�C���I�$��y���h�|*�gO$&�U�dn�#�y�n�	A�pP1fK�� �l\�yB��
q;:zq�$
����FL��y�M���(+e�T({���Z6�D��y4�.�3W/U�y���[6�ߕ�yr���u�eb�Sl~�hxEN�.�y�i��QD��S��*`L(�z��y�KT���c"@ X����j݀�y�Ҏ}��M�sDHKPN�r ���yB��.��@k$"�/��b�թ�y�E16A�2�X�V�&���8�y�n �%t&4 �hY-M���E�B-�y
� ��#� �%�n��c��pŐ�y�"O���2i��C��kdH;5^d�qA"OZ�����2'�=���OEQ����"OP���獧t�PpA�&ǰH�ak�"OV�qĂ�-���x��
�p��B "O2tX��N�%@��3�M51n� 3�"O Ee�FHx����̀y�@4*�"Ov�� �Y�|�*J�#Y�k�ք��"O��CP�
1��<��L]�]��� B"O�5`��;b�&d��
����IR"OL��V�ٸj���S�2O.�A�"OB����:J.@�����2:.|j�"Ot��R�ƒ�J�SLc�a"O3p��g�I�3���(�
5"O"�X��SR���A�U�|��e�B"O���C�Jă��	3V����"O�m�6��|u�7A�&�a"O�q��:	�D����l p2"OB9��,^�Y�t(��/�i� �F"O��Bv`^�X6(���E�d�"O|�4���MlJ�[e�^� �P�"O�rI,6��u�#�`�ш�"O����L�J����`�R�|YV��"O�Lr�Ɗ�?�}��@�Y2
)�1"O�� ��p ��D	/>#v��"O<�{�@ �	��R��Ű	
<��R"Ov��ʃ#�Ι62����`"O��:Q�G� �L�f,0z�U�U"O8Hj�'�/z"�Jk�xy�T�3"O:5��R4�lzD8f1��"O��p�3r�H\��A@�eM��!"O�8��JS����	W*�'�&�2 "O���	��S�(j֩��\��]�"O��[7�	Q�1gnH'p꾔�"O�)�Њ֮�{��C�@ڶ,��"Ob@f�Ȅ@nҜ���!<�-�5"O��:����U��$aRU"O�@���6��ekփ�����jB"O����#˷	,��	����P�b���"O���&l�ߺy�eC5}4ZX�%"O�,
ã��#ⴱ�����<�Y��"Ob��/��b�0��#W��d-�s"O]2F��![��	�e��o�cE"Od�� K�=
�d���K��Vp��"O�MB�ɖje���ͺT���X@"Op��-B�y���ƤI^�u8c"O���5��to,��A�T�8Ke+�"O�]�S� Qt����#�����C"OJ`@�g%��DzA� ���i7"O�TɃ+H%��۷�f�l	��"O�h��L�q)ċگ����B"O�����ѢZ�P,�fMM�8��L(W"O��!�w��h���P�d�L�"O��C��ڴpQ"# �;�($�"O2� �B;hd�DHB����"O��ҐG	���ƣ
1	5d�PA"O@0DK}�ՉrcR;���
a"Ot�هb�o��Ac4���9"O&���Z	V����1☛	����a"O
�X@�s�8�W'�	�r}2�"O�Đ��T PQ�M�p��Tn<qs"O|R2�J�@3���oKtY���P"O���MȩU�҄��\����0"OJ�	q G`�b9�������3"O� TX�pg��I$<spl�5|�(Pxw"O(���T6a��Y�@��� ��c%"O*\�%j>,Hy�Q�K(�����"OH�s��ȐQ�i fI�$��`d"OD��ҨǳfP�H5d�5K�� �"O
�a�Q�����;x����"OF,XQ�&@J�`��_�WPb��&"OFkU,$,�}zd��,1�Ա"O~�@�&�$Q�R�!r�ڽ@!P�30"Oȹ��I�;F�aSCC�.��"O �!5T2qe�p@��l�R�`�"O�����E�j��- 0���H�9"O@��+1����a��)�(p"O�!�F
������֫P3�"O�P
�B�nUDA��`��/(�*�"O:�r��̧l��*�,߱)7��U"O��1w��2<ܘ�CԦB�t���"O.i�#E�[���8��Ȭ{��ak�"O����A��H��0�������1"O:)"�.��1ka\�|�șQ"O~drr	�6�*�a6�	xL*��"O�@"u�;>
�M��]9#V)�f"O(qwJGC�(��-���
a"O$ ��+�-� %V�O�T��"O\h�O,])�ҤӘ�%{ "O`a��46
0X�%��0�����"OF��D$���P#ĺ �JpBP"O�Qu��15M�9VG�6�4%:�"O|�3l�8`tP�#���	|��H؇"O�ia��ڥl�PY�^4���"O�\� ��e������kϐQ"O�t���*u�d�T#!f�q�"O����O�0�0z�!�z����"Ov5�vϭ0��aq��&E��4q�"O\��Q�  N�Q��P#E��P�C"O�*���TX�iïP��Ũ�"Oze2$��;#��run�~�p�7"O������*�;'��bf�h;@"O �r1C�,y���X!�֘c6e��*O�Myvj�n4�zb�ǧ#ޜ��'X�"Si�5�V�;C���M
�'6�ؑR'цh�Er�	XN���
�'~l��%L��jMT��1�P>L�V�9�'��i5�V�L/�@���@�~1��'-*XCP"(Rl��" ��@���'T�P7�
�uD��R���93��a��'��Q��B�q~��dǏ�2��@��'K�h�sϐ�%i�)j�U�,���"�'�� �,țT�H�iTKR�5 ���' ��Ĩ�6f|r �6
"a��<��'��(�Ѡ�T���za/]N��� 
�'#�k�iL*2�@��hH	BU^��'��zvk#~�z��"�ɚ,�A��fź0����vJ��+�=&�N���e�.D�

*y�ѣ:BV&�ȓM�NT�����Z�
8We��ȓb}h�C��!(�>mj���[� m��Xt�E@��/A8��,�3	V5�ȓD�r=�
��(�p�Ï�W�h��ݸM�/�1���E�L�KM֍�ȓ4i��@�7/!�q[g��)(�:���D�`�I�
�fM�(�j<~Jz5�ȓLYԩ3dʣ^��!�)B�+.хȓ#g����;���R�X3p�Zy��S�? Q��u'Ԁ@r�Q�8�\E�q"O� `F��
{}"]:�ژ�����"O m��,��d��� ��+B�k�"OT��n�' �Uڢ�7D�)C"O����]9-@��N\�C%�"OpȫCo�/?�i��_�7��"O�ma����F���q���)수�"O,U	6$F!8In�:��֟UuBȕ"O���6�Y44�\0��7(mĥ	W"OH!��_s�:a�@5lk�ݢ�"OJ����>j��+ں>{�l�$"O����'�tDPU���(�З"O��is��7
n�|"�עu�t��q"Oڰ6a�1o�QP��ϵ<���S$[��D{��IU|�*i���n���J1��$c����W�#�pa:���?<t��	�y���c��ÇC�3I���ծ�y�1.\ع��;i��H�cm�:x��C�I	.�| ���V��
������d)���-q.��f/D�9��ِ��sFB�I2ly@�nH�p�bQ��Zc�B�84.�����Y73�rd��W%~�B�	�4��G�4V ZX2�o��:C�%��7(�	:o>�@e�$��C�ɮ@��`HR79� ���U42�HB�q[��Cp�Em&�9��X��B�I.h��Q s�������B�I"\, (�h4�=01�F�h��B�I�r�i����`�t ��e�V`|6M)�0!K9v$����C��5-��$�%D�D�F��>"v�@#�F��	���>D��A9g�z抁
2׮�(�B*D�s�S7"D~���@y�����&D�8�OE�R����
lq3�$D��2���"�В&֋I�<�!�<�G��>a�(M5�0�۵Ԧ3���@��4D��(�-�LZ�uEL�O�2���o�<��g?�S�Om�Ě�� �0i�ի�HݐP���y2��K��{�('$Od��S�
��O �=�Oj$����[��5b֦�(� R���/��>�k1� #������0�Jb���c�����D�#�t�XÉ8]����Va�'9���˦�Fx��)��`�V���΅-�L(h��ș`�!�ā�H�bШE�ك'���jqň��V��'��gܓZ���K&�]84�E�a%��^8��	�<���B�:���������0��Ay�>i��hO�T`ShXh��Z� a򤨡�A��O��@p�j�OZ�8!��'#���7G8T&��'�L8��N�M�6�T�W�E �'N������qO�a���� �@�ʻL&��"O�,ʥ�X�du��y$����0��x"�iPa{r�]� F��(��~.墠aο�y���r���;�`�3JPH�����>��Op#~B�b�7[�~ȉv�!$���(���V��hO��ŦAE��hʲ�b!O���#�<Ʌ�)�'m�Jtk�&��v88����'*��ȓI��-�s*x{�>X�7���6$�&�$��(/���a�F�x��&��)2C�I��|�0A1^zQ@�ی'G�C�I�!�r�#���ڠ�a�֥}��B�G���*�چ�fQ���g��C��,)�)D�;�<=�W�[8�C�	gBu�$.  6�01X �ܪ!�h��p?�fㅫ��3�KȚ��D;fJ�eX�`�O� LՊ����ɁD��3�h�"O|HQ�O�SF�� MT�G�m+�"O�`��q��i5A������T�HFxb�5~yL�ڠ�W�� h��J=�2Q�ȓ1~�T9RbѲ`�0����g ���ȓl��z`��)�Б�k�-OG��	p�'�"<I�4��(���$�A8��_�r�i�ȓ	1�����+6�B�s���D�'ў"|Z��"qT��g� ��a�#��E�<AV�ǖ+?�Ѵ&M�F��P�dA���xB��b�*� /�,��swρ�hO���I���h���ψ%Kz)����'ݰB㉋i��[E�	��ѡ��ѣo����hOv�<q�+ Y64�Q�cS=2F��Q�a�TX���O4�{�A��d@���V�C��@VS�HmZd8����}�vZ�e����rk&D�8�WA��X�ٓ�-�>:�]n#D��	�.(�2�h⃕Q4��ƫ.�O��5�CBI�^� �Xa, ��m�f�	Z������=����/�haH�(�O��'n�S�3����2ڬ���A1��%^!��МQ�N�B4TF*�B`Í�+S!�DD?؂H9�bT�� HX+m!��]�3eHA7�I�cD`,�%$ہUN!�D Nx;"c�)?��s��E�HC!�$��
2��
s%��o��(2g����!�$��8[��P��w��xp! �C�!�Ă.>2Ŋ�2JX"�j@e!�Ę�I����+�
QJՙw��1da|r�|���`�XRe�� �{��6�y�!��'��T�3�դDn:@��&Z��O"�=�O1<����#TuZt1mM�c�����'�D��0*�f+RY���]���
�'�RTj��R�"�H2Fw����'lA���<s���� �n#���'$��I6��U����a�!^/��J�'<t������h�@G�Qp���'��d��1����#�	�$�/O���N��P\���Q��u���� 	��}�4�pg�5 ��1�/�/:��B��<D��ᣔ8B��ȥhN���9D�8�/ղ	��}ؖ-W4��y��&9�lZ�#}p4�f%��{p��%/ݳR�8C�	?=y��aM�f?<�� A�'Fv���/ғC
1ԭ��J�`q�L�?xv͆ȓ�n] Ԭ�,A�Hl���V�x�'���2�)ҧlmfa��C5N��M��*�X܆ȓb�7�
�[�!�H�0�vYiN<��v=Z�C9H4��qF�rL�=�ȓ� ���F���ܐ�f�A9H|�H����
�V"/Н2q�U�͇�	{�'ϴ�07`�^�!d���dĀ�'�L�R�_ZF:�i�����N��'��C�ER�T9�!,�u�t��',0@�����B���`!�R���y"�)�H4f��$eJW%�t�z�&�� z�'��uY��*�,��ˠeY�D��'���s#�T7b[��A4'��K	8y�	�'n����`�bC���B�<a	�'/��0L��|�{���,=�$�(�'�I���׼V����I�<��$��'t�# LS> ��(i�$@��� �'E��hO�O;���� � \�AP�5��3	㓴����B��8\� Q�r����S�? fX�C!G8^��yhVA��s�"O&���Y(؆�kaȵ"2�a;V"On�@�
�9�xЛ��1#,z#�"OXl����)mJ,zC�1�]�g"O(��桗j�� ITA#m��S�"O�i�,L�H=�' ����qT*O�`s
"%�P�B�n
�(9�'��Ik�)�<Y�\P|`�ʊ9(ҊmC�H�q�<���4L\��aS�[�ut蠴�i
�'{ܼpl��<'�S��ެ\�t�ӟ'�ў擜ٸ'�fd�'E�GLάa%'��.��L��"O�ɫ�C�4m�Q�F�#�9[54O�<)�����"�/j�,��㏏Ad����"O��맫�26Y����6U�K�"O~L����5[6�Z��
n(�� "Oz9B�"0�qI���9_��`d�-|On���шfmЈXj�eL���"O�m���ʩy�8(*1薡��q�A"O��G��l��K���0��l�"O���� �b���E�X|hD"O�@`��ɍ��9�P�K�b��"O��h���4+�A�Z�P&z$$"O��I�	� ��08B�ڠ"O�eR�K"ª���R3m��"O$a�ѭ�2l^��Bhp �"O���1a ,vǼ�5��5�4��`"O0۠�B�� w��7{Mj�"O(�1�N\,�� Jw��6	U���"O�PZ�Qxd�=�C��(��C"O���!N�<ޥ8�"�m�W"O�|;E�L�M�|�I���K��¤"O���nX�j��xpgiΌ*�V|�"O�TXF��3XNb���K=��Ӄ"OJ<� �� H�A�v�ϝy� �#6"O���mP�*)
����і8�"O�5��J��u:���:kĔ�K@"O�-�p#X�M�p]3�EE�'���K"OX�S�l�?�9�#���?`��"O|�Ɖ��A�6�?B	$]j�"O����.[�����=D&�<�P"O�t��K��xE�5�����"O�]y)��J`��x�����"O�@� �I������/�8d!C"Ol�1)D*07d!�1E���a�"O�(A돱R'�<{�����!�Q"O�ͪ��P�&���I6� ��D"OJ�peʃz1Z|��I��O��1�"O���p�<"���a	ޒD�A�`"O�9X1��=c.�}�a�	5lQ��c2"OPP�^�Hzè��d�k�ᔃB����1a#0���0�'�*`˳�C�}#p1B�G�	�!2�'�Zu��/mwDHkTjN�x͠I��'˜`ǡ7�Bmԫ�}�`݋�'���`��V�"�$u��K�8M�D��'mZ` �D�.�f ��&�><���'�����ȋL���9��!bo���'{ �x-�H�,��pH>nD0L8�'�N�W̉�j�b���gY=[���'�􉡀F`:�(�&�]z ���';b��T��F�P �pn���'eZ5ϖP�����-[�o�� �	�'/�L�7��Hhh}a�A�o�� 	�'v��em�;@`����]3f��e��'�I#A���*��q�� f�T2��� �г�+�17��A������"O��iЌ�~��f˅�j(a0�"O�]@b�Z��$�!)�>�%�f"O�����1�N�SΞ�$���B"O�|+��I�]���7"�^˼�!2"O|1��b�3c��\����\��"O���eW�
j�+'�ܕ`�8��"O���-�#���9��=��tZ"O�X�cĞ	R�w�N���9'"O$ �ꃍ^��@O�9L��Q�"O���Gj��E�N@ӲO��a"x�ӣ"O���R�B�i��O	� ��s�"O�ՠ����g�����*J6��"O�T�"
�*s�]���#��1[�"O�����R�48�Т�i\�;��j`"O�9:R.�@?�
�ݍHV�E"OЌ�L�}"@0��l�x���"O��c�.�n�4{�,��R0d"O�9�N
H��ҡI�B��h"Or-�W���*jꔂ��<PM��"OH@8�J��<�2��`��)4�� "O�䠳DիQ��-(#�6z/R���"Oh��.t��wM���0��"Oj)
�e�7e_`��E�1�ܥ��"O��S5爃ij�<ۆ�&(�n(��"O:�0�/ؚ9����,�54�ݹC"O(|r���)+�T�s��V�/y��R�B�V�������,�����C��u�Z-z��4Z(�􄔻R�)�N�T��NL�T��x!�4olB�0��"D��B�!�Oe,M�G�ǀQS
�r�>�	 RY�J5��D���Z���.!�@� ��S�!��pw�@���$Ͱe�R���JH��*�{�������ɶŰ� �̏)4�H�H�_�eTLB�I0AEL�;v���L�`dJ&Z�a��	+��=`$�~/R31)��jS���-RU�Ü�0=i�I|��'���S+T(i��107 ��p��'_f��([~�q&S6m;�p�{�I�7g]�O�Oj��9�MW=F�̢0 
�fB�TR�'g�LcM�2:-� ��Ver��'�4c0��,���',��@z�$�'D�M1��k�B�� Cdz��
�'nt){���!w<�h[�"^���'�����CFB����%��0��'���@֩�"���i`I�L��q�'��a��nQ_ۖڒ�� tp� ��'�d�㦙\%xUё)�
?V"���?W ��f�m�H��nQ��08�6�Z�h
Y;�"O�Hp�	R)l�\�3���/�(Oȩ�F'BO�Ni+���\7H����7@�\��u-�QP!�������[l��a�,��!R��!+�s���H\v?����OL�k���j��@
���`���"O(Ex�I�("Xq!�&V�l�װi.6�{Q�D�)+���
ޖ,��xR��)��0�"��8\C� ��ē_p:� �(!��*�9r`g�	$X94�iI�㍔	C���A-L�b�����Zx��pC��W�K��+S.��V#�\8"o;�	�\&�Ǎ0J��h2�q~�&>IA6��oB�B��:f&I+�!8D�L�/D�
:�S�-�H��w��5b�R�� �8A�ެ0$Q�x�ң|��O�l˵���v�&(p�ōbu���"O����Cy+Fx3 � mkX���?9m�'"E�YT-�ƦQ"���G~��Z��[�,

�F�*G,��0=Y&A�G+X�{��=/��Zq�Q,R2��
���"t+�
� ���'~�1R�8�@iP7�ϕ(�J$Ç�"�X�!~�PI�b9Ӕ,�dB�	U�:�3�ן��ݲ_d���d��1�u�)	��C�	�����Ғiɀ9�$��мy�@�8�&Y28E�P(��m�����;IO�!�'��� xI!pˀm��)�X'�0i�'�}�t��,I^͓AN��DՆx_&��V�� zj"�$�?bI@A�'�S�m<-��� ��O��@u�ԇ~'�)�/Z"?q����d��;R������y�H |����~�x�z����	[����q�p�D$�sG±P@�'HԼ�d�8X8H�Q��X�D4e�#��8@(���'��b�8B�D��[>B�A��ؠF0qțw���FF֮F��T�I��]e����M�p�:�E��hk� [4S��ij�#Q>S-��BNY�
�y+%�''0���[.$㒅A���5V��Y:���~�'��Xr��?�T��L�Pa�xY�j��-n�ѡ��"y���/�=���ْ�J�B	�T�?s���Ң�Ӽss.���eԠ���.��]R�]���$W����7m�6i��D�p�½�' V�6i붊�)L\ @m]	zr}��r���ӗ)K\0��܊|nI����o��E��F��v�r뒟SRn�ď���Px"��}`���R��Qc���r���G!$e��9U7!��$1w@�}X� �[P��yBIL��5V�_?��Ca��wކ�a`/H�	V�����<�5ɑ!�jȑ�HƝ(�>�!Pk��b$�F>�v́"��xi!k�(gܙ�*�4�p���'�00�qB�6N�^��SCؔ�. {�}E��Āؓ����n� ��`Q*���	<
 xt� >}\��X�Ƽg�.�z�+Ƶ:�����$Sh�k��2LO<̉�-L
���cFˀ�f�U"C#C��ڌ�,|��b �ءC�����B�5%~�'/��?D��rk��8��4��֤ ���j�� \+!��,��<y��Be�^��bEۿzl^ɒA�NPb*� 6�+-S����u��#��|���S�T_��  �I���>��G-گGz؆�>�YÅ Z@8���V�št��-- ���g%��Io�x�9O����ɪ|^���Ói�怠B	:,��E-�>"����?�g���r�	A��uZb�O��ب���	!O4X���]a�r0���[�bT�� ��E<1c�J���(�
;cR�k3��3�$���+�i�EIÖA!&��X,��1�B���3T슲b�A�B�Ɍ.~�0Ꚉs��c����k z�1t�;�)�'7p�L
$�Y�B�رB/��:�ȓh���bPo�<�* �����)�HC�IsPP �5yHtԐ����PC�I/ �K � x�ԗ]m.C䉕F����F%S0,��j�ү]8C�I	Z"�����߂$�,|���Q8y�B�	�'6�eX�/�c�8dQ'�-o��P(�év]���>� ��⧛T�<a�f�o�2�S����m�9ÊSm�<��n-L�� Dg��/�@�tk�d�<�x�<8��W�	� o`�<�Wh� �p$�Ɋ.���pUhb�<���#�L��a�Y���sQlW�<� ��1�]��LH�h��9�d��E�<�B%�yD���aBub��U|�<��DM(E#~��I�J�!rmI{�<���@��$��L!o���is�<�ʏ=~���
�L�0URb�i�<єd�oq8���Њ�52La�<� (O�J��q�O u�\���� b�<A����� �ۧ?T���v�������E�I-G���"�*��q33N�;:?�C�I�ʒ�z A�c�q�D��	+Bjc�x�4�)@qO1�ȼ�"�@0x���="�|� ��'T��Q'�w̓x�H`iC+��k9�9�Ǣg���I����YR��|�  I��t[1�� 4����5��D��mjŋ1 :��	��T���3J �3��K6%b��"O��.gH%��[0��#���dc�ԋ����y3��>Y��V(Zy���^}.�猌>0�~��'�*}�F
*��)��L����	��'["e��eB��<�`�%ĥ<?D\:h�O_2��qJ�
F[JD�SE�W�����OQ>;��Ď���
1�_'E_ʡ��(�><�;�E�}���i�Q`��|9J���ɐ�?��K�F��Ӡ>un�7�"��$X�VDԉ��.�<%o�:d�%>�:n���aP�����S�'��B(�j�C٢B^͈�&M�8�`�ě�?��y��)N�)`y�DeC�鴵m�4a�a#��#)��DP�'7��!2���Q��'l2���cO�yʨ��i�1Sp@��'�:ѐa��_���l	?
�ց�G5-� �%-�C������\+u�Y�O�-���S:��k��,����΀('쀷2>��E���\$\X��]1���(���0�� z��$��if��VA�:)�\=�b�G[��wTj�Bpe(��dM�T�������`� �eK<17�I`�di��J�{gj�����#04c>���J�1&H� ����51(�05��H�(K��K��L�%BD7�ʁ��#�XC�UZ'@t{��*����`"]�3F�Sr�DA����#��I��F�<H>���
1c��r"�t31�B/�Q�Z�>6�J���5$��
�r���ӓm�Ɉ`�YS4�59���Z�)��ɕfh@�Ч$�cR��(�7�d�4��y��]k�gB�p�ș�J+D�|#�a�@q�ш� [OPy3�/�$�C����"F&��)A:D�p�賎�qKd	j��++S!�d_�/"%`G*�y���K��ߺt���=��/�:����Ib|9g�R��4�1g$�;�C��$q^���B�){��[�)�=Q8�C�ɖ<�9j�K�2V�X0��G<y�>B�	�!H%p�+����q�sDH�X�B�ɱ&�D��h�h� -��G�XC䉑v^5�FbW,N���� Ӧ@�
C��6&�x�:#n����4�δ"D�B�"�>0k!�.��HP����B�I* ��yK��(A���Wčw6hB�ɽV9��v �h��oK8.B�I�	�<Ȕ�m�|H���>�:B�I�]u�]a� )s8�rEID*�2B�I E���+@�6���c���h/ZB�I\6=����.d�
2(]>I�B�	/h̸gd�!@"����"��C�	�V%����)C�>�m�DZ1C�ɷV�RƧ�=A�xMK7f��T��B䉷b�J����5LJn�xg�$��B�I4�,����N�~WhSG�hC�ɓ"W��X瀂�>�Y"�MsIC�"O��u� �	<��1��_�!����"O��qg���l�ށ�v�H��a�@"O\���@H�e5LHg�XI!"O؀��gX?@��x�@䀱\�R�1#"O� (���p&���柃<���"c"O�Q�4NV�U3p��&h�.�pp"O��p)��}_���% H�i�>-u"O.Ec�
҈0�lA�d�X7.�1�v"O�5`��4HK� ���TF��Q"O��2w���E��P� ���'
����"O�x)�o��<���(K�P���"O>�K�ATT�yXu!�������"O�(aw�H �-!���EӪX�p"O�1�B���I0���0����V"O�ĉ�E�.^�>4�r'šz�I��"O�	+Qb�8*�vA0�H�/Vlz��"O0E �@@�Ga:|��_)3T=d"O~:����X�b40�Fݾ���"OLԹ+m{E���eEؘ},L(F"O�H�gF5A'�y!�O�#��%�0"O6�+��L/6*�����ճe���ȧ"O�ШE���t�\�7#A�r�Z�7"OM�FM�,M��}�򍐙%f��:�"O�2��x ��lE q�d��""OpR�@Z�>�8
�IW
�H�"O&����
��"I���R�	����"O^ܸk/fnU�� <��xU"O��QJ8D�uSEF�>b��T2�"OAS�H�`����� N�g�ZqP�"OLM�$��Ճ�o�,g�X}�"O�qg�	Dp�������)ǔ���"Ox �ƉH�Kθ���;I�����"OΠH�MA�}^�U͇@j< "O� X�+F�;ZP��7LBoFh+V"O.ܨ��V`���c��>����u"ObU)�=Y���,ģ>�ҝr�"O�tr�nA,J�،Q��`�~`�U"O�P;v�͚̄���DEΌ�xs"O��!��	:A�h�B�J_���+"O�S�b�.����vd�zzY��"O2}p�F��CX��"��(
b�C"O�ْ �E�_���Z���$)EL*�"O�ʅ'�"��!�ī\m
q��"O.�q��a�f(�S�ѩdoV�U"O��s)޳S��SjQ�P�0�"OTu��b��%� �㈀4Q<ȩ�%"O:ȱ��>n5r塚�b$�D"O^h�S0n)h`��M5���!"O�ĩw��f>�%'B?��q�"OL(����,^d�K�珗(�"O|��ԤԆt�z�@7� ����"O���b�Q��8�蕃P�Rh�<�y�K�������	��"Q���y��Um�PM��F��H��g��8�yrLQ`�lTF�@�{�(�c�ڴ�y�l��%JUI���|��8�s����y��J�5r3fM�w'���kڷ�y�넨V�B<� "z i�	�yB��bS=�u ֟k�2�څ���y��#}*x�a��1`�L����6�y�ȨO��i�1�B�;z�[̆��y"�Hy#g�=�2�C���y��;`d����B�֑۱��y��U�><���E���Ȱ���y2��/�|L�W ƇF��<x ����y��قP�
���ʃ%������y����X˲iW3�\���ߪ�yG��5�Աq���>L6t���ŕ�y��ʯ��d�B�E�	C��Ò���yR��\��x�iH/�J�A
�y�	��pqд�,β{�Z�2��/�y�One������"�L�t
��y�N��V�V���$�2iJ�����K
�y""�^�D��1�� �SL��y2$�=*�P|q���9��p�����y���f�6D*���]��tC��yb�	 t��Af��rp����y�̓91�(�s��v��H��\��y���$����F*e{F!q���%�y����!��އ$��irȇ��y���]V�\���Մh����O��yL�u������2{d������yr��h��u��ER?����+�y"K%TG
�k� �&R�B����S�y�F�y_
�p�n�M�.-��m4�y���V�`�{��LˠXX'�y���:(xY��ԃs@ � @��yB�D�Z��M�'�y���҄�y�'˚(��"t�I ,�6�sG���y2�  7�|`��1j����DĂ��y()���sPe�:��xb5��	�y�� `�����ϲ�Ќ9��N�y� DІ|�7.�>@����G�yb�94K�Z'�h� 0�L/�y҈���D$�D��j�P0�+�4�y��~�!"E�d��9pGh��y�G0��P��^��ۣ�D��y
� �����VlXy��O�	#o���"Od�Ѵ��I������zY��`q�L��L�=����O�1pӋ�`f. 2�L��T�!0"O��8�`@�Pl �D�Eg�p3Ѹi�@���!��|��݋~�T��� �ky`��H7�p=)�Iڟ@�9��e���BxCz�B�A��f �@��>D���vk�Q��u[3���t�0�ɍŜL�Ԉ��Y!?q3�i�&	5Re��N#��)7� D��K7"0^q�HwD�c5`(!�߹r/:)�EG���!���q��'	Xh9���w�	�@O	�/���Y
�zH,u%o�.�b GEF�T�P�� 7z\���٤u^81T�A�4	��I��j0�F';J:�3���[����7��;v#��pR�NMq�h �B3|�|�[Wb��ph�B5n��3���I3�YS�O&l�!h��KI��ۂ.�l�֍(7�B������پ)��X��k\
w�6t���:IL���*���λ|�~(�r�
rP0=�d���Vi��MF�\�f��)#A?67�D�D�@`��ʑAP0d��C�ź�3�P�t�~x(��L��ɗ(d��qnRk��Q"է��H����DV�I��$�U8-Vܨ@�Q�.T�|I1o�8}G�xc��ӿxY�取񾑓��5"^0��ቀIAt� �!Y :�Ƒ���[�>�nc������,\2�abL�b�#��>n�肅�S�z���E1O�l ��Ι�or��B�M���xҪ�>�}
�K �~ݬ�� ���J�~�S&r��w��*�����ꖃ=�Ajw�@���������" �"ɚ0N7eѼ��rb
n�<a������#Ɯ�!�\,����67
�`��Y>f��Z��3l/y����R���p���B����k��w��� ��ֺ�X}a�2lO<�r���*,J�U��(�5V�����S<ja`3�ҩI�T8��E��y�#�2I<��t�c�1UjԴ8�,�i'�DJ,xc�.�	�k�!"ꔨip�Q���IrCHΑP�H��� G7��q�jű*��0�Q.pB�	�\-<��d(U�<��栈������/J�qO�']����>���:b!��&�6ܰT�M�$���j`"O.D+��Φ8��иC�_Z �P�P��c��!LqOQ>�)A��!��勊 ���)�O1D�y�F��]w<�hԻ�^щЫ1D��ѯV�9r��S5�٥n�
iuJ/D��Z�%�ҡ(1�P�),��0J1D��h�`��4�v`��ѽT$��p�,D�`� ���3��@�f��� 8@��&D��#�!���lèQ���y�Ӆ)D���g,V$ �q��<�h��J;D��4��Wf%�N�y7���J;D��R�a	a���B׉H�s$�!�f9D��&1d�gh\gMXi��ּx�!�_	E�pb�.;na��A_�Z�!����œ1KF%C��D ^� �!�F
5DÇ˞�@�������p=!���"hW���G��ԀA�`*!�DϝaܜM�*����Ta�	!��oG�u�"�C@1�(��L�M<!�d �.��-Q�)>B]t���:(!�dL&i�F`�IȄ}T��:���<!�d�
P>�s�\� ̔��H�^!�I�&̔��S��������!!�D��-j�02�ݤ>
�`�$( 4!�$��T���r7M���<�$∰7!��z�H��F��{�T���b�O�x2�<��}�<A�m�: �(Q⊧1��9b�UkܓX�9Ê5O���jTq�T�ר<=w��+O�\��Z=?uғO1��ɘCꕂn�Bn©d<̚�C2R�T=�
$�O�y�&�*< Qˠ$�(��A:�'�Q�dɾW����,rcǡi��I��IR. W�D���/�u��!aǏZ���i2.��,�1� �s������>M�`B���*�'��>��J��>E��M\��dXj�F�	�����D���Or��)H#W($�K|r&�`nf�:�!L<|h�� ���e��y��4Q��� ��g�GŊ�3�[�<�s���#V��'�P���,��G�NP�O1��-��]-n�b�X���4{P�Q�Э��p��V�ֈ��?� $)�ٴ5H��m�_�M0��#P���6C6L��E�?MSF-F^�q�>���^�Hw0�jV�׀�҃�A ��?��^�M>B��F�I�b�A	V>/D�XGcoL�����<�t�г4}��Z�� ��
�` �B=0L֣?a���l2�	���O�<w�a;3@��.&<5�@�D4c����ONpB�ak����qO|�ZU$�}2���a`p5q2��hq��B
:�>�R�$6�_�^) ��(/�4���
�l�ZaВH� ����
���������sj��Δ� R��hj��ݨ���O]�xZ�V̓O�h��F�O?H2��E���F���z0TD��iI�{��`��j��Cu�K��V������+�O���4	�!S�V̑��M���a�'�H�kA�^ 2��'��=�ڔk���֫ɼ Ę-Ғ"O01�JòvnU�5��	����r�x+�V�둕|���n@̜(���2L�H�(����y2戉}�� Y�M��F� @coϲpa��4��'�x�g�DS}�r�0��z�L�Ҹ:�p��AĄ���,��k`d��^t8t��KT�lX`�Y5V=p�JTƂ;j��ȓi���*`� �	��� �=x.��@������R:��#�+�?f�\نȓ7�j�1�c�v��̃�G�,�N!��6lV�Ʉ3&;z�e�dZ��ȓ$�����;S���X��XXΝ��%�6����Z�&J�@I�le���ȓ[,���BB�Ph*�SӏϘ&<0���D6�єD� Ne\@�ӽ��ф�"�i���[�>�;�N�9I؄�\.���p�% �b�:�/�43��ȓ09�@�{\(�
��Z-w��ʓ ���PG��<���r�'��WL`B�I���	
|����'(�C�+c&�Qq!삓D:�%�Ё@u`C�I18�Q�EΌ3e� �Vd4G�C�ɛ ��TB�H�����c�C�I�NR����J�$I%�A;�C�I3|�p�V��|R'�<	;hC�:N�ұ�c3��4��<A4�C�I3H>��@U�R�$3�H�d�tC�ɗ}�!au��3$DF|� a~C�	1?w�|(���gZl����92C�ɯu�H�z�jD> zPLP��C�ɀ$�H�G`Ҥ2�
�z��\�	�B䉔T�ً��^	=��QHf��?;'�B�I�}�pd"�	8|~��2"\�dC�	..���hQ��oC�� ��۾Q%.C�	6� �9�/2���q�ŢH�B�ɴ#�phr#]D�2A�P�®g�C�I�y#����/B+WN=�"�\�$��C�ɇT�Y�Ɉ�b�\��F!��C䉒�{u��$�p$�a�Y�k,�C�I�@�>Ii�
��/(�G��%t6C�I���{r])XN��Ҭ�2C�Im8m�.�#�V&��T�C�ɂl���P�j�E��؁�G͇O��B�	�ֺ��VOfL��ڕk�F�2C�	�5�D�1M1 �h�f뉾&�JC�I�S�!`,��c8d�B0/lNC�	����&�P�[�R\��I�uN�A���fmY�%��[�Z����2
/�	1��H='����""U��!�I&�6X���Ɯ7�&L�Cg�}$!��yFFT񐫓�&�٢N�T�!�̾VƤ� fG� �䌱'D�=~�!�ė�q6�y����r�!����@3!�<2b�ѓ%m�7<oDԑ�a���!�� � `@H6R!�J��P$U{���p"OX]�O_�"���zQ+ܴu`�[C�����SS��� �����u�.r �V57�hbf�h�TJV��ClQ�`Ø&gt���%d��E�ᓵXd�	�*!��-C���8^}z]�5` ����-��d�
��Ň7�r��#[F&��BM�,N�����=OZ7�_�M�Չ�9����		T��hHa�?E3�-8A�Q�v��D���[$����)�'(^p$s0��$U,բe�,Qi⹊�%�B�BB�m~���u>er1Ύ6?Ӥ�+� �R�����l[�4`���b�aR�^Kt���ӟB�A3 �r��пF���4;i��@£WN�h>�{o[%m���E��;zȢ�:�3����zɠ�2�Z��	9B(a[S�.t��pf\ +��C�I?K}��RUc�$lw�z��-8��|�xB_7y`�h�f�.����ě�y2��kXic�����HAԐ�y��@.eN��P���%�F�%W��y`Ě>��@G�,��;���y�Aɮ���Q��qRP�$��y2��6,�)E	�r���u'�;�y2��6VЈ�P�eɸc����I��yR�2��J��)odH(�@�y�c���� ��Ð(Q�H|Zr	��y�K��ZA��B�HԱQ�4�y"K�%�p ;�/�0/���*��y�n�=���,K�N��aЌ��yZ��y��Qz�$)+����.$�B䉽$g��#W�ϣ*U��[�(@8Hz�B�Ɂh�RL����'Ki&��s	�1&�FB��5v+���J0�*�ddI�h��B�I�EͶ}IE��/L[.��r��+Y��B��#缑(��HFFl(Z�� t�B�I�Q^򄊦�Ɠ$�.��@þ��B�I8n�<�;���t"�YG.�r��B��=ja�T3t�#h�H0���Lx�B�I�=�|�r��F"z
ZyP�Ɯ�+�C�	5ª���Ҝ�`1��h]�dG�B�	�N/��u���^$	�-Z=J��B�I(]5h���и �Y��L$P��B�	- O&l��EF�0������\tB�	�o�&=��B�l݊W��=,DB��MU�!�f�!i�
h�wh]*EBB���@�E�\+'b��#Ƨ�;{�6B�ɪ�<��ˏ�I����3[�B�4_^D��U�`>ʖ�\"I7B�	(
ol�id֖".�RE,� �C�I�a�9���؛|�q+`�
��C�ɼ~Re�b��t��re����C�In�n��Mʶ:��(gEU,B�C�	�H��X��BU �X�o�8X�C�	 [�^hRoW_��0�U�\Z��C䉀���µ`�	&א��u�({C�C�	�o�Ż��Ze�X"��9d{�C�j����$K
=j/jT�(Y5��C�I�[D
|�$�ԣ}�\�	D$ܬsz�C�I�2P{R��C��:�fڄ[HDB�I�z5�}�Ec�T�.qJ"&�(L|C�	�d�ć3z ٢E.��>3tC�#F���s��� �`�+̀LXC�9�8���W>K��؟J�6C�	KKv���(|�@AJ'a�0rV<C�5�X��C�X�9��E�b�C䉲Z6FHxG�G�%Fr	rF-� z�B�	:LIx@�ћuh� �˞�]hB�I�9��jB�0J[<-��]?�jC䉹'0؃�O^���҇�N�l_C�)� N ��bǊSv�kR��$Df|dh�"O��"Eҝo���K�u5�Jd"OVu@wfH�o�le���L�-����"O��愙�"䲔ꁄ%
��"O��W�ݪx�hS���N���V"OX|���f�R�bw��'�r���"O@�R��H�X}��� �$N��"O���U�>Ӫ�{��I�1�� `"O*�1�� $�؝�䨛�(�ԝɃ"O�	��@C8`;��,K��Ad"ONM�6�+3VLᖁ[?�r�q"O
�c� N�/��`� V�� ��"OTh�2��,��4��N�c�����"O���ᨁ�v���-�B��0�"OV�	DD�%� u+qK�8g"�"Ob�ѳ��F�LA�ъ�+`d�"O�E��:s�P���Ӕs\�LK"O:�� �ځX��!�u����0)1"Od�Q֯�<}�(*$
������F"O�Iഭ�9/��	C�#�V�&�z�"OQ��ğ�J ��@�I�x�"O|LzVO|oؘ�j�(}b �6"O���O�k-nLB����N���"O��an��:ghD��$�� �"O<u�ѠΠ>�V��Э�!Xx*"Oޑr��76��b�L�98o0�{�"OTbv�,v�t-��AD�d��@��"Ov�X��ߓ!:Ѥ�[ ��Pr"OJ���m��D�.���Mp��dJV"O�ؙ��׳+�����*b��tb�"O���L9 ��d�V����ڈ��"O>$�*X-�r	�CC��I�i+�"O,�s�	91�6�p��E�i��Ujv"O�L�TG��$���*�Mڝ�<A�"Op9PӁ������1lS�7�2���"OD��B���X{�Yt R�8�`b�"O�U�񬌱=���8V�5�h�{4"O�"N&AĞd�wo@�S�$(��"O��cL#z��)��ǐWَ �7"O����ճ1��I��)H�yo�t�"O(��Ӿq�0Ƞ�Ρ~k>,��"O�բ�n��FX�B��
A�#�"OЄ��[¸�)p��a����"O@�{�)H)0�.�sǮ����=�"O�%�ą+�X�C���|���"O�剧+�{#�4�2�LcM�9�"O���ucI w�� "K�8B���"OF���A�J� �ʐ���L�X;�"O}�t.����B�@(L��� "O"�DP>O�5s���4X܎�rp"ON��"G�OF�t�rC~����"O�8��Ѧ>~�b��I��Qz�"Of���
K�iy��J5z䠫C"O�0�A��cj2H�UO�Y$��8 "Od�Z�+w+�f�dc\�+�S�"Ol=���v�]wDI:��YӴ"O� qd B�&�X8caㇽ!��{�"O�Px�"��)o���FE�8ڠ��"O�4���PZ �LAf+2?�� ��"O��9Ǧޗ1�-���.	�25"O �J�����|`#Dɝ�M�����"O��XF�_�ϼ�+ǈ��2�8=��"O �獝S��(�- 3��`S"O��I������kr�Q >�J��5"O� �H���EVʹ%A"��RX����"OXs��
���1AO?*1D���"O�E��'R	m���I.�4�����"OfM ��]�"�D+#-���T"Op�abgȀ*�p(ҡO$Zb%
v"Or�c��QX���☉BQ���R"O��ԢR5^6BS�.�--���s�"Oh8	�Ǘ�b_�<���H�;���x�"O��"�@3 ��S�ev��P�q"O��K��\�,(蛄cG+d�X�!@"O~��(�"�����
�r��2"O�kk&<�h`��C�K�vM��"OPD!UL_s2~���b�����C"O��1�"�Q����oU	����'"O@R��)�����E+��͢E"O���C��{v�3�� C_x��&"Oҽ�cMS�t���P�E+P��"O�C$.��Ǌy���Ю�aZ�"O$��6g@
k�,�b0̀�cR�*�"OzE�Po�+�����ʉD��у"O�zr��7+Jo�47�V�H�"OV�	�+�"IѴ�S�L�#_���"O��@/���mQT�SGJU��"O(4sk�6m����(�/(� "O���oޢ,�\��ue���W"O�$q��C8qu�d@Z�#U"O�������a`�i�#=h�C"Oj�)U�����$�A��(xQz"O�`�bg:b=!&�O�ƉS"O~����')�]K����F�h�"O�l���1s6��c�	j�}�B"O���k;7��̣��0_@I3�"O��h�*�B��� E9I�My "O�D�g �:BȐR�u)��
�"OVDH�+ɈW��v7n5�"O*\8�G޼�V ����1��"O�D+��W�H�A�J0i���y�"O<`�7�Ď>&�8F�ɤ˲](�"OKW�M:���b�4A���1��y��+W&�}kv�H>��sbֵ�yR$K�$��/����y�톓Oi�4Ұ)�'=}��a�X �yR%Z:�b��I;;{N���ý�y�F�1n$(ʶ� cXvHӃB��y�Q!C���'��*��0�B��y�Ô#J���d��#Ԥ���ױ�y݁M:��F���1��nH��y�'W�{���獟 ��mڷ�_#�y�!X��� sG����Gi���y2獜&�<�K��\�NU���7�y���5���c�FߏR���fȂ�yR
_��!��!ȉEO�l
5J�8�yҢ9R��}@����?��8rCE�'�y�a�?)���΂�>�,Cc`�1�yR��(}�9��/�>r-�B��+�y� ߐK6\Ȱh�jB`1�f�ϝ�y�h��.�*�A�F�bo�y3&M��ybfB&[�
�Ǣ�-S�t;�Ř2�yB�[|4����6[,�{���yr̾)�>�R�^2�y�X-�y"��1>5�iX!nƟV!49�!g�:�y�	�ޡZ1��D���f"���yRm������	 �xY��KV��yBDځ4�� C�� �&%VŲ�y
� ����1!g��Z��"��l�"O̹gL�D���p����씩�"O�y�` #D��1�/�:�P��P"OH@Q��)o>��m�*:�VE�"O�5�V��!�h�3���[eeA0"OnP�0��O�p1��K�TTN!�"O�	X�P/�0��
۞`?�\�"O��p�Lޚ^-���Ɉ;&d1��"OX`R�o*��B��n �D#"O��ą>²�
��T�M��	�s"O�Y5e�&B��:�͕/�␲�"O���e�)Yrp�P1�R��Bw"O
�����y@"��J�hB"Oа:Fn׳G$ �+7�{H,26"O�5qQ G9$2\��C�!2
��c"O�p��I����C��1\�C�"O�H�3�]6"X�d�T�0�3"O�ڧ�P���a"��u��Ru"Oּ0T�س_�	"�N34�X��"O�5��N#{g44��B^�M3�\�"O������5R��"�@~~$�#"O1���\���'X/DH�\cD"O��a!��,ʼY���3�5"O�XbP   ��   �  W  �  �  �*  �5  SA  �L  X  pc  �n  z  ��  Ǐ  Ö  ��  ħ  
�  ]�  ��  ��  #�  ��  �  ��  ��  F�  ��  �  ��  �  % � Q  {! �* t4 �: B nK �R >Y �_ �e  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m���'�Q�XI���M�\ ��cI
lx�2�>D��c�&q��KQʇ� z�d�D�<D�����((�[E�/_���)��<D��8�ǡ��!D�'����?D�����9'�[歌!����=D�L�끐Gp�u�C��:r���ȵ`<D��1b�E�E����b�3&�����#;D�� c��R.0�@�J:=�t��(>D�����ՌJ��]d��	����V�:�d2�S�' J
ssc�+@����!��Y
I�����i�M�+L�u*Yr�]��.faR� Ĥ>���0B���H��ȅƓ�x6�S#VL]A��aרub�'���A��/$2pt���
T���'���c,�.������]* =A�'��k���1}�`�����]��!
�'pP^
DL�q�����S����	�'�`y t�I7��Yy �_�O�~�q	�'��`+p��`^�����X�;�$��'7�[F�2PJ20���\(�ݸ�'k@@����%AtY{'ҽK� ��'<ў�}3jݼEG�!�a0w+:�) �S�<)��*H�@����-w{�M�W$FS�<aE�*�*�����C[D8���N�$��k�XC���`��G]���b!D�t�@NX�Qd\x2�I���c@'*�YQ����i
2~_|�b�씻)^e�U��9H%!�$[F
�(�����8h����'nL�e��'.昉�d 	+��]��'!�1�5J �8�^��F�#)�q��'�ȍ�աQ ^��H�� �(��'l]����
�\��ՌT���P�';������@;��b$�?_�P��'&�3 C�D�^]�6��XZ�'#2����H�'���p��6VO8���'�@��RA�aX���lˊMgP�
�'�B�Qv(���fM�7`��'��Ik��4($q[��Q(=6���'�����Y0w�<P�RŎ1(�A��� �Y[vDJ[t�#��#:h�R`"O�\3g
Υ6�q�J�V'�-��"O
���h��m�`�d*ܑ~&z�v"O�|3`!��3��E*4�G.	�����yBJ��U���� �B2"�Y'�I�yB���G�� %l"�:}:�@��y�@^�**���"�7|��	�ˌ��y&�%)�""�!w���K�J2�y"���i-��i!^�s��H��y� ��_4��.ׯZǊ�SU]0�y�`�%or`ň�DV�x$d��yB$A(ڭpn�$I���Iq����yr��-]��Kc�ٖ>�b8P0[2�y���5^�س���
<%����D�y��F��P�V�=.& �� �Ң�y2g�6$��2���u����	G�y�οq��nc:�W�7�y���f��9)`i˚|�-y��L��y��R�N�B�3�!� *	b�+��y�N�} ���` �~�~�p%�;�y"F59��haVfqR�tR��y"�9*x�c��g��� u����y�FȦc0��eP�[���`�-��yba�a��B۲V�œv�J�yG[�5�|x�D��I� � F��y"�	R0��JL�J
d9Ď߫�y⫆)Cs譐G*Q�ʄ� �
�y���)AB��Q`C�D �,ź�y�"��6%*ɤ��p/�T��	�y"�J�1�����R7f�~Y[� �y��w���*$�0ff~� �� �yb�i2��*bT()s���y�醏�	�8Z����r���y���-G�4(�\�~ z�"�P�yb��Bq~�i�jQ�^�R���ؿ�yR
����'��Xu`e�bɛ&�y�M��^��@U"�/K�4���̸�y���'J���2C��B	zdA��yB���٘�W��N!�@��#��{�-�)87J�3��_lA���ȓ	[�)2�-C����H�&j���+��5 7N֓N�D�JK"`$B���^�����{ �t���BtՆ�z[>e1# �O8�ّ�HAe�$��`Ê(J�'0�=�&�>.��l�ȓ)zV��CN� %X$��.�8Z.b܅�+��)��A�Ky@�5e�2t�$i��7�H谊�A+�L8�M�g�D��I�( �fD�e��k�,T=󾥇�0Q�}��MYMV`��ڌb�Ve�ȓA�J�{���bHLi��C= |!��0̌	GG"&t�'ϛ7�Ҝ�ȓba.��#�!,J�mra���Zs�E��AQ@D�A��E��ա%� �:o޽��
�U��ʤW��-k�&�#>T��,3�۔��}�f�b�
.�T�ȓ'��T�e%I�b�pY$���vy�ȓ$������P�zj>Q����$Lt�ȓB��������s� �q�A�H�r(�ȓAW����W�X�j�*��<��|�ȓP�$�k`��i�.�ңi�|�n���- I��a��qr h��Tхȓe}z�3�MG�f��xZrE��U��S7���c/�,Q"ύ+IX`��S�? Ԅ�GM;e?��ʇ3��"O�̫f�3\������Նn;��""O�5���I�Jo�"�f-�v���"O5�4M*d����͘6��M˦"O��
��U�z,)b��z�A
V�'_��'B��'b��'t��'p��'Qx�Fe!u���1L]�%*a�'���'*��'A"�'72�'���'�l�0VH�,6' ��CS�Li�J�'���'���'��'��'c��'�*����BR6jii�&Q BazU�'"�'tR�'�' ��'
��'��#�%D�I�|�G��{�`=ig�'���'ob�'QB�'pR�'���'/��/<��(
!��Bj���'.��'Yr�'+��'�B�'H��' ��h��\q�-�'*�".t��Q��'#��'��'Kb�'GB�'~b�'-�Ut
d{b�iG�;t�ˤ�'�b�'o�'m��'m"�'~�'�����n15� "QD�2x�� �'"�'���'%b�'���'(r�'�^��GP3qf�9��ҩ�B����'�b�'�R�'J�'���'�r�'��	�A�jDf�ǈ�,����'%��'��'f�'r��'���'+#���S��<K�K��z������'B�'�r�'
�'���'�r�'ȹ�u,
� ����ڣC
a��'���''��'f��'�2�zӸ��O�Ԛ4*į����_O(N�a@ my��'4�)�3?!4�i5�u�,Żdu�L���_EئP�RI݁���L��e�?��<��[B䩩`��W�h�!�((q�.����?�Si��M��O�ӫ��N?c���\��a­J�7m:5ɵm%�	�0�'k�>!�P�Ms��p���N�T�u�aC��M��,\̓��O�p6=�Q����4m�@"�ũkD1��O��j��֧�O��Q���i���=&�e	���K��A�v��2Nq�dz�ȸ�n7z�=�'�?	S"ٜ��r���(>z�-0(��<�(O��O^(o�)�Dc����R�>���0g�תfb䉹��Z����Iޟ����<��OT:e�؎���]5l�
�QC��,�I�R3�%P�&�S9R2�����K�iD1Wä⡪�!X�x]����zy"X�X�)��<�S��s[�1c�*5܆�d�Z�<���i��H�O:Lo�u��|����`��ӷOG�� H�M�<	��?���KVh���4���r>�H��g��&=b<�t)B�C7X�����0���<�'�?a���?���?���F4;zr�{#���|f��%�Z���ċ̦�&��� �	ߟ�%?�	*�@f_�+�1����P���O�1m��M뀑x������iQc"W�H℔��a�2]�d�dH`�N+[&�E�A�L����I��/���X��T勢�*i�
0�E i���D�O���O`�4��|��)X,G�BEYz̓��D�T�ʶÆ��y��a���Q�O�nږ�M3��iբx91�>=L��,�/2�9���L��>O���E��e�bU�2��#H?-)�w.��f � ���& �;��X�'B�'+b�'b�',����"hS�;MT�6�[�D2QP��O4�D�OΥlZ�j)�'i�7�=���.����Ӗ+� !�`�vz��$�@ڴYc��Oհ�ָiv��3(�ZF(_ 6��AR��Y�M`�*p�(d��$�<AE�i��	��p�����	zPp2BEB��TM�AǏ�B����I��'�j7͆�8)r�d�O����|�w"���H�k�$c�:\��k�K~b`�<���M뀑|*��li��8 p�����Z�bϖQl�G�aӾ1�'|���
B����<�;H:�"�ʗ�I������&:�i����?����?��Ş��$�ӦE*�&G�v�4�x�����Pu�M�Sp��	͟4�ش��'b"��Mc�.��W������ ;�J��� V��Jz�I���l���W�Z6m�t�+O�"�kόP^f�)w�[LR�uS�DA���'�R�'!��'���'��ӭ�PY��(�ఈ��2v��4n	�9���?9����'�?!���y�!�X�\A�#1Rj|��.+_07��ԦM�I<�|b���"�M�''xe�W:x��k���q���ʙ'~��w
�y?�,O(�n�hy��'2�	�������BƄ4ғd޴���'�R�'g�ɲ�M3V`��?��?��iהh*4Z2C�C ��Dc���'�d�>i��@f�	$��rb�(C����.I3]�ƨ��<?��U�p�<��49��I��u�o�f?Y��]t�i�)˲y�F�`�MI�?v ����?���?����h���S�>	:�(�cO�G ��*�IT7�$��Ǧa�.ٟ��I��Mc��w�N�Cf �$�L��,K�4̡�'��7���1�ش'>,p�4����4�`e��Oذ�C�*Ey�l\�7l�A�¤Y���ٴ���O���O����Oh�$Q�q�@J��	+ܲ-��@�1Ax@˓6�NA���'i��闀*��!JpDF/�(Da��¥���'r�6�
ԦU�L<�|ʖ遬�Jx�q�E�6+z��4������4e~�I'A��`Ht�On�L���Q����j��;&,񲐤U
)���r�ȋ���I�(�I��Sgy�Cl�R=c�%�O�)+F��|���  ��XW@) Q��ON�n�p�$���ݟ,l7�M�OY�<̒$��#Z(J�X��LW��mr۴���3J�{�O�I��u���� ����wR�i'gNS��57O����O���O����O�?9�pK�RA�u3 �]�N��<����`�ڴcwr��O�j7-"�$�?<f]i'8;���p�&�8�1O��lZ&��$O4v�7mo�P�W�P���ٔ��A1R �R�t��,��A�O���PD#�s������O�$�O���CC����&�&?N0T�=3N�d�O�ʓNě���5G��',RZ>�Yp��"v
��X$���X��y���=?��X����4j���=�?e��`�2���iƗ���ª_���-����?m�N]�	� ���0y�Y����Ny�Ok�ޤj��3�l������㚂V�����O��$�O���ɯ<96�i1^�2�wOV5�iZ��N�3��V�C]�	��MÎ�i�>�g�i;d�mTp��3 iE�!�	:�ovӤ�n� x(n�u~2�p� ���!�剮!(p�"��Y��٣�3���4����O����Oz��O����|�h�0if�s�YE3���G�)���~j��'�������]�2I���� ӔHVȻP鎼-�!۴tW�E2��i5dv�7�c���G�V	�<�L�_*̴��Ko��P(�����iyBB`�
˓�?i���b9��.���2���e���!��?���?�/O�to��D�`�����<�	s`�����_�J�
�%L	#	�4�?�R���ݴ ��V4��C�n��eօ1j�b�C�#j����UԌ�t��G����'�,֝*K�B�O��H!4|��Pˑ
���)Pd�ҟ���ȟ��	ܟ�E��'�J����Q�Br�E�n�=*�����':~7̓ A��$�O��nO�Ӽ�S�@;7���\=>���W���<q�i��7OϦ5!$D�ۦ��'yz�{��?	hGD���!P����Gv�<+�ϔu�ɘ�M�+O�$�O����O����O�`-���f�l��c"@6S���A������'I�����'����Ѧ�<8ê�)�d�=�t$0`l�<���Mۖ�|J~R��MB�NU�%���Lw�Q�W�ڊqC��TOT ����q+����S�v�xE��^�ز>lWN�G��<N�8�����l�������ן��xy��uӴ�rL�O�d���!~Rj�hW)�pzp�Ck�O�	n�m��[��I�M�ձiA46m��
�^��iڸ#x`-��Ϛ�<���rVf��kN���B�|u�,O�=���>q�ԃ���{���B܀'8O��$�O:���ON���Of�?y)��9!6�1����b�:&�Vy��'��7��in��OV�l�g�%p���Ƈ*o����j��5#�PJH<1��if�6=����Dq���K
�ȡ�Gar��C��@¨�5�Z�.�t��W9��d���y�'7��'�R�'��U@B�˙(G !��K�ip���'/BW��ߴ �$Y���?�����"?��<�C%+"U�%	�M*��9��QߦUP�4-L�����(d�|<[��N�;uLp7��- "����Y�z��4�ν<�2��-���;�N�ӼS�U�
� <��n�*lh9ZfB��?��?A���?�|�)O��n��i*P�щ��0GB�ڀ�0|�jĂğ\�I��M�"j�>1��i&�J�IQ�Kw��Dg��2�n���aӶ��_�$��6-~�@H *�'E�.��So��uw�'���[��V��!d`6�!�Q��?[���IΟ�	��	ޟ��OX<m�p/�	��U���$]���`��u�.<3��O��D�O�����$����u�;��$XI1�Vq��M��|J~�`���M��'���:��.�x!`���6'��I�'u~)���ßkÖ|�Z����韠`�������R�b!�Q5�����O����O�����̓K�b�'|�-2� McGA�G�z�������Ol��'7��¦��M<��FC�S�8 ��T�T��(�l~��:B�FPJE.��O�@L�I���ԣ\�İcqlT:��TƄ�sb�'���'~��ڟ����{�X�X"�9��
�HS���1޴�����?	��iu�O�X�9]*<`m�4v� ���F2���O˓.�r4ߴ��$@*ct,K�';]��P�E��?*�@�F֗#M�Q�5I6�$�<���?1���?����?��,�$��S̍-F�5�ai����$J��I�Q͟8��П�%?5�ɰv9���E[�kQ� ����� �Z�O:�8�)��YrP%����R*Z����|O�9�"̛:��'���_x���q��'N�I�f��� ��N!�lS�ۯ)Y���	ן|������i>1�'��7�1D���LW��Q7o�*P9���I�3,e���ܦ�?�FW� ��ryr
�"O�+dΚE�T��$�1;\��i�I�t8ĴR��O�
�&?��G� ��e����WJ]�<�z������ϟ��	ß���\��6|� 3�&�+����C���Zxz���?��!�������'87�(�䇾��Rw�Xd�.[�G�?e�z�'��#�4���O�J���iB��}�6�9�d�H���k�BՉ.P0ŪBJOr]n�\y��'g"�'2��V��Rh� x��H�]�R�'q�ɾ�M[���?���?.��i ��VAJ@Pc���e����O��mڴ�M#g�xʟ���b��Eր�8&N�5�(iB��
/# X�P�.]A�v��|����OՃK>i�O�<  �JSb�;d\���?9���?����?�|r)O�5oZ��:��PFZ�1����`.�mޤ"���蟘�	'�Ms�2ϣ>I�C�,�z��Q�@$)��5���0��&@��V�&��<��.v%�i�<� z�IF+���m���Fu
�`�2O:��?���?A���?I����U�4���67D�a;�e��k��<l�s}Z������[�'fX��wV � c�\9�p��<&gjxe�'��c!��ƹ,	�6mg������N�X`�T��
R��p�,s���$�E�J@��*�$�<���?��,%a�ԥ+%���0�"�?����?q�����\��՛W$�Jy��'��%Q%g|��q��Z|����n}"�'R!-�D��X>�� !8($*t�_e��$ph<,ӇiѦ��H~�����L�	��Zh
3h
���-�����rC�I�����s�U�8�|I@g�^"_,�t�I��M� K�/�?Q�%���4:���<�@(@t��2{�0�d3Oj��O�(oZ��fxog~�D��=L�a�'�TY;�	p��b���5��A�K>I/O�?Ic�4 f�r�+�*@ll+�c~�Aqӄ̛�-�O����OR�?�{��	��&�Gm��D�¥iĠ����d�O�D-��ɏj6��I�$<@�@��>;πM�Цy�JY�''�ax�LJE?�N>y.O̙��ƽ{
�ՠ�@&c@�27�'�X6��QR��d�|X湙��_f��-�!�[�Ip��ڦ��?��V���I��i%�h����V�Ɇ%��,�n��'�t�2�a�IZH~��;V:��z���4�Zu��i^V/�i��?���?���?����O��Y��h��$J`I'(R*3A�'��'��6M�R'�)�O�m�i�6<^Ŭ�6���yw�&i��;��$���OR�4��ջ�u���l$����>|O��:�K�y���02N�]���C�	@y��'�R�'��'9������4j�x�0Ҫ�����'x�	��Ms�ߜ�?����?a-�b>;l@4�01�IK�<Y�OH���O��'��{��|#"�Ռ*����@�M� �ǈƷ1( ۴h8�i>���O�O���A8m�|�	��e&��A�,�O��D�O��D�O1���rZ����x���T+M�l-a�L�,�Jt��'��v��L��O&��Ag%Pp�&B�!&��$Sg�VdI��DE��Q2 �^Ѧ��'(�A��PR�/O<�Y�̑$'���¢'=L��2O˓�?����?����?�����)J�4f�	���\�4 *��.T+�$mڦU�V-�IƟP��U�Ɵ�����;/ىB�H����&Qǌe�ע��?)��*���O[���s�i��$F	Tδ�r��j�����.?�Lǲlq�'��']�	�$��:�jc	�;�^�ySD�8�F��	� �	П��'��6-S.����O���{�i�b�ڣs2@���nW5��P{�OX���OD�'�h�%[������D���5��g-?ysE���ݴR�O*���?a�ŘeCH��o�ftaS0e��?���?Y���?ً�i�O>� 7G�����J�$�f��f�O��lZ^��I�'pf6m9�i�aXeb�#5X�S`G�R�h�b��f�<����, ݴxd��iٴ��$)U�B�r�O�}��ꞇ=9��j�"�����r�OR��?Y��?i���?q��,^�p�t��6��x+Η1��MP*O�LnZ!_����IӟT��Z�ӟ���/�8���q�"^�84�����D���pٴ����O�ٱC�Q��m��
Gt[T�*��y�ѩ�T�|Q������VA�Ihy)R)[�0J��{k�9�wMQ����'��'��O����MAm� �?Y	S�-�~�y(K����5�#�?�q�i��O�D�'�"�ih&7���r�P�`��,���l������c���Sdv��A��ҹcL~r�;T��4j�>>�+�DL.A ��?a��?����?�����O]�}�`+�!2_�-���(?� 	��'�B�'��7-�� �	�O`�o�b�ɬ0;�p�U�3�y�7'[ V�b���IXy��ܴ
�����
�@�?,��T����)DzA��*�*-�Ӳ�'t*�&�З'�R�'��'�� ˇ� C$���I!v
�8��']�P���ڴz$�����?1���I��^Vܝ(�%W3M���@�}��2���¦�x�4v%���IZ
~:̱H�,N��U	�(�/^��0���Őt�qH�<ͧd�`�$ơ��fa��J�9f�}K�b\�8 
 ���?���?��Ş���ȦՁd�!mk�%r�k�*(��0&Fg8��	� ��4��'���ϛF�D�U|T�A(U��d�бЃA�d��lڮ��n�b~2�ǣM����W�^��dѴa� [\���/� oI0��Vyr�'���'��'��\>)��E�o�r��c�	9E��y�'�۞�M+.�?��?J~
��x���wM���H���[㦋�l�$�O�6��X�)���/?>r6�f����� )d�v�Y�@��yٔ�A�r��B�`Wt�MM��\yR�'vdװ��A��$�,W�Ń#E5B�'�'a�I��M�u@��?)���?����7y;r�+�E���^��'�,�9:�V�}��'����]2�<��%�	�'F@=�D)=?��m�����!S�>��Od���	�>���~����%(6q����50kr�'Hr�'���ޟ�F�I�e�Q��*��>֠�S��
韌��4R �����?9V�i��O�N�j2n��J�ca�IJĄ]�_�$�O�6���A3��զ��'� M`"��?E�	� 6�ʠ���X�P�'V'
���a:�d�<����?��?9��?����5'��#��

t�X�QD ���ަqKQ�Oyb�'�O�2&�/g� 䚁�Y?!�:L��*u.�4͛ƈc�t(%�b>Eh[��ثA���`)V����h�Q΋=�������Oj��I>�+OZ�)7�4>Б�j[]E4�B���O2�$�O����O�ɺ<���i�ԙj��'�@�yWM�o2e�HDj����'��6-'�I6��Ăۦ��4W"��$��;<H����>��$��9����3�i��	6~XTѓ�O�> &?!��K�ԉ��
"Z�xXnB����8��֟8�I۟��Iq�'[*Q�0(��'�Ҥ����= �����?!�:�6���	��M�K>!#����t9uoH�T�F��rd�F̓�?�,O�1:��|�2�2��1��C!v(b�D �u�x�WNg�2�ć������OX���O����A���4H�)|���v�E1#��D�O˓���#�4>��']�R>E2��N�6�ɳ��2
���C0?)�W��I\�S���ȒG�҅�F��?�ܤ�V���gH��y���,Zu�Z�]��*�Bh�d�>a�����C��ȦJF��n��	ퟌ�	ß$�)�Qy�L~���Q�A��#���t0�)����1$�˓}����^}B�'R�E�bg]�DY�T�򎚍2�$X�$]�|
"L���'wֽI4%�?�(c\�,�0�<f�X�RE��U��|#ap�ܗ'fb�'���'���'��S�o�(mhC��9%>���(ZEg��{ߴ�|��?������<����y��C�9�je[fE�:����gݬ���T%�b>Uy�ۦ��g@����)����6g΃�T�< 6�˒꿟�%�p�'mb�'*hZ!�̀)	��aM�TzdPp�'�B�'��P����4���P��?��J�V�@d�ݨ]�|hx��	]�|݋�RM�>A���?aJ>Y'K� ��sc��v�pX��@Y~��.i�a��i�F�����'�҅��rbQT�S�_��X`�B�<g��'��'�ן@��?�*Y;Fi��:�^�Zw�� q�4!t��2���?a�iA�O�U�g8@�e��]�6���L�yr�'���'H���W�i[�i�]�al�T� Γ�:1TD��W������8����d�O��$�Od���O��߅u�.䓀eʚ#�b�� �+d�d�1[�eF� [R�'R��D�'�l%J��ٌr�8���H��n	@��>!бi
66�Vm�)�����c� #xU���pHΙ!�؍�g&�-J�'c�,a�^؟4(ј|�S��K�	�2~�:��Pi��Zg�iZ �\�L�	�d�I��Say��p�qfN�O^`�SGG�tM0�@�@#2Ӯ��1��O�\n�@������\�'ۜt�W.S�"�F��f�̤bF���_(��&�i���t��Ec��Od��&?a�]��. �h
�r�dU�ҧ��hQ��Iҟ8��ПP��ӟ��U�'�t(vዃk��j���>-�%���?q��k�Fo�,��IIۦq'�p�ގa���p��R�Q��q)��"�I���'����i�I'QG�y���	2Ѣ�B%��	�3��%L{��P�	ey��'3B�'�BN�7H�:4*�`�@}�֋ĵ ���'�	#�Ms��Q$�?���?�-���w�c#��ե&��`В��(�OR�d?�)�c �&e`�d��r��zS��<�A��]!eF�b-O�铠�?�s�<�D�_��"�$I2$z�I��y���O����O"��	�<Y��i��MxUJ��`5jqH�BfI��SW�B�'�6m)��"���s���#��\d$PA�"�= �������[�44��ڴ���)$ly��"��:R
I�6�D ��B�D�3%ef@Γ��$�O����O��D�O���|�Ug���1�$�P�(̚�'��DE����'"�b�'���T�'|�6=�8� �f��0.�ݺU�>U�������OF�b>9���Ȧ�ϓ���s+6z��!z�'��͓�u��_3�?i��,�Ŀ<!��?	� _
֜yhtゝm�t�	�&�"�?���?����Ą���P�������ş��bL-Y���1bn��M[�7BC�f����m��ē*���#`�<��Ձ��FM }�'}U��(�:��TZ���ISП@ZF�'�������1@
���.��=�L1���'^R�'���'��>��I8����M�*�DY����/#k���I�MӦ �(�?��G(�F�4�!�2�O�K���kr�ɜQx�j�:Ox�n�.�Mc�i'����i'�	�89�L���OPfy� �_�#��0�,�<��в��SE�IZyB�'d��'P��'-�	��2�It$� I4��c���|�剝�?�@��Ɵ���%?��<-v�u��#U�f� �z�Gǳ�t�*O���yӚU$����8	g˟�?i���.	(a�|(1�N�[ `���O�<Y��׌4�`��O�����O'r<<jI5n~@ 1�B�zЎ�D�O>���O��4�Bʓ �&��hxn��k��UNѢТhY��ͫ�y�Kq���Hc�O��$�<y&W�lM�њb��g�n%+���0 �=��4����Ê���j�6����N��7Y�d�d�)�(�05K�����O��D�OV���O���6��Bm�!�+VZ�[$#�Dj,�I�������M;�a��|���`��Ɯ|2i�]��I���ٝF.��r�����'���'�r�D�E8��1OR�D��� h��(7�,9q��s�,K �/�?Y��;�ħ<���?���?��$(H1�-�*4���@��?Q���d�ߦ�ӆ&�۟\��ן�O/�iR��E C0���,ǒLx�b�O���'����?�V��h��\��f͚;�:I"Y�h#�Y
2N�1	h������i�������|�F7N�ip�͠ �d�pQn V�R�'�r�'����Z�,ش]��((�i���a�A�`;$aDN��?��!��&���a}2�|�6}�r&N%��z�j�����b�Ǧ͹ܴt�Ve�ݴ����%O�8�B�'�b�
�����:F��dH��J�l̓��D�O����O����O��Ĺ|���L�&!�<��.�@%̜:B��0����g��	ӟd%?�	
�MϻWȖmR�j�.<y<Mp�'c*4iy�����OO����i����,�Š�'Wm�Mr5��A�d��B�uZ��U��O�˓�?1�zE� KD��P�+���J�D�@���?����?i-O��oZ/H�e�I���<TU��i���?%��g�pr���?Yu^�a�4oK��"<�D�CJ����Ӄ$�T�h�m�>S�����}����)-y��%?���'|���ɼx�x���G�*��Y�1��4�p����|����|��w�O�����<(Y���l�@�3 I��r�e�r�ۀ��O&�Pڦ��?ͻ9 �`J�?#�m���ear���?�� ��6�ӣI&����	Œ41��i��W���rd�W"���Ti��D�O�ʓ�?���?����?q�f^�	P*�De��ʧ�"S�1/OrUmZ�}���	��4�	a�s�L�1N������dZ� ʄ�׮�2><�Iǟ,��<��S�'F.I1��=(����b*$ﺘ����M�Q�(y���T��$*�D�<�@#͏]�H%h��?�\kF��?���?A��?ͧ��$ͦ!��� Ɵ�y��.7��+7"J|ZԑѠb�d� ����r�OP���Oĸl��Z�@�f�,���k����_٦�'z �k���A�O~:��"54=J3Ҿ2��KA���!����?����?����?�����O d�����	��[�f��4	E�'�r�'��7��6� ʓ`⛖�'T�	|bT�&�&Td�GT�e��<%���Iߟ0�	G�Qn��<��O3�n��]���Y��K����C�����$�d�<!���?a��?q�܋&~��s�$ĕD��Y�ֆ��?�����]צm 4ʅ_y�'���T��	v銗G%�Pa��EW4���	؟�IP�)´���!�j��%OһU��a;w�ʘM"��*��M�3^��ӶP��D5�D	�3�b��gk��Lx\Xumݒa��d�O����Or��ɦ<ك�i@H9�c��?~���3%
�d�Ph���<���'5�6M8������OF�6�]�iIgGٟ2�ȵ�j�O����x7 7�.?�;j�mY�O��I�4L�'K
������f�4�IDyB�'���'.��'��_>���-�x���-���!�&�Mst ]��?9���?y����g���ȅEF���@߬J<0��DK��NXl��M��x�O��T�OH*D���i���3@�&�`�
�q&0̠v#�=���Rk���"��h7��O�ʓ�?�������Ċ�D��M0p+K�^0V����?���?1-O��m�z�$�'?��	�3=^ݘ���,� H����|W�O"d�'}\7ME����H<y�iQI�pX񥆞2C���1�^V~�K�e��*�g��fe�O���ɽf."���F�R|��B�:Qώ s�C�jB�'�'���̟0�	���N�
w�T0��b���8�ٴ^vl��*O��n�a�Ӽ����a3h|��Δ)q>��I�A��<���Jfc�6M(?�CX�Q����5E�%q%-�,� '!
.�֬N>/O��d�O.���O����OBAZq��>`W�Y���a�<�PG�<�f�i�M���'�b�'���y�*E4����3+�$�؛���l�^ꓙ?9��������3�e۔k�>ЃE
%�S��0i�	Q�l4�'Ťy%�`�'��$�g)O69]zH)��ߵ!���q`�'���'����X��p޴2V<p��b���a���o�:Y��
֐=0�tw����P\}��'��ɟI��P�`���{=�e �&�O��!8�D����'6<��W'��?Mk%����w�x��f�A��������ٝ'w��'nB�'��'�񟈅�6Х`h�u�ʶna�a��O�$�O�������I�OTmmZX�	Y�� ��CN�<m�x���M�]uP)�M<���e��I�.
7�<?a"+��1]�c�\�:��!���Q�l͢ ��O�%�K>�(O����Ot���O��r���=J�@"Bf0�a���O��d�<���i�^�q��'�2�'��f�ɩqo�00� TJu#čvI*�Vf���x�?�O���"�1'nh�d�P�
Ӷ�s�KAo��t�a�Ʒ~�i>U2��'��$���p�X:*��(BI�g�t�v�������ߟ@�	��b>%�'�N6�W�νa6ğ"*���3���5�n0�h�O�������?�_�\��R�@���s�M�ƣ�')�	�'�11�i��	�/
P�!g�O9�\�'��)3&�9(̡��ɜ#��]	�'f������Ɵ��Ip�Iz��$B�8��V	A�!�&$�ɜ9cyB6�@�b�"���O&��)���O�oz޹h�jŤd)���a�")�4@����L�IL�)��g���m�<� ����(Ÿ]:�=�W��ih�e �0OT������~r�|B]����ӟ�bIآy��ؕ�̚Y���������ڟt��My�hx���Qf&�O`��O�X��!I IeP���1\:X��(����$�O�D�q�	�Y@���h՝N���ӹOz$�:+������M3����jOJ?��(�ڴ�[*#L�8BJ!L`�;��?��?����h�����m�:!Z�)
�@c㜂�����H���ܟ���$�Mc��w�m��K�5k��RIH��ܡ��'��'��6M�	�(7-)?�4$�L���S�(~@P�B<�l���H�Ě�'���'�B�'���'���'���2ֶ>FтF��=%@h$-�myR|�(�X�@�On�$�Ox�?�c�[,||�c@��.�B��	�!���[ݦ)��44a���Om�5�Vز����H������G2��7��q��I_i��'���'�d�'�>uҦ`�m�*ׅɢ5i�����'_��'DR��Q���۴$��Q���`�#GL�s�`E[2�n���t�����\}��'}�	�	&\� �&�.txb�u��'F���Ц��'��jf(��?�	%����w���*���/ 6
��I4EsD���'���'���'��'{�� �^�IB&c�"abI���<	��JJ��л����I&�di���x����B*WX�(QӅ#�Iڟ(�'6�͉g�i��	�VX>�!$�h7�Q�D�Y���\�!��tӊ�O���?���?	�nj2�h6N�G��ĉ�O�^�ԃ��?	.O�o�~HXH�'Z�[>�)!�؝|Q���E�G
]L԰'�;?-����O���'7 Z}���4�x��栕N4`�ybӇ�8}/G��4�T��-��O���=Fu���"����8���O��$�OB�D�O1�����עD�E�G0]fD�ZD́�3���C��'rR�dӆ㟨�Of�$��u�����ִc��I0�ø|��������#S�u�'��i��
�p�*O������m>xi7��xz�!�3O���?1��?1��?�����	�SXEh�*�-S��e���%5��oڒi�P��	����	}�S��r���+�|D����*�[�^f ڿ�?���>����O+�h��ik��"H�Bq*��B9��.иT��D�*6�U��'��'��I�`�	��zi�r�	�9~J��s-ٛ*nu�	ߟd����ĕ'M�6-��$ʓ�?�Td�/Pذ���AH ��0��'���?��I!�'Ԝ`��`�!头aP E _�l=��O�II����!�7�g�S�\F���Oj-#�ǐ)�V��5��ҽq�j�O(���O����ON�}��	�^�bP� �pEH���Q`���U�D�	7"�'}�7�'�iޅY&L	}V���b� �0h��4-z���Ty��¬t�V��ㅘ;A��T&�
���R 4x�޹
�DS�h�^�%���'b��'���'�2�'�@B� �R�a�R:���cTP��A�4&��q/O��*�v�xm��K41���g�Q)�Q�O"�D�O�O1�Te�JJ��l]����,H.�t�
�fAx6m�y¥�T�8������d�z��[5V#8V�
�h�� ?����O(�d�O~�4�&�%��v� ��ČJ*�h#� H�Yd��'����n�⟌��Or���O�3d,���k�D P��W
��Y�`�V�]�)��L�?�&?a��
N��Af%�C�b�C�CU .����ݟ<�I��@�I��I_��!}���У.7��
p��;>t<�8��?��盆�6��T�'2b6&�۬|�昋���� u����*!���O ���O�i��;,7-$?��K�h`YpfҮc, �%��:�� �G*G��~��|�S�`�����	ȟ�O����o�)Gz�t�F�����	By�|�T���m�O�d�O�˧C5��$Թb)�D�t���%��d�'�^���v�f�&A'��')}�c��H8D�~����^.w+�в�'Y�k�~��J���4������_��Or���iU2c����B��;�T�I���O���O����O1�����&�H� �L�(J���V܄V�6���'���m�&��C�O�ilڴc��4ײ��t3Ǧ,k��:5�x��oZ�XAnyl�P~�(ܭ
��h�S-k��g� Aʀ�]E�I磘�|��HyR�'o�'?B�'XR>�)5k�/�U+���yw:�
�E���M�'@�����OΒ�t������]�"���O��De*�3�d��t[ٴ{��b1��I�=
"�6Ms�Ի&�X��Np��)ܚ�s��[�<	�#�	 �.�Y������O���^�+���Q�û0�lqbN@�X�H���O��$�O��r�F�z�'�b�[8���Z,Dz�[�ep�Oft�'
R�iF~Ox�Q��+�F��vhM�w'�lr𕟜8���;�ZHش`�}�Ӽ��`Y�D8fo��h?�(�&Щ=�*����ß��ş����E�$�'����e���㪊3Lv���'M�6�ocX���O�!o�Q�Ӽ;G�اuHl�o��[9:��`$�i?����M���i�$<�$�i�I���(��O�>��R��|��:e�����!C�J�	ny��'���'���'��"^T�t�A��)HxI��5��I�M#�'��?���?�J~�74�zeOʷH��`��
�3�S�D�	ß��H<�|�4K�`�? i�5�#(䘺VN�C^P��L~�N��'r��Ru?�K>�(Oj�kGC��4�<�Ս�%]P���D�O����O����O�I�<�c�O�����O+�!dfߑ>���Ά�y|����s`���Y}2�'�Ie��S Č�Bt�La���f�z,����FW"6<?��LB0���J���߅2'Bͅ����gω�h��K��r�X��⟬�	����	ȟ����ޗQ�&��/`�@�N�?��?闲ij�T��O���~��O|��v�� �>e����#_EZ����i�Iɟ4�i>�	������'<NQ�& ]���%£K�r8#�P�G����䓍�D�O����O��D��V��4Q���b	8��^�[y��d�O�˓b=���� F!B�'�R_>)
���z��&!��x��##?)V]����4u`��#�?�bb�h�U2�΍t$��A��/����;C���������g�|��
�n�l`�.W�Z�1#%JIj��'�b�'����T�89۴x%��6d˻p撔��힣=uPhH��H=�?��(ݛ����v}�Jo�TD�����j�4}珌�`&�<xX��7���%+�B�Ǧ��'"�=�D��?3�Q��X���2Y�}k���&�\��c	t�<�'�r�'
��'�"�'��_��dS�"�<8Q�9�Q�&?�,qܴ��@����?������<����y�B_� *hm��@
�*���i9���'FO1��XK��|�T牬V�(l��U Z���<?�I�q�Xm��Ov�O0��?q��fh^DS3�ڋq깠�H�m�L����?���?y.O�n��L�^0���L�I�S��ȹÀ�{P�`#G޳*���?5U����~��*ܬP�Ӛ�! �ǒ-X�4��'(pC�d�ǩ}���4$�ϟh�c�'���¥�¼q�Yڂ�W��Ȅ�'��'.��'��>��I��6E�1��_z�D�pD�K��(���M��bő�?����4�5�jX�0�RH�E�D�[���14O�$�<9n��M��OJT�+[��µ��5{��dyt��h�Ƙa�/19x�O�ʓ�?����?���?	�D����bQ7w���j�F\�rڈ�0.O�9nZ�� ��	�D��{�S�̡#L�95'�q���.؜Hc���$�O`6��Z�)��� +��(P�_%�P҂Fc3@u-� �n�,�̸0��O
D�O>�(O�=k�W&2��G��l��,�O��B6M�O��4�.˓5l���`��8!��R�Ό1@��ipA�,ZnҨp��㟈�O����O��$ۛ%<�0F��z|lYq�NM������&l�@�4����&�?�'?i�ݲCY�����\�@L� cEJ �X���	ȟ������I��|��I�'C����mû]�P(�'�f�����?��NL���2��	��M�L>�CjNwB89����{�ph+6��L��?)(O]b��z�4�?��T���=Ĵ����J�;g\-j
��=�䓬�d�O ���O���%Pl  G\9�Ԉ�"��-X�$�O��Tz�F�A�6=�'{�Y>!2�$�(B<�g��?y���#?e_���	R�S��^P�I��+@<a'2x䪊�s��H��� $g>г�V��9�ϊI�I�(�d��c�~{�x�#�?�����I��4�)�yy�(lӬySWh��	���d������N�]�����O� m�`�F�����0+�6���F��=��X��ay�#[�����h�Q�@���O8�̕'"PA:�#���4��ǗX�X��'=�	蟨�I���������t��N=kd�d"5�*bȅpůE]�6��[�����O��d'���O&�lz�Q��#Δe�I.]�/NJ��!��M���i��O1�l5XC�d�z�	5��] �SO��@hN�'h��ɴ
<��'�4�$��'<�'�,���'qo|���![
�KE�'?r�'"W�8Hٴi�vI���?i��3IB䱗镡}Dn�	�G�(� �2��>����?K>	�
�@ ���h	O�`��{~Z�Jp1gE�Mۓ����J?�`΀i�֪N .*tAD���
���9���?����?����h������|Y�-B@�X�V}��×1`��D��W���x���Mۏ�wX�2R���\�w��L�؟'��'��.w��&��֝ �N���9� {��A�;	^x�OI�.�#J>1/O����O~���On���O~��P�9��ʤ��V8�.�<q�igp0���'v�'y�OwRl͕�P �!��-:�$� ?W����?�����S�'~����$	<7��+�T,���+�M�S�P�Ed��&��$/��<�'D�0����OU�a��q��Β�?A��?����?ͧ��ĝ̦M�pA�ٟ  � 85k��BǷ	m���B�'��6-=�	;����O��dA�ݰ$�ؐBI��ڧ�0U�pc�O=N��o�|~�i�>.*����䧙���Iwּ)ؖN�/0��(��\�<y��?��?���?ُ��i�2�z9h1��/N�>��N�e�2�'�2�uӐ�򠬳<᷶i��'���Z6G�%Z6�#G�BK�Zu��*��O��4�<x1�Dz���XU�-c#j�+FD�{�b�� ���H� Y�8�,��a�I]yr�'��'6�F�����S�M�+z*`ؐ��=%H��'��	�M�1"������O��'�X�Gg�
 �-��c��2A��'eL��?���|u���� �]���A'dZģK% x\���$إ� 1�q�PU�����IY?�J>Q"��?42�@!)֭m���"R<�#�i�������M#��3hH� dP�pTx��O�(oZ|����� �aD�^��|����.jP 8��П�I2wH�lo~Zwު@��џ��]���Kb�\�9�*D��D�D$>�̓��$.|O�i��-H��b"�F�$
���a�֦1�3�C���I��R���y���=5ꬑ3!��7�&9�N�]R�'�O1��i��Mm�<�I2��|��튜3,����W`G�I�j���!��O��O�ʓ���W~�3P��m���N�2ax�h{�Pm`���O����ORI"!�Z?�h�6�
�f��#�5����$�O���Js�ɜm@��;5���f0@����<,�A=f͈#����M봓��&l?�����yA A"aB�CT�¡x'R��ȓ�T�[sDJ)7>��36I7�A��.w�f�Q {���'N27M+�iޑ����� *�)4oZ�dx�xp�k���	��H�I̤nX~Zw�DPݟ�����=%uNdcV�PD�� �D�<	��$	u�H��N�e�8�$��3R���
�M�4�ר�?A��?���EB� ��DXq�����j�����ONal���M�b�x���&H'2�Je���U�d̢�y�گ*��d�P�'7��I�k%��0J��o�,`�ƨׯ	��˅$G����O�F�l���V�]ᠱ���8 r� ULͣSF�8Տ�6� <�¤�j�<���[�i�pQ���&"X�A�J �N�ْ���(����������/T*f4�L[�'��� '�N.�@���[
dF�K&,�z�Ԕ�طV2��rWeɹY���g�����dI*}I��{�+��q���ѓ	ӡzZhT3�cģm�*�y��7�mJ�_�CxdP��l�f�pX�w�c��EZ���#��I4v,��Z%͊&b���0�N�TF����#G+�9�4l���%K�.Jj�1�&j@�u����xr�'��'��<H��iL�f�Ū|5��'͂�g�8�'
��' �Y��p���ħ�pa��q���'I�J%� ;Ѹi��|bR�����/�	�C󠄪���K���R'A*!/�6�O�D�<��͡S�Ow��OӠ����[�
��%b{��D�3��<9�f�`������J
	�C�̬MR�@���>\��FY�����ǥ�Ms�X?��	�?}��O,����X��`��c��PA�{Ӣ�{��QEx��t��!E\��wF��Gz͊��ֳ�M�r���r��'���'���">���O�qf%G���C���U�`D�4�
�	r�9�S�OH� J<@P�)����fu`Cf��V(d7M�O����O|�2�
\l��?�'���Q�&k���k���.x�ӌ}�(���'���'��G8r���B�G�]6�Yj��TmH6��O��˟�I����� ��5v�JuE��S���{�������^ 3*1O����O����<	��N/]�$�A�(�/�� �sZ𒳞xb�'f"�|rV�$�./N�H���Ⱦ>�NaxS�*�b���	ş��	^y��tʮ�S�wך%�5)^܌���'5L��?������W�>��������
 �x�$����	H����?)���?�,O�1�Gd�Ӭn_�ٱQ�%Uniӳķ��ՠ�4�?�M>�)O,Q���d��8]dԠv*�5j�����/ko�F�'��V��%�B&��'�?���(]�ݚ�o�"�����*.pj�x�W��x��0�S��r��)ƋrRL�X�J�n�Sy�$��>6��o���'��D�#?Y��@^'vPy�.Z3�����Ŧ�EB8(5�'}=:�wɩHСm�/B��D�Iӟ4�'�4�'L�T��q #X<�U��V$���x�$=��DM9PO�b>��I<�^�R�aV� ���j��Ӆs�((�4�?���?�զ[���|���~r���2H�k��j���x"�U��#<�G��T�'|��'�bd����\ʐ0P�m�V���Á�>#�ʒ���<����m�����d؋'�@dr��
�*�S��x:��$�O�d�O(�d�Ol���w"�$P�)@�h�" Q�m~��O
�D�O��D3�d�O����G�jM`�a��#��-i�NNm�7�v��������Ο`�'����!q>�s�^�!��e��;�b�z�$ʓ�?�H>���?�QlG�~j�����9��Ȧ_��ykC��
����O��D�OT�B����[?��ɥ�H�!w�P*�L�ĮW55�����4�?QL>����?1t�L���'2}p�o�8��򲨎�'�8޴�?���򄙝���O���'�����mR�5z����*�d�9R��=�fOL���Ob@�ӯ*�	e�!)�	����Ǐ��
�榁�'�)h��p�v���O��$֧5�ϟ�m��<��H<U8���M{��?iw$O���'�q�fȳWA�.�p �7�^�sP�i>H�	�Jw�*�D�O������'�ɱ
􌕒��,"���h�b�V��ݴP�Z�������OQ�I�0)#��"J���ڝ1�nU�$F7��OL���O(i �$h}2Z�T��~?!�"�-��Y�A��-j�+TI�0]��M>����?1�X���q�Yyk�E��!V�� �i8�H=H�든�d�OV�Ok� ��f�Ջmw�`pD��L���PY�P�C�B������̟x�'*N��$-��T�&�
�,��܀4a�aP�O����$�Or�O���O��K�'ڶmx�qh�U����W"j��O��d�O��$�<�[(J�i�7t����Z(d�|)[��0B��V�$�	b�I� ��78�܌�%��AW�:��(��
p�I�'�R�'ER]��IGҤ��)�O���%���(�9Y�J{����Mצy��t��̟|��*LZ���^�d�x&y=Vܶ`§GE�g��'�Z�� X��)�O���u��e�:��(H"�4z�`9iR/]x�I���I D��l��q�z�"��yVH����3b,�(�O�𦽗'���fӘ�d�OJ�����ԧ5� M�+��m\�e�d�)!ʒ�M��?��ê��'�q�����g؈h�b�U�ݺ�iX�)�a{Ӝ�d�O,���a'����(]Z�b5r$�� �7B�=��4I��@���?�*O(����O��3��+:��8�&G�S@�I��^ߦ�������	��x�K<�'�?��'o����:>�=C�TP }��4�?I/O�,��*�F��'���'�"�8!�|�$��W<
hGᖗ&!�6��O�,PኚA�i>���u��3_W���q�Q.5S'Ů
��5�O��h�i�O,�O����<a�G:�0d�>f�T��Mȃ2���$�����OF�D#��ȟl�ɝ|f '���[��i6�3	�b�3�Ǚ���b���	uyR�'�����ޟv�ca��3�,�jǌ�);� (�4�i6r�'��O����O� d�/b��j3,Ѥ1�q'٦Lx���L ����O��O �:\^ �������pl���l�!�`P�0���B4�7�O��Ojʓ}�"5�����<v��B��(랹�  	%A�7��O��D�<��jU�s݉O��5���斀�S��-L}���gj�+�M�)Ol���On���O��Z��ƶA��OR���J�#�^�!�i��Ib�bB�4��韄������ĵ_���Pi� :���4�Ӎ!��S�4;B�ퟸqH|�K~n��q��
Uܙisj1隽=�6�~���o�̟H��������|:w���.��e��irv��Ņ�<n�������'���L�3?y ��Q~Xuiv���)w>�q�̥W?���'�B�'V�̰�Z���I���c%i[�������!+�	��y��	��pb?)�	a?�2�
aiFy{$����b���ƦM��>U�f�'0�'��'W����A�?9lE��/V�Vn(��"�>i��"NTH�'B�'P�V���ePZ�@`b�d���$��v�1M<���?yL>�+OHAZ���T�蘒s��Q#���$�6}��$+���O˓�?IǄ���Į�0Y|�P`&O٨2�� m���M���?�r�'��?UL�4d<T�w�M¸����O�Z��-�'���'&�^��:4l��'�<�x���p�r��&���J��i/"�|�]��`3�\��`��Z��"H�Q|5�B��� f.}q�i �_� ���%��ԔOIr�'N�\c�v�A�	˪n	�p�pB�4��=�H<����?!BX,MWȜ�<�OV�y��'��&�$�	��Ǌz�x��O.�Of>4���O��D�O@�i�<��x���d冺~{�`y��H6���o����	,
���21�*�)�ӧ?��#A��1�� Y$@6M�!t|el�џ$����h����$�<م@�2��(���|s�Șb:��j�4H�(�Exb�	�O�ȈU��r�L���,�d�F���y�	�����K��خO��?��'[T�s@{����L+}�\٩�4�?!(Ox�rA;O�S����	ɟ�saS+f5�%��Ղ:���3���Mc��@>����P�`�'�^�d�i���f*�*{Y�ݸ�K&$%PKaj�>�+
�<9)O>�d�O��Ĥ<qfŉ�.�$�h�HR�&IreH�� �+Y���'�b[�����|�	�oFX����<a�F�$-=<�f �&!?����?����?�/O8�+'�|Z��^L���t
§s5��1�Ç��'q�^���џ���4f��/��Z�k
�D��Z��4oZ៤��ҟ��	Uy2�"k�R맯?!�*�Άѳ�ʛ\EtP0e�7U��6�'i�����؟t
�&h�0�Ij?!��
�v���-��	�Ŏ�Q��şp�'�r��p�~����?���t���5���Z%���q�Հ*+BU3�V����ΟP���2/��m��'���A>Zެ�B�W&��e,VbA��W��K�����MK���?���d\�֝�1����6*�l|�s#Q�b�7-�OD���'g���OF�$�O��>��^�b{3`F(S�@t� �x������̦Q�	�����?]��O��K�da9�.	0}ML�f!�&�L�Һi�4`�'��'�����:���1" rf<���'t��m�Ɵ���ؘ̟@�����$�<����~���o
�qHM�0%,��Gc[��M;���?���+:��S���'��'.�)��Ar�`�@��W�V���}Ӽ�$Y�"����'��	Ꟁ�'�Zc?: �3"������L�Y꼩�޴�?W�	�<���?����?Y�����8Q�ѨB�Kr����W�
�0a���M}�U����Iy��'���'G�X����W��q�䓿Uh��$��0��'l��'yX�����������"ѡ�k�02�x9T���Mc+OD�D�<i���?��&l�}͓5 � �8���)R���ԎY8 LB�X�i��'�R�'j�	�5�q�����/*> ���[�9Hִ�ǠG���\mZܟ<�'<R�'p�B��y��'w�$8(��k��9u��RG�D�wH���'�^�T�)���	�O������芷 -�F��E�?f�QJG)�x}"�'c��'�X�q�' �'"�i@:f(�,I*{������lo�VW���c�F��Mc���?!���*�X��]��������7�(�r�.6d6��Op��#!��Iyb��S�d�"iJ��½qU������&C��	��M��6�O.���O �)�S}�Y��;��1� ��AAE��(�*^#�M���D�<�����8��ퟬ���0p��Jta��+��Ѡ�M���?���`�4�S���'���O�������Ё�+9S��Z�R���'Q�a��O��O����O6ę���pA��(WJ��4��Ȧ��ɴZ�H)+�OL��?�.ON��ƴq��'Z�l���`w�\?�HP�Q��s�e���	ҟ��	0��Hy�^�h�p���O�aN���N��v�(���f�>1*O~�$�<9���?���^�0x���"$�(ac��2�ENF�<i��?i��?���򄋍c ���'@�h���FN{V��W��#�n�lOyb�'e�Iϟ�����k7!z��paN�ep��NQ8	�����m-��d�O����Oj�m�~-JQ?��I�e� 3�U:��`�H�Z����ش�?q*O��$�OP��Y�T�1��&�� �a'�[?P�����MK��?�/O�����WF�D�'7�OF4l�Ф]���$A	�K���XT��>i���?A��M�,͓����O,�S�h�d8rV�^���R5o�j7�<�Ü�#����'�b�'���>�;U�^(���^�;Ԧ�����
E��n�˟��I�LA��w�	tܧH5n�b�m��"B�W	��8n��򴽨�4�?��?q��kV�	Zy��1m:�U�bo�$4����!�q��6-q��<	����O��X9o�p#L��v�@ڄƐ�(�6m�O����O� �[쓈?	�'ޑy\z�D�Ժ:L�'��b��|r:�yʟ<�$�O8��̣?����"��'kT,��Q�F'BaJ`m�֟��6��;�ē�?i������1
ٖ)r�����C.�\����Q}B�D�uV�4����@�	XyK� a6����`�0�;G��1�N\�3�$�O���?��O��E�p�,Dz񂕟WWШCg�9���OP��?���?I-O�th��|�H� g���)N��>A0@SK}��'�|��'R�ܫ1��$M�_[�SL�	=#�A���Z� +��۟���̟ �' 1!	$���>(��9��Σ=ޢ̫&b�%oZ矜%��	矐�n}�P�O0|Z0b��H����N%w@���i52�'~��uM<�I|z����0b��J���iL$e��Y�J}�'�R�'��
�'��'��	�a0h��i��B�)e�Q1�&\�`�Dg͚�M�!P?��	�?M2�Oy�+�.��Ul�n��q��i��'��@ُ�$�|z�'�" �4��+( ��e�V�fc*��4C4�3�i#B�'-b�O��OP���ezNy�SYrҘ�q��2<jN�lZ*���	[�i���?I筍�"�#F{���H���y���4�?����?�Ef� #�'>"�'���vy�R7��FP ��Έx���|���yʟ�d�O~��]U���r-P� ��ɷ�\�_���oZӟ����!���?�����K� H/T��u�Љw `�W�Dz}���p��'FR�'�[� Z�bÒb��� Z&^�'"�dE4�2N<��?M>	���?afT�C�t��M4=~$�h���6��2���d�O����O�˓6YjE+�;����1�0D�0mq��VΈu�2�x��'��'���'u�(B�'>��BF��V��ylK!�4�"�>����?�����$�+�l%>��3-�3gz4-K��U��d�]�M{����?q��;C=ϓ��g�"�#��	�L� ��P��7��O����<�
ͳ<��O�B�O�"k�*�G�,U6Ƃ1|��t�2-=�D�On��%R��1�D�?yS��<���V"+���0�|���0�X���ib�맃?��V��6F>��$��\��uQ��O�q֘듩��O���(��Jd�����x0�3F�iR]�@u���D�O������'��\��epU��=�왑�oK?M�i��4D����?�/O4�?��IW~v�K�GW-d8*F�L�&5�4�?)���?�bᑤ��ICy��'&�$���h�*sÈH��b��[ϒ�mW�R]��)����?��-��}�%H��MX��*����p!y��i��+	�[]:���D�O�ʓ�?��?t�8�0��2xA�T���;���'<����'u"�'Xb�'MBW����L�c�]�5�/�r��#	��"�O�ʓ�?q-O����O��� c���d��W����Ë�3Y�4�A>O����O����On�ĸ<��m�?ym�G�Vy"���\�XgJ����VX��Ǧ�'�R�'lBʃ��y"��c�p�䄜�6����P���
ꓻ?��?9,OL���f�y���'�p�Q��  ��5�v	��V)�	���d�<����?��ag����?��'ᄽy!�K&bL\r��Ql̡�4�?!���D�<p���O���'����E<m5R�J���jB�U#`Ŕ�{����?���?!�E��<i.��d�?� ��$BA$%�Y��ޯc����ճi��ɋ�|pߴ�?����?9��~��i�)Y��S�U�|9�-� ֽ�`�s���d�O\U2C3OB�$�<��d`�7R��1)���QԼ���ȃ��M��bٲ�?���?����J���?+�<����E����b��Ŧ`rM+���c}�+ɤ�O1���dG�FxUAb��u��g�����$nZ��T�	�fP+���|*��?!W��'�	p�H���]�"�f�O��
w��O����OZp �.�j�@Is�F�*��'H�X}�L[['�{y��'7�' ��:&a_ C��u� 
�4w�yS�c*��ˏ��ԟ��ID�'u��B�̉6ղ�3u�ްPi�]����.8ɉ'�B�'`�'�R�'(h��%Ǒ�X��Mp&�ϒ���S�ѕ՘'���'$������$M�| Mډh�*�����d{�_�I�$�P�	�JEf�>�c(JY�n��7��0�dG�1�ꓻ?q��?��O�Asa,�IJm�L��B�P�,�Ƞ5�N�mʟ(&���Iʟ ��*,�	1rl�pb�	hߚ�E���T��7m�OT��;?�C���ħ�?��'>V�е$3��F�"\��	A�xB�'D�H��OD��08R"�
��9�큃�ɬ&R�6m�OR��Q�q��d�O��D�OL���<�1Hg8�@ "�3Qx��R�']�.
�lZ� �',�B���4��F�b}���ɁU�~�A�$�M�e&,yq���'f��'q��@.�4�"0����
i��� �eP.q
�І��Ǧ1c��s���<��+\�x$��e�lY'* �v�qT�i�R�'��j�81��IL���'��d�)��H�R�E��dx@���`Ex�/!�������\�Y6��5���A�c�d��i�V "D����*9��:E��;a�y��!:\O�)�Nr2\�6/�|G�d1���`\�2��Β�OȢ5x�Hc�Ǎ.��9��?k�|�C&�3m�@b'D�%�� IŸ
���,V�<�^�p�HY*Z�%���<9�
�j�n�I��� cg_���3SnS�(��0
��]C����}�B��N]L� t�ϸV����k
�?i������?�O�ii���0i���+��G�>i�f�����tC�S&�
t��#?���>,б�19[d�()S�6_Є]J�¦3�0(��ǸuH�kvjU�^^䠣�����?�����4oH�Tഊ�!�A��A�a�1O��d�' ��#�������ݞqP�O��m�o亰����t!�Y3��/9\�	}y�f�;!���?i(�iq�
�Oƨ����"�H�ƃ��h�bi�O���C�D�M�1�,,��h ӟʧ���Go�n �eI!?a\@	*��j*q��!t$i�#+V��H�"� ������!�BeP+uѾ�r>y��蟴��h�O���A���D�ͼ48�@U唤�y"H"@1d��r��	���0<��鉂�$z���k��dC^�.��!جO<���Oȩ@�I�@2���Or���O���R����O�1G�Kv*�"v_�Y+�(�4'����)S�@���5�3��ԼF���ꖍ	�*��A+uB�Uj��X�D��I�^��#$��|R�ޕD�н�晥m��aAOO,�r��,�0��O��:�1��5/[�g5|��'6		xB�	U;��i�����$@�C�u@�PƑ������H��� ���A ;IBMṡf����O��$�OL��;�?����4���u���4�i��)�(Хdڲ 4j|E0K�l؞̣�j�$�x�
V&Nr� AGn�}�(��ϖG���'��t�8���@.p�.� ��X&F+:�⅃�g�}kG�'���IF��C���{�"�(<�,I�K�J���xH�U��"|d��X��*x�N��<�E]���'�|)`�z�����O�-�򈅹��-�7B�g��]����Ox���#2��O��S(+²�3���]��`����xb���P�x�%��' *�k��;:4|J�ʰ|��e�����	�ē+T�D%��9�A�D皲1�ȓE��ULU9.\�}�b�R����:=�&��s��5PjS!BH�xo�$[��'9���6O}����O<�'lo���G�6ɣ���Z^��X'̘'S.	���?!� �A�P�B���u��I˳K����|ҡHװ�e+��D��|4RW��l�DՒ4rAiUhzO�Y��-������k��/mB	��`����F��I1�~r�'��>a��4�J�J���i�4�)%'B�	+QXB�������&h��Q������[�'#�U��� `X�|I�@<[�"�'���'v>�;�Ú�)����R0?h"�+�'�8����³
Ӹ,㐪2/���'q\}(����V�1`$[,e����'��)��ϲ��5�皻�F(���� ���9P���� IDx�U"O�!�cC�IRteN�Z b5:�"O���(�*������2BJ�Ѵ"O��A��P�%��m���R:N�#"Ov\[�f�!P~�ia�/_*1D��"OB�1�Az��r�	}!XŢ�'�jlJ��\k��9@��%���
�'o�C3o_.SH9��h6QӠy�
�'|V��t�ש��4��`J
F��PC	�'�@U6�+{�ԀIa��6���I�'�D�G	�+��j��&�y��'��E���h9jl	u$�H�� H�'T4�Woϩj���".��L3�t�
�'�["j�)�`��@��ع	�'&U�cb�i��DȐ��]�	�'h���7h¯]��Z�gN�t�\��'zd�HCi��r��:74���'���7%��X;�u(@hͧ$��a��'�X��i���TmI�(ݐQ��
�'k�A��(��h����BLQ=M&���'��X�	V�kQv��MѼ+G�m��'?	ɶ�\%��)� G�� 08��'� ���E�:O�*0���OW�ѳ�'IpXb̗<F_��Q��J�J#|�:�'��1'�)^M��J�g��G��̸�'��i�_�=-�X���݀'���'�V���>r4�� �׀\��'��ؐI�~���B��/#�'�@��6ǖ�ĸ�P�G�#¬���'d���t�ă%�8�y�/�G�R�c�'^<��E'��c���FDX(�'V2���؀�xJ�#O�A=l1��%��hɚ-x�,���0>�2�+d��p��6�Za��n���a��Q��H��Nv���t�@�Cyd)��#��
�D�3�!���0j�a��+��Q������%�1O���@��'�-���!�0'��
Da�qJ��5!�C�I�1t�3E�޸1`u��.�"��[Ç:WL��z3THG��OF}��'�"b�K�GD�$%��e"O:\B�Lh{��my��D-�hŬ�'0��\�A	ڔcha|���D�f��"�\4���&�0=qE	Oe&
e�d	��<��"K�K�����R�S�\`��YB�<���ܵ<C:k�)8����s�<���C��1��}G���qB�h�FĒF*<�]��yBF�l���Tm�?U|J�*g-։Pl$���ɘ����[��>�kE��H�I�Ic�3*�Q��=G�A�*/-���6��-[����&��ђ2��H�,[1�?O��T����,x�^�2�J0LO�q:�n>R�F9�8O�qڲˑ�&���Pf�:X�"Ol���'N�=J�E�F�'R�<�[��D�%V�,��=u?]9T�(���N_`	�`�g1D��[�J�O��hR�K�Ji>���
����d�,?1�GW���dS�l-������%
b�	�Fש>!��_8;�F1����T�,9��ζs*!��ѕM��6eC�q=�Y�vi�.B䉲"�J���F>�i�f��+��C�� (�B}S ��{f��IE�%"O�u��Kԏ^��S��%Fm�`"OZ� ��	}KN�KPK%2�&P0�"O���'Δ�-�>������`>�xr�"O�p��-�P�'䙌X����ȓ1'
�3��Q<�X�/�c}��ȓIy
����F�q�^.�*(�ȓz�rh����5��phW�}����=9�'�;�j��IM�,�*����c&ց1!�� �e˔e��M�&t³�>F���M@�٦8$�����<i��1-�aA�T��'��A�<V��)K���� 8���i�� %(��r������	
t!Dۛ;��@V`M�U�����ݺ}(�!(���
r�$8Cj-��D�>��<��� y!�D��4Tӄ)݂t��| �k]1S�1O�}�gE3$tm�#ESU�O�-�c�!����*���'�rq;H�I3�������xb�'�AY�0K�>���K���d����pg��E����u�F��� �X�F�3Q� �J�oP=_b�9��Ϳ�N0�ʚDԅ�Ɂbt�u�1mN�]�0I�V$Ѷ���	�J�EZ�\p�����PzZ��u�נ#�Z�8��V��u���,4���  \�HDH|�� �Ha�0�&?�V	�d�����mX�7؄����Oձ��	!�M�oq<=Ap\/mr80)4"O�[4����	��o�9u<��s�!�%S���&C��ox��RE�3�1���PI��RTd�ɒ�C�#�5iЭɃ�,��PRh�*qq���G�$*��s�	����Q�kC�O���rC�j�n=��'���ja�O�Ct�U�^G~���I\�m�&`��'n*�yt��("�lP3�(|� 8և
"g�9�D�!2�z�)q��)����O�ZW�3�p<i�-��!1XI�s�	}�����Zd~�v2�i��͗�(2��1,	�Nq!!��6?��$K*=I �1U�ӳ6&t ۠��(��TӓPy(<Y�
��fo��Z�G�]�]�C��m0�i��%�x��Ӂ��4H��&��I�}�\�O���K�D�p����ȑ
�(�Nv���
�K
�ʸkWK.$hQC�E�$:LPBC��R� �sBf�t�	-i.Z����a�T�k,�N���/��w+R�,�`�b�Ƥl#�yD{�I�+6rF܉$S�IX<ٻ7%�8�y"��hY}3��(m�~��"'T!����7(�����m�B`%��1��Oȸh%�ܒiC��3a�3�����'B�,�0S�P���2U"�mH�k��)ð�
7i�>wm���ą��U*FR�߶�G���e���[�2�$t��'�������ģ��2x�T��  �Y�r\�4�'�>(���B5MN���'�|��R��.�	h�~�)��P*K
8 wNN��a~"/_���A��ݐFn�a��\8���",7Ph�b6��Z�Pj�jy�̄����nBBq�l�}P�@��ސ��`�0�R�F}�F�7@��e�W�lͦ��"�
�?dI��H��� 	D�<|B�K���@�MJ��C���t?��`A2�;�H\�KJ'��@Ye�Mvzz����29�P������ν ����'�V�iי���ϓB�ԛ���m��q��a��=+�69zԻ�G>r�ԥbAf��ja��W�[�p�a�AL�M�W�Q���,OB�"��>�t��B�cwd�,m��Y�Q��ix�x���ȫ��p���B�N���S �>v���c�)h*頦K|y�� ��B���	@�>��_'�d�2�D�ƩA2Jb�'��ĨW	Y-1��Ѧ1�̓� X�>��)"��|XX@A��2FЖtc����	&%�,�0�'�v�&ƈd �k"-F:�ι�hr���P�fRb�a�+Ev�.֨X�N|��7���4e��F<C��	+1�>s�'��L�DC[{Vh��*�[P]saۤq�4e�1o�M+�f#�+.�Ӝ�4�
7�>�ĢLK�����G@I��GH<���\1*�������N�����H�XR��V���YPZ�� ���:䀈a)5O�Ţ���RjP���n�:p{l���'���P���6;ր�gk�8Ob�Y��U�$x�!gL g��3��5�X��(!�0�S <Z�d5��R3�A�O���2br%fQ���D�fu�O;��)Z���!�"�%ҳ�=o��B�	% ���:G��=�r�ˁa\/^�Q ��X�3
����Oz��v�3?�����f��E��B�*L�p�����F�<�U!�)���d?�B�(��R�2�Jː����&$\Olً�	л��p�%�?����B�'�r9�Ɨ�zHh#c�NM��U�H��l�n���ӨJ���{�'!��TH'L\u���`�1f���'��h0n�6���P@G�O�>qig�"�0t�C�9� ��'t������ {�d��f�<.)z=�A�J�o����A�~?I��An���$֯}��=I"�*���:e
�!�ʱ?v�Wd�K(�a9@��!<��y�kת0�𹀪
��p=	v!ХЖ��ĮB%wj|sQ�^S؞Tj��^�/���i�R�K�uұf݇w�0X(c�Ej�	�'���%�F����Ҁ�Ly����$�R�=�5!:�'[�؀P��N 2 ��#$#?����6ޢT3Ѯ֯j>X�wNOc;�ulZ�*����?E��t�? lt� �A8%|k��/~�}��"Ob�E�Ͼ#qV0Õ��hw$�[�"Ol�`_UX�x'����T�#"OFm)&�l��(��zu��["O.��ѦV����n�o��4��"O����L˵v�1��NP�j�b 3"O����ɸC���0�$����#�*O��)��Ѳ!�.���&Pkw��A
�'��Yk�0D�R�p$�s0n��	�':�k�
{�8���M��sL�@3	�'[�����Q֬%r��ڙp@<���'�����H�.��e���(2���' �-H�(	�Y�|����4V����'�lr�)�*@kRe��l�=:�T=��'4���X�"�@��l�Fi�,��'C6�0�	׻4] ���9���J	�'�L�3o(	s]2�ܩ/�4�	��95�F��>E��GψD�����H6�j1%�cMB��S"���D&��y2&!���Tl��|,r!D�2�Od�S���4H�"��eI	>=u�1��'������<1`n&%4A( �:
��I�E�<�'#u�����?�@�ӂ�j�'%،�#F�O:M�T�&�� ءN��*��Չ�'���#�ۗ~;X��!.ְr�M͞97�]��{���'��E��;|�dy�p��%�����eD�����'�v,r�nV&&4U��'U �ĥJ�'�"�p!��F�'�J�Ĝz}��U��;SF@���x���p>	cF�F ��ɼ j ���� `�uKW�h����ʗ�֐}	�?Ii#�,}��< A�8gt8�'ʓgU`h)�1�]X����21+��)>�.0�E��qO�}��rY������%8��zDJӚQlڳ�c�}���i��{�AϓS4b�0��-6$��'�y�#'�O�P���$J�zh@&	�K8�r�"O4�̯_-
d����#4Ȁ�$"O:�1�c�s�,3�<j@�bv"O�`I/ϭ/�H	w@,��1'"O�Es�\5�z����6�d�"O�!:�Iݡ(��]y#�P�1H�Z�"O�Y�$φ�xm"Y� J@��a8�"O��a��S��3��xLeKV"O�����(��SoGp��6"O4����־ݲ�>�"O��I�I)u��)�V��l�h��u"O��k��U)9h�r�aH&Cl��"O�m�$mJ\�T�K�/����|�"O^ՋE$E~})�@�;��2�"O� Y�j��&Rf� Mǽe�"�s�"O�|��-Xp�b)դL��P!"Ojf�N� Or91iN!q���"O�-r�Ge���f.��|g�E:6"O]�0�7b�dA!f퇣Iv�`�"O�d;ѩ�0`In�إ�h��BG"O��A�b�>��@��@�8b}��"O`(�F� rЬ�f �M1�л�"O>-2�Gǔ�<��D�ӽZ��,��"O�(b�.ݠJ� ��чN�Lx(0`"O���艶3y��kA�Rm)��K�<i$բp6VĈc��B�`c��I�<I�� l0-ӠF&"����'�O~�<���`�\�Pf�%[f� ��z�<�3c�!z �xb�-@�֙��L�<y��B1ǬE2��Oqx�{�g�B�<�AR�fH;c"T� 0!ꐧ�i�<i��Òw� ��C�5L�-"`�k�<� ��C��@��%Z��ϝtt^-��"Ov C偧�؀S��A�Y\AI�"O��Y����K���<YzY��"O���6�Ԍ����Q�X�,)�"O<���e>\�!�0�L.~=��"Ou� ]'S����@�#4��I'"O@��c$��Ts!D@�䀳"O���q�Хd��4�G��-D��"O
���-v �O��q>d�"O��*A�^����`��P���bs"O�[�l�;#����Є�"1*��0"O�� AR�v�|���Iا"O�P��e�h��AC�)�%	
T=9�"O�5�N$BQ��K�Q���1�"O�X8�k�6w���(�-X��Ĕ"v"Op��TK�!zվ�@`���fWz��"OH#�����9C��RTY�!"O�Ȩ�`A@E35OW�h?���"O�	S�% | j'��!F;���"O
�Ҥዓe9��:���7jpi�"O䲶�({F�𑠥F�t �9U"O�=��K�<aJ\[��ϸy@LCE*O�ĮQ� Y�I�τ� ]B��'9ހ���_yf�[6+�5w�F���'G�=��`N9W�0����r�%s�'�,��N
/�TPY�&�8�6�C�'m:Dc�EA!,JI� @Wc:	��'`j�Jf��-2��AC�j���'���
�o�	Diڔ��)_MQQ�
�'\��xV�������nB��	�	�'�L�a˞��H�`��8j&���'�j�eA�,����G֑EG�a�	�'p|	�#k�>1�$x��@FO?��''l3feD-�\i�6jۆ@����'9R@yvk��!�\l)�h�(<ڸ	ӓ��'z���ŉ�)G.ኂ�F�,��'Z����  wp�B݉
Z���'���D6d߲�*2�پo!����'�ʈ���'J$:ԪA&�9n�2x��'�@���B]��0���i��i��'%���΍q� �����d[P�	�'�T%1$�'K��m균��LKt�#�'�d)�싒_�hxIW��*:���3
�'�B�K/W�� ��a�\�,5�	�'̸��el�^�Ul�$r(Ԛ�'�l�g�̢V3B���A@P�bX��'>\�_o�T�և�S��u�'nXP���%{����c��E�����'���ACh;f��Da-7���8�'�z�3��C�`�%�S�ޱ��̩
�'1=sT��cA\9������i	�'}�	Ӓh_�}^�Y����`�'�p����а1��UQ�z
�x�'��J���s
Z��,�+\F����'sR�[����,m@�K�6(��b	�'>�)�afV�}��H�q_�=r�'�I�ßMp�*��4cZ��
�'�~س#(�L��Q�툛3� �'n�re<as��w$N*/���
�'����Ej��B���]%��8
�'zd3�n�p�Vy9u�]/��t�	�'#Ca�=M�p-P� L�We���'�P�cW
�\�H�#V�H�:h�
�'��@#�/�1���5��!v26�;��� d�Rc��r�|�kʟ=P�0��"OMI5��K�)�G�;��L0�"O~�h�oX<4���B����}�"O�1V`\�g�4�c�0a��y�"OZ ����nH	ԈQ���bs"OZX��b@�}����!G8X�6���"O�-90���T��'�Pp"O����&�7#/�B�,@7'Jh:�"O|t3BF�e�Ҙànуn����""O�y@ǁѼ"`�c�,W] ���"O;np^)cq� $����S�H�C�!�d�)E:����G+0�j���$��%w!�$��X�ɰ�"X�\�jT,T�!��q̖d��O�g�
1K��.L�!�D8��anF(���IF�_��!�d�:d���"����,P�)ˑ@�!��0:s��bN�b��|�b�U*p�!�DJ�ɑ�T�.�R�S���@!���HM�ak�G]�[��ؕ��s�!�dǈD�с� \	���c���<!�y�8��,X�d|L���N�%4!��az]K@C�BQ�|�E�
��!��4~��y���1V4���7j��e�!�Ę�Mh��V���ʱAr(�W�!�D�E��щ`.;3P��t�!z�!�U'�>�3�ʗFJux�'��!�̆nL��Q��]�87L�+�� 3!!�D��<��yTቝ08�U���==!���?[�� ����>+����Dх!!!����s�a�,h�!!�n&�%{2,A�v�!2g���!��<s�ibQK��?�~0s��V�!�D�&���Q�OW(=��R��T�!���1.��qA�6Q��1�mS��!�D��V�P�+ub��/�L�I�M�S��F�)��e�����Y�@�w,�?Va���<�O��O1`�%�	�0�`�Ň��.!(�"O���0E�
=B$�J�΃:\�h%
��	u�O�&�B�lL�<�e䃹�� �ȓ���a��WB#@+�1<��ȓ"��B�J8�Kt�P�z���Sd�r*סwf�Q!"�M�V���D�@"`$hdd	P#B�5�ć�xN�Di���u<�[WIZ>{.L�ȓV|����F�#>ĺ��d��I�}���h�2�Z�+�)C����A��H�TS������ 4Hd]�<����q�D�S�_�E���P�K%y��C�ɊV�f�yh����@�$D�B�I�L�&��"�΅PE�E  �C�	�!�l��G�1N��y�1$�0B�I�Qff�F�6}V�JW�E1tRLB�ɤ[�4`BC��oq�Qz�=68B�I�3$������Z1��2�Y%��C�	�-��j�/ӑO^�����$i�C�	(8���A�U�x�FaW�(j�C�	6G5�d�`��k�5j0*��^KZC�I+f��D��:�;��	'k
,M��U�p�˅ϝ�[)��q����ȆȓTt�`�^9M�D�c�˒�+Zԕ�ȓ1��t��H�Wy�rb	+&�ZІȓh�"3�g�6Ɋ�[� �mʸ��� �a@�!�=;gd�!u�Ɓ��P<ʠI m �X�l0�T	I�L��ć�S�? `10�,е�5K��R�wb�i3"O�hʓƄ�Q�Ly ��H�>s^@�0"On\��+׌k�-Y%ą9`p�p7"O ��A�Z=Jh�M�9�P'"O~�#���%}C�l�ūH�-*��U*O�E!��J+δ=�V#Υ=ӺLI	�'(�(�&�
X�Tx��J�,G��!Q�'b:�ʃ�2��	QFQ+熜��'X�0�@Ӡ1[�i再���h�'Qڐb�K��R�� ɵ�6��"
�'�pv�E's��p�hD�^(ڱc	�'��h[E*Y&[l`���+��Tzp�"	�'��j�e}��(����T�8�',�x�fX��aث �0 ��/�y�@����Ġ�����ؕG�
�y�ٌ%��beϼt�R��y�� Z>R]�"�	3��S���y�Jɀc���C3e
�x�PwΞ�y�"N����
ABhц#�*�yb� �v��$�g�$V�2�����y�h"BV�t�Є�V9Y�r��8�y��K�+�|K6jԙV���1�^��y�`תi��=Y��_-!=Z�`᫈��yE
�.=�h�����t��A\��y��ȿ��e+�Z4���+����y�)�[�F�Z��X�$PB�" �5�y�O�[i<-W�15�=jRM��y"�G!<Z^hp���1:��� ���yR��H2�9�JP�9��EbPF ��y�I�h�)�A��3.��Z�nΦ�y�mE~���v��=����^<�y2�PHU����J�;�4�����y�N��Ba�"F�� 8��	A�y�ؙ/'�0ҷ��[�`���ض�y�i�Hrv��3a�J��裕F��y�a%_�����b�.I��������yR�B���� ��j��1�B�yb�\�X1��c$��L��� ���y�ފ+�6�{��NM������y�*��3�E�E���ӂ)ȓ�yR��wljԳ�a�@a���B��#�yBf�a�b} `Q\v�a"ٜ�y���6u޴�C�,ϓw�Z��a����ybl�/G.�
��$�\`�1��yb�.`�`R�F% `!-�e�<	ġ¡h���)�}{� ö"OZD(&Q>c��@�Ąd�d\�"O�-3�F�L&�yb`պ�|{"Ov�@��d=.�E/�:%�8-�"OV5�ԩ���L"�#���b6"O�h@Edх-r�Ū"mE8��1�&"O�l�Q�хF�8��N���
e!�dR���U�����~)(R _�/!�.J{�����Y0jұ��,�Y�!�Z,Z6$홦kE?�f�0�.��~�!�C(B3f� '�ǶB�j�.�!�D�v %��dܫ5-�Ba,^!��E�k��#K�:hq�c�FM�!���BRUs3��P���u/݉�!�d/Q2"���;�]3��E�!�Da�$q��V60�깒�@$f�!�d�>hX�q����0�2=K�.אl�!�d��Kx �Z���N\T�#ݴ
�!�J� ��r�'ZOHp%	0K^�!�� �A�Ǥ�1ex|�t�J�n���W"Oz9�bO�7�J�&�*>��z�"O�M����l�83��.H�<�r"O4̱(�	S���0��\~V\�g"O�LB��e��+���`�,X%"O��IW�Z�Rq>̀�� �����y��_�f�l�BQM�2u����Pi�.�yb�3���Z��ܴs[^(j��P"�y�jD��q  ��k�LL���@"�y���тA�$Ǹy�0����yR"�rA��F>ܐ��vAG��yb�ݡ?�Hm�RQ&x�2� ��y"Hߩn�uJ�EZJ�D�SI4�y�EY�9�(�p��ڛ?O\��@���yB��!L���s�	��;���`萻�y"o
:U����&/'(�#�Ά�y�G~�y��G��.����g�4�ybk�?�e�$��>3���L!�y��ҜV��A�"�م>��X���W;�y�JV�u�6��C10������y�&H�Y|\j�H��<@�Y�d��y"$_�F ���,]�7�q��`�'1���e�`� }(P��lal���',T*C@��v �h�!��'���ӁVt*�T����:V=�C䉐�\��p*�2\~Q�P�#1�C�	�~`�X����^��&�� B�7=�X�hb搘xo*1��o:C�	i�¡���@W*M��x��B�?)H;F�Q��"�v�ޅ��B�	>� �(���< Ő�OZ(Z�rB�	�¼�Ӊ��H��ҴM�B-PB�	&�"�)'H�:���J3��TB�I(x�j̓Q)� ��mq��L�:��C�II�,)�!��%vGL�aŕ=g��C�ɾ/�֩!%���K(�B�K�/�C�I�V� )��ϣ�m�����B��.������&�8�p���JJ�B�ɫoT�y#j:l���bb.�N�B�I�L,\�s�f�Lo�m��Z�pB�7������+5�cAH,ZLB��4oG�0��'�28�,e9��R�hB��A��Q��ʔ/���ـB�L C�ɻ<�.`�WO�H�1BKl��B�	��$$��HA�}xb*�F�L��B��{H4� D��j����D��m�,B�I�i�*гS&�=Gr�p��ҁq��B�I�z���V�u�6���QT�B��1/�x���O�OB���B"C�	]���)�OR�L�q%�_7Pa�B�I�,kd+�D�y���s͘���B�Ʌn<���;�찔�	
w�C�I�>�0�`�Gђ fȰ����5��C�mM�	�s���W\)�d�	 2��C�%{�ЍAqɵ{�XqckFhI8C��?e�	��Ñ=zbr�ͅ�H��C�<0C�E��k^�1�a����C䉚��E�"(����K�F��B�	B�F,z��Q��	F�F�RĐB�	�O#�(����Vrq��O͚B�I�[~l[a TXv� ��I�C�=	��j��9r���`��]m�C�I�z�����	x�Zq�XW�6C�I�b�������8ena��#Wee,C�)� Ήؖ��;q޽2�I�G�2u��"Ov��'GG8?_v��Ҋ53T�ҡ"O���E��1W��ʂG\&~�s�"O ��eG�&���I���#��w"OX��4�٤L�`����,l�"On�)U�]2>���b�S Z%^�8a"Ope��˗00��o۽:�՛1"O�K�EB�j���[%�P!@�p"O[��ȸ%y�%"Dm�C�����"O���s=v�8�+%�vq��"O���S��Ac�P1;�d͸�"O|�i�&"��uS��F�i�b�A�"O�Y{�N�	p��� �' ���1C"O������ �pģwD�^�6�A�"OTI`���d�>% ��B�Z�~�!"O:!"��Q����ԥc�$��"O>p��-��D�@�RwH4"�8|�w"O�D�"Ր�<���Ǔ�xE  ��"O^��e��N�`�[�F��LEXE��"O�� *Y=������"$�:�"O�-kA�˦������"
%����"O�p��+��#���D��V*L�"O�4QcC #,�1P�aF s�Ա�"O�$p�B��F���:FT���t"O4 B����2�C�8���"O���o�q:T���3W�:�"O|��-o�٦�A��`"O`a;�c��C��1TM[�q�KF"OP@�Ԉ��T�~��l�}^@�Ib"O�T�EBK�,6D�kFi�.PJ11"O���6�R��U�nМ���(��k�<�A�7)���o��w���0a�\�<��Huc�q(���4��d&��Y�<���ˤ��v�W1��1��SX�<1��*N"�Za)F+4Xb})EJU�<�#��	"���-H�3V~�hVH�M�<ᡃ�����V�Z�D�H��P�<Q�M�9�:MJ�͗	�:�,�H�<�G��Tlr|8'J�k�R��	i�<��JO�A	qM��<�8رKKl�<��b�Ů���J�<�z=����e�<���J�wt�9�3mһ��l�a�<�� J&�x�(�.
�k���8�iVw�<yE�U�b�r�ƀ�?��l@�Dr�<�զ���a��i��S*�)5�n�<�؜6��HwLV=PO���b�R�<���� d��U�I�rHށ�	g�<Y�&ֱs�J�H��O��yT��a�<aq��,f]x��&�"�mÆ\�<I�!�0���0���l|F+V�Y�<i���:İ�5Á+<�`	�ϔU�<sOO�+��mi��+Z�����J�<����L��l��K��L����[�<�@�QF;%Ѿ~��p�!�X�<�uN�6\4F���M�REz���T�<1A)E$K��={�!ǈ&.�ȓ3��S�<y��fD�4�7.�lR|�&XU�<���$i M��4�j�LQ�<�� Ň}m6D��/�n�����t�<Ѡ�Q=)�0����M�dl1��n�<a#B�
2 �C�Q�&�L��V�`�<�\�Q_����#�P��A�1o�C�<)@�O 0ЉD��m�<}Q�	�B�<���H�P_�@�r���4���c��|�<� ��'E@�j4-J�b4y��"O������	Z�jձC�97!jm	&"O� 3��Si��X�J�.84`�"O&��7ƈ,IP�[�*S�}�5"OıS f�nĪ@��f*T�"O(1�v��m��l�E�
z�{�|�'��2CȐ>�P�.N*"~�	�'er����� ��Kt�خt*p���'��A2e��cP�`$䖍p'}X�'�F$K�AF��Ұz��]A���J>9������O�f�qd	X���r�P�h�� �':�SB'�>_f��ҩA*\�>1��'�2��nP�\��щ� �\j�E�
�'�b1��ʙ�X5 3��LI����'BY����9�8�I�J�=�H�q�'%�A�$@`4|��I�
$�ȓ,.0(��L� ���( 60���'�ў�|Jr)�.HN3�c[9逸kt�[D�<)� �0.�l���q��T�]>FB䉕HWΩ�!�����C2O��Y�B�	�c�ڹꕨFn�:պ���n`B�ə�= �酥U�� � �BB(B��46ҠUȗ�<h
����gP�:7*C䉂w�A�D+�!J�a��0BNVC�	�v�PB�(V�yS��$��(��8��C�N�*�c�-�Ky�,��0D�ܪࠋ�INNy��l�؉SR��O\�O��=��F�vBT������hj����C"Ord�樃M�"�"NES�%�1"Oެ�+��w��}H�L*6��ٓ"O>���D
e��p�Ս�'q\u�"O�a��P�n�4��O 'i� A "O���C����i҄(>�Z}�"ORhj�@K:r?`��ed���B��gP�,%��D{�O:��P`$]�|��+S)ܢ*#�9@�R�'f��5��?c�:�M�~_��	�'l������?���KF�\y5��1	�'y8D��lχ�ҙR�ƞp?��'��t�­�56r�;ThH}�,h�r�)��써Y��HP���*�������y�۬68�vΓw�����.�yR!�c��y�rK͍lѦ1#��Y����?��bdsE�I�zw���snM�r�i��07z��������� �D�P̠�ȓ3rIy,˚#�6�6�0B�$u�ȓc,^ X7���L���3�F��Ҁ��o��E�`�>X�(���I�/(�d�?a���~b��2<dx�#����W�4�$C�<��aظ8��8B��8v&E�1��}�<a�m��e�!��@_>M�Ȉjw�Q�<!��Nn���Y%+�8,\�↢�I�<I4��r��{���/8:���Ҭ�D�<����"I&$]A�� �� �B�<9��[>J $��F��8�1*�z�<A���JSN$zH��q��1yĆ�̔'oɧ��֜SQe��hA������(C4���,+D�H�o̜{`�	u-��2uD�h�-D�cBbɶl�e�Ǡ�+ud,(Jb/?D�0�6��)u����c,%+���*D�@���A#.��q���6� ��o<D��á��.P�|��_��IK��.D��2�II�{�H�RŊ2!�@��ū-���O�������&�<��`	�U57,y�ȓ�����`�t~�kT灱��l��S�? 6T8t��r!~"#Ӡ����%"O�c�y�rd��
�/�j�sf"O������94�лB�նIy�ҁ"O�e�#B�2B��H�"�5s���Y "O��*�l� '���C��+y��8� �'��W�Ї�	�`�,	!�eՐ/J�Z��3t�B�I,|�@��;0�Q��1`�B��,���TW=qs���w`0_�B䉛c����`DB�n�����N&=�B�ɢ3����1[��9%BL�w[�P��[>YP�n͔DY򦋆;%^L@�W#=D���&�ǋTX*\c��_�l.|ؕ�-��4�SܧY��u�e@��t���c�f�M�ȓ}�:᱀F�b� J����v ���#D�	 ��N�����Z�����0����D萊� �@��?��d��LP`�����]R��8s��?�ƍG��
�* A�(ŵd��u�7���JB��"z���s	��$���Vi���'�S�OY���5��>q2a�w�(�n@V"OT�6iN�z�4 ;�nۼ5�Z��"O��9��L�-"�rE��E�8�	�"O��h��|�x����&I�HɸF"O<�`0`?g�Y#BB�I�����"O�c�7|�D�"@	�^	r"O����kH#e������s���Q"OX���M����CA/ ��s�"O\�%��	���"�MK	[DQ��"O�h�O��ES�U	�/9�B�6"O�D(6��2?9����q�.(�b�	ɟ�G�Ԯ��no\�en�cb���ʃ��y�@[Kd&�d��H>шD��yr�b�l�TϋW��H�nСjaDC��4��Ɇh�>.�|a����>;]�B�
yA� S���7�� �C䉳y�L����)h�D���G���C�I�;��$��=R��Ɂ*�t㟸E{J?=���DT|ű0�)-!� SV�*D����H�F��2�֟A���'(D��q�	�IS�]��o���]�fn;��=�S�'Z9�Q�^&x���it�F�`h�E��(|�q��Ȫ��0��P�RF����R��H�ƨP2%J��Ā��"HDt��om��is�#G���h�N.?�����W�^((3k�/#��V!��?��ȓ���Е!�#2�5��cª���8�|�k�/A*l��ˁ�;{�Դ&��E{��t��;#�ry�� P#�\%����䓤0>ه�P�hЩ)2���b��qІGU�<Y�C��0�e��1� S� �N�<)U,�=V~��$.w�n�č�U�<���M,""��*.�i��R�<�d͠%���rL��Ku\�1�LEP�<�g˕�f�p5cӪT��0�����L�<��#�&6&��G(_�Y^.�9��J�<�\<2r��w�5FtDQC�F�G�<Ia�הZ������IO�$�@)�_�<���F�z�D�b��S= g@�p�@U�<���r@�pv� �BZ�<�D��j�`� �E�`���/A�<��C� *1��J�P!4�����C�<����?s���Ff�2��H@ȟ`F{���_ 2b�;U��3�ȍ*S�-	4B䉐|������pT��𔦕�,B�)� L<��b��%*�B�L�%0�z���"O�DJ�,U?��Y�eēu!�X�"O�l��G3Y�B'�S��*E�E"O�:�џ�n�cP%�
�0�2�"O��))=^7@�ga����
1�I]�4�p
�E{�d{$�-)Gv#�(:D�{N�5�Ԟ;X=�Sg8D�LJ��[#w�zmpf�E8>� �k6D�d�+�$%QD�����:��5�g5D�ĉ�c�.2Fe�0�5vZ����1D�`�b�7.t���o]�nӴĒU .D��`#Θ�D h���M)b���-D��v�O�<�Hb�' )'h>�k9D�� ��8c �0��o�:,�v@���#D�$x%�-i^,�fX�,D<�l<D�Pa��NE`�vb�H^{ 9D���D!d B�QFJ�;d6=3d�7D�hP4D��	��t�r�. ȡ�I7D�з��wLB�1�i��8�@5D�T@$�[�x�5u�O� ��� C2D��2"a�a��$����R3�1D�t�6�ݴq'|��u�J�}��@��34�
c-�.$� Eȣ�Q1�t}y��N矴�	џ��II��0�o�
g�Fs�� F��}
#�1D����i��/�����/@�{Ē]50D�Z�m,Z2��V��8@G�Y��.D�x�p.�&v���P�&X��5�#A-D�T8��Lu��,����"@d���,D���)q2��C��#*�P-�U=D��iÞu��H��/�10`nXg�<D��;v�O�1��L� �8*���[f�:D��ʾI�*%�B��=�n���9�	S���Ӗt<c4MI�GY�,����G�$B䉻o\T�bޟL��pf��C�B䉐F4 1 #�Kϐd���(��C��C��=cc���f:��;�ݏS�C䉢U>���@*�D�4�m�vq���<9��?Q���O6����K~�Xa@�|ư!�C"On,*��F�;O(�����L�� ��"O6͋�΍.���(2�j�^�(�"O�0!U�B,n��b��
=La@�"ON5xqaX�D��])��Q�sEp�Rc"O@\�b�\}v83�ɘU�b<�"O
$��C©/�<I�#KR
ݠw�'22�'�ɧ��tDHCl�)����eX�t��n�K�<�q�X:9'�@���Ŗ��� K�C�<F��'�$�P"F�
!8(T��A�<�r�ò8:���$��kHF9J�@�@�<� �f��͸����*�� �c}�<9RE�>SB��1I�+5�A�v�<1S"� I�Z���
�#<�q��eHy��'��OQ>���)H`m���D-#r�`��f6D� *�V�0󰭊s�X�+�F����5ړ�0|
T@Z�@�h�w'�1�����\�'�ɧ��JA���"̐���\�L�ɚ��/D�����B?d�L���+3��� U�1D�D�BF_�~~��9b�1��D��<D��Z��J�pg
�it�����9D�0�O]����X�6��,��&7D��H��J����C��G�<�&�5D��k@�D�R���l�L(�����O��6�Of�)�V1�nI�ƀ�W����"O\}��v]d����>9��Bp"OF #BC /���7��h�TP�"O� p�D��_�z$S�����2"O���WGD�Bb�)h3���(HJ�"O�e�3	B�N��SE�S��J���"O�ȣG!�jE�LX�lʡI�h�"�'Z!�� QD�0wm��fD��K@�J�!�$��p�64��ݼ9���Y�Ȗ)1�!�d�p\	
�@�r����α�!�$��Xn�#V�Y�$���K�����!�D4�P�A��H�t0�ɉ"�!򄀠���YbK�c޶���z�!��R�gb�I�흥?ԶL��D�; !�D�>�qIbg��f�n2�d�O!���24ZL*�OS ?2C@c�W�!�d�w�F] ����=�x�#uo�:r�!���>-tx�㇣M���A:��	A�!�ԓwWPY�"�8�r�Qr�	!�dU�m��� ��99��굉N�W!�DB0s�!y�o&y�ĳ�D�"!�^�8j�v� w_�Ӂ�
n�!�	�6#6� s��+?���f(�b!�d�@����R��(E�<�SUn� ���$2x�<xc�D\8|
P�y��.��C��	&ﾉj���W�8�I #K�<�vB�ɹq0��4腆�$��a�L�XY$B��(H������B	kyHc�j�'z(C䉦,dlՉńް�M�f�0Lv�C�I)f���� 9#�aa�;<��C�I�9�����=o��P�G �Q�BB�	�*�\���J]�)��艤.K�8�B䉐z�:����-!���7c݄rj�C��8AG��q1��0`��1�Ì$~J�C�ɷ��U��,�3t�YK�M��(C�&{j�`3��H�N
z�{��B�ԼC�	�V��ѳ������CG�5'��C�	I��pFa֤A�r��$��|/�C�I�~� �&��o���မ�-^�C��;;uic6a��|@��4�ҙ��C��1�ܕ@��ťKN*��#��	&zB䉦0�!��BY,IR�3T�a�B�99gb�����'~T��D��<�C�	2��d@Ч�?3�����K�#�bB�<\(|(�g\�H�Vmb��ݳ 6C䉽-�lq��A�*y� �a`P�,c�B䉹	���P��P6Y&�0�>>��B�I&��#�O�9 x ����h�B��6�1��L�*�`�[q�ʴBSlB�	"m���V�26VH1���2C�	�"��� 5�M-Tl sիD�C�I
0�N�y�]���5��͏�S��B�ɇE�j��ǧgrf����8��C�I#ڨe0d@�:Pm$�%bX�9s�C�I*w�.t�L���.*h�C�	��,Ӂ�^�=�䕒e�'|��C�I�O$]�[3�"�J'P�z�C�	�
�Cg�D��!��9��B�I�]�t��g��0("u;7%M�,Vx�=�ç\�����h�!�$�bE$���k&D�pI��ߺ.B�Y�fX�R����/D�+�g�h��	�g"U���q�q-.D��J��V��f�pG�d���SW�*D���q�0$߬�`�M6m�8�81�'D�ؓ��=$�����G�?�R�:4�)D���t�ì@� �z�EͰ����`�%D�@2��71�D��^&@���j�n.D�� lH EC��W(0,�a�R5v��Ux�"O^Ԋ�N~:ptj��Įr�$8�"O�P��@�|����PI�E���$"O�	hŊ���cu��2��u*"Ot�I�ܑXd��-�#�v���"O��C�[u�rA+Ƃ0Y"����'���S�B�q�j��i�I�pğ�!��D����$�U�p��CZ�Q�!��<G�N	(�O?Hֽ�$��6�!�X7S�0�[Dn�"?ղ	���b9!�D�;m(x�-Q�r�l���%�!�����1$�a�Ĭ
���jo!�$�4ZA�V�������aZ2qh�}��'R@�����3g$W�b��'��c!���v[�� �$�-H`�s&�wh!�Ę%���C�Eʤz/��B@�sA!��*-���a�!���@f,ԐY9!�d���� ���.x]�����^(!��9\T��UM��FC|�	%��=d$!�é��y����_��E�q��6{ў��?��y�Kl���Ύ,H�V���cܿ�?I	�'=�uC��|�L7�9kZ�3�'>�a��V��� wŀ�e/V���'�F��
Wf��apGئdRXqC5D��a����=hP���L�zP�+$�4D�̛7��"|��-(���&�6�*�h3D����W�Xف����@k��=4��� B�&���0��(B#x����v�<�wIY�.���0����[�:��'#�u�<I��n�%BdBэBԂ+�*
w�<q�,�!Gh���͕W�a�aK�o�<��j^�)L��ӖnҶG��b���`�<@� EJ$��O6+@u��L_v�<qt��m�B\ �d
0J
��s��s�<A��Ԥ��H�!��gzt����Dx�lEx�ӧvj� 5��IP̃D�I��y�)L�h��f�@ Dm�������y�G@
��0Sw�S=Q�DtqV�y2,ٓe�t��`ҚP�`���ǩ�yӒ&���C�azeZ<z�e��y"dU�r��Z"&?�ȡqFeқ�yb�¾l�ȱ���ǺY��]��䓡0>a���\��y*��$&��bw�<�pDÐb��jV Ԛb?�@S�/�v�<��@M10�T���B,~-{`kSL�<)�وK�iQ2+� o0�z�o�<�SMݨhz.��ΐ$"A��`UT�<!� ��i2a#[<j��L����v�<I�"��m[�x�d�7h�p���u�<�cC 
�(���ǴM6Z��K�<����C��A��F� d���d%D��2���+֠�Y㨚+c^d�C�#D�8sF4nH�}��I�%yd��w*4D�����/f�4�f�X�7=p�@bf0D��Тφ�ze2�a�
�m�V$D���v.��!]ȝ�,�	y�e� � D�԰��e�y��Eհ�����$?D�L�$���XH�D��oA:e
�?D�����<o��M�㥌�]u숪D#=D�T�D�D�0��I�l[�X�"=D��C�
�Eo��@�-	{���Hd:D���q�
�JR�AO	l���r�-D����F�K�|�0�aĳ��S��5D�<s�'	6F�N�@AҨ��`.D�� ���C���B��|�(H"O�d�PLŌ2�^I8��&9��"O�`��F��^�*��`� �J<2�"O��Y�N�6)pAr�_ Tn\��`"O� �N݀#�`I�R�B�;o�0c&"Oɘv�	�1���U�s�Q�"O��"�FC>R.@)�5nI�!���`"O�3 @�'p�� �MNF�1��"O�a0�4	T�)���ߒChD:t"O$����ɟ_��TI� �a�p�&"O�H�r���+VHB��=+��U�v"O" �� �#@� �J��<E@��AV"O���%Iػ;"a��]�a�"O
aA�ٚ_P�;a� �p�P��"O�E�B�H�@��ح[�P��"O:���
XE��jX�h�����"OFi(�gC!`P��egىf7ڈ��'ڤP�X<�"�&C� ��s�'Z,8���L�!�����hy��'�.�;a%V$Ј*#�L��	 �'�dr4$S k�`�:R��]Ԕ
�'���C�C�hņy�a�ߕQ����'8(��κ"�&�qP$؅M����'��@�W�Cf� +@��4Tm����'�2ICԬ3	����w��Tɨ��'�������Q��Q�a�N���'�$�Jr�-)�,�ǧE�("ցK�'�pI�a�&V���8��W&ъb�' 1�vN�.2�Q���W� ;*�)��� O�uY�ʈ�;�B�)#�AH>Z7"O�E��@D���^�4ʀbȋ�D�!�$�#�:�� 
�P��;VV!�DN8�b�;�K$ �����π-I!�$J�x��%�TC
�v�@�u�۲N9!򄌉a���v��<stЂ��#!�$�x+&t�@�H�ԩ���^�B�)�.A���X`�8�t�̎����'�V1 ��Q�G�ڀ���y�%�/%�ļ0�=Ĭ�����y��ê"������k��x8�dN1�y�ꚉ>U�x��>���R��Ɯ�y�Α�cd�`
VJĞ�@5�	��yB�#q}��8��_����D�1�y�gZ;7.�\�$d� �~�J��K�y@Os��� /������y�c<N��5J�hGXUIq!ɋ�y���K]( ���Y�a�` H�Z	�y2�C��TdYc�ϥT������3�y��8N�nM��EԾ!c�ϐ�yB�  8��&J);���0w���yHU�I4X�x�ݻb���W�Д�y��ZiF-b�&S�b�8��B,�y�L��/5��Kg+ƨT��@h���yr$�"Z�0�P�f��K0`��GG%�y�DL�R0�M�����>�~��&���<A��%^�u�V�_|l����L!�dշ,��XcM��bo2�@�E;z4!�Ę
��8�LM,f��R�B�!�$H�>�������mM.)��� !�䉕
KJ,8%@�sHZ�s��|�!�䔯jD����+��e:�H(y�!�d��K ��J`F�'����TCV�t��{�\N&� @e��K���e��r<!�dցa�Rpk����{��˃R�W�!�� ����U��rX�u��
��A�T"O�eÖB�DP!枧%��� %"O��Z��v�l�`��;�b�p���y�<�FME?{�X"���/��yA@@�<�L��Y溌�Ɵy������{�<i�S��v��dʗ9^�a�Pw�<iCBCKj�bcL�q��qS�Y�'pR�S��0(A��6��x�_�2��C ��	�Ql<O+ސ�эڽw!�d�4��I�����1h��?z !�$Ü��M�<>1CRk�#�^���"O�Ib�E/S.��f��ߺ�0"O,-xr*^�59L|��$��U���ˑ�|��'A��!�_"oap`	 ��"i�I��D*��HD�T"�J�U���6�f ��"OB�9� JPZ �2�� ko�P�#"O�%�f�<c+ -Г��S�bH�"O��)�cGl�b�
ǇV�^�jZ&"O�8j5,^{*��q �X�z�D"O�V�.:��y��-�
}�4yAP"O�,�AU ���ƍ�(^�[""O���r���P�L�,D*�(�"O����G�x�� ��K*�D��"O����O�$��a�ڎ3:��"O���ݦ���Ӿ�p����{x�`�'�xmа"'&�m��.�|����|�'ݼD�	6T��4*�SŜM��'���G��<آG�Um��ϓ�O���X:M��L�_a��q�"O�`kwn�5ː�����"O������&�p����%�e�v*O�qS㊣agR ��J,���y	��ʻ?`na/��M�� s�\"!�R8VָL8Ӭ��X���F�!���D���TVL�@-�&���	k�O��|ʕ.�0x�N0�BC30D�p	�'�(ҧ@PG &|��o�`����'/��9S���D8C��(摠�'�V=�凒>��H#C (u� ���'���4ƈ�dZba3�mߵr�����'��ԫ�m�d�␂�; 4��,O���/�i>!�<A�LE�2��$bwf�Ig�5�'�Mex��FxR��rAMCCdA; "�S ��yB�ˁK?�d+��	�5�>��FӶ�y��l���f ��%�͹fD��yR����8� ���܌ #�ڜ�y���b�PD��Z@��DE��ybΆ(/BX���cIqŇ�?����?����~�`H�>G�~��h[�O*��IS`�<�w$��z�1���.[hM�Fh�<� K�Cb�bt��*,Ԅ!�0.�d�<�VA��| 0T��>>�HY@�@�`�<��0Pz��j���
��	ze�B䉓+]�h£瑯y2 �B�`O�B��$����Ȏ�S�\���d%O��=�����}@$c�3Y���I5a�N_�t��"OL!U��:
�h��I�L6@q�"O:�`��2S���I����)"OLT����,��I !hюs��Hr"O�D���fnXi�GQ�d�ᩓ"O�1��D&3p�"4`]�Q¡"O�-�B�&{��E  �0{����4��ӟ�G�t\�Yl���i��OZ@��a�?����?��<�c{HɉSuq����f�,�"O� vhqt�A�m��Y��!,Φ���"O�8K�̛�{p���g�5�����"O�ZD�V�L��䚷�ΰ1�
l�"O��)DL��\��#��ڸE �X7�'���'H�CVB��|`�Y	V�Ԑ*�����hO2�=A���
�h�@��=�*��P��yrKz�.嘴ʍ G��e2�I�y��үT��#���t���y"��Z:�$@-Ms*ݚ�bE$�y�ɊL ����3w��U�	�y��:�Љ�pO�ڶ"����-�Of%��55���BB�9An��2X��D{��&�`���¡p?n��Lt_!�Ę$j`���3I !a'�@�,V�*A!�$ѯ|r\���
��1�4�`��!�_����c��+7 ��/a&8Q��'P�� �K��bP���˼j9(��'�`�%3/�t<����7c�MZ�'4�9	� ��d`����.6If!Y�'C~Xc�#�j:֝2�
�;/���
�'��hfIV:Z��P����*���
�'4xm�th������¬�j�	�'�Z���.r^���/M���K	�'g<�K���D����)�nHZ��d<�'nh����h+n}!4�R=.��ȓ{�^U�e�Z
/V������?��u��I�<Q����|�� <Y�4X͂k�<a��/#pH���/DIz�hy�if�<qՠ?}iP<j���~�zey��L�<y�B�n	u�c�,e�h�W��F�<YmNeE%)�4�s��D�'�a�i�P�m�A�*C������y�P-�zH�DW���3��Ż��=)����dɠ ��M` l%{X`pvf�l�BO��1l@����3`I�|Rꬱ�"O�{�	�4AU� ��D�n�"��c"O�XS@�±#[|��p������q"OT$iө��|}��)Dǔ�"�#��ID�O.���Ƭ�)���҅®DG��a
�'˼�B��ܠ_!�D�
9��U�ϓ���<q��F<�<�
% �Ȓ���yJS2#N2�Q ��4�pB���y��Rv@M�e�ē���!�d=��'�(��嚼,�AB	�e���a�'̀IąQ~y��IX;_Pʎ�� �&�'���Vm*�c�6`k4OW�<IO�^��1�QH��DX$�R��SH�<!Ơ��c�D�0eĺcoٲ��o�<A�P9��)k�"��Z|L�W�d�<y3��+�.@�C\8#�5	fKM\�<��ǉ���Ai���B��?�NI�ȓ�#�'jX44k��T̈́�F������+���bā�T�0�ȓE��!;��	+j39($A�����G{�'`��5e�<y>0�4k�NL���'�>!��ے��Y4	C"`��'��!cC�۸w�R��-4_X���'0z��c�U�$�Q6
�..����'�5��ˏ6p�L��d�޹19,9�'
Ґ+�L�D�s�!I��R�b�'{ҍ��kS�Ǌh���F�K��k��-�D:���<k��p ��ap ��@�A�<�0�E#�N��MO/{�a+QEI�<i� ���0k�(O&[�@ED�<� 8�;��1�>T g� �`1�R"O�9z�
Cxu�T!��]����%"O� ��&F�%��3�y ��"O����aM~d�
��Z~r�xID�'"�L�S�Ӧ����F�g��L��<�����������t]C��-��ES7"O���k;)�^,�vbY$RlΝ�"O�)�UًO�>}�s,ڶ/Y|U�w"OBD�vi�Hz�m�v��U�\ZD"Of́ugW�CI\�U�N<H ��"Oީ������Nu��A.͔��W�'��D*;pH"�Z/I�����kΰ.�!򤁋p�����C�7T�vH����%�!�DՙK��%��g�N�����ᐝI�!�DQ�+kO�s������ �
��P��@ld �F!�"�(����<R��ȓ�H�*a�� ��)�􂇺/"捅�t�d(�Ϗ/f|�]�-�HE8���	� �''d5x�j�-
�s� �;d�*	�'>�����w/��j�_~�� �'�@���ݗW �DI�L��TH
�'����O�� f���ONP��	�'D�x�P�[e2��!��E�C�4s�'��A���Y�ʕ"�F�w�
�']:H:�Әl�>�[R�@�Cg�k	�'��ea��h԰qS�A�G+Z�#�'��%�S0q$Q!U���F�Ƅ��'L�ar���8r��H
E� 4rP)�
�'j$)�*A {²��Ď�&�]
�'�j-걭��3��t��,��0	�'$�ux5�J	&��hê��*�����')��r�8(f�!)��&6d�P�'�PD��o�S����D��4�#�'?r8�(D+T�F����*;Ax���'g�х@]&��]�4��'Q�t��J[�nt;�˖/UGLh�	�'�zq��;Y~ʤ"��$�k�'���r�*6�X���ΐ/"���'�~��k�oڦ�z�B�}چ�R�'lX`�U��95z�YCf4���'��쓀55�4��+�p����'<<���-3�J��V8? `�':v��n���� ��47��#�'|��9�(H�0 ��T��7���A�'��p	��!,�1�J�_�6k�'�8QZ��`M���@
EzL���'\x��!��%�,bVM	.8o���'F �9"�.B~.�&���0��
�'}��+�kܡc�hQ@խY�+�-��'��dk"¼5� ��� ���(��'���m�<,W��!�J�Yv<|)�'�d��r�>Z "��Lr` �'Ll�q�	� r$nٹ��N�>'
�X�'���y #�)E�~͠�D�*-���	�'p(<��\�	�N0qͲ@���'��1ЃI^=�P��7bm�E�
�'�H�[Ԡ�Cl	��E�+^�`-��'d���UjӖ%9� XS�,Q(�J�'�����D&d��1�C��6N@:��'뎠���/e�0�p��-z�Ё@�'{t{B�8e�qY�I_o��I��'Et<����'I���
@݇l�FP�'ZN�pDA�D�|Ɋ�;o$���'�8�딅P^B���l��̂�x��� �i���=iЈ1�IB�q ��x�"O@<K�,]�JK��H�G�r�c"O$|��+�C
�+�mP,'e`��"O����@D%Ij����m��^$���"Oh=�$Oӟwؠ%�ǌ�
����"Oн�GI�5i�)T-6��P��"O�%f�4`3J�H�vtC�"OfxS��9%N}X����o\q�"O<�2�
?!�Hբ@�0!�,12"OF(aп_��%�ը�#�=�"O!�âN5-4Щbd��.��	��"O�ժ�m�PK�x�'g�e鸽;"OHE�F�4�Q Ĝ�#΄5Y�"O�,� ��'��1�L[�&M�"O8b�hύeK����{� U#�"O|X���< � 1Ă������"O�@�w,M}2q�עןaR����"O@=��l��h9�%���#��5�2"O����!�6��@�WDz52��UJ�<9@�˕(�<��7��E�H�f��G�<)w�-eW��! c79DM�RIJ�<�Gҝ	��L"�ֈD l��mYD�<���-z*ҍ���O
H��ף�h�<qp�L4R�� ����0r�q���b�<7�e��� ������	J_�<�G-�0r� �A�Rتq�J�W�<ɳ�	]��i[D�R�0�y	vl�T�<�v�Z 48��r����O�<Qq�S�+1�H3@��
a<T`　N�<	r�vd��㳨^A��	 �J�<�
�8aԅ9�]�\�\�Ab�<ـŝ�,�49�g���l�B����b�<!�^"��l�	��s��T�<�i�tfѠ4�\�\˔��K�<�˞�H�x�c ���~������K�<A�⌬A�hJ��[�X)�dϒG�<)���{���3C�N�W4�a��E�<���2Hs>��JD���I�s�A�<��D���r���8>���|�<!猌�,��ʗ.�x���x1�z�<q����E�6���s���:��Gx�<���Z)5u��¦�Ɲd��T���u�<�l\�y|�C�,��(�,��2c�t�<��.Q�j@0C���K�b,B�	��5�Q�جvT�(��DY�~�@B�	�%���R3���y��P�i��B��5_N�t�����=���گw&�B�	ow��Z�)��B�L�F�l�C�I�	� ٤D�%��A�eϺv�pC��ZYH��&B���sgc˷I�2C�ɼ\���O��G�v�P��3W��B䉳,^�4�,��(�r��t��B�	�C��w�#�8) N]x�B�I�&��t��:R���P��% nC�I�J�y�(���䚁L��$}B�I!Q!Ф`��0������̶b)HC䉉.}aPa��?�nL�n��@C�	�}ԂdaBJs�<xB݋�B����x�2�I� �h������T�`B�� h�ұ��iB�lxdC��*0~B�ɭM��X
�[,W4ڡKӷ\�xB�	 ����KA��FS!@B�I	�T*�^0}К	���D:i�B�ɒ.����ā/tpT�
�bݲ[��C�)� &q��J�- ���|����"OT�Ⴧ˞Sx�P s
K�h2}�T"O>XHD�)%Pr%�VD
�Kg����"O`8�j�	ꬄk�˜F=؈��"Of����&W'xm@��]?�M�7"O�AX"� � ��F��� �c�"Ot��LD5MƵ*"�ʇs� ��"O.�1,«GQ��#lϨT��Iв"Od]��'�1q�!3��
�IfpR"OX�P�ȟ�Y@�@i���)��0#"O�%"T����qb,{Ԅ��C"Od('F�-26���K��P`J�"O���I�r�������s����v"OJ��@e�#�� qf��kA�L�E"O�CB푪A��#AL�� )zlsF"O���
B1t���`�g���"Oh�mT�]�h<H�f-���k�"O4踤k�=G
ě�%S�e��XB2"OlPj��7_<i �e�;'���9#"O���F�@㨨a�B
�ZP	�'"O��3&��V�u�!b%6�cp"OX�[�Y�N�^tp����VPf"OH9�`�ѯ3޹
U�=��=��"O��)rLJ"k'��	pG!crސ �"O�*2�%��ą�b�| �"O�@�v/�#�ҙx�-ʙs���C�"O`uI�k"��œ�ϗ7B ��"O^�R���i$�L:�L�se"O�}ـcE�Y��q �U�r���"O���ˋ�] ��I�N�;3P��G"O��է�(X�ys�(> �3"O���^�Q2���	.���"O(i[�ː XX���h)%�5�S"O2ԡ$Ӝ]T8��F��&���"O�<҅Ǿc~�Q"�8E³"O�[�d�����AVD�&"O���d%����#������e�<)��I3(�>�óKıdT���NXi�<Ap#��1�������b��=;q^c�<��R�!�$a%���XN�FK`�<i��g�Tݺ�#F�c��!҆(LX�<q'��Bk(9Z[�+Q99�ԆȓV_fԫ��� <�$S2M7d�� ��~���˔�F<U�2P#�1;����ȓJ�mC��4p�\2�Ț	8�R�ȓ��=⣯X�*I~Ź�"�:g����	�@)e� �Ap!"�� `���ȓ2�|��UaMb�V���l[�L����ȓJh�S���9�>U§��}�I��z����j��ܒi��U��f��ȓq%�yGŜ{�uqF��V����o�b��B���F2�Ya"m��#'b���rx�4JX�y�nM	�M	O�F��L�e�e��U,�R�N��q���pbz�Yq�����x�@㒀}��L��Rb`TÎY�0�:�>��2�"O������9�ƱX0�eڪ�m�'Q��[ҮEC	��8KD�?D�����ة+�Dka��1b��8b 8ʓ x����1Vt�@�))���	 �H�o_!��*n�ٗϵZϾE`0��k��MG{���'G9��Ň63�dr��]7/ƹz�'�*�y�'�*��lr��޹����G{.��$��5
�`G��3K2�� �D}a}��/?� p��E�S)V�����fN:��"O&(�P�>�P�k�1'Y\����Du����]���qʌ:6nB� �$��M�C䉽7��(��@	g��]8cKSa��Ø'������dX?�d,>�h���F�#Lؼe�&�� �!�D
Y��Y	" �+%�p�j g5����O�b��F}�,�	��� '��im`��I��0<���DY�(�X������2"%�!��
=Y0��SQCEI<ؙzab5z�铗hO�O���|<��A��tu�F'A�!�de�N��Ɛ�t�$�7g��c�!��M�k���������f�lo��iӲ쫲"+h�()�Dҡ]���"O~���&��*a�P�'>&�8�'�1OƘɁ�]�5)u���[0V��Y�X�@���-<:�d	Gɕ��D��]������#�S�	^x:�y�ᇺGe� �$$V�D!򤍖50H��œ�"R��y�Lr���hO�I�fC�C�ԥ���3^$�2"Ov�a���Z��p�G��|�� �D4lOn�i�N��XxR��� G#7��ɥ"O�Рu�#J�̭��n@�a��"O �А�S1d|i ��:�z;��'����oQQiN�J/���A��]~��d>}��݋���hY�-NDu��'��y�ۙ+x����9%�I9w*�y�&�'�$�q��K~�x���&R��y�N��y	��)�V
}4
�[s���yr�-n?����(C	d%z��X8��']az��F;!C�h��oG0>�x�XU��Px��i�8h���;`,ZР�\�Ql\�"�'*�l�P��%I&�jS�P��8	�'6���a&Z!BUXKs� YEn��'�VR���+y"U�@k*X���~�
W�B�'��d§�K�GȞ1���	�fضD��o���ڂjp���D+�3u�R�:#�RU��	q���ʠI�< ���G�+�Z���*��(O��Ӥg�x����:^1>i��%T�Ok�B�	�j�"���j�&&@$�z0b��`1ZB�	9m\�ygR�"�愂�&�8 �vC�:HF�x�DY6~V��ǧ�k�DC��530iC�$ܐbf1Qq���`B��	yz:�P ��>%J�z&�F&I�C�ɿD�r07�^ܹ���kFhC�	�,o
�Ӡ`�;2�qA���S9�B�	7\�yY�C� ��A�d�&5h���>��B*Z��]��H޵	����FL�'��O�� �O���̓2K 6�j-Ov��A9	�'Q���3� .���:v�P?l�$����D3�'}z�C%"�P"yH���/VRT�ȓC]���u$�2�N�J(�+K��Ɠ!�X��qOL�~��t�]'w����'�ڤk5$	�p�������	<�$�َ��<O�	�Y�HM�J���Yb����"O|e4���]�a-�:��T���i��'D�z2�F7!�,I�TJ��l�����yb͙*8dstF��T��c
��M��'M$�Т'Q���x���fX�'�ў�}���.���`"K���,�f�j�<!w�M�*j��0��i�d9�%��I��HOb�$���QB�x���y��;q3�O������K����(�4m$�C�	�H ,�U��	X.ɉ5IC�d��=	��VI�O�Bɻ�F�KD$�GC�R���"O� �(*�gB�V���;wg�:=j�@��'���w�ĳw�0�w�� [>�1*2'"D���R�j���1�slI�$a;D���c��M��W��$@:��G'<O�#<�����~��xB�^�I��,�"ϖM�<�GH�}���b`� �,La�G�<)��[$F�Fh���m��@���o�<�@BX �2���<kV���o�<p��*;�� t.�w���P�Fi�<9���3$vnR�8QV�
�8x�ȓ2k��a��3��	����@I��ȓq�.�#��*H��l��h^	�D��'�a~��վ��!iE�G�y~�#'��y��ߟT��tBӠ	-<X1��/D �y�E�9O�]��*�,=�q
X��y2��^-	�%�8�� K�޴�yB�XMry��L$0D4�!r#Ͱ�y���b�ff��x��%q(��y"	�Z	��i��Ƚ>mz-�%�ܶ�y�f> iCa�	����D���y���-zX^i�sM�o�@�)�GZ2�y�oҢ;��F
ݻ!�0������d1�OT�Q�ۘ(�ԙa4�@*�e[$"Om!���[���FIV�2��P�8O"�=E�$���V��s猗I�M
�EE�yRh�WzH0��ƜCl��F�����$�O0���;K�=����[(�XV㏩+U!�ݩ��HacS�3,& ^c�!�DԢv�a2���D���9F�D�A��O�����w/��pg�>M�𠱈�3��x�E�,�TLq�ǼR�<`3F�9|���Y��`#��D�^O`���P������.���|1p��ڎ!��Ȗ/P
o�=[��<4������4:��	�⏞�{Ndh�hi���=�����<�d�d ��؀��b����W*�8�y2�'��K�昹�H��m�)?���	˓m%�7m� ��F�ܢ�h�*>�͚�]���'�~���.�X�BE�ɔN|��'`�M�� ɛ�Oq�X+ ��b�`�B.�0(>�b���'�'1��x:#n �)�L���b��9�6`��|�v~J~&����#C�V�h�Y���2��94�L��Ë�x��l)ҡ��dJJ�Q�����x"�К`�`�ρ2JX2�@�/�����(O�0эbJʑvb�	HE��'��(���ɣ�y�)W�W���2���\z�����'��#=%?q"#���fW���&nY�%������;ʓ����		0�R�a���<R�艂e�Ҙx����'�n�{g�đe�x�"��<�6D%�2�S��?Y�"QS R��!P���ݙqa�<��A6�O2�x��f��QC�[`{�@���Od���O�=�O(���`KD�!0�U��J;8G����'Ԗ�J6��6U�胐�Š{��K�'Z�����+m���Y��J,{��y0�'��8R#h04���J�\ʠ��'O���5�O<Q/T��Ǌ�J��aE"O���A	� ���-�Y�$ b�"O��r�Hfs5�����_��90�"Olv�G�m�:�C�N7��)b�"OH��B\�&i�����/6N�	t"O�M�c'F3;t��o�8z��	*�"O�7͓�G\�] 5,��
��hs"O�qdK)a�m�2l;�����"OL�`,�
]F*�k�!ɐ.�t�"O�Re�(uъq�g	��C��y
�  ����8;x�4�_.�6Y"OB��Ńh�,��cD�G�|1j�"OV��Ё�7YlR���!A>z�"��G"O�=�ե[*�Z��b�X*��P��"O���#c�*ʜ��B�[;y�Q"O���#��* {L!Λ9fɸ�"O�����8W����B1^c��ӳ"O��2��B��'%ӷ+y$���"O6<*&�̀*�p ��'���e"O@��QN��Q�*a���.PM���"O�Db#�bG��۱A�)���"O����Ƒ��d\y���
I���""OJ`�4��y�ĉ`ә$�V��"O�	��D^�ajb3�i�)]����"O�@�У��V%���i�Z���"OΌ�B�_�xT����	?,���#"O����1�n�!2�Ռv'�k�"O a�.�<rw\��A���5"O�Z�	|jxh+$MX��P�"O�}�kH�U�b��&fN�m�&��S"O´+��8�Y��G��M�����"OB�ʂE ֌<��Cqp@@�"OFx2D�X?��cDG/O�����"O䰉���Mb���B�o�f-Ơ�?� ,��F�*K�-���'����Q�q��1�ڈJ��$+�'�*`���ag�=��$д6B���'��Հ�&K�,㌹8w q�HX{�'�F|)u��=w�Z�,��i���2	�'��m���(��swa��5��|��'YV�Ul�!Ԍ��E�<i\(!�'Iv�)��[)�d���+N \����'�����̙b��	ׯbhC�'n �BF�߳.�>�!hE��JI��'Xb�HE�In��9ȅhP O����'��m��c�0[�\i�.Ç��x�'�TH��0�fP��Ȅ�6G�TQ�'��@i�&�*2��3�ı.#��P�'�h�R�&�']?�r��Ɍ$�He��'j��ぜ��
YA`�&%����'��A�L�-F+�y�RaD&�D��	�'�ި*��[9@44��Ԃ�%�u
�'��H5���*i�C�	�,M��'5:Љ׬F=3���D)�7<E�'�L�X�$��=��aB
D� H�'�dܙ�C�}�`mY � ��e"
�'<|:���nb�y����'�4����H*Z�piŊZ�"7b�p�'n��Z��ܸO�<5*��_�/cbų�'�Fl����H���p#�S�"����'|��wm��Hd8u!���!P-A�'�$�C�Ϳ0X�����
�'J�@�덜uc��E��V}��t�x1t�Ϭh�`�S��
k��$�ȓ�LQ�V"�e�.1���Rrߦ	�ȓW�NɸR� `��`ȟVC\Y�ȓu�$���?Q��8���I�P���|Xf�ʐ�ߨ]�D���.S�
ͤЅȓRߠ	aT�K�.rL)���:	/���ȓk�����'O�1Lp�#쁶^�b�ȓqF��e�M&*�T�ӡȋ�@Y��=Q��s�gX#s�TX����?� 	��	�
����O>��5�.3�U§�ίG�ɒ�"O8��ġ�K�8���oH�^=�\Q�d.m��
�'C��,+dM� ���9�
N�d�ԑ��S�? P�afK��2bX���G��P�:}j�g��e�qO8����Y����S�-��	ˇl	���T�!D��P�o�j�(�@��ĩU��� �g���V2�Oj��G�@�59T�
�m�L{��'N ��b�[D~RE;OGbU�A��/:V�Y����yIU6 �&8��cǫ%��I�VƸ'�@��,�c>͈��]ZF�1r�j�j'�-���,D������N�<d�fI�Y~J��e�Ij�O� E��O�l�WeW5-5��9��S�`�p"O�Pq��F$�ږ*��z��d��"OЬ!�
� K����2�ޝ�P�"O��tB�5g�pa��T��q�"O�4M&Ch�AI�B��'TX�K'O�2�֚8���y�o�r��Xe��9,_lC�I�vע���a���	􉊈DZF�?�6��nFxb?a�%�J�6R���m��s1&�R�l0D��)��ω	e�h��'��(x!�<���!�6➢|2�oF7Y�P�rP�ʏL2d���Z�<� ��c#0��&�̰����CV��1������'.��1&�`x؈x�ɚ���p�	��)��a��K)5Nn!(��t�4$��B�-��B�D���NW
5#޵+�n�\{ȣ?1�O�^,�b?�[@C�'��<h5��]^�	De;D�5��m�`'B�1b
J��ba2?�&�D��������c��좀!U
h��ܰ�"O}��L�JLʂ`�"@g��U"O�8�c/C�-��#�)F d?T���xRj �|��=�~��%�/w>;�d��|,�� ��a�<��J1q�:�(�JS�7P�����n�N/OH�Pq�J�M-��2��D�v��D���ط
h=3���#.�y�k6	b5ϓ.�\qG�{���J�/5s���4��C� ���٨%� ���b4�	���5*�P�j� �'YY�'�^�2u���0vc�1y�D����-W�t��5���˓)����)�KV
\��^� �朠#a{biK�z��ɛ9�.�;e�Lb�����L����R'�hP6�K��'�J�٠LR$0��В	رH�j��G1|�ͱ�O41'��b9vy�E�ދf)�艀(Tuz�
��W'_��X�B��XY�Ǯa;t}�-O2 J%�]�Bp�塞%*�X$)���5��5��+�V8��f�B�K�i�	*���"��#Z��V�Ax�&� �*�p�I1�na��'J�,�UfD�j���<�UNG]�	؁F�";?�p�@Qo�:<�|��4^���8��
90��
���H� ���|ݡ35cö��E)@�`qBՉ�=��$�#l[`P�NY��0=f��*�Z��4fW�(ZRL�ơ�|��	UIjb��b�&m~z�&^&(����A�EH���hEfG6G���p�^+m�^��"O�(���O����B��>��<�F�g�๡���,/sZ��� \j�8H6�^�M����'�z��;J�������4z�����/�&�����,��$��"\�'��ss�A$�^�d��jC~�4i(�AF��I�[衃�]o1O��n	��xH�u�]�1����I7�n��E�TIh�+�e���A����Ǿm]���s��Y�8"7��$�y��B����0=��n�p�4�I@�C&��eXgF���� M*� ����po��˅�H������|��띐!�@�i�(Rp�d�����I�'c��dE�fT���JZM���(3D 	Q�$8�P�%�ua��3D����y7���.ͪ�n�x�g'��0?���A�J	FP��ç+� �b&$^���C+�.X��̐*dA&��$�~�l�h&�v� q�ީ=��`��Ԍ�4�BN�%#��+�ןXi{�dG��TZP��|�"���"O|���N��Cei�g�(���OB�P��+H|f!�$!�=�#:�E�[�>$ `�?Uon)�b%G��P���צ]�DbΔ��:�Z��<}�v��4L'�D!�3b���o�k����'�8�9�
S���{������Z�4�LqH>���ڇ6�\�y��;:"�L��3.�tN�UH���3�,�O^A0Ј�z��z�U��(��?O΍��o�(�'��ܛ'��i�ؤO��2�-�P8LqsBK� ��u	�"O~��!���7��p��	����r�����A ] �E�=)�Ȯ���+I���uE�&�S�^h�����µ^�JU2���n�*�ST.	s�H�8U��f!�� R��U�\�-��lrF�����Ɋv�����@f�8Iֳ'�� b��CTdB�	����i�1����A��:J�x�	�I?�I�?E�$��r�6�9�܆�t���D �yB̐�CɢhQ7��`"ޙH�Fƃ�y�
Z�g�z��3�ÏX',<[Aiӈ�y"�۷+��J�$��`~P���@��yM7F�q2�U�6,Q�Ѝ��y�ɇ  �p�%K�.*�x�@�N��y��G�/��4�#��$���ku@
��y�aؒNR(-�P��/�p�)�y�'T�/Dad�މ ����*�y�I�%�Vi07�G&'�f��s���y"�Y L<�|����!\h-h�'���y"�c(���N�W�� Ȁ��y��O8WC�-H6�Ċ>��L�"g��ye�A,�%��&EѸ�K�k���yҎ@�J(�ђ B)76��L��y¨��P&L9 I�%~������0�yri�%\�Y��O�eC��3��A��y2�C�X"HU 7!j��le%S5�~Rꂹ;dT�=E��c	�6��UI����]�88j�W�y+F��Y���m���mÇ���	1r��3AK;<O��bf�� ���"�,��9��%���'��1��	
.e��P��sÚ-Z��
�F!�3Hܓ��x�)�/ac1O݇2�>�Adf��hOxi�Af@	G�T�C�����:e	��e�ԝP��Q��C�yR#Ohn�{�D�|�$���d���?��F�quX��)�(N2!��4�x"�8D-zdRƀЁs<��a��x2���F*X��,B�S���Æ?
��  ��LϛV��Wsƀ0���UX����hJ�����ΌY<�ö?�)��#�"91d�3�[z<����׍�� qo�?N��aZ�i";xC�I�'�E��O�ls<Ô��m�H�>���LR 1c��2Q-I�C����a[�N�6-���u��� �������VZ|ț�"ON�[7V�Q��l�'S�Ui~h��N�u�da)��-6m"%�F${��Ox8y
Uf��y���o���K��]�h@ �j��r�'ͥj����1�¸vOZ�2큃@H������$�o+8D�)H0c�+}�#��6�_t��
��0�0QP�h] J� ER�vt�H�4�Y��#Dל8��!�ӣU7�
�Q�7i00�PA��96DY���'/�qc��w�PY�t�,n�i!(O�Mr�!S�b����'F�����Q81j�f+��/
*�@V�%,XA�s̓T؞Ա�EK#	p�I�A����%���C�"�����|/F	H�� JR$��b+���"OX2��@"k����$FxOv(����lC�(�	�^ ���E��G�O/: ���3Kߎ�k�7D��ူ-Ϲj�)����O2m{$�}�����6�Q�v�ɰ@���Fc��&�.l��d��q��?n5�=*,��o6"�{�B]H4�� ! �L�9�t�4��*f=}ԁp��!M�j=i�I�c�|Ϛ+{�� y�a�JUSHD�����c����T�3�Nt�!�ګz��4Yv(
DI(3�Ć��th�j��i�&J��u����2�z�az� �p���BOZF?�R�!-Ϡ�����wY��qD+�����=H-ry+�H,��2i�a�	#4�pڙw���3�gC�o�����k�h�H�y�ICn�v�QH~�O���b`�LLaOغY���6�O6a	���4����5��l��L�0��FlQ��Ą�V��1���H,�$�PT���\��:�(�iX�vt����c�*��S*�����Q6f���0 (ӗ7M�\B��/:wY�� �6��D��<��43�X##�Z�J�,ë9��\�(�0u҆9br��A�,��ìL�?��{WM�#'�B�*l*;���:v��x�D��L� �� �azb��#i�� �B?�1ˉ
$�A�i͎���:���+�����@�����0�߮}���Q�KI���C�z�Vܩ6:��h���
L� �#px����"xl��g������� R�Q�P��ë��}u�5X��M�L�TA���<����'o^�P�G�+C"��5�	?'�\��0`�M
���W�
�z�K"��&.*��+V��v	��t��Hy��O\�&eЦ'`�[����J?� b­�`VyRR�_�4�|2KS�d� ������+�<���DD�=�6-iV��/�l��B�JN��#[�ty� z!�aׇ&#��)'M���n���`K\�����M�h��(OnX �Y���y��:�t�8$�  �/��%�#�i�3�	�&Ŧ��B`��B��;��L&+��C�I�'��� �X2���u�L;7̌�Yk�}Ar.�$!�b���K�p
X���JB d�E�F�õB��x���+#��<�0(��\:�5-�� 1Go�<q��ܡ�B�{��1����&DQ�<鄤�T���ڷ"�/L��h���J�<�v�D<�
����ܕq2!4,K�<��߸d�lAGʌ�{>�$Q#�A�<1��ve�h��E̠dT��@�<��AX�+F���ӣu��4�y�<����ꘘA��� ���psc�<9w`L<n���r�'A"x����Qv�<��(U,{P� rb�8�@!�h�{�<	�"Z��X�P���}�Hy�#s�<a'�ާJ�D*�E���(��bl�<!s���r����b�WW�Ʃz��o�<	��ZQJ�D��$��u�N�<�0�A�0����3�Ŗ>��8�Sw�<�^=S\q�H�9�B��m�<����xrx��f��2CtXK��P�<i�����Sa�|���"��L�<����%�p�)ڲz@�i�r��H�<١
I�@�3|aҡ-BI�<�WM�;��DHN��t��Q�M�<����� ;�S����H�)��OI�<�㌖
V*T��M�:t�A�!n�M�<��+6\#l�H1ǝ9C�����A P�<y"�^�}�`a�4%���fL
Q�<A��]�(���(E0ܔ��RC�Q�<�%G6A!a$_n�ۗmz�<��ʖ9�C>2#>$�Fm^^�<q7�ѾD����	�?McR8c׉L^�<���Sn��	�%�
H8}bi�}�<!�Gњ7���K���35	P-*dN�g�<	FU�8;"II��ҩT1���[a�<�1�
@�p:��P*M*�a��e�<�ׯN'^$\ɧ�_$e	`�ど�g�<���S�T�F�#���1+$Pc%�K�<	dH�7$ج"��B�?��pwh�@�<i2��za��[�#�^
zUX��e�<�AX�����42ăש�x�<�!B��R�T��LTn8&/Et�<1�̍����%m�-"}蜚��Av�<�'��
'�����.�k�Z�<y���sf"�2`�>P��q/PZ�<�⟫U�i+����]�k�V�<�a�ϣs"9V7$��hW��L�<9�/��6��'_�S5Yro�K�<ym�f�81ɡlǯv�~�`�\F�<�"V6v��t.�ox���h�[�<R���SyA)�d�.vlz5I�LV�<9'�߿Q�vX�P�+a0FcM�<A̟m�L a@%m�j�H5��\�<EA޵*�>1b��M�wU�)`&��]�<G�ФF/H�1�j��f/X�ת�T�<y���cŬ4�cC�i0�8Xf�AL�<!�+��E�l�!�'D�7��C���g�<Ʉ��E�8�&�F`���e�a�<�F"ǆ3N�u@ �K�z%���PI�<�ՕR�@��-�2���5BK�<)�%OL�M���I2������i�<	k�gz��sd�bg(��q@I�<�#ϑ,֠�2��"B�8R��/D�RW+�(4>��� �|1mr�l)D��ڵ!̴v��!��m�+����ZHC�)� &+�ߒk�ڣ�´��R"O�r�m��Q� l�X@A"O���f�@�It8���~C @K#"O��QA�@M�z�I�=x#xe�"O��WA�y}8�5g� O͌!��"O��dޏzv� 8�D�C��r�"O�@�3(d�(����z=ڐ�v"OE �Ԡ��	���36&� "O�}���'v|��e���T��"O� E�,J�+�o��+� Ib�"Oxh� @�j��M�B'6/� ѲP"OxY4_�>���W� <����@"O��07!K�窡C���ڢ�b0"O�5�� ~ɘ����_�$5s�"OZ-G`Σ.���2"v��"O:hC �-	��eHU��)I��"O^��xӴ4� '[Qۆ��1�y�ʑ��>ܩ�d�� �
pc���y���pHm1�T((.����P��y��\�n�L4""GM��Ɇ��y��C �TD��h�9����:�yR���g� D�@�$��4m���y�8 �*PL�.x��1��
�y�^�1�h��
R1{`�r����y�7�Hd�pj�?k�D�ȳ���y�Kر!�fȒalJ06Q���؄�y�.�6n�����Lĩ$pN�
d)٢�y�Ո.��-	� �P3���������Q�e��8wK�qy8 �ȓ@���rM)%UM�gQdT�ȓw|�9�KZ�S�Z��qǓ�f 	�'��xP�#ߜO��Я�++�	�'Y ���1_l��i�+���1	�'4���$��<f$�5E�%��#�'P2x{TۮlD��H�h+��'�varA�V�T�L�ިm0��r�z���@��y�h�t���:)�a�b� �V����o�<	�	:d��K�dUV��s�~�`�s�M�Z����K
ͮ��O^pa��.�U!�ݏC]"q8e�߬ ���W�P�<a*K�/ߤ� �*��:mD����'���Â�Z	A��	&KK���"/�6h!�ON�N�>m&\%��gA"�����@5!�$Y$ ��r����Ti���:g8�Ȱ�9*�N�{���UyZw&������1O��Y%Ѯv՞���.Ȕ``v�'�&|�B�c ��mZ�c���9R+�
|�r2� kZH�IXn,L0 cVkazb��2m���"�&�� @�����'�^-�3#9b��'q����~�����}�i�
<4�y#5�GH�<�w�u�=�E��3y��-{E-�yt�1��2^��52B�m�1��@��OE��15����N��-��k�'OM!���@��w�X����u)��)��(�A�Ž|�����A]yZw�H����١�1O�Q��e�J�DS�4�z}0'�'`JTӑKp��Unڈ&�e�6�5Il�{�E�f����@]�q㞲.Caz�L�?��Pp�;Aj�!1
��OB�2��ٍ}��'I���u��3�H(t�c�R4*�N�PW��s�2D�PI�K$��Q�c̸m
�2j4���QbI.�D���?I���;fqn�	Te���IG��'BjA��v�t@�s��RQ�IҪVSح��OS�x�#���x�2�����=�4�ȓcD&�Ґ�B�G��$��!�C�ćȓ*P2d(��G~\�YJ�ڮr2T��$ �q�b��q Dp�e��8��x���*JuX6l]�D �Ņ�3�ĭ��B	�o��8e���fF��ȓZ� ��@�-rhܒ�O@7:vK0D�(�!%D�����ƈ�^7֥��&D�� X�.\�N�J� a�ېi���h�"O-Cgћ
j��%��:�|<#a"O����ɚ�ؔ�g/�43�j�7"Oڴ�㫀�a��s�A)�޸Au"OFjp��Y�p�gΝ5!��QB"Ot���o@�/�����n[�1R��*O�|���qْ`��.u���'�: �6[��u�weH�ao���'
�P��ϖ��
}���F\��=��'� <k�oFD5�Y��{z
�Z�'��uH& <�����Y�� �'~� �,6xPXl҇��0�ؼ�	�'0���@��YתQQ`l��}\���'L�q;@�`?Ri����7be�B�	�ج	RmZ�tݺ5����7j
B�	�z�%����R����9.Y�C�	b,. �C:9�,!KV�\0L3�B�I�a�X (2�4M� k�)t�B�I�A�x	�`H!y،`��ڏnh�B�#ʸY5%C�A��0jb��(d�B�I C�zx+�
�%32bP;���Wu�B䉟�b�C����۔쑃���Z�DB�	=%Y�$8rbJ�#Lt�A��T�,B�	-]����, s�.�Ȕ̜�y�B�	�d�\�s� �,J\=��CΚ^q����
�mA��퓢G2EUL��d�B)Y�B�I;���R�ˬBX��ue�|�Y����GjJ���<��Yi[,�x!�0E����'��Dx���wF*��a��Ǧ�T���ܶ#�l�ʕ�87;!�d�(3f�樊gΌ�@0��0�ў��F�̓\L�!��i�h���T%G[�lAѤX.i�!�dۀk�MqG�]8�d4(t��/v}��r���c솃C���r���!�$��k����$h~Iiq���6�!��i��
���#�|ҡ��2\��L���]�B��7�ܮ@0L�:&K���<�&��I�h��r�	h��KU�'5r�[T�Т'�Y �
*Y��4C�J+$�H���8F.��`@�$3P��ēb��b�"��Kg�E�	�2H|�'�&�q�%8�(�k2�L���hRb�u�K?��¨�L�*|1A�BC#^YD�6D����'T.U�p��
�y|{�lљ/@�z�c�ze�gG5"���ty�7���!��I�NL�c���	b��Q��<����MT�jAI_�R
��)'��X��jM����8ݴ^*��N�\�q�S�'�V|��,:J�]�gՒ4��M�'Ԓ�L�u�7C�O:�XP�vJ�e�vi�@׹r���`)�P�	�V�0?Y�OX�z�l�c�X�~{��I�,�|yB��g��ő���<�->^=�4a&�^�>d��6)lܻ�%�M�`)���D�a���ĝ,d�:�`.OV\r��i��Hթ�cP+�(���:�f�W��1��� 5S��O���G���Q��D�L�H�T`�".a`�4K�WzqOP����*?�*"}�eaD��"L0mE���8�e�h��ɹ�2�2�	�_��	�F�_�*D8��&��H�1;jI��%�3z"�p걊����g�ND�'����&�{X�8�;+�l�r@���iS*9j`��Q�P#^^T���4�䤆�	�V�DQ��Ag'��A�i�4U�L(H��`�
�QV���\X{����'
�W	�4���O,��zt2�,={SMT	,rQɇ�+��!���'�����	��z����r�R]����r_r��s_7h�M��)M�ap7�V91�UÆ���v�ZU��l��&M@1�y�dܕq�
�	bS��B�,��'��%�/ K�UE��$�s���2vC�A
��qa��Qf���D*�-`70� �^��@��-K���b�� �O$Y�C�M+4�1��(�>���ϓ�g1�5�L�t.$��I�&�Xtê�(9ZRa�SC�h�xp���9r�8��ݩKFܛ�%��>�B�ч�s���䁾\�0��&G�6 # �sM��U �0fh�`"4-��5�j�A�_�K��I&C�.h�`�)qO�iݔ)�`h�W';���g@B 0az��K�iq��cP� ?IBI�&t�HԹ��7.<�%֤"��qj���:^�y{�B"_bU
"�[f��m���\T��9�,@��G��^!����E�](���F�uxu� ��ZL �\\)`� �e��td�E8cE;+�6��E�W�U�Y�'[�M�����f����5%ʡ�wa�0��e�e���P��DkB`\�x�y�ұ�ӹ�:Z�FY1��`�'�O�uCrË�p��`��TєPA�c7%3��Q�
���|
� �`�!AٔuR��>".A��O&�Yq��E��cABR�Ys��+� ��G�	���';Z� �`�E�@f�0#d�|���퉌d����S�0�S%K�#D�(���ޠ @ʜ;W�ʓ
fL@� ��gܓN� X�cJ�:?����&ѿHǶq��N�(L'*�30��su��2�n};V�s�Z0��h���^&e�1,��M����I�z;P�@���#H�d̑���
��cP8
q!�D�8~j�ϽOn�rB�N�-!��B*	Ȉq'�ҝR��r�"h!�!��a��B���:!��] v���@Ĉ�R2�iV�a+!���t�\�9�fF|*�ehӗ[!�$�<v��3��&Z��q���!�����g�;$\�x8�Ȣd�!��b<̉q&'��X0��A�<;c!�$Ɨ}ZNУ���#b��j�OF;-�!���\��Ad�u�nE9�D���!�$^�7ȍ��
W�<�*��w"�ku!�dцW�*pQ��D �>�ڀ"�4kZ!�D�N^�5���q�a��S"[!��e��y�GS(;Rj�Jà�C�!���?��7J~�Р�!�x�!�d �?v�C�Q j>�B��yk!򤑬9DT飢+S*Y��1�A�+A2!��E%4lp���Ɩ�Sg�II1� /!�)���[��M�~TԔʐ'��$�!�$�q�B���I�M�R@��l�18{!�D�T�l$��� �H�	���5Y!�D�W�"PF̅�`�Դ;�ö]!���l!'��]wX����(ji!��[ �H��L%��M��H�/�!��C�E�6� �/աa���#���"("��%�L!b��]�%raz��_�3+���㘋84�Q@#�y�H)�D=��EL/3�ވ��-�1�y"����$<9��й��]xb莽�y��:-K�p�Ƭ�/���"�f|��'W��ҡg�򴑡��fY
�"O���iB$ 3�q���4>���'"O�R��5{��Ăт��z,`lZ �'�^Y��.�)�[����e���@��1F�4�(ɲ�J�=_'�'�*��O����r��h@�Iæ�S����(ݜ�E��OT!��:�0|��GS�sꊄ�D,S�:$I�J��y{�I��N	�ѫc�n�s눀���KtV�����Y]d	+��Y�)���HwE{��T�"�ˬa�4� ��~�����x�w�ƅP1F��A3��ˇ{nX U�Q�`�94��<�`m��+G0�!�!-����B�\�b$��2��rj��<���j���Y��M*h��O�/=��u�ˌ�?9���(����Sk8�T�ӳe�^}[ #ƌj���rk�:z��9S�1`Ȩf��g����g)�?�	u�'B
.��2 ���l��OL=I�p�)�|0�G��c��%���?�'���ⓊM�1X�4:֋��"|y��>��0�%#�?q(O?�gCD�I+4|���Y���8p1�>z7F���b�w�S�?�;[�:���̕9;`"�� ^Պ]�ȓ��!���J�1�S&�4b9n`��Zn�e�tB��z� ��2^O�8�ȓG��\�fB  -H��o!zVх�
�$�2�BE�D#�8)�O��}�d���3^ ����B�9p�jS�
-�L�ȓ����E�C5^d�kw@
*-�ȓ_��Պ����듢Z�SF�݄ȓ]A�a���.DϺ�SGkٖ6��Єȓy�r�xB% ���+��=�u�ȓ1
��ZX���XU�όL�tن�P8�A�;�|�]�� !��6D����QN$D�C�V]_d| �.7D�H�gO��}m!&���X�X�!D�� ڄk N�?н�6$�"),��c�"O�l�T��?]��z�e�T
���"O؍�t�� ~��Mh��Т`zЫ"O<=��#T #042D_�֑[g"O�=��c�ۤq1�iuB�iQ"O�y�'c".�p���&]]8��"O�|�-�,@��Jt��;J\��x"O؀CGk���S�Ŏ9Kԍ�b"O��rd"]T��PD�!.J���"O�щ1eK�5E��I`�� �4IB"O4���
�o�ސ��^�ʘ�"OБ!f��H 0���-0�d)�"OD�#q�в1�낏T�J#�X��"O�ݲ�ߵ&+¸��`B}ڲ"OPeЫ�	;~h��#�X�ɣ"O^4e��1�L0!aÖ<<�;@"OJ�q⍒)؁�Q#�_9D�!"O��X4
Ԏ4p����E�b����"O��+���t.�5���]�R���"O�`'E��&���9�́F�]�4"O��Ї��<�)����2��C"O�Y�!I�f�Ф ���Q�����"O����̃0�����#6K�I�"O�9�T��<7Z$pB �^8�Z"O�t�w��@��� s�ʚs��}ې"OH�2�b[$`�>0ڶhښM��`��"OF����M�o� q��(Hz�$� �"O���.�`̪S�\�Z.���"O�q B��nE����̍��րb�"O������
M4݉�	�?P����"O�� �=I�� s���+(o�D0E"O�	�O*|$b��ݕA����5g^~�<y%&�
O$�KǪ����ↀ_�<Y�!�	[JE���K|::�
��[�<��.?c7h�:U�B:�~��ǚ`�<��;�����/�
Q
����O�X�<Q�GE�U��ݚ#� #R�q��TU�<a%��R+�쁰���( �ٰsh�v�<ye*�rtx��`��:�AV
�M�<��	�"[��J +�/��	A��G�<�db�+$�lH#�0��%����{�<��)#�R��R�4���R��_�<)q!��s �-�Q@�2
���UL�Q�<)�- �P�z2�B>L��b'�O�<��&vPL���܌,% I���N�<AW+;n�P�:u��\Y1aɟq�<E�)�ni`����`X����I�<�pL�@^а�u�g��9�tƎC�<)��Y�pd��`dKҼDQ�f�Tw�<)�nĪ	މ*���(`.Y���i�<��E�(}��y��c>{r.��m�n�<928@<�
B �?��x��Yf�<���ܙD���f(F��lpR���_�<�a.�37q:0+#���㧅�Z�<a�*Ӕ5?��sN��]�<�c	 `#fd�,%���h�U�<IC~�����(*����Q�<9qoW6f����%i�F)HǄ�G�<y��ݣOА� ,У2�nU@��A�<!��U�:�KV@K��GLK�U��C�IL�!�?t����-�4G�C�%t3P��v��./�v�:��޾'�C�	Z"d�b3%̤*\��C�%�4B�I[�b�c�*=D�8C���<�FC�)� 
`S� ,�"�ڧܚ)xɺF"O�$@2�1�rTS��H�b�J%��"O�r�fÃp��<��!;���"OE��#�
5��8Ƈ�n���I�"O|�$��f�^�RS\=ˆ���"O4e�3-f��$r����3"O��`��G�y@��W'�I(8��"O�M�#�ņ+E0�9f&�u�I�"O œ憐R�5#DL���ˆ"OL��&��0+?Hi�̙�e�-�"O���c��o���u�K9���J�"O��S�B�( ����	݇��墓"O�	@��t��@��R��"OT)�@�P�*cB���-��bb�2�"O�A���]+�&4�F�#>�6a`�"OT����A�[�XX�̎_�P�U"Ot]I�D��
2aZ� ��9Lm��"O��`v"]�2����)pKjA� "OrC��w�@�� �\�,!p"O4`YaN�u�ݚdiM�;4���"O4�Hr!��mA��W&0t�s�"O��S���� ��AB�N�9"Oz�J��c~2���X�}QA"O�qa�NF�WRQ(�֍��"O��e�$*��і+ ('B�tW"O:I���Խy����
�
62���"OjYyv��Kh��3�i[�Q��%"O�h��c�4���:$��$3��а�"Ox��@��V�:�cힶNh�l+Q"O�ԛR�٭c���@��
T�X(�"O�dX�L�>o�n�+0N��2�"e"O�ܙ�D���Lz�	���L
�"O��3��T����@A���x4"O��!���V~��k�*�j�~t��"O�x�3D��y��9�u@P�oy��"O��@Ts�<JV@Ǥ(a��"Oȝ�1Ϧ]�ޘhSƹn��I+B"O�ڂ$� u���u.�1�X���"O@��@`J#���9���0����"O4)BI�_�:4K��Y�H��� "OBr�&X2|	&S��  Z�P5"O�mIF��XZ�e)�����"O���G�ůG�&�kĊ��?��"Oԥs�.����9��~���"O�)���Y	)�h�$�˗�|�a"O8�p���,WK���Շ�.����"O^iHf�U�I�n�Q�IB����"O�dy�m�9Pf���i�r���{�"O�``K͗1����f���Ps�"O4 "��3��(Xo@�3��`�q"O�܁q���k�"9"e,2�Dt��"O�-+��(f�A0'C_�@�j3"O�=��)݌/o� y!��'qm�q��"Oz� UC�#�b=�"ß�:@�"O�����$H%d�����x���"Ob�
�A�}��`�Oծ6c�|��"O����)N�m*UB&�؉E7(Hh�"O�x2vh՘h�P��b�>qyr"O�� �ͭ	�TK��1#�P%�C"Oj y�N�! �u�S�H
fD�0t"O�Ԃ�$RN�P&�ع(w&�R"O��h�(/i�,4�g픝_2��"Of�,5F��� /��I�'���y�+�3s��)� �$����q���y
� �Y!�`� 4�t�REӨ3���"O$`Z��E�)��a:@�� F(�[�"Ox��g�-MH�3��H�}���"O@�vo�!]j6�3S���X�+�"ON��4�_�{������ |� ���"O��)*�`{.�r���nକҒ"O�	�J��/�-��H�A�D]a�"O��׃U b��AQ%['{��p�"O�dsGQ-zH���ƅ�+W��H"O�|�u��4i�� �^���j"O���`����;Q圲"( ��"O�a��@�l�D�dԖV9���"O�|@�L��_���X7U~1�9�"O�Ց�	O�4MS�薚^/�� �"Ox�ЅO�z) I#H�*  �"Ov�*씯X�t5�4��Y� P�"O� ����tS$,�%i�.�����"ONa��螮Xj��򠨄�?>�A"Oҹ�p邽��-��&&ո��Q"Oj�S�<)Xd�j_�;�:`u"O�� 2k�'<"� ���X��"OF���߃�$�:a��)(�L�0"Otq���`�6<i�lА"��Še"O(�S&eɯ$`�d�G�@�"O�Ԣ'@ɯV
}ٲ!^q&04r�"O�%��@�?3���i��޲fV�r�"O�1"�j�9 Mx�
�6bx�a"O�I���њ#�	�AC'&Dҹ"�"O6 3�+ҝ+��S$��7=����"O��1Qń�"�=�Ǆ_	*J�E;$"O�0a�L�/Lx�I��ރvB�)�"O�}��	��&`��đ�1X<0Q"O� �wB
%P􀐩X�M�(0�"O0S'�~b����3A6!�"O��u���&�Jd�B���H#�"O��BGGT�%�^5�kS�s��DzE"O��±�� B������&JŨ�@"O<`*ugلw�j�H�� ��"O"�@f*[/J���ĕ�:O�)k!"O�"$a�4��Q�����?v�Z�"O� �0��#4���FI:Z�t` "O�����K�4t�`	qh�T��!�"O�	v-J;.�xT'�2L����`"Oʉ�G�� >Մ �����V��"O�ۂ)1���E�=u��5��"O���+�=vzn�Rd�At�aS"O�b
��rg�4�$$�zS��[w"OX�XC�W�Πr2CW�>Jq�"O,<�V!H&��Z�l�w��"Oҳ	lO�A��߲� �1"ODًC�		Od\�ږiA?ؐ��"O*4�A&H�j�Щ�����uYT"O^�����7����,o�l���"O~h���.#���uCW�:7R\9�"O<� kƭ_��lY��7�x�"Oei��sfl<�Շ�*v8L�`g"O�D����!iev5�"�Ɣ7���"O�<�#A�/���#(	! C"O�L�u��,];CКW$uA"O��9'�B�I�6�����`ׄ2"O�-J0��,����H����"O�Ar   ��   �  T  �  �  �)  45  �@  �K  GW  c  �n  5z  �  ��  S�   �  b�  ��  ��  =�  ��  ��  L�  ��  9�  ��  �  b�  ��  �  V�  � a
 T � � w) �/ �6 �@ �G ?N �T �Z [  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8��H��I*Hă�%�it"L�B��AH<��	öZr��r��H+}J����Q�<ᕆ��8a�%HI�Vݚ�;#`�L�<�ǅG�a��P�����4S�h�O�<a���!=�Z;!)��䤒Wo�L�<I«��>Bp�Ā�L��%��T�<�􅌏i����䇺>؈�i6n�L�<1&0E@�9�7Q숨�����xR�[�wb��j\�g�T����)�yB��,�t��܀R�Lex��8YW!�dߟ}�6��-���H�HU�"OJu`�7��⦌�#7�d�c"OJ)� ��/e�:PYq�f�x0��	JX�x�(G�r�q�Cԧ?�Fp@$5D����*�:(�th
��e`)� Nh<�Bg�Np
Ղ�ݼ�;U��h���?!6�R?D��('��d�S�	�Z�<a5�K7�i U��i��U��n�k���OY�)�Ő`m��#@�YifD�b�'����i�J��8	��ʴL��ط�O�"~ΓT J!��57LTH��Q�ܜ��ȓK�p�0�A�/���qGH
ad̅�CS�`�(6`���C7��=�)���>E(�#Զ(�ͣ)�=(v�݅ȓc�����#O�`r��s@·IB ��e�����C�R5"|�d�G�Wlt��.r��Sk_�I�Q"�(��Ic� �ȓ]�~���D4&�p�q�ϧ� ���GS�-M�F���Ck�'$�r؆�)Rp���"Y�R�n����l v���;&eX�%ڪ}
}@�gd���.�ի�o�.Ŏb�Isb��/>��cu�7��DB� �#'O�x��9�{���;jh,j��å �vԅ�S�? �@�V!��\&����dN��Q�"O@Dځ�B�yn.��6�P<;�~���"O��"��Зw7j��IY�U�Xik��'��Ć�5Y&�#���,~V=*X�7e!�č �<�{���+j)�t*#\Q�P��cZT[ׇ 2f���*Sn��5�|B�I.] �X�2�V-���n�:s�fB�	�-���	/�n�����ٲD|�C�00 .�x�/��U����8l��'Zu V��/�n�zů��dH�rǓI9`��)��?1،,���,P�M�¿��B�	�@���c֍U�!9�E���C-]��pG{J?Q��OE�7���A�'�Z�X�[�*O�0���`��UM�-F�J�"O"��##
MD�yc�xT���"O��D�Z2��	84k?cc"��"OFI6l_!j<��rV�ÞN>VH;r"O-��D�%T@�
�(�:E� �Y"O�d�fh�#W.�)�V���
5��(�y�)�Y���і��*�8��K�l��ȓS��,P�(�?�����L��$Szp:%�im�\F~�cĈg��� ֋�1T�P�*炓���=y�|r��,G�yd�J#D�E�ƪ�5�yV/C�r�[ ��$=�����
�$�y�iC�d����#�14��`R�d��y�\� "�@͌0L����� �y��Bgz8�C��!m`����y�@��V؆��+l�H)��L�y�Nٖ?���S`-W �;��Z��y��"Er�rR-�InL�sQJ��y�ɽ~D>�)�JOS/&D`1I��y��= L��9�C
H�ح"�"�y2IɀgJ\RRXC���B#KW(�y����D� �aG�e��{�EW��yR@�B1UG@�V0���QN���yR��7P˺��p�I5NM��P�'�yR��%9���(�<F��xb@���y�%[b�!)A"�09R<u��m �y"�D�v/`���X *�䭩K���Py��4S�4��F�A6�b�'W�<9Ǘ y�1y�A_���sF��G�<Q�aG1`y��J�M�i��%�*_N�<�1�_�.�D9��+U	�~�gk�Q�<�w#m=Ԍ����1	:���#FW�<Q�E���Q�p������Tl�Q�<Q�j)����P�)/�~��!�K�<A��[a2�	��ȼZ��� ɗl�<�L�<q��U��W����`��<i��1 ��Sd�M,�޹xDG�{�<�� :'�`A��N�4D<�Q��}�<���ʠ5�z��ҥ�)?�0�Ey�<��$K�3��̘'4��4��N�q�<Q3�"f�x$(�-J(=�0��'�Yl�<!�]�$d �K�̖�~uCgBCe�<	�i�;���V ��.�֍j���g�<a�ʲm�JLAڿN_��9���n�<)f����s�K�q�gmQj�<��Ʉ�@��`B��E�ޕyC-�^�<I�$�yU>��֋�/#��A���d�<y�Ɇ�ER��R �ح;�6����]�<��6�<�Y��2h�}b�p�<�� I�a��W�b�|��Dm�<���$}L�%aGoU~x4�B�L�j�<�Cǯ>����@Iz�yr��f�<� ��B�!���"fe�="1��r�"O�][��ۚ_���˰�W�f$�Tc"O�Y��8N~�`�V�TD�`qD"O`t���/��=�ҫZ�z6J�1"O@�z@�!R�4�)�'�3��0���'T2�'e��'��'��'�r�'Z���Հ/�����.Ȕ~I�A��'>�'���'���'���'C��'0ԩx�IY�C���e�G?E��u�'�'�2�'�B�'���'e��'�R�'���P�FI��9�#���H�%�'vB�'#��'%2�'?��'�R�'Ä�z�-/�r5p��O�b-��d�'nR�'Q��'!��':��''��'��M)��X�	&��KĥA�9;� ���'$��'G��'{b�'0��'1b�'��a��=��3�h�)��ʵ�'�R�'x��'-"�'�"�'�'������kP����)X�+w
u0V�'��'���'O��'��' ��'¦\[�*D(?TȒ��%��G�'���'���'B�'��'�2�'�����4O�4���eɍ`Z�)� �'�B�'G��'5��'o��'P��'ƶ���֊{� �q�eA�M�ny���'��'cB�'?��'�����7M�O �+��r�/B��^�(�!�O����O�D�OL�D�O^���OJ�d�O��r�i�&���O@�jtı�&,�O��O����O��$�O���覉�	��8+���h�jlbƣ�,e.e`"����O��S�g~B'�O�Cx�\8v�Ŭv�A,Յ8�� �'i66m(�i>�I̟�k�-~j`C��	�{�,�oA�D���""f�m�G~�1�V}��r�	0Y}��JF��%�n��1���c�1Ol��<��i5M�.�!�f^�c�2��0�E�,y�anڭ%>�b���R���yGA�%Os"�æ%�`����R	�T2�'O��>�|"q,���M��'�plx���||�6�&�i�'��d���<`2�i>��y��p�� r:�G�k���ILyr�|@`�D$����>ђe�p֥Y�TEm�3Aɂ�\�O��O��	p}��"���#&X�q2��� �T5����O�	T%_)j`1����j`����14+��ٔ�
5�z	!���G:������O?�ɜU�H�k`�X�4c��̣n��扰�M�CC~r�tӆ��ӼU�H�o�/�u���A\x�۟��	�|q�KA����'��)P�?���&�S�ȼl�h�B^n�'z�)�3�I�X��$��E�N���(�¸Q�|�bћFAŅ��	���ғ ��y. U�4�D{aQ����I��M�3�i؞O1����O:���/��T��P8t��5ܵ���<1C���Iv��������$
.~9�Q��(�$]
B�q���l�a|)g��-��n�O���0
C8b2���UV�p(�z�=O*�oZP����	��M�d�i�Z7m�5FB�{⎓z��`h4���=pY�f�p�!�.ke���I~���}t")1v���-��"fđlRXP͓��?��M1*�����ެ ��PD�L&����O*0m�Cb0�'mP�F�|B���l<Z�L�� c��X��'U��������6���bغc�L3H�&�Qv.T5"*6�Pm?�M>�(Ol�ĳ�N;D��7��0%�<2�2�_ʛ���5���8�O��4�E���2#н���V1 �$1�ON��'���'ɧ�i�Jʌ���&�?������N�Qا�E&`6�Sy�O 0�����0�x���K[^��|��l��9�|���?����?��Ş��
�鲖��1aҠ���#F�:�X$��(T�8�' 7-'�� ��D�O��R�ȦpY$��M8W� s�E�O��Ä��7m??�)VC�f��4���W�`mP��u��X$LA��K��y�V���	�`�	џ�����O[RA��A1���k�k�_TV���|�"��3&�Ot���O�����ɦ�] ]�()t
ǍE��m�Df�I�����M���|J~Ѥ�$�MS�'�е��;B|(X���Qe�lI��'\�	*D�ğ@QF�|"V���	ɟ@��C�9E���p�ƒzX��QݟT��ǟ�	AyB�xӦ�Jqi�O
���O�L��@4uS&E 7h�z���'(�I�������͘ش6܉'��1�s�%� ��Eg[0}��yQ�O�AȆ�B
R���"-=�i
�?�"M�Of��b
p5&��v��~F��y��O���O2�$�OJ�}��'�$tڣ%\!Ma��ܤvz�՘�� ��b")���'��7M)�i�M�u�ܭY��+7���<Ysӂy�\�ݴE���i[d}i�i��	6=�iC��O��H��)H@�M8M���BR��xy��'B�'��'�Iʷ :���Qቕs��<� I�9V��	��M�B��?I���?�H~Z��7@��@"�&q�c�FZ+g"`Z�T����4Fl"�x��$��*�~$!tb<Se�I+7/թK��K��GNo�I�TWXQ��'I8�$�T�'^x)$+��t~b�y�I�S��-Q��'���'�����_��3ٴ@ؐ�B��[���h���I:��&O�pΓX�����b}rFf��u�IǦ��s�6kv�!#<@\B��PHۜ�m�H~	A�B8��ӟ/�O#� �|K�h��
��d�7a���B8O���<N������
����#E7��˓�?��i	,I	̟��mU�wk00�ӏؙk~�A��&�kO>	���M�'j����ߴ����;q��;Ǣ�tB�X����i*�Aq�H���?9'd%�ľ<Q��?���?ɤ��Z?������`�0��l �?Q����d�)IE��D�	򟨔Oj�A'��7m|�E����<L��m��O���'���'ɧ��[! >�r��l�n��FO	W��-7R7M��<1!�j� ���B?�M��xɉu��9,�t<;��Ӈr�B��G�O0���O.���O1�˓&3��#@(|b��B�a�4>���	 )�Ɣ�g�'2�x�"��X�O��$�'�\,$!F�G�]
�K �6%����O��"�L�Ӻ{'�����T��2���<,�)&�F<Μ����a���'X��'�b�'wR�'����]�!_�S������F�d�E�ڴUQl�K��?!����<IS��y7�^=Wr���G�ċ%%���)`�"�'�ɧ�O5��RR�i��d�{=a�
��e�ى1=Oz�`���~��|�X�,�	矠;�.ο[�"A�@6n�"$��J����Iԟ�IGym�j)X�e�<���r�	��M;\���sɎ�ͮy1��)�>	��?�K>���GP(��*:�"y�sd�N~b�TМb�i#<�� �)�'�B��O���q��,Qy��H���:?"�'["�'!���ğ��P ]�[��$��d'3X�v �ʟ��ߴ./(2+OLul]�ӼS�B=~s����D �0�$�W�\{?���MC�i&����i��Ibc���O��P5���6h굁jar��S�IBy��'m2�'0��'w	Sy!t̸�J�fU���"N�d��	��M�0��<A��?�M~�}�&U�˷ub���"����P�]�,����'�b>	A��yG�X��B\(X�1�6[��� �4��D��(�b�'��'��	5'�!Hp-'}�zLՐR^��'W��'x�O3剢�M�0���<y�&Q�xB���I<.Ǡ4W�^�<��i=�O�	�'��'D���/�p(�$n�p��(�
9z9TrQ�i��I*��%3����ߍ;@��
���\�K��4�	b�(�	����I̟|��My��4f E��Q�d+1hR�'���y��'���|�dy1b��Ȩ�4����3񩝵	�Ǡ���8�[I>���?�'	aH��4��d�4�݂'�A�<zt�ǫ��ظ9�'��-�~|�_��֟ �����B�p��r
�)u�D���Xޟ���oy��~�19g��Ov���O�ʧA(��R���E.F�0 S�����'D�5��6��O$O��=-�H���P �| ��K�Av$A�ӍȞ(��� � �Uy�Of���	 �'#^�u��)�
�`�F�"�����'��'`R�Or剄�M�	�:�����D�l.H�dfm�ƨ�(O��l`�i.����M�J�)9 �p�%�>aB�P�JO��&Ag�nK�Nj�|�	�P��T���,�TÄ�<�S�l����\�^��3�dأg
���Hy��'�R�'>��'�rY>��"*�	Sg1hCL|{���eH�M���#�?��?K~��1���w-�%���RTےD2wM��l7�AB���O"�D)��O����O�>��t�iP��9Ef�H)�N�?�b�{�1fR�Ď�*�\�A��-�,�OX˓�?q�1��H
RB�>��IA�T%�ג�?9���?q����Jڟ��4��On���O�$x�fI&dv�r�ٛ<wh�4�O��O`��'���'��'7T�����g���Hd-3�Er�'��[�D��ܹ#`�&����\ő��H�l�$W3/����O�zU.��f·;[8���O��d�Ol��0�'�?I�eE�.��i��fK�gCf@9����?y�'�,�k.O�Im[�ӼG�8l���I�80ՄT�����<���?!��kdT���4���L5	U����'���Ҥ�@8W�����g���y5`,�į<�'�?���?����?�wL�ˏ<BW|tj����P��@����O��D�Op���䅔_��)2��	?H�S⨛�1�Vy�'�r�'�ɧ�O��mKW�зg��h�G�X}���R)R�U��O2�z���%�?�vm"�D�<a�
ĭ:�%bIYY�r�F��9�?Q��?q���?�'����例97��Щ'k�)I06Y��A�i��9`�Vݟ���4��'�$듪?���?ϝ\�� ;ю�(h����'_��`�4��d�����c�Oo�O��ɚ�E0���$�<z��"��y��'WB�'6��'��)�-��ұaو*׎�[ �� mz�D�O���^���B�Mny��e��O�qZ���dF�y'C�?Vk�DY�=�D�O~�4�D�ZT�b�T�Ӻ+�(Q9�幠GY1v	��1{?���'��'�������ΟH�I9�B(pt��Qp�M"�he���şx�'57�Eq $�D�O4��|rE��)y� P�i�#{ߎ�"�+�t~�N�>!��?iH>�O�.]��"�{*4!���ÚGЀt���R>I���Ǳi����|"tN���$�d:���
2���J ���:�͂F០���I��b>��'�6MB"!~p�pUy5(J�G�$1��3a�OT�$��5�?�tX��ɖ�I�T)�p�b��f��,�l�Iğ\kV��y�u�/�<p��i�<� ��У)k@%C�O۔=�V���0O�˓�?����?����?���)ʬg�zmpiڒKJ��Ȃk��3d��oZ�ur"]�Iԟ��T�s�<q����ᜄE���YN��[�`H�f�}���w�ҍ'�b>m��J����H�1�,Ñ+'�]Hg�@��̓B� �3"�O��YN>�+O���O�q�)�	ek�[�)Y&Q_d9RŁ�OB���O��d�<���i�b��T�'��'e��`X����r�-G�P�d����$�O}�"xӀm���V�6�胤ح[�@i睯J�<M�'����ƤËI��EZ`���&CɟxZ��'���8D���<�A�
�6?�|�D�'?��'�b�'��>�ϧ/��d�����i��X�C'��[����;�M�3"W��d�Ԧ��?�;'��L�"�_+�t �7�L�j�����M� �iĂ6-�0�6ma���I� ���Ӵ�Ov&��άT���ǆB�SZ�r6��c�	gy��'���'���'��$�,N��\�d%ۯy�P1c���(e�ə�M#p^+���O�����Ă�jRz�p���J��@9��(V1$��'P�7��Ԧ� M<ͧ��' �"�d S�O�ZP���)$�1c$(?].U�.O�x��̕��?�T�3��<y�lο?^��GX7\�����?q���?Q���?�'��d�ަe��$c�d)��>f��SE��bv�5Ab���4��'���?��?��Fƣt�@��.X�5x:�U�=! DX��4�y�'��`���M�9O����j�A�\�c����CX��#=O����O^���O���O��?y�ū�Q�ڼB��U�m���� ��$���`��4^d�D�.OVlG�	
B���F���W�fu��|޲�$�t�	����"}2�n�j~��tw<QȒd��0��E&��'�(�V�Sğ`˱�|2V�b>牵ZP��,��(�����:��#<i��iv4I�vP���IW�)�)&�h³*�?F��D�$�����Egy��'j�VB*�T>!0Y j����dSlлfc���Edԛ{�0Y����n�П��ԕ|"B�1X؄麷�Y9w��HZ��U3�x2�h�v���.��5+͒lL�]����k�(��wM���DMP}��i�.���lQ�G���1#*\6H�zm���ۦ!�ٴg6�Dk�4���эq�����J��˓j�h)��D�d�*�2�@ݧ|r�Γ���<|O0�@b�ñn�HD�뚣q�I )�ئ�B�	�Iyr�'���<mz��*CNV"`0���䤓	h� ��2�M�MK�i80O1�
@�v���		~bQ���6H�u��C��c��d�=��q��bj�O�����	�v�vJO��L�` %���ax��yӴ�[C��<a��|����O:i( s��I�;D2�2/�>�Կi4�6�UF�ɐu ����/���(�D�3���\ �q��h�"]g��IH~b���O���yѨLCIU�X�ƅZ��݆*Ex�ȓ2�3rg'6N:M� �-�&���?;��$T(I'�ɭ�M���w��{s��G���[sȉ� ��'�t6Ӧb�4N��5�۴��d� z���}o@;�@��fl��wQ�i�]��f-�d�<Q���?���?����?1%Ɋ)��cF%�(���O��d�ʦY�t�џ ��̟�%?)�	�oT���&/I?:Ia��)�2zl���Oz�m��?1K<�|R�L�>��X�| J��T�29�4;#C/����"+���0����O��>�	#S'��;PY�"ʬb~��"���?����?q��|�*OP�m��8�b��ɵ$�`m�`��"w�d���~��	5�M��>ɕ�i��Di�h�+���T��@XrƘ3.����%�B�;��74?ɷ������.�䧛�C����[��Ŗ1I��y��O�<1���?I���?A��?	���j��d��=���"N�
a��=�b�'j�/i����7�N�����'�P�D���_㈅P�F#I��<o�����"�O�$%�8Dd�&��H�D�Z*v�8�5��_��kB�O�c_h�R��'�(�$�ܖ''��'.��'6����E�7ni[3!�4 �����'b�Q�D��4~HL0+O0�d�|"b�ݲu}f�ӆ�U}Fu� @Xi~ⅶ>�f�i���/�?�Qr͞�N�!3d��:�s�yy����w�IsC]��S�Dbb�Mg�DՂ���B�N��$Z4�W�2�� ������	�x�)��my��x�vT���VQ�����?x�V�Y�k��of���O�o�J��G��ɒ�M��"�8W�<��oQ�t0>hʆ�@ o-B�i�H��i���*�����O4E�'E��(V,�4!���h�Y�`]H�'����<�	x�I�H��v��ԭ^?���t%R�W�@,b ��VX�7�;?�����O��-�9O�mz�
d N=v��C0Ɣ�N��ُ9�R�'�ɧ�O3���G�ik�� Ap�H0�Պ:6���Q��`���4)�p�����(�Ot��|J�S-�XI�Ǉ�!n ����'�d�B��?i���?	(O��lZ�u�b��	����	�~�\�-#Zا!�&
A:�KVh&�I&����O��7�䆳H����Gi�f�d��$E�k���O�����\�4�F����S�Rr��͟(�CH�!8�z`��C��c�<��T$�(��������G���'W��`��X�f�T���E�<����'���Վn_��4�M��w���6C@�O�D|�3EzW�@��'�B�'i�,�rS�&<O����,8�ة��Z�� �9�$ �U��黀������8���<ͧ�?���?���?DK����5�F�F�TP�ˋ��$���u W��������&?	�	�GB��Y3���Ts�l�2��<����O��n�&�?�K<�|"Q���R�!'n�:tf����Ʈ$�ވq7O����c�����cPƓO��gM���20أ�lKUxț��?9���?9��|�)O�nڤ-?�)�	�>�aq�ǉ+H����錸c�|��5�Mc�2Ź>��i"���o�d蠐'�ԡ�e�^5ZL��1��w�7�"?զ� <�	�䧘���$���5a�4/�|�RD���<i���?���?����?������,�&KV']����GD2vJ�I��4.���O6|7M5���P��)�r���|Y�Ο�v�!%����4/��'	" Bߴ��$�(�
@#�I�16[$�XuI�dТݹ�5�?��e;�d�<���?����?Q��:<�Dd���;;Kp	����?1���B�E��i�؟H�Iߟ��OU����]�;�\�T-��w�&h��O0��'��'�ɧ�	GI�a�En�p��= '-U�>4���d�)�
ؠ'�<�'`�����YT)A�`��H@i��T-:�t����?i��?9�Ş���YŦm#�LD�e�p0����!xNv	�dݾ�F������ߴ���?Q_�lB�4o�b��r�`G�´ݬeW�)��i[j6�M��6m5?�R#ЖqC��ܬ��d��"2v5HF�T���tc�{��<a���?����?���?�/��t�i�l^��cKm�����N�m�i@˟h�	��%?A�	(�M���`$�I��xsR�-��Y�����M!�i �O1��ܠ��x��扦b��0�Bn�	c}`�+���ɒ/��P�'��&��'���'mV�J�;@
!F@�'��K��'���'AY��rش<�z�(��?����*�JS���O,�ӯ�zU:��H>��@Y�I:�M�Ĵi�O"d�	�~�:Io�
TUp`�R��l��"^�݀d�b��V�����ğ@0M�uҖ�ö��5q|�۳��̟��I���I�E��w�i
E�ܶ �(Upa��m���Q�''V7î+/��D�O!nZI�I��$a�F�ɥ�!�>�����yX��I�M#��i�x6m�N�6m7?�Ń	/ ����(rW�%�CdT1��CTɬ	�j�{M>a,O\��O����O����O:�����>k҂�j�&�#?�L��ʩ<��i���%�'O��'��OE"�ַ���ąN�4��H���� ]�v��?�����S�'���`�ϕS$Py2�ܾ ���2�H�+�MS�^��֡�G���4�$�<I��A?���@@�B!����A$�?a���?����?�'��Ц��Er��
�C�#Py�#��wN�1���|�tZ�4��'���?a���?!QgN�x�� � ��Sk�!!2!Ъ�@5(�4���Ȅs�Щ�����#�� >�tI`���0+L��V?O����O��$�OT��O<�?)�O�l��g���". (J��|��IΟtI�4I.`��'��7�+��V�V-9��D^��2A哀pz|�O����O���3&@N7=?��mYwn0�H��Fb��b��m�p`����X$�4����'�R�'֞��W*�x0�!s�^ �@� �'�"S�Pc�4�����?q����I�*��!Q��ػH�h[���b��I�����O���<��?�[5�)�h��
�@�Q�lݽUu��P��æ1��$`�K?IJ>��OU�5��tX�+ڣ7���0�K9�?A���?���?�|�(O�n�%�����T�u��ԁ0�L�MI��j��<?�Ǳii�O�@�'���L��D+)5���u��&/�2�'���0#�i��	 Zu)��I� ce$���DH�4�q	-YE�Ģ<q��?���?)��?�-������TI��Q��O��j��d�ݦ���
I���	%?��I�M�;B=D�(�F#c�鷅�0U�Y ���?)N>�|
��ɕ�Ms�'>z��욭G�\���3l���'ͮa��$Iu?)I>A*OH���O8}�" �vJ����f�MZ!���O����O��D�<Q�iX�I��'���'�0�%�C�0#��(�R����dMI}"Hcӆ����I�}i�@ 7ܓ0�X}`u`B����$a�$�� -���I~�Dj�O�����<��MS�AшU� -��"������?���?���h����T�HL8���� o �X�珂�~�R�$�ݦ}:4)�Py"d�Z�杽d|(@��4$���B� 3q���ڟ��	�d���
릙�'��| �m��?=�!)�1Zm����O;1�r��W�G��'��i>U�I�$��؟��ɍ\mJ��W��<YET��b�!LV��'��73�
�$�O��D?�9O,=�@���3��X
����m%q���?����ŞH��Ys���,��Q�/8X���m_dê�0����(��[;*��fAV��{yb��q�<�k_Xq�"/۪5:���[�X�I�4�i>�'�*���]�2�J�6\BIJ7o%Q�NYSs�Ԡ�yB�u���@	�O����ON����x��Y5G�ܜ��e�e"���ԩg��T(6� �d�>��]-8�eac⏛)�B�Y��2��	֟��	՟T�I՟��T�'as�8YC���G��׊ݓ�*8 ��?)��c�vh���I��McN>��
	9Zl�$GS &�0���	����?��?yF�� �M˜'B���� �d�&A�U8B$`է6,YUO	��?�P!�$�<�'�?)��?�Վțe��a����SҎ��ul��?����D�⦉w���	�ĖO@���D��ljb	 �Gt��4��O���'@�6�ܟ,$��>��#�H�}8N+�֫q�|��j 8Pӊ��cƷ��4�zU���߈�OByie��U�h9��͗�*�p��O����Od���O1���H���9m�΄en�=&�ȷ�0F ��V�'���yӰ⟴�O�n86�TJ�j�w�`��I�.}q���M;�����M��O&)۲����$�<)���d�l�Jv+KA,*e��+��<Q.O���O8���O ���OPʧV(<x��S79"y��n	*����D�i�p���'���'���y�{��.�X�Zh
fL߽Y9>`���R�jEr<lZ��?�O<�|j1�M�'�"$jԎ�1�8�pc����#�'�hـq�����1�|R^��I��l�#&V12 �:B�[��F�&��̟d��矤��Dy��oӮK�m�O(���O�0�7��>o A�m�*M��;�-(�	5����O���"��l� �@ß A�@� MԌ
;�	?AҞ����߰Fb>�Ƀ�'F���i|��wh�@�l��/_%��d������	�8��Z�OF2�9Ka�a1AɸC�z�BG'�6,?2�pӖ0se��<���iP�O�nAt�,K)[:aP�0�RM^.f+�D�O2���O*���!m���3T3�+��ġ�CL�%��x���\G��ɱ�k�1����4�����O ���O���**b`�!��x5ĝ��HՑB��4�"ԬD�"�'R���'�����I'*tM:D�I�Nie��>Q��?IL>�|�D����<�J�
�dm	N<~��	b"��h~2�"x�Fa���Q�'�剋j�53D@���]�-�g#:��	������i>Y�':��$�,�j�Get���Yf|�MCV��%�y��f�⟤ѩO8���OV���&I���Q��#�t2�����8�s�u�b�{���
����>��]�K#L����)AW�XW��8\J8���|�Iǟh�	͟\��d��Q��a@ט�l��.u��I��?��6}�6^�1+�I/�MK���䊿59��K���֚իԠ��La��O���O.���
6
7�y���I;r0ڒ�ܗj�:%	�� GV�����'-l��R�	fy�O�R�'�ҫ�oe8k3�X6��
t��Z���'���M�֤�7�?����?y+���eNAz�1���6�)�����Q�O\ l�M��xʟv�Ru \�7OޤJ������[���+c��@'A*f�>��|�P��O�ɢJ>�a�Ǉt�H�V�C�@aH�.�;�?���?Y���?�|2-O(m��� Ku�۬`�D@�3�G^°��#�x�D�O��m�F��l{�	ԟ�ZGbT�
��A���Kc���<��%~��8og~ZwkT��ԟT�cs&�f䀟uu+�`��7߸q����O���O��d�O��$�|��V�^yӁ/S/)�0��!�ɥXm���ݪo>b�'3r��t�'��6=��h�"I�>�ݺ� [�r��<�f�O���0�4�<�$�O�e��a�<�Iža# ��	���{�������6|8�8��O�OR��?��vc�(�+��p�L5h�	{����?����?+O��oڤ5�,�I؟���)S2����>��a�ތ.��&��������Oz6�C�z|�I7̘�ͽQ�+X3s��	P��Z�,ރf鲡$?UzS�'沍��Y��UQҧA�����҉0
fe�I؟�������R��y7`$��M��+ͨ+"ػ��<G
��pӨ=�g���ٴ���yw�H|��� ��P9N��u$%���y��'�2�'g0�:Ҷi��	�~;��ݟ�ъA�׸=���g�VX|ةQr�9�Ķ<ͧ�?���?���?!��C�s4�,k&�&qm�x��CɆ��ϦIRF�k������ '?�'R�}h��*KT��h��"'Zi@�OP�$�O�O1��y`gm�(y��ܓ�B5Z��)��R�4��6�7?Y�gL�ZH��IU�	my���k_ ���=&��q�F�3JSB�'�"�'&�Os�ɨ�Ms�R�<��کp���6fÚ �aVc��<aӾi��OЅ�'���'�2e��g��i�b�*�
hx2nT�64t��i��	�Q�������߭�3DL�q"�8��G�V��m���Iß��I՟h�	�P�����
��8�	C?Ja�1 �/��<����?	ղiD�d��O�pnZi�(�}`���3c���Z��$���&�L�I�I&z��n��<���\9���@��Un�b'�>���[�#U�����W�IOy�Oi�')"��'R��c�f��*��\%WXb�'@�ɲ�M�n�����O��'=���#k��4�ڌ��DD*C�B=�'�4��?�����S��`Oh*�-����uPxq$*��=�T���1alx��O�Ɂ��?�6/*��T'4�]�>���HD�
(bv��O��D�O��<��i�́�i�jjΩж	O�a ���䋏����M3�r	�>i��u�}h2Ț�z���n��eY���?0�&�M��O�����E1�K?9�@��J��)`+I�6��'h� �'-��'"�'#r�'~��N�V�;c���l4:S֭JiL��޴!�����?�����<����y׍��/
���p�FAd�|�eVu���'3ɧ�O��lӀ�i��� �XE�W�d�tX�Ղ��e��7O~%�$�ŕ�?y�	?�ĥ<�'�?y%���Ԙ�6��?p���	S���?���?Q����D���3�ry��'����@����M�:2�18u��Vs}��'vB�|� �WD�zv�+v�v������-~�f�0�wĎ|̧R�l���<�?�Ż+����T%P?��ۢB��?Q���?���?��9���9�+C',V��P �$l׆$80��O@Doڔ[�'d�6%�i�5�5+�-s�N�:�tE~ŢQ�`���Iޟ������oZL~"]�_�j��S������`�>yUvMy�f�X���ҙ|�V���ɟ$�	П���� �7}r	�"%��T���Dgy2cӬ� �`�O0���O����T'@f�jS���%�<`B�	ɬ\@D�'-��'Lɧ�O��de�-^$t3��̇aц�x��P� #f��O���j�!�?!1�+��<�ʛ�zcB1zDD,^����b�X>�?q��?���?ͧ������4�џ8�6���,露9��S� U�a%�̫�4��'w���?����?�e�ɓ:g�pXb-��6];cm�S�Y��4�����nPb]`�O�O��#BYf�0�g\N��<����y��'A��'�r�'fb�i�2~��
'�$\�����k�"��$�O ���Φ=@'C�|y��sӆ�O�� ,ֵT�4x1�h_��8�貀<�d�O��4�����or�.�Ӻ��$��Y�2��<b~VTJ�*M'\ �8Q�'D�'g�IџX��ԟh�I'���D	>O��LS2
H�K���	��'��7mU�
�p�D�O���|b��J9D��D�8p$���I�v~⃩>���?�L>�O�$�`Cn;L���� Ȱ�K6����b�i@2��|b%D��@'���Wl�<2��5��!�G� �P�G.�h�ݴ&�� ���F'Z��K�^�y8�����N�������?�\�T���9�T�����<��L�E.��X����h1 /��I�uW��<��	�<�rL�l�r����8�8���E�<�.O����O��D�O&�$�O�'8�j�ҳ/�; �8�P0��)��d	b�iZ�p'�'	��'y��yB�v��.ڷBP��
s�J!)��z5�˵V"���O��O1��i��
yӜ�I-��sb��$Tj�@�j�]Q~�8'�\	J��'�&%����4�'6^��̢eT�8s��_�0\�r��'m��'��T�pIٴn��i��?���K���K��Z&�н�6�J�f夼���$�>I��i�"7Zd�	�:�f١R@<!|s'� y)��9xP�p�'�M�L�M~B�g�OR���)���kRi��}`RcЭQ��:���?1���?���h���d��x8��s��"{n,�V������[즕У��Ly��mӾ���� L��c̨4�-�! 67�Ɍ�M�i��6M�!��6!?y�'�hz�i�#��d7 W�$�6U �TaH>	)O���O���O��$�ON�be� ]Hl装s��P�B��<�q�i(xi+��'��'��y2����#e�T(�0�'��.VǦ�S����a� 1&�b>���kK	�0���e�`�õ�ɿF�-���Sy���'�A�	!@�'��)\2Ŋ$%��Ts@����-p@0��I�(��矨�i>�'��7M� "���D� & �Ȓr��"E$5�V����Ĝ�1�?#[����� �	X\��@̃�Nm�m� A-'R@������'��� �#�W2I~��;l��i
`Ş�k����0�U�.�0���?!��?q���?����OR �2r�%83� ap��8�?���?�ǳi����O92�m��Oby��ģ��Q9V���x�L6���O(�4�J�{�isӚ�Ӻ��&�I���@�/ï����@J�bV�m��'P�'��Iԟ��Iӟl�	�
�v�Y@k��I�����(ռ1?�L��՟�'�^6m�e�����O^�$�|�&� ��h�hE*W)�����P~rb�>����?J>�O���2Dܮ2�H�[Q�3��HYV� 4-R5避i�r��|�꩟�%���F��"�;F�[.7��d�ß��	��P��ןb>=�'�7�������&>����"�� shL�
b��<�ֿiw�O���'B7��3Wj�!�S�0�҅r򈕨=[�Tl��M�wc9�M��Ob�2c��Z�ȼ<QR煃t%)	��!�����<Q/O:�d�O����Ob�d�O˧(��J`��k��u�u�Y1���pA�i�2�!�'��'��y�q��WL���K3��?O�00sk�E,�dmڊ�?�O<�|���J��M��'�hj�mZ/�L v��V�̠�'ئ���ğ�`��|�_����Ο�1�K_0��}�"]�~���ҟ ��˟��I]y��e�|�I�+�O���Oh=�"ͅ�YV$�8q@ϕQ�V�"�E6��+���]�I���ē�Ah�&�'b>^9�G@/hn���'�||q$�I�LQ�<��������l�!�'�uCq�� ���3��3PDN��p�'���'�"�'��>��I' س�aH�Aը�:Q�Q,4X��0�M���Z���$�Ϧ�?ͻ^u>�C��J*#Fؚ�dޚ���d:�F�O�6�E^�~6-=?��d���<�iQ�q z���$�"�y�Ҡ�,BrPM>�*OV���O���O:�D�O�	a<X��`�b�
�,8Tx$E�<�B�i�liI�Q��	Z��؟�#��\�2?<�*��l��u�SA���Ē٦m�����S�'G�@�� ����?n���T��S֎�K���,GT�˓%#�X�6��O4Q�M>�.OD���\�%�~�����1.��@�em�O����O����O�I�<���i̾Ժf�'j Uc+>�"��!��B鼰!�'�N6M2�����D���%���M[Bg�(3a�K3�1k�ޤ!	�����4��DD$l����'-�B����N >�3�Ua�d,�g$�Z��O*�$�O�$�O���6��B�8|����XN���1�B����I֟��I�M+��|��}��f�|��Z��D�W�ʬ0��ȧBeM�O��m���?�S'	mZ^~��Z����ض�#e^Q	��9u��f��̟l���|R[��������I�|��Ň"~�Tő@��-�z 2�nV�����[yKq�*]����O����O˧c��X��l��)L����']:�|�v�O�O�S�b�� �"B��&t!V�- �(MY i�8C,���@kAEy�O� ��	�\�'�<�B��^�w�Xl�g-��VOЭ*��'T��'�b���O��	?�M�!õd���@���8 �VE�7�a�6Xk���?y��i��O���'"�7MO�IA����%Ͼ4ö���HϺ@�4U�	릑81�צ]�'�X%�r���?=x$S����'7�I
����K���e*l�`�'/B�'�r�'��'�哱oT�5�&A��l�]l�tN�ܛܴx�,,���?�����'�?�T��y�L�3`B
q���<`t9@�L0(J"�'ɧ�O,�!�F�iH�Wr�(�HgH��2���@W��x����C��Ӏ���H=��)4�ٚJ��Q��R4�09i�^�H����O����ؠl���� GB>S�ƤQ���8GzP���#6�Ҧ�B/8g�׾P�fI��AO$g�vĐ3e��Թ�f�D�B�����-�
m�p9��O'��d�j�BD�V�T��8�4�$s\Μ F�F1y��Y���# �4Qz[��e�N�˲�7�[� �DgV���P�r�D6J����&��A`NŪ�H�#�b�õ
.��4�)dX��mӭVb����H�g�4�)���g�v�F�Է�~���O�ciV]o������R�����kܥ�EԿ_Ū��۴�?�J>��?	��ݵ��'&��k��������T.(1�4�?�����D�"� 8�O���'����Y�f�`Ă�b��Q$���d�RO����ODekD3�ID�!a�(��|�ԥX'g�0����ɦɔ'����y�����O����h0ק5f(NT@�;�#��G��-"Qb��Mc��?q���9��'%q�H@����/%# �!5��]��x�ib���%d�����O��D�T��'���"ol���i^o����D�	}p���4,�lPk�2���OT:�AY n1�Bǆ"3�M�wm�̦�������� ��m��Ol˓�?��'�,��O�f�l�s#J�#=���}"F�$(�'���'��ҊG�)zf�J��\����
6��O|�CI�R}P���I^�i��kք\�1BP����A��P(�L�>i��/�䓾?����?�.OJٻ��66^l`)6�]�I�\���E�::�`�'���ܟ�%����ܟ�*�_�
	��2�u]&��lv�a&��	؟,��^y�a��T����[5t��a\��,�Ĉ��RR�6�<i�����?a��R��M���"��9��	:�0����+��tk�[���	���	cyB�:k�'�?1���~EZ�x`⍂}�zɊRJ�����',�'4��'�ZLx���6�rp��	�дKZ_���'O�_��G�!��I�O6��៘dP��ڀyk��W%^�X��I g�u�	��8�ɛ:U�L�?��O�>=��k%#  u��q��h�4���-�ƅoǟ(�I�����
�����H�&+S"KfZ���ݹ2�`L��i�r�'��`�&�d(�Ӏ�>�G❮h�x  �/Â6mD1���o�ߟ���,�����$�<Q�!��*�C.�)S`��CU�G@���S?S~�|����O\�F'�%����7��(r(�Z4�R̦�	ޟ\�	U�D}��O�ʓ�?��'�XizV�*dlh�q�N�~�⼐�}�і-�'yR�'3�陛k��u��c�Ƞa�P{�7-�OA9rL�Y�i>�I@�&xF�;�ڕ����iF&(�)N<y�����O����O�ʓ;����t◀0)����w����R"�:$�'�R�'v�'��i�Y��$ݮx���UA%9P�:p�v���d�<q��?)����u��Χ~�Hr1)�:H�.�ca��-k(`�'�r�'��'��i>y�II8rIQħL�%L|��O*VG�O<�����d�O���|��.�8݊���hR�$� ��H��M2��i��ON�$�O��3�b�8C�'�0�"L<o�@��g�C�Z(j�4�?I����dG8A
�P%>����?�طE�7�XE���w��ly��-��<�f�%�?1M~��O��S���_�r���ަ{�t��O
�$��h���O��d�O����<��h$Jf�W�3J|DiRu��j���O6Ƀ6V?
E1O��҉�co H��ö�L�O�,��6�i�t���'�R�'��O��)�cϞ<�^�I�h,H;(@� BO&��!� +6�Py�y����O�(Z��W�T�yR��_K;�
Cc�Ʀ�	����Ij9j��H<ͧ�?�'��	�ڰq1x�8%ܯh)�]�ݴ�?.OpQKW/Gl��'/��'2,�H�)3�'V�J.IてBO*7m�Ou+E�a�i>=�	񟤕'�UӲ����D���L�F8�r����ȅa����<�'�?Q*O��dL�n���r��1�d���0�H��U�<A��?)���'d�6� �P3�^�,��u�EJ<Qb�!�i�J���'�2�'��U�Hp0(�-��īѪ��Չ��^�E�N諕l�,����O��$�<Q���$�"Z:���?&rl���%$h~	:B�#M���'�b�'��X���!͕�ħ��I��܆@v�ip$W^����i�2�'�Iϟ��	�5|��Id�i<{�9�ͥ^Y��!AKŢ:қ�'K�[��5%���'�?���C�Y�it�������K�ݚ�gK�I_y2G��h�2���ПH#f��/����Q�~�L�cW���I�n�	��Οx��͟���pyZwF�5���l��Po
�޴�?����!*��^�S�'H�,����% ���
�J`��n��:����	��8��ПX�lyʟ.��@	�8m��Cq	:.�SR�e����0c�"|���W$y���Z��0󔦍�p���c�iQB�'�A�y�8O�)�O�	�d��ex�iQ1g��9#��ؖ^��7��O<˓o�<x۶^?�I������ 7g?�U��k�f�����Í,�M����©��x�Oer�|Zw�̈�'�@)(z�H�f�A�4��Or��q��O�ʓ�?�n�ʟ\�'�.MJS��%8�m' 8Z$P�R��24]�O����O���<����?�!P�0+�d������|˥ƥ4|� h�����Ov�d�<����XB�O�x ��I0W����Ď�
e���h�4�?!���'��'_����M���M;A�E�z�H&�Q;zx��M}��'���'���&=�f����EL�l#giۉJ���2TE�pAP�l�͟ �'��'62+K��y�Q>�&(�+	�r�A�\%=8��㮁��M[���?�,O���HD���'9��O�$�é"aA�(ڃ�,0D�#��>���?)��m�.�����m�:|�F�Wc[�>vv��K�M[/OXU{��P劣������	�?��O���v��i��d���U�Q�Pw�6�'�҆ϗ�yR�'�r�'uJ�)��)֗E���yv�L$g��o�1�4i��4�?a���?��'q_�	Yy�Mي^���q%
�QI9�r��',�67�����}y"�)�OH�����>�4�Y0��6D�E2am�妙�I���ɓCC�͡�O4��?�'���{���~�L �q�-F�<T�ٴ��tm���S���'�R�'���0l�5��ma�O �|t3xӄ�DG��'X��֟T�'YZc�X���(�eR�Ӣk�n�*�O�X��9O�$�O���O2��<Ic!=
q&� E��)g8���l�"h���c'W��'��_��	�����#���������y!��ZW*��C�z���'ub�'��W�P���Ҳ��T"��2���Z�Η*8�X25 ʛ�M�-O����<���?Q��/W��'���yT	ƚh�v��GF1L��u�۴�?����?����dV�{����OTZcZx���N$ez�e�bB6�Jڴ�?,O0���O �dǷj���O�	&��z���B��$�υ<c3�6��O���<�.Mg��S�����?� �J�LY�l�p+I0(�t�7/�	��D�O��d�O8	�;O0��<!�O��!�`�O����q�T�g?8�۴��'�60o��I���Ӹ����N���g�wW��{G�M>���Լi���'�X�'��'���	O�AUp��$!�2 �� ��ԍϛ&�_�V&"6��O���O��ɛD}P���� w�j���ou���4@Y��M���<J>�����'
 �:��B*�8}�`��\:m8��~N��	���	�E~��O.˓�?�'���H��Ѫ,��A�� �m/�Ԙܴ���O6��r7O�ҟ(�Iݟ�Hʤ�`�j �E1U6��C����M����v��Z��'~�R��i�]�D�G)=��0,�����a�Fo���d��K��O����O��d�O�"+F�����n���Q�!��b�˕Ƙ�p�I`y��'��	���I��h󄑪T���S8�@$a�I�,Y���ky��'��'��:�f!ӚO;�HE/R���풊W!��4����Orʓ�?����?�j��<A���e+'����(���T�Tn���Iџ��	Qy�Ȟ�^��'�?�1�acvş%&�p G��\ n�埴�'fb�'�rh�y�>��Ϛ Q��;�a�m�:������H�'2�A��#�~���?�'c��}y���,qu�%* �?�6��U\���	��4�ɠ8���	x�	o:$*(�Ƙ���E"z|������'�B��c�w����O����֧u7��z8�yaD[�\�($��'�M����?���Y�<�����D-���0��1 �6KH��1,���:7-;��l�Ɵ,�	��$��	��d�<A�	� i<i�����RJ��2�
�V���yb�'A�II�'�?���@�K��ɠ���3]Ĩp4	�*��F�'<b�'6v�Y�.�>�)O��d����ć��� ���7 �Ӡi��O�B�1O�Ɵ���ӟ��6�+-L4��&��K��lNƱ�Mk��@pv�CBY�<�'��U�8�i��01 �1����bFϓo`�,Ʉ�x����aU�$�O��D�O<�D�O�ʓm(�,��ce�>��'��X%Bg�R�~�����O�˓�?���?� dN�DŶh��Ǘ`�"���� .}�����d�O�d�O2�-�4��7�`�2 _&fZ0܉7*Ֆ]E|Cg�iP�	䟠�'Q��'��@C$�yre�:!����������&��6�OV�$�Ov��<	��
,�����aA��P��۴;��M��0Z�i �W���������*MkP��k�� b� �F��+-K>U��J#�i��'$�	!OT� SH|r����@[�Vy
A)�Bٙ[~E�叇�W=�'���'��P �'a�'��I�>/P�����DC��!zf�%Rʛ�U��Y�)Q��M��\?Y���?��OZ͋$� je��Ȇ�_�g��X�i�R�'�8C��;�2����f]�w��e�(�t�b7��nAh�o�(�I�`�����?�'�Z�tq���ʿ��ᇭ׫=t�6�W5L���|����O��)�F��FD	��R�
�K�ݦ���ȟX�I^&rɡ�}��'c���VP{�R%,�x5Sw*C�CZ���|R�=�yʟ����O���A3p��}:'��C#J�#N?c��Qm���P�5ND7�ē�?�����[���$�N�C�'S5�t(�(�S}"	8��S�d�	����	NyB�V�v ��!G�N��Ifᇽ?"�``�>��П�'�\��П
4�0��5Q��+X��T!g�se�	Ry�'���'I�IN�P�O����8����j���O:���O�O8���O2@cV9O`�aΟ�(xvab��ƌmq,���c}��'��'<����u�I|�ߴ��ۀ�C3ZT8�Qh��&�(6m�O��O��D�O~aB�!�I1*J>1c�F��b]��#3
NT�7��O����<�TQ��O��OZ>���E)
j�чʙ@�h�G�;�$�O��A���D#���?!	c�T���X�t+����Da��z�n˓d(�a@�i���'�?���|W���`�;4.W�p�-�W��tw|7-�O���_,y�����}r�(ݏy$|��4)��H��6�S	�ql��H���<�����'�~�0r��uִT�VBԓ�fx�@lӐȉ���OL�O��?9���v���#K��8�b�M�5��i"�4�?Y���?y�"_=1G�'���'s���L.52ɋ�0tܕ#إ^O���|�� �yʟ����O��$��+I�]�!G�1IXT����BÁ�̦���7�P�J<1���?)N>�1#^�4[��"+K<8�Sꚼ+@�}�'�ڄ;��'��	ԟ���J�F,���g��4��`+ŋJ�vH����	����?�����?	�"&�e�GN��,!���T)�8Wy6qhb*�?�*OR���O��d�<��AU�R��iւ;��D��M�`&eY� S�Q������f������nQ^��I�~�T�������}A �[�F8�;�O��D�O�$�<�ō�[�Ol�����:s����B�A	���o�\�=y��8�@٘���?��'T"�2�%)�b�GbG;C>�)�ڴ�?I��������O���'���
�0P���&XO�-������?q��?1���<a-���?jp� ����g��>~�qh}���N���v�i���'���O*�Ӻ2��Og*,sBDӦM�ԍh�E�ަq�	şr��x��ث��$3�ӂ5[�$�#!�3�� ��֢�6-Vs~	l˟��I�ӑ��$�<s�#"�rRl� )%�[G���@�����yr�'��	Q���? "D�ij茀�¢0z�cź0/���'��'�@5Q���>�/Od�D��9J��:�$�� ��E�:��Hw�L��<����<�O�'�Jǿ/p��f-��}���SB-�2Htp7-�O�{��Ms}�W���_y���5�N�1Q��+��&Xu\ĩ��޴�M���b�ܑ����O��O�����'��q*zM�,2>�"�� %r�Ieyr�'Y�	����ş0�"�M`�*wk�]��r�J%\�?���?����$�)y�8%�'h�T��b�ʠd8Tڲ�PCڐo�Hy��'���ȟT��ҟ��BE�~굆�u��C3��$-�����"�O}��'���'@�I"&1d�������Rܩ���U�)>��$�ӆjR�dl���'���'����y��>ӃœN�Daj�o��kF��Ŧ�����D�'�|��A��~���?i�'O.���	Ǌ0�b�LL�
��8Y�Q����ܟP��e^T�IY��'����!O����U4�p�,P�6T�h��@��M�4P?q���?% �O� �VK �K��x�B�p��i\�ɩ|��?�g�/�i������5nX)#�7M��A���n��ȟ���/��d�<�(�9��J�k__{LU lVBǛ-F��y��|B���O@� %��ԁ��#P�����[�q��ӟd�ɞRG��0�O���?��'{��@!Kв ���pT�%r�Rݴ�?Q.O؜�6O��ß����@�$�4�sF���;{������ �M��'f:DW�,�'/Y�(�i���B	`̨q�K�� e�ln�*���9��<q��?����򄈃��0+7�
`@L��I�8(��E`���s}�R�L�Igy��'�"�'q����G"L��e�ɯ��Qvĕ�����O~���Ob��<��.ĲW��i^�9����e-��0�WhG�"��W���	{y��'���'g>EP�'|X�cg��Jf
$9G`� &} Y�2CzӮ���O"�d�Od�[X�c^?��i�	eJ3crk�D�=��{Ѡuӎ��<���?1��b��ϓ��	��U�t+̮K�[��,907��O��d�<��(�}��������?	��*
T�(�ޓ[�8�glݦ���O��$�O蜚6O���<��O�� #�LW�.u����bB=ڮOH�$ɢ3����O���O����O���3,P�m�&.b�j�� &
�t��7-�O��>�:c��� �u�Î�<�&�;P�Nm8�,�b�i5Đ�G�tӪ�d�O����8�&�p�	vG�}K�i̜Kzhс�
�%����۴W�$YEx����O�%X�ƞ)/��r4�Y
/���˝٦���ҟ8��Q�zY(K<i��?1�'Y���P�N��MX6!�A�J4���?���?��؏9$Z%`BG�'	��IqHɺGߛv�'���7�D�O��$?��Ɣ���dVi$k[1r���ٷ[�T�gG'�I���������'Hl�ڴl7QP�&�)1��1N�#M3`O �D�O@�O"�d�O `�a�>�ڨkfc�#|����aJ69G1Ov�d�O����O��D
p���6P�p�+�*@ ��	��ux7M�Or�$�O�Op��O����B�_�֠�'X��d+��.J$�)0�@����O��d�O0ʓ`��ԃr���	VND��CN H(� -��`|F7��O��$%�	;�~c?ћRDAG��j�F�ex�l�DKw�>���O��$�O��0�|J���?���*
>%��AW��d�gˈ�BK�� ƙx��'��Ӥ{h�1�y��:�胩EN��ɂ�J����i|�I�u)�%Jڴw������S�����"2����uI�a��sv�-��4�?��c��Fx����4����gNa*�ũ�J��K������6��O����O��I�_�zI�S��2OԈ�'�A"]�H���i�da2��d/����l�h���sS�_mV"�.�:��f�'t��'�0�R�m1���Oz����4�b� L�[�dͦYѪE%�/��V�Pc�(�IßT�I�u�~��	�8����E�C�R���4�?QV�WR�'���'ɧ5��V�Gw<�b����X��Aϰ��$H��qO�)�#"��O��8����)P^Ls�IU(B�9��'B��s��`´�cR����
���=O��1VL�;#.2eɠ�ȥYQ��Ao×"��\2�C��VY�(A,χ5�^�m%�.%\i�դ�%��,��mȁ�
<�!F��b12�S�*��	��LH���MRnPB��[�@��؄��#4Rmpef.2���D��C�i��ғN
�%���q��9�g��_��FD�P��`���5\?���4O����'���'����(�$@�,��P�Юh1P�b���_B�C#k��$�2��:�vmZ`�Fu�'���
jN�\��!nH��v�[Q	/'�栳 	�r:���7S��
�AE�2��O:��R�'��)�?��xJӂ>ŎXI�oV�`�*�Oj�����;-��{�-�aLY��'�.O^�1����p,Ƥ��L\ 
H��04Op���Lz}b�'��ӞN����џ<�I2Z:^��geY�I�p���KȾH�e#We��M8�}�'�ޱ݄T��S���'��]rA�a��L��%ܩF_ ��>-� )����J:k��O?�$��'���9e�B2�:l��Y�a���ON��%?%?m$�,kg�2T���Æa�
�݈&�(D��r�)Q��J��bN��w:���&]h���' �n8SuMUܖX�g�u�@����?CH?)��Q����?Q���?�g����$�O�I��̡*����O��}��2�NR��\�OL ߚ!�V��1���I�:X�Թ��=L���k[0�8����#N�y�G��&�:B��?�=)wk��1a<�� H�g�茳��[?1#��͟���I�'$�I���d�ʝy\vLR�(]��B��:Ƭ��ӏk:�F���$������?��'^�i�C�q��R%iU=��h.Y�$u1�c]�%��'I��'%��X��'��2��ɐ�D��5d�)�!�e*@��Z��(1��H�-q�X��	�Q"��Q��C �ZT���c��쨧 @�H֠ȷ��q���1�O"O��@��'~�*�*j|PW�_��N�҄qK�ўtFŏ�o*�JM�<g��Q�,��y�FF�<��:��\Pj�8��W9�yҢ�>I*Ofhi��E}}B�'���&MX�[��[�R�P�b�*�/"���������|p���x���j��8b���Z��������P|�l�A��d�n�����/1�Q��k�W�g\Z����4�:����AhKD 	"q���ol��"P(4���`a�j�(+X�������,[7ti��*3-K��da���<Y�	O�=�g@_^5�gc�V����Ɂ��.���q�Bl�Lh��t3�X�<	�dXo��	��H�O�B|Ӷ�'���'�nM�ƢL� D"q۠#G�k���!���RCt���.V����(��OL�b���Q5,�������ՉW�ĸW� 0zV!߰]���`c�O?�$�0=�X�Hv��.Mߘ�!2ꚯs���ӯ�O��n������O��I�[jx�k�c"�]�ŃQ 2C�ɑl1D�#F��8*@i�Vc��e�"<iF��M3�bN�]��n�2j���s�� �>�����?�‪<��Q����?����?I���x�D�O|$A�e�2(��8�i]�Z�2�"�ʃ�+����M���3%��)3�'��pkd!�� ]� �UaP�p��+ �!�ߍ;Di���HS*��䇠%!h�q�oAQ8�����̲FK�M�}
�dfӢ o�M��#��ӈ^Hތ�ai�1LtH��+ �xB�)� x!����	ZČ��'F��\쀢i�m�'���������
�16���Pğ�#��t���W�<)�a� Bz��`��]_�=2��[�<���U�:KX8iP	�3�Y�� _�<�� )	j hzF"�/h\�A��P`�<a�Q7y��� �~ hT�Ha�<ၩ�1a���i卙�]j�hyN�[�<q�FB?"����S�7��-b#[�<�R�b����U�-z���b�P�<��i�8�d �%V1�P�W�<��¶TءR���  �%��PZ�<!7�
1׌Y�N�1�,`!�G�a�<��d�*bܼ�p$��)c�k
D�<A�^���h%�<!�ld���JI�<A�f^<L�B�ϝ8�����H�<IN�8f7r�+2��R�J�J�J�<a.T�O=����*���,e���O[�<���r���&��J�z��,�]�<ɧ�՘J͆1 `�Ѳs5ԑ�'A��<!F�P��tJ%hT�9���� s�<y��G���Cіh��RׯRk�<���lf\�B�`S>J�&(I��e�<��`�8m.AT��b�� �[�<YF/M:q���gjE;��{���~�<�ەf	 I���42�8}�$�b�<iq�_h���qr��4dl,�e�w�<�7�ݛbV&��$�˕ۈ�:REu�<iPE�x��@/NآU�f�i�<1BJ D���+T�O9֐Q4�EQ�<is�]�b%��h#� m����N]L�<q����#�]�-�,��It �c�<�ȓ2ݻA��@/P�D�_�<�b����dcԌ�}Q<u;�m�f�<�Gk�~��C� ^�r�LFa�<��$����H���
�{��-��$�\�<�s��X�����3*��Tc���V�<�w�҃
�I\�0�����P�<�u��<��ذ�[�'f���`�w�<ap+�)H�NP��"�)kkֈ��I�I�<1�I/U{��6E��A�n!���E�<����~��3E+R�u��i��(Kw�<���;IH�]�%b�6B��u@��u�<���Q�`Fn�+� �P����LXM�<y�/�^>�q��'����F�D�<�p�æ4Y�A���ث"v�;q\�<Iq���U�RDH'Z��qf�X�<��mm�6�cK�����V�<q7�8���!�f�&J�58�B�G�<AV�Y�@������% ]VБ�HE�<Q���:��z���!0tXK2�h�<�C�:D.m�U�Z
Q��+�a�<�b�,V�� l0���P�dV�<q����W^�i2�P��>�(���]�<	�O��2��
u,A*��Ԫ�&c�<�1j�.� E!��
rZ$Y�cn�a�<�B�U�7)l��g�]�q�u*t�^�<�	�4e��+G���2*,���A�6:�ϓcB"�Kq꒬!�D���M�l�����I�gJ2ًSJ��-����
�&��E��<�!�=(�5DBÇ9\��R�џ��W	��la�Ŋ]�XSdm�	$h�}��"O�!0N��E*(���L�2_�*W^����
J1IqOQ>�0��Ƅ����֝(^�$�+:D������2z(aCI� |��P��*�I�t���S�? ��!�&�gö� Ö\�JA�Q"O�xT�6̶1��!ޅ���U"O�A5��H�b�Fώ$�VE(r"O��+bn˂C2!D�Ř!�NP{Q"Oİ���L(5(�Y合QO� ��"O�`6��,N��Ew&��@Q�D"O�<���A{?�aA�ņ�r�4\1@"Oh���N�	^`�s��J���T"On��1hVđ�'�rI���3"O� �5�
�-�n�b�GI6���"O�@@(\8/�Di�@�&�j���"Ob飲�@�8p6����1$܁d"O�(��j?�ћ�"���D��"O$4@��V�d����ݣI����w"O�a�(���1�Ѭ,��"O��DJc�tY�KQI2��D"Oj�áC"+e�B�钯f?�P@�"Oؠ�T�вJ���e��-A0,� "OV�2c�@��qT�^���A	w"ON9XC�j�`�IPl��Er�<Zu"O���� �A��,��wE03�"Of�3P�8z��#ۚ\4.��"O�đ��K�nU��PU�<l`���`1!�`���Rb�C8AR���c�(H��y �!�O,��H�O��#P�V�Pei��+�(�r(zs"O����O�2ݸ\���'d��u �	(;h�`��\n�l �|��Pi��ġ��B��ysG�<����: ��ڔ&�-u#P��+\˦�P�Q���f
x���s�h���a���kD�b	>��"Om*��5�VH���!l�}�2¡��1*Q0J�c�S�Q�џ�[ �,E�@�pN
#�����L3�O| KG퉆7�T�BV�z���çB��X��0��D�d����=�`�8�Cݹg⼤��U��4�Dz�i־�r����1���'?݉g J
><"P!�i�9 ���3�"D��)i
4C�-�d�L�1GY���|� lC�n؟El�K1��~���i�hܣU�!��p1��1b	�'*,�CʕGNx I�Ɗ�Q�Ux��O�9p�X�w֔��s����O:Ԣ�� �.�:5U�Yy�|Q��'rE��lQ�4��8g)]�\D����Ϋ$���&�˨3Ҵ����2�Ҭ�E8K��;�	 ݊"=�R�M��V�*�e����D�)���/������'fe�'"O�l��`\�e�0�W�ޘ[���t�i��iҨ�5}��wRs?E�ܴ7�,l�E�p�a�e� |��Ʉ��.T�Z��>��,"`������)���AܩN�$��l��1�6�H�Y�Ĝ��HO�d%Q��Hp���y��dR��I&ɑ���ȥO"�pD��?7-Ȁ
��`����%⑑!�z�"@M' AD�p?Q��
+M<�@q �G���w�  �	:(�H=�2���Tc���=h��ӊ>w̻����	�f���3���4���IMcN�K@�E��4�$_��D����ǒ\���!x��#B�C����&(���'9���O��� ��&ʶ�ZrO�m�`�	� ":,�站�m)���KfRUi��9.%�T.��.L�H��a(�g�Seb���,�o�<��ΐ�=Q�|ԇJ<P���1��2Z2@+m���@IZ#��"��� C4���	��cqy��S�~Ԃ�:���F�1�K��g��$[�+��C��܂��'^�8".R�D�z)�(��!x�m��$�ҏP9��[��Dȑ�[�����y'�'9f޴�s�Z 9���"��0?�ыi�>�{� �������%�.3ܰ��3%jy⊞�d:�q���ߴ\�^!J4푆���y�c[�5��W��X�L|�t�͜ΈO�m(�*Z�xJ5"�����>|�����53��Bc��Aſi��8[�n֑��A�e�F`F{"'�(�R��j7/��MtF��y"!�(a�q����4 �t"���'��E��4ɦ�h�� #Zyai֡R��C�dJ��p?Y@�o�!�����5Fe��A	�5� ���=�ܬj6&�-�~��H,�#�nE�<Q�9���0�g�5G:p�a�ӿsc m�'@6gj��]�n�1�c
1?�y�v�T�<�P*侟��Uσ�%��[�'��Z���i�
A����R\��1*(<ٌ�ڣ-)�@��Ή�aT�]��=q�(�g�? 9*�N�0,,�C��A�0���>ae	��M�,�!��?ٲ�ޯ(Uș�1�� ��t�f�@�M+n��T���~�
���Q7+��۶�.����c��sڰ+V�Z���,�B�E/U��:4�=�O}8�)��D}��Ze�����0i��B�KV���1>��+���1P�)��d5(��(��Y3e���v*�= �}���=jFa|��q~ppĠ�o�qd ؈wy�|w�ȋJb؉�� ���z�/ۇ1���Z���3iD�U��k�?�^8C��1>H#<!��M����φ_�Ҽs� �"���S	<����,Fx-��"F�Q?�����Hb��*��l�dA�k�?c��i���(���2�f��b�j����4��K;0�b�����2ޯl���O]P�:,O@��W�J�K��9��VϏ4yv�E��O�1�� �[�'#k������R��́Uȍ�o��\2����_���kS�.8E\��$��uy��]-;�s![W�ѱ-�k��y���P$ڶ l�'��J��"��?q+a�6d�6 9�iK�-�,�*u�
o� ���)N43Ұ���@PC�(�`�鉅%�Y#��+��'e�X�O��9d�0dĠ(��(`K>q�Ţ,_
)cUJ��U<4���L�8~P-����"v�	Z���(p��ۇ#�-S(���펷�?c���=���0���?)[�y٣��H�'��@S�ў,L���R�ۧ�&�K�-SU}�����O�*\��`ۘtX2�Rף��l����V�ʅON6O�x;��ŕ}Y@e��E6lQ���s^^]�ۓ)��!���K�[�L������Y���BR�%�������Hc呥(j�İ��D��X֤��1f��Y��W�x�&�S�	���I��	�a�`8�47B�pi2m�^	�� �u����+��nj�5$�ZV�6>?��$ŲTjXSgH5C��H&��:zFBEP�@!$,@\`P93����tk��~(c�P�ɖ;kNY�DD@�px@�qb��T�m���h���ŋ2��HkW�p����B�
�X�*'%Ԡt1v�	3��^(d�����V�ұ�t��l��x�EM_4{ Jc�#�,.���#�\�D��i,��a���tQ�#?	'��=*��-ӳJ	�]�L�	F�\��"�?|O�� �;.����lX�|i!ŋ9%LH��A�?I����?��O�5�#�.d�1#e@n�11e�h�&t���3[���f@+��>�!�'C�Y1���	��(2b��a�������<F�‰b�|b��>B��lZ7���0D�4��<��M@#���D���������iyR#+��'P1�+ 	vn]H�o�����k�m�,�q��-!�I{��E�L�f7�����1�A+�)��9��@��+]�,Y��ߔP��T����<�@l��;�RD�W�ƊRF�O��'����&+|cU�=Jh���z���J��':�K�h�6�yլU�"�rJ�/<�ra��~�`Ǵ*�W�Jk �̟���?� �x�(�hq����s�$y1�ɡ0 b��z��Ǐo$��vI��sτXg�t�|��BJ
� y9�LI�q�0��>�|"Ac܋S�ō�22��R3{y�l5��'ڊ���j	9~���O�]�$(�/��d�SL��4���"O( @�+d|p܈sjVv�r�|�b9��v�"����"2�� ,���ˑ|�t�5�F^0��ɲ$<�x���}�F�{��#l����g�ZA�Ð|��h����X�0�**��܄'lJŹb�ĥ�ax�AQ��O
5�t�����
�n
&&"O&� �퀨 �4��5%�����"OB �C��2 f����ҳ#�ν�"O��Q���/^�tA��¨~wεz�"O ��&�GU��0p��  v&0�"Oe�1hG. �� =[G�y�v"O��9Ģ��nQ��ٖhm��"O�\���2 ����!ag�<7"Oΰ`KҎf��I��dB ɷ"O�����1~��#˒`⸣�"O��80��8	Lf �!�]?T(P�jV"O0�:w#��,�����nԂ3By��"O�@E��PsX���-�~p��"OLiy��G�pR�#�1>�5"O@*'�;����h�Q���� "O�$H��Y�dwNyt�{�l}9T"Ox`�睹0ZT�teI�Dʠ���"O�@g��j��P��1�Ѝ�"O\�
##ֹ{����&� ���"O�8i7�P]�����D�>�Ґ�`"O ���f�@�%C���;����1"O��ugǁ+���+k�l�Hd"O�=y�A݋+��`��7}F\��"O�,a�(
T���:��[>|:�¤"O� �u�ł?C�H	cV�'m���"O"��� ���T�03� �{�<-�"O\I�#.Nb����Y	U�&�v"O`�8�M����QB+��L=h�"O�qY`�;<����]4i�*�"O�@(S��H�B��(DJʑb"O�D�f*�2n������*:^D��"Olے�A;X�ՠcG[�=�-�"Ot ���3\��d*�p�e"ObY�b&��<��Zu��1�8�Q�"O��[F
ݣ�Ԁ�C7L��Z�"O����yK
�wgۄJ�X�"O
�ŋ ME������,!"O:�񥅝.f���fb7Wؼ*F"O j�H�Y)��� ��.��4��'"@��$��/� �
��t|hI�	�'�Z���D0c,-yA��yR�A3g�ޱ���	�l)p��'����yR,9)��)F���q��x����y�jN�D���r�� @��]I�'_��yR(u�4�)�kW2wN�����y�'I*��t�r��5Vh�˷����y���y�����F�2n�y��+��yț-,q"�1��]B�C�͜�y®͜Dt�5��ĉ��Hhy����y�ᔚe{t%8B�M�v(��)�-�y�޺8��H!-�]����N]��y2��6i�<,"�G/u�H8�"l��y�8G� �k�"�t)���P �yR�A����J��_vP�P�Ѩ�y�KGm`�fσ(R�X�{P"N-�yRE��'��X1$��FW��(@�y��]�'�*4�����7	N)�yb��[��"� �*hI���=�y��8�`����&Ua�	g�Ψ�yr��Aa8EA�&Ux�{�ʈ��yR��Z�$�"�G��p�1�+���y��Y$&�cԧ،=�I�oV��y��S�"��i���V?Ք�	�g�4�yBߙ{&��x�LR9c6!��k�yBOű�xa3�b��α%U��y�BD���C ħĪ�U��y�N	
7I��ċA�f%���y��Q'"D�E�����9�D� �E�y��6G��@Ї���=S�Ȑ�y¨-Ub��ԭ2���7����y�CK"m�4�S�՘7��D���©�yB�-dX(�1pKI@^��e�C+�y"&�0��X�K�"=�̹�e`���y��&�vT���ǘ5?B%B��N=�y��ϟ���s�U7bl]
�߱�y�ɀb0�t�bU�<�dp`�*��ybm�/Hh���!��4�d��#�y2<���E$�"�髃���yB�/*�J���Ċ_W������y∄�*�TQU"��E��2]pi��'@���L�fG*� I׆z* ��'���h��&� ��|�V!X
�'
L�� �&B�f����H�^)y	�'�ă�샾k_\��7��C�*4
�'"Jԛ0�	>c� +bJ$4�B��'n"�iv�ѩw�8�;� ��WPp���'@��A�<RV� �.I/cFZ��'y�MqV�L0��\#�['b��d��� L�C_�t�v�� �B-IĔi+�"O ��pgҕ�xDS��J�f�x9 �"O��a��Q } �mP$���n����"On�p���g�"�ԥ'"�T��"O4�����3Un���OL��"Oh=ZBC	�[ڤ��%�.��9��"O`2cf�.3@F���s�bi��"O|9{�f�v�&��N��p��!B��'��	4xJ���h�
����C��,{j��� �Tr=����B��#S$�� �� 7n��ȩg�nB�I�?���@��؈q_b!*� OnB�	�4��	���\�d?(A�aÃ{b(C��1" l�b�۰|a���΁�K� C�I�x�R)���rP����a�97�B䉶TafL�fʄ)&в��E���C��*pP��J�0d��p�J��-�B�ɴͦ���L�2wӐ-ZTI�5�dC�I.��c"I
�5��@��;6xB�I!YY�2'�2 ^���7  PB�ɒ!mPr�_Z�~e����18B�I-g.�a�n	
H�07�B�gnC䉬���jEN��	T	�p�:C�	2����T��3��k`�̤��B�ɂ.p���%�E��
pU�b��B��q�~�c���B�����p�B�I�C�p�rp�D�m��=�V�&@�B�10^!�� G�t��
E�v
jB�I�MxU����0�!�6k\�tV�B��!s
r�y��A�Z\�Ȅ��k��C�	�P"Xad/o�Ӷ�B�[�C䉦b�!�"�'Q�@ ��_(�C�OԐX����-8�9pd���C䉀(��!aV!e��6��0:��͆�!K�4Q���-���+t^d���|�&\��lح	R���m)�8�ȓa�����ג^:��0�	D�l���ȓ[����,����Km98�ȓW@����3j����$_7����'��}��A%=j�qc��`����<�y�Đ�58rq�F�яP��E�&J����'��{�aN?t��[7Y�ED.�v��;�HO���d�%i�lS"꟧���C�@�!��@dx���h���K�iٌ{	!�$~���˖�ɝ0�:@�0"�w�!�d�F���C�m�Ä G�z!�ֵDL��N��uflT���X�6}!�Ė�V���Zcł.c�ҔHgf�5|!�L H̵���q��Ps뎆F!��'T�6d��Կ=lJ!�ÃW/x�!��R�)����W�G�2�@Xش��2#!��2Y.p$�e�Y+f��b�I4V1!���-a�4h��I7��i���-�!��Z�����a?D�����[�!�dPpH� � ��Y[z���O.a�!��U5Pj �r�J {���5Hm!���<9��L��n�[Q��"�!�_�kq�ث�&���8�	2�LM!�
a/R�����)��!���;&0��DJ�}��		6
�N��L�2��'d,B�I�&��.��pg~�����b�!�ę�jt��p#BB�*h�Tƕk�!򄍩22�J��,�F9{��K *;!�d��F����g�N/�n1�N#)!�� d���I�tD��l�{�N���"O�q����]��e�:	�@٪3"O�M�T-��"=�-jD^���1�"O���O�G��١L�G���t"O�"N4OӼ[���O���'IF���$Q����fK�B�݆�y"��:n,�#��F�$QyՊ���y�H[� uRx���B�@ɤ
]�ya�~��3cd��"�\䋤�O�y��ƻIKJ���ꕒ�5(����y� �dd�(�%�<,�~e+s�
�yB�Q=X����,��5�&0��B��y2*\)2���K����k1�Q��y"-��V�� �LH<�x�+����y��-���OG�e����D.�(O��=�OZB�EӄAE�DZSi��-��p��'S�Ar� �ZᎬ���]�}�&���'���
�n�)mx���A
�_�Z���'���sF78�T�W�[�Xw��R�'����M�Q�v��5	_�NS
�
�'��-(�`��KHXR�d��7N!�	�'���c�lU7��7�H��'Ĩ�$�&��͑W!P�c��%B�'2d��"�O����h��X��Y�'��8� �'��Q3&O��4;���yr�G�隠���U���I �yrI�W_��C��Fh|�U��yR��� 2�����3@�l�F�_��y�ŗ�S������F9:j���h�y�N�0i��=*�D�d��PR4c��y�$ٌ\j�:�U	_����@D��y�o�H�D�Z��ޮ[�6 sĪ��y��23"�Q�Ц��h-�,�Ӏ�%�yR�J� �r��Q�P�2��P����y�U�|�H���">�@-�W�M?�y�jR6~<u�F�L�:�adc��y��$x�ЈPvQ�)�+�3�yr�ߞ^��@R^2�׋�(�C�	52 |B���,~V�e2�Ĉ�q�C�:ٖ��wɪ5ʼ1���
�C�	&TZ��"Ť�'"��|IŇ��+3NB�)�j�a�ț�w�hP3�-Y�b`C��+>&D�P%8�����2Y�zC��M#�a�H��5q:��d�a|B�"~��U�����> :��+�B�ɝ4�� J�����'��[�bC�I�?�Ġp��yv��t���
.~C�	�*%jp�������y�M�-C�	2|���hB�� y���!)W_T�C�I�4��9�&�(uc�\�#(�;+�C�	�2��<c6jW8K��BBI�m�C䉫���Bw�N{㤽B�eַM��B�I
z �Bb��="φ�"���/,B�ɀw�~XhD��9����B��a B��"c<4���0¸H*cL7IFB䉥L�]�v�ɫ ?������./��گc0�jS΄�H���&�!�D������E�,-D�<�%Q65!�$�� |=H�	?Ӯ���^;- !�`Djm�D�ӸW�b� �ˊw�!򤒘!$
���b����Ң�,2!���@�����&�����6�-A#!��.Kv����ߘO���W�X(5!�D��8�j��ߖ���#cV�E!��  -�@e}�P�2��:�"OбðiY"?��x�錌(��s"OpX6)�CA�5!b��$�d�� "O`e�η/�~ɫ�(�1L�<pS�"O��#��� je���ME�H����"OreĞmz-钆Z1bX8""Of��%'&�=�bh�	j
T�*�"O%��i���%"U�"H
b��1"O����aO��Hi�,�r�3t"O��b�Z,p��x�FNS�n�R���"O,}BP�!@;<�P��Ms<���"ODppc��.��A\�7K��9�"O�m�R@n`�R��֒��#"O>i���ҥ�Ъ��v�Tk3"OD�ir)LF�P�(�3�(|Zt"O�`(�N�.�z�H�*F�D��`"O|�#k�6���`q��-F�<��"O&�J�DR�E��J1[�6TD"O�pC�H�S�lAh���d$�&"O�9cCFF<�� ����6DY�`"OJ�*��$	@@mxEᛧ �	�"Ot��"뉔pj�+�M_0"dA{R"O��q���%
���̛>Y��{�"O��aQGս0Ji��F�=�@<�2"ODй���B���ɰY�,�V"O��y�L��8�`:�f�Z`.��W"O�������)e\�ɂA�D`��b"O�0�tiFs��hXb�-bGX�C�"O|0iAEYNbv,��Q�7'��d"O,1��h�rMiqH[�n!@�CP"O80��X�obL��Թbi<$s"OTy*�'�$~�a��"�\`�7"ON��%B̦<8��I���2"����"O<0�F偵M���`%*s���E"O�	�蚪}6¥:�V�,>��"O�8Q�����8[��Cdx�"OH�f�V�Y%n�@���0P����"O��Z2�D�z��,
/8
T��"OR}��k�	l|�ܰ�*W�r�ձD"OT��-�?!9 ��٭t���"O~��7�9Aδ	�-_�ˆ8�g"Ob�hfAFEP��,��B�Y�"O�� F3�TQ n��<����A"O\L��J�cւ�qL�O,D�j`"O��P�Ŏ�J�N�,�&*�`���"OB�ק]&������`��䒣"OhY1a�y���"���mQ�)�G"O���GN�,;`��2E�f�`"O|��FC��)�*I.��Za"O:�V&7bn��vn��~����"O�aa��'t�n��TL��h�@"O|�9��??2h�'�΂ɨ�"O"L��B�
�P����qA"O���#b[66�.��m�
_�$�@q"O�9A0��h쌹p�P������"Op�2�T:|>����K��d�HI+�"O�����@*.���s͆?r@��"Ov�C%�R�)���3�*ud0��"O�`�$j��G�Fa��i�((�l� $"O�)!�I�N�������w�7"O�m�ʏ.�v�a��H/7c����"Ox�腢�"1�4(f�"X|�Q"O�-[fF�;uԄ`qD�� aG"O���G�L�=�"DQ0/Ӫa�g"O� @8��B��TP��¡Յ\���k�"O���q�K1��I��KS;f� �	�"O&����Z�l2M�6I��YB0J�"O�m��o��H��V�aQ�i��"O�̘�a� vw,(��ܫR����"OPQ�)�>`�+�&�#h�`�4"O|��"�8O������G�l�T���"O,����8*zf;	0LPi�"OQqQɆ4	���1�H�Mu�P��"O�$���5�zD�T.��lX6��e"OP}�E�*\I|t�-)4JJK�"O4]P��<m��aɶ�
�����*OƁI4=,��!��33�l�:�'~�qhF��2������t&�da�'F�� �!S+[�41-Ȧ���	�'s���͇~�@�Qch��+�'�H�$Q�)4%��E���H�'B��xAжU�Ь��E�(����'�����#�#3{����u�����'�0���HPBt{�����|a�'���h�!ÊUf��'ĞI�t��' �mZ��Wm�,r4I�*Kf���'gN�x����*�B!n��Z�z�;	�'�V��g��J�Z�1VBڑf՞��'ր�TC�x
 �cU�4ք��'��S4�ܙ�x�)��2�ݳ�'9�I�`.X�u��M�Ee�r�'�0E�5nͽf/F���H��h��X��'�H�Ҳ.�4N����/J�L\q�'l�}�ᦉ/�dL8x�ڨ�'���� j<
����Ď��@
�'��\H�d	182�GgX,S���"�',Щ�Eɘ1|�@7k�H�L��'�T� A닜I
^��̢s*n���':&�ga^=0��|kW��9�xA2�'�<! ̪-l�-{)ޯ&��� �'����Q,�.��X���D�jv�b
�' �p��fX̘��ć��T1��'3&!�F��$>�&L"v��[Ҡy�'�6�����}�h̩�5'Y����'r�G��@͜�
5��J��h �'X��I�H["AbN�I�͚6{$X��'���0cס8g�0�UL]�|����'5~�r@��,��Pui�?�� ��'NŠ���>:1 ��M�Y�|�;�'׺�����<!�psT�ќW�f,�'����"�׼~r�9XԬKTzr���'�|K�
Q���SCB�G�h��	�'&�E#5�Z> >�`�J2n���Z�'o��T+؄���Y�o��m>	��'(���H�`�0��-��8c�A�
�'���2"NY�y����O�17<U��'��17BP&'\<�y��5�h���'"�i�1ni�T��k�='�l��5D�xd`y-j�P���Қe�>D� �@4Kj�|8$�)	cr�b�=D�${�NqL�Ժ`��(r�J��wM:D�|it�,�����%��x;�k9D���w�Z������E�p���5D��6F�#Ya�0�ʬ�����4D���DF��2�-`�l�=l��P2D�H�6'�){��x	A���5�f���n,D�T�UAE�i��!àX/nPda!L'D��!lH�\|FUP�	tX��q"*D�� a��gX�xB����ʦ\��{6"O�HB��+i�����]3���"OV����A��5X�Ǉp����"O�4I�&�5�v8P�֊ܖq{�"O�,���_�3K �����O���"O�0���P�u�Jyb���L<�� "O
��b���g�d̸2A
 �lxi"OP�<.��P�"\&@��l��"O8dXA�S~!f�z�^	-Aā �"O�\!���t<�e��9���"O,L`�yD�h���=`��D"OL�r׫O�w��F��4�p���yr��-�j��RA�r�b�	���yB�͉О��"�<�F��P�=�yI�#�^1�v�$���!����y��I��}B.����4�P9��=a�y�C�<{��G�9�����	�?�
�'���Kq�˂��.ę7�1��'�&|���H_d
dBg��u`n��'%4�瓷BM$�pՀU�q�
Qq�'���O��Xd+P�	;����	�'�ƌ3u��=^zVq����5J �	�'S������r�Tkv�܎:.�@�	��')�I�6EU�0и��զ�4��i	�'=x�
��ʚ@��%�ĥŲ=+<=��'�P�H�k��I$R��+��'��� m�(-�M�s((ʒ�
�'{ ����Jd`mۦ-Vڔ[
�'{p3���?&�Ѧn��;Z��'�f��2�-�aVEĩk0����8?�6B9N.) ��-U�P3DC�x�<1�JRR������*ʔSD�Gt�<���1..�攪=*͚#fXl���0=i�FS��Ő 
C#bLѠl]�<!%m͒0؜�qG���H��&��<�U5u�V��'�W�3��,+0cC�<�񠅙A$1yt��*����2�^B�<�"�F�9��$���H�=K!y�B��+)��b��[�B�����gH \94B�ɫE�[���=��T{㏊0l���?�<�tL	e��J���F��ȓ�t����
s匝���ӒQ�>!�ȓ<(t� ùJ������7"؅�,+����'x<Aj��E�m��IR�'z@�PG`V'L��T����LpB
�'f�XB�ln���`���5<@���'�@*�aп<0R`�0�8�����'�j��[S8|S�l�2�� ��'��|�u�M++Xǡ,)��
�''j�H�抯3t⬢��W�P2}��'*�3B���kV�I4rN>�L>���)H �J`�Ć��~���+�!�ď�T�Fy�i��D��,�R�I�M�!򄈃F����V<m����:�!�
3�<��DN;T�<y�#��+�!���ڬ���@�$F���u�4`�!�D�V,Ҷ(${��9�ӽ0�!�D�[�B�)RL.A��S�l�X�!�D@0�@3w V.	44`�Yw�!�dT���UЊS�����B�2W��$�"~P*�Sh���JU/�ĕ���� �y��ŋHO�tkç��,A)��O	��y�ɷ�����`ƻ(I M{")C �y���mB�37�Z�id`���։�y
� xd�ց[�|�wk��cf"Oe!�"K�m@�9��РRQ*dqQ"O��U(ּ�go�}3� �%V���	f�S�O1��QhʩM�&�cG�E�)����	�'̝b�N�.��8w-�
L}"i�	�'�|!	��~9x��$S	�'�L�z�+Q0���2������W��y�.�9ȩ(�jF�#r�M�GMQ��yBM��}��Q�(����s�/^!�yRd� ���S刻g��`���:���hOq����q�ja����"E#4�axc"O&��D@=ɸ�K�ᔟp��A"O��A!Hٕ>�)K�K�#���X"O�y�s M�;��� ��E�F���A%"O��k�O�*S��8q���O�ƭ��'��8���)(��ԁ'��Q�4Y�zC�IM��B��+i��R�)��f�F�O���ɸ��yya�+'2���"�>j!��>���h�]�p�D!��yJ!�DXh��7Fʭ���W
�!?+!�d\���p��J�F^���	��`!�C/^B��t��? >��T�_�q!��~�Z��Ƨ`��䲦�ih��y��R�r�ޔ��C�y&��s�*K����(�OL\ �F�r���.�'(C1��"O���2U66 �"&�$���"O��qF�&R���`QA�`����Q"O�]s�"��=��[dj�c���f"O>A��BqI�Vʆ�Pr4"O�q��;L)Q���3^��C"O���@�#c���F�ԗxh��R"O��+�Ǒ+kМ�%^�N\�HҀ"O�!00H�at�[���3PY����"O�-p��T�{�܁(ԍ\�]���"OT�R�)z\�|����4���Q"O&��W�ɬ5��|�r�"���"O�qp�i�U< �#G�C�L��5"O���!�
#�jQx���<N��Hi��d3LO�H[�cYh��
��['7����p"O=����*e�ݺC��i��  "Oҽ�����g��`�D	�t�D�E"O��2%@�H�q�sH�2�*@�F"O����()���2��'&x� �"O�����nπ-t�Yc���>�yb܃����ԥT9sWߺ�y��W ���b�ʕG����'�ۙ�y��>�ZT`D��(���H0���y��k�)Rj\�S唽1f��y�A8B��� �ѧTm�4{���yf
4��BǑI%H9�b@��y��cm�@ F��H�����3�yҤ
'��9!������B����yB#�"~��@���^�'0�Jvĝ����"�O�HQ$�*-'���f��
P�nMc"O|a�'F�,WGV�z�b�=Ĕ��"OF����Q?Wt�*� �^*�;E"O�1�W�h-�Ay��g��P!A"O~�
���?g���4������"O�t�pJ3b�$-���®;�0���"O��C��2Ud!zeɇ�C�P8�"O(�ca�n�[閒#��x&"OJ娀".D�fd��Cqbe��"O|	������*����ePQ"O����[��8�A����\��G{��� ,��"Ue1�p!�]�O;�8��"O^�:Aj��r��r冝�
*Qj�"O�
�%�K����O`�Ȼ0"O�;T�T�m�D��5o�2!�zк�"O�����f�Z��bN
�4X�s#"O���F�;"�J�[`�ߞ[rj� "O�uh�Ղ]%$�Jt��4�bM���'�R��'�Hm(��)�F��p��9�b��ȓ,8�u���ƺaѮ�f�3�J��l*Yʖ�1
����lӚ}��Y�ȓf�hز�GJ>U.��&���ȓg�A{�ʛ�I�8�o�VxI�ȓ{�H�I�;T�^�ˀ��r&�,����ջS��wώ�VIF/9&��r������9�L�5�<�!i��x�v� e� D�x���՝ƭH�c�-RNfeX�%�<A���zBKM�=xR5R6�Îb\���o���j`�T�$�:tn�̊��}��;��:�������kH`����>��Qpr�	\J,��,�9-xν�ȓ;�(Ԓ�	�$t��%U2E`��ȓ�(��qa\#G�a��F
fQ�T�ȓ!���&ŚM#�xBu�ܿ^�$�ȓ��=p�S? b�`2��9AxY�ȓ-.BhCR��=㖵��X5X��ȓJt�K��Хad�1zSjЄ�Z�$[�`U�f�L����.-L옄ȓ]7�����$q.^�a3ᑤD%���37����m�	Yf5�d#�!#��ȓ
y���`ŋ�7Pv��ե�\6*���}�j�(0	P�� �G�5�t��~�)��� �k��Ԓ��;�H}�ȓv����ف1$j����k���� Z�L�5�*w��%:���3"X���Sb0���7� ��I%-�r�Dr�ӻb����l�?X����@��|VB�I (N��U&���ikG�0�C�	�Z��r�3���R�Ȥ}��C�I)5=x;e �b�f�3#�)}�bB��o�8�Ю��00���M@B䉵$s���PgB��F�o��'�B�I�d�ȡS�A�'g��%An¢=i������!ӧ��v���x��bd� �"OfH�2->#*2�a$��+�%#C��y2���e�6���HA$쐑�yR	�cD,�Kَ|���w�.�y�hӤ~p����0o󲨺fM���y��H-�-0W�ȪnM�LN��yr� �b�8���-�=M��ұ �������hO��Z�+)pP`�f�׿N` %�s0D���ǉ�2Dh �P�	v^��g�<و�哼[�@Ly#���g���[ !U�p�TC�	�_�4� ���6��<|4BC䉚7m��̟�e,j\%ҍ�vC� RZ`C	�G6���ʄ9ϢB�Ƀ'���rŅ�`m�D�Di2�$��?����ğ7Zҡ�L�o�hD��Q�!�U$�T�5�Ǖ2J��BЅ <��I����	[�)�'b�vL���&��0�G�ˏ�5��b}(UBA�<U鈙J'�
�����*�H�	�S�N�c����ԍ�ȓ?��Ā��A�E �P����0N����DTj�qr$�/a���ۅ�U���p�'����wf塣�\�_��@��(8]|C�)� P�PG�DW�1��)��1b5���'\ў"~�^�4}���%@<>E�D�
��y�/�r�<Yt@�(��)���#�y��8��bE�0���Xf���y��K�O�`�A�q�D���y�Ï�$O��s!⍎t2V�х�
�y�#Μ`D�8 ���oj�A�c*Н�y�?eC�C�C�d�L���ϐ5��D5�S�O�\�"u�\'��9�U
؆�r���'�N�+���<���(��N�#n���':�#�ɰY��L�����
�'��I�2d�,c��,>n&�q�'M�U�ǣԈ$.�De�N�9�aK�'$���!�V�
���Һ���'��pϘ=&P�����F�kZ� �'Ԭ�ie�Z<�z�X��k�f��'%�`r�1!?5P�� �Z�����'q�R(Z ��҄o��<lj�{�'���ITD63 ���Ԥ�+��i�'�Z�x>��!�����([�'�x Y�@_�[��;�A��^�h��'�6H�PЎ���Cq+D8i�`���'\��9AEʄCa�tp��P�6N� ��'m������c���cA��_�y�'0Z	p5�H�l�H�{`O<%��yH�'w\JPO��3��A����!V|��'֔�C`�Ė5��B�Û a�!;�'�����e��C�J\ID��%��UЌ�>O��X�
��_���s���&3��8�"O���"'C�Q� ���@�6Q� ��~��P�s��܊}��ΐ
�<9��^1�iM�}���
��X�e�8�ȓ(��CMG=`���zd�>Qۀp��"�2p��hr���R�M� |�ȓZ�4�مŉQ(PYr�IԸ�ꝗ'p�	b�)�Oz-�#�E!}�D�3��I�� "O-��P�ak�8���K�i��a�g"O��ٔ)�o�F���K��jA�"O��ঋ
6�����\��T�D"O�(�0d �c!�<y +�6D�
��b"O�H��� ]��L���qpX��"O8�&�ŧ�b��w6�x��|�]��G��'[~�0f#�!`� J��R�#�p��'p$�z�e�%�b�cqV=-�N���'Z �yB@�)68 t�`h3y#�-��'0�u��@G�}�H�_����'�2pXU�Ii���Na2��'|�<(b��
p�:���G�L���'�
� $���<qr��,V�Tx*O��=E�D"��d��)qf�6��l����2�y��VM���%aU�3����ӟ�yB�T��v�G81��l J��y2Μ�
A\$ۥ'ӟ=���T�ܦ�yRE�Poj����I�t� ����ڵ�y� �Xx�Q $�lk��(a�͵�y�b.W����N�dH`�(M��?я��v��<8D)��U���d<=�*���,y�R˛�Ⱥp�M�\�܅ȓHi��iٙ���ʁ�I0��y�$%��>R|��D��E��I�ȓ1-`�b0o�|��!CF\�;��Ѕ����F/�+��s�[Hw	��8�L��"R�J�e�W&��j�a��8n
�CQ��1fD��b��4��'tr��3� �A;pm��>�6`d�T�	�"O�˱O]�b���[ր�4hK>���"O��jƬ�CJzāe��GW\;�"OZxpFB�i�H!�3dE�H����"O2$�nճP�����Zv@��"ONY�P�ήTQÓ�� Q�
h�"O��w��1n�2�! ���́�C_��F{��ɚ��4��띟I��aD�G
m�!�Iz�D��+	\���+���'d�!�DP�9�k����.�4�p���N�!��}D� 0�ׯ26\�`j��!��228��+F�P'��x��hY��!��ў<:��   5d�W"�(�!�� p�T#TDO-u��e�1Z���'b�O�#>�&�
�F�.�i"�ī`\{�l�S�<�*1}.�"4� ��I3� �K�<���w0᱅�ei>�2T	�M�<�GC�)�p��G'�0�:ơ�N�<	5����� Ȁ��8sF�D���F�<� DF�,9R*玌�)uH�rƥi�<��� �E�����B� �AP#��hx���'��A��*K�X0h �${T�m��'�0�	�ÿiY��"/���b�2D��JU,O+:HT9����W��A��%0D�J0.Ƌ5v�(����fe�Q���+D�Y�ҍFM4��"E�Y]|i�l*D�h��M!&�HC��N<��Y��#D�L+6(מU��I�FF��jR$!�D(���'(��b�ݥ�H5 3��+����'��eɤ.�!���[��9(��'l8���晍`}���&	�Ԝ�'$��se[�0H�uCQ�(��ڷ�y��?M�JW$���`xG����yR��=T��L	s�#���W A&��'�az�ă16��*��9F�b�Ai���GxR��??�t��D�\�f�&�J6�P"�y��ŻGK
T�A�#X|�-딎L5�y2�Nk"�,X0Y#X���c�� �yr�M� ��][Ą�]	�d�夀��y2߾a5�ȁv���MP� �F��<��?ٚ'[�ٛ��)�lez�@��^�����=��y�ذ5&�t("` �7�hURfI�7�hO����A�'+�8����-J�Ti�-%B6!�D��
9$%�^@�Xr��Y�G!�$��b��%.�N1����(ڦ !�D©=^�E����@�xT��?f�!�$�F�B"��A� �'$��}R��81"�>�I��܅/�.���9��b�����>O�i6M�!oyY�7�Ո�R�.9��q��M-z���������y""��R�u�GҸ
(��	Y�y���`���۴Ag8�sM�(�y$�0$T�@\6O\�ˁeΫ�y�Ό5P�v���/���c��y�nM�3����P` � UF���yR�L�JҤy�ѩ.�MS�g �y��3-
 i1��#d�c��_����hOq���Sw����,�q���s�H��0"O
�!W!�1?A��,Ð}v���"O>|��Ѿf<q��KO�mv4-�P"O��#�׾Mt9�W
�yV��"O�m0$h�.�Hd�ÃA�W��`���'n1O�q���1	��B��Yr���"O6(+q&�Nt�kglF���T"O� $�Q`d�&F�S��]*��i%"O��cO�a�&��4%��d�*H��"O,������̨�3�Θ_�LX0�"O����H)T�H��a�+6���"O���$��:TM����F�ZE��"O�� PȖ�z��$ӈ^M8S"OJ��R���&�2�ȡ��v^�Ѻ�"Ol|���rl<;�.60E�I��"O�|Y�
�$&�Dq�fK�A��b�"ORa�t	@??�u�w%�0s>��"O@  ��E�nL�C�`3���1"O�p�n�?A��|��$�|H�"O��"��R�f-3s���I`�i@"O�`�%N����1vaJ�{F"O���#ūr��+P�\�`�`e�v"O�d�*�P[�m;QnB\b<��"O*1z3OB<e|[M�d{����"O6��b�/r76���,��C�0�;B�'��d��PK������/Uְʃ :?��}"����"�+@������%L \ٱ$"D��Qd���u��`M�f�=��g"D��y��D-�i���Rf��w 3D���)ٖ%T���!�H�>��K�!<D����'�Ȣ�Є��1"�?D�hx��H��0"ޣS%����>ړ�?����?1��$�κ,g"�HR��"B���:� ���y��)�,�c�L�kIr��c5�y�������H��_WF!�@�N5�yҍ\�Nm�ݚǡ��R|@���`ˎ�y��ׇ<6��
�C	`ؖ�� ���yB,ƻ={j�2šF�(Na����#�y��X�X!&�A&�86H���O\���O��`�U(�djH2c�nC�7"O�0F+M�N����N�b���;�"Orᛐ�\3�lyJ��G.���D"O��b1�W:V��B���?5��t�"O�P��E��U��&� t�"OP8j��#|ZL �A��6?h�pQ"OBu�ĪF����;Q拠0���y�A?&F� JA8.�6$���Ѝ�y���zdR�G8"���cܦ�ybCNN�!����� @�B��� �y��@1� �	��`�\�-��yn�,f��4�V�FQ>��E��yb��2��4�!��E�$xJ�y�@�4D��}0��@�T��x�Ȍ��y�̞xoм�֪O,C\yS#��y�F��s�^�[E�עQ�<��r,:�yҧ��G��QWIȄ3��e���yrҨE�I��?[�ZpYbdI��y)U�E�A�@AEvx�ΐ��y���6����E�7�&�1����y�H�5U�N�x�k�=������y��S�g%�,�� ��z����'G�y�/�'N�����Ԭ~H�4I�i���y�+u��%���ڻ��{�ŉ<�y�d�+�,m*Y�n�tq�um��y�M�ɲ��J�^Jt�УE��yb�0�J�k�]*���t"�;�y���0e�l��#D� ]h���=�y�!T���qS�$X�@`0p�(֏�y��+�< �2��9�!��4�y�mާv��U�#��wV�@�& I>�y�	+1�B�˃�ȓ#*jѩ�ʱ�y
� :��ܗ�r��Ԣ���Q��"O���	�8'0��k�K��`�Qf"O��ڶcF�ތ�H�!"Q���Q"Oะ���%�����N9�Дi"OzLA0�NA\<l��#C$/{��A"Od�ґ�&��ب`��2+�^)C�"O�H�E$�#7_��c���8m�B�"O��!�ݘx�Vj7�T,��x�"Ot�)�i^�W�`[��W��k�"Oɨ (�t��<���%���"Ob8���&Q���0-�����wY����	G���$B�	v|ZP�W�?�B�I�k�B�b�gӾ��Ļ��6l~�B�(�*�hW"8�*	
�f�:��B��0\� �Qa�K���s��x|(C��(!��"A�C�`��b����g>D���u�_:^k �n��q��Qe�1D�ɒ$�(�C �Ɔ*!��E�"D�Xa�Mg�,ɵfZ������?D��
�fM!���@&)](��9�p�!��õpL�C�-A�\�G�<tC!򄍯I��l��Ē�=��e�3�P�!���-��5�B
M
���8��7�!��6<�܋e*�#L��p/05�!�D��F�(2�bU;:�t�A1�W!S!��Ӛ+�8��Q�9�:"�Vj�!򤉁 /|����발�⁞�nr!�d��n��P�j�i���!c
\�!��L�IO�����D��"~!�T�x;�-�8�l��5�3�!�$�=7D�E����!3��i�5Jg!�-� @Nԋm�V���C5F!�
v1�r�U������aI�J7!��IX�����*��a� ��!�<_�t�c휬H�A�!�*+�!�䊧z������Mn�Hz�BQ[�!���)��M����Bk2$´�S5�!��&f=�p0%�Zx�#��'h��'��>��ᦔ�L�0Rڰ4b�K�"C�ɵG��@xs��=w��,j$�XN�&B��#!����*ҫ-�(�[�.ۏ]�HC䉖 ���0V%�<*��! �
�C��7V���e䒹By�{��j��B䉺��TЃG�gNj�����w�C�	�1mp�Z'�<-�)�蓔}<��Ot�=I�y���}�茱�N�}���ˀ0�y�M6B�h2��y���rA���y��'i4��td�0s5Fipـ!���O�4��얥 �R�y��F�x!�DԵh����#� e�:���΁,V!�ޑS~��K �ݥQ��\`�Kѕ6�!�ć;l�>���,��0��)ȟL��'wa|R
ӜJ��1���FJ��(���y�KI�[� 9�,�0?� �C��yR�]'p��Tꓴ+�~��훣�y(�"��e�<7��E�¢L,�y�%�_π�ĩ>]��B�ޙ�y2 |xZ��L�OC,Ē��F�yR@F�Q��w%�K�t1dL־�y�%?`�Ӗ"IR�<P�����y�%�rG��a,�F�
��
)�y�Jv{�,A��K12��J�%Ŋ�yRj�l̲*�˞%3Zii����y��*5�UR�L/���6��	�y
� �8��B�`Tx����Pڱ"O���%��͢%�\���@5"O4����D,��1횄lҦ��4"O �Z�n�X��q�� �x(� "O���&D3�l�Ђh��8�Ұq"O�����'4�b�_=&�����"O9��	�%B���9��\}�t��"OlhP��Īx=L���ĄEg�`x�"O�8�t�QB��CUc˲R�����"O̹���;���c�K�3Pz�% �'i��'�0:�D>r���A�؝��'�^p� �% �$�Q�;qe��'����W��1!7�yX$ЋQ��)�	�'�*)�*�(hgd�b��;RU����'2Tr!灶i�����ڏQ�y��'hX�i�D]�y؝86�Y�H/:`��'�0ḫ;�v�(F��P)�����)�Ot�y��[���N�=b�HKd"O
5a^�c-ݢ�
G�hG�[�"ON��C�[�gj1�*�MN���C�	z>	2���p.��뇂S�o^�CJ,D�P�JQ�y�beA$)Q�<�`H�TD%D��#\d]�Eh�K�0Ȏ�0PA#D���Q�ˡⰍR�Z�&�(�p-�O��d*�O�d� 
 G(h@���d��"O"};-a,���Z(U�L3�"O��F��7��rv��>g=�=��"Or�����	U���C+MOF�p��"O�1�B���$�	�\<�9��"OJ��T��V�Xh� ��	#���0"O�� A��Op6�Q�J�6a��"O��� /�!	��I���NǔYK�"O�	
a�˵5��Y�L+MLb9B�"OX��W ϲ.'v!4NXB�pѓ|��)�m)�]��hX�8��1"��_zpB�I;DA����gG!��[DE�.N4B�	=�^�YQ��'"x���D J��C�ɆP}�D[�.��;� )�@M��C�I$P�Fu�B��/{p��tjL n~�C�	>jy�Ç�+R�icgH�(�@C�	||H�q�R<8�0�#|B�2n�<�� ��q����!gLvB�I|]4������3����e �4)pB�I7N�����R��@ ��_$E�C��3��K��M�	Vʘ���[52�C�	<H$ЁN��)" ��&��N��B�I�M�M1���O����4`0`zC�I�~� �a�J��TՌ��e�dU�B�I�%:��#j�IfL%���^��C�t��49�M�*��}��S�ywjC�	�0�2�����;��yHb��p�B�	1�4�L��w��K�n
#$,�B�I�s.����d�1��a�G�8`��B�I�b隂j1�U�&@�
o��C��l��MP��V�0��%��F*�=�ç7=� xa)´&�!�ae���,�ȓC���g�]E�Ա���6;�Ň�Ht�C��8
 �mS��o�.��ȓ,ްb�	|��K�f�d�ȓ���W� ����{5b<`�̅ȓ �y�
J2Z�";�i>G�\��n��Tq!��I�V�ʣ-����v�����\xь��|2T1`'Y�o�<\�ǅ+D�t���۾A��i+'�B�&�X��t�&D�� b\�fK�E~�80��>\����"O���E��D�d�
WƷ>�.%�"O����E=r�� Eض
}]p%"O(̳Ƭ�I&D�)�.؀uIɚ�"O ���7[��`�k	b��yP�"O&Aa��S",(�2�I�
t+�Z�<�sϝ�Q6�I]|��G��X�<yvI�$Yjdp2��vT��-Y��B�	R)qKƂ�|5��yRm��0���D�ID>���R�BTC���<H6����&D��8�g��k����&ηoW���`#D����Q�0�","�/�	$�*A��?D���Vi̸8t�u�^:@��L��K>D�T���[�*��t͚���t �	7D��`3(�)B`��z���7Gh��k�)D���s��0F�m�m�|��%�'��埄��S�W���hI6ob�E�'+ח)pjB�I��¡H\�B�������b�C����i�ǭ��d3B�R�s�C�I')��EF��RE�,`�f�+i/�C��/e���fX�`m��g+ѕfw�B�I)~B�� ���yybǙb�B�	�6q���G�l���QH\a�d�=qçoܚ6E��
w�%*V����"D��R�d��``f���
-s�� ��;D��W-�"?v�h��jD�#��p���;D�<��E�	v��<�Q��.ct����-D��`�3����߆7L��2�L*D��Á���f���(ț<n�Kd,>D�����Ԟh34� ����P�X�(s�.D��X���<ˊ ��&�&:�4����!D������Cq�F�B�AL�AO!D�� �b͔'~ޕCV�B���x4!D�$b�j��I��!hVʃ5���1�M2D���vVUЄ�3���`��sQ,1D���Z�qF�=�pd��6x�hpM.D� ��-O-p��)0��Yt��L-D��2�7Eh�J��U��ku�+D�x���^9r��Ӏ׻'���@o(D�0�-�tG0*�#U&?&8��g$(D��"@l^��B��������E%D�t�#,]�K�<�*���K0�Ax��>D�He]�M�n � I�?�� q+!D���ţO'i���1qI�c�z�R6�2D�8zi�0JiB|V�̺2�v����1D�t#d�O�F)�z`_=���N=D��Y�0f�N�V����lȊ�a<D���Ԧ�$єؘ�!�a�:�!�:D�L��OަQ�[\<4�1pE9D�����']բL���]*K����  5D�*�*�b�Ͱ�ϛ;�va0��3D��نɏ�"P�e,H�C\	P0�<D�D�Aj+�J��ѭ�.c�e17O9D����k��:�lR���h1�gK6D�L mг+l��p�98nJ���H)D�H�'ڐdd���A����6 5D��Z�dC�3�u3@�gnB��v�&D�|j��Q,&uv9rQ�ÆYV��S�>D�0��DC	��<���N�a.�m{�n8D�����Ӄ+��슶G�x v�3D������p�>8���Ȑ5;`Qqm3D�4�2l�'���S�	$7$�)��#D�����q`A�l�~*�ׯ&D�� r�	/�y�6�@�p:�}��$D�� �p�ܢg7� 3;p*�J�"O����"��]"#��a�v�"O
���	L���AP�U�H�,ɓ""O�\��G�!f�jH u$�K�l ��"OhPrԠ�.i�d���G�Գ&"OA�AA�:6Z�SǨ�?��s�"Or���Ռ�&���I�>��=(A"O��
%D�;&��8���Z��"Oܥ!��<�| NŮ�$m�"O�ȁ!�J�U�^M��,O";p*���*O���l�&Dѵ*�-6��|#�'BT9��@}�ݱ 2 �J��	�'�`@�����	�w�L�g��r
�'�zq��`� ]�����3c,��	�'�1k�K�7e�����v%��'m���6��{��P \3��Cr"O����Ma�H�T��~
 K�"O�t��b����e�ve���4��"O~�yக�S�����2](�`"O8}p���� �!�9X�H-�""O2|��m7Ј��3*Q3sĄxu"OT� ��"*���	���#d��A"Of5W�Р!bj���L<Ai�x��"O��Z���g�b6�S�z���"O,��!���J,�o��yaq"OfSK�q�������/fq.P�"O��jC%�(-�EZ2�C�9����b"O(,��!	5b�<�0�䑇R�D�!U"O�upekY� 5z�`A�X+\��(��"O&造��7�V��E��b�h�#P"O�EpB*\���`)�
Z�`v"O
�2��pҔ�G�0` &"O&MrP��YG89ҏS�Mp�|�1"OV�QW&_>1�d�q�.�l����d"O��쏩,���
�/��4<Ru"O��*#%��%�"���z�"O���6(��~v@��[�����"O�Q���n���)1C��S&NAk�M,D�����A3:,h�{FO�~M�2@7D�l@�#��)���j��$6��K9D�ܸ�S��ɠb ��)����B6D��0�&^kC�}#c��A#bUc�3D��Z�ł�#�:��'*��]�0Ah�0D���t���+r�Q� �#f��-D�|���ݕ�Ta�]D�0E���8D��1-]��I%�\{L��y�D5D��:ӈէ	�.�1���?��Y�/D�Ti�*T`�F�����T.D�hKT�I�d����ˤ(���t�*D���#�U�5�VQ Bj�DP�:Ѧ(D�h)�!Z0@�(��ƓU���+BG&D��g惗|݄]v}��01d'D���D��?]�P��I�-g��h��e$D��p��W�¬Z�c���q�×7|=FB�I1-f�Ec���i�4�' .N�C�	�<��J��Ƕ&��@�3�K L�C�	=E6ik ˸Rg8Y����,f�,C䉇h�X�ҡ+�B�,EǬ�~'4C�L����M^!�4���m ��C�I�t�dMI��\�:⺼��fC9GؼC�kD>�`̛+�F�	灀<�\B�	 $8�y�D�&,6z�ä^�C�0B�Ɇjל�aw��jH�5*w��grbB�!T~�넎k�8E�?m�HB�)� �p�K�Wn��bG� ��,*�"Oz�i�Դ(��ɷ,[�X�.��"O���sd�6dG�ઑ�I�h��(�"O� 	�	KO@L�1�F�EN�xja"O���
V ��S�˛�q%^��"O�`au����@S��=$0��"O
$[���w��`��j�c|�k0"O�Lpª�#�tS��e�X�S�"O�D:D��,<l�E�+ti��"O��S!Y�Ӓİ"�@�j\���"OdĲ��֎"7f�k��X�M���"O�U����"b����S��l7���"OD!���	h�H'჉o�<""O:��g�)e�v��6�чj��U(D"O�1����Q#`�PD-(��J'"Ob��g�F�~L�"b֢$r���"O�EJС��|n|��g�P3ll"�t"O�����PhS��9nX0"O� #�JӸn�Paf_s["��"O��H�iA�Ko�D��f�PO��B"O�rIΊ�&���d"NK�m,8!�dO*]]r�I!g<�(r��[u!�D�2�*e+�<S"���qÊ�.b!�d�90�hbf�57J@�4�@�5M!�䄬&�:q�PM�e���KU�P9!�/r�V�C�eӞ(�"���	�!��:a�h6 �@Q���6�!���,�B�Cv�C%t� ��h�!�8�.$�G-Jf��c��<u!�Ğ�9FN��p�	z�)�t"�9c!�dF�N�J}H3J��h��(W, <qb!�ĝ�>�p*@,�Ύ EȘuy!�$ٱI64�P`LA�X;�0���c!�S�����l�b��9ТEAc!�+��I�ۙ/���1�%�:`:!�dP
�X7d$���bO�0p)!��^�-��̀��VRlj#n[�w!�$�2c�`է�.f���vM��~o!��2R�VIz o��+��8�4��1�!�$[ >��yjf�G.L v�`v��
q!�#$��\A7&�r�8��	ȓ}S!�d	9��`�A�S�i���̖aD!�ę-H5$!z��c�t��H�SP!�$�h��9��*�Zl�c�%�4|�!�D���d��U�D�M�?`!�dR������� �z�2r�@�E!��>k�J���b5d�����X�k�!�G1I�X�{U�%芐Bk��h�!򄍔<��+ ����r5:�i�)!�$�9Y�� �ЄY=:�J,Ҕ�[-N�!���"���T���F���֡�y�!�U�5�0����ο(��Ě�2S"!�Dg��1�J0h��-S d!�d�5?LFb��P>��Pg�kT!�D�$9��y 0R|������-cM!�GV��@��O�
�z0�|2!�	� ��B':��[���na{B���b8����E�*�r����G�1O|���˸L�hp�*	,Zi��Z�_�!���O\!s�5�v��PE[>#/�`�"O�����\g��AtI��;&�2��4G{��	D4KQ'��2�@?�0P�	�'\�ȁ0Z'���
��^}��yR�'U� p�OZU��Aʃ�
�Ȓ@��� 5a��H;6��1�A�9%6H�c�7�Ip?�~&��˶g�[e�yqA�:H��@�� .$�8�#N�66S&�ё��. ��x#��y���&�zTp%�Ģw�����^��y� �}�"M�-�$^ ��B�y�@�v,ޅ;�d�p��r�ة�~��)�'��g���>z��Q�)�XX�ȓC����P��(Y�xbg
C&6�,����aKH|\<�䛨8�q%�D{��ԧzqK�Gq.�`s�?�y���$i���ˢ�y�V���Ǖ���'��%��Ѩ�0	ӈH������3�l+D�h��^�r;��C֨W}V��3n)��?!���}�&����"�h��D�'q�!��X,�)������]z�ٛi)��hO���;��Z
n;x�Șqt���'���؂t�C� ��bd
2RLd�"�>����f�z�ˢ}٦u�*X�5�i�0Ϛ��Io��ħ<]���gi�a�$�e��1���C�)H�y���0T�� �A�T0FX�ڕ$Q��Ov�"�4�<�D�	�#0.�i��R&���&"4���%�İ��@��
�r��@֍D�<A5�n�P�I�/H.�s�$N�<��G�=mR,YF��g#��@M߹��x���m���x����L���
��F��ē��'t^��Ja�$p�(��ۡ`��j'To�<�5ꉄ���3n]�|R���&[l�<�����w���sn�m.|�U�S�<	�];4�����OwFAT&�h�<Q���g p\�4,��0P��xDI�fX��Fy��Z�s,8BA��á�L��y�ؓ��,Z�A:�U�*E����hO��ʘP ��� �0��2o�I��"O4!��+I���V[Ѿ��V��+;&!�Au���6�N�>�B閡a7!�
0kt|�k��e�B�R�,!��҈haCb�����ì8�!�d��jl�f�̴��
.R�!�DC@�q�U�,�Egֹ)�!���(�>Lx0� =B�tt,YX0��'�B����C�(ھ�!��_(,0���
�'�`�N-g����m�Oc:���'�6x�q)ϩx	�I��9;����'s��b�Չh^�iA�I1iH�0�'rR�Bԉ�8iv���#����'��� Ю��F�L�EmP��
$���d)�'m�����ն�E"��7��d���R�����*~09�i0$m���ȓ�����D�"E`h��S(�o��ȓqE�<�u��n��$+��U���ȓj��d`Y�#�)!b�޽b^��ȓ)^P��º?o>����I�&�>q�	�j�3&��j��0�a��c���ȓb��Գ��D(YlB�r�c��u�ȓ0�Re�5#�8h"~��բ�:+��чȓOR�m�UG��X^�zQ�_�&m+�'�� k�N�}�ɘw˛B~2L��'�Ή{��"�2�a���7B�l�i��ē		�!)M�EpF����>��a��hO�>9k��2F�`7�@ys��	�C^v�<��X�k�ҠS�m�1)T4x"HH�<9c�,X�[����y}�� `RH�' ��8}��>��E��⦪Փy�"�RdA6S�(��	^�IS�2aJ�I�!H��7�Ig6M�O��'j��9�~n:� !��-XG̅�����k��ਔ"ONu���R_"
q�X�PL.p"O�h[Ќ�@ ,m�!
EGl)ɔOB�REi�L�Z�r��£r��� C$}R�'Xx̀qOD�r��ڀ\�i�����'W̱Y�έt-l��LP/~��'����c!�o��x�@R]���RM>��'ț��i>�	F�i�E�х�	�=८C�#�d(TO;�$"�4,��w@���� X�VI(Q�'Oў"}�c�Ƅ3��E*��No�R�B���8_ў��G<�(O��Yw�]<��-3Q�@�v�B4�>�d��O.�� �NJ�"s���q
AjQ8�aB}�x�I�F-���E��s�=�OP�DY���A<�n!+QI�St�l��I@�'��*�OX]f6Q*ƨW�����'kZ�0!ǹ@t2�е��~���J<��4�O���3���2��I
��z���"O���r�0	J�a�5�`��p�D(O
��b�쵋P��>]��0��
a!�',�h@�"�)T+���˞n�!�$L�{�޸���!�irQ��(��z���K�+a>�
G*�6t9@ɘa�!�>��}p��4���D�`I!�d�^�I��|s��0�DG-
S!�dQ�����Æ��� 2��*ga�2>O�干o���(qA�GL=�U��"O6��*\�G�Z�kJF��`��It�O0�iӰʐ> C���l#�⸠�'�R�)`��5��"/�; �D<A�'����g��l�81�ÒH
�Y�'.�� � ����H�"J;��+�2�I{�dÏf�T�BJ<]��A�4M\9@����f���ZB.{��H`S�O7�a��	Z�O�n1�NB�
�4TS��m�2�����:d"|�%N�Q1$8�G-$
sǫ@�<���$%f�jgn���T�A�+�VC����]�,��qf�;7�B�	�N�s����gkB�k&">���iT7;b@9)E�����Y��X�y!�䔵���C�A�pXb�`ԩ��T�'{1O~">r�%yp� �c̋l�8:ul)�h��
g@���MT�)1�H�I��&z\�I3m���Dy�O1OX`�P�Ǻ'�X���$��cW��Q��D�d�>	C����3��D�؅1��Y	h�,����|r�]��(O1�`|@5�T�fFD�0��'vݺ��?Q���\:/+\`#ʛ-h'th�hO!d�!��P*�0T��<T	b$J� ��	-<6�<Οɧu�kٱ)�\l� (��Ô+�/��i�v��a������;`�Iġ�>�-OR�=�;{��0�e��>kb�'H�3`�T�Ɠ.�}��@2�3�E$l�:<��y�ͅb���O��:���GG8�0T юg�6�`
ӓ��'���q W�1ڎ�%C�*5>�x
�'���A\�\�,�I��@	C��	�'cN��%ۈ����ga�:x,��'�XE�/+��1�F�/n�@���'�D�*ハ�J�As!�_!X 69X
�'��E��Sk� `q�X? T��'��eB�jڋqb��*$h8׾mb�'��Q�� /v�|7
H+>�*=�"O0$�u`�1P�U;�-�/D
$��0"O����-D�"��A�!��E˨�:6"O4�c*��Hm���%���z��"OP`�0�^�o��	Rp�T��5��"O� �x���al>�J��Զ�1�"O�=�S�K( ��(k@��?F`�"O�e�ܯ �R�j3`�

��p�"O�@[%��n�tX���AU��"Or:7���Nђe�C!�;7��6"O��4�5aB���S5��"O6�P�B��KԈ��э_/�"ORK3l�9�=�r��!*��u��"O�ܻ�i�/�D���N�H�lm��"O��2&�C�+���`A��_�*P*�"O� ��&Z!Đ�Y��^�a�"O�(cҨ̺�h���S��`Xj�"O�H'#q2��� �*N�xĉw"O@�+��Y���*WO߀�6ݩ "O"��� �06ld���>@2"O\��0d��$���K\�6�RQ�a"OX��Aع4.<���z��6"O���� G���("��8�: ��"O���W)�=��p҃H_06e�(B�"ON��!&]�H&C��"sXa�C"Ob�����l�F�6�E��@"O~��!�Oh�2$Xba��s�N���"O^	 �ؚh}�q ��Y��L*#"O�Mr�1$"�h&�\$�8�� "O�5h��+/ @r��,K����7"O5�S�y���cr�@�6�|;�"O��6�ɟ0tPr䈉��2}X "O8���k��JH�Xj2�CV����"Ozp��"��+������	u���b�'x~H�!c<�|�{0�*H��b��?��u��'Sv�Ya���T�q'�����'�I�DnZ�,�F��j���H�'n�@ ��>)��9m��rD*��'�0�PF�>f:���GLl���@�'r���E�rl���ցo ��'�
��נ)
���sf� Q=���'���@C�r��\#��R�Ue^h8�'t����/{�ft�j݈L{��+�'ɾ�ʥ�\(T�RY�G�I���	�' ��D�L>= �1��!F���s�'E0����� T��510��kr�� �'7R@��(��v|�1�#��R��'r\�*B�Q�u�̑H�.D��'�4!i��Y-#�D-�v��	n���'F�$�-M�)��&!��hr
�'-8 +`��i0$��5�4etR�'�%�$��z��ܙ��	�T�$��'�(!���*\g�%���2C�}��'�#򣃢�d�д1N�e��'��i[@"�,q�(��蛖ZH����~ƈd3��	A��(����F�(��f�l�s@o̢m^.�	�k�+�b���+0*�+�͇�O(��ܟ�����T�DK'�F%V��p��t��y��L�S�$x=Jx��A�U!��-��\��û6�E�'MZ-`�����(*��R\�><�tA�8Ɔ݅�UG�I�����J�"�0O{(����*�1�nͷB(^�@`	q��}��|�&-���&�0���^L}X��Cr�=
�e :x\P �B�V� ��q��D�f�޽??*��%FҼ6�l��ȓO�(�!���R�r��v׾x��хȓn�~��0-ʹ�ҕ���L�q����S�? ���I��B~�}�"���d��"Oʕ7��;�5���@Ǭh��"O�q��˚|7�9��f����%"O��)7��|��R�)5O�>P�@"O.�x��\pu���ԩHS�05"O䡺���=.�l��'�!)��#�"OV� w�Lx`�����z��5k"Op��E@�<r@в�e�,5��ɇ"O��ȶgL�S�H��G��P��a@"O�Ms�F�-L��h�5]����"O�TQ��2o~L94&R2f�ļ��"O�����.FbA
�%�!hẼ��"O(ݒ�a��i^1�7��3(�x �w"O����%h�*����@ތѣ�"O|��H� 	(�DA��ӛ=�X�c"O�uA)jV�1:C,T�����"O��Ӷ'U!��|�᜛B���&"O(��Qbh�j^�d�����"Ó M7����L�!J�hH�'�vAI�N[S�����)>��Q8�'^(�x&/V9g��k hDI�X�	�'ܮt����Z.dT��#-�Hy	�'�ri�f͑�O,��ƪ����@p�'�
��e;���Jvn��KD}��'Dp+Aj��j�V��(�M����'�� ��BJ�Z�䡘��T�w\̈R�' �5����FaƘ{�+	;kU6	�'�ؑ�m���cpm�m���2	�'^����Jl̩�2�Xm� =)�'�h��8�*�i̦7h�k�'#f,���ڲi���ajQ�>�u��'{�l���B�K�n]��������'W��Z`�	76����P�"��'�x��ʉWҐ�td�=Ft5��'����� ��S�*ɋ#���'&6Dj띡��!cdǈ�����'�0d���`i
��� �9b���'�J�`�&K1*c�!�`�/L�PP��'�áBK(MR���ە;�
�!�'�9���-F��9g�������'���R��l�y�F���6$���2,���aӞQ��[P�ΰ���� A�a�F"On�kG)�JB�iCS�e>�3T�ɡk3С��Ae�O���Z2������M�/����	�'8�-c�Ǹeݬ�#�O��2�����_�4�p�c�m���)����cT5#q���uB��rlD��*D��s�ƔS�r�j®�zL�Q�3쨟�z��v+��C��'咸S��:6W^a#O�6t�	1�p��-H�D�;'���u�ݧ5�<��`jI0]���t�1D��$L��(�:	�3�5s(2�v�,=a#��.�,#|Zg"MT<��
AP&R�zGk�f�<a��}�`,ِ� ��|j��,ŉ��Ǒ� ��O?��C&)�D�	��כq'��!��C4�!�䝠bxl�U�A ner�^��$S�A�� R�듊�0=����*���L�$ "O3\]���$�k�~i��EE3UZ2���^�0~�����&w':l)�'d�Ѥgi�6���ʖ}���#����7�|�+&ʧ'MȬh���u�����K�2R��0�ȓ(d�(KAe��%�<r�F�+ Ĭ�b��V2Kb�O\	� Ŕ�(�T��K0�X�B�0.�KW	�W)8B�;�e E'�� ��	 =,��3�Q�Qp��Q��\w�u剨Xm�EAJ;<����T��^
��$��c�4ɋ���y�*{P�Q��t��@��M� JQ���g�ٔƹH�	1}����(���֦C�e��=y���0�Bm�񨳟Lz�Cۙ�X�:�� p1�!���W0���W#F1�d]�s"O� �M�7S;�#���=q谝q"Mtհa��Y0#*�;�NZ�3*������y'k6|O)�DخsPL�qo��yBA͟[J�#&n[�@0D��U���e��<h,5�	�A�d�iE�XR%؋���	>�*��E�Q�T���JJ=3l�zr�T5P�&��"o��B"� �EQ%��]�����R�@��P1O����	�f|��ꅲIe�cP-��L"��8��M�$Έܰc�Q%�ej ��o�d}2a<����CG!i�f4qa-\4g����"ON9��Y#;�Vy���w�� ��'T-}�!�s�U&9���!7j�M{B-���)H'�y� W:e���h	=}S�ђ�X�y�f���H��ð��U��J�?u��X�\�>�7��*�Q�[w9�U+�	 ��x�SщaY��k��J,�����Z�^�̺`�Y��Ĵ��D,$�Z)��.̥y��\�g�@(7�@�R�����>��&ޭ���Q'��|�`���j�'�V�£ş\���'>�YA�*H��`�חv�"%.D��р�7�.i�0gԗR�Y̣<���CRXD�GI<}��)ɞ+G�0b7a�&��dZ� K	!�J��Ҥyf�s�΀ b�S wX����0��+dF�y����ɌN]F�;#�g�P�2�@0^�������P��d%Ƨ/!�Q�G�$N��] ��	S:�D��}%!���7�J{�&��w�{�E?8Y�O\p�oNE��P2u���OV6��E�0}^���eƁtz]�'+ܤ!ǥ\�|�jq�p�|�()�B�pY�A�*ַ���"�(��	!�,��Ƀ�*fp(WD�<,�B�I�8��9PR"4U�!$R�8�pt���s��U��4F*i��@͢�P&e]y�Zq[� ;{����<W���s�����dZF��2��8kC�
3Z�Н*�J��Xm ���7��8��.�h��۵���S�"X.؈��<A�/ߘ�C@΄n<�I;Q)�97(��B���?uq�62hul�"�4<���;D�t�f�.HE�Ak�;{�,��E��h/���� ��ʨ�'���Z�m�F"(�)A]��]�5��	$LL�Đ�L��KC�	=5�䪧'� V
����F�]�=ʱcK�zun- e �.,7x��%�P�1���7gVB�'�ܰF%ԺP��$t�n	��	�P��09��Oh��iƈ)b�l0:���.�+�:X�.=�eIF"@�P�����0>1����ln2(X���[.<���U��_$ �fh�Tv���F&B*�d(qÐh�ZUͧ>3�u� #��WbA!�l[�&Ѻ�ȓ:Dl��b��S~�,�Q�P%.��G)��iEG�AMb�?Cf�$?QH�B����Q��2O�v�Y�������7ʟ~�������ƋHn<�ps �%b���
ТA����$��0.�
�b��.�
=:���Jh,�0��,r�$�x d�0��r���##K ���3ړO�
QL�3G�ZeÀ�INI�D�tQ,�U��̔,T!*��l��N�*4H�хI�B�zeB�~������C��$z�1�N�23�HHl0"�.\1yz�̈G�ig�I�p�IE�ҍ3f�O�����Fۧ���xd*]9`�����5v($�$�zs�!c��$Bc�.-�8�I*O����M�z�J~�=rA�K�0=�$�*cИafD	#� �DҐJ�p�z���ئ-�b>iZ"IS/Q����#���N�b6h"���)k����J˒j�`X�A�fX�)E���#��ݘtJ�&�d`�QIB�=�����^9/���K�4�0�#	_�;R��ʋ8&�fh�1�B�8����t��%�1d?���+1�6�����>�HO��2dٱ���FOq�V�K���,M�-SČE
q�z�B�|$�g�QD�\0�`'�d. ��g���t�=A���O�M�iC-!��I� �bLY��i�*q���>1�ʵ ��(^h�ҋ[@��}�1b�Ԡ��*CxhŐF�R9b�r���J,�r$��m�<����nF{r
Y
)F�`�P%�_x�YP�C����R$N�Q�$�P��'��4y�i�l�A�B��E�������$H��qQT��. �,��F*d�jİ<Q&��!�L���РaI��#c�Z�koR!)T
�
��I�sרXs�:O\@H���"�܍mJ�4���͟P\ �<y��@)��(S���"`��\IF�n�O��HB��&n��1�И�Ƅ�"�'��]�A����Q *����r���F<f逖������\��y�#ikL��=E���=|al8����"S��U�w,\�&����Ǹb,^�|��=y��hO&���ϱ-ڦ�� �Ѩyhat�'��	�Ed�
$��hA,�JB�I��(D/���p��Q�<�oǾb�ؑQHۑr�f	��N�q�'��Ѡ��_�W�Q>�z�%�[�XE��G�<HJ0 (D�H���ڑc�f?P Q��rq���Q�;�a�{���)��$y�"U'f"H�����7�B�I�<��D�$��"4�&Tht�^�|�.B�)� l����
���AX�E=���bv"O����	7&K,}�p�IGt2�*�"O��C��K.�@Ǌ�m 2�"O�"GE(�e2�Z*TF�!�"O�pF	|L����6f��س"O�$���+�B��b��4hn
�"O�H��4�TP�&ĩELؽA"O�T)��Hx�o�#<0j�kQ"O��FH�u�|A�J�J#�;F"O �5�<$�%B#m�&{�$:�"O���˒.e��Hv��.b����"O��)��G&f~PceJ��.6����"O�8��C8<r�$�j1W*j�Yt"O�u��V�4�0���j�E"Orh{�@Ф^4t����Ǐ;i��"O�P!`��%7u~����Ʌ`4����"OaA�Oߩ_|,d�7�ӈ��"OXekEh=��̀��ͯ)��t�u"O��P���k��IQ�� G��i1"Ot��5·.����)��(�pТ�"Ol����`�����6_�&9�"OV�2k `���_ҴTg"ON\� ��h�n�H�[�-���"O�MZ�̅;f����nȗ��e��"O����M��[�,둃�g����"On��`$�F���hN�B���"O�m`$F  p�r���$���4"O�A�1JQ(4�r4��J�r}PE"O���
Ξ,!��)�,��&s"O�y��¼CWTD��i�? I��"O���t��,Dh�ڱ�ϟp�+�"O��!m�"�g0%/lp*d"Oh����Z.�Ve���
�"O���'�K~,�R����zS"O��*F��v�D�'�Q� 搊f"O��#�L'$D���$*�Z�Ӣ"O��8�/.@�`��:6�8p7"OH��ł.��V�\�)6�Pcg"O��S�È	:�l��a"�<fr4�Xa"Ot����v���Cv$J��b"O��A��x�Ju�ݕ'��5J�"O�=�B���dX�!Cq��"O�-5��"H��@�6��d.D��"O<�h�
5/4��	!+�0�G"O�}��*����(��ζ ��W"O`aD��{��	�KK�x��h�"O|<�ܛ ���+g���R��i��"O�4H�;Or�B�	�ݚݰ�"Onu�S��=��ģ�� �:cڵ��"O\� e��^L���glz�"O&��aa�i�*�0(p(��W"O�ݱ2��;ț��ԮB
N�X|��"O��ز`դaQdĹ��;Ό�i"O*Q��L˳4m ȱSIŋV�ܜ�"Oh�R%�[:���P�۾i���ca"O0�s�]X(@<J#a�73a<M�"O�m�#_�^)b�{��S�{j��)T"O|1�p�r�d̉Ao�|}p��"O6hZ���hE`T��(Q�tI	"O����24���� ��9n��`D"O��"`���g�J���V�bP�8a�"O�E�3��3G ��R�JO�a��"OH+"���qzx�
��*1
D"O��y&`��BG�Q3w�8$�n���"O� \!E�,�.u�s�Łr��x�t"O�-��&k"��g�t��k�"O*a��H0
z�(3&P��p�r'"O���¡Y�����N�r<{�"O���oϥ(r������
k��L��"O`��V��i�JQ���Ϲ'����"OJ�W�b��i�W�χ]{0H
A"Oj	8 �"e�`a��6UZ��"O:ɱ�J�E��⤓>4��P"OD����ʳf�xk���>s��:�"O�(�Q�~���A����8s��iR!���
06IR6�ʻ�(<��폽,#!�$K1��K�Aӵ�:7mMs�!��hk4�H�g���{d��/]�!�ė2��q���Y��\�{ Z�b!�$Ԕ���B�b����{�� �l!�$	7���A���]v�x�-��"o!�&f�Z{��P_�X��ȟnI!�4�@2팷V���A��6!��W�0��+#DV���(��K��*�!��43�d��
�y�R��u8l�!�d� ����PL�2Qũ�'V!�d�_V�,�R�� ����x�!�D%4ӊ��¾`���g��!򄙓" N(���4	ug���!�,���mS
�4j�i��!�D�R�}y�!�MZSM<6y!��R]pJ1D{�z��4iT'!�@��0y��M��hD�X!�W�*�*%�+T)84�Qh��:7!�䌸\�� bq�-?����$����"O�)3GtH�a$[�1�D��"O�|��� ]�����:7�:���"OX��f��xN^HЗ)�M��Pp�"O.(Ic�Y�+�D��hF�>����"O�P{@K��y\�YK��Q�Н��"O �Z�&P9@>D2��P�<ޘ	k�"O�u9kK�9q��RP���-2P"O�9�d����8��Q�_y���"O��R���=
�+f�)Kc�@��"O�I��.�v� �Fy[��H6"O�Ͱ��F�R7�|3)I���"O���샴RL]���H������"OpՃ���r�t۶�H�a����p"Oġ���α[�t��K�90�Z9���'�^1��\ʦ�C�˃�3[`�����G�`�9� D��3�
�r҆`�RU�N!�Y�� �f��Y Ϲ�(����+��DܴP!dJ�{,�\��"O���B��#y�;#m�/f���R���.�d	���2��S��?Q�S!M���3I�m�0�##q�<�5�U�Z���k&O�6O�q%��s?Y�^1| ,�Ib�(LOr����-'vI��ʂ:\RJ1�'�'�zUyH�����r��;��*D��5�Q�UC�\�<	�`ô����s,�1-�ٳ���Z�'�d�Yp�·���G�䊁�N���r�	�����E��y��^�P�!8Չ�Dh`��(�2u��U����H�"~��F+�I��EB!p��"De�rC�I<G� ]��+�.h���2�AK�o�t���]Wdi��0XazR�΅h��XC#R�m��#��2�p>Q`/��|�>��Sڗ`��Z�l�#wLh!��ٖLdC�I�~&L�c,C�zS�� �,bV"=y�"	�=.�9��Ɋ<��͑.�|j2��'FX23�!�$��zzP�X�f�aX�"�o;u�V���G��$n"��|�ܡӵ�$�'�y7jR�j��P�v�2�: � %�y
� ��+0
O(2]d���`p�J� ����ѢS������#���(Od��5�5ߺ��FČ>p��Hh��'`���<-�m�&������t�p(	1��g�|a�(�0j�x�O�R�P��d�gH�}��OQ�BȠ9�'��!fV��Rg��&)��>F	��$9���kă/�f]���´*>��"��2�yb�<v6�Lˣ�q���+��_t��/g��ѓ�Mr�"��8O��}��}�!�u�ܵ�ŉ�Ly8z0���!�-!V��h`,^}yL5Ra�;b���B҅���������#�t�v���#Q���ɖj���  ��5/��:6$�9Yb������=)���YY�=Z�(A������5fX����Nɢ]�<Cp)�8-t�Es�WM���A�}�x��B�3-͎�=a� ��c͔܈�(ھO^�7  �IY6Lh>��c"��b`���ceB]��(D���Q�G���)'�9��,�l�±��hCֹ2 PyR��A��-��O�`�̻?��є�^0^YL���`�b���3p���a��= ��G"�#	ENaSg�;�\�s z#6ꐤ�Ǻ�΄�(O0��4Ɯ�z���eҖz�
R�'^"e���� �:���� .�d��#��+�8��f�1�2�F�o8�����[��P�*��U?�M��D' 4�?a���	�Bݐv	:�I��<�Ji ��;A��"D��$!�L�P���ZWf�6u��.�  ��	�P���Ad F�I�S�O�>p�UfS��V�p`���vG�Dr�'8����!�(wܣ��j.�p��|�h+�`���y��J�Fi��`� ����q� �Pxr��#42���>4�jm�E�Lt�V0�`c�I<��^)��N"����ɝ���*D65b�f���`�/��y�ȓEƄ"�l�M�( �$dV�SY���ȓ|�dM��[�{b��+���x���NY����Ӽ老as,�Sz1��v�%"%mBn؈�p	�y�@���:4�q �"�|I��_�o8�P�	�$%" �'�.1
�&ߏ1�$t�!��= ���.7�M�� ��~"�P�]X:�a��U����h�b�1�y���s �4��2��@:S�7��'w$��3c�n@��G��&V4b��-@����LM�ub�)�yb�ߧ:>.��	H.x �e�H�U�c#���	�:*Q>˓_�J�)q
���=f�ӡiW����ɝO��U��2Od�! b��y�a��'��CJ0��B�� '2��W�=xa|����$�R�B�#
Zv:\�C�Oy���I>'K��ɔ��D��L�8
�L7	���95�:UH �A�tx4��'���!�KP.7�������cǆI����a�
�ZSo�O�,��r���1���>�t����V8?0�`�O׮i����@�'W�I0�㞞g_V��bM7R-��$	�|��ir%��,��Dcu��sJ���X���"��5V%��!�D)�DDEW���C�@%.(z�bj���=a"�#)�@ȩ���9��P%'n6�ó2I	���6�%YM5>�88;��Q�IV$Y� '5�\�K�8X�F!�S�N!��h$cM�~��]�qJ� �6D2�kJɾp�,6¡u�؊������T.߄�.���5�a�S�����D�x�%`U�+|h3-O�z�mVV⠒�qO�D��b���±�`�NSVA�É�/'~H�N�b@�de�p;�@ͧ�Α%�<��%�z{b!JvA���ro�<��Y�g�g��򤞻rh5�Pώ�qF.9����8��ۥa�	�,�4&[^�A�Ý�{�0��c�HJ��r6�	�W���� �lj��+�'3���z������484�O�1����5�i���J��P��ԭ��txQ�It�n�[S�L J���0�&���q���:2�ДQ��]��?Y%�ͻnG�]:��7<��qt�ئ�Q��	�M��Ȧ�'���1��̚v�Q>�ػp`ɤ�O�C�~Ec�B�7\��C�G�M��j�V�E�8��?�=���E؞0���hÄ��ƣB+�49I��I"(ٶ�Ƚ�y�OM��I� �����#HFִ8���
G�CR�� ��R"̉fA�P��'A�=�E��Ȇ,K�LN#� Cc��p$�a/|�(Gx"�`ŀ��Ңğgo��G΄p���U;�0U9���$sC<�{�#O�hO�}P��,NW"|��MP:�Z�����;w7B0�/Ĭ	���`.T��['�D�<�@�F��K�L���H<r��뵂ĨF`�Γ
j�̓g9�)�'ZGf�۵	%�B];�+��O+�e�'��)2lU�g�Z�ꔢ@`F{bj��:����mH;���w"�p>�6�^�rG�N��:����,or}C�R
%�B�ɹ;4��2A�7"�V{&��'�"=)@f��t
l���� ��3��أw��)����ǰ]�V"OdUj��1�4в����R����'�s�Cm�S�O�@C�@�M�����A�l�R��"O��z��͠C���g��XF"OJ 
��E2@60�5	��Zq��c"O�XA�VY��@3I��$�4"O�}��� �56�Q���,����"Ol�8�۳\�*qb!�{�I�"O�h#�%�)f�pEY��;,�6`��"O�����&�h�� \)U��<��"O��!$�P�֩x��7h�*䐠"OV�y�iP<q�꽻��[�a�(���"O�ѱ�`��r���o�9}8ja�"O�`+�h
<mݮM"A��:E�p�K"O4Q��Y����Ic��}SP���"O8i3�O��Ca� �� V�)M$�Y�"Of	[�GH<M:F<���.z2��t"O�0�2$y0���4Z�$�$�S"O�0�� ��.0\�ʷ��>���"OiK�BW6be(y"��Y�Cׄ��"O~m���Еh��8kA�Ə$�bL�"O�Uq����yia�
�"��Iz�"O 4��凡Jؤi��X�(� 岥"O$a��a��48�����G�Mr���"Or��dU������z{^�T"O���@�fP<%��8���ZB"O����ܲ1�.Ę���/G+͐b�<�B�`qSŘ%�)��]�<1ѪL��Xyp��$`(Q�C�U�<9���n,ʉ�2-�#�x0� P�<i�(�Q�dȂ�� g�p�5"�N�<A����!����6K�	 ���H�<!�H�D��y����>~*��gUD�<ɕA��y�h�#��K�7 �YC3�DF�<���Q�i��� o��Q�W|�<�#�͞���,M��F�3���<��#��#C1{�
	db䃃)�v�����Z��� ��;Px5JaD��@	&�R�)#D��i�l�*�.���,�}���a�>D�x��� �9$���딪'���O<D�� �ޚ~,T�'��8.�hC�(D��K )I�G'&�#�F����`!'D�p�WO[�pW�1)�3,E~��1�&D��G_&Hr�PJ@+��|��C�	�2��%"�*�5P>.��,�2��C�	��h�go��a�8����Y7�C�ɻa�nѫ�NH�d�6`�RE*f���r�yN���B�^ P��,.�~!l�6�Z��' �K�)�m��;��������L�T��F��>c^�t��yR�O�����ݚn��Tc�GʰS>t��pO�o�S?v���'NLC'.Ȯ!�x������4U$����(�"�6QD�����gښ?��b�T2?���3L��~�P��]�a��m���C�>���X�o�P-3@��8��p0�C�Py�Dف2����I�(	Lk%P����Ƶ0��OȴP��OF(���'��TZ�fcaAc��Ē'LR8Ù'l�9fq�(q�T��}R�)ڪtzp��F�!�0�0�Ϝ���Bw��O�Z����	51lIX�`�A6е��dQ,�T��D�EF���1n�}��Rs  �,�ee��(򫐃{@.Q8/O��Y2��/B�b>%�,M�I3�T�o��^�D!@RyBm ?u�xEQ�����@���O�v�ߢ�
XB��_o���JR�v6�)�����t������ ;�&�cg�~�)�)�'�0��䃶��ytD˾3�py"aLӟl�MQ�?1�YB���Q�2��ԋZ.u��͠`AN�t��O*\��O�r��Bc�a�A*�o�'JD��'��E�cG�r���GB�*!}��:��� �8b��~�zQ�b�L$f>�q8�"Oyb$�����q��D�D �kb"O�����Й��(���ܲ(.�1"O)S�˞�q�Uт�$=6>!��"O��S"�N6G���;C�3�Y�c"OB<k��������-�@��aÇ"O̅KT!��A*�īZ8v+�"O6Y�����i�D\�:rNi��"O$�&�P^�X�7%U�m��"O�Q�C��a)���'EFh���"O����)�p(ر
ڱS4 ��"O0��wʈ�7{TH�F��0{�\r�"O�h�A�(}�n�cg+G <�t��"O�(H��?A�H5p�*�"X�TӲ"O<�)c��9+�(�7H�.u���"O<��2`T�|A֭��ȣ.�6�R�"O(x�fG6AlyڵmX��x�1u"O�:��	>�@,�+U _.���"O�H����C�R@��k� ��K�"O"0
�i��]o��)_d��;"OQ�
ݚ/U�h�w�H�UV��	�"O� x����
|��SV�<AX0K�*O2p��#V��$l�a��c~<	�'�m�b���B��S/]U�!��'\vS0M}}�$ʃB�+X���	�'O�yQ�R5\tx��Q�����'�`�[���y��:���!��h+�'z�� �/C<^p��
��A�q#�'�tıe)U�@�2�4c!C��X�'�6�aef���%
̦B����nT�<!a!���U���	 m�	���P�<�sÜ%4��,����	`��X(4IO�<��kX�s�](#�0n��s@D�s�<�1�!6� h2 �c�d�X"`u�<�1噢UD�Qn��"�I8�b�W�<Y�@ (c�ڄ���F�"����V�<�q�K�8�����(�~�c�˛T�<��	���!;��:@�����GT�< ��2#u,���V"�^D[��L�<� ݧ�9 U��zF��b��a�<Qsϓ�q2��"��r���۷)�B�<Yf�B��&��#�n��\���x�<٧,ʦyΈ�j��C�K��!Nu�<�B-�%��:V�@3[��B�B�|�<�4�ĒG�XtX�iQ�� `�N~�<y�S_��U��J���X8rO[C�<�PO�E��
'��:�6Yc7#M~�<��� �WdB��#$C���t�_}�<� �?@QP1p��P�oJeo�c�<�5��2|��S�-^�$$�a�E�<aע�q������Ҋf-*|�6- A�<�R�Öl���z$�Ų$V���e�W�<ݫYp��鶧AUnz	�'�o�<�4��\��SW��.P��"G�D�<Qc��
a��P[��5MHA!t�\A�<��ʅ^5.!H��

\���b�UX�<�D��.�����d�'�V�+E��U�<���ć��{�Vv,��B�w�<����'
��T`�:.�R�J�j�q�<�R*���%z��3+���j�i�<�� ��|AΡ"ЄE�Q pA�F�J�<�� }y�(���%7*x�A�M^�<��ˍ*gx�xD�Δ2R�y�4�J[�<ɢBP?I'�k2�	D)�"�FX�<� 6�gh͎x����@����"O�|Z4�	�j��[� 
&%��<(e"O��"o�6a@)3c �7k��!2"O&�rTl���V�t��fx� "OZ0SF#�T�t(H���|�|���"Ol(���*`��@���`��"ONѣ�+J
>�� ʥ�%�@��"O���Ӧ�<��xڀ�ң�
$�"OD���Ə 3�D���?{f"OlpɁA�3u) �4�H�t���F"O�Тl����%d�C��"OR� 4jYK�DX�u�	F��D� "O��xՆ�	+���K����W
��"OR�
3χ�(l��a�N_73h��sp"Oؠr�\�ˆP�tM�72t���F"O��e��n��| T��.XKP���"O�H�#�0�b��@H:��&"O�!+�UOu�W(q"O�TE?@�e��.A:y)���t"O`�!� ^��f�A���R(Tj#"O�Xa��K��9����>�
�`�"OL�ڂϨz�q肨�(:��H0�"O�Q:�dP>P���b]�Y�3���Pyb�B#|����4	� B��L�<Yă�>%2�*���t�$%��+�G�<Q5��-���-��:�f��`M�@�<qR��:6�� @�����+�g�<�����>���Ⱦ&��`CoVY�<y�ə�>�F�ڦ��4$<�9�H�\�<g������򌇶r�\q��iTt�<��8\�H���핈UF��F�o�<�5C�&и}�U&A��^���A�A�<Q���UO��!�^&$R��Da�h�<���U�0�Ccǉ�W�5Ba�H�<�����	\h��fD�!P�r��Tz�<@Viݜ ��d�ty��R�EN�<����)ʅ��B�=$p���K]F�<��ۏQ�n�&�E!JZ�`R����<����-b�,��Iʵ}>�b�iEU�<id��\$*���zu���gf�Y�<��e�cժ���$�c��E�U�<�0���vp��K G^� u��D̈Y�<��dO�p�zQ6��\�`��,|�<1���)PJ�	��
� ��m fKz�<	�;D�n�x$ƛ�7�m��v�<A ��
	 y ��$�����o�<y"痣�D��5��l��F�T�<y���k:8��dQ�`8�r���k�<٠�E+���Q���<P�J���GQ�<!Ĉۼ%l4�º2H�<���r�<Y�Y+LH�ۅǋ�lj��3rD�n�<�I�vfȍ��+��k��ŋĈh�<b�Z}���#�x0)��m�<�NN(8m�!b}	�9)2��j�<�A�����4�%A��yX��^�<��*���mҶ�V%~��q�b�D�<9w�WM�N]S#)�*�|哓D�<)��\�g/6t�ѝdZ
�;w̅�<I��V
	B<d�A�J�v1�Ӆ
d�<��Ҵ/�Y;W�}X0c�"L�<����a���+�$��$�:կ�Q�<�'�!�v��&,�.�z ��X�<�eI�'iy�=QF!U9gXP��F��|�<Y4aE�p`K�+�	t$�ee^~�<� ���Br��gY1B��""O�9xqhA^�
�jC�lۦA�T"O&в.�G�\x�򀄡cɈT��"O��ze�		=�<y	r@��ޙi�"O� �cP�.F`��@��	�z5A�"O���D"ɝw��x�+��"��"O�AFER�M�r����K�\�f@r�"O¤�QI5+8�!"P[�D�w"O��X#�%H�B��C��f�"O�h��B�C� �#�&]�nu�"O�.�`񸰇İ"�&�XG萕7!�D�`�.��%�>2�F$0A!Z'^!�D�~����F�G�h�Y6�M9�!�D�$�P1���8���JV�>�!�Ē\�
�;W�ǯt��A�ЮU:�!�S��ʘc+Ր<b��p�n�t�!�<_L����1p�]�FM͍U�!�C)c
0�)K8>�
���N	!�m���r
/�<
��Z;�!��\Z0�����w����R,!�Ę >�8Q�l�G
���F�O/!�$�:�ѺweQB���*�
!��		�9�̘�������
���~����`8`����Q�LW���di�ZƄ�.�Br�#VU`1�ȓji����E��ݩ�(��&{H1�ȓ)���0��&��D���[�c!.$����$+G2.b�h�&.-�&"O���W)�<>&�����Y,���"Oh�r4���q:�⟙/�H<��"OF�R�B��D�"�pH��q�(���"Ox� #`�V��'��?H��:�"O�|�T ؿ|���3F@�8�4J@"O�iF�ߙ^�@�k�!D��r@"O�җ��MR��F�Db����"ONY���*D��
�.E=�R��r"O��Ȅ�*Z@J|JV��#f��r�"O8 c��Z%O��y��U�E�\a)�"O��(@�Y�923LR�k[bT"OZ��Q�	dY(���D�3XX�a��"O���0�l�$=V��t�G"O.Ѹ`-[6pr���$��#-���˴"O��ѡ�ۓ.���i�'M5!�^,1�"OX�S�,V��5�7fR��>�g"O 5(� ��l y���J�N���"OXH�E��.&���0-�`�'"O�q�)�Y3�P&�ӻo��"O�`��D&h��	\8Ze���p"O���R.m���;s�P,0`�1"O��AFmY�]��4�Da�D�Lp�"Ov����
���9b�0��kv"O���B!�\<@Q)R��+�*@Pw"Or0Y5�K�0��a��L�.��-��"O���0"6C�a!�*أJ���b�"Of)� I�
[��)pCD���-Ca"O�8{eF<_� 3��C(=��"O�
�I�9Z(dZ� �{*N��"OL�T�PwH|����
o9�*"O�ı�ßg��T1��?/�8+&"O����)�m8Ĉ"@�B-vt�4	�"O!����8o/2����R���3"O��B���0�e�5�7B��0�"O�Ũ�fP�<'�mQ��596��"O��C�.�.���1�F5H�q"O� |@ؗH�%4v�
�d��k2Ҹ��"Ov �Ƃ��LҢ�^͖�R�"ORp��
   ��     G  �  �  r*  56  �A  �M  GY  �d  Pp   |  ��  �  \�  I�  ح  4�  ��  ��  �  U�  ��  �  ��  *�  ��  "�  x�  � *	 x � � �" �) 0 j8 �@ �G aO lV ] d Mj �p �q  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbE�X���Ț��<��FU0ݰM��E2<P���4��v(<a���%>Cd�e��O[ �E�D�yp���C
Or%��J�H/�L�%h֨k�� ��'2X#<��'vJf��u�� ��9b�w�<�+8��uȧㅕ!Q�$H��K�<�R�H��T H�|�1R�	GE�<!F
D��&0S��*X��QӅ�h�<�3+��~U���Ó2^����b�<�TE���ؚJб�l��C�R�<g ,�dZu�M $Ւ���Q�<�ծ�'�8��'^7z��$c���K�<ЀQ�1��M���B.<@��΁E�<)��K����1�[�P ���C�<�� �+@�`�UGB�X�>`���W�<Y�.7E��4�P.��~wh`:�Pn�<��'S)"��%ʚ�6,�2 �l�<	aN��8��끇ݳFM���a�j�<���B�5ܜ����;q���Sk�h�<t���ER3Κ�Ua 9a�\f�<��%�4AZ���&Nc��ʚa�<���� �F�+�Y0:<����JF[�<�R����� &g��!�D�QgZ`�<��,9h�2�F���I����\�<�peJ81-@<�A&[a[�D�<���q�"���`�8�U�q�B�<���\�%еi_�vI� dPc�<y�)"b��@Q/C8�d�B�i�<y k�$<�B=��j��?�$Ei�b�\�<��υ�#]�A�)T":����b^r�<�SjԲA�c6�<�,va�m�<I����a�>?h`W@�q�<���{��8�Q��.�SEc�o�<��蟿{��X���B#p���Q�INR�<i�
C��JD��M�]���\N�<�@a\Yq��R�v��@��DTH�<QB��6�.�bb�űEU�A��DZI�<��b�F��2�슯�F�p��@�<Y 8v�l��Ü/l��DK�|�<�$��
I���{��D*���Ҷ�]D�<)�C�]0�� &o�����c~�<�#ԫ�2�$$H�f��=B��L~�<��KZ5z�8)kd�E,U�������v�<�3�ϡk�z0D(R�~f<zWm�h�<q���0e:<�S��άI,��qd�g�<���f7�01B��(Y,U��Fg�<qPGG�JM:yd	�A�Sq
�H�<��fH#.�"y�"o���Cݘ�y`�"`�x��S7�p�ч-��yρؖ�9���ã(��Yb�ė��y�CE3r��lZW�8X�nD3����y2a�S��帑���Aj�I���y��oxD�׎C�R�~)�F*���y���c���ud&~�n0����y�����h`"��q*hD�#�V8�y�ʬ*4�P��֚;VQ
ώ�y��ۡB{���N�2,�5Rb��	�y���/#A2$+"$��'�����Y�y�lԠ:�
�вH�q~Y�i;�yR��&6U�h U�Ôn͔D��F۟�y��K:�|K�a@�e�\0��yr�M�>PA�_;sy ��/5�y
� �(X��	7����V䋣{�ԭq1"O���E��T�nb �H�o.D��)��ʏDfda��2�ES�i,D��k�F$+\�� ��Q�r�J��+D� P7�E����KE��YW^�ْ�Oh��Or�D�O��$�O����OJ�D�Ot�h�Í)-��yz]�|��1h\�?����?Q��?���?����?���?�c/�?m?2�ck�ZDp�Se��?)���?y��?���?���?I��?Y�!��khr1:�(�.Z��@�@�?A���?���?Y���?���?���?1Vh�Y�֠����%i���K'�I�?i��?I��?���?��?��?���si�)��^�T�X\�p����?����?����?���?1��?y���?��@|��X5� ^�&1Bf4�?9��?9���?Y��?���?��?I����
I�����!R�� �����?Q��?���?����?���?����?��������W!Ǳc�d8�3�ߛ�?���?9��?����?���?����?���4X�#� ��,�p�S��?����?Y���?����?���?���?��D�����/
��'$P��?���?��?I���?9��?y��?�&�[�6b���T�*ܼ Q�ۏ�?���?����?����?���?q���?a�	�YIZ�R����d!!2H
	�?a���?����?)���?��O��F�'c��R�e�l��E�*V�B�Q��3.˓�?)O1��	��M��I�c:��w�0H,����!�(@�'Ξ6-&�i>���̑7��$�@,�'E�<�� @E��̟�	�'!��lZh~�8��M�Sc��1-�=Bf��FD��P�\�1OF���<1����
G�l��E�=1.`au�G4{�Ҥm�f�jb�x��d��y7b(xJ��A0"�*D1���.Yc��'6��>�|B7���M��'="��잦(������.�*���'��D؟�2��i>����Kp����5��I#�E^_3�	@y2�|bc|�|a��V�.�*�喾z�+�䜮`j�$�O����O���o}"���6!3)�[���ˉ8����O�[���q�1��S�q���$ǦX �0�R�jyTa��d�pʓ��D�O?��if�B���tҺI�`�)���I&�MsWw~Үz�0��^%Hy �e�,���J�5R�x�ן��	��H���Zʦ��'����?� %�E�:��TI��_��;�Ǫ\ў�S`yB��t䋻2a0E�,�Y��u�B�������)�v+�Ip��C��(�����U07���KG���d�O�g��&>=�	؟�����CVdܳ@� �V$
��Р/���9t��>iQ�mӸ��b�'V��'�t�'2��@-M +������-�>��5�'��^y"�|�Dl�dȺg;O@t�P-GDFh� #�R�0O�L��<O.�lZM��|��?)���?Q�j8 ,���  d��H��E/�ߴ�yҠ̐���O�?E���"���/u|kl�>*(�6�ʣmwd�2�bA�]���O�����S�;�2�����a�
�(�&Ǹ9Vc�8۴! ƨ�'ƈ7 �dK�!Ŋ��@��� R�	�db�-l���X}"�'Nb�'ւ}�i��d�O���^
����t�;nn�ȕ�F�ZT����I�\�=�'���ORi�$O�!�D{��#���ɶ3O��O��lZ�{��c�\��?m��ʚ�P��x����?t���"&?!�\�����<���'�?Y���;j|�G_4[��	��k��?yf���C}�]�'$�����p�|�'�!W&Fɹ#�� F���u��YJ2�'S"�'���W�4Y�4K\��dX���53wb��>~0%�@M
�?��  �����I}"kf���j��ۈ!��9:��({l@�����E���TJ�nZ�<��k#p$��h����'-2�z�Ԭ�^4�97F~��'��I����	Ο�����D��T��!�'Vv���/��~�*co�[,�6�Q�S��D�O���#�	�O��lz�Q�4��4 �� �^��Hh����M�2�iɧ�O֭�P�i:�W�t�(4RuI�m��(�#� ��C�h�����	>0�O���|r��Q�=Fmݘ�:mЈ��X,:��?���?�)O�Ynڲf�4��	͟<�I+T��9d�D�֬����3;��?	V���4A����|�?cT��8��\���(�@�����9=��*�% s1�ؐJ��h���u�HIQ�Q�]�ѧb�t���D�Oh���O@��+�'�?aI��>����1�G��Ɉ���?i��im:����'2"�rӖ��5��}���S!*��!3�E��r�ɧ�M+0�i	��G�s������������_�4��QT��r�r��J��a�l�%�������'T��''��'��5#� ��Hde��!*,ܡ��[����4��ey���?����'�?��Î�C�j�S7 �u�<`SH �[8����M[T�iaɧ�O�Qpc�G�?h��k�A��2cؙ�u�B�%�~8��OҰ� ��?ɕ+-��<)�Ė�L����O
`���k��X�?9���?���?�'��$��9�"��ٟ��-�  $D H���z���Q���:�4��' �r��"dӞim4�:��ѧB�~�Fm��� .-zX��ƦM�'�����?�������� �i��닖�`�;����;�BD�A0O���O��$�O����OV�?��tHY�cs�ԓ���x���(�o^����I��p��4�p�ϧ�?�R�i�'V`X
�N�-5�@�
(mZe��e&�dn�~�n�?��ᦝϓ6��y���9,�L;�'W����&3��a+���O@%�J<��V�D��Ο��	՟�R7!̑8'�d �戝B���4�����Ay��{Ӝ����O�D�Ol�';% �a�M�!^�&e@eY�H�X�'D�X�f�d�u'��Mm��[�uYf�y�L���DH��K�F_�D8�EE��y�ȅĺCBoӖ�?�Q�1}Zc�Jq#Fd@-?<�ŢUƘ����	�'_b�'D���O^�	��M����*`g�b�D8+.]�A�ņ	����?�Ʋi:�O���'�7�M�\м�����+d �H�j�bb�m���Mӷ���Mk�O��K�̗����j�<鄉&� ���E�kȲy���@�<a(O����O���O����O�'1�J�a\X��% ��N�mb!�	*�ƠϨ���'N�����'�"6=�D���Q
qp�۲���!���A�C����S�4����O����v�i��$M���0��:A�ۥ�ׂ�~�/��=�9��(��'�	��T�I�Xxa�Rv72,:#���Dd����؟������'T�7�R�9h���O��d�bw��bs��
`��N)���-Ot�do�l&�`[�JW$Hrs�
^a�IP@�2?1���;F������'B��Δ�?�u�V d¬����!&��C͵�?���?���?	����O��r�Jv

���%\$%�XX1�O�lZ97��	ҟ�8ߴ���yG	ڶJx)1rNЕz�[7����y�w��n��M�����M��O6̡��I�V�69�i`#k��=��"
xy2�O���?1���?����?y�f�`�{1�ٍ�n�I6,V
B���.O
0oZ�P�I�����N����Xх��4"�0J��m��sp 
&����ڦ1��4r���OZ
����	���+dF��V�Գ4���&Ȟ4
�_�Dy��R�BB)�o�IsyR
I�**!�b��&��Pr�F4���'�B�'��O剠�M�w/E�?W�S�y�$l�P�P���?�2�i��O�і'�i�7�o.2="Em�$TZ��<L�1�Bu�$� �4�d��zQ�I~B�;Ӹ|��f�%�6��\�n�1��?���?!��?I����O��ђ�/\#3��rf(_';��-��X���ɬ�M#A���|���N@��|2�޲&�
ե�=[��8�/A��O~�m��M�'`� iK�4���X�iL��p4�Ê�~)!L�C��;u��?!��?��<���?A��?�*ʲD:X�$f�7Vz���bX!�?�����$ۦ1SAǟ,�	ɟX�O_T���W��깈�����Zȉ�O���'T\6�_ʦ%�M<�O�̺`J�'w��12���1��*��� \z�i>H'�'�	%��"1"���2���;��i�$��ߟ0��ş����b>u�'r�6��."�L�V!!SΰU(�Gڰ9�H��0B�O �D�ĦQ�?�VQ����4I �(��H��a�l��h��%�D�i�7�BB��6Mv�H�G�.G��tk��O|�@��?1�V��h� ���e��\�Bb�O���'u��'"�'���'�.(nHȵ%�Y{�1��	�;��9��49{>�����?A����?Q��y�Y��yG��3r���`M�1�7�K��q�N<ͧ��' d��9ߴ�y��
��xU/Q�omB�)B���y���W���I�"u�'��	ݟ4�I)6n�0�sD�:A���S�Ɖ2����I̟���ϟ��'h6��b�z�$�Oj���!7���V�>��(�ۧ&N��D �Df}"fmӠioځ��Q���*[6JFDĲ!��c���ϓ�?)eD,K�T�����D�� �2��p6�d_�_�Z�Rt��*�����cӒa.���O���OX��<ڧ�?����p�δJ�æ�(��ф�?���i�&i�$�'`��kӮ��_��A���q@>��%����	��M��i�z7�] �6m%?1�KK9��	R;c�`%ے�I<ᄔ)N�L�;L>i(O�d�O���O
���O��@��OB0j��0�3(h�s�
�<�i��Hq�'��'��O�R&ɍ[=p=°�	�+��9K���H˜�M�&�~�(%�b>��sfY*�ҍ�`���nD�S�^�Tl��"��hybO/{�Z��ɾ��'��	3�(�O�::f�3���Y���Iɟ�����H�i>�'�H6MԜb���!Bƚ1��K"K����*X�����Ҧ��?	�T��ߴPa�֤pӒ����փ��59��>R@�d�/:�7�/?qѹ+�&���.�䧠�k#b��=kh%���8C�¸h�n�<���?����?���?i��4�,g��)qA�da��"���5rP"�'Rq�4��T>���$�æ]%�4ـEK V���iV�wOP���.E�ēr�V�g��i�� ]t7�.?Q�ȖVkθ��ߎ����*��D�h���f�O��K>�-O����O(��O:)1�`�x�N��7� <�p�x��O����<q0�iP	x��'8��'<�S�G�ЅȦŎ`ԉb��y��j�	#�M�ĸi)�O�'`�"�;Ǩ!N������=R1�l�	��~ d宏��i>����'�B�'���b�)9ꥳƢ5	��������I�����Οb>��'�66�0'��pB"�	a�|�k�_x�	P���O��d榝�?i�Y��3�4L����y ��ϙ)_�d�q�i�|7-�&^<6,?��A�v��)��� �q�8c��D
A-�Yr:�6O���?���?����?)���	�"^�Isl��9ۨ��ߨT���K޴8�Z���?Q��䧪?A��y瀆m׎PA�/��^"�a#"��2�n6�ѦٓM<�|�Pi���M�'a�B��y����w��XB�'���'A��D{7�|2Q���I֟�y�C�Dr2��'��\�ԽI��џT��ş��Sy2by�Dir���O����O ({��j��1���	;�hbf"��������4|$�'��Y�Ԇr��\�� �_��yӟ'�H](7�N*K�z���\4��X?Yw#M5�u��O�Q
p×�Q$����G߁W�l�!`�O����O\���O�}��d��؊�N���t(r�^?c���������AB�'f�7�$�i���〚#
�x�l��?t�	1fo��ٴK�V�o��H�@pӂ�I�p�Ch��u����LY�{���:[����^�~.�$���';b�'m�'���'��ٷ&R#e�8  ��2s�f!�R��ڴ_x�����?9����'�?�F��R�����BLX 
�ké�8c�I>�M� �ie<O����)Q yؙi�D�$!r}{P���X��<���L��	�Y$�'��'���'r�p�e�|�X�e�(�̡��'B�'�����U���ߴ#���������f%�h�!��(�'n���?Q�6��U}��q�T}l��MÇ��j����e�Iؐ=bA#.$��5�ܴ�y��'ht����?Uy�O$����V��L��S�)�Ǯ$	�.A�:O����O���O���OH�?B�a�Yk�o��c�"}�`��������(ܴw�"X�'�?���i�'�����U��]rb�D[�II$�!�\ڦm���|2���=�MC�O>=p*��0��p�F
I�+�@��r�F�t��Y��g���O���|:���?y�XKޠ� ��	�͏�uG�t����?�)O�lZ�3R��͟L��x��)���1@dD^�pt���II>��]}}��i�4Tm�1�?�O|z��H<xs�$ θ�2�݅Yp�<Q�d���r+�����d쟶����'8����`�%X�0}aM��2��E���'!�'�b���O���MB9?,��ʎ � eaģ�+�#?9w�i��O� �'N^6��	hx���'ӿh� �b��\C
�m�M�#��M��'O⃝�?��u��+$剛'd���AA3MG���'
�&��	hyb�'�R�'�r�'q�_>I��ÑGˎ蚥+� P\��E��M���<	��?�J~ΓF���wےH�0oP�`U:� Y;	�س�Ai�f�l,�?I�O������IH-w�6n��8h��	V̪�&Ǿ-"���s��H@Oż8b����<i��?y�IU7y��2+E	Vn�dsa�A��?���?Y����dP����V�d����0(Re�"~�x`@0"Љ9���ņA�t���*�M���i,����>���I<x��"�g�T0+�.��<���~,8��	����+O���&�?��'�h\���U�Y+Ʊ �
�b�DB��'���'�B�'��>1�I�o	N��ɯv,�y��gK"� ��3�M�3�w~�{Ӗ��ݳE]��3w怀z㮡����-��.�M��i�(7��G`7-p���:J���3�O~�� ��̢2����HZ.KDp���8��[y2�'���'w2�'+�/G1L8�a"�[���[��	��Mkq��<���?!I~�8�J�RRF/nU�P�;��-8����M�f�i|��;�'!����N F�MJ����t|X��͍*��)O��2k�7�?��{R^�����.b�n��aS�d1{
�Ɵ���Ο������iy��iӜ��8O�L	��<붨�%IM	*�����6O�o�T��R��Iȟ�nZ��MK7�/���E�0�V�Շ.C� �۴���V�`e^����V��މ��I!��2��ր9u���� a�μ͓�?I��?���?����O_~�kX�P����V*t����'���'(�7M�~���M[I>yG-�J�Z(�N_�U��<{� F#r��[���ܴ'��O	�%zбi���9jtZ��͟�G$�,Lc�\�pՠ�"0��� ��Xy��'�b�'D�,�=3��wg�
7耫�C�M���'X�	�M{� י�?���?�)�b1�У�N�椳D�U�<��]�×�ts�OLnZ�M�0�'ﱟ��&�T�+�i��oY,I��y1f�� C�L#$E�69��|�cM�O(�PN>!�rSj�u䈊O?������?����?���?�|b,O�xm���3.�v��a���C)�0k��M@y�mi���a*O�6-͈��B�S�>��}`w�^�iҜ�I�)z����'Ja����?��[�|ppj�mL�=p둃~��k�p�'��'#B�'3r�'�哿Q�4���'E�.��h"�]v� ߴ��H��?!���'�?	ջ�yW��85��X�(*<�H���cϱ*E�7�R���&�b>�R�HݦMΓ
�&Ի�J�a ��D%͓H;����D�OX	K>�(O��D�O�t���ɥ4�$݀�DO5�qx���O����O:��<yS�i�PX��'���'��E ���?���T�J�i�c�ċby�'K��x�	��;��$F��8Q�D�^�y��'<���C��.@���`]���S�0��������3z�.-*��Ȳw��) G䟜�I럈�I؟|F��w;���w��6[�^Q 2��3r�Sg�'W.7MF-A��$�O*AoZT�ӼK�]�'LP��ר��1l���m^�<y��i�7-�ۦ��P��=�'i��0�/[�?�K
� p��[Vy�  ����:��>���<����?����?���?y6�	%e�"�У�R�v�R{'S��	��s��Ryr�'x�xJ�Ǟ�7]HE��m�Q̄���E�a}B�b�&�m0�?1��X%2#ᰃ� �8��ΠS�<�:ӏ	4���<��y��+�O�kM>�)O�T�Ta�2<K8��/�/{�z����O����Ot���O�ɸ<aԿi����w�'��T��+A-x$��Bw�'/r	b��'6-$�	���D�Ox7�Yݦ�+6*��[T =��hŴ0yH�P"H��zI^�m�Q~2C�7Ђ���@C�O���ػi�X�	��
�$��G%B4In���ݟ��	��(�I����	A�'.�R=�A�A�G"�F�������?y�kf�ƀť��D�'-`7�:��U/�B��q���uf�C:�\+��xb�~��lz>!�NE¦��'�zr��M-Cd��U��e�x�D��w��|�	�\4�'��i>i���t���$��=�P�P������i���������' 7�Ь~����O��D�|��@��;��	�E�o��;a�[~�h�>9D�i�6�AN�)Z6O�Z��X��!�`E��
g#�Ukȗ?!D$�����H6�|LS.rJ����g��\�2/�'���'���'���dX���޴9�@�B���+6tkd�ӛg�iZ����?�������$�a}��cӪ�0�kݠ~����6l*ni���Hɦiܴl�=��4�yR�'�%t,��?yp�O����$|pnL�t���~l,!�$<O���?i���?A���?����	S�bxQAڿo��0s�E�1"�\�mZ"R]�M�I؟X�	d��؟�����V�^�H/�E{�b�A\�8R����iٴ-�����O�D�@,��6:Oj��		YB2�G�.-1LZ�4O��1�� �?q�!��<�'�?tc�
kg�W�x�� �̉�zD��������I�(�'�J6�ӧ}c��Ov�$����@���6^v�(pD#br�[�OPlZ�M���'��I u5̤�eկF���b�b5�z���j��%f*QQ�o@y��OՐI��v?��	�?A�|�HH�e�Xa���?����?���?����OP��#��*��L��X�rT��!�O�IoZVٜ9��ΟJ�4���yGE����L9���۱<���Q��O6M�Ӧ�3޴"��iش�yb�'،�4N�C���QoX�����˷ ��9˄�H��䓢��O.���O�d�O���[5n �pp��(-`B!�����}���=����ˏ] ��'pҔ��'��ba�̦&��!C�J�TC�u ���>��i4�6�{�i>����?�*��,�#Bӽ}��d�2�@�<u��0	��I�'Ҭ���P?�L>A.O�qa�^�5D @���jd@����O��O���O�	�<���i�`��'�>E����@9���I�R����'�67�8�	��$�ӦIH�4N��&�W=36M`��Hb#��K�"Ï\ôTS��iJ�I��r-��ӟb�����B����"�in-�V*ɷ:��D�O���O ���Of�D?��G9굂硜�{�dQ��*�U��	�L��8�M[�E�|r�z�&�|ҫ˾C��hiQM	YK����K���O��h��̶nu7�.?��%�!!_.�:cK��f���Ҥ$E6�`���e��&�l�'���'-��'�=��ӶCG�����^<̓c�'bV����4����+On��|�D�U�d-z�Y�OL�( aE,�@~R �>aS�iW�6MK�)j���n �� ��0DP�(x���$ު])wGș�M3 \��>;F�$1��T5��,صb�2�Y��BC/a��d�O��D�Op��<�4�i3d�����7$��	I�M��҈q��?X�'z�6�:�	5���l��1j��|5�(��@!F��牜���۴l�
��ڴ��W�50��O����l��� DT����8Y�V��Wy��'��'�'�\>y2�+Z�^&x�81�ϭr&PX��*�M��.I�?����?�����u��Ƅ\�b�9&�=%
P��҉�/x�HlZ�M�w�x����ޏQ;�6=O�!�D㜜#�F�[� �x��� �6O�ɩ$���~��|�S�$�������K  v�m����*�4-�'"ǟ �Iߟ��I{ybGh��`�w��T�ɚm�jP�VL�������"im8��?)Q]�Ј�4."�6��O��!�X���m�<�jI� kk 	͓�?alL/.Sf���f�����8\���~�D��?�D`���]�P`���J��']2�'m�Sӟ��'���s�& ��ә1M����ڟ�)�4|�8|�'��7�/�iށI��R�5��)%g�+������ym�֙n)�M��Q��M��OZ��T)2�RTI�EJ���Ʊ �R�b���1O^ʓ�?����?���?9��g7��ؠi���-�7)�"���	/O@�nگ~��	��H��G�s� S%IE!;ab�J5�S�&�aȈ���D��eq�4%�铿?�D�����i%�\�SG��=i�\���F0:ɠ��'�P�smɟ��=�.O|���(BH�ak H�l`���!a�O����O���O�I�<�g�i,$���'O����E�x(|E+��@Z�jȟ'�^6�%����������4"ʛ�i�!N�����-�&��F�w�,`Ըi��	d�ys��O
n('?yR[cP ؅Ł7ڝ�1靤Z�~�')��'�2�'r�'S��	 �C�3�0tY����u�?O4�$�O�mZ�Y��[Z�&�|R�P�Ih�M��,�?���غq����>���i��7����@Ғ�uӖ����#D2� ��3�#J�)� �CEW�@&����8�?��{b[�8������꟔��a�#��#�(��b�xճ�DٟL��oy2�j�@�"4O~�d�O�˧>������^�ĒG'�).�'��6��A}�(l��x�S�?y��� Wkx��;J���� ��:s<��4d�(����'*�d��ӟ��=i�fʵAm���L�"�6�ꗤ�?	��?a��?�|z(O��lZ�L�|�˗n&i?���e-�l��$���'?9��iL�OR��'��7MS�X���G�6�Fp�6T1YKr�2�lZ�,NmZ�<��;��!�$��-Oީq"cż���p�!�G��L�3OZ��?����?����?�����ֻ|N,��Xwe�8"�R��E	Ժi�=��'B��'���y��~��nQ: �9"H�1 �l�����W��m��M��'Z�i>=��?5�S��ަm̓&�PY�Ӄ��u؞p�Q���x<N�9=��@�m�O^➴�'�B�'��2�B1:�)H ���u��7�'���'S�0�ڴ&� ���?���Ȁ'�K-����'d�?Io\(;���> �i�
7�P�1f���\� ��9�FHT�3C��tA�����rg���|jQ��O����NZL�CI��&��;�F��3������?����?���h�F��H2��!�bŪm��R$��2��$���͂�J�����	:�M���w(����pTJ�z�Z�4�D��'Nj6��ɦM�޴G����4��Ě�vi4��'¶}p�AS��J�T˅2`��dD;���<ͧ�?���?���?I��V�F�d� JO�q�pla���&����-��D����I��|$?��	�#@�a&����-�Ф�52)�(On��bӼ�$����p�$�R'��D��;+�8Uq��[/��u" ��d���߰
T_�qy��@X8 ��%/p�p �'�N�3A��'d��'��OF�I.�M��H��?���7kʒ%��
�b[&<�fD�?�Ӽi��O�)�'�6mLۦi��4<00I�܉7��H[c��w*T��%����M�O֩�T+������w���3��ʢT6�d�5�(��	!�'��'XR�'�2�'�ؕٶN�!SY�ıH�)MIN�@���Or�$�OЕo�;b6��Ο��4�?y/O�Ӌ�>B�A������Z�h�y≗�M�7�i3�t�:���:O~��N�j��<#��
H#(����&w��i'a�2�?!4�2�Ĭ<ͧ�?i���?� YF��T3�F��(���?����ަ����X�I���Ok`@�Š�d)�����' ��O
��'�6m�̦�iI<�Oܘ�I�������&��𖍙��NIˠh���4�t����X�OM����p�d��V�)4�bM���O,���O��d�O1��˓[ћcF��C��	S.��#�Ϝ N� �'���k�㟌�*OB7�)�ڙ�fi.D�X�Ǫ�%_�:�nڻ�M+JҼ�MS�OΕBDi/�B�*�<9t�_3jXPɘ��^�[%�H��j��<�.Ol�D�O,�D�O�d�O�ʧ=��	��Ђ6����u��(��5j�i��8S��'���'~�O���~��n��N��9z��_�F1@̚�IN�i��Mn��M�'�'��i>����?�j�]Ǧ͓,{�4{C��GF����#N<Y̓3TF�� ��O�9�N>�(O����OVH@�] d�|�8�&[������O��D�O��$�<mx�t�J��O��D�O�}R�$�G'n�a%�#z]¶ =�		��$�̦]J۴!�Y��b�S�(T$�f"
�N�VH��g�6�i̠���
~tRH��T��S�5&����l��H�
�vq���=h��@r�]ݟ���̟���ʟ8E��w�82��Ä ���4[�:hC��'d�7m4G>(˓Tp���4�&�	���7G�����ۂY��)�P=O�oډ�Mㆰi����%�i��	5�8�s��O�4(·-M��J���BO�<O�q�j�q�	Dyb�'l��']��'���b�Ĵ
1��,~b���J�/J�I��M��D��?y���?	L~j��V����'�-al��!eV�},��Q���4P�6�/��i�3>��qH��bl�vȗ�s$��WaV/A��.�� ���' ��%�,�'l h�!G�:�8��BR,^��7�'-b�'2��TP���޴k���C��O[���$X4�
��`	�+�*��Otm�N�JB�I��M�F�i��6�)��Q��b��%��8O�Μ��T�p�����;���?
\����e�S��5�cY.o�GH z��["�yr�'J�1��G��F%x��'�ƙD�$tq��'z��'��6-�	O�Ӣ�M�M>k�(BmGä*��!� �@��R�ԙ�4"��O�>�*��iU���XG`�	t+E�c�F���g]9I���a��B��oj�IWy��'���'xbLN�<n��3��J�m�:�*c�	7 ���' �	�M[ n��?	��?9(��A�LH73>�h�F��Da
����,�Oʐl��M��'ܱ��D`���}5�0�@Ÿb��qg�Lh���ʔ�#^����|�b��OD1[I>�)׹i��G�/",�l�d�Ԁ�?A��?����?�|(Ojxo��-V����O8J*�ã�`7@
"	������M���,�>11�iM���@NN�` %��*^'q��$���y���m�@�F�mI~�N�`9 �Sb��V��䈥('H�&�I�mW#B��D�<���?����?���?�,���j��2D�L2���Z{^(�����}�B�џ@��ȟ�%?I�I��MϻD|r�kAA�ZJ��Ц� J2J��i�"6�Vҟ�է�O����C�iG�� ,xPǫ�#ch�� �ȥ5��<�1<O:9��:�?�S ���<	���?I.�&W��j #�
}�~I��S(�?q��?�����KŦ��IE�� ��۟ذ����fsH�$ma�~hb�L�zE��'�M�D�iB����>�U'ʜ+8bm�w��u�m�E~���;쐔-f�
E�O~:�d�O6E���pd�1����F����A�[>��B���?)��?����h����M�|(�R� �1m;ġ�r�K+����񦥘BI���|�	0�M��w�HXҠ��gv�@�;�\�p�'��7��Ϧ�޴.�v0C�4���	7X����'D���t�����)� T�eV�]CR�2�d�<����?I���?���?�J�(G��q���n.A��I���ĈڦQ�2)˟,�I��%?�ɷT��ث螁f�D�q���$A8��q-O��D�O�O�O��H*PE2EԵ�jL�h�C�ݷ;/�qc2U��a� u����F�	`y¯ۀo���N�5�j���N׆2�2�'���'��O��ɻ�M����?���AI}���� �NX�c`��<���i!�O2��'��7-����o��8(�솆d+�����ie6��E��ϓ�?I0����	�����<�n��.�L��e�jM:��l��d$�D�O��d�O����OH��?���X��☁L�8 �%-����	۟4���M��`P������	Dy��Ƙf�Ts ����["�=4(lO�mZ��M��' cy�۴�y"�'.jL�;n�|�yӢk1��'ˢ|	���'0	'��'�"�'�"�'JdS���v�^I���:M4�:��'�_����4's������?�����'c�m�p`z��AGaL�\|�1�'Z���f��OO����y`�B�����)nrP+'��_DTa��?7����1E�O��M>(�)Bh9�a�%A9F��"
��?Y���?���?�|-O�	oZ�8���C7�B�I�X�ɡOրU9;�jO}y��g���ɩO��l/�by���ނe��#��
N5�u��4k7��C�3���6O���5�*4�'
��ʓS���0ѯ¯H�4�Y���l��4ϓ��D�O��$�Oh���O���|��D�H?Hd�.�4n�ݫ����u���^��'�����'[\7=�:�C� g=P��̕	��ݠ�����4(�����Oa��+6u���2O�\�"i�/F�L�b�!C�{D�M�0O,���W/�?G�;��<ͧ�?6˜-�t�õ�ܛ���(`9�?���?I�������H��MCyr�'�" ʱ`�]t\I;���,4��Q��DSX}��n�h�n�?�O�Y(@��h���w��vҵ�R7OZ�d�UU�mX�$M#�6˓����O�̲��,b����8XF�����C`��b��?)��?I��h���D_�Q"���ɹ3/����!�*d����Ѧ���QyB�e�N��
'��x��,8!���
��	?�M�õiN6����V7�s���	�0t����O9��i�▮p��Ek��$;AR-�r'�K�Idy��'���'�"�':�EJ�G�r��PE+�m�� p���M[�R$�?���?1K~��O:y��g����u7̟9���Q�T#�4�g�O6�v�i�����U"MJH�`�h6(^�	X$"�-�<IP R np2�DS6����DLa��˵�A/@��s�撈t�����O��D�O��4���:����'la�I={G�a8��I�c����K�!`�R�{���,��O�Qo'�M��iXт�����k��9"�����O,<����ĳ��C�C���I��*D���_�}����s
��V�l(�;O��$�O����On���O��?"4���P�Q��!l�kG�U�����ӟ�	ش,� �Χ�?Yײir�'�H�2�D<e�(�S �������$��������?�A�O����'�H@1�cAx���&8b������F"����/U�'$�	՟��՟l��8�~xâDB7B����f��BC���I��T�'D�7m��a>��O��D�|�$���siF!:G�7���V��g~�d�>�a�iy"7��ڟ��~z5�Ld��U�6�TX�R�F#S3� ��Gu�k+O�į�?1�{��U�D�G�ϣ`�
�Z�M�J8��'d�'����Y�8)��7���A�w��a�C�"io0��n(?��i��O���'6mЋI�Xp�R�0l�R����J�M�ưl�	�M��ײ�M��O\x1ElI1�����<�l�>k,|P���co|������<�(O��D�O����O����O�ʧ�(�K�'� 3�L����=y��Z�i�$T�'1��';��y��o��.
�g����U�2a4m��'15"W��śF��O4�S�'��Ѱݴ�y�O(�b�j��+x��y�]0�y2(v����I���$�O:�d�3[wH�[@M�t�����b�T�$�O����O�ʓ[�����)mK��ɟd[����w�b�[0q��b��Vu������M3G�i7��D�>�v�1g�91E(^3$d����F]~�P�gW����I�Y��O|���ɍY�2.L(�tU"�:1�d+�$!�b�'6R�'��������5D���a�K�y��u��I ܟ�S�4�@q���?�&�i��O��9Z��@�*M�N�&�p�Q���Ȧ�8ܴH�&�����f��d`�B�P7��
��s�D-��"Ȋ��ܓ~�|'��'���'���'v��'2��`+�$Hl`%LDDP��7R����4-�f� ���?�����<�!�=o�d#c� �{_$�z�c��	��M���i-z��"�'o���� v�;�J� 5�X2"�?{����R-ֺ,8ʓO�Tm����O�|�J>�/O����մ{�t�H���+r���s��O|�d�O���O�ɰ<�վi�P��6�'s��K�H��������m����'-z6M2�� ����¦��ߴ8���s&.�J� �1���i7@	_�xzԺi���%LxAb��O��%?�J[cuz��%S<+�l��I3�|1˘'X��'���'M��'��V�zAͩ$�t��Ī��*3�,x���O����Oj�l4L!�۟P�۴��.���IlO�6H�B�c�4��2�'���6�M3"���h��F��T�7��e�bPaY�eS�݉�"ÛP��p&�'�A%���'QB�'R2�'����`�_-r@�� �i��M�'�R�'z�	;�M������?����?�.�d ���9K����4쐚7r�]�b����O�Xn���M#q�xʟ��' ���Ć�=N� �g�M�@ITB~�TQ����k
a?�J>ٵg�#w�Ve2˃0d�:�p�/��?���?��?�|�.O�lZ� K��r�P)q��>04�c�qy�.}���q�O�m�4U�k3�L%9�,%�ᄂ'o�RyJ۴bl�V�U�UG�&�� c��9��ɺ<qD�ĉ&��pS��H,�ı&��<I*ON���Oj�D�O����O˧[�tP�
-G��$Đ�~D 4�iWnDK��'�B�'��O�2�`��n��?�8Ѫ�>��8a%�,�6�o��M#t�x��܌F>7mk�����R(,�f/�[+L���Do��A��k��%��<I���?�#��,� MK�m,�z�ᨒ�?���?)�����-s�*V���IП�£'�6{�,���B�'b�=R�h�������M{��i��O"�
��J+�v�pE�P"X$4*`���h��T0i�dn���'n���	��Y�&�:'�2EKpa^d6HaF�ٟ\�I����ş8E��'7��k���6�6E�WB�q�B�`��'܌7�3_�B���O2im�w�Ӽ�g�T�p�(�gl�K��X�M��<	E�i��7������ڦM�'�hٲF �O�u�T;!�v`��J�j�8+Ѭ%����d�O*�D�O���OH�ɛC�­P����S4N��q�O2�ʓY ���P+~b�'����t�'���E
�ʬ�@�^�#"Ȥ�S��>p�i$�7M�Y�)�S{�M8�������5b �9˞�jC�M�Sr�s�<���O�ZN>-O`u�(FGH1R�n��-�4qr���O���O����O�)�<Yǲi� �B�'[�e�C��ɚ��ƴx�MB��?9�i��OR�'�@6���m9ߴ)�|��߫o:t}�@��u'I�MK�O(d��b���j2�	J��"CU�0T��+~��h�֪�<���?���?����?���dg����`&fT(��4[���:~r"�'o��e�ڹ#�O�tӴ�O�k1�ˊf�� �+�v*���u�Y��'�7����S�I�el^~R�X�p>�0�E��>7�"$y�M�,hX3Q��П�sß|bQ������I�J��asd�Rb��
zN��5a��� ��~y2���h���O����O�˧DX�%rfE�'����%e�u����'�D�E����kӄ���h�'r�����7�2�@�E%5b�`G��N~���� ���4�l�����8�O���0��"�R`�0mȇc�R����O.���O,�D�O1��ʓ9����</^0xj"�tP Pɔ�r&�Kî���d�䦁�?iPY�$Bߴn�2�#���>*:y�ӫ#�Bq�!�i`b7��`��7M)?A�*.&�i#��DF4�p���/%�@�c3gA%&�<	���?���?���?1*�$����@F�D����_2�;��ۦi�D�H۟\�	şT$?U��-�M�;L�<E�sdV:���5�ǊQ�Ұ�`�i��6�����ק�OL�x�C�i��d	�NI�A�q�KQ����A-:F��40e�0`��T.�O���?��M@�h��ۘaL-pWL��1�(J���?a��?i*O.�l:����ӟ �IO�f�R⎇8b��MH#���,P�?IR�LZ�4aś-��"D)25�W�c��5� ŜG�I��0��]�O~�p@����ɳTcTP1�1$�x��dB|C䉪���Aeѹ@�ȤSf�fZv���&�M;q�\��?q����4�^�!�a[#3��#�傸|QL���O��|�(�oZ�a���mw~a܊(?�m�'B~�OC1wќٰBc�:Ef�9jN>�*O��?��e[�7� ������܈B��_~"�o�F9Qd��O �D�O~�?}��dI�AP�0�Cğ�bh.D��,Q����ܦ9޴)�R�S�W'&`(�lUa`@���[�_M����.N�2��Ĕ'Q~E�!_��4k×|�Q�D��JF{T(���ڹW$�(KSk����I���I��SKy"�}�RL&L�O�0k$����Ȣ,��G
2Lp��O4�o�W���I�M��iN�7�X'�=�F*[�H���St�^�_�����d���y��3EF����>���=b(Չ�*�0�*���Cr���	ݟ���ş��	����	E����aIYq��L*& ������?Y�}@��Fۨ������'���_(W�v��bț8y���YVl��?y-O���y��ݝNf7#?���F?��t�A	�����	�C�,�S�OZ�ȕ'��'�r�'�H�9U
D�EJ��1�T�*�����'��W�h+�4]�L����?q����)N-R��I���=*����i�M#��9��dV��ł�4o���� ���G+� Ȋ���z:�Z���U~���A���G:���|Ӈ�O"�H>�d��fP�䫜
G����	���?9���?���?�|�.O�(l��5�d�A����K���c��L5�F��WoVXydqӾ㟸c�O��oZ^-�x����z�8 4oޫ/vu��4.��vI�� ��V��P���x���n�xy���t��+V�E%�����*��y�Y������X������t�O����V( v msA��rS�ع�jfӢ�xD�OL���O*���_ئ�TLj����S���IP���7�hi���M�R�'�)��K._�Z7�r��+3��Ya��a2HH&"h�5��|�\����$�bp��Uy�'�N85�5h3�)O�b��$ͭs�r�'{b�'v�I0�M;1'�'���O  r�
F	O��!�DC����, �I��Ȧ��46RP�� V�݈jВA:rəIl8�� ?�td�`�L��S���'u��P0�?ʹQ����BF�����F���?����?����?Ɏ�)�OpT�ax�	���hUX֨ �1�f�D^���{��lybIb����Gz� �TDZ	D,[g'���	 �M�d�'�F��t𛖘�4Cg(�����q�����l܅�ҷ6���7��$���'/B�'0�']��'{�$9�m��~�p�H�mQ�A&���U���۴	��?������<�͞?%@$*�L�f�2��gll��I��MkѼi����:�'Z�ܢFˋ*�Z�ae� � ����4����(O� �&%�?�B�*�D�<��	���N���τ42��	$-���?q��?Q���?�'��ܦ�2��ݟ�)v �B�2P0�� A��d�m�|�4��'�
�P���o��o��踹���	<q���È&c���*��!�'���rb��?�q��Kf���S�Y�4w���E��P	��A&}�@��I�7�T��!��:yN���L邅�I韈����M{��p�Td`�0�O(1�BQ/S��������Rc≇�M+����$��'N�f��Dbͅ�Fs�i�%�ˑ1Q��S�;U�L�bt�O�On˓��'_ܼSd���g�%��*�	L�@Dь�ئ��j�����	韀�O8H�g#�	�4�P��Ce�,��O�t�'%�6O�ѐ���O���2!\�Vݲ��G�ܔ�ɠ��+�"�Jf&s��i>Q���'b��'�l�ve̐hnP�3'��4��XRHS�p����L�	ɟb>)�'�,7�|u�wǬ bd��3.x���E�Ot�$R����?�a_�T	ݴ5��+���<�R���$�8v�[��i�6mZFX(7�0?y�'H<�N�����d�5D��@«A�7$ 5ó�Y9 ���<����?���?���?�.������'6���@�g9��KDj_��	Y ����	ҟ<'?��:�Mϻ���%�w�|uN�>]p@���i|�6�]䟘ק�O��cױiV��
6|i�9�C�K0*��/�$HU���F�0p���O�ʓ�?Y��xb���%ܗs �:���^Ű���?9��?�,Ohil�D�Vy�	�p�	Qe��+�(%JKD���.��~����?�_�t �4:��N�O��?@���V�y0�TjE� ��8u�'�`h���V�G�*	�0��DE�ڟp���'�51�'���HB��n�"}1��'B�'��'��>��I3`�XQd��#Y qPԬK	�`�	�M���@`~�/l����݅*0�-t�G�D� p��>���ɺ�M�R�i7M�^;|7�!?���_8�i²wp^�s�gO5s�F�"d��
A%,�`y��'���'�b�'�f�#̈́)�qk��`֞$�5��I�I��MS�B�<Q��?�M~Γ1Bmz!c�<0E$]�R͎�K	�5k�Q��I��qZ���H��E2t.ET@LIc�(f��ҰO��/��Yd�<��>��5�	Cy�97Mr݈���0��j�]�R�'�2�'��O�I��M��e��<�C�͹X �t��l��n��\
�d��<�p�iq�Op�']H7-�Ӧ��4w���dK�B:�PeO�d��&��M;�OZ { U���L ��]�k7 C��0Lh$D�$�2U�쳟��I�L������ߟX�
EhZ��s���=�����o�J��O,����Uc�M^hy2�b���O�yд��F���v 3 艘R�\G�	�M�c�24��'�M�O�yP�Mٍ:2�X¢�#o�ܴY�@�Ԭ�,�M�$���<)���?����?	5&�)X��=�QiZ�b��ŃӮ�?����$�ߦE�Q����������O�|���?�dͳ2���\��%8�O���'Ϛ7��$��'(F(X���$&�j��w��,$ׂ�b��%V8\i'+����4�`����Zf�O�yҕc3q��I`G�ږE��@$��O��$�O�D�O1�*˓aܛ���-n_<����	)#0��X4AS��@��U�T
�4��';��x����G� '��X�`H!@��K��z��oӌ��tdw�4��-�Pd��q�/O����qI��S�@�v�Y�>Onʓ�?���?����?9�����5 䄸Q�F�S�=C�C��o�Tn�2�Ҹ����	]�S�����Sǖ!W� ��7(���H�M\s��D�O^O1�Vyɤ�l��I�YM�ax���'�漓�$3��片g;(�J��'�(d'���'���'�9!�� V�\�s��xߺ1x��'T��'2\��!ڴ!{ځ����?!���ycʃ�Ui��� q�����ĵ>y'�i����=�� �U�P�� ip����
,~*�u���%&I*���8�*Pm�,��+��\��Ӫ
��e���BL���qV
�����I̟���ן4G��'в�	Ê �\\�4 c�//Xz��'��6��/=e����O�xo�f�Ӽ��/����ɜ-r:��vF?!��M��i��a0�i���8��!�"�O�X�Q�Q�*sfq��\��"!��]�Yy�O��'\r�'L��tЭbb�ګ水.a5�\r.O�Un��p�I�4��w�s����E���g �^1��!І���զ��ٴcP��S�%Y,Q2 � Y�FpIы��"� ��N>% �'���{����=�+O�X ��X�E\ ����Y���O����O��$�O��<��i�rD���'av�7��%9�ʸ��E(�!`#�'�f7M?����$�ʦ51�408�%T:��$��gN()����A��M�p{��iv�	?�z�)��OW`�$?M]c�Hz��L2XH�Y"H�.e��+�':�'���' 2�'Y�:(H�hM3m>yP�E�!�l � �O��D�O&LmZ>D���۟���4��2,��$��(D��h !��l$nY2�'#�	��M����T"� f<�Ɲ����U�o�bhY���Ve��oQ��Bោz��|�R� �I���ğP�&f� >������x`-0E������Hy҃|�D,a���O@���O�'[y�R䥋T�0�
V0aG��'�AA�f�o�u��a�'Ga�p:QᎦR���6�)S��t1�'N�������4�`�S��E8��O�M��eE��"��bӂ[�V��O�EnZ#W.`r֦D�3�2��Bk�/�4���<���MC�Ү�>i��i�D$O�լ�)E.�5���	��i���n��c�Imk~Bo��̮��'���Ȉn���E<p���a�W�)�D�<1�b�������$���լM��� �i���1��'}"�'&�j�oz�iC��L�*Pj�nϙ/2�����M���i�XO1����VHk��I.H�B�)��8<�� �K�6lHz�ɜ��ہ�O$�O�˓��D	bH���KЌ/C �I� ��:ax"	dӄ��!��O&�d�O��`�b=49���o��]�!�(������O�7mPu�ɍS@B�жI�� �p����^�������ӈ۶�M����$F^�S��$Z�j ꈓ����C!��y�ƒ5^rxLC�"�3o>�H�ա��9ZD�C��?B8�hS&⋳W	�h9cÙ#r*�,�G$�)[^��J��-�Q�Ɖ1�0q�p�#9b�\ UJ�/�>< ��5ΰj��΂]����شE���cRd��9�!�Ժ���FQ�eb��P��F2z!: .��GRl��g�����p�d"���X�dDT�I:�����rZ��{c(G+`+�0�3�]�r�L��UlU8}�*���.��(K�RdJw��;_*� ��U���B�GO:L�TiZvg$Q�v�4cAi[lyӊP�{ĐDn���b�=���?��������/ӌ<��A�������S'�u��?��������	ޟ�����q"ŀ>���EE�	d�듢�9= �I��$�	���	T�I����8F�>ȐP抑xՓ��K�EF.	���F�v�P��?����?9��?�g�%�?a�N�.��t�T�A�>jޗ�/dQ��4�?���?YI>����?��Q�u�Jm(%��L��V�H��0
�U	~H듖?	��?���?�$��I�O��f�,r%�*Fj�"D�8�$j��	�	v���ɨMmѪsG(�!w��!Ҡ{.�S �ԮUL���'W2�'B �@R�'6�	�?I�sπ3Y��l��)�1���[#�	��ē�?���l=fI���Fg�S�d �u�P=`��9BmL�y�����M���?Y���)�?Q��?Y����+Okl��!��P�q'��&�[v�F�,��&�'5��]�D40,3�y��tN���%�f��X��jՓ�M[�۲�?�����d���˓��D�k�����yw�D�peT�W���mZ+:q �`� 1�)�'�?Q���t�nh� nT�WE��ӓޕ8w���'��'bٳ��.����`����Af��G������-4}�>1��R[̓�?A���?	G�^4>���z�h��
(�t�.���'����/�>�*O<��;���@X�P$Ѝ4���5��n��t�R^�dH����',R�'�BT�0[� ����3k��e���ekU	^� �OV��?YO>����?���
�	��BJ�
j]���@�~ƒوI>A���?����O*ϧ~���m�&q��8v͟&��ElSy��'��'���'��j��O($yg�˃_'������6��RrR�<�	Пt��Ry�&E��맧?qg-D�b� c�Md���i�(O�O���'G�'���'V���'�A��Ų��L�!��X���NT:l������Xy�/�W2d맳?�����KH"���q��),��(Xg���'Y��'������'�'0���7�@q;GM��;B`�pd�tÛ�V�\��+[-�M���?1����sT�����c̊j5���mG�}n7��O���'-�����}j�&�C����U/Ι8v@�¦���!��M���?Y����cX���'x.�q'/�,V�����ǸB~����z�r\@É4�I|���?Y���2:oJ�ɰH�I0�1����4��&�'"�'R�TY*�>�(O��D���7�
�#Q��F��8����9��Fq�}&��IƟ���*�0�a3�īU��g��kU6�޴�?��3���py��'/���X�#�R!��c�L�����dזs����b2��k���I�8�'zN� ���P� h�H�
�kQ	j��m�/n��	yy2�'��'�"�',:h;����LI y�U"I�(�Zb�V�)x�'�b�'G�T����C����tA��$��͋T.�*8�D9qP$A�M�+OT��-�D�OV��܆*/|�	;>��a��dňT��b T��듈?y���?�,O� ���Q���'���֬�;����(����iӘ��0�$�O��DV�CF�㞰R�nˣt��H�F��T
�y�UOeӖ�$�O�ʓ
$h,;�U?����ӳ-5�$��+�x��
Tq��I<9���?�dné��',�i^�T���&+�*Y��LB�cG�0 ��Z�lX@���M�R?u���?���O���X(��4b�J׆0�:L�F�i�!X�4�	<�ħ����bN����PC��>�l+�JqӞ��Èۦe��������?�jK<ͧs�|a{��8d�����O*W}���i�>�pD�'��Z��%?��������\g69�L5���J�M��M���?��!��Z��x�O��O����r����r�L��F�i�B^��H�*�>��9O����O��D؊i����a̒3�$�j�J	��m�,�ࣜ����|Z����Ӻ����@ ��C�T]@���b�R}R��<U4�P����ڟt��By�L��<�j�RA���+�S�M�F���³�6��O��+���<&ˍRl����hȏW�`� A� �M4�H�����?)-O\���9�4��?N���w�3�P����
��7��O��D0�	ܟ�I*�
��`l�Vl��ɐ%ov^��t�Y�i"`���x��'��	�8)ւ_e���'�6��E�2S<8�0�!�'\�*����a�
㟴�	�4�P�8;a�O���T
Ҽ8K>JT�2(pn-�0�i�T�D��!XD~\�O�2�'V�\cr��T�@�Q��`� M�B 6̲O<	��?�u�F�+lT��<�ORXc�Ɨ�^T�A�W��<1~a"�O&��cYZ��O����O����<�;ɼ!00�ܦ@�ZR^7��o�����I,s�<P49�)��_����aoM�4��H": r�6�1��D�O���O �ɸ<�O��娡e�:;ݺ|��O�t�)94�t�zB�F�(
1O>I�	��S2vK��	7H�.s0�+W~�2�D�O���1_��'��S�x��9%��Ar��Z��i���M7��o�ߟ�'�,J��'T�	��������~�fx�Ђ�*i��� v��Ja�7��O�)�7�BP�i>�IE�	�~�H;��Hs��Yq1�@�=��K�O�`2��O�ʓ�?I���?�*O�dPS�Ǳ!e4�(Qn�^�ܘ�����'������T'���'G|���c�&��1VmD�3�@)��P;'2X�x��ןl��`yB��/��S�	�\��CgN����ڱ(�86����?y��䓻�ep�D�T'�<� �ȑ�%�X�@5C���>1���?������]�V'>�y�&�i�� �a	Xf̀�t�Ҏ�Mk��?))Ot���O>ԋC�O�'7'z<q·��T�L��	������'��Y��EƉ���'�?q��fe�&?�6� �&`�x����p�IVy�I�=��Tܟ(\8��R�2�؍��G�8\1"e�׸i&�	���M�X?��	�?���O�e��_*lߞk�iD66/v��p�is��,Ox�	�	���'����ɶ� qY�1R�	Q(3���4�sӤ@�6n��=��̟����?�9O<�'}���F�P�����/8��6�i������'P�U� '?�	��"��l�D(ЏH�8�h�"ə�MC���?���$yĝx�OF��O�� ��>=�h� AQ�H�2�u�i	�W� � �����9O.�$�O���Dl��� 8Ȩ!X�"	�=}��oZß|�"����|�������!�޿BB�0vM�R	X��_�$����� �'�2�'��X���TCT e&d��\��@�k}`F�I�O�ʓ�?Q+O��D�O��D�&����\�i�������#A�	����H�I���IƟ��'��]{� `>��eE� �(a���T�K54I��bӮ��?1)O����O�$ߴx�DʊwW��G�ԜIa��q��L�*�o�ԟt���,�	ey¯�10 ��'�?�)b8R�Z�lG\��P!�NߛV�'��IƟt�	韠��H�t�OҴ!wc�+� 9.%}(CY(�C۴�?9����l��O�R�'��D�Ʋk�*`I!��(�`��2(�}����?���?��Y�<���?������KH�]�\u W�A�������>�M#/O@\��φ̦��	��p�	�?9��O�nN�_`	ؑCS�~!z��̍ho���':���yR�'��Mܧ:z�LYրQ��4��P�>~tm�����4�?i��?A��|�Iay�dʙ"X����fV�['LpG-A�7Mфc ��O�ʓ��Ox�&]+�z�gȈ),<	�p$G;6M�O����O���@\A}�W�x�I|?i&.��\І���I�x�X��`�����PyRk%�yʟ��d�O���8�*�*��I"~��-Z��X�j�&�o�ܹ�j��d�<�����D�Ok��@���#P=&N8Ւ�QF��	��Iݟ8�I������Е'���:��@K�,v�C�!��,B	;c�
����O��?����?!��> 

!��*_�`xa�U�l�������O����ON�#��a9�ވj���>�4�"P�B�[D�#��i��Iٟ��'���'d	��yZc��Tq��7߶��2M���0��4�?i��?!����YEZy�O�Z� 8���!d��Q$�0)�h�R�i�U����ן���!g���|nZ�(������X�a�`Nߘ6m�O��ľ<�%�`�����4���?��K_�x
���
�Ԁ�2�Y"����OT�$�O�騵1O6��<Q�O�h��.�7^R!��DQ�5��5Q�4��$ ���m�؟���ܟD�ө����~��aL͝$rd�0�K7M�x����i=��'�}�'2��<)���	�.jH3� �t� �R`��M���4%�F�'�b�'��ɤ>i-O�����g����Q��	��5��aR��y�%i{������8��b�'�?�f+�7�8)��ֶq���Dc�l
��'�"�'���S"�>�-O��d��<#�ɚrji�R�Ӹ.	H�� kӺ�d�<���<�Ol��'�	�l��0�0�T�TB�14@7��Ov��Y��	Oy��'��Iϟ�)�.�K6f��&�6ݢs/I�
�p�G��̓�?Y��?����?�/Oޥ�s-���><���B p�t�Ѡ� ,�҅�'�	ٟ�'��'er�fRv�8��� =��X�BL�_4�ٞ';��'��'F�S��� ����B�)#��9!�
1�*Hq#Nՙ�M{-O��$�<q���?�C�<�TFN9)%�VM���c0*�E�Pq%�i�2�'-��'��0aґ��N�Ĕ�,�0X�i�$����S�%M���l�ş��'���'�U��y�Z>7mW5	��=C&E�!$����߭����'��R��	掚>��i�O�����:��Kv U8�KŦuC ,��F}r�'+�'Ԟaj�'��s���'
�2��AC��[zn�����Z�unFy"�E/��6MXg���'���g)?��Y�>.�l�3�H"�E(%*���%��ݟL�4n�X'��}Z�k��j���S疛z�ԋ!GY����U���M����?Y��Z�䜌g]<U9�IF�SA��Ҵ�uڶ�o�&+3��\��g�'�?�V�I5s���� �씢BH͂v���']�'t(PPA<�Iş��U�j�y�i��T�U��+���n�M�	 w��)����?i�w�	¦�7�}�p˛lz ����i@��#o��b�|���i�)I���	[
���`��?4.mXsa�>��m�U��?���?�)Ori�T���7��-j��GX���c�~�j��>����?���ܹ�IҘ������]f���
O�?I(O~���OD��<ч�� -��i�U�̉p�,	�uX�QKuE����'��[�����,���jml�V��M"��׫@���RS��4�:��'���'g�Y��N��'k����
��v��'��R/4)��i�|B�'����y�>�@fV-zF$$Y2ƎK��������џܕ'U��)��6��O��iT��"��ʈ�y	��[�B� &�������P�.r�%����h�t�&�r�n�E�?AZm�NyG�r��7�Q�d�'����??�@S5@ۼ����7k@�5N�m������Wob��%���}�r�Q#;��ɢ�E� p�С*Z�%��!�+�M����?������x�'���&cA2l�1�G̀`<B]��r�@�#�O��Of�?��	�*�P�g�OW����=��\cܴ�?1��?��Μ���Ol�ħ����:B�K$��o:.�0�Od�h�O�U��7O�ݟ��	��*�)����nŘX���� 	#�M���g��$���O�Ok,�Mj<��ĭ�74��A��2/��:̪�IMy��'��'4�8���w�PA�M����Ь�z �u�>a�����?i��<Y>�9��6��;�e�%a��II���<y+O����O�ĭ<���ݔ@>�iۍ;�� JS�	O�8@wG�-.�������I~�����ɇ3K��I�2�5��S��\�H�(9�vD۫O��$�O���<a��Y�=�O|Dj�ԶE�p$��D2V�m���x�4��5�d�O6��X�W�X��*}�b.]%�I���7_r�h�7l�MK��?�.O6�s!
Jn��Ɵ�*]�� ���"��|��0j��i�L<����?ѲN��?�J>��O�z� � RK?��ఠۛq터��4��D^�~�@�o�?��i�O��	�x~Rl��s�hl�  ��3y�e#�K���D�OpiD��O���<�~
�&�+
��[f�N�-_��BDIѦ]ZJ���M���?A�����x�Ov�h)�	D�Q�M���=3KLQ	gӐ	8���O"�O>���.�vȀ��2�^�a�]*�d*ٴ�?Y��?)��^�8&���D�>��d�"K�l�x��Y�gM`�@�)������My�g�cc� ���O��D�"n5̑H##֓#���j0�ӞFn���d�v����p�I
��	�O��OΑ8��� J� 4�M����H+`�U}�d��?����?A��?��o�
[�@]���nn\+g���b�� -O���OH��6�$�OJ�ďH�(��`�u<�5���)VKq�&�T�1����<�I����'xK�1��i
�-�ve-+@1��o�$k�	�����؟��?)�
F}�D�I�J����׾}ۂ��Ǌ��D�Oz�$�Or���O�1�+�Ob���OnTr�nT)vM���p��?�u#��Ϧ	��[������w���%��ؽT�)�,Q�H��!A,�,�V�'�Y���"�^���	�OJ��r�����N��A�G�?"X]�2�Va}��'��'2髎���?�,\76O:�b��A)uل��wCpӀ�4p���in��'N�O���Ӻ� ��Ʉ��?w��X��K>,��Y�i���'U���'M�Y�t�}*�fٿ�H�A1r#�ن���[��M����?����"wT�З'��Q#c�O�qT�X��V1gj>!�Nt���s6O��d�<���t�''���S�]��A���R�>&42�v�����O:���l�.��'���ߟ���`��S���^q����<\���>�pM�Y�����?���^#8�����Y�tI��E�82��'B~m�A�>a+OF�D�<i���)+���[FMѼ]?|�x�e[�G�IrgF���4�	۟ ������'N�UC���;Vw��;�J����!��^�d�����d�O���?q��?aF'�'&����BNy�x�k�O@�q�����O����O2ʓ
��p �?�}���-���6�ѿ8Jxu���ix�	�'y�'�R�W�����)A,L�v�RЂ��qc:ne�I�����ٟt�'���*�d�~���Ab䈄�Y�^i�)�d��� B�be�i��Z��I����\���������{��a���4���	iܹH;N�l����xyR��(Kl���?����fǾa�PRfE��_e��A"Mʠ;�����IҟlB�a0�-O��Ӭۦ�G�B K�2�X"]��7M�<�q"ڱǛ�'�R�'B���>�;lBZ��m�?Qe��j�-ۆr���l˟��ɫ`������9O��>q $�z���2��a�b�B��Q��)�Iǟ��I�?Y�O*�<Q�ؚ�j�J��89A�D�"����iXY	�' BT������P�H�Ӱ�ݰT� �Ҥ�~�AH�i@�']R@������O��I
�p�I	�c�.��.��$�~6�6�T;"(�?1������	-\pb��v��� " �T�8hn�i�4�?�Q�N���	_y��'
�Iߟ�X4=�<��!+�^c�p1��2NAX7-�O�x*u?O@��O��D�Or�$�<�r�䕙�&�# _�=s�jHV�:��\� �'��P�$����0�IO�]Z�g
/����*�un`��u���'S2�'��R�Ƞ�����t�Ծ����v���s��I�F��-�M�/O��$�<���?���z���'�M!c�;L�I����:���O����O��D�<�eΒ#���ܟH!�*)h��*EI�*AH��*����M+����O����Olԛ?Oh��y�gD�8߲Qr�`X�����s����O�˓��s�W?��I֟���=�� p���mHH�B`\�-(�O��d�O�����+b�+��?ݢ�a��'�I��˲c���D.n�:ʓp"<���i�R�'���O��Ӻ�seܒXV)ZM�v�v��V�M���ꟼ�ƈs���	xy���Gll}�BQ�6��= �5S���
�8/�F6��O���O��	H}"P��bs �X��o��re�+�M����<���?����O�r!�9u��x1d�Y$u�B�2��r�7��O���O�)"aB�{}bP���If?��߼w$���T�d�,lsEU��'����dz��'�?����?�7oG(=�yy���"Bp�C��2��'��hY�g�>q)O,��<y���%`	 P�C�ǕF9RbpE�d}@��yҒ�8��G�ϖ�$��Q��
��͓B		�"�t)1eb�<Q��A,5J��`��	�X�P�Nw�'@�Jㄋ	9�p.Ԉr��8��B�)zVXq�i�=h1شp4C+�Q��}��m�WOM/��Qr! "�8�l�+DY1�E{z��b㌆_Ƃx�&R�v5G�^�n�$���wx��q�U�[n\��l�8�0�#�ٔ#Ӵ��vᚒp��)@�	�,p��sƍ�VMBli���(J�H��G�ѿ�?����?!�iYH�}�u��l,��ֵ֥v���A�z��%i Ja�Ds,� `��<��G�v�:7C֒,���E�ط{.��`O�)��cg��6C��w��w�!���?$ ��'�� 1b��vV�(8�����,�@=O6�����g����S���V�V(R^a|B� ��.d*�)�NLa#J�`Z��5���'|�]>��U�ş`�����f�����5�^\�6ً�@y��3rJb�v!��h&�?�O71�bc��x-@��Ɂz�:e�
:6Vt*D�
�V��eh����O�I���]�M��$ydnǨ��V^
����O�S�SM�I:.)h��$��7Mٸ�
R���rB��80�b��f�G �F8"Dl�(IQ#<���)B�B�$z��P��͒g�V\�1����?i�N�F�P�ۥ�?	��?a�e[���Ob�$\�8����w�ݚz	��e�
��IJ�ؔ��L~Z	p2֟ўL�X\�v��kQ9DTi4+J/�?AG�$�V)rgB�	v�p�3ړ%|>��H +������Dl��kD���ҟ�F{�[��J@\����S(yE,5� &D���6G�.��C�i�ha�lH%�HO��|yr�!n�6mS�f?��[���<b�A@�i��5���O��d�Ovy�VC�O��Dq>9�NZ_��iwG�'"	C@�t��@��22�N� ��Ix� �U��)�uc@M2y�r��&����ȧ�E���4�ʦ/����>E��'��GH�(��x/ך��,b ��H�'�BI*�E�:�L+�ϖvs�IQ�'�0\tb�t�l��!�7l�dHX�'�X듂�ף{����'<Z>� NEI�WF����� �0(�x���ב/�v���O�����;ͬ���ZGZ8��k��0G ��OjC2�N�^��Hc�K���R���2k��B�gBx�$�bcG&��Xkw&J9^v��ĭ�<X:1��П|���q�Zb�&c�X������ZU����M���ƭ�*�I���<�	������%���J�h�dz�<�O��$��(A�ԄE��hr&��h���$�{�H������M����?�)����Q��O^���O�@	@��	86(�[�h5��ɀ4�J��@�T�Z�b9��/�i
��'���<)�Cԏ}Qy�JW�79�HǢɘbk�AIT�ŊD���Q��D^�9�eXS�Ͽ+�N`1�"%��q>"�I�� �^ÎA7�[۟x�I-�MS����i=�9O��Da\�QxA#P/q��`�'��'�!�@��%&�cC��bqr����)y�4���*��f�)�4b��&	ryi����wT����'���s��A�-z�1�@�w�8��	�'0�`r���/�ȱ���	�u�۲
�'h�4�u�
v�",�D���o�<�2
�'���r"	4c4��8cꆚY�L9	�'�����"�*��)`�E��!t8�q�'�0c���0~(p#��/�<�X	��Uq�T�
��:�*�
A�t<���$D�tId���-�f�c�,��l4i#c"D��(`�ƾa�FAV�O%� �0�$D�d�q��)1İP�h�7E�����$D����$���^#0 JPF("(B��' �uQ�)O�Xր�� ɈpH	�'�ƠѠ#�%ܼ)B�[�q����'���`��M� �� �cW&�|И�'�*-�g�մ+�Mju	�+ �~��'�v�!wH�,.��PE�ǁ
��(y�'����'��e�dYJ�%�6��,�
�'�9;���
�� �SIƧ&
>�!	�'�ŉ�E�7[���@�K�-"���(	�'"��C��6�V�I�EK$��	�'nN��P�߬
xp���
։g��ɺ�'j^q�n_
t�vU�Ѐ�\b:IR�'$>��7M˥Pv����a��X��y
�'�N!�"��Q��ɰBߠN[*L�	�'���6蓪o<�Qb���81��2
�'P���A&��8�k�,
ƠI	�'R� H�J��d=���AME�'�Mk�'$Z�m�*�l��5b���X�"O���&GL�75ZE�3�[�Z��v"O8��Gރ\}~�#%R�tm�p"O��#jS0
����ԫ�� "OB,bR�/S�h�X��U,T*r"Op��SK[�Amΐf�e�� �"O�HQ�#��t	�كQ&�-_� ��"O���(�8S���6�չ�iXR�'�$iVmǲ@Rx �eϘfA08�@���������S�)�s?�-#�$�B>�5�5K	h��F|��F�a,�������v�cɟv���Κ8D�<H��H��SQ"O�|�w��K����T�"�v���8O|�����iIP�j�o֮H�a�$O1A�d���T#;@�K�Q��yr�ȩB��tCg�:c<��F�׃_��j�'������B�<Yȟ��4v��I�EW� 0AٍC?�1���O���䍏#����&�UQ:�SR�ӜTЎ�CN-}��b+��'�rq��ɶs��;���
�p8� O)-S�#>��n]�|/`�SԡC
��O[t�K�aH2Ɍq\?F��X`��0��a�L&�Ya�NV=U��scLN��|��2�t�5�=3��d����X��'h�ZE�f��B���C���R
}�ȓ�h�C��V�r?�ƤĻ�n0	ю��<iw#PhDZ�)�'���A4Or� @��6xH\@u.�kr$��5�'\��#�����EFX3��7�٦>dT�X�'l�epK>�	݈O�Y�g�G(a�^��CMϸUm���b�I3/���H��ѩp��Y7�,�D�6�δJ&KU2Y�IŚ�0)�Mi��� Xh���*��]*��� Mb�H�<O����ڧf�H-��F�0���~ʟ6xa��πԩ���H�!TȠ�"O�䋀E]�uLL=q�gB�beTl�`�I�P���Cr6$i��Y��1����A�a�E�2�F�"5�İ��7�O�Q�@+�}���98�%xₘn�X��0O:\��|R@ٵF����GF>5 �i� ��c����=�V���'�5I�Ҡb�s�4/[�g��P I1w�|	0u�U��yR�0?�G����C��V1>�X�����<��P> �~5�3���;�!��ә"�e�����9sT]J��ɒ����c��`5ۺJ�$��PĖ,l��q��<�K�)M|��B��]���d�B@��˂����}(�bą�!�DYT�e���J�2�rE��!�R"�*c��V넨�C�K�)r!�D
U`d�b��'�Ҥ8��>T`!�Ĉ���J�J��f���G8E�B��z��1��(�cP�(a.�4s���$�6{�,�\#���X�@�9rԉ&D\�Mo��
O�4#4��F�$ ��Bɫc�R%B��I4:�����8H.��|ʇG��|�� J+�[e�@v�<!"+K�O[��s�]:<@Ȩ�Q��ן��4e :�̅����xy���Ήv^@�Ѭʿp\��Wj��8��B�I"�hH3�Q1��$O�&���C�p$b�8e��b
Ó?}@1�H�,¤����5�R��	�1�B0�S' �	��Z��_6o���!��Ò_�(���Ni<�vQ�
>��R��f��E�c[�'d������D������J��h.��A��,8�0�]��y�b�@�@1��,�3W�=�6�D��y�1=�2b�"~zBA����
��R2M�"�z��_�<a��=��b�G�,Y
������[�<1�/O2�ԍ����(O����kBa�<y4�@�
.�Ԫ� #��(qf@�W�<)�$��F@qan�ȰD��\�<�+Zp�x��ǜ����m�[�<IgOX,r;�p b�
!Ԫ\Z�O�T�<�p�D9V��� ���/j$�5-�H�<	1@[�S�^4#㔞J�f��-�H�<�H!;|dX�@����c�G�<ys �H�IGB�X!J�rѾ�y"d�k��1 F�^�0%p�1u����y�C!�q��P%'�$��7�y2*B"v�� AD.Lo0�4���y"F->l8&�FX��	A"X��yg�*,]�mzp�$8B�T ���y�B�,� i#�I� ���3l2�y�)��,����P���큕�
��yBˏ,�,�R��<̌]rkR��y�+_7nV$�K�'8�L �K��y�
�&�<a!�>/��9BA��3�y,�60��q`K:9��1��^0�y�O��tX��B��YYda/W��y�A�5\��O?ac4F�1�!.�5J���8V,+D� #�&zp��"+�J���o)?WIN&Oa{�͓R��0�K\�A�v�0�����>�g(]��xl�=�4����d�aQ�Ʊ
�PB�ɵ�"�գ߾&z�X��.�&�"=1G��24Q��D�4M~������Ȕ5 B�Q� ��y�n����t�F��~qfh�p��:�M�2Oʧn��<E�ܴ4_wꃗZR����κO�^���H�@�_O�P�� �C�	�'��&k1lO��2�ⅰ5��P��<���Q�'�j����))H�ULQ%5_N�ؤ
Į]���ƓID\��1'UN7$DȀ
]�~��ɾ=!�Q�?)���6�F	2���BU %l�x�<��"҄V�E���UT���ՊΠz�"L�I4=Cʤ��
�-�7����� 0h�ןQ�t��.�`cM��"Ot��D�jg���K�T��`A�JG�<�r.H�� �	�$&h�Ώ3IP��t�KZ�y8E�)�x���)�+-lO"pG�uE𤪰�Iӊ����?}��5Rb	
:y���2��-�^���'BΨ9Tn80��}�q�Ӛ��$Џ}�.�{��;��H� @9����9.��7]?��� ~�
!��'..����6K�!��&SX-���h*����k\ �b6�łOZ`�@��y ٺı�O��ع�=�а��	
 ��`�t��qOl$ŭ��t*��Љ?"�L9�NU*q���dQ�b/���%֤3(Ԥ����?����X��F���C%�+ ������5,O���B��L���E��t�V�CQ]�D�Pi����_[���-t�P�I� ����>I��@E4��h�1/ʠ1���l�ɾ#ޔ@1fN��)Tk���'A���:�����\�lA9�vj�\g�Ai���y�l8�a�T]�U�B\"u'N��P�˂�+5P�Y#�5r7�%��t��}y���1d^�GIٙ%C(��pF.��x�a�	`��h����'�ԑ�gi�k񨨑���&;�y�E	V�L���z�'����5+����oF;&�H��
�*��,�3�Ϭ6�z��� [� I#��=���ӬƥC���P��d��|�����#��^��SV��M�'=�,����	-�@�_z���S�1yj�\��$��F�Rщ� Me�C�I�hpV����J� ��\k4*�oT~t�o�LL�	ԅޕ�?�B�7�ӈ 4�I:��]��y?��r���C�pC�	�<}��rR.����!��ׁ2>$��ԇ�geB��e�?"�~*�KҪ	�џ�(��;ܐ�5&�w�Y0��=,Ov�#�c\*6o�<�dhWXź��� E�u*d�Q�W2������.?�R5���~k����BKplh���<�&����@�-j�y0��S�|�4�D*=P���ɤ@xB�	�k �����<O��cv&�).��*	j�I6P�R]��O�4I�o�P�|�"$-E&R����"O�]sG �76��[�N�_��`�aN�7�2ya7A!�O�u��U(Y�L�Z�-	 �LȂ�'.m�@�h~↖4T�t�� ʰ�^�P�@N��y�b����"�kJ�>0@���yB�ΰk��D ��`�bb���yB�F�8��4�N�(zb��sB���y2��S`�Fm������M.�y�#_	H
n�2����a�����yr�ق!-���LZ?4 �㖣ۮ�y�7\`IkB#�r�� 1�S�y"b�tp�e���-�@�����?)�b�px�A1ĩ["NH��i=��0�G���ab��e�����	�p�L�9���=Q"��jMW�� �?q5�	4g�T����H6Y	*��D)�%S�zy����%�xrE�v"q��'��P��ՅY���k��0*p0-Ov��ǯ�<^�����U� *��(����"ph��P�~�XD��WJ.C�ɧ]��R4#�~�xĪP�.kN]
P�X.A;�젇�F�}`��fD0��d&,0hT�� Z&@�C�Ɂ'g!�d$(8�4�毟5L�6A�Q͕�QU*Im��y��n&�|���'���ʀoA	t&� �${����d�<E��X�f�����]8�	*t�L�<5n�:�X(�GO蜰aC'TD�<�W���(�\0�b�)��!hs}�<�4"�n���]�k �)�G��{�<ɢi��_*P��O�ari��u�<�� �x\�� &��c���*�n�<�ĩ� h�z�ch{��z�,k�<aq�Gm��B�	<n��x���N�<���,!b����X.\ذ�mI�<1���|tL!v�Ȃ�0�p�gZ�<��@����������5P-pDA@L�<Y��
`��C���l���5�OH�<�5���f�<���OMA�uC�G�D�<�1�$&�t�AEO�(��܁��v�<���	'���I'��
*�Д�ao�<� 0d1�@R�zz!�EB�`L��"O,��a�*ߜ�s�M�(O����"ONMc��@-+���Lsg\ �b"O�E;�	Σ'�p�V:Sh�ܸ"O���F'���z���-D�<�*�"OL�q��*E��u���_�@��њ"Or�P�ˎmش��F��TKV"OIb�L�< �:!k�#�D�#"O��� �<�F���:T݀��e"O 0hrȄ�SQ4A:��@�3ɴ�E"O*4���"<�dh8�O�<?��E�g"O65�£F�C�dB�n�/�.\t"O�����~ږTyt�bR��r"OB�t�M}�l5ʕ"Аm�Tj�"O� Qd�@�$7�H��@E>.iH���"O�M��	 �,�*`@W41R4aBf"OVY�A�A�B�BA��H��pC"O�#�A�&y:UDF4{��rP"OjhQa瞂GJh�`$Θ%��Tc"O8ј�"�:��4Z�W� ̚#�"OX]��KB0Z2	{��
�Y��"OQ1�О�4=�lڥB&�+w"O�]��c،a�:���J�R���"O�8�L�#aK>�cף�	*D*�"O���ɖ!uA@Ta��Ƀ"O����)]bTq�X�9�Z�"O\�)�g����;��M�ΈA� "O�!"u�T�_�.9�`�N��X�˃"Oh��H Y���
���v�J�"O���|G�kr�Q;���G"O��R���Hb�^)q�<ͳ3"O:5p��;̨����U�b~�ر"O����F%C.4i��;a�e�E"O$y��嗴J,�X���F.J0��ѥ"O����(dz�t�`�K
[����"OL�	E[�)���i�8m� �5"O�
@NEL2�h�)R6d01�"O��x� fJ��è�(G��q"�"O�Ia�ā<^���B��D�.�5"O$y�P]k=B�K�M�����"O��F+�<	���\�(��d"O��k�(�b\����[=���&"O$�+�'4m�Q"۾7��|�u"OB0Y�F^�#^�@'I� A�"O}��-qHYAp�ݓg>}+b"O
I�J8�h�CG%k\T� "OX�b׹9HqA��K�Ns�"ON�b�N7��" %Q -j�az�'�t,�1s��1j%��[�֠b�'��=0�bD�yhٴ-��S$Ψ[�'�^�	 �Rˊ����0E�>�c�'�欉��\�CI�H�#C�+PB�DX�'!�Y��MI�2�@l���ƣ~,`��' �t����bO�pc^�qX���'Z��CЇ�R/r1�%X�f��l �'�����/[69r@r���Y��yR��0}0��T	
}�B1�!d�;�y��/j����B�m-@�X�gD	�yr#P�?|�k�
H7hZ2��� ���yNF�~�2Y��EO�ڽK�N0�ў"~�Akje#�bÁ{�4
a��.KX��ȓt�V$X�
ˉ4�Hx;!KV������z���i�4�Bq;�<T��ȓ4�F k7e�lZ�����2����?����~� )�"�I�ذXJ6�����"O�kD��2$]��pD�R>&�R�"Op�����/�����C��'O��"O�ܸA��t.L�pq�i�� �\��y���� N48QnAJ��I2�n�y�h�&\!A��3I��v@B�y���+k�\�R���S]������PyB�A� �4��Η�D��� OY�<��LˤH2���>��p�NQ�<!�g��r=�xH�F������M�<�� �(o~�����#l<R���O�<��BU8j�4�2Aa��M��Dv�<��/�%��3�`�άc	�p�<�3)����qDț�x42���l�<�7ꞹh6�ҀjY�G����i�<-�@� �)�v�`TJG�_ʊB�	h���i�F�A[ZD�R*�M�|B�	�}��\*���`�F�k��T�U�B�	/d	�Ukv�ѕmdDX��
��B�ɀ d�(�$��=�`�4F̖ �B�I+2f��'�-����w�J�CbC��.D�luY�/��
8�x���5K�C�I6b��"C�>�hf�:m�B��%Xz>H;d'T"� ���烽^�C�HZ�)1��!X����9N��C��HU��	ڼf�J�p�N�>�C��0�0��!�E�s�[�y'zC�Ik��:S`�2=F2u��GƠA_DC䉐VV���A��q�4��j�'Z�pC�IW~��W.�D2�s�ܟ@�2C�I0&�����
 Ϫe��"�0K��B�	k��H̍�fx����X�Y3�C�	�"8B�i�gLCv� ��ʎM��C䉄8̼T�U%�{�i@&T(7B�I�y��+V5j)4�JQ�3��C�I,r4���$�c1��M��C䉑N���EJ���"�ɉ�-=�B�A"x]��%Y�)s��x�)HJ#�C�	Q'Z���,�������ǢR�FC�I��ibRȇ�~�Z4;E/�+w`jB�	K�mɢ�5g�24�'��i�
B�=w�H���<.tX}�1h��C�	A��ɂ�!x:�
���O����3?c�E�ݖ�]��@�"���m�<���/꼈���?2CF�J"dc�<Q��JQ�ͺ�%N:� ����H�<����(`�Q��T 8aJq.�D�<iE����`���I0Nx��@{�<)�
p�T�Pg���pU���A�<q����-�"���M��!�CFc�<�ag��J�\��,ݛ����-�C�<y���,i����ǝp��= F��}�<�Tf��W��qʱ%�!"�Ό�0nCx�<#H/<�(�EX�Ic�i���p�<����
e�x�y��e4�J��wX��Dy҉K����4��+|l�A�+��y�A� {6�S�oP�{�����ٟ�y�ťZc���M=H���6L���y����U����";�*��aG�y�o�9C+�u��΍�7�<˵�*�yr臨8h`A�d�%m�)�#��9�ybF۲!]hȀ�өq�0��[��y�L��VR�!��
]��j��A!�y"�F`c������Ia /S��y
� l�ٶ�@5A�D1a�]	�`e��"O�m��G��*,2S���j*��"O�l SeJ[��<���m���
�"O�ɲ�⍙i��a)ㅅ��� [&"Ori��ќp|JA��N���oׂ�yB80����r؂���-���y�
U8u%b�ȕ阔h������yB�����T���ǚiW���Ц 9�yҩJ�M|�����0@4=�'�H9�yb�X39� �b4�Ku4ȳ�B0�y�k��8[�K 
uR�LF{+TI��O��=E�cR:m��5��%�64Ƣ|�$�y"�( 樹y�o��|��\[�k�	�yRoP.0����C�g`��[ņF��y�D��������:X��rd%���y2�ҦwBޔ��&��?(J)H䂁��y���)4� t�OnRX5�sl�*�y"���U�\��P��;_SfZs	��y���# ^��уպa�������y�C`�8qɶ�T�6A��W�y����|�J���	U�`��#���y��/�I�'dG8�
1I���y�GC,dm\�ٔ��41mt�z��Ԧ�yrM� ��i�� 89���S���yBDE+~���gA�d���3�+��y�\WP���F:5:�y�V�)��T���9�t�`tG��yBjX;:1^�C��6�v-I�+���yB��C�T�� �5����Q��y2�J�G�S"9��I+��yr�O�_<h�F	�b�����yr@�&�V����^\��@�U��y�O)&4��EhL�i�vP-҉�y.�7"���rD�0Z=|q�'@���y"^��$,2�ߣh���(��W��yb���f�����3N�PŁ��+�yB@Z�drF110G�����*ɑ�y���Eb�ӁGY;����G���yB��na�a�B�>A4QbG-M��y���^��r�ѵ:xF��穜��y"C�Sک"l�v�=�����y�덅�x����"h5A�����O&"�Skڂ1䖩*f+�6e�����ZB�<ī��>L��F�<��C�g�<�k
:Jjh0stG�"����"�J�<���M�a�|P���a�=���C�<!�'G�o�X�#F�1(�V,�@Oj�<�&Ꮈ+�D�h�**,유��m	A�<�J�<B����ˢ� �� fX|�<)T��qN�#���xL1���\�<!c�X�K�l��)�q˃�LY�<���S{��D_�I�\�k�� A�<)�fL�F����@�&&M�b��|�<�"�/#8�L1��\�Nq(��O�<����Q��]q�,M	H�D�#�u�<9d�V�'f��At�H�I��p1� l�<�U��d�l���C�'�)���|�<��Ɩ�JJ�$@�!r(v����N�<���.��@�S�H)�0� D}�<��ᇑN! 3dm��qg �s�-�x�<i7A
J�dp�Ѓ��K\��C[|�<A��V�0g�	S"M#eJ����@�t�<1�_/MBL;aں!�z%H�u�<A6�=�H�S��3t�l�� �t�<� H� q��'G�5�)8��Zb"O"�2�݋>�p��VH�	Wk���g"O��&�3zy�`Z��[+@.���"O�\�$�L&9� ��eH,Y-H	�"O@�����OvJ��9	ڍ�c"O�ɠ%��l>����X��J%"O��	���-�OX�9C."�"O�5x��a:��@��CMdeJ�"O*��hU�I�MZ�z�XX�U"O����Ǯ��T*�LȀ&��dQ`"O��PF�5`3n�3� �Ws����"Oԡ��%O#$$��lRT9Z�"O�@:5Ɓ(����q.#B yjP"O�Ԩ����.�5���b.����"O�}�5�2|�X�$��P.���"O��g�O+Q�V�0��X@�U��"O�uR�ώf���@�8����"O��``��k2�����K���6"O�5٤;?�����)�KoH�k3"O}���JA<| Ň� cj��b"O��{�cP"uE��`�ty��"O
�3�aA�͸0�}��H��G8D�Ae%1�:�� N� 3����`G5D�̘�ŀ�I�xy�)�-S2��0d5D�4:�"�h�	��W;:��B�)D���d����axR#@�r�N�Q�,:D�h�`�K3Hv���p�/5��L2��9D����*7U��P��҂(��Ȳ��7D���P�S�lq�AACP�v���i D��Y�́h��1S!BZE�̰��=D�@�'EV#M�P�@��"h���[/)D�|�����3�d��v��<| "`(D�txBK�'V��e��$x���PSc$D�����3��LѲ��D�j���#D��s�B�7r{��K�B��+8$qu� D��:L�2z��ɠ�T�T�Fܹ��;D����"�xx!��R;,���,%D�tjG���U� ]Z���:�\�(�.D�\z�o�$w$D|�@��<��7D������(B����;f�
8�k4D��ʶF�c2�Qt�BX
2٘�3D��lS�A��2�`ԎUV\ղ$�2D��!�oJ;?�,� "S�>t��y`N4D�,�&���"�Tx�!Z�zd���1D���%e�|�x�Rgl�h��ǁ"D���#��V�$���:z<,T��>D�0�'�B3_S���dOMh�>�M=D��P6h>'�^u���K�=�t`V�6D�d� �H�M��0�B˹(3ZĪ��4D�4�V�Ӡ>�:��V�-p�̛��1D�x�"^H)�%Sc���	����B�"D�8��3�n��u#��%z���?D�H+��p�v�t.r�5���<D�X�2+�
69�׏N��X�� ;D�0 -Z�%¶�x3"²c�:D�X�WhU,n�*)���Lxb� �6D�i��� ��ɀ4a
*p�6�{�5D����'��Sِ|R7��!"�Lt۠�4D�ܘ�Ĩ/l�87�R�@@�C'I.D�P����'|���U��T9�a�
�'��@w*m{Q��bI�B�B��'g�y�J;O��	��·Q/�I��'{Z�{"�ĀIrP����G����'���faI./���a�+��`i��� N�cwmѽh�60�U�مF�\�"OȘB�B�Z��u���9`ݙ�"O	��hE�6�(2PK�;/���Q"O֕Jv	���)�u���Bڂ�p"O& �pi-A�t��J�ȴm��"O�L�M[���yh���:$��#4"O��ä���9�
����TP���D"O$Pk�*V���DمXx�J�S&"O$��S,!L�L�ӳ ����$��"O.��I �!p�[�V�%#�"O~��G���4	��(\� n���"ORȑ"��J,ʣ�q9�R�"OJd���ԉ�۰EG�(n�y�
ҹ�8��<*�e١���y��!��k &!�������y"i��_y:� ���M�v9`�mN��y�,�50�<�*P����a"�ǅ�y���l����a`<i��
� ��y���6���H��@6�T�0-�1�y��E�(�f����PZ@�YP��y�!8�b�CD�NF\��0��7�y�N�֑[+T
K��\ �	D�y�̖�г�B�!�J�8A@X��y�͜V�:�p��݊8n���C�&�y���3Rz6 I�NH�0 ��$���Pyr�P�r:l�8��Ϫv��R�N�j�<	JՑ
6zɃ��"%,QYU	_�<!@E�w>)8$oN�U���EY�<� ��*�2����A�O�(��iFU�<�sA:.��X�B� m�e��m�<�'F���� �ڽ���Kf�<	�1>Y X�C��=и��HOd�<�%�ǡ=�1�$郟|�ҭXe�^�<!׶`��0��LW'�(��A˚]�<���T�P�,���@�FM�4'^Y�<��m����c��?8m<`�A�<IRN����C`�A=P���#�c]B�<G&B:��E1��=��ۓ��w�<�0T�k>�[a �iz��2v Vs�<h֦+ۂ(�h�'Y��XV�6D�����	6(�(5)�~����A�5D�pإ�>;��S���#dZ	�C�'D� �0�_�v�,]y�hʀq�\�`�$D�4�Ǌ��R��52���P�ǆ!�$˄\�t�����Y�j1��$v�!�d�y3~蘃-�26�]3S�7t�!�^�&  C�E
�Y&JAbg����!�+>m�,e �$�< C��t�!��QaZqcCE$.����E���Nz!��B)'��=)*�9wZ�	�&@��PyB�
dxqp2��t�ȉ�� �y��~�ˢ��n_~��  �y�n (��l��,�T�bT
�G�2�y2��e9�t�¦8��u��yb��J��a�.�_��dB��y�I�A��Mp4��!l#���N���y�4(R~ �3fE?��8�F
�y�o��s��E�ѧ�6E*����(�y�`fikfaS������:O0$�ȓ�#�+\<Jܘ�[F�V�m��Q�ȓ$+l�S�Z�)�:hSR!�s+(��M	��"�СwW$S 
G�y��(ܰ��T�����MU11ƀ�	6"O@p��.7~�2���/��G"O� v��&�΁z�up�e_�#�NeZ�"O�4h���6K�h��B}��;�"Ot��!��.l�@!a��sn.�°"O��Ơ����Ʈ1��ʡ"O�$��%w �HQqH�,N���3A"O�-��f��l)�8�ǁ�C�9k"O� q�'Lm�lT��&��n��"O���pEڢ'��`���6��l1Q"O���B�1R��1�1��)��9iC"O�e���I�X;��?�t�c5"Ob��F�=llH�!ƭ
W�&���"O�<� �'Ȏ��֡�)f�L ��"O�Cŋ�V5H!��Y�^,�wO��q�!����A%fX�`��-<O��3�1D�!�w�ہY��YQF�"�B�	&s&n�{Μ�c*qx�� M��B�I�"R�K�(1`}���#%�B䉆Nxv�3Վ�--*@��f��A@C�ɴ�t�����)n����%��H� C��;+������7�
��Ђ�_ C�I�T%��+�� �9�~�	4T�2F��E{�|b�)���!k���\h�����D;FE!�\^�e1A.QKP�9T��,T?!�ѩ���{�m��X.B��u�B�C!��[�^�rd��9CHq�!��2�.�rF	V�^�����ʖp�!�D�j����橖�'���0d�� �!�Ğ�\x`�i�k��!v��3��75�!�D�=3C�3�j.||�3�*��!���}A4�"I��{�,�a2�^��!�D׊�t��\$^(����葫7�!�$�1Ab�ԯ�r�0m�`gD�(%!�D^"E*j���$�4�֡�S�+!�䑙3��Tym�S��%р�Ú���$(����a�>����
PB�I:�ȐR��F~&�R�$մ
�zB�I7��(R��ϗ|�}r�.��"�B�	)!��ձb��pJ�l�G��QC
B䉮��qq#�)a��8���O���C�;xҮ�B�woV ��c��e��C䉇\ � {���$&z��v-̌l�C䉾7�0��M�6d�b��ɱ���d$�Ĩ<I��d�w�����V�XZ8U�D)�q�dC�ɰ<�m1���0��@�=#�<C�=H�Z-X5A�8}e����D�F�$C�-��Ɂ�ŭE��py1���4�>C�	<����c��6�Ԭ ���%,6>�=�çX�lH���ȥ3�HA� n2�'����ן���""���We�lȢ0�į�uǺ��8�Ş��dL�D�|`�w���]3F�ҵ�^�!�$:	8pW.�`���[g'���!�$�F�<�Q]y�����ul!��G/#�f����l�J��+g�!��� �Ɓ��G�C���0��|�!���$���RBf�sZp�S���S��O@�=���L�S)Iv�ŁfI�
�д��"O����A� 7Z���È76��A-D!���CӼ,����q,`B��C�!�$D��:Wɉ8�����!\!�D�����JPހT�����1�!�{����H�a��Y[�U�c�!�ē�� �����:��1(4�1��'�ў�>�8�%�,rj"�%D��{zْ�"7<O8"<�r��3=~q+'-��C{�B�Řn�<� :8R ��� 
�HsI³4�^�R�"O�8�,��QQfePf�X�r��t"O6x���,�k&E�a�(�yq"OfA����=F�:�����/e�Tݹf"O��a��[:I���ʂ���!@"O��2��\]SpY�a�	��gr�<a���&o*�����6X�4)���kx�T�'{8L-ϛ7�NYH���C�\���'t<��J��H�B��e�ǧ=���'#��nٖ�BP8V���=�;	�'�01����-�y�O35z�xZ�'�<d���]+JD2���DF�1UxȘ��$(�'T�R�3��	SșKî�);� ���vL0s��B���E+W�_�@z�܅�hִ*�-�B�PMx�m����3���J#k	J���C��@u(vC�	�u! ĴV�Ű�N+Y{0C�ɢ1QN�U�8خ�A�G�f�dC�ɸs��@ɳ��LO��ȼBc�C䉱x�X� Uk[��|�b�X$A�r�=����?Y���?���?�e�f�"�"���:�VCU5�?����������"�Ġ\����+>"N��@#D����ξ~���`�յ*�<u��!D�,���^�]L��QO?<.թC�?D�� ��H��	��!����-#D�<:�a�p1z}���'0#b�K#D����m�L��x$�����0WO.ړ�?)���?���?A�TH(�Pj�e���ӯ��&O������?Ɋ��i¨3�h� 6h��z��h�����pC䉋m�4����6^^���c� MjC�	�&���H�
c^�tR7$� 4PC��(6,���"T������*
�B�I�$�t*�k�*49� �B�ۂB�	�h\ �a H܅x�z���I�v�=����?���?���?�!B�//�Ġ`g�-��	a��]����hOq�~��ԬF�0�cO�l-����"O,#��.'z ����N�i��MzT"Oج�RÆ>C���#$��Z�q�"O��Qg���hiK��A5X���P�"O�S�3 ��h��}v����-����G�	h�:ݑfö\oh��06�}���R
/x�E
B�N�����@��I
�2R���ڜ'�ԅȓG���_�7�P3E�� ��p$0� ƶqf�0uj�,v��� s.T��5B>��'���<�Ɠ��8*�e:=Kxart�՞[r^a���x���+�&�(��=��r��P��y�'?ؼ�@�G-��`�G�$�y�)��6Il��T�m��Xc؄�y���<sȉɦ,��/�8�څm1�y"�X:^�.(��Ī:�P�(bE\;�y����)��D����<��ɡo���x��
b��š5���A��5!�d�B� Ek�,M��ҁ�4�џ(G��ə	�~䲡�H�i�2A;��ٷ�y�*� �0a�P�or}!�c���yR�\N�P� 0�ڊ3A$��a��*�y2�D7'څ� KI�T���g����y�	!`6�5���N8inŪ׌T��y�ʀ?�va��c^$m���I��y���9a�-���ޔ�f(��a
��y�F^�u��q�i�x#P�A�O��yҥ��.����H�]% �B�A��y
� ��5�D�~S
��A �,G�q��"O�{4jC�+y��SH�))��H"O(��p��*vR�P2�V+$��,b�"O�V�E��,cd�Y�.�,I�G��j�<�Ud޷r:��� W$14��AwfGp�<Q�@�V5n��.��tAă�A��ݟpD{J?�:R�>y;R(��B(�l8�*D�|0@�=P�
�pR��k�01�3D�l����!�i������+S�/D� ��a�!���v�P(D��t
�I/D�@��GQ���Tq���k�g2D����kR,E�t!+a�"*��C�1D�8*��V�(�X��@>!��=)Ê3���x��S�=���i"�V�N�ح�f�Y*7�C�ɖq�~!*�JQ�`4���MEj��B�ɠ+p�Q���se2���-ȃ8�B�ɞ<��([����%b�	j̢B�	(U\�����X5����B+w���ţ|�FDX�o�i���@��I�r@!�dW��R)2����	������1d_!�!�`���	\\���W�^O!�$�5������^�}�Z���l��;!�d̻ �
 �qJ�#Az��!��j'!�d��{��9J#��$]T,)e"
_!��2d�Ω�G�c6P5c���%+�!�$���h@1&bT�o&�2�~C!�F�/S"�P-�^��M#Ό� =!�L�cJt��`�<��3 B�(�J���r�A�D��z�!��y	�Q@5�7D����j��cW�!H��Q�jn�bek:D���T�A�fdd5��+7r����!�<����S�C���3�o_�sx�=��c��hFC�Ʌ&ɘT*ъM�K������E�nbC�� 1��𬏪$~Μ�e��l��C䉨^H*��� 4�����/Q3]��˓�0?1e�����UDӳ!��ȹ6`�_�<�F	�@����"���&\���N�[�<���;.ʲi��W0e���a@�o�<�`�I�p��4s��^�z�mZ��ny��)ʧ7V�$��Ɉ$]�A�&9MԖh��-�1eK�'d�<�PB��.+2��ȓ%�%���ޤ)-\=��o�J$����	%T"(��G� W����J�q�B䉫H�d��ӌ܍r]����28C�I�5��lpq���O�^�T��f4JB�Ic��k��ǔukJ��'$�:��5��o�O^��� 2�$���?}�D�b�"Oҩ	&mK�hѨ�*�3%��Uڠ"O矠)�8Z&ʖ'H��	�"O��Y��R�yRCei `ya"OZ��4lQ+o�0���Ƒ-Q&�'"O�!��(�Z�=S *3F4�QU���IX�S�OϾeА�
/(ruUk^�9 �-�)O����O���>�@� #c���av%��@	�k 	$D�p;AN6(�4J���Y�p-�Ө"ړ�0|Z@��]U~8񅮌HjȢDBk�<ل�3����	b�0���k�<�ԅߖJ��iꆥL6'U}!E�\�<�L��N��%t&�19xAС>?Q����<`�̙����^�N�@��{&L�<�I`�T�Ɉ�~���y����9��|��C�	`L]��7�-����J6��\D{J?͉�G0lN����P:�hd0�,5D���O��(�� ,��+�2$h�
9D�� <� 1OF�b�8w�8,��b"O�1�Ǐ`����φ�h�a"O ypg�æ)E��`a.�� Ъ<��'Oў0E{b��Ny����T�Ŝ�j0��5�!���:HX���A���Mj4�P�]ў����+WVuµ�T&�Q�/�9�̓O��D[��*LrƮ�o�{���G�!�ǿR
њs�K7@ȂVN�Y�!�Y(d��qb0�5���!򄏯�b�hf��,m0@MS,��DP�����+�V�˵%�yO �R��F�$4�Ich�6�hO����&ZJ��r��!���J�V�SK!��W�7e|�Y�m�4<��h�`҅w�!��̙Yk��fjӮg��0	Ɔ�"4�!�iv�����+xn\�d�ĭS!�DC�IS��IҢ�j�xd�@*U;n!��n�,�R��<N0�ҥG��=!�$R�t�tl��;zA"�a ��!��C~�L2CZ,- ��Y7j8\S!��Q]ҰZ�)Y�z�N��4<�!�dV��8#��K("mta�O"#�!�ʡ1F�%�2��,S\Q�a���!�R1*9 AHխ�
#۠1�`GkU!�D�'B��0�T�C��Iz� @T2!��ĕl�.)��,�5?P�$�鞠U!���؛oU�[2)��B"|�ޅ0WVC䉘oH���f�5(T§���pVC�ɫ:[��"-"bi�B(��F�<C�	�F'��x��S�'.y�`��0�JC�S����u$�q�(�A����0?q��G�c7��T��&�>�3�XX�<�����$�g�r!\l�#S��$�Itw��x�.�4O�L�f��P�|�����Ӏ.2�����d� $�pT��46L��ّMJ��ܘ+h���ȓ'� �A�J!No���/Y�L ��Ho&���� ?4LptZ��A�؅ȓF]
	�6�)ɒ@�fծ;s���l��1��N�Vu6�;T�ÕX9$܆ȓbf��r�*.w�<#�b�P>��ȓ}ð<�'�;X���C�$]�H`�ȓ+Z)@޾d�Z�c�Aנ+g�]��,���� �4?�KS�["S̈́P�ȓe�L���Q���s��L����M�^ s�ۂ~"q�b�M�4#%�ȓ{�V< �@֊}ݎ�r��O�
Շ�	E�'R��4H ��nʙ34����'��`�)]��|:dɜ� �Z1��')���M�, y��c��=ӘH�	�'��X�1��^��qp��	�G[����'�<5X�A�CJ�9��Q?�`�M>���I��n�-�$JY(E���h@���{�!�Dȵ5�JUꅠV#	�| г�P�F�џ��IM�O�Ped��>)����j��`�'�\Y�"�#Md�)�d�X�yu����'gl�"AN��!R(�0F-F̴��']��c�  �lHL�O����	�'�����Q�HN��KI'>Jd�r�'a���"���/��9�E�0B�(�c	�'���  ���|iKSHC�8ͮ��ߓ��'�=�a�ÜO�n5�s �,%�Z���')�����Xc
�{F����e�'��ҷ#�z{�	���9i^@�
��� �0{���CK2- �2@m��٠"O�1E��'L%�ܰ�(�-o�"E	�"O��P� �$`mT�pqe
��Ԣ%"Op�����."� 8�D�v�1q�"Od ����+`��q��C�j=��"O �h2A3|V����ߣ��9Z�"O��K��5��{1�6�ҍ��"OPZQ	�ZR<�+�E�<����"OZ�ӣ��;m�P��oG*E��$�"O i�I�5|����-�/2x��kv"Oz��&�hŎ]r -��8<�+r"O ��%�S!Yf�)33���
n�9E"O���b h�t[��	
�d"O�-p ,\!WK��0��X���"Ot��J=t���ٸ�5R�"O�-��؟b�&H)�E	S�,�ʁ"O�Px�Ϝ�q��0��͋���	u"O.��2�o9č`,�"U�����"O�e*F�U��z������Z���"O<l�t$эmL8�?���5"O���U#y�H|���5	�,��"OP�s�!�� �ct�]/���(u"OR-�f�2���6Q�"�xRV�!�΄\A"xZa�lFLQ�'�i!� z��)��Mu���u�E!@f!�D��JbӆS1Z�={w�1
�$�4E{���MԈ+M��c�h��i6^�s�b
7�y�NS�1�N`����"c�fXbG��y��p7*�q9Y���Kt�K6��>��O��j��بr愽 �	;��d� �D�O>����#���j�Q���̀�y�!�G?¥���ו�$eIR+��-�!�d��@aC@CO�	���ˠ��?0������?E��[3R�-�4@�Un�"�C�yr(��i�6���+W�Pj|%�4�G��yB돣a�����a�	P��M�����hO���<M1|�	�	�-�h�i�Xg��`y�'�?qcÊ�u���7����h�AB-D�0馊B��>Y3�FI	R��@�0D�\��/� ���p@��3�(��.��1�Sܧ=�17��CҤ,@�HD�Y�����n�	�)�(k�T�3�	�/T��Wˀ����K����J�C������r~��2q���,n4�#��)�y�/�i���4�ǰ= �DI�nљ�yr`ǈS[
a�!ʰ#�li�s�F��y"cA%?,y��I9!��m� э�y2.ҏ=��ѥZ����@X��yO!`��e��8)��5P��$�y2��"����8Ì@�RL��?������'�7O�X���H7u��93�\!p? �iS"O����2�=�p�RS�<�2"O�1 �m٠T�B���(YnE���"O��e�	P����VED�>��P`"OԌ)���l�}����&N��d�b"O�UB��
Y�P9H��	\����"O��ԣ�k@6܈F〉 ��X�[��$�4��C���'C��]�B,$�@�^(d��`̞@�jC�LB��	nV�F�`تM�Qj�B䉅%�8�ԅ�9B�&hC@�S�LǊB�	/�D�P�޿9��S̱�XB�ɍ�*H��D������p�	v�B�I"YK@��	ٽ}�v���Q#5�B�I!o"d�']3tL����52x@�$�O:�"~�� �@�VoA�H`�@@��6�C�"O�("�>i��i@��;p���`"O���)65��1C�8�P�Q�"O���a�$�@K�õ%�*`c"O i2&��tl.�����R�a��"O�2KV�9�]k�^�dPj��"Or��Վ��Ԅ��v2�U�'�ў"~j'D	�gef�k#n'�[R���yrnͽq�ȁ�/�v����F��y��F�NY� ��� 0bM�ď)d��br���V艐�R�ER��=D�|Q2j�*O<�0¯_�TFB1�6D����牗G�t䱐(��9�����2D��i棗�@�y�W�M�PY���&2D����HG���Ɋ�>C�X���-D���E�^��LE2ǧC�Ir^�7�-D����A�Tr�K���B�2��R�*D� �1�ީXaP�qF��)+��ĩ�(D�D�2MƝ�������?2㎀�&:D�����37��/�5X��E�$�9D�,�4�	:�ab�6P"<�
#�6D�t%'ߐ
���C����0�Py���2D��1VEF�uvD��n�@!
Y�/D��R�$�<��ᦌ�Z���cb�.D�`���:ofdyХ�{m��1�h-D�|PQd�&��hE�7��0c1D���AIM�p{Hhؚ[��l1D� �V��Ib~=��
W�vFŘ�/4��HC��u�%[�Ma�tBpe۟���J4�	@��v񺌚d $`����M̓�qB���[����'V�<��2��TzGE�$|ҝ��#�=b�A�ȓ���p�]NVe�q���\�H�ȓ6�F=��]�j�`�A¾W@����Qg��U��8r�n8F�0��)Ζ�:4c�84>V��`�cJ�(�������I,%����d�KyR�b��/�C�IwsΨ���{�0�8u�'v$lC�U�rA�f �8=s���lH ��ȓ�����D�61*$��/͖]lp��b�zl�B
�#v����+a`Z`��2�E*V��.2İ�a�E�||pY�ȓBF@���+۴gE��2�O_w�|��>J6$��n�bV s�8Đ((D��)U���3��ݸ���8$&D C�%D�@`0d��~%��1��0!74���"D�Ĉ���B��)(�̅.����3D� Y�KI�\���(��W"���B1D���SlT!J��4(B/�a�0D� Y�([�8�A(	۠%<��[TJ+D�8�� ަch�i�F"/9PP��6D�� k�B`�<�E��FD���#�3D�@��KO2缌Z�MF��(�&D���Q��+Hqo^<��HʅZ!!�d�
6.*,��Ȁ�W�X��B+Z/!��C��:��lD>X���)[��!��#��4��c�8�t��F"E�!�dX�"ndz��T����R ��!��˂jG��z�'��`'�U�-ا��yቀv��\�5�Y�4:�PK�ذ+�~C�	,E� 3h�Q.�䲱�X�Y2�B�	 �hD��J'�|��$,�@�B�	���xV��*$l��V U�;�B�	��Be�6/^
(�R��Q,S�@� C�)� ���ğG�*c��� iu�x�P"O�a#��r�m� L�G|�xx�"O�Y�U�R3"��i`��s����"O�]��YS�L����N��@)v"Oޕ��Ȓ[�+NU�I�YQ�"O$��щ
)T.�c��08���#�"Oܠ�l�+Vj��6�ɹF.���"OX<�T'#!%����Ҋ1��\Hc"O`h�4i����mh���%vꬬ��"O<|Ƀ��D2�t�!��f��x1"OP�6"Z<['zԹ��LE�q�"Oj����,쭢��&B��I�"O����(7��]@����\s"OT���%*u���J�"�
R�<��"O.���)W�1���V�	�l���"O�������2Tda�O��B�Z��d"Oȉ�v��.����/ED�}X�'��xjvS��1�#�ǚ'>N���'!�钣��/U�H��v�R*�B8�'$|��J��H�� �%�D����~h<�c	��<�L�z��Y#YL<,���E��y�%]��R�0C�@jR����y2m�HK��kA���ZȪs�]����O���#LO��q�N�)F����ƞ
ƴ�0"O,��Uă��2�9RD�\�X|B�"O���2�_�E�*�a��y�hDP�"O���c(�3Z�<\r� Q�,ʹɫ�"OP)āF� �LR/V�w��Ph$"Ob����ZU,��l������S"O��i�C�*�Ը۴,J�/�t5�"O�̨��E�ޜ��e]*)�F\0"O�%��야(����e�o�4@9�"O��%��L���˧/f(1�"O4A�����6�x@��H�f���"OZ�9��|}�<���ҹ|�H�'���'�ڔHE�їR�"�-����'ML��C��X�B�0�a�#y��9�',����$Ҟ�S��v۪-�'/��9��4_&x�xDe�mA�X��'o�025͆W��-���['m��)Y�'%�8!�I��]{� d�M�
�'�´��IC5͂�����6H���?��
&X�gO0)��}�ŏ=���ȓWh�QHE���}1�	]=xCH��ȓ8v�U�_,k����BL�I�x���V��!�'����Ǎs\�H��j�j�_�7p�8$�]� �fY��x�0��㝌Q@8`�L{�n���M̓$TLu9gJ9;F�x�χ ��q��I<!`��|��`�E�ˆ=92	�)^�<ѧK(�l$�$lB�{�B,��N�X�<	���G��U�ul�>@�Ҁ�`-�R�<�*X%��ͫ�����@�f�<т��$U�����E�f���0�͙^�<�7���^1�
�`�U���\�'^�h�OhqX�Lϒ$��	�!D�8�-�
�'��x5V��#f�P�'j�@	�'ڬ����1Cp�|{u�#��Q���)�4K_�� ��bJ�
I��2d^��y�ؘB"�	�P� �P�u���9�'�$!BY�kaq��
u=�A��'4x�O�2V
[@�O�VS�����$6�'O�Jm���I�I~bT��!�x�vH�ȓD>"�Y�͗	�fl��Ώ�h��S�? ���2L�,��ș ;�Պ4"O���k���\���\�'X��w"O�a9�cĘ���&oU�>�2P"OR��$(�>4�h�vO���J�F"O��ۦ$֦&��Aq�B�z��E)�"O��q�T6/h��;�ެ6J<��"Ó�B�F�`�+k���P"O��8�D_�<nnI�U�L��Ч"O���@W�;���2u�O i�0��$"O���3���bQ�]I��4���:�"O"�#�ݠR� X���]5:�����"O�QB��S�!�������Ee��2�"O\���� �p�na"1# U
�qd"Op�!�̟Zh$�P�A�xE����"Ox=�`G �B@�2!ąC0��5"O�-uG���՘�2X%`ՙ�"Op���^(�P����T��j��"Ode�r��G�θh��[�M͠$�'"O�3P�υ.(���nO�����"O~}��5*\����ʎ{�F�X�"O(���P�0������,t�1�e"OR�#�Ί�?�����/.W�"Onp2H��o�T��8,LЬ��IQ>U����^P 8���>�Da�@6D���`.]�K��y��ȝ�!��z�5D��"�+��u���C��^���i4D��3�W�B��P�JM��b�a�%1D�8��p���1O	�tYT�RÎ,D�B�o�!Z>t� j	�>�2�tn?D�<kW��HL�a�l
)����H �O��	�xۂp�&[��Ndⳁˀr��C�	{�PpZ!�Li.TC��}?xC䉷R�ଲ#��h����5*0�B�I�qҩ֥@f��i�橃}�*C��-3#����F�Sx�����ޢ�:C䉶����ʠM�5C���,C�I+p>�y�nZ)�T!�r@�"F����:?f(w
f,�6� �~�J����IW�<��#�<��"R#4�6�C�NCP�<1'G��2 �R��8S�A3ǫ�J�<A@a�M�u00�C5���î|�<iEAP�O���@��}���I���u�<��IQ�'pd��u�O�iFC�s�<�P	�o�9�$Μ	x����͕o�<q���&7��hXd)�"�LT��IGm�<q͚#����7J��k{���g�l�<Y!� �P�&h�v�)�ν�P'�}�<�a߹�9;�	�~`�u�5o�<	�T�r��4�� ։xc@b�<�R�u���G晩Y�4�3GX�<�u��-L��)�eI�.�R���g�N�<�`��V Dȸ!�³_�6@��b_�<9%������ �	&�Q���R\�<	D�_0� �HU��?:�*��&@EV�<!6/
�ܢ�E��B� c�5��N��h�@h�7.�(DƝ�w7���ȓa��8�o�+t�U��F��B��(�ȓj�R9��مT>��A'�=NrT��[�Ą��0ƭPSi�^� ����l��h@�+�$t��·�1����ȓ�ty�̽'v����d�Ȍ��0��kT/&�<q1��^�Bt��ȓ�V�k6K۷��5��JuJ��ȓoў٠��0���Ǣ=��ф�S�? �-�fȁkl�T���Z�p�`k"Ol��)ޤWt�ਖ"Q�m}�%"O"�S#��"2��� E�'\<}Q�"O��I�,%:�@����U�"Of��g���P�ջ�(P�ƴ��"O��1����D�ԬsB.L�d���p"O���O,|,(�a��*��
�"Or��cB��`]�KE�eԐ��"OX�ic�>d: 
�i߽&e<��"O|,�%�K�LB�xgk-rc�� "O����/��M##��aK�y$"O�\3�"�4ঀs�JN�Bv���"O��@J ��#"I#t�,�A�"O�a�� ؾi܂���ؘ�V�X�"O�%�:�"Ż���9}h�3�"Or����A�Er |R4瘊bz���"O�(G+��0�X���=M��I:"Oz�rr㊿L�0x�^�<���"O����� 1k��
�Cѩ&/���"OްJ@�2{��]Iw�8*8�"O��	jU2�>��#�Ű!�.Y��Y��E{��IĔQx�zpN*S/��a�ŀ6yb�)�'<��p�c�OP��a[�
�	���'��h� F�S�����r�z�J
�'�~����^8٤��@�	z�`	�'!8�[sԩ<��L���;��Q��'�V��IN	618��6(('�:D��'�&���
W.�X��!�^	��'i�4x��0j����A�D���'��S��\f�P���
�$g���'��Q)��>0�F��Pc��'s$Q�'�L��b�� ��%�O�N�����'��12vKF�L#��4��A�s�'��鷅�^_ΑS1�F�4(%��'
�Z������i�c�H�'��2�+�>5G���eJăW�Z@2
�'sb����;3L���%+�!z���''�A%���(h���K���8�'c�yȅm�1��ei�n��Hw�B�'�r��d���*E��;� �'D>(H�'�0t+�	� �ܫ�☜5T�-��':�H�*P�x|�JA�Βd�]R�'D�9�Mv��(b�_�����'e�(A?V�Q�a��	��D�'H�y�WfOQS
�:!�0�: �'p�t F�����D����6_(B�'\۷D8���'��v�D9
�'ը��C��O� qjGd�%7b��	�'����=:"�*�ϫM���	�']4` Q!�A�
����UE�E�	�'��͹!�si����j��2 4p�'�&Q���"~��3��&�0-�
�'X�a����:�����F�d�
�'�H�CηMx���O�1|�z
�'���QO�_9A�a � ����'���ȑ9X0��U|N� ��'9���� �2�����so���'��-;��� ҆�:r.J�,A��'3�	[a���K@�L�80�d��'@`�{bH� �UH�ۭ)D�z�'Ӡ�۰�(O�h	x��$V�|9��'r�x� �լW�.Z�A�Cb|8�'YJ9c&g	K�D,�s��?�ִb�'�
���DS�v���I��_6x�=��� l��m�rnt`�!��a��#@"O\�C�X�}�~9"T�ȿ"XPU:�"O���,J��$B ���\�c�*O�!c�E�Qd4���J�b�d���'����єS���(͓Ѐ4D� ��
J.?\�	�� (<����7D��B���?���!�!�(	�t�4D�<��M�!1Y��iԠQ�;���"�6D�p0-�==C,� �Q�о9���.D����-
[)�6e�*;���pL+D�0["��4B�l���d��\0uC&D�H�4mܞ6���kC�L�(ҖXYB�6D����B% HХy�nֽ%�Jِ��5D��1"�Qf�SW��%�F�Z�(D���Ǣ^^�20��M�kl�]��('D����搨6��"gL֦V�89Ug#D�I��Ѽd�ڸaRO��1��Srn;D����$~����7��!$ԁ�C8D��ɧ�C�O(�@aO�a3�@u�2D�P��cP�,6����9�����<D��c�L�)):�g
:d(�*�C5D�ĸ���,����cH&j�0A���=D�0���@3�vq�e�²Y�aC�&)D�l0B%�VZ�{�e����%(D��ʆ_4#Ρ�'#7z"��'3D�,	4�ʪL��9C�F�\��w�+D���Cگ"���:�L�&/'`�T <D���w ��M<tZ2bW3o����&.D��aB��9ZA2�'�q-굸$�-D�(��(Ǐ����F덗C��9p��!D��(�!ǠK �2m�(��I[� D��ar�D+L�\j��=V�A�G>D�8�dJ0I2<zp�w�p�%k<D�4��د9���%^/�b]{�9D�D�
4����N�(U:��*D� ��Z�=&�h��V8Z��$��*D�b�(90	�W"Z1i����c(D�x�cc�zlH��e�p�*1D��H�-��mG�]�*,Y@D;`A!D�L� b �!�,�⅀Ffʈ�,D�8f�F�[�r��`C�$|���� *D��j���0gf
i�Q
7>Ђ�a 	<D�X�S�_4�nq0L�%�Xt�=D�D���4�J�X&��q�:D� �6�X�w���@���?,RD[Ƥ#D�@PM2-S&��ѫ=q�s��#D�`��)F�F�U�S�&6 3�!/D�X���?)�&C�H��Ib6�'D�H�Å�j!p�x#�UJ�-iu�&D��y�X,[���S.A02����%H1D�К5�ւ���(�J,^9�� Tj*D��;�GWyU4�{"gó1��!�&D���BT�S�n���+{D�X�Cj$D�T�0DȞIy�!�&I�`S� l,D�xp�O��X��a��+N-�nx�C+D����l� j�>�hȆ�lx�R�4D�LhU�H�P�d	EM
�\>9��G1D��ʔ�ʰ 8"e����$(�����"D�<1#�&��	�b��0n�����m+D����� �j��D��(��$D�,�gT8T�G�]�	����e�!D�p��2��9��B��e\f��� D��@1�ۙ	!�h7��Q`�ҕE*D����פER
��#V3k�:-z��(D�� f$�B
�rN��!��& ��D;�"O<���I�tS ����Һp�(�Ru*O��Q�M~M�Sp�G?(���' ԙkЫ�_������)=���;�'fft�5�ϑ@�&��N�l|�		�'6X�D^�G�Vq�Ė+e(@�
�'z�}p��i��xA�-U1q��d1�'�� �\�Z�����U����'|�����%F�8��U�yUn�3�'\����1T��xХ��[�|=�'�H��w(��o��<!�ŮOl�]�	�'�Ȳ���^� `���G"T��'8��(�#�.���uz��`�'� <��aٹov�)�@�Bޡ��'��H26��
/r0t
�e���4��'�.��-Ҹ3w�����T��*���7�����H��|�6��w�S�3ӎ��WĘ8���\���k�C����!�E2�m9#l8�t�3|���ȓ��}�$�O/I���!!5H���ȓV�l��T C+&��V+�'"Bl|�ȓIlၕ�Č5��y(�#1(e��R�x@36ņ'Op����Ƙc�rY��;�<1D�X0�Ψ�5��`h���xg��2��`��#��F���ȓ/�R :�#e&i8�߀��P��J|ҔrA�[&OD�h�@!&���>��� ��wW��5�V�K>��ȓE0�q�ż" �q��B��'�Y��j����b�@b�r􆉄�i���P�1R��Bc�O�0)��'P��B�݀dD�$�b���u�j2�'�.�17�I/g6�Z��J}�:���'ޜ~5ZEB�W�\gJ��'��y����Y��D�;"�ɨ�
�y�.�8�.��5�_���z� �y"�Q�r(j�۵�2e�f�`�����y�[�恻�H�,\�xY:uL��y2��X���@4m�6[��(�*��yB�U7X���!!�0`�rl�%g���y� Wn��b��B�[�>�a�+��y���X�/T>J�A�Ԅ�'�y�͉Q�X���=5�Ke�Z��y2hM�¸�a@�CED��)��y�C��B���IVBƄ:�B��̒
�y���. �\�YIt�a�H�K�fC�I�4��$�:F~��b��@�m�FC䉓^Z�1��B�E��t�U��(J��C�I"(ڼBD�[�Q����%�V3
C䉪9Ț�H���$e7��s�X�C��T��u���Y�����iƛH�B䉢&���`v'�] 2,�d��x��B�ɽ^��Ʌ,�Q����1m��(G!�� ��T���9���3K��v4!��U.X��ȣ�� Lаs��A�!�ɫC	z�r"�q&&�#G�E�!�ćTԈLk�M�|��2�f֔D�!򤛕$���r�L� ����EC!7!�d�Z��A�Dj�O]�X�f��i!�ĕ�y�0iж`!>%��h�E�V�!�>ȄP9t�[�LXd� JM3,�!�Ą {�dYx��O-��T��I�{
!���sbp��_�-ޚ@��g�n�!��F��-�a&O�*�H��6IQ1W�!�� *��� ��hŹr�"y�D	*"OV�f�&1c�����þ#l��bc"O\	1��8b��A�I��]k���"O|�rG��u�@���Ŷ	W|����,LO|�ѕ.V�,c�`����):��� ��'��m'�d�1L�+>`���F�Ιat+j'�yZ>��q��J���5#b�1���>�B@��]ǲ����t��?\J6����G�@���`$"O��Q6K4\�rl�#'�2��i�6a!�y�	/�g}�L3VbQ3AQ
N|��@�	��y2ɒ�d��Ѡ$�!ܰ �����	pX�L��7���Ui�h	�"&)�O�q���%.F&��=��
V�h�|�Dzr�'���y�G�#J�]����xײ���'L�;2�]�r���7〼k�"ɺ���6<OVm ����H!���t�|��v�d5�S�	�]w�h4�4><�Y%�X�{�!�֠3�2\QC��;�h#d�ڙ�!��,.
��c�+)u�荒��	�qs!��B�wLRX �
��e�j���ς�i���b��H���Ӡ��vri���- �P�v"OT��&j�<I���R��7�¹3p"O�%�*n���9��F;t�	0�"O�� q�G�����pgE����)U�iJ��D�9/]@աu��?)u�pO�,l!�J�0�(�ʎ�D������
�pP!� ]�tT@bK�-�Tѐ� �O�!�$�s}`��2.�&�r���2�!���!x��Z��B��$m�)�'�Q�x��	"��17�GheYRr�R	F>r#<i
�S�hˢ��Jd���B�*؆�c��l2�^1� uq�j؜rA=��6����C��d7R��/�?|�r�ȓ0H`�����T8�˺.GD���Z\���L�<]*tK�1!���ȓv�ab܎:
|�)cB�`����aȃ��-���b�?RŪ(��%?��Ji
@"�H��^iU�Ia<	$ h�es�M�#b1BUJT��a�<�$UH�Vy!�,�^�H��m�V�<�0�	�k� �����|3�q�d�L�<٦�I%Sn0	��G���%�TI�'�#:��fT��� ��1���:aɗG�<��c =َ���]� �����!�*=�S��M�T��N\�p���xPtQ� ��h�<Y��8qM^	!'+��T\��
�b�<)%���'�9X#	Ւi�� z��d�<�*�8RZ�����&���u��E�<!�ǕS�F���N@f��% �L�<A0��!)�䃶	\�*��x��B�'��yb�;i� -"��>Q���)�OR7�yB�EΜ�	�$��O^�-#RI\�ē�p>�!C�M�`�@�CP�wRH�H�g�z��hO�2S{ba�}���"��+��5A��U��?Y�'�2e(��O0����V**~� c��ޢ=)!�K53�����f�� ��,��<9�{b�'eB� CG�$4-�Wi�$z��'p�IRS�xF{J?%����4��`!^�
2LD��j4�Ih��ħ|�(�b��N�l7 �{��+��G{��'�r�q5,#	�֬1�%�^yћ'�qOf聉�i�?�т��Q��P�2�:R2	���0D�xB0振&v��dQ���s��c� ������x��s�� o(��fH3b��ʐ"One𠣊�xZ&�y�̑H�T��"O� ��9�ꕇ]8��3ƠN�?�~��"O��R#,�V�T����=bg�q��"O$��o��	���$X3(�\Q���V�'��ӵnUPe� ��5B��ӳ��{���U؟P�4��C�@�*t�T|�	�a D���<]��<�2�ε/	���S�<D��+Ӌ�����|'�H���A3n}�C�IhDV�'r�(� ��:h��hO�O	�� +r���q�ܭ
)p�Xu�G�Y�!�Ķ|6U��t�ĩ�#��|�x��˒ � $��y�����ybc��BY��	�Լ�3+.�y�K;uj�w��	0�H���n��yR�j�p�I�5hA�cB�y��H�Z�<����zOM�xA$��|�������ca�U����0M��m��X�"O�,���	��dcCb�gtPbA�	y�O��*�"�j\����74n~�
�'l�|�)�V9.�� ��y�p��'�ў"~�0�WXی�:�Ã&ɰȋ,IY�<!�CQ�Zؤ���ϔy�4ȳp�\�<�/)�"���V�x1ʥ;�c�V�<�ň,v��V�ż ~8��$�O�<w���!�zyf
���|��J�I�<1�ٛ>Щ�$�F*{�����+�E�<�4
7�t�k� �,u��P���j�<9pj	a�t�t���AM,�h1�[~�<��f�<QX��V�9s�Ҍ�U�<Af� �^��g���\!XDp`.DP�<�X/$�ZTa�K�(&���B��U�<A���.��$��9Ԓ�kTG�P�<�0FV�:���ڑ-C:�}DmPA�<���F>X�ɐ�C���e͑w�<є���,*�����>R"���r�<�SGM�{��9��ۼ	�BCfpy�'j� ��#V�"��fF�0G�b�{��>Q���'Dn��1��+U"�)�kE�'u�#�*��0�%�P?O��Dw�|bV�"~�rW\Az��ό���b���<}��
�L��`ʬ	2�]�[�D��'N�}�@��4r �g�JU�A+0϶��x��ڹa�(��A,g����NZ�kC���)��=�� Z� ���4�N4/���#�),O�T$�x��w����5�St��|����.����'��~�mZ8L��y1W�*k����d�(O>�q���J��4��0o�X��U+=D�l#� @bU4���C�5@u[֨:����������o��2��
aX����Iiy���MI�<s�!C�\�H�JaGm�듵��C��S��>����m� X����A� ������3��s�LC��"lD�!��I�X�� Z�,ړ�0<)�톯ag,���"Ok��)CS)MG�<y�Q2h
\��a�.[`-h���C؟\��Fh����
�+4�<�c��;\\��G{җ|���/rj�C�@�/5������!���>d��k�������ָ}�2�O��I}~��	ܖq�u�c,Z1<�1�!���#=�	ÓZ4�q���y��*�U���ӏ�D5O6�ڵE�~/D�A�OJTA�&�iʡ�ǚr/]0��=.�2qsTD�+k!��6���W��^�hpW��9iZ!�L<�nq{�a�)=���9��+�'Oўb?U��Z�ժD��S��c�Ǡ�l�O^ҧ�g��!zN��@*Y����ֈ�WS!��'7z� �hr�@U�K����(O�	PP0�4Ou�Չ�0O����I�	:Qr��=G'&�;$K̅Zp���	�M��%'�4e��q���l}��R%�׊"!���1$(t��㓈P��ߖd�O��3R��qyH4(���\�<���� ��`)s�^4!���U�\@�l��F~F��F��|�!���U ��/S?��:�e.Y.!��8t�@:�iνB�5�R�!��8�0�Y�Q2��Y�.ׅJ[!�X-jy���pDD9-ub�i�@ڐ#E!�d��Q`$�Ad�_xQ��90�!�DΗjԀ	�N1O�Lq� �J!��И)�a�4A���W�T�i!��a���+� s�,��y�!��ެg*���#S�P����E�!򤄦kG\�1��(gڶel\#KoJB�I�a�R���e�EP��#�d�7<B�84�$�� KHI�"A�#
� C�I+Wfl�ȴ�ߓ0�8���'N��C�����@�KɁK��"0���C�l�`	 &������(���ȓ��LI��F� M��q���+%b�U��ݦ��I�xH
��d��f�Մ���V��+��Y���C�c@TzD"O��!�J�f��;CN�.=�Y"O�tB��R/IF���D�+�mA��yj^/ K�鐣F[�5�b�  @��y"��0
�l1⋚�5	h@Q�C�0�y���I�y�X���*�O��y�o�!�pݙ*�>Q��Ia(�1�y ]6{���f��K��i��ֵ�yR .}Vq�Wf
$Y>r��G���yr��22�ehEkHz�<����A=�y���P[R!k��.lR��Rb��
�y҅�u^`A�.�(>ɱ	ɓ�y��Œ[FJ��B�;��Q�G��yB�U�l�pTK����:�����W3�y�&?�<��d�#��yHяF��y�G�4^�~h��I@ μQCBF	�y�?���EF��7`�!�J� ~@ŉ�A٬�0?���OF�ਘ�Qb��yI�(�x�<���|����
��,q�H�M�<u"�<^Q��f�)�d�h�q�<Y�����ű#i��&`�Y�adBQ�<��� Qg�1�`�Ιns�t ��K�<���F�F��DJ��r\����c�<	�Y'
�E��0�:�6�\�<��O�N��d`����3�Z�H"�^�<�F�F�P�;A�K9:2�9�US�<�6�Śl�^�����/D x���@�<GF�<��)���1[i\�3��VT�<��\)`s�ܲF�U;=�9�5�Q�<�阥<P�ӆ*���F"AI�<�$��![�L�
�[-�
y7Ň~�<���юXh�HC��P�:�[�<yFŖ��4%D ѻ.͚|BeN�{�<�ea�K<������g�&����Fs�<) ,S����Ó7/�Lq�ae
m�<Y�R�[����d�1��5�w�@U�<17k�'_,������Hi��C��[�<�����tڴ��bᰑ@T.V�<����25�F���%���ޤ�!#Q�<A�N���q�Y�Zv`�:��H�<���2���i���	+"8�7�O�<� V�S��t�űr��6v�mr�"O䵢���g��i��[WL�P��"O�I�UO��_xDh��ѻx8kb"O|Pb%,V=;� ��>�������xSڄ��'T':��T#=�0�I�$�:(k�=��)���:�.F-jHR@٠g��}����-ߩ��|��E��Oh��3�g����O�Y��H"O���JG�H=�$R1@[�6������ěc�b��t�#��>�v-�+Y|�=Z��XoD<sV��@x�0b���jRKfP��*! [�|1�XH��9u5X�%�?D���FC� Ĭ�R���$�v��3�:�d�1!�`���⛚�ȟL]Ya(�.䖌[�"�#d=h���"O�0 ��0���X���;v�*���́ED>�O�I �,�3}r��s�(��U ��*4I+��xBb�S��a� üi�$�v��2 ��hJ��H>���I+�����I.5�����(�N���	�6������N���DQ]�y���5,O�<�m�(z!�dƺ�%KsN��@@EB��M�1O�L`uE�O�b�*2/�74O��Z��ժ۴��c��n�<1�ʆE2(x���):���u��i�<Y�a��fB����R'W��#�M�<�נ��ƀ�t�W2%_�y3�*8D�8��i�>�:��ӝfS�ő1$3D��y��F�~���)@�xO@�!��=D��J��ݬ[`�����;_��ѣf@;D��!�	�(L�`��A�����9D��rD��^��uFP��؁C��7,O TB�,�ɯ,hڐ�狆3;�
=��nG�.C�I�k�`2�HT�𪶉�#��'����%͓I�S�'�\�3a�ǔM����Ɉ�I ���h��e`��)ǘL��/h�������Ó/��Ubs����LD�K�\ߘ��F�<��Bn�=��t�o) �a��	Z�)�~C�	�O�d��$�Ejx����K{���D�MW���yr�� ��h0`�B@3�뇧ߣ�y^ f����NܘAc��W-U���	83���;���i��5�sCO�=Kg8�j�MW*~�!�d ���*@>k,˰
Y�WױO6�b��5O�����	*~r,�K�K׀6�<Y�"OQy4Lm���#I�h(�xQ"O���вS\$�#���y"���P"O<A��셉kc�<8���� �"O�E�V�k����6,Q�%�J,�"O�t��(9)dP\r�lZ5OI�4�"O��0�b�"*�K�%�DmpŰ��>����	����?��f`Ʀ1�"5q��S��J.D���w�\_�\��GD�xq`�+e�k�I�yuj�%�.�3�	�I����ʌ0*����$ާX������*2���3,O�$�ˇ7��r�'C���8ņ^�{�~`@�)���?QM=hL��#�
R_�`-S1K�W~R�%4�J�J�R�أ��=W�0��%����JT�]y"��%٦ �T�8�y��F�G�����J\-Ld
��"J��i�hi�	X�*�������+�1�N?���� SPJ5�'�B�k�`BSQ���kF�x[N�
�-%�T9u�ܙ}|�C�Ցl�|`E�R �D壧@A&=�R	�6 N�Tc<%y�
��x���Yv�ڃ���B�d �@��dI��1�t�q,���"%��C��|a�43̚i��h8k�Ԭ[Vm�V~
D������V�'����-o϶I;0�M�3�6Y�aL\�S��V,��Ɯs/������O���V?��> ��C��Qe��X���A|8C��h���vHѕJVv�DhT\ƤA��k�I��֌M�T����쟲���I\n����U���E"f
TA��L<	6d��^>>[�{���'T��ͳsED!c����͋��ia��
f�������{ۨ�p�mQ�4ۨ�@1���-i��?1B
�Z\��``B��Fк���^^��3Z�髣��-����� �Z��E�1g��)%�ʕb��iZu$YH=�B�+�T9�9�(0".�^�QA����O��X�w@ك �
�@E�Q0m��+��z�	 bn1��� �Кq��+0 �[�A��_�b���*O��1��"�x@��]�sN�ڤȋ�നA�
�O���Ğ*��a���O��vMK��M�u��s����'0q`�GI��� �V�� �}��Ka��Y�`�U�tu��!���}�L�)�"�bCD�z�hB�H|=@��?A��)2TX]�����?٤���5�x�{���B�?)W�詃��D+�!�ȓ&&��&�0@B���� o lx`��*iz L>E��'��H�	R��Z�&�>Q��'�f,30�@�d�kg�7��4��'��[� �	�c��sCJM�l���C�#�O2(�)]�'N"��J�j[���V��0s
�',�Mh�ԀQd��א%��t��d[��F � !�O��icSH�.}-��C�����'���2��ݠZ�V��đ@HFi��������,eJ�D��"~2��=!$|`y�JC�&����0�yR�9v��С`����@b�}VĜ�Ie��9�;!��ȯ���8�)Q�y�jH�+J��S�L?�O��#�&?D�,9z�(ǷR�lxIF#���(4�G�D�xl��&�O̅���٧K
6�C�v�<�jC�ɬ7�đ���إO"f��w��S)0���%�B�c�V8
B䉊'��m{�ԇ/2����d�ҩh�	��$ZY��CX/D9aVj=��dQ���.]jja(a�
Z6Ruy��4D�,��%�'r�:�#��Mk(�"�CU3ZXFy2�ÿj8P���S�6Z��g�'e,�����,Cx ,Y!���=����D��I&FW7�HLʧ������� K��h��)ZyP\|`a��=��>9�6(t�h�K��+��蹅��H�'�6�3&ǋi\��
$P��b[>ѐC��1ɠ��B�Βb�A�wG"D��qb�;7gB=h���/���^�&�P�3�FՀQ�����hT�E��w
�HRg��i������<e$u
�'G�Tc�6�ތ�0��7�R��_�@5�yK!�L
?�CND���D�	8w8+��2U���2��-ٺ��dW	e�d��vm�����\i2���dK�8j��bA R
'�2� tcʽ��>i�P"4�bȓV��A�X`rT��N�'�n���	"@bh�ȇ��)>����X>5P�*I�v�l|�7G�c:
�҇�$D�@�U�2
����7/U�?�LP�4[F5��ύy�FA�SDh�4�~���.m��D5fd�"��D}��C�	�R�x1�1̈�	X<�q����P3����x�pa�1�:УQ��?�=�N�b�� �π����ErX�!pBˊg�ε{��21TI�Ǧ[��əg�YI�=3�!�t���qJ
 y�����-��B~�9�,+�f[��u��=R���ᦠӡ���;U��0�F��M!�q�wBL�9f�B�I�N%�yA	C#���"H�a���^��6T�q�ظY"����B)�0q�0a���7"��q�%D�8kr`K�;2��BnU(m�c#}��\*Q3(�$O�F8��8�����q�*Y�]��ɸP�'�H�0�(T^e��T_?$�*��ũ/�@a��JZ�)�"��/]#2�(po٠p���ȓ(4-3���-�ܤ ��P�y	zE��V�(���0z�	՟{M`�ȓ�������k؀�)Ej��R�D�ȓxi����KE!\>)�굆�eŤ�PR(Vc����y�4�ȓ��hʖ_ҡ�ԇ̟?�Յ��	"$쓌-h���(�A�����z�Ĵ���Ǫ�L�cvL'p|�ȓ6+6�i&�=�*��e쎕���ȓ\򴃒��&A����4���
� ��J��3���|�L5��I}���ȓ��ثTeZ���KD��mޡ�ȓ|����۶a�w�Vu�O��eǅ���䌩�Jt���BS�<��#�'�a~���kbF���!p��q��69�2�a�3_���=�T�GL>�( �'��E{�'O%<�뷀�g1� t	����^�ٺq�P5zo�X��"O� ڸ�%nBcΔ��E�K*��2��'�>9`���;NT�0��R�"~�BZ�9�^�$��!L�z4� ���y�-N61����.F��s`'W2��d�;?>  cO _������%Ag�K9�UF�a������ f��D
�ܸ������&�Q�H֌Dm-b�ik<�0�Ϝ���q�Õ����
�Z�'h2Ы�'�$>�t��P��zx��hR<QKR� ��G4z!��O��:4Dԑ=U�Hq�N3+X��GIP5��%e�)�F�� �GB�\����¥?U3
�'1 ږ ]�n�<kǥ��2є�k*Op���L�P�\{�)O�m�qt ���ҍXG��9��'X��ϓ�>��Dg��̀VK %;�! V�^(<�Ҋŵz������3W��aJ��SI�'�\T��I�/P��^qy',�pV,�jcAG�S�\L�E"O�<�@M41:��3��E*,C��h@"O<�ύx/8�� ,D��h0"O��Z���.�#@� �l5�p"O���hB�>3�F�!pm�Q"O����<=v���e�7u��C4"OP�@CO�i,H��b�cf�V"Of4P2m�5Xd(��1"�
���"O��@��9$�Ȑ%a��
�]ȗ"O�ѣ�bX�N |�����X��&"Oq)'�%�
�;���4S|X��3"O�`�		.k(0`���*{8�"O������K^T�
V�\]l`�C"O�xtǏTBK�j�)��'-�y��0�Jf
�f�vQA�O���y�ƅN���S�ݝC���:�B��y��G)���_FD0��Ǐ�yra�fA�a�%aON�\aq H��y��̞/��D��&�@2��AO��y�ο-�tٗ�߄Mv�(��^��y�⏞%:B]���)C~8˔$���yR,��b
��X`��(S`�*�3�y2�x�ҕ�fVB�Pe��&���y�A�uYސ�P���*�`�cƷ�y2l��V�ըM2�5(c��y�h�p{���a&	+�.�
�yrH�:'��)JR�� �!"�@��yr��3K��!ӓ��4O� ���Ű�y�N[�-R����
�	*%�-�/(�yR�՗3�)I��Q�Pvʈ� �#�y�i�>ȶ��Őgi��r���y� JZR��$� Y2�Tzu��y�B�2O�y�WdL�!���eH��yb�T�=�Y"7(��\��Z��y�D�����-3�ݰ�DS.�yF�"h�(�(�����ӵ蕐�y�KS&D���( ���,s�Ï?�yR(@�Z��w�E���������Py��j����8o�������g�<�K�*�.�bfD��_�Ja���U�<��O����1a^y�6%j�CW�<ADˋ".���������Q_Q�<y�䍜�Dh�r@���u�<�Dl�4^'���	�.�)_T�<V��`�>�¨� jӌ`�f��Q�<y�!��Ā��R�p�H���`�A�<u�,"�z+��@�"�H�a^K�<tO�0�� �6."
k<Ex@��I�<QW����*��"r��d�ŞK�<��
�3Z>����4���f�[_�<Y�Өf�H`���V�j�$���l�<� �q�����]5�a�D%̀cP� "OʘQ��9%)�e7w�0�r"O�����;�DK��+IPb�) "OԈrC��4����4�ͨC� ��"O��8�'Z*K&����ױ\��8u"O��� E�L!�؁0n���3�"O����K4`�Έ87L�����x�"OFL��`���AC�K/����C��O�p���1
çIm�`jA�3ڠ�#[7t���ȓr(�J�G'`�š����T�g`ҩ���Z�D��Od\����&��|�'V-A�8���O>�ô*\4:�����_�|�a���O��m�qA�˰>�F�48W����摱EӨ���Awx���E�P2@ܾ�:�[�DSF)�2OhΙ��ǅ�sT5���9D���ā�1�\8�k�Q�2��� ���8T�$��vk�=�ȟ���5b��W�L�k6��7v�8jr"O�HJC�A,M��Da�>D�53��N&3?d�O��3�$(�3}�M��\DХ*b��y%��0a��"��x�k��t2\� $8���R�I��@��C,&D��	�p�I�	��
X��˞�"o,��D���L��+ވ���.}���HE	V�);����)!�� �Ur�處,�$p���#ߔ<1O���$c�>
��G&No �m8�J4N�.� �_w�<�W�X/!������M�� cF�K�<�2;V��a��:C�����A�<�r+э�V��@F69�*u��~�<Qj	������iO�̖�,�C�I�0 ��<|Ռ�$t?�B�I�(1P�&�1'_r�Ao��n��B�	$]j�;F������X��� P"O��٠� y����+5A���t"O�C��O9a6�$-]^�=��"O&Y�����?\���ҭ��,^�1JG"O�P���V��d�u!��Pm���C"O��!sO�D*��k�Q�H�"O�Xw�K��v�adE�m[t�S"O>�a@8�~Q�����^��"O��b�45>PS�dT�y��3�"O��$��X� ��g��=
��T��"O~�&o�g��[��E�3��9"O~	�B�n�����DF�sԅp�"O�EK勝�i��9�g˵2>�!q"O�̛�iʈF������ J"O) ��F�i&q��L[%j�j��D"O��С�
�&͜0���l����"OV����"li
\Z+X�T����"Ojq��d�J�:��
:F�<�"O�ิ�H3P�h���o�(|2n�A"O4p���V�e�Y�G�ǀ0����>��ώ� c���?թG��n0вL>?�f�B�+-D�<'��,^hX`���vKR�i�ΊC�wOX�AՎ*�3托e82�z��!,l��Dd�5<M���ĕ�;����-O��q��C#o7��$��j�&�`��J�C̐(�cѮΰ?y�>*��o�D�j-���Y������	��z�k�>�G��~6}p��6�)��'�؅i2����#����O!�$U�1􂽣uYqf��*FH-V	co�;ZŚP�F\�d�����~" ���\�5��OUs&�U�F ���d>}�r��T�'8�I�gh�1 ��%�ֆI��xYю��AR%� ]�dy�Jϗ�Ơx�eѐK4#?Q`R�%��$�9�"��'Pf�'|mB0ϒ&�-���	:�,���i�i*Pf\�&�Du�@�X�A���Fi�-QR4�OΰH#��f¦\�\�����*"Kf\�9��1dY:|�"���M�6	��FEp����<��sޅC��+W�����]�� ��1D��!�(�8N� QF��47P��	N$�x��T�d���#�/���	V�L�.i�a�2=H!��O�|� P�mb���aNB�/���r�'�,��RhI�.ˎLI@� �T�g��N ��AmP5M�I7��|"h��AÊ�]�Ĉ�r��?9`c͸���2�l�XDdQ�ˑZ�K8l2�@G�w����Y�Y����t��"4n�	G���w�HI�IR�j
@��t卶S�� q�'�49x�H'e�^[�I��1��e�$��a�Y��D�f��(ބI��9�S�{ŏ�]ݬ�q���a�soF`�<�#V�Z�Z��3��Q��pƈ�>l�5�D�=�J (�O�f�|���X�N�Dx���Tmj1��y*1�C�����=��g�8N���b��b!) �4Z��;�ܸiQ>w�����Z�X�������e���K%I:
,������p�O�|9u.��:�N=�j�OPPa˗�����l��Q	�F��x����瘀X�!��X�]|��5�A�Wф�3�F?��=����!_��O?�I��Hi�`��|;��2E͈�w�ZC�ICe�\󃬞� xƵs� ������e�8�#�'w��o��Q=Ĺ�v���)d����'B������ 6�$���B2� <��'*�mabC�3P�A���B5�j	��'?�[�����(L� `�-u4%��'���*�[,m����RW�j�'�y�NDB H��wß=@�N͉�'�D*�hn�YWM�*l�l�
�'�@�ӂZ�'��Ԋ�Y�vD�`�
�'I����@ԝK$�mǀԠ5���J	�'ƌ��u�G���ѓ�[,���;�'�~�q����](�IQ!��1k�9�'�H���@%?�vp��@	�|k�E �'�pٲD��5�q A�u����'z��APO�!ׂpp&Ř�h���'%(²@V��!
P�o�3
�'� T�WH �-
�87F�K�n��p��JMށ$�:Ȱ��!M�8A��5�`Q�+$�#CC�����ȓD�<��/G.��(*7��Z�ȓY�=P5��|Ǆh�a��e X�ȓ?%е+�喃5���{ Ɖ��n�ȓf���&�
48^��H �x��/yA�P�t���Z��aʙ�ȓg]�J���pe�!Kg$��isf<�ȓE���bnFQ����%O�Lr��ȓ���5
����="�	:`�d�ȓ'Q��RABb>f幒���X� \��1�� oJ?!DʔQCoOg�f!��'���h�(<�4���+i2�K�'�Z[��1 �>��'��4	=�%��'u{$T�Z���8�N"<�����'2�j�b�&E��%I�
o�mj�'eƭ)�
Zx(e�����(�|��'�NX�JŹeװY�v��J�+;D���E��~�b�:���: |�y�7D�S&JT8�^�J$�N��d�d�&D�胇%ޛ�h#�<��8$J$D�����\�9�|xF앁��e���$D�H)5���}�$�����J�2>D�\����6k�]�2��.NJ�Ir��=D��z"+��k�
�8s��6|�"v6D�$&��
5���%�7ִM�Sh7D��z��-��P��
F�)�
/D�\��%CL��9!�q�f� �B/D�H!��ڛq��-
�ݧ\��t*O��K2'��GV���u��L�k"O%3qG�&+���(2�K�	�݉g"Ov��럴kj��&�Y����R"O����L�Fz�4H�`��^�L���"O��"U(��|y&T8�oyll��"O�)��B8/7p���7�����>钣Ol4	�	�S�? ����M�I�[3��*��]K �'Ӫ5�g�߆m�X˗B>[�$�Xv,ɔ�5Q��u(<)�
��H����ը2��8�Ću�'����Ƨn�)k%�I�u�����JP����EI '!��Y<�Й����,���f�I�⣋�p>x9!ȓ�-i�)�'�����$�"�0J��J���m[�')&���E5`����GM%qV&�S+O���G�67��q��-O���a"�5&�����8x��4��'��(@0E|��∦X�Y8��Ǻ4+P�Jӽ Ԛt��O⍸����o�y3�Ă�ED,����	6z$z$n��jن4�|rp��B�r̙�j�������.�q�<��F,{����(��0�@	j4
��Ȓ���H��aIӎ`y��	V�_���c&��>[Cl40B�N�<[^C䉥-���a���tn�)�ȏ�-^&˓^6���GԢ< �p��_0�1p��w(1!�j�oؔ���7mN���-AL@Pd����8jظ�1d���
OR���˃�H�p�!eDU"M��8��	:-�8ИTK]�'�\����)6����$荅ȓK��|��x�h�iů[�\��e���`�.��V �ͣ��Ӏ����g�" �Q�D
n�X����A�5��3�ȼ�GjïQ�Љs���%}mp���YxTd�we[�<J�),)
�X��3D��Br�¹�P(@$���*��ر�I<D�x��C	CP�4I��5k�*�c!D�|
B��.dlzEqA��� p��8D��Ұ��^H5öo�5 (��v�8D��ygG��q�ԧ�?�.H�0�7D�8�n�-8k�0��г6�
\[b4D���` H�8�FX��7�>-X@�5D�xӮ�
��j��K8���9D����	�!Ƞl'%��~y��b�	5D�d����:���ӢU�o���.6D� zw��c��h�%Q7B��A�V�4D��k`ݟjm�x( C�~��!� (D� ���Իc�QkW+�.�jukg�(D��q�Ϛ)J�P�1�R�~�,��'D��áD�"WL�7/Q�@����O>D���j�x����͑'����=D�j��0J��p���+�
�q�6D��Y`��6
IEp�e�=��P�0T�,��H��6)v�ZE���6��"O*U;q	�LZ�������a搑��"Od�P!	���ȱ�ޕ'��lj�"O�pK���2�cJ�&O&J�"O�!���8����5�U�"O��"k�Jd�Q
۳!��	�"O�|QQ$��V .4���:"�0��S�
�J�u��'?���ŌQ7&�f�
TM�%�����'j����O���`h�4�H�M���S�'�	yև�O�:\
�f �-|�=c�'׊��g�A�(+Fea�o�&$�}�
�'A�u�¥]�|<7#οI��
�'u�4C i[�h�l�`��3�UK�'W�I ��Im�Q���8�0m�
�'ԙ!��0g�� ze-�(?B��)�'�X�[��m�����<�P��'J�C#�wS^mp��4$@��'8X�:!��⽑�D�*�$U�'.���C��W���eY�(�2${���5OJ��RE�$�v�r�&H�p�P�$D�(O1��ap�f��I�
�ڷ��=�Y�V�x#�K?�S�O"zx��/�$����I%{Ǌ��'�b)Dy��4��7m�4����$���)J�}lӎ8(E�P�OL�X�ΓP>� ��CB͒�QǪU�2&Aٲ����ν$�.�I1آ��5�0|
�n1�Єa�,{�RqZ����~r(���d�ˆ��
,�)ҧNV6�Ʌ�[Vv%�C�ڡjP�do��4�rtc�j�.dwjX秨�(h��%3Vb4��K�ut��KV�¦@XX:sc��:��1@a��:MFF�H��R?l(`	da:�I�,�.��	��6�l�v��M�fm���5@�!��`XB	IP�ث��C!H߫.�!�_�9̌�#�4|Hш'Cp�!򄌏 H4�Q	S�k2P��D���P!�D�.(���0l�E���*���d;!򤗔U��P��[ d@��GE�"(!�d��v6d9bB#@R	2����'!򤔬Q����l(��a��'!�$����h �J�5
���ݖ�!�D :��X"�08��0J�%��}�!�$�lT����\;7��A�ꋰ%l!��:Z�� U��8.����Iߺ&p!�$�+ecpٹ��V:EC0XDC� ]z!�D\�zrb���Mo������5\!�d�&7��I#�!S��!���5=!��QUft����u|`�x�oS�$%!�DS�|W2!*E��Z]�U����8P!�d��u0����k�X��ر̆Q!��ӝS�����L'���jG�M!�R@����vF Kש[r�!��Q��ب Z��F�"y��	j�'rܨz�
Y�y�h����n�f���' �H�s"��q�@82b&�.+�9��'� a�sBt�Rcd���Ys�t��'���d�Y	N�Ã�ёE��iȠ"OƠRQAT�y�h�N1��"OV��ڛZG ��t��.�����"O�0	��K@X��$A>7��p�"O~@{�O�),�k����R�"O�W��dh���:�Cƭ�@�<!��Fɹ0O���A�%/B~�<�V�H>��jek]������v�<Qd�[;y��%�b՝s>00ˀ�t�<��D��p�6�#��&��w^J�<�Q<������$ HA%,@E�<ᆧ��8th���ϵ�J �f�<i�k�$lz�	)Q-ϵfʶ}I�Ε}�<���0]M���&�uI5�1�\y�<�ă�>C�T�b1\�d�0t��y�<)��]�S�vL k�!@��|3@�r�<����;3=�����p�t@W)�o�<��eޓV�"�A5���g^8����U�<!��|+�x���o�nP�.IH�<)��̎3��a*�����*]z�mUH�<aï�:ym���3,N���)���D�<�C�����3�eĭ"qX�Y%��X�<�V�/��h�搿	隀i�FW�<�p%�z�p��AP�)�UI0O�Q�<a�'O�[� �{ǧ�$/�D��RC�<!�C�G�p�B��k�PjW�i�<٤d	u�� ��j.%:Wc�i�<)�@�(\��s�?�]Ӗ��M�<��l�1_W8h"+-:��3�I�<B�]+�|�a�(@$l�GE�C�<y7C�&;50��n,oJ�p�%GI�<9�� M���µM^$e �0!G�<9���#ڽ�D�ݸr-6���@y�<Y�L&Lt��b�'�K����)^�<�1��8��D!��f��8���[Z�<� hz�؄<ꂥ�%�>]��ܚ&"O���ՂJp>$�P��]ߔ̨�"O�9�J&�΀�堙n+@��"Ope�6�ŕE�u`JF=U��Pg"O��;D	�>��ËA��a�"Ov��Gi"AY�3��V+h��eb�"O��d��`m�e� �0�X��%"O:���燽d7n�;P���ڪ�� "O4������_& h!�̢Y��"O�t ��׺q����L� ж0[$"O�a��Z�ay��Q�����q"O$�8qJ��~,8x�4E_�"��q�"O��r���FG�YC
���h�"O�-Y�EN�d �1ܧ7�n���"Od��k�1����)Q�:¾Q	"O� �5䖾4l�c�c�7����"O⩛'e�p��itHW<n��8 �"O(���/!�ah���n�6,��"O�\1 �`��sW)C:��"O�Hwݲa�Ń5p<T�"OaH�"�2hS���>R����"O���6CE�h���I���&Tc�PB�"Oހ;'$����0@�e��z�"O>@���lonib��W�.�l%��"OP����EPh��J�EIZĳu"O�eҳN�-[�PX��� �
�9"Ojq�Q��Hܩ�*�[|d]�`"O6a�/'q_z����/[G���2"O(싦�FAaİ�F�h2 ��'"O8�x�'w\�Mb7䖟b�:e(3"O�`�AS"r
>���#����Xʧ*O��Pނ����J���K
�' �á� ����;� I��'���EԦ�� ��׊$S���	�'� �`�.)`D#f�Ȃ����'�h�sᑐ@&l�JŬ@�\&��'����t�"|EO�t���'��qD�P\t�Y!�	�H�	�'NIZ�g� �4�������'DЄ�Ѭˁe�X�pF�g|ɘ�'�P �l\�5r�d[���-r8p
�'®�� Ć>�4�`��4�pL)�'>=Aǎ\�}I8mB5��}bH�
�'��8�2o�/+�
`�&�?y�a��'u�U�h�ܦ ��jÑ[��{�"Oh�۷�W#�i��	N�<���t"O��[��ռ{Ƙ+ G�{#�Ī
�'d���gL��8ʥ�ٽ���	�'mh���B�>l�ȁ?d�Y��'X��z�$�	� X��*w��3	�'`�cet��`	"�jp,��'��y�A�m��l�1Ȋ0i�H�'&�ʆbU�uB %jq��'u�B��
�'�T�c��&%ң@��kr�Q��'f��DU�8�`h$�9��8i�'�ʹ�2��!,�z��Ç��86
]#�'@Fىe'O�8��
�M�*����'g6��eӚX���ğ#)H��8�'`2P����rN������D٣
�'����i�6�$E;� �>���C�'�̱/֕<4:\{���r� 5�
�'�e@DO��T���'C�s&J��	�'�����C?~(�Y�i�f�0Q��'�� �A�7�M�k_ �4R��� (uB���~%�����T�ʰI�"Ot�+�#�K�`����^�]�@�
T"O��sk7b�9ӀIπٺ"O�x��"֗�	(��S�L�y3"O.�8D�_�\;0�;'�<7���"O�	Z��U���H�D�*��L$"O(UK%�U!Ft楁�c����12"O��*�摭{�>� �D��"�"Or���	F�m���a����"O��W� ��%	QJW.���[0"O K�e�*x�8�D'�1�p� "O��B��ĥ�&�*�C�D�	�e"O����/Q5u,�وUlv�~��"O�t�����6O8��AH�&���t"O�a�e�Rs5$��"��9)�>�@S"O�E�!�܍t-�	{���}z��3�"O�]Q�o�2_�~�
�%�a�ҥ@$"O��9R(�6�ؕpx���`"O(����]��T��S>i�ZD@�"Of���Rd�����+�"OYʤ�D)�.mӓ'�
����"O`��@	x1Y�&T�kv��3B"OʉP*ʝ>���%q^�"�"O��@�U�t���V�S�T���"O���4C�`�ݓ�I�\?N�"O�5����!dZ"5z��d"O|x���S%B�;!b�>]4���G"O��₆N/jlx1kt�ɽ1)�<�"O樀��Nj q�$$E��}*�"Oh��2 ?�Aӑ��,C@�F"O�0���]j��&ȔR�"�b"Oxt�ǁG!;�̌J�/8����W"Ot�	�@	6FҩH��>"��R�"O��
��w�!��L�$���"Or�x��K�B�a5	�P��"O����mM�R�\�0�j�H�|��"O\ԡ��
4;�j�)ޚ���"O���\�O,^��aȆ�\>��"O���4L ;�4FeHdq6"O�4q�f̱Ǵ�#掆��+n]q�<�Ǐ��RG�%{ � �������Lv�<QS��2�9�T�
�xK"��Q�r�<1�-��9]}�儉-7Kr�x���U�<��M�29\�r�ݫ�H����S�<��(Y�.|�cG
&Y�d�;!�IJ�<��̅�"�"�h �6C��%��C�D�<AYM���(B0kq0����?�!�D��l�
P�q@#
c��ҳl�4�!�\�)��B�$�9\H5���!���\�$ ���,�XU���Ѳ#�!�D�'J�"���ں{(�X�	҂�!��D�|��urcj��-��}��H��'�!���8N�|�s�䆦Q"��%�4�!�D��&�N- B��s�<hv�B+oQ!�����c<|4��ヒ�!�$T�W���H�"mF�Q��J�|�!�dDL�,�!Kcd�DH��!�DQ5=!���)��
.tع�#F{!�d�!���3J�q��$U;A�!��ݚ3h� �v�F�"��9gA*V�!�d�(�hUQ�-0	�j�˜zX!��U>X߾��Ɖ�"���QL׹`�!�$J`R��+?l�s7��"l1!��"�D� ;p#t0��I��:�!�� [��ſI�q���f�&�"Od0���7����aU2"w~H��"OB�ҏ�Z�A�I2��l�"OH�Ӱ���$�@�� d
�0s��cD"O�y�)՘i5��hFj�:�"O���ؠ&��Ȫv�O:��`pv"Or��n�+���Հ�0�"OL���?X��	+��+S"O��z!�P*e����j��݂��c"O�A�
�7h�@Ptj�2(�D �"O(�A��B:Kɨ,�eM�X����"O��ȁJ�|x�2ph��^E2#"O}0@@U�*�;EW�"
h3"O0��   ��>�2�'����WS^��g�47����A ��Ox�'��'��'u.EI�c�-2�"4��k�);B:���O�E�e�Ea6�BO������O�p��DG�0��RoͺLPdU��f�O����O@���O
�}R��V�N�P#�J%7t�1�cN�
� ��6����fFr�'��7�$�i��[5 #u<0����Y h�D�S�ee�0����ɌLz��nZS~Zw�D�[�՟Jt�QA�&��:!K� o�0(�-�Ī<i��?i��?�����1)L �{g.�Wq�iP2^�$�'.67ҳ|�����V�'a�O���/ � ���1>kL��	\�k���?Y���Şd�V,a%-A5[d�9#.^ߪ���Bл�M��_����c����6�ī<�'�fb�u-A�^$��-�?���?i���?�'��d�S��V�h�b$כ0k�T� T��$�jR����۴��'f���?!���?!5`ֶz�(���(a��|YQ�۰n�JU+�4��EX�V	��O�O�'.ȒGQ�+�{A�qju ��y��'�b�'R�'���	ѽ'��7�'0�dR�G��1���O���C��3[���/�M�H>A�B6��gl�4/߼�����$��'������A�h��曟0�*ۧ;v�ZW&ߪ٢=c���1
O����'q�&������'�"�'���[e�5u��Q�F^�8�z s �'��^��J�4_بΓ�?����	X�k��@ZF�J�O�H�#�/��Ƀ��$�Ŧ@ܴ?�����^�."�-;֋��q�xl��H��!��H0� Z�|�`�����&�2WO��!{�(C7 B*tn>�hT�<_���I��l�IΟ�)�Cy��aӬ�s���T�H��PC�G�֑K�ˆ�Y�����MK�2m�>���i�p!+�K�h��c����%kw�l�o�%dƎplT~k	h,���\��qAk��{<��cgZ� v:O���?���?����?�����ߦ+(�Au�#<r�1�T�Ƨ-0`�n�V5l������	~�s��i�����nZ�1nL �S%{s !�� 	�6�m��P%�b>�c��͓b߸���.4�2�	De�ER�I̓?��TR)�OQL>)*O�I�O���AIԘ;�����K�yb�O�$�O��$�<v�iEl�A�'���'�Ber������X D!�2kѐ ��O�e�'86�	ͦ�M<	rU�m�V���%ɥ)�VԁH�Q~"�KK��DRS
P��O��d��@��Y�6�z��I������Q
^�r�'���' ���c��nx.�(#m#_�n�����ҟ�K�4����'�6�=�i�i�3<pa���<��(v�X:�4n��oӼ�JG�y�z�x��/���J`-��x�a	v���2`b�,��A%�Ȗ��t�'��'B��'T��TGF�:�IQ
	'Arj�@vT� IٴH���?������<���ԧP	h�P�A���=!�-/gI����M��i/�O1���YQ��5���`VK�-O�E���U�����Zs;�{��5�O �L�ޭ�F�~d�8I�Lx`���?1��?��|�(O�nڨ|X�q��(j���;��M�w(D���.��ގ��I��M���>���?�;r.��Tl�7�B��#ˉ�{�(� �T�M��O�M�h݋��t���w7�=�FNR8 c�=�%Dou��B�'��'�b�'+b�'�N��NCH1�(v��<�Ju�wn�O>�D�O�AoZ�X���ǟh�ٴ����C@�Ь)4��㠣ٯ`xɫH>����?ͧ)�bSش�����chϦMx�ͣW�$��R�HY�3���Io��Xy��'l�'G�T�\�i�G1N�����-cR�'��	��M��eB��?����?�(��-J6+͗l$�ib�9a�h3@��,��OF�D�OԒO�S�rG�Q To��b�	J��	S�Y+�B�	wְo�)��4�Z���'��'DM�1���9���󉞼�D��'iB�'�r���O�剂�M��J$���J�Ä�%�| ���<"`@��?�0�i��O�D�'8���;�*!�U�EQ�t��Af�%	��'VN$��iR�iݙ����Xb)O�i�Rd�ܠM*f��5,�
�3ON��?���?��?������e��
�F�٪��!#�oڜ ���'qB����'!Z6=�d��P�T�}ux�E��+�f�A�O���7����-��7�n�$
�!�>Z�x�raڏ-BR=a�Kb��S@�̈́/�� �$�<9(O0�8�f�hB5J��<Z���#�'��6-̯�&���O(��ʗ�n��vQ/k������m����On��O�%��2!��<5�NA�p�0[$2!*��,?�Da�h��h+�4��Oʜ����?a2H f$ "�CP>mL��ʵԶ�?����?)��?�����Oy��/֜�! ���)�@�ë�O� n��-� ���`cܴ���y����R͘�R�OڠH���h4����y��'<"NiӜq!�jӐ�pJ�4��n�?� h��Xn���D���q,���?���<��D� a� x(�7s`^	 p�(+���:�M;,��?����?	��$
�N�H@P#�;%�Y���R�T�1ݛ�q��I'�b>a����|�Ȁ�bn���	h)�0���\>v	��_x���� �O�%I>�*O6�)�"��SqV-�2��b!;���O2���O����O�)�<�D�i�H����'N��ʵ��:5n=���I?\��`i��'��7m&��0���O����O�E� BD 
4�� 4�B]b�/��>Z7�.?uI�?v�8�SS�S��Z��0Ri��Z�K!:��L+�Nj���I;I��B]=5�h-��}h�����������MÒ�P��
o�
�O�hb�M2w4����/��1�"� I��韌�i>-�^Fb7m>?)P"�1}�x!Y���� F�I�oY#Zr��)�� %���'I�OY�A�F%<�X,3q�b ��F�I�M{B���?i���?a(����G�9$\Ī�fĎӘd������O��D�O��'��[��-��HF�a[��yV���m�H����עfm^LJ�4 ��i>Ys��O��O�����D�&#θˢ	�8c��b��O���O"�d�O1�l�Eݛ��Ob6 ��4�&@����L� &�|"&�'@�yӞ����OP���Sֈ`ȑ�ǀV�P嘒� _Gx��HƦ��E���Q�'D2�IF jz)Oise�ւs�"U�HB�=
��3Oh˓�?a��?i���?Q���򉂚P� ,���5Fx܅��M�>.x�xm�`���I�����D����I�������j��x�f�?i�Cq.�|��i�ڒO�O�މ�Ǵi�$� 5vL*E*�8.����k/U��Ǥ�\����v�D�O^��|����`��-X�����'�ב@?6����?��?�-On�o��#ZA�I���	�-
\��K�,-xCi�=TVh�?��V�ܛ�4����-�DU�b�����J�]�.a�CC�px�ɔd2�]�2�H�*�'?թ��'�*����:����ʙy�z-!E;���I�����Ο ��o�O�R�sY�uᘤW�.U�1k�!��v�����O`�������?�;i)*D�-N\�|
S�Ӎd�(ϓ���k��\l�b�j�no~R���E���h�p�rL�&ÜH��#
��țp�|Z���	���������Iៜ����Q�N(a$�M����!cyB�b�P�c��O�d�O�����>s���%Y
����ʬ"���'+��iVb�O�O�<��EGFx��3�ʇ�i���㮒�pd�)#S��k�$��H��L^�Isy"�J�a��kg�
��X�	ŋx���')B�'��Ot剮�M�� <�?W���ʌ"s��0a�C���?�ûio�OX��'���'�2�	�aT�x�����|,"bK{���ųi��	-q@��`�O�q�H�N�Ƽ��, ���J�g��D�O����O���O��d*�S�N?��e]#��L��!_5eL���'�rex�l!�=�V��Ϧu%�d+�C٢+4����ʳhQ�ٺ'�Uw��ӟ��i>u i@æ��'ۊ�Q�9�l�3ǆZ���͒�G��Sȅ��8sm�'�i>���ӟ�	(,��ܱ3�Q����b��V(/�:A�	؟��'��6��Xh���O~�d�|��
�}�Vp�MH��`�H}~�f�>����?�O>�OӠp���Ĝf�Z�@��6M�
�[����Ԩ��4�fm��!r��O�y��E�+07�#��nm�M��O�D�O �d�O1��\j�AM�T��l�C�-�A�`P+]A@�@E�'&R$c��pX�OB�l� 4Q�u��[�1z(�DN8O�>�S۴*��a�!����@�D��3�T�~���҉&����A�6Ge�T�7�X�<q*O���O��O�$�O��'!�֝�lD�mh��&o�=H8M` �i��8���'�b�'E�O�2Bk��.Ѧ[��5�b�!':�`��=hnZ�M#w�x��D)IM3�V6OVb%f��^G�ա�/4bɆXad5On�p�?��L(�d�<�'�?�QޛM�v���tm��raJ�?���?9���D���i�,B�<�	ߟ(kvl�pF]��@>:��a��s�l,���M�#�i��O\�ꀣ�#D�
#˵.��1@V��P	�M^&r[�1b�%��rS���8" oQ�T�|(����"	|(��B���I���I���F���'��@PlǬ�*��p� ��2a��'�6��l���ORAm�c�Ӽ˗b�]Z�<P�lԼQ�LPR���<ѳ�iʘ7�TĦ��%����'�"�@���?]��$�HO���'� w�6|r*X�bN�'��i>��Iן<��矈�����Ik��^ 2�k�@.pjy�'�6��12�t��O��D)�)�O�yU�W�Z�9�VMF<;v0-�֌�T}��iӤ�o'��ŞD~�����/�����B���01G��,,�l�'-\�`���P��|�_�0zv��3l�K�;z�P��A��B9d���O&���O��4���l�/�?�#�_�o0��z�˂�߲-�����?Q$�i+�O���'ü7^��ܴ���WC�'��]:"/�L����B�MC�O:���"?�b����w�~8���T���K1@�)<ԸS�'���'O��'�2�'��*�(W��y?���"��p����Oj�$�Ob�lZ *���'B��v�|�d]gޘb�U�z��D��K$O�$n��M�'�x�	�4��d�$N�� 
-�� ����Eo��brf��a!���?I1N;�d�<�'�?���?ys��=v��pyS��_���	lN��?������������(��쟈�O�$�HS�F� I�\H�,��'��XX�O @�'\��'�hO�i�O�}3�T�:L�i`��q4V4�4A�7?����u�ݖ'����i?�O>��V�n����.� �D}���W�?���?��?�|)Ob�l��:B|i$�E=��T�T듯{��@,�֟ �	0�Mۍ�	�>��~� ����� xY�)!Y�5�������%.x����`h���N�I�<�&�	�<i�nf�q�NV�<�(Oj���O��$�O����O�˧Bb*X)��Ѣ�P���#�*�Zf�i�RŰ��'��'��O�R�}��N' d��mG�u�H��Q����D�Or@$�b>�Q�K���ϓk栵��mR�o��P��U����xخ5 f���H%��'Sr�'��	g��'s����ǫ^�9���I3�'V��'��^�`޴E~�C��?y��sD@�Q� �AT�KQ�њ_]XEY�b�>Q���?YA�x2�A04h��a��hߪ��u�;��DoѰ<21Kd�x�%?a4�Od�V�-	�0c�e.OX�k�
��\6 ���Ov�d�O��2ڧ�?��n̺$@�x CM;&���W���?!@�i�Pj��'��h��杓>h�A0��2 <��͚~�,�I⟬���M�!S�M��OX �dm�?��4��.#�z��d�@/4�ʰ�4˯/Z�'���֟T�Iʟ��	�T�	�:wXlSH�5l@H�O7\נ��''F6�0���d�O���-�9O*�u$�4}!6(�%�0-��ԱÄ�N}�qӘ	o����S�'}���a��]'@�<�B�$k54��V
P�]i���'�j�P�,�⟼��|�\�`���F-6�@V�( "B) �ʟ����H��ڟ��{yfӄXBB�O,��(^�	?v��g�M�܍a��OHnN��~���ҟ8��䟈��±@��H� �6K.p�3]�|qx�nD~��tv���Sgܧ��S�lT j;p��4��8��G7���O@���O����O���7�S��U��!N~�Z�i2X���I䟨�I��MceN�|���P�V�|��љ�y*��S3�����F)�'�����iQ�u!�V���xt�D���L�L^a$R�)3 b����'���$�ĕ����'.2�'����#��(I�2����l2��'0rZ��hٴ,�,đ)Od�$�|�Տֆuxjћ�� Ojl���
y~�h�>���?yO>�OM�Ms �-)�n�c��8YH����d� �p�!�V���4�����qa�OJi�aK�"r\i�C�$]�N�@�O����O����O1��˓u��'B�i�e�$��2�aX~�U���'IBjq�6��ˬOZ�kظ�a����h-x�!4Z����O�0k��x���-f�) t����O�( ��$�
%y��+�L	����'H�I�L�I�X��ҟ\��o�d����� �_�7:��W�
,XP6�ڱu����O2��"���O�mz���Ԭlj�Q8E��RIʹ��П��	D�)�S�yL�Il�<i�A>Ô9хd�m?���ӪC�<�3L��TI|�D�����4�f��W&*���qnl��'�d�O��$�O�ʓb2�v�2?��'��+�f��J0�P�K�ćO��O@��'��'��'�\MSU �7qZ��gcE�f�D�r�O��KA�EH���@5����?5H�Or)&��?�t-@�.�6D��-R!��O����O
�d�OJ�}�;[�)B�@�v���4'z)���3<�f�����;�M3��wC�� ��2sL�s<�@��'�7��¦���4
n���ٴ����v�J���'d�-��H~�D��`�^�.แf;�ģ<ͧ�?���?!��?�I�9ܒH��м���be
����Dڦ����ky��'���c�Oڵ8g�;EM[0{~���d��{}��}�4o����Ş��!��\�<}��'��2+�@�ٶ+XS����'S�QbC��򟜣��|"\�X���ͽ!��=�h��!8�X��L}y��'R���]�,�۴���͓$�|�X�\�T���f�;��H͓S���DLP}RIl�,=n��M���? [��8`a�"�ql<��@޴��$A�Y�<��'��Ͽ�&b���v-�Aƀ*3j5XM��<��?����?�����ɀ%���Q�(��a1*�g'�Iʟ�ڴƦ��'y47m(���=`�\�cvd�6s���A��/
��'�T�ٴ���O�	�#�i�	�{�����-�+��q�$�L���O�"��Yw�Icy�OJ��'��#�9�޴��Ç+8<�+bN�L��'�	*�M�C��<����?/��4��Ɔ�-��Ÿ%�^9C��җ�0�O�o5�M�q�xʟ*ɠ�S�(<"g��-'�\�6M�\��ңu��i>�� �'��U'�4�ì7ybq�(_�{�z��V֟��	�x�	�b>�'C�6�M) �e�4�D����$F�i�Z�ۖ��O��D����?Z�4i�47x��!kVQm��j�J���@r��i6`7�B'�\6�*?��@�]i���<����BO1K��)J�&p�-���y�T�@����I՟����ėO�BB��S}�#��V�k����4�b���`b*�Ov���O���r���Ԧ�L ",Y���&ۖ�����j�@��d&�b>�*�f���S�? �h#7��u��5(��� �°�0O��!Ĉ��~��|]���	ԟ��pd��Ny�m�`��W�ʁb��]�����<��cy2/uӆ��j�O���O�e�PiԜM�Ts��� ��׃=�����d�OT��3�Dx�z�Q��:�pT���֪@D���ub2a2e�̦�PN~�t������i�ޡ�����0Dy���Б~=�!�����I��d�Io�O�"M��M�*A8C+,\t���� J��.tӐ@��OD�d榉�?�;zA�A���:v�(ᄏߒB����?q���?ar���Mk�O�N�C��S�g�0�7#[��T�H��S.l�� &���'�2�'b"�'�b�'�ʄ3"K�Hh��Ч[�w�z�õ^���ٴ6�����?����O���{%�έp��I�p�>C}�LS��>���?�K>�|�2�F�|��Œ0�Z&u[&(V�V�2��4nZ剰"ۚ�h��O&�OP�IV�����O9� ����2*��z��?���?	��|r-O��oZ�`3`Y�ɱ+�����Nֈ��t+<[��I�Mی��>���?1��S���˥e_2a&6٢1A�,
�|ծӸ�M#�O�(��������d�w{�����D<w8�:n�c���p�'�r�'�B�'U��'?�@}Ht�%(+�<q��(uȠ��s��O��d�O\\n1sw���ޟ�ڴ����%�q��|�9;����i �xrbb�>ulz>� ��Kܦ��'	��A����]��Ix��[,g�5��`�	,~��I�g��'�I�@�Iȟ �I�}�z�k@9v"���(/_�����͟4�'�7�������8�Im����Np
9�r#GX��E������J}�	qӲ�l����S��Lli$���lMD���ߌ�,d�T
t�8$�uP���!Rb�S�ɨ+�03�`�Z���X:�2T�I����	ɟ�)�Cy�nlӺ����58a�l�.PX(�� ʊLo����O��nZH�G��I��M�Qc�(~?�8�$nد��[Vj
8_7��g��i��q��|=�=�e.����,O:(§�޹��!�󫄻Z��['?O���?���?��?�����)�lX�(W�o�dAz-��n�lZ�w䨠������^�ퟠ����3ШD] �5@�&�~H��J ��i��O�OV����il�O��~Y`B�yJ���̡R�$GA'J-���i�Z�OB��?)��G� 2�J�A ���eԪS� �����?����?�-On\o��e  ���L�	(p�8�Y7�Y�e����2�� (�|��?�"T�d�Iɟ�'������H�PmJ�gK�w쭃��.?��l�"˪��4��ON�]���?�V�K�_.�9 @�#0i���?����?���h����PWȕ�bO(GL�!��E=t��T���Y��HIy��i�T��^�贂`,۝(Y�U���1��I3�M�0�i]�7-��r�h7-#?�"��Pg��I�G9L1�� �>�2k�*��/��XsL>A-O��O���O����O ���(��9+��Rg*��J$(Sg%�<�5�i��8��'�R�'���yb��1W�&	8e�!B4�`'Ծ7�,�
�& s���&�b>�[w��Fid����l�B�����<k��;?��	$�$�7�䓟򄊁}nq�QÃ�=-�|��e3(���ON���O��4��˓(�f�HWb㟴gA�"�D�A0�q��F4BAcӶ�4A�O�in��M�ѿif��f�@�f^��b�@X�kBz�C���g�����a��[����	��99'h�;h�0��6�"w�V�p4O�$�O�D�Ov�d�OD�?)��lT�r"��>T$+1�_3@^���OR�����9��By�}Ӹ�O���P���O0X�`m����V�L���M�ĳ����3��������@1l0�Q����A�����o��q�Ld��'\5'�p�����'B��'Eb�����IV�J�☪c����'o�V���ݴ\{�Ub��?	���i[�?$�<���ւX.-IBmJ�r�����D�O�6mKc�|�%�2-/|�J��	
ɘ��FAMP�)S �,�-��D�ן [R�|rFҶ0#���MҤlXhz�
�!yQB�'���'����U��0ݴ�,����(�"�طC2F����G(�?��W)�����N}��'�V�qvI�e�����A��N�+&�'�,���f��DGdY�#��d�~BFJ*���;F�ؒ7��'k�<�*O����O����O��$�O�˧d�8e	�[��\�HeJ+~�:��i1��#��'��'��O�R'g���
�r2�1g�����"ȎS,���O�O1��4��z���"J�p=�֏�R� �P��B���I�h�x�)��'?��%�������'윈EM�1� "gC_̞��6�'���' �]����4�@����?y��{e��"sn��@'�ds����B<�F�>!���?QL>��������B#31x<S��t~��F<f6��G���ߘO%���	�_UB��
$�@�p�]����Q�ZQr�'���'���ݟYƉ93�ˡ`@9H�ժ�ARҟ��ڴh�D8��?ᐽi��O�N�wu���SM�"辸x����<I��?���0�
)c�4��$��_���R��ru
��D�o)�:7�
J�X��Ɖ0�$�<ͧ�?i��?���?�G�Zt�P@@ �<�\]CA���̦��bȚ؟��IΟ4$?���8fkvA���"Ep9qc�2����O��d�O�O1���2� ���c׍v���"ō/)g���ǎ�U�	_�(c�'���&�4�'�t�Ői�����E�i�F�'I��'�����tW�D�ݴ4L�l���#�����͐��������2�Uț��d�v}��'�"�'(Y�7+�7���6�݇	=�xt��g+�6���8P��F�������A��Dֳ@��ؔ�Z�E�mQe5Of��O��$�O���O��?��C@̏1UL=pu��>6
�9�*�ܟ��������4@��ͧ�?�»i��'�V���͒�r���$˕u��Y��|"�'��O�^ݑ��i��I�U�d#���o4r�r��:����#�Բb?�#�o�Isy�OJ�'��&2L��� T�;�\��	�B2�'�I�Mۄ�J�<���?�)�l�!!H�.@�#w�|(@ ��X	�O�l���M�g�xʟ�d�ߜ(�R\Q�ex ��&�L�K��Qjӕ2�i>�Z��'
d�'���t��	� m0�_���a���I�����ϟ|���b>!�'�P7��:Qy�Djv�
�sʼ��S�J������8p�4��'W��N)�V�@����Z+Z��a��`ӧI6��h��Цe�'�M�4�Z�?]����qV  �/�~e��ʀ�4�*)؂7Oʓ��=��X3l��CF��3)~-R�
�vn�f�tb�'�r�i����@]�H�6ʞ�0�i�6LP����%�b>u�̦-͓8D켒�^G��q�فj��͓x 4e0�ﾟ%��'E�'��I��hS�Q�|EZ�l��d*&�'�b�'�B[�z�4O-r�`��?����X	!Ԯ�9[�Y�AA<Y��Y+����>!��?)J>��ǒ7a:d�@-�V���F	n~Z0ۺ��V���Oɸ����j�b⛒R�X���h�z�D���ɺh=��'���' ��ɟ�ZЩ��v*���T�_#������t��4GP��'�26;�i�}����&�h���k��>MмH%,h�l�ش��օoӊ1��'h���-|2��J�����3U����HD��ũSFK�h��O���|B���?1���?���/�v�1ԈJ�C��CwC�?���(O��n7{���ğ<�	a�s�\�D18^LS��F��Y������dRʦ�xܴW���O�:A�Q`Q-�>P�ņ=~�����C(�	��O$�y�m ��?ipc7���<���_jҥ�C�C�=���$ؓ�?����?���?ͧ��������i��S��]ƽ���V}�����f��Iݴ��'1v�Z��f�f��-oگ]�9b��DZ,�sA�L�w�,�g���I�'���$I��?e�}��;e�ʽ�����7��Z�g� R�Γ�?���?����?i���O�A�����f�Ed��f�����'X�'�F7픐s��S��M�N>��b�!��"�fS���ӱE�=*�'��7M_֦�7a.�oD~B��+xbqkw.å[bi�ӥS�Z�2h�ƥ���`��|�U�D�	���ß���l�>�܃g@ˏE �,H��۟8��yyR�w�H ���O��d�O��Rt�'� g���rCG�`��	��8�Iv�)JVˍ5�N��6�T�g��Fe��e�|X��%��;X!��t��B�|�j�/m >d����Y�!�.�2���'�R�'����W��;ش}`��5�Ш~PB����&��iY5e՛��d���=�?�Q�,�ڴ y^�Z Kр@��*��C�
x��i`7M:9�7�+?1 �� T��.��+G��DPꥤ��y�´�(���y�X�X��韘�	�L�	��d�O޴��0��!g;�v�r)ae� k��7m���p�D�O��D;�9O�lz�!TD^ز�VJFIl�A��"�?ٴE�ɧ�'+��9i�4�y�Z�l媜)3��X�Lܭ�y�ʴ2ψ��I���'��i>e�	G~Z�j  1p[(�;���)K6}���|������'�r6�*`�˓�?�t�R)~4�`	�m���	�ʚ&��'�~˓�?�޴�'G̐H���^���pb���U��i�Ox��Q!�N1I�R �?���Od�[�c^iݱ@$A�q��!
���O��$�O&�d�OP�}���	�y�ćS�\�� #�/cX\@��jH��Gc剘�M���wt:6E]�c�yQa��i2����'��i>n7�O<7R7M5?�qٴ�P��ұD_�$&��ژ�� �af.�AL>1-O���Oz�$�O����O쉸C`
RR}�r��=6��m`�μ<9��i�4 x��'�"�'��O�R�,7�FeK��HB0���B�?}�$��?���S�'>���!p�ړ1�v�*�D�?TE@``Ʈ�M�R���@,<L�a��J~΢�P%�8���i�e����a"+"GU8]�f�	�t}�t�*0�:q�Ѣ`�����J�(�:�p1-�5h�1;��º_(.8y/�ǟ,Ζ�>R��j_?u���g�.�I0]�*�qTꜯSj�h���:l̼s�.�I����!�}1r!gD�pt��S�J=�	q_'^�)�� G$�\�@>$e����$�21`1eC#\�U�"�ON$�F����A�5s* ���4gx��q�:���2���i.�����,��YR�+�v ��E�(��a���l��CV�L�B6��<�����OB���O�Ģ`l�O�[`��#��Y���;W�}j�,B]}��'%2�'��0r��[��(�$��Br`���� '�:E	���$%�rYm�8$���I��J���gܓJ��
3@����j�+=u��n��4�Iay�L�Ib���?Q��RU�ަJ4d�[����\��\@è���'���'z�P�G�Ĥ?� PY2W(H�I�hʦ��m�����i��I
�J�s۴�?��y�'m�i�-��N�/������%?���)�
q���d�O��Cd�O^�O��>%y��ك#�NE� I]�l��4b�nӞ@�bD 馱���@��?);�O|�g��%1��2t��%ˑ�8a��h��i��T8���$�SǟLH�IОFK�=�2b#[߀�	B˛��M���?i�'_�}�a^�8�'��O�CEN1�N�p�J@(����i��'Ȇ��G	<���O0���O�Pa�S�kO����nޫ[!bT@ek\�q�^���`�O���?�H>��J��0�J��*��C7�� �J��'@�#��|2�'\"�'<��8ϴm�R�ńXŠp�A�_�u�8�diۤ��$�<9����?1����R��J� H���R�O�Z�< vhֹ���?	��?(Oj|���|���	�.����ː�Sf�1�c	��!�'��|��'�֢^��T�d�����ȅo��mRNJ�E���ğ���ן(�'��|�p��~r�d�X!iq��F��q��}�����i�|b�'�ҌX:qO���fd��,xl8 B&����M+���?�*ON=�q�|����y�'Jk T�@�	n��U.Ѿ~�1{��x��'����:.�O�S�`�T�@�i��_���:S�5&�6��<�����c�6��~������X#�ϕ�zw00S���2 <�V��M�/O���O:8'>��O6��;t��$:0j��L%����!ݛ���i�R�'C��O'FO�)�n^�A��ėdS2E�@�Yo�ƁmZ
n��-���8�'�����ڑ4ۘ@�-;.׬��$��2�o���I��w� Cyʟ��'a���B]!>���`�3`&��I"�I$r��9����'<��Ց�0HN�hb$-RV*���'!B�kfP��R���⟠��F�-�	צJ4L&	�����g��'�B�'2T��z�Z&T�~DѲeÙbX�4 .4~���YM<I���?�����O ��2K�b<@si�.y�:��4�����7-�Ot��?����?�-OTaÇ��|2A���7܈�0MޤB1�Px���x}��'���|�V�|R�IܟD�%iI @�xv��T0t�I0�U>��$�O"�d�O�˓"Ѱ���T�,_,�h�F�[s6����Q�b6��O��D�<���?�ˍ��?�I?9���7��$J��C!=�tGw�F���<���?{zUq+�����On��Ƹ��樏U�(��e�t� �xR�'b��'��y��X�C���Y:��Pe���T	0�( ]�������X��՟Ȕ'��tY���P��h8r��2�X�p�^�T�d7��O,�d�$0%f��)��j�<P;nR�yM��𤃓3����K�jHr�'��'���T��'j�*lq� �6a|3v!G���MAйi�<���c������d$���e�b��S��āY�nC˦���Ꞔ���P8�i���i=}"�P&З`�lD̉R1+N,q=�b��ȴ���'�?����?a��յe�L8[��	)Ά bch�~���'���I���>�/O4�$�<���cF�ŬpH��SC�ǭl羉�E������2;�����8��ş�IޟX�'� |B��̡�jś�TT��+�%�ꓤ�$�Ol��?���?9�'	xx�׮�2/� �"TC�^����$�O��D�O��(��qp�<�΁��	��6@�E��(΀}�R1鵱i��	Ɵ��'���'r*��y򭓭^0��RC�=\y�Yi-
�5\���?���?�*O�EJ�+�w�T�'_0�x�� @ s���Gh H��}���d�<1���?��[p\�ϓ��i2����I�ـ��[�:�Y�4�?	����d�����O<B�'3�4B�N"�i�A��%Hu�k�R�<����?����?�i��<1���?���]���`�ٗL���$q� ʓ} `�r�i[��'���O��Ӻ;�h�=
G�|�uM֬@,����Ԧ��	ޟ��A�m��	jy�I/��
A�K��;F,�'6�v��C�&6��O����ON��	D}r\���aO3>��(H4��S |m�Enޢ�M�"��<Q����9�S��S$����R��X�-sR���M����?!��m���6^���'�R�OxLj�Ň<#�,#te�z��ҡ�ih�W��R�@w���?q���?a�L�i�>�	b��#8��c�%��1_�&�'��h��k�>Y+O ���<Q����֌71�U���P6`���Ċh}Ҁ��yr�'���'A��'f�	@���a���Z�(,�󦗆 �������d�<)����D�O6���O�0�eڏ3�r�i�R�h�����_�$�O$�$�OV��O`��1A5�X�2�n�:I�x�����0��)�i����ȕ'�B�'��nZ1�yr.��8T�P�B�j�p�F�#$��7M�O0�$�O����<�CJ�AK�S���P��.[��l��`W�o��C���M����d�O���Od�i48O��禍r�7O*@a��X�ȀU"%�{�F�D�O�ʓ5o�ygR?��I�l�Ӆ?�"@E�.YWҩ��&Q��X�Ov�d�O2��4&����'�f �gӟ#�(�W�V� �fem�Ly�+O*"|,7��Ot�D�O��Pe}Zw\��&��;g���E�شGR$��4�?�C�B���?1,O��>����O9t���Y)���Gք�M+�LW� x���'�"�'���k�>�-Oh�yPA�^�L͂:7����������{���	Uy���O�8� ���!I��+vPc�4v������i��'����>�V듫��O����`��j` *~��u8ӈ�"6o�6-�O�-�D�S���'��'����J5��!��Bk�0l��`l���dÒK2l]�'�ޟ��'Zc�����NM�C��÷�۫|�Ұ3�OF�6OT���O����O��d�<14��/m���Ҁ����+�H����V�ؔ'h�^���Iϟ����T!0��gC
;6eh7�mXi���w���	Ɵ\��۟0��Ny�+́E�~��y��sG���Rz��*V�ץ!8"6-�<�����O*�D�O8�h63O�$�c@�����MR�3�H���æ���ߟ��Iܟ�'��=٦G�~z�x<Y଎�73���7�C�O��[��ij�W�������	���A�D�c��$�~�3&�H&(�n��|�	xyZW��� L|
���vͦ%��E:��^�<�Ͳ��R�
l��џ���͟��.�ҟ%�P�����g��9~���a�hQ o�\pm�|y�e)F^6MW��'��d* ?i"j��vꞍKS�ô9�
��aC�ɦI�����"B�&�t�����,m�ʄڱ�Si�$��6.�4k�v\P�07-�O����O~���f��ȟx��h�,%^%@�I�6Yj�P��J;�M���];�?�N>ً���'G��B5ׄdDH	%m��xxn�b��tӶ���O��*Y�$�&�L�I����eJ.�Pb�"c���n8��oZE�Qg�HqO|R��?1�'��L"*vP����.���c�iV���, ��b����`�i�-�qn!�z4XB�Ń~WI��J�>qb@�<�*O���Ox��R�f�8K�<�;��^L���VH[*l&�'� ���&�$���\1F)9�|��V�v��$dđ)Z���Wy"�'���DJ�P�S�;pP�:�A�
I a��ɋ�Z�듅?A����?I��Df�%Γ;(��AV��Cg��(t��W���Iӟ|��Vy������i"a��1p����ޡl?�Mx��Gͦ}�IJ�	ϟx��
����=Y�j5�����苞H�
�{Q��Ȧi���x�'��b5�:�)�O��i�+V�����{HQc!L�mլa$���	؟\�T(Bꟼ'�\�'O��,�Q�
��Α �!�/BIl�_y �Dp6�D��'���k'?�E��?g0%��G�i��)S�ڦU���4s�,��'���O��D�1:܌�����(�D�Q GEV���&9$�7��O�D�O&�����͟���"ޢ6�t�dH�i,,�2�!	��M��m̀�?�N>Q����'��,���hv ���%00A��p� �$�O���M���&��K�P'�
��4&C�Y$A���%*����'��	�>��L|���?����ԩSP��qr,21%�1*|~,��i�j�EΠO�i=�T#�2�M�!��<1$ ��R7���'�|�[�'��I�l�	ԟ��'� (����<$'NP�d	�=
��)%�B�XdHO�d*��?�6]�����Ǡv���Tm�J �y���?i��?i���?.O"�a���|$)T.~�zE��.Q��H�u}��'�ў����5�Q���\��У�h@�v�Z\xm��*	2ٰ�O&�D�O��<i�%��O��5��'^�h��)V[�\@8�5�d�z�=���V�݃����OxT,�FF��#S����BB�$H6M�O��D�OX��I,D�����O����O��	�
����55P��J��K{�E$�8�I�����n��dc��'R��]��/�(��2m֘E`�aoyyR"�hx�6��O���O��	�X}ZcMx��Ț$Q^�|:c)S�4�u�M<�������'����>�B�m�:A9!�;��B��]�QIƢ��0�	ҟ��	�?��'L�S.Z��Ӧ�*
&��ϟ�E�b�ܴpH���.[\�S�O\BK�e�n�hu�Ȼ	�a���Gؤ6m�O��D�O6X)�DԦi�IΟ ��ޟ��i����YW8�$:4hˠ0�֥ `A}���O ��3O����IJ
b�0g�TؒP	���B��A�Ɍ{�h�@�4�?a���?��H��t?���%;���1G�X<?���Cn}�b��y�T����ٟ��ҟt�I�>��8bu�	�o&X��l�)�t������MK���?���?1�Z?1�'}�Q�|.�hS����n���ؑA4�D��'��' ��'n�Q�$��G�����شBP����/G*.�&�
P�Ŵ�M�.O��$�<���?I��)�����-ՒO�&�C�.9ul�������	ȟH��ݟ��꟨)�*���M����?	�ě�?��l����b�Z�[V�UU���'B�'4��ǟT��c>���j?�L[�b(`S4Ş>c~�6&��)�I՟���ϟ�9.��M����?���RB�Mt�I���A(� �2ě��'��	ٟ�h�dk>y�����Mk
��B&@)4.�Ur ��q�����ğL�hN�M���?����
�'�?����\�A��,�!9���2.]=��	�� �������ny�O��'O�Ȱ2%��i1�6��'�h�n�@	��"�4�?1���?��'%��{yCF
fhMk�c��!� ���b�'v`7�,�$�OPʓ���Q!ӡb%�bQ��[ 퐢㗆g�.�Ɠ��-I�����a�*^RI���	Tp4���9��`��b8�oE�hH�sP+YM���P��<���.���T.�,��5H����i�݁�g��v���jdJ�4��Š��C��hQ``�]�L���-_p�Fdj���!mX�Z�4�C����n4�!�$�f�;� ��� u�I��Z�u���2���Ol���O��I8)����O
�SB�Z�� C�	��tlX�fD�M$^�T��R硇�{�Z�k���Oj�GJ!R�\3�$
K �D�ĦY�7	�0��D�
)P���F$rDmG~�ќ�?��U��i��#�"o$*l����W�N،�3��]6�^�M�f�:2S'�Hp�ȓw�rlx���8^,Q
�Nm�\�H��Ify��9.� ��?�,�^"����)t��T������똇\N���i5���d��\s��Y2˖�����O�S�^����H�� Y�-ʡ'���<�p�i�Pi���Y�<� �`M|�cI�CV<�;D�6BR����q�'̪���?���t��F#.��E.�<������
�yR�'���df]Y��5pV�
O�DHk���'i|\��_���E���DD~X�'����I�>����I�V����O�d�(�64XC��z�CBh�_r��H��T���ˢ�Jt��|:���v��y�VC�@@T�ⰣOq�$a(�*YZX�sgBѾ>U8tad����"�֬G�Ps�gC�%�Xy���qbb�z��'Mr����&�O��� b��Peܵ�`�������"O�����N1	���U-gN�c�	��HO�SZ�t��d�}�Rܻ�fעo�~m������R�O�3�v)��П�����Գ[w���'�jMsꁟ����� �81��J�O�D��486��b�������::r�=3��&?M��PcG%4\0���9x���!�%>^�s�՟%��l���'��j��Ae�"��@�F���'
�(�����=�f�T(^0�
E��Z����S�<�B���4;���r�<m�P	Inґ�"~Γ��kc��� ��q�&�8 �ȓ�88��)K�B��J96�������d�Ԭ;��d��2�z$�ȓF�3"��!I�4�`R�b�=��dk��1�CC,1O�|��E�
���P܎�h�h�j^Mb��ͷf�*��ȓ+�,�҅D8'��l����&��1�ȓ���Yc�F�Nz(qq�U|���}V��{���6XzQ r�JM6	��#�����HI �Z`gS���ȓ!#.T���e��@��?H����DCԹ�S&#�` ��>o�8\��N�}x�	�$R ��S��"{T���J����7B�l��U3PB�7o����_X��rǫ��Y3��jF�@h���h��L��%V����$�U&����2TgW�8����L��f�ȓ��Y!�BJ/�lj⠞*x��ȓ���B���$��{�Ĕ>n�dt�ȓ`�8�`�\�U58�3�⛞T)⩄� >xR����Np��p%�0+���/���Z/r��«�T/�m�ȓ�Ń!�FV$N�`3o�r�$��3<�Pjw�\?v��pD�E�<���A�+�vP��X�V��%�O~�<tA_��АېN�T�p�2�z�<QmISj�iE�����!���A�<)V��A��}r$Z�`o<���z�<�`���Y�̑
FH�?l�I;��Ey�<�TI�Y7���%�Ua�ʖ��o�<��VxD��T(�?�q�t��n�<aK�i���\>ODL�9�g�<��˙�#>D��	����G�a�<!���ݸa�EG�8R�8i��_�'�H �Q�4��OP,yspΔ�6��i�W����UZ�'w�����#�vLS�kH��f���'��<�5c��YKɧh���OH�%���	6�C����"O����D5D*�{�M��/b��4�>1w��.;W�˓l�R��aA�a��e��? Hه�	
V���
�^3�8HP�Y�Ԥ�=v��e�ē����v-֢r���aTbԱ?�D(F}rl�i�rj'�� 
-�JPy��P�Q�g��iQ�"O��S�ДNٲ��ɧI�J��O�T�M\�d@1O�>�rpJ
;%˖�طm�����fH-D������Ai\,)1T�Yt��A��7D����֍3*8�ҹo�حu�*D����8(BP��Q���I)`�5D��H�C�|X��/q���ȴc>D������#U��r���	{Ѻq��E>D�$
DgB�F�kw��]���x�K:D�$��(\{Wb9����bC�ԙv�;D��Jv��3[���s��aѪ|{a";D��ڄ��2q�P�Y�F�P^p��$�;D�4ÉSKZY)���)z�6X�CH9D� �%���'Ϭ����w�����a8D�x� E]�`J �B���:.T��"8D�P ���.I�l ���_; �q⦯(D�����|1a$nʚ)r��U�$D���c���J��aG�@�l8�?D�T8S/͹l^�j&�E�/ʜD1�<D�,�6M�K���c��ǎp(��&D�ps�Ě!@�:���8r���):D���!�MCl�(ӣk5C-J��Q,+D�l�E��nL놌��f�[��>D��h���[��� �/��m��ۀA;D�вKЊ6Bfls���/y�VU�!�8D������m8@	�&@�]O��Ib##D�d�S���Q�$A m��!t#D��qTBBEn�񶀞(�4��$ D�|��'��"��qj�엄��f�(D�t�poC:3�`��I"�:���1D����
V+_yt��	@���F(1D��*P��]��;�(�.[�0��-D��Q��LXs�	�a�u��H��H*D�8x%i���̚�(H2*Rx��,D��q��k�$�!�N�QS<�� +D�HP�͘
V�\JƊ��oE�ڶ,,D��8q�;]
��B��!�̹�!O(D�l�'J��7�x�XW N�-�ܸ+#�#D�Pj���'G��D8��͇B����i>D�83h�8$��E$˳,B��r4=D�\�������8פ�6�6D����` <-�\m��O=�pi�N/D�`rg@�y r,��GO��IR�//D�$�A
�A�:9�t���$���- D�t[f��}hi��m�!'sP���2D������2K5�(p�UWSpEɷ�5D�����7�N�"5H�QO$�Ȗf2D��Af��>�a��
�����*}�"5X��6�8.��?�` �B>`������Ҭ$�6#D�,�c��KZe�GK�${��0:�
�n�&�'촐��\��Ϙ'�������{18,����vGȡ;�' ���^#4������0pc�p�B P@ �4@��N)<F�3.��0=	��#V>����L�}��j\���ޏp��E�s䚥7�`����� y��ȁ�f
V��h)��ܙ���Ɠ4�B�RA�^�_�����U8��H�'Q~X���[/7!��0�)T�p�Q��t��P��@���f1��x�%\�lb�q��X�x�bf��4��� $N�J)������MPv��R���� ��B�S�Y$�'HHiWo«r\���N�o6p��N���fUS���G�
%L�[֪��wuV2�S4���VΌ�m�󄗰���yD��"Q�@X���_�8Y���
�f�*���J�G<����G@� _h�)�!%e��J�$ߖRZ���Oƀ���Q��тΛe�d!x]�� phH�v�^-�#��@	�҉�ئ�?��λ� hѠI�6#���I�8D�8�� ̹!#"�4|��o���@�4n��?A��P8F�x@N>� ��H��ΗfK������ ��C�'��J��ºm��:@L= *
�Z ��:Pߨ��@R�c� ��ȉE�����C�� I�I+��X"�l��m�ax�X27�zXJ��
���lH�)@�:>�#�O�&��K�*ТOpJ���O�92OÝJ*4�zr��9"��0���hj��B��P̔�UÎ��t��j�O�R�Y��Ȋ!�d��C�8����')ҭ�B� �s��*sAO<�<d;P�F,ay3)�v������S��?�F���y�CܭB6.�Qr���b����!Ƥ��O
غ�N�b��'bnxG%��o�D �CS�yJ��ԏ7ԛ���*D�x@�GX0�0=!Ṙy^�YB )Ȯs�~��fkUM?�6��:�q��/2Yl�S�t��-6Q|��Ŭ�-3hA�Uaʻ���#����U�"O,I�C��;3��0�C��?�vH`dɂ�y�@ ?�@ȓ��09�N��]�zi���.I,�"+�L2tE4w�ԁc�?%�����RxX�$�/&8�C��. ��]p6��<kb�I,n; �s��0Ks����Y'v��	I�P�5��/�����$˪o��D|��!J9��Z��<�e���yB�P7�Sg��*}ܼ��n��;t��qKP5l��c��[��0�bK��&cRز�Ks3���SFi��j6.�m[��33+�}�bC#��2FқVR�]@���S�F�X.�������D�;&z�#DlK�~�r�3L�f�$�a�D�O�!��v}r�b3n�,Mf�ݿ�FD��lϦJܘ��WEF��^����#5��<�2ʐ�,n�¶���)?��#�V^��ɞN��@4�xT0 .��?��i�/��/�왳ᒽ.���jSl�:FȢMDy�$�$ob�훷邝n��hWd�H��	/8ՐM�V�� �RrVgʢ��W�,�X�U#� '����$͇e.�B�M�<T����j�Uk�}Zr��
_�A��\,1.6�R��'R�4{�E��Q7j8�c�ƄM�"O���ʍ5/8p��#[�>�nl�@��q*�x�-��,M��������%��!}	>4q�䝄n�Pт�x�t�̐�V��ȐG�06d ����9%v��%�O������/�̈́�#�4l��(�G�%�ݩ<���R��߂E���i�A�
��(;D���PH����E$h��h3?1F�?|B-��$��G��h*A��c�A��/Ăk�{�'����<!�Kα)��-��e�3N��S2>��V�͒zڦ9�3�ԉ� 1���be"l��-Cr�0CTC!��Ɠ2Tx�	uC�_�����m*�}��FG`	pg�U|����+� �ص�lS;m�h!1����������4��MB,�S�&�jr�K@i�:%�a� Kѧ�"�ؑDvP�W��M2|E&���O!jpD�\m l2$��(*(�`�j�)�d� �F�t����"1O��&��N 88P0g�,X� ���.������jT�����M"Q\Ua���-����B�Z�X�%��E5z��G{�f��hn���7������V����+[T!�dM�>���e�m�����}�ў�ANC�O碅�aN�[���ah���s2! �7R��G�~���7�1LO΁!��Bqd���`��I��e��`�e5�5�2�G�VPL����'���RR+M�h|j��N��d���$0>,���&W�^�D��1O^�@�>R?b QT�ӂ|1�lp��$#|�8��d)"x��)h�˅)-[�0�c��:�p?�ҫg�l�+&�&}1��B�3a_(�x��Ɯ�i���p�'B����4��`b�M')�F���="1��s�"O�M�IԵh�6i�1��.�n����ɿ0S�iq%���d�#e�[�[�&��()������Dw��LjE�H�U���$��&��t��
$�DH���D�,�f��IH��͂���?>�f�{��	�f�;����T��O<ɉ6�[F� ��%�Jʘ��s��W%L���bA_�uF@�0��=m1��򢌻"k
+#�Z`˦��6hXJ�z��k2��06�'P��R��I�5�4Y UԠp�M	w��7G�5 ���SA�?E��w�
�QW�&� �`�3H�}j�'��%���J�ך|�V��Y=�?!���u�p���eU���$��e�'Y(�[�Ƌ��r���� ;�L��(��$�lۍl�άb�#]�l1�$rL��>��X�f$�6�Ҕ�Y`G������r�Ї+V1��I�G������4i���P�G�~���@)�O�IN���!BV㍡1�p�ե��>!�բ�f��&+�i��I�F$Z,h�dF�+2����T�២|λ�/ 2n8�Bf+ޝw݈�������˱.��s��]Ք|�e!�.���d�gA��QE�wb���ƄX���j'�S2������7�!��j���;M#p7D��ϋ�'�!��O�X�aJ'�	�z,欨V�E+/!�� �P��|��u�@��h���"O +t��3H�E� �
]#"O(P� �WkZ�2��0�l���"O�e86��$�ST���|M��1 "O��I]�*5<!���x2A[�"O~���h����,*�&I�ލ��)D�8��S�Y�&]:�	�^���T�&D�aCC�&<��aNۡP��%�5E%D�`���W���b�V#"{޽�D�"D��Kd�K=�6�Y�j�m}r��d+D����BD;Bo��J��<w">�K��*D�HPskӾ9�=���φ _"EE#D�\!��2GA��2�BK~��#5�3D�x$Z�R��R��L�U���4D����"M�zr�<��ȋF���d�,D�l��Έ1_�ӕ�ɉJ!��ӂ�=D�L�o�*:��ˣ �.њ�C�(D���g	��Z}�,��.��%(D��Ð���ε�$!�(4��]�*OEOC-[�|Sf_�<5@�"OF�F�9J�6mr����t�"O.y�!�H�`��JT����x u"O�Th�F�1��� �BׅW�F��"OH����u�ʈ��*��%�<1v"Ofp⫉)�6��3O�$Ȋ���"O���!�Oܜ�H
7h���#"O
=�1�1tI�غpgw��xS�'D���pɉ�`?d����+F���`�B D��B�˾ ���ɸiC�Ҷm0D��B�I�6J��ZP��D鰨���.D� x7�5@옔���P�z�+D���Ӯ�gm@)Z�(�*�n0��'D���cK�-;-x��U.�Sml���	1D�e� %�B*��D"53����0D�Dc�X,�гS
Ɵ6�����8D�ܛV6y���p �!J,�8� *6D�,���T-]��3�!Q�/�D��Ն2D��r�* � (p����4z��<D����,B[��UB�I�� �ѭ'D�(�e��L��{DC	���3 �%D���׃C0f�t��f&�d&t0���#D�88���8][N��C��e
��ai,D��[��Ьy$���!k���2d8D�����
5"��X�DT�V��:��2D�px���6b� �rS�n ���0D�Dh� ��*�Q@L�}��o0D�4�V���J�kӏ�r�\}���:D��ر���u�xB��3^�2�7D�h��`��!���M�<�$��%5D�4�*�0�As�)�8a���3D�� ��
�/�Dm�dn�`�ّ�J&D�`qv�9�9"�A�7�I�W!0D�8qAd���}�hU	x�}��,D���',�#�l���@�{����)D�8#�/%�r���D_�ay&1s!�<D��B��E*l�� HcB©F��Kc<D�tq�-�0,VY�6��P�h�S�=D���"i�q*6]�2�%�~���<D��DM��S�`'�аk�F���'.D���%����JŁA�YB.��ю7D�\um\�'�N�J�����5D��{���)�nĚ֣�k��RV�&D�|k�� >���ťO��(�Q6!&D�D�3� �t �kN$������1D�� �����ޯ�Nx�P�^�Hj��"O(q���8z�rz��ܛ!N���"Or0!�*�/,��HԌ�^�v���"O��	+j�@rPP
r�&)��"O�I����g>P��91xlXC"OꀍN[~Z�JT C���u��"O^���í0�h�Q�^�fN���!"Oh���O�4_K�l˜e��'"O��XE�D t,�%�C-��r�"O@ ���Z�t� n�=`oF�[3"O�
����Iܚ�,KV�
�z�"O�� A��4�u�*q$�y�"O�q�D�<r�Zu�FT~DYw"O2bc`B<v�X$;�IcȌ��"O�!���M/#Y�xi�f�5�Ȅ��"O���3���S��4�P&S�p����t"O�hإ��U�F�6�
�{Y"X`�"O(�pH3,�R@ZD��A�xű�"Ot}j�k���l�V�<rz�4f"Or�����z�-k�B����P�$"O %�Z��(р+�5Y�Ĥ��M\�y��_���|��O	�O��`ϐ�y�FT4O�����V�}Nj�c�����y"�� 2~q��jF�rN�B����yrm�`��%�D� ��m��M�
�y���5N������z4akSO���y��?N\|��IM�
�EXSbџ�y�BфM�v�*�����9����y����ig��O���r"+�y2�Y1s���KQ���M���y�m�;K��,�ⅣD�S:/��1+�'tq����!7ݬ�{F�!P�,�'=�̡�*:x����^!����'�t�ç3;W��$�"PF��'l��pQ�$Qw�Q�f��K��i��'�(a�$��B2)v�ԯC[�h��'+x{7��F�4�+�a��&��Y��'&6XC�gɄ�Rt�P4$mHMA�'�y[�)oe�8�Z1���@�'b����J�Z<�]A�����R���'E��K^��4ev�ӯH����'I� ��"� �E����
���'Ǝ]�Wd��*[���Wx4Mi�'��H�cnB*i��Qcʀ^����
�'-&$�BJ�/ �Ԁ,�Hc��
�'�r�#2�R�d�@X�A�<?�}�	�'���RiÈ�Ԭ1�:��:�'�Rp"
 >g�*Ax%�4����
�'�L+�)X3>v��*� Z<.��U3
�'����T��;����3��z�>x�'^�I֡]�w�ҭ�RKֺ^�����'-�e���S&l|>=eD�*p���'zҵ����%^\�a@W8'T 8	�'��U[�-�*��b4���N!q�'� ��&�L)/`$@�#B˦e/���'p8eiƀ��?t�m
�fCW�v�	�':�P�@�G�
�'i� x�� H	�'0|d�� �=�.���������'���;폣x���Rį\��`���' ��#6G�;0j
��C�BҒ9��'ް�P0�̲!A���"	����
�'�Z`��&I(4&]@@	V��	�'�ĩ�B��e��Y��%.N͚�'E\�u
�F��� A�< ���� l�k�CA�<�c5ό���)�"O,Q:!�͜~fn����_0j��Z�"O"�H1,$e�#�Λ]�T�r0"O )C�B�)��))�L�_����"OP}��\$Qd���-υoth��'z��HV*�Z�ț9,��tQ���Pu�C�I<Y��|;�n�1A��ɺ�
)��C�	3|:`��'χ�H�So��C�ɒ�p��@I'a�`��Cµ:��C�ɡ7/���@N&rMP�8F�ñ	R�B�I����l� �Ϣ�X��'�<,�V$�,%�*E  b'#7Ni�
�'��4���/.�@x����) ]J>a�4,�HѫP0<�k6'V%�,���v�i��
c�ݺ��`��M��KLbp��3`'�L�UhK�����������'E�u�`ڱzpL���
�,0I�N��lJ�5@�dQ,�J��'�i!�׈>F^������]�ȓX� i�UM��b9�@��D��K,�����a���K?��b�f�&hR��ȓ �NHkrS	v��,` �λI�NB�	�sPD���W�T�5(��7#t,B�Ʌ*R)��i�%u,��� ��B�	�&��R%ŗ .8̨�M0�B��x�2�k�C�30iޱ��' �c��B�I6S�2�z6I��eqdU�n�=*�B�I�1��|+P)�	,S~d��JT��B�I�4�*	����<rQD@�Ǌ����d�`P�-:D�fY8� �ML��sJ7D���riF�;��AI`�.���J�n5D�@#&) �ԝ����X��@���3D��3��T;N��BDՙ�&p��3D�Ly�K4C�a����"1D���A���X�;�4h��٠�#D���Rd�t�0T�W�l���'>D���0%ܖ>X�
�	\�Nu��E<D�t b��P�^,K���5d��8D��sP��J�q�I�f�8 Z�(�y҃�:��c�M��8F���y���Yfc�o,{@n	�y��w�<�e)O�mo^�����y��I�P��s���]� �A)ݻ�y2�88l��O/&���)4 D���'y�z���qa`E�5��id����?ѐy�E�xYVT*�1E��|Bp+6D���D�>)8��pS&X�=��<*d"6D� r�N]�7��Q��J&���&4D����U�)��j�!E�%լ`q�(1D�l��`ՖF��J�E	a݄�E+D�L�R-�#<R�L�B�Į ]��Sbc=D�j���<*�r�xb�h9���W�9D�0IW���(�04Z0�B�Uc|X�2D�`���Y|� r�F�	C�!�$	1D��&��-��4J�Ćq��cm.D��`��ի)��<���)^��U�H,D�@�E������K/f���(k%D�<J�n؉)!D��Cb[;i����b�!D��c#!<bo�Y3���N��At�?D�l��R�<��=I�GF2"zy��'D�$8׫��A?0͊�i�	l�@�Ǭ$D��B�(=A�wB@����	5D��*�Q�y6�K�K�ĘP)-D���E
*rH�a���O -�H��@%D�� LzE�N;(�T�3投o��͢�"O�s� � (�Z��ɫm�$Y��"O�%Z�G��$���2�	8q�R9��"O8�� π�2��E�1et��"O"q���1�:iɢC_��� �"OB�i�Jزs�p�uț>HR��"Oְ��Ɋ8[>�Ӥ�7s�^iS�"O���Fi=J��X#��Y���(�"O�h`#��6V<a��rV���"O��s��]�M4.X+�@�G�E�c"O���F��RA*1���W�!��"OT��1ϒ 6�zUa# �u�"O�y�4�0	 ������k���W"O2����$le� �7�D��PT"OPJ$�P((�paal�;I�xT��"O��a���ZC�#�$�)S���I "O�1�*>7�jU�2��)Cy�@�B"O�3Eݳ^�~I����!�X��"O`��ڻOZ�X��HV�o����"O�p�"��Vhy#'�A�O�d���"O�A¦��F�X�zB�Ŀ�|�c"O$�8�`ڲ`Zv@s�Q�YR*Hu"Oh-��{lx�3�ͨq"~\BB"O\h�JH�wA�p	�e��c����""O� eo��M�X�r�Ԃ>P�"O�|����j�땉�P(z�"O�E��=��`K&Ґ��"OB� V��g5R!�匓dZ�ĳ"OP�j�B�0�2\�cڅS�%��"Oܸ�s���|y�C�RJ<�"O��s�1�j'X66�`�1D�Ԃ�(-[RtD�W�p&��U�9D� �ؑ2�cG�5#F�Q�g";D�t;��
yf͹�`�+l>�Ѫg�6D�`Q!���e)��K�C�U ��9�K4D�L9QO�v�44�tC�,mV�	Ơ$D��Ip��
����#V��h��v=D��1��%���a�^f�+t	:D��Kq�W�#a��Հ��>慒e%7D��`�ԯJ6��P��d���F�4D��PĤ��6|$ZM[�I�Y��'D��q���&lo~��:a\(���)D����NޏV���@�	��Vر�4D��c!Ս}x�+�D�~)�.D��2PK��]��(�c��O�ލ-D�9��O�hv���v��]X�3P�&D�4�5\<A�p�{�J��G��p�P1D��ZF�ǬRp�e���*6�zUK/D��ba�U(	��m�Wj�!R<�q�K-D������0{����`%�3w��1�5�-D�5��e!x\�����ax��-D�h�3�H)�0�v�Æ`�"V*,D��(Q���V9�  D>L&=Q�c&D���U�àeP	i����,�D[0F#D��"�j)^�$�@��.<}f��, D��YU�٣0�ʅ��̓N(�2�>D��hr�Q�Q�DI�@"0Rn����:D��Y@�B'�s�09	��8D��A� ������3_1F�Vu:�(3D�0sE�P�V �	"&Ș���I�D2D��Q@K�<e���C;[w�};P�0D�DK��)4����L�s�*)�b0D�ذV��/nȽ��Q�T�"ъ(+D��çb���G�P#T��U�C�&D�� �P�c����G� �:أ�"OJ��މm��d���]v�Hi��"OV�E�	J`�h��ON�{�����"Op�� �D)���sS�Ԑ(�&Ļ�"Oh��%V?E��P;de�Q��C"Oृ�H \��P�q&5�:�ʓ"O$����/VM�D��c��h�S"O6iC&$T�NID�i0�ԏQ��X�	�'���b�]�J�Qb��W�_��
�'9��A�gO;:8��ދ��Y�'����c��+�m�b"��~�$Z�'���Mԋq���' L���
�'��h&E8��M�'J; �K
�'P��G�_�c��-�fJ��`@�L����=�J�.4DI��^ ��Ʌ�F����3s�B�ؗ�X[��8��'�lt2�!B�Sb��L} ���96�0c&ҧuP��!��QmK"D�,`��)w��F�H��(L8D�\�3�E�>8b���@ߐ"�Hڗ!!D�D@�Ǆ�B�X����V���d�)D��⦢�m�J�8P��Q�%�&�$D��Y�eA$f��t� �M�kO����4D��
!�ɵr��)	���,�b�)�-D�T����l��5cް!N��2�(D�$1#��-e>µ`'�F� D�g3D����h��Z�P�tŐ�kz�� &*0D���gωe>*�BCȍ�Qa�e�� D��@(W�C��L��+9v �q���>D�\�B�0v��d���D�P`Z�0D�xp�F�*T�8Qą֔>�e�-D�\�6C��C1����,I�� ��&d8D�lp����M��5��L�c��XY0A3D�����n�d��e�ʪhR����E;D� 0�`
���1	jܥ�X\i%�3D��Q���3a/ �h��]�B@aK<D�����A6�����Y8 CD�j��;D���d��`.����Y4
�b��6D���AНa0��IE�	(l-J�фf)D�x����h�@$ ң�	s�R =D�@YF��3\* �[�hE=Bb��b&�;D�<B�JV�,����n�H�d��I&D����8!��8"T�*����"D�x"�֑Mֆ�{�L����.D��'(f�P��B�&b`��,D���H��
P#jN_�v8�)D�<&��_�����	S�A��(#D� Ʉ#r���0��L�t:PX�&/D�����?�$Ջbˈ\���j2D��9�o	�_�Z(�^��� �N/D�l�@O�$Lz�XզݠMn����.D��ԁ�*<�])cb�1x�x��S�+D��h+�v���0�^;>���f7D������BÚ�Ca�]�<:��:á3D�4
�LH�G��8���-���ڡ�/D�\@�狴&��}[EA��8
� � �.D�� !�=(���{�C�$h
d@`�j)D������Pm�I��F�n���c�%D�(P�FQ�K@b�TA����Qc�#D�@�j���Ͱ�e�|���x�>D��bC�Ǔ@��I��I+��ؠ��;D�4�!dFɣ�G	._��49n:D�$����,���7fF?3+�(UL-D� �O# ����dQ�<b!�� ,|����c�"�� �[�<![�"O�<�b%��/ĆY�Ь��P�Q"O��	�'���� Ǧ��|���"O>��Aq �P�O��J�z�"O�X��>�uH5� |����"OU�`�Q���Q� ŤaeX���"OV� ���>�Js�ƁU]m�s"O�����4u�l�RwNK�qK�9�"O:���A�5S�����OJ�ɗ"O���Wk��7�b��UM�=|��"O&���@!N?
�"��R�)��K�"O�0�\�Uz`��@*/p���"O�I�5���-Xz=yP+03���#"Ox4�ǯӂhz�#����*̨�*OT�Q�@�B|y��K�����'﮹WN΂(\�m���O)AP��S�'&谱�M�z�z͢��J5�H8s�'�t ��*ً5+a�f �c�!!D��9!���W@JQ�š����;�O=D� kse�B��*���aF�qr3!D�r�\��4m�s�ط]8ty3�,D��3H�)Q��8�,ՠۜ]�H+D�D�A��*|�2'd,�@��B@)D��;�i�M�MI!(�D�x�"D��[F��T��Q�ԯ�Vu�m���+D�xk� ��	<ɓ$*��9����,*D�x"���&13��x�e^�r�l�s�*D����V!�d��6[	˔tK�D&D���R�f�P�$:/����o"D��RBo�,0^DArO�z�����;D����$'^��˕�>�x{��'|Oc���k^<t�i��b�k�tp)g
2D�����W
�~�S��(#�Z8p�5D����̍3ƆPbt�I���
��>D�����i��j�W�ve�v��<�.O����,V�I��͇g �:U"$!�������l�le`dX�kN;k!�d5l�¡d$��kDd���N�!��.W\K�"Ó*Bv�g�%oў��ቄtƪ��o�L�|��4���C��	t�rB���<� �HC"W�f�C�:`�H�7��j����k�P �C�I�FLn��UDKb��ly#ʉ�O�pC�	lNhpq��O:���*�AFS@lC�	r��*��u�D|��C#[�B䉆Q�t)y!���s�@�J����DB��q}���lȽ[�Pt����9�b��D/?�&h3*���0�	c�ȁ@��^H�<�I ���fɟ�����,A�IQ���OuTT�a`�6Px�� BQvCR���'f��:ՠ^�M/�8`H&pZ���'oHy�V�҄[�����a���'5�cW�T,���ǋV�����'ּC��V;� ��J��9l��h��?��yҮ�sk<B���:��@3
��yBb� أ�,�u�4]�S`��'gaz�!��(&�]z6.Ui��`�u	��y�-Ӌ!�v]�4� e�BL{���yDF0�X\HǇ2����(0�y��ޟ=��T�ń�/C~�s�Q!�yB�.4�DcjҎX�}���ޅ�hO��O��O���7�G�w�Ҽ��*_�W
���8D���H�"���

@��SRJ!D����ʈ�xTz���)�-�p;_�y
� 6Q&"�$6���f�QxI���"O����$UN���7*E ]ո�"O"���k�E�08{7G�.2K��'5�'�az��I;9q.%�"��+�BIX�LM�?��R�s��y��F�|p#F �U�X���HG�<idD��d��&�Y��A��I]k�<	�LO5|�H:��A�t�Q��K�e�<2��2+�pK�4#�]
��_�<�p�J/1x���Eѹ
*�`��DUu�<�vO�:�CB!�Q�6 ��Z�!�D^&M��lЎ���%�S��Z���=O6rCJ���8u	��M��5�"O$��!�)
�(ܒ4�\����r�"O�1CE�5�n|���:.8��"O�� ��	a�q��Ę�SB -�"O<�	U��.Yq��#�c�>F�flQ�"On9�c�ܱ7g��p�$'.�S�d�Ot��͎h�,ɹ�(�m�b����=~���U��\5�%��ɛ��J	�����1�^���c��B�,�@�D�}
�B�Iz��
��]�H�)�0ԗQT�C�I86hp�J�&K�e��(���C�IG�4c��"i!�� 1͑%~�,B�-��9�GlJ.c8��@���0�O����O��𤟬S�re�n�>~�Y@��<�!���]n�eȂ�Z� ��xR�~�!�$
�NӒL=&3z\@�%��G!�ül ���I7H풥��H/!���]b�DY�`C�R�x@�L��l%!�dϒ~�	j�*�>1���1����!���lt�Xv��5h��ĂG��IꟐ��c��S�e��b�*�F+],�ѣ�.=D�x#EȣY#V��`�+3���"gi<D�4Y��\�J�b����
5Pj^���O����S��{r&�W�xq)U�JXR��ۤ�y��:"*��0�+�A����W!�y��2}vIkCC�'5ٶ�y',���y�A^$-hV|r��8*ƌ(�fƔ*��-�O�$"qL�A �a�+d����"O:�� /�vʖ�a�\�)�ȴs��|��'6D��$ڋ	���Ӂ�޷ ax��'��p�7��VO��p� �E����ʓI��ȳqJT%u��T��C�"'`�Ն�>�q�r�$�������z��
/�dұ��1��q)v=dx��v�p�ME6M1�=�d��?�䄅ȓ�
%ab�L�b��:��O ��)��dl�Q��,T" �H�����ȓlҤe2�K�qP��Yul<`L�������Y���&��C�4����"C����*�u����4(�ȓh�P�Ԧ�y��MP�Z2���	O��ea�8)fdH�Mډ3/�����8�5�ђ;36��@+7����l{�bʣ7q��+GJ�'M��i�� �L��"p���ۓn=%�@���GȨ0򪁀L���{E��0"؞���_�E����s:*(�5.	,a�m��Io̓����࣐�[��dS�"�*g��E�?�ӓI��!�d�L��ʨs"N�;DB�ȓM��)�ԃ�?1��x������	\�m�,9u�ä()>z��P_�8��ȓ��Lf�O�N7@<�(K>�Q�ȓ{|:|j��D���)��.F���S�? ) �N�%\:�j�K�8MN(�V"O��  F���D�����>4�����'��d����I��C
m����g�;7!��rj��cȝ�l�> �'�30!�$��]�Z����ڜy��x&J��%L!��<w6$E�w35�|���"1�!�䞾l�p�1U�r�e�� �SV!��!�&��� ytp�1�Ј!�D�_0���� A�O�f9`�]*"��6O�!c���4i��h���\�����"O�������m��y
��$J��!c"O�c��)mx,@+%ڦ։�'"O�PR��Ih�(����-y.�"`"O��j��W4z�VX�D��.2���"O�)t��.�`Pig�ѪB�"OΡ�w���l����NƦ�q�'���6a��=�׬G�����k[�7�ў��ɓqĮ�6�Y8�\uaԮ3��B�71���xF/µd���QҮTel�B��:��|q�,֤B��ku-H�d�C䉄&~܀�1LV�,��=s��I�C��4(��y��5u��E��	�,}�B�	�ro�8[j� 'n�<"D��;�˓��<��O��p�jJ�]X~�r&u�@�"O��j��H+/�r=�D�_�&p�"O>���F�9+v �i�Ɲt�^T�E�'U!�U�+ttiH� �L�"��!���KFZl{�kLu6ȉ��,�+t!��Կ%��x�&�5Q��ܻ2쒳a	!��5F��a�˫zJ�����}��'2��~~���g��@#��*��#���y��ǧW�^��1���̴@8���yB�������b>x8���l�8�yrDѪc���d�ن9���)&���yR�G�U���W�#-v(H��G�;�y� l��đ�Q7#��A�d�B�yRd�	[�P�[���.�)�d��(�y�Q�2b�JB�ѯ9P�M��y��r�$�#���X�UC�BY�y��)e�n)h�ەg���&��y�Q;F����Ə�8Sȁ<�yr��`+��"S-L�|��\2S��yBBɾiJx�5�F4f@���2�§�y�E�e$�oK=P�F�s2�M$��.�O�l�u�P��2��T�44.�K1"O`���&V7�8�&���L����"O��0��ɾw�>PaS�Z�8^H�T"O
B��n��q�V-W�W*J�"O�ZF�ϧW|�����LV
`�`"O�T1�M�]J`�j��6��ђ�'�1Of�K#aAlyV88B��s�z��t�' �	M�hy%(�-W��͐r��O�<��h-D��A���+Q��]�poً~�"=Avo&D�x���
!K����U�¦Y�D�e�"D��C# �;�flPrg LI����'!D�$�lּk�2�qa,^�%Q�u`o=D�P�3!�:��(���]2a�ΩZ�a=D�$(%��y��%[!�H�@k;D��r�AΜ~�5 NسEW��2GJ;D�胂��CMva�����m%|�rg7D�,�Ӡ�!QRܡ���B�\�Y�rC�I�<�"lᑄ�8t���S�H�M�JC��,e�H�1�F�"	�0x�&D�%B9C䉵r�P̢���6-��m�TĦ;�B�)� ��fd�he�艵�\�Avp-r�"Ox%�f��Cd"���L�-� L�F"O���ïҩe�`r���4�N��p"O�10�I��2���}l�أ!"O�Ѣ�K��@~���BO�+Z
�`�"O�� ��;|�Եyb�:e0:��"Omy��C!`�P��CPJ���"O�y9��%�z0�b`J'��l�B"O��s�Öc\<8��Y��9��"OD��w�D�=,P��V�;-��Ac�"O@����ˆ�x1.��O{��"Oڼ��dJ�d����m	�pzyA�"O�X�%� 5��0�*}�G/xY�ȓO��Y���0�L�ɤ��nI�i��	��IR~�Fj����$K&4�6�[�S�y�1h��Ԑ�,G8�����y�lҜ$a~���x�|�@=�y�cIH���(�%��t�l]S �9�y�ː
Q����S�@�8�����y��]�^~>psTk��38ш�aO4�y�Ҏ�0��J�*$�X��5�9��=����D��rc<����/3�)p��'Pp!�d��бD�=T��6��^V!�����z����{�& � 	p8!�D�]�X5	�d�������7�!�Z�Y�����Q&�H����9X!�d1_0!�P���WA����HMU!�bF���(��4�t�tGŉ6\!��Q�ȉW���ۆF�"O@���C$Ѽ��N�g��iˢ�� R'��D>�	ϟ@F|BB[����`	�0}�^�)&3�y�S�%����y��lZBg��y��R�Yq���:X.-���%�yR�S�G���rFI&|D��� �y�Z���F��VTM��g���y⬆�,�� o�+���P�I��y�i\�j 4��Q�U����?)�r�'��y©G����dҷX�Q��<D�l�c�� }�2������r���3��<D����a��.��T��0aV�D0�:D�l�!�DoP=�Ex؈� �7D�h�H�^��e�!1�����(�O�=E�$+].M|�b&��r򼼐�n��%�������4� }�����I�@w���d�-D�4˴�"���;C�F�IXmP�,D���s������oF6i��1���'D�4�����v�R�b�-h��YcH1D��B��Q9v�
��!��
`#�m[��,D��a��moh�-�s�u9���O^�=E��n��D���"�;��-0E�'�a|2���#��]�	.������y���!Ar%�2mI�yfN ����y��/ pi�S�Rs�6��� ć�y�&��T�&�Pa�؀pJ�L��%V.�y�`���=bA��Z��� F���y�ic�|�rd�>f�.� ϝ0�y҄@/�� `v	�B����
���0>�6�[�Y�~E�C`K�4��=�$��o�<aD-]�X���(y4�b�ǐh�<���W"}�r@��D6�,�K�a�<qa�٘ptD����ɇ ����T�<	��{����Gˎ?���2+Wg�<q�nO�[b�H�*���d�#����F{ʟ�b��S���Ls,d�� y��!%?D�� ���3�E��"�9�`� ��RT"O� ���۬VP��B���R��A�"O��kb̀7/9�ܐ��VR�TxJ�"OT�`���#Z�ژ;��ۮ����"O�����R*�T���`��[k�p��"O������.�*0�ѯQ��@Q�Ic�Iܟ@�O�Lrt-K$:I@��Zgʶ�;�'9FI;�bL�NT�
���W*8�ҍ��=O�x�-^�6T$!��
̈+uT9B�"O��H�ԉnR~u{o]�B���"OV}�ª'8FD���(�2�xT3�"OF��uP�
�݋E�T�>��l�B"OD���"C��a4ɇ�-P,00��D�O ��)��7U 2$+��u��2��9!���Wd� p5o־tX���9^$!��f��,��n�|M,���N;S!�dO i
�- ��%LR-�fC�+!�dd���㘸(]|9c !�D�2���gf��Vw�A@ >Lh!�D_g��Q��{c�0�aǓ��O�=��
,Y�J�C�P`4Yp0l)�"O�$Bf!D�Yb���S��5mI��"O��p4�N�z	ČI4E�AO"u��"O|�U�N!������e@TI��"O���F�P�$�c@ɓK�,�ɂ"OX)0�D*fg,��^��!�"�!�S�~�z�Cq���<�6Y��N֩lS!�D\ D=�p����j�dD���/45�}��'=�C�:602�X1(X)krN��|%��j��<�2.���؆�f� ,�d�$D�$Kw�%���T	/V��� �!0D��Wh@4m;������d�v��/D���'�Μn�����>0yl�R�,D��Be�]7`��yb��W�33lѤ6D��qBկ:�`���F�T�2�OT�d�OB��g
.8��DC����G2x)J��O�B�ɔ A��`��:�<�ӌU�=� C�	AhhI���Z@�XA�_�X� C�Ɉ~+V���DI��(�����B�	%a� 3��̀'M�;����B䉬�&��	D��0���({�TC�	#���"�L3&�8�G 2<���O&�-��\���@�,F��`N,�������>��'L����n�w'��;�k\;Hn���'^n	�w��"m����⎎ED�l��'bн�w�kN|԰p���A4>\K�'K̽�rc^�!�Z	�gl��:�l��'� , !�
���\B��H]oȅ�'T^�z���@]���P��x���?ɞ'�P�KB�E}���s���W�t�����ϓq��DX��D�&ڈd�գ��RQ�ȓh�8V�0M�PD�B��LLI�G"O~��%R�$$�,K�ƅ <���"O��
��6X%P����/ �1�b"O�����y�01s�B��N#��'��ɦcO�k4��B ��P
�ds�M:��M��� �L>w疱P@��{y���Ā84�tPB���\͢A$*6�ҷEBq�<��0�6uJ@̀e�ldr&��j�<1���*��%�a&� ��x�%�k�<���U�y
%�a�֔\�����`�<��JM�m	r�kS�*a����T�<Ia�+��Xr�;O��H�i�Py�U�����RM�FL=P�����33<�O��=�}� V0C��^�+�t��lȁ2P!1"O٪�Lݲ,f(X�L�8�b"O��j� �Dw:9��$]��x�@�"O
�0�?����#����#"Oz���Ȩ�
dc��hN�4"O&��UG��چR�'ߊy�pyi�|"�'MJ�PQ���o��Y��j��x	�'B
d����[C��6d��!"Ol(`Q�L	"��	�UB�`#P�""On��g,1z��ª� � u"O
)�N�����1C҂ :<(a"OD]9f�Y5w����S,(��a"O<�`�(C.+\R4���t!�j�"O=Q��� V;�H����IAp�@U"O��1hXQqPtɲ �5nͰ��C"O��9���F��@A%�"�҈��"O������/�@�D��H'��[D"OLM�Sn]4����b� �Er�"O��8���$T�"�p�m��Q)�"O�Dkt;,i�'$(��"W�'��	�<�N���Y��e B瞷O��C�I�N�
E�]�:�j�c@��V��C�	,3qD���j3��T�Uk��<B�	"cx�8Kc��QFB����"+#B�	ql���'�&:�>E8�	Z�y%B��{O��!&k۷WVЕ����>cB�I�K����.QA�Uk7���Jyϓ�?��yJ�;1��ie�á%Td�#4�A��y2��K
���H*,�P1�H���yrɅx	��E � E2rA��y,�?_��mBe��aAh��y���/w�4ВԁV�M4`���O���yBIָ2�N�Ju&ŗC`r-��ڑ�yRlM��J�i��@���d!�&��>�O8uaq�L��r��F��N|J-��"O�����H�����9`X<�%"O���H�)�r�*`8("�-B�"O�9�W�Q-
(̱��G�KplA[�"O���G�&+rP�q+ R�p��"O������b8�6K�4C>�+""O�Ȼo��t���K�)�i?-��"OV WF93*�y���W"�*�@�"OМ���(r���[!OxJ��$"OHy�Ĝ"H����!.q���p"O�5xn�)yL\h�2m�3n���"O���㗢l��1�ҩ�TFt� "O!�!�N�L�X�'	UE�0�R"O2�k�B�I�DXWFW76�hH�'X�����8B -
ӏ^���ͺ�'���h"T'�zlc�i_�5.#�'Ő݋�c�7F��T�Q#͡3���'�(�풺;�ႁ�@3�va�'*XZP+�e3f���ͧ+6̚�'���v�֗G��h�M�8�<ؐ�'�\�֌ �r�b����4\�e)�'
�b�L֑a��*�˕-��)�'&�)ce�������C�('+��j	�'l0�Q��
�zJJi�4�^$�`-`	�'c���Ԍ�,HR��8qA�}q���'4D|@R�K]��ī��C�x���j�'����L��M�X�I�āC�<I��'�J�S%P�/{<�[uI9q����'��bn�.��a�M�2�4pR�':���敋yWDi��D�W�#��� � ������m�-\�9�A"O.Y�Ў�pqZ$Z���w� ]�"O2���ɏ�bk�E{�H�&�.ɘ"O���G$�m���aW��vخ�p�"O�z�M�cH>��(K+44@��"O�����G�Q� �1�Ҡ*y� ��"O8�Q���i�����t��"O��)��\�L+h�Z Z9!����"O�������t \�1#�ԝ4}��Z�"O~i	���@x�3Ų[
��"O�` �f�U��e�߼+�iW"OIz���-4[ �00�|M
5"O��R�@A0AOj1{'��rk�՛�"O���G��"���������8b"Ov! V�ɉj��magd#}<y��"O�l#\1
()GML-V@E��"O����"�Z��0�4�i�"O&�ٖL6�����M�4v�Q��"O�[!e�wD	(���	��|�S"O�rU��)�������4�b5�B"OhT�&��H�F)R�;���8u"O��5@FT���@���]_���"O��2�Ǖ7E�8���}3S"OLm�s!Ɩp����QHae`]�#"O�@Z�GQ�5���%�a�H���"O����M���(���K]�zT"OJi��I�V�4��	�.�(�QC"O�d��GB�C���@�:y�\�Q"O���`o�:qcl��n	IM�L�"OTEK��'r|��x�,Wt]C�"O�y�AIT�}�Ҋў��� t"O���4j�{M�=�	�E�u�v"O���pǒ=��%�TǕ;S'ּS"O�l�1j��x���VeF
ڭ+F"O@��c,N7>��0����S�$���"O��1,M�p�I�B�ڹ�Ƙ��"O�Y�Fn�9j�lH��2�~���"O��Xf*�"$�J$xR��	I����u���1+ٟ1�J�C��܇;�¬G��'Y>�S2G�;g�"@\�|PY{�e!ړ�0|�A��X�09J@ X�A���Z��~�<�,��_.�(Dl�;)&PʂDX}�<	�ߖai&��@�?#�lqPfͅy�<Q��
�N��y�L�:W�0(A�Tt�<iU(ͥ\J�A_9��Y+'�r�<�.�02�z� �)ʊMJMc�^Wx� Dx��B��)��cިA�|8�RI(�yr�M��L�At�K�;C�0�a%���y��[��4��ֆY�8��T1��ˡ�y�ԿAǒ]Af�=+�������y�"�bj$�W	ˁ.Nb��6�y��Pk��q�VS��8���y�;9�༛#��7ER�`�G\���O��$*§J��
.Ϝp��+��U�?��I<�i�����Dl���JgG�ȓ ��R��4K���Ǽ �t���t!2�JR���~�%ꏐsS�,�ȓ[��)�A�$1�\��N��qq�ԅȓ$Z08@v)QE�
n����ȓI�Pp8�Ő�#��)��&Ȕ�E{��O]�eϺJ��P�T�C&�@{*O���B�2�\�O��,r���`惕Ei!��r��'�Z�&-�#��L!�=c�LS�	�3�\�'�Lk`!�� *d�g�R�86ڹa��M�9)|)�"OH B��J%D��9��c�(l�r�"O��C��L1s�
i�����R<Q"O��G%�z�í>$y�"Ov�y3@Ř,&xxq�I�f��(�5"OF���ݑC�TI�c�)��	�P"Ov�zR��=t�h�F�3L�T��c"ON�c�B�g�漉�c� p�J0��"OT-PI_T"����I�T�M�A"O�E�OK�U�&e�v�0oʅ["O��ȵ��C�Hpv'ɮ~�>Y�R"O��	�A�o� �� ���p@�G"OD�hPA�>��fQQL��E"O8y��ôs
��[�#�	(�61J`"Oh�pf��/�tx�R��>��ժ�"O�,:�	��NЪ��Q�^mz��E"O��
�  �<C�����M�2F$�"O���C�^+`W��D�w뎴)�"OniR�S�������85�`�"O�\@�"<�e0�"���N��"O:�!�$LL!&!W5���hB"O� �*h�X��
E��IRr"O�����D1|�H�/��|����"O��;Q��xj��B� S�"OX]kg���Q��;V����"O�`��G�t�(r��	\�d�k�"O��F	rip�h
[<���"O�|Iq�
�$>��[0nM�^���"O�ؒ��K�I4lM���΍��!"O^�c�Mqm",���G�\��\�S"O*`! ��:G�+㌇�`�a�5"O"��R�� �AE⍸-	~�aV"Or�f�[)E��P�Q;,��(�"Oh���$J�rp�y� �F�l�Flp#"OJ�넃C�{Ͼ�8�ʐ1�&u�""O*�� D�	X�0�*�u���1"O�r��@:Go�ːjL�Nu�I�w"O<4���I 5#sf�ӡ2s��s�"O�Ŭ�=��1!)�*\(-�5"O��1ׅاN�b��0�B��!@"O��x�'�]�L8�Gx�Ti�"O&YG<N�Q��,yq���0"O(DY��2��I�D�]v ��	�'�>����N;7!LZk3�ٜ�y)�n�p�d聂�$@$+_�y��ͷ+fp�;�(Td�93�Q��y�Ö��4P��	�FBL�bh���y҈�8?�:�i���@NЙӆȎ*�y"�,%x���>�F4у)�yB�[@�{s�#l�m�s%��y��gx�MB�*1��P����yb��B|�yyQF�!�P,�E&�4�y��ٔcV$tzP��;~ɢ���y�oįK8Ų#�X��*V<�yBΘ�#��W
�@��BF�y2�Z:"ٸU��$2�,���G��yb�H=�Z�ccc�>����)4�|k��,.rf�Y����;>b}ˤm;D����V1p��e�ЁZ�_6$ R�8D�<;e��
���ue�+����,7D���v�m�R5���	����h3D�����V�^�"L��b�J��5��*%D��Ir��]qCj��?�ʥ��/D�l��	6�*�`��iL�r�j)D�� ���"�R�?�I�d��2 ���B�"Oʅ"� ����0cD�$ii\���"O8���A�aў5Ó�:�ᱲ"O�(0��.�ɆC��+L�1j2"O|�2�ʈ(y떅[���<s�N�R""O���ub�~H �������Y��"O�Lٓ#Z;z�)�3���B�(ʔ"O��'�Q�.(a����i͈1�E"O<%��a��!H�����K�bD�"O!ˢ탇~����4
:B���"OH��R��Q�&���xs"O��j��]&[v���M.x�N��f"O�	�r�?�b�	�,Ƒj�(��"O�؃Γ�T܌���Ꚋl�
�U"O(����F@���*��S�F��"O�HS�!�kH2);�H���� �2"O>D�l
�BP|��$.�z�Rp�v"O�"si��sPXA��lP�8�{�"O�)�	C�E����ާǤ=��"O0e���6g��gK��Q"On�;A�$k:n(Hƣ��%1l��"O�X���HC,�TZ0��3	5�)w"OF4c��"G.4 cM��z�xd"Ol���L�m�ꄠc�A33{��"O*�ڡ�ؘ	$\@92�J���Bs"O.$�JZ<7�\���k[7��bV"O0�( A3� �8a͏r��3"O8 �m�<Y�ݻ�@�%!�����"O���Ê� r�	��mX�rQV"O��򷃑<+Z:$��	uA�=�S"O�ᢡ�X�f(*sH�5)$��f"O��X�D�#;��Qe)�8���"O�AR3��F�u��-�>m��M��"O@ #!Q7ꠁP����w5>ҥ"Or�0sgU�Tڐ�S�)cTX}P6"O�%�����@L��ѐ�>y8��1�"O��s�!!�ԛ��G9DL2٨�"O֭��M,{��Ec�(?Jv��"Ox}�s�� !N�<����;E|��"O�ت"�ǰh�JA"�.Y'	A|�!R"O�� qeJLq���E;���"O���噓��!C/�Q0��c"O��Q�f�>j�ibGZ�`ߘɢc"O�E*�ĕH��3��ޠ.����"O�� �	Rt��a��*�&��a�"O��i�!	f�f ��,����"OZ�Q"Z�Sv
15�8'x�"�"OX8�H8L�N��㥆�3*��V"O��z�d[0&����Ą~��8"O�U*`�E��8X��E���`"OT�$IZ w�ε1���Pq!"O&0�u"��C[T�s��-C�v��P"O\��0�ͱ>��rC�<#Pn���"O>�����@u�1;�G��N�����"O��T�y��i⧨D�����"O���F�$5����UH �({�5��"O6�+5�i�"�k��G�[p;�"O��x/؛;�T�b���l���"O�r��F_�:D�S�O�Fh3"O�	Ɇ3쪍�SM\"8�>�"O����ĕ/�����)�	�ؼ�"OR�B�ʙ R��<	��G(/~r��@"O� aA$t�\�s��y$D�"O��3eS4 �yf�,q�%k�"O� 8kACE'3���X�@ :X���"OH�{��й`�~�p�ɖ"��}��"O���R W�q��/����p�"O�;��K����ܒHb�q��"Ot1W�%��X�Ώ/>\��i�"O��i�NR�@d���,g�L}�P"O�5�gM��!�)�o��V�~��G"OʩR3��EȨl��g�"Z`^� �"O�	�]RX	�ܝM����b]��yr�΢E7~�d��;V���1�P��yMǖ9��)�%|�����V��yB��8ym��%.t��$�y��[2d�Ȁ�μ$��a��?�y��%O�X�W�(e�x����y�D/o��@QJ&Np� R���yR��z�Bܻ��MJ=��)T���y�,W�a���@@���V�T'K��yR�"y
p�h� E�[�PtY"ٸ�yBL[�sP0�%O�8O��`�᠔�yA��ez���f��F�B�@�'�y��Q5V�J��*D����ތ�y2�H
kh���Wb:5|����#�yeT'rȉ����3R�1`���y�#ǡse�\B��Z�,Ϥ���B��y���5;@LtѲS�&y�јV�G��y2P�M(���H-g=�����PyR)7%���l�SE�� x�<�Â����$��<2����!XO�<Q�΍~����l�����b�Q�<yĦ�0qn�"7%�s�\��3F�O�<��!T�9W��іCX"�l�EE�a�<�a	�^�1�%�[RZT�h�'H[�<�A��'�N`2��U�TN(=��V�<aA��
�~q�$��##����mP�<9E�:wD�ks�_8x�B]���GP�<YE ]%
�F�����7z�JL��Kc�<��B	�.�btYR�D6r=��YF�b�<�TdE:Հ�`ԣ2 c|*���U�<!��U�Ip�R�A(�d
'@Jj�<�EB�L(B)J%k�`�`�l�<��� �MSt5�W�!Cg|����i�<1�\<Aؽ!	B5`{� �c��<q �ļq1!�		�Y�XK�a�u�<�o�/$Ej1���R�X�� KԎYW�<�	+GR�)�wM�Q�<�w�ݠ��y��C���b)�K�<�w��N�����������lNI�<�hLX����Գ7��QRD	�F�<!V��B�*y����/Z����kP@�<�p��%d}��	�t�\ �Vl@r�<���W�k�zPCGS�=K��aJb�<�r��-(�;������W�<����%1n`(�J�������V�<i◀]K
�*�k\�J3����^P�<1de S�I2��,rS��a�Yv�<9�W�W��X1�H�'b�=���y�<)�$�BBPǉ�n1���I�v�<QdJ�95P�sn��]�tI�h�<Ad��x�y2���=e��1���@c�<Y@�/p�z��%�F�tlĝB���F�<����>.�x�.�n0���U�<ᑦ�]���V�|�lk�G}�<q��#Kq,`:���u���T�LS�<�P��0��p�ЇCv�}�u@DO�<� �dy�B��i�>d�7ӠF�hIS"O���1�|��-2���"OJ]��`�	)�6 ��L�?X�TkF"OKѾ&Xma��2o傰�O��y��!R�I��`���A	�y�&�w����D͖g	�lń�y2��S��yK�J��0��F�y����t�֑��'!�eq�)�*�yB��,�b���0qh�=r�ȩ�yRe�$2!y%&�,m�����y��J%� S���8QX�����y�3if2��!W�*��i$N��ynViK��ban�)"Q��TG�"�y��
�!}�t� ���"��
�yR�7 �(��h��H<SH	>�y"J �ƨ��*�~�x���,�y�F[ ]��}�d��E��܋����yR�X=^H ��!ƚ89����2 5�yB�����%�aE�m(�	��y�cK��z����R��8�����y���<AN�*���K`R��siF�y"ϭn��P���'Js�i ��E�y��X�h�`k�����'��5�y"�ݝP$�Ŝ���*,�yr�	lMޅI��"/����J��y��NN��z���*tw\��`���y"��OvxX�*�s9�Х�;�y*�f���BE�zp~�"N���y�,_��Y�7��H�������y�b�4#~B���k�$U/|]c���y�e�v��[����S�8��QkL��y"�׃G��hEl��T�4-�e���y7?�p��� уL�8���	��y"�[��z`�S�>B���m�yg��KR�I;r�=%�ر������y��Sz2�@�%�"W: �d��y�͑!�rp�`�+�e��Ǔ7�yb�A�aF8�i#+ߘ'�Z�Q!W+�y���uCnh�rɥ!�x40 gJ�y�l���)9��
!� e��N̳�y�855x`���*����I��y��'k'�M�E� ���Dl�y���h�p�*�X��
E��iG��y.�&Q!vɅ�t�a���yB�Ea%raQ!S���Q�ҭ�yҡؖ&�b���3G�hp@�1�y�b:�� B��6NP\p�A�3�yBh�Y��5�r�|������y�ω(f�t����dX�p���H��yB+շO86h��DſUD�1�AP��y�^� �A`C�]N��X��D��y"%��)u0@��IU	:u�P�@��y�kމH=��f/��1���"H��yҮ�1<����R���-{��z���"�y�X<E�=!e 9�
��q�ת�y�X�w������dm�� ��B��Ts�IО �A(��C��B�	�]�����d�!G��)&w��B�I+$���P�3�c��6pB�ɔg�a"�D�#�l�� ��-4��C�I l�H��!鑥hF��UO�~'PC��L�yBA�>]����5� ,�LC�I�c|X�����0�8���	�JC�I� ��i0t:g(ȫ����P10C�)� Lݢ��
�_$ ��N�1U��y�!"O HRKԈ#�`y��u��ň�"O���j�*��=��mc� ��"Oy��! B��� �-�<9Ǵe�a"Ou��j��m����S�u��"O����
Z�V�8���E�0�!)�"O��9!o�+z8r�����Y��Z"O܅3�n�3���U�o���c�"O�}�4Ԉ;D�2T�!����"O x�m�F�M�b�!֦�"O|�S˚�h�]ї	F�:��h�"O40z"k�?tj,���&���e�'щ'��T��w1f �r%M0im�x�M����I�v�,*v�����e�V�a����{��A�ب0� )���ַ�8Q v.-|O�c� ��!�~�A�#ԇ1[(�9e�(��ȟ4 [#� �B�	��F�&����b�I�:}�>m��D0��¤i�<]��L)�F���E{��)6b��9���9����ѦեC'�y��1M`1�#�=-��p���3jb������@�X$V�J����n��1?A�C\6�qS�L�-XAT)"&����B1@tK�ڗ��-	��x�n�ȓ='������<9���P'�kz^������a!���H��e�V�U��ՇȓWD�i�HCʼ����
".7�O�O*0��
k�ȁB ���rGx "O�i���k^�j�A�1O%��G�'E��-�ĀfJX-6��0�DH*{!�C��	D�P)�R��V��P�n��d0,#>���ƻl����fE�6H�]���T�!��O���#)J)n	�A�u�>dƄ���"O� ����" �R98��GM����'�>���.��n�P���6�y��,<��p<�$L�u�p`fJ�	�2��#��r�ɕL�{҂�3p[r����ԧ���#"¡�M��'��;��%T�8�Cʉ2��1�'�ў"~��"��2aׄ\N���"�Li�'�?�P��{v��R�fS������0D�|���2J�J$[ԃ��M=���m9<O�"<��!�,�Pq�1F�\�����l�<�"�"U���4�2�� g�*p��	v��M�?i����<�N�{�,^�� �sf�*P�!��j�J:�R�u����H�~�'�a|�.#A�a�5N� @�ҕ���Px��i��ɗ�(B��Io�k����'C���iC<&����sd�.W�-��(O<�s�����q3'�R�!	�� "O�	q���V�(ysR'�; P`s�"OvG��:Fe��5&�
���W"O���&�Y40X��&@6ۀ;"Oy{�֢Q:����P�tQ"O8�+'��u0�j���B��}KQ"O\Yjw�M
-S��5mB�D�6�R��;\O� �n�p�����i��q��"O�ej0J�V��y��,'w�I0�"Oz=���)�A;A�޳bl�(j"O��q� N?�,H۵(���"O����g26�(����2�$<��"O차�\?o��|2W�E.;ٱ�"O9���]�{���� ^/Q$>�S"O��0Q�Q�<mh���]�ʰ�"O@���>��ԪW�֞}�2}��"O�9�SJ
����mG�^���"O� b��g
��J1���Yv.1�"O��3f�Ӛ0t��b��O�<o�K"O��`$���g�pP�Q��J�$��"O�m��H�p���G�����w�'�Q��u��u^b�1�O
�*>�(	ׂ8D� 1����|���G���Aq�)D��Ye��_U�\B �+/����f,D� #�	�����Ó�'Rw�Ik7cn�ڣ=E�ܴP"p;���aÊ��K_;mb"`��e�j�#G��0q\XakCI��8(:1���?!��6#�r-9��4+ zm1SM[e�<��'��poba� ��g��`p�
K�<Aw�]��A��.�ZY��lI�<Q`��!�|�"�)AJ����F�<��;5�^��â�?L��9�G@�<�샐L(�u�'/.�%b�o�C�<�n�V�u��	;#vy����c}�)�'*G��`�+�Pa,����L��ȓb;a�&���3����EƗ丐l�;��$!�O��Q�0DXM�#�C��\��' ��O:-B�"�tR��+���#����e"O&x!t����yQ#�\�\�*d"Oq�PAV�@h�"������$7�S���}���Qz&`�uET��B䉒Qg"�;@H�y��q�Q��:a*#=��4�䓱��O��t��F��JD����|�<�
�'K�H�	�(���ȿ-2���'1ў�}��'E�l\̀*t'�e�ȃ�Q�<��/N�|GD�K���:EHalVv�'�?��@*�;x�nat��N�N�7D�2�J�,�F83�B�>2,]����O*�$,�)�'+����Z�]�TTƌ���pH���hO?�*� �0Tq�Er�?,(xx�c�n}�(ZTx�PUMӘr�(��t�	�a��1�9�O��?O��I��'UT ,Pv��x]~���"O�x"�if���K�a@"���I|>a�W-	5(�ب ��W�g�~<)T�;�IA?�{����9BĚ����7PI�1�1��9�yR�֍x*F�q@�+F�,YaI�y��6�r�j�D�D9l�1�V\ �X�L���&˩'f��	ވ-���I	��d�<���Nvd@����<�r�k(<q޴R��5�R6L��< ��� C�*�Ex��)Z�Ѳ0��Y8u�9jE�O�W�<�7��J j$��i檀�s��i�<s
U�8�]
�$S�$U`�[%	}�$8�S�'*�:���Q�&��3���?�<��~66��wBW��Z�[ ��-=��=�	�s�QDE�(%�r)۳RB���ȓ�nő��
|L���]�V� ��e�yc"L�Pzؕ�'N���1��aM�t26'�}����(���ɇȓ=����`/���K0�ȩp=$��ȓK| �B��&D�� {R�N 2�P�ȓ[n�O'��z#���F�؆�>B-��kU"B���։��}"px�ȓ�Pzqb�K� ���Ɇ1�2@"���s���A�=I����$��L.�O(�i	r�&�N_^|U��.X�o�༅�g��E�`&���$a`S��>5W�Մ� G�a�$m�/ X�H����=����i�$�E�_�̔�1��2U��H�=qۓ+|dj��1�ԙIEL�$cr�4��)����*��	ڤ�_�v��EnZD������ L� �g��cܺ���G�;!d杺��'-����Ha�c'ڟ,Z.�Z���eC�ɣ^�B<��[1����*Z�q'�#=Yڴ�ȟd49Bc\$֖�HfC��0�)p"Oh��͓ a�����\3X�D�!&"O����+�	ǠaA%�?\�h�@�"OR������aE�v�z��F"O���� ������Ôo��8�"O�<(�%�"�S��Q;���0"O�ۆ�D�ĭ��		4p�q�E"O��k�GY�X���(IOzf��"O�u���  yDXB�%z��a3�x��)�S�sl�������&�Jq� �&(o�B�ɟ��Lh��wp�H��k
`FQ�=	����~�q�FS^"4��ɜ�.\�ȓaw�x �L�s&�a笎3m���ȓ$@��S���C�¤P�@��$�ȓ$�ƭ��N�Q,���@]�;鰐��[Yn x� ��Z�p�X����P��i��P򷃑�D�@����B�� �ȓ ����6������ �k:fE�ȓt�De�Jܿ=�2]PSQ�U~
��ȓI��(��g�+!����F�@Ϯi��*��h*�R}� �!%��91����ȓHz�]��T����WA+bgnU�ȓ'�.��.�F� $��R�p ��ȓ欙���=��X(�h�L��|�ȓc�*�s�QҀ��5�S�Ax,����ė�kh�ӗ�U�K�|�ȓu�0�D�]��(�T#Z��]�ȓ R�xq��A)�u��H"1_���ȓ<���0�������Z5B��h��Dp�;3Cb��VTnm�v%?D�p���ε8���a,D)RN��)D���a��o!�L���\�PF6�`�B5D�Py��ȐU�B����[�zLU��d0D�t!T�;�Q8���5��L���2D����R.�(8 [;ene��I1D��gE^$�r0��EAb�k�:D��ࣄS�j���R�B�S�(��;D�V��U�q�aE�|��"C�\$�y��ٶ-�����M�oD��R _�y���:Y$��%k:g��uR��$�y�X�\�D<h!G�))��2����y�_&����0]�!��k��	>�yD�/�4��Z��E��y�X� ���  ,5z��U�yO�#���c���Jq�,�$C�y )r2��� �N��!�⅔�y��LvUr�L�#9��Q���L�yr#ۉQ2c�N�;93@��M���0?�֥�P�*��
��u0��R _�D�eOQ�<�Nv"� ![0Q��lQԫXy�<��XK[���g��&m�>Ѣ�O{�<�R脪EA���
mP.�#c�r�<6�
O:���fZ�c.�)�fo�<�ǾV\� ����^���I�d�l�<	�c��3��vF�"X
���f�B�<Q��Ɖ:�I�LÊ�AW��v�<#�A�*'ƔHÁ�n�ހ����w�<IV����(RJ����[$L�s�<qU��?p���N�+�|;���f�<�4CFe�faR�i�9^��=���`�<1'mX�a:("�[�,�e��x�<� �)QAR���(
6ʤ����s"O������ 5��X���G"O,�����$�ҕ��<��K�"ObՓa՟D�H@Yj̕K�̱(w"OԠB4 :]�l��ǃ'�Z��5"O�|��)+�.X��4a{`��"O��@wf؁Z�� hP��q{6H$"O�#ՌM�SB5�2)�nj�a"�"Ol`�f�
*6�d�y��V	<\��"O��qGƶBb����"S	�`�"OVdzC�S�HQ`a��9Y<)�s"Oj�RDCO#$hlx!��H�!H�uv�'I�}V��)D5:�R��ANgʭ�� �#(�T"Of9��ɟ�o^F�1�a�1:�>���ɵ9�lʴ��6.���p��c�1i�0}b�B "O\i[T�i�M!@H(V �9�նD�0�����������F�)�й��/Nb������yB���4I����H�1#�yJ�I�<�~"�C2�I���#Oay��U�H2%�B��,ɶ�2c(���p>�+�Vʊ�uȒ!�DaH���+eD�;�ͅ!�2M
�'װEj��^p>K2�-!��yp��߆Dݨy
� X�]u:b?�&D�x��#���#�4T�S0D�T9��F�~�ݢqP�=<�ڶbU�r?d�����.��j)O?�D]�/q�h)PGS�u��1�4`�w)!�؝(���?J�hx"I�"��Ĉ)��y�� �JF��W�d��}K�����tC���w�|�M�#A�u���Y�$p��~�s��R0zT�0X2O�`0�M,UCǋ�mW��Jc�	j�B$�6AI�'���s� ��M�ϓFa�E��"O�)V�Ä}���Ƀ-�%Y ����'�>D�JY�=�ɧ���5�
�%y	"��s���eG���2D�Lb6��	QPe1�̭�� ��c4D���R���L��hJ�^��c!D�|�򪈥7i�� sn��C��%A�0D��QUȕ~6dD��k"�)��n/D���Ҥ�*�Xl�P���ZeH5�-D�
R�* �Dٕ&#-,eY,4D��ӳM��SpiS$�F�!2A?D�8qe�00_�\z0�О/|^��w�:D���CK<Y��͏�B�F� ¦,D��
��M8@�Vy��G�@~28��Mt���gx��kC
�%Z<��A��&`�Ť4|O`����B���$  ^���2,��7#�b!��K/lv���3�!"���ee�O�0�s�M�ȟD`9����1�����\��p��*O��Y���	}�`Y��K�l�S�!�`- ➸G��'A���+_x�r�ۗ_@��	�'Z��W�Z�kA���&WJ�9��2�)�f� �O��AmF�Y�RMK����|�4�a�'����@}򬈢J�(|0��݆w
 ����O��y��Ut+���+_e<\�[�hҀ�OA:�F)��3d�L�N�$��T�A���ȓ5{
@����@+B�zr��pޤЄʓ^��D��-�T�"�xtj�B�B䉵(p�J1�G$&���g�B��
q~�ւ�10��Ha�@�FB�I�(x���b%5/��Б*P�όC�	Q����� 2nT���ĕ0�zC�	n�f@BE�֭E�J�K�ă<zB��|�
2��S���#�.`��C��+P� ����-"�%�.�[ C䉢W�m��đ%���	�呾s�8�g.��E��?E�5�̒l�
 ࣈ͆\��3T�(�O�L��L�L�f�����ۦk�qP ��`�'����Y�� Te*6�<SNa� 	�6Y�p�w�	�h3��2J�D�'i�z@�O�: �Z��!B�=xPHyu�Ǵ|�\�#�Ʌ�#����ٴ~wj%2��2$	��=H,��n
�� @��D��Ir�Lz>��`����h4(�͢�#�>��������M�X�J�dB�I19���(�C6s�b	�B{���]�.�FN�'lq�r�Ԣat���a2O��X�`��.�B1�;_a��	WL]8���N�j$��	>Nh�����\H⑰6j�{���Ab^�uH8��U��k�����;'�1i���9^MF�[�z�1O\Q���!0�<|j�)�pV �p�I�g�(zC�&t�b�Y�`�ś��Øq��C��S�����E耥$���)�j�2f(q���)[�
���N 6K8�qs	�1GZn�:� ��>��Hʖ	��K��ԅ���P�$�d��)�|1��]�p�I"��?���"�J��?K��������$�n,u�S�6iTY����D&���B�Se:�h���Z�F��B�j$2E�ӊ4oDq�eF!�NDQ�D9Ĭ��rtvl"���_�~2��JJQ��`��wk>�2��ĚF� ��U�O�/ !I�&S�ULN�i�P�_�(���S�rg&�b�dD��d�𸳎��+� 5�W�L�>��Gx��O����.ο)�(-���͎:��KpfJk��d���@B��uB�W���F莤,@4hY�gt��xϓk�b�(#
�,�6h§#�.��O�mɖ��mj2 9IX�`�z�	E���i"ѻf&��E��AV��;IRPC��:eU(W���,4��u�j|��J�.��|hD+H�	��q���j����B뉆E��lÐk��p�x\��������y�ƍUP8�A`}�.����T��Ig�I�zj�pe,J�^ʰ����;a����T̨4ɕL��*i�+&h��xEl��uw�|�7D�0�M��Y�D-p���&�O��=�'KԐQ�\�K3R�7�Hm��BV�N��a%�0T,�YC�4LO<!�B�`��}
�&ڲe�|@�'�����X�lÆ�s��@$M��s7��o: (�-͞}�E��mAe�<��#�7��)ɇ�XC�<04-Z��19�mPf���7�x�2�Fz�O�@�CEi
:aHC	Lo3���
�'�����_44'��0r(�v�F�	�Jٞ2�U[C��͟\p�
�����{V0��.��=��`�T�V0z�d��Ɠ�^��/H�.�<�a��O����ǭՀ9��$��/ ������m`���a"U$�(�A�JʫO�z�Ĥiֵ��*��<q���RZ�̓�K]'r^���K�w�<Y�	9E .�K�Q�dϪ��t�t� %��)�'���a �vg8��f�?SJA��$��,9!	�'Y��YF��0�ȓk�,p�Aǣa��E��C?�\Ąȓ���r���~�
����ϙ�����`t��*}P\�[ ��+E֙��I�H�U��P�b�%�䵈a�>A����7k0D�L�נ_#��%�*��$�4(��*�0�tF�T�O�Ι��ɟ���Gh
kӚ=
�'/�1��̕y���a�K�^�^TY��/b��'�L�����>a �
��p`F�� �rLBLh<!p��un��ր[x;Fx�<Ӷ 
W�h	����-��`6k�I>�2��؋@��y�E&�b�-XK}Bm�;'�X= DhW �Μ� ��y2A�'{~���F�"y���e��;��#|���-A�u�#җ38��	�5Dȏ#����gA@x�<a�Fo��L�d�8R�XrP��-@�|x�v�>��@�#����=�:��q$�%,B�x�̖\zC�ɧj4R<k��M�U���4R�,�&#D�!��ye�'�\�� �%;b!ꆫŒ  t�i
ϓ;h9��KE"v�uhY�#ꅠ>�� 3�]�16ԭ�ȓv����#
�p��t(�!�>����<!�������b����.;��1�s�BH�ӒH�5$�!�d�K�����]�mB��D��%F��x���Ē#�(���&'F��rV�H"Hy�a;��J8]��B�ɬDDm�B\�{}��F����B�	��XK&� =E��Y�C�1&����)���],�?%�e�Æ ɔ�HRO��wa���R�+D�,��V;�$04�Vk%�%k��`U��|��&�g}rK��p���vk
no`���A����=��F�XF��ZU"�&�)9<L����بS�����$1h섢��o���(�
�]�T&�14� e��<�I$A�<�Wțc}b)̥gb4)�ԡ��|� ��t��!9�2,�éN� �H!B�"O���p�ŌN���(#E߯8�DpP��8P����Oz�Q�"�SR�a�������Fc��U�~�ӣ��.$���7I�^�<�d�؇ ���C!j�B��,iGLD�M�U��?�>��c'�D" ,CLr�#<�G)Y�$i� ��+Ӽ��D�x������7)(:�$>OV��5B�0Y�T�p!+")�PmU�Y$PPhSE��a|���G�4�i2�B�z�!�N_4��'ɚ�*g�B�"5�Q:�	&�9~�\�S��d�W��I��8�@�-0�ZB�	 ��\h�ᚒ_<�kã���6(��JM�%�O���C�@��n�:���Ǽs��F�{	N�󓃖j�u�A
�C�<Q�◒)Q�%����m��\����w)|%���ܰ-n�͓:���S�b�-[ʣ<��61+֝���Ö?���;R�t�����%�u����#�'ِ�C�>����db�6�R�KY <S��� �X����?c�d�Ǎ�/j���ʧ�:�I�~��}�6���<�e5c���ˇj�~´͋��J!�7ҳT��sA	�s�<Q!�̚?e�U!J]�&%S�	1P̤�s�O6����K�����x�EZ5�
�|˰�c��A�s/0����7D��IDKؘ�\���ؤ�
�2'IX�B��^C�䀪p���?�'�&Aa`�_:��0�â{p�a�'��V)Z,o��crf�F�����ݽd����F�P|X�@c�G^�N�8��N���B��+<O<�+0
��N���O�lS���!?(F���D��Eg"O�|�,�0ZK�q�F�Y��[r�|R��Z��k"	�g�Ow���D{᦬_b�R��
�'�4��4)J@u�ٴ�F*4t\�"�әM��'uX�:���rb��Hȓ�i�.g�����m&D���E��s(�a0F� �~��q!8_�T ��-�O$�@p�K?=�P�-�z��("OV� ���_2h�ڐ,I�
`䘳"O�hС��	��b7KP1���
�'�@���PI�Z�d��a�D�q�'=���fN	V�]P�b�b&\�y�' ä��6B�t���'X��"OD����މ�H�۵C��2@�lr "O$����͗2����#��|`�)F"O�U�F�� %o�4�� w"O:1���SY�QA��	%���b"O��*�OE���t�f�+Z�K�"OȽ,��x^�0*]�?��a�S"O҅±�R
\��Q)֠�:�@�Ғ"OB\��Q�_>�ز!���c�4�p�"O�L��F(d̴(Em<65dH�q"O*]�v��$�eӁM�{+P܂"Oĝ�ŝY�ĸ��P�|���$"O(0K��Щc4���kH9:��"O�' W�s9��k�JK��dғ"OT����	|Zȸ��o�&y��"O"Ԉ�
�+NclP���77��"OFD�M���R5h�ÕZp��yR"OT�S��'� 8s��ÓD(��"O|8�vf��XTʑ��[�/>!b"Oܽ�6�^<>�l�D�Y�X�Nk�"OZݑ�D�X�M0�	Tk�x�P�"Oz��##�[c�	
pΊ�g�v�S�"O:1��J��PQM��OG08`D"O�@��L4+��u@���W��Jq"O��xQB�
�����31��D"Oz	�gjZV>���8/���S�"O�9 ��H�	%~���v"Ob�s��f�Z�YV�J�m{$ᒗ"O��2"�� Ҁ1p��MG�P�+�"O(IRu�m�~;���xCV�+c"O�[@	�V��z����PB�"O�A;fJSM��Q,��I�"O� ���OĬ��M��,�H*0c "O ���L�BX���T�=j�2)`�"O11`��,����FO�\���"O��YAQ\l,����V݈T��"O&���FK-�-YoU'&��j""O��,6��S�,���$y��"O0����r������9_H9��"O�t��eF�أ�	�W\T��"O�%z���L��� ��R�i0�("D"O"�u���p�'�_EF�j�"O��jƓ5c����7���Y7x "O���$�ܾ9�1��
D�I�F"O$��`e�>[� ��P�y#��-�!�9�$�)R��ZA<�P��9�!��D3A�X����
i3X�נ�>s!�D0��aւK����OY�`�}�ىb@	��*>F�,�K��	�(j�@�h�Nd!�D�8/��\���Ē)j� 	VJ���Bb��XE���w���dTʭa6�L�]S��9!oY9�!�d�>0_���Eg��YL�{�l.>�F����(^s�t���py���'r�\qU�Қ7u4�����(z�'�>̪�n�d�:�)B(�s��K�'�f8�u	�G���K��'}l)U�U��
A��;_�h�o9�T�c"LQ�/$|[7�X�YH�0&DL�c#~�:�'��t�Ə�)�ڰ#��� #�H��d�g��H�6_�*��b?�(ǫ�=6Ac΃XY��b��;D����Y�z(:x�c�
w��$�7��I���G"�4:�Ҵ`/O?�DB j�0��Q�3Cr��V�y�!�DؤH�^%�,R.Z0m����"+c�d�c�f���(J&���d�\ڥHiϙ�q˳JZ��|�m�+j2^��-E�~���
�r� �+̡D����7O*���N�X d� �%v$e{��+?����RX-3�n�� j�&r��τ(�a��"OD���A"`����oB 
`���'�,�A�B�|���&!^��M��&��ق��\+0�xC�	�\~�\KT��'���Yu�čz�LC�I `a�Ү]c����Q��D��B�ɏg�<�ː�,(&L�򁖗k<�B�I7b����/S6�:4��W���C�I7{�%r��O&�P����(wsnC� M���EOύENi(���B�It�<	z�iŴq�:�Ə��r��B�I�v�� �q%M'e`���@[;O�dB�I������ƽP��L��ݠTVB�I'p&���7��X{c���B䉾ZG�50��"F�2yB�b
$��B�)@0M�fb@�k���˵7�*B䉇?_:��S�)u�����4h�C�	/Hc�x{�J%>P����=��C�	�f��҅i/Q�� ��� ��C��Z���9_.E������C�	��Z�Qv��by���GG�|}�C��;l�J�D��	7��l���L3X$C�I�{��Uf%���Ƚ�C�	/ ����5�ں�(21�K%�B䉞4(5ic�ܑ"ܜXR��ˍ��B��,]	H�)� U�j��p��I�B�	�LjNXX!$D8�@�:4M-
�B�	�\�\X"�˅:j�~Q�� i�B�I�%�l���M�I��0�bRm�HB�I:������\(�xP����7Mb\B�	��FUɧDS�g[l�"`d�i�8B��)L!*��nV�8�hm(�MO�m��C�!2A�	W�_,N�� �X]\�B�)� �QP�$�01X$���ӃY�t�
�"O �
�/��)�t�T�H�;��Pr"O���3`�=�tX�aE�%�z�p��'�����Q�)&¬�ԫ&9Ā��Q57B1��-`Us�P���!@�MB0x(( E~뚢m�H�kF�韚i�^�)&@�,D��SC�.D!�D�/�!Ѝ��7rڝӵ��O!�$ l�
���N.]�\t�-�'I�4�;3)N�Pnn����H�(��1��c�&8�4��9äq!��ӏF�=��¢O,6-�5-ljP�Q���3�ɣ����ݑ0�(�R��>������"p�H�d��[���e���v��n�CĀ��"k r�`��'ބT�2�Q�g�4�P �u�ܬэ�)�	���
4�	����de� (x��i'l�.�J�S1̇�y"�\�d���Ï})��y�FP�~��H&r���M�3��B�r�O*�uZp	�9 ��MG蛶
�LX3�'�r<�.�����	-*�ɣ�(����΀j���PbR��3�I��<@s�KQ�]I���	BA�����)kt���(x��Dy%{�9�݅X�����ԽNt�����Q�x��l�(kf$���ڒJr�@�"�f�LMs	8TІ|��Y�)ʽn:�6ᙖM���O/!��K�_��z���8 `�Ǝɯ�剪�
���[:%���«�F�O4�)���#n�<��mJ�� �#�'Hȵɲ�B����Mȿ=��$.�:�$�而�Y�0Ɂ��!�$B#�SY�4`P$1D�Tr*��s�,��ズ)i���Ҍ�O`�+���!ΰ>I�ńh��@B�L��b~��&�v�<!� ��(�R��mзak���	i�<���L�LQ�-��ws�EʓM��<9��ƺQ P	ǡJ�H�R���Wa�<1��A4`�$����ސ���[�+Cz�<�5$��K|Y
�x�h��"�R�<���	�bJ���R^�;�I�<9D��T�(̡2���]���D�J�<�C %F=m['&N�M�R(@
_�<�D�X8`7��y�,�6�1���Y�<�'ہ|��@	�MMMZ��O�<Yև��Z���ZFҽ� �@�<ad�ڮB�Լ°OD�Pc1�	�~�<����.<�4��L{���I��u�<�f�ɆH�8QhsCӫD�t�)7/Al�<��L�&Tb�k
�&RʈS�bBi�<Y��Q1F�p����݂c$��A`��hx��A���=�sHG!=�"�Xt���B��B�I+zjU�d��\�5:����b�0*V(X ���F�4�I�1�����ɵ?{�q��)���y��XB�����]#!L�Xi��-��M89}¦W',]��O�n,w.3r���ʝ����ƓD6�`��7? �j���D��`� ��SDDX�C �O�!`�U�pl��V�	�dp��a�'rf肖�aw��'g��Q�?�4��h.6A�@�'�� Q%�%g+�$��T��R8�O>��DԤ�J��+�'���!B?z����鞾1���ȓ �n�Y���S>|q�Qm���>�kЮg��~ dUb��L����肨G;����_�<�r�`�':4�TXˀ1?���uEW�2[� �'����0�#o�^Ua}�Ȕ��S��L�c��@8A
��<Y�g�?`��Xa*�>��l�<-�P��1�6�z�;�e�<鵪��?���q���&h%˄�g�&`1�Ԅ'��걛#E�h��s����l
a"O������>'�()���%^��t���ʩ)qO�P���Y���F �R�	J��Ц�P�C�&D�tX$fwF�X��Q<<Z��kf�$D�tJ���BS�H3r��	��Á�.���p:�����/5��%YS&P�=�89B���#r�C�)� �A���.��'��!j�9�B�^%_�t�H>�b�>�¯�9�J1��3��m9���v���)3	]�R�I���k��7r����Ɉ�@���ѪL8^ndg�(�OȀ�"��cyx,�P$G�D=�T����5&�#n�>I�aH��n�� Iu>)�d���n�����.Ɠk�W�2D���M��ANZ���D� �Y���Q*]ܺ11Ą��T(��S�p�J���)_��y�'3!�6(�Q���x������y`�?kr�X	՘�~l���]F
��㶁։q�\�i�'�8,l��D�Gx҈F	$e|�x�Ip�P�X��S��p=A��-+N����m��r��&�h�� �a�N�CS(v�&�rG����D\��ްz�Փ`<�)���BRqO؀2tN�"/�L���'M��p@�բrHA�'��୕*y8!b@��T��ȓ~lK~����J�f%��%`�=0}V�w��0;G�) k���c�	��yW��9Eq�}�ե�?Q��A��R��y"�J�)ޔ�H%��,U�jĉ�J�#G���"MH�Q�4�B�'� 	"�J�*ր�Dy�eS�B� ��Q�ZA2����p=�"��*UW��	���Om0tJP�`�J*ғe�l�#)I�A�
�2��Z �>�r+�6,����N�
�ꬸ��L�:)&5QT�J-�y⣔<�>���b�R���8IN`��h�K�Dy���Ƣ�y2��&�������.@|2���T��Yy�￟��a"�>�0G�ʼoV�(D����
0�M��y�ǅQ^@�u�M�<�,=֍��bt ��!}"ۦ ��l$܄����)z�(��Nƭ�2�Ɠq��H)���aq*���Eh�8p����B�"F�2�Oe����i�ף�*�XђR�'�q�w�T(�P��'t@I�+Z�nl�Q1��^bdԍ	�'if�1o��"��̠q
	�]�� @N>�Q��.^��8h�F&�'m!�M��FA7L*�8RTGL)���r�`�0+�+w1��I��N�
�J8M�q$��W
*�g~���t��D(�I9&��P��&΋�yb�� �h�@"��{�d�c�R�-F��p���0?�cȟ+L��3��h�,�	��M�<a!/O�i} �*cR�I��a�m�|�<Y'.I.��ҥ@y�%���Q�<Yפ�Q
���9�L����N�<16L�.� X�K�M�<-��·q�<���[dtI�lխ?\��!o�<1� �iጰh��Y�K�k�j�<��&���+�t�HD
�ȓPs����Tg?��$ꙉ>ܩ�ȓa������!R�*a� O�qT$��pP�|/�--2�kҵ*�����
Xi��Ħ�:T�I��v�t0�ȓ��@���׸ tN�*S�­SM�������#`��Zq�&HMA4���E��2&%�:!�Q!��e����2l����̐�{����߼|h��ȓuj�Y�-�aV�놡�7U���ȓ<=��;F��mG�	cn(,�Fh��u��R�LD:-���;WjB|M�ȓt��e ��H>dFTk�'��x�L���$U
�U#w&�-�+Kt��,1�)��$J(N�Vh������9�V�a���A�}z�J�R(:���o�(����uV�����*L��ȓ(��h$��.H����c�b���RI�	�N.D)��@]�?�B��ȓ 1�gkS�s4���恕Y���ȓY8��I�`�.4�@H���'tNم�	�=����M�p��|����8R��)#���6b�B�%z}v��s��D*ve���Z,O�B�	���uB�K,(V$�(V@�B�	*ct��!&ƌ'_�r%��/~B䉼!��=��Ġ0��1$���I`B�)� T`pqbU����B�InЉsG"O^���ċyS�a*�/JFh�]��"O�m�pƚH`��j�m=J]0�"O��
sn�d�
�aE'�Qc"O�P@��+�����I�M	�yz�"O�p)T�
��  ���#�2�
�/OB�qO^��ç�`|����2�6Q�C�u`��(�����En�<�2�'k$ܠ�4�ۓQ�&��oضT���'��IR�	�0m��ᓪC�J=��Oَ\N�4B ��z��I�|�t�zR�Q�@���S�O�"�yt*M�wn��NGKO@����G����a���tP��4O�?)!n]?s����C�{����v*����;GJN�z>v����i�L��Or����J�L���P�'%�U�&H�� �ܴ�V�����8j�� a��>��)���2q�D����.�����*��-j��(��˩�?E��DT��dʕtquQ��>I��IU��0N�^�IG�O��	�'0wH<�'.�R6�QYH�Te�0vJ8�7�[?ys�&*����)EZx��	؅�F��!R�^h�B��7*��Y�LT�a ����O���iF`�)o�����W�}���r-f$�����+^�~1�'̎��0|��&O��$��KG.�V�����Zo@t�4�"{�v�:�I:[޲���S3E)h���U	z)H9c�i]>(�x1[�����Q'u����çz12t���M~>��Bn9F�v�S��x@BJ9I�����OA>A�DD6ސ�2gi!j�+�'�Zp`����7�$�ǅ�f(fh
�'Ǌ���C��p�Ҧ����8K
�'I��!%G&z�0�E�.3=s�'�\����4?ld"Cc��#r����'_B������lh8"ʜ=K�Y��'b�]����'N����镎EW6�c�'����Ū�;&�ˆ��?Bq�(H�'��в�Fr�E3�Ǻ5t��'���*@�$ϾX8��4s����'Î=�I͎10�d	U��ʐ�'�=��\+u�q��ڶj<ة�'���y0�	�_j��2T�Ӥ�`�k�'�d���A�5�t�#"F-0�ܣ
�'r��r�OÀ}�<�#È}3�t��'��Ġ爋�RB�<�aM2t3��[	�'r�D��H\�� ��.�n[0}x�'��]АbZ	R8n�
��˷Y#�=��'��P8�̀>g�2 ����6Mn-�'�l��k�OU�L� F�x7���'@p(�W!?� ��g�@ l����'�0
��S+�h�*�L�&8g�j�'븘��EͻN�;viҶ[��Q�	�'����& �+܎E�UnH[H����'�Fd'����@22�ȶZ*��
�'��@y3K�9�8h�1 ֽB�<���'OR���R���HR&˗<N  ��'I�H���V�%�a��9C4P��'�p��reɉocD�ɑ��=�@5��'����! f��Q�!I��*�j�X�'����gV"m�t����Q$(-�� �'� ��2*Ϋy	~�X!gH�1/T��'vF���b�8#��ː��6)��y�'׆� V%X�o�D	����12�QY�'DsĦʖ}9\BG�As�����'r���&޷|��yS��Q1cp���'G���q�M�r>��Z"+&&�����'?�x�5EZ�Av�Y�d!��2�'���JF�S4xC2��lf�S�'K"��D�Ѽ*���(�,(lČa�'`���g�S�}$�
�i[��Q�'�d4�e��(b�� �a�5MOJY)�'�TT�D� 'Ɋ�CI�<L*���	�'��W	H2/�& QcM�U}j
��� ���]�$]ֹ��g 7*�hy0"Ob�C#�=�Ɛ�fZ�0����2"O\�����(p��Q�BE�?|���p"Op����_ϐ)�ecJ*'2��3�"O���V�Q��	#Bl�@!ʃ"O^]KW���4�H@Rq���"B"Ot��$-IR(b@��ꓠo�b5�G"O0��҅5}�h0�O����7"O)����|Yq0o�	��Mx"On���(ګ&����'P����"O��2e�ܡ�P�Q�n�q�*��U"O �^y�(m0bm� ����"Oơ�㄁5  n|sT�N�U�~�pP"O��+�bةJr@	pN ��d�9 "Od����2
&�E0��G�4� HH�"O"�Q1��B4�-h��&E�pd3%"OL�"#���`?d��A���f��t�!"O�kg�a��IB��9�RdS�"O���0/�#a�����V�_]���"O2��e�H�>�a�G�ʂ}J�� "OleH��@^��܁§�./xh��"O`��ɸ86�Hq�'��4���F"Olv�N�
�q	Y�35J�"O����IH
d�G)�(���"O2 ���V�Y �g �U����"O��JT��bFq %h۷E ��"O�t�'GH�&��0���Ч7F���"O�I�I�y��l�L���I�"O�l��J� �*}:a _TNI�"O����=`���3 N41G`cf"O��d*��9��؆�(*L�+0"O�������F`N�y��"O:uP�ʆp��t���5ɶ�"O��k��_!�!��Nc[�廖"Of�BEf�M�� ��g�<I�)��*O�
P���gj�C(ĬP���'�ޭS�̖+<7��*E�T�h�Ԝ
�'@B`1Q
�����$.��e>ly
�'�&���j�P �7J��(�r�2�'A�<gk�yH-8��� (����'v2i�5C6�{vk:+�Ű
�'#�ЋT�ݮ�V��$H:<�B�ɕ)Ύ$CMQ�
,�DȊ ��B䉅t�S�O�7� "��)G�pC�	��L���.��3�]�(JC�I�^2
��&e�x��o;1xC�"O,�Y:!��dH��e�7�B�	�Ed�l���P�#-����*6>B��O<���ㄓr�6�p�N3	�B�I8�~=�j�+G���C�	�-�Q*%c��4����LwzC�"H�`a[�9�&AnN��zC䉞`�̝
��еK�V��g��>sNC䉿n�P8�-[."�іK6&�(C�ɼ&��  e�F�\c@�"�Aw5C�	�d��(��C�|A�b��^�,A�B�I9m����J�#Zf�p�g! ~��B䉯j}�` nB�����&R(ԦB�396��c5��\Yd)%焐uX^B�I�R%6�[&���G�@i!�aX�n�vB�ɦ+��ʢ�	W�@��$��jb<B�	���r'ҡiD2U��FU!4�HC䉤e��̨���O_���E��	t^C�I�y��&m�01�h��Gg|C�)� ���0�ϴ[��T�7��j�<c"OVq�C�J�[XZq$لܨ��"O�1��_^7��y�I�\�
��"O���,@l�8�"�?7�p�4"O�S"*5^Z�0����t��Q�"O��)��Q�v�|h��"_�K�h�v"O�9���b=:�����v��9��"O�$�RʈB���BH�z�R i�"O����FD�1�Z� `x�"O�*V�̔W���B�e�Ջ�"O���Ta��l��$�Aפ+�Ȉ�"O�<a1�W�5� ��E@V c|P�"�"O���2�_8H�p��mRdal-W"O.�q'��50:š0�ƎvU�-K'"O�⒍C6
�^M��.͘3M����"O�1�R�k���K*Q��X�"O���L_�$���s�P57"h ��"O�9tG�C�>� �'F�\�&��0"O202��.��X��gCu�h�`�"O~�pg���ж�G�
-x ��"O�Lh����j_���s L�w6\�q"OB��RAY�E�4���P8��yA"OͲ!^�,ZqIc�Ĺh��"O�� �F��9PI
2�����"OT\�BU
�u*Diß*�6��"Ol���EhL�S��G�t�[�"O.��'�r�V,b�O���ˢ"O�Հ�P`�XyQBo�*�"O
x�Ed �1��ajg �=%!n���"O�H
S�0U|V���Ů{K܂�y2D��a`)!��6�D�8 ���y��ż%&�8�Vb�0��I�c�L��yb�
��X}�(��)L��hf��?�y��Wb
F�����+�b�9V%^)�y�̟�a���MЖY4� a����y��;��@&°O�5Z �V��yRm>O�h2�	�p�.e"%�y2�
1Q4L���CS!��yċu��\r�IT�A�@Lړ���yb�FY�B��wnK�$�
Q� �1�y�iM�g*Ȱ��ϕ�M� Șv�_��yRI�p�m��E�F�ha���y�I�"&�^A���Fc��[T��y������>�P�y�I�y2N�u�>ܱ �.f�Ȉ�2��yRќ/4���ǗR�0�� �ӿ�y��݈1��(Rs	�)@��]�:�y2M�(�	6 �?(~���U$� �yb�ɗl��Bc�ȞL$�bg^��y2�	10�L)ɣ��K����D��y�	 :x���6K���[��yBiTAy�nB��*��.�<�yR֕4�"x���%{�d,[G�>�y�יTI����Ĺ�F�[:�y҂�e�H���X�MQ�l	�g!�ʘ��iy� C.tdn$�7��f�!���oDųvKt]�YJ"��C�!�d��|�p�%�W�mP��gG9e'!��P7�$�cO#{��h��DS9M!�d�@��ٳǏ6��\; �?!�١c���qA�W ����%r!�$�&r�pr��)|���ҍL �!�D��Ǩx�@Ia��M��B�-�!����Z��$����,QƌD4I!�� �x��~�Nx�
O��2=b�"O@��ffO�ji�`���������"Ob��7L�!� 	�jH	m�t���"O�� sߝX���2�P�<�Y:�"O����R$wپ�
�IT�j��;2"O��[�+�0��ٛ @�2��"�"Ov%b�/l'$4�r�p�"�R�"OBá%�(�թ��@�d��0І"O���d)���Y����#"O�E��윧Y�
��6g� Խ�3"O�t곣��>�����,H�L��"O�J���֙�tj��`�n`��"O4��u-�@N͓fi�=t�P6"O��i�ʩe�d� SG�1rp�@�"O a�G���;n�0"Ve�?T�#�"O<�5������� 4��Ȩ�"O��B2,V$1�Rl�4^�B�	�"OB�y#oP1N5�Ě���U��`	�'�>�"4���k�r٘�	�	;;��q�'��5��!���=җN� ��s�'�<���I�����4@�L��
�'(�����H�����A�����'����i�*Q6����@Y�'�}��'��4S'�GT��ض��wa���'_
�"  ���   �  >  �  �  M*  �5  :A  �L  6X  �c  o  z  �  |�  �  w�    �  ]�  ��  �  J�  ��  +�  ��  &�  ��  ��  �  W�  ��  "�  � p E � $ �* �3 �: �A �G <N Q  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#����!LO� ��!צ[�n�V��G!��~�҄�b"O�%��$Vݞ�x�` 7${l�"O������$|(�bE� ���`�"O�4;A��c���A1�R9�\+�"O��:�E�M�&���B��C�"O&��T�Z	/ �x O"g�<!z �'3&8lZ"i�L�V�У#��)!%`'VB�I�`$���(E%D���(H0�?�t��E_襲ү� �bEx7�ͣ �B䉙s��u�"ᖵ?�z�P�(c�h�'[ў�?�v�g���ԯ�J��xhsL8D���D�,{�TͣE���&�(��6D�����SƸ�6�f�8H*f2D�l:�ЧZeN9�2@�PpT@0D�n�X�\0*nJ��{�/4�4KbIߤ*�pQ�͔�-K��)�r�<%�1��E�o�%V��n��+�-��&��C��L���5�	-0.24D���%
.�����AG�R���-}A/�S�'}Ѡ(�qk��j�����R	al��d��)��  �d�jDeN�mFM�=��'���i�<�*E��#{N�Q�	�'� �,�x4��`(���^Đ�"OJ-��-��h,ч&�9`�n�¤�'-�O�y�JW�����w�b}PEM�+�y"挤$(��B���p�L1���^��y҆��!}���B�x����mÙ�y���l�f��wpu@�.A��ybD��~`h�� � �څ�F��y�X�\�j��#C�?�ج�Q�R �y�V\QR.�( B�TB.���y�aǟJ��R��#'ABX{��=�yr�L�o�8dpe�;!=�8�3�y�hө&�$�R���zt�����y��J�aA��b�<	u�Lh��H�y�+�9�4��D�X-��\Y6 ��y�)�mv�pr$q�M�U�^�y2d?��̨�G Р�)����y�Ǚ�hV,XLY�Pu2%��/�y�ʊ7S���c���޼)P@���y2��=`di�'MUy�V�ǥY��y�fT<a���Q��� �v���.=�y�J֜'�D�;e�� l�x�����]�<�#�:c���ۓnծI��M���i�<I`!�CC�="� 	4騜���o�<����7)"^�c����8Eok�<It��/NQ;Gi G�Z�k�P�<�hX9
Դ��P.Ż. Yy�#�J�<!�ŋ3��s-Az0�+�^`�<RMڤC|��'Δ ]沬iQI�_�<Y�e\�6�B5�w&�$W�$h����p�<ydiO5�d`VN֕$X��aF�T�<!C��K�fec�A
���AS�Ke�<���@�>���y�b՟P�|��F�F�<����	��������.m�3��w�<���	14��$C�k�2�b�cl�<Q#l,� �P#K�,eV�i�Kd�<v�!}	PV)�Y&�Ih�_�<�KU�3F��9�ޜv`���KL^�<�F�C���ڔ�.]Ʈh��nGZ�<����]��	3�Jۓsq��� �m�<�5 ��7�Nx�&Ï4&��b�Ǖm�<�`":._Zt�"!Ս0cV����o�<�Ɔ�*o'��z�*\/��1׉Ai�<� �	�����iR�JM�1��І"O��8&�?s7�����I��Lx0"O�rt�S Y*P�a��$M�Ms�"OPɘ6���^;d)ې��*Jp\`�"O�e�牂��^5;�I ���)�'��'���'vr_>����,�	!K\j��s(ԛb�SL�D��Iʟ����	ӟ �	ҟ�	ß�ɉr"���bM8����R8,�I埨�	���	�@�I؟�	Ο�ɦX�\`x�aZ!�p}��$Et���IҟX��ӟX�������$�I柨�I�lT �(�P�`뤈�ƆC :�Iޟx��۟����,��ٟ���ß��	�m�R,���1v�\9C�rq���	��d�	ӟ�����D������ʟ����^wp�I"���i=*�:4DZB�p��I՟�	������@�	ҟT��ϟ���IP�]����X�|E�A�	�-~�����I����ٟ����,�	ޟ��	���|�/�̑җo�>8�)���|��ן\�I㟬�	��H�	Ɵ �	��n�`�#÷_8"�����9H����˟�I���	ޟ��I���Iß��I���`ūR�5�v��ՂH�zq���I`���P�	ޟ0��ԟ,�����Ɂ+h��A��'(���DT�Yn��I��	��`�	ޟ��	�������ɨl�49��+]�Y1<�C F: CR��Iܟ`������	ܟ�������۴�?���Y}f�å��/;z<"�b�g^HJ�W���	Jy���Ov�o���,���,`Ԅm���
��N�Y��"?!r�i��O�9OD��H�:D
��Q�^b��P�^���OlM�Q�e�D���d��*�O�^�blG�\m��BR�ӟ�t�yB�'���q�Oi���3N�#�`ґhW#:���b�&��E�-���M�;y����DKӡ �N̨`��D�8���?��'�)擾�IlZ�<��b?*����?%{P��F��<��'{��$U��hO��OHi!�ؚ�
���N�5����v5O�˓��A%�V�\
��'��P#΄82K��ʋ�u^d�b��$o}"�'�;O|�2B<CEfW�Wl>� G�4�~��'�b��` @����d�Zӟ����'��<�&��1Q���dc��d�����Y�@�'���9O6��A�Rv������B��I�:O��&;V i�O5m�S��|z�>���"B��uz5�@"�<����?1��c� �ٴ��De>�@��\���H�B��.&H��2�0�&�>���O2�4�V���O��D�Oh�d� J'(Pz"V;� $�,R2�t���OK�̜&��H����O����A�3?Y�B��~�a G�|���!���?��0���a�f�m�k��D�O���fn�hҢҘS[d59w�ź<�lt��Ǜ�L��Ă�OL��sF7Lx��J�tݱ�M<��^��±D�r,ݐ���`x�@��N�@�Iß���ʟ�Ky"�q���b7��O2M[W�fT`�E�i=F����Oimh��T�	럤o���Mk7	T5 `P�J`I*6@\�5 ��"�Y�ٴ��D� A:�A:���������A9Y�P�Z�����gΈ���$�O:���O����Oh�$7��h��qJ�=Y25���چ4\\A�	ϟP���M[ת��|���Cu���|��D�7(���g҆BcLE"6N�4R(JOƝnژ�Mϧ�Zyc�4���ŉ�� Iʵ>=�p!d���e��P�H�?�?�Ӄ"��<����?����?id�V�*�pQ��:;>Z�R���?����٦Y��.�ly��'���aF@����g�����ڶrm �@����M#$�i�bO��`�5��Ȟ:��};p�Y�1������>�ec��Tey�O3�����S��'�j��?}�t�4̋�[V�8�'���'�"���O��	��M[2a�k�ʕ2G%�,s�J��ʕ��$�����?�3�i��OԵ�'֛��2&�|\�tj�TX�Lq� �.vql7�Ϧ�j�ۦe�'�x4����?YqsT��Ps� �3{� Sn�\%�PRB|�H�'g��')��'��'���B �mZ2�͈�s�ʍ��[޴5��	��?������?)ǰ�y�ˆ�4T�:�i�ҁ�'i�_�n6�ʦuJL<�|B����MK�'R���:t&z��aO
1n[�}��'. �A�×����|�S�D��ҟ8�QN h�NqI��Ą�ȴ�5˟(��ߟ��cy��s�,(Cs�<��yX�d��(D�h �KZDO��O>y�A����M�Q�i�xO"��d&I�4_�� V0��T���*�@���Q�b��v�&�2��D�RiĂ>�x8Ȁȋ�~�� C̟,��˟h�IßDE�d�'�VP���I����SRŤ��7�'�@7-�%VQ����O �nb�Ӽ���o��3��ِW� �i��<�7�i�t6�����Ō���'�&ih3I��?������F�.`�!��ڌ��'c�I����ӟ��������A�ܔ2�O�h�z:�HMn��=�'�>7͝� k���?YM~"�|�����4_6 �h�A���5C_���I��$�b>� ƫ��RKPi�CE�W]B�p�&�(N])�Ty���$�\�ɒo�'��	(u��)��l�Q3W�Y�9�*���ڟl����(�i>A�'�P7M٭@����$�R�`M�/��eBAZ2�h�D�ϦM�?)S���4Y�f#r�҅QP#��H2��K�
Lն�0��V�Zn6�(?����{b������'��� ��{���_4F�
�;<��PW0O���O��d�O���O4�?A���F1W��M3TΒ�L�$}p��ş������޴;��x�OL7�6�D���`M��$V��
#���9���O����O�)��>��6�3?��;���i�%�������|2�i�%ǜ��?�A�6���<��R�D(;���#V΅�_�����U�O��oZ�D*�(�����I@���ѥq��ÇB�P�B!i�c�����S}��'�b�|ʟ�%� @�bΤy��M�)3H:db"�X""fy���]����|"Ł�Ob�L>9�kGQ�|T����	SuC�l�~<	�i�xUj���X�`�����ݒp.�v���'�7m2�I�����OqD�ϸ"Q��� �-t��a��O����R�>7m ?��+
Y���(t�A<ڔr6�ܥ#��Q�ah�\΅���&|Ox�R�L�Tw�ŪP�p~pec�@���)�����<�	���:q��yW��3=�\���l��?:�MS��6S��6-��-�M<�|�	��M��'B<a�#g����03$��&G~$'vֈ��Oɟ|j|�Z�4��ܟdX�*O�A5�@˰�p��#`�ן0�I�q�J0f��zy�$o��X��������Oz�# N�9KjUb��]5;F��/�O�ʓ�?y&_�ě޴�r�xB,B�(Y ���,ߓ��J��9�yb�'���Q,	!�����X�h��7&�B.C���t �F����ĨrVr��n�ܟ��	��\�I��4D���'��p��@2s�x�&�T�Z²@���'��6m��`�d�O(m�}�ӼK�\�Ta��MR/g��R�eI�<I��i��7����A8҉�ݦ��'�<iE��?���FP8�:bR�UKB�kT,"$�'N�Iɟ �I�D������
n���8D
�0œ� �	W4T��'N�6-[.�J�d�OR��!��9d��hW��\����6!��1�O�$�O��$�b>}����r��Ձ�.Q+�]�6��!z��+��3?�&-]3K���'�����Р{Er��f_%$=؀�*��4�L���O~���OZ�4�>�.�VMW�l�o�p{2@�F�gT��D0�y��b����ɨO��d�O��oڐo��щƯyZ�-��� ���	������'�F,�v��?I�}2�;5��9Bǉ�R9�	��A�B��?Q���?���?�����OV"JC�(Ht�`Lq�S�'���'��7m����'�60�$/
�CG�<S.Lba�0LB�&����4'���OX.Y���iY��
^@$@�&&P�Ub�`M¶g��x!�FǑhe�%L�	Qy�O���'���:~��m�:+�|�hT�[����'���<�M����$�O~˧B)�Y��	�48-�R��]H���?��S�l�I���'��K|P�k� ��萰i�W�����G?G̦���JI��4�>9�� M&�OB� ��)E�*��4n) "�OR���O��O1��ʓsf�vJ���)�'#��5b�1?�pI�T���4��'/�˓�M�����)2��p5`Ns�|��!�;���ef���K�At�"�,3>����b�O#\T�w!޾{ Xѡ�C�1���A�'�	ϟ��Iş��ş���f�� Eצ�Q��(�Lԋ� �dO�6��6L��OF��!�9O`9lz�aq!i[�B"	��N�/+6L��d�����Ş7�ڴ�y�@��L��X�D_*|iC�Ї�y�@ț%_���I5D��'Z�i>Q��e�~�SW �c�9�æN�X�>��I��$��ğȗ'�H7-�,�"���O����z��L�Ң��|n�Zш �& �lR�O:���O~�&����.+o�(����K(/�Xg�&?�ס�\|�� .�P̧W~���Đ�?Q��ȯM��9	G�?z��Q��MK��?���?���?��9�0T�F��XG��ܬ*���&��OvTlZ"���'�67-&�i�ը��D޸��١EY� �|���I֟������m�B~ZwN	�p�O{�d�T��'��Eh�!�1!��d�t�D�	qy�'\��'�R�'
�%N8B�z�A�+�(E4��Q�H�^�ɾ�M��D��?����?�M~��L�j�c�:���`s�9�%]�����'�b>%�e��:HN(��� m��#�T�p�� �py2��"~1TA�	(��'4�	��e����$k��y�K9l�\�����H�	̟��i>U�'v�7�ΎJ�v�$�	r6|���M�*+�d��eeV`�f���ڦY�?�EV�HݴId���d�R�ƎW�s5���X�Q�h;CGQ���7M(?ᣭ�^���	=��߱p�$�
��5F(dzdhZ�Ol����ퟀ�����ڟ���v�W0�R���;�����ˋ��?Q��?�Q�i�(ؚO�R�p�`�O����W9a�q�g㗻b �uĈX�����mz>%��$
��'M�,�q�'��eR�!}x��"��KV�}�	,,X�'S�i>���ğ�	�x� d���M�I�.1;��c=�Iҟ�'@7�_u���O��d�|�&�K.p]�r�&a�r0��.H[~�,�>���?1�xʟ<�yS�"�@�� X	
�2�����Ud�0�o�y{�i>�r�'�� '�T�F�B��A	��
5 ?|Q��k����П���˟b>�'�*7�
5eB�����(^n�B+�(q�0�AF�<!źi@�Ov��'���)e6�)�AL�`�P%
A�3�BAs����eӪ��f�y F��π ~p;�H�$L�@䃕.��"��5OR��?!���?)��?����I���YP�K4u��@�'KuNX�m
t�hd��ܟP��[�s�����w�(�<d�%	�R�0`qP)ّ�?�����Ş�z��4�y���2��vM̉0�!��K��y.�7j����� +��'���� ���j\��Hso�*�(@��	~�:H�	ş����ܕ'RN6�ľ9~���O>��X+4 0�8��^
G�U��m����+�Op���O��O٪/ӗ!c�5���I�&�ra��PkB���)������s�S�(�R����W �8��IV�ȓP�Y�������IןxG��w��S�"R07:Zec�G�C�9B'�'f�7M
 )-��(���4��С��K7B��	�ǃ�q��� =O��d�O8�d�H6�7?��\ޡ��'˺�ʑ� p����/l���U�"�Ļ<���?����?a��?)��;+�`�d(_[!�\��)�;����+�ǒߟ��֟x&?��+0�y� �"�^�K���3�r�p�OfmZ5�MCR�x��D���p�X$� AH	+@-��X46cld���7Z�I9bK�����'	�D$���'w�=�WC��G����C$4ڔ��';��'cb��DQ��8�4G�Ha���k���׬Ҫ�bP'��;�Ԭ���4Û6��^syB�'�F�~��q��EvB8����V"K�|QJ�^���6�&?�EiN�t���)�����stk߶Co0*���G�\�% ��<1���?!���?!��?y���aš�%B C��2X�W�X_��'>��jӊ	 �;�8���-%� x �N~A!&���'���t������?���|�7�U:�M��O<�cg�}� ���h׳z�<Q��R>�,�������O*ʓ�?���?)�l�RѪ�j��/oҖ/x_,	��
�����	YyB�bӌ�Q+�<���IJ�&]�Mǻ�B]�C�?n��I�����Ot�$2��?5*F�P8RZI�g	ɟ/���֦Σb9�gD\�z�~ܔ����^ПX��|b����=��F80�C�Ծ8���'iR�'���TW��R�4> ��P��$���BR
V�1���A���?���m�����Hi}��'N�S���c" #f�')"`���'��6M''j6�$?��O�;��	2��fI�~����B#n- H鑭��y[�������������ß�O�.� V%�2M`�(�٬�xٳ,{�zp+W&�O����O �?�y������ȠPc��3��vCp��0A��?	����ŞS��ڴ�yc�;�&��g��;^ɀ���D݉�y"k�}ڡ�ɝl�'�	����	.aGp��Ƀ
6�90��A��d�	ȟ,�	ş�'f66m�+�,���O*�$&l� ���&LȤVE=�㟼�)O��ds�D$��꒦�Y.�(�,�Y�hy%�'?�Q�J>x��d`��Z���'v���DZ�?q�fN.��kC'Z ��֋�?���?���?y����O�}�f��L��څO�nh�Ը�K�O�umڹ:����	ן�ܴ���y��� n�s�n Anp�?�y��v�inڐ�M�r.�2�M��O��0��X����E�-4I6
Z��Q��%�29�̒O˓�?��?����?���>��B� �����FF4U�*O��n�0.��8�	ן���I�Sן8��*��V�\]a׋�G3��kq*S����Z���q�4z/���O�t�J�G_g��d+�(s��e�%���3%�Aɕ[���7L��R%�|�	_yB ��tp(��MB�c�ME��$C��'��'�O6剹�Mkc�?	qB�)ErM����Tۀ͂��Y�?	��i��O��'	�'"�$;��e)֣�V��M�EE��j��1�i���!�)���OS��%?u�]'2����n9�n�H�S	,���I̟���ğ��I���	v�'P3��t��`��9�̓�o7` ���?a��`��6� �剗�M3N>qУ_)�H��Z*_ܴ��'��;���?���|jDHT��M��O��T)T2�H��+j���bSE� k����c�O���L>�-O8���O����O�X ABFWd�O �S�
�	�/�O�D�<b�iI���'�'0��'�ӖM���|��E����m{���OT�'[�6m�榉`O<�Oq�U� ��Z�%��%\_�D4�&��	�d�뚡��4�2����D%��OʠG�6�B�+��_
1�d���k�O����O���O1��˓���̢qyP#\�t�ٳ��
�
�"�x��'4b�x�T�$@�O"AnZ�m9��B�"��6�����%/����4_��v�Z�v���R4+7���wy�I�!p��a�� KDu�ЎU��yRW�(����@��۟ �Iԟ̗O�vݛ���2&@�;!h��u��z&�~�����d�O �$�Ol�?)8������/'	�Ѣ2���a�ʄc�h��?q�.����O*m��i_��3�}Ĵ%8�J�T�D�$��<YFP�X���dN�����4����*d$��*tH��ˁ�D�::���O��$�O��G�&�Q�$R�'��f�!R
��# 9�ysF�S�=h�OvA�'���i;�O��0�ݕ( ���%�0	z���`��f���OF� x�ԟ�YCL̝.j�d��O�|H��'LΟ��	��0����D��w�D�.�9w��k��,H 5�'�>6-�w��$�Of�n�i�Ӽ�P��U\،�T	_+�H��A�<Yֵi�(7��妵j�*N�}�'P.���h��?C� B�P��}IB|�6�˥+-�`��B-���<Y���?!��?Q���?�Pc��u���\,���g�>x�'��6MU>)�˓�?�L~���!4xƎB�W��U!E�
�|��S���ܴp�v�0���4[��k `����"U�_¤u�e�>w�˓V�JK��OܑL>a.O�X�ÊY/2Ά���@ŮY�Tt����O����O ���O�)�<1R�i�����'W����lVb�����N��t�T�']z7m1�������Ov6����*�([�(�l�)�h�iT�x!
�t� 1mZp~�>��<�Sp�'ڿs@�E�$*������}�$s�K�<A���?����?i��?���)ۼE���y#i0�
�����,���'�bji����%�<iP�i��'�8t���3b�(��
W�\�0�#�$��{��|Z�ɜ��M��O�q8���]Zm��ݗ�h��)Ɖ.^�����ؓO���|����?��7��)Q�g������qI��R��?a/OJl����%������Ix�$�P�w�Tqy ���;g�Ѳ�Ρ����V}��'�k5�?9�6?k�i�OC`��8P�^#k9Tc	Wp����|"���O���K>���i@F��qH_�p��v��?I��?����?�|:,Otxl��F.B�j�+3q"�s��J�E�XK���8���MK��Ͻ>��
f&�1�	�Y��W�j�������G�f��6����$�ϩT���~�w֩1��|طn�51\�S�hC�<1+O����O��d�O����O��'�p�{-�R\�O
;Sz�M�C�i�jI��'���'5��y��n��� �*�� b��Ђ!ԈD�1�����H�4{���O��A��i$��#`iA���;]�bJ�eF!>�d�i�����s\d�O���|J�F�t�`�IH�.�Ȉ�V!�Q�@1���?!���?�,O�Uo=0F������I�g�J!&�	l�|�ʡEȄw��	�?a^���	���I<	�N�8�c�-��YRi~ǌ(J�R�Т֩�O�V�	�i��ڋ'��0S%U�Nu9@g�?h��'l��'MB�sޡs��ݫL6዆&2����W����4H|�a���?��i��O��K�x� U�)8D���i�F�2���O����Ol�Gg�"�Ӻ��Ƙ.��g��a��gJZ�W���ե̖jS�O�ʓ�?���?����?)���2�p�T�Q���0��;^D�)O�)o��e����	̟�Ij�'qu����
�%��Y�%��B?�	�W�ؐ�4N��f�'���,�p ���rN��.Q7�!��Z�R�ʓFe�!� �O@q`H>/O�-��g��H�lś��אg�����O���O&��O�	�<�ְi(�ۅ�'�܅���f�h���B���4��'`7�>�� �����5[۴u��̅�@tuJ�Œ�L�P�0��"U��P�4��D@�z�:1K��_�����N�	h:�������#�a��~b�'���'�R�'h2��o��Q��04�� 1@ �M���d�O��Ąæe���w>i����M+I>��(��m���K��H���-=��'�67��˦瓫/��n�q~��nI 	�����z��ژ5�U%�џ�Ё�|rU�d�	�L��ޟ�r���D,Q�ƅ�x��(�c���X�	Zy�fy��d��O��D�O^ʧ�^CfC��f�<��Q:#��D�'RJ��?)�4e4ɧ�)�9�T���R�g�X�x����)m�a���!\^�P�ʼ<�'l�~�䙫��}��"E�H�y>�b��Ԟq�(|���?���?)�S�'��򦹱�H�"�~���V�_H i26!�5I��%��ٟ��4��'�~�K���A��?��
bC�QB.�A�D-_�7-�ݦ��E��˦}�'����?�AsW�X��	I  ]����p�T�k��'���'m��'���'|�+�vTQ���4L;] @��S�ġ3۴Z' P���?Q���䧊?����y���G�(媔��7؈�y��S�^���'�ɧ�O�zH�V�i��dR�>�,i�աGȼ��g�A�󄒖sTlY��y���OR��?)�������I�O���� B`�T���?����?�)O��m�51�j%�'2�-{-<X
�l�>bVp�@�M��'≬>i��?�H>��D@./Ʀ�[7�K�*�5b�!�s~�n��&��5���Þ\P�O��)�I�\�+՟|;H�X�̓%1�D�i�2�y�,�="��@��ھ�X�
.�REu�8����O�����e�?�;a� �t�дAG�,�qG\�����?1ڴu�V�M_����Ĩ�'̊J��	�#�p��uA̖!��� �O�t��m%���'Zџx��mT Ux�$��Ǝo�& �!=?y�iS8�� �'_��'��d���<��p�Ù3/!MS�Ryr�'ϛ�(:���t�J�VP4-F���t���ɬ"�)؅հz��'&)
���'��I'��'J�Xp��<t�h-��KQ���E�'���'���4X�#޴ � �r��W����U�@:D�ѰHK����`��˛F��Vq}�)q������������v�ӓ'A;��Rei��j��xm�@~2J����I�S�:��O��!�0�,�VD�*25�bB��y��'z2�'y��'�2�I��*.��!��K k5���� }s�$�O��d��A��On>!����M�M>Qe$�k���N0����T�UD�'@�7-�ş��Ƅ@|�7�'?qe$�G�? ĩY�KF0,��q��	�|�"��s���?���3�d�<���?����?�EZ�$���"�%
n�jT �7�ZX�����d�Ҧ�@�ޟH��ǟ(�S��M��%�ip���P#h�6���id���I���d�O,�%��O�����#1���g�œ=���L���}�X a0T��S�\?�B��&Uf�����GK>���@�[�I��H������)��yҍ|Ә,�P�
-@D���+Ռ)μ JЏS	J��ʓ=�����L}��'U�AI2Ŋ�P�;%N�>n��.��'��D�e�i��i�KQ@��?��U�D��h�;oB4���������z���'��'���'�'f��=D�h�䐽��]�sH�/;��%��4%���/Od�� ���O^�mzޡK��P̺�H��N%~⪡y��ʟ\��O�)��-oZ�<Q2�%��hÔ�D��J�D��<A"��6G�@�D
,����$�O>�d_�i��X	0.Hp���CߢS޲��O��D�O��?�&cO�8�I����5�� +��9��ʞ�D�p�CTz�	ܟ��O\m<�M���xrC-!�����L8!��ק^���$ߙGp��x,[=B������@��@�l�D��`a�=+�q����=V��$�O��d�OV�d%��S�.DK�(t��D�f>����m���?�&�i*�b��'��+|Ӡ�O�9�*��ł@�[�Uf܌s�B 20O����O��D,Obn6m+?��^�j#�'[,:��%�˨G�NU���%x�H���*�D�<���?���?����?���ȕM����2��B\��C��[���B��1�Ԭ�ҟ����@%?����g���ɗ ^֜B�A4_�,�
�ODlڹ�M�ƛx��$l�nh �$�FCX���� �*�҄�c�F�t��Iڋ��?�n<�d�<1K��.ѷ-˓���$R��?���?a��?�'��D��I�#	�ПH�3�D�x����
;H�Z��Ukk����4��'n��V���J�O�6T����j#C�d?�!
D� KNQy�vӊ�I�L-��N���ȐN~��Fݴ�B+�"`��P�� & ��?���?���?i����O�f|C,[�0����I��C2�'��'�7�(pI���M�L>�ը#{)��MO�,��!r�I^]��'�l7͑��S�+$,<l�y~«�Fy0ɗ�<l�ԵQ@f�A7���<�q�|rV���	֟��Iȟ�p�Q< �,���:�j��ß��	`y�ohӨ���h�O���Ov�'v)^=4j�U���E$\�t-�'4�'��j�OBO��W����i��@�ִ�a�˄s"�xe�O�3r��
��Cyy�O�����1��'�z�Rq�*Qt #k�� ��p��'x��'����O�剭�M;S�Z&>."��m9W_�ݰ����`����?��i~�OF}�'o�*�;qgr�z5�A�g�i��I��R�'�.{t�6����W�8��剏3��u"�s�wB� �N�	fy��'�B�'���'p�[>]b����[��I�۝{^�d{��C4�M�5EP��?����?�L~�#���w��d�4 :R�ر�v��C��'���=��)�<<|6�r��c4���)�԰'��#�.�vh�ěB�	zE��a�IHy�O�Bl��^"9�"�����T�g�!���'���'��I��M�rF�?����?��m�jq ��� D�ˆ��O\��'��'�O���J� @���f"��g�<�#W���Qu��?�΁{�N,�>�BN�ٟ��!&��j�Us���m	�I���I��|F�D�'�l����h\ɳ��YG�$%�Q�' �7�RS���8�f�4���H6�c�U��Uf� �'��<�ѽi|�7M�٦��E����'��x@�$��?�G�*BQ��k�� ��lCSg�S~�'��i>��I����I՟P�	� ���kW��z6�Ջ��K?6pD�'9t7�VT^����O��d/���O�T�pB�rd��흯NC��N&g[�Ɵ��	W�)�iHY��CQt�a�mZ�d���ZW"^�7K�˓k����V��O�,M>�.O������|��xb̒.D��)#W`�O����Ox���O�I�<�G�i^�#��'{йz1h���dz��4t'p���'z6�=�	���ě�����M���,R��)��I�Ą|�c�ɧ*i�H*ٴ�����b��4��'p@�����[��U�ȃ:L��e��k�����Op��Oj�$�O\�D!��� =��`�'��D���A���� ��4�Ms���|Z��MA�v�|bK�����/�3sx-��&Q����Oz�q��)6v��6"?�%�?MvVdTTbU�e)��2M0�
T��OJ�yL>!,O���O���O6�W`W�b�lz�$b�n�׊ß���Fy£w�(�E �O2���O�ʧn3�����N�E<�8���$����'d��?��m;����P`�P�҆V�t#J��蚇[E�TJZ�In3G���Ӱ3���
i�	�E
z��N�*��Lі,N �����՟��ןX�)�Ry�xӾ���fC�H�<�'jķvYP�a�⁕&l0�Xћ����w}��'!D�+a�'3��Hs�(��p���i�'�7��q�6�2?��ȘKF��)=�T��!T�Se8��L�U�
�yrU���I����ݟ�	�ܖOT��R��{aD)s����P��2��|�ʡ�d��O����O4���č��ݡn:!�����E�q�0�	�%�b>��e�⦽�S�? �ih�C�*��!��9�$Y�6OP��CmO��?�S�)�$�<y���?�
�$XRy�'B˹kJ�ygې�?���?1����ċŦ	0��៸������E�	����'́Ih����)KR��?��I�M��i"Ox�`j
�i����U�_oh��T��TQ�ʝe����wI�}�d�"IJ�H����0H� Z�,G':J�Sj�����I�������G�d�'�"�"��+�L���𩅢�2��+�l��L���'>7�.�i��dIH��|a�'ƢBL���a������"�4n�@M0ܴ��!l����LB��3����<���atȚ�u�����,���<ͧ�?����?1���?��¥ ��d���r"�8y�C���P�x����	ß'?�	#&N�� M�mȚ)г�"nM�O��D�O�O1���1��I`|�8)e�C6`�S��ό�Q��<��bG�8�t������1x� �x�h��
c$�u�_�d���OR���O��4��%�FK�w��E�.�bls5�>-�i � �tY�gӞ㟼��O����O�Ll�B��QY�M�3MY6Hy@�S��Wc^����' @$0����?Q�}��;|S��`T"y�
��! ޴$�����?����?a��?)���O�t\�R&�H� z��[�\�Z�s��'dR�'l&7-�y�S��M{K>apĜs�,AR��8fy����*5�'�t6�[����¨>�@6-!?Ap՜F@>\9 �&6�1Y'��cֈD�T�O�`*I>�,OH���O���O����E�i=���c�Y2���b�O,�D�<yҺiq�"�'mr�'�sU�'��.|�6��d`Ƞ]|�d �OZT�'<�6-���'���H�ET'(���"�(B܂��������F����4�D�;��x~�O:��U�W	y[�<�M ��� �O4�D�O���O1�Fʓmk�FMχmB���&>��a��Q�x�|y���'mr!}��� :�O�n���،I��\$|(�1kY�L¤9�ش0+��oʕw�ƛ��Y!�ܣ}/�dk�Zy���h�a���>,���sF�"�y�^���ʟd��蟬�I��O�R��%C-ngR�!c͚:" �x1�lӾu�խ�O����Oܓ����S٦�]�mŞ�����2<hV��b�łq~�t��4F���L/��7-b�0$ڵ	�8��$�zt:�`�&o�L���S�aH�CZ��oy��'���?����	��,Hh��� <��'���'���MGf��?���?���ٮ\l��(t,��o�t�ˆ�ۯ��'FL�m�V�xӺq'�����c�r1K�JiSP�#�<?A��-����CD�$��'#���䕤�?���ܨv���U'�)2(�7�� �?���?Y���?Q��)�ON��]7�6(�$I�*�Z�bQg�OTMn�G�&��	��Zݴ���y���!U��@q� ';'�8ʁ*�'�yBDj�.lZ	�MkV�[5�M��OBࡐÖ���*�Ӳ��O-/�P:#�^�%�<��|_�,���l�I����ޟDk�K_;��!��LQ������	{y2Ba�z�����O����OΒ���<
�U�޾2b`8�g�ˈO��)�'t�7��q	I<�|C��z̚�d�J@fhI����V�>X"�I6����b����&�F�Of�B!�H�L�X�B	i�GQ�*ޞE����?���?!��|
*O��l9� �Ʌ 洸���J/P,��� E�Y�I/�M��"�>	v�i 7����y��o��S������q]�TxDN��a9V,lZN~�1@����'��O\w'�<G<�ÑD�9:��S"��y"�'z��'R�'1��I�?'�|s���rNv�1c�&r�`˓�?ѳ�i���+�OZ��f���O�8c�gշQH@�s&3���Э	s�Iןoz>�r��]�'K�Y�Ce��4��|YU��?��"��V�`H�����U��'J��럈�I����	lþD�#�!p�$�G,�.s������Ė'�P7-a^����O��D�|Z'-L�a��k-��4�^��	�o~"�>��i��7-�n�)��l��n�A�U#n�8���̲L�w�LX�V	a(O�	�?q%�(�d��e��ha�/�6 9F�8�	yT��d�O��d�O���ɷ<�Ŷi[����� ,H`�� 4e2C΋k���'�f6-#�ɞ��d�O�1&�F;e@�BCb��#<�å��On�$7.6m)?�;eh�z��&<z�R��� �8�:� �I�6K~L���$�O�D�O����O>��|�tp��q��̈����7�A3l���N�2�'�"���'i�6=�0�*�n��nx�@�j�#����O��d)�󉏑i�07�w�D"u�� �>��CK^�vX�7mv� �1�<=���UX��}y�'�RHk Ȑ�l��mh����!	���'�r�'k�I��M�tD�6�?i���?�@�Z�fr�����/<X(����'��듖?��8Y�'���k7���>�\D����,9<Uq�O�XR)M^yҒ�醞�?����O�=c�	ð�\�(��@ Hjp(J�"O,А���.kL�Q5i�:l�̹FC�OZ�oڇS�$%��џ$�ٴ���y���g�湠U�^*;�l���@��y2�X�*f�i�h6MX�^<�77?�F�͖	yp�)�3)�l)�)�>R��$��㘓O���H>�+O0�?yf�O\.)�G��37U\I2�`~�Kw�Xz5-�O\�D�O��?�zs䖻U������W���� ������̦�xݴ���O9�B� �A�2A߃�(��P,p�j���i	�,d`˓n� BѮ�O���O>Y)O��*�jJ	!t�%3�ꂿ'r�����'Q`7-�������4ڜ��2���"�qB敥5�~���ۦ��?V�D��۟��I�<[�1�G��2 3RT��cL�}ߖ��R'Sզ�'�Zk�?��%��TꀉT~�z��;d�j!y4M��ar�%x$�ߦy�f��V,�Q��Y���Y�YV��:&�5x����O��uZ��8��԰UmC���B 1���_)\/dL�e�8(-,�uCV�s�!�D #�ͭ��B΅ �>��4�F.x��`�eV ]�dx��j�-^_2T"6
	+@��r�̀
�NlB��A l�����	S*q��q�(�&������<LΔ iFH��o�z�)�<�Dpc���x���[W*�:��iac�2X�Ā)�J[�C�Ψ!�@����q�R^@�us�۶�Mc��?���^��t�����Of�I�@��С�vm�}XSF�o�c�x�&D;��ҟ����QS��2 g`���6a[�`�b�
�MK��Jؑ�x��'�"�|Zc�4��ː |+
�I��)��O��B�{��'�b�'�u=�QJ�� ���T�V�A@\�RfM#���?9������DL:an�(�7[
 ����Ԥ=s�?��'���'y�P��3BN!��t�N�w�LQP�lO��ԧ�>��$�Op��2��<���a}"(�(.�К��+Ae}��M����O:�d�O��
�l91��t��J``Q��L��xz����.чR�6�OؓO�ʓ7�T)�?QcZ�䥘�����)kӤ���O���t�q4��$�'|�d�p�M�� �=`��9#  ����Or˓Io�Gx�����,۔7�5(�!*Az��i�ɮ�jLٴM;�S��ӆ����-����g`�����/V���U��p��p��|&��#��,���1%TX�ԅAFnӂ�Ñ����q���I�?Y@O<�� on�q��(��#n+�$�� �iV�����Ο�pQ��k����EѨ]N̔2��
�M3���?9��r��5ןx"�'e"�O�,q�(4YMXup�d�	&KFTcS���: �1O^�D�O~��#b�$�� 
.�E*@l�T�Ul�՟��d� ��',�|Zc��ic��}b6����)y�۬ON�J��O$�d�O��9��,B��@�	�I*���h�k�F�"P�''��'��'&�I�c�4ڢ "~0�k�0�`L��"�	ß��	���'�1���j>�9�*Ю\�m��� (���>q���?AH>y(O~��'Q� �"O�\+b	����1����7)�>����?q��?��AL |���?��'����Ց`n�u(�nC�TW{ߴ�?�J>��?�e�9q.�'�x���i��E(��\�D���If���$�O6�d�O�<cB�O��ĳ<y�'�lu����?1 ��Q�ϟ�: �C�x��'� �*l�y���a;Po��]@���UG��%�iB�'w
h���'�2P���SzyZc-�����OP2�:��,�ƽ�ߴ�?�+O�����)�ݦg_6d:"�4���2$�Y��CT"L��'C�	�?	�'G�I�/F�FO�f@"�	�n�����O`����)��`�BQ"r\�����D/.� ����\��M����?��@�Μˁ[���'��O���a���6��$�}zm���iS�'X��#!�	�Od��Or؉"��N��P��"%H`��%�֦���;AVĺ�O�ʓ�?�L>�1[��	��b71��"��";W�Q�'�̜Aї|�'���'��	 ���+̍?��,1#�iz�t�`&���ĩ<������?��y�Ĥ��d.zf�%��J��|��T�?�,OH���O��$�<!.ҧ/�	̏+��eZ'P�,+�-H3@���&U�`��R��d�I:Wbx�� .�ͣPJX4�d�@���3Z�.��'���'�bY��8ɔ��I�O���i &t\٣#�PC"�J'�ܦ	��I�	���! @��=I$��<tYft�be\6Ț�Dʎ��	ڟ��'� ��D�~2��?1�'n����j����"C [o>آuZ�P��ş��I	
�@����?����>*S��sӬ��\q�|�pr�ʓ����%�i���'R��Or����᪂3w20dL�pZ����I���Q�	��dA'^����O�,,��H�b���6A��A�ߴ%}�(!t�iTB�'���OL�듸�D�֐l jBv�h�´H�?Xj�lZ�a�4Q�?Y��T�'~6ٱ �'9���/B��(iB`aӸ���O��$��YM�!�'8�	ޟ��QU�\�5Ŋ�U��@���Q�l�,�>�LM��䓪?���?�s��j�@S�B��lR�퓬mP�V�'�Ku��>�.O2��:�����$^�	,�A�)��ԅ�>i�����?	��?/O���1��?������S5m)�B�g�J��'��I�$�(�	⟌�Wj�*�D�Z�Љ� W,j�x=1�h�Ox��?Y��?�-O�Lj�
�|�V~�0�!Wb:�LI�d���Ŗ'
R�|��'�DR��$�W��qxq���t>����(ʺi��I˟H����H�'g��'�U�K�p���lD^�A�  \'��m���'��'՞$��')�'W�6�H�_+L�L�� ���@mZҟd��iy`2j�`����k�WM�E#I�C.��J5��f>�'��3e����C��s� .�� �[�N��cf��?X�� �i剡*����4R���8����D2-,� ��(Rh&,3QB�(|>�VV�p�S�T�I|:M~n�Y�h��5��g����%ć[L6^>?�����O���k��i�<�O�h�����D*}P�����< ��tӶtk�i�p�1O?)�s%L�7���Y�ں	o��Y3e��M�����Tc�)zI� �s��;.(���`B!XH�Ԯ�ǘ'�<��'A0������p�Ud*�F� ��-�"oE�Yo��<	uMCy�ͺ~����
�Nb�Ec'�X�g�L�rύ�rWh�j��ړj��?*O��D� �f���#�nDq�*ðZ��)�2N�<i��?y���'��"��U1
]�e�C~9+��.X,����3=(���?I���?�,O�Q2���|�¥ܸ;᱒c��\l ��Ԣ_G}R�'�2�|BX�,@��H��8w�I>K0�}ai__��!�Š����O���O˓?�������}B���L��*�5J�� 6�OV�O(˓K\T�����7U_ҙ�F�[�]��9�g�D��6-�O�˓�?I6��*��)�O���kܹe9`	�H�.���;�!�>�']b�'���E�ؓޘ���	�J�ђᓪ ��YP�F�FY�,���0�MC^?a���?�(�O�`6AOl|$d	�
�
#���D�i���u�dP�I,��'��禁��0|L�M���Ӧ)���!��Fɗ�|�7m�OP�$�O8���w�i>qk�E5<�B��B"�"t�������M{�)
��?9�����:����Ã� �Xj���j�pTcD���M����?��'A4��(O�e�d�����B�	�c�r8慯Z��d�<A�c8%S�O�"�'���;���[�m��K^���c���7�O��a��_�i>Y�	��'���S��,q�:���0
�n��r�w��d�	C��d$�$�OT�D�<Ab&�'HkzY�&KC&s�n%*��C~}�xb�'���'���ɟ�I���(�J�\I���(�'xl(�b�g ǟ��'�r�'5�R��p�����$�;�p�b`.� ^S
�����)�M3/O��ļ<9��?�f��q�}���[>i ��1(Z.lΕ�a�i���'"�'>�th��l�$җ~ǆ(Sh<|�����ն!�No�ȟ��'�b�'#�C��'�U:�i�#�ڍȗ*�)�����4�?Q����}!��i���'�b�O�NU���N�]Cy�U�[3H
PL�>��?I��u�'f�qs� ����³M������Ŧ%�'��5#0�|�>�$�O��$韖�קuW��
嬄1�nW�N�l���<�MS��?ye�\�'*q�D�0�8?�&JF�%��8yP�i��dרwӢ���O�����'�I�9��`P��A����`��eְ,rڴ�t���?i,O6�?��	�(��%$��0c�J>XB\�Kݴ�?����?	�����ey�'�$�r踨Ck��T����ڪ|ÛƓ|RD��yʟD�d�OV�D�5���e�L`ҹ��ʗ�+F�Ilޟ,��,L���d�<Q���D�OklA��4���<��e4��& �ɭX���4��ɟ���ʟ�'�$Ű�V�$�irÇ�.~��!�&�����O~ʓ�?�(O|���O���[���1��Zְ�q͘�4�l)57O���?���?�/O�����K�|
�+�Z��(L*9��#I�Rʛ&X�L�	Ay2�'Y"�'�@Iۘ'�H����)��G]�4���'oy�B��Or���O�˓H�x���^?��i��L�[�=9�� "�z�Su�B���<1���?�y����?��g�����V���Y3t`�4�`1��i��'�剎�������O��IY�V4`���օ4U���v����:��'�B�'��N���yR�'F�GR��^���a��6E� =a��@�՗'��q{�iӨ���O��$䟌=էu��׃X4�� /�a���9r4�Ms��?y��Bn~�P���}ōM�
Ѱ��oY���A�禽����M����?�����FS��'V��#P"��B&�<o�v�Rdʚ*pQ7�c��$�<����Oh&!7D
A��/9Q�D�@�'Q��6��O����O��S6J�P}�_���IZ?��Ƽ��dQG�̇aVb�s�IK̦���Pyb��8�yʟ��$�O�$�<��Q �/ƈ����`�`�xl����� ��d�<A���D�Ok�R�v�<���;XY2�{0���Q��0 ��ß��	����	y��'U��3�AJ�X�l��K�B�@��&ªs�����O���?1���?Ye�#q!\d��D��dV�C�)|��\Γ�?A��?����?�/O�� d
��|re�!^�����W���$��Ϧ}�'eRT�x�	����I�oe��ICeP]Y��>��(!A������՟X�	�����{yBJ�<7�N�'�~��0:+�cЬ�<IZ]; eN��M������O���O�y�T1O��'�kԲ��b"3���Ǎ�M{��?I,O�����c��'���O�A��nL�D"$�c�H�Mr������>���?����Y�<!����D�?U�5�ڸ]fY���J*1z� y��8CJ�hg�i��'\��O*�Ӻ�Ԧ�= `���"��@�2���EAǦ��I�����~���ϟ0�	a�'j���ǧ��"XDb�@T&ߠel�!��T	ڴ�?Q���?���VB��hy⃆�o#b����;�Dq(kU�&6m��4�$��Οĉ� zAH�l�|$�s�I�  |aſi��'|�·/T�����O���6[ �SCnO��j�{��͐H�6m�O����ORTC�0O��蟤�IƟh���G�o�;�i �W���'� ��M�� 	�ÚxB�'e�|Zcnr�3�IĊ�
E�cs�M��O�`N�<))O��D�O���<��%cX�����&
A��c�D��0��!��O^�O��$�O�]��)ثv�:�)D��2zʦ������<���?IO~��KQ���)��d&bE��B�옊*�g��'��|��'�"b\�y�, 3|���T!N�{�2m���݆up8��?����?�+O:��`o�f�8C�U��i���D'B�qE�D8�4�?I>����?��!��<�I�,��2PMl�[3�޶FAhy�Cm�0�D�ODʓ^u�����'U���]�M( Ă$T����=?�O���O��@�*�OP�O|�SA=��X$%�|���ը)�6��<�jɬa����~��������u�!.�	XF��#lr`4���t���D�O|�	Gi�Op�O*�>� K�,r���R�\�!�N����~��eZ٦-�	�8���?�0K<Y�[Z|h n,l'��W�l��xsv�i�nM9�'��'���S�?E�!W#ƒ��dFv+��o�������HyCNE���?���~2��c��[Q�NG ݺ����'����y��'���'��%��+A�ya@��
��|ZΉ���z�p�$�/Y�,�>A�����a,񰴑p�>V�ڜ(A��q}RbE�/��V��������[y�-¯ r�:����I߼���ÞR���O7�D�O�d=�d�O��:�	�h�rt"�1D�P`��a2OJ��?����?!-OȠ�Ta�|���"F���ڐ =���\}b�'�"�|r�'�R���y"M�5F�y��O���P�����9����?���?�-O8<���J⓼d^�Iud�>=#�Ya$`���Q�M3����?9��bHۍ{R�I2}����ԢT5@�ҥ�׏E��MK���?�.O���$D~�S˟��S6}>R�
��\6|X��g5vW�K<����?qQj�<1J>q�O*8A���<W޹"E��	k��`�ش��I0a��Uo������O��)�u~B�עp�f�YQ�v|%�֏G��MS���?!��9�?�M>�/�p��t��9[�m��4>����K�I�p7�[(H
( o���	�����'��Y+U�W�
��WW9����iv�V� 6O�OH�?��Ɇ^fE3�_q�}yi�`t�$xڴ�?����?�g�pL�����>9�e��B��`��* xq�M���?�����'/��'*<�`�E�qh�qA����brӺ�$G�:5��&��^�'�� F'�z<!�F�5�h9L<������O����<��C���'�Y�$�~��Z�KP5q3n�:�?A���?Y���?�O>Q��~B�F�b�;�@�/�|Z� �M���s~2�'��'��ɝQo��O=��V��(��y���Ҳ
��pcO<����䓑?�{��P�b���;�!!�������O����O�ʓy�x��W���!�),��#��]9#t���+E�,7��O^�O���O݁1�$WIp�v�)K�ԠRH�E_���'�rY���⩋��'�?��'_I�	��U?Y��#�)��rz�ɠ�xR�'����O4��"ऍ��)Y�z7����Æ�]Ubd�I��0���D%?㞄Y'�*C�� ��[vX��9D��sц�Z�WQ�,����U�D�Q��TpV%hb_� <�x���cC"Š&�W�8��������I�4`�Ƃ֒ld�H2�)]'=񸱂��-hP��h��?e��%rS,�Ќ"F�݄@< (�g,X-)����#tc�����i�VD������3�ٰZS(�Ie�
 ���rA�=���'��'��֝��x�ɍiX�Q����=��,i�y\I��ǋ*
�����9b���;���?� ���֌b7���<3th�"$��(`��Y)6��:�uB@e�2R?4�ٟ�hDy"���Z܀��]�	�)�	��~���?���hOP˓:� g�#W�D=A�F�
[����#[^t@A;GE����o�:���E�)�,O2��U�����!��U#�J�Ȁ�8X�L���Mݟ0��ڟ���1^ܐ�	��,�'p򤸚�ǉA?�}qC��Xj���+��f�d)r˘ �L(�ϓN���P��\3���݈��"��j�"5��\��X`�M�rx�:5o�O���84px��(<5^���n����=ъ��M�O�|������d,r&I�]�!�đ�o�t{RL��TOZ��@�w���H}B[�蓁H%���O2�'F�\5i�ٹ!���	� ?g>�-`�K�?����?��ԟr3l����+�|$x����i�t�~�꣬�1O�	�P��}�Q�x�dHCŠ	�"�&>�&>��!NJ���R  ˷y8�`��>ʓU;���(����_�O����X�O�����<���;<���F%g�z�І	�t��	$�����~��a[����SR�����<u��X��П��O$6����?1�a�hm�"�a��|� M�8�ȓvo۫JG� k���9������I8��O� $:��ӻH\H�u�W�0;Z��p�@6�ڂ&=N��i e�#�֔���,<q�w�Q:G�1�J	�_J1����f��s��'�Җ�����OL���$eB̸���©D��)��"OX4Rg^7-/���r���`�Hu�����HO�ӷZ?��Ca`� \�DۥC�k^(8�����k�%�S�0������I��L�Yw�r�'s2�q�J<=�ȑ�nC���5
�'<9xT��,C}2��׊=O����nK�`yxc�ĽDn����O¹
3.N #I"��be}X��8&�8� �����(0��Oȥu�'=�Yy�'�Qq8Q	�h�kׂ��y2������@v6��gZbr���@.�S��V�����:X���(]�]P�(F�'?&9��$ѓzA2�'���'�d���'��'>���V�'L��^+X[��jr)�*&,��0U.L��p>�e%� ��Y�䬚02���+�����-�<E�2��$�P���'���bB4_ ]#7�Q;MF��pp��B�D�<����?�I>�O��h��O/�&`!��Dʆ�
�'К��T�8[��C�O�C��q)�'�7�W����'��M�5i�x�D�O�˧ ��!0���V*x �w�ϕ`z������?��?���Ǖnx���|]>sGS�$��hqU���P�:y�v%�B��ZDF[�>"|jc�СQ���t�1�D�G�' �p���P��Lp����|�r�Q';r���(�6m��L��̚��?A���9O��*"�P)F�6����l��!��.-|O� oZ��M[��,�`}��`�-y��=����:�luϓO2*\B7�݃�?�����iݖ����Or�$���G�	7a  {a�h�m�"�Bn�F�&��'���?���\b<��,�:�Y!7�Q+�9�e�*f�ɧ��R�B� b��X�Ov\���+a* 
r�'���'��OL���IG(@Ud�WYd}�4 c9Oh��%�O $�T	��b�R�qaZ2)iٲ��ɞ�HO���V������h����I�Sot���Q	�(R�)����%JQ��B!��+�t�ѡ"�<[��[e��z"�ц�X&�
�*��͑S�ْ+���r�@��fй<x��) 6Z���ȓ��%H���63�}y�X�Z�<�ȓ�a��i��^��Р�) : y��[��H�T6꩙f�Ġ_bd�ȓ~>��7�� �@�9��	�����
�L�R�ȋP!��95/��8H��r��Zc�ߐ4��t�G�.�j�ȓfn�@��!Y�(���t�X��ȓj׼@!�Kߘ"�r�i�`YLF`��,��� �N� q6��P1H�f�����2C֍��+G�g�n�pӄJ����C�F5+A��b�!�҈һJ��ч�9Y�=��$		%�5�ׅF�<Δ�ȓªX��&0�����^5[��ȓ~�b�R�g�/uz��C�A��4��B,��;�O�l x����S�:�lh���8P���R���� ��'�`H�ȓ;�d	3c���;~�DYE�]�XX�نȓ|D��]�W��`q�oj��m�ȓ����\�
���SS���u��4�ȓ�M�� �uvv����x�'/0D������)r�h4�1j�0?�� 0!g*D��� �8 ]��%��RaR�J��&D����L�-]G���e�O��M2g!$D�(�늦y� �����)p�ps��!D�����
[~>�āݎ���5`4D����O���h �Z>pVr3a�0D��:š&LV"�Y`��\�.��@�:D�D�D/C�%�� ��W�� 8D���D�0$|�
Ԧ�5U�$AX �(D����c�*�L���<Hg��!D��%O�XH���q�84+��1�"D��)ЂΑB�|�����\$�a%%?D�� ~dZ�F�0N�&��j߇I@܋"OHH�%��֌��b�S�|a$"O��Q���>rhy��ǐu��˃"O.�$U�6P�:׏�/,$
`"O��
2�G�#b���V!9+�^x2"O����*Lp����%t��}
`"O��P��81��Ǎ@�L �"O̝RD�!���d��<h�8�6"ORh��$�%;L�ꎕCn�ͻ�"O0��74sF�8��CXiv�y"OP�Qt��>�F�+�
��\ �h�"O�zuIH-����^�r�l��"O�L�f� �:�n�s�?�	�"OD����EN�6�pg܂<�q{'"O���Q�,��@��ݷ�r!��"OR�0��
Q���ے�܋w�d92"O��y��\/w�,�0�Z)G!�9�e"O$�0!�� �M�FH%N$�sF"O�B��ÝW��b3m�O�*ԋ��		|AB�,��2~�Z�������59W4B�	�OE8I�"F�U|�(D`\�{�˓�Fѡ"@���S�O"�=;wLE�j��P�fR3["
x��'�0�أ,�%RS����,]�FP*M>��.Y�VpjÓ?2�M��Đ�Mp i��fI�U8E��I�;:�m�t�D�_�"���)�~�"{��W�H�^D���)[��.�y��8揟'�B�E�Ź$��}:���؆5����� ��
�K!�$F�&*�Q1�,�=	�*�	�	�7�ɱ,�4���'�e�)�'SI�<��*E����fJ�n�l��ȓ=f"a��7'���&Q�^�ܸ�<��P�Z�̘��	�~o���!�֓���V��}��B�I' �i���T:9m��c#�]x	�B�IN��q�i &?�L�X�ZG!��$�����D�.$<b�O�!�$��#��lQ������3w!�d�ji��+��,�X�`�o�,Q!�dۜ�z�A����E���^&HI!�ē ��\�e�0X5z9`'/Db�!��yĆ���iڵ- ���4~!�DH>�q[���G�J�1RMط%f!�DM�[$Z�)���>�>ј��&eB!���|HDr�&V#,�h��E�Q�!��L\���p)�)h���g�4�!�:N<�qH�Zoh0�3�Gr!�+I�bdXr�X�n�F!��@.�!�dۚf{�4�P�D�.�j����!�Dן5m<U�@"�L�feX#KS&*�!�D�@�p�Q/�2c|�h�B	�rz!�Ѫg
���B�3uy���G�:(w!����r�F�zs.�w��7F׭	`!��cJ�!���*+�� E�3]!���@��%�I-��t���T�d&!�dH	p\�2�@�*!��1���t!���']��J��N�4�cƒ�Y9!�d�C���".���aTFI�H!�ݼ&�>��&��=S�B�;Pl���!�$�%�*�#�>~^Dˡ��F�!��Ɉ)rdQ3�Y2l�����Y�e�!��&Jв��Ή\j��&��&7�!�d
88遀��0¤@��U��!�d�2�������3QH��"�n)n�!�Ė#D�!ʵ)?��r̓8`h!�Dt�zy:��ˌY3H`81L�vt!�$A �n`���Q�` vJʴNG!�� ��B��7nD��� 	{����"O����J�d�����N$��5"O�lIS�Z�i��'�[�Z�,�"O��rv��+-|Q&'9D���"O"��E��\&\�FEռ@A�`�F"O
�X��)=$f��U�%E:-�"O6i[��-#yh�Z� ��nԠ]��"O����	�YO�)�d/@)��SA"OP9���62��;s��
`�ִ�R"O��b͗1`��8kQ�%�@�'���т]|��
"�Ly�W��m�F����Y}����<���&�����O�u���U<2���)v�F'v�X�t�d	T�����ة��'V ܻ�%,�>	�% �N20z��aH����������c�Ȑ:�ʘ+T'v��f�Ƀ5X��p���G����O�yed9Pq��ԮR[�4�*Dqb���|���aݸ0:��@c"O�d0�*�Bm���d/f�r#�'�:���"�4�^MB�j��~҉�W����b"���f�N|���(�yaH�� !��	ܦ`G)R}�>p�H�o�,�uG 6��S�8��\��)L�/����|�b)M��~冀N��<Z3�]�8��`����0?�a�Uh�u�듃.��v!V�k�f�aA�":3.J�1��A|v|p��$ �#�uI-/Z��sXY�\4D|��1Lp������H��8��UE@k�n<�pFE�6`:�&Q�U���v�'[�}1I�Y�y��߆f��k�'䁛�Q�7*�ljbDA���S�&�Dٙ�'Ͷ��f@��9U� �1Ȗc��q��cd��a� F�+q�%Fⴵ�ட�Z��[.h��˓� ������@���y�g�1�l{f��i��� T�J �p>A�@�j���L܂S�d�QĄ�
��i���,ry:O�Y׮��,:AA�9̈q�L|Γ_�̱�$�!�fX� N˦Z�R$FxR�M���!�gAY>u´̲"	���?�'E1`8�f�c�9Q�턅�,d�/�� 2�3YNYڤ�2Od4S�
��st�&���tA�BVe.pX8C� �,B\��F�{�J?�O\��kI�%�ҭ:SO�7��O� :!�dYI��O�;����F�_f����,�O��1�A@�-l���֟���sRZ�L8���2�.P���ç�߳LGaybX ���G�#����*���"����E�� �]SZp� B��RXx5nL�w@�	7K����1�m�O��J�B�5��� D[�0 �"�$XA��dHZ�aF�����BӒ��'V��Θ�)���ǌ�_T0�C�����Y9��7�z��a��3O�k��&(k���̋�H[9� A_�_�M�6��U@�Y�4�x�i����x'?��R�v�1x��#;�1���1IjaZc���� ��`*\zr
L&MіeS����#���hR2�"(8?1���+t$eM@�)��1z�h���496�B�'������a8�����ȠJ�i��O�B�X��ŦN�Tth1�G�#\*��V`��M�F_���dY#2��sbR:�:���!Nϖ4�O��q�&Y�\x	��-Ռ5 b"�>��K�Y�jA:�L��v��iCE��F,�r�j���b�W,ڪJ+�� �ʈ��6��V&N�����-@.��J�7
Vtx�!�x��-�rOz.�s��r�M����$����O����h[$c0lX�N�d�<�D�S�d�&C���c�,Q�@�����D��dZ�x/��굨MH�ܭc�K�>y3�^�a%�`�djx��Z��U�0��b04��`�&z�x�p�)U�D��$e��Ӻ����;)z$  G� i˼��RM�$4�}�mH�-)Le���'T}I��֕Y����,����S*Tw.��2,ݶT&����{���)Oٮ�YnۄY��3C΋b��	�-�f4q$�o���0��B�/����iGQ}B`��3^2�ZA��rD�`�I܋�b�Bnțu��8(#H�(&ļ*�!F.hd�x��^0�(A�o�c�2x)�K�\����0`r��s�)�����_0D��X`ːt�S8h_�P�aU�ƬB�K{������'@�l�z䪰 Ih�Z@�[�u[�T�TY &ye���d�� ��)Hl2Jaʇ�H�����C�Q�b��@9p"��R!^��0ǒ�#��x�ЩH�J�z�G�>Ҟ�p��H�4*�-;�L�)`��?h�8I��!�/H_�H��Q:U�-@�ĸB�h��H<)/�H˦�)W�&}�&��"�d�'�R���&O*A�L�W�z�L0�S�R���~�l��s��y�=xІU�<Q���Qfb �q�_���[;E��S�.�\��xt	��%`0��)��R��H�T��j@��E3Qb
}�<���D. X��@�R������P����I�10�*q�m-<�'� �<1ǌ8�.9��+����t'�t���3�͆1��aB.&�L����c���!�ڋ#�l�`6��1j�j�3��'T@J��N7P�;2�M4f�*���DM�BT��8� �_n�Zsl��(L�O���w'S�8�΃VTp �
��� ��;c�B�M��rT��ԉ����s&.5؀b���Q��A��
ٰ�E���BZ��EO%_Fl�g���z�Մ�=z=������Y����Xe��\�U@��v�4B���|����ȓ)�� �Q�C*2�q'�6W�r4��VBHql�®�2��3tHJ���*~8�s�E��~���QҬ]F��i���[w��
�Q
��ݱe���ȓ*x�Lk��}�a�M� 1���ȓ^k�� �G�A�X���D4hȰt�ȓ��y�������X��۷
\d���$���ѕ\q�,u�v�^r�� �ȓTn�8�`��P�n05��m0�=�ȓp�j�1�腴��t�OZ<+�tH�ȓ�@��% �*E�:I�c�� ].��ȓX*,PG�V�2p�S�298@��p�����	ހ6������@��ͅ��`��dA�1(<`8�II)gfI��&�����AN��J	�p�B��ȓ*#F��tOÊW>0�3c��#(# Ɇȓd�H�t���:��n��j% 9��g���D��2���ϛ�R���p�Vmӑ���Q���P�jd�ȓ+��	r�ܺ�@�cኺ;pb���i��L@R&�����"ߤ���kTىgN�G�<��#K�6"�ȅ�n
@JQ׌A��Q;р�(	�d�ȓw�up5�G�:�Qۡ��lXb=��Eb�չ!�ƴwE��ʓk��} l�ȓ8�쥙��#	����.vذ�����9�-=T��bG 	LLh��ȓŎ�I'��5�"!H�"ЇU��чȓ"�e	�]��}9���h��	����Hd2!�(��o��>T$�ȓq��%�̖#������z+d�ȓck0�Sen�;j�Rү�9����ȓ[6(p;��-�D�� 4g�谄ȓT�����c�� � ���X0��p��{rn�@ ԭS����'U�!zхȓ|�̙r�V)|n|�Dj�)k����ȓ ��y�7L�H.�9B�g�A@�Y�ȓVHJ�z���˜�+�)A$ډ�ȓ�a���_���1��<C
�ȓJIJmZ�L

o@2�:P�-�ȓ&���b�:3��(S��h�:P�ȓ@��|��
��Ik2�c۞rb��ȓ}�Y8���8@,F	����w#R��ȓd��c��/OhHY�cO=5ΰ�ȓCO����*0��286 �ȓ4�a؅`B���pjC�[k$��ȓ5� ��,�&L�4ҶY�6#�Q�ȓ>L�T!���9Vr!�βxl��	�Dr�"��	��("�fY�S��	���J�h��\,7n��X�J6�RC��8�0!q�� ���Hم`U�D�C�	sI��{"a��-"P��d�7y�C���I@��~�l�X��Ӷ	dJB�ɋUn����dK`5t5(f��48B�	�=C� �q��7m`h���%>�B�	5P��YxG�R�^L���P)En�B��>�*�m]&�N�x�`ϴt%TB�	
 ƌ h���,%>��F�˥chB�	�'�L2a/%��4��I�I�&C�ɠ,���Q�	
������B�)� �p��޹T�R��2HO0n܄d�%"O�����;�*iȈ	�h�j�"O6咑F�
�c��+i��4B"O�lY��A�C>��@͍c����"O�4[P X/9��bg/��QV��"O X��"P) )Ҭ{#0�x�P'"OX��um�A�W,��H��ݳQ"O�9���>��F�-���"O�Y�f��8e�m��#c�6x;�"Ont����0�H�2��+Zz\�"OL}{b�G�t��"QGG��"O:���+���H;wa�Z8*�j���r����^�"uV-���7 D��%�I�!�ă^P���p����0`�1|!�X�~Xl�K��W N��r��S_!򤃠P�����&\=��`[�r!�)�^�H�M1)v�Ɇ`�:M�!���S;Xt���,&97F��6�!���o���XT����z���04�!��B.r���J8V�zŚ6AV!�d1
�,I&mU�8�ys���H�!�C�#F@��c �":�6�3b)J4v�!򤞋�Nd!�����`�
V�1�!�щI8�aHa��:��dz�*M�!�䖆Tۆ���̐+~� z���'J!򤑬ܬY�O�p4�2�H��J'!�ыu�BIP�ų1���&�F#!���z���)�p�\(p!��g|j��F�.��B�G!��?x)����:>����%X��!���t��2K����r�#Q]}!�R�X(��&�B�9�� �T�	�(A!��\�A�Qq7͚�W�~ ��n�-E=!�$W=d��e;o��S��e��mܘI>!�$э>I6%�$MtFA���G !���	zH\�*֔|�Y2�
G�2!�DQ�Yu��"�`�� i
pP��C!�D�<"f� �q!T�Y�A9���mE!�z@�;��H?k�� �5��A!�C+o|X��TEϯ���R�Mټ(�!��]	 ���kg'O:��TP ��(�!�$�]@��GG҉H̖-���>^�!�dV h �`&�X��`�pѢE9Q�!�Xw�MH� щ+�N�aW!A��!�$ߎ@
$%���]�y�V`c���<s!�dgS@��K�1l�1��iИm)�B�I'K�aiF��3��}cS$ӥ:�fC�	�y3d�S���Fz�i:�QnAC�I�6`1#4Ǘ�x);2aʥ1 C�I�+����� ?[���i�Ǌ0x�B�	�[)��R�G�@}�G��Qu�B�	�-�9x�gD�;�D��+�W~vC�8r�V�i='l-���4N:�<��a[0�C
x���d�T�C�̜�ȓ!�aca�C5�̴�T�\�2�܄�x���j��J$%04�ޏ�谄ȓE�h&���E�`��6'�B�ȓ`����\�|�*�"����Y��8��y��ԧ�b�h�j. ���}߮D���*.N�����7�@��ȓR��U��� ��q�`�Z*g�%��AE���G��u-8dY����x6p͇�Q���OG0?,6��P�8H���ȓb"���%�2��+ܽ�.���S�? �5�����[k@	Y�N�-��X��"O�1Q�o�#e��$ÍU9.��\�3"O��;B�ĀPQ�Pv���v�~,�"O�h�c�8g� ;��T.��i�"O��)�\9z+�G�3]���b�"O��A"d\�O���	�fŐ.�̨��"O6�v,�a�����,7�^@2"O*( fmU�8��
�jT��R݁w"O��FE�Hcn�����L�<H�3"O����F'~���"e	DN���z�"O<p�A�Q�b�`�7�@�ސ(�"O�)8��L'8���6�¹�`��>���Ҷ�G���	���.,Td�� �4A���Ċ#PD�ER
� ��I� Mfx�4
�:i��8��?R��<���T>� %KIC,;4�_
o:���$D��y�ȃ�lȨc�Ɍo'����!D�X�3A�,�c�Bc7�)`�L%D�ء��W�xLl��QN��N�)b`5D�샖kJZ_4��F�g&zdrƆ2D�����-hU�5��E�0���"D�"]�`y���/�y��m6��hO�ӨxA�Yr��-<V8�ȧ�A��B�
7��(�a	=BJ J�ƛXi�B�ɫ<�������~?�U�&KŮN�B�9Qu��at��4�ؙY��<7��C��<`�1Y&��X�ڨ���&�XC�		("�#7�Q�]�� � ��/�BC�	�6_4��0-�6UV%8saWX�LB�I�S�����E��QHԻIBB��b^F���'��y����?,'$B䉎r��"g�գiD��)EГ/L�C�I5l�xRe�i�P�����s�C�	�y����ӋJ�E�8��Bƒ�[mdB�I&� �0�)65�����P&ku�C�	�jY��W�[n��Q�L%<�8C�	�G�4���B�u���@��ֿ5QC�	|f4$���Q�D��wo�B�	!s�\��s��P�kBbֹ|MnB��� !�#�a���#'VS#�B�	�$bT웁�¦uV���'�FB䉛c���h��:^��a��X^B�	�s��*�I�rW�qP.�%S@(B䉬s��{��̻n�^����$�dC��!����VV�%sfQ�`,�*G�2C��B��d�ʲ|�,�'�7>R#=��T?�狞�9Y,4�$��fe5D�<[C��;��Թ��7&�� �ҧ0D��k�O��H��o
0(�P����<D��ca
�0v�4c�ϒ�
Xpk8D����O�!�^����O&^3���5D�tC�� �Hլ����&M��jqi2D�x�@O,C�*bJ�xր�A�C�I�t�^���)K�G�x�a�Á/B�	�R�#o�;rL��ת��G�R��ĵ<��G�1a�qB��ÿa����D�F�<) �:�6�K�gH�\9Υ+��H@�<�2U���sQ`J���@R�<��.Y# @A���z�i"�Ph�<9Ab5Μ� �G
?M@��w�P�<Q�m�'�raj��u?�t��e�<���T�B�B��&D�iq��I]�<aǠ�k����B�e���d�@�<I7�S"=�0�!Ì�:��@B�A�<� �@���>������dC��`U"O8 �D�G��nu�����=6.(q�"OjASFC��Y�0��F!�F��5��"OnTb�M�
I���{ �	0�N��"O$M�g�T>bzmK3�Ñb�� ��"O��9�ašPͨt��fu��P"OHD[6N�>�%i@��;
\r�
�"O�y+%"H!$�x(%A�z{0)Q�"O��h���\�.�hQ*�A�B���"OB��L�*�ڵYgU8l�Qٳ"O������2 |�b�F�%R��٠"OB��WI_�I�I��̩>����"Ob�ۢʑ8mB��M$?�B�i�"O�D� &�B1�"�mK|Q�"O��	G"_~�� go^
R��pV"O�xq���Z(�p�̌=� �c�"O��S����M��lR�I�#�����"OP��Ɉ n��%k%h�
��� �"O8ш��Q�p�^|1�Gݚ~z �y�"O�)r+�cjlX��G9v�8��"O��ٔ��j	C�fH�#p܍�'"O$�":_���E��F��|��"O�H"s�G����OĆZ�f��1"O~��h�1Mh�b�Մ�Jd�G"O� �T�¦)�&�.d$�:p(��!��7`Tc�\T�5!�F_�9�!�J�X���C�m��&�,����5R�!�������ϛ�y�2�1 �BQ!�ںZ6$101
�m� 3�K�r�!���D(��K�]4f�B�1.��!���-�6<&��J�V	���R�?l!�D�� H #U�O������eZ!�$Mf�F�[f�ɧ/�Fl�� -eA!�dř<c�,x��H�]��IUo4~�!�$؄
��uR$�?R�l���GUd!�$�ps�h���ܛ�r4+�L�kS!��0�t�h	d^y�!��,#!�D� ,�  �"�+%bT1��83!�D]�b�l]��hQ�� ��$a�!�B�RUAK������n��ITb�H�'�y���R��,����Cn��:�'[���Sḷt��%z�<a��"aK��^5�h�SJ�s�<iqaB&ֈ�u�;J`��� �d�<�u�T�^dQ�M�:-%�uӃGc�<�M1(E���%��ta	e�b�<a4κ���
�Y�O�b�<���ˈq�Z�����z�Jህ�c�<Qv��V�����T��IPӠ�G�<)"�yC�����^�0�H��N�<��ڃk��mxRg�d8DB�p�<a"�Ųi�Bt�1nԏ^ʂ�����c�<�%L�_���k��KA!�w�<� �F�F�mS��W:X��Bp�<G.ʮ6T��g¨fW�ґ-Fh�<Q&��?s9��j��Z"0�q�?T�x(2�:b�&��--?��c��?D�T���Z�.�r��]��H
�C+D�\Z��ĿMl��1'ѵ+|�)�#D�|IuĐ�h�^[W��d��'"D�D2���-*�"� #D}gb�;��4D�Ӧ��$oT��V�&�DlSa�.D��ib�6��I@�Œ�7�RI�ǈ*D�hG-[d�hQ�&�Q3-~���N#D�� N�b!��=T���Z�%Uu�F� �"O*p;À�4'ܐ쉆�L%b�,��"O�X��G]61��[�/y	��"O��#Vj�g�}�tn��J���
�'�"�;U�,�>Pk�R�"�'�V$r7l\�W:��p2��J����'����� �r���KR�I�=f���'�����8 �$%��g��	�'���H��$v�D�C'b��D1�'�HԒ�^&r���.�e��c
�'�������;rI���\u]�ɩ�'�r!Ru�\"@&�,	��Ա�f�<a��ۯ$�4�
u�ѽ9xz=�6�Bz�<	E �/װ]H�Ը�n�+���{�<��I̲nji�1B��[%ǖx�<a2	R�(3��C�J41ve[�@V@�<�у�Y��J�/	�Lc0�a�<�D�;��� ��'D}�UT+�D�<	� \�v�� �6�RQ�qi�t�<�T��Nnh�#���f�v P���p�<���11�}xG	�Zӎ@Q&�G�<	W�D�Y
�Rp*M���i�<QC$A&1JP,bB@�icb9�!c�z�<��kK "�H�C#�I	'VT"a�x�<�+���"���܍0-H�%��M�<�4��<=�Ƶ B�e�|P���Q�<q��#��dhV�>$����[P�<9�jU�ǀd ƩW�y�踰dHI�<	Я�2�ƀ���4{��@RL	M�<@�>-Ѭ�0	&q��T�pJGL�<	 �ҍ{:�}��̐#& ��RS�D�<	%��`E�y�'O�8\A�S-�w�<A'�[9Q��1gɟi��x�e��X�<�3�ݠC�$��W]�~*ĤBe�V�<a��j,�8����=+H��VLI�<�ƚ#Q�]ydO�>;o c0��F�<��*��MQ�����i���F��\�<)��8n�^q	�����ɐ�[�<y�d��]ú| s�5�	�d`FU�<Q��.N�QíP�n\`��[w�<Y�dh����[M��+T��p�<��̊�Iw��(2cԋv�a�#cT�<��bׂ;�J=IS��� 7�Ԣ)j!�?��X��#�1l����ч�%=;!���2�0��@��U�� {�&�>!�d�E��E8P��A�Rp��T/!�_N�489���7[wHLK��Z�!�$�7 �]�֫cZ"�˔��M�!�D��0(��ቜXv搻B瘸*k!���$R𘱦+�c_�����L!�Ć���R�`��J�>E�֤I4�!�$��p"<�f�� ,Dl�QrCυuq!���D�y�g*Ӱ2���VI1a!���	U���C�mE�O��Y�`C]%!�D@�$0��S�I�ܜ��^�F!��F���s&���p̂w,E/!�d��	S�P�uǕ�N�v`ʔE�6A!���;�@˲�� ���iQ��!��P�Yh«5k��9�e/Ǣ�!��/{���a̵�R�Kc��!��)9��@��-��r�J5��N	!�C�ASx���{��ኧ
�T!��<p62�Cdʣ4����QC�&cC!�����I�L%��j�a@>o*!�� ��4N�:`����U�<����"O�\{Ġ%���R�Ǒ�S��#�"O*-��N�-Sz*憊%w�� "O�5�"���Lvjy��h�4|d�i��"O&�����٬�y����0e�$�C"O�UpcY5Y�4ٚ��:u��9�"O�Q3�F�hL��S����=k�"OZ%�R ��w��g��i$t�F"OdM����=1Z��kA4Pz�4�"O�9KP�X�b.H=e�H$Td���"O�iء�߷�\� E�ӫoL�9��"O��J��ׄi��� $�6/�i�T"Om�����0��\hr�K�V�� b"ON8��,B�a��dh��\�Q"O~`B��#~\͘�G�=�ҡ� "O�\�FI@� �D�[�X@@�"OE�R@ �c�c�7����"O����i��W�Z	���Y�r��G"O>�7�E�/4N�2�=x�Z��s"O�U	A�X�6�z��� �}a9c"O�4��^�\����̬I4(�"O �z#Hү{�<m�b�L<Ұj7D���Ќ�j��$J4�T�pP��2D��ٔ��)
 yGяԜe�U�:D��
%��4��(���2�<��c�+D�3�J��-Ba�9��%Y��-D�ؙ'�L*'�H%斓9���N*D�T&L�7CQ�����V^�p��)D� �>�,x !�� U��:g.'D�Tc�+'[������H���1D�t��,�v�s�6S֙�Wd"D����
����&^$At�� wf!D��� ��!xh�2bN1U�l��f.5D��"Se�:/��I1���b�k��4D�bc�f�z\KqI�`VM
0D�8�u�c�, 	d�W�{� ��1�-��<�O��KS<��ň��K4oq`HX"O��JEh]0"	ș� �+>p�`0�"O:h�/�S~�١��� p�a�b"O@�3s��#j�F	���G*;��"OV��q��$�HQR�O�\6�9�"O��S%Ɣs�Z�a9�^���"O���7�E)	Ml��G��%J���"O�4�
+N�B89�Ä�sq6!�W"O�@afT>�>5Cc�Vfp2"O�	r������5$�薤%ar!��V����h��\xqq1n�e!�Q� .�g�7k��XІJ#U!��C�/����G�ep�EpV&��L!��X�Q�X��)bm|0Z�$/{��O>�=��P��G��*#����k۔Ө-�"O�bG=o�2d����ϴ�"O�A㤚�1Ѝ��gҖ�T"O4�hte�7e��6Aѳ�@�@�"O��B�tRbDˑ��>ZA4l��"O��8� �]�	R3ԜR"�$�q"O|����p&E�rN/�HbB"O0 ɔbX�_�W�%F�$4��"Oh( �9ռ�JS 4�9��"O�$��O�'X�Ī�N�!���	s"O�d�EY�H�����R�S�L�xS"O�| � �>x|}��k�?+�"�0�"O�8q��),�P$r ���9�"O���S*ؖ-���p�`�:ie�Mˆ"O� Z1�d��O.LD 2 Y/eB��"O�!�C�˯.(���@/m�hDAp"O�M2q����M�7��-�y��"OU��M��:�0`�s%�^���"O��f OF�)�j�[�
q"OZ��GL&B�F*�(�pa#�'��Ă�6�N���"N��zA��j�m�!��p�����ϡ+�P�u�ı�!�$2��P K�Sx���ÿ*�!�D؆-�*<�D�X�s�N��!��-�$B'ׄ>�*���/��q�!�$���I��(֧?��Y�aO_'Z.!�䑊U|�����%e����" C!��	xP��F�LGes�J1PG!��,Fe��S�
i������!�$<�А�DdRs��U�+@d�!�� ��m����O�EؠKJ�Q4!���0�Ubf��=	��3�Ō4!�d�'B���+���ę���X�W)!��� �xYS�dQ(������<(!�d�9b8�7�ɿi�\�:7ʂE:!� 	`x��)W
ޞA���,!򤘛L��	��+C5=����͝�	+!�
���$
rN^)L��QY���D
!�dS&&�X�c "KJ\(1�g��[
!��[�E@��?_�,�v(�,!��BiXRU��"������@�/ !�$�1����A@N{L܃wM��%�!��� N���4�Zxph�l�2!��?A	�l���r19�,�!򤖻J�X���g%��Ê¶
!�D}�.�H�Dͽ2��*6�^�b!��.�B;q���<� 窎�N!�d� �Nh2p��tĳvʔ�dd!�ҕ;�����@).�,P���ѕE�!�Dg2 �P�}��7�)C�!���9Y�1"Ħ�a)�;�Zt�!�D��_��Y���+|�����!�����y���]3Q�P+aE[�!��*}M^i"�gR�x`�Y�'�!�ϡF�Es �@	� ��Ϲx!�ě)8Z��g	�P�DUZ�:08�'��D��~b��J�����`q��G$�y��#��Mq!��]�:e`@hH2�yBbR�|*8��u+�&~��D+�bS��y��2,��|zG��)�La `���y�/Njj8�$��'�����iج�y�ꒈ+��x��'�&�f�yr��/A���i��T#6&��F�����!��|
�y�Ò�~��\8��M�lTr#�]��y�k�
Tnu3teH�����G��y�i�%;�h|�%#�BW,��y2Ǌq���+�
Ě z��c�K��y���)$`"��ΜM.>��E]��y���y|��QQ%�!=�R$�G����>�O��Z�mF�C�}{��6k{F���'I�X�����w8��쌝0��L��l$D���'�����"��5U:���P&$D�h�Ă�0+%���e�n���R�� D�h��Hñ`*L"�(LA���:!�#D���A��4�"I�Ӄ֕=��i�CH<D�$�*�"�������0i�1ʐ�8D�L�U��_@�)s���>V�u��5|O�c�������o�"sR��9�(1�3D�� �h*b�ڦv����U*,{�T��"Oti@��SJ�Y��J� UjL;�*Ol��5��Zhz�s���x�'pF�I���8t�eRc��1$%�q��'�F�CW�ϣN���	C�޿ �`�@���'H����M�u��` �i�	Pڡ����$ ;D�)^��mXä%��/�!򄍬n�-k��q'6l�#G�u�!�D��;R����G�k"p"I�l��I䟴��U�Iy�O�,�I��Yx���0eƳ>�����'��`[�(!I�g�P�0іx��'��Ex�Y(y.L	�@�߲��
��?A�yҀ��d�Pa�Y�	Ҕ�K��?�y"���k��U�b����y���yR��k`�����3j�d�sdJL��y"��	=��R���[��	��@J6��3�S�OG�0�`*X�U+�96,T�6[��P�'��d#���5u��IEE��+ڊ�)�'�t9��LT)�#��e4|�
�'e��c�dT�a_Z���aɚO^(`Q)O���䙼{T��Cg��6|�,�h���,
6!�_�|F�Qx���l��M؀�Ey!��*\�|q��¥���8k�	�4��H�)ʧ.���
2��hI��ɱ�^���t���M����A��|����	 �2X�ȓ{Y
�"�B�
u4,с�͇Z;&���)��asOG�JV`�д�	/�����B̓E��Y���� 0�h@���S�Lp��E x�Ð;y*(�3�lčm��Q����<��FZ�0l�+ 2G"��˴��U�<�b��3-�R��ת%9N<P�k�S�<�
2{�<�[�%V$<hǴ��ȓ�����_3c�8y W�[ �n���=��8����v}� �B�!.�>����������$��"uk�.T&P:���8�}�ȓ ��53���=�*�3třk�Tń�	�<�!U��dx(��M;�z��q �q�<�� ��DAX`�OL]La�l�k�<Po��n��`ؘB��i�VAE~�<�JW�,)�i���tLt�P�T�<���p����.".��BIP����F��9j$(\<M��A��p]���	u�'i8�p�fP{2z$nڟyp�Ń
�'�根%#�7A"�t�ւk��X0
�'���qD���)�"@a��Zx�Rd�	�'�����F�m�z� d̕?kS�@r	�'{�lqR&�aD��(�-�8�hp�	���y�N�"*� aC�<�>dR�h���xBa)I.�)�Tŝ�{Nl���燰Y��O8r��۵ ��kT�wk6��P"O*lb�ɃG�Y[Bb��,���x""O�'E�kTH�pNޑy����"On���m;rlP��U�V�%�8�+%"O�]ʁO�u��]�D���H��"O�i���Ψ좥�C �.���(�"O���B��`��3�ݑ\c��Б"O�%z�X��6���ݚ2mR$xD�'�1O��rOݿm_��aoQ�D3$ @�"O�Rvm����yr�rOp=y�"O>��A`4_�x�0�K�*(QR�
#"Ox���ظ]�^1aqj��|5�m��"O����6 ,1ŉ͙J�>���"O�����]�J��T�$�^��"OF|S ǎN�h��g�#'�P$0P"O� (��ń�,�PM	�^�-�����"Oh�R��� P�����!f�:�jf"O�X�c*ƿ�Ƥ��)�B�	�"O�9 %��,, �R �Ic��]��"O����< b�����+[��q��A>��ۦI)0A��"!N�h����"D��@��S,%�0]��)��y4\`2� #D�P��h���AP0o�hӐݚF� D�0��;N؄[�.��%;�� D��rq'ڗ�MQ&	N*C|��l=D��� ,y���
.eɜ���@;D������/����ĝ&nyr��O��O �=��`A��K�'z��J�O�t�����"O�#S�N<�2���c��d�R"OVX 2�
FՊa����<�����"O�m f�w[<���=F�a��"O�x�OG
 ���;$��'VX0�"O]�1	���z�!_�rRHI�0"On�3��14L;vR}+HA"O��%��%V��c���	}@0�T�'���������`V�H�� 9��9D�����e���Q��U�i�v��F<D�0r�� H|̜a�شwb4�#W7D����&�T$�e!$$�K��5D�ࣗm�B,�b �ة:�|�`/D�$����hI˕CY�3��� t�-D��� �/5�p��nˉ���6D�<��,��A����2|~����*D�ıF�=�(0Wㅘ|E��@ӈ)D��yc��?�=K��6k�rh��*O���"A3pN�� �/1���"O��b��c}�����-8k M3�"O�T(S�^�,r�Z4	R��f�#�"O�|T�Gg��r�H�$�i`"Ov���
�㓨���Ib"O
8��I�jM�萀7	
�	w"OL�Y���q|������0�"O*4um�^'��Q�?P��1�"O0lC'���V>,�m��$�dy9T"O�y�N�%8b�ԙDL)٪}x�"Oı��J�kW����?�4��"Of���3R����壕�w�x���"O�X�t�]�n���,�Д�"O���Ԧ�#d�`MyRcU�F�@���"O 8Jլ]����u�G=_�p�@c"O���ʙ%U ��O��M�e�1D��ZC
�-\�te��(8��ׅ%D�d�b�\����� ��YQ4��t�!D�X`�Uw��[Rk�1M\@�&�=�O~�	��xh`�D�x��M*1 �^��C�I# l���@����y�Aߩd��C�/�\ur�dY�nj�5X�I��C�	�N&|���N�2j�x���-ȱ4�tB�ɑX�I��� �	cr���"�XB�	-4���C�Z+V�J�Xǋ��#2,B�?F�0�y��V�*ٰ˙\�B�I%f�tz��Z2��HjP!G2��C䉗;+�h��&��ox��S��	|C�	�j��]��X�a��Z��R�w<C�I�������%gF8�2#/a�B��&����`���S�N�Q~�B�	4F`z�����_-"0���
!h���:�IX��~R��v;�혧B��`P��P��y�jڰ;u��2�Kdx�0�l�y
� ���B��5Q�J q�1v;Ŋ�"O̙�2%Y7z��� FR�6�V�*�"O�x1�gE���poM�
��L��"O@	��s�Yx�Hޜe�0�"O�t�RX�Q�	3��=*� j��'rў"~�����K�xcRmeGZ��Q:�y�L&@�t�S��LC�lJ&i��y��v����I%���c���y�!]��0���B_�ņ�Y�Aи�y�$�QG(� ��}i"�V��y�)_p��y�3A�{�.)��M�y���5c�t[@�zJ2Tpch��y�z4j��0C�t�>}R�,׏�y�	HT;�e#��=��E���y"B��Y�D�PcޅO��,��-��y�FF�s&���]0�ș֪Ȥ�y�)FR%!�cǪ�ceA^	�y��87���e	4b��!J��y�aY�<��Q
1KJ7$
2ՙ��̚�y�"A7.ZX$R�k\�3U�,�s����0����'��HB��<WA��H�HI.�����',R4Id��;1�Rh�7	hd���'��(�Ԍ�/���*��-{"\��'�<mâь����i�|�.xK�'�ހ�p$Ջw��ㆎ�
��pz�'�`�����1��%(s�΢v�䀚	�'m�I�RSN| � �7�x$S��$2�k`�@�C�_���q4)�3W���AD,�H��*6ZiS���V��ȓW����$�Z���]k���{U�5��kL���ܿp���O+w�!D{"�O�T<q���{>j	���@�'v!���M�;y,)��y��T{�' ��B��!��c�B�(le�x�.O�����X��@Gʈ-8�,B�L�!�ęH¬� D$�&�,�'N�%`!�$Q���Ы��n@�[�?2~!�d^I�(����WQ��ɳ��4sf!�D\�s �Չ�NR�|�X+$�+Q!�ښ'Vu@�G��D��Iy����^J�O���$͔Z�ܠ$o�}�V A����>CO�)��<BPjh�b�;"����"Od�"�:py�YYW�]($��"O���l�5e�y���̄e����&"O2�mU�/�`��♲&���yP"Oz%I�� �_�܄�����f��Ȓ"O�t�$�D�, D�(0-�'5������j�@&و �4_^��e3D�j���<@^�@: ��11!�.D��+�GG�p��h�ĕ=b���di1D����ãT��8c��Ba��ۆC0D���.�8����fH�pd~�t�:�����O.��,IɃ�A�w\�e��h�0��q.D��8�g^�I��1A�������-��Fx�$+RE#(�l����[@�h�'fFԟ�&�LE{J?�b�Hmp�L�q&�nf���5D���E�GJ�DA$#9�#��3D����Y�{�Z�Y ��[�f �D1D���e�9{8��hс��"
M�7��O��=�O�1O���ꂅ0���c/�c~���0�'�!�$�<}��(���,M�ш��btBOT0Ӆ��B��Q&9Ip����'�!�$��wwb�b7M�Da�e9�	�'�'Ia|��P�]^n�"&�kXʴR�jʪ�y
� �Q
��� ��@��#%���zD"Oн�efӗA:�D����=�dȃ���2ړ��č�Wd�sb��1�0�[d�/�B䉶z�$�!�F�k,麃�2B�I�[G>PRR(��P� ��eb]�0S.B��<���� {�]�ʙ8b�B��+Ly�(�ȄD�BK�he�C���(i�CKO�8��$ʎ<XB�(`����F��&K�H8U�	�ZB䉼�B07lLw �IyPN�mTB��7��J��]�d��{a�D3�
C�I�~& 	�d�K%b=��� [�Ң?����ɟ/[�u��<`8Cq⇌%�!��M�����̈́�7fr`�W���u�!��.X,�:�Y� ��1��`Q�lk!�d'�x� b�P�z�ָ �aǌpN�R5O
��#�׋J@IyGH�&$sj�"O����(�s�D��M�xo(:AS��D{��	���rbd�?&J�����4�ўP�ᓾlhP�����tct�6�%	grC�	�m�4̑!��:�Ht(��Q��nC�ɩ>�l���A-j���a1o���DC�	[�IK D�V��P��X�pB䉡8H�iB�ϫQ���`���#Q�$B�I�xy"ܚ�n:I��P�gXʓ�?q��D6�I6 ]
�	�É�	�0��b�'^�C�	=�
=�0��!6:�;N�C�C�6K���PE��Ԅ(d!S�"O�m���t���1X�y:��G"O(�ą3p�ڔ�%�̀:�!'"Om!q�h�$Ÿs�S�hj���X��D���7�]"F��Fh@s��O�C�ɣ\H���݁h�N���ĉI��B䉖Tx���m�$ dZ�I�(�p�O@��ē�N��0��,>;U��[2!��A�unlb���X@�J�I�,#!��Gl*��A��Z�Ƚs�.D�l!�D�XسFg������[�1W�O��􄄁9D���̕
k�D����Ψ+-!�d�5_�U���47�-FB�G"O��:�L\�27�5���O�)_�y�|R�'az �;/� �CN<+T(H��I��yB�d�Z�&R��0��$I0,�ȓ2�ꔈ���o�n��F�^h��ȓ(�j��F�H�e���1�h� pR>��ȓ25~�@픬`���V��2]8BI��P�a��,
�L�Ӎ�_`��ȓ�r�K��TZG��Ge&��'~a~b�>]2����_�@������yBOW�$�x�@V�9�\�@�A��yڧ�T~�|a��@;F�r���<D� ����	������@�r�6�Y2�-D�lp��Nn;�0�b�߃^�Z�l'D� �B�փS�\h�D�:2���(�%D�d9`h��	�͈U)�4*Xy$D�,�1'�u�� ���V��A���$D��z4 Æ}(� j$+�'����l D���
-w�X���	Є9Qx\	��2D�!p�O�W(p]�!�a::�[�g�<i�D�R���H�=݀��@��<\`���ȓ5��ؗ�Yu�]�p��y�����J̓l����)F�ĹX�G@>*E�$��\��Y��LٿahƐ��&ɷ�(��ȓa��I�D���ab�շ)4���S�? �qz#,]�����MY?�&��"O ���6����?v�|{e�|r�'
Nl� �;+��BӇ �-Pd q
�'�$(X7̑�1@z�K��Ha
�'�N��dJ/$����wɦ-k�"O��Q%���m�M0��B O�Y%"O0����ȵ
�"��n�Y�G�`�<9t�΄�j\����Ps�P��f�`h<��"��i9�DY��E�ǆŘ�y�\�m�d�IfiM�yd���Q�Ҽ�y��\�X� pš��"8IH�
>��?y�'��H@���+��%y\���'�P��w��\_���q&�
Vui�'>.�b��H�H�{��W:T�\D��'�yB��HԨ��Z֜9H�'T����*_9f~�0�gS����x�@�o�ƌpw�'%¢�zV&L��y�E�Q�����+ �"�����y��D.h��9;��}��8#D3�yR,Ɛ@�h�Ǫΰ7Z�U!�)�y�ϏDH�S'�V(S��DQ��y�dУ�6m��.���\��	�
�y���!�L�3�Y���)����O�"~ʑ պw�ЕA�?j݂U�5�~��hO�L����)5`Dx�(�<\�؇ȓMF��]	t���g虾2D��ȓ1}`��#e�.@6��η!L����}0Q7dіD���@�ʹY����ȓG�dbeִf<��B%PVu�ȓ<�D�!f/��`e"�"V ό	��q��]���)E�}9z���N�l;���ȓ��S�	E+]���26D�[�݄ȓ$�dM0I6��
��ߨB_P�ȓ�Ɯ�0[63J�r���=✔�ȓ(Hlx��ƴJ��b��C3�E�ȓ{���P��I�b�E\~�@}�ȓK���)]�r D���Ǜ�H�'.a~���a5�X�����8� e��y"/�f��2���Ж��d�T��y��U!x|0��Ҿc�A1C	W?�y��D�_�*,�PG�VT�S�"�y�A]���PVbހX@��Sh�9�y��Cc��A��ƈK�@1c�H9��>��O.�ʶǊ���ш�8'j��"O�l�b_'�]� �R/3h����"O�q�E�A�ɸ�-�O0��@ "O�-�'GG�~�=e�Ƀd!�t�B"O�}e� � �
�̃�s0�#"O:Y�%I*"�����*�s��s"O@��d_�dBFM����+px�$�!"O�僧�]rW��M��pI\�z�"Ony$�!��-Q2�z���!�yr�	�:|�uJ�T�� U�С̭�yR'�c;B�����?`���)1�y� �p���AV�ڍ�\)�'%��yB�J@/p�jrO2N�q�E�7�yB'�'G*��mu�f�,Κ��>�O��%j�	������D�}��Lr�"Ov��`ז+�T�s���n�Jt��"OZ�1@$X b}���M�Q6�y��"Oniad�2�rUa$\(#���6"O��x�J��o"�!C�[�eU�}"Oԥb�.�:P0$вۦwI��Q�"O�-b�FZ(�HXV-S�=�\zF"O� �p:�`<!�0��g�I<����"O���uL�	 u��C��K(��"O0P�)��um�(Z�i\�ȳ"OZ�#�lG��L��d�_	T��L�b"O��#���BDT�D�?J�tɣg"O<�&AI1xNh�j���B'T�Xw"O��`�aPEz�����"g>�)� "Oz�"��ǒj��� �T�f�@4"O�D���e���C  x�Ĉ �"O:X#��+�\��s�&i�6tpB"O��� �?A�@ {�H\51�V)��"OJ���&QsI�gσZ��y2"O��'I�&,�ȉ�׆�IJ�Q�"O����)U� t�9}3� �r"O�E�q��:3�p,9���$.�"O��{�eøl�n����4]��X�"O���X�����Դ\�� bV"ON��D%���ٰ�# e�[�"O��1�\>N���'��-�X
�"O�\#,�N*�(B�K�~��z�"O2Q��O�>6��M�aS�J����F"O�$�U�]>[��d�ĝ�u�"OV9(�c�2$v=0��\Q�\ȳ0"O��!`�ڛ'�	
4P�.;�e@�"O�q2ccL7s�V���'�:+$V"O��c��h�  rm>7���"O��Yq)˥����թF�{���;�"O �cc�5$=Zxa��\�sF���!"O���A
�;� 1��Ď79~�F"O\$3�ɪd%"��s�P�(�"ON!�P)�%Z��V��B�Ш#7"O�ɩ�C�G�!������ �"O�Xbpm
�+�xab��#xf$AD"O49����&2 8�K����村�"OH� �mނ<_B��ȜQ̙��"O^	��*�����E��W�*�"OhmBt.F 3��ЂZ4d��#�"O2R��]�/��+�����N��"O���!δ4�b�RãX�zT9�"O�ͪ�락(-$��I�T}2��t"O0�3����3a�ɺ��Q]�p��"O�}��L!g�T�b�O�)�Q "Of�õ��b�~��5�W��"O:eȖ,�.J��7N!H*t�"O��AQ�n[t��N0�2����$��l*�z��#��uh]�&�^�{A��V�<)��Y�F"L�q4R�M�Zqc@XS�<�`�'Ğ�;3��M��k4�IN�<���hi��Ei��3~R�ⷍ�I�<�`�D*a޲���&�e��	٦�k�<A���hh� Te�5���v��f�<9�&��K��	�"Ӿ}�b$��K��0=���7k���CK9	�"���N�H�<a�<�pyCmɫv����f�A�<9���05�<s�)ԿF� Г��I�<9A�F�lƂ�C�:o]xx3���F�<��ē/��9�N�ҁ�6��D�<�v�K�g���q�^1Ew���o}�<	r��&>���GV�	��
��_�<���	�n��T ���W��m-Y�<���-4VjE�rh��v���Q�CW�<YăQ��E��C�N+@d9�O�Q�<��\B�2QSC���&I)�%QM�<�t$��t�tU���� �Xi�6��E�<� yÇ�2'c�=�7�<�ܵX�"Oz�Ԧ�Db�#񧄎/dՙ@"O�lxj�F F�I�~ld �"O��!2�R+�R�s�M�"_��Y�"O�,�F�,�PhA��#5J�I(�"O|-�Q�.I�]
�
/�؄��"O��ӷ�<]1�,�4%G�vp>ͣ"O$�(r!G�OϚa���+4U��Kp"O���*$Q[��_�wb,u�R"O����9�X���nǯNK��)E"OLPP���GQ:�ZŇ�J@B}�"O�H�+D�pg0Ԩ��˞Uf�H "OV�+���z��6f��%^�Q��"OԄ��d��D��Ъm�8	b"O�Y���M7��h�SRFq�"O��[��p���Z�	���p�"O��H��,��x`�޴6Ī �"O��	WϜ��X�c�`Q

$@ݡ2"O:tIG[�X����"-:y0"��2"O�a�$d&�H�a�,#��"O���cERc(�)�2��`�t1��"O��R�|授�M��^����"Ob7H��@���	
 ^6��"O�AA��j�)&�P0^L@ (�"O�͘�"�1't�L,3O>�m�"O�%��
D�V�Bu���ڰe=B(��"O�(k�#ʏ3�h��'�"6#.1+�"O�(�g�0	纀{�'J�F���J�"O���aƀK0Hu�F&�6T�>3�"O��S	����C�%f��5d"O��BÌM��0Q�&p��"O -�U(��wm�|�s
֊id��@"O�x�-��a��d�T��+�)c`"O����l�I�����A���@ �"O@%�֦�C0M 	��Q�.��"ONձ1��LXL�q(�`�֑s"O��c��.Q$�Hbj�/ ��ʲ"O�R����'0�X� ��^y�s�"Oh��*дA��0vϜ o�fU�"O�h��.҄�>��B��e���"O�3�MՕ}�lM '��2v��QW"O�d*�'�r1Ѥj��*fu��"O��z��_'K�H���݀�R�`C"Ov�!riې$�V0�T~
=�"O�9"E,����e3W�U:�"O�X���ѐ\���m	�O�,�g"O� � �8�f��&n'2��}b"O�Ъ�C���a��у_Es�"O�aX���GR,Y�V,؆bpv��"O�`��ۛm8*�p�)ָE�0���"O��k�U�uH�a�7h���c"O��!#��� @2 	<��"O�X`e��Y��a���:��u!t"Od�
�+�%;����$��jВA�A"O
�l�6+�̰E�߶P�"Ot���#i�yP�> y�"O�z�(ɮo@:�0�l�h��h�"Oz����L�g�6�²��CJ��Xg"O���$�Fg��
� ݌4��C"OJ����W��4�1.̖j���g"O��sʗ^r�6)����tH�D�ȓ2��rv�C�.Ve'�6X��T���
�Q

:z��aaA�W��!�ȓ>��
��:�4����y�i��S�? �Q(�CƄ^G�@��D�S~(�(�"O�@h4I	GDL}1�c�Fq�)��"O��K�,L���=��\�eeXEj�"O�� �AXT
X�@W�^�jy2e"OX	�#K�LB��ҨK%ote�"O ��ݯNMt�󆚿+z�s"O��X�&Ѡ`�~A����>g��(%"O�u��"��VLx+5iف$yC�"O�D�(�v�9���ފEp��"O���('!~�S2jW><6��"O ��b�:XDd�!�I̕�4D��"O�Xr��Cz9��.˽U��ŲC"O,��P� vJ��g��w���yS"O\C�*H02x���(hԙ��"O(�ks��2eP�B�hߚRN�a "Ox�c��Э7|�����*pʴ"O$݉�l������@8���"O>�� �5��ɚ&�'F(]�"Ol�-nX�����@FI��"Or��Fw$Hh5���s)�h�"O(��ኼ;��M*��X$���"O���_���ᡥT
�❈g"O��RF�de�f�\r�J""Op��o�11���;��¹ d��0"O@�0Ϝb��T�������"O�E��	V�9t�Q�G��p|z`"O��`WH[�v���cHo�j���"O:�k��L@�Lp���H��"O�u�3dG�������>_��AG"O�A��F�@&�/��+T\ɳ�"O"}Ѝ�;b�Jy�O[8u> y��"Of	jV/�Q�ޜ�7�FV:�
 "O<�(�iR-AΩi��8:Y��"O�d� �S&
���ǒÀ���"O~�on�<�Bs.Vr�� ֆ,D�����wj|9%�{� ��7D�H����t��Ё3��&��27/*D�([�c J��r�'S���(#b(D�h����p!�p !��J�f�&D�T����5>X�U�2� w�/D�0c�I���#��2Y �!QL-D�(x'�	�T�6U� �T:��s��0D�,h��4S+�$yw��;� 
!D�H�1`�
O�����La��Rp`!D��vT�~��]� �L�$����#D�����|n��!j
? ,��a"�5D�,��l�4*�vh�˕�^T��1D���1k�HT�s"Td{کs��/D�h:���{���cH.e�0�:D��Q�J7^ș"1��}(�� 7D��3�	�Cl��9'/�K���F� D�@��*&v�q������A�*>D��S�ж?M�@!�đŜQ�т!D������ I"t�J7(D�y��C!#D�4z�拶U���h0�T �t� 4� D�|�BF�B-H�SR�R�b�����(D�b��k�� ǎҲÆ I�1D���u�	m0pA�T��%R^d�w*<D�#R@թBo�y��DQ�F1J�+��&D��9�(G���rR�Ɋ|&V(��8D���OӼ{16D9�#�
L �1H7D��HB*C`XzmH�JD�0�A�:D���S㍷#J)"vg���Li+��6D��cǌ�� ���ѵa�b�R��3D�� ��W�Җ-y�tr��/�f�0a"O�Ġ�h�ft-@AAV[�ʭ�S"OPu�#K�d�����OĒj[�"O� ��DZ�}
 ;>�|"O��c'*z���Rt.����f"O&|��o��1	�<K"-�}f���"O�(��M�< ��0+O��`�P(""O���sC��0�IE.�e��z�"O�pذnL�q_-���UR�p�"O��!�'�v�l�"Ƙ�`%�I�"O�%��2<ʼ�p��(v.l�a"O<PmӀ_n�S$V�.=�A"OH�x��יmv���*I�b�b�"O��3��ж@�c�m�� 6"O��*ĥ��P i�U����� "O�� �$e�0����[Vu �X�"O�P��:E��Jڠ���q�"O���'&&N6��U���;�&�0"O�Ř�gۇ{m�<�A��!mFV]{�"O,%��Euz`�ұ �,d1����"OF�Fŝ�aҊYY�@��x*�"O��(X�jW�<
A-��,�q�<�&�5�D[��:���+��F�<�D� rz"��S� ;/������x�g�5gf0�*%�Q�#ϔ��$e�͸aB��
��ub���A�T5��p�������'O�,�g9v����ȓHኴ�� L'Rdt1*B�4u �݅�"tHct��4`� @����4L���N:"Ӗ.�/,NtX#A�|����ȓ|� �`��M(}���e��%����ȓ/X�e�r�Ǘ3I>���ū����w�μ�Í�"�2�`�l�,P���ȓoH�S"�V����r&���J��К��cm o��q�H�zR�1�ȓ?�6҅͐�D��$	��CO�2�ȓb:L	!`���a�0�,U�;�$��ȓT �,�v�H0W�~�Є�Ċ?����&����{�X<x2��s�-��mE��c�!
t`��fRr��c �%�`8�,�X�@� �jt��s�XM tEBf�a@����eu��ȓ
h,T��ǌY, D�ʵa6D$�ȓJ�tya�R�N�y�@�43�x���j�@�!/C`F�k���?�����K��m(�FШ/z8���Q-F�y�ȓ�2uWFLb`%+�V-l0�L�ȓ��"j�o�h��� )�$��=0J�:vk�p�D�J�L&N�$\��)�����I�#�Q��#��?�,�ȓ{z�����ӊ@_���R&W�-��Մ����SC��N��c%�O�̙�ȓj�RH3��IN��!B,�<q�ȓ%^*Is��+69�9!������[�N��V��-C!��Hdi��$V؇ȓ!8��TÀ�lD��H��ƥ+�����7��u�������<���"6D��� �B�Y���reZ�m��tKCN1D��0���J��a�Y !:�!SM;D��8��Š`���P�ء_î8!#<D����Qn2IP�*V*qƌ�R�6D�l�P��e�n��6��U�����c(D�ԡd�,v�p���xX�v�3D���2�
>���Z�/�
,�8�0D�<D�� $��!fJ m�-"� �z2}#�"O�Mq5%�p�b��M�2Oa�PH"OPmZ�M�{?�Xs�͗�vH�8�t"O�5���1��pDmͭsF��"OR����y˄�4�ʙ[���Re"O�AB"`)����J�^��1�E"Op<��"U6T��P��4�H���"OPj�1KM�|�#�O�4���"Ot=�B^���L��/�y@�"O� �b�D�}�4fљ%����"OtA�@ꊺLx"��!f�D���"O���J�J�!�o~cƼ�u"O*ܰ�k��8��H�;Zp��a�"O$Hu�  U5D������T�1�"O�1��.K:,Ȳ]�����"O�d������
�QI�j9�"O�MzQ(�	"ԩ�\�Dz��0"O���!�%[�x=0Q��7FuH�"O@#�>=�D0Ps�U,W�e
F"Or|XiJ0K�$����M8?����"O�,�S����H�P��V,8!�Ǖg�J��4�s��Mpt+�?.!�$�1���е���f���jF�!�DЖy�6Q�O��Z��t"�)[�!�Vl�f��V/�2f��"�l�!��Z�i$���s#A�/K�|BAE�)'�!�M$=��	�	::��;e�(5��HE�D��?��t�W �p�a���E'�y��J7O<.�S��T�Rta�D��y2%2:n�8WG��F�n�x����'>ў�O3�{S�ʹ�8m
�o��,8��p�'~8ģ�.%#v��K�!����'�0i#F�� ^��������'�0��By�~5 5�����0Ӎ��)�t��J�(q�bH��c���yU�g`pEMB�E9�8�h���yb�ϤM�"p*�62�X�X�ޥ��O�
 Ǌ�:������"@�`#'�D�<�1�R$O]�A#D�_�h�C��@�<�w��}�DL��F�-x�!'I�u�<9a⬻��8kА��
��p>aa��x)��647>hHb�Y�=U6���	8LO��'���Q9 �X�.�Cʠ�cI�N�ў��e�'�>!�7�/����U�����T�0D�@6E���@1�#LR ��0@h0�	E��$�3���`l� qlܠ�G��qh!򤖻
�9��R�h���i<|��'����!\O����(-,���_3�u��"ObT�#�M�VB~d��Ή�ڨq�"O(���/BȂ�j¨�ɱ�'���[g�P>�p���E'~�Z�%����U!c�J� +h�
Qd�r6�I�<Q��_�{�(Uҷa��M���Q�(D{��鄪]�|���?k�T&fQ�V!��9K�x��%R�%�DY�t�҂!��'�a|b�ɭ<	D4i��D�M���@��y�N \��VhL�[Un��۰�y*҅Y�����P=X��h �T��y�D��f��� �ɾ��ˊ�ָ'ba{��1	6t(�-o�(:2a���?9���>O6��fcX�Le��q���L���ȓz��k �����	��/v��-�'O^����;4Մ���Ϗ� ����\;*��~�[�Ęb�S�Քy���/P�T���<D�� ����--I���ڤY: �#B��B�O6$�y�@-l���
�}�V-q	�')�k�FA�H0��V�H)n/�I�	�']1��/H �=��̫5�V��'�xacQh�KI�\T��=KD��yB�)��DV^���Y�A�p�DMZ��<B��$�H���V(��x�7��XG>B䉜�D��Iٜ2����ۿ\R
���<��/�R� �	�JX���u�<Q�%}	���Q�蕓go�G�<�g
�����yDdӔ	>6�p���i�<	Pi�#�"!ps�K�D���b1Uk��q8�Pi炘')'��S!oƘ��U���>A�4�~�ޤ��a�B¢(�f�#0����yb�֞T������h�Fj���hO���I�K����eމJA1E-A�!�$<����'C�;�Tzu�̸n���@��(��X+	�Y�J�!p醷:T	��"O�Q�kA*%�Ii��ӠcXI�>Q��"�S�'�!�6.��o	%��"(&�1�ȓOp�l�&*63���eg��{j,�=�0�0LO||�!ɓ}9�!`B+�2:G9��'��	9jl��§�Y0H��q�F�E�l�	|���s�H��m��KC�O�X�����n"<O�"<1u/
s+���f�%@�!����<᳂;�O����&l�4�"�� K�fMȗ�|"퉰��"�4�H��Q�.��qX�Y&-��U��Kp�鵀YH
�y�N��&�X�ȓq��dS��l�����'�ў"|�rJX�
�,�㶃N9WOj��R�<A�F�"����-�6@kJm*% |�D$�<q#+�!޺�{w�^���<D�(@���y
�q��D��M����`����&�X�<	��,�3�0��0�	P���Հ�y"IXB��<�v`�9Ř�б�P��ybގl۬���`T�0D��ِE��ېx&[�k���D�b3�8�A��(��B�ɍQ�������Ԣ�#+o�DB�	�uR�a�vkGA��i�.��D��C��?+
�-;�o�`S��Ṙ�JG��'�Q�P�<yU	����ɪFdՅ"Ɋ�(�NYu�<���~��`e�s�X��V�Eu�<qU�%�t�y���]!���@u�<	5��"��� /Q�r��t�<�e'��G���� ����RG�<�o[ <5��FޜC �y�I�B�<i�N�w;,M��.^�_�|٦,�g�<��ҽ[�~�����){�(����J�<��aJ� *8zS��y*̠��H�<�K6q��	ZW�*@�r*�lA�<) P36��A&6|��zy��'ܐ9r�V�6Y�cn%+ĩ	�'st�Q�O)�K�$hPi#p"R�<Q�E�!hz��W�Z;�%���hB�]�� @�@�vL�af�>��C�ɚ5}�A�CװNP�!��P� U��'4��JN�,�r���dU>H��
�'�
�ؠ�S
:lz'ě�8)>(b�'�VYru%�,&yBW�3�$��'۲�9�dvނ��'إ'mb�I
�'Ö�R�� ���E���4j�2��I�̊��)�S�7�~����U:P�
�c�%�3r\B�I�l׌�p%�Vv�)���?u6��'��$2����yuB[�����V�	4�)��'��I1�� ������ri.�#׍^���R�<o�b�'�Q>5*W`L#��H�b���ۤ./��Y�ɺ���>�K�<��U��#@x�[I�'�y�F�)�<@M]�{��ڃdA����j�'ט ��r�a>�S`L*k�|`S�%�~��4�ȓY�&���C��{6�͛s+�����y���9E�DBx�'���b="��h�4���~��h��If?1��ze�\�s*�0?�̃Ǝ9�Jh#�{��N��<�p_���k�m_�V���NYP�'�ў�B
����8U�����Ҿ&�<S	�'1DXd�;�T�95��
H<�0�����XD��[�q�P5X'I��D5��x%f՟�yR�@/=^T!P'	2CԁC��H��d"�S�O��Th@dX^kc�U�R0���
�'��|��J��'��0�IK�D	��'8�PvÃ�\�l�P�1P�*@��'�(��� �^��Ń����P�R�'S�1���z+(=P���#�ny���>�H8�D��TtA`��Y2:\���"O�1���
9H�����P�3��h+��'�ў"~��h�  �#N,�y����y"B�jo4���'��U�7�yrN
�$���ꣀ�<g���׊���y��Y�X�h����W$@�U�L��y�@=��)�⁯M�P�x�lɃ�yr��%J�+�+C� ��!�P
�y� Ś-�����? y�F�?�yr�Ҩ?�>h��CI�14�!�yBLZ�n��0����F]h�h�yr�Z0C� ��M�?/�n��.��y�אd �hW�	8,lv}�b�K��y�m�/���b��2��W�+�y�P"/�������b��(����y���C��(E�Q�l�.��受�y҆Q8Snrk2�!:���9����y�Ҳ��(S��˛,�\����,�yr��*s��Y[�, R�^<�$N��yR�/:��j%JO�:����m��y�
K�w�b����,��h5A��y�[<J6���@ ;,snI�q�(�y�,G9&����C�(_t��>�⤇���" �ЍT)H$i��Y�pم�`(�e�Tk���ȁIO�2��<�ȓu�b��w��4r4�R���v����g�qP6�"`:��@���
;�h�ȓ"�*E+Ո�%g�FABQl�7Q�vy��zQ�u�āԙ5M�ui��B�et��g��*�D�n�F�ag.)�.�ȓm܈RțQ�>����Ndq�܆ȓ�҄�!�̩Mæ]r7#Ă*��؆ȓ �<�y�.�0zs;Sت��&��Բ��T��Q����~�T�ȓ8;�H�c���N��	- �X�ȓt�`#���#���ˋ�C��ȓ0��OJ�*+�ͺ{���)�"O.�!�A�9���C����@X��e��[��'�Ȕ��X�
�Q+<m����'f��!���� .)�mKP�d�<A��E�N�kv`˰D��|S�L�`�<9��ǉ.Hp�q�3m���d�_�<I�`��xM ��m�1>�������V�<Qr��~.F-)�I� JT\	���u�<!򨇇8 �P`VMW�"�Ƭ�&��v�<)�"�6,>œ�H
�6��E�n�<� �m�Ꜽ"����[�y"Op2��V��c[�7�ZT��"O���pB�F"��3b]9�"O YȄ�F�e�2���_,���P"O�@6٢^?`�n�0U��-�"OnQ0����-E�*Ha�A"O��f]NC�PC�j�Q�w"O|D(��<�f�0�»D�"�y�"OHa��K�%%��ԀXn���""O�i�/38$Q�e�آ��"OI�1��2c��2��(�P]��"OL��BO���$Y@��R34$P"O�Piĩ��H;0�KY�����N��y�m��<R�׈	 5��2�yR�.:�9 �f@~֬�؆JK��y�$bq�]�EA���3g�L��y��k���ؕo�
E���v_��y�mW�
|�)���#"�xs��%�yB
��{e�B��<��D����y�/Ƨ]3r��QȄ�B:���k��yr,���z����5�����	l?D��K�+T���'��l����9D����Oĵ�����䎐;�v�"ԅ7D�p� �ۿHA~�I�>X�bQ(��+D��k �U�3v0��T�?�D�0� )D��b���E\���� ��%w
�Sh(D�����"/�b�"!�36�VuHу<D���d��<����a�J�.���&=D��9E������0m����M8D��k����V�Y�]�ܩ�Q�8D�ls7�ܓx��;�)�*	���Z"(D�xr��ƅno0d�"*�4F�@!*D�4��(n��
0g�:�L��m?D���5��T��P!��aj:X[!�Ō88<�TJ��@p~pa��U�x!��R�T�󆁡moDP�F_�r�!�O'HW�����U�`��1S��EE�!�^?A'
x�$�а^����c�/:}!�D� �ʬ�r��:9봉� ���h!����ع*��_׾=�3BK�w8!�ߌp�D%�!m��7�8r'ؐ!��d�4�����-6D�	׍S��	$)Hd�1��Q��H�Ӄ��<2���S&�ZB��<`�J�!R〨 4��Ga��7�J�'@l#a.�'hnay�Y�[߮p# #Nf��L4�	��0?��$�'ʤ�Z���<8�󤉁-=d\`f
�'��B�Ib�
�@� $�,m��d���R#>�L_��40��3�ӡ4��Sr/��L�>%j����N�C�	�+;T4r��Z�g8�0A&Z-(>�ɣE|�5��ƒ�f�S�O�\��0�a��Mpd͉�V89��'�����.�8��ǇAy
�@�O
�I@	N�� �	�^\(;�	I(6wH�r���)��	�z���� X&���  ��PsKM��Py:
O�d�5A �A����EV�Z�`���I�n�6 p��~�q��4#2)a���ί$v��2H��y�ϓ�
�%��[օ)uV+�yr@�nF�\��!X��S!�ީ��Y._{\'-��1�C�	��I��G�%�>y��Զ,���'J�mn��Qٰ��$����\""���+� $4da��̮ �	�+>w���4�0+�p���Qh<y�ܔ��Ԙ���<R̨c��U�<)R�@��EyS"S"98����h�<	7C�'U�P��&aNP0���_�<���Ȼd�T�
��Z����M8��id��*a1O� �u�7I�[�x�@�� �$TF�+�"Oh�3 \P�����fJ8u釚��ӡQȐt&�"|�aǫg�T��&/�5L�h2cGg�<�����S|�@L�)�`*�"�ҁWU�@U����'/>��g�'�K��@Kivt���)<+��I;^���p� �F�*�_������OV"L��� �.��G���
	��C�ĸ�Nޑ1����wW]�a�?��K�O�^�Yg��%oUc�<���.A��%P�RJt�t0�
�0q�!�$�* �R��m�&o�4�)ROB�*�ʴB�j�zݼu�֫��'�.���� ���I�]��9T�W�=����3D���Bɶ:� �)��:z���nۏo(�x�S��$�bd�'�X���	Q.B�8��04��C�HӥIs����ۿw�,a���]R&V�B@hA՜�S%	���q��X+�d�4�¸z ��>c&��Q"�0GT�(0����*d.�Y����~�@(������?t���l܉.�<�3 dI��y��ߚbq�$��G%0���p �U~���y��M�#�zD*��#�������� �hXWbPz�t�2 8D��!�N�B���:��e��eP��Bc��	t�
,P�$Y�h�t�,�i+�>�X��L�J�Аǝ� ?�����9��q�Uߟ��:w���i�h�V( 1���I?KkB�[�h
Yx�<3$���y~������1\�r��)��Q+r$A��&��l��cE�n��R?�
��G3=`0)�&^'^ز�`&D�t S�5d	r����P�C4�3E.K1�Nx�ǩ_=5
�Á=V�d0��ik�����	:hh1Ӑ�ҥ=�)"m4D��k��CryӠ'�pE 
�$��T�ᑤ�4p|9WD�!CFZ��U�HO��XuĚ 7w���H�)Mk�I��'�n��tƘ���XU$�0����b٠SM��"���-JvH��	�J.�����~���#W�7,`8HƏ4h���x�v�[�$�{u��.2hL�P�ޖj��S?
�&�Q���
��1+��� �
�'��}cu�

�n99��U��r}xb��5Sm�@�p���RZRU:mօ%��|j�w��<g��	$��'mY��F8C
�'�4��X�w�h���Q#z���Zb�S��Bl
:m�L���葽d�L1��,&ő��B��Q�Ze�9�M?O����f'�O�q�T͝�79n5k��_K�,�7��u�tH5���
�͑�h��z����=K6�(@hƬP���YEa��UXQ��K�E�<N:�0���Q���IU�?�Y'[,LnP�Cf��1_��(D�0��D��#_������;Wj���"��ٲ�ŷ+m�	�r�>E�d��M���2 JX*/m:-SR��#�y�ę�^��%���n�ZT.M���	�:8��u�P5ax�!h�4��d��o�akdK˒�p?��D�E��%h`��;Jr�m�eb��|8W�� c:C��l��"7���k+B[�I.db:�>�� *t4��b4��^��M�� �36���CE�c��C�?�0�ŭ�3Y�-Y�
 :'@���(l���J�hH3U�S�Os��au���t+��)�@ !,��'����d�o��b�)��u/p�yO�$�����V�R�"��'z.m����9���	D-[�u�Н��3��H�c;���;�a�Ow��h2��{��{�O�l{�D���<qs��&�jD�clU=o~�ʅ%�h�'�<P�1��qy�e�6�|e" '@�c�t�aC>���EK��p ��L��$l�:���p���K~XG{r,S�@"{�mC�k�"&>5K�C�jՉ��Q�Z��H�s*O]�E�R$�4���AX�5U� D�i�lY���v�8���
!�H"nZ,	88�s�*�La���T�s@NB��7R�L͸2�]�ͪen��^�\l;��'�V��Q-Y�a�UM�~Fz"��>X`�@R��j� 
���=�p>1�H�e�.h�0�
����vm٘UFR�h�^z������lՔ��d��t,����0	��5*�j���Q��,?&��#�,�P��UU/����)G�Jx����9h����ׁl�!�ğ%,�@�!Q��.� ��\�u���I���I����B�?ҧ�yG�:$+�q+��:o� 	� gD>�y"�@�	�xI�ஓ:9���OFK�������,�� c��p��\w�"`�ui�J� �$����E�6St8��� O�&���+,\O� �W S2J���R�oJ�_�t�j�⁌A�i�f�
A�4<2�-�*� aDY�i���(�#,O� 4�J�*��\�h�ŬY���!�č�@�n�@"AְQ-ආk*b2���Ȗ�"`	�]�O+�9���F�Q墌���wY�C≙O>-Iƈ�-]�杢��>!�ΰ�1dR�`�N�u�ߪ���+��LD*6�,��	�*�y�皁EƸ,3�"$J���I2�A��y�kZ� ���;�ˆ9_L�+��*���m��| t� "gJ
{)���EW4>(e��"��'x��$��`E�J>�B"<v=�eJ"\O�D/OH`�*��Ն�~L1&镇A�:�"�LB�F���F4f�Ne(�ïq�2�ׄO��ay2	U��&�@�<4���\�k�48ێ{b�T4s�E��Mv�L-�eA��~�DU[�!7J�� 8�A	R����d�ZK�A	q����xr��0U�Hթ�#�%��
A���k%m�i0�a�J* !�P���T�@ٹN?9R 1��`W�ͫAQ�c	���"O�[�h��V�"6"��{���ё���}C���g$~�j��M�N!��D�)��2/(�$�G	�("�4A��	�}��b�N��N�YgN�-1��$U�(��tҶ�w�<�
�a0�O�
��T5L��Ɉu'I�!p|!8��I�=���� e1d�A�����,����pݭ,��BD�L �y"�Q�|����P唹$�Z��ЏZ�yB�Y�VH�SR�9���0wgf�x�a��n�d@�CA/'�bC�ɻm��DӲ#%hHCܿlH�Ol@c�?��<9ń�24^ΑJe&�Fpv�G˚e�<9i�B�zm���� 
�T���b�a�<�PB�.$z(1c���!ZT�cNG�<	��g&1��� W�T#��I|�<)ajG$?��l��$��$h����{�<I6B�%��Hx�NW5�ZӯM^�<!�
�"H�v5"%�
��Y���Y�<� �f��Ss��	$�� �@2T�,����)�]b�='�Vh:�(,D���$\�\�r�U�wY�0�,D��E��n�� A<_E�铴�*D�� ��G�7rfe��&Y��-E`"D��ѣϻf>�\a��+g���&�#D�Dv�oO4��`+��S�.ah�%D�$"H�Xm��&J�0wkD)�F D�`�b�B����6lm:��$D��x%=	��<��j��69�B�$D��:C��f-��9���q�A��9D�CG����(%L�<"���� 6D�4�%�[�j)�I��&qI�4(!D��sQn�,a3ĀP@�\�H�Z��l5D�����5-���+ �I+�o0D�A��O�pnŃa�ٔ/�f�r1�+D��H"fZ�'�%���>�:���k'D�P�ra �I�`tA"��]��m���.D���D.S���G�D+m�t���/D�X��ቁa< ��@VN)���!D��:�H�G�L��S���q�X�S�H"D�0(d#�e�郡��a�����L#D��#щ��~ċdMߢ��I�C�!D���mZ�A@��<��-��<D�le�S�A�3A��`��l�`o;D��He�.P��E;c�V���B�;D�ఇN� �̉Ai�
k��p�9D��І��("��{�m�=w}�@�6D�p �
T�Lu��)Q7e���7�7D��[ �mF2�`��(w�e��6D��;��]м{�Q�I��G�2D�`x���qO��4��&Vv�)�0M"D���h��?��E�e"�)FL~�sT�!D��G�6ޥc�I��;�N%s��-D�LS��1C�\��*j�����<D�ӥ� �Qj�@�Ɯ�Τ��A1D���H��aU� S\�h1�i,D�Pa�V/ R��)�/�ؒ1c�L!�� h�rC��B�hU�$,W�l`$&"O�尃0%�ݨ�̗��$()�"Ol�)v�-k�Fh�u+�T�|�` "O:���K'T�8�@D�5�hY�$"O�I��Z�iԦ)#�כC�r��""OZ��Ĩ)�~����:�R��q"Ob�q+�)�Պ��ʤ`�^��"OHp ��\��1���'.���"�"ON��##�o�^ �����.1!�"OK��NXR0��œ|g����D��y��ez|��$�$!�"\Q1��y"��/jl%*0/��r��V��yBW=�&��@��. ����yb�˄G���a(<i��yWl���yrJ)%G��+d ����#f̍��y�!�5�<ㄩJ��Y26%�	�y2��0�H�J!��.�}!���=�y2�=��0o��W5�qz�)��y����k�����_	G4ب$���y2��S���D�AiJ�iE:�y�(�;>|����8C�t�����yR�ް;�u�7bV?
�L��w����y��U/z6iɧ`�} iS��L=�yB��}����� �~K2<a���=�y2kˮd|";�ԇv��!�Ť�y�%F�N��Ȅ�X?Ѱ�Kd,މ�y­�>JR�XW�+h�K�G�:�yR�Z�j�Dyj�E�1K���EBý�yR��5�1)�"_&�S5N�y�j�6�T�3 Ă�T�p�ā�yrfQ7`�v����Z�p��T��y�oW�-��@���>1`siƗ�yB�X�um>ݑQ�\�A�fۓCЇ�ymJ=o1��{P���	U�u��5�yrʂ�M�$�%: �2�_o�<�0�Т[��Y�Tj�g}���C��q�<��!�9=��`�N
?��,zg�e�<��C�y �`�g9'�J�Ȧbg�<�mG�vF���94F 6bGb�< (ls`c3�ˢ$�Jh�`�e�<Yd�?r4\�G�X�O�X��+Sd�<	�aϭ`�h�ƙ�SB`�5��K�<��jT)w\A�fÊ,*YT/�K�<�a�܋�2i��h*
�59���D�<���S"�Nᑅ,%v���H�A�A�<��o���3����
����V}�/5.T �=E�T�đWzF�{��<����J�y�j��AZ��JuKѳ����F[���ɢf4$+Ao�vX����fث}]�c�Ѯ1���X�$�O`��"_<7�ސ�;�"q�ݠ�sfB���PxrC9q��k�a�x�-rQl���Oj���4xE<����k�84����Th�$�K�LE��y��!%���"Z�~
�ɇä�yr	�E$�U��@Z���9-G\���-\6'd<�Q�ڰ��C�	�DK,D��Wc6(C"�D ����D0v�׷%�D����
P�@t2���m� pfl�+�a~�lE�H�N������]��H��ҹqB��ҦT4T����xl0A�S�ʃU*��a !�+d">F|"�',~~}9���|ܧdɦ]IFFK,H_�!CE��\��u��}��4K�o�cin �d ~�t���,a���K$�ӧ��м�Q�J#xԤ��F�E�^��"O(%�s��3h���i�ESD�p��%�>Q��'6���˓:j����b��2vL>����I!pp�2 @C*����f�H�aA�mH;��� l�C��3)$�M�u'
�Hڦ�	Q"O��rQ�r�`����`��h*2"O��Z��W�zBХ�P���6�ֹ2�"O|;U��C(t�Dp�ƍ�'m
���KPy̓F@|$�3��<k��5�#��p�ȓ ��)�TH�JT���r�ã<.0��'�����E��Fxɧ�4�6�� *,Q1�M:;m@q�"O��1Q$�=j4�2 �E2:#�E�r�ߟس� �(�^0�C"�%)B��I%�:Ց��R�M��Y�i��`����B�M���P$� W�~�3�쁡:Y�8	����N��pe��?7����7w�>�A�BնF��"��(H�TH���(l�Li����k��9�e���EJ�+>��/��y�F�1���y�/�29�P �d-X�K��J�EЃs��	�H"Nӌ]ۄm +[ =(���O�|�� !P��e�#�U\iaV"Od�����4���N���e(��V�>������4�����\�G����������kb�G�N�.5�6s��{BO��T��Pc�
���	+7+�Z��q����}|�)��v��D��	�v�p����g�$RWGG;X����@wk�-���4-ǯ:�4Y���4�F� {��ߠi�Q��!�6�y��	0�������!dK�=�Pd���ԸP��ʪ\�j���
D���*%!7@|Q3���	j<B,'D����I
oǨ��(�%h��S���+o���lڭ-�H�Y�:dɈ�i1����	�ɗbV��4��6�B���ɤH��V"�̟8��[&-R�Y��"S�����ɁRߴq�b��ux��r��:��X��G���:��x�\#t%^�"u(��G�1�h��Q?�Ȅ���qM� �����f;D��Hq�v����v��"jà(9bN��/��0'̿l��8��L�&�L�X��	d�%�O��v�+e�6,� ��G���y�NP�R��2$mc�m��	����Ġ�,S�D�q�6'ظ1���O	^"=16���@����G�V�P��
ZC��̈��}��)��E�*�"t��
-Rx�CͶ
�H!s���E{����'�R�QR
/0���S��8�RJ��r� �tA¢�v��0�J�@���κ�{5��X�I�Ο�y2iLFZD�𨖱�p`bunQ�V�ʤ���D�	�n���$S�Ju),ʧ�y��fF驵��ch�S$����y2�;G "Wʁ�y��[�kȟԆi�s���q�@a��ٹd���!��;E
#=y����P��D�&MΠ2��PK�0y2�ՈN�^,q��δA]b���U�k��bƭ�/8�\��#KZ����^��MS�D'Fdā��IAB�<i0dD_��Uk��ĦDf���'�)j�NG0:���!ÂAʷÜE�<I��]�6�$� �[zl����F?��a�"4��� 3}��I�$N����Ʉ�\�E #j�'6�!����`�I�3i�RXY ����f�&��r��#(���F+~�q�䍎1�DZ� F9��~r�N"�^��@c�'>a�f�'L�Np�֊��	3l���r4� �����~�iҫ_�I��aE}���	gvR��J�Z�'9�T%�w���"�p�� N
�B6��$����2\5Wt��wf�;Zּh��䦙�㌌�0w�ӧh��A�p�P8#��Y3Ã�P�<�`0"Ona�%X�][���Pb��g�*P+��>��D� �fM�v=O��
T��;�a��(�|^��!�'!�YIEʆ5�JI���6E۔q���&�6|H�
O�Rf�Ǻ�X8hd�:
������=�z$s��	�v+��gH;"�T�P���!�d��w�j����N,���L��!�fݸ��I�8"
-X���5~�!�� B�����:@pr�K�?V�!��s-�LZ��N6$�P�H-b!�Ɍ Z69 ��D4̽H��H,h!�D�)s����i��(��	%��<W�!�$���I1֡�V5�}I5��!�0��%�� �s��s��!!��	�:C��!���cw�$����*w�!�d:8��6ȗ�_m�p�%I��z.r����Pܓ�h��� ZD1�Řa=�t*����	z"OX�Y�"�_���i�N�����iJ^X(��\:8r�&���JW�usb>���mTK�A9!f����B1��K���Iu�6?�\��2O��2!�@Obt:d�G6s�!q�W�RbC�a8���PO),O��P�o�s]��s�Ŝ�0�;���X����&���'$�k��ˈ �*`ܠR���0Q��u+�5�B���͐x⧔�O����dhۛ���q'��tR�������37$�*QiUu�}�'jF�g>M3qiM�d�
e�6LظmEBC��95����'�`_Z�Y�!�,�C�i��	�,J�9H�	�f��5�䘖��禑�B�Q�	r`�Ҩ�h�|u*`d3\O� Rg�["Y�ɜ'	E��^0R���v��6Rr(<1�O��zFG�^N���c�'g*)Z�"�g�D�+2O��Hv�{F�%1��y3�QR�Ӥ<��#���+(��s�O�&!F �e$S!l��ĩ
�'�X|�QE���	�U�I����nS��I���'݋>��R�4�*��t�T�e9�I���W�nl�E8�"O452��y_hA�F�g�2=���i@�	cO#�a}��(蜱�O�K��2��}�����A/2<�	���P�QE �Ty2G�B�,B�ɯ+��XS�$/����`�j�B䉿C ��ѣY/ml�u���򄆕2��b����"&t�qC���>v!�C��4��%N(6@�^�dz!��j> ��IN�W(�Qr�cZ'F!�$�8�\=�Q�ʉ*���C�	�!���.l��T��]%���sKO�R�!�W$L��8 ��P�u-*�Q�T'�!�ė�DpN1#��
C���H�f�!�$ѓ=��,���RN���GI<`�!�ʯE�~���T�,&�!SA㞊x!�
�	QFmB���#�l��B�=FI!�$�La�\�6-N!\)N���0b%!�$�|��#��٪D�ؽ�7��<�!�D��#-x� ��r�*�Äb�-@�!�J^*!�\$s�Z��oް\�!�d�5n�M ���"@�Rl�#�R�w�!�ć�Q�,R��>v�u�n[�2|!�$G�h&N"�Ȁ 5{䐃���~f!��[N+�X0C�������ˑ�{!���o�X �A�Z��$�Ѫ��gS!�d͋��@�h�T��I(PC^8YV!���i���a�+�[���@3!��z��8CH��H\�1��3c�!�D�{50A�rMԏ]Vh �`Ȓ|u!�$D�KT��h��_�?��B��[i!���|��("C�7(z`1���
+$!�dX6Q�B��sր&����C�!!�ֻT�~y������c'�(sc!�d�Ǌ���A�:U�.<c��L<mg!�Ę�T*7N�7}������x!�$յP��gH��#~(tC%��Xk!�$	$;���4D�
!,��!dܫ3!!��2�Mr� �LA�͚�!�$�a깩S�b
�h�BK�!�$^�>B�R-�����@K�@g!�.,�����m��ht+��Q��!��"�铧��_b��j��ݜv}!����x�;�f�D��-��,v!�d :���u�X�olJ|�1�A?R!�dć��-�CX����� ~V!�1Wfy����0NF�j�Q�;B!�[D@�������7-��I�!�;bi!�dϻ6=��`Ā�`	ʴ�L9R!�D���nDa�(«-oH��a���Y!�d0ֽʒ\K�0��9S���x�8f�a~
� PQ��*՝4ąV�]�a��Ex�"O��ӕ�լ�wJ@!U�@ �B"O%��O)B�j�t
�-�,�"O�)����>f�`9���t���"OjxN�2d��Y��3\���*�"Oj%"
�(�x��&êK�H�`"O��z��#RV����%��$F�(3"OTE)E�OL��@�J	�� ��"OF�B�\7w'f�X�Q�D���x5"O$IB��ǦkV|3eG��<{|Ēf"OF	�Ϣ&�(;7�)zy�x��"O�)���֖��R��L	S��p�"O̸��GX���n�2[��s"O�L5�U$d�Є�&��)��ZB�'i�A�֩�@�$ӵk���I_��}�U�Ը|X�A�a����S3i����вS�}a7�ʆ,�.�6�K�)'� �Ҁe�ş�ݶB�D�ƸLWRh� �9�vh#4�xb��d��y�L'�Z٘bj2U;N4R'�Ǥq4����͟$[�4�y"��� ^~ם�ӈ����O�	V�@�H���2
�D#!�Џ��Ղ:~�,x�����Ob�q ^*,QY�`�8��eK�OPe�p���:�E�ş�"}jcФ�"ѱ�d�$	
�:Q����:w���4�>E�d��/s�M[w�2���qd���>����"��4u��Q|���OW�D���B¾. ��$IV�@�!�2����'pL�{yA���O�������N����M����'.�p��$�<i�0�_��}��h-[TI!���6���{2 �|�<���D�>l���b�=YĶ��ȓ.)�0rF,O0�Y
'�ٝ!1�u�ȓ�$0p#�G�J��D�$Ohm����0�چ�jخ����J�Τ��`춨��@��f��� 0AK�y�ЅȓD�b��#���5���F�����ȓ
��˄>u�N�`k�*C����ȓ-V��x�n㕓��A��e"O�u�T-W&Y��5o;�h8"O�!Kk�0��0	��0"/�i�*O��I>�t;�c������'g2��Um�}#ZXぇV�ssJHc�'�čaR`Ѱ�FY`���4< �[�'��@yCω�p�a��6.T���'�t�ئ�H�/�RT+&_8-�~Q�'0�$�Z�_E��kU'�	�X8
�'s$���p��1��Lu��
�'�U��R�S�4�6��.l
�'_�����!'�{S�;M|�y�
�'Ě�83(��L\R��"s��0�' qˠ��gB�yC���j����'�hx�f^�w(B����1c�԰��'G�U"�@ڰ&.`;�E�S����'C� ���őg`9ȐK��E��'�h9�^�X` ��J�rp���Qc�<ɷ%ho��s�j��EW�<�Mʼ^V0 Ӷ���pt��O�<Aw�(��(�ܨ;��u��[G�<ٕ��S!}��"�-�D��,�C�<1�m-7�5�!A$��w��@�<1�dX�mJ@����"=�Z�W.Yy�<���#k��k�v�4Ǩ�J�<�a˕v∅��[ �F�*�n�G�<91ʅY��X �i �>H	�� �o�<��� �z�b �eE�$j��u)"I��<���R��Ep��#	� �cs�c�<�5!W�DԮ�7eƥU��p#G�Wa�<1��G� �!U���K^�@��[Y�<I@پ�<��em%%���ZqZ!�� X��b�V!���52P��S�"O�SR�^�7.�8��Gw'vY��"O�Q��ƈf�
����;
");�"O���E�*`���4FD.�윩�"O4M``KәO'P�!&��3c����"Ol`qf�����9���d\I
�"O�)��'XƦ	q�3Pn�}j`"O��q�ߞ3o ��Aa�\Apu�W"OeIh���<I���m]�9��"O��+&nG"G���y�F�T��"OVXi��u���pd�D=�b��e"O�\)e匂g�4��D|�L]�3"OH0[�dЄX+��:P��4���U"OR�9�X[�Xhrd� G����"OrH�hT)zLm�u�S$T�B�"Oز�n?J�F	 ' �\�b�"O����"�A�4�Z�!=~���"OBL1���4����Đ
/2=�'"Oi;`��	l�Ҳ�I�H��"OZt2�J�W�t'���z���!�"O��Wcʊk-�-�F��vZd ˓"O�aK�B�p�|�#%5YG���T"O��A�'7���:B	и6��A�"OԚGh��^���#�� <��	��*O��Kp�h�6��Ƭ��m}���'(iIw �&Qt�j��eB�`��'�f@�%��-�p�u��S>H��TW����yI�Ă�W�1�܄ȓB�dC���h[ԑ��͚;L�x������[)���^8<�f���`��HynH"�r��X1�<�e"O���􂓋D�e�@�{n�!�"O^����+�vQ����8X��1T"O*�֦Ȇ|����$�;�@˰"OT��e�ѡ?|0���^:%4Ҽ�"O�M�`�|Vٻ#�	 ��9Q"O����D�!mj*�d�#qR�*�"O���@�ӛ%�!���
^�D�#"O���jN�mN�"Sd����\�"O���cC!�0y��b�y��1�"O�-�@�n���!���R��"O~i"�'��M(A�����^0Y"O���C�R=I��\a� �g���!"OT��4D�+/
���iZ3g["O�q4Jʐ!�\�1�κ�X��c"OD����A�! �@���"O�Ia@yj@�� ��f.�L�s"O�m�"m��gw��e@6BD�s"O"�:凘�%��/�6/��k"O��`�h�(k�vI��J�,��`"O�|�n�	|��Ǥ�3ks��f"O�Q�%OA)pf1K��$����"O�����0�����4}S�1r�"O���Q@��7NHHgDoL��0"O� �N3S"�L�#�.-x̸�"Or��W-�.c��*dC�<2(X܋�"ODyc�/R!7vTz���'z&���t"OP���D)_@2�c�@\�S� T�"Ox@Qa�4%���Ʉ���8t�G"O�y�� ��ψ��t Y1V�(93"O�h��.d'}r0O^�P:ʥp�"O�,p�ψ!V����Ӕ+�R�E"O��פ��Z�jQɑ��%,��"O�q�� 8�v�8��4#H)��"O� �YSW�Pw�v	�AX;5�8�`"O��;��O�:jE�d.�~��$��"O�t���>P���L��L�\�r"O<`�X"iY�X��J�=ip�"O��x��&l�� ۧ	�|:���"Op�O�9��]��F�:�ҵ"O���V�2E��0CK�x#ơ �"O~� �+�� ��x!u�D�JE��"O����B~�lB4�,=��Z4"O��DZ�+F���A�ųv�~��2"O����&AL�8c@I�!&��9I1"OX��4��6i������7�����"O�p�m	����AjK�Q��"OJ��coD�#�f����)+>nMF"Ony�`�b��h��ɹz+hA+�"O�(�c�H��Y�C��!b\��"O��)+ɤQ�� �	R$�����"Od�挏�dB�`�X�q��8�"OZCO��K�d���n�f���+5"O�k�*�H�R5��c�Ȱ�E"O
��C����ɐp�3z��a"O4��4`��$]����+�!_żA"O�9��)N�f�r J�[�q��"Ol �d�P[V ��Ɨ8sZ����"Od���'N;2�i��Ȃ�4�d]3�"O�Z�%ƍN1`H�v��V� ���"O6��n>K������=Ȁ�C"O�J�BY*W��K��3E��#4"O�I'�	'l���E9[� ��"O�mѶ*�jfUS���B�"O�����)�ۦi	
ead� 5"O� �+�ּ�+�57_*�I�"O��S��^�:���@�	%#\B9:"Od8�v쌵0�z� �&eIRq�"O\��eч�\�p�Ň
P���"O($�b��B�F|�dg$su"OF=��DK�1���# �Z�6�Ұ�U"Or1����23�d�{�D-����R"O~�ѓ�t��� ��d|�U�6"O�,��&�K�`e/�Bl���o�!���5V���d�Z ]Jj(y�f΋ !�7n���@1#7	C��R�C�K!!��O�$(z�H��-/������'�!��9l�\$���8~B�cD��y�!򄈯E8v-yÅ�$8��P$�ݺ$v!�D_bqAba�j�� �O�"!�N�,M��s �=�����2�!�$�j9���P�K�H'�E�e���H�!�d|���Z�f?��S*U�j�!�$N:n̪dy��	;�uH�X/_!��a���0��Z\�+6�G� `!��QdRR�&BR�`�P=�%���w�!�D�9�(`���\�d��OZ5�!�D��C���Y���a�Q�G$ՈSy!��S����
AjP�pȴB\� ;!�4%�,����Ɔ�5���ˉX!�d9�^��Tň�{��xVϕI
!��M��P�0�M�[���i����!�A-2I�	�݃,�R���(˙�!��oY��#E !z�A)CHL�w�!�
��2�[7�[�4zdȐg ,�!� Rfb=x��|� ���hL�p�!��(mfI;�N�Z �p�bGW!�D�Q�C �Շ,=�Ց�$�6B�!�� ~���h�GJ$<�Wb�4V<��{"Of�0�旤r��hXt`��'���"O���'#�-Y���ZQ��,yzݳ"O*��VoPbVF%qeU�<�B ��"O,x�`��;Z���U���\$�yP"O�dZBAY>�tH�ry�6"O���ƕJ����T���_�5!"O���q\R��9�ț�g:P�"O����Q+	�tbČȲ1MLH�"O��FI@/}	p���'zX�� "O���Ac� qHh��+��$W��"O&�YE����f抧%�QyD�k�<�T)�2R������@�E��A�<q�aE?&>� m%)�4do�f�<	d ǭ��ʔ.ϫ,B�;��Xc�<yf��y+�c���vlM˰^�<q"#M���0z��$z�$aYA��W�<y+	�Q�J��@�і;�-IQJ�I�<��%�an(�)a
f?���$�\�<b�!�
�z���=����SY�<Q�]�1[F,��M������T�<iV*�e���c1M�Ue,P��NN�<��o�@�¬Y��>����o�<)tH�?E?� �㋒�|�<ͫ� �o�<�r�á
q��'���1rs��R�<��`�R��q�X8 ���%'�Q�<	ƭ�7=�|�g.{�.�ءN�I�<��h�*]R�m�'��!4gHC�<�4�
�����U[N�����W�<�Ʀ�7   ��   -  �  �  �  }*  >6  6B  gN  �Y  e  �p  �|  y�  ��  (�  ��  \�  ��  �  9�  }�  ��  �  E�  ��  �  ��  R�  ��  @ � � 9 � �! /( �/ �9 n@ (G �O :W �] <d �j �l  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o7�!Dy�'�L�{�5� p��*кKDX��������8�\�`UBY����Z�h�X�!��oV�y��:�Z��B�%;�!��3$y�TΑ#9LȺD�\1!��	�e���N�dK�ٚA�H8%!�dI.k�e����&,�բ�0!�d@��!���&�fH+I g!�D͋�@�BB�/Y��$��,3!�\
F���+��UN�R#n��V��-�O>԰�H�4U#��C�N��i�B�J�"O,P3�nx�Е ���i�\it"O�$�P���t���4���5"O̤ �&^�$��	�3dD2����"Of�:CH�3K�t�b�����#�"O\����9+Ϛ����@�6�it"Ot���,EMcx񱡡S���8�"Ot��	��K�8-3�ݣ.��i�"O�PAa�;���!aE3rE(�0f^�������L�Ƅ�f��>\�Rrǫ˸C�I��
 �A�K������'F�F�bc���!�X��s��9�����6S���u�'�qO��	dA�i:aB�C~
�s�	(e^���p�4�⌘��h̊"���C�B�:Q�,��Kð=i�����[%M?@��ȓ]V�Ӄ!��P�D�P8`���?�
�j��ү!�ʡ��C-p��r;�L5N�b�ǃ��uW~� �!>D��@B�~�%ic-͍"Sxx�6c�<Y���?a�'I ��n�R�����~A4H�'�$9٠�ޔ-l��t�Ή yVM[���=��eJBӑG^�#&럅n��3�"O� J�D�N�䕐tʔ�.J I�"O�iS`�,�f<x%D����s"O��hQ�T?C��c� �+[�M��"Oʁ�c�נު�P�/G�t����"O�� 	-i�rx�M�Р��2"O<XIaH�2/N�3-�)�vuY��OR�=E��e k)|J�L�i��Y�%զ�y�L�>)<�䃕�.���@���+�OJ4#eC �.6` Z#�F=.�*Oޠ����*��`Z�!@�m6d!�	�'�2U�Q�E�%4<�/��l鄐1
�'�t���B�zSBA� h669	�'����!J�� ��@��e��x�'6�aQ' �T��)B�g�>���'bxY2�X'm��8��[HH:�'�2s�-RM5@���D�:_nl�'�����ʟ!(Е3# #VC,�
�'D�)5�@CLB݃Ir}�	�'eb���ӓr�F�	Ո�4���0	�'��M�����|�qd�a��5�	�'�x���\�c�C�Y�F����'�,<��l� #�d3B��=Y
@	�'�l��ǆ7:�� �r�S�G��p�
�'6θ*��Ť,��x�����;�Н
�'�،�
� 9rAȝ�:�~�	�'H^�2@�/\|Q���(+��(h�'�&�£��3]6�0��
#b�P�U�6�S��?9ҮA.��pt`��9�6쳵͎k�<�"�)b~^��d#Ŋo�%Yg+g�<i��U?�������*Xp�� �\�<�6薰jJdI�Q�w�����WY�<9A�"jС���K��q�HT�<�M"m�b(�#��>z���B�ǂQ�<i�`Q�U���ǎƽ D�-ђ̘W�<��h��<ѐ5��:_��6�Z$�y�g��5y�pc�BM8|�H�8rH��yR	�;CE�Ѫ��֙{�,��.D1��=!�{�	�4*6�:�l��&�!m4�y�!\�){ ����A>�u`@GF8�yrcSv�"ìL*s�0��DL�y�!��T@!��*��XnP��W����� �)�矼҅�B7T�&$١%NY�� ի!D����NT5d�@)�Í͸~W���2<D�t�CbT�i�X� kQ<����©;D��h��J�m=l����J���8��%D���^K��ue7�X7$?D��zso�%4��<9�삚�080T)/D��a���iՠp�!��"¹2�3D�H0!�*UID��Q����h�6D��q!jK�4��q�����c����1D���墓#e �L ͌�K��1C#0D�P�Q'�t���颁��I,�(�G2D�8Ce�,9u�9 ���)4��(#D�x�3�,i�[�!� ���!D�,���/{b^���BG�c���Wf+D���TB�T�@P��.8�Py�E*D�����:R=�&��B��0�7�:D�p�]�sx����(¦�� �P:D�0"t"�>B�tx�1k��؜p��8D���$�	PG�f��?~X��#;D�P�@b�'p��z7hEBuT����8D���o\�F�
$!��C��~�I�K4D��iC�J�$��M�E�B��A*4D��a-�{`����,O%P�4�Fc1D�� l�2��U)Ij)�d&˧"��"5"OT�����pr%M�!6�p�0"O�� �(9߈�ԉdǦ�I%"Odl3�잋�����6X�J�QU"O�� ׈I=mr�@�M� �A	g"O�h�L�l6�A�8->D#�"Or`P�7olA�#���,a�&"O:hٲ˨-�(���<v�:\3A"OIHv�վNjZD�@O1d���iw"O��4"�F0�h)��W(9r�d(�"OE�C
)v��I���h``m�""Oteɇ�
 @^ą"VlXmn q�3"O���7��&;�R�*Ǳ��})�"O�����K� �	�f�A.n�80�V"O|QZ����ܘ���Gk�}[�"O0��A�K�&k���ef	�H�M3r"O���V$�7 !T,�q�Ɣ�D�I%"Oh���N#��x�eY�GFX\�t"O�X�!��DENJŕv��X�%"O❚�`S9�j@�ȏa$Uq"O�0���_�N�%I��`��@5"OYS �B�Rb��J1���:Y���Q"O��`
*������N=P@��"OP��w���*e�e�)�q`�"O�	Sٍ@��d �Ä�'TA{�"OT� ��ȥ=�$�#t,�N耀�d"O��3��r@�եo��Q�"O¹`��5�h�K$�>�"Q�"O�H��D�g]��Z��:؞!P�"O�����Y�K\��B��� �84"Ox�	�#$W��]+e �!�@)&"O���z8^`���B##�XA�,D����8�n�2��
kE���=D�8�I c2ܩ�������f�.D�L�!$�	x�2x��́۠}��-7D��iٶ�y[W.�;�V���5D�L��Ћ0+�ݨ3#?��q�5D�#%��������:Vi�4�B>D����T6o�y!�+�<g
t�ǧ;D��h"�m�� �+9򒨹3b9D���"�@+�:�#qV�?�@}k4H6D� 
`=�4�E��$��T
�/6D��{��ۀa��5�WԸE��PQ�7D�h ��ݒ
��zdD�2lKbx� #*D�X��=^�AJc��Jq`|Z��)D��HOT�]1LI�����V��v�%D��Qv�\69)rU�����60#��$D�Xr���	w"�z"���EB��D�"D���&)�w��� ��G�АC&D���C*S�
�y�T�-�`��W�7D�``q�o��i8��*Kj,hҫ:D����P�:�LѢ��W�J��N9D���"U<t����

;|��y�7D��{��x��e���]"el:D������]��5��j�*[��q�v�#D��0��3�T�`HXOGd��L&D� ���!	�Eyg�U,�(*%�7D����2w��H3�f��@b1C�!6D��S�W�Q"������ �)D�����$��9�+N�J�T�<�Ԍ̹~�b5iӂ2�@s���b�<yŭ�v�� P�e) &+6\�<��nZ+i��"L��q�����`�<�`�A[�V�� �)z�-�£Y�<� ���f��'U������ZF����"O�*a��!!0AY&�çN �"ON�;0d��fOd�)��@:;��f"OV}�aA,P�`�-�Tȉ�"O�l�D��. ��h�H �RT����'B�'��'��'/�'^��' �K�m�]����v,]�;�`��'��'��'|r�'��'�'��Y��U]�z�� *˛j>t4���'E��'���'}�'�b�'4�'��`X���C��{�o�"M'�){U�'�"�'���'l��'m��'-�'s^p�C�3�\�ʢ�ڻ8G��X3�'�2�'���'���'���'M��'�.T�b̨r����ri�.u�$�'6��'�B�'�2�'��'2�'8Z(�A�F�ـ�J�z�t�0`�'k��'���'���'�B�'H��'e���7���1X�
E�S�3FB��P�'�'�2�'��'�"�'L��'Pa
�mPaQ�)g蜛w�B�'"��'}��'���'��'}��',� Ä�ZP8�+�G�7]� d�'��'h�'���'�b�'��'�z��b��zxj�n�*hrt�t�'4R�'+��'���'�"�'Y��'�pP�T��D��A�.�P���U�'R�'���'b��'���'��'
`�BT45^�Xkg�:.`V�:b�'U2�'R�'��'��Lz�@���O.9YV��Vx�Q���֥W;�u����SyR�'��)�3?!p�i���qcJ�B?h�`C��x�  uᏌ���Wꦵ�?��<���P�ĈQ���H�g��9v����?�V�B4�Ms�O�S���H?ё�f��}�L���f�f0{!�ϟ4�'�>�J��M�\����V�v(l��`���M� ��K̓��O�&7=��,� a�~��,� ��$J\��*���O&�dm�D֧�OZ�Y#��i6�Č�t�(�ǋ��&��#��To�s�!��8R��=ͧ�?Y��J  e<d��A;"
��JT�<	*O"�O$mڅ��c��KׇA�B�b1	alP?z�^(��x�b��I��0�	�<	�OL���<>L4)`ԣ.B��a���X���2�>�*�`6�02��`���"��cV���O��8�43�ŖoyBZ�0�)��<у����P��X��1k�L\�<��i���O�-nZU��|r��q�x� 7�6�%3UID�<��?���G?�Cش���n>Y��?�\��L�1��L�s�G_�ޘhrn(��|Z)Ox�������E5~��Ӆ��J��󕚟���4>o�,�<A��� �>L�64�I�q8���@K�t��?����y����'�"ض^DΜ7d�'}`��	&l��[1�����V,Hh es��OΠJ��Y����/�;9*�0�ԋ)�l�����韸�'.�i�	��M�f���<��Աڐ:�V)(�L3��L�<���i��O�9O ���O��Ą���Ȱ�U�@�L2T+e_�!�-h�F�I�j)���4��џ���a]L ��XG� �d�#;P5�C$Hʦ!͓�?i)O"�S�O�P��g�?i�İ���+��9��ybhm��@����3۴��$z����:���@��K��`�'��	ʟ��i>���E�ަ��'E��<)j�!)�)\d�8rk��D������ў�SWy�'IB���	�����W�k�;�'��'!�7-1O��'O�Ha�G�;1�<x"hS��X�'�Hꓼ?����yb���'�"1�� ]$]����3��øo���+bȩ�ON�$���?�S�3���=-�1lڌ@D6@�AS.�j���O�˓�?�|r)O��m�,f����cd�=|�f�bu��(%z��E�yb�q��⟠b�OT�nڞ�] �o�
^X����f�N�2�4�?�vcޒ�M��O8���ۄ��K?�J��Ԉu��
�"5+����e���'���'���'���'�S�(�μ�e�4,�ss#PM�>��۴�*�����?�����'�?����y�%.�"e�a�8u���Y���p6��]$�b>5
�g�٦y͓zaV8@��7�1;3	#�̓�|��b��O�A�H>�*O���O��EӍM�6�0�JєD�I���OR�$�Or���<��i!��`��'���'ʨMJ�&�-C��HE��=+�Y����t}�,h�>0lZy�3�4A��>G�Z��f�5B24�x�7�M�
H�|*V��OdHy��@��l��X�9[�1�Ц� 2bN����?A���?����h��NƒhڡPfQ�f ��Ĕg�t�$��͊�Cy�m�N�杊&�HA��N7GXs��R<C���	��M�u�i��Zd�ƞ���$K� A��%R�`�ؐo�y`tb�g��E��U�|�W���P�	џ��I��D(���;^�YKF[�2̮��G�Iy©l�"exb��OL���O���J�䑑F���C�G@�<��iC"�94���'BX6�ئ�%�b>9S�!��T�,�KT�R�(}2�)qx��I��;?�dl��M�����7�����A���Ls@��O#�* �c*rʓ�?!��?�'�����9�fdEß�`��UĘ���VL�<�2FΟ���4��'98�~+��hj�`<m�!*�.	ر��3r�<Q����<<Q����Ԧ=͓K�8)�'I=LP8�I�y�'ax��s�{�? �qieD�-&]�:P)��&!F�370O����O��d�O��d�O��?�(���&=pX7ҩC�Z{d�ɟ���柄[ݴqO�E#)O0oZ{�	�`����J�`�mVhҷD�:�1I<��i_7=�L��q�hӊ�?%<�B�kP�o���Sb�B\��8���I�����D�Ox�D�O^�$H�c��oT�,�6�ɔ�*]h��D�O"˓G��f.��a�B�'"\>���h��S��,�အT�rU��*?)�[�T��Φ� M>�O=��d�E�����1RrʌP��9A ��E��~9�i>P@�'c��%��Z��S1ڴ鐕���f���cE���	�����֟b>M�'��6�ɾ4=H!B ��7'�\�P�;4��@���Oh���Ħ��?S��lڲi��ơ� ���CW؟NƢ,��4$ћFY�B�����<�F�B����Oy�bF8CD�Z@��5i��U0�JϏ�y�T�����p��ݟ��	�x�O�!1F�}���UoF�*��(1�u�(P����O����Oޓ���� צ��9�̨���wtpq��� ~-Z�4E4�F�=��[�j]�7h����`P�R�p8P�Ö�cr�;�
d��*�*6b!l�	Dy�'Z�Ď�-���Q�}	x��&L'x|��'mR�']�I��M+$�>�?���?�H+��Ix��Z=v`r�'fŬ��'n��l���bg�ȍ%��F�U"3R��8��� �Y�1>?Qq�ڷ9::@C.��2>"�d��?�T��#"�H��2Y��)�$-�?���?)��?q��9��̳WY�&
�]���h^ryQ���OEo�,4m�	��4���yG��x۲�I��'����W��y�Ek��ynZ��M�d "�M��O4C�ß���[P��))�JU.:��a-�&�2�O*��?���?���?y�����CȔ$FJ���$���DJ�(O��mڻV���������b��D�X@���q�T���۰D��8�[����4��H"����Qdb�Ҥ:W�9He��/Y]^I���+-�˓ �Tq�e��O��M>�-O�ea���3�z�$U��� #��<)��?��|�)O��lq����!�BeH3͵.��`�f�3qw���&�M��R!�>ჰi��7�NЦ�:$��>-~�;r��9�.��gn�=8މn�N~��?Y�y�ә9��O����?x�˗�ǥ_��	�&
� �y��'0R�'�r�'@�	ΡEZ��@%-P����)�I����O\����e9#�#bu�i�'qi�7ŖBF�0�ƍI�ڑ9�'1�$\ۦMp��|�2���M��O�(RO�#02�a���r���UH�);�(b��r�
�O���?!��?���R<�d��4r�Ձ`/C������?�)O�nZ�A�0���̟p�IL�l�#J����..�=Ir���ęi}rib�@o���|:�'a�\RV�
3���i�8����l��3�K�r�ܖ'��g؟�Yb�|"�ݥ=��3�cP�Т�s`�I+��'2�'����^���4���5At]:!�S�[2�r����ĞŦ��?�SS�8��4���zq�[�B�\�"oB�h���ihH7�Y*O�6-n�h�	R���0B�O
rȕ'/������o��ʲiƂ $�@�'R��`��ş��	矘�	G�4���T���⢣�32/٣G��t�7�L�]r�d�O��2�I�O�\oz�y`Ɂ@8���̉$*���B���M;R�i O�I�|�i�'հ6Md�ĨE�7i3RuX5�	f�ˁ%x�d��ՂW/�a��@yR�'R�N�`4��^�k�S�j�R�'�b�'y���MC�����$�O�	4bJ3H��2�a	�c�0ɻ�?�����dN��1�ݴ!'�'2��7C�/Z�����#	}ZH���OV�#!]����C�)��_��?YC��O��y�͉�w}����#)������O���O���Oģ}����&��"��/CҘ}�Fr�>���n��MBo��I��M��w� :$���D�,ɐ��H�'�h7M�ئ%S�47GF�:ݴ��ę�-6!���N�&�Bա]7"@pi��N�|��
 J*��<����?����?Y���?f�	2e�����3?�u���/���Ѧ	�g�ȟ�����$?��I9)�JH.D%����'L���Ț��$����4T!���Oz^d㨀^^��i6.�3ؒ��N��
��Q�|K�*�8���W�Gyb&�t�xP��k��4����_�	ៈ�	���|y��vӐi��O������0��U�U�%D[֯�O�\l�W��d4����M;S�i�z6����|�#��e89*�9p���� nc�4���%a��H�K~��;Ob6	�^+��R��L��?����?����?�����O���kȶN6����g��4�UIS�'���'?�7��jh�	�Op�o�M�\�X��EԱw��S��F�vC���M<���i��7M�b�z%�tӖ�I����%�U"U� ��k�a��H�h�)�x|ru�'�FU$�\�'��'���'1<�a��l��3���'T�I=�M���I�?����?�-��a���rph�,�R� 嗟��-Op��k�%��i��HX8�A-K�B�PA $2���Ȳǂ�O��
�m��L2˓�Jë�OT0�N>Im�e׾%� C��J3�y&OO��?����?���?�|j-O�o�}&U�1/B;J�B�C��˽@�r�y�O�埰����M����>¾iĢ;D�Ϝ|�D�&޽-�*4�JzӞ�m�>V�l��<!��}}��� ���m�.O� ؀'(W�{b�5�����鹣3Ob˓�?���?a��?����iۑE7d1vMaD�X���,P7"�m��9@�e�'�����'b 7=廊SSi��+D���=m4h��DN���j�4������O��)�	~�V0O��8'�z�4�X���TV�	f9OҰa�����?�e�1���<Y���?)Ф>:�:��.�9f���x꒍�?a���?�����Ā�=�$����H��̟�{&��[^�$�SGZ�dF���|��:�	7�MKжi���?1�?�\AbM�2\ߞ�wo��<ѱI�O�H)�$g�O�؈���\w�
�I��r݉:��6�bE����N����$�*,*���?���?����h���đ���p�jS�Y�(�cL�T����Ħ�I!@by�gӘ�束~����s�6���� YAL�I�M�i�l6�_�{06�n�t��o�8ۂ� ��k,�95w�Dسț��]@�%�#��I8ʓ�?����?����?a���!� �"8� V a$�H+O��oZ�g� ��۟X��F�s���0�Ȕ��q2�2K�,�(3�����[�!��4d���Ot����e�TA(H�jL�R;�U��Oހ?�P�@X�O��{�-Py2CyӼ�l�m�'΍5Y�"GY�%j�\Y��?����?���|j,O�xmZ�S?� �I�f�Hb��y!�dZvB{+���!�M��� �>� �i��7-�풤�U�BĀ�Æ	+z3�����ȻL��� !*�	�*c�`�T�O\Ą�'K����ߩ0������i�pIZ��zT �	{�l����0�Iן�����,�*D��2VNe1��0k��1�ʛ�?!��?���i��pSZ��h�4��<�҇ᆶ2�>��ˁ�L�����xr�v�n�n�?�#
æ�ϓ�?��E�Q�� %G$X���b+B���� O�OLD�/Ox�n`y�'+��'��NL�R��M�t)�N�x �`nA6D���'��	��M��
��?)��?!/�| ����1��p%��30h��������O��l���MCԖxʟt<#�%F _�R����|X�]��H�3vXhܛ iȮg\ʓ��n�<�?pƭ<�;P��%�C�4]��7"��t8���?���?��Ş��D覥�V��u<�3��&�X0��_�	�|t�'6M#��%��$c�L���V��!�� �, ��@���S�4���޴���B��5��'/׮�[��M�f�v�2=��ʃ�Ax=��i��I��I�h�	�|��t���9���P&�� %
=⡎D��7�@2�@���O���7�9O�lz�#�τ$/}�t��IĽ����aڑ�M�p�i��O1�NA���z�6�	&6�Z|8�@���R%p�bM�Q���	S! ��w�'2�4�'N7-�<a��?aB��!&d��V��&3>�#y�u����ߟЕ'@V6-N�Z�����O"�Q�+6��Hܲ�4xP ���� :�O6n��M��x�
 7Y�b)H����;�2E����?[uPE��*�#)���6�����?a���O��M��{�Y$g�.a3҈��$�OZ���Ox���Or�}���n����X�0��6bΌUG�U�����_#;��ɔ�M��wN܀��&S7�9"'�	N���'^,7���Ձ�4�[�4���+ڴ���Pn�%ɚ�Ѱ���#��A�A�<�g�i%�����	��(����d�Ic��Q��G[��x�{c�ӯk���'ߦ7̓�k�x���O��2���OR8S�E��F6
.`�T	9���Yԛ��b�,-&�b>])�킚3��X�D�$,�Z䢶N7 �t�:#N�Vy�Z.P��T�I;�'��	�yoL��%�2cTtZ�lN^��������Eǟ�R�-+c~�[R�ǪL�$u�����Ԩ۴��'��ʓ�?�ߴ\B����!�=2r����=jt"�T�~HZ��i��O,���Ƨ�Rd�<������f�D<Ky�
���,$ԡ�n�<���?����?���?y�����=�@��r+�4���@�H��_LB�'���z�`Z�;�J�$�ভ&���E�ʁpSNҰy��i"��>���?I��|$i:�M��O����Zd�b�l�B�6$C2�T�"��x���ܓO�˓�?���?���0�L�d#�{�������g�$����?Y.O
}oڽI���	�|�Is��Ɠ�bQ�L+e L�K��7
���'DF�z����O�O�韎�����6��g�Gg`�r���A�t�;�+�v�p��.�O�9�O>�P/�I7��BV��/b�bq�fnF��?�����$�O1���.ٛ�Q*Z) �z�g��TlV�!��ƠA���'z�q�Z⟜Y�OLMoil`	IR+���#*��8Ix Q�M��(m�#� imZ@~BDI�<�~ �S�$t�ɤ[�m�B�
$/��a��ƄQ�P�	fy��'�����Ŝh�t�5��<<~���uӔM�Ob�$�Oh�?������cc�y~ X���V�F��X�m�*4�6�o���&�b>�� ͦ�Γ�h<A�d��/Ɋ�	��X]F��FJ������O���O>�)O���O<�x�&�e�^�!R���v�ӆF���'���'+�	�M�'��?I���?�H
�')XӴ�ގ^��0�uhە��'4H�,���{�|�'��(���o���a&��/bX�-#?�ƌ&�h� Z���5� ��[�?QE�N���#�V�)�����B+�?a���?����?!��)�O����%�"����6�y�2��O��nZ�
��'�>6�-�i�ǢFghƵ"H�
G*pU� .v�dX޴vᛖ�q�N|HA�c������c!��F�� &�zV';g_��9�ÆJ�Blr�;��<����?����?����?Y�͎�AE�xy`o� ����c׼����iP��ݟ��	�($?�I�x��	�3�>7��-�OL�Lh͑.O��DoӂQ$��)����ɃA�f`I��/�XejՎ�1hD�D!��S��ʓM�^9R��OR��I>	*O�]�vhE�7~uj��B���!hi��$�O��D�O�4�6�4���b[:4�2Nܗ$������xB�E�H�<�R�~���,��OD`o�.�?	�4�F�j���X��R��E!+A�R'�/�M��O�`� ��!?����$�b�+i��ؖ�Ai��Ɉg6O��$�O��d�O�D�OJ�?�K�
�+6�f����$c4��$eI�����ȟ|S�4K�(�/OB�oZv�	�j��!�ɋ�s����3��Xt��N<釷i�d7=����D�a�d�r�~�Ñj�T#�����X�uC6�i1!C���D�����4�����Od���%Pf�0��T�$�R��Qq*����O��c��'�%b�'�rX>q+���1yn�����li�VI#?1�U���4^G�&l>�4�,�)�^�9���
9^�&���{�œ%.$\ ��(���KTB!�k�I6%�����C�6s���צ>C�)������Iʟ��)��_y2�`Ӯa#R����ؠ�1�X���1���-���	����pyR�iVpA��� �e���rN�yGw��l�%1��ToZ�<���h-x��(�����'�8�"�ˌ�b�r�R0��A�4��'��П,������X��S��j�`Z���N�v�3�N�.6�0l��D�OZ��5�9O^�nz��)�՞��r���	�Th��)�?1�4R�ɧ�''��1۴�yr�߁wzi�u�.��p� �
�y�g��Z]��2�2 �'YZw��I�O�QS�ދ+�����߃&�T��.��J:�@C���Ov�$�Or�	����0��<����?���
q�0 �	�]�t@�UIJ�?!��?��ثGjZ9Ou�D�i�D���?����Y��IТ|���Ğ#+�9�3ON�D�:�D@��7x���2A��
�u�g�O6M�g��U�r�b§v+~X��E�O���ON���O\���O�h��m�O�� d��O4=�5�!u�A P �(r!�D�O�!n�^V�20�09O>���?�%�їx�ZH��L&;��5g�#�?��iP�7�����
_�]̓�?�CJ�a��1�%"���\�@%Z�	z3II�L�qJ>Y+O���O4�D�Ox�4לּ�	d�`]3v�|hu8��<ѷ�i0N�:`[���In�'Y�*�����Eϰ�Z`��%�(T�[��`޴U囆�0�4���I�.Y+p�ʍ=X�q�G"��ґ���4(T�(�<	G� ��d������Y�&�H����#�0|�ed�'��D�O��OZ�4���	��oʫX�2�	�&jE��>Cv�A��V�y�Nt�㟘	�On�n��M��i��5���+7=���à*��3t/Wi�f��hȂ�P�q���_����E+QcG4�(r'� O#LD`��p�@�I�\��ɟ����t�
��]�D��$G��{�uX���?a��?��i.&ى�O�!j�z��<��c1���ַ���a�(��]���x�)c�l4n��?�)WNFզϓ�?��#�1
aa�?4(�,¢T�\��#���O��+I>	)OH���ON���O,�i%%�%�>�`	܃��|`%��Ol��<�1�iF�q�R�'���'|���O�Rt��[6aي4�Ԩ�!<`���O���'h6�_˦��N<ͧ�z1D�3+ 7�J�P� �# �'#p�P2+O.����?	@i%���eshd� ʆ/|4(;��<*��d�O �d�O>��<鄼i�2<�c�#�r�iF���{Nֵ��/<e��'s�7��O��O���'����
<B�t����d��)�FMNͪ6MԦ�0�̦}��?� �Qn���5����:�� 3Lp��6M��y�P�4�I��,��Ο���ޟ,�O��4�Phc��su�8I�C�kl��I�r��O���O������X���]H���k�c,�0�1^�Y��E2ٴ`>���8�4���i��8�"d�c�d�0�1��4:��m��L�����I�8-�ٳ��'���'�̗'���'��iq�?4V�}�����o�$q�'��'�S��ڴ\O�y����?����� 5��"s]��z��^S�������p�I��M3��i�zO�Ȑ3E�24ll���LoPr���?On��&Bk>�0�ǋM�ʓ��%��O(�*��'���Q�G_�V z�`-�x���O,���O��d�O&�}r��W���ŀ���1�[="�M!�	u�F�<�b�'!v6�"�i���J��S��P�ĉ��F�����z��"�4z��i`�����i
�	Gr��*��O��<K� BV��}��mK6i��iy /�a�	wyr�'4b�'�2�'��D+>�P�e!s�\+が*3��	��Mۓ������O&�?�!�d\��'��A�4З��������4����O������yX��W �uy����v �EQ�|�����c��`WV�	vy�
1���r�R6Dr��Ew�2�'��'��O<�ɍ�M��"̻�?at�ƙ~.DY��UF���&�8�?�ói�O�}�',�7�Cٟ�m�3�`ѻ !Ҡ>�)Ӄ��<R��tmSʦe�'�@��� L�?����T�w��5��j
9w<�Y�J]�:h6�'�"�'�b�'��'�R� ���A+�!p2P4]y@��s��Ob�d�O��oe/,�̟ Y�4��P�څ�D�ˤjV�T˱d\;��8՜x�!i�Ԡo��?Yk7�צu��?!ŬDh�? 6P���C�_��H��ޢ ) 1�����?1�"���<���?y��?���\�*ap�M	4hu��B����?a����D��=�w��I��4�Op�p��v,у�M۳S��p9�O4��'�6֦�H<�'�"$��-w�P�@@�&��B�g2x��'��m �*O���\��?�##�d��=6ZYbԋ�$VTe�d&]h���D�OB��O���<	�i*���VK�:B7J��*;v���DM�j�B�',t6-&�������ڦH�.ؤ��EJ��� @a����bR9�M���iNX,���i��I%f�=RE�Odౕ'��+�Z}'x� ��m���'3����	��x��ş�	I��E�5r�#`��"{Z���CD\�7m�Ud���O���+���O�oz����4PPzm[V%(-@�K��Q��M��iٔO1�2�	iӌ牓s ���4|�zEÅ%�>i
�	=L;^�ӷ�']Ҕ'���'���'`�5��-1�<�4(vbrE%�'u2�'�RR��PڴW8Q���?I��y�l1���
�:7@ܢu�й��RF�>R�i�7�@�	�	ʲՉ���'6�8��R3��7O�m���#O�xt`J~2���Ofth��V��J�H���@��$�����?���?��h�6��_�*��3�O���D�u��	��D����'�V֟��	�M��w�>H���ј�M{�D{4HX8�'h7����4Z��Q۴���H�Q�T����nU�%���[��ݱ�lB?:Ԍ���1�D�<a��?	��?��?Y�Y�%��Y0�e�j��
Th���?��D@:��0BqL�)�?q��?�3�i��s�$�"lS�2��PJN�<�u��IɁ��D�Ŧ5bٴ
s����O!�T%�<h�b+,_8�"R>p��=2��.2��8 ��bv�'���&���'ł��U*�$^XP)rңF1f_@�"��'���'q����^����4.n�:�OA��#�H�)wJ��g���V�E�S��&�Ec}rGp�ZXo�+�M���/D���ڥE3M�l�r��?#���ش�y��'j� �F��?��_�����q;�Q�=���Y��ԪH�*�(��e�P�I֟������	�������wz����$ :*�;�ɉ��?Q��?1b�iS\y��O���}Ӕ�OXh�u��[�zD�#)o��h�6��v�I��M#����O,S������І���b�� *=�<``i۷�f`Iq�/V�%'�p�i�7�O����O:��_�G��RSjZ_h�LIAB�sw
�䜞JZ��d�O$�ʀ�N�n��	�O������3Q{Ҕ+�ˊ0?i�Z��Ul��Iɟt�I�<q��Mg�i=Y2�S>)��F��1��C1^���DTv˘!j�)�mΐ�3��My�OP�C�����%��&��̚���oGw@8�I�+[��蟰�	՟�ǟ ��Dy2+ӊ!U'�!\X
I���3�x9��;{t���O��D�O���|����y��i�p �k�[��d!U� ?ڠ�¥�`�am,F��en��<�޴ ��(����R
Hx�Y� yd,W�,;w���\A ���<Q��?���?���?���?����?���BB��,�)�L;�5R���'R�҉��A��On|����?Q7�i���O��f�O̕I!�Tax=z�m�{��&�Pئ]R�4<��6�;Bf�O��T�O��Mzշi��$E�`X��ďQu��A��<8}�$��Z�f`Uk	ȒOn���V�'i�&
�+`|�e`�c�p�{wa�);^��'3��H %�I�M�Q"�����?�4�!(��&l�08�� I��D��䓸?1-O ilZ��M��^�h�ɳ>8�Pâ%|k�b/m�:��ٟ8aрW�?�j�Ж��cyb�O������9�I<�rr��$Kh8�"tbŹm������h�	៼����ɘ4��ؔO������p�S"-1=d9A
�B6�On��376O����O����O�ܦ� u
J|H�h��Ѣ�D	VޱZ	���	��M�iy�7���7�m�,�Iam䑃e JbH�)�����}���]�I�(
3�O��My��'/R�'�'R$� ���Q�&�h��`�m2j�Ɉ�M+�"��?i���?AK~z�.�&�0�G̘(J��F-���e��]����4���x�O����OsM���՟.���De�<<���Q:\���^�\��/�Dg�i�IUy\
��L�2`̢Bvt�z�ŉ�0>�a�iP�Mh��'�^`朄I|�,X��$k�j�R�'�7�/�	��� 㦹��4h,�&����L���.!�(@!cS"-���P��i��ɎM۰y��OO�1'?��]�r� �W`�EM�(
���>�|�I��L�I�,�������[�'C�b����|	6��7$˃u��A!,O����ۦ�3w+*���i��'|�C&���$@r�� ���	��8�D�ʦŠ��|�*���M��O���Ҧi���c$�&<�zAs%J��,�i��7FP�O��|Z���?��q�t�{q(E
RTJ����'4��J���?Y/O`lZ�r��m�������R�$L0a�d�s�T aS*AP�(�4��d�`}�e�,o���S��玤v��Q ��*尜*�uy�h��H�X��O��Б40���� 0�I(t'V$�r\x���� ��?I���?���|*�T+��K*OplZu�
H3��
�ae�I0IK�(� ty��'Z�'��T�4:ܴNHޔi�ʎk�0zP�J=P���ɣ�i�X7��%�6�w���I+V�l ����*A�� �D���B-�Is�cѴA+ ͓�?I���?���?���?q����* �"B��=2T����g�Zn�t��@Ь��d�I�?��Oy"��y7�Q�"��d�����C�[3�7-���O0�4�*�I��ByI�`r���)� \<9t%�P��������ai��7O��K��?���(���<�'�?A'+�!8��31�P�D�ʕI!��?Q��?i����ŦI���Hjyr�'U,�Z��\�U��xTg�%G��B1�$|}�!|�j��	z�ɦA� 1b�Z�9��Q�@3m{��s�"O�(���N~�p��O���'SBp�����Q3&e�"PZ���?y��?	��h���dA)f�HL��R���!�U ���女#щ�����I!�Ms��w0,4)>%NzIC\��]�֮x����47�»i�U��i��	^�%���Oل��!��2WU>��/ʀ,\pbD��M�IAyb�'�b�' ��'�L��KF�����p�T�D�>�剆�M�d����?���?�J~��<�%R򂖚fKL4pa��[�0��R�4z�47�2�x���,��X<8��Լo�(J %W�W>�T`6���[a剕\�^�2�'Bn�$���'�e��o�g�&�h��Lm^9�@�'�"�'������]��b�4A��e0�j�Ԥ����Z���sa�F��VA�ߛF��}�r�Ƥ�	�!ؓ��'�"�R1hv��7f]�da�InZ�<��
�&�������Ep/O$����\ڀ�O�7f�tHE�5HN�r0>O��D�O.�$�O8�d�O��?���������+�(UV�Sc^����	ٟ�3�4#)�ϧ�?	�i��'��`��-@�8�x�^��j-�$�O��O7����i���)4�h!���^$�B@�@�ۯ�H����B)Dv�ey��'�b�'�"!�. H�h�)Gb�̈7�ۏ1]��'��I�M�NЈ��d�O�'Wt@2�(5�eKCmH a,��'�v�Q/����OO��!����D�m�L�$m��b�N+Z�Y��vy�O�du�I��'��e�+�>N�q�ќL�����'��'�����O��	��M��%��&\��43(
GM�<�����?i�i��O���'X6�٫6�%���ƞ<^|a�m�+3ڱ��¦�`�-�]�'�������?a��R����Q2��P�u�@�-��qd��̔'D��'���'E��'哼~���:��شf�y�z���4~�F�p��?Y���'�?q��yG���*�������]�V�a��֨�����O��O�On�(��io����P^ll[�H��}�<�@�O=(�ƶM��j��h�Oʓ�?1�'�V�AP�
�Ș��)���5����?a��?+Odm�P8NȖ'�$��`LDtBci�����垲yO�O�Q�'�@6�BĦ�BJ<as�D�"�VQKK�b��2V��l~b&��b��lZ5�L���O��L�I�}m"�ƆY�ԕ!��G�TRm�����y|��'��'b�SٟD!R��_��s M�+ �$` ��֟d��4i���k-O��m�V�Ӽ����R�t�����H�QB��<)��i��7���u��-^���'�ف��H�?�,IN��qWbE�G)K��H&�P�'���'/��'���'��x0�&��5��ܙ���&'fBe�P^�`��4Y�T=)+O��$2��hYrdvl�\�N��RM&p�/Oz��~Ӕ<$���望��ҍmO���'��C:�� �(�5�bܠv@�<�ڢ_`��dہ����D�[h�
�F[N�25j ���@J��D�O>���O��4�2�g�����%Y�A�=z��㵎
�P����!ĺ��z���̡�O6%m��M배i�M��Ĥ>"��c$�� �pE!��V3O~���&2��'N}�ʓ���;k�M�1�ʴQ\B��	J�����?����?A���?Q���O�����*�V�H��ĒZ<��8�'�B�'v6�МF�˓!���|�k��.^��$��#vu�4�5m�8l��O�m���M3��� ��4�y2�'����,	�JDּS"b�oJ���*Qd���	8%o�'��۟X������ɵP���P`R�&�bU�p-� �^M�	˟�'HH6m�v�^���O����|Zfm�+�F|���
-b���A�j~�ɱ>��ik�7-�|�i>��S,ݰ��ψ���Ģ�����B�H!�f����Fy��O�lX�ɥ��'��<S��I�GV�ɘ���O2��	�'��6M̴&%3D��F�i�'�M��{r��O��dA�?)�Y�H��4?�p�o\�g�̭J'�9����4�i�7-O�!�6c���	
}+�E���O���'�48��Ϡ<�P����M�XY��'�IK��ܺΎ�H�Uڵm��A��y%@M��MS��Q"���Oj�?=c���SR��%w.���W@�z���b�*�u���e��$��S�?9���y��o��<�6
�1R�.�j���OryB,F�<i��تF}R�Ė�����<-Þ�s%g�D��b��?Z�t��$���:�������ޟ�3q��$4��	PG��)5���@�y�������M��i�rON9i�LK�u(D�zB�: ����e����u�'=�Q����{�Ӄ&4�˅���t��s�*�ك�ޤw���Ӧ� 蟀��ɟ,��韨F��w�޴�@k��h�Ne!�E�('�4���'�N7m?0��˓6L���4��uY�̩l'6|��!9I~�3��OF�d�O�6��%_Ǫ6�$?�rDP�P�`���\�HrgEx�!`e�ƈEO~�*J>Q-O����O��d�O����On��D��0�y��j
6ʢi�<q&�i(�[��'���'��O��O��D8�f�A�vW��W�Z�TT��+	�vO�O�O����i	�2� Ș���^� +~���|I��q�i�	A�|�c$I��O,ٺO>y+Op�r�Q,*ӂ�C0J�M
����O�$�O��d�O�)�<A�i����'/N�S%��0<���AA�)����'׌7�O:�O���'"�'$��(��
�PLBꆗ۰��  [6! %H��i��O�`K!��'�:2��<���ǿ[�>9�`\c ��	N4< �`��<����?Y���?���?ي�$��Bh0��d~G����j�����'F� yӪ�x!2�4�dަ5$������'L��f��R���� ;��_���-�O��N��b�������
��$��G2bT|z��ŦIF0��Q�'5x�$�ȗ'9��'�"�'ǠܳAG�6i|�0��'ʡ\�Z�!��'DRU���4	>V�0���?����iӽT�|�qQ` X
J}�Ō�i��I���� ���4n���)"��Y�W�	J�)�䝪K�:���-O2��8 ���Sd.2A�@�I"J�Y�N~[q�p��?^-<��	П��	˟H�)�SAy2w��@��'�"���3 R$"�!7��� �ʓ	2����SD}��w�	���[�@����@���Y�/��A{�4���1�4�����|�������	"I�Yk� Ԋy���bK&U-��	uy�'���'�R�'�r[>��HځJ�x��r��_.�)�̟��M��oU/�?���?iH~�"ޛ�w���r������b���jQ�IB��x���l�?��Sܧ7� �o�<�Q�̨*{Z� ��h��s�`Γ({" A��O��{I>Q(O�)�O�=��j5d�$�B��e�Z��T��O����O��d�<���i�QB�'���'dL�*g晄��܈�^�]-�id�d�z}b�y�,}mږ�ē/��4����C��j�E:@�`�'��-;��F�V5�I���D�F�����'@����+	�7~��2 ǈ\���'���'$��'�>	�	�{h�b\�\'$ف֣j6��ɨ�M˗�΄�?q�Yԛv�4��@橑�-���1� ;�<��e8OZ�o��r� �¦��� ڦY�'$���?�T���
EiA ْ{�������;d�'��Iٟ(��ԟ�����ݧS���1��[+�]J�k�v4�'�67mM.q9��$�Ov��4�	�Oܡ���8(���2���fq� �r}�J|�Emڮ��ŞI�����	=B�>���Z8R�Ι*l�-'���".OFu�`J��?y«0�d�<g&��!*r����|�U*W���?���?���?ͧ��D���y�	5�'�ؤ�cgI$���eC+�J|+t�'��6m1�I���ĒƦ�9ٴ_o��(G�y4���%�>>ߠb#��h��Hĸi=�I`��I�Q�ON�h$?5�]N�t�"�sb�dZv�H�=�l�	��I�d�I˟p��G�';���H#�^�g�>��p)I�xD����?!��-��V�L�����'A�7-*�$��"KD��4
ߝ��T
�m�<ϒ�'��ܴ���O�`��i���y���P���J�P]bW���sH�7�RDMu�LyB�'8�'s�Å9]��I���X�sܔ-ԅM ie2�'C���M��.�?)���?�*���VD��n�xa��\u�Q%���/O��tӤD&�ʧ ����J�!B��lB��V�T2 
�yT��1n�4��4�2��2�ғO��3�M�\�<C1@7!HPjOdo����h&��B�lJsh�%��0$-LKy�Ai�2�HJ�O�n�
B���`��kL�E�lE�M��,	ܴ�6*�g��6���x�HۑjE��lEby�J�a�t8�왢-�,� ��yb\�����L�	���������O\T��
x����J����b�`�(P���<�����OR�6=�B�bE�b@xٳ��<+���$����4\����O:�J��i�:|�� +L�U����u��G�������!��V�O���?	��>��P-�8Έ��$�G�r���Q���?9��?�.O��oډn�����	�'A�9rAʄ8vu,�ybc�$���?q�V��h�4!��)��݊���`؏2 �� H<I�ɲM < ��(f'?��P�'x�I*�.-���p�0�ȫ|�f�Y!N�������d��ݟ|F��w�pQ�F��	J����Q���b��'JT7�j5zʓ6����4H7o�;A�q��C�6����:Of�o��M3��i%B��i���;l0x�1��O��%�B�L�E��9W��S3JRb�Dy��'or�'r�'��f�)E�"Y����R�6�b!c�%?Y�I��M�q-\�?����?�K~�	~:�r�!��uV�%J�/ǰu��	��U���ڴD����;��	ڄ�xWF (j! GM/5޴z�mӘ�
$�(O��8�
�6�?ِ$*���<Yd�:u���Є�-{b��V�S��?	���?A��?�'��D�Ӧ�A�Pڟ8ZWǒ7g�z�F�I<�p}��&m�piߴ��'Ҝ�$��/v��o#	`�(��Z�^،aѤ�U�`B�c���q��?ya�ϗW?��5�������+��!��̆�s
8�'MZM�$�O��D�Ox���O:�!��8�RT��#��֍{f��5�$������I��Mc����|��:���|����3n<i���g�D�`C -��OX$m�>�M���'��)iܴ�y�'��99S�,2��|�p �/T�|A�Ҥ(����	N�'+��ӟt��ڟ���gZT�R��$=f��s %Ow� �	🨖'g�7ʿ),����O��$�|Z0�G�+c�ۀ!^t(��P���Z~Ri�>Q�i+�7��X�i>��3� VЋg�E�bXe�@�<L I�$�&��W��ʓ�Bw`�OV�3H>9'A�na�l����$���P�A���?��?	��?�|�(OZ�lZu-�-R�K�r�a�%B�{=5����cy�	r���T��OZao��%��Y餇���e�e�ӈ(�H�K�4*��VR�vڛV��@�$���4��Zy��Y
aXXQLG�7�<%����y�U���I�����ٟp��㟄�Oce@�jD6�
�,T!/�����y���S��O��d�OΒ��$T���%fe��Em�2Ȭ@��ɪb�Ph޴2��F�,����__�6-a��37�7��I�fH�4$�[R�d� pcA�#i�B�y�	cy�O�Z�9|fŠ�/�#M�r�1 OL3~�'�b�'��ɂ�Ms@�&�?A��?�Q[�G��ǀ��T��� ӓ��'�D�]E���a�Z�'�p��N��V�<�KG��5*�Ҙ+�/3?��U-S���Q�]t�']���d_��?b.�.3iV�jg�'*�0��-�?����?a��?���	�O���C�2@"N��HW��Uq���O��oګN� a�'��6;�i��i�������ϑ�0�C�e�������!ش���4����%��'>�(���b�?Q�f�Z��Y�^z�"�$�<ͧ�?)���?���?�Z�Y�D� c)\�hP��d���D��u!���ΟP��%?�I,)U��&�)�V�����8J����OH�l��M�x����yq-�&d0��=G�@�pF���ٙ�mKUy2�z D��ɵ-�'%�ɋi����G*�e�Ƹd$� B*������)j�˟��X�B�*�)���tؘ!�6%}��2�4��' 
�3웆�z��lZ�o�*�f˟qy	�d�e�Ua�KЦM�':����?��2����ws>�r�F�^߆<-��a�S�y��'�qqWI��CpV��m����b�'���'w�7�I�VU��?�M�K>�0aY(�2��B�Q��D]K�@��'��7-�æ�S8��nZY~�aP�N��.;/ThD;��/p2hEy2�����ґ|[�p�?�d��(	�80B敟5��m�%,
S�'��7�E�v�d���O����|��([�Q�
���'0�Xk�,H~�-�>i��it7-n�)���ݒo�	�Uj �21\j#��9nlN,�G�S�3�j)O��ݥ�?@�,�䑘!r���s`�Zk���1
�G�B���Oz��?�|�+O�9m�!��<����ny�L�$�Q|fn\Z'�SyB�vӺ�h��O�o�a�P�B�C�w��)���u�Pp ޴Uk��Ϛ+9��f���Z�Ov��D�\y2� e�xX���4y��4�y�X����Ɵ�����I��O2>���R>5�B����3=���gvӾ0�F�<Y����O@6=�6X"��
-\nE:^w-}�bǺ��F��O$O1����` f�F��#r�N�8 ���X��G[
��ɍs�0%(��'�x�$�(�'-��'����t�]�L @��9N�~mS�'���'��^���40��@���?a��{]�% �!?L�HY��B(����B�����M�ưi+O�$��B�=�U+vF��#	K!>O��Y�gE*��0�b���$��OR����@q>��Ɗ��z�
L�ʊ!0���?���?!��h� �Z�W����5G��%p2�"�䚨@K���Ŧ��!NǟP���M��w=��*A�P�b�4���RP�I�'T7��A��4I?���ߴ�y��'�,��aa��?�*��C!HKL����)7y�Pxb���"��'z��蟴�	ڟp�	��i=4����7v �i�b� &���yyR�w�`����OX���O�����\��Y*BD0z���w�_~J�u�'��7M�Ѧ�cJ<�|�W�ŤGL���ŝ	��1�5n.]�J� �d8��׸y�L�b�G�OH�2�hE�%"�/]^��r��H���l���?���?Q��|-O�Xn��h4��ɡB<�U����&�R<��	�MÏ⬷>Q�i��6m�Φ�ya̅*���5�2}k�R�k(�<o�E~bH��u\8��xܧ����([�!���h�����ųu��П�������՟���A��nW��k��]�l�꘻ �	(v����?��/\�F�E> ����M�J>iuK]��J���ʶ5#D����]�V��'�N6M��ə=�V6m2?YuKC:I��Z!�	_J4�홟`�*�p��O���J>A)O���O�$�O$$R��Ȧ2�s�+��4��A�O��Ī<���i��M��'S��'��S% ��j1i�8vyB���U�B�hS�	(�M���'.���	]/��0i�HZ���ڧ8\��RV	� p�$5 �
�<�'���V����� ���E� �ڄ�"^l~�j���?����?��Ş���N���B�:2��7���00�X��(<.d�'��6�'�I���Dߦ��Q�pVf�9��e3�h�H��?�4?&p���4��d�8S3�8����˓<�
3$N�:kjpU@�ADTΘ���$�Ov�$�Of���O4��|J5.ֆ_:�ՠ�j��2t��X�G�qϛ�/;�r�'�������݊k��T�p���R}( ��%l/B,�޴:b�x���/¤j@��6O���p�2J����J�:	P�JT1O<(#�ꞁ�?1 !���<I��?� ��XH �u�J�+!�U�bY��?���?����dȦa�U �ޟ���ҟ� �!�;> p�3�ϱ,���{��AO��1�����M㢷iŰO� �,Z#��$U�)tƍ�K�Bhу�� S���5������A�S�5�(=1 O�~L@�a�)ߞ���4vPZK�K�
D@�nO�~"ԙ�F&Ӻ���z��#�ΤHgß"Z�}�"N�9b��RDB/Gl.� e�?:���V�"\�Ld�ǨO:��3��h������Z "�a���
���Af
V�Ģ�,Br���/��Ddg�F8r����躑[R�JJR���G��G��r�
v�L�9�)ՊR�<]���� 7�PQ��K�	�
H$J�@}�� b���裨��}��ـ� {��W��90��3���6�jR�i�R@Rv��O����O �Ok,�J� pӨѺQHx\�_�5��f�'b�qh�'a��'���'��'l��ϴjȈ�b�E�,i�\@"(�������]���'���|2�'�����\/��R������\�4�I�}dZ��������OR�d�O����O�m��Ϭ?�!��|���oֽr�:�X3�sӚ��?�N>����?�$�>b:�o��h��beB-z�f�@��E�z�v듀?���?����?�wh=�?����?�GK�b�����E�P��)��\"��F�'�'!R�'�f ��e���ēI-8h8�,�eF���0�$]P�nӟ���֟�ɵeZx�O_R�'��@Ö#z�B�&��?ʄ�kP�7�XO<��OF��&��'�1O�$B�|�q���iZ�b��"C`6��O���ԅ$��$�Ov˓����?����Sb�]�3�8���I��B˦I������oX�HH�b�b?�"GGE��Ny3�����b�b������O��d�O��d�8˓��I�
hWJ�Q��̳|Rt��`A�IXH�oڋ�a�a�5�)§�?��gH��(|z'�u���Fa޲-ě��'���'�>�R6�8�I�����r���/S:>R<����i��>Q�aU̓�?����?��F�k��C���A��pC��+g����'�ꐻ��>Y.O`�-��ƒ�+�|� {䖸cY���V"A�	�����Ɵؗ'�@ex1�.�]i��s�^y
�B�����d�O0�O��D�O4��n�Gk6�I��L�#���1ⅉH��O����O��D�<ɴ�ȗ��t#ޫm V�ht��1@�`��⃱�MS���?Y����?Q��pɌtq���|����L���=N���QZ�`��؟���Ny�f©\�d맟?���?(��($,�j@�SB<��'��'��'��j�DB��84�"o�%[،��� n)��'lr[���1�M���i�O����JX��Ӭn,dj`Eɳ)}jF(�B��ҟ�I�,�*��~�$-��	#`Xك#A13ʠ��ڦ�'y�E��k}�z���Ob�$���ק5�,�+H(����,m&�iK��Ս�Ms��?a�b0�?�I>�-���"t$�P�&U "��a�ň�6�
�J��n�͟<��ǟP��2��D�<����z���sÔ�T�`y۰F,H4��F۔UxR�|B�	�O.�q��Ƴ rl��ȂI��oNݦ����L�	K��A�'�r�'��O�����?��X%#M%k�N���i?�'�T�-�i�O���OFm&�ͱ[��QAf��g�8�d)�릱�ɍ"Ɏ���O���?qH>�1F�6]�V�8\4`C��~��'���|��'�b�'��6#1 ��@ԣ�� z@�&�|��#©����<�����?��L��u���Ɂ3"̄R0�h�dǞ���?��?I(OʅX����|
!�R�UJ`h!"\]��$�̦M�'`��|B�'aRA3k=���?��2���n���p��?:���ៜ��̟ԕ'F.q�Sc>�O�p�L`��*�J�k#��=o�8.��'$�	ӟ��Ig�%��e�iX"ؑ�%X�I��aa`��/V�V�'�"Y�pj	���'�?����m@�
���q�R�OJ��xp(�զ	�'��'��y	��'���ԟ,�s��i���$9\`(���"Fu>0mJҦa�'+zmk�cӶ$�OX��O8>�k���!m�Qʘ�)3(�4*�l���h�	2:g�������'�*��Fk�qdH�#'п3�AkG�Ǖ�M���F)*���'�2�'�ċ<�4����ŤU.=����H:�l{#��]�f����L�	֟����?A���].7)���ʇb�&8�C��g��n��\��ş �������|
���?QU*�/>�.�����.x�j��2k��'�2�'kJ��o�~��?��?�#L�.�΄0%��L���w�בE����'&��{>�4���d�O��.�"i��l��VY�d������2�ipRgA�T�RS��SП<�'\��H�74�����$Y�SeD�g�$qSS��'��O��D�OV8؆�޹����@��l������L�`����O|ʓ�?�nF����J%,dj�ZB�;x_ ���� 	�M{��?i��'�� �ۊ�x�4MN��1�ݢ'��u��Һ:��5&���	jy�'� ,�]>������ͨ�+9g��Q���m�֨1�4��'k2�'��i�n����w��Ԑ�c@$V{�R��șZ%oZɟ���By�D^/^�l������klW�rc��(C�5$¦����F^���I��̰p(E�8�O����5�i�a�D��5mF��)"�E
J�7�<!t��/��/�~����ƒ��a3�X"v�a��+�QkB ���j�DʓOЖ�+�
U�O���M�e�C�T�lQPvjI�z��a��������P��<�	��,�	�?�����C���ɪ�K	F�u� ��2���'��������ON��$��$[�U��'��ِ��I������� "H��L<ͧ�?1꧀ ��� �&����2		
���R�i��T���랞��9O����Of�$X�A0�A�0a�t�`e�Je��l��L"�­���|����ӺC3��/c`ЪA  [,R�"D�L}2��1"P���I���@yb�ΙH]@=�����#R��1IT3w�ЀTk4�D�On��6�d�<�*��g�-r��׍t�is���%��A������O ��OH�7��)59��% C�׏J� !�Mě��;����OH�D,���<����?YB/���t�Ɇ(��,Q�a�5	�' �Y�@�ɚ2F��Oq�!Z65S�eyDA�=�H!�򈂫Qi�7M"�	ڟL��#e��t�r�5�_�3uV�C�JQe�Ё��ǫ#�V�']�\���
�#�ħ�?1��S���7jԭ*p�T�o4l�K�cw�Iiy�͋�+���П��!�������[������i��([3�TH�4ao��ɟ��S?��d��r<j���IH��`���蔛!Q�F^���e�ϟ��J|�I~n��`9��I�[�����ҀXK~6�2��uo����ҟ�����|�����@�bhG�d�2�)a+N���i�z��'�BR�($?��ٟ�P��U�G�A`W�]X���Ug�+�M���?�a�ͱ�W�@�'�R�OTX9 �1;��E�g(E�7�e�5�i�',)������Oz���O @�'� 44P@�cUB�$�P٦��:vLq�O˓�?*O���"͂�@nN����k�P�
�S�T�,4�{���	����	˟���iyŁMLj����.�vi��H�`��D˦>Y-O���<Q��?���<P*|[��_�1Д����K>2�r��<��?)��?�����y��Ḩ6���`)�!Y�E*�S>:��mZwyB�'��	����I�l!G�w�֘�\��'j��XG>|1�Ȑ�2n�6��O
�D�O���<a��\�W��ٟ��

ZZ(�Nd<Ti����B6m�O�˓�?���?Y���<�.OJ�x j�O_�1ы�L� �4n�Ŧ����t�'�d��$�~����?���YZ�BL�M�{6iEl~	h�R�l���,�I�N����0�'�i�&���2��L�1�d`��ʏ 8��T�(C/C��M���?9����U���Pұ���Q�xR��Y�J��g�z7-�O���_��D7�$*q�z�s��i�)z��H�-:�7-O&bum�џ��Ο$�?��d�<A�k�Imf)�� X=�f�`#P\I��\��y�'m��'���DU�Cl+�I� �� V�v���b�J�D�O
�DǇa�Q�'���֟h�|� �G���mn � �@�wB֜l�ٟ�'
k���)�OF���O� [���?$�����ab 5�`�æ���

���O���?�-O�����	@g�@�[��@�T�ܹ+��`�P�hY7�z�P�'�2�'�RU������}y�h�S&Qz\�EN�-|4�yïO�ʓ�?i.O����O��$�'>�"�p��%u)Ƽ$�٦s��;:O��?1��?9(O���0��|��X�J��A���g����b����=�'E"_�8�	���'�~扱Pl��ӃD	Y,��s���K�pX�4�?���?Y���%i���O
�..WO��HG�Q^��\ٳjq}�6��O���?����?�BH�<q-��� ��.#�=�� J0lv�z��˅�M���?!+O|���O�W���'���O�����~l�i[&d�n�\X���>i���?Q��
F�=ϓ��9O$�4-��1x1J��T�� J�Mט.�7-�<��O����'�"�'��N�>��v2qP&�4g�Y)$� 5h�5o�P�I�d��I��h��ퟤ�}��F٤NX¤� F�WtX��K򦍹5(�M���?����V��'�&�Q�֎ )��+G�ѿxK��u�<�q5O��D�<1����'}n-8�l�f^� ��a̠��w�����O��d N�R��'^�����?�@�����%��)D	R�A�0=nZi��5���)��?9��P�f=��(�3�>�i��+2
����i�b�Y�;u������O���?�1>�~��N�G
��@䋽Ф��'�Y�'[2�'�'��U������2�Bde�mQyR͕Wv���O���?)O����On���!a��ы�#�fM�`b�j�2h�9O0���O"�D�O.�$�<��FE�x�	�1	ATE���,��e(��U�J���Q����My��'}��'�b�����)�҃�g��p�"-�u��`Z@�i\R�'oB�'
�ɑZB�􊮟���LU+����K|:�ʁ����,��t�i�BX���I����;��IJ�����4��o�+���i��7�V�'�S���Å��)�O0���ޑs���ZV`*�
�w�Ir�h}��'���'�L�ћ'"2�'H۟$����q
h�2�]6#u�TK%�iy�ɿk�U�۴�?���?y��6u�i�Qɡ�Ηa* �@a�m���d q����O��8p8O �O.�>S$�ˆ#y���Sb�d������m�6�)wD���䟨���?I9�O6�\X���f�G.�d�#�<p.�!�iA�aȘ'}�W���j��Vlm9����s�"=z��؎L��i��'No�)������Ol�I�@�bAY� \�4L`!���վ'@�6��Oʓ�.X�S�T�'��'�b�ÎޟR� 8���3@/*A�V)d����]{g°�'����ȕ'�Zc�c�K��mW�4�D}�O<~�$�O����O���O�˓{W����g�K�@!�cA7e?*0bD!��Fy�	{y��'��I��,�	��H:� �e㥌^	/d(;pb<��"w�C�<)(OH�d�O����<i��D+d�I$#H���+�V��)�BH�YX�&R�0��]y2�'=��'Ef�'+F �֥̀$��0i��X��(jת�>���?A����L'>q)�k�D��ݣ`聇hB�� �J��M�����?���1�������I�R���a�D�&O��![��A�L6��O"�D�<�)2I�O2�O��tr3B42;l��`��@Z�����#���O����P.��'��?M(K_%L��6��,`�hŰ6�`�b�k��{q�i
�'�?1��k��	'l����Hs�=�妈	M��7��O���8����}:�gK��f�@D��({��x�����W��<�M��?	��Z�xB�'_�թtF�=���!�L'vK8�-~ӌ����O��O��?Q�I	aLn-��+��EH�(�UJ	���X��4�?����?!�7t�O
�䯟����J�>�A���PN��P qӲ�OFl�ց@b�㟬��ןx���
C�D�P�ֲpQ.0�"�K��Mc����Ԛ!�x��'L"�|Zc�j�ē E<���(q.��O�Y�g��O"��?����?�,O�1if��<�T�'i܎;����ШP<L�h��>!�����?)��#�1)�.S�> ��)��۟tzj$�᫩��'���'��W�D�ɷ�����=0��Rao�&�4hY�$�����?YJ>����?�GM��?�'�1����!�^�fˌN��	���ҟp�'�x�3o?�IL�q�$`U Ȥqļ�����;mX5l�ܟD%����ܟܚCu�|�O�$�`�W����{h�}��j��MS���?Q+ODk��_Q��֟d��#IZ���,Ќ3��$ `���\��H<A���?y���<�I>q�Oe��cn��G���
R�4/��K۴��:|�ڨmڵ��I�O���RZ~b�3�0:��
7��x�r-���Ms��?���P��?�K>Q��t�V���u�V��73/��0��
�Ms� 99Л��'7��'^��h:�$�O~P�n�41�0lcHI0G�M�`dԦ��uaUƟ,%���*�� �F�ڰ/��@Z�d�PZ��铳i��'�Ǖ�0�tO�	&}�N�=y� �� ��&t��"H���Ms/Oz��_�i��E$>%�����=y
������G������"CĤ@��4�?�G�63������7f�<Q����(�v|���D�?���"a������?����?��?A*O��kΗ�2t�҅� k��ɸ�` �<��$�'W�؟T�'V��'cBg��+��Ʀ\�,��)I�K�4�Nr�'i��'�"�'�V�� ����.'�peYf���͡�M�-OX��<���?i���'�^�T�W�o@��{@* �*3~h)�O���O|�d�O����[���$�O���H�p�QS�K�[&��V�<)l�n����&�������s�j;m)�O|��dր@�����X:~A12�i�b�'��	�n�
]@J|���z�d�(ɖ,
pf�:*�T���}��d�F>)�s�h����9��BC�Ҿr��$K�i�2�'� ��G�'A�[�$��yyZc*�:,��z�株¤w�nA{�4�?y�(d�,a R�S�MKt��0*Ķ�LD��آP�f�WB�>ߴ�J-��Cbh����K�?�>9� JF4I��Q� �}�S��l�<9#�\����o���z�ʦ�:����~�����/B�z�2�r�Y��qHl���
$
'�.3�XVBH Env��6�O�UYFQ) b��S1�T�$�ԏbG�Ju�IAᚐIԤ�u�R�sa�L�4�S�yy��O/y��|����6IP%)סS�t'�Q�S��H�vm���?����?����&�d�O��S)EP �uZ�IEL1���^">��tP$&�;n�~���`X�i62������O|͚uѩ���	!�`�idK�({L� D��'5�r(�r���qѴ)��w�}b0�ʛ��'��}�@��(�(D�AƘ�}<$��@��?��hO⟘��^�P.󶣀97�@�Y�J)D�L�M]>B��y���:��&:�ɹ��d�<a�OX�q{�I���&Ez,���'��A��'�0D�b���O(Õ�Or�$j>m�B��*k�ٱ6��(r�~To;.�pf ;A��˳�Q�n�N��ē�;��Ѳ��Êb x�s&hgӲ�R7��(9r:Hcr�æZ��0��'�������?�/O�E����0+������/&��R��%|Of����{��L
�G"���Q�O�Algx�`�66�����~����fyl�9WB���?�/��0a&a�eX�ư��0�T[�?< d��O���3}:f�`�ǐv4��! �d�ʧ���G]@dS��١	@N5a��� 7T�b|^0k3b͵bL �.U�O��0v��n�* Pq-����n�j�D� �rh�E��OZ��B&]2gV�
JK�'���tO"�	��F�Oi��#�N>S%�!��'�L"=��	:8��I��;RhA���yqݴ�?9��?�e*�"}*r���?����?���(����� u	�����'z}�T#VE�$,T�3E�8۔`�.Uu*b>�O��K���W�h�P���:r��*Ԧ4��X�J�ן �`�@+�q��'.�@*���\$��� gςR}��b��'��	���4���=�m�'^
�Re�ھ5:6����T�<� ���6���>���o�1��MӐ��؏��?��'v�a�Ɋ�O�09#��J�;�D�ؐo�j<�U���'vb�'���z�e��ٟ�Χ%�B1��ɺ?��VM]���b`�B)6��ʐM�P�����4t�g�J��$��EǁA@������&d��K0��!�&���`�"��aI�.!��}y�DX֟@��S�'L�O�@�m�u~I���^8C��3�"Ob�ȗg�3+�<��S��t��pT�Di}�Z���'限�M;���?0i��,�N���A�q���F��?I��z���?��,���3��A~�'x��Q*�3Rs�Ur��5�� 
ǓH��y�t�I /��"I�����]%z���a'�c���%+&O����'<�7M馑��X�2�����<6� ��b�.$ i�'"��%�ʡ��B�T���0 ɸ����hO1��Pl�=���2Hܷ!*�� ��#zd���ɔ'�Ը#�a�4���O��';�ɚ��	(�{�.ܐ��@R�C6��H%�?y���0�C�����򙟼��-w��I3�Dώ��E��f>}Rfă�O�I�t!�%Pb �I��2/��A���>��BC�`��� ��A�'2�4��V�=|��Aŏ�'�\M�<q����<9DO�#�@�w�
�$O���+�A����"~,��"�BH��kB��9n��	Zx�H���95��Iӄ��8S����?D��U�ŴC{f�H"�x0ԭ�*:D��!BD�*=(��B��h��+D�8�DO�$� ,R�!4Y���@�*D�P�G+k��`9��Ҳr�8�U(,D�X�A�3�&���^;h\� �5�(D�$+S+�B	�5��2� �	��B��	E����Ԗ_;z��c% �l�B�I4V��`��I	��I6�X>B�C�ɤ5�����[g�2t�BGU%m�B䉇#�`�b#!�
Ai���a��6C�	�$��qbbC��A}� ⤂��a�,C�ɸ*}�I�G'G��� ��ۅ-�B�	�lh�95���q(����� H��B����!֏ӿy����ޛkM�B�	M��r��;`��R�k]���B�	�t�8��L+9Z�J���
76C��T��2��̀f�LY '��:�C䉮!X��1J�v���i�5��B䉅��M�f�$^�s��k�C�ɀx���ps'�	^�4�Q���~�^C�ɍB�eR�I�>�*�)���hC�I
"���Y�c��A�ۦ`rC�A3ppц���)7�� �K܏J� B�"2:8���C�:+!�	���#t$.B�;�^�pgG�(G�}1$�B�n|�C�I�k�$�Č�>����G�-'�B�Ʉ=�j��p`�D���6�ܭE���$'&��8scA$}��ͩ��	I�:i���s�邆퉓5l��`��h����ė+d���Ia�G4N6Г�Թg�1Oҗ�ę'o|�@2#I�T�|E�`[����t�z��G���)�h��6��6˸C�I�|�N�X'G	XU��z$���uY���s�ԬU�r��Q�Y���S��"�m{�)RF刺^3�M:6�Œ5B*�*��;D��7�G�s��j�&S:+kF=���<���i�����k1����GyRL��9�b��5 	�j��qQjS��0=��Y$u{ƹ*��W�",̓eT�NDF @���;k����v@t�@l�A�M���'h}�{�S����k:�(���V��A�P���'���E�@�D�
ٳ��ӭra�jI>���$���{�NL� �jM��㞌t0��K&"�Z�S��y�F��$����6s��6�^59�d0ȴCH��a13�@���S�i��*��V��#)ʝW���R#��y�dR��{	����M@R��kB�s���Gxb�>8�"Y[G��Z$>�;֌�	���?%qS�W�'D��"rJ[��P���3b@f;������b�Is5�M(����,۔:�ay�bػv�PE9A�I�i�z�B�I�+����78>�[��E\JTb��Y��U=�T��&�O�����|�&S�sAJH'h�}�WK�8kx�'��|�SC�+�Hl0�@W$��s�{
� P("-���RN-��Q CF�1 b ��'Jh�ZH>���H���'�5�c�TY�J��*׳o=��y6J#|&H�A��p.r<��I0zm��N,<�b�1��[*.� �Ob�3��+<Oz�   ]�Rq�歖��@qC��*LO^	�RC�,- � Avm!@hr�(�Z":C�`����'C,Z���'äa�����Z�	�$W�/�Z��:h����fLW�~�,ڢ�DG�>,ئJL�%J적��8.F1O�y�Í(DS�,���7Nz)�И|���z(�Ԁϱ�܉@0�ߢ�'v�h5��>�~��򃆢RɎ�bi׬��ad��i�h)(��''���à�>TH>�����
J���u*�>~�*�A���o�
���I�@.���JF@����d��m�"��S����a��.��$�77s�`
w��-����i��!7-
�{� \xf̓Dy�'G�<` �/�8L��y�/W�|� �'�@�=J��.\ꄁ�D�Q��6�*��ٰ�O
 �d�#.8p�F%)Z���&CV�����c¯�Jwx,I�E�� д\'�,K�MѢ@P�]ADf|��p�7�I%[�0�z4��B�ze3���c�u����1*P�G#j�1;2�Zf0�D{rb�=�\���j�I��@!��ϛ6��\��E�J+�a���9lO�X����=T�Nx2�N_��p�pΚ�:��A�'o��#�7Ng�^�x0�F_��P���K���+ ��T��@�P�{���W���As�[�,V�u����_>���d�ٍ?��Y�]z��'�����*��u��×?s�4���?��FcI�S�D@�#
�5S�YrS`�of|�D|�kڹHhzE��n�
�0�Ŝ�?� ��yn��إƁ�U��k��D�R���g"����Y�D�IZwx�
ao'�)��m�� CY���E�Jh�x�F��ȶǟ'm,Q@Wϓ��6�`�O;|yӤź>���9~H]����p����oS�Lx��7֐�ȁ�'�:�#�e�-��h�cj@�"��\3�}��P^L��ض��%�� M����>�u9�(�o����fԪG�Rv"O,R`�ə5�T�D&�W��X����e6�[�E��	������H��Ʌ2����S	� ����b6�B��\�Eb���>�4)��G 7��(�������%"Bpϓ�X��4b�X;�eH�&�/)���퉗L�Х򣩈�$w��(�hLy0ac6�X�$pA��7Q��D���8+'��!`���ñ+�#:��Op����=PJ!�礌���O!�3��Zo�8�&��\�`A�'�@�ᖓE.Z��dˡYWz�bȎ)T�~b�U?��9�g?鴃��=��l���B�#�(�:�́p�<�'
�Ҏdjӊʽ|h"�2 ��a��Kʱ��p�U�]��yB��!acDM�f!�!����۔ϰ=��*T�Cq�Q�t�#����� "���J(s��t	�'34��a��W�L������0��5;���!F60��3Ñy�|Qz�ǜZ�'�)��ŀr��+ �O��4�ȓU�t�I��ҨF) 0�4�T� �SD^�P��)�)�Z�"�ڨQ�d�	�ӪB!0�L>�a��*!�$�R.M�'B�r��e��xi�֊�N�Kq�lF�ɀ�)M�R�p���-r�qZ/мL�Ι�#M97�h��'KWx���B�1o�~�@d��:x�vn#�	�2X��n/Y)�9���)����g���N1.�ipŦ]� �*99��Q�{.B�>#�:50p͚�Z�m��
����sүR߼���I�&- Q)��Kuq�(p�>﮵� ��� ��B�It�&"O�1��ЇS�V8!�ڛ|4�Qd�*g �\{!d�1&���IS-Q���q �хW�F�>iqi�6EF������E��j@o��D��	T@��t��V�OӤPF��}YV�����-8l�
e�!%��ӓiU����҆�'Zt|�vH�������XEP�yB��He%Eƕo�da	 L�^.xc�M$�t}�fN#h���j$[5�JU�w�� �y�d	��|�)���Ut^��(��¨�8[r�L�Cd��|�&�ͳej��~*�ET�����1�(Y���޾���r" �\�<I�� E�|�RD�Q�R.�	2v�ӷPB�)��VTke�#7<|	!�"A�l���0�	�!���f��0B��ʃ)��T���%�PŁoP"h�HU�I4U �	�S�תH����.,r�EQ���x�z�����!�p=���	��h"�`D�m+A�dL�Mk� �9v��"dl��f�x�B̖r����n��� o-�N@�'� cb� T�<ѵ�3U�FږT/:*�BU��Y�`�dŃ)aP���)5X=��t�'P�Hͻ{�~1�T ބk�dh#�J�xn�|�ȓe��Dc�摍<��5���wW�H��^�M�u�:<���9I�h��FF��O���E#�"+�~]q�a���7�'���@���8���� U^p`��3B��ul�@GJH�o�H�RF�9��و��+�0>�gˆ#hl�C���+?��s��K_�7��1�Z=%��Mz�Wd�*��-�?�R7�� ���b��YK4;��A��ΐ� "O� ���/�dm�`k�Xm�ӈ"&��8�&AǔI>�i��дx�!`V�i�
�]�_n���.ٮ-���c
�|��C�	;&馄�ƅ(r�,�`րh�7-ʹ0�عA抣%��e1O��W\�]✵P�g��� d*�'J��T� �%b�)�����C��-ܔ�e�%v.\!)�
ODu�Q�߯E��]h7E�p����$�b��эW)??�hs�������߷H�5��,֙�Py�Z�1с�w�@;��߼Kܠ���1]�@}�'s."}�'��r��cR�c�h\�UҼ��	�'��2  <R��`"EI�Q�HX�C0 �!�@T]��	�
P�� �:S� ��7�$o�1��w��Psf s��B��!����S�u��\�H3�������� ��Q4�t	C��}�:��I-���'{�t0A�R��d�G����#V
� ֩[05�L��,��=s �f��́c�@���. ��8�өǾ��:rlh� L�"~Γ
��Y�m\��$ k�'p��1�?���Z{���Ӝeoz��e���j �L?0��m��!S�`؞dr+ޔ5Ʃ��ӣz���U�I$%���~�$�_�*�2�O�`���J�q�2ՙ2A�P�!�.x�T�k�Y�b��f��g�K�3��'�p��!�\�OA���Hן}�(�I3�<B26$�
�=�1�'�N�Z���^e�� �H1@þ-:�O��(�6�)�'[��̂���$�6��3�R9zX�ȓ�Y w�Ӛ1�d- �J=9�b�����X��)|	�E�T!�o�b$��y3��!$@�k+�̈fKЩA���ȓ	�ࠇ����\�G憼��B�$�"��Y��1�3�^��6��;��I�5���?�L�AM�8T+���ȓWd)fE�9�E!W���a�ȓ2v4�@�
,w@\�I��Cj�ȓ3ID�A��-t��b�ߗv��Ʌ�*���r��W�B!C��^���%� YÇ>\O�]��	(�D�r��hR���'��}[u��*��Â�]5�J�Ç�b�!�D�(_��Pl��!�ʢC�7"�џ0H�#As�OJƉ�#�]޴HZ�APK�	��'�,�b��Il�a2"��E�2�Y,O6���)�)�'=��E���8�ـ��C@3�X��z�~�smAt�����Tigl�%���5�U]���ŉ[�Tƒ,I�i�MҴ��gH,�O��PE��.&Y��z���6� u�V���54�B�	�78`�:3��\5�1�"
�>uwvB�	<?�:�8��Ľ2��V͂�%LB�ɡ����1J�Ғ�1Zm
C�	#e!\%32K�*
��
����1!�B��>~��Q��B��ے��� ��B�ɴB^�xBbw\6Ƞfl��oN�B�|�e��R�%J�鑢�L�h��B��G MB�K�7T�ųt�ʸ%q�C�>�q��G.戱�r��&N
B�N����'�/ ���Nנ)��C�	!dK���V� �~��iħ�3YbB�	<<�a֏Z&c0�3��K���B�I�_ZX�I���H:�E�g`�;U�xB�I%~���Ұ��V }�����Y�bB��.B�0A �Ћl���IU��2��B���(Kq+�s*8�q1�	pD�B�I�=�2lKI��� $kMh��B�	�m�Lа��9d�r��I�.��B�	_L2=x`ː�bTk��2�B��/:B�+�ň�Y�ɉ#�L6^�B�ISul�ST�ڟ7j���6(�;�C�)� 6���*�ثS�Q�6�h�"O��3䙡Dv�h ��� ���"O.}�*�<Y �٣���C���bS"O���V S�PdA3b��\��I4"Oz����mV��+чD�S<S"OJ����1��!� ��}8<D�"Of�	�
	`���)ˎv�Q�"O�]iVAżz�\�S(E~�l��"O#�Ԅw?��z7'�;�ظ�$"Ol-�v	��6���{߰���"O\��F��uY$D�W%*4�]Г"O0�sbk�7V�ݩ�
�P*���"O$ٳ��S�s�Bi�sG�!&|B�"O����"�8���CӅ�6�xL02"O.����
�K(��pb�
�:�;�"Ot\���:Ws�}�Ύ&1��HPA"O�	�d�� xa�\�ez�]��"O��R�FV)�Y��X���@�s"OP���P;��TP��Y�[$ �)`"OĒI��m@�Ȅa@�r�uj�"O\p"i�����CK9VHP�S"OBd���..�в2��j�`H"�"O��1�� #�@�C��<�v�R�"O����:[3\��#�66_��!�"O��P���(Jv�Z�Ē�"Z�|�p"OЀ��Á�-�Z�9���=�����v�<bh�3h ��ëhC�T2���yB�.U��HY��^d1	wč�y��Y�o�Fu�)�(j�x��v�� �y�'�u�������p�tq� 	�yb'\�U@T��F�<�Z�h���9�y��d�l��K*g���AɌ�y��(�޹�ֆ�����x�'߃�yRf���p��=b��<9%\��y��?�����a>����*�y���7�i# V=(����$a[�yR
T$��p����kA �[E��y��'T�p�z�J9dh%���S��y"�~���[�!d�j�2�iD(�y"ā7�=�t��hzI֣��yrώ7C���M %d�j-�� �y���) "�Ez$��2[��ps7���yb�Q si��OY�i���9&�ވ�y��	���� &!�X��ʌ%E�lC䉔/�:��f�@�ee�8�MЇk� B�	�T���P"/�V���G�S�-�2C�I��<��N/V�dX�4��U�B�	�h���y���"�-Թm$�B�I��(�3ތ(1^�Hc@1iӮB� [12	a�M�oL �2��3hl�B�I�B�p�#�8W�d(�g�TւB��������	3e=03���\B�ɲA���#�"S/I�����_�^�*B�	��� ń�kɞq����]��C䉅6_�����9"b;���B�IW�t��"N�#3< bQ�֘B��C�	b4:� .��3JT=L��C�	\��)z���#���[�.�I��C�;z!��B�Q6ID�̪��$_R�%D� 8E�U�@%�"�V��"�<D�����x�Đr�E�a�L��#�?D��a0�M�Y�����R�k��yC"�<D��I���*M�0 �!Z��m6�9D�T@d�rh�+�Ϝ(] �	qԅ8D�� ��5�>��Zd�V�& �V"OfmY@ON�>n^��wLX��x"O�T����Le1�����*t"O�����U�_╰f��=R�V��"O�\Z��n)�q2E�.q���"Ox�z���o�h�(��ط,lN4 G"O$�r%M�\>"d1��Ye8�"OT�R.�lG��zB��} �M�b"O�a[
z��`q�ϙAz-+"Oy&��@��k�SN���"OD��g9�<�R����z�:f"Ol9��
9L�^��G]?c��4"OrHx�G̘>�D���h��u�"O\�+E��83���TG�t���b"O�x03�@'N����'��>����"O
�W.<h\!�7f�!R����"O��ub�'�HիF��/o;�D*"O�� !���E�	��W!P�ɶ"O�8�u!Ϗ5Ѵ�;�[�:r�z�"Oe��!�:!7pLK0��+����"O0D4��+ш��	1c�n%:�"O0 �,�>��	ʔ�>|��t`�"O��8�ME3T	$���.S|4"O>Ũ�NAB���s�X2*����B"O,�CpO��t^�y�R��qx�(�"O^=�'��}�ʔ*��@�c��ps"O�鋃+>'Ԡl�r�E���H0"OV�	���6>ɤ8p,ڋ߂����A�O��d!b��iWNܫ"KC�n���i�'�F��b! �4���@���:9���1�' ͠�AN,ir^5�4׉�:]b�'�d��ǦY�m�l �t����Ƒ��'3�����ǒCoĚ7lL�\P���'��Pce��&�
�1�CG��3�'}4� I	�r.��dW�䲝��'"(U���;Ţ(�F�/[&���'�%�pn�`�:�*��(N�
Mi�'�\MA�	J!��;��7����'��!�Ǯ�h�����'�4O��
�')��Pc(9��\K��Ga�<��'�j!��O��D�(āf ]�ȓ`[>�3�)�*�(���4r����)� ,�$�ʒc�IB��T`*��ȓh����/q�N��!̑�aHe�ȓN��z�O��,��m�#��A�ȓfS���DY�}������ 3�� �ȓno~��6t��śC抙\�4\��3�!`�����&�{�#�W�z�ȓ{�\��P�(H�u�ei�.\��ȓjcz(�BM��M1���c�hL����(��e��0�d΅ �N)�ȓe�� ��̤{z�5�P�Z=�숇�	�С�9[R��z��]�WH���ȓ\���!�( �7�в䢂�6نȓbH[֧����!�.j&�����E�T
L9P�{���;� �"O.��P�%Z���S�g�J�n��0�'1O�-�PBR	}�|�'Q�5��e"O�4 t�K������I��!H'"O��[!�ي;���U�_^�ѡ"Ohi�@�j-��+d���Y�"OH� 7�C�,��� `��H�:$�W"O����w�8	��>hqb���"O��8���m��h`ʗ�VQ��+�"O� VJvŵNh\;3*ĒLP u�p�OL�=E�tG>�L�r᫉�Q$La����yR�*s�}��ƫR��l�dC��y�CȄ4�,�r�"�,D� 0i#�X��yrm�90$ ����Bĕ�"�Q��ybcT�d$�`3��F8"�PG�Q2�y���(#�����A<�'kB)�y2aՎVMF5���GO]h 𱇄��yƎL�D��#ջHҁp�7�y��S��:������%Q�3�yҧ�L!L!��ۇ]�����Z,�yrJ8� �ȖS�>����O�y���u9���C Ɓa���ٖ� �y�(�;H�`���$� �&�
$�y%4O-��o��0���G+�y�Ǟ3,E0��Em&8j�Ö/�yR� �1��I�5k�3Κ� ��ɪ�y��BL���@@��%���+G��y�Kfv4q�gְ+�v�2v.�*�y2���M3��$$*Dc��� �y�dėXv���,��p��'�ل�y�.��I��LI�lN� �����y��'"2([	�PI�����y�*ױw	���D�(G��`�@ǆ�y���,����^/�\�yՆ:�y2��5����#[#R*լ�y��� �h������h�N���y�#	�*7֙)���0�D�.�y����-�2xK���
�|��G��y� ��y�&%��FA8���G�S��y�J��P4p H3�ܫ%)�U;6d��y�T>Nyx�cp��6iQ��i�p<��z��]�A��;C �U��M�!�$��v����������sP�C	a�!�$����+��Ǫ5��@rP�os!��]�'��aF�3�R�Bm�<KV!�����;�ɍ>o��I��+B�!�d�������%�v�TL'HC�H�!���YUʽ	A� ֶ�A�&�!�D�40bL� Ǖ qŮ���A�*_!���L@��x��ȅn��,�E��#Q\ax��k��+�KڪH�����A��qH�B�	�gg�hwLNk��|떆B&.�^B�I<q��걍�'}�x�D�@�Q 0B�ɗ/�-�b�f�hdQ2�;@�.B䉀'(]�GG�,�qc�H�B�	,xP��HI%P�@�?o0�B�	��,aq�J�sB&�����M8RB䉘n�� P�H@Fg�ЧR�-XPB�	��� R�	q���F'N> 5"B䉎 ]�D���5m�}�\��Y+D���ҧ�"�ʰ�v 
<�$�c�-D��ZuNj�5���!�6�Q1
-D�T��T;oX��"�Y�
}3-,D��!@N�j�Y���>%V�|Z
=D�,�$d��I��-:���"��;�<D�0�5�P�(P"�8%����qe8D���q&��O��$�	iɪM��� D�d�BM��F�9����z�l@ǁ�>A�z$�9c�/*@�x��ύZ��\�ȓ-�4�Q�8�F��(����z���:di)+����hM�� Ɇȓ_�V�b2�+�pK$@�_���ȓ?���gՅ!�`ɺ� C�1]T���S�? ��+�LͶ!��{7�ڿ*����"O�I#cFT�X�g)����"O� {6,ԙ�ʭ;ǌVh�ٗ"O2�jUMSQ��b�J�'>Tt��"O�Pq��ĮB�"���	�w1�p��"O����I�b���?`f�C"O5�c�<�r�� X��d� �"OT�����!7&Mi�A���-��"OF52d���:w�5�`�����""O,QQ���	 �Ύ�/��4h�"O����%��3����N�0ʀ"O�H)A��=t����,��iz�"O���`�1o�L��jH-X��L�"O��ș�/y�I��I�?��2"O�P�#D
5���m�4Aڥ9D"O^�AAGH�+:ꥋ�C`�:�"O�d1�	�`���%%U�R�Q�"O��Ѵh҇(�ț��I�
�����"Oֽ���_�Lr���+����"O ���Cʞx�l�Kچk�jl��"O�A
f|Ϙ@J��Z�"�a�"O�	��L�&��; N��q�#"Ob��H� v�m���U#S��M��"O��84�R/on��梇�t�H۴"O��v�Y>�D@�F�P�� �"OnL(Ş1꾥 w&�� �Tͪ"O0����Ĥw�TibF G�Ԉ�b"O���A$�8EF��!Ň�(�����"O��Ұ�X�IK����7��y(`"O�{�mD�'ɨ��"� y�r��B"OJ�ӂe��t[V�ʱaX�w��@"O�xT�T��f�:�Ȃs�&�Q�"O���� ~�S�+�t0��"O�����B>u=.<��k9�`��"O���e��y�J<�E���|����"O�Q�@�N�F{j��$
A���Ʌ"O�}[���
o�A�N�*fK���"O��k�JP���U��i�Q�"O��8TF�3y�a�4��Y�~��"O�x[�d_�:ڄ��$�W&~��MKp"O�1�ʉ�]���T�^$�R��T"O�]Rтʎqa0�04�@�;|��qR"O��X���=XE�]�Iz�(2"O����6�� �ƚ9r�}�"O�4Є�V���@3W�F�P���F"O|�{�i�|�ʡ�$�@4q�""O*xQPn��|��i`�.��6	�T� "O��ߦm~�c�M���X�"Ob=b�)S�l����c	�qլ�Q�"O��E�^��SB�	:G���a"O����=t0,)�U#���8E�"OX8g*�qL0ى���`Q8"Of���.�k���Jŀ�.�HD*�"O�D:��=�ұ*��+L��"O"	�7�_�M{2���l�E4�-��"O��u&\� J,�ABm;�8JR"O�m�*ЁY�T9А��;:xB"O.�k!C;:�s�bY����"O�}��-��c����_��RL�&"O���7ˏ1}Z��ֆѶA�^d�"Ot���o�?o"9��Y�&�De��"Opt��֠�2�SBK���"O��J���<�~���|ޠ�(G"O�9[�$�"�`1��(�;�b�3b"O� ����N��[��a�1��1�"O2���g�2 '��Zbƙ�"�2`��"O8uk�C�tO\�S�C_���Hq"O��"�ӿcKj �'ň�Z}��R�"OFy��蒠�\{a�C�2�l,0d"O�Ej�#_	%��}�t�_�rޒ��#"O�T��]<*�"��#��0�"O����U�s֎}�oO��*�~�<q�V�F��4�e,��8��q@�<��Q�
�xkd���'�je�z�<���ޘrfv��P/L)�H�!co�<�Q��������o��S�b�g�<�����Uӥ�E�f*�3��O�<9��  � #��2W⡹֬�O�<Aԫ��n���'Õ����t:!�$�\�"�қ\,u�УO8E'!��)h���w0h±q㖿!�@��@z��,S$���[[V!��=w/�,� �N�D?�!���ѤwA!�DJ�Q�Ș
a�V	�J �fa�w-!��14@6�SMX�rGT���[�-!�����p��['([ d�A�O!�D�/&=z�@�->H�8ŏ� yy!���(X�I2�G (('V�Q ٓ{o!���H�x��-5��!�GA�3pi!���V�a����W澠ɕ�	�zR!��K
�-��I��x��I�B���!�T<2x*b�W�Y�f<H�%�4�!�䟎QV�B$gA��$���S�!�
!ȪA�A�?n��t�QhƘ/�!��TG�B��*n�0U9�e��7�!�䘷k���Raˏ��b�83n��U�!�d7n;,�*�쒰<���c���!/�!�$�Q�0�rƘ�v@�K��Xj!�d�+}�t�� ��@�i�*͍@�!�������ⓡ��D�2��9�!��?$�P�#B�����D�F!d�!�D9%�8���������Ș	�!�d��w
� e�D�>�D�p���(;2!��]�P	s���K�"�E��*�!򄀽n2����"Z�7@N��$��	 �!��πZ~�Qq�"����!�t!�ą2	�n�zɍ��,�� ��U!��$��5�o�=�4�e
�oP!��B]
�Irk� 	���(ؔ!�D)zyx��C�N�h��	�!�D�1,����vcW�ƒ�Ǡ\�`�!�$�#cS�|�� ��o�Z�!��O�;�<�PaĂ_N�y�h_��!�8AoV����K>M>iF���nu!��D�65�="�O T?�<�䪄D�!��9�� �e�TK X�a6@��!�֦s�|�	6���Zz�!%F\X�!���J�=r`CT "��7e��/�!��өMbr���V��G" ��!��Q[:��0e	�:8�p�꠪X�}�!�dC�"e��͇l�h�Z�j�-*�!�dոq��%�����y� 4�#I��w!���;}@v����%R���J��@Qd!�DU�X. ��5N̳ �R�3QL�6H3!�D��0o�@)���/a���3lT�L	!�������E�\����R_�	�!�D�0=8꽫�&�ܥ���D��!�$�i|� �F��?`��ł,�!�� P쒕iW���\rqm�6;V��"ODܐ�@�)}
�H��.=$zq)6"O� �-8/���YbL�1UB�ib�"OA�4�W"�~��"�L�8���w"Op$�pg�2[� \K��ǌ��4(d"O���T��s��)�)�%4�\�t"O�-E/Κ^�2��Qi��G���7"OH�z���o���KiP�{b5�"O��R�
Qf�*�r��Bi:a��"On Uk$9�>�0���vfɨ�"O6����E}8���i�`j�"O�� .IyX��bK�m�&��"OMZ�N�'[��uAS�Dl���"Ol�˫� �Z⃣N�h��E"O��b�h�`*U+�E��}z�"O�m�"D��S$�d)�v�`�F"O6�;� E�a�L��ݸtl"=rr"O �xC�N����E�rl�Q��"O��[�W/5,���
��'I< �3"O^LشA109��U@Z��`|Cq"O��`2�˴=Xpgώ�Q2����"Ob�a��0M&x(;5n��dKf<��"O�Y����:^t�R�N><�T�B"O����^0�`�җJ�%;�+"O,I(��q�Ve�@LU!Gb���"O�����n-|�8��	���q�"OLp��e�*�Z�I�0n�R�'"O6��Q�)�2R�Y!�H"O*�
�%H%P9j����go:؋&"O��X�&��d�rPB��ufP5�T"O���A�f���u�OxF�X�"OP����Z��+� \�4d�-P�"O�����V $m� �?3XX��"O��!%�:�f,� :QC��%"O ���aߨR�\��m(d0�B�"O�����[�
U�@�˪$�$ %"O�X �XxY�EiAa�,ut���t"O�����&B��܉���+J���"O�3p��Fv�c�t���"O,D�s��P��Y�t�
e�"O �P�O1HM)e,ƴW�P��"O��rQ-ݷ/C.(�P!��Y�B��f"O2��FC_/�ҍ 0]�ZB#"Ox���Fc�^h�p�Vmʲp�*D�{�^=-�0`�g�@�E����u-D�0��bK�`NP)�nߚR�ȹ%J=D����$�y8zX����$�Af�%D�XC���%X$
@��d��g��HL!����� '5٪�g/�m;!��6#jb��J'%�N9�-�,!�$�&ߌ9(�H�#9q��웊1�!��٦by�<Y��(>�Bu��#�!���7v��$⍉1�9	W+�+V�!�DO�*�� �灊$ZI����?t�!�d�LtEc�d�'_�j��񬓬m�!�$ն
�:ڀ���<&8�+��.�!�������)R�Y�ƫR5�!����P��\L蘢�,�LG!�����m�T��"0]�)Sy�!��H(��9qkX��(J0G�!�DM'P���$+�>'`n��H��)�!�^+q��"'��9��Q0�䅍i�!��8oJ���� ,���;�fü7h!���ss&e:�K�9c{~�Гϔ\T!�� �
�"ܛ ^@H��A�v���a"O�i��ǚo��y�&&Ѫ}Q�'�B�P���n�R���Θ�^�Z��'���+���#F�1j���,�p��'Ќ�HeI�I�VbU��6`S�',8ʷ��b��5M�x~q��'/�4Qw��؁QeI��	�'�J��%]�@�R�����L��'Z�a��͉_ բra�'X<h�0�'%@�U�>��c�#÷I�J=r
�'e`m�S$P�+S��hD-��=���[
�'t4QTeŷ`�\شj@�;ߎԪ	�'5�V1es����H�7���'�eN 
];֜HF�1 uPtZ�'��5���0�d9x@���!��$�
�'�=yg��k�Xs�l���
���'����1 J.z>����ο\`P��'�hE9���ڒ��τ�pon8��'>��J� ޷fB>1�Q*�oU�p�'b���F�K �S�"G$Z$60��'���r#lY�*R0�bB�/J�v���'����I��xw.["���
�'.($SU*�Ce��#� L!���
�'�H}���͐\�TT0���7 �Tm)�'2z�c��Zْkv�ʜb�!b�'�ȥ�c�S"|�:2�*ţ
�*H�'Р��g��b�H��E]�y�~�'0L�d�"	�>��LrzZ�S�'��T��M-B�l� �άg�����'+�� �@Y/�����=k�!��'Nf�J2��s����#�?mE�1J�'����ʃ�?k��1P�T�]�ʓ!&�`r%�';�h�S4�Z��ꌅ�D�Р��M�mnHK�&?�ԄȓaU�ݚ��M	'����P!VG���:L����ʡ&�֍(�@!	����|�H]*re@4�P�A&�I``��ȓBY6��J[0�BڕT�X�ȓhM�Tk�h޹2X�K�	Z���{< \�PI�8]����an�H8��@P�=c h�8fv�|�Ɯ�0�݅ȓJ�4)��%8�t�4�$b~������h�LT9��!��O�"Ė��ȓff�(	6H�=�@hň��V ���4z��ꐁԵW�I�P�V�� ��rx.��lX�q��}#2��"=F��ȓ}r����6�`t{�k�\�l1��}��*���
&TK��Ή_����ȓV�8Qt��;Y(Dey���w���ȓ:�ꁺ`D�2td�� o�b`��ȓvd�J�KJ6�|�p��(\p����J�J��$s������Z$l:�i�ȓff�"N�6%�<գ`B$1��ԅȓg��B5�\?u?���JT�\&��G�p"��R�lF�U�A���(\���
�a� �>��d���3d��U��.Nd�#e�Q�(��8Zg`�+
�dH��Et��.[D������#	���ȓS�ZL�f�Y5�\ٱ�L��U�.���1T �l��
x<(� /=/���ȓ.R�Q��� 7.���O�,a9̆ȓVW|�$*צi�f�S暩T8���uq`�MZ#FTV�Z�N�$R�p@��Z��� @�	�"�zCdܙ ��E��S�? �0!�F;��Rh��0M�}C�"O����B���C�֭02&X "On����C��a�)�4��"O8���P��4Rч�0q[TQ�c"O��I$�����u��	�ּ["O��X��ӚV�9�N�0���"O��y�;Mt�ɒ����ʤH�"On�k0��":v�cUdR�BW�i%"O�k ��k�I�!d�9@;�tp�"O*�!��<#���<+���$"O��i$ʇ�g��V�a�8�LD��yB�ߣr^��&��+�p��l���y�D֙w2��2�A�*s��0!�>�y��޻Z�rP�� m˾�2�A��y���#����h8 lb1A�;�yBDM3W#b0��@n���SE��y�C1m�@�
���R?��*#GG��y�� G<�C"��ZD�������y"ҩ�)Fc��(������V�y�	�\+��bw�]�'�()�f��y2"��{[8D�gK�M�� �+�y"�^fO@�
3f
݅ةyC\E�
�'�	����1:TE��'5j�l��	�'<N؀T�Q8e��5� $gf�C
�'D����|D2��`)Ӫ�*,x�'7R�gFG�{�D@�n�*(�r��'b�9�ӊA*{n k'�)+{��B�'+pS��[q
��Qb��rqX�'l���
O.|]2ta�G�]�r�'�,ذl�1+�����<`&���'������ �H~�$c�IW&C�IW�`҂�*R{Ҙ{Fct�<B�I�~��L��
*�XG��C䉴>��Y��)}�Y1!����C�	�}=��1��>��l
�Ѐ{4�B�I-T�Bbu�
>L(�p��3�ZB�	x:���/V�����F@��.���D�5
�r��6b�>M�X��ST�+!��V�)�S�D9�<qɑ��1�!�$��J�(d.O\L�!� 5%�!򤒬�SK]���A .ʐXo!�D����|BF:;˸=���C�!�䊜5��x��k�
ze��P���!�=~R��ʵ�C6�W�]z�!�D<D/<��M��F!�(��[�q�!� 6Ӑm�ң�6	����eϳVv!�֔��qZ��´1�p9B��%E]!�ě�e���.I�Z��0vh��jG!��[P��Ĺ���3���S'�cK!�d S�@3��ܨ��'˒2!����ؼZ�hQ	:�Z�� �ٔs"!��x��I�D�B�+�n$BG�ǥW�!�$��W�M�s�їU J1a#J^�p�!���-�>i�Ơ0Lh�s�N�!�D)6��1)2��9 E���X!�$X,`�����H�7�8�b�F�,!���2+ud6*n�5�cͩ�!��:
Q�C5c�j�+Z�|t!�d�3s�$�R���I��Ꙥgf!�$1O�b�Bg�C�H� 	S$3!򤔣}�j-�`<p���q�K9l�!�Prp����� 0��-�I��!�_�=ӌccBF�!���r�A*?|!������.N��`$�M-ou!�� �K��	���)��ܱ+~$�"O^���ϊFĜ�����{�"O
X�`ɉ��PD��,�'�2Xr�	E>1`A��Uh�y���>�kg�'D�Ӷ��*�d�1��.(Y�Tk'#D�H��I�n�R)T�P��9��5D�D��<y�<��kή�Xn3D�����BvӬ�y����7��F�+D���O�Uv� ��B�f�-z/$D����C��Pa�3�@�V��)�0D��1��o#�(H�g $�`�
S&!D�p+4k��}s �݉xњU�d! D��I��[��p���LҢ[&�<D�D�����W�\���A�g��rc�$D�x9�Dݺ<�!�CJ(�z8+/D�,+T_�"�D�K��H�\J�M���?D�!&�D�Lm���%@�rGF�y�*<D�\����9>���[��Є4D�ph��"X�rۣI#@�����1D���N�vTE��Ά3^\���*D���s\�K.�T��h��@��6D�06/J�V� ��"���(<�s�3D��`B�3�i��F@�K3�\i�G3D�<�󈙯9��N�
+�����;D����&5 i�aV�״
�2�O��d�O���9O�c�,�V�0Yf�Q�e&�[c��)��8D���P��/�(�3'$dPu���"D�٦�-;����B�6��E��� D�X{��Dg����c�"���c�#D���d�:�-�S�R�*Wl�x��?D�|i�	�R#<ɓ�##Y�{U�>4��{d �1h������8��3�.�_y"�'�r�'��	L�'�%���[/h]���#�<fS�-C����'v�>�I0g{��X�I�m�<�M� ,C�I�|��F"y+����5_�C䉺J*$R�'�8_������ UbC�09��E+���%e��%���f<�C�
,d�f�OzǴ���&tR�B�	#$�h�l�9��2�i��gd���2LO����@�6�>�7cж}���"O&Q��(XW�sQ��/P�BP�"O�8 4�:�ȱIp��  �8�"O��rK������0���v"O�˒M!��-;q@]2���"O ������ҁ* �=�,x��"O*A���*G8�X�s!Z�4�d�)E_�ȅ�	�{���8.��L.>`���F�T�C�	D.8Jd��6o��T�QA�4B�	q x�0��_ҹ�T�#G4B� �j�Õ �)l�x�e�_$�C�I3c�4�` f�F F����l��C�ɉD�촃F/�+=_l�q��L&�C�I��l(��A� m�S�o�/W����'�S�D��ѱ'h  �,�:����e5u!�dHP��)1��n�.H������B�ɧh�)C�dd֘J��S�8C䉣�\Y�p�٧h�f�c`�O�tjC�I�q��S4%�2	�!�ś�W��B�I91H&�Qc�*����٢(�ax��o*n��2�$.�z� � �#*x�Ol�=�|��8]��E�d��P��I�7�;�0>��ET~2�W)�X�T�6dܘɐ�U�Py��I� a� �j�J<\�n�c�<!��\�d�I�啑�zq@Hc�<� L��!�ݮ`ǘ1��rʴ]��"O���� �a�̱#d�-p�~�T�	ʟDE����:P���g�:i����%��y"Ǘ�_ ����Ch6��,A��0=�uN_̓S M�mO�?����#ТF��d�ȓy�6��c�U�a��U��늺?T��ȓ(��L��ӆ3쒐1�gU9~�@M�ȓ>���1ע3XdIa�Ʈk�l}�����òGE��IyD��F�RM�?i���0|RgK�]4��r�&�Ś�*�Bx���'���9��)w�T�Q�l�M���00�ץ�O?�ɕI���dM�% �c�ІL�:B��0��Aaf
��sp��d�C��C�*'0�4��ʩ}�l0�倊WN�C䉄Q�>Ԙb'ȠH1��� nI Y��C��;4�H���;|ޮ�UeH/%�F�OR��'LO:�r�X�Ҧ(R5�S	����"OFk�''NVak��Q�Y��܊��'�O�q�!M?�Ӽ�'�,X���
>^p+�)�S�<��`��H�`'JO�E�C�Q�<�����RH8{A B�6%c�e�g�<������nq�%�ʸy��UK�(�X�<q`E٫0I��+�� �3��	Nx���p��B�V�.�%-o�l�ȓE����9��A�V��+��Dx�*I#�0|��b'}FԘ�eE��>:���a�O�<yШQ�`s�X��Mų4������XL�<	�NV�&��`���.H��@[�%�O�<�ş)J��"�P�AP��#�(Pa�<���(f�؂��T'lU���f�\y��'ؤq���A�fK�����4c�|�
ϓ�?���?1��sS&�X�B� &l(�L��`7�����?�
�#�jy8�ʇ�s���1��m�f��ȓaT����
�.�d�W�
�+�@��	�b!ؖ�CR!�',�iT�H��"�d͐4L�?���ڔk��o�Xh�ȓ2����s���ӣd�(9%����ɁC�ȕ��9�4��B���M����d�O�D�O����,2z� �AER�p�`���9$B���Ob���՘��܀��j`���r'ڸB�!���_(�����~NJ3�¯~!�ē1�>��j
�C6-Q�A�+_!�V!Xnt �W�Ə*Qس�`@�hD!�d��X��ӖM�;\�(�/�9!�$�1v��<b#��7�p0�(_�!�y��'��' ��.���&i1�Ą!��D�K�B�'�X���'�I�<����&D�<q�L�2�LI�l��yr�Đ�~m�S��!H��ǭ�!�y���+@�0�띑����gn�?�yb#�!y��k=q�j�n��y�(�1.� ��@*y��@RM�"�y�N�$
��r���@�Ց��'*az�#�����ӯ�'<�	��U,\����y����	�'e~�YHФp�4��GW5G1VC�I�.�
�#AjʗB���#�0`NC�I  Szq@�e������=%��B�I�J��(�Ż���C�Ǟ�>��B�6@����B�3V��!���jB�ɍ'������p�����L3 F"C�	�^0�tA��v����!	�>cG���+�	e��~����9�x�;�a]�B�X7�=�y�BW&I1CM�X��Z%.���y�-�ܜ]Ð([�f%��hŝ�y�IB�Q���(Ӿc܌�!q�У�y
� bd����\��A0%��x�!�S"O2 ��LǠr ��CC�M�N����'1O�����1�R$Ã�L��\�4"O|�ȅc�2�g���ft��"O��:6C	4N��a��
>E��k�"O8eچEB��X���	�zH�"O6|Bu�D�U���ɝc'"\!�"O��B �Ԑ,���
�?i%)��"OT��6W|��[�$��"ON��6�.h�,SrfK*TX"p�'�ў"~�uL�!4�Z�yW�"C�=��` �y�*�Y�\�9�FïG~�Dx��p�
�'F�h3V�\9(��Eb�#��A��'��t��[��R��:Te��'Ƭ�{���-I6�� �M�|�<p��'��!��˔;IN���%�EzR���'���c��z(eK�E�40�
�'��h���;U{P8�#�0ʬa���',���<�����Ɵ(��)�R� C�I	nEV���͸DK�-��e��2C�I`}���7����|5A���,�B䉎i|L݀PƊ1,�Pm���PQ�B��##��Wޢ�T�c�bס�" ��'j6�YS+@�=q~��v,����'Ny���T��� ��pLJ�'�ȭ�� �=o9R��tȉ��F�+�'ۢ�
J>3�*	�E�O�*��'�"�2��ϔ�YАBy/�DZ
�'E8!ICM�rIq,�m-�	�'�n��h	�	��a��g#Bl�	�'�<Y�G�f 
��S ,�h<��'��1�
�J\̲fˈ��P1�'��pP�'\�-����DI��'�����+�U(���B�_"����'d�	�f�Z�2�zr��Qc����'����skÁ~��|��KQ){u���ϓ�O�"��ڤ"�d�B�P��}8"Ox}q�N�H��j�@��
���"O����4u\@����}���A�"O��+1�	�r�n���ҕK�yy5"O:�i�I���Z��B�	�x����d"O�� ��^�v�j$@Q���"O����P]���ƕ(�0y��	̟E���0b9F�Fnm��@��y"��0����lN��zq��@��'�ў�O꺁�&@�)�Lp�g^%�dD�'��=�qJJ2o���/R�!��'� �x�M?X���X��R�f��
�'!l���M�i��\:�m!}]��
�'��T��x=�h;��[=]�qA���'JbI��Z�G����0G�[z���'��	��]_�|Y�@�U!U8�����D'��	�� zx� r�@���8�"�'!�$�[����T��^�Xa��K�^�!�DP{�j"�E�f&�]rW-O�2�!�޲.�Y� �
1&��H�L�X�!�D7Bb��3T��<=���x�W�+��P����I(p!� 
��P�)�� 㔾~t�C�I$O�hTHV��$**>�X��$M`C�I�=�~�Y��OGp$��A �� C�IO{��C�H�n�@C�
T�6B�I"+���@/��XTcՐNh�C�	�H�p�����r��&oH�a�*C�I��l�U��)>$#)%{|(���O���� h3q�H�t��A��!I(tR"O��	5(�3��@밡7?������s�O�졲� �K�L�#ˋ?>0�H�
�';��kK�
*sr(�ҥ�� tJ��
�'n�)�2�$(Ԝ��3��%��K�';��3�F�|��9JÇOJ��'I��{&�����&(f� 0�'ޤ�B�J�h�8��7&N�����hO?]��@݇
�"��`���]P�Q�i�s�<��B$��@�F=<MB!NJ�<	�H1ax�����N�v=¦�l�<��g��S0\�p���*^V�)d�i�<AWD�w3��ADޙbp�YV�_���hO�x���Bƽlծ]��゗~����C���t��  ���b̅�c�ȹ��Y�����JWiU$H���4�ƾ$ִ��@4D���$bŐ_�X�)E�Oo�h�c�4D������xu:ă�gA.!:`���1D����� W�E��L�g��Mk�0D���e'��>"����iG:N~Uh6)D��@H���X�hF1���a�!D�4R�o;@rR����e�H�(�O˓��S�Op!S�°#���&�P<o��;1"O����A�B>4�T�=r4��"O왑.Z7KQ��4B��wZ"@*�"OQ� $U5^���Z=[Z
\A"O��g�ל!�Q
a I!9q6ͪ�"O"y@��-2�u��O�.DV^ D"O��p��)M��I��B�hW,H��"O�`��a1V�*��0$0^��"O��DG.'O:���_N<2#"O����F����bK����"O�p��	�tp����+�:���"O�CԨ�<6΄B!,*m!�t�"O8��S�T����LT������"O|2�<E��"����5�☪�"O|R$O�;A���qI���I�V"O0�:'�W�5��Ye��*p}x|�A"O�����@�*©Z�F"io� ʖ"O$a!)b�M�!����P�"Oxm�7��+n�Ӳ"9�B"O6�[F)@�/�4��w��V'���"O��mII0}���
	}���I��|E���
΁�͒&$��!c�[��yR�V9��� ���:Gn���yRo	�4?vI��
Բ%��Ӄ!�7�y"Ĝ�]n��S ɝ	�:��cR�y��4a9�yj ��9 D� ��̊�y�k��oI�q!V� =ru��WO�y�&R�VL��8�N1n���ևO��y"�E]��%�@b�mkh-`Q���y��hTP���	�d2�����)�y�+�?�^|�"�Z�]i��Jާ�y����00l8��-T/��
�쎊�y��R�N���EυJ��;�+�y��
�Lb�}H�%�Hv�X��]��yB��������&
�N{~P����y���)>6����Pp16g	�y\�}����i��|:dsŉ���y�/�L.
BF
*{��1`��yR>�x}�dz�̥I��ʹ�y�O͛65� sC)] �EXV���y��X�'%��r�$�Z�D����S1�y�j�p��93"͆W�m���y
� ~܂�L�<Q�a8��T�7<�0�"O^u��^,��wN�u$+5"O�m@���J�	#w��;9�~m� "O�ȃgM�BM��J�� $ƺH�#"O�H1B@ R����Gu��uv"O���2D',tՠ�,�*{ަL��"OjP!���(32���_�*��D"O�4��J� u��Q�q��A�]�TD{���?94�K�m9/� �nһSxC�I�o$X��r���6��*eE��R�nC�I��8��VJڒu��]xRk�ITC�	' �P��d.�1�(�1� M�
�6�OZ�$*�)�t���ӫ �-��&
2�C��Ku��3�.F�-X�`��jv��:�S�OZPH4��AHT��*�Έ���|�|�R����x�$��>Nr��7OS�f*�}��E �yҋ�v��q�DΓ3N���4���y&S�w�&��'FZ0��  I�y�j[�;,��,�>�����''2�O���qU�܄�r�s��v4p*�',��;�II�z��gEU���`�'�A�6�B�$�Ժ�ؙa�*���Z���	؟@$�d� &
�h�j��e�%Y�j�h�\�<i���[m���֪��?A�e81��Y�<�u��Zɖ5��^�
0���Z�<y7�0F�bD�F��0\zp�f.X�<1$��o��1�Jh��]���U�<�Enŧ#��a�e�B�>C��Ii�<YD^:-�r4�����uA�H�Zx���'{�I�o.�8 U%�"8{\![	�-m�B��$|��ta�I��jV���S�[. ��C�I�p�y;Bm�q��2C��Dx�C��#x�h�j��P�^�����?F��C�Ƀ=�ܬ����c}�����ۄ%�C�	�cw��	���3dw�E)�Aĸ��B�O��XY�֍X�tI��D j��B�I�.� �E @���H�L�#�BC�ɤI�1�̹`f%��S�C�
#���;eJ�r�^���'N0C�ɵw�$�����:;4�[q-E"��B䉭j�j<��Z����C��.be�B�I�k�H�=Y��Pؖ��8�BB�I�fʡp(��*Ġuc���p�NB䉽	����� !JY�qۗ��M�.B�	�S^�A)I�&+t�"T�ݗ| B���Y��$lbp��H�.1��C��<b���h�>�c��8Q��C�Ɍ�"�(Ad|(%��.#D�C�I�'����#� c)����Nҡn��C䉅>8s�Ο֤51�]��C�I�}���cI3n�4Ճ���6B�C��0�L���H�v�q:F�׫,O�B�	<S((��-�o)�i����d�hB����E(��
�n��I�����e{B�/Lr�k��w�^%�vk�	��C�I�T;��:Aн^�*�XT!�	�C�I�*�ؙa�f_�mT���ԭ[���=�Ój�����:QnM�섑0�J݆ȓZ-�hS`ۦ�Pi�lBJ����>�����&E�h��bN ����A-&U��d��W�����Қ@�⸆ȓ/�\��ʍ6D݂�pub^�*�Q�ȓ"|$�E!�jx682M
S�F{b�'�ᓻO�RȰ��k��̓�
	�MW��<1+O�qO� ��S�E�!�.$K&��4�b<�A�'4�'��)�3�ڕM�T���/'V���&Ԅ�y"�΁	0�xD�D�'j�3�"���y��ngl\����(+؅0�⊗�y��q�`�xF�K�\��8�y�I4OҌ+LVxQh�O��hO����O
�x�TBۣ9�¢�A' ����4"�ҟ���M�IO��O�l^�C�<�&8
Qd� ;䰖'��'��>��:YZ9Z #]�uZ2E�QFLi^"B�	y�Q�G�>�ix�m�5.B�I�z�b�0�J[�6;�R�'w��C�I�+a� IS���I8�K!n�1��B�I�ii�d��E~!"��Z$����d2?q�K��~,*����@�$!�Gy��'��h(�"@	%�0E'��Z��e`�'�$T��)��8��$�E��;����'�x� 㓢}y�ƣ�8G3��8�'�ԩƯ��$�Fb�CU\���''�������TC�jԌJn6d�
�'�Y�>5�P�k%Äݾ,�ʓ�ؕ��,�',Y,��RiƀQ���ȓmmrH�F�ߤ2u���r�9i���ȓS�-�cT������%���X�ȓ挡�Gg:�Z�G�e�ScXI�<y��L�kO����#[�cQhEr�E_�<��T
A�Ђ1G���}Qr��yrkā�@Jf�S*)}�	�1$ڕ��>)�Ot��÷��!N
`$�5�V"O��w��MJ�Űĭ�18;F���'+ ���� 3��V]+^�n���'��\KP��(�lȲ�l�X�tq��'�D�� ˄[����c��!U-��'螺��䒓�6)т	Y7M���	ߓ�'�����S%���b'�1S�r<3	��'�<�I�T�o8��Mts
�'3$[C
ŕG����
� qu��	�'L������Hy`(i���a�ҥ0	�'N���G��g���ӭܴjy��	�'J����J9{ؖ�k�˖�c�Q��'Ռ`�v�ԧ/���bǀ7m�p��'&�����dN�|�#��c�HL`���O�"|��#0y|8�4�`��Iч�^F�<	񮒜�^�I���A���I�<�&��9R�4�ѭ��
�R}�V�P�<���0 m)B��3j
8Y(D�g�<I��_����f��.-x�{�L�H�<q�\�1pL��.�&1h��KR�QE�<!��1�r�*��b7���T�]g�<��*ϋ�ni��\��c�y�<Y�@��0�H��(PT64hH���x�<a,:p�Mj��Y{`��dr�<��Δ�q�`�93-
R%z�*��n�<��"T�~EZ�ǈ9Mz�8a�Kc�<!�*M�!d��� ڌa�:��f�\�<I0�Ur6aqƇ	N%�f�L�<��J��_�A� � {l�AY��E�<A��9a��X�C&s� ����y��;{~9c5o�3�8��#�y�$(_ �:��$zx�y�d�;#�0`�ce�'j<�l҃�Ԣ�y��5�Ԡ�� &`2�e�v��y��ҺB�P�*A�H�%�N��F���yRM��#1�����s�����O��yR�2'����hI�W[Tp)��6�y
� MAfaG���Ay��WM�q��"Oԙ��o/t@�v�O�.�R8�"O���a]5AX!P��ҳ"j��!6"O 1��Y���ؙ�گLJd9��"O��0���0���[�e�:l$���"O`��q���U0<9���/a;4���"O0t�����$��p"�˄:����e"O6�U@�T����N�s|��r�"OQ"&h�	07���P��Kg�Y;�"OR8hC/փzj��p�˗AqXpv*O6(��@�.h��x%��/�z� �'1�d�S�Rg�xuH� �:'��2�'D]�!CCC�Ӣ����'���%��&U��(�Ad�=���H|�"2&.��p�5��<ÐI�ȓ`��y�N�$P=¬��K6����l��@M62��M�]����ȓ5���2�k˝W!�m�T��*c$���>J���3�Lk�t0o牜u���j��E-y�`y� �jM�� �ހ�
��2)FU�� ���\��2i��:��K0yR�c����*C�T��"`�@����8����T�k~z��ȓn�H��VN�*3��35`8x���ȓp�Ҝ;ԉ:'	�H3����]�ȓ.�� V�M�p���
2ތp��$3:� #a	7�Z�BTMP�+En���Ѡٲ7BH;jކ����i�f(��s�L٠���{z-��F�?:t�ȓ[5lrr,у|�L<�b��v��ȓs�^�1	V��1h oԍ+M`L�ȓGh�s�D �@&��3�����[]�!S�H���8�B*F*yf݇ȓ(����t���y�ハ� Ү5��d2��;���Lư���R�W�(�ȓD���R�KP�(Ҁ���x��L�I;���&�f��b�[�k��9�ح�7�ڧ)aN�0���q��ȓb5\�b�O���I��8h����
�!rw!�]��v�O(���W&����]5��;�E#UeNy��E�j�ɠ��!W�ZM���Һ:4��\>h�ː��0!<�*f�ҶkR��ȓ8�|�Cǯ^��1єh��<���z�����%3�Q0%σ4M*�ȓ3J4䰱h�_s̈Q�יzl,��G�Li��v����(B�`���ȓմ�����h�`C�ﶍ��-F���0%%}��!��׸_y���f�R���D���R>��-�ȓrX��Ə ��ݨ�e�1KD����5�2�"�oñr���x�Z�fT�=��&��i$���( �U�$��f�����l�P��j"^E*���C#]�ƙ�ȓr#،+�ԥ<����%I9bt,y��h؀8K"oD�:�@X*u�ĠP0��f<\�R�f8f�"�ȓ�<�(%lXEd���`'�5S��L�ȓp��Pg�/!0-H�H7�|d��G�:	�F S"_�0�B�{����vy�5���X�r�� �Uh0�!�ȓ]^`�U��y)K
?)M��?�m���#X���@�,�vi��|�ٳ卝�a���-�0T`Մ�S�? �@�-�p�)�)�Z��G"Ot�䊙�g��I��-�^��X��"Oh�)l�7oq�s�Ѱs���CR"O�KU]#����fƌgd�a"O�#G�
�*<\MЅ�� f"O �3�b
{٣�Ŀ	!J���"O��lœ*io:YS�$֢Xj��W"O�q2���#�ܰZ�P�iR �t"Ofܘ�@���ʂ��#�bI��"O�I�u � i@�,�fl
���"O����N 2��[��;Jxy�"O���ai� ��AB��
-D �"OJ���o��D��	�(��"O��DW
}lyӤ��
	�J,"O�ms3#�eBE�
UH��bU"O�Q��)3XM<� mBoUJ0 "O���	�%5<!:s�:s9Vhy`"OH݃�Hm�����&$	a2"O����暤?�������Kg"OX8��E:>�>�2pj{qI�g"O���c��V����
� �@��"OFe)BKT�tE�q	b�%�$ę�"O2��cH�F�6��B�RN�A��"OB���'R%'\^=�@�!^��E��"O.A)��4
R��Tl�e���R"O��@RJ�c�pM5>�^"O�u����	X �VV�s�ܤ���R{�<�4�C�|[У�v��9�⭘u�<����;׈�$��=;X���Ko�<��M4h�2���偔�^�
�� n�<�&�6(lm���v�%��c�N�<��枏Q��ik�G��|�\yC��<!`'�.(��3�/V�^��}C��Kw�<I5������*Uj�XФ�s�<�C�*2�j�`Q0є�����r�<��̋r,�=x7�ɺ�� �C��s�<�c���c��Y��ӹ> �3��U�<�+C	K��h�F��;��S�@Q�<�"��2:,F���З5<�h���w�<�Յ[�\�D�FfNI�,�&Gt�<aK�O5>�ٓ@N�q�*�xq��l�<�Q@Z�'�6	Z6�
$�2�ԊO�<y��Ɔk�\ubT��[��X@"�Td�<q�A��s6-BF����i�6�_�<�P�OKt�����#�N�R#��r�<�m�x��B	 M�ag�s�<qbƇ�D|�Q�;>�\�Df�<�4F�F��4V�@6p�&cf#^�<�@�Wi��(B�M.(�}�P��A�<)��S(E�rM��G�$�ze�X�<�`��.~���eT-Q��뗮�n�<qnߤ������#�]�+t�T�ȓH��M(�W{�ma�׺����ȓeN8�2�j\
L(}�7�¸fmJ��ȓ<����� �$<��y�]�+��E��	���t�
8Hy�%������ȓ"��ǏƭX(xyҁ�ה�l�ȓ6�|�R�hN���ha��[M�D��xP%(`�]�嘘�'��]���eZn���kZ�Ji����ȁ\%����W�V�S��
!n�xq�çK��\�ȓ�����"�����ũ,p��ȓj��3��3� ]�cU�]6���)N���T�58�X��@�y$]��S�? Hi��A�KH�AIs���5�B"O�L*�K�8o�����ET�ԙ"O�h�4�ņ4��`��:�R[S"O�h�w��1W�R1�����\}�3"O.#&=���������˄"O=0 � ��t��E�?�xܚ�"On�3�̎0��kp'֪=rf��@"O ���● ���'�L!XXrT���'!�޹<��i�EG��PY��w)w'!�Dηy��t�L"�t5(Ĥ��!��
0i*`��
S�j� �"
)3]!��L\
2&��2z��cA�ȓ�!���;�.l3�@�tC� S%�M�(�!�X���rn��<M~˅ �5Ka~bS�����<��٦KG=S��Pb)?q��uT�-C�xu�`E�I�v��Ixy��F�����eO����x���yR/�	���� d^�
d��$a@��y�a'@K����Ĕ� ��|ـI���y���gux89g�=K�,aB�*��hO:��DR2^�H� y�=���t�!��~��}�Ƃ��BZ�M��N��&��O@��5�W�O�2T��c�;�����	D�����N����uc��C:�ha���%$!�dE�U3F��nG�Y+J���j[�@��=E��4k3Vu
Ch�� p�\�b0w�:4� �D��4� ��@�
�z+���@$O���*-�ɸ�t"P�ӹg�p�pMЕf�B��7lk���5��Id,(7o�59_��'`���3��~���S�Čm1tQ:QC��>�K��'$��:@��%#�07]>Q�7��Q��O���R�_�Iͬy����q]
�C��[R����:�	�!$b���ΓE�R"�h�(4I�C�IJ������@�l���B��M�˓�~���~��Z���5t}L�೩�	P�B�	�(f�J�ٗwW� W�Vp�p�O&��d�/.e�c,��^-�x� ;)!��bF�A��c*
�*�/F�+!��1��L��e��!��m�ю٫f���`��:�L�^�b�s@��^�VȠ�\�ȇ�	�>C���e��1<��ER㖶_a�C�	�%��P�`�K�aک05o�W�C�	:A@��ę��|��WԻ]G:B��6?:��!��5�@�D�7"�C䉣J������Y�|y7�,0��$G	X\kBJ˧yh���t&T<1�a~�R������yo�e	��J*{�T1�DL>D��򅏨(x���ʇq2M���9���ny�h��r�ؐ�jR56r	��"O��(.�7��D!5�_�\�Ȉ�7"O&��0�C�erf��)�,�����"O�ЫT��q� -�D���&�d���"O�*e��ǒ�:'��g�LQ��x"�'t>y�w���Xy��#&�U/uXv%�	�'!�9+pC�0S��"aD�d7�A��'�M�7�ی<4�Y{�:ː��	�'���Pѯ5hj��őx��(���hO?U��o�>#������:��3�`�K؟���Ew��X�v���+�K3q��=��"O2Ҵ��Sh�͠��n�.�sr��4MY?�*��¦q3�$��Ȫ?���B7D�\���%FC�}��/G��U���k���S��|,�R	ŕ\�vPJ��<C�	8X���(�F7[S�C�� T:C�)� V�2�"_�����M�&c��x%�	F�O7j�9 �Z� ��X��T�o� x��'\����.L�xr���U%�k������d;�Q0��0�6��,}}!�d��X���䁯k6(�"�
�~o�I~��H�)�0'
��-A�J*.<�آ"O��2ņ*����G�e'2�63O���g8����&W"q��Cg�"�z��)D�H���T���⢈�3 0"@�<D�\�Ѣ�A?�4�A��t��鄂;D�`Q�Y�"Fb�)�d ��8D��:��Yq�6x��jW*I5
���7D�t3���H���:�*;&pYB* $�,��E���LH(�>9p���E�y�	?�V�a�0Ԟ�@��yo�,(�"Y�#*2�4��(�MC
�'I�����?n[Ru�Q�I�Ap(}��0�S�'���E�[�p�� �G'L�C$�3bX!���JjD ���S:�@u�M�In��6�I��HO��]�~��\��Ս��<���,o�!�$�,��0�Ah�4&��Ma�Nٙ�!�Dz��0�����8*4�C�!��Cb2�;�aZ1{�&���.�y�!��'+�r����	�d�F���g���[�����`رe߆�Rrh� U�����I%�O����OPH0
;7R����D,;��Ti ��L���=��I	��2L������j#>9W�i*�>���*D-���6O�'h���r� D��`��9D��H���j����\F{��i["vJ9���'/T��� !�$#
��I��&-f�`��d9�A�	Q����ˣT�<� L<hzVչE�"/!�dL�s��Di�3^��bUC٤~.�FY��'���<�! ���	�6\wH�`� 1�8���^}���7T��.��>ș0#I�MsO��O�Ϙ'Cj�АiT?��M�����c�|���$Y�O�>�*��
7��-�pk�'g;���'���� 	5%��!Cό6[b�����x2*�{/f�F%�>^��`eE��d6�Ș'�!�קd���V���I�l��'�=�!)A�r4(X 1��	v��Ɂ�r�x���?g�ڹ�6�E�Z_|�s�e���C�I�h�����Y�T�P�C$O�^�
6M�<�M>E�ܴ2~hB&i�v�xX:$bK�(l}��U�@�h�M�r5h1�5���`9D����R�1�c��mL�Ѣ�Q6����@y��E&A���H�&M<q�4�'�ў�u�I�E\���2�%D�T|!�Ă`_�B�	�=�Z���2�tP��;(�@�O2��D�)4~��$BI�V
���"Oa��O��%�'"�!���#s"O�����=jf������?o��Pv�	V�O���ƫ�:l>����+d4��'��q�J�f\(�#q�U(*��D-OmDz���I�dh�a���F�$��B�Y:��|�g }�+��o��!p�IH�΀���E��yb�K'3�`��N�t����Ԧ�OT��D�Oz��b�ɕ�uJ�S���3p�#�'͎�p�ٙa	�(��R�{i�̃\�����i���*!�g��*F�*���yR�Qq3�Y�pGC	,���$�*���䓕hO�nA��θ8ң�@�MjwN�T�!��G;8� ��@�i��ȓ��uߺ!���'�ў"~"����A����,�c�#4�y
� �@h�o�Y-�����B�]�l��i���26IB#1T���CJ3[!�D�J
��o8>�yA�"�!�Y5s^)�O*L`p#O�!��Nl�xx6	A�Jhi��,m�!�䟨=k�4�鑵|���+Ǣ��I�!�ĞPd�����]�`K�!��!3��3�h�p�������={�'��|2�:*)\���5m@�X��<�?A㓁�dՄid�1
�ڷRij�s�-]�`�!���RI��jTL��5C^���<���9�ɫ���(�ωR�B����J�JQ�B�I�<���[R��(/�(���
�a�n⟈D{J?�#�O.,�ݱ�-�+<a��P�%D�@�b���@�K��[��j����$D��Ha��%�<(ۂ -\�&eh�`-D����i�=#+�5 �\6�d97.!D� �/S5L�,qE%>T8��:D�1�aQ3K�*m��n<6��<D�X�@�Č:^����$0��-:D� ��� �R�JPL�0���P�6D��!i�.u��������� p�/D���w�S9U��Ux-�0��S�+D�d#� K�>@i��[�p '.D���(i�<86cG� �1�'.D��qq So������lK4�X6N>D���SZ�-���¦�Eol�r�O.D���Q�K� !���!/>���'D����qo�h`d�@/y�D%��K�<������9x���E�&"|��:�%p"�Y!_`p��$��Rx�ȓL	zmq1�D�
Ոfo��d���ȓJ���I���`��9��8fl�9�ȓ"b⼳Iݦ.�����09� \��w�� ��
%8@��E-%�B<���<�!�a��^��˲�Q�6@ꕅȓDM.�[�.7c���A���ȅȓ\�Ȕ	��]#���`H�z��h�ȓ_z�P��ԃ�)�.��H��ZK.���! )|�yr3�Kx�l��ȓipp���!v�-*���&ń�%�����(e^�!F�� ���	|�Hv!��Yyּ��S�0�ȓ"���]i�����G�@&��0�6)�Ɩ�S��P�g��k�}�ȓhp�|��ƇE�h,�D�:	�Ԅȓ �"��4�D�T���#˕�
/��p�Ƀ�IT�3u���e�BU��	�OhVi��o�7Ѻy�dB׎1�C�	�6*AD�g�pY��p��C��^X�]3B�4�I�lC䉐G԰�s'L�!�`���� N�C��v�Ջ!@U=~lQ�j@�Ww�C�	�!�N���Y�`[4X���@�8�C�	�q�~Qu�4G�0l2�⒡P��C��xw�,��ˋ�+��x�W��`C��1@����ң�v����w+�QdxC�I�-N���j�!������nEDC�ɛn:l��?9Id���EV}zRC�ia���_3�`в`W9{�j��S�2D�T�K%nԼ�b�#��6�����6D��k֋�do�K�G\�=q�HЃ2D��`��=��M��N�!��ie�7D�xr��C	1�4<����y0l����4D�t�1'�z���91;�9��'<D�� tH���П-B��B����SÚQ��"O,�{G�ڨi�"�b���JAX��W"O�5#�M�d�^���mC��"O�u�N��HC�<��@�Z ��hq"OND*���o1(*v��1Y�r��C"O������"戳#��
ɶ|�"O��P\
`9A��x�L)�E��y�KO35RX�ӂ��f\Ĉ;e+�<�yR�Z>c��CUoX'R�
�`T�,�y"NR ��UJu%�>�����y�a\&Nj�8rF'(j�P[󮛮�yRH؎=����"�'p�#2��6�yR�ٿ;r��@J9��G�yR���1���?��,;A���y"�N,L�\�)�c߽ZoN�Z&��y2`ыj�z���G��^�B�������y�I�xL)���7]'T� F�(�yb ^�iC:�ɣ��%B��j�LA��y�\5}�AE�:E2�І��y�I���Cd�4D
@[�A
�y"�W�Aj}��_! ��){��B�y�ޒ/̺���G\(t���QS�%�yf�.z��f+I�Ƣ��[��yB�#�@�"�	?'n\����0<7H(rH���)];]�rP'ˁ�'�3�(D���,A�|O:x���_y��(���<��)�|6���K>E��"	���}��mn�a�@c@.�y2+�H٦T��� �7n|d� +�50��5j�А�!אhe���'��\J6(.+M���!%Y�O�D8�	 �]�$�Ǔ^�b�s��x�� ��W��d��I6�O��Y@Έ&�����!G�c��!+��ɃqM*h��=�O�,l�Ѥ˳>�j�� Ǜ�^�֨#�'�:���5Rl�i�OA�H����O�ɒ��{�YjL�"}:篑:_Lx���Dݱy`X�Àz�<	�՗3S61;cKީu�d*�N�7��I<P�,����.��g�'Z�KvJ)8'���Tv!^|`��J-$]уԩ��S���q["&�&��`��K�T�*��� #�o"[ �A!������)�a�!P��� ��O�Ll{#��RL�Q@Eݾ*:d=)�'Y�̃-ǥP�(�1'�E0|&���'�N	�ɼk��M����s|e��'���Ї���WW����/�#t�y	�'8�lr�0YVj�:�+�36�	�37�
�coӞѱ�/�R������CdH��"O�Ppp�C�QS�!��E#���	�9�\h@�ëPR>�� ���q�:`����>A�X ��� D�Й��D$B�H�e�	]y̹U�K��LT��5!_����'^�>�	CiR�j� ��T̈Eh�*FآC䉈|eޱ� ɿg��Ш�7�L�wl5�GB�qf���<O�p$��F�(*�/�=Ox��r��'$�5���Ͼ\	V�9��J�`!$�C�V.��e`��
��5
O4 Z2�ük�ޠ�t��l3��j2�ă6Nx-�%ѐu�E�f�&�O�"�It(�gN�������
�')��:p���sh�S� �"��J��.!kw��;FhH���*�(��	�]BRMp�V2J	�q�m�&6%2B��#$p,�+
	%*�T�A>-�m r�G#	�����R#���<.�iD2��-.��ak݀p�č�(���0=��� 9o�T  T��t.�Hidi��iXx(ۤ��uKP��E����Q�,�Dgǌe484��!­Q�D�<����,R�hsUӏFb�`�3��+�H�����f����%l�搅�W���A�b�(1�(@�҄*�`I�/	"��rs��Ct$A����Uyr�.�Xpg^T`e���,�y���7X<�<�r���uH�D�T���Κm��cI�.�A1G$�6N��1��Its��A��4(�|�!�L*n�j��dڔE;ܰ�F4E9��3� ��)��x�nX�@h��2�����dFKhP�# ��3x�EçI�bL���> �nZ�i�>��@�B-�� �`��[d�4ϧ:杷rVeb���)��Z���2C�		�R�"�[�fߚ�gkӭ��P��e������s�2ݪ�@N	�X�
V�[*dڐ�wk3?�p
�)~�Ĺ���V e�Xx���B�:�Z4��
���r�`� 	2t*ׂ5����b�'��ღv%pӑ�K+��ɵ"�� � (hvB<)4K��RyВOF,��Wq�|{�J	2��6펈%�l� %�ϛhCB��&ʛW��L2��ŏm!f�0���nk�B��n��2`�[�6��Bs�*����V�/��M1�/54@�Bi��l�� ꛖ7�7�F�	S ��;q�H����!66�&��8U��y��I=N�"�����But�1�E�%eo����L9[�Y�GF�bR
i"F��.�?��ePDzl�	f�P&ce�O�����6 E��	�EM	,��]"��Ɂi�Du; DN�W̤���&Ds���hF��b�'�5F���ؤȭiR�_8x��=⇥F��0=�D��<d02���g��4y���'�U?��Ǭ:)���S��?D}�L��!0x�'?�ѩ��n���`�@�~�L0넄[�N�5I�F,D�T���C��8y��c��,s� C��$*6��j�i>����犐3���O�x�<�cRd����m�0f���4
�_���*�'N}D]pE�4G��B�"�>U�#�eU�\S�O �&���#
�a��=���=���$��EY�xG}��w�ӁZ.HO6�y��7`��Y?~d^�( ��H��H� ���D�!�D[���IsCF�'�*��悓Z���1��9��M6�x���M����|$��b�^��i��^���%"O�c�Ď#s�̛� S�'��k`Ł 9�X� ���H
>y@r푾W�g�=��\ ��]�EJ�%:0�u/t���."~���b�&��	2��;0�9�@�.+2oڶB�x3�'����DA�B2B<��˂�_�tђ������ ��
Mj��5+~>�x���!��y1���8t@�A�)D���-d2*��	��~���)#ʓ�<�+T� �d�1�rț�Ԃ�hűW��C�$�
��%+�I1v�X���zI�6-�2�`�#\�-��'��Y3��/��q)1��!N�0�(D�DAV��X-����3�u�[��j��1�|b�;�g}�ڥ"TZ����֡~��d���7c��Y�=aC�q���	P5��2���/�������ЕcX�0���2�'1���T��;(p��D�����m*K  ɠ����C�P���?M��D���Sǅ��Zȸ�E�jgay��K+|��!��^y� ��x JM#5�ͻW�䰸��W���'pR@8'�]���G�4@��0�2a���E����E� �ē(��AV����
Î6��ibFcD�%�����	��5��1#f��S��(��	FLଋ­��T���v��-�11��Nz���4X0&��~&�T�3��(3�E��
�=���]%=��R���6=�������C�R��IlIr$J_!s��d���1��@��ā,J�P�{����y2�P&SN�Ћb�
;f0M
�����<�G%�z�H�Df�<�O]/d���ǧ�\�؝��[ܓO�Ę�s-z�x#~B����Z<�6m��x�"��p��_�I�_��u2��=��?ʓ)I/p�c�H�$��y���O!>��4��|��/�g}ҡ��5�"�ׄ�^S�A*��B�*^Dp#�>��Ç<Y���'����So�M f�C�E �:@� ��?�R��$@&�O��	�ḑbxHa"�� ��"�W�#E�Tz�@�%��>�phȈH���{�ɵ��P�ƮvX�,���h
����]�,q5�o�� ��((l��A�8D���!�e�5CGK�	Q�� sf�3�dW	S��4SF�3��['ˀ�V0��ëX*�Љ��"O�b�A�aZ���UȚƈ%P�Eo��=)� �V���d	E��!w��^���۳��0YP��9	V���I����Q���6�p`�� ���d� Rq��k�'��Ij ��X�)���&��@��'��z�*���I0�VA�p�J>A��@�t����!��'9��n�e���=	����5�̠%�Z��$� �CU��"��D�1i�:A�=�Q%S8V�@�S�IOeܓk'�>���^Q&�3c��6�j��w G�Q�x�E��0qLp�I��@`4��P�:X�l�;���٦a��P�}|d�a)ИQ2 A�hZ�o�@�J�ʬ¡!	�G��ҧ�i�51���'��#���5���b%��{Ԥb��� \�b�)ϤlX��W��e7x8e�>��O�.�v� ꘊP�ODϧ~���e�B�&(*�Y�y�Ɇ��~��[� �<o��2שANax1�� Z���fOJ�i �ۢ�Y��&H�\������IU���	PZl1��<��Ш��P@$#E/W�,QҦ"OZeх�H�*��E�v%��g5 ���O�E��l÷.�,�I��}�Z�9ܘD+Jp�`�&'g�<Y����bm�$�7ǙR�hA��c�D����̏��0<���^����1�Ow�,e�KS؟tyB�ߦN��R+G#B��
�华P���A	�{(<���@�Z"bU1� G�\8�(�F�'ln��u��B�'�FQ�A�X�Bܢ��V#D�������{�ң�lJ�J<��(�ȓQX&�r �Q�J�3c,3�쌄�Q(�m��H;�`KB�.�&,��nd��F�\�Lؚ�,��B�����~��H����#x�pb���	r����ȓ;���"c��:`�u����&�"y�ȓ&r(��+�c
l�x��?cs���� �P�4�^d3� D�8'�ܬ��X>j���n�E�xxA��;��=�ȓ:��I$��I��A�	ּ��o��;�-J, �]�Gt�5�ȓ#U��A��٘2<܈a���N�h,����Z���$n��la3�ƿ?�-��|=�@�W�K=w�� G�J��0��ȓ[
����C04����1e·@���,��9�%L�1i��!�u�խb�ڌ�ȓ�>�ۣ(�U�֙�'C�w��Մ�E�F�	ef�:��i�a�^`U@��Q���BS�L�pL��.�/2�؅ȓ)�X�S!"id�������'}hm�ȓU7����]VILUI�ϩ-�1�ȓm�n%cA�Dx~�PM�'n�H�ȓZ
6	�Ɛ�LQ!�wJt%���g6�`��F�Z���J�dl�ȓo_�=��BX3l9�U���l��ȓc
psdӞ�L9樑�x��T�ȓO��cr%��r�&�bU�=~f��A  �4˜�)��<���2Q�*��ȓ{�$}�vB�1����&���F�V��^��@Kp�_�H"�p"���A'����!��L��.ɠي�J�"����q��QeB"s�zt�ggA�,Xąȓ[j�L�Tg�%Q�z� �Q p�&!�ȓz���)�����
�Paߠa+̥�ȓ ��,�`�ŸS� 00�ݛ%}ĩ��qA��b$���-��;Egؐ&8�ȓZ$��h$钟'�蝃1�KkB1�ȓf���)V炋N���H�WՇȓk0�q�bӯyB`��J;c�T��lFީ�'�_[��L�*v��P3�q��dD/V0�A���B]d<�ȓf�1�"x�6�'���+Ԝ�ȓf'���`�=6�̊uf��n2>���;)e����}6؄��a����ȓ#�@�QT?$�V�+�jܻq��ȓ&��%ʃ	�� ��u�N�0n�ȓb�Nx3��ʅ![��!D��.5�.9��:�XB��7U�I!��і��a�ȓw�PP�EFƒwdJ�O���Y�5D���a=6��X�ů� ?YD���0D�([��V���3� ���.]��#D��+�+͸xv�U`�/	 m:�D�V�:D�� �a���إ��@�%�B"O��Pa�), �K�O+:�Y@�"OHQЁ�:ZĨ1��º*T00"O�H��nj>���呜����E"O��Б�X$4��qz�@�RRȴ�T"O�D��Ga)E�q�W�8���"OjQQGԵ��h���V�zL��"O�:W���*Jf^ .�*���"O�#%�M#68
���
=�U"Ov�H�'�+e�&TR�/0q�f��"O�,�ѩG�V�|]b�,;�j]Y"OIDX�0�R� ��@s܁�"OF�[���,�B�B�>
~�'"O�=�� `��CX�R�Y"O5�6a�0��K�+��W�(U�"O�q�"RDP�� �gA� ���2"O؄���m3�@�f��=�xm�v"O���m@��
����R�*l�"OB%+0O�tE����M�� f�I�"O���Y�Q�E ����l��1J""OFp�'͡5m(ԪC�-9��f"O�i2�AZ�Hr8�j���8 �숙"O�5��Bҟ_�(!"��\���C�"O�xk�EJ)"�h�� 	%Ҙ�#"O���pf��ʒU�D d|���[�<y"�ړR���q6څ]�p��'�V�<1CT26(&@��CtkECFP�<�P�Ԁr��Љah^Kw��aE�D�����N�B�qO�]�7>�^Ͳ�		�����"O���"�!1NaZ�ѰuD����Q�d���E��%��|jg�(u�,T���ȓl���ȓ�C�ǉ��%!�'\�%A�$(I��c2h��@��aH|�>�s*�daZ�`�@�N���g��e؟x�4��� �bЂ�4�吅*�;/@��B �.�2�E�nZ��C��d���'���O�h�"�_��9;H~b����Jn:Ո%ʞP<"]xG.WE�<���/%x�a��K<��M1 �T|}�k�:T�mD��@�铍6=Ҡ�����0 0�)�v�C�ɱ	�(�`#@�aԔ:WSR�O<�y���1��4&>c�\p���0o;� i��K�I�x�$�/�O 큐B��*|4Yq�3L��p�Fחv���� ���?�"	(��< P�,لm��HLH�'�R���@�^21�"<�#�Q�0�!��x��"Op-��)
�@� �A�G�k�(�"O�����,��k��.�.���"O�@�󊐘C,�( �4���P"O���a�J&jXƌ�G X�v!H�"O$dqe���*�C ���-hX��u"O�̉���>K�r�Q���8���T"O�4a�l�7�Ԃ�aD�1)��9d"Ot�{��D�LMj)bsb�y��R"Ov���i��l�̩ڴ �*=�nx�"O��t��K���@�n:�69k'"OR�Ƀ�	4�D�0�-�Q�`4�G"O18#`����Ӆ.�8i��-�"O"��&b�k��Y�a'#� �
�"O���&��.�q��&��
�f0G"O�ɠ��ćNfmSq�]�b�!s"O��yGL�!|�Q��2(����"Oj�RW ��_��	����r�ܩ+s"O萺P��+?=�0�Ѫw"�!�"O�A�`� W�� �F�^�{&t|��"O���#�Ϻ\�h5��JJȣf"O�4�4-��w]V)���]4�:���"O� qp��:xYF�XB��f`2���"O셂�K�c���p�`�'Ͳ��p"O�b���q[��#!��!�6��"O-@�n�=XR\��ɧt��}�d"O�ay�f�r[*�19Ħ䐣"O̝��:>}����o�8^_%�8���&��I�a�Q>˓W)�xhrɌ��� ҲlI6bxX�ȓm����W��,x�!�uDL1v�"P�&��;}2 ��'[�^E���d��G��ӑ�Ctaʁb��UNx����*��wfƕR���"����q�� hu�;iG��^ R4J�I�<�r@F3M�����㛰hD~�IW��E�	�jBn���W�+p�t�]o�O�n�C&�-�l��N�=m/�1a�'��q ��� 5���B��Z��u����#�=2���*�1�e�ޅ��'��'�	 u�+<J��Q���
�B^$h;P*�"7�\�04��r�؝rp�߈Ah5"�)	F4|�Y���azB��n��d��F7S��ٛ&#Q?רO�&N�7Cf\S��?j8
��OP�oc�cFi��9��=�wKYZ4��'�4a�)�	D�1+�i��H��yB�'[F�`r�سH��mB�̒�o�$P��eH�O���V�?�N4�է�7F�$�C�'F�r�f]���Eٖ`ݙ4��9a�Яun����ț�nέ)c�����6*�1O��y�B֍{�`ű3)Џwn$iPC�'�L+R��"����c��:�"ѱ0�Ԏ òT{2����EN3Jq$!דBƖ��`��,�6x � ��4G}B��.:��R���Š	0	;t��>EP�&�<?�����P3hp�d��"O�|i���\Tð�Q�{�d�k��O2��d⛄(��L��}�#�|�JY�N�d�� O�<q��
14���ޏXK�)����a�d�=��kp#���0<�P�@�))�#�HG�[�d�S��v؟�6 F�V!s��=L���	�v��[�*Ur(<��M�B��8 DM�2�v�׫�n�'�J��@P�$<�5P�$[�y�(ё��^
q+Nć��T�
T�S��X
��
(�Xl��.����^�)�H��Q,�=Vm�ȓ	�9Q�l:M��@�̕#���?�R�Y!;�#r%'VSW4����Rrzju�3(�l�<�p`�.{T�2�iڼ;r��F����ʒg5���a���dˑ�d��P�bH`ѐ#��'v��{�S���	18R�0!��u�6��т��P��Ӈ��ն�p�M3|OZ1s��no0	��'M24I�ǒ1)��&3�q�]��B�Wx(�I$pcF`!t�7��*���򤝻@��8�e�ʽ��D��A�����C���!2@RqO$�/`�ڌ�	
�`0 �M=U{�5��D%C�'���+�L�N$�HE��j
�{�8�3�	U#>d6D���W�����gj�?��	/N,Q>�;��*u�IDl<��&��|4���S _���ɶs�|P��L<�C��:�H�A�(D�(�<�� Y�:&�U�c�1�H,���7H� ���ś�`P��2�(�;g�8���NA
S�%#&�	3P �(G���1X��W=��
�V\�z��F)3ay2��2#�0�����MyH�p|MڒΘ:=��%Z5�$��'��*��E�G��B��B���|���^(R
H�I<�EY�V�,���%��`� ��e�7"��ti�� �(�c_ԒO�D��O��ʣ)R�~Q��@��A'r8f�8�.?�&�'�zЀ��#�3�$��>�ʭ۵͟
UY��	b/W���\�\�����ɟD�.�)��ԏK�JE�ݡG�f냚�\�d�'b
la�HJq�� ȃJ�n�+˓�4ڄc���E	�����ƹ/������'����ȓ@=��&ON�=j��ه&���'���ǧC������S%6`	��G�x��\�Fˊ=�B��!re�E�$���Ƞ30kJ�+�2G�\j>�o�\��+
0Z�)�f�,�J�ȓ4��t�kC���sf@?v�ȓ]�k�f�0��s\<Y��i�ȓ:B�u` ċ Y��˸M��%�	4�K�Lay�H�s��S�.��3fhș��?1�C�3n���j�(e�1WɁ0#���ѶbƟ�Px
� $�SՇ�r��Rc��cB ��9Tx4��QGO(4�1��k�J��2ߨ��t�~nDQF"O�hb�l���@a�c�=K� 2�O�|��J�&�I:M��}r���mG��s�b]��5�Pe�I�<�΋�s����#E�gD�ɳ¢�K�dŐx��e$�0<A�/�kܜ-Z�7Μ����p?�%᝘{v��(�BJ �2H)�'ѬkU�A��X
A,�B��%,&�y`��ǏLL�qB�a�6�>�2�@�f��$.�/��T�*I��H8F�I�HC�	�8:r��OCGܙ��6-i���}:�@��""�S�O�����&J]�X����f:YC�'L����cE;Vޑ`�"P��"N��3w �F���[U�'Iĕ�'��<_
����їK�,��ߚ�5�
�L@ǨңC�x��v��R�����'R ��a,ɞ��xAb�^n���;����%yr�:������AY������k�R��L-�y��Ja��SHLT`y���ވ�y�!�2�a�Q�T�H�Ĥ�i��y�Bɦ` ��%,��K � �䑻�y��A"f�`�� E��'[(�yBa��4��x�'M��B�"�$T��y��P�w"��R���&zSdИ��y	k�t�c��B!i���f���yb�,/L���ީ?N����yBA	�\��Q&���d 	��"ڙ�y�!S�oLY�2�'Z��p;eC/�yr�'��es�`U8ڠ�`%�ܶ�yr!�(f���E�Ȅ?֦�g�̘�y�<�ހ*g@E�y����Ǝ��y2HLX��̳Ņ�8uLc�O
��yN�(I�/=P��vnWPN��'aNpy���(t �uc�PH���'�P���ީ(X6��KM*-��'*z�A1�f�� �S�Ah
Ȓ�'�V�k>��=�Æ�nL2���'hd����?�v�RO �r�~X
�'5|�j�'� �$a��G�C˚�

�'z��!e� >�H��A��D.@�	�'�>����8�%A�qdj5��N�<���ǄO�L(���U���N�#	�'�z�F��s��U�b�{�"�Q�']"1*3�KAd ��wa�6&j\�
�'�B@�`�ЁV�����/A���	�'`�p�B�-���'<2pe�	�'��m2��I�c�}�uL�L|	�'���c�F�s	iƅ�9*�-	�'M���%��LP��`X�>����	�'B�Y!d�oLa�sEF(-�xS	�',�#���������*Vb���'�^���gF3eJ�]�U�'=�C�'D50`g�}�����!J��'�!Y�˳ϐ��d�#|�8���'0zT��Ą0����F.�-1��(�'e��A��M��| �MQ� ɣ�'��l)E�9q�v�A��8�B�*�
�U��cשFS���������o];N4��z�&�_�4%��8]3`�J�K��b�ٖ]RP4Q��OXX2��U��ᓺ!x���b� ����0�	@D����2 x���Ѹ��Oy�(�3G�)5V
lCC�[(B�2��� c��Zs���4eqO?yBt�ز%+�ћ�+[����ŢħD��)S���O�4\�#�_1� ���Iع:�"�k���'�*�'@�`�����������
�V�d��<��*��V�f��(6�'<�)z3�&\�(:`������'�4劐e��kF\츴l=�'u9z�[��І<���g� �S�θr�-����F���y��;��*xz6�Hr�UNc��v �)<���	C�0tc,�)�'�� �0p�-O���G�h�|*�H� �X��/��)�^%c�$ �D�U2R� _�:�(���fJ OFqrA�)���`3��+��th�@'�b�H�|�# �'�`�@�O^B�x#d�%C��I� M�/l����+Oɺ6�ô!���n�h��򩔫�dd��� �I�'�F=xRH�"pm`h^��'�|�����zW��q�X�0G��!�� d�+w$�y�'�NвG�к'������S�F�D2��WdM�^�$I�ҝ>�Ï�$�M�<����9w���(�0<@T��J<G��I�D ���}����h�tM��j�,b9 �cծ��y�m����O��'�ZXb���Pk.KR�ʃmX$��'���`�OG$�h�C�!��Ԇȓ0ؒYSS��-
J�6͔" � !��'��5��R�7~�AoJ�m;tP��'����.��1��,1���������'�f8�ԃz���宜"�:P8�'>�&�7e$$`HUk��4���'���#b�,CuޕB�
̴e��B�'Ԛh�̙�N��ġ�叉}�.8��'��e����2hP�@�n��'B(ikD�X�8�2[��=u��8�'5n� �/'�l�U��*|P�9�'yQ[&Ȋ����+u@`�'��T%L����BN� h4D��'��DH�eӁw|��Z����J���!D����,� ��c2�F�f��@�"D��[p' 2� 4ir'ڳz���9�!D�p�&�Y3$r��%��.Ӗ��4K3D� !4��=&Q~L���
gq�(���2D�TH�l��
Q���6k��.Ԥ��5�:D��[�*/#,��dG�=��k�"9D�dZ�(8|�i
E5\�Zؐ��9D��kW	�k16���&3�0�6�;D�$�$�"���#�
%�^�x�,8D�,Ǟ.9\I�q��������4D�4�׏�,V2Iɒ�gM�(k��5D�ದl@Kii!G��Ul��{I D�\�%�ж���B��8t�8��d>D�@�H�:$���Q����YW�1D���4�*��0 �⍸r^f�a@�.D����
S,��­
<q>42.D�`9��x�ث�d�	B
�q`0D��0U!7�hiI�ON�HՐ�.D��1��;C��P�m�t^�my@k-D����q�"a9��N�QC�+*D�H�ڂ�C����R+�,b�x�Al:D�(�S��F�>��$#K�r�~��7D��n${������
<f�� �S�5D� f#ɩ]�|�r.J!l*�5D��(�ϙ�}�lpQ��E%,���ц D��bc��[1|y1t+N�O��:1�!D���b�8ab����M��xc��,D��2�P�?g�݋���8jn"')D����,��ī�̏'w4h�@G'D�!mM"}j	{�J�(t���e'D�4�%3�VP��
˧,Z�Qb��&D�@B��]w����	5��a&)D�ܺ��'�%���I�cո�Jg�'D��:�)N�qO��q���0bZ�81V�&D��+f��y��٢����>fV�ɴ/*T�x��dE`���ڋM8B��v"Ov���-2~���) ����"O�J������������5�2"O��j6��`qp ���5p�"O�@�׏�%b��xx��B-2��Z�"O� �1��c^�zQ
s0m��k"O���Q˗�j0��-��AI Qї"O��[��ļ$��`�,�ҵ7"O䴫���{�n����G��0��"O\@�F�ԓc-.8 a7*uv�s"O-B�k6غT�����PjN�8�"O���a�	����²MƆ�Z�"O&E"�!Ι)F*!j`��S�DL�"O.�S�M�v��"��
�J�Nu�"OJ��k�x�l�9�K�(I���y�"OdyC^9a)J�caAϺ]�|��"O(%oC7A��݉�����"OV���G�4HPލ`B`X��0�"O�]x�Nɔ_�N�(p(� e�x�a"O>āt�P�g��5�T�P�.r�٫4"O��� [	��p3��Q6O�B1"O��U�F+M�b �e_�'�pt��"O�U�&��{М���CF���q�s"O&��8A3z�0p�ќ#���"OVuj�\�$H��H��V(�"O�����j6d܁�Aȑ=�d��"O�جkc��wk��r"O�H#�fR�.c���O�74f� `"O�|��FR�9g��u$�f"OT���\�L���3/J�X�
 T"OPDS}_��mܔ���a"O�����4t�A��:K��"O�+��3bD�p,�����"O�	����2��S�гsd52�"O��ɦ!�$U�,8D*ٽd^v��P"O$	��_6Ea�ٺI�8Q�c"O�@����Lp IH��7,�^�t"O^�:v�¿3�R���O$3��YK�"O�yc%/��(��9`��Z�]��tr�"O���A��63�LA��ÝAQp��D"O���v�K�l��ܡtOG<H���"Oީ�"�_n��R��2j�&L(@"O^�K���X=
l�2�@\�-�F"OF�I�?)�V�c�;iߒ�§"O���A�+Tv��[�*�;0�(@s�"O�8)��R�^5R�pʅ 5`�]��"O��k�jȺf��'�c3�9� "O\=9�$�d#��q��4[���"O�@�2#�%V'�A�+ߜ-�셈�"O6����`��B��V�w�.AÑ"Od-ˀ���UE��c4n/9pJ-�P"O�T�3�N3��L`�"*n��*�"O@���'Y���]����-jڽ9E"O��P/d�aA��\,]�B"O�����lX�Y�Î�W�T��"O�B��7�T���`\\���"O�����-\��#ρ"3��@"O�p���*|�BXq�����թ�"O�1���;��5"�8�"���"O�EPq�N�=��l���º����t"ON���b!h���{�#X�Ζ4��"O�g"�	���X2cJ:-�	$"ONuaV�X	���a�>q�Ѐ�"O��@��P/5�L��A�ƢRV�%��"Of��2�� �HEH�.�QR�4��"Oj�q@'[�)g x�a�tH�(p"OX�1D���)�x���cB�)�U"F"OBD8s�[$Z���#ޖ6�२""Op����A�N*��eI8�"O� dys�)�Y�Z�[u�=E䀲u"Ol���
X%E�H��NW+�A��"O6mp CR�CQ�$�P�M� �(P�"Oq�&��� =���%mJ<(	<1P�"ONh�ǌ_2uP�X�ɫ�� "O�]����/Ov>��f�4$����"OfU1���
Q�"���A?e'��"O�ES� :j�85��+K.�L�� "ObĘՉIw�xE���)�Nt�b"Oh�O^5O�n �w)R;3���1P"O.����I�k�aQ���}xV"O2=z����ZH�"�I}&8�7"O60��k�[s��I'��N�<�"O�HD[�}��0Aԗ8�֐�3"O�`cdk1	T�=87`������"Od�D�e��բ�.�L<R5"OJP�Qʒ�2��yd�Q�d�!RF"O���vD� �~��4/� ]
�"O@���f�"(�!HU�"�TP"O��+�>L�ћr̃:MlZY��"OZ�PG�I��dH��L��S�ّC"O��P���.Ana�k���5"O�t�FoS�O01XcoYb�<�a"O�y$��:y$(�� ę9,t(�ٶ"OԴ��a�N����� L>9"O�q{��X#/���˕(D.8x`96"O�������/N*�Z��A�R��2"Orx��ե=�$\�&,@��0q"O<�E���p��EJ��5�����"O�Z��\�d��xxt�X�u��kw"O�� Ώls|t��(�3v�"=��"O&��U䋜2fx�*�d�����$D��k�ͷv�>�H��_$��$�#D����K��R#p-F6C4��i�d-D��j�K��F��5��DB87� ���7D������ ?�e���	$Xŉ�� D����l�B�V127�;nvu�Q�#D���Rd�2Xa�ܠ�/`�F)� #D��0�IN*s��0	B�^�U%�HRà-D�4���.B{J�8qϻ"렘X��7D��z��PGl��t�O�X��
3�4D�<����c��۠�N�h�ŸqL1D�H���źA>��8s�0%-zep�C.D��Ib�V"*�I�ToH�E���c��-D��;��F�T̤�Hr��Xuf��E�&D��+���5^d��P$�8w@���1D�sd�ҹ_�z��N�R"��� 0D��҆,�,� Mh��K e���.D�$�fi�<s#���$�]�N�X�@ D���Tk��IC���Bg�>��1R�,#D���K�,��� Q�U����B5D���#�Т#J4He�� P�s�k3D�� �^Qr4Q����&�%3��1D�� g/B��!N:[%2Pe<D�|9� T�T�*�˶Q�~Ж 3�4D��ӆ"ϯQ5"DzB���h��2D��` c�1*�x9��K�U�<Bq�/D��Jp�L�Y��pˤ=K���A-(D��t��m���P���~��:T�3D� ��\)2�8 g��`8�+�n4D�����'m���q����X��@K3D�x٧'F�g�����"9b��rE&3D�<����.��H�RŖ.&����$D������H�f<�u��=�%H# D�� :�Ivn��m뒽y�ʔ���}�"O���c�ǧ�fx��	�(� 1�"O��j .�&$��$��L�Y��"O�`{���^`Di�r�G>+�$h(�"O���
l������&�H��"O>�1U*�.(#�X
dS�8$X�"O��Y��W�f\
�d��*F@�۵"O�h"'J�%�j�F�" S�"O��0��W�O����:{�D�F"O�����L�
�����P��0t"OZԓ�JS(�a�E����"O� %l��T��"�`�+%x���"O���j_6hra@*u���?D��ò��;�^ �Rh�	=8m9��0D�l; fO�*���;� �/R��B�0D��B�k*L�5NU�M4�20D� 0!�_'`�`�FU�=�LCsi,D���"�dN�0�����g�&D����ΌDƪ%����J�j4�sb?D�p{,��Y�J��=%;�tV	=D��S�C   ��   �  f  �  �  *  h5  �@  �K  WW  �b  �m  �u  �}  Ć  n�  ��  ��  N�  ��  �  D�  ��  ۿ  2�  ~�  ��  |�  �  U�  ��  ��  ��  P  �  W � #$ �, �3 �9 B@ D  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1��2*Q��'/�ܱ�Dnٲ�0�rG-E�ws���ȓC5p�yaL�!	:Xy���J+K��X���N}BI$�dH�ѮI�4�S�[��yb�_"`3�a1�$�H��5p�+Ϝ�O�"rl�$RB&��JW�z����y�<!�c��rrY��/�t/�u�e#Cny"M+�S�O�t$8��:���ӇԢYӮyz�')�T���܂f�l�Ë�Oې�s���x§�)9��Ź�.
r}\�K7)��y��)�N>�͍�_B�FG�>S	���r�<!���5k��y�h݈��`Hqy¿i���&�S�D�ˑ>�����F6!�ѩ�+�yB��$�xRP�K.~Z�CK;�yfΥK��p�&
�ۼ�� K	��y�ggd"|�ãY�V@�P�Z��y���� Vb��aӐD��Q�������c��"<E�D'S!&��L����
Is�UAO��yrkǴ�;���/���tH��y�:~ls�	R�(���)�N��yRG��U�X,�d�!�*}�Pf��yr�gq@=)���LÞ4��G �p<���8����ԓ�f�	6 
T�!�$�9-"�"P�3��D�ׁ��$�!��B/�haB�88�L��A=gU!���21܅%�O��l �7P!���J鸜@��%��@��	��w4!�Ěe:b��p��{�,�I�D2w!�d[�-N��AҖ_KtP)2'�h�!�d
-r�ZP���0I��9��Z�!��H�s �^�v ¦	�!�D�Җ��S%O�`�9�V�Ҩ?!�D��\��i3�O�Ih؂����_�!��U%0����HAzTXȐ0aP,R�!�D�~�$0�%��|K4Qj�@��!�A��4�Jt�"3� x)�O�!���b�ѡ[ t��{g>�!�Q4 �F�"wőjrN\���R��!���V<�
c�[C���P�J=Kw!�Dξ9W�Q��E�|������W��!�X"M���[�sHȄzDG*T�!�V�@uمʇ*�m!F+�!��V;������e��"J�_!�d��)�j0�V��QВ�
�˵q�!�B:�nQ�Q�̇D�T���MZ(}!���t�}Y��[�:���Ǳ}n!�dE�1���l�>E��#0tW!�$ �GҼ���HU�̘0b221!�dY�b��
�,�!�ڜ���9�!�^�:�D|JT��K�m3�@�g^!��>[h�QsG�e���p{�!�� ���ր�$OK�]Z�hB�1*Q"O��@�08��ȓ#K5����"O.4Be<* �7�Ȫ�n9�0"O��SD�I�#��;��=ڄ�s�"O� r�xu|�[�/K�*ר�ف"O<@�VV8y�P��$y��HzF"O(�x�Ō2gd@���V�3�v`+�"O�V�E&\h����8|~֠��"O ш�C�NX�����e�}�"O�Y�wm�*H���C�ei��[%"O��Bb�  �M��C\&VP�P@"O���ŋ7lP̢1�O�$�|��"O�<�+ �}�^�i�`��*9K�"OTR������G���Y���$"O��{����d�͌]���@�"OX�Kŏ�56��A�D�0�&l8�"Orܪ��έb��%�S���iia"O�ᆎ&7�|��Qܨ� "O��P���_�D���=n]-S�"ONP�t�\-6�=HR�#Hĭ!3"O�[��קBy�a��`��)84��"O�,�6i�v��������"O0��A��"P�a�� ϗ �r<�#"ON��D��ą�����T�W"Od�hG�^b��C��.L���"Obh����n�$��R-�.wb1�G"O8uA�,̎k�D�%��ro<]��"O�)�T+J:Y1:����ªT�[�"Op�K#�׾4\ʔ��8HB� �"O���S��'7��Rtm�^�j�;0"ON̡�o��%Ⱥ��&�N�h�Q°"O
�B����qZxl#�k��KA�31"O���d�ȎR2�1�,�%	�y�+��X "N "�B���yB��=hq`D�[(K~nQ{��9�y��$e v�a��2Q�0qi��ybc�2N4��cF�$�Z��aR��y�	�;�� ֬�%D��b�g��y)\��lt3s��a���X��y��S�4hA'MG:z�@��5�ybJ�?Q ��o21Ëն�y�U�/t�٣`�Qo;�4;��]��yr%6c$c��d_q�A�B�y�Cr���D	�Vy8�"N<�y2,:p82� g��*�֝B�C1�y��9fkL|���Ͼh�>��⮔��y�g	�Ґ�Y#����@���yR@<O���7��+5x�X�F��yI�
k(��^���J���7�y��(vH��`�I�Y��d�`�&�yZ�1���%F�K5�u�T$٨�yr��)Ph$\���=2��h��;�y��/�H8s��ߕ'���`�щ�y�-����P�%>"�z���Ԥ�y�ͅR��%�)�`D�����yR̎Q�Z|84��k	}K�˲�y2�.  9��+�c�}��E���yb�L�@�T\��7b���ɖ��yR�
�t�E��"�6������yB�W� ��A�5oFz��˰��y�B$h��f"�%��1�L��y��'=�v%zt &�R,@0)Z��y�+�6Ы��U�R(q'!B��y2j�!
w�eZ��D��zq�ݿ�y
� @k�N��:*�1�Aͩj �-� "O��CE��7!�VLbb�ǿ�"Ud"O���#� h6��!`�+s�yH�"O$ȡ`�@<'U��d���'Fm�"OjL)!k3+6�쀡HY�C��ت��'���'���'nZ>�	柌�I6:w�M����i����?+�n��I���I����Ο��I͟4�I����ɨd%��7�J�s�2!{A
1sib �����������՟���ڟ����(���m����f�
��jQ�>[�\�������I���Iȟ���ϟ��������)4�HP
����0�h�Q��%AI(�����\����H�I럸�	ǟ��I矀���������T\�t���]�fW�a��˟�����矨��,����H�Ʌw1tc�bN��2�vM�[s�����p�	ϟ���Ο���ҟ��	���	(E��p�Ŧl��k��$DX����ß��I�� ��ڟ����T�I����1ް�M��>����r�,m��ޟL�I՟��	���	�`��ʟD�	�!a�((���n~��P��"'�Y�Iş�	֟4�I�@��T����p�Ɇ\�D�a�9I�z\�Œ3=�¬��џd�	۟,�	�������	��InpM���s��Yd,��S�Fu�	�d�Iܟ|��֟$�����	��\��0�:i��Iܲ bD�"�#o6���Iɟ���ڟ$�	ߟ��Iݟ���4�?���s1B)�� ů�X�B���I�d�S�l��wy���O4n!���``��X>�Q��G��qc��)?Y5�i8�O�9O8��E�DD�$1eiſ(��ck����O�\��`xӄ�����O;�e��X�"�|�P+�1��}��yB�'��	D�O�  !T�G�8I��p��׆%5��8#�e�:� �$9�S<�M�;r����$I �$��Hc���*� #��?�'��)�ӆ,x��m��<��Y�qVf���υV6��0�+��<y�'�^�d���hO��O�y�AJ4�kQ��L*��bB:O�˓��uV�&D ʘ'�h20,�F�@���B�����$�V}2�'��8O��"Ş!�O��j�D��Pr����'�reǒ	�X���tE�ҟ�A�'f3��ѩ$����B�λ
���Q��'��9Ot}��j�5���AK��(�`��0O��nZ�j�?���4�.�ˆ��"&�x ��/w���K�0O(���O��
#%�6m#?��O�P�	2\�\��DI�M��k��OT���M>y-O�I�Oh��Ob���O��A�eX2*JH�ɑ-�		���׫�<�Դi>��2�'v��'��$'[;.w�ɘ&�VH�KA&t����@��]�d�P�O���2�i>u��Ο�e��+F�� 	H��=I'�8���[��Ny�$��Z"a�'+��%���'h�Q��Yl��bm�6Y-�ak'�';r�'�2���TW�0;ܴq�(�;�(8x��e���Ū@g��(�E���U�Ɛ|�O��ꓪ?���?Q�>X���U,a�����ȟ.Pyfd�4���#_�|e��O��O���J������hϤ{���PЂ�yr�'�r�'`��'�����r�Qz�k� �"e��B=�4��Op��U��8�q>I�ɽ�M[M>�"$�A\�B��]2X9H2h�]̓�?I.O��KŬ{���-B��A`H
T#����!�'3A�P(֢S��������$�OZ���O�扅	PDE��^��i�'!�`��$�O�˓%,��ɗ(�r�'�W>5����$I0�P�@!=_����>?a7Z���I�D&��'�"��0�S�K�A3EC;�Ƭs�/)Ԑ��ڴ��i>����ON�O�h�6�4�2�� U��e0Th�O �$�O����O1�4˓ ��Fb�M�z��' e��x�
���d��X��@�4��'����?�E+["
ӚA�%ñrX�pRn̼�?��640R�4��D´NPR��'���w����Tꝩ�h9+s
��F^��IMy��'���'2�'��Y>�"g�N n�"$T,D>pL�Λ�g'ܴ�v�d�O0�$5�I�O�$lzޱ����p8\��� ��dY��)��@�?�|���9�MS�'�8%��i��1Z|a��9Y�z�'���c�W��ԙ�|U�D��럼�gSht�P��D��в�K矤��p�I`y2��)�Q��O���O\	�a�C�d����̫>`b51��5�I����O���-�J�Y��|�Df�LB,p���r����+�d:&�����|�d,��D�	�Z!���ɒq�*��r���%8���ǟ(�	ݟ\��j�O�Mԣc��p�W ��{<�����ۖ�ҫoӚXJeϧ<���i��O���^�0YI�·�C�:9�@��,��O<�$�O�9�2�~ӎ�MC�-����lQ���	5
�ŋ�ȡ$��a�����䓦�4���D�O��$�O��D�/uq"�Ѓl�|Z�@a��*��˓d(��E��{���'�����'����;S�[���oR�䫵��>���?�J>�|Q�@�  ����И�Di��tF��������$j�% ���O��2���x思�S� ��Z��p�����?I��?���|�.O�nZO;@��ɾx~F�VG�1s��A��ĹQf�����McN>���e��	����	��s��
����$�3F�<�zG����@n�V~r띋s����S�D#�O�� $u²(�$;�±*���Dn�5 >O0�D�O����O�d�O��?�S/Y&���#�Rc���NX��(�I۟�@ܴ�ϧ�?)5�i,�'��-�CT+ !��*V"��d�|�'��O<�x÷i��)a 1�%�+N0>ıĉ+���ϕ�ZF��\��@y�O���',"�$aFfQB@�Kpp���ᘩP!��'��ɉ�M�Չ�0�?1���?�(��8�d�� �,��F�M�@�zD��Hq�O��D�OғO�/������JNk�l��G�7nք���$UF�lZ���4���'�'4��1ů6&�}J%gD5BIŠ"�'���'�OE��M��ڠ>�f�)%��
&(H��D�^��	���?���i��On��'���29��Ъ�@��z�%D˱Mx��'�(E���is�iݹ���?��P�yPfM*GU�D�`�!�Hl��Gr���'Z��'T��'���'�S�/� }@f�a�8�pÕ|m�۴'X��y���?����O�|6=�����&V�  !T2�@F�O<�� ���b��6Mv���`c$T��hU��3T)�]��e�DB傈V�2�E��Ny�O��BA2�U��K[	!r��e��1�r�'�r�'��I�M��*��?���?1�GԦaY�$����K��-+�ş���'��ꓡ?������.�����=e��S#'?�o�;|ca(3�z�'{b�����?�5ȏ�A0��4�ы5��Q8�]�?���?����?��i�O���b�5ep�D�%aA�7><)��O��o�E�&8�'4�7M?�iށ��ΩK������ C�.t	��p����˟�I0b�	m�h~2�P�I���'p�B��,A6K}��&�l28�IM>�)OP���O��D�O��$�O��2�h�A1.A�m�e��5�Ƚ<iŷi�0���'���'���yc��d��7⋙2����r	��t��?�����S�'r�9�n�!Hՠm#�I�0@  S��"Q�'2� R� Ɵl��|bW����"]PT�P�ۺE���ƀΟd�I�����py�)bӾDXR�O���*4R�h7n���=�b9O�doZp��Z���؟������;fr`��͎�L�����#l.(n�z~R�_2�p(�[�'¿+25rZ��A/�?F��r#�Z�<���?i���?���?A��d�YJ:|1DJ���(����"�'�"Lm��DA�¶<3�i��'th��eό�+F��i��ƾFr�d��|��'�OUzH[2�i����f�C&�f*CƐ%�Zd�ĈL�L2i�a��ey�O��'��
KyA�x��K�B|hP�n�0���'��ɵ�M���ʼ�?q���?A/�R��r%�nG��e�ƥQ�)[a�����O��$!�)R��ʰd]a���s`��5��[7�&��x-O�	\�?a�<���@>��c��7�e
𢊆���d�O����O��	�<��iw�E`hq���d��o���؀,�D]����س޴��'2���?   !�ՈfO3+��Ԁ%o_�?��Ww���4���FE5��s�O��I� :D�`���t�-���r�IPy��'��'2�'rP>�"� �����QΙ����f��$�Mc����?9��?M~2�9ʛ�wa��'+ئ�b�:��M;?ɼt��'�r�|��D�L!
��8O��%��<`uNƸ  �X�A4O@XC ��~b�|�Q�\�	�`BQ�ɍ��ip��\&��9xã�� �Iӟ���Wy"#`�:�rDN�O����O�l9#�o�z��s�U�C�t�0J/��?��$�O��@�Ac��#o:�H¬���0C�+?y�D_�0[f�Rc&R#��7Yl��R��?����8NN}��Qv�ڠzO���?����?Q��?1����O^p��'X�;M���cǅE��黑E�O��oZ)/wz��I񟬫ڴ���y���;Ȳ��ƹ,"-�����y��'���'��1��i��i�E����?���вN�~(�U�\� 52��Ʈ�G�'1�I��X��џ(�����	�Z��H�#"ƭ��FO���T�'�6m��{���d�O>��7�9ORh�$H�iz�\˧n�����4��T}2�'�|���k�)�������l���ö�@);�1Q�.IfG�I��\����'3�9$���'=�r��U�54^PisF����]���'���'F"����_����4[ۨm���=N))��P��x�GJ�]�h�����V��d}��'{�w2��a�$[<k�:�(1a�
"�Ȭq�͗&�V���#Å�bu���Za����uؕl)~CxQ B�9*E�V�y���I̟��	ݟ4�	�����F�$ZI�)2隩���W��?Y���?�R�i��ȣ�O
� iӼ�OxɂX��q�a¯v4%�L��'S���$���R��擟����	-�P�BDg��{�-	���?����"�O�Of��?i���?��x7�r�.J�0;�ol�D ��?!)O�Un?r���'l�]>EۦFS�mdz8#Q���'�ޠp��)?Q�R���IT�S���ёz�5����aҩ�!'��iy�(N=g](���L�$��4����HRS�	�Dh��#��Ei��aѯ�"wg�����x�'����R�x+ݴYt�kc�D>/kB����[�nD(��>�?�������$�c}2�'
&�yG!�	KEnX"A�(i�ȣ�'�'�*6}�&��t�1��[�d�~� ��I�nNP�L���+E�f�R�5O�ʓ�?����?����?)����6U?�4� l��Й2΂�5ݾ�o.1l�Iݟh��x��ݟH���s �Y. zb}٥P�X���	�?����ŞT3Njڴ�y���`Ą#Y�\a3�]�^�\̓FL@1��H�OΕ�H>�-O�i�O��bP�ϖ� ���+�<� a�On���O���<ip�i�J����'Kr�'�D1�䛣)�V�� Dn�� s�Ds}�'�"�|�#���1��h�A8�[cM���$� �$���t�J�%?	" �O|��щbz��E"�Q��`Kݼ�\���O2���O���9�'�?�a��8U0�a�R��vs%�S��?I��i�&]��P���ڴ���yׅ��b<�zi�V�T�Jѝ�y��'��'�4�x��i�i�q��?�(��O�hH�.!Fl�� ���99�'�	Ο������	�T�I�2!��¶$Y���cĈ�61@���'w 6M�Dݼ�D�OB�)�i�OL<���*]1�Eم��C�T��D�q}2�'��O1��;�'D:T0��u��x�,@�1�F�VB��k5�<� %�(�P��8�䓟�Ĕm�vds�`�&�H�)ŨB�t�f�d�OL�$�O��4�XʓE^���l��f�>b�`�H���~�������yr%g���L��O���O��D�&D�<ZQ�̘<}���2��=�|t�"Nn��O�V43���B�>���MW|���F.���
'l��h'j�I���	�����Ɵ���J��cLH�"4A%
TQ����ߦ�����c�4e���Χ�?1²i��'�0� ㏓�FT�$�� �>Y�ğ|��'��Om���s�i���?�$D�w������r� �هbN�{���$���<)��?A���?1�͠��"6��\J���"�?	���d٦�³FP�� ��͟��O}L�`χ_h�dҠ�R=6�l��OX�'T��'�ɧ�	��rS.i���K�n/�X�T�צCodX�5e��2QV��Ư�<ͧ&����?��I���dD jv� �
8�X����?A���?I�Ş��G٦��$G��V�={�\6_�<��j͕"v�����X�ݴ��'�|��?y�
ޱ��ܱ6.C�&E�$����d��L�6M ?�ѫ�n�8��R���dɏ
���x�tsN7 @pI͓����O����OT���O����|��^�g�����s���J`k�5Q=�N��R�'���'�~7=�IZ�![�x�jQ����2Q�\u{ n�O���6����	��7-f�,���ٚ3��p�F=��C���$�%a�@ ��6t��O���?��P�`� ׻E>�H���A<������?Y���?�.O>xmڧ1�V�����D�I8|�1p���k�(	�o_��*��?	#Q�0���%�!�x8�dZ�a�m�6�1p$?ٴ&Ș^�b��`�ϼ��'U�l���<�?!���V�hj�������7���?���?���?��	�O� �G�/L��K�e�[`(��M�O&Mn�n���'��72�i�a �h�-����Uig8�QR�w�0��ʟ����M�x�mR~�C�f����M!�-�' ɔ5�<S�O���e[�|�_��ȟ��I����I���� ��&�x�0+ҨM����ƩTMyg���"O�Oh���O��|���x3N� ��Zr�`8�>8��}�'�"�'rɧ�O�\�� ,��:Űq(g�0_�8�p�E�Pzb@3�X�tiCeC4V��q��ty¡_4i�4@�2�Lb� ˀ�>"2�'��'��O���MӲ�F�?��e���)7O�<\_��	`�M��?)�i��O��'X^�h��*[&��� �E[�δ{P��1�F�mZI~��������7{u�O���?�n��v�KR���1NȽ�y"�'���'���'�����0{�xpSH��@�\KQ��)?}R���O�����ԇo>�����M�I>91��9�&��s�טUs8�cr�����?a��|����M��O��(���I�҃Q8X�4S��(R��U���z�IQy��'vR�'a�c�G2���.�?�&D�үM4ob�'��ɱ�M������?���?�/�t)rk\2&���Hu�	�}��tJS����On�D�OO��<Fql�(��?*��F'�C�L�c�ƙpY8�oZ���4����'��'ݔ�#�䜞y��p%���pܑ�'2�'c���O.��9�M{p�� b�8�@ԟX�T[g��#XDL���?�i��Ot	�'��(�����Ҟ.���zadj�'پ�P�i�	<}�>������j��Ǽ.dL�c7l�%'I��<9��"hb٪��?A��?���|z�̊�/՞����O�v�$be���֊�uj��'���Ou���'�n��N��_F�yѬ���L���
�,.����Oj�O��O�$�Eq�7������* v�q����#߸Hb*e�� �[
�R�KA��Ty�O��2DH�82è�|w�$3�ɚ��b�'���'��	��MC�I>��D�O� 9�$M��SF�ThlT�� (��<���OJ��5�$X�}�E�+���Ʀ0j �I�b�"�:7m>擮)w��O8@b��7�(@��$NE���$O�OZ���ON�$�O��}J�*Ia� NF�D����cb!I�i%�F�_�"�R�'�>6�:�i�q�R�L�E�.,4�H����a��������8N�Lxl�m~Zw�꽳e�O?�� ���'o։yf���N�TD���	0�Ĥ<	��?i���?	��?��[\C�=�Cc�3DS�(��点���	Ʀa�Ce	ݟ��I��%?����N�����h�Lp�d�C3����O0���O��O1�D]3G-�(��q���|�8�0���kV�ےC�<��|y��$J�����D�1,4����4z�f�᭔!Q/b���Of��Od�4�V�雦��)�r�C�g,�Er�J�� Q���1+�\V2�|�^㟜`�O"�d�<A���.*7�}��F��6�8k��)QȪ���4���	�4�Dd��'rߴ��Z��S����WN�:��P($�X���O����O����Ol��!��/�[L�>Q�آc#֏(]�d�'�Rk�n��G4���$ݦ1&���ª�"�CC��)F�� %�H���t�i>-� �ߦ��'*�`�1��;���#��L;Cv`��i�Z=Z��r�~�OX��|J���?��%�j@"���C���a��̓_�6E"���?I.O
�n�Qy"��'��[>��C.�>$F�p��A.^`��7�o���������O�$6��?`A��_�)k�F�w ���FH 4���ƌ�ݦ�k*O��G4�~B�|�\�b��A+!�j�`��r�c��'��'`���X��Y�43Ū!k���Vbũ�A*6���)S2�?i��^��$�F}��'B���
�
�4h0@đB���� �'�ïf��H�B�$	���<y�lG"1ҭ봀ξ^X��t�H�<q)Ox�D�Op�d�O��$�O��'�Hh	�*��<X}2o_|8� ��i�&��W����C��П�������DڿLAR�J��6V��cp`��?�����S�',��a#ܴ�y"j�������R�2�����y�`�:��M�����4�6��>*� .������7� �f@����O.���O��o�� ш_K��ڟ�e�1YI����*�c�K��������џ��?i3-$U�"� K[3. �Ek���U~b�f��|G�$B%�O��h�I%Bl�ݦEAr% U��c��A�u	7;�B�'��'S�����#��E-U�Tmy��v#�
 ��� 2ܴA��.O^4l�c�Ӽ;V��,�v<s��-S���@��<���?�k�8i�4���7Td�8x��#V�P��9G��=�K�HBJm�VD%��<�'�?Q��?���?�qޅv�`�yAM_.Y�J	��B�����jXƟ������$?��	�HNP����*)AJ7�T?&����O�&�)����:�g�9�D����~�tO��cй�'9 0�������Aw�|�T�P "�pN(zv�.}��*��͟��I矌�I��Ny�n�Ѡ��O���.�:ap��4�J�9��@�S*�OB�o�o��r��I����IП����]2q��$8�GX2ʨ��2�Q�5��me~��%Gf���oܧ��d��0#�r0o��ھ�Ab)��<Y���?	���?���?���T�[(����!-0ƍ�	%���'�b�yӂ�ڱ�?i��4��u� :V��; $�����F�AO>����?�'e����4���� B%�0�4����!�JPP��S���������O����Ox�Ę�3�;�OI�M�T�K@ ��D�OʓT���Gg�ɟ��Od���C��G�x�*�`Py� 8K�'����>A��?�N>�O&�x����Y"r%��A�x�$�b�gB��l$a��i�.��|�t���x'���fiP���hF�N���)�⟨�I���	��b>y�'��7m�}�U�3�U=tp�Z�ѯ&���b�g�O^��^��?��Z�����D�2�z�����3Ј�`����I!Z4�}n�n~��]�aJ��}�uHL"T0K�pP�95�L�<	)O���O��$�O|���O�˧�� �mG�-�ݸB�KP�&�Hn<W� a��՟8��N�'#d��w@92���{i��Å�
+U�=��'�|��+��Vc��:O�E!Aʙ4�@�w���A�n�@�<O��YFL��?I��6���<�'�?i�S>\����I�B�jȫ�?A��?����D�ĦA����I����B:}V�\�S��>��D�5ʞn��
��I�\��W��B*0Hs��٢V�ы���3,�|�E��q3@��/X��|ZP(�O���Q ��h��>?�ޙ	�d��u�:�*���?����?a��h�@�ę�Ŷ��,~R�(U��Z���Ħa�Oky��m����].`$���U'Ç_���eſxچ��ȟ|�'?�1��i��	�^ Pԛ��O!����֐BtL(��`���4�iV�IK�	wy��'Zb�'�B�'5���|�~@�M2b:���r�����9�M������?���?�N~ΓL�P:1��8,�"��-[SG
(�WT�`�I���&�b>�H�f]�m�!�.O�(q�:NH|�`�ض�+?t�5�v�$���䓴��(v*����蒜R}�š��_0<v�$�O����On�4���s]�v��'�ƘH�xP�w�ӀF3��c��y�f����O����Ot��SYl�D���o�(�4k�)��cCdӎ�0df���>���7�qX�h_�4L&�� $�Iǟ���� ��֟�Is��H��d�a.T`��C�n-�XU����?)��(ƛf$�+j��	��M�J>���R��*�Ⲃ��L�N�Ҥ�4���?���|r�޴�MK�O��YE�? ��t#MH�H$`e�
3wh�`J]��?�$�-�d�<a���?���?�5��B�(��u��,~n.��*�$�?�����$U�!�C�����	��h�O���g��=|񰄉�5榁C�O���'�2�'�ɧ�i�/W��XǗ:]F� #��5C�0�pE �m%P6�My�O|����b���R$��PNxd��Ō�'R����?���?��Ş��ğ䦵�E-^*& "̃a���	�L�<N�I�����Z�4��'u�듀?� ���Y>�YP��B�<ٛ�ݭ�?���V�z��ش��D��x�����e	�@CjDIvY�� 02��T7�yT���	�L�	ޟ �����O1��������<�l\4}
��u� �f�O���Ov������?���JB�צ4H��M�v������$�b>� �MD�a�y�Qh��
b���˛�@P�̓m�q����O�iAH>�(O�i�O��U�ܳ����%cO�&�3F �O\���O���<�4�i:D����'���'����,���#��n��pP���S}�'l��|��:"i� D�:-G&X#1�M.��d��bZ���Bs��c>H1�O����~��5�ťZ�`Gl� @��,s����O��$�OH�:ڧ�?Ɂ$ �U�D#"�^ �t��ƴ�?���i�� ���'��/h�z��]�mg��pREu9h����2qB�ٟ`�I˟�Xw'���',hy���L�?��R!!��1 �% >H���CL�'?�i>=�I��I��,�I�v�x|8�(J.5�=�a$U8��'��6�Qeq*ʓ�?�M~r�bRI�b�D�T����k��We�%��V�\�Iş�&�b>ɢ�'�;{�� ;��C$G u飦�O�`m%��KE0|*�'��'則-]�x��C�e��+��Dd0��I�h���l�i>��'�6mU:��ɒ
Ǽ=�t��98S��f�1���$���?��\��	���I�Dd��S��s�f$�3안+�=8��'#6�&�Q�O�KF�9e��{��3A)
��1�yB�']��'���'V����')�&�1'G�'"nޱd�Ԗs}���O������X��o>I����M�N>��F�RS��
�
ޜ^^y9�㚘�䓎?9��|� f�"�M�O�a!P��S�vxH$$�bV�qW�L)�����AB`�O���|���?i������Z�7�����8��TJ���?)O��nZyhjE�	ȟ\��]�ă�=@�(!*`�
Z��<�+���D�W}�'�B�|ʟ>)z�B@��4=)�DÒT5j=if���*+x�I'�������|b���OJd�H>Yh ��Q �O	Z�ΥxM��?i���?1��?�|�,O��nZ�>�j���� :o��t ���;J!x4ò�V^yB-a���@ �O��DW?�F����{�^�Q��S|t�$�O�p8�v���Ӻ[�%���Q�<�#��(�1 �P���pP�<�*OL�D�Od���O��D�OZ�'�5 1��]h�1�t`�=;�`���i�dс�'���'��y"�~��7)�������U��q�h��n�
�D�O�O1�f̑lg���/|�~�ٲm�w����jOz�R�ɜ-��y�'��@$����4�'�a  F��`�Ʃ��.Y��(0�'|R�'BW�qܴR.Zq#��?y��I�� ӂ�R�k��Ց�J*� �ی�m�>����?�I>a�a[�k�\S`�L�$!k�k�C~���.��P�`W�O����nMb�A\���
� X]h3O��l���'���'�"����ؙs�*����#��&`����Sߟ���4~ML����?���i%�O����x4��ꪉ`wZ�Um��O����OD���w��n"�����?i��Օq�p�7-*t�
���
�V�Ijy�OJ��'���'G�E>q���Y6AR"+FUР���X�I
�M#�/ˆ�?����?���4��v�Y �$req��$Z���?���S�'Q#-X�G�U���B!l¨Q�A"�a,�M[0^��ʕ��D5��<�C�ݢ)�hI�6(G�w@D���ڑ�?I���?��G�R�������֦rҌ��	�!Rĸ0� T���#)��+$T���M�I>������џ��'ʰ�����/�p[F��Z��{g �>N��8O�z�i���'_�˓�B��Uj2��e	����ҨV?��	��?����?����?���O�DY����*���1��q��%�'9�'}@6M�q��˓����|�R
<���!�߱cА�1f�ј'P2^��RbDѦQ�'� }�3� ~H��z�JYFx� �8(��	�7��')������I̟�ɀL��bJ�c���p���(�ԟ0��Ay"irӔK� �O ���OZ˧7���pF�ӂa���F*Yw��'f��?y���S����W^f��@K� Uf4��0JI����Wt�9 �iy\��|�G���%�du-�.�l̫Ҏ@�q�6D��ȟ������I�b>��'#7M�=���u�![�Jq��oªz��i� �<iS�i�ORq�'r�E*Dmh�猼_����ٮG��'�ʤ�F�i����CKڥ1s�O��'n�n1рh�l���Qk�>sn8=Γ���OL���O���O����|BJ�E��-SR�����A�*�)�����%eHr�'�B���'lB7=����R�T��1�"cP9�'�O��d!��U
f 6-u�� (��^��@|��Aӣt$���t7O�U���?G�:���<ͧ�?q��֙:����E6��x2���?����?����˦�	��Eȟ���ş�����0
"	ބ� 42f�J��$���柰��E�I�=-�H�E�@dʶ�T�B=����4mCd��Jz��|�t�O���DrH<�ˆ�$���NT
H�P����?���?i���h�����
J&л�M����2�䁂z�
��������Rٟ4��2�MK��wh�Xq�i֊q�(2u�ߵ!�Ԭ	�';�S�<������'���R��?Mq�L�1MK�@'L�}�n����H	$��'��I�T�����	��l�	����t���	a�WJ�'06�}�t��?QI~r��$MptK�m��Jki��bn��GT���I۟'�b>��1,X�Q�zO��{��� K�&��m��dx��4Y�'��'F�I9��8;w�*]bn�q �!63�������ӟ\�i>��'uD6퉍?�����MY^��t�ȴt�|z��������Φ	�?%S����ן�9K�¼��`F�=+���'�W�L%h@����'	^2%��f�M~:�;,��	� B�õ)�!VHΓ�?A��?q��?���O���I�4[�(k��B�JJfyR��'�r�'wp6MZ:i+���O>9m�\��G��͢�a*4Җ�j�'�t���$�8�����|��lF~bÑ�v�X�c�n��
լ��R��$5��UR�Ez?�L>�-O:�D�O����O�]٣b
�'�:\��̌m0��p"�O���<��iAN\[qV���	@���J��(���hz �(F�����Mu}B�'�r�|ʟK��#�F�p�@��Ji�5˃��Xx:bC;��xc�O�	��?�Ƭ>���]E�de՛-^�$l܏D|���I䟸��ğ��)�By��o��qz�II�gs��/�h���J p�����O���_ئ9�?��V���	�^aM�D.�(pBt!:pdԗE����Iğ��
�ɦ��'8��a+�Q�(O�����<)�W,��8�{P:Op��?���?����?����5F�|�A��X�Th��6,-mZ90�
��'U����'��7=��-���"=ހ�pi�H%"�K0`�O��,��)��{B6z��ؗK7H|s��>&����k��q#��W;�0��<�O�$���b�x�T��5f���	Ó
7�F/��I��0+@A�_�1���N�	�P��%�s�3�	ݟ0��M�Ʌ� ��5j\>XxH��f�'%��}������ON^��J~r�l�OJ���i����"h؃Y)f81�/V�D��P�ޑ�7
��S�����U
��b�b��vB,P�	��Mk��w/�E�t��`l�{k���ĸ�'GR�'�R�ӆ��֔��Z�� �<5���.c)
l�dj��w��r�8l���O����O��������2����68��������4[�x��+O �"���D��̒֫�+ (|sd�M ���O����O�O1�@��c�G���I H��%��.S�7�RKyR��?)_t���䓭�D\��A`�� ꀉ#b��a|��y�lDY���O�l!R�%g�0$����^r�Q�6O�yn�F����	ޟ���ҟx�1��qc4�IS��	z��j��?lb��mZr~R���'
p��S#�O'�(0� ���+�#Y^p�a����yb�'�`Qs��^�$L��־NH��]� ��;�Ms�O�_���`�ΓO*�����&+p��"p͘� ���6�"���O�4��a�~��
�4y��(�N!��JEN_4g���2�Ib��9�eR1K���EO^B�xU���}GedhS�Hؼ�P��B�I�@2�W���U*R��&�n1 ���_�ո�W6�^!SPJ��ejʄ0�0э�D0]����W�S�����$�k6	���J
�.30�Y�:^�0ya䑵V����m�5	?�5ɢ��zf��D��N$�xDJ�*j$ ����)�|��Ì�}��\C�N&'��,�s��1&�x9�L�0^|�����?'�@��"�	�t����F�G�6��U6�d(�!o� NنȷK33ƪ�`gB��K���'�r�'���Eތ��"l�9hN^���N�>BLO����O���b�1�	C�F�\" �fQ����?3*T�Zu+����'}�xRq/u���D�Od���~�֧5���5g%hE	LT}��U{Tȅ��M���?��O���'Vq�^ZW�A�lL�kp�}�$��!�ik:�k��iӄ���Oj�d럮1�'�剶RU���b����1��;WX���ݴm+��Ӌr���O6x�G � [�jBjL�rl�x��覹�I쟈���N��X�Oh˓�?��'����˹1FUy���:x�@ћ�}��Q�@��'eR�'��'7%:���224����c9P7��O�؁A��_}�S����w�i���Dm�F͢�ۃO���	�/�>y��Ѓ�?1+O��$�O���<!3��4V�]	�ԁ&^�8a䫔�.M#Z� �'�r�|��'�b/M	}'Ȋ�
��J�ӥϕ�!��(1G�|��'���'��"�0�O�j���gK/x���c�J����z�4����O��Ox���O2�+�[�8�e��BuFL� A�)|��Yef�>)���?�����ئ5��Ocr��^���3�Ȯm���"��=i�7M�O �O��d�OzMrG-�p���T痾&�np�'h�0>�
6��O��Ľ<�K8*������	�?q�� z��!@Iv�B�bҗO �8"��x��'�LE�{=��|rԟD�v�T�PH�dp�/�?o�r���i��!	�xߴ�?���?���g��i�-� l�)�pA劚�	�QӢwӆ�d�O��#��#�Ik�'ug���S���aI�0c2D�D��nD�
|�ٴ�?����?!��2��|yRƱtzB@��Y#q��ј"��	8x�6�X�� ���B��!�ؑ����ZC��D���e��iH��'����L�f����Or�	�G_�[2K7Z/���uKևOFFb�|�w�YQ��ǟ���ߟx1'�z���D.�x�8G�*�M+�X!�a��R���'12�|Zc��|@���"�ΡQE�7vºӪO�����5���O����O�˓W��pX�K�Q\���#����#�-�a��IoyR�'��'B�'� ��>�|���I?��Z�eE�13�'>�',"Z�|�PeA-���O]7"l �p���Z�P�2����$�O��$4��<�'�?���غ1�šU�Ο�����`_~���P����d�'��(���7��C�m�ͻUęE��}'���b�`lZ�4'�Ĕ����'(�'d���Ъ� 
PMz	�/.�zyoϟ�Ijy�ɒK��"����kX�2E���B%�#+��qC��Z7}ʉ'W�I��$��\�s���?�"EhaG�d�g ùs��6-�<�߾Q��̪~���Z����3 �)A��R�C3\t�-J�Ji���?��@J�O���M#'٨ΰР���,�+ae��[��Y��M[���?	���C�x�O�F!�P�]Ƅ 3@-��ؽ�`�q�,��O���1��?�	��y��
.D���{G�(��iY�MK��?)�u=�,�U�x�O���O�	:�
T�x(�� �*ID�8�i�|��~�'��O@؀gm�j����=~0�i���K�w��	����!�I<kO����*15.%�B@�'i��J<��j_q̓�?�)O��DF5�����HU�b����t%hEɓ�<Y���?��b�'��$��
��E*�HƵ�A�b��7�����'\Z���I!/}��'vS,���79�H\Y�Ξ!�Ql�ğ��IY��?!+O,����i� �av��"d��y��(
�88�O�d�O0�Ĩ<Y��0[P�Or�UK��M'+a�\3���Y�u� �{���D,�d�<ͧ�?�K?}����Ҁb��[�xzf�l� ���O�˓S-��7���'��\cf�]��Iqc�d�T'R#'�hK<�.O�d�O����'�_��R�ɇG `�U���ɫg���	ן���̟���oyZw�����)[<z����Y�4h@ڴ�?)-O�0�S�)��7$(�$�֢%vıp�٦E;����$\6��O^�D�O�)^K�i>%AD��OE@hx*B.7u�̹
�M���?����S��'y���;o���⨌4���h䕜o37��O�D�O@�c�m�c�i>��	v?���^_�t��G�_N H�όƦ}��n�������	G?y�$�2c~�Yn#4T���΂Ħ���	c�i�'$�'��'�,x��(�WHt\��дF���hZ\�'q����O�$�OR�d�<aiE�G�"`��e�?$h�-��C�8N��;S�x��'1B�|�]��ݞ5g ��u/�%�|��J�U��7-�O�˓�?����?�.O�ax�J��|b��Y2{N!���Zj� "(Tv}R�'|b�|BZ���㟈K&O_�[��(��	^L\H������d�O����OF�]�6Y�Q?��	�[K2�yDJ�*��Tج�{���M��jyr�'�"�'j��	�'^��'v=�1�2F,�@��J��1sg&�����O�˓Wߒ���Q?��	����0,��*��p��DJ�,�i�Ҡ�OL��O�$�?r��|Γ��4̘#S)X �`(8������.�M{,O�X���\즩����I�?y��O��#�L��@�����R��զ��	П$������zy���׺p��U�『�CL��`��؋b���S5j�6��O���Op��C}�\�d�ŏZ�w�h� �2ox2���.Đ�M#@L��<I�����,��ޟ ygi�\�2ɱ��lOR�B�G0�M���?I�*v��ȱ^�ȕ'5��Or�*$Eʸ<u����Я|��i��W����Ov��?���?!$�D�V����&M�8S�* y�+V�/����'J���%�>�*OV���<����i��@�s֧ [���z�&�h}��t?�/O�D�OL�����#%SW"Phy�_0�S%��<S�x�'�џȕ'��'G��߭[��$�UgEbw�P9�m\1H�"qП'wb�'���'�bW��(6,���Ċ��X�BlJ�Q�>�v��M�.O���<���?��g�܁�h�4�EÌ �D�� X�#P�W�����T�IpyB�G(8��?	EC6�S$��� c��H�s��v�'��I˟���ٟ4js���	��8���#J{�1���M�N�
�ZcL޷�M����?a,O:u+Q��e�t�'�R�O�(I�Bmߤ�8�`�!֭,����Ʃ>���?��q��P�'��[2����K~R���ߩa�a�5�Ϧq�'7{�cs�r���OP�����a֧u�O�U�$Ft�� j��7��O��d>!�D=�D"�S++a@��c�F���̀"jL7�!x]��m՟H��ڟ��S���D�<�� ĨR�� !S���%�^S� �iM����'�[�$����pR�[��8�f`⒇�4$|�`�a�ii"�']�M˙,�j���$�O����s�b��,F�f�,	CPbPn%�6m�O��%�<�S��'b�'�bKM7!��h�aP�n1�1�kӠ�D�*,��'���ޟȗ'�Zc�!;�-إ{^uS��z��� �OX�{�<O2��O����O2��<���-8��)�r�-�@��db���ġ<������O��$�OؘIS��v�(�r�ԏ4�(��Ӫ�u���OL�d�O�d�O�AG�*�6��A��E���0��ۃ1Nν�Զi`�����'a��'��#����	ϩE�H�J#F�[9�(��;��ԟt��ßܔ'�E��E�~��E��H�m
��%��L� -�8��i�BQ� �	՟$�I�V��IA��|b�$�Q�@j'f� ̐uJ�F�'R]�8�v!���'�?q�'tb<�ql҉+ȡ����:kQ�I�xR�'�B׀59�|�П R+�4L�bÀ�1Z�$k��iE�I�J�b��ڴZO�S��������W\z�y�ݽ<.�Bu/��gg���'�B'M�O��>�#,
H�^@Rs�%W�A`�k����˦��	ß�I�?={�}B,��F  M���V����͖�O��6�T
���3�$ ��ៀ�dI��@�L�KfiI�`3 %Ƒ�M{��?	��v����xB�'y��O�y:t�S8�9s��\Y"$��i��'�ެ�	,�i�O��D�Oݰ)ԛ>�f8�%<_��A1�Ԧ��ɼiK����}"�'�ɧ5&�_F��0y����֣�3��D��]�<A���?�����y1z�#ۑ0�LQE��r?~I��d(��c���It�ϟ��	�k��(q-ӊ+���'^�,�|�X�g���'���'�R�!F�0��d&W#����K��w��I���'��$�O�d�<a��?Q�>Pt��E
䪰bņ�*#@��\���UU���ӟ�	lyB�*^��(l�����Ҷ�7NUس�,�ۦ�	P�	�� �ɌC���@��Ap-~m�D�e�i�nG�l����4�?Y����Ḏ2�$>����?�k�"�+P�\((a���["h�A��	�ē�?���-=8Γ�䓒�4B������`�b�U�ֹ�M�+O
�K������������'�x7��I=P��ǿQ;x� ۴�?)��eKT̓����O\�a�1�F& @���1#H5��xH�43uܠ1�iG��'��ÒO>���c�V�aeK�����ʓ{�Hnڨym�e��q�J�'�?q`��9���c�$:��T'-$t�F�'���'�hP��.�������m[�5���u��T`"���L��Hl�@�	�f�<��H|���?���;��0�H;XI3�O��-��}9��i�CO�i��O �d�O^�Okl�>P��]xb��0�Pd�EI��;���.b0���myb�'���'��	6{K��A/�X
S)�A{�y��>�ē�?����?�s�� t�%O:�x�^n}��؜M����fy��'I"�'���'[v�mO*RD�Q�Ӫ��,2ҋ���q�O\�D�O��O^�d�O�4�T��O�Ĩ2��s��%r��H;��1 F�`}��'x��'c�ɚtC2�rI|j #�B3��J$� K3�Lp>T�V�'��'}B�'s0��S��V��pa� �46�Z8JV�V'����'��V�$CV/Q�ħ�?I��^����d�1�93�ϩb��t ��x"�'�R놁�yr�|֟>	�%�T�s�����ǂ�t�;a�i��<Q��ߴ��͟H�S��$T�3邵+�N�R�$��hK��f�'���4e_��|2��QYƄi`ʫkD�*Eƀ@l�v&�0�*6��OH�$�O��i�E�i>Y��j�q	�(�DÙ0�>�h�bT&����O��b>i�ɱq}FP@7�,(8*l�I�yg�(��4�?���?	��?�J~��~Z/��9���Ԭ!@�K*̄4ʜ��d�f�Sߟ��	��0zW%��.���Z�Ix�Aq��M���h)L]��x��'�"�|Zc:0X���ҎK��L�#/[��h���O�m�d�O����O��Cr���G�ϰ^��u�è��_
���$S
�'��'�'��']ʰ*��"���!e=0[sJ����'sb]�dA��̢}Z���@x�Q�#��V8�A�5�JL�<�5%��b
�����~�� �OH�J�؀焬-��83��Քgi����dv�zB�Hl�A��$;s+�%ؔ#X�c��taF��'RZ���Z�{UZ��u�G
X����a"!OSx�$W�W�@� ���W���H�V��a�v��?20��e�݈jtX��0hY!eX�E26D̀g�4�i���3�jͱ�%"h��L�	z�B��3'�>a�J��E״K�rA��🨓)�'74��G�^M�B��0�ޠV��I�|.��p�%�O�X�����6h��Oı��훳$��g� .� 0��͛�ڦ����!Nl֝�G�©ŉ��|,���ф_�N���'�^4���?a��	�ODh�@��.y�R�p��ѣN��"O4�g�;U�T�aF��Q׺�2��'h&"=YD/Z�2�*�@��&���4oռDu���',b�'&*�7���|o��'-b�y�\+m�����͝ %0�G-�y�1O����'�́I2,S�$�\���	B��8Q�{�	:��<� (ze�Z�_KJj2�t�*�$�3�ɒv�"���|�D�O��L�T�n�t8��ڬ�y��ە(�2�#Κ˨�͟���CJ���Xd3�c]�r`j�0Q7�HI��X<`7��� ��O\��O��D]ٺ���?�O�^7a��a�$�^F�j����D|:ə���/%��',�h��ý!Al]	Dۡs^�]b�'�82�\cq��R l�K��'�\+�,���q��.u�~��Ƥ¼�?1���hOx#<V�ϔy0F�zg�1%���PK*D��$5{\�`1��S@&p��#��)��ļ<����Rٛv�'��)�+z��,�צ��~G����V��'������'6r<�*���'M�'�,����,ZP���w���rH�I�	�,ܰ��?!��;l���Z�5`;
]��FF8�"���O��O\)�0�	��-��+� �"O�����R�k"��'���FO
=oڑ<���(�OG>y�$��ǀ�nc�@�����Mc��?-�LqRs��Ofy���F42��ؖGV�8���V+�O���Z��D0�|�'�~qxaըL����$�v�[L�TPGa%�S�',ZbA	PG̹h���P �;!J4�O��)��'G1O�1�� .r�Xx��o��cu.��"O���dZ5YK<e���}�鳄�',T"=ѳ@S�U����!l�S%d�ӅA�.<���'��'���'hW�>�"�'��y�AY�j�0�
�;+���D�O21Ov4��'Ɏ�S���F$X�f�ͣO�x�ۈ{��<��<�&b�dh�tI���81QX,f���'VP,1�S�g�+��l��F�f��	j����7�$B�I�:���) @�Q����K�1��X]��"|B'N��*��Y(���2pZNt��%�<P00zU��?����?���+5���O���i>�9��)F�X�E]5v�~(
ud�vB�I2*�A�nO�U���,!/N��<�ˆ�X�^@Y)���?�B���gC�2����1�OZ��
�0��!�1&ˈ|B\�"O�X ���;�� b��Sh�YH��di�J��V�i�"�'�r$�!APU9�x�D�,"6�� t�'�^�.K��'��c���|A�*[��86�G,P��3�@�p<�d�m��}���1�iW!����� �*�9��I�_q��.��6e+�h��/D�QZ�d�.�!�ĉ f�)[��σ%P�����Q!�$V�-!C;l�.�épg\��$�(D�8�ks��2E�X<a\T��s"D�����	��2���!�1{p
 D��j1�%kl�yX��}�U�un2D��+�D	\�<��v�
�&��	��,D��!f��D݀�9��I�:�(�r�l D��は�8���J�B�U<�
�)D���d	'v�65����d�C� (D��+ �X���H9`%�6*�؅�%D��)1,�u8����@7H"`�S�!D�ؑ��+j{v���(��0�⽀��;D�pK7@ߗ1?�h(�H�{vD��I;D��w�J�W^@���I�7&2)
@�:D�Ġ�	�<�8��.B�c<�\���4D�,���!n?♈3n���@�P��3D��چk��w�:1���܏$�4T���1D�LP�'Ģ}�8�*�-�R��j��+D��Ѕ� q&������&��9�#>D�dqO�a~RL�E(I;OH$,��k<D����O'Hv���f�ڋf4� %�:D���d�Gc���-T�5�R1�6D�Ѓ��ų��d 0!T/-eT��%�'D��k7�׫XǶ4i� 7����I+D��*�j�X��Pr/�z�ڈ���>D��P�}e�]��)�^�f�1�=D�,�b��9(��X�J��xi��!:D��d�vZl� �(W$�ʹ�c�6D�� VmYa��VVh�ak�B�l�)�"O@��&�\R
NI1�㊇HА��'��E��bL�T�XK�Y�Y32�)�'��D� ��(7	B�V#���
�'��٫#?;j���pb��E�	�'��� w�8�0n��-��e*�'�(�a����\�"���ې��'��M��A;2W�8�C�Z��ɓ�'�����ʀv��|���q�r���'���(6@��*� �"�a�P$
�'e��\�6.��"�;'s�t�' ��	�FB�{O�u*�Hq��pP�'����)�$l��������,h�'�j���'�8?�Xy�gW��4y�'�p(��ޞCSf�v��,��'�!
뒝s�ݒp
���"�'��zM��3�0ys�ix�B�y2,�3=Jvu��C�t�lL���ƭ�y"�]�4jH0t���rv~�K�#,�y"��:J0-�R�U�@�Z�vK���ybb��m[uJ�=f ���֭��y��"FGz��և5�(Df��7�y�fE�j0z-b*�4CT��Մ��y� �[�4\p�T83�j�rEg�y���*[���j["&���Ǧ���yb� 8dY�P��}�f��ɟ��yb�Ӗ6�yz���f���[��Z�y�R	v�Lq���@^%��qr���y�耀YY�H1�k�$F�݁�ǂ�y�O�Hb>�*��H9Tø�
 ʗ�yb��5u��V�J Hlb��V��y�	C�Q�l�;�Ɯ�V���s��>�y�B�"Tk^�8��$��q@Ci	-�y2J�*��h�0��1Ǵ��R���ybk�(7����2lۢ�Y��yJ��	�>�9Q'!yπ��2��.�y@�/#HHX�B��pO�4���?�y"�P��� �;*��C�͞��y��HZ\�Pp'��16ȃ��-�p=	ec<扻=���U�NBq��Qu�R�<�HC�I���kլ76�.}c�m��g�L➰�2A5�S�S1W��m@Ӣ�v�L�
�/O	4�HB�	�U4�1�@@((&(àZp!�?AD�B����	bf�*�|���JP�!�dD�U���!�R�7c�ػ�Ğ�K�F�Y��?| �z7�'��x����~r�ئ
7�l��h�,@�H�@�d���{0i 8�$h"V�۟�IqڤGh�E˒�2gD(�3&'�T��L�=��>Y6N�W���d-F1dɂ�Q䡓h�I$I��S੃�%c�=�L~d������	<B�<�q��Xp޹	WkH���C��'v�}rFĺb���a��U��9�v�B�D�)�Y86 ��Q�k$�x�bL���N���i޹Pt��8P�U�&��,��p{a� $��"b'U?}��9BRJ����qX�(�'����T?	z�I�1��*d/E=W�����p�����0�q��W`���^�C�&�0�Z�=��  ��%�~@)t�
���MQ1������Q׺|��j�7V��p��l�=LMt�L<)V�YO{ܱȢL����YS�Y}�A����
�:E
5I�a�Vٔ扨A�:�ѠX�dF�@���c�b�i̦k�KHC� ��Ԅ�A�
��0n�}ay
ʨ5:�U���!�������� ��X�I�{�*���'��xҘU�T���m?�O(�i�D�>f7�-kr�ݪ%�����*�O�i�`"@��	z�jK�R�IF��$f���䐰7�6�(Rȟ�AH?mW"�pI(p{��T�b����P��%�(��k �o.p�Y�'˔�TF�A(���o�{p&բd��w{���7���<R��
�	������j�/7�ƵЗCR�<A�`�C��9N/v�p�cL+=��'"�"s!��	��2��G���K<�7mL{�x!�R�.ZT*Q�\�F����'��E!C
�2>��ѫC%Q�F�"�*WF�)���Q=P=:Ue�rQaz�gX�Pj�"@�sʾphF-����{���6�5;��{�(���^0Y�Ң�<�'��� ����M�	4�7Sl�	SpOި�0���9Ju�"AJ�>ؤ��Α�-�Z�+��\�&Ih+O�Iuݕ�$M��V��H1���u�����'�t�`p��,�-j4���g��c��0	w�
-$d�{� �l����d�;9��5X��) ER�8C^����ɺO� *���92���K6ʍ,0���=�r&;O��뷯J�s� �# Rܓ�M�'�h���`(��>{��8�Y��!���>�.��f ��h�Y`�J�ZQ̓*��Ȉ�I�%&.43d��~H.�E|r�&ţV��H�
�h0��B���cf�A*�l삐���FJy"Ó�>�貦��!j�`F;l2}���n��i�q��f��K��`��!�YM�y�)	z8�@
E�ş4��5ﬨ�`��F�J��qM�;D#hx0`�'WD�A0��'CƬ��d�_����{�`Y-*�)���Q�qO�3sb�O�Z��EKziS� _w������'�x�i���%F�`�  ��2cb|��}��ȥX��D�1��&7d����ē�A�1e�"H)��V�ָnSv��P�'��-���>-�n��m�Om�@���.�("��쒔3�E�v��D�2��2�&Y�Dk�y���ص&�PTx�+V�+�HpĞ�h��|)� T�W:b��dC�H^]�Dfч(��a7k_1F6�����E�dƞ"��ԟ.d�G�f<�V�_�~X��Y|1$�t�c8�Ē�g��K���,�%<�Jɬ(jĨ�|"]��X�hT�'�"\��ñ���Ě������5�A�&H쉓�@+8�laa *ړh�r�s�2;b�$R��~Γ������(�Kȓ�=��n�6�� ��*�8�xP��L6�>�3ғ+9�8�C��� ��b��\(�RD�'��(��.���6曞�?Q�*µ\���4��);2�C@ȅk�ĠEa��q��+�Yx���֫Aj���@uB�=755�r�7��7�4�v��:)=����.�T��'nW��Q*� ���'��p��Xd�����hZ����FT���5{��[-8�Э���<O�DD*�bH�7�Ԁ�ͪ�ȟ��M���R�AB�<Ȁl!��X�y20̈́yIr��w��u[�
0s0��dw�1{�O�%���,�Q���bȔv���DK8ή�� 1D�9U�)��������a��o*D���r��%op�3���|$���*D���Bԏo6�+�$U�q�M:D��&b��c� 0���-b��Bb�8D��V�@
F�"��F@�[|]Ʌm8D�d( ��+ Z���&
��D*d�:D���)К��f��q|�0:D�4�R*�,��5KD�7����5D���D� #�y�#tVvdA� D�h2��˻_�.H3fE\S�F8��1D��0�،{�N�b��5Mu��ys�1D��Ԩ��2g4��$!n�K�/D�{�%A����g��<��(�	?D�`ôD^-ihTًCh0���1��!�	V��8Ǔ�VA�EΏ�a��8FA�2'�H��z���F�˽j�ZeC2�\��#o�B�	zw��U���[��`�J�M�\��V�j�~uJ�yRfO>p����Ŗr�b9�A�P�y��VF t#���?�2ь���	/w�aC�}���b�R���SѠ׍����5KZ��ybG�*5���&�o"����$14~d�&�$i��Hf`q��'_V� O�S�ИfH�@$���
�'�R�)�BS!d 6u� BL�hu¸�Ӕ%$5�b2�O�9�p��;a�$@�
��ZRM !�'�uӀ!�(D�"�'Þ�*��=ZT "u�&��Y�',@X�h��F|ܐ1�ラ$8�LqH��a��WA`�J<����έ�v�*֨ʮei~�WL�j�<��0w�iB��.y�Xma�J��O����$̸��Ҿ��� 5{�v�*� 'Q=���mWX�����K�l����T�cd�`�)�U����4�':vh��@�=��)H�H�/Y"l�y�x�' � !��_�(Y@s�8J%��13��z�(��z�x;*�(e�Aq�ceYA3!2}�c0F�0���O�����gUQ�����r���A-.D����7}` ��R�_�	j���N��'��RT�s�g�	&8p��P��c�"�#��B+�bC�	0� �E!�	]3v�-#�@ִAor����^&��3��'�
�y0&<=�:�KdK��8�DYǓx�� ��.�/z��m��ѻ�ΓJ�ҬyG�GT����r��p���S�~���� N�hP�0E�D��'ٰ�!�	H�S��W�Ab�h/YvQ�R�	���\�O����O�0=C	F2Қ�"s�G�h@f�Ltܓ'D$ ��&;��?�ᄣB8?�"u����>y�Xې���~��Bቝa� �##"�M�x(��	�|��)u
A:6*Q��)�I�>�����s>���M�-�xQ�v2,OlIW�@̓eRz�I�F��R���;P�F!r�p�'�T�rd�<�)ҧn!JD�tAZl�^�ه7z�؅�W.�ݣ��\�jmc�B�}v0��"����k����H�Ԅ�"Їȓf���K'!&��\􌕀m�:��ȓ	gvՓ�脵9f���$ͼ��8�ȓ,+�E��N:$K�Y0'YaɌ���h>���s+C V��F�Dz�=�ȓH�(��](W�)��C�yWTT��j�@����ɤf4�@`fb�F��!�ȓ^W�P����N�{ �UL�@��&�F,���&G�ZW������ȓG����S�O�B�j6햞n�|���]�乂�Z��<QR%�D2{朄ȓ(�t(b��2:I�A��G'99.��T�f��4!�����N�إ��^�6UQ�c�8Q^Tx����w-��ȓ7��T�$[4�$�:�胝0"��ȓ<[$٪�N��{R0�ӎ	��J-�ȓ4x,�&��H�v
�D� ��5�ȓW���E��� ��0K��z���>��P���ɂwy(83��4`�|��Z�[S��jƌD�A�Y
�2�ȓ\�����N$NL�% �&�eL�(�ȓnTc�o��T��q��,D�3��x��$R���+J�pc����%�0�M��JZ<=�cʮK_bH�󦖍-:�]��g������,]}y�I�4�dP�ȓuj����̦9��0i0g�0;���nTU�A�ɒ:�2�F����ԅ�=V0��+�}|���$ƋK�
��ȓH;���� �b��|�(��2(B؅ȓu�x�gA*�.��V�؄3��@��:;8[cf�K���e�U6�(�ʓ>�:<)N�;(��c�#�;�B�	�>��
Q��RE��(��Dn�C�	E��+�g�8�5�E.xC�ɑ?G`����-�����Lܹ+bC�	,��=[G��|E��9�EY�Js(C�ɹV�Ԝ�w�՚� �0�Q��B�	m�8}�d�'��Ҕ�6;��B�I�q��QÇ��W��D���ކ+��B�ɸ~L��H@L��}�	r��^+� B�I��$���
,A�`���׈Bb<C�1wP8��,�?0�`2�Ԯz C�S!Z�PC��5h
(�B-�d�B�I^x��P
,�8��ץ�.=��B�I�S�4��(єc�ƌ���N�m��B�>ؾ@j�}�\5��!��bB�Ii��D��> �V�"��c"*B�ə;d��a�30�V�IV�6�*C��<m���1�@M�R!���
D� C��!#��Q�D�.ɻ�D }_�B��1-Z��@ƅ\�<���`03m�B�	�nq���BE'e�A���jϚB�)� ��gO�%^Ͳ�d�V~�QB�"O�����7}RN�X�&d��"O2�Y�E<+T��ƍ�'K�x��"O���.�M�|�JvŽu�X��"O��!�b�Ɣ�9 �'-�J��"O6�y,�8of�i�*�#MD�x2"O�	
�H"8t���է̵(���"Oxt�T��!h�d���eҩ�pl8`"O|�*ĘP�%�&�هX���"O4%qC��Cr����h]�w��"O^�SױT�
���=/`ayW%K�y��A�	��l� ��3�|�w@C0�y2N
�?_�(�!F�ܕ���T��C�	�LOVE���96��;fO��z|�C�	�QT�%�2�łȈ�K�	!N� C䉘7��8��OM��<�Õ�m��B��:/�))�G��0������3p��B�	,H�A��)M@���7N��EO�C�+�Љ�mO������2iT�C�I�'xډp́ S^<`�3'N�RC�	�:�T��hK>)D.���Y%vB䉨ap��%.Z�p�E`բɡaSC䉄;�]���D������4B��0�qs+��0�<�+�� |�TC�ɴn�be�H@sk�]�%�N�C�ɫ���b ��-g(	ԅ،2��B�It­�E�N�`���e�Q;*^�B�'%� ��U��]@��9�+\5�nB�0l��p����1V�!��%,B��>:\"P�����4�'��G'�C�Ic1~�a�P m���+!�K��C�/a?��:%�9)48�3.گ�4B䉆0C��0�
��n�Vl�p��o�$B䉀?�2@j��ʜK8�K��L��C�ɯj�,$z���h2f��f�T�a3�C�	�Ne��Ą.
�8�'678����#�	9��m�*��3�h2��	��C�I��Ę�Da"��A��^�fKLC�	4��� ��?jz�(Q��\�,C�I�:��1���@|\��a��?�C�	}\|!ٖ��f�8��$`ǻ:�*B�I*;YΈI�<$���+i�.C䉎ԞU����Sܥ�"
�v{C䉔:����K�4-n�0`D��R|DB�I�2�@]���ƽN��D�r�P�C�	j)Rwf�YG�����F4�B�ɦd����A��Y���zЭC�4�C��6j炍3�9fF�Un�S��C�	9��PR���_;d���Z��dC�6v�ts�K}��� w�p�)D��@ ��`H2@I&Ñ��~�Y��(D�ܑw%
�e��&�z~e��*D���"o[6f����Q�'���r�-+D�4
��ӢC[���#��H1\�t+*D�����(��A)v� �9t�<A1+(D��xw�&���E4�:����(D��)ªԄ*w�Ua�Z7m(�\c�h2D��Z�`��e� @͍�e�l0 5&=D�ܩK�DQ~��v�K2�,̳Ѐ<D�8q�7��iQ#_;^��`F�:D���C�G�U�V�Vn��~��ճbN7D�L3�-Є�nU!eM����-K'A+D�`C7쌖t`LGł�H�x���/+D�dq�G�4u�Y���6g��5b��4D�� pȹ���<J�l�#��]9q�$��2"O�X�)ޟj1��Ԫ�8h�"O�X�,R�I�z���:�<$�"O���t��.U\ C��J=���(7"Otd*���fXm�MI"C0��d"O�9�D�4��X��P�;�a �"O�aQ���:�ūP���5"O��{��F�u�ej��e� )�R"O�M��E�n��Æ����"OJX����tul] �FW\��e�"OxH��P�J�L��8|PQY'"OP�pb��JU��q�)�#UF��"O
l�l�d3����ǊLZxʓ"O���3$J(�$@C�'=[�j5�%"O"��1i��:e1�<q90�H�"O"���"ð}h����

S�`E�c"O���4���U�����4���g"O�����#NƼ��� �lM"O��b��Iz��a%"]�w��y��"O�!�@(	_Ա�a�-u�U��"O�t\��gLN��h(�G�y��o�������z_&��B��y!�:1� 1�%scz�8����y2)�"a��C�e�=c�BIi0�H��y2��I�2�s�̌�_u���
�<�yb�&&��Z�.`:1C�L��yb�NL�܌&�X�����ɿ�y����F�h��0�C9!�(@�%և�y�h��V�h��*�vU)�(��y��@�-,����+�j�H�A��yB��]\�JL�#X8��$_�y�H�9�bI��̟�ȖDSNI��yb�H0G�a�����yRE���yR�K��x���	�%$)-��dl�Q�����&K�(8#6�8����y2���5Gnh�W$J�Y�8;4X��y�.�M�̩��D�W1@�"�i�:�yr��V~\-c���Q�4`0A�
!�y"闍qM�81O3	` 90�֢�yr�d�+�N� t5�O��y�^�s%����^�x�ndY�d��yBd̵c 8���R�@,.q	f-צ�y��V�I��OR�1���[lҽ�yh��KU�թ� O	&l�@�  �y�ǋp��|x`�,#2q��H���y�jT�_26Rpo΀�����y¤\�$Š^/���	p���yRʙ�8^�-��X;q�\ى����y�DD�r:�qO1xz���#JC/�y�O�� �%!GoЖ�KçZ��y­�$V
����Ѱn7��HS�D��y�A11�r\1+@ j�6��"!���y� )C��x�S7Z��@��^�yb#H�o��]�f�\�T�&2r ؟�y"����(�)i �M��H!���y�ņ\Ѡ�zR΃n]f|�a���y��ŭun�U����{i�-��N�/�y� ұR��Z���'��"�����y�F9��4�f)���I�I�y�⒮kft�S��̔	UxS���y�g�%��S��=0.ty�s`��!�;�,}v-�=', ��F%o�!��H%���ۥH�<TY�pm��Z�!��?~^	h�@6IXM/T�!�� ����� +�pCpޏ"��a�"O�ܲ�̊<�X��#�
nL�PS"O�rFX�t���'Ϙ!U^��R7"OnS��O�N�V��Ut���"OL��B�8�:!b��R�
�"O��p�Eܿ#o��륅��;"Z���':�F�D��L}��O�4"����a�`�!��\ n���	�'"i����F��x����?��R��Swu���B�&D�x�b?D�PH@�8l�`dJ��d���A	#�I,�p=�`V,$�(]���� �Z!i���I�<����$Ai� �e�;J>Ƞ5F�]�<�eHݒ�M/T8F�em�S�<i�L�d���� �(Q�H�MPO�<Y�g��ؐ�"P&[�I3&$�E�<9q-��d�>X®��(����~�<ѧ�:/(=��/��\AՇ
F�<�5{[6��(,omT�2i[�<�e��#e�X�k�!T$_K�(s*�n�<1��7ߺ:P/�!-d�}h`��@�<Q�Ꮔ;lflڤ���0���[� �t�<� G*y�zy���X3@��8�p�r�<�s��\B@��hJ��sISq�<aF,SV� u ��F�,�Z�9'Dn�<1q"u����Kƫ3�
���k�<��(B�� P��C�%}P �&�q�<�����{_\��8�u�T�@m�<�?O��SU���ڔף�B�<�TDG(�\�����;J�XH��Oj�<��(�U��9sf�lܜq�[N�<�*Y�l�跧6�T4��H�<��L�1�f(b��݋v1(��[B�<�b�\��>Ժ�AR��Q@�A�<!PM�/]�FQ� �=q�"Ys��E�<�#)֓pv̐�\�m����paf�<�+�/<�<(P�4.x��G WF�<	�O]"d�7��.lm���RF�<���#D" @��&\�>H�5�A�<���F[�\�&��!86�Ѱa�|�<�0��%*"D!�6�Ȉ��u�<���=x$j�+��0���i�<�E'E�TƝ�C�:t�A���h�<��G1?ј�U�0qg&-re{�<q�
.[{Fd)A$ϭY���� '�{�<�"�J"F>�"�a'D;Bp�U/�y�<�gF�iDF	��+��1R�(m�I�<��N! �E�d��쎏m"DQ�ȓp�d�:���=ҀS�,H�7����ȓ&��$U�L�e����"]�g8�܇ȓ@�K��ߜRp�J��T�-�ȓ>E�Y���p�4�bs�3r���X}@�+��!_e�mڄ��$8���QZ�L��A_܊(��J�z��a�ȓ��c'\�4��ɅƔ8�ȓs�����?h	� �	"8\����<>
E�soѕ(�n9c�J�)X"8q�ȓ ,�v��'F�b����������A�CJ
(�
�@֩o
���4�P}sG"]�l��Y�w�I�-��,�R4 G�ޢ(��D�goéOqH$��e�"YS§��`�D�6BX�+gD��p@B��S�'݊|[w@D�EDr��ȓ9Kz���LO5r�ܥ
�`̚W���������"j�0�)rB�Yf����S�? ��s/ȴ.�x�C��{�<K�"O����m�c$'
�9�@hT"OJ�2�/#�@1�r�\��<e�p"OP�;�%[S�
[bL�v	\�{W"O��;�
m*̙��̕�S"���"O@���̅�R)�d�_�K���D"OD`�/Ǒk�Ơ�w!�F�("O�Iq�H�u���J�Z"W>^�`t"OLLq�F��T��Acdo�x��Qz�"O��2�oߒe��[@n�m2���"O ����r���"��V3<	:"O�i��B��LӔ�A�S�Z,�ђ�"OdiA�ÕH�J�1B��e!�)+�"O�� �m��/�ʸcT!y�B$"O��ZqjD[���Xv�J�+�`��"OH�� �ʴ*E^�p ��}YXa��"O�Bu�L� �c�j�bGpB�"OFa�­	m�\ #	LQ@r���"ODŻGźj�A@ S��	�"O�IC�S�^X`Z�|�X���"O\1��_&ex	�]>`��U�"OhI�`8Y�Q�`�B�v��%"OtePc��{{r=j�e��m�w�!���'j��eE�4�ţy�!���_-v)�œ1܌�w�]�1�!�	N����*V+-B���@�)r!�D�k���f�S(6P�0�ؠ�!��
�IP�x�Ӫ��#1��UYy�!�JGn�b/�*"�1q�g!��ٟ4aJ��Q�I�V^��t�Q�!D!�$�0W�]0�B�6���3(^"xB!�$�R�tԓ�	11��5�&�[9!�d��O�Q�a̫���f��#t!�d��XG�(ba%֮u�P��N��!���e���Hp두ej��7.K�q\!�D<�n�����z.L�:��߫�!�D́
��,�0�C��`�4���8!�$	|xnQ�7�'mЌp��ɀX !��ډ:G�E�Ԣ�R��2���Q)!�dα�P(Y�C�[g�Ċ�	��!;!�5/�~���ɸ^�2��BbN!�DZo��a�����iY�M?!�$F9 vd��&��"03�e��M�
"!�/+�\	'�A�App/>ܔDR�'����q���g��9��X;�'Q�@���7i���W��/�����'&�xҋ ��ua�,Ϧ/�����'X��B�*�f>h#M͓:�� �'�8��%�I�_
d��qAŎ{�0���'��m����%�����<w���	�'�~9���Õ?r��*P#|4�
	�')��C�X�%�L��0��)��'N漑��B�D#ΐ:@*�Um:���'�v|�@Aɹ��$�g�ߚ�p�	�'��Ha��s_.�`�ƈVz�A�':@h�E(�T��w�G���8��'f�%*�ޔW�V�3O�z�z���'uzp��Y�Jδq� %b���'�Z ��)j���B�$(X�'�-�*Ϧn��	1S���Р�
�'��`r0�� Fwh0�a��9�e��'��"a'�fR������{	pEB	�'��P#[�Mʖ�����]�P<:�'���E�� ?�� �������� �y@(�t��k�-��'��u2"OJ=�(ѢY��[��P�f����"Ov��fl�R�� ��I�SW��i�"O�\@�/S�oW`hi�<s>�I�"O�1��Μn�N��� ėq2�8�"O,t�PdD�m� �q��@'�@q"O��Ha��C2���g�!?"<�:2"OF����Q��D�Dy��KQ�9D��ط�>&�(:um�}[	���=D�8��(�+L�k��ƞ@_�@1��=D��q��BR愡�P#J��"�$;D���k�yN2M�F��;vPS�M3D�l���G)��@Sc���>��Q��6D�`��(�5/�*8˖ ǒ��l4D�P��f�3[�!�T��#bA��`-D�|���3� )��V�l'6[�-+D��p��y��DA-�"N�rţv�'D���3%�>q2p�c�R�I�"UQ�%D��gH@,@tܛ�&�;3LtU�#D�`[�a��f��!�"
J>]&"���N'D����h����DJ3$��j5)!D����)��y��ć�s�¸���<D��`*F*w���S�hZ�jǞ�Se)/D�(!4ߑ4,M�WK42�T��&h9D�d��#�.B�<D��[�7)(�j@6D�P�wDߪpI؜"�S[� 졇K(D�`�!�\i����$��8�Lܹǋ%D�\����h������,�2�&D�����I""��q�&���(D�z �˽1�����G�\dI�&D��a����8kրh��E�� !a&D���wnj�����ę���FJ���y�&�9�>��aҒ[�Փ�
��y"`��ϖ}��7������y2"W~©c`KJ-$o���p��y�o�����.�!�"�:��ɳ�y��U5����������u��&�y��N/kVrH�WΆ,	���j��׌�y!��>$��$S�x� �9Ū�yB�P�3�k�Jt4�r3�[��y��� 7"q��1p���T-ݦ�y��fK<�x��� >�l�J�"�7�y��FNx`�)��a�@�cN	;�y2DD XP�������S�,�yr���2�<�r�aV�7��Eł_'�y�I�Safh�1�W/9�.iä`[!�y2�A.JxF��W�M3�\@X����y��l{�� �ᘔL�`5�����y�K��$b�'"
B�Ჲ@�<ABA��/3���j�P��a@Qf�<��X7]���r�!�H�r�+D�g�<��$������Y�UTDB �Wj�<yV�ϋ���>F���Ŏfx��Gx��1��0�smO�~�z��C-���y�`8�Q����wm��x�����'���O�H1�wI�b���v��)BSP��
�'V�����D�+�\*gGՖ=h���'�l*� E"e��!�х�4�	�'�X�(p��t~����K�RgTmK	�'�np���[�LEr醀ϢP�&Q��'�D)t�	>c�tM _�O�b���'����CE��];j����uڹz���hO@⟼�;S�<��#(u��f^7Ay�P�ȓ��f�U�NCD"���'IVą�S�? �͊�Dڼ8&`��F(����P"O֔X�oO�M6��1�	(sx"�{'"O�\�DM	
t�@Y3,!pzE"O��'i!��i2�����[�T�p��I�\lɒ�֏�<e8$�ҕ>1���$7K��}����r�T����+��t��A<�@�N�M���z�L_�jQ��a�̐}�<��È(?3N�rd��t��e�dOT�<YC�t ��h��om��@� �P�<!�`K%DAĹ*D��;���ȴ�Kh<Q��G#LW��Dd�?-�z4��I>�y2�Ց6X���&��%�0�D��yBC�0[o�1R��P8*��E*��!�䞅cvh����+~Lι��ϛ�Y�!���� �q�J\h0�ဥ�Q�!�6Sr�1�%F�h�a�%]q!�M�~�pH�&�¶>M<�I���Vf�yB�	�������ӆ����	-Q C��.�~(F �v�09s#����B�	.@��Bd�>k�����M	)��:��/LO��rTF�Vx�0�� kdAس"O*	�6��~��ɪ�F���޴�t"OX���U�W n;�E�!����"OvUE�¶^�Ȟa��D`�P��E{�I�gC�� �N�8z2����"|7B��f�BQ��ޚ?(00�
�=H� C�	;uo�ie�.}zdK:1!��O��.LO(u��m��N����AE�FS�x%"O��pCT=e�pȋ�ǋ�YH¡�"O )�ɋ��HE&�y�mA"O r�E�	`�<+�?��q�"O��ЩԱAښcЯ�]ָ���"OK���\A����T?ǲ�G"O��Y�'�05  l�A(I�?���d"O��2��]�����B�z:!�s�<Q��W$l<�ܙ���.@��|p3��q�<��΁Q݌4" &ޫr�~=�@ F�<I�[A�0KΠN)PH�<�tI%6<&��#2��`T�<�dhMt���{G�H	u�ڄ�bYu�<y�G)E��+�M� �kP��n�<��̋����Dj�2,^-��O�<Qoų	Q��=
�L<�-�N�<�a엖]�|�'/�7�����M�<A7O5%�"�y����S��`�J�'ka�Th�0S<�"��--��u��G̵�y�B��/Zt�]9�� �
�V�lB�	3c��8[�@ĿT����8��B�9'�z@�"G	b�6�����tAdB�	�=0�ե��(Jfl�bIA�BB��yCL衇܅)�LЉV ?�tB��b��)�̜�&��*�4��	(����k���S`_"�젆�9�L����,��ȡN�{6�I�ȓ`%p��ϝ9	�v�٣끍Zk ԅȓ
<�Hs6/�;x�`�� �ȓ�|x�&�Cv^�)��:�`��5L�$j�ް'>Ht�3eŬb�`X��4M>11�-�xW2����$@l�M�ȓ4|� bҠ�1��*�N��l&�l��F�z����E��a���O�m���_�6�P	��^����i����J��xۂ�ԐP����EǏ�
܄�f�\1r	W
Y�i*D�/�⁄�S�? �PI"-��L[ ��L�#?	�"O4��`@�#b��+�c0 ��`"O�T�-��*[ڼ��l�9"6�bG"O��"���8p�����Z�s�5���'���b�8xZD՚G#"���9}�hC�ɄE���@@�N�Zi�+�G	%2}4C�-tZ U��.]�H{�ʇ�T�TB��.�ȠK���0����W-�6l�8B�ɝ8.�p)�0&��o�&e�C䉼=]�񀆪������D�%�B�	�z!8����Y	~��8!�CE��?A��IA�x�T"���bF�����%!�ӟM��ū�M����उ��EX!�$Sr�Шa �V%ڈ���ޮ�!���k�����J�����6�?
�!��?b��ڀ�.���"�D�%6�!���Z�\��B�����W䀃/U!�䇿>;�0	%#��S��)����k!���	���[r�r`ĒË,Vџ�F������i��*1���H��Ղ�y�C_�p�9�*�4X #�ѯ�y⬒8s�Z�[vk9v�H`�2d�	�y�?n� ��1�6_s� ����y�ܒIA�L[Ã�b��8!w.Y��y�f��qm9��1Pޑ�ևٙ�y�D�#Ll��ڻ*�p}�����y����
p-��"Ɠ\z����yB��:r!Rĭӝjr��@LO��y�o�/���s�&�#"��*����y�Dn�����!{Z\`@LL!�y"�B"?	2�����(H�C�,�y��#JG:�S5EV�XJ�rB&ѻ�y�HݖrΎ��#��+��Rq�׭�yb.��FԒp��Q�w��p��K��yb��6s��"I=[�^�Ď�y"GA%v�0�Qn\(���Ǥ�yk+\����"� �)���y��E,eTfHi���3����G��y2l��4�6Ș�}��ڡ.�5�yb
_�J��(1lؖ?�S!)�;�yBɈ�[�r�$�2�� ����yb��'I�q3`V�"|�30�y�B�q>��b4�J�wr�qc���y⍑�z���a�W�@�D#��N��y��!�$*"`I�>�4Y������yĈ�F�`l;�'�5�%Ð����y"��kb�]�L��$�Bu�ؠ�yRi�2�z�)#�� ��$)$$[)�yr�:P(Lq��I� ���p)��y�%Bp+`�Ӓ)��bQ�BH���y�Y�(�Đʴ�+�|+l�"�y�#ڔ<�R�Pf+���[���y�A֓1P�K��)�lP����y���RPX�Um�,�E�GC��y2�S�lq�f"N�4e0Th�h6�y+;<<Vt@�nзƚq���״�y�M b;.������4b�e	<�y�m֨ �����
.~D0��ō�y�,�&9�	���̧|u���3/_��ybn�?Yڹ�p ��+�bȹ� ��y"���h��V<�]20B���yŜ�PB`�j��*��u�B㍧�y"@N�9� jӂ<_f��O˕�y�h�9_��U��!B�`H�aD���y
� r�[�g��Hbpa��-�!�ȁ"Oԁ�B�ڐ�d�l��~��d��"O��F� n�x�bJ
���t�"O�uF�ϨS�<�)��� 8䈀�"O�go��Q�(Ps�V&a���c"OH��F��,`�]؇�\�	ǰq9T"O��A!KC�U��D#@ν��=�T"O
U�#�%�@Q��oE�3@��R"O��+����M�1�!U�g�S�"Odi�d֪w��'�\Sv�Ip"O��+�#@:o�D�TA��f4n|��"O퉵L���ybA!��v,\�
'"Ot��WpfQK�mF�����e"O`ma��<02Tұm��^�(10s"O$8�l�#~iHmA1���<rV���"OT��wg�&HV���2D�H�pG"On$Sētݸ��
�Vo`�r"O�=Y2�ڋM���K$�"g��:@"O��֫�3K �D*�5b�ؤ"O�L�C�_6r��醈#,w�%"Oda�G+ч+k���F��
���"O$��萵��eJpc��T�2"O��r�l]>T������/;ޙ:�"O�h��D��jh��ʶ#r;e"O~�p��5���@5���J�"OZ��T� %�$�	�	4�R��A"O:]Y�-Z�al��A���a���pW"OHȇ�\E��z�%�m���X�"O|1�B�$0h�ϱM����u"O�`P���;[��KV�I �8�31"O��c��E�Q���[*S�,t�P"O`�eVy�6��Tf���V�ۑ"O���.ZBI6o�,Lf��JS"O����ٜD���V
UJfx'"O��C�[�p[a)� �Ԙˑ"O�z������A�E��c��A"OA�q�Շm�&��gS*%��	�"ON��e�#(L�F��S�P�U"O�P��'��3� ���e�Ay���"Of	��dy�ICW�
�(N���d"O8�I%*Z�X;:��t��p���e"O
����ǐ71��@�.l��:�"O���R�$`��JA�A�2X��H�"O�u�$S7u��
��XVP"O>|h��u���Zf�Ɋg�x@"O���C��(L�-%Vو�"O�L8�1W�h��[x�;S"OD�9E$Y/���L\����'>أ�C�rl*��`$�<EF`�'FFmɆ��1f��Y��쏞"�n<�
�'(<�ֈ�w]$�	g��(i2�X	�'���yCEP��6���E�����'�hQ�!n�J�p��-����'�$�õ�*,8z�АP0�m��'�<�N��8����'�+KB���'��Xy#��:��a1�ɢ4�*���'���Ai�sLx=��6'�-�N>9,O�}�\���5��.c����d�	E"���N���HM��wq ��}*���
$��=Z�pG�K�Y�@D�3D�9���v��p�B��4�����5D��b�H˫/|�:���7�MIW-/D������X��q�3E�3u����/D�h0BD�S��i���X�#ך��Ћ.D�� %�'��C˘��cḽ1�>��V���I9�C �H�ry�"dŔ�oJ�B�	�~`�85��T���'�� ӐB�ɛ�*��a�N�Z!37�E�;*|B���ppG�)�"��!%@�ifB�	l3�M6@�/k�P���B�2B�&(â�Pc�ğL��p�Q�t0�C�ɏ>���VFM1Q25
�b��i��C�I�_��P!w �\�e�Q��h��C�M�z�Is��ܲ�!B�QRC�	�P#�Q'K�R���׭[<bfC�	$��9��.�)W��P�f˙�	�B�		MBv�[GO �e�ls�j�B�	�xq�Uy`�?z���A�F?�$B�I&l�`P������8cP�B�I�'���3a��>�i`B��C�5u����X�53ޜk6b�:g��C䉑S��們�S
Cj����O��C�l������]�����k��B�	�p]!�G�1�m�u�J�dMxB�	�Dh!B��{�TMA�����b�D0�X@��K��}B�ΕH���)2j#D��J��ܙ3�lz%NӢ`l�-R�K!D� ��̎�J�v�K�i�(M�����*-D��F�؛/�|�s��)�Dk�o)D�`��b7z�2|�g�*a�`���&D�D�&΅W*���ğ�9�
�� �%D�H���Q1'�-)�@]�I'���)��0<q��ʤMcJy�ˆ�.�j`��^s�<i1jr�"d�	�6ܾ����W�<9�؆'�� cnժd!F�˲��M�<i���07�J�SQ-Ҍ
�"�K5HDM�<I��
�N`|��P��Ft;WQJ�<�!�E2�c�i!�pCO�H�<I3FΛSj0��Yc���e�A�<I ��.o�����_�h×S}�<ar-�4p�p"�g[��];O�|�<�G�~z��G��@��}�d�{�	j���Of&�ss����	��d�8��'�Ș��G�� Ƥ=�g�υs�A��'Ƽ-�ɒq����Ԧ̭6y��'�ٰ��S�A���{Tŝh#��I�'���g��$�قS�O�
6�x��'��q��DF�0ZIK 1 p��'.x�����,�(�'6{.R�'�����i�0�x����ib��
�'Ix���?[�ɷ"[1K�(A�
�'�6 ���*� �P�i���
�'e4�K#(�aP�	÷A�b��a�'�α��`�� X��U���9��hO?�#��F��ljA���M�SMV{�<��Jֲ
D���ቤM���SMAx�<i��W4)q�ޟ1���Y�`�~�<Q�k�.SA��s� � C3m�{�<�Ƥ��܉�KNY�]V
}�<������u��}i��8���N�<���̊3�`P$	ז#�)Aլ�A�<��ɛ�(��`���D�����e�h�<IW͈�L������mw\��f`�x�<�4e�Hd��J�LM(φ9�PE^�<14`2 ��E�X�	��ы@ș�<�p�$e/�8��LڠT��l��LU�<�`F�%n�dxF%ހ)�tY�gZG�<їn�u����"L?��M��W�<� d�z.��?}��p#N�9b����#"OИ�S��:R�@"�n��6Ɯ�#�"O��A��e���qH�0��ѫf"O��ؖM�e��H�'U=	��i"Ox!�e��R�� �"�U&�,��"Ol᳃Ze�u�f��6�i�"Oph��V�`�,���Ԩ��|S6"Op�U�	��%��v&T!�"O�	�EG���0��ЫFm����"OT��ϛ���5�t.��7<�0�G"OXI�U�W"Z���#n�C;T�R�"O�} 4��4pQ��H7|&N�X�"O��I�G��O�x�r�+���"O�P�a��o��SK�6���yrF�<cd�ܛT!S�Yr4
M��y�Y($��֯�4� \��'���1��DY�V��@ ��?��pi�'G��0�iD�=Ֆ���^�� 4@�'�������z� ���QЊ%��'���:��G1>������ "0���d0�48�4/P�Cz,T��$
&i3���%"O9A��;kڜ@��"V�FG��"ODݨ���=�l@;��ؑ>;��e"Ob(k��,Yl�0�"D"��1"O
P��G������ąZ�*��"#"O4��]$J	h@�9�����"O���p��r����@C�7n�ت1"O0h����>b�=��Ģj���"O8P����'�jMC�IB@����"Ol9�snΏ{;������v���@"O�E�&#΂�n��p&r�0�"O<���ݸ{����
L �L�" "O0����<u�mY��A��Eaf"O&��mB�b�(hp���+��"O�����d�+�F[� �ѓ�"O  	��ʬ
��|���[��j%��"Or5��d�<8�P�ϻ(���"O%I�ǷdB�STN�'3	چ"O��12d�H����A>bU0G"Ox������,yDlR�Zn��V"O��S��$}�̥¡P�2��C�"O�����-s�6���E?�x`�"O�Mb��՚x�b����ő;���B"Or Gʗ�C�����@�@�|��"OH�ۢo�������K>lN�#"O�] ��Ҟd!.�#B�3��"O��A����LT�;�/J�*~Z�"O�I���$<����L
P�8$"O��D�_1
7Pi*'M�/Q԰�B2"OpTŦR.��d��V��"O�c��:K<��.BxY,�y��Vl��v�ŇWFK��q/@��ȓ�vx�N�&ޭ�lRm�.��ȓ%�&Л�'��|�&ac"�a��i���F��%
s�pvlN,�te�ȓW�$��b�Z/s�h
vD� g��0�����Gi�%\�]���
27�dŇȓ��0Rt͜2s�B�ər�`Q�ȓ^AL����
(:�/�x�B��ȓvg��@g��5*��Q�K�[�=�ȓP����߹Us,y�g�K~h���4�E�3�T�u����`�isXi�?���~r�B�Q�"�	�b]�)�dl���zx�T�'Q�{����t�hƥ�eNhл	��� �XR�֋�I9�
9�d�"O�ys��@n#��!Ɛw[8p�"OS�`�)&�񦭖 B3��+�"O4Ӧ^�i���JD-G' /�""O����ܺ_O�<ZÂ5vs6�(��'+�	^y���au��#q��ŐoWe����'D���.������V,��@X�$D�`�Ce�"{f)3&�WJ�Xb*O�Z�M�&��'�V;tZ�r"O����oB�5��A�S(�
*Y��2"O����*H�j�8E�T�ʔN���K""O�z�eG좁�C�^���"O��R�f�T�N0��e�3U2��"O^��Ն��4!x�qd�	4*2��"O��	������Z���
 ����"O�� ��aK��2��÷m�iB"O� aA��0
���b�3f��\S�"Oz�y�,��Th��@Y�+��(p7�'��	w�ʱ�UR�m���X4�XE��C�+yа���;Kzr��w	�=@ ����0�IFZLp���Ƴp��0���\��B�	�6xjL�uNlc��cV�ۗ)�B�I%vcш�a��k�L%��^���B�	�n΍��V�� }A2͜���B�� 9��"ЎN�&Q@
�;!�B�I�+�r����~��U����0Y�B�I�=Ғ(��&:P��MF�!�P�=�	ç8�x��Am�꘳&E�SU���*uРRw��J����C�w��_�L�"`�D3M��e���N�z�����j&�y��k�%":5�E�ݾ*였�ȓm��+���6�&�⤠�>8�r��ȓ 
��2J׈*�dy�"�>}U���'oa~��JE ��į��C2;�e���O�#~ڃFÐ9��X�Aɝ7�B�@��Kb�<�A�Ȁ='�=&#��sI�ehUKDS�<�t(��v>:$� K�s��#�t�<����S����/��a� ���Lf�<�����45a���:��Ԙ��c�<��hD5=Jeq+Đ|<(A��Ib�<����"o�h[�YK5z��h	E�<��F�\��0G�]bDD��g]B�<�w�bd�m2dlO	�Z��r�LB�<�W<~��
�Cٞn0�#��ӟx��!I !���U�}�Vܹ��r��t�ȓ>�lP��R<�&Щ�F�>���ȓ�Йö"�)dj BG�5f��'�ў�|r��N$6s���$��%7����K�o�<	s��7{4�$B&&��8�	!��g�<������

)��	#�X_�<��� =:xL���"��(����c�<!� �,6\�3/ĆBM����A`�<������8�d�:Gj��(Gp�<�BL#z�t��➒0OP=ɠRC�<	��[�?KB����mRذr���Tx���'a"�3�=�� ��mD
I>�(
�'�b]1#bZ�*�@X׃4D{�e�
�'��c����LhRР��:�6ٱ
�'�n����V�w?��Smĳ4p�	�'�İrW�Z�*�����:Uh~0�	�'B6�taX����L�8I7�
	�'��<�D��I��9��e�;d]	�'}`)ɱ��$x���C7-ֿ4y�p����hO?����6��=�k��3���Yf)��<� ��G� Ab4����@Yl�,�D"O�9��4i��D5e�#�"O1K�mށ �̠����R[�p�"O�Z�E�{.���G\�i۪!�T�X��ğ�&��D�4e	�l���`�<Zᇜ�y���&2Ҹ���X������d9�S�O`
����N�(��8 ���'"O�̪��M�w���0c˫,����A"O�h����XED���J��T�b,S"Ojj���#H(M��`	��$0�"O2���%�.rD�p� ��7]���3�S���'�ɧ(�荨��ʥB�"q�� o��Y�"O��0V��/0��!�V�-4���$��H��� "
X���b���|ږ"D���N\�AP����S�2��=��d;D�t�2.�*@aJ�mS���҄8D� �&��R�@v�S =�-��0D�,Qa�N)V�����g�#�H�dk�<����?�I>E�4B�<v�՚#*�mO����y�D��@ip=y�ϋ�x~��X�l����&�O�(�!��)h�lifQ�͈��!"O��Q$ԯ0N��bP#�?Gg��X�"O�|)�	$���1r�5 gX �3"O�����>O�~��ASǆ��F"O��Z�=�hȊ���+����E"Oz�*�k�x\(#&Ǣ*���UO���aL��7ˤ�d��#�-	��mJ<!n�6R�NQj�ψ z��ec E]�<ɕbȑv �'$%�x� ��X�<I��57�p5�Fo�h�/XE�ȓ;\,���n'�|�ã�y��Ԅ�؀��+�H+tep�-{�$�?����-?��KB'��x���Č�XQ!o�<Aq���I�
��V���$�Q��ԇ��^�X���G{�z,XE�,/(,��W�He�@��x�C5��V�zl�ȓo�"� VC�)mR���)�&fIZ��ȓy?�Ր�Iʷ	�p[�+�W&х�
{�\� %T��)�EX� �$!�ȓ5�BT��M�;o�V9@�M9
��D{R�'-��֏@>=S�4�g�8fB�H!�'��չuGT3	Y7J�V\J@A�'�b-`P�S�@Ӟ�q֩T8h:`�
�'�\��G��<|E�ty�/����
�'�̽�G��hv�d�� *���
�'F��C!��7��d�q��=)���)
�'Ap����2=���X��?���0	�'kRPz���r����X���\3�'˼����,�`�p�	̺Q�`�ϓ�O�K
�e�e��Y!V��yP�"OP]�V��=b`��Ѓ{�2hj@"O��v��E��Q���b.��"O���pmђ��Y�Sˀ�6,���'���e�Ǯc���A�`$�0��M-�d6�Sܧ?�\Jp��~�0�˓fS�5����?!��0<��@
��~qc5.�#\M�UQ4�X}yr�',�	����J=Y#kE�:����'�V)ӷ�Ǎ1w�hFm�,L��;�'+1!7j'E>�}'ߠ4&��P	�' ~�eK�g�<�R��(��c�'�h�E��,f@�
���qFzm��"O&H��J[�tV@���ؑ�<���D9�S�I�ɒ���' @6�dthMR6�{r�W�� ��1��'`x9���		2�!�� �m�PƋ-+�F���m�1kDH�`"O��&ld��1�©3l X@�"OŒS,�7bծHysD[7Uj��"O�D2�GWPx��Ȑ��iEz�rg"O|���-�}%�X(�]�#BPd�5P��D{��	@-u[.,��X8�Fq��.��Wc|�\�b>�'2>l�� `�Ѝ���5�NA�
�'���*"A)x��Ô�Տ.��C
�'�D�j�	B1:\���\+�Zp�	�'���SŁ[�JB���'��uؾ1�	�ј'E�8���4�T���'T�=�@t���hO?��G�!� X��,�'{� ��� iy��|��OK^�� �G'4ҥ�S�PĜ����'�ў���X�����aM+Fs��8C`0>�B�	�*��iRA�N�r(X��%�1�B�ɄVK,!��)��4����ϦH"�C䉟`FFp���9��}ذ�S5����d)(�r;$o�d���F�7VZLL��~�������
� ��qRoD�N�Y��m8�'�S�' l��K�-P�H�hb��f�t���'���y$�J�<�4�x'	^(5�لȓp̮urE�\Pt�` &o�*~��U��\��EC�*B4�Z!��"1��y�ȓ&1��)���2a�=ZU ˜|�"��ȓMNa��*H�s��`x@�"���I�<Q"kD� t`9��J,X�a�B���hO�U�hl��l
pE��Ι)$�6]�ȓ.�P��^4Z$��$gG=3�L=��A�ʘwE���$C���a��q�ȓP4z��$�@�Q���>��)���|���A��!�,�B���k&���>� �'HY�@�����f��ʓs�����0Ml�2o�����=��Z0Ұ�u��":����@�H@'�l��Q��@���2�`M�Dm
��e� ;D�L�Ę	"A�5�2I�x=R�g�7D�̫�#�#j�P��ҰP�����8D�T�Cc�=O��L3�9Jގl�l5�d+�Sܧ%��su�B�m� ��T�<mp�ȓ6��aA`��g|N�!��ʋR�=�ȓ)�x�(��ͺ0�(pt'R�ɼ�D{�'�|E����0b����gL!``(���'��|���PƩs�n[��@�s�'�l��G�W[���e(���D��'���SS�g�`�����=�����'�Đ�ņ
�V%d��@���;@�L��'�x�� �<U0@�[�2'�|�
�'X*����O;:�J|h"I�)~���c
�'�詑�.Q@&�����$o(@ٻ�'{�4Y͙�gzTq���f��'-=�h��ˮe01$�.���	�'�4m��h_>0S���@E�V��'�J99ЮN4y��[G��U��
�'b�L`���4	8���%bLʤ����?Y���	�W�>���Y�U�\�F��e��C�� �>yq�ٹ!��(�J�E�HC�	�>�@K��3}�h�7�l�xB�	"^�� ��?Ϯ�"Q���b��C�ɚdl}�&�υi+T-{�C���C�	�iv.�:�_�-�D�rb%ӈaK@�O�=�}▊�&k�L�@em�&[4�"���`�����Ȼ�+C-1IĈ��{�$�ȓWPl�(�/�~D���B��H8�ȓ�����B�0E�ܐ�g��-t+0̈́�S�? jY#��λ'����Q�]b�ɚ�"O��S�X$|�uPEb�'�ҙR�"OB3�d��d ń9���E"Od`�g^�1i�5�V�S�v�-y�"O��
��#v��Q�@Z<���"O�1�B�Q��͚ "��T��"O��y1d��H�H�(��	&xy�!"Ob����&�
E�e���)�"O�c�.A�{�@���P�-T��KS"O��Xd�*�8A:��<gA}1s"O���Ʈ�=BF���B�7$��I%"O" C�I&����I[�#�%z�"O���	;�����E$�	�"O����*��U�k*j��q@4"O��W���2$��Q	S^��}�"ODP�6��@��Y#\�(, �"Ox��i�7�8|#��Q�Bwġ�""O�aD'�DXj �@C
�k�"O,���] �\�P0kI6[$\��"O�8���D�3�ŕ5C�4&�A"O*xC�&�|�9����-Pd"O �а*p p�Ӂ �n�.�J$"O���匦. r��Ntn�
3"O��aB
�5i>иC/:;sp4��"O�4��%	@t��x��V:$>����"O�!�T��-*��p"A�� Z���F"O>E{5��!*h@�!u�͔|=tR�"O�( у�%8�z�g@�=��u"OPE�B�	�n��j�H]3)Z �G"O���D��&x��1��]B�I0"Oԑ��ש0��%�-�4 1"O��1���@�N�)�'�1>:�k�"O�$aK�$rH��c���@�H�B�"O�yY��ZA����j�(a�qb�"O�yc��N���{�&Dz	� "OR`3rF�>�x��6��_?�u�d"O*��3�
�ye,X��!L�ڠ"O��2���(]]l��fiXp9�Q"Ozm���: UX�S�9TaJ�KQ"O�uz��'��!B��ں0��<�"Or\��nШT�p��H̥3��\q�"Ob�*�	
c `�e'ڀ0�q)�"O�]!G˒H��i�å�@�D傐"Of���N�[A2\�F��+,�$��"O�����^�u12�j Ý�Q�\t�E"Op,��$�52�ʩ*�a�4Y��i��"OLĊba�d�\Ju��Z|�
"O���j�<�t�X�ꀪ^M��d"O�5�3$�"�TX��W98E��C"Op	��J��j��\�%a^�Y��z�"O��L�|��Y鵈��|YprX<C�I<C��$cAkU:.��yx��f)C�	�?�r�X�$O�н���N�X�B�Ʉw\ε;��ۡ3pqcg	_�:g�B�ɔ3���p ��g� u���G�pӦB�I5w�4�Э��-�&�B��! M�C�=>{� �BϘ{�H�!P���tN�C�ɋE�ݩ���I�֘�0,ٺ1B��'r�-��
�ĕ%�9_�rл�'����V��/c��1��[R�V9�'�}��I!+��	�f Q�K2ĝ��'�lh@�L�R��y��l۝0���Z�'t��C��5���
�e��,ؖ�a
�'��8�Re	u,�P#Am��*�m���� ���_/w���r�
�D�A3"OR�
��"0W�0����96Tk�"O�8�t��6S�3���l�z�YU"ObI��F� ނ�R�j�2�"O���(G+0JE�d�yn���"O�9bS��y j� G.J^뤅�#"O�	�Ƥ:X����/r�Tx3�"O�D�E&ʝ|���4�Ǚ7�] �"O�8���.}��(&��78̨F"O����U�D��'�� �\H"OZ�Z�mM�kvf��^�
��"ON��K7wVt%I�k�{��y��"O��F,,�$�Qp�M�����"O��WJV�i��RTj1p�*=a�"O��	���!Z͘th�
�����"O>a�W�5P$x�J�g 3�F�k"O�a��AT4_4!pe����""O�5@C=7x�dö��l��u`#"O̥�R�J+kUt)���'�8�x�"O�p
3
�bվ�*!Ϟ-�@���"O�����=a6���mP�N�b��"O�eA7�ѨUF���v�5*��Y��"O���2M�6<�*�;VPz���"OV�	p�m>�U����S����"O6	�$ȅy���b��͞�@p"O�� $�դ�8UIq6����U"O�B�I�RIHi�IT�C�"��$"OJ,1�ۢ?�Y`Gj�� �*�ID"O�3c��~�֔�AI�g���+�"O��� �!�M�������"O0{��?fBRyc��-_��C�"O�(b���v~�\�g*�d$l(X�"OTPp�Ύ�R�p��ƨ
���a"O^hj�AύX�ai�Ȕ#z��"O|RT��4:�Nl�P��\]{�"O H�@(H�%m��x�G�+�Hu�"O ;r��51>Z<�3�';�EC�"O��BA�^�D�ZR6�Ҝ6���q"O&����Y�+"��0_b3�0�a"O��X�n�+n�<�چ�]qK�%��"O^�2,�g��@��A.B��Y�"O&`���¨00r�4��P7��""OJ����@�Y��Q�;Q&����"O^}q��,@�͚3�	�
��`�"O�3s�1rq�,�c@�F����E���"も7�"ła/� R̈́ȓq��ī�iضk:	��9XF>y��i�BJF֏KU�ݱp���iML=��nF4�,īQ �ܹ�HE6R�A�ȓ8x�� �	+���aF��8]䱄ȓW;.�9��!|�A��߭D\5��9�T��Ŏ�#��s#k��B�B�<i7&M):4E�%f5\�~�yD�H�<�&���&�Z!)B.>	�c�YZ�<y��e]Z4X��J�#�����T�<��u@أ�&HԛVcGu�<9��?�����%]R��I@s�<Q���'8B%�`J��5���1��Tp�<� '�%[�8��V�ћDb�P��p�<�0�3#���a�*��:3p��'F�<yGb����b��ʠZ-T�b�Eh�<�t�j���ف&D�Z��A���`�<��B��[�9%�ܤ$���э�\�<YS@�%���-��N|Q�A�Z�<� ��� �: ���(2`(���	4"Ol�P�S�s���JD�C�(m�ɹ�"O��yvh+�}� .^�S�g �y"$�I���kG�bIf����yr�L��3�@V�����&�y@W���q2KW=J�ļ�%����y��R�H��5��T-�yRN�i�r�#��#�8%:Dm�<�yB�Ȑ*C(u��-ƣc)�D��(J��y�)��? H�҇ =è��y�	65�J(X0C4\�y�k���y� �t��[��X�� V�
��y�E�:ц����ا<�\����y��N
��{��\>1��A�bV�y�ɺ-#�p���0�ʉ*��	�ydֻM�<X�bE�+j������yRBD`p��7�'R霁3a�W��ybJ z���W�D�,}2��>�y��*�d1+A" ���y�π��y���������>c 6�[�+��y�iZ�;���!��X�lTI
?�y�s� ��o�>g�eKv�/�yr���.��
!Gȇ^�Aڥ�F7�y.� 84A�P��PfpUz�̂��y��0E3���P �
3�m��ў�y�M.[���S�#�������=�y�B����<B4	7w��iC��ֱ�y�A\F�A���twb��H���y�@�_��`�� )h}١ī�9�y�؎�ؠ��i?L!2�+T���?1�'4HD���C�^��26�]#�	 	�'ՐL��jˊ][���e%O	��	�'yx��"Z2TYd ;�D�H����'�UҶ$ǈQ�|��Dd�'mc�k�'�h��A��>f0�b�
E$3Kl���'q�<KQ�[�^B6���ˌ�(ǒ,:�'�N��2��u��2%�xV\Բ	�'/v�@���r�����Q
p��@`	�'\�I�������� "��]�2*���;,O|���$��"H�a�7�P3 ��3�"O�Mp��ҰK��4���
t�\�c"O�4iS�	k��r�f�34nBuX��'��O��k �޲xE�ŝ�KT0�Ǵi�ў"~n�e���{D-�nC�P��5��B�ɗb9��@`�ˆ&�5 3C�" ����M�O�YHHE�Ϙ���Ѷx$�ȓ9��j��Ʊzv]�e���&͊̈́ȓ"�9�a�O%�-��)��iy\���+EL���Y,��YŭS5��X��)&D�$��<
/�m�EGމG)�ȓvTf�sMF��r��n�Gx��B���	I:~<�y0�̓�r��"G��!�M�`6,x�i_�sR!:`��- !���O����N����������"O�j���#{����·m3��X�"O�)�ĉ?�LH�BW�,0:���"O��0 �Y�F\|-�X$j��"O�%�� K8n� J#\�HD� �"O��#�rS�tpfh>��8�2"O��wF\�+��ip(��8`��"O|)`3��4!:�K �ř?�lH"Oixq$$�J� -��&�M��"O��k"� ���ul� l�j�"O�\H��ؕW��!8���0"O� ���s��kY$ձ�C
j�F"O(��L޸M �p�bɟV�  R"O�U�C)@�!8>��p�'�5h�"O�,���]���!��6� S"O< ����͆����H�G�5"O
y��AX�lUX�ۋ1���p�"O�(S��$���ɷ�R�*6�G"O�l�猈�)����'	L��1��"O�󱪊�Av<9�(J�t�~�Y2�O�O ��䑄x���תz�	��Ưf�!�ă�=��y `X
}j" ╏�<.�!�$C1�V� bᗼ$n��-� 8�'ua|�ń�!�>a���5nD�H���yb�^�RC>�.C�t	�Q:s����y��Q3�^���06n�;�.M�p>)L<�`x�M��!��Z�أ��V�<YQ&��np��ɚ�XK>@`�F�W��M��O��|����99�A3��3M-d�P��P�<ɣ��i?
8��e2M��2$��H�'$�xB�[�aT�-� ���a�0��Z�'g���j�u�훥$K&�"t�'�ў"~��J7_�ʕ�2�Ҳ6�n��H�|�<y��P*��У���a���6��'�a{R���=�̐�'/�L��g�/��$����I�����d���!5�T�&(S>�m�t��;M!�$0Tm�W� �k��
fFX9xa��,F{�����'F
���RY"�u���Ȝ�yb��:-��� 
�h7$Ix�˕4�y"e��е�f��3e}X�Kbo����=�O�Ʌ>��kՁ�1f6Y��"ǬYm����>����u������&
�b�
DY��hO���O�fNëZ����C�/F5v���"O(���54|͉R�F!�8hG8O��=E�4�O
re�qЕc�u��ga���xR��"J(��{����rv��|��p?����=b�0��"A:���B�RK�'M"W����0h4�J�T)@�&��'(�X5"O����Kf9Y�d��hQ[�"O�Mi���bV99Ј̦i�ԪAO<���7]<��P�Ӷ$,|���o��OQ����I�_�$4nXl�*����9o�C��?�:�pE톥(>	P +�I}���
�'�|h��u�%(C)O|2���{r�)�)��AQ��jG�="kz�z��V5!�$R���
1gܬ�E�31�Oz꓿ȟ\U�P�ۦ���d%R�(v��0"O��%K��;���c��2�"�je��v8��Q6L�1=������%� !�2;D�`��H����IAB�5K뾽Z�&D�`����3�0� E/ٛZXf���	#���2�GH]%-K��h$b

 �ܑ���'�ў"~"��U(?"0�5�� q�̑ 	���I��HO?)�g�Ѣ�v}��lޢI�D(���-D���K�5��ه��;5XD�x�!,�d-�OX�q��H�7��e,FZ��]ڢ�'�d�`� M���J(g���@憋,!��7��yH��7�x���F �
 !���{�b}!#�" �p��r��T����H>J9��蜗.e湐sK�;v��B��&F�����h��-���j �Y�8F�B�ɭ)f����]��'B3�B�	)O*8�
K�*�:! �i^8��B�ɾ~>�m�U�3ng��/	��B�0>�P+g	�:	��$n�$qo�B�)� ���bjN�&6���3��P 6O2�O�S�g~Ҧ]�L�dZ�J��������d�C?qӓN�1IӠ��^LR�n�v�<��IP~R�P�h8r	 �^+:Z`����2�p>�J<�el�U��� u�D�V5K���M�'`����ؑ7DRal�!&��� 0B�"O�Ms�/ (�B�w�Q�P�����'�Q��ɷ�ݠ:^ �2!F�?㞝a5�:D�L�!��BXjR�	�|�CB�9�d�M��}R�ēB���!aO�n�����@]F�!�dDG"V�2�%�	��J�o_�fyqO�7�3<Ohh�i���=1�h˞Z�dM���'`�'0���3�S+�Z��$��5�f�Dm+D�Hy�B� *���s�,R'�3<O��}2`�El��n�;�J����y��LA(r-���	�	6�Zr�ܠ�M���sӮ0�d��}���� �K'@���"O�09�����s���&X�P�"O�uUt��1D� 
>��w"O$���B�1{l1���]/P� �"O��#Ύ���0��N~�F����'
�'c��N%���s��	*SPl�"e ��y��Ɲ3�P�у7YghYKN�
�0<q����&G��Ɉ�K.M�"l���#!�r�V|u�T��r������8�̓�HOz#}*�iJV����4,7V����{�<Y�B�b]�l��N�>�`�ia�L�	B8�t	�D�V Q��FU�j�`���$4����'E-힕k �������V�\�<�O��y��ඥV	��БT�Bx��Exb�Ɍm@z�%@/�~�C�M��y2�+i��!S%�<Q*H�l���yDŲ)Al�j�AN+g>V転��y2LҚq�8����D b��y��-���y�o�1x�س���]�aBLS��y�`��GN�j&(�IP�h��c�;�y���	ox>i�,q��� -��y��.�X0[&C�q�*D�� @��yB�!b�� �Q�T>e��rƐ��y2(՟~T�q����K��`R�j�%�y��.M�9&`V-B�x���#�y��=�֍��
A6p�����y�aNB#��Ɂ��Dd"���.��y�.��:p,��IƯ5��̋'�B+�y"�Ԭ��hQ�d��1��G+�yb��8Na��p%$O>cZ����T.�y���#GS�Qm�=.h��рM���y���*;O�	�O�,�~,YPb\��y���^o�p�b��TJ�J�%�2�yR��2B�2�� ����<	�F� �yҧ�����sf�,�LX e!���yª��\����f�1!��J��-�yr۸X��=�d�+w�|�0���yҌ�57�raY� ��D�fica���y�L�$�������Abd�@����y�-��b�V�k��%A��ER؆ȓ.°5K�'�$-3��x�)�?Rzb)�ȓN����[�F��*����5f"$�ȓ��	фM��_�N܊���U �ȓ<��([�{�FLP�f����'G�mb��6Q��A�[��j|�'�֑�d���P�y�����O�}��'�H��B��,Z�t��P
$݉�':���'�oH��y��O@.Ĉ��� ]�#e��	_����@�$g�p��"O��J�)�MF����A�,G>� ��N�xH �x�.#�,p���Yl1O>�#f+�r�ԕ�!�7���7"O�E;�	�)y�0u`��ܼ`����"O ԀTN�8s����T白ln����"OƝ�v�&|��� f��-+��i�"OD�BT�y"�C�HW�D�H)�"O�a����L�'_�P�"O��& �0R��ph5�R�	*'"O��P4 �:z�b4BaΎ`��8kT"O��q��ڋU��H�a�91�D8u"O�̋�EO�5L��A���!`$���"O��"�H�����#�r"Ob<�k��.�@Yphؚ��%٦*O�yB���|A�S�]8`Wt���'G@��2,N�J.��i�(����(�'N�h� U	}8r�&�K?q�9(�'�Q�#��>th�@B\]A�'�������m�����J�J�yy�'�J]!d�(��ؐ��ѵ�r8	�'��������0�m�Ђ���rA��'Š��'�͢'��� ��]n�
�'T����_> ��C�'n��
�'$I2��
'}6=S3�����	
�'�a*5��;P�0���O�1xʰ)r�'� ��'��=�@�I��&xѠT�
�'x`�b�ǋ�d|tiw��NI}�
�'詩�f�0>1,uQV.S
��4[�',�%��$���{���5F���'������ 3��8S� 9:�p��'3b�Cf/ �-�.pV눀;�D�	�'x���4��Y�G]Y-��'��:�Gŉ|�:%i�˕���A)	�'"�Ui�1KVC�2~�V]b	�'��ۤ�0$��XA$iu���`	�'�����MՇ�zhC�Q�a��%Z�'V���G$SV�-���mW�س	�'Z-��ܲ/�pp�1�њ)A�4H	�'�>u���N�P����!�'.Cnk�'H�$�o�/8̒u���loX���'sny���1��Ŕb�^��a�TF�<�wB�� P2J$�27I�}�<�G�F�&��ԣF�U�a�vM�Ԫ�w�<�7��"'��Lr�`F&A0B���p�<�*Ԑ��0�b��"D��P��Hn�<�6oԶa���Rvl�XX��s3Ac�<��!� ? �J`��$�x�c��KQ�<��M
J54qA�O�������R�<I�ϊ�/�pH�B�j���t`QL�<q�M7Z�ad爞X���C�U�<i	Iy-pS���$�>��A�k�<qB�^�d��㓓C�4)3F�o�<)�&�.N��*pW���A�A�<��㏮p�ƠK�"�6}XTJFˉ~�<�3��W�5�� ��U�ƍiю�|�<ɠi@#�bB�0D��kQt�<Q��I4<2�剴��4���C�OH�<��$�`E�a��ϽY�����`�S�<���P�8x
��?�	�Pl�S�<���"?|b��5�N�*��}G�K�<)��N�N\��!O�N6�\���O�<���זb+dq���ɮ/�F�r5�Fx��z%�X]<�����g�p��/A�Wp��jU�
%�y��E��\����N��=���'�(Oy▢D��T���� �50�	ǝV*8�k!g�R�\0d"O�ٻҫ/X��E�S���	w�=*���5��$>wʄ��h���	2?�dA�Ԉ@�^bv\z�H�!�Dڥ?dhܸ��_�� �cj�{�������TH�kћpJ�qc�'�Ā�C�<&96�1 �Z��u�3lO���6�`d����J�4ir�f='l�SUN��0� ��i3��5�R!b�<�0h��� '$5��JA��#�
ޯ5�S�aE�@r1��!��#K�<�R,\�PS$᪂"O:��$&*��������H��	/r@`H�Bi��}�l�4�ފ]�Q>�w�"���3{��T��C���ȓx���3��oX�)�$�$ƪ��-�8䎉�����w@TB1�
;��O�¢����l����3V*�Q���'I0ES#�X)�0�;6�Q1�t�pFT
̞T!2�H��,Q�D�W�f��R��Q��ڰTd&48����'e $`č?y��xe٭	\J�Q���F����sS��f�Ja�ᅣ�yb�].����#&�[�*0��e�;q̭�"�.9nT��";[�G��U�u�Y1g{�]	���*����r�%D�Ӷ��T���P�w�	@GΔ�l�f\+��^>!�+P�v�JG�՟1=��C�@"%�(l��U�0=�S��V��)A�'2��9V���p�D�� ُe, �٦ �`%��yCdE���/_ܬ�U�W�aTfT�<�u��bSvpɇ$�&	5���M���'Y�4{�ke)`�9K9��;C�6D���U(8��ңgѢ-�v�#×�X����m�.9}9�"-�;1tc?A��O�R���?<�(�(�4Q��}�"O�<ҔF�28|$ٰ퀒yB��Ώ#Lj<<�c�F�	�4)��k�axr-��$h�&Q�u��z��Ұ=!�n:A	p]�2*ڏ>1a �o<RFPa��n��{����ц�Px�ɖ&��&�*`���QE��'�rX�ǡN�Yo��Z`�Z�b�q��=�#�;6DrЬ�,0�P0"OLsJ�g�| u��5or���T�V�L=P�M �SnY��h����8F�c��1G�my���z�!�dޝ������w�X @�����DFA'Z���B��0=�'��p>�9��
0@���SE��mx��[U��-{�ƣ܋8��|�⍚4��l:�〛�y�)؉u���b7�I<5�E�e-�+�yb�H9.�0E���&$h���a -�y��'<�51���ؘ�j]�y2�O��`x2�["g� ����V��ygL<|"h��V���V���y���Z�]qf(Q�Q@Ż�D���yBoȼV� Y���`txx�%�*�y�l�?Ay��Pc@["Vd�tF�:�yB致H�XHl�H�^���ڂ�yr��!@T��e Q�B(0I���y�̗�:g��I��:� 48$
�y���3$�9��)92�K�'�yr�4z��x�CR�P��yY���y�¼	��� �ōK���(B��y�&��Q���(@�|)C㑻�y2.I�Y!�@+D��s��1Cd���y�G�?2$+�Y��rhiS/A�y2�����$@C���r�V��y�a+8�Q�G��i����%���i����9�)�S)Q�>�p�T��̰!n�K\�B�	 S{�Cg���E�`����.� ��|��2+�c?O=�1K<kc�ay��,@R(i�s
O�0��§ǨЙ��T;$n
Mhe��J� `�,��0?�3$C7�,�r�Ռ�L��qF�D8����DJ�R9r����Tq�τn!n�e��^�$	b�f%D�th�h�]��C�,-��(�� }2'
TB��!�����E�4	ԩ0̭*f&_*'����e��y"�Q$_�̹g���%�ܝz�'�Q��ϝz�"��(Tp: ���y���EΊa�s��/J��dʛ���?a�a�F����V�B $��`Pf��Js�� �[.k�&xR��g���䗷]�� �@jp��mS�I�D�XP��р5e�$��O�A�"-�9l��1�J�5��܁\w�vhjSK
S�L���+J�h�j����-+QF���>�/J�ᒆ�	�\�!���S��'	|]Ġ�8BUX �x��#}�K��v��A]�+Ӕ\�A��a}�@��A���JN��G�
����!^M��W�47f$�I�+���դ�x�tæ"���,�|}ba�	,fwJ�f
3���X�ℨ���b4����q#��+WGʶE�
`����:{������,XV>�;���'-
X��	�ckaxҡ�Y&���Ӆ+e�1�Be��Z����VB�,?�:U�'�n=��/[l���)B�6ьl���R�C^�MK��ߺ�Q��?���*�`S�i�P�:��r�'4��e/T���D�'�l �1��N�P(�A��Y`  �I�4���nK�BpL�����PX��O�ȅ�ei�E`�%pR ��m�|���O9:c���kbx3�ObI��(�s�K|bEG��TJt����1�����VvLc!ė�?�lͬS����|�<�IQ7,G��'���Zz�@�p�8�p�j�z��ī�<�N|�5�B�R�q��&Dߒ���KX�O\<a4B�E�03n��h��1꤁EG"ay2&�2�xEZq�P! ��D�sO �Z�Z�ۤ"
�' 2<�
ա�,�D~2E\"�[��<x�p��ǯ#��OrM���U2���fVɡ%�L"f:�)��F�g��C�C Z��Z��.�O�l"��bm@�H�6�*����Z�c���6�t�j��
�ǉOG<i3�Q�cK^p"gg�a�ap�'��C�L5Q��,���H)^��!X,OF�j�Z�!�r�zO��|�ƥ�+5^0��2Gα9O��<2��B�I�$��XSuÒ-�j	�͒��bD[J��2�g'x3��$?����,N�V���JU�0��z��$�OH�e���z2x�)�D�\��%kJ?��X���߰?� (��)����Q휢:$�d�S�'d��*f*F�v��$>��T�:�Vu�"<dRT�Q�%D�jf`Sm��k��iX^�Z�c�<Ab���'n�IA�+=}���{#$<0Qb�6yhиf`1!�$��J���k�_��b���4�!�O|�Bc!��lJ��qOR����3����*�%&�����'�V��K.q+6�R�l@|ef�sC��[���"�"�j؟ �1��%x����:�
�j��5O �3'�d�ҒO��S���s��-k�ǆ/��TzC"Ob(�N��]ɼM`�+F��h@c�>���׌E)���?��EB�m�dA����"�!.D�\i�HM�8�td��r���z�/D�`�1f��J���Cg����`�"�A*D�̙��P/Rd�2�$��؈�+D���$ʸ.�l�al�D��}��(D���D�N�t�p�sDE�u����g(D��VG�J�ͩÇÕJ�|�pF2D� ����ڄQ�����w�1D��!�$�D��p���΅JӐ�B��=D��;���T!-:q�"�3<D����b��"䚄�6��xX�(D��&�	;�9A�P�e\蕘7C)D����*6.��
�B}h}�'&D�dv朁#��%�a.�J|�0�AI$D��+fCV"*Π�d�H&at��"D���4�J���|���6�ʘ2�<D�$�ō޿@C��G9��h���&D�#����K�`(*3��H�@pAE3D��ĕZfr-*���h4<XA"?D���A�2h�x��s�K�%tFq��*6D�p�a�&Ą�W�E�JR �4D��؅��bm��b��
�&�y�B4D�T(�EYi������J@Fa���3D�8�t
��K��T�p�d1a!.D���W.�1���Éܙ�R-��/ D��� M�;<`}�3�֙���b�+ D���� 	�l��3񋋯)J�5�",D��q�AJ4�l�x!AF���g*D��(���> �ջ����iHZ��Q:D�h�u`d�C� P�E���@!L,D�� ��㣪,.��1@g@�1�ҵ��"O�@R�Ƅ/]h2P���|��Y�"ORe3��A�fZP2*R�('�25"O�PJ�MC33U�) $� >8O�qrr"O<��A��p��Q3�N�D>I�""OL�P�F��@��s:̅rU"O�P����k���beKC"bk�"Oz� ���$�, ���7�Q�"Ol˳+;rԬ��%"[�F����#"O @S���4��(�e�G&��Q"O��+զ�0��a�<�F�*V"O����J��n!�98��l�d@U"O@Pئ J��P��9P��B�"O���aݜp��9�/�)f��4["O�bVFթC4��1�[�tv��� "O ��!o�b94$�".�2d�k"O,��R�?%@�D�Ӎٌ;��M��"O�q+�Ċ5'؈y字�5{V���"O93+�}�UB�GǶ1Ujؘ�"O�З��'�5ñ � O��Q�"O��{���C���(B��%���y2-жhqn�C1E�!b~�sf����yb#ʽ{X8l�A�E�Q�N��%��y�� E�S�Kك8�D}ᅊ�y��>��q��M�e؅.�*�y�F�A�\((C�H�sS�,Rd��yҨ�*8�A��G�:hr�u�B�L��y->�@�ōՊh�8��#�y¤ظ<>`	�鍕b�����C��y��;5���V�Ϲe��a�	Š�y��Я)�} ��	!U�LL� ���y"lКM���Bi�&H�������y2e�"d�X3`��8N�̰!��ݼ�y��B���E#��H�ȁy���)�y�`�-95ƕ�D�E�
�Q�'���yRE�,p���JZ���鈟�yBF	)����6����	M��y �_����/����A$O�yZ�
��D��}��3t*�+v�"e���&ucf�ʄAϚ��<.T�$��RT�u�h��͡¥��1�݅ȓ8ĺ(�ڨ= �t2�H=?.1�ȓ� a	��ˬe���1�i^�Q��)�ȓ3��x���*,�V�A'�N�krv�ȓRSBHiWA���	�,^�Ƥ��s�`�Jգ5޸�����[`��Tђ��b��	�$z�c�a����ȓ'F
ň����R6��jƈ �&X�ȓ>LJ Y�%��)kR/���`��}��L�Ɏ7+�Nj�D�#}˶,�ȓg��(��O�/�M���GW��ȓ#.��s�ۘM��YU��
!�����*.6�V�Q [�l�9%[fS�-��y+�œ�iA |�QV&�2�m�ȓwC���)аO�@�'���``(��\gvs�bŰ"�
���k�G�(��ȓw�\��j\"`ߊ��R�
�ZU����faQc��Q+,�ӷ�Ͱ!>y��;�^�ۥ���'j���,HI��#�ܰ��U�s, S獷2��ȓ&Rx��Ɔ�t�-0�lʭX��h��!�.t��j�1c�(- �	ѫ��I��2�X�B��Ɍ*F��kR�A�搅ȓE3�  ��Sɔ��*H�����S�? X����1���1hs>�"O�=.���QcWj9���{T"O��!��&^��0��{f��"w"O�����lm���5���4���S"O�����#;j�Pc�ƍdި��"O���/8|�I���@(9�H�7"OB��)2/ X���Fi�Δ	e"O��HG*����QS��."�"L�"O���GQ��	��H��U���"O����8}�ޑ�@Te x�4"O�i��ý�x���aŲt,lL{�"O��c�CZ�9�|��@ɴ7��T"O����%��LES�)¬9�,}��"O�1J"M�=%�m9�M90�����"O�A��;w;��bB,,I����Q"OR1��m$l�t�˄&[�8ш�w"O<܋ר"N2��fkݳp"��p�"O�8���?K^�����5	����"O
�j���]ٺP��AH�=�r��r"Oj��u��cL<i��� J�[�"OtY��С8��4��F�� ��"O���� ��3e� #勵���Y�"O\�i�� �/��d�P�9G"O2���^28��xS�� R�a�"OR�9��8'}b�9gFU�a���Z�"OpQ`���1$� ���>�H	'"O�R�
'oV�I!鍫lxf}X�"O�aD-�N�-�� �H찲�"O�*�' �
X�M#s���j�"OH�F��t0f�3&oCn{�8� "O��kdə�~���[�l1F0X�"O �ôN�*k�T�9 �K^)Ba�B"O�D�g�D�X��0bD
� {�i�b"OX��� U��HD�/�X(�P"Ob}z�/Q�?k��ȗ3���"O�4�'���S�n}Q��RP<􄂶"O�L�O���S�O�aJ ��E"O��� �M+�R �Rw#r���"O�Q�E�9�R4����]M�p�"O ���d�=Mt�z6�ޙJ4�	�"O`a1�(�ZZ	Y��"'���1e"Oh0��Bߏb�2h@�N�.�a"Ort0��S�h��u���?���)"O�Xrt"G�}�������"O��ۥ���nS�as ���<ѱ�"O"U!�nؤO�M!b]+b90��"OL����1$Z"�Pv�:#$�i$"O��r�7k��e��DL��μC�"O�!)�ӄb��!y�#O�o�,�B�"O��1��d�� 1˃��F��"O� �a�_vĘ�rJ�(m�@���"O2Q���*]��s��y�x�t"O�tH ��oL��I@c�l<$
E"O`I�t��>g�� صi�3�<p�!"O���a�
B�S�����n���!��],[K*��aM
:z���"���!�$ܴD6	�ƞ e�:3@�?I��'d�* ��SܧZ��6��<{�έ�`>~7�}��'n�lҶ&ݽ�ʨ���H>r��QR�f+���>p��E�~&�|�AJ��	����$B���p�0��0u�Xo��%���$�U"d�kj�y�F�P�[�a~B�Ln�Q��եY:Eƈ�p<q$��S�r�hTa8?y���m�6L�7��R�R����I�<yq��:5�<@D�K%�6h���TI��ZI$�]�Iɨ-j9P��� 0�3��W�-&Tا/�7�v�Zc"O����C!��]�vG+2��;��[�N<��0bk�O��
���81�1O:��F���B���S�Aǥ,ђ���'>��6���b�Z��uii�b,�l�n ��j�� a�F�VX��P�#;3k�-*�%�>�R�E�=T��#��I�G#����l���JR.Hԙ��j/�Y%�?Klj��'*0��9F$�-�&�����&Z���1�+�d�V�s��;��I..e�:����x�,<�u��(?w�>y�%M�F���b�K(�����>It���_�N1h��-}���7A	���l�{~X�JR�_#PmCT��,�l���'U�!y�ua2���{r �u��SV*�8.c�M���T�	�qZ�x�g8��Oᰔ�)�O\	pa��,���ո$�pL���Y)y,����ΚvF�+��0<qA��
y8�V��YK8�(����j�3�� n0��v�:t�N��M�!��� �n�y�NT��ԩ�#�`�	�GO^�
wdA^1*E@*:��"?�w�V��\2�ʱ>,��z��PB$J ��K���q��`a�'F0�$�:G��R0'��0|R�nL"(%��
�oSY����Rm�P}�̕9{�����L�W}���`��ٛ4Ŗo�ӻ^����#��=xCHȆBLz�+�E��(�����6��x ��'�3�Ʉ:�4P3�C
{�q����6�tD�'X�K����f����4��&l��*�:�H�V�YDyNh1��Q� ��3@jǞeI��R(���D �
Ҁ!#�яF�z�q�b�,�V� ��Zc��`�O`= �ǳ
�����W��[�
,{���*��Ō[
џT g�ͺ(�荖'$+�!V"b T���L�
�.I��OF-{z�pR��U؟�ce�[�Y�`���6W���n#?y�D�"o��o�j�G�G2��Y�q)�6M��p�mF�2ea"O4a���1<��mY�X�SAR�0�d�Z6fRjta4�>E�+L�l��(g�Q��f��33\*B�	� u�Tee0,��o�2 �H�hx��^8.|$?��ۄ�`Eܝ����&HۚT�ǈ,�O���$����Z�!��cK���$�h�hZ�KU���?!��ƹ �x��Rj�=B�q3S/�h�'����J�`��'>Y{Qa�/0.�9
v�\l�d�pE�1D��ʑD�\�l����0�zݐ7(�<���9m[ظ�%>}���ܔ`�^��Rk/ݰM[#jԘc!��*h��5���]1�
!�P��O�����.J��qO�z�ɔx����l�b���pU�'t�J�I �/-V���F�uκlb�Fmf
�ɂ"Ux؟\KG͕%]P�A'��$�zPcG@9O ���O;3�f�O昪�M3C��Rb!L)�l["O�M�V
@tT���= ��ƛ>��e�;wy��?qhd`i�\x&F�r��㵋8D�@�А��T��B΄i���z74D����l��/�>�!��+8θ\��(4D�����9iL��2d��t���8�5D�d��'��tP��qt!Ǥf���"`�,D�`hB�O>V����Dov[��	`g>D�D�K��&���m��d���1D��iV�a�H�!Ɓ�:�l ځ�8D�$"�-Ʈ&���31�\iTD2�9D�{2��\h�%�ݶ�+"B�y2�D/�&=£N}�Q���:�y�kD6|f~��� �.~�A�A�/�yB�ۻ%&�QX�G̦�dt��b��y�9>|X���(DFxs��ȣ�yR�Z_?L!�Ǡ!=+��C�����yb��d��䫷�	(�z�ȶIǀ�yr/Gll����K�
#��ؗe_4�y���H���ZWFK%���/Φ�y��)[�,�)TnV�.ܴdղ�y��<Pmz�����|��Ceá�yj�Vt�1�`��`�c�D��y�G
�� 2a*E��qflE��ybL��8�l"1�R7	_^<*�m�yb�G�8|[����	 D
���y���O�~E����k�R���4�yҢu1Xو @��`p��1���)�y
� �p:�)�zH���@˄�7bT1"Oh*"�R�+h�d�a�ʦ~�IH�"O�U�$W+*�� �Åu���J�"O��㷂�Y�={RK�V�@�S�"O� �N�3�EGi�'k��s"O��:ԍ� 'o�l�g�[�_%�1"O��
%�8N������13�x�"O��׃������Ks,@��"O8\�Q��*U�\�p�G39e��r0"O.Ps��ѶfղdCK=T�	 q󤊾[�5x�ö `Q�͊5g?1O���斖"�^}�b� �#HP��$"O��x#n�,��C���|��TA�"OH���jf𬴁��
�.��@�0"O�}Qe��.>^��J!c��A�� �t"O.$�$ ��n�qC� N���"O�Ei�H�Q\���$�#�����'����'� �*�)�0T����%� K�(�J>��ԠJ�,�O� �t�qx
��2E͓Na�4j�=*X�ߴsV�	�F���)��{V���<삢7M&Р�GT�!�A�Aa?a"�F�=�l� ,A�����O�����b=yF-N�u?f�2#��T�� Ϊ�!�·;B�)ڧDH�ez2�X2J�5𠎅�BK��K�D&'B�!)����Z�	b�O=&���39���[�w���C���4�����h�7�П�?�韠-���� ;�z�� Y:X�<�
w&��y���s�7?q�,�������sN��Q�	�*�<	�фY)8�,�'����4@S>�
����9�h�A4j��I �R��,��$�蟄&h�u���:���O�S�>�,�ȧ�ثL� ��U�p���J�$T+�8�g�)�iW�9�¥q��S�r t0�Pk1!�d���*dcK��M LR���{!!�����0�'��~��!��!��K�;���mI;h����f��+(!��2���)�l�rdi���=j!�D�-�ʕ�S慠R��!J@/J!�_)+T5����$&�~�$kI!�@jG\y�7��ٸ�:�*(I`!���:,�!�HD�d$0���)ea!�K1V��mp�H�-�tMi*̸EE!�	�6 �#L�T��jc��.V8!�ޝe`~=Q��;H� J�k�1!���Y9 }�'&@��MҢ�C%l�!��(�Bb$Bާ+���YG�9�!��C�L-f�A䧗8t�h((�E �!�$�y��96��(�=�u��,!�d	8('�b��(_����)	i%!���0~��ّ g��ĭSB�F�/!�d��`�PI�J15�%����A4!򄔰\�t����">Ƽ�%(ɝb!�d��s`DJ�kO	 �©׵ �!��,��`�@3|z� �emS��!�P�?
B�����u[��xr+9l�!�$��6h��#ǀ U�顩��j�!�$Րs*�"� WC��+��#�!���+�x�A��&:�%@+�(�!�䝩N���2v��p�|����Q!�d2v�V���@�xiT$�F��W#!�$Ӻ?Bi���2cp�2��]�h!��6of��Ҏͨ6���.W�)!�$|�#wN�t�>1�$�
!�ąGbX�a���:���D�A�!��$��r��� �dd!��ع�!�3A�D3ĭU�g�^�:��.�!�dG;Ҏ��1O�-P��L	2FU	
�!���4o�)7�S�yy �	 k�n[!���s�i@���JB̽�@
��a2!򄔯VO�sӨ
$s'�H�	�=gM!�� ��!Ȑ� n 0H�ǚ2�\ "OR��[�wEB���Ϗ
P��A�"Od`hS
�{OD��D�K� d �"O��ehД?)n�{G&H�N��"O���q�ʝK� ̢�<��s�"O6����Z�R��FD_N��u"O��Z�ā�d�xtH�
�N�S"O�=y���d�0�R�AI=����b"OlpP�.0�H�#fp؛�"O�]p������؈�E��_f(92"O�@S�0/,�zs��wep ��"O@�[��{+�ᴃ��n�����"O~�(T`A��L���8�NUh�"ON	ۑ+Oez��A�՜}��i7"O�mq(��6aV��@�4-��0s"O��R�KȐF7�� b��c���#"O���Qor2fq4�ACMP9I@"O^@�sC�U�B2��>fQ@P�"O�Q��;*� �Z6O� *J�p�#"O�8�$ą���زK�<v���"O���g��U����@ s6$�4"O\��§+5��4*%�R`9R�"O�9�f�!A�>�X���'��p3&"O�d(�(�,: ~�$]�N^Ԁ#�"O��r��J�_�d���e��iS�]�"OJ�"!��+ר �d��	rr���"O�r�M;9�t���C��#���D"Ojq#R���-|d���<���c�"O���V��8�d�3VBX�K��yc "O`���M��w��wA�PwH�K�"O�hz��ͯ���P �	�9Ӂ"O��c%B�C�	�#oN�BF�"OQ[֧ŸR���G� oTI�S"O���a���%��-M��̺W���y�̚�[��UK ��n^�y����yB����0�E�4iBl�ɓ��y��0�pt!@	���(���*ժ�yB�R�h�9&���.���4�yD�/���㌕� *���9�yB�[hq������Cc��y�jP ����a���]��@׃�y�FX9d�L�P��Ź}��${��H��y��!R�^աV+W(w� a[�Ť�y�n��l�T[6FE�%r��hu�:�yR Yj���RA�34	��&��ybC��e��ӥ'l�����yb��.���à��^	s��T/�y�(Z� E:yy�.����$��y"�T�1W�����I�X�3D� ��y�M�-�tђ�G�6�F����y�lU�0f��J� �)�9�����y2OD�,F��U $�S���yrD�b�e[��ׂ�tP2�l�/�y�+���3Ɵ4H,Ԕ�"�_��y�� ;M�R�����FXf�B�eÈ�y�$�	EPȤ�0�E��L�Q�C��y�G_���7N<hY�!���y⇝L�&��2J�iYj�"��T6�y��,(Ѷ�� �݆g�
u���$�y�AZqm��� H#6�$`a�m���y"�ުH�̜��J�* �d���dΟ�y"(V%x*E����szQ��˅�y�M],i$ꑹ�EDR��$l�-�y2� _F��q*,k���n]��y
� ���.�&Z��Ƞ�bYY�҂"O�����3)�Pq�#l��� "OLt�0��\ �X9��25_,ĉa"Op��tg�.�$���=N�|�1"O�;q�M�+�H��7쌹�"O$+��$�����#�#2D�R"O���Ǭ�e)�TV��S�}"O� ���KQj )���G d	8�"OD(�/�|�Kw��n�byJ%"O.��0
F�.�r�oQ�_���"O  P��!����a+B+�V"O�Ut�х�N��I�gΉK�"Oh�{�K�>2ς�b�"Y~��4"O�$�al�W��듍�F<��Ӑ"O�l��sZ����>/�jd��"O���L2f�()x�hR�g*$"�"O���h�A��i$
^�+٠Ec"Op �R��E����'<��U"OL�P���)�b�Zw��Z	a�"OHqc���a"�aQ�5]��"Ojx[�����va��J���]rS"O����@�R3Yt��� ��V"O"���X7O<D���A�c�Np� "O���%C hY�C��Zo((�"O
�GK��@0�%��4z�*C"O�ɐ�i�J�����&[�q�"O���dT�Y�$�W�>��8��"O�	[��q�Z@ފ�Q���_�!�d�=F�&�A�G����kɖ�>�!�ȿZ����Z�'�*q饂��/�!�B*�BLI)���b	[��F��!�$� e���^'T� �Qqh�;{1!�Ǎ�0Q����-`Ď��P��?I%!�d�0f$D����G%e^��JdJ�'$>!�^�TG��!H]�IM"�# oQ@C!��N���u�#_C6�����ѓt,!�$D�Z���Z�J��p�BW�[+!򄟇WHPp�iX�lp�{��@"�!��	m>��gႬbR2D��QV�!�S�#j�Tj�Y(O�!;'�Ce�!�DK9#K��Pm�<==����&�/�!�DA�$`���- +�nl��k�)�!�C�7ʴ`SE�����&�O$%!�أd�*�!�Ǎvr&ly$cÇYl!�D�""��83á�*g�%�U�P�`^!��#_V��0b(��S�
j�?D!�$I'M�*D`FǞ�X]�E�ɿ�!��_h���+\�sR��EfH�Q�!�dճA���"�d$�pEݝH�!��� 5jT)��R���A��=Q�!�dS)e��a�c�=p�L���9!�$�z��4{u���fX��6�L!T!�dU��6��P�	�?�X�*�GŐx
!��UޢmpD��H��@$̘?�!�d�&k.Ԥs�K~�cM\�Hg!�Ӂp�*}ӔfO�&�� ��o�!�ĉ=&��9� ��*�s�	�s!��Q~
�I��-P�	W�����L�!�D^����p�;X<��iuBW2o!�䍩[����w&�=[Ϥ-�!��d!��oalݫ`�S��H��*�D!��F)SI�)�#�OA�,Ʌ��0V�!�D٣3)N%�2�]�WD�i�!�d��O�xZw�	(?:���8n0!�� �y9�EQ9�|����zG��e"OP�!��NUu�a����v	�0T"O�̊F,/xw��P֥N�0Z�ؠ"O��C�f�lՂ���$� ��(u"Op��qBF�(@��$�,,�pX�#"O~Ѫ��X�s"��Yai����� �"OИ����>����Y�)?A��"Od� ���	*���pG�'J^�)4"O����!�sD�)C񣅃V8���"O�aA$K��:T.`��%�D= �S"OB��4�ޟnהD�A_�q�J��"O`��6M	TЁ�a��	U:�"O��z� Ӑ5b�2�*��V�0�"O"��&�'QtH�"	�>�Ν�"Oti(M�;>���`A��'|�4��"O���'k��r��W�1eh��G"O2E�0f��&�$�/�-R>@y�"O��!(X4� ��smӦ��@ T"Ov�9��)XN�[N��*��(#�"O~�Uj��7r���bf@�x�t"O �!T/�1f���sǮ18�@X�"O�����O<}�,h%-�<�Bř�"O�)hq/ϧ�H)��W`��\�d"O�!4h^�|u����C�(����"O�T#T"��A��i����8\i �1�"Or�q�&�;)?�u��`RM� ��"O�X���#}��l���J&M.!"G"O��Q�ቾ\�<�$�]X���"O�Lq�F?�|2s%�4j�\@�"O��8T	 TӶ�@�
�qo��t"O� S��::B�a��A0dY�D�7"O����K�^��QI�aLJ4	�V"OHU�Sy9�iRT ��>B~Ey�"O����C�Z�#��ەq1V��"O\X8"��&vn�0%m�("/�	�p"O�� �E��Z���-�=  ��1"O�P�QH,�TPJ��o���"'"OᘕI!��r�훑�4r"OP���mR�p�v	+q/ظJ���Q"O���
   ��   �  P  �  �  �)  [5  �@  #L  W  Ec  �n  az  ք  I�  z�  ��  ţ  �  b�  ��  �  U�  ��  -�  ��  �  W�  ��  �  f�  ��  	 �	 � � � u) �/ 7 �@ �G =N �T �Z  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8��H��I*Hă�%�it"L�B��AH<��	öZr��r��H+}J����Q�<ᕆ��8a�%HI�Vݚ�;#`�L�<�ǅG�a��P�����4S�h�O�<a���!=�Z;!)��䤒Wo�L�<I«��>Bp�Ā�L��%��T�<�􅌏i����䇺>؈�i6n�L�<1&0E@�9�7Q숨�����xR�[�wb��j\�g�T����)�yB��,�t��܀R�Lex��8YW!�dߟ}�6��-���H�HU�"OJu`�7��⦌�#7�d�c"OJ)� ��/e�:PYq�f�x0��	JX�x�(G�r�q�Cԧ?�Fp@$5D����*�:(�th
��e`)� Nh<�Bg�Np
Ղ�ݼ�;U��h���?!6�R?D��('��d�S�	�Z�<a5�K7�i U��i��U��n�k���OY�)�Ő`m��#@�YifD�b�'����i�J��8	��ʴL��ط�O�"~ΓT J!��57LTH��Q�ܜ��ȓK�p�0�A�/���qGH
ad̅�CS�`�(6`���C7��=�)���>E(�#Զ(�ͣ)�=(v�݅ȓc�����#O�`r��s@·IB ��e�����C�R5"|�d�G�Wlt��.r��Sk_�I�Q"�(��Ic� �ȓ]�~���D4&�p�q�ϧ� ���GS�-M�F���Ck�'$�r؆�)Rp���"Y�R�n����l v���;&eX�%ڪ}
}@�gd���.�ի�o�.Ŏb�Isb��/>��cu�7��DB� �#'O�x��9�{���;jh,j��å �vԅ�S�? �@�V!��\&����dN��Q�"O@Dځ�B�yn.��6�P<;�~���"O��"��Зw7j��IY�U�Xik��'��Ć�5Y&�#���,~V=*X�7e!�č �<�{���+j)�t*#\Q�P��cZT[ׇ 2f���*Sn��5�|B�I.] �X�2�V-���n�:s�fB�	�-���	/�n�����ٲD|�C�00 .�x�/��U����8l��'Zu V��/�n�zů��dH�rǓI9`��)��?1،,���,P�M�¿��B�	�@���c֍U�!9�E���C-]��pG{J?Q��OE�7���A�'�Z�X�[�*O�0���`��UM�-F�J�"O"��##
MD�yc�xT���"O��D�Z2��	84k?cc"��"OFI6l_!j<��rV�ÞN>VH;r"O-��D�%T@�
�(�:E� �Y"O�d�fh�#W.�)�V���
5��(�y�)�Y���і��*�8��K�l��ȓS��,P�(�?�����L��$Szp:%�im�\F~�cĈg��� ֋�1T�P�*炓���=y�|r��,G�yd�J#D�E�ƪ�5�yV/C�r�[ ��$=�����
�$�y�iC�d����#�14��`R�d��y�\� "�@͌0L����� �y��Bgz8�C��!m`����y�@��V؆��+l�H)��L�y�Nٖ?���S`-W �;��Z��y��"Er�rR-�InL�sQJ��y�ɽ~D>�)�JOS/&D`1I��y��= L��9�C
H�ح"�"�y2IɀgJ\RRXC���B#KW(�y����D� �aG�e��{�EW��yR@�B1UG@�V0���QN���yR��7P˺��p�I5NM��P�'�yR��%9���(�<F��xb@���y�%[b�!)A"�09R<u��m �y"�D�v/`���X *�䭩K���Py��4S�4��F�A6�b�'W�<9Ǘ y�1y�A_���sF��G�<Q�aG1`y��J�M�i��%�*_N�<�1�_�.�D9��+U	�~�gk�Q�<�w#m=Ԍ����1	:���#FW�<Q�E���Q�p������Tl�Q�<Q�j)����P�)/�~��!�K�<A��[a2�	��ȼZ��� ɗl�<�L�<q��U��W����`��<i��1 ��Sd�M,�޹xDG�{�<�� :'�`A��N�4D<�Q��}�<���ʠ5�z��ҥ�)?�0�Ey�<��$K�3��̘'4��4��N�q�<Q3�"f�x$(�-J(=�0��'�Yl�<!�]�$d �K�̖�~uCgBCe�<	�i�;���V ��.�֍j���g�<a�ʲm�JLAڿN_��9���n�<)f����s�K�q�gmQj�<��Ʉ�@��`B��E�ޕyC-�^�<I�$�yU>��֋�/#��A���d�<y�Ɇ�ER��R �ح;�6����]�<��6�<�Y��2h�}b�p�<�� I�a��W�b�|��Dm�<���$}L�%aGoU~x4�B�L�j�<�Cǯ>����@Iz�yr��f�<� ��B�!���"fe�="1��r�"O�][��ۚ_���˰�W�f$�Tc"O�Y��8N~�`�V�TD�`qD"O`t���/��=�ҫZ�z6J�1"O@�z@�!R�4�)�'�3��0���'T2�'e��'��'��'�r�'ZJY@䫋?��Q����}RȈ��'��'���'LB�'���'w�'��h��'��4�ؠ#mB� �'�B�'���'u��'���'6R�'��̪��
"%�9`��M㐩�$�'���'b�'��'�b�'YR�'z
�����"�����s�����'8��'eB�'^��'t���ٴ�?�'�D�*�6eء,4.��1�d@S3�?���?9���?����?i��?���?!"��m�C��ˊW�x��b[,�?i��?���?���?����?Y���?v�Vi? ����M�hRf "q�M��?	��?��?���?���?���?�U�CI�T��@	\X۲���?����?���?q���?���?��?�f��l����
PFJ�Ҿ�?����?q��?Q���?!���?���?���P�XI`L{-7s��@��bQ�����I��@����,�I�@������	 u`d��ԱcD����S�O+�Oz�D�O`���O.��O����O��D�Of��
��x��p�ÿ0�L�S'�O��$�O����O��D�O�d����	ğT2��S#AZҝ�r'%�:� ̐����O��S�g~BAsӲY��$d��#UJֿn�*Qh�"�b��I<�M����y��'�$�p�+;�d���K�U|(U ��'���[�q�撟�ϧ��D�~
Ł[�9h��8s�K� [��QCPz��?�)O�}z��7�v̸�l�p���`�޶n���K]��'��\lzީY�OZkm��y#�ƹ4'�x[�f�ʟ��I�<Y�O1���@Ӝ�>��Ac��;1�B����$f�	�<�'!�G{�O����2w�����	t, ���#�ybW��%���ݴH�H�<ATnx��h�ހzB����J���'��듷?i��y�^���U,���/ңi�����??Y���j!�#_^̧�h�_�?Iul;00{��Q���8(L4��Ĺ<1�S��y"�<(9z	�eɂH���0��8�y��q������H޴����TE	��%j`NԘAd&�p�E��y��'��'��7�i��I�|j�O9����H9['��3í�tm(6b�H�Ivy���y(E2I�z�1��щ*�@]RŅX���d��9 �n֟�����TE�9]9�D��&���X��^�mD����McF�i�PO1��� JEW<$�"KK`����j�� ��<9�eMm��Ă�����?<���;�-�D7�p
p"
�u�a|��uӒ�R#��O�pG㖔)���2CZKmt	��L�O�m��_R����M��i�6��0>)�$��؂43\��aE�hZ�$	�Bx��z#xm�5L�.8xL~
�;<�n!Q1l֢v�-hbܔ���̓��?�֏�#�v�[��D=L�D�P �_��?i��?iF�iʨAbɟ!n�r��7FMؠ��:��R�M�Np'���	��S�.e�)m�A~Zw#�� F#c�)KaI�������៹<�d0�D�<����U� ���^_����@�P�Ol�n#5K�O���O�˧ �X�  �
 �6QC�J�LЙ�'���?	����S����/;��}��н)sȀugV�p).D��H�e=�fm�<ͧFD���\�TБ�<{S`�T"I�lu��ɟ����@�)�Sny��bӸM��/�|�k�T E�$QG���M�&���O�QlU��U�	���Q�n�?kS��BA�V�Р�Fş��I�~�l�r~��ڀo��T��A�I�g��Jc�F�.]̌�WA�3I8�$�<9���?���?���?�,����#3{^�K@f�����$!�U[r�K⟼�����%?��I��Mϻ4�,D���ۋk�B�Y#�5m��Ks�'^�FM2���4��{���7OpP!�&�0=pĈ�ņX���BD?O��G�8�?��J3���<����?���ҹR�Nq�u��(������ȯ�?���?�������i��`
Xy��'P
��!�p�X�a3��>e��(Qe�DWX}�kw�D�l0�ē�j={2�^0NX���G��"H�P�'��|��ɂ d/�@����d��T�D�'��ڧ��}�
@*
)�li{7�'���'�2�'��>	��*jLJ�M�#�2i�dAt���ɵ�MS`��$]�A�?ͻ�bQRAщ'Q���e?lRd�����O�6��-�b6�8?9�e?j~���;�J]��n~K��s);w 0�I>i.O|���O��$�O��D�O0@��R-{�4|Z�J$wj}Z�m�<AҺi�����'��'�O�i�iVL+ K�9o�Ppi��C*7�T���&��O<O1����Q*��32x��d��0�"�Є��1Μy��/�<��]�0���>����с
��QOý@�f܈��	�����O���Of�4�*����X�Rlʭq �d�e%��K�XM�Ӡ҂B��DiӠ�,تO��nZ�?�ڴ(� 3b�]�w<L��P���ABl�.�Mc�O��S&���ʗ�4�I��� ~h� ��7�,��U�����36O���$�#c��)@��|���:0�${����O����a���>bV�i��'!�c�+��bq��Rgn�:?��0�0��O�6=��X��}����شR��3��;��M�I���ʧ���0�䓄��O���O.��H7>�p��*c(�D)�&Ry����O�˓i����F����'BX>��2'�T�4�L�X�	��+?q�P���IП�$��W������K������aE�X�pMpش96�d��ug�Ϯ~���/}Zc� �7l�+x,�i�ᔼ_�Da��'�"�'��O�I1�M�N�8�~ty��t��t�`Ak�JU���?��i��O�!�'����-�J�wȅ�/�Z�J�J�y�'O�z��i,�iݱ���W*/O:�.I�
����偋m��q��?O���?���?����?�������|8�臋&Zl	��Q�'�|�l� $��'����T�'͈7=�t��g̋e
�����&?���R7*�O��$+��	��*�7�d���a�-}�:�����N���
t���g�*I{��.���<���?���̀!@'��~ȩe��?����?�����$���E�%ϟ��Iӟ8�0�	�UR��:�E�Q��t`��q�/}�	ȟ���t�I+CZ���.M9}�
ٸ׍%[m`�s���2c��2֦Fy�����OZ0���y4D
� �,A������O\�$�O���O,�}R�'����7�É� ��U�U��;�Va��A z�r�'z7�5�i����޵QBp"�,W=�lP��%������I��4"���Bܴ���
i7I���}�:Q(��,k"�G�Ʀ6$�����:��<����?A��?q��?�t@],�Т��N�7�������Ĝ¦�pr�`����̟�&?�	�W��۶MK 5ź�9��_��|��OB�d�O��O1�F���T/hH��b�V�2Ӻd���
�$7M3?��N?%m&�II��Ry��w�Б�bU,b��ɺW*�Iş�����Hy��xӤ���:ON�{%W9n�'�_���v:O��l�o�X!�	ϟ�	럸C�#�����\,��5���O�rG�l~~� 
?��D���w�Tɡŏ�=l� gy��p��'��'�"�'�\�b>-c!E�Uz̛'Ü.��U+j�h�����p۴ �A�'��7�&�d�"Ip.<cHΒ0C�����5JВO����O�iD�G��6�8?��(�����=;�Qa��_�$�x�c!���%�̕���'U��'Њ!*�A�mp1%R6��7��O��$�<a��y��#�'���'��F��1{2B�� �<`G@�$2��	��M���'L����Ԉf�BP3-�|��M�b�Ff.@���.�vi`��<ͧ*a�����O�Zq� �5\@���+D�d����?)��?��S�'��Y�А�?qܴE�Tj�3]�.�P1k8,����ԟZݴ��'�t� \�F�E
v�`�������	B"6m	�®���a�,,b����t��Z7�y��g��@{d�F���s5A�rd�O�1�'�r�'��'72�'��ӈTV�"����1�DO��@���4Q �P��?���䧺?Q���y�L�%/����D�A��L+��ѝʜ��OJ�O�t�O'��L-T�f:O&�kqF��S����TFX|J;Oȩ�:�?�e�,�D�<!���?AajV8:����͕"�� ����?����?���@�����J؟x��ǟX!� 7�|lq�	�����Q'�ԟ$��a�OB�d�O�Ox�Q-�*a��A;�dZ�y�IB7O��$�+Mz����G�!����?�
W�'I���	%%��eq�L�Hd��i�����Iٟ��I��X�	j�O�"� M����������BЊ�Z-�OmӸ1�� �OX�D����?ͻZ�J�k%���j�eY���Γ�?Y���?��ٯ�MK�O�hٔ)�)�z��%� ̻�e��ظ�T�0�L�O���|����?Y��?�\�C�օ_�X\�E�!�+,Oځoڻb� �������n������eqf1PѠ�"ZI�r�ث����O��/��)��@0Uʒ(C��ȓQ�M�5�qriV �ɛT;0Y�b�'�@\&�H�'^�A#�]?pBf�Y#�SuU�ȣ��'��'�b���_��b�4q:�;�L�
�d.5wv�ea�2Gp��ϓl����D�y}r�'��'x�z��C�$.x�` @�*�P�k���/;z�Ɯ� CQ��^���&�i��@�x@Jbeڔ*�� �T9kP>O6���O��$�O���O^�?q�!fej�j����A�V����� �	�P�ݴ)�bϧ�?�ǹi�'��|�A�
��`dխC���%�|�'��O�0�{��ii�i���'Л[I� ���g�8�RB �Pr ������$�O����O��dP#m9�*S��=[S.�2-9��d�Oʓ��K[-��'��W>UQp.H�%��c��� ���Y�n&?��W���I��8$��'4*n��rHW5r��PD_�yPНX�"K�z �L3�4 ^�i>���O.�Ob�j��&m�v�S��O
cL�e1d��O\���OB�d�O1��ʓq����7x @�p)K�p�D(�ߢa��ŊG�'��j�J�h�O"��½C#)��B,]6��+3���f�*�$�OvtR�r��Ӻ���,���T�� Z�0�I�	~�.�[a#K�W����;O��?���?���?���	�8P����D�A1'(�p`3e�T@o�w� �	ڟX��_��ڟ`�����aL�	�,)i���[j�I�"� .j$�6�rӞ-'�b>ik��Ʀ��=�[a&<��H�R�KA4�Γf���m�O2��N>�)O���OI��ݓu�8�3s
A�k�0����O���O �$�<!շi,hp0E�'���'�Zl��C�{\`z���:=1�]��D�u}��cӶ�l�>�ē����.�H P���z vm�'F�
P�#� ��֗�4������f�'*f�{��R?6��lYp&�,�P�3�'���'L2�'�>��I��Z��`X2})Rk&(=F�� ���M��c
��?��'8��4���g^qz���2(W�q���a��O�6m�٦�4$B4�Qܴ�yR�'������?��c�Ą5D!I�������L�r��M>�*Ox�d�O|�d�Oj���O2|�P��\�(e	���$=ʰ ��<1��i>����'4��'��O5�A&R����=�r��!*_�`��Hg�<,$���?��S�\��iB�����#��Ǫ�tؖ���&�TՔ'�����ğPR�|�S�`�gH	�>l�;K�i�J�hec�Ο��	����I͟�SIyb|�R)p�<O��)*K6.�˓`G�N�h<O��ne� ���某�	���b�"��q�=r��^=Rk@�pB�?=@�m�<y��`���f%��'��4�w7�f���+D*�*o��q�Ξ*�y�'���'��'�2�I��q�z�is�:0�화NH�FO��$�O��$PҦ�*��i>����MSL>A3 �^��gY^�$�SBS���?���|���G1�MC�O�Ha�������K�/	��3���@LzX���]���Ov�S��<��I]D�8�BH=bZ��)��Xs�'ג7�ȁM ���O���|"'�,b�Pi��,O�?@|D1q Uv~bE�<!���M;ƚ|*�.%��1o����TƈB>�HCR�)`فW��O���|�t��O4�;J>i�.Q�"7��Z�
�
:^�І�s<�Ľi�H��4��2���ce�\���l�&D�/I��'|�7;�ɏ��DȦ���
�
u.�m�~�̰�'���M�r�i�G�i��	�,t��O���'��sd�N�H���S�ʉ�2� ��'��k��|*g��i>RU���	45#�U�c�R��M�S���?���?ь�dMl��.��d��DH�H�F/κ|���l��Mr�x��$�~�&1O��Ec�3�,����x`�5O8LP����?a��.�D�<�+OT�YS��Iք�I5��u��(Xf�'�6M=x�d�OF�D�2`d�P�&X5������n�l�O��lZ��M�כx2m��^q�{����f?�ً�[����U1#�`��*6b�2��V�(��`Ȥ���2wހ)�l_�^�H48��1"O!�DŅߒ��C�ڶ_�ua��C�o7N�����P���|�I�Mۈ�w��t E�p��H���2��,��'�V6����mx�4U�iٴ����+!7u	�'%���+0&L&w�tMHv-�8�Z}�!�D�<I��?����?	��?]�Y?
��D�_�j������iu�����	�D&?��ɅP�+�I��9r�- ^�L`�D�>	B�i���$���*۪I�ȗ}F´ �G�=Њ�hDC�G��rZA�6b�O4�M>�.O�]�V�J�xnJ�9��A�v%'%�O����O���O�<�$�i��R�'���Q�G�4=N6�X��ĻQ�p���'4�6-)������7��Xo�7g�.yh�JG��T�Ю
������ӦU�'�*���?��Ґ���w��S��!�.E{)��p���c�'���'���'���'��~ps� ǜq�`M��@�Z�d��d�Oz�d�OҴm��"q���'�7-�D�?�`i��U�^t�B�	)H4M$�hB�4?�'4���ߴ����G��	����-�*�8A"�=#�δwސ�?yB�+�d�<���?a��?��/[�\�d񠬅�a�v4��/�3�?������ᵋ���	�\�O�
<CVCZr�"��B�ʏgV8j�OL�'�^6�O��D'��'A��rƦ�3���U�[�K]��!d�V! ~ă����4�����Anz�O�r �Vl{�!��I���(�O8���O���O1��˓X���ɡJtm�D	O.h��H�J^���P�)�4��'h�_�v����\YK��]>~L���D�;���u�L�� �eӠ�U�L$0�n�HU1(O*��U�ۏ?	�!��P?�M��5O�˓�?Y��?9���?�����)��b�h��H*@�F�3'�5<��oZ
�P�	���`�S�0;����"����k�	٬ ��E_d����?IJ>�|�U��M�'LB��n=~�rȢW�[�\Ѡ�'�&���ퟬA�|�^��S՟ ��Pt�:0@ń[���Ή�P��П��IsybD�Op=��^��I�++��*��G/y²���S>O�l��?��X�$�Iǟ'�|��\|�Ex�	6�:E���r��I�W�`����i� ��%��O�A�w[�xq�环IP>�C�@�-����?I���?���h�|��@y>�����w�H����7��dYצ}�e����I�Mk��w߄� �E�<�*�F�7!��P��'��'[�`��>O���:GBT}���d� 8�ڕ�Ґ
�ДC#F�	-(U��3�$�<ͧ�?I���?���?�7���=�
���9=��M��%���$�æ)ÔH����	ܟ�$?�I�x�2�c�M���qP�*^�� �O�$l�?�M<�|�co�P�t�Rl�5 ���ڐ/�[�.M��ȅ���C�`oV�
����OP�(�H��j�������H�3j�i��?1���?���|�.O2�nZ +��P�	�Y,�%I�
%�0��U��X�|��I��M�"�>Qջi�d�v�\���O$t9��`2�I;��1��9@6�7?ipǂX����_���ֿK���;V�8C�	|��X���<���?����?Y���?Q���ĝ�E�R��o���p��%�1ZMb�'��Oo�~�!U�?��4����c�/�$>Ъ-�-A��[Q�xR�z�D���D�bvb�b��j���U�bR2� ͖�Z�>��E̴�v��q�'��'H��'���'L���hЀ(٢��E��w5���'��Y���ݴ��Y����?y���#K��b�
 w���Ϝ���	���d�O�D&�T>�p�O
M�J8i`�[8.>�bR�W���0ԃ�¶����D�ʟXۂ�|�OC�Ve���ʘ+�fD��n�"��'���'����Y��BٴdIn��5Ex,v��'`��it
pȑ�I��?���e���|�O��,�����N��H�i��M7H ��ϝI�6�ݦ��F��'��B���?9 Z���vh�T�c��c�zz��`�T�'}2�'gr�'���'���L�j��Ş�y? ��&?J���Z�4_��݃)O��d<���O�nz�q���	L[��X`H�)���M;��i3O1���q��|�*��?��e���]��ՠS�#YN�7���E�'�'��'���'j��S
���h��U�l8�!�'6��'��[��۴7���j/O��$3�JKD&��*{�0�R	�`&�O����I}R�x�rdl�ē�Ĺ� &�-t��A��a@���',�ԩ��P�nn��q����@���q!�'�����dE��r$D��7���0�'��'2�'��>��5SF��&�I<k�qC�v�e�ɟ�M+�O]��?�2z���|��y�.]�9E��"/��
6��j���yR�x�$amZ��MFc�*�M��OdB�c���6'4aX=3�ɥ@I���#޴�O�˓�?q���?���?���"���P`� j� gA��rmh��(O��l %N��'B����'T���#�� C��9�kZ�u�XZ��>���?H>�|���
�F��Qd��C|` ��ӹ���:�4p���9=�΅���O�O@�pL�
���v��8 B��*�T����?I���?���|�.O
l(����"b��`z��.�>1�G̻D���4�M���>a���?��;OD��Wh�=0���c��9
�,�9�M��O�'���(����F*/P^�'�B:0�v5)���=����O���O��d�Or�D&�SLb��b`���&����O#�V�I�L��<�MK�j~��b��Oٓ�H�p=:uKP�sg���*0�D�O��4�,�c*{�d�D�hd G��A�� :�Ń54�����#au���A��py�Opb�'���M�&Z�"�d�*^p�u�M6<"�'o�I��M��<i���?�)�
���ź<�ft��B�w�U�'���a�O���ON�O�P�H�C�˙M6��U�Ó;:D� �g��w"l�G~�O�ܑ����ic��Լy��t�%J^q�]����?Y��?��Ş����ɦ]ha���5��AUw����C��En��'�����{}��'��H�ch��&HP�.ӑ%��3�'���!O��期8���� 	q�<��6CL�u��ͰwJk:��cG<O�ʓ�?����?���?��������D�O$��ѻ�� ��m��J��I��0��h�������c�EA 2����3�I�H��tȱ@_�?!����ŞV�����t��5�̶H�n��A��!R\�w��<��.e���o�IMy��'��F��<|�q�E<X17�n���'?r�'��	:�M���͢�?Q��?���Լvs� �C�,��&Z/��'���w�V	�O*O�� ��U�����I3v��=���<� H�aVpyb��f�S�b@"������7"U.w�����)Ǒ?|��v��ǟ0��ן�����LD�D�'f���B&Wݸ5��M�u�L���'17�3'����OJxo�M�ӼkA���;��q+��EE=KC'��<i���?y��T�[�4���Qi���a�'�q��MW�oN��C�nG:
!��K��1�$�<�'�?���?����?���� nS"�\�ٔO���D���QC��O�,��Ο�%?)���/�t�`�����8�:��Mrh�r�O���O�O1�TX�D�`�l�qQ �;q �{�b�	6��[֕�:��E�d��M��_y�H��=ٖ�3��n�v})R� ��	�����ȟ�Szy�+q�丘�O^�Bv��IR�SƬ�Gc��9���O4mlZi��l
�I��������%1w��y����Dgxً�l���n�R~B/^��.U��cܧ޿%��=�(hr����H�-D̓�?y���?)���?����O�b��5ɝ�'˂AÑ��3����4�'�r�'MX7->����OAo�R�ɷT�M�%��(F<H�P��0~lm'�H����x��+RA��l��<��n�d� ��H����nX���[:�@Pf��?0�&��<ͧ�?����?)�*��QV^� ��ρS��`�t��)�?����dY���H������	�@�O,�!+���]����ɝ8${��
�O^)�'��6�]�$��'.v|UCA�?��Y2�ݏ{0��b�I5vl����ޤ��4��I��q���ObqQ��4#$�0��=j�jr@	�O��D�O&��O1��˓qn���>�R��A�K;Ix�P��cē,L� �C�'�o�j��I�O��m"@�4������H�@�0�R���M۴IK�M{�OJ��p�׃��N�<���M�T�)��<��U�aF��<�,O���OB���O8���O��'!�����B)~w�!�ӏZ�F^��иi.�!��'pb�'K�Os�Lc������6-����b�*Ԕx;��oڑ�?iJ<�|R��>�M�'48R��S�=.�S����whɞ'�>E�#J����|S����ğ�K3��+=VN0˓�q	ۥ[��?���?�����$Ҧ�C�l���H�I󟼉&ĩbd@&�*h�n1��ʖY��g��ٟ��k�I0ܘx���C�wU�%ӂe�+���5�V��tE�^�']����?1��V�R�$���4C]JmJo���?a��?y��?y��I�O���
R-��"rL�g�i��O�nڙTG�a�I�l��4���y�L�(p#B��@�2��-q5H�y2�'���'dB @�ie��#t\]ZS�O���!��R `�hՃɳ �<��O]�Isy�O]2�'�2�'ir(�_��93J\l5�d
>]��I<�M�pʉ&�?a���?!M~j��Mޖ�A�$�p�8��wG�����\����ߟ�$�b>myg�	]��(e���K���w'݊j�P��qE,?�#�D�԰�����䓟�$�,,��H7/Q�O,�� hQ�:�*���O@�D�OD�4���,��&�W�B�I*:9�\(��޽E���𭚀%b'l�,�Ԁ�OJ���OB��Ψ�ԉ�D斬ԍZ���o���;Js���;C
#��:�>��]�>�Ha�Sϒ$;�n��p��/r��I֟�����	֟���i�'=���!!sN��*����?Q�aț���!��t�'�6��O�ʓX�v岤O1NL��+0��"$}�M>)���?���X��k�4�yR�'�ح˅dF	j���7χ}�0�aт�(&Zdp��/��'\�i>%�I͟����TlR�)֘te��b�K�h��h������'i�7ͅ(+ �D�Ov��|:E��'e������8"(Dm��D~�>�i7-n�)��t��gO���� *V'�=��� ���F��M�+O���?6'��E�mkG��d�33`���D�O��O��<���i��U��K
܄�DU����Yt앞	�剂�M���D�>9��z���E/]��RUC�e�'.������?a�ͫ�M��O��P�V�Ey�d���Z<��9����d���yr^���	����I��I���O��;Ї�A������$=���w��-�"��O0�$�OX���d����]�i*���7��:k+$�;3C� ���ڟ�'����P���CE:�l�<��R,R�Jڱ�£ ��`��<9ulɡ
(�IU�	MyB�'��Y�(�v�bШ��Q�ΉȀ "]�'���'Z�ɴ�M{Q��(���OP$8'��'T��P�I��Uj`0rB$�$�O$�'��i O�dQ�.�'OxX�b�8:!2Q�����R!ĄV�Ġ��AD�S�\ρ֟h+��-A��b�,�k��QJ��[�����@��쟸G��wF��P�ǉb���#��s�8���'D6MU}p�I��M;��w�˷���9801!B���f�d��'���'�B�^�$��Ɨ�p#�� _�	�@�2���_(�(�q@j��g�b�O*��|���?���?��޴��4��nb>-#��=Y8iK(OAm�%6���ßh�	v�s�$b`&]7(��ElU�o���*����$�O���7����*H�JaR��\��W�ȁ�ZP��Lz���#��{Pͦ��&�8�'��A��(�hZhx�A�Â}�ܼ�E�'���'=b���$Z��y�4q����r�����W�2���5�8h�F��K�6���F}��'��'u|c�)�=k �����),��!��^�柟������Q>��ݎy���ԡ�'FRD(xcD�7mH�	����Ο���@��k��x�(����O�dXe��g)����?��W�������Jݦ�&����FM�~�X[�dK�hIq���z�I�� ����,+�g��y��?wG�{������!f \qVkE(q6����I��%�T�����'��'9�0�#-;.v^1#Ν2D���0�'��U�4�ڴmw�!���?i���)��l�X��Ǒ*��闧$��	����O���!��?���߯[b|pE��D��L{�nG���5"�NLW^ ��|�TN�O� �N>QA'���Q����q����ބ�?)���?���?�|b.O��m�^��i�VL�o{&�Z���t�(�bLƟ���8�M��j�>���34��sQ#�-g�p۳�_���`8��?�*�M��OP�1ŉ���O?�B`��vzN�ra�Z2
K0�R�@��'�b�'�2�'�"�'�員
���a��!f�2U+\�7��Q;����'R��t�'B�6=�~�'��4�p'��;e�J7��O�d.���9<7�j�� �u�GjE�9�j@���^a�<�f;OR4�kD��?�F/�$�<ͧ�?�E��n\�C�h�R�!�(�?��?�����$����!
����	ü� _�~p%)�d�n 0���H�@��p#�IƟ$��E�;m�ڜځ���+(� -�Wil�W�P �@�����|����O��x���j5b�kR%�>1��!tN9����?	���?��h���#a�\	�`Ν_iʜ�և��5f��������ٟ��	��M��w ���O2t]�I3�Q�k�JM��']��'�B�/	m�V���{���7R�� 5d�n�pFb��D�lsDD��T'�d�����'"�'@��'jn��Nʤ.��]�G�4h�a0S��c�4MZ�E3���?i���'�?��j�=��h�G��%� u����	��Iݟ��L�)擷)�(�K�����XC�G֡5>���M�!��B!�|�Qe�OV�N>�)O��5/M��H�0�]t*H�pf��O����O����O�i�<�4�i���:��'������o,0a$�N;H���'��6M!��0��D�O���O8�iI��zt���&;�PH��ЙS¸7� ?�B�ľI���S]���ѣd"�y(�[V(_Eqvpr�hw���I�� ���4�������"D�|Ů@`�Ǔ14y����?����?�a�ib\���O��
x�b�O|D��2]�ph2�Ҥ)�U�s�'���Ot�4��bF�uӶ�Ӻs��ǽ��c#M=h�
�ZJ��n��' �'3�Iȟ��	�8�� ܮ}�f�Si�h�X�iG+p����؟@�'�6�ɗY�����Of��|�7摠]��P$n)n�.�r�o~�l�>���?�M>�O�)gI���@G^?�>�P�N�"2&�Ұ�im���|�!i���&�X{�JT}��!,ߛ2Z�p���1���4B���㟁D{]X��A�&]#rOD��?Q��Pk�V�D�^}B�'E~u�G�8�|aA��'��YhU�'"�"�����֝�7�t�'���R�ɱ׃�wqq��:Q��ı<a��?Q���?I���?�*�$%��k�څ�``�X�Eڨz���l�"!�����ݟx��e�ݟD����c��Y";��+TΚD��DY�@T�?�����ŞT�dA�4�yR��!<`x����)SH=��Y�y ��y����IxX�'��i>������a���F��C�%^�h7���Iܟ�����,�'#�6-�b�����OT�$+w�"�Ѣ�ԍV�����0:����O�m��M��|ҋ�	F�<�0L�T��qȔo~Ba�6�v�v�P�;�O�~<���p��z���W�U6N��ۄ�&���'��'"����Tk__yr!��^�c+ր�,S
2��bq���e��O�������?�;?Xt��,b�H�R���1IJh�_˛Fj|Ӯ\mZ�9P�lnv~�J�/@���ӈ.��{�ݥm>�3���`�@��|�Y�4�I����⟤�I��0`U9�^ض�
�p}|�B sy"%}�؍8���O���O����$�$~`j�"ݙ+B�9��#��'��6�DѦ��I<�|�u�КT,,�3/��Cx���j���e{�"���(}/.���K<�O&ʓki�2�ܪ^�Nu�5
�?�%��?	��?��|�+O�Enڞ^�M�	,)a���d |`z0�a3}zh�(�M��>a��?��%���8�⒳I����`l@�]$��ě�M[�Opm�c����������w3�e�E
M�AaPKɊ!-�L{�'�r�'���'.B�'�������4e��5�K+U#ޑq3��O���O|nچ������ܴ��V�Xp��O.I;�̣�7v�rM>���?ͧd|���4�����X��r��L{�"H�K��pPp��R��'��'�����Iş`����獓8������	v�H�r� �O6���<���i�H�r��'C��',哤SjU%�(Q�h �W��[�R�p��	ßH��U�)���ץ��lZtO׎h}�&�J-X{�]c�װ�M�W�據[��&��_-#�0Z���n�:@�r-D�����O���OZ��i�<y��i���� ���>��	}Hܺ�&©��m����?�¶i��O6��'��7M'dI���G�Y���� �,6dyn�"�M��(2�M{�OA������`�<AUO8p��Ap T*ƀ��wA�</O����O0���O|�d�O��']5܀3s�E�m �c��4`�\@w�i~H8� t��'��Ow2�z��N�kp)��H����"�!\��`o��?QJ<�|j�	֘�M�'NIh3g�4(�b��$͊�2�o��<��H�B���Dā������Ol�$�*e����EQ�.!��b�O��R����Ov��O����������'��}�4��q�ưS�H�@�c0�O�U�'27�J͟0$��0�̤B��yS7c݅ "��Pa(?��nغRw�-["!����'\q����1�?I�"��_�����4�MH3L���?i���?����?ٍ�	�O��"Ag#w��[�˄�}0��ĉ�OD�n$^�~���某ݴ���yWD@p=$�ْ�XB��
����y�)r�rp��Ѧ��-���'D� 	PD��?%�LĬ+P$@�dV=�"q7+��'��	�H��ԟ8��ʟ��ɬ<��l�� R����V��"��'P,7mڅF��D�O �$ �9O�)&��=�օcQn�\��e����f}�L|�v���F�)��n� h���	8i� 9��چ=�:��jW�u�˓i]���O�iL>(O\�cw�O���RPfRd�2��Z�?���?Q���?�'�������SC��R��#�@�$v���ɕN�����4��'%��v��O�6mC�_j,�Kt��.t�Q��B�#M�Xc��`���	�n5)p&��:�1K~��� �"�ч&"�`Y���Yx�̓�?���?Q��?����O�\�ԌŸZ�ƙA`�M@���?Q���?q�i�d���\�<��4��n�L���D(�ЛԃL&fA*<�F�x2�g���"	S�mq���mpM���'��B�擎(zH��!/P�(f��]������O��$�Oh�dM� �`�#�_N�	�([�V����O�ʓE?��b!��'r��'���L���7"�KD�(��޾)���.����!�����S�tF�z=�|y����b��ݹ���[adL�gn�g����^��Ӿ"L�h�	�*�������&|x;L�H�T��	����	��<�)�zy��l�~�O�4L���	Z��%iE�y�|�5���dI}��gӰ�q���c��x�vϏ�.bD)҅ߟ�l�!���o�y~����t0)�S1��I�$u�(�̣Ux�Z��H$�v�IAyb�'�R�':r�'��Z>�!��<)�۱�	N:Uȑ�eU�M�U�]��?Y���?K~R��s���w{P��A[�h�vM�͓�d躱�'�"�|���JF�/�&;OD)�p.�?gd��9uW�w6�i0 3O��E�Jl;����$�9F��!s��fz4`���ER��9#�$��D����X͉Elג>1d�!�O�w��h�؇n���HP�ٯ'~��4�&�-H�kڈ
Y��ڢ�D�[�p���	: �"�PG͢M=>x�@b�X?1IH�8oq�a���@yG߄e��h3'��  �];fIjկ�;���҂��):*��q╣\�"�2-�6��L�c$7#S��V��%+�:=���36R� S�瞵p��<�� <f@*�P�&I�)��kd�ɴ1��b�=v�8�	­z�j��pf�Su����4�?���Tf�@�+>�jIa����4�iI�|R�'Hn��5qO̽��*��fW��9����.��X1�i�R�'�剿t�\ly������O��i�vZ���6�2)����go5A1��%�$���Hs�m�r�����¨i�>1Xv	R�s���ҫ� �M-OZ��V&�զ!���4�I�?%��Ok�2�lii����ٷ$�=j�V�'����+��OD�>A��eE>f��U��b��i1�iӄ�Ռ�����I�8���?q¯O˓5+��If�G970�y(%*Pvq**G�i�ZX��D9�S�����ԏP��| �E�?J��-����M����?���rnѠ�R�x�'�r�O*��I�{`r�*�)�z��@p��	�(�Oj���OR�d��6�L�1�N%}��`����/!�-mZßx�$�_�����<�����K��~4������kF*U{�,K}b�[,M�'d��'PBY�����@X` �5��=�����EH���O�ʓ�?�L>��?⭗g��M5H�0��pS��ӓM�fqyN>����?����D@bN� ΧP3�=�u¹D�Nȱ�����mZ}yb�'��'r�'�`��'�����H������ {P��t`�>���?����d���2��O��ybP�L#;k�ےdA�\��6��O��O&���O�o�[�%�Lh7,�% ��@�U'��6�oΟ@�	Ry2�� �'�?����Z2a�4��qjWm]�)M��Q�ָ3�'R��'�0����?�г�� �� ��'� ��%� -v�4ʓrG��ÿi���'���O�����@�L�?Hֵ�Qꂳ����`Rݦ�����
��y���O�r�(����_#ԩZ#�ڕ1�3۴S�b�Ļi�2�'���OH~����A)QpJ�5>_z��'T�
�Dum�%3]���R�I�'�?��J�=��r�'9���yeO 5���'j2�'笌 �Ϧ>y+O��仟h���V�
| ���eo@y�,%���)�j%'�����\�	;oj0j���Kx��R������s�4�?���Ϟ/i�����'\�'���J�%}*��P�
B��Q�v �d�O�˓�?���?�.O��)��W&6�z�)���}htKt�ŧqJ�h&�,��۟T%�(��u� l��`�T#^$��h˱I���Mc�����O`���Od�#:-�#>�`q�W��*YS���Di�#W�h����$�l�����'�J��Ό�dϺ�2���rԔ��.�D�O�˓�?�POܱ��	�OҙI���;z��C�P�Zw���)Xۦ��?��?� lY�<*� &���aNʗg��W�Y�1}�2Bj�H���OH�mH��p���'b�\c!��sc�ؼi	�n?Cv`��2�xrZ�l�7���`'?Q�'l|���/t�fq�E[y�*l�'m��^-���'$b�'��D_��]c���� P���a�r�G T�6��O���"xP�s��i�|U@Ȩu��F�<p	$c���_��r�'���'���X��|U:�3π��D�fR3k*r��6�ik ��g =������dƼY-D� D����	*�"(`�e�<�d�OR���mn�$���ß���ȹqkO�l�ܘ�{]"ElZ��'��H�+�~��?����?)��R=O��
rm�/�S�j�����'��Uc�#�4�p���O�˓O���ED�|�a�V?�:�2�i�"�L%8RR����'Q���b��xF-X�u\�-	Rf��P�d#�\���۟P�?y���?92� ���Q,�A��H"��,����%@�f:|��'��'�"X���� �>�����K�4���/�� �c�X�����O\�d�<Q���d�����Č%<펵����F(�$yaj�E�-�'~��'E�_�Ҳ(�&�ħa�޸CUD��;d&�0�C�1Y" )D�i�R�'�	០����:���t�i��W�T�"��N*�8�$��OC���'��Y���Rf��ħ�?���ۓe�:�hI)E.��!J� ���q�	Ny�'B�,����dП�Ш��Լ�q)W���jyS�[�@�I��*���ɟ<��Ɵ���HyZw�~]8�m_�e�űT�ݢ,?����4�?A��0��c
�N�S�'x6�U"����M檙����&C�vn�]��I�0�I͟ �Yyʟ�U���Y�r��&愐FQ�����ۦ�����i :c�"|"��U��3e�=n����V���K�i�R�'�r�C2p��O���O�I�d�ԍ j=CH\��OH�3NP7�OB˓~� �Z?�Пl�I͟PS�W�I��h���[
��l���M��1,�xv�x�O""�|Zw�6@ 0�Z\��� ��<^X�ӫO�h�b�O�˓�?����?.O�iXՀ�'@9&��b�Y�r\U�V(u&���I��X��dy��'�2o�>n�
9VCD�2����g��6q$�`6�'��͟��IiyR�'��	Wҟ�՛#�� 1���%Ґ}P&X��iiB�'��O���O�{���
���O�-.��q�F�.���11ML��D�O�D�O�ʓqb,q�U?��	�-��E���r0��	���1��)ش�?)+O2���OD���&tp��|�2���w��
� ��� ��l|H���'�bP�d!f�����O��$����bB�;^� �)�.�l'N]��K�L}�'�b�'��h��'��'1��
V*��̓u��:�__���_�(���#�Mc���?	���[��ݤ��	X��'Fx
�	����O��6��O����?-���Oh˓��O.*!�po �'kL�׋�.���۴4Z4	Xôi���'m�O�������B����铔�r���$��m��<���d!����`��

ĈIT��5ɤ���@&�M����?���[g�SY���'�"�O�z牘�WԊ5��cB���!2�i��'|�\������O����O�y��3(k������J$��Ǧ��� 1�� ©Ol��?�,On���b�a��Y0�!R��j��NP,��3�8�I矈��Ɵ���R��'��$�Ǆ�(ک)���,Y���`փ�}��ꓛ��ON��?y���?���]D�:c P:�8`��P,Z+��ϓ���O���O��:%���2��Z1Ӓc��I�T�
�:U�E�i#����'"b�'���%���&$�������(i��9��c�1���'�b�'2V� �G���i�Ok>tJVt 1 ,!�̱��Z�y՛��'3������	�(�p)|��	|?)�n� A� A E]�
�f{�O��!��러�'�!j7�~��?���u���(�n#��xW�2`�L-˰Z�t��������(��w��'�i�=?�y+EA�0,̱���	3j���W� ��Ű�MS���?!����V�֝�;~�HbSGl%���I,%�tс۴�?���r�HD��?���?���d�p��p!�g:�8"�k���MS�*Zs'���'���'2�䁤>q,O��Cc�������0� $��"Ӻ)W�6��y��|��)�O^�4JQp'��X����nx�E�Ӧ-����x�ɑE��hk�O���?I�'_��RE�F�e!L�Rˏ�&�@��4��D�O���$1O�����	ߟ�R�"�F�8�b�ږ2lԋ���Ms��$�xX%R�<�'([�8�i�A�F��%`��4��HB�p7 ~Ӽ�d�)<���O���O&�d�O
�Z���w�֍�*����h�䉡`�����FyR�'�Ɵ@�	ݟ�#�R�7i|A0��	.8� �N\s��IFy��'2��'��*L�Ƶ+�O��J�KC4y?�X �IW�P!���4����Od˓�?���?�a���<���/
% �S&@0�:�sJ	���V�'K��'x�P��K������Ok�"(,2@Y��ȆY� Dx���כ�'��ß �	̟Ȓ��n�$�O�)��KG�o�`� �^0J�J0@%�io��'剠k��⭟.���O��Iɯ�� ��_5'By����e��\�'��',�g��y��|2ԟd����4�DBJ�ԪM`�is��4?`�/n��d�O4�d��"Pקug���Ⱦ<r0䝒 �v�_{��7m�O�DƱo��$�Oʓ��O��5Kg��O)A���g��T��46�v�A!�iB�'�B�O�"���^:/�$��b\��Ūr�ėQ+��mH�	����'	����G�=8�����>�D�
7���HemZ̟���ȟ�e'���<����~�B�5p"0�DAĲ"z����ӣ�M�N>Y�i��<�O���'�rܜ0�.B�8���2i��J�,iӨ�d\;(���'����L�'�Zc����R�S.r�����Dʧ&ʸ��4�?�N�<���?)���?�����=Hx��F�V��9�t��*+J����@}�_����Sy��'~��'���*�n�6Y����ŋ�~�.Uر/�+�yU��	럸�ITyRf��Sw�ZYR[�xQ*f��z�"�9��i��	韘�'���'�r�� �y��U|nD˳gV� o4�!E��!�7��O����O"��<Yc��C��ʟ�؁G.��p��
B (�Te�+k��7��O��?y���?�n��<�J�� ���r� `��< ������zg�ig��'��bR�"J|���2rDީu�ڽI�c��"D kÌ	�H��'��'���'m�'����6	r���h�P0�����0?���V���D�$�McsX?]�	�?�I�O���H��xg�G�9��0H�$�M[���?�aA'��'�q��z���/���������D�iJ���e�~Ӡ���O8�D��'�d�ɺGۮ@BdA* P����� �
���4FVK������O"RQ)�d�	��Dk� (BEA ]Q7��O4�$�O(��+�`��?��'��Y���O8��ش�Jb�։��4��i\h�S���'��'���ڦAG��k�e�s�pZAr�<��F�u�J�&�l��՟�&�֘�\�m��&�7I:��v���v��l=,�A���$�O>�d�O��~"�p�7���kݵA����gB+|D�O��$=�D�O��dPx�:���ʀR0e:�BDD �Վ�Oʓ�?���?(O��RTO�|Jc�ӻ0�AJ!�ΉS(�|Q�#R}��'ҕ|��'��y���A.p �eLw�\��	a�xꓭ?����?y-O�:�N B����5�T�C wi��2Dנ7V �:�4�?�H>����?1��\�ָ'�� H���]:��!�ϡ(�`�զ�����ȕ'�X�N%���O@�	C�M��dKu�	�>f���i�42�ܸ'�������Sp�Wܟ,%����;���QٸK(��p)�.4 ioZpy���K!�7��v���'>��>?����T�*1�C�م\b�@@����	�,r��S���O����F�M�L���	*�z ��4� �Ã�it��'�"�O�6c����C���I��pWN��j��MۓM��?�I>����'}���R-W��;��Y�'Ȏ}�i}�����O2�M9Ҡ'�p�I���(�;��z�r��S
j%�Io�d�;*���)����?���J��A�g�9`ԜId랓2ێ!üi�"�� 3qjO��d�O��Ok�G�2xD� @U�F��iA����	�s�0�Iry2�'����\���6ǅb�6	��ϻ^��Jvp�'���'3�'���'�RAq6U�B�� $@	%�ؾAbU��������UyB�P
���>�x��s� �+FNڜJz듞?a�����?i��|vݺ�L�[3��%P��+�)�vhd8��]�X�	��X�	Uy��הt-0���ԧ��V�� ���٤]Șy�� ��QD{R�'��HA�'�r�Od�qH'=Ղ)�0?��Yռi{R�'Q�I lm0@#����$�O��	ša�	�3��< �ٱ��%R1�'���'V�Ɉ��y2Z>�jzDH�/Q�xq̳'���ـ����'J���e�n����O�D�<�էu7S:c���v-��an��J#쏟�MC��?Qe��<�3\?�Imܧ|:5��/�18*�,�eĐ�pG�n�-L���"�4�?i��?9�'&���ayb��5�V��l��	ځ�S�_�V7�S��d�O˓��O�k�	j�� �ի 2tI�D.�sĆ6��O6�d�O(�{p�P}Q����K?�EV�^�k�h�R����$�զ��IkyB�<�yʟ"���O��dV�Rw�(��k�`) �x��	RK.m�џ�A
>����<������Ok�%=<,�G��$��AS+%�F�'�^is�'��	П�Iڟ��'j$t0��qiA��¸BhY�l[|���$�O���?��?��Ua08�oϿlޤ��$@�e�'�B�'~"�'&�Ig��@�O��L �᝽h0���K;5L�aiش��D�O���?����?��`�4�R)c=��B޵"��e'����O$��O:��8��aT?U�	)cv��H$'�� C��y��ʏ(-؉��4�?�(O|�d�O���4��'}�ƙ�uK�Es@�[���Q)��M��?�)O^���z�d�'yr�O6�9)7_�:���� "T}D�CT��>i���?i�n,����9O,�өk}r䣄��8�a��A;��7��<qe�O��ξ~����Ґ��ɢ�D�*�&nÈ Z��p�V���I���ē9�]a�W;���YW��Ot�mZ����ٴ�?����?���]5��gy���9]�����".9Y�L2f�P��6-K[���+��7�����J�KEY�\H�d�\)P�0��X�M���?��fK�T�H�']��On¶�h���pb�����ɦ�i�]�<CaAl��?���?ɶ���x����4����O�T��v�'*u�Fʹ>-O���<	��s�̈́�RLr����
�2�)��_����	�v`��Ipy��'���'�前�|ɑ�GH=�0�w��	��q�藢���<�������O"���O�x����	���6�6Y1���Z�v�I����	�(��Xy�)�?��/:=�U��OD*0z���t�(J��6ͦ<������O��D�O�uC�?Od K7�wKN�q�j�(y8�}�Uئ�������I�ܕ'ԒU	�!�~����s�A:��ݪ�8/�N��G�KӦ���xyb�'_��'Vz�˙'��>����B��"\�EA������Ox��<A�/Cw��Ɵ,�	�?I��n٪V�d���,ϏMe��"�^��D�O|��O���3?OH���<��O2n��ֳnv�;4�N��t��O���R�Rw����O����O�ɮ<�;_�ࡹv�<ZnD�9��X]�,lZ��8�Il�`���D4�)�3� >�@������Zq�G!*�:Ř��i��UZ�q�����O�����4&�H�	�=�]{ō�
Iz�<(�)��H]�yڴS+��Fx��i�O�
#�ةK�	ᑢI>��az��̦M����<�	:�I<a���?��'�r���dDx�(��'���Rۓ�?���?9�2O��9�Gȏ�:QBVሐ  ���'���q�:���O���8���ܩ��GC�d�F��6��"D�R��R�T��- �I۟����$�'h�EJ3-�M�z��C��1)��U P�$4+�OV���Op�OT���O��0%?/:��6Ԟ��;4�F�/1OR���O����OB�
o�n�����AT�U�n
h�u��� �L�nZޟ��I՟|'���	՟\��GS�"�$6��54�L��fK�)�n�f��	����͟4�'g(8 b�/�ͥ~*���\�?=űP���xEnZݟ��	`�v�^I�~*G*�y��\*����(�	��ŦM��ş��Iş��ǫ���IΟX�I�?e�g��Ϡ�����S�͆��ē�?��V	T�[��K�S��!�]ܪ<cL� �qH��M�(O 2�FϦ�h����韜��'� 5�� _�1�5������]��4�?��Q��yFx���T�;���Cr"���E"�d��`�=zQv6-�Ox���O��)N���z��$mH�R��0�ṳ�i�Ҭӌ��-��͟��M��G�(�RH�4��K` ��M+���?��W���Ԛx��'���O���M��h��������㈬ZV�����1O����O8�d4V*uò�;x5���ߣ[ �mZ��{���ē�?1�����We/s�А��ǣj��A@�a}�*���'¶<��@D��d���G�����e^&���ȓD���[eI�Z���4��rHuE}BN^>T��ř�mMd�P���M�̵e/V�.�pYzv��-h� �e�N�
K���qc0�yB��	nJ.�I�*]���9��� �LAeb�r���ڰA�5"��������P�/L�S��^{X� �`X"� �HbA4S���x� �*~r=0���&C�4��"�kM��E�\�U��H��l�,(l]9��?Y��1�艉q۝T+�,+V�R���P ��?9ʷkP�54jL"�k>�`8Ke� ʓ|����Tm����+pM��L������F��};�fFx�@q��)È�+Bo +��'B�`��?و��-�#z���D0^ ��r��2�y��'0T���Q7����ڏS���*�'T@���c<	˴�ЫD���@�'�b58�>���򉄄���$�O����!3��U"��������!�"��XK���>u�$h�QmC!)���|���|���X����o~8��r(�:�����)���W�����������ӇX��ݹ� W�FF�����רN]0q��';B������OR@r
�84_�嫇hӈ -�|8G"O�ŉ#{d�V�ϲ�ԣT�	*�HO���u�fԋW��P�7#זh[�T��ʟ����<�r-�I������\�[wZR�'g�3)<��5i�Gߎ �⒠�O2}�r�҈v8mH�ܺ�����ɀ�h��@�)�N�XKխzs@��I9If\��
��U��Yˤџўt���G>\�JC�R?6�!�fc������O��$7���EU������5��Y�T�҅"!�D��b��l�bƣ{���+$gڥEzʟPʓA���`�i���qn��oҨa�Kb���x��'���'8�ܰw�',�	�X��zfG?�p�bi��6��|I���Y�6����i؞T!u�4���8�!��lQY�HR'
�9�
�%0�p�Ysی5�����!U���'U<Y3�&Z"��PIڦFzx5h��Y�'K�K�옄jDt37��&�8��'M"+@�\7O���h2M0��'[2���B�!4�d�'�RW>E�� A7S��pw�]5/tV0ل!N,>����ʟ��	�ew
`� 	�sh<y��жt��x����&���7���l6Y4�.�! hfK�(HO��ʲN��j���c�e�@iY5G�)u�Œ鞍WĊ7+B�c��O���P�'�2�)�v���E�!F$�� ����1�Oʍ�P�X�v�K��\&����'�O:(UI@�o2x�񠋯`����3O&�Z�AWq}��'S�35�@��۟���%U�,!J��!.ܥ���_y$���ܹGjT(� U8�,��|ҋ��p!Hiz�-��?x���:�2�'�:@�Z�����I�n�S��?q'��}8Mx���U0�"�\w5: ���ٛ���<%?���Qyү�	8�l�Ke�	 ���,�v�<1��E�x/*ؐ%�_5)�>L��IK�'Ă#=ٱ�igbf��*�^YQ!�]�1u���6jd8��ą�l_�Mc���t��P_���%"Od4#3p#�`��(��4��* "O !j�2\��৊�%�LJ#"O<���u���	�_�8bw"O� �}j��A� ج�H%(J�XU"O����Zu@��I=�(�0"O�H���`���K.�!D"OL��!�P9V3n�b�.&L<��&"Ot��!"��\pQ7���1>���"O�-K�MԮR<p	�ꏄa"�J�"O�SUG</���iN�HD�C"O�X���.z�La��)�= �nE�%"Ovp��F��V����ȜP �0'"O�I�n�E�v%A1�B��)9�"Oh�Y��ܠ(�L���"��R"O�t�z�Q�d�����"O�5h��M~vL��dV/g�6Er"O�\��B C�\Ej�d;/~���$"Oê�=a�zY�Ei�3s:8��"OR,���ŭ|[��F�J�"iC�"O�a�T��8�"4햚\h>��"OteB�;X��)�%�ƲR�dY#�"O�Q�L�7<�t	���+
�2-�b"O���Ս�%a�� �գ.����"OL�"��:}�pQ�5 ��"�"Ot)��k��6u�T��Y
JE��"O��Zs��&d�­�p͊;U܆Aq�"O  ����L�	跋ߙ ���X�"Ob�C%���{���  ���\h�3"O&S�gK<81b 
�dؘ��4"O���0�)�d�\Ø���"O���
�g��0�E-Z��b��"O�H΅t���M�9A�f"O�!�̥H�l�(6�i&�I�"Ol�j��,1��=�f�<G)����"Ohe��OX(4;�r"7U(us�"O����7v��i��)O���"O��"qd��n�|cEɍ`^,�q"O��I��Y�8E���Eh��m7�� "O�d��<+"T�y�'��X��)��"O���r�˪V�غ��_�X��0z "O���ӄ�7S�����DkȂ���"OH�"�Έ]Q2�pDŀz��(��"O,]���Н��Б)�$Qnd�A"O����޺~%��+q�K3eJ�r�"O2���K�e?�h1�?>�p�"O�y�[�V�Z$��!�Q���t"OLᑆ�i ��i��a]��j�"Oj(����XԤHr���Q>dS�"O��3�Y,w����hK�g��Kd"O�X�T��RK���_69[��kB"O��B�'W>X�LH�&e`8V"O�����߿n`F���Γ/Vd1B"O�U���~�Ȱ@T`�p��eP�"OB�����H]�H1��ض# ��h�\�T����ا(�8h�(M���Z�.��jA &"O�e ��Đ`�j1׌��Zڽ��|R���^ʝ��I;�~�����w�X) ��`xb��$G?�n8xܾ/���H�TV1�5�#Ą��x��($]6���
��C\֨�������O�T� �(��Os������n�T��F/K=�Z�z�'�$�s��64�X@�f���D�&�8�O*����e�S�O�@�A`Iӽ2j&�)f*��e�Δ��'7�i��(�$Foʖ)`(���'�~L�� X/~BZ�c夅���M��'�n-{ "��V<�+��ۭO�9	�'�05�lC�?�XK��y� 	�'�$A��͝&jɐ�H ��b��� �Au�I�t��"���Yd�ru"O|P�T���T�@ߖqCf�X2"O,�0��Q)z�X��F*i?�H8�"O�jw�]�o��鰤��"@ɑ�"O:ɐ�玌U�|#3��
�~z�"OD�`��4:��BG�ӣBzF�x�"O�}Q@.G0P�"�S i��?kp̲T"O���`f�<v��i����=\R��D"O�A����2?Xi�@�%H*�s&"O��B���=S'��!m�qC�"Op���R|��Y��݁֝�"O>KB�>~jh4b����H��""ORص�!j�����>G�r"O���/��snr��&®4��rp"O捋e�[2`�B���uDH��"O΅���_,�fU��o�(6���"O|��� ��8]��oܠ3�d���1O x��2�)�a�$�3�ѫk�b`�Q�^1@��XeP<h$�D�y�Ĉ�V���'��1���'���
��<��ҸU�����q����a܎`�1���D�(;���҆�
�b�r'�	��x�fu(&� `I\"��=�PmC<�HO�
5��pS�� �1��U ����?��(2�&�7u&��ȓ0~�RB47*�,P���3��|o16� �`J�e*Pqg�O?7��<"x�c'�G�+a.�a��u�!�$�[�"Ы�IZ��dI1��5`B�I-/J�Cr,S�aĩ���i���aȈ/Z��� � [�}��g��XY��"o����I�n�6�r���8JGX(��$�_�������jh���Y荑�"�pֆ����Z�gtpe���0�I���V���( G<i+�Bk!�DL� �$z0�VpJZi���3jG�V�$�f�IBQ�A��}�S��M���E9ԃ��I�o� q�tS�<y$"��%��ԁR�C�W0֑�C���~R��Z������-"�<F�#Χv�h�@�,U'1��yy�A����>����������	+����1�]=5T�U���/X�`���*�Or���(`���b)Ղx�>;��ɱyLTKmQ 7x�M�����%��R������&Kt�(�O���Px�BV	}�	��
1JG�e0��4Hx`1�3� O�,�r�M&SѼM��?O?7mP�x*��צe�ӡ�ׁN�џL����O����ųi����䉛mb��0靆&wH�I<^�����.�L�hjv��q�'(� {".{N	AÚr��Q��'�p؁t�X H�֕i�T�ā�ë'� �	�N��!y�B�:}b`)q*�������	�*����#�q��� �+O�|�j���'����n*������h�Ov�+�gK����lv�]4<�@� ��L<K��qd/AE����$Q;�E����OB�{�ʽ2@�@.+�)Ҕ���)l�&qF� !���B�y�?5�7�� �~�M
�f����a�����-��O�H����}>���Q���	N1.5(�惛�nD��ʠ*n��K�,��(*�V_a���0*=�>Q�k�L���9"�8���J��<�0�I�c��q��ٟ!DL�|�'Ӕ���)SHB�Q�3�KS�`��a��� P2ԃ %�p?!�	�/a�2���,PO�@��YbϘ����d�x���<�-�#���}M���/���C�l:+<�񦦚�.ߦ��DJ�/S }�p���]yW�%	<�A�')V>�2��)K��(*�>Ho�-F�\{���~�؄p��?v4]��DK	J�b�E|�G�P��a�Ϟ�K�i���!����P`�9��c����a�A?�?9�3�I2"�_6�3�
v�����O$��{AO�:X �y��E��Wt��1��r�g?AB�UEhQs����W��ڠ`��r�,`P�W<���$ �hg�,� o�zݞ��&�a����'����,՗pQ8�ɹeK,��g?2�ĝ���.)� 0ۃ#ǹ*�d��'�'g��5*�$1�d10&ָ`����e$Ȟ+����\ S�b��c��]��@}2&H%����4FR�#TT䙢�!Q��}Jt	�d���!����JǨ��7M"������O���	˲�aF���r�TVbV�J�)5�[�����Uk~��C#P<t��M�e��TP��n�( ��S7o_d Z��^埢|��nN�B�F0IJ �z�� -Q @{���4��$�'{M�	tc������)__�x���'�F(�Ġ_
.�P��=���c��	���O� x���h�*����
m��H�5�'�Pi��NC�=<��Y ��~'~=q&D�28��VIE�c��'�$��U���`q��ԏgN��XJ|���Z�s����EB���}l�OeY��=�|Ȓ����>P[�E@�eL��ԟ�肢
Z�,����HmHș��h�p`��ڒ~L��Ў��Y�����YX��{���~��u�C�S���p�I��W.L�S���W8�81��*G$��~&���*O6[�;!E I�XxB���]!�e�1�>(>6�K��	����%����[i@x+U��O�	�D�'8Ha�����ɧ��RZ�1�P�x6@[�
���'�<d��i�:�r��ԟ�o>r��*��^�p68���l7�*�@~�ў��Ӣ�Mb�k��-.��9���@���!h�9u�. P��h�̨��X�#̫'xd!��MT9'ƠEic���A�ҝ8�Ob�ɣK���`-D��(�3��*4�@�D�/PB�5 �|>�@� ăHQ�1VB��L2p퐄�N,x�$lrsi�0#��)� �.P���G�Fx�8*ơ6Aؖ�[�lL,M(�	b���"�jaߓ$��hB�Va�Beʃk4r؀-�.�IT���8,l� �L8:-� �J�d$��S"�v"l��K��J�yF}�A�.9-b��6L9�����$�$�0�EI�M�.��FƖ3 3j�Pb͌Z�D�z��Ŝ:sڔe��R.�l84�V+eV�	 F��ɱ�Ќ=��g�*#���Ę�h��yBD9)T 1H`�_�]f�L͡��I���󁡌�  �"��z4�����_��)

�b��!�ǣX���O!R�`�:=FPx"&L�@�CN%�ƭ��k�c���RD�pdџp��X�}�|�� � mk��"3n�8՜E���'�i@�9�*���)��<!�9�EE�^V�Ǧb�6�җ/Tg;��O&Ē/U�Mc����f�^QT`��@��"(0�WI�s�'%Tq��O戩���tZI��'Ov} ��� �6`f���8�$�
2hvЈ�4i����Ǧ�6~��yb"� �i���� rF�����C$�'k�2�^+4X�Q��"������8b�D�6��P�L�1\N:��4X�l���<*���y�H�|F|b��0�6@�DÓ	>~L�$E����-��E���T�NYx��?щH��A�	\<%���ElI�1�8Q�u	�������+�O�Nǹl����d+�
l�v1s�*��y��ɂ��6���3��͉p�?��vn�ēO���B�,�PY�]4�Ϣ)�B D�L���'��`�H 4- i	�\�5j~�كχ	A����P����$SE�h�mR�J�v�Q��Z8|F�	�M�:#<�2�I��)XD%^?1�+,�i9�(�Bs���c�Q�<���#9Ѱ��V`�S�I�W��J��W H�S�Ū�'� �O�b�C��)�L09���<����'�r�P㌃%?��P�jL�@�ݙs�ަ�y�faV�}���H�w�� Ȳ*�&�y�N�C�Ph��׸g���Yª�=�y�㇀nB�	ee�nQ �R�K �y�gӯ.�
��T	̡z=zyȡkT5�y�G�K��]���l��!�1���yBK�X�����n��-�e�y��z��Y���8m��p+�%�y�)ܘv���
U)�}���y��ֈ�&!0�J��i�t*碊��y�oK�s+(i�P'�2|�vb���y�	&ܝ;�
V���M�W�y�ꅻ}���)�aOl�T���_��y���[���_¾���،�y�޴h���QqN+F	��SU'���y�	@�;nR�AAɵ6	"�#�a�
�y�M�nLM�!"�'�<Ễj^/�y�>�p9R���^��Ƨ�y�`�pw�932�T�B%�CE��y�o� �6xb*C�j�h¢��yҥ�h��Zsb��04T�"�=�yG��Z��j�F�4"l�����7�yBl��Z$@M|X���E?V[�C�	c�<z��ևれ�j�8ҼB�ɩj�X\[f(�PP��"0`�6�~B�ɀ6��S��,lK��u�ߓ6sBB��0�����Fð`cXm;�aL��B�	�	:=�C�V6sD4�&� ����	"�.)F7U��AT�� *Q!��P=X�dL��`9��K�R!�� R|h&�\<մ�.ޅ{1���"O�5����)I5@Q{��
� 1N �a"Ox˄����YIw.��x:��D"O�lPv��lxB5-C0s���"Ob��	��TЃ�l^�`��̈�"O8�ƥz6�P��}�N��"Oh�Kpc�sD�C3J��7ò�v"OF�Pc/
�%���!�]/n�^���"O�$sҊ�=}�MӰ�˼-���S$"O����`	(Z'�l�tb��4��EI�"O���'AH�~M�hEpg��5"O���#Ö&_
)�c��>T� "OX����5>�����dI�:���"O$��@�;�r�8�#�}6�1��"O�Y`�P�] ���B�,Q�d��"O^�0�&L�l/=uDx�`"O��t$^,G��.�	=�����"Ob���gU�|,��"�(��Y��"O�\�WE[1O}�;e�[�ֵ9v"O,�����sHV=���@99z�l) "O�QA��#[j<=a$O�;nA��2%"O�� f�Ǻ]$��G��W1|��u"ON�Ɠ31�,a�P���Zy�*�"O4q�`��\�H\���C{s� 9�"O�0râ]-���M�_Ȱ�0�"O�����Cx�� �Z��"Ͱ�"Onܰ�(ސ6ܙ�Q�L9X��@B"O҃�%��={�m�����Q"O�$��l�;?,���mG�T��4��"O��
џin�Q��K�}���"OM��'��J�Ҥ��LOF,�T"Ox�"�l�{�1B*E%v��E �"O�]�śA�TH�H��it$�y�"O�I*5,R�����X]Υ0�"O�%	�i@]��@&F�~n����"Ohܣ�+C�|���a�ƲzX����'	4�Q%��P(��Ei^�Y��'�
�2�G�%GI�*.��4�X�<i!�9S9*�.�)՞0�fQ�<i6�M�MՈuh0L�I�����G�<��_-K��)�N�vF�R��n�<A4�3��ՙ@o_�P��Qb�`�l�<�O^,@���r��|���ǟm�<�R�O�-��p�ࡒJt������A�<!�\�Y�$ �jɄ/0���I�<aw)N*5���G�)zI^�Zn�p�<Y�肩0�=�ь]�C �1���q�<YU��lY)W,�c�B�Q�m�B�<�2�\�Q�`�di�� ����TB�<��Ǜv�6�c��A�4&I�d�d�<)bJ�4S8��%�	^R�U��g_�<1��v�5R���2�-:��_�<��䊃�z��C�ƾg���J:T�A�/#!��I A�n��#�-D��
peƸCƌ9���Xԡ��$*D�Dy�ɔ�(�HGC�0Ť��*O"�2��$j��ai��%���h�"O�)�È*z��X��9�P�P"O��+�i
�(*4ʄL�"'�2h�1"O� �+\�6�D�)����"O,�c&�y��k�D��ޢ��&"Od$K��_|��CD��8��"O����'��x[�� 0�3�"O�y�dà-�X��%�#�~Q�"O� p�A�@��W�<Hs'Q�
�dmi5"O�gKJ	uEֹ��F^0Z�p��U"O��t��8n���;Ŗ'zsN x���l��ɏ���	�]&tD�jW$B�	.��� &���v4H�U�9+B�IMY�9Ja���>r�k��3�C䉻m�����վ&�h9�ޣDI�C䉽)�8���ꄆ��:����zC�ɝQ%D�Ǭ�u��� ���<C䉀d�DD{��N�b1�3OX�p�jB�I�(2Z��Ҫ���
ѫ#�< K4B�I�Y�^�(��
�`��E�Ͼt�nC�	�*��pC��H%	��^ 6C�*j ,v���R�&�:��#:B�IS�@�HA!K"
��Ѱ_�$B�D ��� �H�c��\[u�\?>w B��
9ź]���6h1�HP�ȘO B�I:N^DT;Vƫ{6��(���z��C�Ɇ�xp�&`V�"a���gT�	��C�H�Ƭ´-H=/f]�rDԶkʔC�		FP9��D���c���[�^C�I*]9�m�����p$� !��H 2C�It�h`�%�5PI:�s�|�C�ɕ
��51�W�(�,��h�?��C�	X �[B+A? ��3�ʱ9~C���. ����[<ʤS��0�`C�,�ʀ0�Koil<�g�OtC�	�0u�9���<o{L(w�\?#�4C�	�p����q��?A�K�-�6\��C�IJ���c�GݨGB�`q�IX	s�C��$ʺ!�b7�v�{��Cf�C��(�{�j����x!�K?&C䉕mR��N�!4�0��h��ھ�Ic����^\x��<uD���#-A�^HV�ۦ"O���L< ��L"e�C@��� D��pD{��	[#�y�1DΜ:�0��g-�O �=%>Y:���ctXفDɅ7��,���>D����(���0��@_�iIʜ�f�<D�X��Z�!���p�"Y<L�����8D�l�THE7z�(�؇�U(v��H�):D����kV`|��W'��<+D�X�r�G�e��5�F�E�N�x<p�)D���혞LH$xJԨE�gyDXJ:D���%CI�:�X�x�l�
!Y��d+4D�ԫw�GX�@��&eW�&W�i�	2D���왹p7J��"kY�5�mp�-D�p�1��j�R��Ɣ�L�3��'D�lj�)Do��9sG�'3H`�,:D���i���%�N����  �3��C�	�F��5���ˬ2%@��p'�Y��B��^a^17*��*q�@���"nB��(~*T���ͥ*>I8r�ִm�B�I1̬`qhM�G��T�����L�xB�#3���#g�\�
�HfAU,/PJ�\��	6�M��؎%c����B�A�PB�	
�D��� t�aA��ǰixB��g��M ��j�$M3ǾX�VB䉛LR��@�k��p��1
磈���B�I*՞�R��'�ܠ15�J�%z�C�	&8Sm]���x�ԡD8bX�B�	^U����'|sv��'hò<�B�ɥݜ{�b�{~��B�	�|�h�����n���W(mB䉃#k`m�:7��	bUY�L�.C�)� �MK�0$qFG�%5�����"O����&�M�\�������"O�8�)��u�])e&P4y���s"Ob̑�)˅7�Ƒ��,K�H��"O��i`��a2�ZciDVQ*�:@"O��	�I��Q�F���\,?��@�"O���dJ1��IᔄћLHH��'x�"���$}ځs" �'��	�'v�L� �B06����Z�R��<�	��ē���8$CB�F�Ѕ��N�t�*��ȓ�l���'FI��	�EH��ȓF������4G����n�Y�L���L;������)X/8���ύ6l!��
`ڬ�WC��RU�S�\NVȄȓG��TG� �DI�{G�U!�Q�ȓv�2�����60��BU��E0t}��B�����W�20��b�I�	T:���.��2�߂]IZa:���>ײ���NƔ{�#�P4���OP�L]�y�ȓR`dxK�DM�"����2q���6��q��a#{�*��w�0G݌A�ȓ^��W2?!pp`��@�f��Ѕ�Oψ�E�&���)"�fp����`XWnD��h�[�D�"X�}�ȓQ\h[�KYk�S�&BB��ȓTx��;�e�G+��ʳ�{8����,%(S#�=>0,�͕?�^܇ȓ'Z��B5��*�p0"���0�ȱ��uI��5'��Z�"!ҥ��.o�"��ȓ~���y� �4KZNl7�D]^@���ptp�bI�M
|q��+V ���h1E�T�֮P���׉��}�t��p����ʂ)e�$�LO�2��D��H��8)%ϭ6���q$��.C[���v�Q��C�(䡑����q���� �FE�rMF��=y�f
Vͅ�~��+1́/���Hp㞸D���ȓk���T�
�*|��c�9�X���(�za�A��p!�q�p�ݲ{�t��ȓL-zL�UN�<Dn]AW���q�ȓ�@����؉;\}8E�V����9s��f��ћg��.�ބ����<�We�7V��K #�z<����A�@���<3��x����1�ȓrzb����;C	�9��eY�5����{o�|���	�R��}8��K܅ȓ�"���O��@|H�[�v� ��P?� � ēi��C@M��(��c�`��� �X��fٺv�T��u�4yB%`�a�E �˶L.���ȓ;D�4�ΜS�&HS�Ȱ%�����J�pGIUnL  s��3_͘m��xSR-�'l�Z�x�ҠDͲL�*E�ȓd��EaI�
��8C%Ҭ<�h̆�P8���%�1Am���"��)N ����s�����_ "nR���&!@,�ȓ�łuG�3h���S�����6\�p2% W(Ե��I�!�F=�ȓP���Sm�Xi� �9U|-��$>��񋁞Rұ"eBnڀQ�ȓ ��P��)��	q�Y�J*�q�ȓ3
�tĭ .x��A�O�u�t�����ɴ%�$���Y�E(\C��ȓ}�~�(���1B�\��i�#/� ��S�? f��Q`R��4%�NH�(t8�"O6ճ`lКT
�<�E,_�lͺU"OФ[e�G�t�v��AkƗ|��}j"O�{�K4�	�%� ��r"OJ��BC�J�2�!ċ�%x#=�2"O�I�F�:�L)�w�{���s"O��ksD����@$�!Z�xͩd"OFPs�O��~�|mKB�M�U� �X�"Or�V�E�v�(����V 1ւ!�"O x�p��
L��cT��z�	Z�"O2M�1.�?`��CN@>a�Vhsg"Or�`�"�:�\|�aʟ=U���[A"O�ؒ$�4�+ ;x��%�En��y(8=.�]R�W!r
%�%���y�I�47���G5'���YţM��y��Z�c[��R2+�)��rM�6�y��W�*"�ha�ݠt֥	R����y��> �(c��<��{!��3�y��*/iZ��)Q�4�0آ%�3�y�dԈ�T���\�%���(fN �y�`�f�e��BϢŁD ��y�/CZ��J�#P
=ae��ʵ�y҇�dm���'R8��)���y��1s#j|����+Z64�b�y��M�b�����gF�U�n��� V	�y"��4*@ά�&�Q�N,:�o��y"���*X"Pn� vg��r��Ԝ�yl�.q*2��g��cPF[��y�)��l��YQ%
�g�xш��y��t�	"�,FZX3wM��y"!�8Rvu��AZ$��E��lͩ�y�P�]���h�ǃ�&$CO7�y�['�4��rCY����R'E��y����t�=Ya���j���Z9�yR�IN I0� �h��pv�J�yR��%g�֝Q�Œ#aA2@ce�P%�y⫀"��� �̛opp5
���yҮ�W�.17g�f�����`7�y"��8l���s/[�Z?�qI�����y��2[�>����jT8IU����y"K�)��TɁ��a�.P�����y�E�8/�A�%��n�@�K���'�y�E�?0T�y�Ý�hE8�L8�yÙ^��fĢb��lR�j�3�y��J~�a��ݾS����iS+�y�a�dm����Me���)�y�+-xP$�H�C�R�
���y��;7�L�s�Q�I��Y��K	��yr�E6-�椁Q�ގ/�~A؅�7�y�OO-4�l�_2������4�2�ȓ�f��6A��|���D�d��ȓ��@@�H��!٣�\=p�
���4��q��В|4���*I�>�مȓ@*�y���@D��C�p�x(�ȓUm�A�1o��A�
Ա�!%j�p��h�$��&�=+�(����I�D��_(`���N}�v�aO�~�6D��5U&���/޹"����4LT!����ȓb�ҡ�'��� ^t�F�D8T����9�"A���<S ���NP;u�I��)��XP��!p� ��Ȇ�N_��ȓC5*I�� څ"��	������ee6���C>c�*�����h�p؅�a�X49-/��f�S ���S�? &A����<N^�:E'J)G<b�a"O��2���܌X��C�h(4�Sf"O`�i�jT�_Ř�(e%R1*���S`"O�1�E��6���ö$�`��pA"O�49�CT��l�ا�@*!~`�۶"O�}��C�a�zM�ai��>ɶ�"O�YP�C�H�����NH(�"O��6�\�e���#GHY���%6"O<�9����z,�P2��#�:��"OV�s���uJ��$��r+�)�`"O0dibdQq¥+"o�%�h��"O����ʁ�E�ݘ#dЊ.W��7"O�yh�F�/[k*�r5�N�qLm(r"O����g�	
~@��tkȎ�V hB"O:q��eX8ˤݸe�P&x�F��"OH�3.T�?˰hP��U�p�l�I&"OLqC��CD��p�(��D���c�"O^=kϺ*`8�����L�S"O@<��+K�vVh듊Q�U
G"O̹��(ː�*I�s�ܴ��}��"O�����^�(,z�G��ɶ��"O�(�(֔mabT�T'ʩQ��9"O\�%�3�nM��H��n>�\�"OPj%�#x�e.Y$�t��"O���*�xcCn��jD!YS"O4d[r��U��L�@�K�"OD����L�Fu��I�!����"OVm���S-��h���	-Pi� "O���$]d��L Ä~u:]��"O��I��݋5�����c�1r�`�4"O��1V� .�(f�I��4l�7"O0��`Lҝ]l&�"⒗d��<�"O���kN�I�� Q0X�e+F"O8Hpp�ϝ��@��Α�9OH���"OV�r��V�0���{��˯>��kS"O��F˅�T����Ĉ�"�y��"O���D^�0Lf� �˪E"a�"O�����&MH��ܴX��X 0"O��g*cj  �4�Eڣ"O2���_���RD�s�Ii�"O���&U�Y����B�iȝ� "O�4#Ԩ�*+V��`�H)^0`ň�"Ot�ðH��x˰�ɫk22]S"O̵yԀ�𼊠o�i�!{�"O�[E�ޑYk�@�f�#`9�"O��E�ȿJd�0�J��F%x"O�x���8��h�o
*����"O��P��.#"����N��� "O��* b��g����"�72rL�q"O$I�"K.q,�yK�!>�`�"O:(�C�;�PP���#�t�%"ON���g��L1�Β'?����"O<�$O]f�X�E���N�lyY�"OTm���*}���Rr�e/�0P�"O(A�``��"������F�{$jD�"O�IubU�E{�i�'��7`�,X�"O>��@�%^0�9u�ջ;�TMӦ"Oच�)F�!��:�.ɨ"j��"O"���"�X q�M"rB��"O���"��x+bI���<b�苧"O,)@`
���j���z4@4c�"O��I#��J�������}
!"O�,j���7� ��m�a,(y�"O��Rh�%%�Ap+��i6l��"O� f]�c �$#Yl�[ժZ�d�4��"OfMjQ�[4io�@K�ɕsX����"OR�2��S�0�i@���/�N�k�"O0|[eH$;Z�Ba�Ж ��|c�"O�
PJ[8��j�N�bYF���"OLQ�𩖣y�h�֭�HS��"OVv���9�,��56(pQ"O��v�'�<aK�K�|�X���"O��a#�r�P��6>���"O����fL0d@���e9�:�"O�,C��6|R�%ّ�Q�P��UK��'^�O���@�6��2ա4�����e��N[!���7Vx�3�'eN��1k��c�!�Dڑ4o��j��H�#߰x��o��v�!��J=M����I̼J�\��LC�!��R�PĀ4���E���ҭ�Fn!�dQ#	�!�A��6 �и���W��!�$��r� � .��y¼��!�.sRO��2d
}�
q�1��Fm	"O�q�FL��(��8&�V���"O<�#�B���)���9Nx��"Or8k���L�3�K��Ah�ѧ"O�yI0���r�w툸#'2��"O*x����!!=��Q��6�L%ږO\��Ʈ��Anh|
R%U�BLU�T�bʓ�0?�$�ݧpn� ��o�-1JZ(.DQ�<�AM�$ �t��Ā't�&��#ZI�d���OrTbb�/k�yH�¤*��E��'�����?i�B@�%��"M��(�'���&ζH��9ɒ\2O�Ƒ��'b0�s�f_�B���a��E�����'��e�%OȪt�"h��ǟ|�<��'�?V�A;���t�<tAfx�<�f��1�D��ɋ<z�aA�M�H�	x�S�O�L��A
�Y*� '-�VD��K"OR���
�6�yE�1I]�Q��"Oh@���F��}9!�bR�[�"O���h߰x��U�%F>���JO&ђϊ"|�RYB`
�,%����#D�����_|���D"��|ƒ�Hd&D���矋(|(��T�ly`u�@>D��B�a�/ހ��&٥a�p��d8D�P9�K)/6}[���%R��:��5D�\A�P�'�Hu ��׍7�~Xr D�� �� ,j��'*�B�2Ç1<OʒO,�	8~Vd�F$�% h8�R�OE�m�C�ɗ',��(1��r��R�̂�-�JC�0W���΃(aRLQq��46C�Ɂn
�=����]�IS�M;3�B�	�M�QrUD�;E�:�)0�B�	�5<��*�eM&:���Y����"bC䉫}gdd*���7��H ���$TC䉜L|��S&�(���R4#�5�8C�	;@�&�Y�+�yy�<�R�=F"�=/O8"|*5o_�Y���6鑍�(�W��U�<�,���|j�ˌ�}I�ڦK�z�<ق�٣s���"�#���BB��Z�<����Y*����ۄ��i��mCV�<� @N�=j���g�>p��Ir�K�Y�<��o����u登7��1e��I�<�$��nX�(����pe���M�'�B�,J&�#R�Նv�P�e�ȝ`�C䉺54��i��}8��V�ƽR�B�	�f�N�R�C�(A�r}맏�4rXC�)� �ua�	Tq�EC��_�%�, �"O8h Fnߝu���b��xE֡qQ"O���3�E?` `Ѓԁ��;���R�"O��Cg�K#5��y��'X�j�A�'m�|{5/Ў+b\��Ԫ�:DTcC;D�,��<P�PPT�I�{�u��-8D��J���p�f<���ƛ7���g�6D����\.8��H�2f&v����)D��z��)m4�Y2���p[���v�54� �Ħ��{ܮ�g��73L����`�<�6#��e ��� �ݥL��إ$�^y��)�'�2���+O),D ��@l��|��ȓ¶q(`��u�~%���N��R�����1�΂3}� Q{ի�<��ȓj�u`$N�?Ơ[�NޅC8���Gx�r�E��d��$���E4�4��T9���O��.���W�(Cx$�ȓ<�ޘ��Ş�:�0�Y��W�6�l��IPy��|ʟqO����W&?�H����	`�|�%"Op�#����p�<��N�#�R	J"O��!�D��(�� � MƆv�r�`�"Oz��n�!oH�z"L�= ��&"O��#�(5���6�U#H��"O������B�����ˆ@�xH�"O|��B<H"�!�o����"O(��Y��p�Ӿspt�����y�/$�F�LMr��qt��/�y"��/�l����lB4S�o_�y�������@/�����J	�yRe)٤�+2`�S�-��yr��G��mh3BL�h��bA�yR+��<�i�~�z��-L����hOq�X9@��F�Ƞ�
m��z�"OTu��-[-q����a�^�J�N���"O����]�Wj�fY�0����"O�E���çz``�I�S� 8xC"O����
�Kt���	o!�ā�2��}{��T�o.<��ək!��~$��`���L|ݸ��b!��Un���E�HK]32�&�"O�б��=�(���Ð� ;tM�E"O X"s�D(��� �S�6)"O�0�c���ͰF!ŊvQЀ"O�{�垨\��5cd��<�6��"Ov�㥢��h� ��Q�J�$y��"O�U�EfI3?,���Aʌf��LC#"ON�R0��v�,�"�)�t�A�&�'�ў"~QJH�.~�DR��8A6(�.��yR�^�>jDz5��6���@�&Ȇ�y"��H2��q�\�_���{���yR+E�*�L!`�A20|������yR 5x��(��Swl�tY�	L�y"�@���@ b�M0���aIL��y�Y�T�W	^�z�ڰ�A^�y�e� ; aۜJ�xWL	f�&���:8��;a��A�xA�D�\:g��ȓ+���g�6V)��
շ.l\�ȓR��6�o���R���:�G���/��S�AL�6��Q����C䉘w]�����Z�]��8q���	��C�	9Vԫ��'/.�@P�L��{�xC�I�S|t�d@ԣx'@�D�0:W�B�ɦqS��J*�,��K���>u��B��+�Uj���;��{S�Ɋ' �B�)� � �ą�N��QG�É�عq���(D�Ԏ��u��l��-�`Dr��A��yҩù��\�@��Q-��%�K0�y��l��@Z*JH=�4W��y��U�)#tP��/�o��:!���y"@�-.�Hd��o����KR/�y�lT |+x��UŞ�t����yr��j���q*B�e�⭀!���hOt��I"��Z��ٹT�4�q�K:�!�DW�H־���N�������#~v��)�'k��[�oX�4�]���0h��Hy
�'jv-�1KT:+H� �Z.6�X��'�x���I�O�а���ӯ&,�!��'�8�֮?kΆL�&��Ko����'9�8h �G�QFąB0BC�s�D��
�'+,��Ԩ�1�y��n��$�
�'���Uaױ/�������iLt�
�'8"��F��?~*�xBM�h�Z�1�'�t��f(��|a0�pAHZ�H	�'�0�V�|��=Q(ŧB��!	�'���0C��(߀Eb�L�2v&��'YV�2Ƒ%a�j���H�/s�9
�']b�(��H}���P�^*L҅�'��H�1j� 8Jb�*U�q�+�'z�0�IKT��I�ԡM�bT� �'���ҐhTC �h�N���{�'��q����W��s�Њ4����'�� �.&Z�ЕnT�; ���'	~���N�<��y&�DZ������yB�,L�hje�H�d�I��C��yR�ձ<�(��H4XLl����yh�]4�(;���U�
ܰ֫�,�y�&�'�lPU�ڳ_��-9uF��y�c�'TPdI��ş�,~H���bL��y��$t5�}�1$d)̑�y�3{� �օ��H0B� s(����>a���y��-Z6x�S�G�U�X��y"�Q�uY�lQc,غrFN�{p&�;�y���y�8�rr���X��E��y�H��Oibe(0-<ޢ��b)�?�y�ȡ*P�D�"�C���37��<�y�à(K�"��G�,��b�/���yR�
Y&I��ȉ�m㲁�BV����!�S�'�y¨_�"鸱$ʬw��Lp�Ŷ�y��Z�{hu�AɊq84i��B��O�#~�s`�0DUTB5ĲUm,ܸs�c�<a5-�P�ra�-ɷ��%�s��F�<�#ʖ �F!h���-��p`0��C�<�����Q�.��FجY�,�:��C�<�vN�3V�� ��\7^��@�j�'mr�SQ�T�n۝8�I����qK$C�I/b��43gB[�#�>��Q�R��?A��?q��ԇK�P�s�5���5d?�y�4t8 ��킶h0	R	ځ�yB��4rIH��E�C'*<C�@��yR��XX	:1'��$(u��0�y���	>�TRB�(-h��ө��Ob��-�'�5�f�N9f)� b�P��H�ȓ~��yCD	�>��"4DȨ
�^�D{2�O���7�J7H�X���ԾPFL��'O��bg�=Ӵ]���P+G�@a��'� �С��b�hh���:etmP�'w`h�6~�F�3��6.��P��'
^M�'�_46���B'��}���� �� G��v�)�O��>}@��"O�����"S�,HQ�I �4���b���_�Ooh��l��8�& <L�e��'m̡�R��I`߿"�����'GؘC�N�o�&�qAâm}�X{�'!� /M��`�l"���'��3򢈌pD����]�zE��'lt�D���W���JT�Z�X�L(�'��a��L�<<���C�C�T{ʭ��'@���˸7����ΒG�,)��'v�Ȼ�⋥d#�0�M��
�'l<B�HI�;�aIwH��tD�-�
�'&��e�h�sl�l��k�' �����D�j����Jں��J�'(^�����C	(LsA�"Ъ6"O��"s�Q�+���cF�E�J"O�5�l����%� �Z?p'D#�"O �ޖZݠ���V);ޅ��"OpI3��]�:�R�/@2.=q�"O&){�/
�~������uhDeC�"O�9f�$;������LR�zw"O��ac�������+O1Xh��*��D �S�	B
���j�ЃU�X�!��U$�48�#�4$���{`��!�dԷS�����h}�O1�!���(����[�@������Y�`�!�$(�P,�j�-!c�e�&��:�!�$٤'��퉧�]�SK�x�'�ͨ�!��]
P1�(��;�Q;��V�/l�'P�'f?X�X�O�N��w*����� D������&ʘ)�'D��D��!"B�>D�@���4ת��e�Ҹ���$*D�t��+F15D�Z�n�h�	-D��"�Ɨl�ܑ�&b�t$�D�+D�T2D�W�4	d�C��$/���`J-D�� �hŲF�)a��=v��U�V(��`�	u�O�:��1�j@�%�~݄��'(�}K�-#&q�p��yY.���'�\��̶w�@�v@�a�:i�'�8�A��5؎i��ƃ�.v,Y�'E��� e�4�&e3���*�b4��'�PŻ���A��(���#�,r�'~��k���UDܡ���J؈�x��3�'\Ti�����@��`�Ԇl�q��Tx�4	��HF`�a��9Y[�A����}yt�X�it�-�+�/Zc�ąȓOxy �	�7w� a�0���}�Յȓ��h�mI�"�Y��L^�لȓ|i.���
N�*�(�냉H�`�ȓ;��,�WDӴ
�h�e�u�N�D{2�O֐��U��
:#����(�����'����U�[�0�ehC�~�|���'bɑ
���Jݺ��K:u�P:�'�ۡ�9b��@AF�
m�,��'	� ��K���5i�8���'y�=P㏍�<xņM�\	��' 	��j��+�S�� ��e:D��렄>qv��@��K�3F,���?Q��;W��`$��ct� ��
�%E!��p�*d��+�*cz3"ꋾ�!���q�� *��:x�¼H�ס�!�DT/;�s�Üd�,T��ɐa�!�D�^��æ�B�x��͙��õj�!�D�(-.`q���ll���K��=!�� ����ӿi����To ~r�x�r��_�O����/�"�ړ�ڮ+� �h�'A��胩˱qyB���N���^���'��I3s�,=�ب%IB����'s:���7�p�e

�]0�	
�'Z�R��M+��M�T��$Wc�8�	�',ȉ!E�.����"cZ:m��'H:5p�	4����'�7g|0J����'��?9Z��S6E�t�`ѦH�o"Ѐ�S�n�<�Tm�%#��z�HKt��XEi�m�<��
۩s�za��n�8�1��`j�<�%)vZ�@#S*�	2���Rf�<�����ˬQ�pC�`����l�h�<�b�@�E�|� �F(L��kd�b�<��o
�"�
�A�	�L�r��U�<iɑrd��q)E���P��WyB�'��X�C�ˏsh0r �:��9�
�'AP��ĸ/Â� ��X�\0c
�'�QO%[d�i���OM���'�Px��0ո=ȡ�A�1VD�
�'+~]�s�U�JA85`@�
gKU�<1��16����1���?g���  O\x��Gx"�]1,^H]0�-J�x�bv�J��?Y	�'1Ѻ���;TP�	��^/� �
�'6�%:���-�����D�	N��i��'�0`��!كr�����أd��'p\l�׆ۦ/��a��X�64�`3�'���Z��(1Q2
��\�z��K>�����	:D,��&��	7����fC��N�i3( ڔ�ʸ;�\|�2M2U8�C�ɛW�v����̴�V�W��% �C�	�>�("$��JH̒W�N��~C�Ii6�Q��3I&Li1&�I2�*C�ɿ�4��eߺ7�2-�/�.�DB��%@	��0L���<�ARo��[�2�O��3ړ��@�t�ԩ�nP��:�撒o��}b��<��
�EFj�ё�C�t�hxh��6D���E�d����@�s!4��0�8D�`Q�a�m�P�B�(B pg�5D�|�$~��LY�
��F��	��m3D�H�㖎ZB5��DQ5��,D��[���VMBi��j��\�1+�<1��hOq�8����K�B��)�U�љNd┰T�'����LJ��J@�,[��s�Oȍ�!�dA1����4�E�S��B#Y�8�!��C2g<��)D�07��wl�(�!�$D�b��ܘT�?M0-�"LߢE�!�Zfˤ���&O�A�2�i��Ȥ_�!�DE�x����_�0�f����!��>�.��ՁP� /��a%�I�!�ޓ"6��Rg�J�&"NĠ�d�"��yr�I@ֈY��jS7*.�q'/�lW�C��<Z����Z-\�j�hd
�?y�C�I�E$d���C��EQ'��9I'TC�ɲoz}��c<��u�I%��C�I(G����P`�	3@����(�B�by�c�N@
^[9���/	?��$4����&A qK�1����*�����`1D���3L�;r��z���:��Q�U�0D�<
�m�;��8A��o��I5�/D�H��݋5&: j�
؆f�}�B�,D��A��(U�J��b �'y��I�%�)D�z%lO�}�(㡄98Hjy[E&D���F^, A�T���7�2E�f"D�� ���׊$(�����˖��pH�"O��J��f�d@Л�FP('"O ш*��:�a ���*�B�"O:Xc#�ZT0Q #���I�"O���!���<K�#�K�����"O���ć�d�����zz�hkd"OdYs�b�
N���7�
*\D�b"O�e�候	o\����NEz��V"O�=��cա}����#�C�T�Ѕȓ�h�$`�tw�c�c\y(Q�ȓf]Q�Q���,g�Us3�ćpp}�ȓj�*%c�A�Ԣ�2TH2��܄Ɠ�P4���?x6��u�P=������xҤ	�;o�-P����! Q�&���8�O�A���B<7�8�-O;&Z�J�"O�V���%��u�G5B���"O�1��m�0T�$H��*D#2v��x�"O�cq�� $���/�p@!�	�B!��8	2���Bh� p�@�*�^��}�'(2!ɚ��P���0q�ƬRu���e�Ov͠S�L"/lx�Ş]$��`$"OU��ΉY)0E;s�Z!nv�hS"O:h�2Fc0�I��Z>���"I�x�<��RQ���b��A7_���"�l�<@폻m"�-�?��9Hǭ�f�<��D V=���1f����^����&*rtss+�lt�89��<v_��Iy<��O�<w�a�vv�CQ�Y�<y0�J�zE1-C?. �H���o�<�wo�).��IC�9ki4�sf$�n�<�Vl�:X���r���C%��B�<�h�;R����MX):}*���D�<�/OP������]<����X@�<a�:
����Q?o�f�(a��|�<����q1���
O�WX��Qd�<��
߽J�b8A����G����cU_�<�H�2Z[��cv�ǍEx��C�(
T�<9��U7����'�
��듏P{�<� ��]�}20
�@ s �n�<�UA=K 29N��@�Ƀhb����U&�s�m��#� �Hӊ��&�T@�ȓ>}�!p^�6��hأ�V3^0H-��}-T�u��G��ʴ�](0�(��~��І�}���À�u�Ld��b� u�1�� ;t���d��$��ȓ%j�J(Я~�̅U/?r����K��Z��+K�BA�d#��m�p5�ȓ|�x�+6�ڗf���gܑ{h�m��XY���� ��J�0I$.M4FB���g�����^�t��T0�:���,�qDD3; �H�"�/Q����t�0�2���;�dX�Bܬ���ȓ���3�T<~��*� I�d�Y�ȓTÈLJ煐�x+��dRQ�J��dQ> �m�	1���1.Z?).��ȓ.\%{e֒G�����A'|��ȓeM��x�S���t-�63����"U���B!�f��û"$��"O��3	;��\S4d+wV}P"O�� q'�
'���6`֡	�:`y�"O� 	ㇾ�:IP��JJ讁H�"O�}2�f�(TI���JE4�T`)B"O��� �=T<��%#
�`�f�"O
eo�2)�2U�#b� �$19"O� ���S��(�@7�^.
��	p5"Ozl(��"p@�YP�[���4�"OHLX�С:��T#�0Ĺ0�"O�< Ba�-����O�+-�q)%"O���r	ArY�HI��y��'�ў"~���M��&�Ç�0B��m���yrf�T�+�%>�:��b� �yrd�.\�H�����Th�P��y�������K��	?"�ᑆ�y�HOv�=�vas)���Yw�4܇ȓj�2�1坩5* -�*W|a�чȓ>  #��Z�Xu�u��L>L|��ȓc�l �ʅ�{T1aqfպZmU��2zݱ���1.�
0�Üa�ن�W��d���o�ݠ&$��@��ȓ,��Qs��B�F:q�����ux$�ȓ�I�e�%x�4ؔ�0T>zy�ȓ[^p�R�
_��TCe\�k�ਆȓ35���+�v{6��tbמ5�ư��|���ʙ�DD�$jA:p֌�ȓ(=@M�����5'��	'	}�h�ȓ 6�0٥OQ�;q2�9a�
wԲ ��fF�}�,�GBF�3fS�
e�̈́�'��)s��X�F����ˉlY�I�ȓ����vD��>����BI��y��/�2�)��Ν?���ВaJ=qm��ȓs��Q*C�xL����;_4.1�ȓcH��)��P�@���?V*���c椘��i�&���b$6b��ȓ1#r��E�(S�������>� �ȓ�h`�똱]#���0#�Q_^�ȓ3�|I��1t$�T$0�v��?�N>����O�ށ�B��= �Ri�a�]�&|bD��'��@T�׺�"��!�1��m@�'�e���ҹa�͑k�_!h���'+Z�;1B�
}����o	�b��܂�'R�!��[�9�H!{s��=#�6lA�'�<yS�W�U �ϑ-���	�'=�=pU.�<J\j�G�'���/O��=Q�𤒀B렴�3���?
f���κ�!��<*=&��s���Q�HŒ}!!�)��1Ң��F���)���{!��uqL�0���8P�:�t���l�!򤏀j	�1�G�WM��zR��0�!�@;,�*�"���t�N���B"bj!�D
7�(�t�T�<�$�呟c?�X��(��3��1
���W�֩[/\�G"O�@�M�U�@��&B-�:G"O��b�i�@�4A�D%ۥ\z����"O��u-ӧ>�]��&
���""O� ��6V�}Ҕg_���u��"O���K�z*��g��sX)k�"O$JS�%?�~��Q�V����G"O꩐���jB�+��ҀY>x�_s�<�ӨG�."��0�7��!;�C@r�<��L��[x ���U�DI�j�<f��"rV�S��ϤV�F��!��d�<a�N�5Y��Y�V�@x���`�<�"#ɤ6�((Тg��G(@�� T�<y��h��q�V���v�)�䏉N�<��$Sj#�ũd����I@ I�<I���@����A�[�"�S�F�<��%R��ْ�!�1�^�c'LH~�<! ��1|f���.uc����hWx�<� ���@�N�(0nar�	�)����"Oxt����Hv���󨙢8!�Y��"O�Th��C:4�6Y����=B�~���"O����˞3S��%�Ґ&	2�҃�';�O��}��c]��@d��PPЅ*�*	 Q䵇ȓs4�)����(TJ��NPP���ȓC)�zw@�=ws��	����S���(l������@s��Is#�'1��ȓJ��������= �P��4��4��L"�K��`�2@�K�wl�9��]x$�S�\�Z[��s@HR77�蘖'$�'.�>�ɼTl@�+��T5},�8B��ۨB0B�I�F�ïA3��T �*�u��C�I7d~T��	4*B��Ð	�	|�����=?��)I�(�`���@ݏۢ�4@�v�<!Q�G�y��ș3���?Wf��h�<4�D�:u�az��::}:e�J�<�S�r���Fkm*ū�&z���	k���h���e���!­�+t���Y�!�D��a,��,Z�^�
���l�[�!�x��bC �95k&�`7��z�!��B�R��l(�j���P����/�!���Cv��ˇbB�)�"%��#��!�$�9�6y��E�
E��I���:#!��$�l]+���&=�`< �@'I�!�Ĭ-�V�i������i�􁆎�!򤞆1�(Ac�.Џ@UU���.k!�dҼmI�<�CØ����0IK�zP�y�ቹf��Xq�[��0;@�۱plB�IL�,`��+e\$y$�W�f{PB䉒\|��D��"���(q��D�|\��9L|a���/s�����^ j�
���&��t�/�]�]x���iu��ȓ	X2\X��\���[@��I5�\��U����j�#J��ATO��NUd�ȓ#���PP��k8LB��ֶD�ȓk���;��Y���qR��G���ȓk�c󌝯���Y�����ȓ�@U*v���h�x@�ڃ4�F��m���GkO�#�r��C���,]����.F�5ё
��N�:䙃�L�h�����l�U�dW8��� 6x���v�R!��@�/|b���ۦ4�v|��u8X� ���R�q�R��z��|�ȓ="r����@�So�`:�Ɵ�����	r�V��R%�X%����HsV��7��B���9�S, �ȅȓd�.���ؔ;�x���>I�`��?�PqaT.�1w4�$q��Ñ��Y��Ir~�EQ"lR^p�,X�AN�0	A��y��K�b��Z�&���y�,�&�yb�N�u��sc)� t������y�
��p�4y@g� t�b�)N��y��V/z�hب��!e�D81��Ǒ�yr�.2��u��B9`��D2�Z��yR/W<r��Yc$�&ֈq�!�L��hO4���Q- :X90RML�͛Cݳ"X!�$U�P���7�aI|���`�6m�!�d@�oν�"g�/nX��/˞n�!�Dٴ׮��Z,P��o5F�!��R�2̰��$R�K�ХM�a�!�$���$�W�='P]$̓-&�!�dG�-��J��T&x���mȒc!�Ē�����4kW�	�,!l��M_!�� ���J|,If�@�D�BE+�"O@�I*H���Dx�-�{/�Ё"OV�+�@��[� ����A�"��Q��'����p��#?<x9�`!`L�f�0D��Q�.Է������$�Ӂ'3D�(�E��}�2� ��9��2��>D�@C��=OR�8�Ul\$6D�e��;D��i���ĢE�;4�M{Ʀ7D�`t��Y�q�Y(`��\/btVC��)L���G�ւz:�|ڇa	<��D�O<�qu�37՜: P�I��� }(��ȓh�����X�h�Ƒx§P`zl��f���6�K�<�:	��f��m؄���*�
�d
�:O2D��T�P�ȓr,M�ҏ_���hH�e@�T�ra�ȓ7�� 05�	��`T	K`�Q��.����a�o'��(�Q%Ύ-��IU~�nQ�c&D���	��G�F�yBK D��Y[@�3�����X��yb/Չh1(E�V΂(����aGͩ�y�(��HrB�"� �� �y"ψ3
-:��sM,pJ1�v���y��=��rB!�)n�zX8�n� �y���CR��AEO6Tf��
��y�J_'�.YjWD�`u��#�LZ��yB���#44�� P*/x��F�X�y�Y�t�4�1�G�( �Ÿ�iΉ�y���-n<	�����u�~�I�*B��yb( "f���'֕#�tQ7Jր�y��H0o����Ęu01jUoز�yB��/9���+J$<�v�b��	��yB,�#CVR����,�R%�����yH�2sn���N �,��)w��5�y�H��J�q!.N�V��6o	�y�cАa��ȶ�4��q�geY�y����m�̑�d�B"Z�����b ��y��?�D4��+��L��l
&GR�y��ĺ$ ��Ɔ�M�����"���yB,
%2Z,��0G"FD��Q��(�y� ڧAL�geO�p�l���JA��y�`S=QV!�F�<[YHq�cGW�y�+��*uL������J�k���y��f,Ԋ0�D���m����y F1�R�#�[�v��1��`Ƣ�y�@-�Vy[c7vҶ1�C���y�@���n��ȋ�E���2үC:�yB���c@��"��-�M��@ԋ�y�O��H����"�$�����y�g�;p��ӕ�Ы�yʆ���yRjL�V��$�P�Ѵv�򴀘9�y2Ύ�d���aBJ�
`�d*d�[ �yR�I>���1�-4�jaH���ybaT\|��\)%3J8��ϋ�y2�]��CJ�!�Ra�@���y�o��4z
�PQI� <�y� U�y��O�i�pг�0f�`�����y��P�W���%,Y���ɸV��/�yh�w���	�"��|��u*��<�y"	m�t5�)H��ȣ��8�y���Z �mY���P��jt�N��y�O�r�(��,[�Ȏ��nU.�y��Uz����T�+0<���T�yҋZ�����
]S@*
5���yR��7Jx� ��ĭG�4�B���!�y
� ƈ�B�{׾L蒧�)o��q"O��U�I�@�AF ljС�"O�����W�r ��Xr1�E�T"O�i�A�V�Lݜ���۸N.�"O� u�B��C@[�V���d"O���l�5�z<c��Y&L�\�Z�"O(�"jG(xf8H�bg�����"Ov�@OΞ��LbR�
�W��bP"OfJ4�&%���Y��\7�|A�"O$0"�_"���i�mӃc*!�"O�+C�/��!Ǐ�!w�{�"O��t�P�{�ؐ�&��;l��y�"OJ��%0<�J�q'ђY��i`"O����͓8�0���WO�8! "O����l�E?��C�k�
p$�=�"O<0 �h�c�@��F��UA8��"O��2�/�b��aP��>���F"O.�3��_�2ڼ%ےgO\��)�"O$\ďZ��䓣�ΌRE��
7"O�J'E_.��0�F5XXT�Q"OD*$.��%s�9Hà��D�i"Ol	��?1W�LK�.U&nG�l�"O*PK���&8� #��5J�}�B"Ozl�2�eM:mr�A�B�LI�E"OP�z�̎/�]ۧ햗I�2��r"O�a�w�]�\Z0:�ș#M�Q��"O⹋����@("l�tB��b�"O��)!U��������p�FT*�"O �f���Y�<;
�� }F"O��AŌ� D˞�{�/F��N�0�"O������3"�1/����5$N!�D��3��"�c��Ma<�`�l"ac!��V��P�MS=3�k	Z!��_�,�b�ȓ�ˍ9�<q��
�sF!�D 5D,�ib�Hs�ХK� T|�!�$�%[� �$G�`ȑsO�?(V!��c��C&>}A�h�`��I����k*䒀�I$ۚի�F�>-�%�ȓ|�<`�gG�i+Z}KT�U`(�ȓh���ǫl5�г�*M�۴��ȓ*������̯v�:x3�M�d��v� Xȓ�An��i�.K�FD�͇��D�yV�T�*pi!��O��ȓy+���fa��k�Z`	a�p����c+r5��N��B�&$р�ŗC>0�ȓĴBQ��#k�]ے炚;�,������@=)�\C��Z_S�a�ȓn$0�E�lT��!P�H�.��ȓa�9���C?N8Ti`2���9�&h�ȓhf�p�O��Mho�$3*}�	�'OZ\#�/�8�mH�O�}Gx9	�'0�� ���*#�Ř��û]��A�	�'�>9�Շ���~da���P��T1�'�(td@26)�bc^�D�
Y��'��� �n�"i�Fa����L{���'�z���  �X�e��&I����'dHx�QH<yb@�A��Dh�=Z�'E�Y4�L��݁��:2���
�'ʠM�f�.E*�*2�̜6����	�'j������9J��б ����c�'��k�mطf�$cQ'T�m�\i��'8% ��T>C�x�r�!A)n�~h�'�4+N:xZ�R�� �q�'��FmI6$E�� ��X�R��� *���m�S��$c��ޏ44+�"O�4���@�e:Vi�G�X�VY���s"O�0��W�a隸1�H�>�S"O<HA� X�2"v�Cf�@�/��-��"O0p@�9`M���W
9봸6"O����Dց�ܭ�!jJ�Q�<YR"O�6��V0��qaH��`Zw"O ) Ɗp4 ٦��9q�Z�;"Op�*',�$W�"����S��@�8�"Ov)��W�Z���Ҁqz�hS�"O��إ$����W���=����"O�Q�񌓢P�lP�f��n�`��"O�p�K�J[�W��X~��j��q�<�� �4:����힌1.�q�ABT�<P F�P�$�;c ��J�����`�V�<��`��@�����(�mE���WV�<�,�o��Y��O�T��rc�K�<i��	#H 9�N[�w�pC�H�<�h[$PB/ٴa�9�VGH�<�Ӆ�.�ڄ�bG;0$�� F�F�<	��H��@��歃���)�,Lx�<�Go��q'F�"2��#"A��	�p�<Q�@@�N��y��.Η3�(�05�i�<91	�0 ��$Y��.cr��a�Zo�<����U=R��~-�Pxq@�e�<qč9H}(I��	�B.�)(p'�`�< �	ɒ��1lȖA�m�Sg�T�<!�$W`�(�sFF�s��9�3��N�<�̞�S��Ȣb@ۦ*�h���@B�<����8���+�%��9�!��<!0�)YC����W"!uup�K�`�<IP��7�f�c)H*6��H��_�<�RF�g���!��&�>��`)[Z�<i����b�l��Ǌ#���[WU�<!� �;|�@u�cl�n�+X�US�B�ɤ"ݔ���^
ME�`�ҋ�{�B�I�1��� �]�V6*�5�A#J��C�9!4
m�D
6��1'�B,�C�I�O?��"�©t&�T��m� ;!�C�	2��9UL�� ʀ�C��~+b��G��\�`G
+#@B�ɼd ��%A{NĐ�I"NB�I��n�1%ۣ��ĉanZ=E"C�I&�@����T�D��M]���C�1d~uc�#F0T���".�H'�B�I� �9�s�?*Rp����"�B�I�U*�as�� 2����E�
~��C�g��Ti�؋YJ��%��1��C��(j�!p#��+4̆�t�[�2B�B�ɇOKFQp��D�OTH	Q	FP�zB�I�c�fmx$�4@(�v��\FB�ɵGP�3�Kr�Tɲ���1%�R6-��xG{��)�-��X�J�	�1aI«L�!�:E�SC� h�b`��͈�\�1O����B���)�E�q���B*vax��IM�~5;���&?	~�	� w�(B䉋v?Z��e,|�`������lN��hO>��i�l�jA�q�3@@\̀��4D���c*4��!k���|��1 T�2�D����=�~�l��_��)���(2B���EAb�<������� M��3��Zg�UZ��p=��Yf�iPˈ�g� `8B[�<�4B/�QEHӵo��C��W�<�u�-8��1��2nF@��'�Q�'P�?� �DkUB�sچ����I�
���"O��Pf��j� (l��W�� au�9D����Ʌ�t�Er��ɼ@-�@1�9<O�"<�Q쒳B���G�M�.�d�dF]i�<���E�/Œ%�P��#'h������c��}���Of�5ru%�)E�4���M��Ј@2�'��� �>R�|�CV�R<��-�ĥ��0>����Ĝ��%��� %U]Ѓg��!��S7uj�ۓh2k/�\��C���x��	�&�y�Å�9&"�Z�+�	*B��}i���y�F���A�,�썁��<�$�B{��(� q���3=����7���f�d�Y��'����ue�ozH�Ј�c����r�8�䘥c��z�%�@m~Y��Ů]xna��.����'
ў�Oq���P�o�X�(c�٫Gc*d���C�<Y􉗺>�HAIS�	�fp�1V��B��0=E���p�(�'�;�H4p��~�<��|]�53P���L��Ow�'F�y���!��e1D�?ջ�L����<���B=N;��9A�����!�N��p1�<�ƓR=�5I�B�4�87��l̨���D����3A�0U:R�ݼ#(���zy��Qs�:2TtscgǸk����ȓu{-y����y�����ֲ#eNM��KT�𳦆�4,^��6�:��"O& ��
=K��3� �<d��Z6�'�Q���@�P��e[�L��pvx��q$<D�hAA��\���Ȧ� QI�6D�`�Ā7Z�( 9�)��D�xe�D4D���� ��$:e�;x��%0D�xR���-"�u���"�*CA-D���"K�`Ru*cB%eƨH�4	,D�D �,ȆjϺ���Btd��ʀ�+D�ځ�0@���0���	 К1�!)D���Wk� ʄ0�"J��`BJU���(D�\ʤ� �T��BS��*ū��*D���E⓭{�p��"�ȝz�L�j#)&D���e	Ǵ4L,�Y�'�c�ت4�6D��1��Q1JtD2EA7H�Ta���)D�X۳��&�v�; A7r� �%�O���mn-@%	�2֭�B��B�I��hz� ���ʃK��b+�C�08�.騳��wF��H���4��C�I/]����`D�(`��	uh�=D�C�(,�B y�hS�v8�4���� �C�ɰc�D�#�kޙ7ݔ�i�*�1�O>�=�~QE�1w-H-���Аt��D�i�<�$��0{�����?4b��"���d�<��O�O����ږ2<�"p]b�<�t"H<pr:�	��\r>�4P)$��<i� �;𘭰��X7H֞9�2�n�<�F�=$bD��T�2r8��(FUn�<���"/�L��w�['\�:�j��f?����韞e��#^���h�	�<c�<Q��"O��H�,�����7m�<��w"OR���5�hS��\	|�~�S2�d;�S�T�O
-ce��-6.�x4�Y�R�`��9O(���D�6�w�ʹX�F�E���S��f�i�1O���gyR�~n������^3#�Qk��D)u'hB�ɧ ��0Fʌ ����5HA�4B���c�GA668��򮀁E�hB�I$,R] �
OsZhLڅi^7^� ��b��3}J|�O:�rR� N��c�����@"OhX�6 A&X�~�S�G�d���p"O� ��l�/_�<D{�N�?�(x�6S���M+M>�M|z�'�=��FH&S��rF�;""����'n��a��Sf��y����9k�y�#?�����+�� t@��0�@\�`|4�k��Ie���*�3*�j5���ڮv��<��+G`��~�d��&�)ڧS}",kÁ��05�悀yI���&`D���¦E�q��D�[�x&�T[	�'+��6>-
�����a���A����I,����H
�[�˧G���ȓ�@���NG樀s%@�&~�Ȥ��	Ϧ��>�]2:
�12@�5p��H�r]�<Ya�mj Y��O0v�����LW�	M���O Er�>.!p��5J=����yr�'H@ЅΙ g<\�D�R/y��h��'6x��%-.�H�@�F��tQ�'6��YAkF��j`B�)
��d$$��E#2fJk��Wh,(���1D�dAEn��I�j蘤���{s�0D��8a�~b��	�kSc�}Y F;D��B4BG�%�
L`h�\�����9�$$�Op�2#�F�)��AtbA'P��S��'��$C�t,�zZ18��u�_3�n��*x6\���:G��3a���l�v���, jDz���K���s�p�ȓ�di�RÌ�=�đx���v�$�E{���n�:8��Tsg�X���C���d6�O��g-Y"E>D�`Emצ2Ո]r�|���2���'6p�p��AG���*�{����X6 �H ��|�U��'4~b|��f�����O^��G�[v��X�0"�'����� T�<)`�EU~��@��L�!�#$u�<i���#7s
��e��7Hh���Bk���'� ��#b�C�Y+f�L%1�'���1�e�70܊�oN��d�i,Or�=�}��x\~����q"m���x,�ȓW��8��(D�4	��S7)�H�y�xB���$PQ�8�#���]�������2�Li{��ٟ(��	�<��́QXX���R�ʍ��.�Y?��by��#�{biP<Ѹ'���rbL:������=��p
Ó��'��A�K�z� ��0�����Θ	�ybi��><�4��	G?%q"]@�mV���Dk�<c���|Z�',ⰀĢ�=A`6ܛ!��s�ļq����p<�s�G-�l��$)�QQ4Md,�Y�IJ���	��0k7�[��� �	�&911)D��@ -i�P݉TID	N��&�$��c̓5���ɀ P.����#�*�D�	"D�p��`�@~�5���|n�*�(�ch<���� X��H��R�0�T`ƜI�<�1��!,���K�	�"ѓ`��i�<�ׂ�� ��:��\�b�����Zc�<����(m���r�c<@x������H�<��Fޒ6V���BP"3����k�<a�A�8�NM��ɠe
L����]�<�7��P�@�2��[�X9 U�<�Ԉ���X��@�(��t��O�<!��Q�1�����S#cvŨ�`�<Yt$��|�V�� 	�88�-�\�<�����^OV� � � 	�t���)�P�<��I�Ǫ�j �;./L}9A�O�<�ňp���nI�PZ=�p�OO�<���\�kwB��a�G� �DM�V�<���Ŀ`u�u�􋜴1.� Q��R�<I1o���nİp��X0��P�<�tHՂjN�l�b�rpF*�J�<� �U�U�ׇUN�Yg�\�T,��@"O�#�lϩnZ�!&(9P����A"O�h���[�a�� ��Y�d�`�"OV\)����#�ly�@���i2!"O�Q)��Š�tɹVo�&X�a��"O8<�_8���+?��*5�X�!�d�:{S�h��+X��j(4�ҠM�!�Ĝ�me�L��HF�/�j�J&a��!�D;G^I�j֊;�^)h����!�F�m����L�Є��7&!�DQ�x�X�Ň��,���*q!�$��~VZ�K���F�����md!�$Y�P4�� 
<pڀ̱��а'\!� x��P�2�$Q�]J�b��O!�d�p�D�r�/�<%�lL�6^4O/!�$���]PJ�O�½k0N)!�$M6x�1A��	m�m[�#G�A!�T2>�Y@U.S�H!P�"֘d!�$B2�x1��!F�J�
7��
D!�0���m��lxT�����!���@�� b@�˒-kP�Ҹ�!�ēu�F�{e�E]2�cB� �"2!�Dד=|V��v`�'SA�@�68!��_�@<��m�.:�rG��*��U���a~��R�PJ1e0�Pq���+&F�B䉁xX�Ԉ�l^:+�֤�r�18�B�ɊH6���ȦM�P�+GbW7 �C�	���]�p �h�L@�T�fB�I^���!��[�k,��UJ�kDB��	
��F��:A�v�"��O�kx\B�ɒa)x,�g,�H���u��m��C�I�Y��\A��N�Z!�0���"�C�I�Hs ��r&�7��1xR�A�dC�VP���|�v���G��8�$C���z8R ѰUX�#�Kk�B� QX�CrNǼ	�u�eɌW��B�	>+ݪ��˔~H���JƮ5��B��d��@��lרXB"�b���F��C�I�4eڝj3�Ň�8��q&�W��B��.o��o�+t��0/ i�C�	�o<H"fC�xZ�9�a��p�
C�>����BN
��v�μa�C�I�7bݻt%]�6�޹Z��MT�C䉬d�dH�&d˜y��	 b���b
�C��)P�v�@q&�/L�,�$P1T#HC�I�S�lh%n��f~n, Wie�ZC�	�>kX-��Kh�\*�
X%doZC�ɡ�H��0��2T�N�cjY�D�&C�	5'�0�� K|��g�T<E~vB�	�X[ ����X-AD6����	��XB�	�u6L���B�
�Fc@��}a�B�I^�����^/{�bU(c�#,?nB��0oy���N/jD9�ҍ�.��B�I��T����D
��H�gP9ɦC䉑{�TB�Y1��a�ԈN���C�ɍ-��}�FnU0bѸ�1 �9)��C䉻{��42H\�>��q��윖D�@B䉋420��WJ�����'-��^HB�1xO���.R"D��٤k�+�B�(6�qxwi������u�&C�	�aYKg�@S����^��B�YN��V�%��SgÜHpB�Ir��QK�菪r%����F��\�B�	�Q�i����0�{Bi˞}�"C�)� ��;�위L�V0`/n+��I�"O��3�HP�����ψ,�Hك%"O������%�@�b�)P�l9�"O6���#��G�콨���9g!��e"O�	�N�5d��!�k��01"O������(��]��g�/)v4ѡ"Oh�&��-d���委:x���"Ot�
0�Û5>p�I�ews�i5"O�QzDk�u�l�D��H1z53g"O�xy#×�$�P|@�FR�x�E�s"O��ԣQ*0��yj�%K2.AIx�"O  � �E�a�>ib�.�#��4�p"Oh �&F�,�ћ&�0�n���"Ox�J��N�Y��׶;U�pb"O*�f �"R���׿+;�͑B"O����O/�t0�D��g2p�0�"OD����=-���cHm>��� "O�QaX?s^nm[��Ńe\��A"O $�����i�	P�cg*a�"OH��VB����ER&b�FA~0r"O�W�&�&0����^��dEx�<Y���6Be��R�t+��i�c�\�<�$�$J�U[E��[�ȁD��^�<a�e�.y�˳nR$]3� �U�<yE�D����3��8�z�cA�N�<���,h/@ڤL�:�<�0"��E�<��z�K2~�PDё�����=��'�Jb�F��Dӂ��
S> ڶ�Q�'�
\I�BQ2-�и�W+	+$d��C
�'�"ܹ6B^�(�>8�%돏Bd�	�'�m��I@�K�Ju�e�TJ:Ȝ���+� ���4�)�'+�8*��ǐs�̙�$9=Y�	�'Ҽ͈#M��n0^ ��H�0o���'�|��b�GЂ}��I����:��͚��P��eٽOL����M�zZ��ۄ�N
��UŦ]�2�a#�2��P�(Аx�n�5��3��M�)�PQ� �>���О7G�  R��֭�W�b��ic��ħU(Q���/c�qB�^�,@���6M�fM���J%
�2��p�-G>Qz��*a�=�v�<A>��$S�ul�����H��I�D86D�
O�ji�dO�$t���<I���\d&�'~���ST�]4xތ"Ͱ����'�<G �Y���*fG�˰On�<	2�G-��a�b!�<�؁�ԓ!�r�biN(2ӧ����O�x��#�VF����Da~)�R9Gb�����^̜h$�'�4�`E�w%2 �fc�P�$�����A4��� �!5��p�C9U�Qm�)_�ӝ/>����ϛX�1�BM]+RT.���K�v�Pm��K�^�\D�ؼv�!h�k@�j�P8�����D_���a_�"�T�h�"�� ˓^쵂uK0}ޔ`{%	��H��Dy�d[�R����p�O��@#l@�ua�.U|p�qF� #f~�Y�b��Y ���לf�џp���J�:{�@� �&)0�/�x����#�г$ҧ��|$y�� y�����U�8�Cꉩ3z�;�=C�n�p��3�O��#�T�S����톽$���[��OP���,�%m0�=a%�_�_���j�/��L�cޒ��I  u�8�!�n���ܐ�H^	s�a}2k�=�"�Ζ�q���.d_��Xcb�6=` ��'�F��f�7"�p��&§���zm�T�w�Y�FT��M�1	;�O��+!�>S��T��'P���q���M@�Ь1  ľ|�4 7%P��ظ)d�͘V��׀M�qU�Ȁ���YM�x���J��i��Γ,�⹰�䌶o>�ɇ;K�ܲ�"S��� �82�12W����1 *D�P
z!{�G�8�^��0"N��D���]�r�Qg(���Q���#;b<㕏�u����OEa���F3Y�f�!gK�哎�t��CH��E:'�F1Q &i���l�zr̔�MP��sԅ�<�B^�)��A2��S�tTZ�36bY+���2j]'T�>=jw��O�)�b�ު-��ir�K�b��O�<qd�θc������<���#��K�|�t����"Zt�K��ܴG��Б�(���4�Ä7<�xS�,4H��Q�� �M���Fj TH�%F�X8,�Oz~Q2�l�$y��I�`���6©�d&6�\D��(��49a]8J}tY�O8�3�$p�4��eI��LC���!,� ܸ����p��͇�V���AGeal'(��3�V-S����gď:�Ly���=3�f�z)-zH�O�Œ�j��ۀ ���,�q����ڊaZ8 �A�'ﲵ�"
FnX��	�@�h·�D-Um&����bҺ [��A�xpX���O�	'xqZ���D"@�J�����5,x5`�"��qO8b�(�q4	�➷��I٠K�"��� �O[�Mk5�y�6qA�e��4Ԡ\��':����Yx�AT=�:�����ޔ�է#;X���c>���1<�-�+��2E�9�	�&b4��"O��Y��E�?�.(ٳ��QlƵr��DK^��#�=�EK�](R�����O�'�,E*2�Q?v
����(=/&�9Z��T� ez��ӟ9��	��R$�B���A�y�,ݩc(>�Oz�y�e�[ΈH��_-W�jMkA�	�h` S�]3~��O2���GX�'D|�Qϊ'�ȇ�ǖ]�m��7D��:�ǋ8$l���'n�d�%�pIɧ�8jt`׮^�N�1���2�h4"Ob�Y+�cΔ�Ç��탵�������ÓH٪x�ы��E0��(��P�ȓ_�dz�&� ���J��%	�p�ȓl�<iBw�˟V)����MG����ȓl,�`� �V+غѢ�&�D[ܡ����eY0&߾ ����{D�t��'.��P��H�&HN�ڢC��`�ޤ�'�)!���	4���� n��-��oSS(�HG��'R���؛c3P�;�	�c	�}��'�"�F�C-[��X��"
,\{���4�`i�5Q��p>�4�.�����H��e`8hX�B��<6�ٙ���0O��X�DѱU���1���J)����"O���`���� !h��I+r�!R��Υ��8����������MK�×���?i"Իf"ON�kb(��!�w�|��q�ž �fɁ`�2~���̚��T�E�'�ƅs��oV�q ���d��h �\P0+ƃ)�?٥�.[��Ӥ_r�!xЩO�]�V��rś?H]����]�"�:�Y�7�(���޹8�P��+G��&�hQXe�'m6MP���vvx��'q���9Ca_ s���s���%6��9�ȓ]��+E{h�C�A��T��E ��B(�ǖ>E��U`ʳY��ͧy�aj>�5`�D��8�M5	90��k!E<](`�K���zRA�M �£�ym�E#P���%z,��D�N�fL���4x h�!G�0��Oo�QS���7'x,�J�hq@���!�e	 �C(Ԃ��5ғU����q@�O֒6M@<I0�� 
��u!��`�zfi����yңn_��Ms `ZY� q�%@ԽL}����R�(���7��?PN�� ��P��Z��
8?v�6-�(TY�a�j���M�R.�?�Xe �j�?�9��Yq��"���h֋m��Y���yJ�J0 �X��(�����$Ϣ	�3ʓg{�]���׉x3d̊D�ZB�Z�[և[�j����ǯNn��0�4����{9�$�A�P�S���$��}8�KP�n�р#	:J��#r�ڄV.���ɢs�|ه�4����U�[?Q�<��U�#:�׻i�m�Wj��D2���	'y�v���+�x��1�#�*D��亡�G�G�c�4 0��1��#=i�\=t�H���O�AX�E���i@;SC<a:B���S���&�I��UĒ�&�h���h.���!��O2H9rEH6��hRo�03yNI�iE�)af�I��%͓#Kfl�R�*��×+��O
�����9AD$؁�J
x��@���]+,��C4D%���g�'R�p�F���N�'%���¨OXHm�5w�6!��Ě�'������E�4U��ǝ\BL����-U.��"��)&v��ϓW&��rEO�@F���'g\/T��� n_�(O�!ɢ��.*�>i�'F�4cb�姟����ߚ8C�DRK�L����ɗvֆ�K�So�̔�N��q�<tђ�a@�U�L4�Ј(W��,k<��S��?ɑ�31�J�Ȣ�Q�{����� �}�<���(yB�8���]�ށ4j�W?�3�D�fO"���.4LO(�
��l%:X� Ks�YQ�'#��K�P�����в:�|`!�/���(%D�ao��7G- bH�v[�LP��1ړG@�����-ҧb�bI��Ι#q���Y���yY���ȓG�2����b�锃�)�,����Ř���2m~\iae�@z�8��0�@c�CI"�(V��U���h�[`/Z/F�x����El�a��:9 @� �нXe���gH�+�!�$�*e��
���A� �U
S�6�!�նG#��c6j׾ׂ9��@�t!�� �d`��F? 5�=l���"O��ZS+\09�p�BB�	^��E�s"O���9�h*v�²}j� �$"O��{u�]���5��h_J��"OYr�������d@���(�"O̐s&`�M�$p{a��N��3"O ��bI��]9ٖo^h�t��"O�	�
(x��P`�
�G��=xV"O| !�Ǐ  �J�R���0�@�bf"O*a��˷%��07�ސ��p"�&D�\
�O�<|����vB��∵@g%D���b�J	HF|q�g�?i�x �j5D� q�,Q��PIWH��v)�X A3D�� ��L.K���2�A�(_l�|AR�0D��u�� ]�hx�/@2L�d�@,D�4�1(r��ػ�J�2S\��pE�*D�L�� YH�R�����@!B̸��"D�8��*P
Y����}�z�K@l D�@!Gk҂D6�8��;$�d����!D��kL��q;э�Z.��A� (D�t��7�*A��3'L�� )D��I��H*p8q"'FʳBZ��3D�ܪ�T� W����M)?[<D�a.D��DD�m�0�3b�7M�}��0D��҃Mݎ\^�×g��&zJ�a4�1D�tX������0�#ʵ <6� �-D�<9�停~�L��%�^����p�7D��qC��[��"G+ͺ!���5D��`� �+B.�%)�{�Α CH<D�����[�Wi"��� �{�D��e8D�D��#��r!q*�v�(���%9D��AcQ m�l�)@��^���a� 0D��0��&o�ؒ��M�q8���Q�1D�p��l]
�r8`��5�i g�1D���C��8%� �9��<h��R�,D��.�ZQ+"c֑X�`�����0~3|C�I3|@��UK~M0-�*V~"C�)[��i��ў!#�p( �W�PC�I�?:�١#X���E�E�%r�C�Ƀ3!f0R�I�8H��Ĩp E�b	�C�	�Yd�#�G��y��F2C䉓�Z��/���A� A]�OPHC䉪���+'�U�C-
ss�Zp\C�Ɉh�PL�A��pRIq%�~�`C�	#;�N��O���,mH��SB�IFlP�$�@#����D&�C�	-z*Q�勀���Ԃ#�ֲO��C�-��p�*� Y(aq" �6�nC�	�'l"��� @>�x'$WJ�^C�	�uY D�GGB#Z��Ç��b �C���F�Kd ׋?��x��Q:"r�C��=�pM��V`�!;�AZ��C�	�E���GbФE�,<�� �lMB�ɾ"1ph���T:(�2i7#��B䉞K������n��D�Ez�B��x��=ig��	9E
��ul�g��C�I4BPƴ�E'��W���[�I\��C�IjؚMPBFn�EHƨ1 *B�ɧS����L�;(U
]�ǢQ/}�RB�	B�L�C���8,����l�B�I	_<�	
g@�pC1�ʤG�vB�Q����1�C-ɨ ��I��B�I�:N5B�� �l2��P�zB�ɒa��d��g��@:��57&B�)�  ��Ţ��"
���	�=2d��"O�!�V�H�:y�(�nM�F�S�"O��+A�"A��J#.ҨY�RY*�"O(U�2`_�m��005�ʲ%�P�xW"O�ԙA�5��5�BKP+�h0� "O��B�F_\��W�C#��("OV�b���>�(ТA*
�8<РYR"O���aϖu�:�¦�E4تg"O�=��$@�uz��R���v��% "O��@v([�=)h���G�y�"O\�ks_$���!���^���(B"O¹	0���{�d8��(*�jP�d"Onqؕ��C�Jy���23��T�W"O>� 0@�[,�;�Px�uS�"ON,R7(��TT<q�D��B��H$"ON��ӈI�wE�F��H֛��=D�H��lL�|E�\Z����Ê�ya�,D� +�;�њ�K��F<�h�	+D�4�D�*R�B��;HS�eVl&D��Z�eM�.)@ �c��s�αz�)6D�<B�IʞF}�����7��hî(D����,n<E�ࠑn�h<x�G(D�`8v���
��� 3A¡?7l��O'D���`� �w���EA�~@�Z�	%D��CU� 4VF�3�^�6��+VF"D�[�jK#9��Q�5�]�k;�9!Ġ7D��v�í:����V>=Ւ:��4D� ��&P�F�I1%?n;�0���0D����(�+L��*Ɲ�5O�]��/D�$S�Ĕ�l�i�#�o���RtN-D�P@6 �[U p"��Ѩ��M�'*D�DP���|��jY>�} �?D��[���hh� ��/$t4YZ�=D��#J��[�r%��_)uvl!r�?D�8�5#����`rDB˦VJ��f	<D���®ա���ۀ�	3N	���pJ;D��ZDB�d0����ld��7D����B�	 ��p�T��]�t��'8D� �o}����v�J��4D�<i%�J
:�2ySk{��D�<�$�ͭxV.���C�Z
�$�SE�W���1+ș�a}"#V1 �i�DK��D�hX�O҄L5.��ΐ(
1C�	23�l����b�6���CB�h���<��H��0�b�8��.�'/࠶�g6*�GmW���L����ls�,�$	\���l��vz�i�G	L7CĆaҠEJ^���O,L��ޙ�t������k�"OD=��Q�>ؐ�+%[���G�O��TA�7Z�&�Bӓ8���1��\����&��/�^M��	�x_���mϬ-q���N�cy�E����=B�衵"O��[3BȐeļ���
�(�4-!��I�@k�֙H��8���i�<���e��q�l��!�ĉ�#(��C���<j�z,���;?��P���<!�jЃ��>E���$N� (�B��&��-����7;�ن�l���1��M�7(c��K3&)����6m����"_���Ă�[�Ӄ!	%'������'�a}O�:J*I@f�ۀL�������
^@i6A��#C�I�8;��ۄ$!!�&q;�O�=f���L��lS�usrp���O$y+������-&-"m�ӊ��M�\�k�
�-X!���Im�80c!�!4Ƹ�w�\�w~�������^�qd��Q H2��;�y�#ީBH��tm���F@��L�&�y�AK2:�� #�$f.tQ��>�0�COQ6�Aj�'�����eYy��Dx�k�9��5�S��J�j�Z7�j؞�X )܏Y�yq57Op����Q�5���`���'c��L�GY,M	��Xd�a|�����"âB&�1rf��5޸'�%�A,y8RH�D��1	bA�0>���g�? �tñ#5h�*eR��/vT��g"O$�A$C��=����(�*n�s4
�C>�4�sN���&/�3B�0�i�I�"�y�'��Jh(6*	R��7�Ը�yb�S�>
2Xm3|-�C��a�X@BdG��/7�!Ӏ��<�&*��'Bz T�R�	�1�@U�j�/�)SG}0~�����~���k��^ ��SŃѕ��8��D!se(�#��<I6}i�(1U�F"�`�P�5]�wQ�p�pCЃA�=�HA!�+�j�-j�*���e[�2��p>�
�iC�H4�j���@P�h��N.D���%�C��b��Q�Щv|�+���X'4��h����
!�;P-�а5�	E߼��=U
��3w�Woz���U�<qbI��lJX囐��Jh��&�%� �ʖ�վx��녅bF��өmH����!G�1k�ۆ�)DB�]R�b%�OR�#"aƘK��ԦW�r0�)P��[-������?�QG��.����ν��' z�'Q&����Ӟ8�*�&>�8�C/􀨨qG�p�xp�4:D�t�r�ΣA�+M��d|h�6"9?)w�ڏ���H>E���p^�鬘ecЋ�-B�j�RC�I�o��IJT㑜N��8�@�%dr�b ��28�axR�	!B͋��,@���q���y����4>�k1杁4�H�G�֙�y�M�.0�ĩ��֢r�@�d"Y��y�*M<�H�;5l��t��H�I�7�yE�+1�`�b-�=1�� �e��yr��V��[G� �8�E��y� t�� ��jO�x1JB�\HP�`,�H��~�P�z�&�����bPȽ{7 _��y�aށA�r�fn�4Q�� ��ǿ�M3��s��ř�Sb�t'fQ??>䰒$�)ۢ���8�(��4���)��O�1m�eI� 2ts�\BRlײ �!��4!��(�$H)w�Ё��h�qO�а���6pЪю�	�|tN�s��'<���`�Z�!���t9�A(ٛ ��}�"؜抬!�����`�O�x�OOrFx���0x,m@ЩҾ<�������0>�V����hK��x�S3��#�}y��ݞ�y!*�:0�}`QW���&�k��8doI:%Z�p��;�	o��aC�N�h�qF�T���_�|
7�D�^VJ�Y����Fw�H���Xm�<A7+K�t����<^F�H�&�v��|)��@(����e��d�I W���|���'D�t��\E�R 8���8d�̦5���2d��/Q6*�3�'�	H�딌K���C�nQ�c��9!gI��I��T{�	I�W��yF�w��a�	�6�����d��YGi����-�R�@A@�8lֽAƂS/!^^"=��B�p.F��d|�ҩyf�,'TPh�Zw�½d��V~P1 �%CSnݹ�47����
ϫ'n@����:v�I*=��>a����"\�#'(V~��ز�mm�P�p��J�~�՚ڴ3�"U;Ci����)�❡u9�k�6��u&��ľQ ����fSޱ��'f�Q8al�fQ:�U>�<�&�J#5�����Y.���
 mԾ#� _���Ґ
��M�����U9O��:P�ČmպJ# ��R��,:��/0;�2a�H�2J�y��LbX�4��_i���a�77ذ11e�4I�4�@N��F[7%�b�v	�柬p��!lh�i��G�l�Tq*R�?�e�F�-Z$!��I�z��� �,5ғd�Z�R��D�.����=I�zx�j埪� �[�3e��:'"���#��b�]k[�z�sQ	�b�ԅQ���''^̀��]��P�^���۴��Aq����I>wJ���s��j�+���qB�g��1c'�����Z��_+��Cf�1s(��3ړz��(��\�oh�3����l����'�6i�0�\(¨aGx���4i������M�O3�}��B�c��@b!��^�"��Dc.( ���ɵ_�(��#^Yh�����V�$��C��@�DGy2�1\d�����T�.��c�+���C+70h�kS-Z8	8.01�IΈO�qx�F��(�Tp���2��}���Y�,�WH��N\!�\�;�X˰���"~�	m8�����"Z�4�*��H��"O���t�s<�Ș7��..6����Oj��a�=:s~y�	ӓ X�c�� v�j��v W�Z���I�4��WDK�0�Ԩ���*9���pC��. ����'\x�(���d
���I��'
_�'}��q` C�O��Ǡ�
x��A�3��( ����'3��6�@,c�`��.&?PA��'� p��Ԏ%��+6ا$��\��'y6�hA�<�6}�E��?�5��� �u���8 �<���I�/l��za"O؀@6���L�:g�ס_ֲ�s�"O�й���� �1�äP��<��"OJy�THN�
Ϥ���L�/q�� QQ"O*!�jٴHxn	c�( @��3L8D�L�� �
���f��=��`�;D�Ђ���1[Q��b�hKr��E�:D��
5Ñ:O/l���D(�z�c/D��Y��ҶFs�8�.��B�<y�Z�R�6�8Ë��`� �1��|�<��+3��Q�d�K4H���A��<^'P�l�T��6-�X0�
g�<��J� N������ ��u 1�c�<�撢��Yx�o�C%��I *�r�<�u��M`�gܶEB&�E��s�<�B$+#�v�{���#) �ۂom�<�R'�=@gnY��{�Me�<!�H�X0��GL�!g�!�`%IO�<�h��Q�j�7�"9L����^�<a�lC�*q2a�v��������M�<P��Zn$ڒ"�(�b��'dc�<Y��^�? �8[�l�7.v����F�<q�h��t���Ì�\���+�YU�<��R�c�l	���W�8�HP��an�<��m�`���ˡdNt��-Ɂ*�m�<a���%-��%+��o�`�x���Q�<�����sb[3`����%��I�<�s(�z��K'T3s�ȅ�6C�J�<��nYE�IZ���MJ̨�	~�<Y��1K��A��B���:�OQ�<�p�V�l	F0s��
XR�tS懁Y�<�%�4):sWȐN��J�� ]-.�1cBBr������5Oޞ�h��^:��(	a$;D�t81#�8j�4\�w(cozY�f�8D�����V�W*��ْʌ"�,�C3�8D��	��܊rp>tڤO�9~4,���4D��V&˴���b��*n�|C�*7D�����)g��J�]�PQ�(!D��ChB��8I[u"D#r��:pF=D�@sU��?�@����p<�S�;D���ע8~X���7kޤnX���!�8D� �C�	���9E۪A��-�p�T��Ol��;�N4���۠,Z�Ą�b��e�4�-z��	y"+��z�a�t�I�#�q9�D
�4�`�8��O$��4�b�0��d�S�'?�x��L\�*`٩w�+�ԕ'���Yt���̘���5?ɷ��C7x���G(��i�j��|�2dC���?��Z���<�;����Fl�
h1�-�l�o`��� �OjD�A�O���
�'�B�D/2*ڢ���h�"|͓Q@6���mV@�+�j��� T��)�'=�
�AǄ����"y0�S>a�2�B]��IT�x3���"`\�y���X}r䗗��i7�t�?�r�HפL�.D��h��=�:����N�w�vI�''�X�`C�OQ>��C�O�D��ϊ8<�D���LX�(9s_���&G�Ed���,��<�j˞\������Ɯ"/B�<�Ѕ���>D�WH����ᓘWZ�<z@��4AA���D�.�n�� l�#��H�J�/B`�ڴ���~:L?��0c�-K��1Ч4�V]2�����?����|h@+0O��#���hb>�{���r`Rt��F[>���U �$A,�~�����	9+b�*Ӂܒ+JT%lٳ
U!������[~=�xP���!���=�L���C� V-{�D�e3!�α]v�'X���82E=a<!���J��H����ҕ�Ԓ �!򄛕7�!ˆ$+s�Z�x�1�!�$:�d�a㜁�vd	��$&z!��O��JM�V�W�j���S�Ї^!�� ������ ?o�p�CM��r-(u��"O����b��jOV����̈́ �p1
W"OT0����w]�M1�!����,0d"O2��v�A1s>�k���`~̠y�"O�R�6"lܳu��@:!�"O:�sK�4H����FH���C"O@y�"��9"��z`M&/�*�"�"O�]��j�.-�.�ql� ���{�"O ��%��S�&<�s���I�"O��Zf/�t�$A��I�xN�$"Oz�Sq��V�V5"�	�b�*v"O�Q��I8|�(,�C%V46�"pɢ"O�q��h�0��[7��F�$u�W"O� �I�t::��0�tW
��5"O�\�����v���2> Lx"O�yJZ/%'��{��P+V6�c�"O��a�=�qs�јT�C%"O\���G��(@�W�"`%�Pr�"O��k��Z�R�p�
�.[3�"Od�@r�����c���-���I1"O4��q�ҝf#"1x��j���"O>#WǍ	a[�y�=o�V�;D"O �)d�_�^o���Iܨ�P�"OdtA���x�!zw�� ˘l!�"O��c礚~��,	�G����*"O�pn)g:�y�K�/wK��8�"O¬@�(�>b��@j��&N�D��2"O�e���Kd<Ձ�[�\�^���"O\�!
ttÀ`W|��-��"OH�g�]{�*u�Ԯ�e�ܤ��"Oh��0oK�26�MAw@ꍨ"OJ�I�Kɡ� 7K�6%�=��"O�����=K���bK׼d���"O��"(�Xp�j����Թ�"O�����$�l���H[�@[�"O�@PT�n����	�jo���R"O�ႱÖ� vP+P��cgd�a"Ox8cξ;��<��%��a�� "O�Y	C*"kL�C��\-uφ)A7"Oڬ����{�X*/�b�lը"O�9k�m\�`z4L��&m���1�"O~X�"ȏ%k�1���{$��"O��*���fޢ���ӱl <H*�"O�$׀��+`Phꠌ�?7
*T�e"O�Y(d�Ϗ
0�+u
[1R�U��"O��k�A�����`B*ƙV U��"O�� �o΂l�V�g����hӀ"O69�f ��7|����Q��i"OBM�Nԭ}d��"L�kFB1�"OНQ^t���ʔ�D�ޒlP"O�EB!Oھ��Q؁���Q��"OL�Sc�T*\�H� �|�2�Xd"Om�/�vx.	�����p�s"O$����R�sJ��ڴ��49�|Mx"O��K4���Y`Y��0?�4)`3"Op�yc��tm&����VV/�l� "O,Ra$�"��}�PaY�`�"O�PqF�F,Q-�	*V%^�s2���"O�u�v�*P����*u\(h��"O�����`�U9[& ��"O< �W#�6b�A\��x¡"O̙ZtNJ�	���\�'��R�"O���.V�Rc�E���"OvE��#�3$�z�P�"rZUA�"O� �i0T*L �(@jd˜@~��@v"O�)���>lƄu�Q�˾FF,��"O.4IF����1�@Y�*�}�`"OPQA�"K�Bo��Ţ$�z�"O��;H�>�pϏ"񠁐�"O�	h���8@dT�C<|����"O���@��.\�=T�3P�(U$"O(�	4=T�7B�#-s.��P"O*�bG�E�i��\;f�ςUxn�+"O(E: -
}�li�����0O2H�3"Of4`A1�l��m9�H��a"OFA[����kNH���L�\Μ� Q"Ot!�ǯJ�H�<Z!lE #ɢ�@r"Ov��� �`��|#T˔M�0xg"O�;�"K���X����Pt�"O6� � 8�dEz�҉xT�"O�{Enɋ$niC�
'��ځ"O��D.�*�v�(ag�A�n!�q"O�%�U��Sd���d�R�"-�!�"OҜ�	E~��Y�W&�3v*� ��"OZ�����`&��B�%J�)X�"OX�;�̼W�8h%	@nM	S"O��H%H�p5��+��)x�ð"OT41�`á;̒��b�]�*(���`"Oxt���@Yf�.j��@�"O �z�d�B`\���V�`r"O�YI$E"U'����a�x&�R�"O]�t�X+)���	��3W�-IV"ORliQ��1F= !;��V/Yk��*v"O��Ӏ���ltm�g�_RLI�"Oѳ��2
�X])��o;�a��"O~u�B$�
>Ta+�勺} Pd"O5����,A�J@�]��e`�"O�hy�푥	��� Iݍ`nH �"OX�$OU�D�1���Vn��3b"O��J#��QAja� !7����"O,P���ԗ+N0�뗈�3s
 u:�"O�,hA�K�KyBi�f^,^(T@6"O��n�����˰N�.�	"O�ș	L�N�H15�ǿ$.��"O�-	�Q�N���sK	*Pl0�r�"OuqSnD}jt:KNU8�� �"O�L�f'L�bR޹Zfk�)oV is�"O�P�Id�������ʸB""Ot$�Gg�zP�#�I]N�P�13"O��8���%S�ꘋ�f֫J2�4R�"O����.��H梨��D��L�:� a"O�@��C6ޑ��"L.QR��r�"Oh�k�!אX.hi�t��]Cp���"O���Z�\h��O��v��"Oީ�-M<
�B��AC��4 G"O��2�� }Մ��JB�@�U"OV� �?��8�%�2G�}ڕ"O�ٙ�(U?$"�U* �~��[b"O�)16.P�^�舗-��<�Ȭ"O��bd��*�еʵ��9���"OH�Ɗ�>|_2`B����~H��"OT�0���1�	����"U���"Oj���׍<�������L��"O�+��6_�K�)}3����6�y��^�̀9��^HR� b����y2�$1V�jp�>�tU�1
S�ybBIn-�HwG7;�5��"΅�y���?�P0��AX�6��]c���=�y
� �iص��J�R�ŝ��� ��"Oـun�8U�@Q5�ӔW�^L�"O��R����a �1Ft�%!�"O�IIV)���B�n��R}��ء"O���Fʙu-N��T-�8�]"R"O��#�J"c�2L;%�
�2�"O��� U���)���X�I�B�(�"O�쁲���<�.I�B�ӆ�Nl�"O
Hrr����dc�E;(����""O�9��G-f�0�d�	�&���"O*��vϏ?9���!"��j�
�y�"Ox`;��H!}p����`�:U��R6"O�!�J4,�j�F�R>V�"O�ࡔO��He1%&�,a��"Ol��L�?K�d%P`�	q���˱"O�Us�K��.,�hw�C�b�T"�"OJ���ܴZ$�(���f	5D�DhRF9����צ$�5�ק1D���kƏ��\�Bb�]�����"D���O�-rݸԻ3��'Ş�)F�"D�S�Z�_���e�[�@#��c�,"D��[� ȗ'�v�AAFY��\��v�!D�\��4P"�{`"Y Y1L���M+D��с�	~rxr�dC�Qx����5D�`��:M��D� 2q��P��5D�|kClˬ&�Mp�(�*����/5D���G�0q[��e��:a�	#�8D�@��
�s!�����Q�$\�G�)D��� o��l��H������@��)D��z�B�)
G��b&�8n��G�&D�l���79a�`[��Ū�4��n8D����AX7�ؙ�/�L�R�S `6D�苕E±o�d��Ѧބ!��ȔO4D�$ �#v쬠�1m�0g�c��1D�@��"�#���A1E��b1 4D�����Z��[�c�e�a`P�,D�\rҚ<��Z��	�'#�i5D��K��o���`�:3���(8D��q��V�khJ0�ԬIKD��a3�6D���UML�
 +A�+���p�n?D�Xɠ)Q�6n<i�NF43��j�?D� #�T5K��Ã�ȂZvd��;D�2��M�R�ݻ���/�V�ae�9D��ëW� ���e/��R�,D��Q�EA¥8�k
$I��y �/)D�L*M9[=D�y�j��%M��A��&D�����	@�=�&�@*C���j�9D��W�V�@�[ �a��"C,"D�,�_�p�"s�<�` ��
�$�!��ء;5ԀB�޿U� �HeZ[�!�D>^_ZE� 醶l����eH	{K!�DҖS�|ȥ-��4�t9��J�m�!���x5r��+_�<L�RCOJ.A�!�ā_t�舀���g�%��BG�!�ܔ} PIA�FN�
J����R�\�!���K|���B�X!4Ʊ� �î�!�*Fِ};����42n퀷��:p!��:|T��Q�	��!��I!�;/Ϡ��c��#]�I(���8�!�A>>�Z����?L��fmq�!��=~�~�S��$��I�a�I��!򄞘_L    ��   �  W  �  �  �*  �5  OA  �L  X  ec  �n  z  ��  ��  ǖ  ��  p�  ��  �  D�  ��  ��  R�  ��  7�  ~�  ��  /�  ��  *�  s  � ( � � B! �* y4 �: B �K �R 2Y u_ �d  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m���'�Q�XI���M�\ ��cI
lx�2�>D��c�&q��KQʇ� z�d�D�<D�����((�[E�/_���)��<D��8�ǡ��!D�'����?D�����9'�[歌!����=D�L�끐Gp�u�C��:r���ȵ`<D��1b�E�E����b�3&�����#;D�� c��R.0�@�J:=�t��(>D�����ՌJ��]d��	����V�:�d2�S�' J
ssc�+@����!��Y
I�����i�M�+L�u*Yr�]��.faR� Ĥ>���0B���H��ȅƓ�x6�S#VL]A��aרub�'���A��/$2pt���
T���'���c,�.������]* =A�'��k���1}�`�����]��!
�'pP^
DL�q�����S����	�'�`y t�I7��Yy �_�O�~�q	�'��`+p��`^�����X�;�$��'7�[F�2PJ20���\(�ݸ�'k@@����%AtY{'ҽK� ��'<ў�}3jݼEG�!�a0w+:�) �S�<)��*H�@����-w{�M�W$FS�<aE�*�*�����C[D8���N�$��k�XC���`��G]���b!D�t�@NX�Qd\x2�I���c@'*�YQ����i
2~_|�b�씻)^e�U��9H%!�$[F
�(�����8h����'nL�e��'.昉�d 	+��]��'!�1�5J �8�^��F�#)�q��'�ȍ�աQ ^��H�� �(��'l]����
�\��ՌT���P�';������@;��b$�?_�P��'&�3 C�D�^]�6��XZ�'#2����H�'���p��6VO8���'�@��RA�aX���lˊMgP�
�'�B�Qv(���fM�7`��'��Ik��4($q[��Q(=6���'�����Y0w�<P�RŎ1(�A��� �Y[vDJ[t�#��#:h�R`"O�\3g
Υ6�q�J�V'�-��"O
���h��m�`�d*ܑ~&z�v"O�|3`!��3��E*4�G.	�����yBJ��U���� �B2"�Y'�I�yB���G�� %l"�:}:�@��y�@^�**���"�7|��	�ˌ��y&�%)�""�!w���K�J2�y"���i-��i!^�s��H��y� ��_4��.ׯZǊ�SU]0�y�`�%or`ň�DV�x$d��yB$A(ڭpn�$I���Iq����yr��-]��Kc�ٖ>�b8P0[2�y���5^�س���
<%����D�y��F��P�V�=.& �� �Ң�y2g�6$��2���u����	G�y�οq��nc:�W�7�y���f��9)`i˚|�-y��L��y��R�N�B�3�!� *	b�+��y�N�} ���` �~�~�p%�;�y"F59��haVfqR�tR��y"�9*x�c��g��� u����y�FȦc0��eP�[���`�-��yba�a��B۲V�œv�J�yG[�5�|x�D��I� � F��y"�	R0��JL�J
d9Ď߫�y⫆)Cs譐G*Q�ʄ� �
�y���)AB��Q`C�D �,ź�y�"��6%*ɤ��p/�T��	�y"�J�1�����R7f�~Y[� �y��w���*$�0ff~� �� �yb�i2��*bT()s���y�醏�	�8Z����r���y���-G�4(�\�~ z�"�P�yb��Bq~�i�jQ�^�R���ؿ�yR
����'��Xu`e�bɛ&�y�M��^��@U"�/K�4���̸�y���'J���2C��B	zdA��yB���٘�W��N!�@��#��{�-�)87J�3��_lA���ȓ	[�)2�-C����H�&j���+��5 7N֓N�D�JK"`$B���^�����{ �t���BtՆ�z[>e1# �O8�ّ�HAe�$��`Ê(J�'0�=�&�>.��l�ȓ)zV��CN� %X$��.�8Z.b܅�+��)��A�Ky@�5e�2t�$i��7�H谊�A+�L8�M�g�D��I�( �fD�e��k�,T=󾥇�0Q�}��MYMV`��ڌb�Ve�ȓA�J�{���bHLi��C= |!��0̌	GG"&t�'ϛ7�Ҝ�ȓba.��#�!,J�mra���Zs�E��AQ@D�A��E��ա%� �:o޽��
�U��ʤW��-k�&�#>T��,3�۔��}�f�b�
.�T�ȓ'��T�e%I�b�pY$���vy�ȓ$������P�zj>Q����$Lt�ȓB��������s� �q�A�H�r(�ȓAW����W�X�j�*��<��|�ȓP�$�k`��i�.�ңi�|�n���- I��a��qr h��Tхȓe}z�3�MG�f��xZrE��U��S7���c/�,Q"ύ+IX`��S�? Ԅ�GM;e?��ʇ3��"O�̫f�3\������Նn;��""O�5���I�Jo�"�f-�v���"O5�4M*d����͘6��M˦"O��
��U�y,)b��z�A
V�'_��'B��'b��'t��'p��'Q����=)��X�#^:,t4e� �'�b�'%�'wb�'��'���'��8@��T�᪅X3#�4<p���'W��'�r�'v"�'�R�'z��'Y�� OӾh����� [\A��'T��'$��'��'~��'Q�'�������$�m�t�[�?Ȍ9�U�'���'���'�"�'rb�'���')^Da@E:]��kFJ��gs舸��'��'�b�'���'"�'y�'��s%̞PɌ,�u�;gj�8D�'hB�'�"�'c��'��'m��'f����L�;]�汃���6�����'���'���':b�'���'�r�'�9�7�-:�.XAଏ
;iR|It�'��'5��'b��'�2�'��'TPɻ��� oY�e�Q�].�#��'�2�'��'Ob�'��'W"�'�E�uC�n�:8�7��4:���'���'���'g��'�R�'��'�
�#�a�
H1>�0p%P#u���P�'��'L��'"B�''�'��'x�j�ȃ�s�����E�*pP0��'���'#R�''R�'Irn}� �$�Od0D�M�!S���Q�[�@��MCy��'j�)�3?Qb�i�Ե� '�5�H�� �!29����؍��$�����?��<��M��1� �@7y��B���S�|i����?��2�M��O���bK?�+Fl�$�Ԡp6�ƟW�h��3�ߟ�'��>9c�莟�"�<�x[�)�`��m�-l�
b�<�r���yg�Kx�.�����S�p��s'A!<���'��D�>�|b� �M3�'&�Ļ��B *P0<�S� 2��4y�'��$��4 C�i>��	�?X��r�žI��H�e��=a���~y2�|ҋn�f�
g�__r�NA�GR�!2Cӑ{���� �O��D�Ox�P}��U�a�H�`P%A��&�crA]���$�O��q�"�:G1���y��G��d� h�L���$Z�:!���mBʓ���O?�ɉZ���i�H�
T�1��N\$I���	��M��A}~Hv�R��0l1�%�����!�������d���I��I��`��,���)�'��I��?��V��fsҵ�s��(5r����ў4�'4�i>��� �����ɹ<sZ��ըUJn���/�0Az��'/@7-�(M����OJ��-�9OЍy���W=TY��\�EtLi���	Y}��y��Hoڪ��S�'06��a
ćI]��J��C�v�a�e.�$���1�*D[7�
G����Xw�$O�(�'7=JUG3�^��(�.<��{Q�'}��'�b��TU����2�\��ɻO����%�'�|b��F8�I�M��"/�>1w�imr6�]禅C�g]@���J�$L䛳�A~��l��<���~s&8(���	��.<�4�A��%P�C:8�H��сJ=?-�-IF�}���	��p��ڟ��I�P���iI�!�0�hR�U�uL4-�AE]��?���?q��i��LCTY��ڴ��X*�<��#�5���p�MKQd}���x�"zӬAmz>�竗ɦ��'�T�x&��s�8���ּ��ܓ�E��#_�����D�Цm�'���'p��'�<�3AiL7�~�s�.l���'�����iy2bx�ԴPv"�OD�d�O��'Du@��CӳC��)JT�2`�' �˓�?�۴,2ɧ�iҀ�{2�ϝ)��D�#X""�`R�D)�6�MEybI`�9���O��Ӽ���>h<���,Ôe�L(�م�?����?��?�|r/O*�n��3@�Ȱ-��A�|���G�8g<���ǋ͟��ɤ�M#�BC�<�ڴ��scö�����7.��i�iaj6�%	X67M ?S�k�\�'���U?Yi	a$K�Lɓ�l|tT�o`yr�'Y�'�"�'�U>!�p���_!�`��Bz�8ٴK�p|����?	���'�?Q7��y��*d�ҙ�3Ǎ$&�<�r �Ս�6����aK<�|����"q�{�pC� L�7�HA"�̣4��h��z�xqc�T�J�d�<��i������	-^��R�F����R���i�>�������� �'ټ6�ۇXU���O��Ϟ"���,K<nrHB E�U��⟴��O�nZ�M35�xr�ÜM(;�N�8"�`P�C��D�,qxѢ.p�t|�'�f�݄._���O��;�%D`|$�Q��F8���d��Ov���O�$�O��}λ[	L%�GG�3�\,zD��j�P<��9D�v/�E+b�'6�.�i�I��%��m%^pK�"L���M��N`�H��4���c���q��w����ESDŽ?��c��`���R�
���=+���hy2Ck����?a��?��?1��l	�}�wf�U_$A���0�l��/Oحm>o�	�I�����j�'�ƤqH�B�B�R��cy�^�C�44�Fl/��I��ӡJ+к�+v엩��V�gӆu�'�N���mOu?�*Oz�nZvy�D٧'����3�8XuK�$� am�'jb�'a�O��	�M�7c�0�?�������rcI(8$[riT��?i�iV�OT�'9b�i��6��H�ء�GiQ�#��dq5���)T��y��{Ӕ�sV.Paá�?�'�֝��� D8
荣klZ5�����Q�:O��d�O��d�O��O�?�{&F.)�ԙ���&1�.ab�L�����I�X��4�fM�O�6�;��¹=�9�	7��9CJ~1O��m���d	�7-}��1Ï�soz$���ieqP��)�2!&� ^Q��P≵��$�O��$�O�����ЅOյfuBD���C�)c���O$�,��&�Jd2�'*BQ>I�U��:)�.(�J�=r�Z�B�,?%P����4y���.*�?���b��XXe�֘��|���9+<��F"E�S�Ԭ�ɳ@���0��HQ��Ԉ�Ok�����È�viP�
��K�Q���O����O���I�<���i�.#Ds��I�_I�u�e�ݮBE�	��M��I�>1�i�� ����6XI#+J�V�$�u�j�p�m�%z�n�\~��L6R]��V_�0\���ĭ:y �i�Fd5��4��d�O����O���O����|z��61u�hidׂs�<QP3&����&M�-ib�'a���٦�0wh��,\T�����*C�	��4��&k7��E�qi>7�b��ac���ȸr@Ї
���(|���.̎*b�@Iy�Dc�p��?��@��e�f�=��r*��pػ��?����?�(O PmZ�)�,��ğ��	�?fl�8�l��1�I ѷzz�Y�?�#_��2�4Cb�FF-�D��l��wD�5J���[w!�?i3�Ɏk��-&ͩ�ک�'5�ם�ae"��؟(�U�3LP:'�0q|�D�4�ğ������	ҟ�D���'"��@C��*K��HxE��(����'Ub7�)5���D�O
qm�T�Ӽs�D?e�4L�d�Q�^t�{���<Q �iW�7��ݦa��YƦ��'��<#Wb��?���^����v�� Pp��%⋾w��	��M�*Of��O��D�O6�D�O�x�I���T� s��P���<��i��y���'}�'^�O|RHN�Q���	]�a�	T�R�_"�ʓ�?aڴc�ɧ�'G̸�jg,�Fjlbb!
B�F�)�$X�j��9*.Oq�����?I爱<)Խi�I0/��y%��-��D�GgJK��l�	؟���⟐�i>a�'͞7Xp���J�sJ\�Q��@1��H��L&ru��D Ц��?)uT���ٴs��FEoӰ�"$D�3M�^T�"sV��g[�/i�7-'?��OXi���ӹ��d��?����z�P'��9j몤H�d�/-7��O����O��OL��?��o0XJ�*��ł�J,g��\�'ҏl����7�*���Ԧ�'�\2� �{�l�S,��1O���ON���b�f�f��Ỉlt�7�#?�d� �쩋d�nN�lY5CV�l� ipn�O�Ѩ,O�Yn�CyB�'��'�nֻm�.MP�
�F���+\�f��'��ɽ�M�䒶�?Q���?�-�x��1��/bd�\���\K��1���X��O��m��M�Ûxʟ�H�;T}�!��`���U��4����Q�ݐ��˓D뎚��?!��<�;F���h�E�>T`�[C�H��M����?	���?1�S�'��D�I��T�n��4�FN�҅�����B�'T��0��>�M��¥�>��i���K��W�jj�]���ɜܸH�v�oӐ�d�&Q"�7�~���/A_媕���6�ug�'���mC	����$�͈�C��?�[�0�	�����h�I��T�O��qr��3f$�tC�)��فdz�n��T��O`�$�O
��b�DF��$z�J�(Ԣ�����
��U�2H���M���|J~���M;�'��R�G���b�0b�� k ��'|� 9�H�ȟ  �|�X����şd�B˒*�f�թF,O�@�y�S��t��Ƛ��My�!lӔAF��Ol���O�8�$g��DV�������D�x���)����d�ݦmy�4�'#LM0�Rs���1_SԵ��$+?�׆���ڄ�Kɡ��' �����!�?�2�F�Zt+�M�>#���'ˀ��?i��?����?��I�O��*�L׿KD�� �6�%k��O�-o��`op��⟐��4���y��ǅ8G\E�A��wo�`ꂀٞ�yr�'��IqN� o�k~↍�.�����8��!sDd�|�$�2rFQ�����q�|BV����ݟ���՟\�	០å��0�Ұm3h�k`��?(:z�i��ƅB����'�ҙ���'|�d2���9&!n$p�,P<��|Z���>	�����O�:Hs�P!ɒ�b��(Tz��DG) �X�X�0��DRr��hy��պ4)�W�J�AzM�-29�'2"�'��O1�	��M�$�Y�?I�Й8̵1�)[q�֠jh[:�?閰io�O�8�'"�T��[r��v�"Y��I�8Wv����Z�VOil�S~��:k������H�O��)�o���*B��C��X+�aH#�y��'u��'^��'��iV�?G,�B�]�E�,0`�͝n�b�$�O����Ϧy��hw>A���M�I>�c�5@9<M�a�S�8?`i�`�?>�'|6-�ݦ��;�4�m�j~B�G.k���#�,+�5�u��y�x�������|�Y�����X�	���*�M�w�`L8U,:1���ٖ���`��Ty�}��X�O�O����O�ʧ(���J&�Kj�R�1��-�i�'s�=��pӖ�$��SF帲^Sr�Ci�=yx\%!Ga"%)����4�t����\cO.����1SGd��'���E��,�O����O�d�O1�,ʓ(ڛ
B�Ux���Q"N*d��ԧ)1D@Q��'&�Jb�x�(��Ob�$Vu ���t
��I]X��aMDb�ɦ�	�Mڦ!�'BHX;��e�*O� �`T��8{�@�hc��9���5=O��?Q���?����?9���i�N��YgF�-
]h8I���d��6-��)�����O���1���M�;B�d$IS�S�es�����n'y!���?I&�x��
ڳ
��8ON�AB�F&.�v���NG|�.��3Ond ��~�|"Z�|��̟�a��"s�i���͊Dz�S4%�ӟx��ޟ��	py��f�d���f�<�LxT�p�K����Sp@�/O�m����>q��?A`�x"�+���a��._V���bƜ1��D��Mh�dӠ�%?Q���Of�dZ���U��kyD�T�7�R�c!��+���)�)Be>`+��*��զ�2����M���w��Ճ�g�J��Q�Z�X��'�B�'�6�'_�>6�5?�@�-~&���xF�H��IDo*��L��0߶m&�ܗ'�џD��O	_z�:t�� F*����4?�7�iO*���'���'���w=�� ��e]�|�42�H�_}��'�B�|��d����0�7��.�u�B���:ʬ�i,6ʓc�p��@&��H%�l�'�~Q�sj�/4�)��d��=2���	�g�&ƕ�b ڜ#�1j1�(�`u�q�C�h}Ӯ㟨`�OB���O�΄��:e�a�;r�^�whĒ0v�A��fӜ�K��H1��?m$?��9D	�!��j�ܜ��ifl������̟�	��D�	A�'/�T�%E��y��MYCd��Hl����?��p��\����'TT7�%��	�~��m@�+�jx���N�3��D$���	��ӌ`��om~�B.{�LE���=1���w�]�9��9h!�e?�K>�/O����O����O�pr'�['y� �8����{z���O����<�E�ixP]��'��'���M��ೃc	�>4���BO!D,:�Az�Iџ������S���WShX�"IR:=AQ�BV*A8�XpE�\3ٛF*�<ͧ�P�	P�	�;�ܐ�-Ƅ�(e��Ɨڐ���͟����0�)��sy"jh�@D ���$�2��D��(>�X���Li��O�dm�|��x^�	��D���I�S�`sb�8a)&�ɷfFԟ<2ݴ��<sݴ����)+	p��O-�	�Zbl4kfԿ�b�BlˎGD��Iryb�'2�'���'�V>}���:�*�A�G�q��Y
\6�?1B������ݟx&?��	7�M�;1p�I+S��bW�]S%
7K��!���?9f�x��4�F_ۛf1Ohp(WOWN:�h	1,�5˪@�e<Opu�������䓽��O���5-�0:P@��y��,�Ѭ��TW���Oh�D�O����ơ��_f"�'|���.Tn!6f�])8��E+K���O&x�'�2�'+:O�#�˽���;����F��V���7D׈8���o�.��'r\��џ�ږ$^��$��EA�7?��#������ǟ �	���G��'��H�]�G|z���Yj�l���'��7�L"A���*T���4c�	55f��Sd�Z�,�4�	�:O����O�1l�T��lB~B�A�YƐ�'TR��*'b��Z���1�ǆ%41�O>!)O��$�O@��O����O��rW���!ڙ�DE��9as��<Y%�i�}[d�'k�'��OjB͉�p�Ih#�d���-� �I�OĐlZ��Mk��x�����>k��S�T�D���Ō�v�6��G͑/W��I3dځ�4�'�\'���'|k%囁v�H� eCD�����'��'���Q�Dy�4h��3��\?���tL�2D­�&�ʢĆ�����v���qy2�'ś��g�0�B3DY"Y-qqdثQy*p�A��y'67�0?���	���)H�䧍���Q�A�,p��4v0�G-��<���?	���?Y��?������<���g�˖x�$r��<b�'mdm���23�.�$֦%�l���_��<Qj�fܝ
L���&���<�')�P g�i=��6
l�i�D��(h�,a�
\���%aᣃ�Nr�BC�	Ty��'�2�'B�ȵvb �[���8��0i�N�>Nr�'2��+�M3&J��?���?)/�J��҉[)tMC �hҶ%6��t��O�!oZ��M�v�xʟ�5R��P�+��C�	5J��8Qp�Y#H�j�J�@P�FA$��|J���O�J>Y��JR5ȕ`�6P4:�1�OC��?����?y���?�|/O�o��l
6؋0�E��=X`��Y<)��E����	)�MS�2`�>Q��i���#-P�H�@�u�C�=�e*�.nӠnZ�P@*Ml�u~BmЮH�\��w�	y5&lzf�PHu��Ԥ0��Ify��'��'�R�'[�]>�����*+�j=A�97⬺dH۞�M�"+��?���?�I~
����w�����E]�Zq���4���8���O\6��K�)��P-yiR7-c�l-nJh�u�*'ܠ��S�c������P �JI�	lyB�'��'ֻF>�I`����l)RJ
�y,��'3b�'��	��M[��?���?�$,�9熄q�H� Yڽ�b��8��'���N���q�l%����R'K�4�*�o�,d3L��2o"?�U&l��qȠ���fm�O��m�ɼf&���T�H2�Lȧ���a Eb?��'���'G��˟Ԫ�a«j��A�Vc��oY��r�@�4h9�hb���?� �i��O�J8�u*��ӓQ%�tK������O�6�����Jt������'s�Mb���?ՙ� ^�b�]�ـ���
uט�ᢁ<�Į<)���?����?��?�Վ�����ÇF�ƴcd	��æQ�`��cy�'�O�B!�!H�� �2�Y�q��#��#�\�)͛��n�D5'�b>��"�<:��'�)2/j4���@� ��q��cH|y��^] �	�!��'_剋
�/ED4Q!~�Xika��O,���O��D�O�)�<!E�i�|���' 8`���� ���\D���'��6M?�����æ�޴�VÈ(a�t��g�t9��,_�x�� ڂ�iN�I�|��(�O� �$?���/@~� ϒbMTkf�ϊZ1���ȟ4�	柴��ߟ���A�'&�:��֢���`�R��e\�C���?���a�֮��zL�.�M�H>�3$s|�J�g�8����T��?�-O �kf�z�=ÌA�'^�K�˶/W�uJH���E�{p���i}�O�˓�?a��?��$���0��N�za�S��HY0��?�.O�|o��y<�h������IK�T��0 ��0�׬5���Kŭ	*���n}��'��O�S'n/��#�ϑ�t�dʍ�%��q�A_�M���1��ly�O 2���92��'z�����@ֺ���oxD���'"�'�2�O��	��M#Ǡ�&6�mT	1m�$P�TK*OD�lZ]��1�	���&E ��I��珚f�Np��&_yB%P'6����d r��8y�$�UyB�M�BM�PgPA���ŏ��y�T���I�$�Iܟ,��🄖O�j�;��6��EZ���
��˦-�OT!a#�'I2�'���yҊy�󮐆^k�eiU���B��F�	Z����OʒO1�ر[�Kd��w#Np*���cKtuJ��Іe���ɧR�1��O��O�ʓ�?Q�w�������h�j��Ҹ~�`���?a���?1-Omn5!jE�I���i�A�A�Z�d$�㩊�y.ԙ��$Q{}��'�ҙ|rU�1$�f&�	E�=iT������L2)�1zEnuӖ}%?-k��O,�$��XP�"Om4����6��O����Ot��?�'�?	֥�'7����G�?z��[�J��?y��i�v���'
bFk�P��]js�ݲ/ŤJ,8�6�!]�����L�Iß@�/�Ҧ��u��Y�]��V�n��̡Fn3�͸�b�5e��O���?����?����?��tG�m�6��'!1� e��-OTl��[�*t�	�`�	R�S韜AW���t��o�%��Ug������!Qڴ|����O-��K��'SAI��>P��_� 
i³P�``���}�	P��iyr 2�;�N?�<� �*�6H��'��'��O|��-�M��bԊ�?yCl�+j� �Q����P�z���B��?�øi��O�-�'!B[�D`�'Ɠ9��H#�{r0@�-HiO6�l�H~R � ���?~O�OWEe(����cE'Fz���"�y��'w��'�"�'g��i���zp�Ԑx��Qb�C�o&n�d�O\�DYצ��t�$@�i��'�>����d��*$?��{�y��'�剉}���mx~"��,���n^�4����dH�� A��ɟ09ї|�[���I�������Hhs��I&T��V��0zͱ����`��KyRC`�0P�c��OR���O��'w�F�����.`%t<ӱ��Wּ��'gD��?q�ʟH �V͊�zθU���Z�
�9A�w�]H5�W5
<��|"T��O"P�N>a`j�M�-0��G�7���Q@���?!���?���?�|�)O�HnZ�r�ͩ�O��+F5*D��5.8�
 dXܟL��	�M���<�454(;1�,��El�984ʴRS�i%b7M\�h�7'?	K�/��Ɉ9��d�) ����a��k*8����!v��D�<���?I��?	��?a+���c7̗�&���dN;V'0h����)PU#_ܟ���ğ0'?��ɯ�Mϻw�^@Sc��q>� 6�v�Th{������Opf�ʐ�i�S�7�ȩ���R�~ Kp�j�󄌜!+� ��Z�O���?�����Z���[ai�,��͢d��џ�����	byB�e�T �+�O�D�O�`s�ᄙO�Rq�ň6c+d���.�I�����O:7͆v�	�Yg����gM�!
�J)~�>�z��X��H~����OR���J�n��	Ic�\X7��Z�����?���?���h�$��ܵ{-@E��-p:����w���d\��%��$�ǟt���M3��wƎQ�)@�v�m�B �0p�v�۝'� 6�����ߴѐPݴ��D�<,�R���(#PN�4W�����U��y��	)���<I���?����?���?�nV�.J�I1 	_�U����A������;����`�Iԟ $?e��+xڌ��̒r��i�o�� �/O���u��x$���̕���S8%�@
\<��j�e�7pHq��Ⱥ<qt�#����B��䓢���9�)��� �m�ph�v^#jZ�D�O��d�ON�4��˓"�v��-;rl!e~0p���.L����"�y�gӼ㟸��OT��<��N˹�d����\�x0�T(�	~j#�4���R�_'*����(&��8�n�;l��<z<���S�p���Ox�d�OH���O~�d*��- ����WO`zb��KЊ[�����ȟ�I�M;���|��uǛ&�|�l�M|�e���f�!��A��'h��'�2�1&w�&>O��ِ"�� ����h�*<�#��G&y{t��?���+���<����?1���?I6䏢`�x��f��ADB����?������W馱�u`����	��O�.��4>we�x
��ϊH ��O���'����?�c��1K��X��.��$���B:X*�8 m�%��(���d�����3�|r.�����P�Q�~�"8�2���B�'��'8���X����4<����ɓ�w�dd�B��!�Da�W���?q��|S���U}�d�Ȉ�q,���*���=��8��ئMs�4^�­��4��䚳X���'?�@�r����F"���(��)^�e9�q�����O���O(���O`��|:�E4��8�L�#��M״ u�F�%�ϟ8$?}��$�Mϻ:���>Qʾ��V�'�j������O����$�ib�#�ԅ8vL��lY|�A#J��d]�x���������O���?��o�K׬N�F!0a�l������?���?a(Ob�oZ�bͲ0�	��	��� dPy������1 ���?	sP���ش>�V�/�� e�xq 蜤測�qƙ�cd��8I�̥��%(�t�&?͙��'�t��ɿ�!����?o���R��R�&�R��	ٟ�������t�O�����% ��UFNuk���t�'G�6�96���D�O�(nQ�Ӽ�LC�-{��r4%Ѡ��|���Q�<���?ِ�i����i7�I�D��K�؟2���*�tsZ|Rǀ�-o�v��p :��<���?	���?���?a6�Tm#� �lY=pNX��Td������a�S!D柀�����'?牚)�P�R��IJ�}�C��4��O����Oވ$�b>�0�	�%J�n��ώ�V� �*��*�oZ���w$���'��'�	@�4�c���?R>)�AN55�@�	˟�������i>�'@ �$�=X�n�=~[�s�	C2Mu�,���X��yoa� �\a�O����O��n��5&���@�4�jAt̘�z��ߦ-�'w�!brgCErK~Z��~�r�RQ$��~f��9�n�9{���̓�?Y���?���?�����O�d�ڀ��&f5��ڕF��j��!a�';��'-<7�7%$�IQ���'�I�l�D0$΂.�p1H�%��N�"�%����џ��	�Fd�m��<1�Ox��
f(�>P�+��Jf��#��/`���5�d�<a��?���?��ѽ-�Ρ��g��'Cx� DĂ�?a�����
ݦeR��Zyb�'�-���W."��,2���4Wy��kC������Y�)jb��G��	Jf�Xjt�-���W='ւ��`�V0�M��Y�擅k���:��mA � %#�Q{��:z����O��D�O��$�O1����V
�u�v��e��x-��d�
0R��'^rfwӼ� �O�dC-�����ņ5�)Pɐ=l���$�O�m@�oӖ�Ӻ��I�����\�4�5�ۦ%�����'����H�gp�d�'��'b�'zB�'-哹.�� ���w�Vt����!L����ٴE�n`��?Q����O!>7=������<�z���0@�x=�Vȝ�e��6-�Ʀ1�I<ͧ����/�m�ߴ�yRd *+	{�㆗>�Q0f��y�b�g!hd�Icm�'#�	۟���(U�Z1�5��
��d�U'�(����������ɟ�'�7-��crJ��?I m�D�9��j�V�(4*'�*��'B��d�6�u�\!'�,7j��|ƜIPF��j/�A�h*?��h���3��P��� ���P#�?IBb];Z��` ����,���!ݜ�?���?����?9��	�OLy������d+2eR�����O@Po =�ܔ'�7M%�i�� �I<�1��>U�XՊDn����^y���˛6���S��կI�T�ɝ��9��%�F��0!HQ�(��$�<�'?2�'P"�'�"�'�R��ao/�ndK�N�D�VA�1Z��ش4� ����?�����<Q��ٲhEL]��H�
6�i�&j����ȟT�?�|dˆ �����f��b�:&� H�l�����X��Cb��O�ʓ_��T4�Ӿ7�䥘A� �_��A��?A���?���|�,O� l����ɵ��y���Bx�z���.gC�Q����M��R�>�����䕗8+���A[/���84�@$+��I��wӜ���(ŅA�L~j�;0'&�Z��K9f�!jF)I�_��L��?Q��?I���?�����O-�Q�&�]�ze���D͚&H��z��'A��'�6�'y�	�O��m�A�	�j�@)PU,LX�<���+ �N<yS�iD�6=���8��w�r�^�D�� ��7ɮI�7+��Pj��]�
��D�4����d�O��$�O��DU4BalX2�l�� L�D��):�f���O�ʓ5���*?0s��'urR>]��=H\f��FI\�WN`؆#+?��]�`��U�S��![%��Q�5�[1 �j������%�P�DŜuX��[��vR��|�p|Xw$ŝ�����`c>4��ǟ��	����)�Syy��z�rq��/5���K��L�	��f+��S�J�d�O�	l�s��7�I�T�� ߾ef� ��w��!�a�V}y�`A0�F���[��"|��DL@y�nT�Q�4�R�F"�Q#0lZ��yBU���	�����ş|�	؟|�O�
e��
�
Y���Scç{�>�Z�,�O���'02�'��O1�s��N
ej��P���Sǚ�I��N�`9����O^�O1����t	a���)� �!J��.+������7��UQ�2O,��a����~��|�\���	��X�r�8���'���W�N�X����	ϟ@��XyB�hӸ=����O���O8ب�]�-�y�{�=
v�#������OL�DFC≦.�U{��Y���gc�	��3�$�3lI+�M�!��d�S?��C0�epd��+i&���d$/(zX����?)��?I���h����d�$�������*��ۮ����ZǦ!cB��џx�I�M���w}��ض�c�,$*F��@@v��'{��'c�6mV�&6� ?	��X�,8��pSER��=����jJ&O�2�$���'4R�'��'��'��e�� ��':�lj�KI��,��Z��)�4,�8����?���O����p�2p����w���#ZIr$�>	��iG�7-�k�)��Y�$p�d��M��s�a�\�l哑M�O�4��';pY�E.����Ӕ�|r^�L�Ҋ�<JȢ�:A�!�WA�⟜�	����	��zyr����p�'Ũ�2&cťj�rպ�L�.��	�A�'�X6=�I���$�O ʓgI�xb�n��B��̍�~�H5����M��O�U�Ԡؒ��*��������.Xv6�C�! �"0�:O��D�O���OV�$�O��?���*��x����	�`��+���O�l� f\�|����|r��0�P�zE+�'+F��RC0�'�R_����C�ͦE�'���@�c�MI� ���'�0Ut���4@�'�IПP��ןx�ɲ5@>x%��~kx){w�߁I�h��ǟ��'AN7m�$4ʓ�?(�"�ɗ��_�
��jlC��R����O��$6�)���+K>f=�G�X<.62}yԬ��a蔹2uK	�9����(O�	U��?1��+�Ď�4wи9b�Vo���AN��6�n�$�O��d�O���<��ia��;���H��P��dw읳�6#���'�6�.�I���$�O.h�6ϝ*9�����N�*qO��V��Oحn�AйoZd~ښYaj��'��Wc�=�%�%j/�D���+Y�<i��?!��?���?I,�ޜ�F,�;d'�:�!�18
�q�!�䦥�τڟ��I�%?�����M�;i/�٠A++ u��H��F$�	���?B�x��D���:���=O9�5>w:����ςK��(E>O���q�~2�|BX��I�X�������Ņ華�e��h�������|y�eb�����<9�m9��)$h�/dh��)��U3�`���>)��?9�x��LO(f�(C���)��E��(���F!iSE��Boӌ@$?I�b�O�����8j'�P(Jt`B��/M��d�Or��OT�D<�'�?Yr�%^�-��)�
W<$&� ��:j��-Ǧ%���'��6�/�i�%���25y~��)�5�����Ad���	VyB�]Λ��<PsHX�<��臏E=��	�I�S�%]�ܩ*��.�D�<���?����?����?�b���7*����4i| AN�����Zͦ	J�c Hyb�'���԰oք�"�B�k[쉈`p}��'UR�|���j*��1B$����ӠiP<D@�Ҷi�ʓL�.��1B��%�̔'Ӏ����I�Yy��8��.��ɘ1�'���',����[��Y�4`�lȸ�����m[(���k�IW*�@�ٛ���w}��'��w�l5��ZO��QƠfC��"!!C)<��6M-?�K�O���A�����&L�Tk�|�+V4fS09��F|����ß����|�	����sѰ@���h��9xI�'KH8�?���?遳i���O6Bhq�j�O&0��E,�|�02_�c�U��"��O��4�Д�b�vӺ�Ӻ˖��5C'd=0Ť�`Н�ˏ�Y#�'D�'��Iџ��I֟lΓq��@�3��_�ʱ�4de��U����'�7��Hj�$�O@�ī|��_�P�,�J4�H8u����iLo~₰>��i�p7mx�)D�~�b���O�TYץ�C�M01Y�t�* �.O�I��?���3�$� AQ'k �ThStg��z��$�O�d�O8��<y0�i4
�j�[{�6i�'�#��J@�\;Vk�'�l6�#�	�������� ƅ���kU%2=!�J�(�M#��i��З�i��	��ȭc�O8 �'7d�8�+R%b�^�[�!� 1l��'��IƟ��Iٟ��	����X��O��0C���bݣ� �&^��6��(gl��?�O~*��Uߛ�wDV-� Gk|�<�6kW.{��� BLu���o���Ş6+�]C�4�yr8i����Ě3e�L�X�ל�y�kМyP�%�I�u��'R����� zmn��v��@}T�2J��2� D�I�T��ݟ��'��7�G+��$�O���G�Ⱥp�ްP8x%k�ծ0��(�-Of�Dx�|-'�P���7V�~�:ǉ5mؐ-j4�/?�u� (c\	+��^(��'&`R�d^��?���R�=n8�f�����%*�����?����?!��?9����O�����=EL�L��PP��*�O�	oZ�[�@4�I�H�4���yg,��[��p�tH�XP���~b�'	��t� J�(i���
�x-�w���"�
YL2�w�V"�(��P�������O���Ot�D�O����J�����I!X{���v/6������ǃ;{5��'O����'�h!�%����b-!&
�q�>|0�e�>���?��x��T(4ˀ d�!��.�Hx�媐�>k�X5IdӾ8�'���XSɇk?9J>�,O��y�H0y������U������O��$�O6�d�O�I�<�ַi��c��'�6���k��½h�Az�dl�'�7�=�ɬ����O&��Ʀk!P9�ݢd�P+J� �;0cѽE�*�n�I~R���E�\\����'�#5f1Od�a�9_�͡S�Z�<i��?���?����?��T
�:dh=Y��^.Z��P[��I�3�R�'`�O�O��3�Of�,~���Ob��Ql�N:ebcJC�E�4yf�&������5C
xl^~2C��bª��Ǌ,_B5�$'�j$� A��ZQ?�H>�.O.�D�O��d�Ov`@c�ŷclQXQ/�ck\�SL�O���<Aӽi��8E�'�R�'/��7(�,��i�|��Q���P���X��	 �M��i�pO������B҄F(���p��Ha��&�K@��{�r�����M�蟜�q�|B� mN��I��~�X�N4)�B�'�2�'����_���4 kh�6Kܿ�0�A��-!B}B�(�?��DÛ6��q}��qӐ�T��c�>�Sd�'LjP��	��2�4&��H��4��d��.��k��%L�ʓ6�,��&��s��p-Ƌ0�2����O`���O����O��D�|�%�K<���)Q+�ZBh�~d��ω���'G���'�7=��3�B�&y2��r��ac��BՉ�Ot�d�o�)�5JH�|o��<Y
��&����7�H���M�<���Z8:
��R��Iy��'�r�J"	����f=8)���	�R�'yR�'N���M�ĀQ��?y���?���ɂ0Z,I:1#�}����S���'����?9����87`�VI.XZ�Qb�4����
G��A��ւk�D����i�i���d�d��p%�HQ�bt��G��L�$�O����O���!ڧ�?�CRdux��V�ġE$���!Ӳ�?i�iΚp1t�'�Rg������ Ѵ�ˑb�l��#M8,�n�	���'u�P�w�i���>	Ҭ�"�O���x!%>o�1y�芨W��@��]�	hyR�'��'���'I�
�������L��"�z���:(��I#�M����?9���?QN~2�A
�"�M�%>��D� �WK�d�(�P�`��ȦQN>%?u�`�W�(���MB��ica"d������iy��-����	���'��	� ��U	�jWy���T@��9|�`�I۟�	Ɵ��i>ŕ'^\7͎	<e���A���2� K}ʾ�sCG�DP����m�?�F[�|��ޟ4�I�9+^iuG �Q�x�����w՞�����q�'Q��z�HNJBN~2�;]69 gHӻK��"cN<�~͓�?���?9��?�����O���7/��L3��y4��;A�P��'���'�@7-�"#��JO�V�|�_t!M����
C1*���FN��'��Z��2G��a�'y�]@wn�82��a@h,:E꥘���h�"�����'��	������@��"W�]�̶��0��k�
~vE����'I@6-��\�$�O��D�|*��O�j�)d�7u��p�Oh~""�>q���������]���t�ưd6�so&u�Yk$	�5�\c�m�<ͧ`�:�$Y6���L!�M.doҨHC�c.����?���?��Ş��d�Q"���6xn�K��׈K{�k�.R������<��4��'(.��?��/�k�����A��Yh�(΃��D4=.�69?���ڡ��i����$�i��	���.P���Aᖻ ��d�<���?1��?I��?�,���0 DC;l��X�vɚ�H��e�r!l�
�N��I��X�	}����	�����H��Z�;�Mö_4�+�O7/��r��d'�b>�h�c��̓K�������/�F��(]1.�Z@ϓK|� r��O��H>	*O,�d�O.D�↉�C����L[$� ����O��O<�$�<q"�ihJ��'+b�'d��� =en�X��@�#8���6�D[}��'Ґ|rdճR� �X��)$�>��DM�����+dH$A�FzӞ=$?a���O����5~�I�c��7:0)H��ρ"����OD���O��d6ڧ�?i��`��y�OB��Œ/�?	T�i{P9
!�'��}����>�>�J\�$�+y�B1*9O"���OX��M/��6�"?�;N�\5:�O�P�i�'þ@LI�`�E37��P��|2W�x��՟P��֟���ퟰ)���)�ؤ�糊`�c/XC"��;�M�cf��?)���?QM~"��s
���IĮi�H��en6\l��P�L�	͟�%�b>Y�DoI�/Kr��ǒfTB���g�|�|�mڙ���K�K�'��' �I�:���ݧʕY��L�B��	ޟ(�Iޟ��i>��'?>7
�=G���� �<��(�`�^�u+��_1����٦��?�V���I��ܴt%d,�0	F��L=J5�Тqz�X��M{�O���3���������w���c�^�u�@9A� ɝjn>0Y�'b�'.��'�B�'��@c�iB(&�Ќ��E�:���@C��O(���O��nڲ Q*@�'��7m-��۝a��ݳD@�?zŴ��ǘx��%�h�I���ӢM��l�F~���!{���4ȗ+hzA
Al̗C��趡N?	I>�(O@���O����O~�ꆄ��>�,�I!�ϣ!|-C5��O.�Ķ<���i� �K2Q���	n�4̝�#�ؼ��+��{����8���M}��'��-�?� ��쁋gn�8b%�	i�-I���3�"	g�r�E����y?�J>�@�
g��jӭԟ8)l(����!��ͦ-��![8p�Vt�4���}���bR�φ�����`��4��'�듭?����(p��H�p�	s<�`�T/��?����t�4����H�`��?u�'_b,c��T�rߞ�!��5�du9�'���l���R���/��iFjP�Bqa
�?�M{�CD�?���?����om��N�6����K�1���:d����O��&�b>�`�]ۦ	�e$�<PS�A�N2pb�	�4ds�(�4��T3ф��&���'��	6@����س^�����7/[���¦}yD�ߟt�	Ɵ��`��/�2 ��(���ĉ��N�k���� �	�ēJY����T8�҉�ba�
KV���',�т�0�V�;�)ƃ�~B�'P�|;��K
kL��a�CQ�X�#�'ā�@ʄ4~0�r�I����'�$6�E�#V����O^�o�x�Ӽ3!��n�HQxs�Ӑt(��dJ�<����?Q�sE	�4����N�b$�?��V��(���aŌ�01�x�UG�H�	py2�	�]�TJ�>)�*�!�럕;�>�_f�f�:T�'��IK�`"�I�k�X�����6���'{j7�JѦ��I<�|b5%�P��=��&)����#��:-�9B �^�����F�@Y%o��Ei�8P��ǖ� I1� �_���T癷u��u+��r��A��[�>��;�k[�8������^hU�#咡Y�N�jp�F��H#T�1Fizu-ǬH��I���M�0���G'W4D��TA�,��2�44����-T֌�j��Ȃ[�h�@��A�'��%j���(����W�lŹ�$V2O��)[p�	�&l�NT�$��R�o��;��mQ��k��%x#Y,{�n��$\�Eab���Q⹻�oJ�\`���T�T-5ݘA�P�\�}�ztHᗦu ��@�ֺ786uKD��1�M��Ŵ3�ސjѫ��Oq�����bÉ'��|�R����h�>A��q d��P�]�L+z�� �s}B�'���'Q�Iv(�J|��휭�Zp��#�u����hƛ��'��'��IeҲc�\	1���+_��㟀P5:Y3��p�����Ob�`�d�X��t�'�4�SEJ(��j���`� y�!��:�D�<�0����I�!,���h��,J�p����+q̛�U��s����M��\?%���?�`�O��8���Hi(��E/�(y�� �i���R�#<�~���0��Y��ᖶ9�J����1�����M[��?����g�xb�'�����#z� �
����c�	+��c�
��c�)§�?Q�E8R����$�0s��H��՟#���'��'����� �IƟ���3^H��Cw{��� �Ǧވd�>��]z��?A��?q�95�DT��G��l/���	�$ ���'���8�%�d�OT�$�O����7F�]�X�e�G4�@�0e|}R����'=�'��V��r��	��ݣ@l�7����s���o�\q�H<���?�I>�+ON�1�dH�WMܩ �CBi��1r�/ 1O����O���<��E�!`��)�I�
�B��[���p�EX�P��	�����C�IAy�fD���̏^m�1)@%B�m����B�\��	ɟ�������'}*�5#4�WYe�`K2�7,bA�JDz��n��%�0�'dD��}�D��%a&	�Ba�1Ba�(q�X��M���?9.O����BR�̟����%g2肏�5<D�@�����O<Q)OX�(��~���
�5s��'-�2���S�,զ]�'RfĐ� ~� P�OE��O���(rl3��Z�'0bA�@創"f0m�A(<Afmmђ� �	�*J�i� MǦ�`�"��`�	hy��O���'��I'<�hesBƅ��X�D�22"�ҩO��2�)���tr�����@��^6���"֠&�M���?��1P�UR,OTʧ�?��'����&��>LabUZA �� 3h�R�$���O���'n�Z2�����A8�I7�G�6�����̘*O˓�?J>a�睳SaPj6�O.u�^�g	-|�'
@��O����O���O���A=(Ѝh +��#ovh;�dH�^;nE�B�O`���O����OԓO��亟0�dΏ�:1|��(�)rXZ��p�2J����	ן��	Ly".�$�
�Ӗ/�D���N��t)���#@e�6;<������?���7�`��'�Ɯ���'.�u"r#�0u���O\�d�O����<q kE�:G�Ꟙ�a�
o��I��"0rRH�M�����?��,�D���{"���P��v)��y����"�M���?1+OT@�GD�h�$�'���O
B��pgW~!�5�����k�F����%���O��#P8��4�'�Bu�F⃤
2lpUCK.�>elhybIF)�t7m�OH���O��Gn}Zc��e!���s��tG �g���4�?��������ɔQ���j�Ɩ%-ĉ��'͛&` �]=�6m�O���O$��^[}"X�Lj5��~?���׫Ӟ��0um�*�M���_��?�O>�����' �Uy)'��Ȁ�]�"��Ds�Z�$�O���ߟ`�e�'��Iߟ��}���PJ�b�x��C�D�}�>�mS����?Q���?I`ٸG8��Q���N���!�"�)pu���'z")�B�>)/O���.���� ,��%�0E�9H�jʩZ��30W�`�L�[�ٟ���՟Ж'��fΈ-(^H;�K���l-��`.����$�O�O���O��c�m0n�h�jf	�5o3�I�� � ʮ�O��d�O����<Q�'Z
tS�霶G#�Ȗ C5|�F�����U��X����^�	����	�q�̹��r�Er�*��u�'.�K>��'-b�'��Q�4�%��I�O�E괃�'(���&ٻ[6�����\����m������ɳ3m���W���XK��ʱ�"�}8���3lw��'o�S��ɶ-W����O���"-��Oʗ�*0#a�,MȌ帇@UY�ӟ��0�i��e�IjzQ�C��t�@!ԪA�T���צy�' 
"�'d�&�D�Ov��j�ԧ5v˛,t�@�r&�*Q����a@^=�M����?�V
�1��'�q� �k��`nHp�
[:{,���i쮼� �m����O*�����%��3t�.|C&��^ ��&`�����4m�n<���?�*O����$�O.!�4M�	��p����Ų�+P�����<��/�~�QN<ͧ�?Q�'���kT@ҷ[�
Us�B��H�>x��4�?�.O<�So��'�r�'V¯���6p�G��J�d�Rc�6.��7��OHd[S)FL�i>���L�	�Ŏ)�%G� ���HQ��y26m��O�xk�o�Ol�O����<��=T^�iQ(�4V��c]�3�<�B�f����O��$!�	ݟ �	�z�!��d��k!��A�LɈq� c��-v�xc�(�Ify�'�$3؟4쉓cX��t��b!A�@Ѣ�տik�'�O@���O�8�r��f"ψF�����H��Z� �M-����O��d�Oh�S�D����1T�cSIC�PiXl���A��7��O,�O�˓P֨:����Ӫ6B0Y�j#1o�x�d���`�7�O$�ĭ<I1fU��OE���5V�%w�l����~a;�(�M�,OJ�$�O��b��O$�������z�'X=i��
`��bm�y��in�ɈL'�,Fj��O�2�O�����H�f)P�4���K� ��Nmn�_y2��93��h3�)=��iL���R�*��s�E�{v
�q�4i��E貲i���'g"�O�PO�I�i�05�# B�`���i���n�6Y��؟$�'����Ė
r�HH�ɍ�zĐ�Pu��q*n������ӟ�Eyʟ��'�JQ��H�;Z�9�d؞i�*=@U@+�I�W����O}�O�|�
תuZz|K�!m�k��i��Vo���=��I#�I�U�R� Ȅaq�Ax���+i��OΩ�u��p)�������'�j�"�O\>8��XV�x32�a����Ob�$�O"�O`��`�����=PP��P������"����?�J>����$�O��k`��?]u(T�n�I1w�ӽ|P#$@q�:���O��������îX�:�6M�57���1H�=��P��U�z��	ȟ�����З'xh1"�0�.X}�ɒU._�"�ɓ�)^�X�m�&���'l�����'�S��|��C ���Uy��mԟ�'�2�ӼUe�Ɵ����?ט�rD��*`"�6gX��D��f��O����O.ei�nW �1O�Sz�2�#K�/��\��i�!X4r��?��h�?A��?���j-O뎃x�r������.���@=}��'QbKQ�;�赃�y��d�,c~p�;�]a?�H�(��M���D $���'��'����>1(O����"����&HZ)l%�4� ����q/>���O�rm�3,�UAg �E �d&7��O����O�`��d}b^�`��c?��K�#p3�E�.�-�)��m����I~y��R�yʟ��$�O��dԣm1�I��ey�]@CR�oV�n���l����
��d�<����D�Ok�؃`
p��	>H��呒o{�I)<	6�IEyb�'���'��9dcF�"� �j�LP��"(�ڴ��CĒ��d�<a���D�O���O쥰'A��.y!�%\�9^��c���>y6�I��p�Iɟx��by�K%|���ӡ+LP�gE�nB�Ի���.6͡<������O��D�O $�WT��#'��<u�t ����i��ّ`%~Ӡ���O`���O��2�x��S?q�I4S����A�].�tBr�м]D�ڴ�?q(O��d�OH�D_�	r��O�	�|��8��DM,=j��$�KӀ6��O��D�<�"��
`�SğL�I�?�n]�~�.�CSNӚ���h7�$����O����O���8O���<��O?�X��bC�Ij\0� b�D;�M�(O�9�������ǟ0���?Q`�O�nM�,}	��M�?�0֌�.����' B폴�y��'�2�'|q��XJƥ�g��-#v��3,��ճ��i(��AFq�&��O���8%�'X�I<.�p`�-��~\�aV(!xn�4��ϓ�䓂�O�B�A(+$���nH�v,><�&e�QX6m�O����Oԭh"��K}�^�,�	e?���DG{���V�|��Y�!�Ȧ��	П��	1��)����?a��5����.vdixt��;C�&MH��i~҈��w(����O�ʓ�?��g�̨�s$�(f��)�f�	�R�p�l�����G�~���Οp����x��Qyb��G���w��1z(�0� E�#|	p%�>)O:�d�<��?������h6U:q֪-</��<�bJ̓�?����?/O�᠎�|*�"Ώ9���=YtL��BE¦�'�R[������0�����扟�� �$(R��8�n)���-#Gx�ҿiG��'2�'T�	*"�e������H�<#ִ��L��=�Si��b�xo���'R�'2 ��yr�'�$��7|���U��@��рޓj��V�'�2S�|i��ǡ��	�OD�����1V'�5�(�e��7:> ��iF}��'���'�h��'[�'��i 9X�>A�da�*��sT��)�[��°���M;���?����UX��]�0�4h[6� +OQ�uAB���6��O���5]w�	qy"�)��b@��[@θE�L�Ն5}��F]�w�.6�Oj�d�O8�iE}�[��r�Ȼ{�J	����!]Ǵ�r����M��'	�<����=��� �w�T#	�y�#W)\Y2ء ��M#��?!�S�\��Q��'��Oθ�g�ǟYv���JƧ#\�90�_�Ė'd��`�O�)�O���O♐�H�3���J�N�'"T[�-�Ʀ���;��	i�O�ʓ�?�*O�����5�S�1w9��S'Ԃ([�KsP�H��lt�P��ڟ(��ϟ �IUy����o���L�
{ب����3
����ց�>�+O��ġ<����?��e&D�7������t ���������<����?!��?q����ܗR�hϧoW���5�P$�FxR�����9o|y"�'��I����П��P�p����7if�q@��N�raZp"�Eƕ����O.���O��b@ �	b^?y��7iD@���OTxdq�Uj׷/��]Sش�?Q+O����O`�D]�b�1��&�V�u�VP�1䇁.�������M3���?9(O2�ZD+z���'+�O��1t��.|��jQ�ӲT'�U*�ý>���?1�YC�x����O~�� m`����*OF,u��Ĉ-L�6��<aF"��5#���'g��'�4	�>��c�J��K�Cg����Hǅz��mɟd��`��	A�rܧ9��eȣE٣@�qi��2��mڃX +�5�Iǟ���?�{�O*�kn�9�N�>����坭�lSq�i	��'k�I럐�z�q>�b��8Rz�B��\�݈�ir�'�\'ɤc���	v?a��JFY^�aSI�#XרY�L��M%����av���?���?�R K>��=�ဆ
Fq��#ЭJ��f�'�dEYAG.�d�O���,��������� �<-x��]�LI@Q�<���'9��'��[�P�ե:%���"�W3-����Q8�AHJ<y���?	H>q��?�̪ߪ��4�ɞ\�<��#Ʉ
M挬�����OH�$�O2�H.���S>�|�2�_�O���-�w���%W���I���'���	��H1o�o?	�����x��)1p �T�c}��'�r�'���9Q�>%9N|*�g�7b�8�R�L�6T�c�C2^�V�'B�'eB�'A(DX�'z�PU>9�@�ˤKmr	Aa꟞0_Z	mZ��	ny�1*w�����9R�`XgO����E҃ Z�YH��P��䟜���DR�	S�y
���sQ�tÄV/�,�pr�T�Ֆ'Yr�ІMd���OJ�O B�Z��l�#G��B�xL�s���(�nm�ߟ��I��`#<�)�l�ɶq�6��!��'J\����]�R6�N�&�	lZ������\����ē�?��)'X��iY��h@��n�ƨ�5�b�|��i�O ��ʎ�@�h �6���Ww����/����I͟��	?����O<!���?��'��!(V�M�4Ϙ͛�MP#Y�ߴ��,c���S�T�'�'	��A4��-u�DQ'�;-�d���{Ӯ��Z<\#	'�H�	�p&��؆}.�yD퓫I>��
*ů(���Y���I>A���?!�����]�8�� 1��ŬLr�LE	x:���0��R��˟h�Ik�˟l�ɸv�|Z���[xz����l4Pj&l��P�'��'�RU��U`��􈘣	��zC֜m����C�����?�K>A���?��MO�<it��U�p�Yd�E?@�ByIE�y��	�`����̗'�x�ᇦ6�IթO�I�b�A ҝjr%L��"�oZ�&�@�	HtIl���O���Ϧ������ݾ<�p���i{��'��	X\
x�L|:��2��B����2V�Ŀ=�n�!R� � 7�'zR�':��s��'��'@���4k��]I�-�q��`��I2;�v]�0�&Ņ�M�S?��	�?yk�O��7���0t^d3�eX	ܺ��dR���'4����T�R�k(J�ӄX����6�V��M�T�
�����'p��'K��M�>�+OT\���
n��5��gR�'㘰�c+��Ԏs�\��SyR�	�O����]�����Ǉ|�R�K���	ן��I��r�;�O���?��'*̴��
w�֬;0I����yX�4��[��S��'�"�'��1A�۬Ko���g>}V"Tih�����5baA�'����T�'�Zc9XPC��U!_Bx�{�G�3	���O��Ђ<O���O����O����<!��٥��P���H�sS�&KcbY��Z�@�'��\�D��۟��	�u*���m�%`_ ���FY�z`�%��`�H�������t��dy��ia��S�my�(@ӊ@�<��#�Ѿ��6M�<����d�OX�d�Ol�x@7O�D1�T��:�E#N䰙1@	e}R�'��'K�		�"3�����T-�2���O������>\o����'u��'��Eڴ�y"�'���"�8�b[����V��l�ݴ�?	���$�����O!�'��d��-�U���V��ݳ`���4�,듞?����?A�� �<�)���?� ���D��x�$�H���-}�y���i��	�9�l�0ش�?���?��'`�i��'�A�w�������4C�F��aӆ���O���6;O��$�<���Z�/��#�b�/a����sT��M#����?9���?������?	)�Z|i����M'P�v��s��U[``�E}r��	�O1�
�$�( $ �EZ�1��#І��!*@�oZ֟L�	�0�da����|b���?�����
��d�\8��1{�!���OVMJ��d�O|���O@���f�J���+�WL�M�pm�d}�JB�_c��Ay��'s�'�  �g�ݠ�:��'���q��5���.񤋂|��ٟT���'^�̙  D4�R��f�iR�FH�	�FO����OГO����O@y3�[�{G����U#��lr��5^K1OR���O�d�<��`�N��)^�!T�dh�C�y��(+ )�F��'�b�|��'�"�����D!�\0zBMo������|���ßT�I���'7�<H��-���31� �D6�Ђ"�5H�Q�ش�?!N>���?qҨCy�qjf*���r|���$d�:Xelɟ4�	pyBIѹ5������Frbi�K1��`. �.Eʕ�\�	ΟX��>j�F#<��Oxw"3��t�qc��	�H�۴�?����-b���?1��?��'���-#G�	6[��F�ڄ+�@�0C�i��V��2�:�S�9C�H�P���+T+�I�g�?im�7͚�5+*�l�ܟ��Iڟ��S���|rD�H5F��e�PO�"є�����Sכ���3�O����O��rC��=#2��,[� �r�l���i57��O����,�<�/�r�$�� ��'6bj�`�a�aKT��=�Ot�&?A��Ѩ����-D )�6I�^�4h��KO6�!�$V�:��ih�%�\�v4�c�����z�&W$	��J� �)]E����ç v����צE�P���-+�V���dG����%j.kڰ���ƭ^^4�@�ܰi֮0e��7܆tΝ�.\�3En�"���q��iӕ��<E��w���WF8����1SuHh�l"M����V�@�n�↊U�GC��ā3KĘ3G�O/c�2�'���d�'�9��8W�T[hs�C�W����lȼu������ʮ2s����H��O�XtF~�+ʳ9��XH�k�Ǌ=cK:5"%$�,R��!Y7�PK�iZ�(;B1\h�*SLp�ORij��'��[��#�GЅ]�l ��*���y�K=�	B��LH�T�^� ����K4}�Z!���0����4+��rC@��P>���똣w����������'W�Y>=�u��џX ��5�����]���,���@���0f6�2���-�b�	$��?�?�O�哰H8z�񂁘��rm�rAΙ@c��'Y\5�A#���8�
9�>�J�����t	V���00��Ц�'}b��?!��h�v��>y�zeJ�K�6}����+�H�!��R(,_.TY2	ՕE��I�6�Ⱦqax�N5�Tv`m�2�S2Y\�qP�!�K>��Qe_������<J�L9G�$���(����(.b�3�Ά�+�r��aJE�wў9�!�Y�������5ɋ�_�Bc>�O�YX��K�9�,�����<��o�%�t`�_�h�����q��'�b-�B��8�RiI���)<DQ1��'���<R8�4�Σ=�'��H��`�d-P�8�1���V~�<acM!T| �Li��� ���}~��#�S��[� �Ƞ�`y�ċ�FPєN�odd
�	ҟ��	ȟ��I��u��'v4�� 0�Κ�i�^�6DS�,��p�Ёɀ�r�7)ٖN"���I�+�� Qal�1��p��Q9�@b�@�	"��!"��<���s"O@1�ɑ�s��
�Ey�P�tͼA�����柠E{���6^`<@���KE���e[�d!�䃼Sw^� @f��r�(i�^xh D�dMI}bP���cf����Or8ks�ΛV8왩!���N[�Ћd��O��ě�f�.���O��aLn5%)O�^6`�gdɫ�"-ٲ�ތ{����d�9I@l�6�'c0���ȟ-H���[�FpSQC]��ZPZ�R�|]"!�g	Ęqs���D?�������>�� ��Z�2~.%�7�)@�1O �����Z�y�>V�l���8z�!�DL�-p`�<O�i��g�a�(�ǈ���?E��'��T۵!?,1́�1!�$4]޸C�'��btE���𓠎�~�t��'�Z�˅bm��f��
x�<�	�'��P*���5�\(��%7t��![�'�Vq�˃�5�Ha��$�1s�. ��'�pۅ��e&lѴ�L�e��)
�'��$�"d�w���[5N��*��|��'r������0>���DH]���9�'� �r!O4P����l�2 Ud0�'nn\�k9q�\��6������ (��BW�A��+%S�@$�$��"O�%�4$��\�j�4J��A���"O�m��,�$>���U(�%KژX��"O�p2  T� tX7hgq��D"O4��R�ΪlD�Y`��L5���"OzHbE���l�b �B4h'Z��"Ol=
��2x�eڐ$/aê���"O�M2D�VdP�%*E�E�n�h�"O" ���]�d�B���O��'[8R$"O*L����K��L9e�^�iV�exg"O�}(��;+V���-�?M���"O���O �4c�X����9�0� �"O��ԫ�R�T��e끽3�H���"OVl���3���)�}��1��"Ol�V
��y�����&�?[z���"Ot(�MK�f;^	Ps��=zT^|2a"O����MPmn�U��d�&E8}y�"OLe+qء(�`|���ĝ�ru�E"O6��`$*x^f���ŉ�"�6�І"O>�VB��PA~|�ÎE�J�f�z�"Od�*�	�mg�!:���(�"O$0x@�{�n��THB���h�"Ob��P�N�.*6��g�0`z��	U"O�dSG1v>)Y�^sh0�5"O~�J��u����gP��ё�"O��;�#�.7u܌�d́�x����1陿75��2ӗ�ԫc3�g~r
"�N���P�a�p�.�"�y������R\�<�ħA��� � A�5��`�5&���d�ME<e�IV
.�v��� �"���+�^3X�	߄P ��W8-�0չ� F�@B�_�j���#ɀMy`���؇ ��b�����م$��X�ժ7�Ĳ�A7��
2'�Z:�,�ȓR��I���Mb���/+ ��iu
�� G�!�'H�	��𙟔2�C"`��	��,���S,7D����&ҧv� uy�����4�>Hf2]*Q�����D��@��	R� Hk�,����=�azG�1B�3q�Μ�y��9"�$�ޚ1>�1�p�̠�y¨�,F$xH/
�x���WJݕ��'��=��Jܗ ���"��)��VF�Z&�	J��qӵ`��-S!�D��1#�X#�MR>�N��O��~a$�[�b�7f���"_��"|�'���˃G��!�҈���]�nj����'�tܺ#M��`(��AƁt���NƯ?�Q� ���0>)`�@;��l��Gr�t�; k�s��l�#��N��=���x� �2#��X��AZޜ[���{'L-D�P�0»Bp	"K\#M�E�6�-�I!I�e���7�0"~B+ًB2�ڔ'A<	���sC�~�<IL��*�``���T;`)��o�O�<�Wk5Y�x�@�4`��б&@u�<q E�#��	����
V�d8�%�x�<�FO��X�P�'�"�b�ۀ(�}�<9d��_gHi��n�^OX�+1�
O�<	a�ǘh�HIHaM�*?ĔK�CXf�<��ύ:�5 ��O�˜����Ql�<q�Ɲ*M�F��+ۢƺA�2~�<�V �ښEKR�ҥ'�*URg�~�<��?��I#���p@|l�RXn�<� HS�T�:���f�Xm�3�Ip����#�	���,up���U7iYvh!ΐ�9��B䉾h��-@�kRY�D�#��b�[�T�c+�鉊�II �l��e�+Jt(��o�>�!��ˊLZՍ^k��)0�͇\�8*��؄]�I�O9�"|�'��<��HC���k��X[RPm�
�'�z<�F��k�e�F�
(5(5�W�׃~��"gA(T����@�!��db7	;���Ù�5�az���=Ks����˺!�
K� �ED�
�*0��Z��"H�Ni�"O������#�6S�'����.g����J�`��	8��	+Ā��֤�$/��ǈɇ]@!��2�$B��m���ac��3��)�(L���ۢ_v���8��)<�$�:���'�2G)th��k�!�$�2z@��j�MYc\�ѺJ^&��䰰�ύF]��3�m	�k!�d�%].�p<��p�����'���:��1��m���#��{Yl��с�)ml����<�l�ZѦˏw�lu���G4ulN��
O��Di_�,le���4(fXa�����ҭ�-��Ͳ�,�<(�i��Oq�DM�vM��R�&��oB״��"O��"��8|K�E�r�1`Xb���`_bڰ���lO�mw-��]���O���	�S��F�=dz]H�ǖ!��B�	����d�;9b��x1�
����t,X`l�y�ʓ)�9�Od���,��	���z��%@*��W�0*����ĳp<> 堔�2��PS�ϨI�vu���5sݰ���ř ���xsfG�p:�}sW�OP�T`I��p<���.,wx"��C������[~B�"x��;���#v�Qہ���?��hؽ2��'W���K�+�T���C�yxqM�H(<�ǀ�8x�t�g ߧS�v0BAK& �Y���Xw~,��hHqOv1@I[Ƽk���"6�,	��\�4e�hx�d��fN,�m� "�	��ݟqV��ŌЭ4�VA"��`�ɍP^�8$��k���c��L��->PH��Bޗtw�}c�o�>C��=!v��#Tr���-ͽ6_X�ٵ��p?YЯY+���h���,s��z�FZ�5j�L
r�>Q��cV��I鱨OC�'"Y�&"���t�sb�ўAyi�'�����D�g������Q�X��Of8��dא\L����R��P�s�ϟ?%ިi���HW�(��y�����sV��`L>$�j��E$`�h5o���I+Gn� ��L�Y�ei.�����Ls�u��%,�; *^�yh��yb.=�O��I�i+D>�hVOS�E��x��0	Z;~r�iTK[�e���'����'�I��0��݂J��ŀ��O2���LJ�G����#��@UPa��I�.M��x d���	P�@N2�D�2c�!�ddۨ;�ԡ3s�ź$?�-22�6��eB
SZ�I�K�B�' l�V�՞��bŪ���ʅ��i�L��FX,��D�L�A�m�R�žUaդ��e�1����P`e�6_��!Ǻ�C�I�|L�)5�S9p��8�gP>���ɔ��,�A�ݦ���W�|�'Eh�O���Я�DHd�#�H�H�e#�O� eN}*\���WS�X�� �;�I �5a8�x1�<)�.]`��JG8�ݓK��� �ՒBV9R$a�4 ��R��6�_f&�85,��HZ�(c3�-��n��p�H��'vȮ���*ai(�Wi�	B����(v>�#���CPjtxP"���	;f�ޡ; �V�G�"<dF�6��!��ڦ�>=cե��K�nI���C���d:�.4D��XFg8f�E���L�m���s�%���a�)O$8z��dk~c>��>�%�V&x�y@�
@AA@TE<�!�F�:RR����n�|�BwhϮhZ)�'-ś���"�˂lߎW�Z���:�v	0�-L$�X�6�����x"Ȅ�p���f�˨vzRu�C���O�n�p���[���2Bi��OՓ(�N��5x􈛹��1yr󄋙Kw�0{vDAi �����j|N q��\���y;!��1T�!��G0G�z4�)żp�D����|q �W�\R�)�'.�<��𙟜1E`��%׃!Fl3�.D����@Ť
ʜ�0WI�r\LhR�'ȩH�TM����,3$M#��'�t��G/״D�\�fC�2u�E�	ӓ<�P��G��O~����k��>ȂmJ���2X����� �9�� �+$I2 �
��4O�i�<��	:t��hS%Z��|B�%�JZ�Q�t�� o���S��l�<�)κW�y2��:����b�	p⭩u폗`�~�VcN�|�'f�q� ��1�H���H_�b����'�� �ц�V�H��r�@�I�-��4@<�q!��P��ד�Z�։ӎ;F �k�)�D#�-��I�٬!%f����J:44U)B ݦ���¢ D�H�pF��uh��t�O/b����=ғfn$U:����tT���-bZ����X�'����𬎎r���R� �,�dE��'C�h3�$X�Uପ��Q�U�}��'�8(����{K��Z�����"@��'j^;T�@� 4tb��
!&Oz��	�'g�%��T�lJ�c�����x	��� �UWg�>Ac�|!f�J 11���'"Or�A HL�mt4�B�Ŀp-x �"O,I���L�FJv�4�W-$���"O��R�S#z�d��c�gxt�80"O�ՓUO�\�*B�bեOp��w"O:������Y����a��#w>��"O��
�M�b�#�������"Ob5SSgʋT�0}S��
��Ct"O�M{Ċ�R�4�P��K1�Ҷ"Oj-������2�����h�"O�TI�E*6ZHԋ'M|^�Ӈ�<y��t	����/W�p�1���X1g��!� i��Ks·�{�읣��,��( �ͼ0�qO?��
�\�~��P�x�^�'�!��Yh��I�E)U�/S�q�0 ��D�-N�b]�
�#~*�P���"XuB4�L��T<ą�I2"B%��7O\퐒@�	ǚ�+ңϭz��c�"Oj)� 
a�d�VM�1w>�`�I
Yz	C"��bY��h�h��.?r7�%#FAb�,����'��>�	����wdƼ]py�""6V�`�8���Ov�"~���)h��H���gCTY4'O+�4��� B�|0�L0�<(!�XY���6oٗw5h������F>�}���r��>�ՠ��AU� Q⨺� �V8�h�#��\S�M�t'��.i^���	Іj��O2!����ȟ<�����+i�ay���au�s��)r��}���i� �|k DV1BLD�[І��A�v=A�`�u�S��y�ިjд��v��:MP|\c��y�½��aj�V�@�ظQ0!ެ�y��ң#��]�b�"?<�X�#��y���C���G� �а�k���y�k�!aD���@�+je��b�(�y��R&m��ʢ�K[��A�݌�y�O��!,n�f*ݦ�0�g@��y2
+�^��2��<��7n7�yRo�!=���e5:���#���yBC���p� �F>�� 
/<�y�'O'S�*1 eƷ	�J}�b`���yR#��?+.����ON�ʩ!��G)�y�cL�tN(��-Z<Ux8���yr��8u!�I���*�<���ѻ�yc�M�HM+�l>�a�4E��y�D/���R�hſc�N���	 /�y2��}��� 2�
�dǦB)x��ȓ��ݸS�%�<��� k�&���+ !k��5?h8! B�p/p���tZ�H�T��"y��p�)�}@2I��u4@ҡ�	p' `���V�dU��y��Ы�G�Y�\����*_8���R���[s&�7��,xV��	7�̈́ȓGm<��_�AQB�¯	�Q�ȓ��@�*cȂy�3[�H~��ȓ:TLQ��p��86��)J�޴�ȓv�H$8�eQ!o���b*?��}�� ᘈ�6B�'��\�vb�c~d�ȓ,�
|�"��8Wۄ��A�Y�y�
�ȓ[�U���H
B��,bɯ�l��ȓ'�ɣwʐ�'�H9��큠�U��5��ŉ�-A	3~���m�yL�݅�x7p�H��@���ʂϖ�]�� �ȓ.��(R�ͽ:W�=�LB����ȓ	p���gD-#+���H��;!�D	�`��iť@�L�(<X3�!�d��w��8�U�a��,�¬E�9v!�$˖j�lb�	M�8YX�L05g!��  I)��E ���`H�l߰y��"OD$�p�	�]�����ƒq~-�"Onl��Ns�ܣ�
Mvp��j"OꠋbB�=rS�lG�)A��-"�"O��a���|}\�#P��
LѤA��"O�Qb�MW�E	����L3�HQJ�"O��$�K�X��3��!ET�"O��`��Л�V1��-`@Ե��"O���EX50�˴�x,b��"O���D�7�Dt��A�x�"O�Y1B��P� ���Y�&��(�"Or)�CnO�'�ιz�N��9=Nd��"O�12�]$����F�!�1��"O:U���,"H�����*-��"OƌaELX��|���ϰP��� "O�Mё��|_��Gᗘ(�:�;E"O0�I�(^;n_4��� O�4��X��"O����I�q~��u��4��i��"O�3���v(W�\*ԩ;!"O�	��V59M$� �I�8�X�"OXl�F�Ն5��%��S# �b�[�"O��Z&�̈́.�-�AՋ;qf���"O.q��M�%��dA�F:}D���"O�m��O���F���e	j���"O��!/5\+
�ʄ"�0�\	�"Of�8�B,dnr�����&��)C"O�I�S[����S�fT!+ֺ�iF"OB���L׌$�u�ыx��j"O� pu��6g*�����)a"O��R��l.��Qp�ڵ4�n`qv�$4�z%�?!��Bbg�u��x{լ/D�D"4��(!�Rz�F�3Dؖ6�7D��§�U((���ݧ`>j �'7D� �ǁ�a�@D��*�+���(b 7D�D�q������e�&z����W� D�xqt�ҫ6㈐˥�
h~��cV�)D�TP*����\�a@H=;����	2D�X�Š:(�y�/H�4R�RM/D��2�ǘQ4�IU �Y� �(��0D�j��$8"X8[�퍄d����c3D����PN� �z%AO�I_���3�&D��rTaX7yy�8C� ��ӡ$D�lVDH��5x�L�!N͆	g�"T�`k7���H�K R��"O|�0r������p��+P���"Of����9w��e!A�:4���"O��R�
�tĒ��Q�.;��#"O~=ZS�[�¨I��E>y�c"O�c�+I��D�U�Q�0	"O�9��k��0���B�e���q"O��Ze���b�K�SH.�S"O���ć�	TJ��Kw,@�
E<�E"OJ �q���;��t�Ѕ�*@ʹu"O ���
]��Bd�O�@��"O�d q�X Wk ��` ߪ<h�z"O�\X�!ɥe��S�@�@I���T"O�{�e� ����g�-|&�$�w"O�͛�ʘ �@�!�	�ej���"O(
�P�/\�wkC�	V1�D"O Yz(O3 �ɡ�lދ^ps"O��Y��C�	�m��b��<�xh(p"O&��r�
2�~A@#!	%	�v1�3"O��!��X�7Ўtd��-���"�"O�����ݎP��sFa�5��S"O� ��j�ހw��!��+}R�L��"O���ӉNz��f%D#]�B���"O�L�Յ�rX5A��(@3`t�c"O���̤q:ii�f�&@h�s'"O�ǣ�%���*WO�@�@�"O�����T�,���$��$��T"O�m[5�� h��i*T��0�<\i�"O�Ȉ�W�+��Y��O��䘧"O|�5!o<|id��$|��zR"O~0b%�ϓ;ܘsL3/z,d�"OR�0U%e��M�PJ
K �!B"O*X!��{�f��	�l8t�h1"O�q4.�0m\�b���0rҌ;�"O�Ј��֑X��`�'�%O�
��"O�P󢝀�p���D� ��lzW"O0Q�c,Pyh���޵��P��"Odhk�hSij.)�J�^���"O(�@�$��蘷j�� �J�*c"O�`z�V~jp����:�d���"OX����k�Tp���`�
� s"O�3ƪԛ�y��iF�(��<b�"O��S���K�Ψ u��:�hP�"O�hc7"0mk~��#��r"OB�[�M�j�`����e.J�"O��Ӧ�Y=g��1	�`I�d�PȻ�"Olt���`ɖo�~�LUJs"O�!f�͟v���h��k���e"O�e�6� ���Y'��=x"�"Ox�	ͧM<���q�*��["O�T��LZ�8e*�>�R�q!"O���T�'v��z��[Xr�=OB��d[-z�eQ��;q
P#�o��D��~�\�d{Rd)�-�#̞&��e`We;D�(�Ջ���SA	�-@��� ��5D����)��=�lL@7a�-6�U��1D���u��9���bRBڼ礁[&@-D����/�r�l2�Y�hQ0#a-D��R���W������b��)D�|���ҀN�x��l�3a(%�3A2D��B�A}f)�G�� lV����'2D�pI�
E-&of���;�,#t�$ⓓ�н0���3�(�Q������U#!򤑛r�|IR1�[Ed1.[4k�!��Övf��3%AH�K�� �tJ�&M4!�d��ę#8���bIҳ5#!�dW'�
 S,{$���嗺�!�d
5v-��"�\M����K�!�ɧR�r!��·:����E$Ϣ~z!��*n"BՈg���W��H!̍\!�d��4j4�Pg���6x���q�'BF!�ݟo�^`��ȯQ^��cղN/!�d�������y<��1DM^�f�0��I�4ԭH@ߖ5P�iRB�	xv�-�sh�	EK�С���@B�I-���;�b��=Ʉ���m���B�IO�\1��QbF����!"j�B䉄��䳴�,kV2� � ��T��B�+:ӈU�� -\+��עO�B��'L$*rM;ڍ�qn�8	��B�ɕePZ%�	�+c���KW�0*۠B��-5��9���!�8�B�m�A�fB�ɋY����E)��qC"���Kʄlq�B�ɃX�݈Q�f�ڵ�̫@�
C䉾-(`Z����,�HP�\�B�)� T�qT�3t0���_�JH��jd"O��f�\!�Vp�|+�	J�"O<M�ń�,C�Լ���N�
P�rv"O ���]�B�RcB�'|��L)�"O4I��B�9�Θ"�Mg�l0� "O��He"M�D�����ڞ�r�1c"O�;��؜2�2�(�i�1�<,��"O>�ڷ�ݛgP]k��3R����p"OD�$�ՔV�FM�7i��|��4)�"O��[��·M��D�w�D�"O����j�V� � \djy�"O�TP#
�:<~4H!�O�J45� "ONZ�b�$}Z����5�P(��"O>5pdfN�~�m��47j��Z"O<j�ǡ_��	@g�4Vc  �"O�G'20�bp�3�M�TDy��*OTqf/xaDÄ�B�~�ѹ�y���3|<��q�P-�`D`Ț�y��I�d���T�_�k0cϦ�y��DS�f8q��~�u��m
��y�EL.}��ٳFN�}��Z��_�y��PF��v`��s�j4����*�y����>Y���_����Z0�y2�/B7(�+G_K�:�g��y"L_'�8�3�d[/H���Z�@��y�=P$�c!L�A�&���A�y2�÷xZqX�/is��3D͡�yaCxc�� ��l�V�PP�<�y�D;��l#���;*��,߬�yb_1U cgLˁ-�dH$D��y������QWQ�V��aP�ݭ�y�kG�6�yْĊ���3�*���y@Y�~�Чd�b��Q�U���y"��҄��� K4W��|1u�%�yr�ݠ,Yt���Pf�@ !��y�n�%�P���
��8�7@�y�㇜)�p]�>2Aǩ�,�yB��X�l ����@��W��*�y�@P9[U���ń��N4LCG��.�y�`͕|���s�DG�D�h� 
�y�	]C�-����S"׊	�yҭ�/v�(֥�%@��J���yҬ����3�ş�
J� �M��y���,��|�� �,����C���yrć	��ݓ"CK�>�0�y2W�D��1y��W8j���7�N��y�#��qwhpY*�5S"��b�
.�y2ˏ)����%D�H�l5r��y�!����ճw��O��u�%H��y�mm��yj�O�7LNpQ`!�ө�yZ8u1���ZC����i���ֽ��'R��B�K�(aj�(Y���"+����'�h`;���E.1!�MX4 �;�'��YoO�`�ڕ��i(J\��'I�<D��ju�S-I�Ɯ�+�'�T)�@E�&�|�$�J���2�'R���a�5h}�� V�g�4�!�'|�JC .ց� �^k\�r�'��yY� #��D����*��Q��'X���A�l.�x�''�y��'�L���#Z��1"Wd̨4_���'eT�R؇15S�m\�u�HP��'�r�Y+Q�S	^	F"X8 6P���'֤�1�=j6ȸ%�A��@���� L�[����@K�$��"O��g���6c�rXf̰��"O�Y�"�@ TP��e�'A��ʒ"O�q�u� �J�d����3�Dyrs"OD]I�K�2w�# Ҳy��j�"O�s₈��B��1�ÏL@3"O�(Y%jg�XۀN�';�kF"O�U�s!�Ӭ�A�'O)s�48 �"O>��Ye.����߸��d��"O��7G�*'�]��F�0՞}��"Ofa@R�ȪY�kS�T�	��Ua "O��a�Ɩ:e�9��Ȅ�tT�I"O�R�CE1�XI'V6nG����"O��p�ɝ f�`g��R+f-{�"O��`�K�{X��.tQ�"O��1�m�,W,��T*���~��"O~p١�ן�&zGC�-]���"O�h�l�%g��T�1CK:�$iY�"O��LU� ə3b�� �U�"O��*�h�S�|	$b�BC� 4"OP�*U�>z�֍�0jȆD�b�i"O��U��!*$�QCh�#2Ӓ��"O�0���S'G��ೂ�����zs"O�Y��$G1��H�#&D%0�^A B"O��́<)4���DH�Df
��"O�X��%�:�(H�J��\^��"OHX��H�1 ��(Ҷ1\Z��"O�����sb䐑GH�7kp�x*6"O<|���P%�	���@ F�1"O ����<WvU��FF�M����s"O��+f��*#�Yʦ��~(��"OD$�g�U�_X� K�jE6qz�0)R"O:��'�J64z����˓d\T��"O&E�CR�������p"O��[�
?`��NVrE`���"O�
m�`z��-9� ��"O��xci�!S �����H �Y�"Od����_9��xt�>H�踛2"O������@�U<?�>I�R"O�e���Z�x\��҈6F�qg"O:����ݦ4I�!h��+��yB��n�H
 ���=�d�pW��y��X��`9�7�`��&H��y�C��j�6a���!2b	� U0�y�ùr��B�
	BYhT��F*�y2��=w��8T㈐�.)��y��t�>��F/�
�\��ۡ�yB @�ec13B�
�2|C�˔�yr�/@�
Żc͎�qP^,�C��&�y�FS�Y�q�5˚�hQ��2	�yrI� 5��RSL$1؁̜(�yb��.W��!QD�@��|��ʋ�y2 Afj$�; �?D�4�h�K΀�y"*Ģ ����S�6C�8t�0`.�y"M߆ Nذ��n�)f����� �yB��uK�yy'LT�~�\�SK�y���M�bգ�E�2d��Sk	��y�CX{9�Di�Gہb>,�abkR�y2)#L��
�(m��j���y��f�(�(��3�P�I�����y�ܩΖ���R�+Sl
�+���y
�/o�>h�􌜹n�dt���y"�h-�<ڀAߩ;v�2�B�y�W�uh�Рт�6kD�j&`�y
� �@��78�DJ�JͺGc҈b"O�� OA�Cd��HO�XIԼ�b"Op�k��W����E���p<"�D"O�@�dݒ=P�ig�)��Y�"O��٤�<�|P)��R�{Ux�@�"O~p�B�Wm�0-@%m�� 7b�S7"O�-3�M<C��Ѓ��{4��"OR q䉇�!blx�����O�^��s"O\�[bF��s���t�ч>Q���"OHp��Q=����G8\��"O�80L3T$&X�5j�52J8�i"O:�#�ʖ�><p'_�]as"O��0g�ʋh��qS E��6��(��"Of�s&�۸)ì-K�C�pB���"O�mp��G$��$� ȭQ��1�"O1ҧ�1$qD�ω� U�b"O�Z�AϿ����N��So�e��"O\p P��*.�GC@=~Q(�ZG"O�ي�K�8+
�9�cN�GL���S"On���+m�ä�EWJ����"O~��'�A�����-��h6"OhIz�@�1c�����kn� "O��@��P#葩tkX~RD��T"O��c�R���",׫9p��zS"Oa�Ju6��t�ͼsO^,ز"O(�۰EF 5�yP(A9E��	��"On�Р��=����ג���!"O�Q�e��$
(�SV�K�10�U"O��`+��w¦�8𪇱y��0"O�@G-��r���d��d_`���"O����N.w7hZq�Y�e���c%"O�bPhD�i�\iq�D�`��ݳS"O�x֥�Hp��Ҹe���a�"O�l�6�X***�� &M� |J��"Ov:�C�5�)�n�"i���C"ON4ň�^�R ��,T�Mq��+D���T�����&�E 0�eQ�(D���RM Cv�Ku�A�r�+Ť'D�p@"�<)}�1З��J��u+�k$D��y���� E�X�gb�d�R�)-D��ҡɟk�5@`A.v\N��֡%D�Tۤ���t#s,@�n�V�)�i%D��5��(M����D ����!D�ܨg�����-�v�B�t��زM<D�\�*�jX0*c
�a4���Ѯ8D��21�ğ	���z���6uSI8D��"Aɕ)�˥GȽ�dؗB6D��(�oO�[(L�K�b0O���Ď3D����'o��8Q�B?y�SE�5D�4S��Z:�%���?�rm��/!D�08��6C�樃�*��I�@ir��>D�t���M�6�Æ6z| k�*;D���b�Q:(������p|@eK&D�в5�������?_l���J0D�����J,P�\Q�����ZE�/D�|bu�:�<�اk͹�����.D�P���
KΡ����0���9�9D�\Y�ǆ�RB�Y�%�A��$f5D��i��ٞL�x��L�;i��K2D����?[������$���%.D�����_�	4@P���'0��h�Ѣ,D�i��˲�j�9���z�|̀a�/D�P����&�J��ߠ^�\ms�1D�`�2+"\��{���j��x���<و��3� lPb�bw�LMI�؅|N"O�`�U&�*(րT��`_�Re���"O�9�'"A.P�B`�5�Q�p4DY10"O6]s�S�H��+�ƵD2б��'`R���eW�U:b�V[�]�C\1v!�_+΅)e	ӑ|>RY"5#�9.�!��A,A'�<�2��#'�y�0%5C�!�Η����n��f��AQ��=�!�d[�H����b��S�v��Wb�!��1'���<W0��p�!���Z��}��+ũ#|4)*��џtF��oȤg�����.<s@���Q�y2%�"���#�aF�2��)�s���y��ۥ	�ʍP���%� ��s�+�y����.,h�tmΐ-�p�b/�y�a�)1����H��P=�b�_��yb�B3�<���
�Ax��]1�y�$ͥx�v�9�LN�x6��r�ܗ�y�4Z4�7M4i����&hH��hO���$�Z�Q(#R+s�P�(g��a�!�ؐUd|�%W�K��(�Y6ў%���<�T��24�$}��\8$�֯Y�C�Ƀh4� 
4�٩wx�m� �ԔT�^C�Zі��f��"n+ĩ;�ȑ=��C�I�_�F���n(J��(aR	L�{��C�	%.�P�y�/��
X~����K2�C�ɞ!Ѧ��q �M�� g`�#5�C�	+i�^X+rAK�$�Dh�I��B���d+�S�'���J;��l�RG�'9윚c�kW�'yў�>i��Ε�,�H�!!m�{�j��!*D� S(L)mc�!0J�0&���-D�C��0Z� {1�/|��s0�'D�\��lG80)|E���_I��E`b )|O@c��fG��?Z�� �OP�^�fX#�#D�zF��K:�I����SN�CrA"D�\`�)�+P긃��?�ƿ<Q����(��]ʧ���^��	M���*T"O��X7ok
��W	�L�6��&"ObycID��[�(�2/ǈb�"O�Iq���s�̙C7.�>M�U�"O��;�m����k�*T�=���a�'�1O,�{��ğ^P��p��?y;��)�"O�HZ2�^)D�,H��:3^���"OفS+V/[�rB��5���E"OriX6*J�O���t/9�0 "O�XE�� E����g�1P�Q"O�͡��ѶO�PT���Ѽt�=�"O
��AO_����Q�[�g���"O��[��O�o�BT�҅p���z�Ify���%��<�  �N)	ҋT!p$�B�	�L�zd�树�$��x��N��xB�	��je���Ȣs~���$�M=hB�I�a[h�c�̆�fq��i��L�U�2B�I;O[tYQEㄜn���h�bJ�2� B�ɱ.Ĭ�R@øS��
�$֫x��C䉅sBs��3}��	.@+~˓�?Ɉ��	��Vf����N*y��	�oтE�!���"�8�g�]Rv�9I�o�e�!��,~��zG�^8`c �����k�!���	�m<{CMÇ6Wx�q!O�9�!�D I��4
���|U��`�9I�!��5w�茠FeH�=�i��&Ղ}�!�$�w�}�(� v>�T�V��BW���'��>��
(�������A�p���B�)� �I�0��&UU$ȑ�ԓ.�i�r"O�}�q�تS���qEВFR}�5"O�=x�,��T�h 	��3rD���"Oj$���T�d^�
 �� �x�'vR��B�BC
.����9_b�-�t/'D��P�����Щ�p��8<O6#<	f!�6nt���I�\]��`�p�<y��6g�3�-P��(k�@�<YՈ�Xǚ��*�'!��y:���@�<���Ǔ<!0:R)ŊS|ڢ�e�<V�� 5����s�|�(q	�b���>O��ir)���[6��02�X��6"O��j�����1�`�LL��r�\>�/T�O�n,Ə�.l����!D�Б׏��� ��M^I��F�?D� �c�����A�0���E��yUC3D�� �"X�o��"En�ux�ax�O#D��7�K�79�ڰ� dE�q�׆6D�@�W�Lg�J�s�&<��� �3D� A����NȨ�� O�����+2D���m�oN�m;Ud�����C%D���F�Vk�B��!W�O@��+�&D�����w&VPH4��-�l��P�#D�����V�z*:���� 6*����Oh�I�u�U��˻hX)qH��k�C�ɦ�,M�� ��y7X�Yr����C�I�<�V�C��%E4�� 킨j hC�	�Z�� �`��NYl���]��C�	1F���H��B,0@�P�v'�q �B�I�3��J�@�p�R�Qwe��z�B䉎5SLБ�I��E��a(&��^���:�I�k܎ ��m[�z)���F��ϊc� �e�ya���S�&�qu"O��e��P���$X�b�"���'��xB��ېA�H�g-�9,��m8!�-D����	�%G܂����_.-����++D��۠k�%7�X�QDR@����t�#D���&��/��I�V�U2��\(7�4D����#W<��3 �0+��H�&+2D����Ċ7,�d͑g�T"#p�|zo4D�89��3��ظ7���&�qg/<O�#<�NQ�~�d4�"���&UfX��A\y"�)�'L�2�Ǉ 9�Q M�?5��ȓzR�W�+_t���#�0�MS�"O
�-�)J-���Uc@%U��d�$"O$L0s��"=j����=�J`��"O�	RFG�%J�qVU��yҏ�$v0��� g
X�)�����y"-�@�&@�d�щ|;r�Ȁ��#�yB�܅;������xgx�2 �^��y�m|��\�W(u��Y��%� �ybf]&���7�M�l�,�Q�/L�y⪍.�]�uh��d
n�Z(W!�y",9;B��Ã]����Iw�@�y"��=1�5PF�5���2G��y�E�!<�<�(S�?>(�Rgd�,�hO���)�f��U(���26b��f@��z�!�"|���&[�a��kf!��_�%U�Õ
�28�~L8���Kt!�:X"��/XZeP�L#s^!�$���6%�(5b���@#0R!�䌁/�XqG�Ь6��#�2&M!�$f���XE����x�GW <=�O4�=��B`�M�!�8x�*��Ps�A�"O� ��I��M;#�9�v�ֽ0r�E��"Ob�2 �KH��q1���.]�I�"On�B�%e��J����Hu�<	�"O�,��'�^��Y�䎞��UQ�"O�X�a��>R�;r�Tr�0�"O(l��\5�z� ��sK椡"OX8��)bQ4"Z�R84f"O���cfH{L�A HЮH
x��#"Ody�)�I��{r�3b��hT"OX�ʥE� ���wQ�R��xK@"O���UGI�����B�1?X�x�A"O�����
�>�ɠW-��"WΝ�"O�Z	ۚ��T@�KT�;8Xpd"O0�CD�Z�r/�����v�0�P"O:�4I 9��h�q�4eta�"Ob0Ѡ�J�IR`JF��&`��1�"O´�F�Ðlhf�`CЯ�l�@�'!�'L��'"��,�4��&�pq8���"
*���ȓ�>X���?^�iH�"����V0��#�1Д9�+�$���ȓq7~��S�^!�ԩ㠨?*�h���ga�Da��ǳx�VD�� �o��Іȓv]��#�=A��%�Jm �ȓ~Y~�X���L�"�MV�!_^���W����,B1:)�v�X-p��ȓT���b�h����p�D"ؿ2Rpd���Y�k���5b��1�ņ:���ȓP��0 ��տ}#��{-ۉ'���mt�Z#`�aY+�5,�Qm&D�H�a���&)n5�5����pA@�8D�pr�t�M� ܧkԐ��B"��؟T�'���	G�58�PD��j�0	Jt�R;�!��,Q�]8RW�<ܴu�Sb�+O�!򤄇)��;'(��qxF�#���!�$Uf���?S�A��j���!�6y�B0p��0N��P�Ȍ-i�!��ow�)S���\M��H�'��:�!��1��h��\�B��3�ّ�ў��ğD���$'}���eC<,*
�"M��yC�f�t�b1L |zB!2��(�y"�K�\��Yu��<D�����y2�:D��=���Y,�F�۠� �y�	�Z�ݲ���* ��ӱJ�"�y"��aw����(@�p���J#���y��̜7��5��X�lÂ1�[���O��!§sx�M[qL�25��jB�+t��d��v\�ň���!;�\�"��P�aT��	]~���Z��h���أP�@��$LK+�hOp˓������U� ��G�� ]��5��"O,�����!PY��)K!�V��"O\���o�1��a�	:�h"{!򄛳:`�5��H��4��ԅHS!�9}.2�A��,-��\ELʦ�!�ÁKl2�!�ʙI��\�%Zd�!�D����@!$��>рm����u����2�g?�F��X������,#�Y���j�<�P+�Nk�]8�޼0u���]d�<���>ɮK"�7,Ȇj���{�<�QB�.K4�����+Ec��c�)D��`���/k z�k�L�����+D�����&DX��Sj��-����gB'D�x�!<R7&#wr����S�"��0<��G�3P!�X��I*B�l!��&U�<�M� k���Vj��_�Z|��GDW�<� �\�E�	%>��=��" �|gdtj�"O&���Q){JJ�`B12�J�Q�"OZ$�-Jk-��j'�Q�t�[�"Oh4���2��قeI�d|���"O.8sB.	�i ���*jd���"O(�����W ���R	�g�����"O>�9��Bx�JR(P=Hxe"O�����&,%J���d^+w�h�"O�X��d
C;�Rqe��M��<��"Od$����`����t�ֿ.�.)�F"O��8���^�����-[��P�C]�<a�X҈���GS5z��e��Y�<a0��w���`S%�:�0��Q�<�g���S{�0�ÕG��$K�<ɤD����S��R�{�R���L�H�<QU��e�ֵ��/��pPz�N��0=�0)�)%��p��Q�we���MLG�<)W�^O���ȲD�U~�tY@b'D��k�L�6"��(AŪ��(���rs�%D���J֪��qB��vA�[t&8D�P���JJj�4#FDQ\ܼ",D��k0	1^ݻ�.�IlAB.)D���^5:�n�H'F��O���I��+D����nZ�-4��wo؋GY��y�(D��sC�I�A�аdJL�Ɯ�Y��(D��:�cR�4�!��3mO�͈Ѡ9D��0�,W�fS`�$ʑb[J�f6D������<�Q(lF=���Y��>D�|��B�H�Ɯqd'ҀU8Xy"@�=D��#Ӈ�%���{����TG�aCf:D�p�eF�;L�R�D��F��(�W.D��[s#�U�Lu�ႇ�*1��X3*D�x�nؑ/c��/R��RE	$D���c���1!��!onM���#D����m8d@�P�!��u�H	(Q	!D����%}�0YÊu;-e�3D��e�N�F�IQ�b�93��$3t 2D��
D�*u��D��	�Dr�'.D��1"�=2�bԆV`�ܙʰ�9D� ��αHеB��� Y�I�U7D��2�!�~tzv� �)��o?D�X �W��!I�qzn,�TH8D�<ц"'%�� �ʼ)�yX�8D��K�DÅft2p���4%���2�4D�9q/�%Q{B��S-�O�@��N.D���0��"F��qD�%5�(ST�-D�4b%R�y���P�d�a��-pQ�+D�"�c� f�B���0���A+D�|�gJ&0+��ӱ@YF�a�"
,D���G��U��A��Ul�f&�O��Q�^0H�;3Բ���;�b���rhz�ܼs��Ё𭊕0 ���~�pI���H+{a��j�AW,v��q���64Ц<�'�S-�nD��<]B
�dE�E@>g��	�a�EC�<	��K�J�
DY� ��e@J��e�|�<y m���@8+�50j�P��v�<�JDN�h(�#��¹0���q�<a��6`*d� ���CZ0h0��o�<1Aoɩk/>	�sAʹ5���r��h�<) Y�/��(�� M�\�rC!�@�<�pA�f6X<K��A�G�DaPd^r�<��EaNX��E:}\�`D�IV�<�6O�u1�	�� �3vA� 
�$�O�<� Hl�����9$2f��#��i6�|R�'�azB,D$y�*����@�dd�F%���y�l�)h�aD� _t���MA	�y��6s1@��1�\�������y�o��{~=���x�9�3H�yReқ1Oĭ�X){��A�ă��y�Y�d�Z���e�)$h�XD�;�y��;K�t�Qń?u��F"������OJ��8LŌ���̻�. �b Ų��q�p"O�e��ʊ6V���C! ��`��"O����.tl �����VSt���"OH�8֭��)�T)r@H7T0]�!"OJ��U���8̱���+FA�s"O,�r�2��4�S'�*' ��'V�ɃA�w�
~���87��<��ʓ�?�+O��� ����8�j�?Ne�hQf���
o!�^���e"D�F�-h��xw/�J�!��W2_��qa�"�;'���{�矢�!�,ߖ���3��911̟/!򤌄~��<+��aʆ���Oy!��ւ�\p�f�N�A�T��kل>�!��$Q�)�%�?�\p 7a� 4��O���3O�Z'f��xt
��`eAW�!��A4:�
������I�2��/(!�Ě�/m.y@LݿP��T@k��!���+�$p�Ѽ�![�c
$_Jv�`�'�İ��Ԓ%��H��,*�h��'��h�%���@%��r@*� �'�����c�ip�cZ.n�����'
6���J:�i��&n��$�c"O8��mJ�*d�eHƗr����"O����C�./q���@��lp��"Ox�`�o��[y0�p�R�X���"Oj�
E�3p�d2 �8�j Є"O��i�-��{��(�^�H�4̉�"O`��"�� d@�ҧ���N�hcR�,D{���g�.`!��!�A��i�}!���8}���H'�õB�nBhՓI!�d�U��|	7NM�9x�`0�A >�!�DG�Jڄ���A^�DNwo!�d��EN�s��{ą�ѯF�"`!�ă��Љ�paU�"XBY�n˹q!�D�m�d(�G _���aْΉ�7G!�Ou�2�)���5�~��r��1!�99�"�P�p��j�|��3"O�uآ�ů�0X��	'���x�!򤚳}Z�� ҥ�.�4YY �U!���S,�(SE��T/x��3��:�!�d�&:&��
��́'(J���*�1�!�$�mM$x�o�p�,�P��
G�!�Z�zR���U�Z=8���%G��!��/N�EB-�Ɋ�C��;�!�d��%��ͻ���C��h80��!�Қ%��,
���,z�`=Y�C׋2!�"
�B��W�P�N�ٰ!$!�$٥&�`� ���M����&#��!�ĝ�TqpF�Ϙ�1���G�!���ޘ16��W|�)[ ���!�D����9yVbD�G��"u�֭v!�dG=;�<���ܞ��8��C!�D@{0|$��i�	h�BH�&!�L�rVt
�F[�6�"��d!U�!�$I6��[�`� �laAͨ]!�іx=n�È�,����4�D!!W!�� aWg�@��mRV�C���T��"O� ���.2D9���9*�V ;�"O���<�N�@���_�0�"O�hǢF�!�� ��,,����"O�P�e
ǹD^J:�I�2���;1"O@Y��A�%n2�EP4ኚN ���c"OD@sd�6��ʀ ԧ5 �+2"O�IX!.X4Տ	[(U�7"O�ib�mK)���"t-_��@f"Ol9%��6���W/lva�"O(�SB�YA���ң��7��5+V"O�)��"���z������p��A�"O���Ʈ�t�>|a�S�f$���"O�˥��I.��t��o�@9�"O0�9�
ܺ}���Q#�T2Bc"OZ˄�W�Fh�*���&@y�"O�d`@�ʆ,d|]��#��#��҃"O$#��ߥ[�F �E���~m�3"O8U�gd�1���pĢA�7��0*W"O\ܹB�L�%��K�O��!*�"OTy�D�ƺ\X�X"ŪK	a�Ҕx`"OZP���xd"���.�5��"OP���l��.���o�v��@�D5�S��R�a��"bk�!q���'?�!�DE�*֎=����<E�Q�ɑt!�D�2�hK�=p۔9�w��NN!��,�Jeh5�v`�����B!������g(G�'cdi#�zA!�
�v�8�ۃ��D
 �7�~B��$0WL�� 	�CJXm�w�4�\�=�	�'b�N ����yj5BD[bO�a�ȓW@T�zu��L����2�μ]$�ȓ/�MT,�/g©��J�|T������%�34�*���b��~�B��ȓP��o�+��ԋ�"�b�U��J�! �C��o���p�\�g��ȓR���A[�1�=���5����'���i�J 7v-cpn��Z��������"h�/T6�b>|`��ȓV�K��&�JIK C�<G� Ɇ�\���fI�5��a�.���f���L�'>Tt���>I-��ȓf��F���5�d�H0�F	��akZ�RC.C�3��)Y�ʃ�5rA�ȓ�&� �!پz.���2EY`��!�ȓg��T2_�[K����A��:�Ņȓ|�������B���`͵JT���ȓ,4�|��g��G^�-Q:pթ¦>D��`���J��2u^?o1:���94�LГ$��iV�T���7	,X�a[n�<iŋ;S�MhP�'�
�NVe�<pK�%� �S��f�X��7N�c�<��/X�U�̼��%7p�
�w�<1s�Jf&8� �F�47��
5�Zn�<�s�"@� 3aO�*�����S�<YkZ��Bt�Seϑi*8�e�R�<���� %W,��Eѐ:���B�j�ן���P��1I/	s��0�UF��D�l\��v�cp�U�L;�S &X��4���E��9��. W�r!�V!mpD��ef:@�f��'��Y�h��D��ȓGE���eAֽ	�V�	�iضQ����d�T��+_�t��ay!��{0,������5��{2���<����S�? p(��,=Td��вc�%��m
�'��D�~�0�ڇd;)ڝ�G���!��;Bz������p��D�%FB1UG!���j>u��1 ��)��Hs!�$��c�~yBSE_�C�� ja��!�/7��챂�P��B��{�@��'����=9�	��
M'��*Op�=E�D@���$I��[�� cT�P���>��OҀ��c�^��D�I�,G��I��"O44*���
sf��r��5'�PtC%"O֜���	�q��KP����4W"O��0���8p5��.}4��3"O������H�F/c��I�"O�Ux �ېL�
�dڌM�ȉ��"O�l*�c_�\��T.J�kpN�!�d��T���#7�G\�� )�#��7=!�I.K������ C��������!�D�!#(��:� MWx*-�p�La�!��2�"!��E ywLh���g�!�DA(�$�@ϒ`&)�a�_6<���ayb�|�ቮ4��X�F��6p,عa�ڷ
�6C�	�d��L�@�w���C�:Q�C�I�S:9�Wƌ�>��K�/	,kji�ȓ�r�Br�Χ*W��s�'*��q�ȓ �v�Yv�;�j��@�d?\(��6�p��Q(� ]<��S	� Q�ȓ8����υ4.r�y1�]
1�'�a~��K5@���
� �����T
�y"MT05�ԽT�^rTrx���L�hO��=a�'������R>�N|�#IV7_����
�'��]#�6LQ��!�fQ��d��'\F�8e�JΊ����0F����
�'L��Ar�O3d�>	��ŎEv����'���"I�<CvD�#4�߽4��!;�'Έ8*�!I&.��3nVV��)O�L�IZ�O��]���#F�2X�N."�Q��'��Ru.��B�z���&��-�x�B"O�DR	Ơ(ab(a��O	-�XQ� "Od�	�jL�� !��D�zv���"O���$����X��t��/[�`��"O������"T���w�	V�y�r"O|PkT�����q`G;-uX0��'j1O�h`�j�,F�QR���T_���s"Ox��f��.F2��/T*VR���"OB��7$[�8�\��"@��{`�L{�"O��� B;�vl�@�~b�Bp"O>%)���<	W�p�Ai?d|�к�"O��(�[4�R	��獘*hl;C"OBi��#܌���g��-w`Mq��'r6O�cV��u�z�Rr��9b��""OС�1��� ɰ6�0Y�pس"O�mڳ���u�$a(�$"����"O�X`�ԫ��xx�W�p��
�"O�00BC�w6XL �-G�x���"O�h��k�1�Lx��,�9!�x٧"Or�A�y���ac�1���v�'xBJY0Z�j-���V�԰���ў`������J"kZ�X�<AP�-A�.���'��V��,v���5�����f�#D����*� h����>�ce#D�P�t&��$m�@
�b����ї�5D����]�b�[��Ȕ(�ܐ�Cm�4�?�����ӷ�߃N�~	@U焎Z�欨�j!ړ�hO��I1(RX���S�c�4��q�̫Q)B�)� "l�䦏0C���q@_�r{���r"O�a2��X
6�T���s�c�"O<8���u��i��-
B��"O̐�0'�7�����. �Z�"O53��X�B �`�c��.��L���'�ў"~�օ�D��R��P�p2�"�*��O�#~�Fċ9b.0X�(�8��d#�F�v�<Y�FϔF@^Y�D�[��t]���-D�xs��D"�a�rĻ�Z��59D���$�Ǝ��a����	����Wi*D���
=O�`C' �%��B"�)D�,2��E$v��C��7���&D�|h�P=#���0�o�* O�����9D��ْ��z2�a��-Ð �$�F�6D�X�c��.NH���˝*����5D�p(����T����˝��@e'D�h�4僷1��%�v鎩 Qd%D�d	6�� �-� b�2�Ћ��(�O��I�S��tC��Ȃ0�8)fBݧ�lB�	-x����P��y^����Yx.B�	�U�NqВ,�81��a�]�9A�O���D@!*~�M[�
W�L�>�Ç
�a�!��(rd ��3�*Ea�N&j�!�G�V�D*wjۖ,̹�4Ό0�!��D&"-.y�D�K�]"�D�T���}� !q��;b��;�n ��l�JeN)D�<+��T�1t�X�S�ȣ{�TM���;D��t��.z�&M9��fr��!Gc�O���:�D%OD � �+R�H)�P+6ڜt[�"OZ�#*>I�F���ۆQ��4�4"O���� �wE�m�å3p��A!�"OF2��
2ē�S�"!������'���p0`$���+?�\���f�!�¯*楁WR�X0��ْ���8١����m���V���1s��{C�G6��˓��$/LO��qBAޒU{��Z|�IW��w�<qՃ͌O-JL���S� F� T�Jp�<���i�"�ڴ@���e3��r�<9�]	HK���F �cOʰ��H�q��(�:��� S*7J\�
�ps���'�a~r��u a+dg�"��Dȳ�]��yB��*Oհ�a7�B/ T9�s���yrkP:��Idf�^J����I��y��.p;��y@	���@�aǮ�yr��2�4k��mo"p���;�yҢ��M��� ���;9��k�m�4�y�V�$�V�R��!3չq�ܷ�y�iD>\����	~�\�9"�����'hў�O V\i�/ϞD�>2�����>�*�'钍kf��r��4�Z�p�'
�}	WG��F�X�s�l�D��y�'����p��.:����C�;;7��`
�'6�������H���R�� 1�,�z�'l��FE)>j�z�E�+%_ X*�'.@q�o�+f�|x!QfղI�p�z
��y���_Y�'-t��(4�T���7�O �E�+Vǰ�R��T}��*�"O�|j��]ʽ�[�T|�"OL�rm[�a�^�Ґ������"O��-Y� 51�G��6g�}��"O(���ȁ!X}�̨ ��v-��b�"O���+�GtD0y��4�.��tO��� /	Vݼ��P�
�J*6�Cӆ"�O6牯~&��4��mBh��p��2��C�)� t��a���bG�e���g�lt�"O& q�ȝ��R���`K�q1vY��"O�R��W
4��i�NXq"OX�F��E�t����9��J"O� �q��1|��9Kf�ϝn|=I"O�)z�[�G=\ qMܨ�"g�|��'�x� ��g8y	E��7f����
�'�yCFmo�����K�d�� 
�'�0�【�H�hͫင�jh@#�'$���,?3� ����E0���'�*(�4�5P��4� �
�'ن���(YZ,��Wi�1CL4��'�D��UNӪy	h�9'� �����?I��Py$b�����Ɔ�s	�'u�y�EM�X�p���3flr�'�z��K�p:�@�F
��L��'8
Q��-�I���"� ��%8��'ڐ�0 C�d�(q)�dY2B��	�'��v'�'"`p�.�Be�	�'ўё#��	A��`��)'�`%B	�'7@�4��0Z/�!��艣#"2İ�'�\=(��;O"ru��r�Ρ�'�H�gH5H~ܷ$�y
"��
�'6��s"��{�ƈr�MP�\��	�'��5���x`1�fA�^J:�y"J&D���C�6g���(_�A7z *�� D�<�',v+��ެ_}B��`=D��hH�.˦�2�D��a+h�b3�%D�89�ڽ:�� �2b�Ix�(�>D��Qb��)2S|�(��B+�
��0D�4��-I���Ke��g4؅
�C/D����h	�S���p� ��F�)3�!-D��'��	�i  "��*�X��,D� [0�Y�Z<�T��(����F-D�$Z��ϩ)��H3G��*0�<�+4�>D���%kZ/y(*�J�T�Bí D��P�g�8C�蹠���h]��I�=D�L�5���,IҴ�Dd�2F ��<D� 0�)0��l◁�&f݄�u�;D�z����f�j�3�K^+R�P���4D�0" ��"���()�p<��Y�!��S�̞HkQG�!e>���j9e*!�LbH<P7��,�4��e	ګ!�D+_%���X�z�z�rb��~!�d�'����.��^��AעW{�!�ѥx�(�_��{�k�!�$�(1���Y�,X�w��A��ږc�!�d�2h���%BBh�jx��VD�!�d�i��D#��W�.����U�Aw!���	��b��ߙh�$���?!�䛝}�����H���}��c��p�!�Q�N���h��Ԉ]bD8�M+�!�d�( v��po@)SR24�E+�z!�D��Kb]iRn�1�R��JN��!��QZg$���3U�:�9���'y�!�D��J�b�·�@ڄe��-R�"?!򤑃Ȏq��V�~�*�;d� !�$�+6X$��ȟ�o�Ƚ�Ӭ �]2!�?�e"'i�+� �8�JX:.�!����&����s�rX����<�!�䝢nv� ���R%.�k���0!�D�<PfB]��hJ�]!
���<a}!�
S�b`���e�����JO�!�V#j��P��O7���vM�z!�� �=f �f4ː.��?�m "O*X9��G�m�pa9���u��}'"O��J�#�d:Q�W �w�ԥ��"O��*�錱U����Lؿ^�$�zE"O��0E��y��u�fJZ��a0�"O$n�� )��1��ʈ6]��5"O�UB�.�@�⽲SO�*_Edd�V"OҶ�2Z�g>H�vy:"O����ςf�b�gH�L�D���"O�,�F�	�r�6T��=JrȘy�"O$��jM��4���E�/{�>Xb"O���c��;�`䄘1�H �1"O�u�S���ļ�A
¶i�.�ڃ"ON��REW�y��iF+<�N<i�"O�A��V�== �,Lr�a�NML!���t��8#g�1o�I�sm
A!�d@	Bx!(4�F{�`E��ֿO=!��;R"�-Rv�1gYq"e�f!�$6F$FXH���T��4� 'D�Z�!�dϰ\h�HԢ�};,0heE�<q�!��,�\��V"Օ76�e���L�!�$�.2h`5n �Y�dI�,[,Ac!�r���;��&k�04i�FD!�$,{T��&I�Ljf@�-�q!��G�6���@��Yg�0T!�d_�F�s�% l՞�h���&�!��{�H]�1n��b�����'X�!��s��ңi2r���pa�$s!�$�H�M�h�I����@��!�d��jt֐�q��9URa����&S�!�D %t��H1ĬP�_��#��]�D�!�Wv�����Lv�� �6�!�$P� }��㦍�j:�PH���!���U�P���-����aG�t�!�S�p���r�Js���ɗ"�63�!���5t�E3 ;Y�x��\�\�!�d�y�2Qy �JLT����$f�!��ƭ?��b!�߽b��'�L4R!�$�UZ����O>0�����Q�!�Č0m���"�+Z�t�ވ��g�*!�D،"��= �Ä�.~��:è>u)!�dUG�vxX�AI	_����F�^!�^
`Eh�q��YEJlH#+�	=!���_ j$b2�Q�v�a�f
�j!�@�p�j���/��tl�B�k]!��[/ �>X�d*��K
Q��ϊ+3!�d�	x�8Hp�'Q�zY�%��]!�d�
q_����)�8唰DoS��!�d
�$H���L�R�� �˸�!�dǷ%�&a�dm��<���4^\!�ͭj3�]��E87�|��v�^�!��!\i�!D(ҖN�6d�6�M@�!��0@�����7�b9(�H�!�d_%B���1�I���]膠Q�L�!�D��t���+d�Vj^4���iь>:!�C���� �>��U2�I��0'!��E}Z8�2%A�v����Q!�d�v((��ȟ����ԬB��!�/N4�2�l��$t�!4�M�
�!�%U������ {n.����݁R�!�d�u�v	0G�(,a�80�$pG!�DSwFqh��W�#�Pi���))/!��(���y��	D�꙱P��>!���
��H���N�b���G%I�!�� �}I�n�Fv�D�E(�F@�0D"O���D�Jj UKG��#VJ�b�"O$� 利8����1�K�DZ��q"O>ź�(X�Sv|Ix&E�&BEJ�	�"O�p���c�}�D���2%��"O�X�bG�ea�����C�8�"O~�s�⅓� JA�4�$���"Oƨ ��̩W�V K'fH2�����"O�9���w��AJ�E�+���Q"O4`�rb�z�x�У���-q�"O�1R�Ç�OA������:|�> �"O�d�sۜ;����g��nΨ��1"O^\�P�e�j�[��)|�5R0"O��"P��P`�\YG�H5�Ƚ�"O�U��B���\�"E8)�nxP�"O���3�A>X|Xe���!� ��"OP�B%���5X���d�#"O��J��M�}���K�2i���B*O2���L�-�J��ҔP���q�'�>�pW*�ik��9֏U
t�0���'�.u���5��= ���s{`�b�'�6YӉW6J�´�f���j�'��Es����D�:��(P��l��':vHa`D��h�y��Dq"��'������?uu���N��N�Y
�'�$Z�C�o��UL �𾅹�'\����ɍYWΘ�� ��s��j�'τ\��`�V,�P)��P��;�'�FpA�!�= Dqv���ȹ��'H�q�a�Vq�b�xV�ޙT"�C�'�HL�����M�MCq'�?s��Qh�'��3�a�1���T����'	
�ӲH�A�ʀ��.�HSv�J�'�F�xP�̯��ms0NQ�G���Q�'n)���ΒRk��;Ю�*���'e4�it������o�4����'���
CX�A����h��.�ޡ3�'�6l��*4Z^�	D���#1�e��'��L��� bb,I�s��f�1��u0� �F�r�"0`.�v�~���n���y9�4;NL�	���ȓW4*= �j]
i�����=�t�ȓfĐBb,_;����-ڣG`���ȓS�)GFP�y��0B��υts�܇�G��W ���]{w��>�n|�ȓ1�DK7f��.N���$�6�B���L[�U��ǥC-��#�Jω_D*	�ȓ� � �/�*0�,Js`��@�-��?t�8匝�D��}1��X~�bh�ȓoOx�*��P�J�p�K`*ON����>�X^��C�A��	tpС�/�F8���z���l�4_��:���QQ��qP"O�`�P�Dd�����67V��"�'p�(�'���2u"Ch 5�
D�F��'v��d
0oV<�CŅ?Z\�c���*�S��&�,YP�g׬!���JÆ���y��B!Q���%�R�j�@�,�`���<	���O�|[6�ϩx�fj1'�1m�����"O��I7�X2O�̭#c�B���̣V��C�IfQr��T)N�F���O֦���	��0�th��� ,�h�Bb�Uxu����\YR��e2 �J'�ʺ�0�$���'��$!��8���/p^\Xw�ܔP���ˈ�y����I!�OO���2�.�?��}r� �g?� �DG^nW�%C�/GGԜ"WO��DE?n��"ǌ�K��0k�"Y�t!��cB�hڤ�k��@��@_&��x��ɰ@��[#���l��]�d��6�ΓO~��d�*'��s�GX� iarM��!�D��n�B�A����l ��a�Tb��Y�Y.�h5�L.A缁� ��(��'�a{��V7���*�d�7?�*� 5F��yLR4MQ�웡	8
��d��MS'�It�'��	�Aҵ?�V|)#��I�,�1ݴ�hO駆�'IJ1���H���2�ˎ���'?�M( EJ/'8��(��6�lek��HO�5ˇ퐣L\�0Q"̟���Kb"O���%��F�|a%ԱG"��Ǖ>������)�
a�1*�w<��@$�	0!�D�".��M�j�j ȕKD�e!�DNG�a��W�i ����÷`!��Y�F`�F)S�Kg�=��Hϴ> �ð>��m�Y��芕m�u_xA[qo�B}b�'Eƴ����ns����b�U�
�'�|y�`�7}<�z�-�4<,��	�'�"��,wD�!�ܮP���	�'��!��[�Vp y�N�)��MJ>�����U/$F�H;O;�U�ź!�$(6����ʅ^*pjW�ȁYqOT��$^�2��"��U#ƙ�q��G�!���&�8�Ңʼb�/sL!�N�Q�����mE� ����T'��Ď����0|����N��E�:}�y�#�(T��Q&2`xc�R�&��W��Ob�\��'��TA@D;V�ʐ"�$QBp��Vg!�O�˓$$�����:�0�&��I���'����)s\����B�Q�V����E l�C�IQ.n�h+R:Q���X�$`c B�	�t�9q�)�|��p��ȂB�	���@��<^�����nB��(Ќ�WmV�X�(�#�dS�sLjB�	�2��Q�@� ���� �B�	�XN~4�a�9B0�����FݤC�I�R�  �k7-�჉�%�.�	S����@P�֭^�	،|pw�Ӻ7f>���'���5]j��0�\�Z�.��D�>1F��>���\����z��&
�a9$�w��~2V�2"m��n�py��i_�KB�2�@4D�� ��d���Cr�?�(`�5�=D�\�w'K&�y ��̡`@lX�G�:�IA����2e�k��9Pg��h,iW:����ħAAN���fD�\p|a�c��+�\��<�$(��SR$A"�"-��$���'�ɧ�Y��sE"��Tcʰ� �: �$qf>D�����M�SZ��#h� H�)�p�;ғ�p<�^z�<����;�	cb�=	}ʢ>���	G?w]h����	jg6������'J�+�,ھx��(Ce�E�u�� �O�iGz2�/�Ɣq�#d>�,bc�Dd,�C�	4�v��� ~��8iA��u��'����߁B1�İV�V�d�ΰr��$D��}r@T��~�ǚs�����S}\�9��ۢ��'azb'C�-h4 �:~�b�Hջ��x�&Y�b��4�U�,��l�U��VU!�䌲7O��Q2��#Q:��PST'c�!�L6[���T�M|4��ץe���� "��\˧n8(�@2hˣp:*B�	?i,�t���,A#��'b�:`��C�)� �@J ��B�hͦ;/��35"O��aǏ��RH`��'g�a�ve�Q"OlH���'~�����ՂJ�J���"O8����"���z���4l���QE"O���i�A�8�ζM��4:�"O��YjV� �������R�:<��'�ў"~
�7T�y9uE��W���A��L:�y���ђ�F�Ȇ���=kB�4_:�"�h��fHK��S'}�<C�ɡ*(0����	|���84:C�	�"�!Gn�(X(8��O ��
C�	P����&�G����1jY�C�I4\�0as�!�2׬� 
ݶ}�C�	7W��D����h+��{�B,C�B�	�m��<!U��%��a$C?+b\C�	�_E��C7�ǽ@���gZ��	t����Z��'n�����,�/|�T�"O��� �<l��3FӠ^[4�r!�	T�O�H�D��E�8YB�M�$r:0�Z
�'� ��pl��)g�\$]#mJ�"�'����ӌN*B1��cG�KZ��Մ�B�	3c�`�b��5����"˙�i��B�	3<qP1��`�ԋ�+[o�O��=�~g�U�S��P8���v�LR�<6����L�"V�-�v5��'����xR
A)��"Y� � ���0?!.ONyS���53z�z�E���A���Iox��a�B[��z�A���0r�i:��M?��{�~RU�աaL(Q���@#a�T����C���'���>���U�<��	I��A\��$�#L�pH<�'2 �~�jV�C�D�Rx��)�%q�&7V��?q�Ȫ�����h���y����n���g��O0�nZc~�, l$�1h�cB�s%�`���p?9�O"�rV�N���r�����*��xr�����	�R�"���(P\�����-��B�I�4wƝ˱��78�[���lZf�4ϓUz:}����B�UQJH�~.��n�oQ�"~*�mJw)�\{f��p���цW�,�jB�	5y| �`W�D��I��h�
`i��DXh��$�S��$o*���2���gt�a��ɁZ��	8#�`���S;i><d� ���\�6O��0|��S�e�!���Iτe
V�g�'fў�'�=K�-�u�.e��)w]q*��>�S��yb-9���Bt�%!8*}"�bE�X�6�a����|�J�t��sI;̥�& I�yr��02�Ta:�#;��6��y⇁"e�Z�R3	E�+�)�*�5�y�j	5��S,�1��)����O��� ie����eA���
�bHO*!�
�T��9r4)�]�l��B�>!��E,P�)� Q�=� ���LBG"!�A=V�ȍx6�N�Gv��ibeML�!��Y�<\�Z@Θ
Zb��g�L)n�!�$$j/މ���[#(�B)* �Y!��Ijrt0d�Гl�0vhO7X�!��׎U�x��O0gydAfb�!��<e���#.C�TH�S%	k�!�䊬��4�����|��hH���[�!�S�V����qk�N�����$+N!��ܩ�<#F�-��|�R��,L!�
\Ȑ���T�.�̽g��+h!�T��C��#�:�
�F��FZ!���L��\� �M=Vo�y���*�!�$��4��$�A:�+��ȃ�!�� ����n� u�M��˺d).	"�"O<� #ho�r(�c��G�l(�a"O�Lj7OF"�\�BWRۆ��"On�X���
�������O��!�"OL�el�!n�Aj�".����"O�yzlHN�6��*�E��zr"O�l��H�F��R���n 
Da"O�4p�b�	�h� A�C񲑨U"OP�C&\�3���#���B���"O���DߪB5:H
U��=���"O��ϒ/QJ>�3�n�>(�(� "O�-�v�BI�،�w�Q(S�>�v"OB �����Bx>��1�
D�r؋$"O�P3�*�tx	pbق�*�qF"O.��܈>*�Bt��cYj�2g"Oh�7΅%�Le;�BC�c_0�0E"O|��ve�V�rY�(ɲ<��a�0"OdS�h�*.�z҆Բ%ɠ=�`�d1"ƾ�B��2��E�Q, b1O�u�fL+D��U{��P�����q"O����֊�PӤ�O�$��"O�ti�N�L�bؓ�Z�J�t���"O�����ޑSV�Mx�,0^�����"O��b�I n��%�
G2W�|icU"O���I
���3�C.o�R��"O�I�����HE�W	�A�(dq�"O��J��n���k"(��"�>H� "O� ���̴A ���/��Q�"OT<{��A�$Y�ʐ�qur)��"O$����t���a�i�r�va�"OX�˂fS*BC�!9��D�x��*�"O,�rt�#k�$(�0�ߤs�8ͣ�"O��*�g�,q�h�STi�E��a�"O�-k�l.(>v�k����w�H�!�"O^�C�/Ŕ5K�l���,���j�"O`A���nk �)�*N?0Mxe21"O���6�H�#���`�*�7"N�z�"O2  �nWA�ε�Q��-O�e�u"O�y����/MF@�j]$��S"O���t��+t��hP�1e�f 
"O�څl�>�`)J*>c ��' �ѓ��2f�y����x�n�y�'�(!邲_��azS��JUT��'�A�,L	.�Fir��Z��`u��'].�㥦Y�zC�Xkg��
J����'��`['+�V�@�Nɇy����'�%:��˅H�ޝ��
 �q�
�'�����BF:��!,�3�:��
�'�mCoI�""�̣p�G�;��[
�'��I`$���	0���J=k
�'P�M�⬃P�	g�]���4�
�'��d�w�ŁĪl��‑c"Z�8	�'���z��ʤw$pm���۸d�Rm��'֦��ăړ+�V ��(̮�b�'�vbEBY%�T���K�/�|�'�P���9���L�.m��X!�'��E�ƿ$J�)K-�����4R�@����V�ޤp�dN" �\Q��W=O�Ɇ�	�P��u���Cү�f�Up�`� ��(D�芴��ss�ف�U�6����%B�����OI�Qh�
��Pψ(`��gfQ��'�J���+	`��#m�UKr|ZE�ը��'=0�F�,O8�2�o�#eR����!N���"O^݋�Ŝy���r�W+Sl [�=kP����'��h)�랚X���E͆6~�EH�u �|i��-?� d� U�S! M*����^:W�A�"OTQ	!hȋ#�Vu�"��46^HQX���MP����\�s�[�+�Fq�����n�V�A�"O�XZ �O`���S3(h�0"O2s�?k�Fa�#B]r9)�T"O��s$!@@���Y�x�ܙ�"O%
�(�B�&��ddĽVT����"O�	#҉�
v.d��Õ	<16���U	>22��ǆe@7�ΈT<��d��	S�� v�����Q�����w�0u��b�@劦�̹�p=�WC�S��˓Lh�p�B��W�(A� ̗�d Т?y��˫:tZc?MhS�U+T�)�ӊ]�|��b-1�I1Z�����?��h"bܵy֘�!�ҟK�r��e;�(�)ʧiq��+��J�lK��Zw�"<��ɡ��>Q�qO�}��Y�x�"�O��^����.�@�%��*E��&-�D���p���I����"'��3hB�$��뉚04<��
T�mm(}�`�~�B8ٵ!��^�F��D>B&��ʨO��pa�/"�Y���3�f��p�'��< ���{�Q���O��3(Y����c��qFxRL׾O��?AQq+ۨ` �Qk�j#��i�1?��D(C��"|��8[�(��i� ���K_�<�(PC�����Y8F��劲�	Q�G������)Opm)���f��,H�lڬ"�\�7H7�	+{� #|��,��H�@c��=L�h�R8L<��R�T�Pxk��v�h����@i�
/��S�V؟H����|��Yaȝ#dv|�'a1<O�	ш\�����2A-��s��|ӗ���U�I.�όw�i�U��\|�"0�����J`x�(cf>�D�$�8[��ټ�qO�5�C�_
K�X���&)��I��l�d�"'ڕT��$J�α��*s3�zҪ�8)z�D�����@8fe�� 4����Z��AU��]�C�'���K�g��Yܔ-�v�X��_)L�q�hR�4[@����d�֧�L���ڂɔ�1��A�銕or�|�t�	)-�HՐPC�&��P�'���'%��x����5w�AI $���8�1B8�0=�Iʆ�����`��T��DFm�����M������BLf<)�f��?�8� �@��<9��X$P���GDҭJN�� ���@��Ԃ�dY�G�����$wW:a!�œ\8$k��ˑ.���S7�A[2E  eB�C����	�	\p-�0$ѡ_ä�A�˶@�j�t�fHVf��rt!��A��UK��Օh�h�PF!�.N?���A�#t��5�@f�ܶ���/޼ъB!Ѫ_H"0���Ђ͚�-��u�� E.�!퟈+Ԩ��"�Qj�ʼ�E�*Z?��->�<A����DPB�I�%�*A�3��[��(#��2K�4T� c�Ѽ$�U���韦s�U�0��'����Ć���gL
wfn��"�)�OR�#�sL��[2��sш�jf�0j|�!)\���p�퉩 m@�H#�>����S��pِ���6R��I�%}Q�DJ��Ӕ	�rհ��4Y��b��٦ u4Q��� ����I�=Ay����'��5[:B�ɏ%������M1�I����R���jث�o�.'�44���7QR~�(���lϚ4�BIu�F��`QQ���0�yB��,!�[�ꊖ�&���K5��z" ��q��x!0	�LΠ|k��$�|"/
�-St��g$H�H��H5�x2O
!/�"���2m�����J 3���0.��V���(��'�h?`dD���&X\Q�`�|���8 7�O��	5��u	zDa�Ā)�L��b�ZO�@�AG3�R8��S�����(P禡�T!�G�t��"�.PҢݐGC��	��\��Q�Q��F�����ӏvD"|����<���ٖ��)v^La��gp�'��	�6|�O�܁�ǯݐw� Ą�2;6y`&��}��QNL�@Lz �#���� {V4��Ŗ�S�f��Tn�J�-�MYz%c�&�)�'�XM	�+밌h@�V}�Aե�l�jY�J  1k�N���6n^�V���j�E1l��d�'.?��J<g�d�O4���d
�e�n)ᴥ��B����R۳m\��8|F���!@������0ڞ�I!���:|
P�����q_����3��ܶp\��msA���H�H|�GW� Uyj��ɕ %$�Ӡ�I'?ur]G��۵� ��JQ�gxhL5�A�J}�Qc�N�"��{�Q>�@4MA�f^�u�D=�g����U�ȓ3 d���C�yz�h���$Q����^�<В�֧� @A�G���&�Ω�DN�-\p�T"O��I2�~�1�ݙ��(��=D��C��3: ��@F*E�(q��!D�|`w.ϸ[�L���%u��)�qj+D�����M�*g���D+R���I3�<D�X��Ǎ��2�:w�ݕ{@�i�AL:D�X1B�_�Z��Ԁ��݈z���C�:D�xv�WBE*�6�9��w�:D�`���:�P���n�%AҔ�IE�8D�ؓ�šU�<�dG��1��h�6D�p�A��$C-��R�ґ�D����4D��b憘#_5�kîҸ�|�A�$D��j$FX�*�p��A,�HRPX#`�6D���������v��(:`�5D�� `e^5_(Bd��@�����A!5��x��/ Q>=�Â�ta+�#h�>�(h
L�<yD�9/�0Y��m�|�����G6��˲�S|x��O?�d�G}����ϝ ������G�2[!��	��3�z�HN�kp`�']6��vk��Fu^�H��'Y��Q�F �lu����% �@�9��([1��lmX�B��ځ$AN����VXb�0�-��x"��V M���]�<=���B�����qjra�<����L38�~2�=� �i� �2#F�����y�<9��R&E��s�Ꞧ}όk5�	�&y�!��`��u��L�0T�(��|�לxR�H�H�X�¯UQ��CV�͜��?!vD�K������2.v��l�ktڄ.ޜ~2�8���O�~��� ',Of�
�'F�:P��օN,G�r�a������H1��8�Iꕆ����qU�/!�v1��(�^�d(�6�'U'��2�)7�O�|)s�G8SKfYU��PI��W�$�)U2B�RPj!ʟ:Zƀ�a.Z�L	{4�Dd��G;3��U�Uh\T�蘚@�u#!�ā F�H�3��8]��YҦ���t[ n�hs� )��9K�cA�+��T�H� 31�k�(��^�1le(e��?U�lq!j&�Ob<���� g&��^��\�R!Kl8�U1����?ap�ը�ʗ5Ĵ4hC�	������8�j`p��� y�.�?	��C��Th���m����
F;t�>=5l��QBlو�#]?_r�T8ЉV�� ������!V���A��(>�l�o9]�$�;��^`;FE0���O������8F���afc�����&�^�h����\�j��
��zR��8R��
�P��3��_�$����s�Q� �X}��L��<Y�*89�yCb�U'Oȴ�;M|�6�W*M��a�;I n�QՋF��5Y�`��E�<Q�$��c��]�$�6ҧ ���:U�� a݂@v�J�6�PQA�/P�P�`��
C�˗���*u�U `�Q��{�-[ v_��Zw��d\<��D\�RӢBו>i��z�+ݨ�)`��Ғp�FY�F�\2�E����@K@H���r�nX>�,Hj�#AG�t�t�Hgs�����¬|0�]���ǇI����'���.��g#$I(vt�\wn���>䚧�ڧI*x��2k�ޤ�֫Y��@%�FCW��6���O��m���~�σ�v�l �0��}6,�[�#��N�(XX'�F��y��cB8!5V��/Æ����uNr�rw9����e���h$n¹Yʬ��$�8Z��1ȲhO��� �	�a�4x�� �'��&J �¢�-H�hۇϋEr��zB��-+�źt O�{��ht�;n�S�+�#3]�\��u�lXi� �f���'�f���'r�|!��
��L��./%�8g�]�	v��N����gIχ������ �x���(�^Y��y� qp��{"+�X͆L��ō�Q* '��!�fI�,	]^��	5��ps��+�k\ˎD�'z"VyjD�H�eW���2��>�zL��I�)��]I���|?���[�-B@@��=�`P����	s l1�%Zb?	vÊz4Z�k�k
��	X�)��P�Na��B�E�J���rj���9ٕe0�� ��%��P,5[>����(�J@흳 ���z��6���2��!��-0[��`'(O[	9���ɉ-��@0�n<lhS�'r崈Ї�����r��I	;���FƷ7M�u�'H�U�@+B�aLXH��bm� �y����&<	���tX����,@�X憝r���s�0IqӘX6�0R�Ҭ�nP'hb�$�'�L�?�� oA=\P��E4j�M�g((D���ƌ[E�����@���M�A�����'�3�I�7	��〇@��pÐm��Bቛ��,ȗ���%�Z��� X����J�}�!��� g�tE�0�ζ�je�V�C:.�!�$@~�2��7z�܍�wN:*�!�U�S-vq�v��A/r0�wN�v?!�� �tB�h��6�2��πX|��"OP�[��	 ������Tpa{U"O}1�g�	� �Z%ét6bPB"OD����� &DҴ��=�
-�b"O�pG*C0,>(�s �Th� �"O�����X}*D��#R)ג�`�"O�Ԫt�7V�LR�!�07����"O:��q�A�P@ď�� Z�"�"O�݂��E6M��\h���z��Yڶ"O�`s�+E�`�[Fj�I�~H�%"O�b��D�����Ԉka:(��"O2@�'�ՅVt����i��wQ��� "Oܥ"��ͬs�����O��\ݑ�"O�i#��L�O��0!� C�H�Ƀ�"O̳���8EM,cEN\�x��"Or�AE��K8� g��-)
ΉqS"O�=+�¢j�"��O!i�I�0"OȩK�c��5+���W��cx$�q"O�ԓ��U	�q�7�T'#Ep���"O�� �*ᖤh"��#F�`�"O葱J�o��殜�6݀���"O�ԏ�B�$U@�g��]�d�Y�"O�X�@�W�AOX��V��Y�)�s"Od0rt�F2Kl�	b"���b"H��"O~�85�X�5~�`@��zf�)�q"O ���C�'�(��d ӰZ$iۤ"O.�:�!�.z�)Q&�)	MiIR"OT/�>f]ΡɠL�+��A"OY��hB�Wt�x�
S�V�N�Ȃ"O���Q�D4y��)ʒi�0�ԅ�"O6�8b��Y��#�X�0{�"O ��՟phtIҁ���z�0X�"O�I����R���இU0�5j�"O>�2�(���X�Ѐ-Q�?�4��*O�J� ��Y��ȋ��g�L��'KX����¢W�|yǇ�l,�7"OP�ӊ�/R$�豑�X� c�IY�"O�٩�#Һp�x��&RP�5��"OĤ)vh˥?�4�R5�@%kN^I��"O�Y1Cm�PϒDr�+O�'��t�"O�A9!K�B�fT1�)ҼF#��a�"O��S�ʐ3|�U��S�R��k3"O���H�I�)����3?E@�"O� ���@5&���@�fY�?ʅ��"O,��W�\�U��]����.~�<aWH\	|4�X��^�i۶�z$��x�<!��Ȧi���ѲB����h��n�<�T\)e��J�(J=9�U���M�<)��Ԇ2B�
�l�}���SdAg�<��U�)Si����=cqf��g��a�<Al@,��у��|��1
2�BY�<�Q�=tP�)T= ��p���^�<�g(V�|�9���C�3B1�	�U�<���D�TU��DF���QrtQ�<����'UN0�`f����~re�S�<ѕ��u��\�p�G�%�����`�<��m��(�ph �������k�`�<Y�f�:��@f��a���)f��v�<A��L�b��#k�ca�1�ՇMn�<i��ŭp- �Cً>�!�h�<YĥK7<�����G n �)Zg�<9b�ʁ~�IQgŤl���jd�<IF@�)$���H�-*�u
�cg�<��G�W�ƙ`�)� ��8*�)b�<� �(��C�\ 5���nu���"O
���U  X�}ض�ْ1p��A�"O��"���+&�:��8%xFa�p"O�l7k��C������SS�F�<ѧ�����r�'^�SD	�e�<�W�rM�fڀ#O��І�Gz�<G�
o�� �u�X�Y�	���z�<�u-֪�8�B�h+|~yʔC�<ٗJ%!Z,�0t�>z&"e�#�t�<!�@�<F�Ĉ:�n>C͞1q��s�<I�ȁ�AN����лo
�	Zl�<�f��0�J��d�Y�r��̙��Ns�<��&W�jB�#�M�`p|����q�<A�gɭq��i���ҽ�pܑ��l�<�e+$5�qxRI>TӤX�4W�<��FS�ui��kuN�q�(̨��][�<��X/0-8@�)��y���W�<A���}'��Y���1J�>� 4��M�<y��ġ.z���qȄ�P?�(cm�V�<Q¡3�����A&�҅R�YL�<��"��*�4H�bK�;:��e[N�<����M��\�@+PTۄU
�g]@�<i��^�{���Ơ��/����!��}�<9��ϿeE�гE.�
n���F�l�<���՘D��b�D׍>z�5�Q�G�<� cʛ}TT�g&��l2����)Rk�<Y��������	1��qK�g�<�3��][�s���XMx�	u�b�<Y2.6[�.��-@;�$����f�<a`���*��ׄ��x��ؐ���c�<Y��ߖl�<Q��bXd�L�wg	ߟh�F�'(�q%�֝)N���>I�b�RClISD	��M�L[3
�r�h�ŚSD���	"-2��	FvF��&��*d��0JH$�c����p=!F��Q����X!ml��N�a����1l��4��64�a��(�0Fm����*����{(b��.$D�����&�����eI`�
�
��1��0�Ȏ���d�hP�(�CI �䧎ygLٗM�}���Z:)�I�c��y¦�����  Y�*�>��NlX8���Y����<�; �������4��'�f��u�2
�<�Y�Ғ���kߓ$.�q�;e�b6��Ⓖ��Ƕ;�eyУ����U�$5����ϋ��0=�D�Lz���Q�JX3�R�qB�f�$@`��	�'�@�],R�X��R�A`��;�"�"v�b��"C�E�,D�4i2�J��8eF
�hb��DM�%kz��t!���7E���%C҆��'�yGM!�,��(F�J���yR��p�^����_�`eA��.%�U G�E-|���`*�<��p�T��� ߏ��'�	 `'T&fV�9#%�э:�Q
�q�f��pM��?)�N��9��A�a����N�v}2�Ȑo
��e�'A�@�C��Pm�c+�>�da��D�WC�HJ>�.�O���l#�j��߯\�l�r3�J'	>C�I	l��I�D�)
`n@���"�$B����}b�+G?>�j����X#f^B�		�εxů�01���d/Sk��B�S�����gFF�vԘr
ەAѢB�I�oJy*���5UX�����ܪB�	7TK2,�u.	3�@x��%�.w�B�I"6��1�	�ym� AW+��w�VB�	�L�����?^ʸ���' ��y"��	$���!Ċ��I8xa�k� �yr���:�h�3ņ�1_*@i ��8�y��N35h��Qȅ,�P]���?�y�N�O�R8 ��@	
���� �ʗ�y�@���(����۩v$��Ú��yR��<L���}Z6\A`DϘ�y"�V�z`h��]�m�LT0wK��y
� �l����d�X��S��6(G8I�6"Ob��V'P �cFH�P��X	u"O6(Ҵ�W�t��xj�nI�_��)��"O�50��W9���U�<�$@�"OL!"�f��t;�y���Qzʨ�"O��Y���l�,�2�J�'BV��0"O��aa�K�R�zrQhU4OH@�F"O��⭊|�4�Df�)v����"Ob�RaP�)	49��%X�Sf�䱗"O�����'%P�!0���lg�Yە"O����#�K��E"%4�*@�"O�ѳ�膥g��g�_�h<��"O|�	�LN�&�!A��9��i$"O,L��W�x�R��Ё�s� �"Ot(�UG�F��r�#�.01�P"O�����̈�A�'À5�>�إ"O�4B��n���I ,�2-z�;"O� ����8	"���E�΀&o�#"OH��7ꁪ,j�X��9�a���I�~��Z���( v��ԀgGt�ж�Ph�C䉩��؇h��>��
$��I�|��� �[�)�l&��J���.1���2�B�<#�2��ȓF��;�`Z�� ����S�R-�'�2�3�JO�LpfL���#|Ҩ���9�`THgƌ
���Dƍ���M��T�z���г
�<y"F�A�}�Z�'{b
�Z�&R�H� �-�څqK����a�Z�Ə�Gmhq����Z�'�N� �kܖx�C��\�ఄ�~,�\����yl8FN�-;:<�ߴj��93��D���5���O��O8J�'L"|~}ɠ蟖
Ԗ����'�<z�F�z��UNJ
$l�p����An����� 㮸
t��`��-s��Sh֮l�0;Qc���$�?A�GN�\���˂�D�XJ�ċ]&&��ġєc��X�f�Qg��Y�!¹LE��I2eB���2V�`
����ʓ?�bp�C��BT\���C�޵��lƔ:��49ȟ�¤���y�2�H;jS�a�"OB�b1OL�s��p��^�&Sn :��覍Y4�X�m������Cʸ�����w�F;�	�?�8��r��8;o�TQBJ�A�*���R6<� 0B&�$c\����J�Be(�i�� i�Y"�}�ʙ�Dϕ�g�p%P��=��ȵh���.=���z��#^`tF�"Q;;���*&j�<q�I���
D���LD�q�1"�$�� w��&G�NԐ��W��T�q�	0x�x`��ױP��9jr�lӬ8&�ޏM���f�_:FLb��b��ѐTi̬f����Oyʬ��߸c�b}�#QwAZ�s�Xh�`�A����*Lm�eP�]#��rs� Y��Ɇc�B�h��6� ёE�j�ӼTj�(�ck��ʆ@�f�ވ9���*8;�-X�F)��*9>�1`��m	�>aS B։���[�O�H$� �h^7j����<~�L�� CV����%V����K��d��n����N�U�&�V�D�CHbp����)��I����)Q\����'��M�+Rp�<�Mظe�^8���dJ��;xd�V�\�{-����ɸR��uqǌ%%�xx�G�څ.J��EKYq��@R��ǖyc�A��	�S��ם��e �*��p��i>ѯwT�t*6�A�g�2�;#��;�0=	�@_1F���� ����x$��8 �@	�p��Xp���ad �Bd��˔�MN����I�B
�@t�6�5�ΐ?�$̻B�Zm
AI�X�����R|��<�� �z� ��5§a�t���e0Px����	~n��t�ÞHU��'�,j���MQ6�餅�2Vtݲ��d߅*���P�Ύ�+��q;bJuE���!��j<�'��B�'Y�~ǇD�|̠5	�
/�$@����<�謠b�?v�:Q��g�);����	,�n�s�!�r<��fB��yCS������G�|f^P0��42�DP�Q�
"�|�G��C��Q�M������'@��n��f���-Ďt�p��ɳh�ݩ�b�;t
�$ 
	�Xu�NlȆ��6"�eX����I?YFL6Q~Sp ���I��;�^X��aޅ�fh��Cƞ�{q�I	P���))�IH\�۔�	)i�>-!u��<25H#�޹N�Ш�bE� ����5�����P�h�G݂J��j�Q�ă��� s�tñ⒅?����Ѕ�JŀJ>���9���5#"M�Ӌ^\}BLز�(�����a��$ȁ��"��)[��>�����
T�;�
Pr��`!@���7���~%R�n��o$|���y"+��o�����G�}�Ը)!�بd�C�I�N�z�z�j^%ծdkS���Ų$�`{-���c>c���CDќli���`��G����-7��1�� ��b����GX�!�m5e�k� )7�!�C�M��%���3�6�j��� A�!���!sz]T�U+����� k!򤅄]�&�C���(�2/;!�^�i�pQXh�'M1v�XEN�A!!���of$���(�d�C-�<	'!��340�[� Y`>td[b^y !���*�Z�(�n�'�mx��!�]'#l��ĩi�Z|�t�X!�F"Q�.x��固�~عC	
/V6!�:H�K����-v�3Æ�jI!�dQ�1�X�5���l�ti��̖G!�d��DW*`y#�ѽ'�d�1���&0!�dʵ&R�� 0���cЬ����ئ7!�d��Z�2�g��� ����#�!�dG�쨘�ŕ�p�H���a��n�!��mtҔĊ%k�Px⒍�((�!�ű`x �Y���_s�A�䃄h�!�ۮ4�8kuAd�V ��,�!�$P�ur��*�d����ӄ���!��/�J�覉�0`�<� b�x�!�B�`4 �I�����X'�j�"Ox�F-<~9�U���Ƶ\ֵ;7"OL-��ܸ,(@Q�6D
��9�2"O>1P�iΑ���	�&0��s'"OX�1�ҁO���"��o���#��8h���[�d�4�>!�t�ܭ&]1O�`�QɓbIx`@%�T(Jبi��"O��#U�ؤ~�r��ʠ1��xP7"O���TLO�0�HJC�]�"�h�"O�=s0)�/%N���Q�+��|J"O�5+т�x�8V%���q"O���*�=DQ�׷�&Dh!"O�P�p"�4F�� 蚞!z�\��I�!�<� ��)�]��ӃG{���c$X�q��ٍyr%q�q�h��O�V�p$�T!A�6)��{$JqyBEĄ�>�����h>q@��ː.�$x���5M�@��`�>9� ��d��mBb�Oy��I��Rt�qg�$u�*���/t#rp�Qi��v�LZg�B� ���J'G�佬���?�	�jF��;���53��b��B�-"X$�v$�>#�Y;#���v���OD$�a�'P�j[���aS�6J��JPd��Vx ������y�DO+�0|�j
�\F��G��R�P	�A�9��D�e@ĺ.q�FJS�=jd[�?��AG1�4�$�B�j��݂�,)���F��@�(��&˚�*�Ś��ZΟ"~��	"|���Dm��G�64���lNĘ(�'L�H�d�qKS~���ia΍I�8y�#æ݊3�T��ʜt:2����'m��k>+��YLظXp�L��p�Z�3���1rn�c��;��2����3T?Z��Wc\�y�)���/RJ���bJ��`⌄�}x���c��H��%" �T���F��� fT/7�Z��E@^�Z�/.HHRCخo}���ȓ�Dq2� _��K �ݣj���ȓ]�T��BX#�Υ��=kR��n�����Z���yCoҾR�4 �ȓ��m�b�K�P��dL�7y��E�ȓM����)	�<�X!��N(�XՇȓwt:�a�n�m���@���
G�,�ȓS�����B�v/4��J�?"�x���xh��u�
uK��k�.ŐA���ȓ;���iu�҆s-�P���R�r"nЄȓ0���6"ܿjN��y���30Є������I�Mj��P��+�,��4�ء*V�ץ"�����!Z�rs�8�ȓ�v #�(�p�H��I�~��ȓ]^H*v�:O�%u��VB�X��Q�j "U��
q�&ᢶ$Mnt�ȓD3� [���E�����Iمt� ���S�? �=��dY#ZR�д��,'���J7"O�q@��WF���5+�|�"Op�����V5 nU%R$(5b�"Ov�x�B�6/��X�L�gE9$"OVx�O�"�`m��hU�`�X�Z�"O�:��X���j��&8����"Ob�Q��Q�\E
H�`OH�<!�R"O�h�f�ڮf��u��M�'z�<�"O��҅�^
2�`B�ԗ;R ���"O��� ��7�ҹ�c�R�m��mX�"O�Ÿ��.pspE�&� 0�`-��"O������![���G�;D�z�y�"O�!t*4 �-��EO�U��\��"ORHr�e��k���H�l��k�"O�d�&oX��)Hf�U�M���r"Opx�` ��F�V�����P[�ܛ�"O����(�L|[TF7+���PS"Ov��k��V�	 "Ś�:@��R�"O���,xzLm��Ê�59�@G"O��1��#`�4iq��F֝P�"Obp:�#V9=�PqG� mx�'"O��WbM�&m����U�
4��"O\�à#���`؁��If"O����o��<��MQ�> fQ��"O؀��@�|&�8��<.� a�"O<� *H�OlEaD���f�T	*�"O��`v�@��$�R
�;Ubt���"O���t��W���bFۭk�&q�'"O�q�ӮȈs� �3⥟7U�	��"Oqx&�8�<`(�N��[HS0!�$ٽ6'��RaU1;�n�h�V.
�!�d˄I��P���^v�0m�THBu!�S0���{��ŷL R"'��6`!���TA���˒n"�tbq��~;!��XN���4�':�����v0!��ɐ�����K�t�r$��%!���k���q���fЀ�%B9a!�:f�T�c���!%-<%R��]!�U>R��< qN,`�1`�e�!������ЭJM�A`��T%9♄�@"N�Р�\��TH䁋�P�N,��e�D	�#U�N�,�����h��U�ȓA��k��a���u%^��F5�ȓ���B�U�|��R��Q�K��\�ȓ�<U[�`I�L}6 ���4xT���4�����ca:3/I=>lZ�ȓA:�i�2 �[T�J鋺����lс�����f��QP�@��U�V�"7oŝ�J�YbHe�*��ȓ6�B�#�P�	�i`�l�Ԇ�c�^t��ư�d�F�ψq�*���d��R�D9'H+eH�W����#,����GV���L nk����k����F	q�Ȝ�E�6 �t���O!��s�X!%���0��H����;!��:Va�{���(�
J$}~ąȓq���զ��P�t���YXb(��13"�w�׭AyH���
N�r
�I�ȓU��pAڨ�\Q!�_j~����1i�!"^� ��آ 
�6�t<�ȓ_�����ќ;�D8Q�Ϛ�d�T%�ȓqA�Ԋ�獭qN�8 �\Ay�ȓr�t�c�V9��k��l����+��}�%����
���A�X!�T��S�? nػuŘBŀ�%΍2>2��"O A���M"5��e�{"̴��"O� A�I�O�\�d��>*20��"O8%�Qb2 �X�@%A����"O@(�@f)�rBZ��8Qa"OP�C��G>n���W�Cr@4"O`i)��V8.��ړ���JcR�t"O"Ek��0 �*��hїkC�\�t"OĀ	���&"�L�,KFz�q�"O�U��GR�@s��E��. �Ac"OTLpr���h6"�1&���C���"O}��F18ׂjp)��i	�"O� ���R9�R�B	�77ޞ(�q"O.�r6lL���(�X�{� m��"O����G7	1t��t��h� @a�"O�xB��|S�
(�\Q�"O%#�':RX*�j􀃼jV��K�"O��d0@��4�6��8/n��� "O���hݱ���+4���{N�)�"O�l �9zu8<��B��?�|H5"O@}ժJIA�]�a�'+�a��"O�	q�l݀S)�}{��Ũm%�!W"O^�ۂem�u[�nߺq�V	�f"OHԙ3&��~��`OF&{�pl�f"O"|2'JP"b�4+tl�If"O��r#_ 2Ґ�jv�ؙ+��L%"O��d���:��@;�ƌ�U��8�"O^�b�BP�Q���[t���Ѻ�"OR)��� �7��	��U O~�Lڧ"O��h�H�x��຀d�([�1XT"ObiBr)���42BiNU�Ȩr�"O6�"�E��r�Av)=Ԕ*�"O� ����>\��d'"��A�"O���Ԯ�@> ��+Q&W�)y'"O���
�I�tf)V"}Иݓ�"O
�u�A�O�1x��Ղ3�ġ�b"O�MX1d����{$��B�v ��"O�`d������JS��k�4Ȣ�"O"�3��å,+n%@��B���#�"O���s�O>v4Lb0�Z��8s"O��+f-�(5`�n[�|լ�I�"O��"�;X�A�'_�skJD"O��1�+�+xؖI9����L\^�z"OԸ��$G�u�� ���=��"O:�i��]�(xJh
��rLC�"O��T�Ǻz��A�G�����S"O�0��ΈFD��h���J�V�R"O�B�N$��i�q �H����Q"O�X
�/�9hL�a����K�,�""O�q���
� 4r��]�d�2�*O��C�§��P�&"_�W�����'{��	�&\�r�١�
�C& ��'|(q��ш���3g�̇6St-;�'��	�ŗ��r����Y�-~M@�'ڸ���B�\�|�S��ƵR݊�Q�'�pQ�BI�84d##@�EuT��'9x(U���/��b˖(;�
i��'�TP%�@���kr�V4qd���'���i��v�`�.[�G޵@�'�0$��>�p��G.�cq���	�'�a�dC�go`Ӷ��&&�s	�'����"�d���B�#��}
�'y��x����(��1 0�m�r�'���hUg�BԤ��7�>������ v��Ӫ�%����0ML�YL��a"O ��F	F�T��L��BW#;1���W"O��	6*I�1;8iy��! hŐ�"O+%��ff ����D5	="\��"O�ɺ"�R #X�H��>B.R�"Ox�P�ɟ9>������^.Jh�#�"O6lc�&� MZ;S�V�\*�	c"O�axvִw�:��.��ZI���#"O<P9�b�^�F1�_B,�!�"O�$� ��>M"����)\'����"O�0�1�X;y�T�i�k�5z���#"O�RI	"R@�Ck�*Z^P��"O�]�CZ��x�i�0��%�4"O&��U�C9@u
4�Q�!�rC""O��-S�*�*"$�#���}z!��ҭ8����N���Xi�O��B!��>���3g\�Q��p�O�=!�$�]>Bi�䎋EDL){sO�v8!�E�*C옊�D�:��[dn ��!�Dö���C����H����s���*�!�'�p��Oӕ��亓��&�!��R��YA+�f��D�k˫@�!�T�PPDP ��q���IѣO��U��C�,X���"�Ke�KHd쬅�jR*%���.���'O�-_z-��5n���
��+arUC�^�c\��q����(1ex[e��� �����!�ڢm���B��&�n9��sk���*E���(�o��d<��&�&�����vn,8sr�ðkc��ȓ��[BI'���ɂ�Y,+�=��xH�
7�Q�Xɰe9�C*@L���#q�ِn*~���Bcݚ0�d��ȓcni��f�����"���E(d�ȓ.�$�Gϝ01l�j��K�d�J��b�ܹhQÔ�Qg���D�d��M��Цb�~��Esd�	i��ȓ}�����N�d��%]-(aR���;�� �Yu����g�W�_�p�ȓ-�J��1���V	iA�#W�4��+�1;q!]�֐ ���Z��ȓD���`��פ7����hκLԄ�pg��� �\�0ɶMZ��
Uf���"�r��+,�.i�2�J�z�T��ȓ����� �q�Э*f�
��U�ȓ&����W>{�@P�&���@Ѕȓ �\y����\Z�q:��9�*��ȓ<x�!�F�ЇF@���E��dY�<��:��a!�߃7v^A�+GeN���h�����[�*8��G�;�.���BH�<{p!��"�f={V��N�����w3�Py�]�<���)0���_2mc'd҇!�$�h�郆Kd���a3
���9��cWLFv���ȓ���:����j���-�3D��u�ȓJ���  @�?