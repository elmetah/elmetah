MPQ    ŉ    h�  h                                                                                 �bI=�dʎ'Y��u�l2uWɭ�zڜL��x����L+W��C��&����P��(N� *�S��Y�5y����c�s������썵�Ů��a���6��8hf��D��<:9�/�ii��Z��*�F����,r�`��A��P��\�d�f��(�H�Wh"^U�f�~�)U�
r_ǰ�2�I��d��T�����C��y���>��X'�5#��Ș@�l��$��p�ª����Nw|�/�G�p��Y � �N��,�m1s��3D�:?D�r/��@��gk�F�a���}����6���z����K��\H��ƶ��ޱךOc"����|��.��2��s�E�s!�w>�_)�K�<���񋝴8���_󽰙U6tIh�Md���%/^�y���T�ˣ���GZ�?2�'?_'���ߛ%�ѾBT�o�8[�s��8���7 �_�P1��tRu\���t�˻^|-��@�(�<ac�O���ލe�T�Q����vZ��2��AaS�c�X�]��W����,I�X��Wi��Qy�S6-mwZUSb���b�M�k/������}��<��򄃁RaKN�Y\q`{�H�N�e�
�?�9�D���)����qS�����ǲo}����(�E�S�%�@:ʔ*v.Qt%��C�#�{����xߴ�{�%���[�5�9���1l
S��&�����������}g9wI �����XI�G;~��=�I�r¿4q����NS�X��-Y��S�T�I�P�g�9�}�b3��=�	�+����㫺(x���}��?ӛ�!��3��	�0�\���}�'s�2y�KK�꥽&��H�KN@�_��+���"UѠ[ќ�p�G����+����]��"��Y���R9c_DTuQ��+�����'�����UGd|��FCoj�%����<�z��*i�)�e��xW�tc0s�E��N��ˇ_��,ʮ��j��v���07����iѶodxo^ࡁ#Ϥ�x-�>��s�G��������t��H٣���V�H=��P[i1L�U�������<N�'����UB�y�q���������%:< �S�$fǧ�3�qOI}6���)�r�j��6�x]�Rz{�XN���S�*G(g�$i�*�T�cq��_i3���Z^�����If�����(ꁘ��������hՉ�.NU�IN��3�J�����V5�/kS��Z�ʃ��ըY {�c��~�k�fII%��As�7c�B�6)���l��!�\࿯�uwLRdY�Gh�'CFhB�WV<���r�-�#��5F�"�:^��s�w�+�Pc�����ؖ��Ԏ�}C0� !Қ��Nq;���������E3���GQO��1�����_�@�{�/L ��k�S���|����65S���2��;^o��O����-���T����#�
��#M^�l���&k�����o��*'舸	�QC�o�����J�$e$�E�U�1����"E�����8ۓh����u�S���������+��Cr��b)�uLž�Cz����E�G�9���ŕ�)�tj��*���O��=��1�W"�'�TJ�����쳖��OM	�@`�1\��Y˵Fp����C���gؖ�j�R ��������hף㹹�pLׇE�ݥ�]j��a���/�������{�m�����y�wv�%*��8VP4:-K�Gݕ��1�y*�{�37nn�&
*yFYe�����J��zڑ�w�$��砘�Ώs���~�fevr��:Z�'l��D�E���c�2�����R�3�^��TI{��XY�DQ�3�s�R�FT�$���1e����$�"�i*�^�Kx[��g���W�d=��4�V�D20�n}VJ�.z;ϸIs[,�Ճc���ܻ俜.S�=�1��X)$�KR�"�Cڂd�	��_��]�_ysOA_���.c~P&�A?�yd�8\}�<c�͆D
li�F
�����2�K��u����92 ���+-7�	l��/#����������P��K�7{w�`Ѭ}�(�@�h&u!1}���]�L9���k	�.�I��9�#_�߅�-P���*�e�߁��Xi}��d�]|��݊�%u���W5e�pA��,���� �1U�u�M�x� ��g�K��'Ϸ�;ר��Ǩ�OcK��&�]F��p���lD$ۘ�T�Mu���Qә�
���2bMo���as/lEi�L��-��\���ضVL�X6�%�̝��?bV���+����G}��$��IKӂ��5�CHe,zD+ܶ�Zjw�Ja�A���,~�&C:��i�h���1}���4����G���D+��u0_���j!��\;U	��s̓�� W_��� ���Ƌ$8�iO�1a�K���sLV����̥APjD��_[�ҷy�]��"ӈ��.w�7���WMT]��B}/~BB�-Y�iK�%��F�P�7�T>�,�c��OA\A�9��[jC�.��b�_�$%��@uFo�vOQD��S�`��.OB��%\�%�:��>67��V�	K�R�#kTE[t;*��U���+��;�~q�9�34�
�� �%��κ��Z�G.�)������F8��'�-��>�����O����7�.�K0�����3*���*s�d쫤� �'�����T�Ȟ�ް���鹯����g���h �&�����J���``]_�����w�۩�Y�����x�u�(���?m�����Y�|%���I7ɲ(����)�ZֶƳvr�OD��O�?]������٢�8l�x-诸��s�/5�q��3�|Oc.���1�e�H��RA��[��'�E$ɹX���T<�Í|`�߹��xOk�E�N��;J��y�V �ڔ��j�'�5D������+$�T3�E�'*�ZzVσ�B��e`�u���{ ��	08Z,[�\��X�y�qH̓��f
��"t��Q����B�i�ER≴F�-&D����g����M]�e3���R T(�'�)=��M[�,��QT�=�P�7��s�u2QQ�
I v�k��>8���\5)�����x���aI��\qp��_��i�2�,5/���F>*�)�f�Xh�M3g�k/�|��r���֭ܰ�_K�k>)���! �C��n¢�M3�ϥ�H\W�9�9�̔�HK��7{Gf�{������zl�>	9��BA�M�CY��w'��SV��,#������T�Q_�F����x�w�@�/k������� �&t �m̭'���W�����-(�Q�ŏz;�!x4��} B2��O�&�8��B0�7F���fE��k�񧾂GɊ����Onr�-��7�|Et���箍ZE%�5�r-._��m�����
�Z�/-���~'���QU�Zh�dm�0��S)��{ݩ�G��~�)�?�<ZP�ȉ"Ŀ'�A�VϺ��e�Tl,0��,�T���>��h*7{2�Ɋ��uu����_����~|-�	�@�C<�ݛ�
����
��Õ�y��v�!�2aw�aNli��� ��1o���,�6��f2e�����3�mr,z%'b����,��M�cOk
�ţ�گK�$����d�<��af�hY�r�{|y�N� 
z.9����b��b�_qnE�$�����+o�$��_g�E��Z��):�>vIe�%?�C��u{
\e����v���qf�[v=p9ۗ1��nS�5�&Y�a�����[��\g��*I;��܋�X$�VGv���p=��%��C\o��Nn������x�S �^�䉫�b�����"3��cX�e	��X+�����q7���������?�ϴ!mȴ��0�:<��}Y�M�-ME���h�`|Q&�+x�Ƨb�:LA+>-����ĠV�)�G�T���ܬ]��M��{�<���M�|_���0&,��*�s�R���	�4U�eQ��{�ošA�Z�J��q����Q��d��e�ZxR�ot�/_�S0*�i���Fq��a���mj-����.7n���5�ќFd�?��|a��ߙ-s���}	�G��!�\�3���nd�؝ۑ��=��8PV�#L=8���H ��	��v�.��|�@��Bn�q��(E��ǋ� ���<{���F���/<�K}1�  �rf�Q��]NO{��i����xu(bQ�$Ġ���Gq���i��9�5>�^�0��(IaJ+�#B�E� ����4^�����{ݬ�U�<�Q�JJx�p����56kS�_V��\�p�k v��R1ky46I@o�Acpz�6dт�!�!�J=�
Ppw��Y���좶h��W�z��Ux1-�ܚϐp"��H^�N_&6.+��~cKЍ�q��ؑ<����C�7I!���6Xp;�
�jk�`���@����uOюQ1���B�t@�_/�_3��(}ւ��QW���6Po��b�tQ�;��-�z�b��Ў��
`edF�����j��5�o���� Ѽ�o�Kq'�#�	�C���0[�@�96e���P'�&����j��鳽)�n�d�_>u�	���Cڄ/���Q;�^:/���P�P��Uz�z*��@�TG�i}�|e���~t��/��ߊ��=�]��,g�W}�<���!Vʕ%#��q3��L�M��`.�\���p�}�#R��=�>ë���"@R��;��b��gG�^�n��w�LR�ȸ�+��,�IkQ�.�/ܛX�I A��L\m5�ʋ|��òC%�e�8Q'�4�4ߣЪ��{�y�S��tn��*�vY`f;��1�H���� $Y�s�m��u��^e�tC?pZ�0M�e�EMc��'� �Z��.���T��{���Y�ODQ�sy��F��=���1��
�d�:AiEP�٥'x6�g�i��8=��߱zF2���n�7=m3�;�Lys�;��Z��ঞ��jS>r�1�e�)�s�K�k]���� 	����:�Z_43�AzEGԩ�P֛?����(��X�(��
'�wF%\e������<K�W)��4]��&�+�	�U`D#gJ�2�`��Lp�K�^a �76f���F����(�+� �Wu�>���o�����W��j�������P#������������������s��ٔ����(�d�G	5��:�W�F�@ro��eׄa.� ���U�^M������g.���[=�V�ߥ�n��*���'��]�i�p���l��q�S͌�h#��$���t�E��1�b蓓���/����Q��H��\I7�ؑC�Ǔ�:%�<�+�?�8�LY�����}<n�e�Lӽg#52
H`z D��&�#�e1������[(~��:��i�[�ku���549�İ|5Q���\��T�u+CITT�j��*��U�`Ds�Z�[��"S �|�u:�ߑ_ijy�a\ �����VڴJBs�AK��L����y��|1"�o��w'կ��MO�A���B8��~]��-���K�C����G��ON��k;�c���Aw�9\�[E��.ؙ����/ ���o��Q_?G�04`j݁O}�����~%{��Ǚ���MV2�,~�#F�[�1D�TD�ӆ��j�;�Y��b3�d���»�C��
����G�-F)̖��8y8mó'�9�� ����@�H���C�@.�4U݋������3e�v��ͨ_�E�q��mdo���k����������#��ޜigQ�&#�=Axp�H�Tx���@�\]��w��Y�w�B��ի0�I=����2�#��m>���.|�N��V'��ͽ�+���]�:��crU�١�M�?��Q�dc�ٽ{�l`�l芫׮%^5#���.�wO��o�ހ8�c!�n�k��%E�IOX��T����H�Z��D��h � 3���BJ.Ǎy��+',Ϯ��B9�D�j2���v�$�7T���zo�'�
�zd�]	&e�=̃�ݻ���H��03O�,�X#�Bxsy/,lq�,��/'fE6�"" Q�l	�� ���H��kȘ�͇��R��,]���S��R��G�B�/=[u[\�ɓ��=�؎m�r���ysD6�Ql��I�Q�k�0�>sQ����])�
��bZ+�adB�ח�p��_(}`����5*�m�*��*m �f/1��_q3�'kj]B�q������c<KNͭ)�"�!{�OC��������Z�'���̪W��>9����\H&��7�[��G�؁�	�6'`�>$���r��j�3CP6���N7W�BD5#`���,��b&�|�%��v���vt��[�w2�}/&Ch�S�O�	 a;L�mg���nG������@c!���
����w>Ԕ}������-w�y�A�Ra�R�N�f;��,�!���N��>O���\��R�]|�������dE����m<_�uO��:�%�q��A���"��3��Ulahޗdȶ\ӛ�ر�Wu�J�Z�Y<)�z�%Z�׉i�'h8���T�-bT��|�������!0���m7֡������2�?uR��:�"�1��-%QB@�~a<x��Ń|����J��T9�v�l�2�)AaIrK�gC����Ġ�,?¡�A-ї=����Q�mm�E�{b^ٲ�G(M:�k�% �7<?�n��T�n	��?ka��\YR�4{W�@N./

9}�/׽���q��i�hp���to�����*E�޽��i�:@�5vd��%��C�Q�{E�ݮR��q�����[1e*9�� 1b�QSb�	&�|�52�����td[g�LIV���bLX���G����s��xE��5n*�	N��@�y>:S�S[=�����]-��3�B3s��s�	z��+uA� 7�^C���?�3c�?I#!+8e�vF�0j8wN}��@�(A����[-&����A!���^+y�w�X��Q`������J���M+�f���5�w�ǒ�Ҳ�H-�_����,�$)��"ݎo�DsFU}����Щo �]�c���舭����v���e9��xM�wtOk�;���H����.۲�~���*j�wt��y�7�X�������9dn0L�Wa����-䶥x��GGZ�����'R�����H�̸|="~�PQKL��R�h���-{��)����{�B	�;q�4��j�F����!<�e��G��K��v�},��v��r!Α�l��]�k�{��U��A(�(]35$�ғ�q���i)dH���^	@vRd5I\���~�/� �[��cL�歐e�a�/��G�QU����$J3ay����5�
Sq��@���(6 q2�����k4"gI[�Ai��cK�j6�$����!�Xv�e�w�#iY�G�J�h��eW�� ��-������"M��^�R��+\T=c�9"��،��DnC��!GX���;�c�=������;���T�O���1�e�Ľ(�@�c�/�ް��bVx]�2�x�n:g6k�E�!�O n;�ch��Ք��& ����Ý� ��������\�EѷX�oK�'^�	�UK�e�6����{eZ���K�����Ҙ�����ɿ�I�B*�u&��ܩ����"��y"f�X�d�+�w��0Iz�ef�;'GJ���7]���=t�������a�=F��'c�W�s����<̕��3�L�1�ǨM?d;`�|\9��+
O�>�����3Æ�$�F��R6EЁ���Q9���yL͖oȓ�Y��q����/7�������ˈm�J��WL���0~%`��8LOR4�[�������y a����n�)*��_Y[YD�_0Y����3f$�Q��N�\��x��A/e��Q��ZFY��.��E�SNcjx��[�+��v!�P%���{WD|Y�z�Q�0�sT�F���0:1��b�v7J���i`*��T/x�g8�ō��=����y2���n�8x�Wd;� ys�j�չp��ې��uφS��E1�Q�)��K�����ڸG�	�G����_��A�_�$�P��?-䦝n�귃e�
�iF@�����|KOkޭ�%�/���D��+��	� ��:#Bm
�m-�I��F���7��m�p����(�6�[�uWl)��P��5�;c���P�?�S�҄S#�x��3?G��.�#�U���%f�1e�����K����-����W뜳��a���ܪ� �)��c�MH�g���g�.L����q?�w6L��\�b+-]|CLpﻩl�\��ɹ�Rs����O<��1ύb��>����/"�f��{�c�k\Ĕ��lP>��f�%A�#�
��?;ϒ�����}�қ@�����5�%�H[�D��������!(�7�f�⽵~�B:,
�izX�aE�&�!����4�逰WC���"�AEu&G����jy�ئ���U��(s��ϫ��&~ �K?����i�*�a�Ԭ�}�V���9�AF~/ߧ�H�yv��As�J��wb�
�J$�MJq�M�B�.T~x0�-OH�K���<	���J~��j�cl�oA��9�[ ��.����f�+��	5or�Qz���4G`E�$O����[!%%v��� �uHV5zk�ɿ#!�B[�Gҽ������4;F�-�Jr/��3��.-��V�y��f��M��G�t�)純��Z 8H�'fB�t����m�������S.�=����{rY3�`;�Z�;��ި(���Ñk��#~L��&�4�����Y�g�@�ޯ�\Wʔ�K�S�*�{�l]�Ց���wZ�\ʐ��&�n�����	^$�m�[@��� |� 4�%���rG��)p�8
�<Z�r��G��k%?�\��(���l۟��e���� 5����)�nO��*Wޛ�/���I�r�#�EZ��X�>oT�2N�������n�����o�Z$8J��3y�4��w��i�,�]�>D������_*�!��u��'���z�%�xU�eV���c���4��~!0.d&,���yJc�q>&�ƙ�f��>"�nQ�L$���7���c��jV#����
��52�'�]ɛ����Rvߪ�]��=�%�[7�O��l{�s�b��8'Bs�lQ��xIM�k��*>�S��0�)�K8�wn��sa%`�R�9p��l_cN�h��5%��ׅ=�*(��fJ�[^��3��hk�9�����d5�f�K	O�)�۔!��jCt9:�pV҃���v����Ww�I9b�̊�]H�
7�D��5O�Ep�d����>?����E��C�3U��Pu�Io���{y#��������W�!r�|����^�w��D/�������_ <6R�~m����<�K��ڣyZ<ѠŅ����)y�}V������5�4���m�V�̓d�A�n�g��}J+���yO$�7S�g�m��|���~��$�"E[F�hk*_:��m��@�Н%vλr�&�n>U�yhّd#�h�V�k��Su��&Z�4���Z��]�.�'Ü$�̎��"�Tb�U��� �����hM711t�?`��M��u���c��l-���@��b<r2����@�/eہ�d��/�Hv�22���aD�	�iLƷN3ʙ�H�,�m��H��xT;�$�/mh�[0&Ob��b�M}0�k��ʣr�b�4���D���a�hyY���{2;uNi��
�9xy��T��0Dq��C���w��o.3*͕D�E�0}�6��:�jv�5%5��Csw{����I<��l�:�'��[��9��1��S=�\&�)��І��i���Kzgj�Iq�;܁χX��xG�Fz��L�+!�EH��Y�N��`���\.��S� p����X��Ď9�3.t���	���+P{�<����� ����i?��!F#
��#0EV��'}��K�#U��\�c��Y�&ѷOռ�+��,+�����7S�L?���Knx��A�K�kY�ֲ���*���C��_Uk��/�"Џ�i�^��1�mLU�c��Eo{�y���������P˻f�ڗ�e�>_xH"tt����en���Ĺ<x�ۍ+!�0�jc�����^7$ø�O��W�d�@u�2��U��-�fI�s��G��<����B���d�������=�k�PL��L󘑻#���4pk�l��������B�#~q�'�j��$���O�<qW긵h,�3��B:�}'�Z�0rܯ����]D�2{i\�=Cw�V�(X5�$z���{�qї�i����^D�����IW�����@������Rj���@������۷U����J�㥆ԄY5,(oSL�݋{\��� l���f�k�/�Iv��A�a�c&JG6ڗ�=��!Æ���
�w}��Y��2��fh��=WWݵ��-����F/"!�^)eN +7"�c��Jŧ�؇��ԟX�Cau�!#��,��;i��xrVʖ��6�}��2�OG��1��M�8��@n��/�}�<��sj���dz�)��6��Y*�;���{���>s�����
'�{�B�Z��t�� ѲHLo�
_'�z	��K���������e��2�F}�����S��P��5�$xpeֹu�Nn��/��M��\�є*����d�]y��zz`��6x�G�*P��؏��t�n��&� C�=�Nz�"�W3H����W���F��'�K�³�M��`�|\�����Y��3�t�a{�����R�#��¦F�*���ل�)��LHΦ�n�w�T�_��/��Ђ�O���j=m+�ϋ2S�(>�%���8G��4K�g�xA�&p�y��՛�M	n?*JYVl	������S�Nws$j��)Λ�$���O��e��Y�Z�;�I�EC�lcEK���q�#l��n
NE{�Y���Q�3s/l)F�+�~�1�`���*M���,i{`B��xcx��gB|��(�=�/�g��2K��n�Y�c�K;`�Hs���T���֚x���S�;�1�]�)�r�K�nJ�Km�S�	����Z=_�#A��ԟ��P�	�?hIf�	"�����
��~F[ K����QK��୍�u�*
���C+^�	�Ϩ!�#����M�����A7���7���(�wO(�a���u�s��Q%�]:I���E��ͺ���Z�#
���昆���vn�Fᩳي�'���Ά|��}0]��H�WF{���18��WG� eU���
�M�c��e�g��e�X��������@������ݸ]=Np���lU)?��\	�����/��*��l�Yb=����/}��ǔ	�~ٵ\?F�G}��	/�%ܻ���?s]�����1��}2�Z�q@�3�5h` HVvD<d'������1������@�~Za�:ǯ�iu�N�����\��Ӥ4/HI�2qi�O�|��U�u!k
{�j4�*�ޮ~Uz�9s^�������� �:.+��U�hi��aR� �X��VP��x �AA8/�쟗��y02J'�e�%�w�����usME���'B���~�ׇ-��gK���w&��!�?�E��!�c'6A���9���[�q.N�g�0'V �Q��o-hWQ���&UV` O�� ����%q�T�O�_0�-VP��"5�#��i[%~Խ������p� �;������3�PTnc��[���⸏��^G_�v)�˼.\8#'Q�'�����ן�#1�*.gw݁RI�VN�3�r��y��U�'0=�=��ޥY�a��Y�Y�aGi��V���6�g�I���wV��>..���G�]0�C����w�q��K��������{ӹ�}��qmt���R�|6Ӱ��B��HB�!�����w�:r������(?n���ڔ�����lVc��@��$"5Y��$�aOtG��>0޶>/�Y��$�	�^�vE���X��TM��þX<�0Q������$����Jd�y��6����$4�x/Dv���[%ѯ�������p#�';=�z��K����e�����B�,�)~��0)��,lᰛ��ye�~q�`���#f���"EۚQ�L��S�Χv�ډ���V՘~Mw�F��t�]�f��	�R1UR�x�=Q��[l%�H��/�~�|js��Q��I�h�kt&�>��=�-��)��u����"�a�(���D�p��_�?
���5 ����N*�fe�٢<3��Zk�5�ͧ����[����5K���)紀!q��COŀxn��4����Y��W2�897&����H�� 7,!�L����گ�ή��]>Z�
�h�H ��C�PҥH��D�-����#�:}4A��X��2�B�\�j����Ӂrw�gL/���=�E� n��9�m����*���4��^ҵWAg� u4��L�0}��~�Z2�7�t���و���HB��7�Ƣ#�����&�O�
��x|�N�YV�_*�E�!Ľc��_��S�(��[�w���[�M�^�mrU��9hԫHd~IU����oݩ@���:�����Z!F\��'!�߇���=�T݋�Ф*��MW4����7��e�����h}�uH3b��G2˧��-[@�@�T <�"�;�H�JB�@�*�
9vFc�22�a?ޣ��Q��	���D,59�����������umc�m�V�b�0�}n@M�F3k��%��^����$�Ńm�^a��YH7�{�YN�Vh
KNj9s ��s�F���\q��f���R�voi�:�0�!E瑬&:�G�v�a�%��CN��{�B��E��g:삛r[��9,U�1XT�S��&
���k�|�q�*S�g%I�Z��\oX�RG'{���h�����zR��vN��H�o�K	iOS��v��	��SIC�閣3�|����	p��++<�wܒ������i|��S�?�*8!a.��lr0 ��� �}*�n�����X��x�&���7t��˦�+��9����G>��X*3~e�-��O�F���M�ş��>��_�t�ad��=�^��,������FU�*���� o�ޕ�&� 7��$�˖Pp��eo�xC�\t���㄰F��l���]��h��k�@j��R����7M0�
Wt�"�xddqj���ϐ�-D	��n�oG��ښ�M�]"���v�i�f�B%�=XyPG��LNyP�ޫD�O�c�������B?��q�,�Vv�Ǽ�ɩ�v<�h����n�]��}"3b,C"r��?��-]��{DH��x��I�(SW�$�d��@Mq�wi���ƢU^����IR�r�4�R�v�݁b|��>T
��} �U�i��bQ7J�����~�5�esS'�i�����A'� g-�cH�k�]�I���A_�\c�s6+��ذa!��|��w8u�Y�F���h��WB�-�&Iv-��yϡg,"�d�^D R�1{+kc�k�B�n؂�����CD�!>s��4v;Du��&Z�1 ��1/?�
��O<�1hbĳq�@I�	/8=(�׏�n�%��\���6��H� >��;Jع�K�n��?��W��S$��q8��	����X�o���XѭXQo'Գ	��[%D��6z�e�l��AXd7i��_AJ��jw��g����u\�'�����@��$>ѯR��NQ�����z����1�G �y��t��'��t��(�;D�=Qw���,W��=�@%��r�G��+�����Muk`�\�f�ˡM>�t������<����Rl"��x+<$׏�D�"L�%J�I��I3+H���/���z���)zm�o����ckx%���8B��4�
\�3hA�y�����GnzG*�YZYQ���5h�y1��iI$��?�+�_�r��vXe�TQZ�
I�d�aE�:wc >��[*�����´e6D{��Y1;Q���s

�F@Tf�"1��g�,>��k]2i����J��x��,g}��Ûw=�m�����2�<n��� ;;��sG)<���:���o�+�_So�41�X)�!�K}�Ƹ���	�çK�_e2�A�*'���P�S
?��9��N��|�9Ċ
XT�Fv��Z�^FTK�k�(�~�%�%����+N�	ؼ~��#��{��4²���<��r��7gH���*�(e���A�u�'���r���z���aT��5��P	#K�m�iО���M����"��a����z N��8�tŹ��XW��q7��L�R��� @�����M~������g?�_��&��'��m%�û~.�د8]�V�p�5�l��ۄ�M�������`X��i9b��]���/���炗�ə3�\����"���D�%w�[� t?Ο�}�<�L�}�ǯ��h2�n�5�oHQ$<D�ѷ�F���a�-򈫘� ~�_:buUip*�$��� ס�04����͟��j�w�Iu��e>�j�!���:U�\vs9�˫�z\�Q �IY��y�_�i��a����3CvV��'�A<��]w��
�yKM��È 7w� �Հ�lM@1D�DBi��~���-E}K�����[M�}r�@>��|)vc�a A�I�9uܹ[�o.��&��n�Q���$o�M�Q���䡕1`�l[O.���f�%l��Ǫ�-�	�Vkj,���#� [`�J�%�ę��{�;��c�c%��3��i��}�.��~���Gb)Q+��}j8�U�'�����n��j|�Yj��t��.0�t�����1Jq3�ԕ���P�;���������ٯ��r�4zޜɑ�U ���3�gbY�T߀�u��0�	k�����]����Q�w9��dl��d�Ӕ�!�4�m{����9|��m뇀�=��:���9H���$r&����?ɪ���]"���l�F��D4�_С5�e��POϏ梠����	7��L����0�L}E���X��T��^�y7#�K��duȻ��P�Ќ?J�I(y��8�r��t����gD�W4�6y��ըj%oI�k��'�azB�V��M*eLY�rA�g���0$�",��w�s�Wy�1�q4���|ͥf��4"�g�Q�l.ﮭ��1�u� ��]�Y��S���]l�]�Q��d5"R��=��k�=��$[�kK�=C���V��4U���su86Q��I��kO�>$��ȫ4)�-��-���*a�K��H˜p�W-_�P����5eN�;��*�D f���Tt�3p��kR��BA���r���RK��)��!�ǄC*q�Z�Zҹ���m@����W�@9R
̀]�H�0'7gP�����kX��>u���Lc��VC�c���N�??�SJb#���O�-�Ӿ'E���l����wC
�/W�O�⾤�Jp ��p��nm8����8?���Kur��{�����}�ސ3v���3����٣r�� �����݌Â�K,��ʚO��}ɨr�mA|+D�4��皞�E���^)_� v��'�vGg�?5�(�f���zU=5Rh��md��!��&?� ���������Ǟ+�Z�Ӊ'y��B�:�XBTX�����@��p�����7�w���Bƃ��uÈ���L��?�-���@��<(ϫ����e?��������	v�2��a:D�w�Ĵ����,�$z��ݵ��V�Zj�m^|�wb��A��AjMs}�kv���f�ȣ��&�(��a��*Yø�{�|�N�"�
��9n��΀.�N�8q�)�nˀ-S0o���ˡ�E�4��}�:qDuv��%+��C)9{�$��o��bh��ݗY[b�q9G�.1ӶCS�<4&E��������zg�$bI�l �w
X�|[Gb��D�<~����$[u�N�C�����piS�ѵPt��Nl�D�3��K�J	��+������/d�����D�<?z�!|Yl���0��U(:�}�*���)�,��L��&��ղM���+*�(�)o B]圳(��Gr�H�D�
t!�E�(�Β`���9�{_�v���X���_�nK����4UN�Vͽ�fo13��F���;y����qZP�e
��x>9t*mP�?C��.0�2cp�Cu���&�j�֙��~7�����L!�=��d��+�� ���F�-����i�
GXzؚHμ�x�M�Z�D	��}��=�\PB��L�y����c�jVd�b})�n�҆,�B�4Kq�ؖ����w1��*j<g���k
���`�x!�}�����rR�<��`�]:�{T���1^��(N�5$0�ߓ���q �i�Z���Y^��#�+IM���3d�1�$��>���������ELU�A��(qJdIk�
��5"�#S�%������ b�u��J$ke��I��qAڒ�cܙ�6P���s��!�BJ�vEw�M�Y�B��nh�y>W}�����-� g����"~ȭ^_�]p+��c75X�݇��}���U?�C�2T!Y9d"�%;.W����{H�,�<�eofO��n1!��.Fw@$/W/s"�rV�i~�C����6���	 ����;��Н�b������[{Q������qtKj�3擄~�-:FѨ��o\I�'�ΰ	.LD��ڢ�X�qz�e+t��<S��f+��Am!��	k���w��̅u���͛���8���T�ʚ{��M)뼲̾A8z��1�,zJG[k#�h0��B�t���q�w�veN=쿤�wW�Ӫ�k���ݶ��8��MX`
1\JmI�\\���i�)���Ӱ��>�RA���jlbm��Js+�_�L>�Y�$h���u���N��ac/HMI�5�G�	?m!2��!5Þ�%1x8=�h4�p���g�\��y��Ûz��n��`*��kYL���p�O�4/�����$�����}
��B?�A�e����Zw���%E9�mc�P���W�Y������>�{�Y1��Q��s���F{�j��1�χq3�&��i�,����Ox�g@g�d2�^�=��W�4�2���n��Y��;�Xs���Պt�����S*��1�\)y�1KX��I`�ډ��	�&R��� _ roA�a�ԕ��Pm��?�s!�?���\G����
F�$�����9[�K ���G?� I��U��+ԣ4	��R�a�#�L,������7��R7")�#�-�m&�(@��u(���۳A����lF&7BͰ$n�cf�#�����n�|��,e�����/�ـ�0�U���슳�e���W�_J,���g�a�M�g [�A��M�b���g�r9���<���ͥ�LlÖ����]M��p��l"�?l��ԟ�����!Ԧ�f-bTfё�9�/3��=��ɴ�B\5mm��6�>%����v=?)f�8P��gz\}(�Лрtө�>5�5�HL�RD�^��F��ѱK��E��s��~�}�:�Z�ik�r��W�w�	��4%e���,�����uf�!�j�b���UpF�s�Q�G��P� �x��Ƌ�8�i��RaH�	V����M�A7C߸>.�yo0yf
�`��ۆQwkg�y�M;���^i`B$�B~Ʌ�-�G#K_����Wz=�;���׸�c��.A��9��Q[��	.�Z�f�\�ܷ��o�S�Q�sU���`���Oi���,9)%g���q[���V�ilp#��[�J5��IXп�6���;w������|3\�_�P,�'����:D�^CUG�8)8ϲ�$��8��'Ǫ�E�m���]��Е�/�$.K��wK��f�3Q���1W��KFF��2Y���.n�WJnA���k���	s��P�g�m'J���4S���u�,�]fsp��9�wk Z��6s2ѵ�}��o����m�:�ߘ`|��j�Bު�9R��������Cbr�䡡���?$��PF��)��lLJ����$ך��5�>�)<O*�:�[o���F�O�
�ڰ���%E+��X{=T���46��f�������I�qQJ��vy�q2�R
Ϛ����}�Dl<���k����E+�fW�'��z��E����e�;`�M`��W���0c�,"�>�.7y�ȱq�5%�W�Ef1��"{vQ���	�\���4�;�K����4⇎
����]�\����R��m���=G�[ȋ��x^-�D�R�
�I��s0y1Q�J�I��mk*��>_*p�c�l)���ǈOF�LaЎY��q`p_�e_��9p5�&ז�z*Y��f�)�e�3K�NkV�b��.�~���w�/K:�)�0!g�C=~���T�n�o/��W���9m�����H��7������5zL$�u�'�>����^
ֶ�C<��~���:�t���#L �j�U�N�J� ��W��Mu���'�w��/���@�;�* �=x8 emӲ���f��\����������!�h��*z}'^5��+����r�e��پr�>��Ҳ+�w�N�P��UO5��W���2|�tf�(,��2�E,9�Y��_KoX��a;����Z��>��WUػ�h�?�d4\�Ӈ�~��6e��ŷ��f�SZW		=�'ԉy����s�T��(�Z�7�{���@��ؔ7B���p��ƞ��u>�X��q� �-��d@���<�!���Z%��\Z�6F���bv�َ2h4aa5�l�z������0p,+0E��X�)w���mY`�A�bJ$��4�M��kQ���#FR�zOڶ&���a�Y>Z�{�M3Nr
��9i���)G֏	��q���Z׀Ϲo߸��f�yE����Go�:,a�vЩ�%��C-�{1'����]��8�@[D<9bsN1N9WS��&���Dd��ѯ���g�W�I������BXk��G�/����y�V?73�N��q�e�����SG
�����I�pğ��3_���e�	f{�+�������Y��蛩���f?5�y!��)�b@30�o�cs�}`���Q�m��&"���-G��ض+eB̍�:Π=�j�G��1C�c3ᅸ��t@�c$����4�a_f��-�s�4��+�I��0U�M�͸dHo�����x�V������L���g5e�\x9��t�����c��b�����J)��'j4���e)75���b�X^�dZ2��à��-z��dׁG�o6�o�֓r���ͱ�4u۸V=���P=��L�N�T����l�݃F�I���g{Bu��q�x��2�.�E��<���F�§���E�}A%�Gr���ٷ]��{�%�����(I��$������q"d�iB��|0�^�H��IH����u��Vp�:��r�e��!�ddݳ�zU�9
� �J,�%Ӏ5�@�S���,U��w�� ]~z�m�k �I���AU[8c�q�6��@�N!���ђ�w�F$Y7�&�	��hd�fW��+�\t'-�YP�W8�"9LQ^z�q�Ε+�K�cr=�x�Z�x��԰��C�A�!tc�g;��)�}�g�2�'�v��=�OxO�1<�cĩ:�@��t/���=}d8_����Z�6����_L��a;��۝�ϰ�)��O�B�w�(������E�[�Ι�����ѣ�/o���'J	�	I�<�Q����Z���eƛ��7n���-҄�<����_۵���iu��"�ȁL�����4��S�D��뗍�|I�z1�e�'+�G�;M�#/�]<�tѦ�Lx߱�_=�(޵��WD�	����Ld���ҳ���s81M���`�P�\����>��߉��. ���2�JR����|	�����T�z�lL�4����r��׵P{���>�/�Ʌ����m���S���%�%̌�88/�4\9���m1�w��y�<�U�Un��*95YGe��˹w��L����L$ys���:���_� ,�e�	b
�Z2<����E��Pcփ�GX����|�4g�{CS�YLgQ|�Os���F�fh�`l1�|������)i����@%x}�g�g����=׋F�x��2|
�n}5�)�;��s�g��%��xr�ᴸS�Y�1)B�)��+K3�!�,�$��	�[]�x�_��A����PHGO?9��N�\I���
�	�F�f���D��TK;� �^�������+��	�St2#�,-�Y˧��Y��2��(k%7�)>,��A�(��G�u�b#��ʏn[��'�&A:��+���>��#�}-���V�w��A*J����6w�0���7��N[>����WW6R�Z��c���ܙ ����|�DM�{f��Kpg�s��6�ݏ�c���q���N�]��$p�/�lfNt��#��Nѱ��5ӻ`��5b�*ݑ��g/�q�������G�\�J���cǺG�%��s���+?�����΂��}��������'59ЖHG�EDM�������!}�#�[�N�L~��:�`if|ʹ����$V�4�#�úF� ��G�u�3% je���/!+U�Ots�����p��,i ��c<�Ӌ�25i�.ea�fE���kVQ�I�A2&W��ŗ4��y�&���Ĉ�\wN��ն*�M6���|B߭�~��-;2SK:%C�(&����6~��2h�cXwaA�9k'�[���.��A�^t'�b�o^y�Q�P��vL`�l�O���+0%b�o�`v�aK�V�ڍ�7.#��~[����[��к���16�;2�Wt�937���n��UD�������G��)Smb�� �8�W 'W������{�Wh��AH.f�G��� ���3�88�����F���8�:t|�/����Ac�'E�.�����ōg��ʎ�������n�gOw]����A�w�'D�|)�3|Z�Z��J"�J�xmE��kC|G
���[��T����ˎ���('�r\/p��#[?EI�O��Dܯl�m���I��Ռ5*���#O������ _��	$���.�GEƬ�XvNT^@���Tݡ���Z��g�FuJ5A�y�p��0b�U���^�D�@����K�[<e�a!G'L��z�+���5eB�Ӄ(�λ���OE�0�,}����y�q*�A�2��fl�z"��Q���dLT��2�V3��s��߇�6�哻�]���*'Rbv��e=�'�[�ˇ������{�� ��<$s�ِQ��5I{(k��>�p�����)����/r��a���>80p:c._O�߽��c5]�� *�f�wDJw�3&Qk���x���y ��2�K��X)8 �!�`�C�(5�M���*���z�jsVWc:_9�2��v��Hm>7�q�\u9���Ζ;>�����=��hCwh¥#��5���	��#�#��%������������Ī�w���/��-����;� ���s��mn�+��ۇ���ڏ� �Q+�q�z�C)Ve�U}�Ä��D�H2� �W����ѹ=4�5�S����̍��r,O�zD?&�ٙL|�ݴ���G��$E�tK�Tg�_����Y�/�I��̻�5��ZKUsb�hŹ�d�[�BТ�6����d�ˠ�7���Z�)��1'/n�߸�����~TN2�5�j����(J�����7����+�Fƹu��֓��2�X��-,��@���<�[�l��������&��v��U2�a0p���!��:�1�K)�,�[����~�dmB���mTь���b����G�MiJ�k,C��^���su@�5rǃ���a�|Y�K{�>(NU
��9d�yׄ->��7>q�~g/��jo�e��E�碀:�iv�}�%!D	C�s�{lIdݵ"g�X� ��'[�9}2�1���S� L&���<��I$�;)7gV�VIݠ��m�.XF��G�g��zt7鿱щ��NN�������S�M������D�Q��n�3W��	���+��}�(g�eog��d:���?�`!����0�_��%}�i��ė�2��&=P�ը`��\!E+��#�_&�8�+�i��d;��~Si� ��h֞�M��C��/��_�P�����;�Uۈ$i��k��U�*ͳY�o�;�¼�'�q�x���'�_��e@1�x4b�t�ˉ�P��<�(����>��'�j�-����7���;�G�sK�d����@b�A]�-��_-�G����/Z֮J��P�e��~���n=)b�P8��L_ڍ�/.���}�X�o�$�ކ�·B�xqߐvgX���W�`H�<]]Ǹ!,�������}��=�yr�v���r�]0��{��!�)��Q�(D}$�HI�qnWq=��i�I�W')^0#Y�}IC8�E쇟�ο�UO3�Br��ñB��N.AU�Q��s7EJ�.��@-�5ވS�L.�g=2��� Xa;�t��kۦYI�-A�CXc�i�6Ƥ��`�!�~y�, 3wi_�YR���'h?��W�ص�9t-��5ϲ�i"��x^��M5+��hc�'�����s�b���CMp�!�%�1	;���d���U�"��,O3	1W�P�$OA@�Vb/�:���Cc_��	B�RX6�Y���u�J�;��ڝ���������	�b'�Cg��g�� ���	�آc��ўH	o�'dw	d�ݜ̥d}�����ea�*�2��H{p�?�TW����ې�HQC�u-Yd�ÇĄQ�L�H�� �ɿD��r�ྷ��z̹��"��G,����x�qt|�|�'���="�/�/`W��ߪqY��ê.�鳓8�뮤UMF�`���\ ڃ��"��(��q�ͪ�m�R=�ၮ�0����b���-L4��ڕQ��Yi�D��;!/�e�.�8'amk���W���%g��83��4� ��d ��،y�Db�0�$n+��*�ضYB�v�&�߯�����z$�������i��6�e�g�e�Z�ʖ��E/�c�֙�����iw�nv�A{��\Yg2{Q��s��F��7A51�p��=8����i�x����xX�wg.�OŔ�=�Jq��P27tsn:�O��;�c�s�6������~�<~5S�N�1DΝ)o�K�I��Sڿ��	���\l_�Q�A0�ԋ<�P#�	?T-�u�Z�|�J�P
�>F����v����Kv��������+J��	)D�" #�,~����P�(�-O%��X7�J�YI�c}0(�L7��u^0N�ѕN������}�\]�ͦg���#��k�:W�rj�����`T�,j�v��ä�r-���N���W�,���\W�C� �D��MO����-NgP���DH��s����H�L#����p]�cp���l���۵�3�
=�9Ӗ��X�Qb����	�/���_���p\+HEسp����x%H:����?�&��EΝ��}Aw����{E5ԊnHB�D�٩�wʑ����L��)�
~F1:3�KiaU�(�U�ͫE�?�t4䰞h[�;���H��u;vH>j `ܦJ�_Ufy5s�Qn���r-(I �6C�0��AL�i��a>����V<�Q���A-`��n=��y�b��g���Vw�_�Q�)M1����B�ݠ~���-�<K��c���ӛ�1N��7Lc2�A H9�|�[g��.:{��D©���ko�QN��`�O߶��b>%]d1ǻ���V�#�#h0f[�f��$�е��̌�};�`.*	��h3��@�E�]>���@��GK��)n+:��T8��'=#ƅ{6��_՟j���/.�K�mī����3���g�#�AJo���O�p+�J6#�MY��.��MĚ&==����gs���㒅�*�� ���<�]�|���i�w!ON�7<�N拵ո��%.��8m�ʀ�^�|�\%����o������&�c*�r������?��4��w�_plB�H��U���5Ũ׭O�(d��M��"+�E�I��L�J8
Ea��Xq��T��ê�����L�ա�B�K����J��y��I/z�r���_�Dbe���4G����R��\'�"zs�ж���e�������V�ƒ0��,�r͛��`y�Vq�����f��;"�ͱQ�����k�b��q���� ��`����.�]��U�uԉRl����==xe[~+������z>��s��s�ZTQ[iI}�k��+>��r����)�pD�>0\��au(��p�_�DO�o��5	,�L�&*Ϩ�f��Ũ�3mk�f����tw��-�*K��`)SY!]�fC�4��Ҋ�	��!����W��9�v5��S�HH��7���5}pF^�+���΍>��>�T$��Z
C����g
�0g,�dp�#����Dw����H�T����ٿMXwT��/�5�H���1� ��w�FNm	Ƞ��"�*��Ju�A��삿��9�i�}]I̐�}*��_q��\����W�4|���Ǝ�������vO�������_�|yg/��y�K�gEb��O6=_�]�5����坌\����_�*�U)�h�Sd�����Ԫ�Q ��,���{�מ�m�Z�L����'�r]�sF��w�T�u��R���<��Y���7��m����ԅ�u4I �\�˓�0-Ǟ�@��o<9�V�'�����,'ƣv�v2�p2���a+6��0������fq<,!���c�������+�@mOb��W�b�_u��zM��k�2��#��B�p�]�M�Y�a#�aY4��{yO�N�GL
�\�9_�<��3f�	gq+����Ӏ�&=oU�͜�1E۪����:���vr�%���C���{����P���S?��L[���9�&1D�"S��&�k����������gI�jd����X!S�G���n	o�q����N+��[q uH�S��۵!t��?�UL�3�ߔ��	\�E+��s�cջ� �-��MǇU�:?���!͚��X�$0�˻�E}����
���#f��}3�&X�(�#�&�7��+�*/��1��3z)���Oe1陴��{��|���K�1���*	B_�Mw�����Ъ��'��0�U�Gͮn�oB��w���S2���a�8%�e�}Rx/Bwt;�V�p�&5���3���S�W��jj尙~��7붏����юXXdPs8�y >�|�-��ϥZ�Gi��y?��B�ˤ���C�.~�=���P3�WL�:M�ʚٙ����������ݟ(B��3qڜ���-Ǩ�$�{5<���A�Z�dI�}���\lr��̮,c]���{�7�d���Z(?s$A*Γ,{xqX�iq}�2>�^k"��ZI>������bf�p��h�
���X@?N��ҟUʉ���n�J�Q��[��5��=S��z��E� Sd����k�T#I��AKLDcm�G6��Dۚ!�Lۿ���w$��YmH���^ehbW.�����-�k��~"��$^�L����+~�c�P�Ů��nX_�f�AC�W!�K��=;�Z�7rʝN��+��v:O��1r�ğ�@� /$z�Cj�Z	�TC��ж6�/�z>q��;6AΝ�����)��R��^N���s�����D$$��ϟљ�~om��'�ސ	b&�G��XG�";de�Ju�-Y�5����.ru�z,x�kg��.u�+~������%����3��:�:�M���<zg����YGl<!��#��Bat��^��)�'�>=�Y��	��W��U�, ���(!��M+�n���0.M��m`�>\[@AˍTN������'/èƍ���R�\��� Xs���{IT��$WL��ȵ\ �5��.���X:/Y"��fv��Sf�m�9p�y�O`^%�8.��4�n��0���y�3��#nfhl*Q��Y=�������e蹑ՠp$o�Y�pu��K,��Va�e���LiZ��g���\E���c�I���Ԙ�*-r&��A{�IY��Qr'�sv��F,��A1ل�Ϙ˽�W��iO^�68�x3b�gi���/�=�)��.W2��nU����E;�׉s3&��[�]转��g�S[c�1_z�)�dK��a��o�Z�d	}%觷�v_Q�A7���P���?�#Q�A�ɼ!���
D?F�J����YK�����.��
�fo�+e	D��j3�#dL���ݲ�>��(%��u�7S��t�����(���du�q��6Ϗ$�/�I�w�|�!����g6#7�=��ro�m�2�=Ǆ���0Z��������!έi3����uWC�]�$�u>��5� � ��.M�v��/�g�������xťY�Y�'���8�]�apѩvlC�p�%1����q'����b%����D/D�b�n����\�e3؎=��0�c%�l��?<?:�=�i�θi�}����b��Z��5oeH=�DǺ�2���"b�� ߫�8~��#:�ˍi\N,��?���r�ZlF4� �y6 �v����u�"ы�j�c�e�U��"s����x��Ca ��^�.����i'�aa�oڃ��Vwo���A(���ɪ���]dy��i��v�l�Aw�	Y���M,��oV�BU-V~�-1gWK��̓�p��(0/�,>���&)c�3A4R9a�"[B��.u;-�7���|*��o�$�Qk�ח`g�O����p�%X����%��V�ʏ�.n#C��[Lm�����аB���|;�� I� �3�͡{����F���.�o�wG��)�	:��CP8j�O'x0�����Fk���M�`E�.�;�谂��yb3���<����D����e��Ȑ��U=ވ����Vɻgg�
#@���1��z�u�Q��Iu]71��Ǳ�w|�x��n`ipe�P��� ����,m{9A��q=|����s�!ɊQ����f�Z���Mr�$����?5`������z|l���ϖ�K�U5`�����O;�8��!,�=v���F{�k�m�qaE�M	XlT�e�'��ꯙP���T��ݿJk��y����MR��[ֱ��Dݩ`��m��%����WM'liz.�k���e8����|Y�Sr��h�0��,3甛_�y�M{q e�贅f�Z"L�3Q�,��k��(K���)�9��5k�?���Ɋ]�=K�О,R؁����<=��[Y��)p��!��L5Z�sa�{Q)�I��ak��>]��4"�)�qnǙP�w��a!��4%�p��o_��R�
:75�Xק!�*�_ff�s)@�<3��ek^ͮ��oo܈�GKk�,)n�U!�yJC�`F|T�%(��5%� �UWٳB9���l;CH#̡7SY��S/Uks5���]D&�>�`��VGgܻC��q�O�#�+_r��g�#}hG�#�����y8��PQ��rٺ�w��3/C��c�v���" ^eo�Am���ְ�mwx�n\�Q��g������Gi}�����^���0���0���ѯ���c����q
��O�֚.OF���#:�F�|����R�熯^E�K��J%�_\z����d�����Q������)�U�%h��dE�Ӹ���l�����5�V�g�x9Z(�_��k8'���.����TD ���+ �,��^�ʕ�hY7S- ������.u�֓7�#�� �-bƋ@���<�0��Ko��s⁧Gk�Q�Mvm��29��a&���L���7>���~,�/�>��ڹ��Ơ_mJ�R(�b{;��bM_��k�.^��d^#��k�H�o�a>�nY���{T�"N˓G
R019ZC<�:ZN�:�SqFM��À�7o�^��7�Eּ��X�:]w�v!��%S*C�a�{����U�N|�I��[N��9��1���S_D�&1��r"4�y���W�g̯�IU��c X�/bGN8����j���gV�G,�NF؋����P��S�3���^��:?�İI�3��u0F�	�e�+r����c躛����VP����?f�!�E����0g��ߢ}1m��mЗ~�W�8�#&s\�՞��r+�]B�.c�b�ڮN�5���E�������P��%s<_w�TL��x��K���q���vU���ͩ��o��$�2a����խnp����<W�ev�x*B�t��C�+��Aw��1ۯ�⮒�j��yf�7F�G�c~ѩ��d�C*�T�iϷ�-Ks�U9G���4���Z��F����tS�id�=_�P.R+L����&	�֢��NW���*��]BF�q����)�c̕���<S����͉�����oD}	��2r>�ڮ)%]&��{�Ê���PI(:�?$�+3��}qsP�i����u^��7�I92���$��k���H�G/�bg{\�݄��U���)ƙJP���vA�5y�SnF���m�H�� N���*�kQ"1I�A�t�cH�6<�p��u�!�:��:�w��KY��C�zҏh�D�Wi쎵-%�-�$��ha"j�T^˧����+Y�7c#�d�I�q�i�w���jC�-�!őP$�;�Q�ڋ��8*C�z���h�O���1���;@���/_�R�ް7U&h������;�6(�m���LH2;q���R�䰍xR�`��=b��yU��]^���3�������є��o�F+'{y�	�T����3,�]�e��w�(���ҵM�R�����F��9ucp���H��^�W�6�Iɵ���(޴�-�%zUҩ�G�l��T_s��Xtr�L��e��b*=X"�ǹWUSl�������;�����I:Y�$ݺM|-�`��j\�ƾ�H�|�����8Ã͖�[BRs����r	�r��6&*�˘�L*��ȐC߷p��!8΍��/��;�!ސ�nţm|�T��Ê-J%��	8)�4m����f��L�y}?����Rn�@�*�w�Y8~���o� f����.$�ޠK]������eԃu��Zc�i���E%��cg�@������m��,��{t��Y�(yQ��sQ�dFg��mb1Ը���~����iE����9xKog��=��~=�({߉�Y2��lnp��E��;�k:sn5������v���p�S��1zF)eo�K�j5	���Rx	x�g���_�9AR~�ԁQ�P٤�?�H���<��� au
���F���l����=K�6�/fs�5����R+�:�	_>�cJ#?��
������#�9+�7����YTO(�1�`6u�+����K��D�X5��K͜~����)#r��p럘hbr��ҵr.U�K���lT��$O�������rWhy� t�Ӯm�9�� ���-�&M����Qg8b��A~�.�=��*��1%���]��4p̖�lw���+�@������Lid�Λ�b�8���Y�/�7��)�S� �=\!���i*y�k��%~9}���^?�˰�$G���N}2N�= �ӕ��5
`�H8jGD^�+��h��=2��������~�6�:i1�iWg�����C$�u' 4��T$5�����~Yu�D,�Zj�ݍ���@U\,<s�cK�3-�c� �t�M-|����iB�La4$�zVuV�.�(�A#4��$d̗eB�y�:u	��G�w�ӑՇ�UM'JP��:�B�~5b�-��+K˒+��E��ìZ�'N��C6&c��AO��9܇k[/V.���Ҵ�Wg�s�o���Q7����o`B�]OUm����U%S�H�qF��2V��lZ�#F�[�ch�,��Ы���B��;cxrd0K���3�����o���j���p�G��k)�b�x8E�o'�N��=���M=� �`��J.����c���x�3=����7��I�E�5�x�C��{����4��\��ɶ�g)G�����"� VP��w]�����w���ʭ�����s��ۘ'�Umyp�ˤT|Xa��.��ɥ����5a��ِ�r-�롢�J?�,�<)�ٕ��l8���b�G׆%5��Q���O�ٍ�G�X�׍;��Fhe���LE��_Xg�.To�� qC��@;�˴ݻ����A�J��y�-����φev�¼DX*�}�b����,�#�R?�']՛z��5�Se�9������$ *<0w�,�{\���yeyq�_����ef��"�NQ����u*���Қ���n���*��z��d"�]����+�R��Վ̓=3y�[4K��d_��#�����?s�QD�Is��k�p>KF�Ϗ�)�������2	�a<���K�p���_ �꽥�5����S*E6�f"��k�3��xkB���IS��j�u��%K&[�)�k�!S6zCq�:�Ce�������{W�W���9�^X��B9H��X7�+V��H�f����x��>>��	�J�B~}C(�g��Pո&wT��#8k�}��:��T��8���s�ٵ�w
�/�0y~��'� 9]�$�m?]��^����^���������ԱPF�}��C��O��Ypp�Q�c�*�]�*YO�>*��{���Ա��YO�dpRF�*L�|oڨ�{K����	E��˽E4�_�hc�������M��e�o���IUD�h��d�B�s>g���ة"#*�13�R��Z�/���'@�A�霷���$T�����%c�g��ӕ��}7����\;��
�9u*X�E��	A�-�	@���<���1����"�ܣ,8�v�F�2�>a!"P��޷k�ڙ�a�,��������a�vmE��b67מA�M�mBk���Ǝ�3�f��Fdj����aY[�Y* j{/�'N �
�#�9U�wו����qaW wL �t� o����:JE����t�:v<��%�
�Cp{pC݆+�Id�e�[	#�9�/1:�S:�h&lfP�WT�AįL�g�b�I._���M�X�,\G��ƥK�*e����Hj Na�$�Q��+x�S3׆�Wi��5��g�3KQ�K&�	RI�+M�����6p���Շ&?!A.!p�N:G0B�%O��}�M<� a ��,���� &�2�mY��+Q�b�0�.�)�؜z ��0��ּ�q
�hM�O�g� ��_�L|�@@��Ʃ�����)UU�ͤ��o��A���M��!��b
˸k�w<(ew�x%b�t��P��O�\ٺ��^Pۊ�ծ͗fj��0�tQ,7�+@�l�����dF4��/�����-�x�P��G�o��15���҅��	���ۤjq=�jP)��Lp[L�@Ҽ�������3��B)�S�&B��q�xZ������<�q���΁�Э�@}�|N)�r�[��D�.]���{fo��ڵ��(5�h$�Lx���fq�4�i ����m^�Q�*�}I4��Vq����Ɓ�\^�ߐ=i�����|%U�Y��=tJ�І���5�v�SI��\��$m I����6�k�I3�nAA��c#6w>)�z0H!�H3�=&w�i!Y�H���e�h�GjW�J���J+-�����Y("%�^�"y�\+4Cwc^���T�d����3C~��!����M);f�� 7��%�鷗,�>Od�O1�n�ĕL�@k/�Xq�y&P`#�
	�F� 6C�p�z'�W;�5���1��}9��Q`��O��|���hu�/��.��4)�яX>o#�'640	�f��=F�1��[�e2z2�#�Y
��p^��O��pM��!�t�Cu�0:��YU�b���y(��Q���0�8�9Ǿhb�z���/�G"��������Xt��F�kߝ�m=�
���W��"���Q��~�x04�$�C�_��M��`�\m��o��ۡ����^^ܖ3=R�ځ�)D���"��,�L����kJ����<�aZ����/�x��em��Dm���/[���J%88$�4��������iy��ڛ�7�n�8�*�w�Y3q �7C���ۑ+�$e�/�&e��+�e�A4v'6ZЖ&�E��cB�<�3��`��h�H�{/b�Y�SQh$�s,]gF�(� 1��NR����i8[��,ˢx�S�g��B�e�'=�GZ���2hq�n��t���;]�s�dYՑ���`��M��S��d1�2�)��LK�fbpC�ڐ�	soc�m	[_ǐ�AmUB��bP���?�՝F���j�[�7
��F�������K'm��ʽ���9��`+{0Z	z�)30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�%ڜ4�z^��2�Z�n�;:�|͚�<���͟E9F�_6���(�(F��Z$����8#lfuP��Դ�I��O����Ŭ[:v�,�82�B'�l�(�,YB��F�2�%xd4��o����C�ƶ=wS�%һL>[q
�\�������� �1}?M6�h0&�	 Ic[:������  Ll|�A5E�Rv�/�h��]��
���Y�������le5H>�Q�핥�'��Li��?��?�.';.���Hs�o����=L#����ިa0׊���[�1죪Q�)�0����m���獖l]v�%���6騌 .�~
�J~ :��J�?ą�@vW1}[I���Y�G���w�qT2n���_Hw�V��Ԥ�M�z��ް؛��eB���b]�=�o�f*�.�_��e�b�Lo��n�|uwAB��R�k*�H�3��<�ێ ��X=۔�,�͠����
Z�#9Q�`N�\�&�K+Ď
�Â�P����0�&Z&
�
�4qg��^��H=Cb�&��Ӈ�JV�WK�Mۥkek'�x��s�a�t���&J��r�8/�sW|%g�B�!!u�is2F���in�^�����M��y�����`��s��DP2q,-������t�M$~����/�Qy�'���������)?��\�o᳋��4��8UiqQ'��,U(yVY���X2>�S����4��[g��2y���s��a��u�yM'�F�mr�TR�RUq��:�j�xfˎ��csb�Ѡ�˿ȷ�9/mۃ�>`�-�!��U+��N������{ <�z}�ْ��B)�#4�o���z�������XpՃB��)�`T1'�&�����M�������f�Y�� �lBi�2f*�4��?�A���.$l�8�L�'WΓ!i���xh;��=��IgC�&D���j�ۢ�Z2�'R*Pa�J�m!�CE����J�e�nT~q���Z^��PO)ju<���&�cAiwU�̊ڋDA4�����[����-�oc��w�x�Ş�t��"��
�[ȟ�U%���//�1rI��ӈ܌�ѨNM����q���t���u���^�Ϧ��!�ч����ꣃ�"^���]�Ȭ���^�e�CS{�p
�kc����Y7K�v��0O�����M�y�)�q�<~���ȷ�J@�u�����/O�Ĉ=�|J�UWuM�V���_���U�p�{wuw�$��Z���!l~46�.!_��dH�d�����,X9����a�l���D��V�ݜ���sR'�ʪ9͛/~wr��O����l��K��w>��sj��D��E�? @K	�&;�Șl�e,�$��>��.�~. ��)E��\��q�fezc��[�;f�y)Y���v�l��j�����LH�%�z�OZ�M���e��+}�h�]V��W �r�V���(ZX�nO��rb**�ԏ��y�Pf��Eu�.�<�w/A�����٢�sr$X�&��{@��|274.�����@�K�_��'��T�)�L${)Y� \���7m^���U�!��1�a�}ĭ1?�M�y���VRv��HU糓Ս'�n&��/��w�����G�TZ��k��B<��k]7B�/< f4�d��#��qK	���z�<�3��	��IfЭ�S�Z������	�X�N���ۑFZ3���ٹ��QŖ.�{k����G�J��޳���q㪗�h
�5�Q��\���?���)�l��I�,@�"E�J�v+�c@��Wx�_�{�����I�0��&9J߄�N\����0Ҥlu���ŗu�+�����u(���q��2o�n�IF��6kV8��u_"_�vq=�w��`C!�7¯��K��L/<K�19��t��mq/us�XV��pMK��&�(8���cI\ث�%M7f�M)X́~}ZG�J�I)_o��j1�&g%�u�Y�$��e����#��5y�Q�����w��ĵ��c���@- ���Hf�'Q���η����c�90�����J�����}��/f�K�B������ �<*��I�\�^�Օ8f��vKUHxZj����=�aؖ���� 8�e6�B�Ġvg��p,�h�����K�a�RO�Ա������ֹ���k�R�B _���^\�g#]��r^ �W~D,[f��&]t;�ӕ�uZg8��lH�`��1?�N<�Ai��t��t����x��$m���7/y��A�����N��MX����Fy����ΈS볥!N�|���](�����;���mŏC,�\+�9m6[B(�mMC��̋�!{��x�c��l��5������2��pa��ĵPA˳���X�Xf�p��3�]�J'���mq�������!51�`?,-�fڨj��������nownM�9�6h��Q��÷�U��{oE��������r�6�|�fu�H�H�g�->�\�1�.#���$�<� ꞔ���]�������^�ߌ"2Ot��	t�k�ˇ=A]�e�"�u/iY.�ZO7���75ꏞO������3�9Dʂ�e�847���<%��(��ȟ'�A��8�Dlw������P'������C�����ՖVX�i�Bnbo��hu�h'���B������mT�~�W��p-������U�pk�=�����5�����F���D�Њ�Ӭ�!�R;|73�`/ŧ�F��Z�p�m��W��W{? .C7R K�x~�d�s]�Ł������w��$釤�j}���0p΃y���:�uT�C�Q���>�(Pr�a�gR��y�q���K~�ʭi�S�ūT��,�'��6Pp�&7��m`;��THS�\~�PVB��FSd"�1-��Fn��"`9b��h����Q�	�>J ���-%E{��F���F+�M�	I(�L������
��P�Ck��**Z5ʧ���UY_�˘������K������~��L�c��>\�nJ
P�z�Y��6�&�q���.2�W~�Kw���nv�SGuO��D����R%.i�,��t5�@AS�9�������քD��8L��T0�ZNaH�_�"�u�و�� Zh�g�M]f"�|o����ڸ�"RKꇙ,4&�t�R�{|�Ν�ϭoGB�t8����7 a��I��Y
(�|B!@!��<����f�u`7̘I��ݎ�ԎM�/�V٘#e*�$���։����6��6\��X0گH�g#vs�=��uNY4�W��$n]>��0���U����7��!��3����k)���o
��r�]�&���f���{6�X�b;�5���52�k?;E���'�d)
� �z�>�)V(�h�����r8W�i�i����v6U]Uk�}>��ֱ�����Ϯ�\�NS����~ʌ��">e�#�cJP]o��r��/�9熶��ڲܔݹV��[ e
t֦9R�����}~�*�tS��7��d	��^>e=�5*�w�7�96��?���G,��X,kWz�!ʱ���`L�]Sm�u�?*��Du#�y����%�D��L2�L���-��G�佩9������.�^����fj������j� _׋����E�ע� 9Ec�;I����x�=�E�!,�(&�_c�<,� �*�%��ĒZ`'�@�Z�h�;�|�z�C�����%#ў?\k�n
�(&�VZ�X��NklFG�zz����կU��Â�;8��f\8�^���B����Y"j�F���%XB���{o|���#jvƖ<Sˤ�қn[Q�\_s�dV��] c��?-�h�P	 �j[F��hfu��Y�l\ji5%�lv��h��S�f�����Yy����Iã��45(���13�Ϳ�ԍ%�n��t�c��'�S��-�s��E���=,iO�hraa�J�����I�1���y��ǔ����v��v��l��L�^�.��.�*H�:�!�*��e�xv7�[)�J���f�'��W�q4��ە�HW����Ԅg��Z~�ސ��������E�b=��Ox�*��C���EFb�k�o��n�"�w!��2��*����U|<���n�愅���P�wF�|p�Ƀ�*c��Q��=���g>%)[h��8������?���Q^<��+%�#������5+t��,����z�����]�m+��m�8F���dm+wE����}ǒI<�� ��F�8e��]��V,�)�����$OsK<���6%�k���L���"K�`a�����{a��V�rC�v?��nu���/p�.Ӂ1g_�p� D�\]�z�er쾗ꑟ�5~�]YdF��ŧ�񁹣���uX�9?-
��J�-{���=�F.m�+�o1X��%wlN�6��A�t�����b���%�m�D����tJ����2�ݶ�Ln�^��;~�mм�2�+?cVh>1��G����Ҧ���_TI:<�I�#��TԠuAG���L�����s�&!*���P�?T��_�S�P�.�5�q`��3:~�!Y4�f������rmO�V�� ŮQ����A �8��߶�7�Q �q���m��Mn��n՚�ح����-x;��У�r��b��C��(�=�r��ǧʈm��v��um�0y/b�Jǜ��t�f�&c�#ؚ�}9��R��G~ct@��v�g�!J;lb��j�axAN�4+-P��u�w��)�~���R�/[L��y�c��vd�1^��O���D(F֦Gqs�p��f_EcA��p����$t�.2=�%N~z4p�:��T�LC��a	"\�p���l�=���y��rJ�F�(�����8��/U+z�V��{��$��E*����,��i��ۨD����a��Z�$e$t���ؕ��m~������R�6��×J�B�q��ֲ�~��c��y���|��Y��L�qy�y��2*�P��Hե(��4������2��B���� j���3T2D����Хhj��w�-v~�j�՘ {�2��c�}e�D�;H�z�Ō�K�F�5V݄�y��T�UU\�Y2I`s�|� 1`��=�\od�7��G�Y-�G_�+�n����3s�W4�c_�[Rw���Y��|_6��@4�7��>3�BE���0\jD��+˱xNH�@��e]@�erj1��.��*�{]��&[����ߠ���"�*�Zh�礚Zm���1��K��<��ޮ���N� �.�19h�(x՗����F��-&�X�������e��~N3�3�N�����j�͓XH?-ɛ\�Ĝ��lN?�03,�?`&�@���j�I���e�) �W����S�u�6��Q,͉�:���l�];w��}�uS�*:�IwGȨ&F7�qO[�zЧK��7hg�gG6���{\�k�}�@bO���T�i����[��>K)�=��DR�\�j������)�����Xs})tUWn�`:��LzXW�Y�0���v���E�ۈ��x�S����/�W��Y0U7������c9d9n�`5&�t�HE���j^A�K�������>��_&�����l��8�j�{ϖ��|������@�;C���!����	� �H&�ʑ*<�R_��ba�i���V�h�58Z)z�*�����9��4rc5�~�G6�k%1lO2^V�O�F0E�O���x�w��'kX�K�h�½��|�`�E�N�6U*x s��24�
��Si��E��(ֳ��E��C
ʙ�g�h����v����
�A[�7 ��Vڃd�,0��M�;S�$��qB2���N��TW��1J,:�т
1�8���|���9D�X����1y>q�����UJ�g�Ӹ��Ե�g���k�<ݘ��J��' �1N��Pqm�yGX��!%���(���;�x�௎����r��ѿ��:�����{�Zr�����
~�؇�:����:-�B��c�L'J�v~ ��s�dB�����%���7��aU% "�,��@�9���&��:��O�Fač#�S��3$4���;bU�<�^�,�����c �I��ZHIڧ�T��;G�u�����L![���V+�0H��zm�"��d�79f���hЖ�_:yi��ڎD������d�@��pA���4�"�����S�8�^V!#�]ھ���AY���@�P(�N�:�8��[t6�+&�m��V��3���i��}���X��E��{��k�V@]�;Nb�hq�g��װл�QɒL�c
(�!O��|����}�8Q�M��������BN���|Zp
L�Q�6�}ƃFB�YO��N-�LWw��?��
T��o��0B���Zdd��ŅM�Wp�\�ݩ�]���1@t��(Y�d`�k	p������� ��Ga"�1B�vh�4����1/���He���9�>Fl�n4�ﮖ�Ȓ`��H{~��B�]�P%bCE����&��F�AP=��P���2	gr�mgSp~]��8��I��B��l��S/?@�v-r��׀�����#N�g�M�=����@g��[��0^ZP����1qZsʟ����q��N^ސ�=��&S����P��wޚ�kkRҤ��s�7)t��X&����5c8��W���/��!B"s_���P�M���Ä� �M6\���?�M�٥ zq��q���bH޻���M�\��S��e�'yӨ��J�:?�?��u�� ��4m_nU��B'�_�,"�'y��丘��(��-��4�\�����_�F�����ξv��V�aF=}�Ag�R�#)�g�#�E�pnso�4����Sp������۰n�`ϡ-��b��k�TH�����h�z��:�_B� }#Ap%�~��zX<Շ��B��z�&����BBVɧ!p�T����b�?����r����S�X����$ 	��ih��*X���ve�AMq�.Q��ݿq���W�u�i_�>�O;�aT�.jVCA��DL�<���ۯ���8'N��PN8��~CCr��Ƚౕ��T�ͭ1�=^7��P<&{u�J��SʧA6��96ʋQZ�p�"�k�ږ��F��@�x����	�9��!?[-����%_<�\�����I:�~����UCG��
8^�d�!I�����uk�p^�b��q��4�� {�pa�"�cǫ����U�^1�iC`��pĺ����V�
Y�S����0߰��蒼#�e�֧�Ɖ����g��U��Jm�C�|�7M�����)��J]�Wb�BV_��C��2��~w��6$-R��7l�lk8���C_F��d8N�a��9Y�9��>���l���f���s�i|`��/F'܈9z�~����P���D�r�����Z��������$ -|��IE�٘�<e� �$,�T���.L�� �.\ERiڲ���3�zЙJ[�0��&���"��Y�R����*� Hf�BzHt��ZZS�̄+�"��J����H�ǟ�_̛ARq�`X��顀��bw�|�|:yCuf���E�9�.���[,�/C��&Ds_���^{mN|�x�.`nZ@�Vn_����ľd)8�{V�� )��ͤ���uUq���~��jŭ��`��CyY2��K�"]�U�xk"��'��&L?./O̰t�^�#�[G�t��g/ߓ��:<�0o]Ġ]/i0=4��ہ4�*N-	�9��a�\<�"�>�\�vs�����ǳh����	U4�N�#�~�LZ��Z����ŁƖ�1�{� ��*�ǗR:���Z�,����^|hז 5 ���p��f��� ��Y�1��c�Y����n�J's�+�4+�qJ����^������]!E��Jo_R�[��\-2�>v�Yd0�pLE��Q���\�gh�(�I"qk�A2�3�["�I�ʭ6�K-�L���_%�`qꎢ�;��CL�<�DK��L�YP���ぁa�W/¯�XCδ���VK��`���t�X�\�-�%��f3��X��}�ح�2/I�v���{m�3X%%�����n��e�D����I��厲*���r�b2�c!S���h-���K�UϺQ;��p#و�g��`fs�]��S�)�C}�n8fnm�x����,�ë��*)�g���2����fMuKbLx�Ɨ\��*f�ae���*�8��g�xĭf��bNε#���壏�R|���l�l>����f}�|�URg_�ox^�6�gP:Y�?�V����,��s'�t(<��geXl�ѹ+��[cKA����Tt�L��+����q�iN�/�x7Ae R�j�}ҝ����s�b���������|�d?��f �(�3�ɩ ��������m2��,溼��=*6�Wz(���MЙ�5��SЂ��c�������
�Ǿ�L��:T����P<��4e�$0�[P36���7 ���&��}"�˘j!�؃`L�t��jk�M��+�0�n�<M��K6�\��^Tj�JW��{\x�QXB�̈c�?��6I^�s��H29g�3��Iּ1^�_�=���C��m�����]�B4�
�Đwˎ�l�`"_�9������X˔�q]G�"6v�/Vce.���7R�L�����{O�������h6D�)@e��M7��0<��E����Ȭ*:��U҅�DY��鄃��}��>؞�8�������fV��1�#5b�mO�E�5U��s:��1��o�m��������/��>pϽ�=����5���;Ug�����U����]{ǖz�,�Q� ���R�%���B�d���ʬ*:��b�j����7&�|O�0��y��:CI���QM9>S@!!��)ygc��y������K�=��>�6SS��T�%��P��G�����7*>M`�)��8S��{�!�ꥸ�d3�=-�h�n#�@`�|���n��tdQ��h�/5Z�	8�-V���j�XBs��aQ��S��Ժ����́��k!\Y�[5�4��Av��6YP�ט�?�/���M��e�������D��Yn;nϋ|9���&���l�2[ė��uf�v�=ngXSX�~��3��9�ä?i�<�%U�@�V^DY��+VP��A1���aȩ�����Z��p�P��"��'��$�CL�Z�1Mg@��f�Kao[�`�P�"C�{����4W^�ӣ�s|Y�ɝk@o���t	����� r�fI�
yރ|�$+!&�FCQ�m���f��7$�tI��3�Po��[��KA#�@$�.g�z}x�؉��K�W/)�0Kuѓ{�#'e��g�u?o04�+��U�>��0�QUBB~��!g���k:#n��^�Òϗ����,^�X��Ԋ��������;�V=�O����ױ	����)Ga�h�^��W'rS������:q�v羄U<p�>���,���ٗ����������	U�s��>�_�#ɼ�PI|�o���B;v9x F���1��Zݪ�w�l��e;�5��������Q*BAW��=���!3����enp�*>�7_i�6�i�?n�0��Q�IJ�W��R(}���LHom4�X?ۯ�DF�j7��"�T�C�ڝLr���-���޽z_�u��s�__�^E���L��jP�X�eA��uv��p�)�|������1� ������`�yY�x��HE��+�͐E1�Tb H]�%Kcܒ�.��(�Z�k�;+<�ͫ8G�(�&��6��~��0(��PZ�4���0�lwkCˮ&�g���@�0�tWw��Z��*u8#_���irBX�Ǵya�Y��WFz�%)�
��>o�g"�TК��7�S<[Z�,�[�d\0`U�X���l ���?~�:h�'k	�t�[�}�9�Z��AslmPQ5V�Qv�k�hc�� h�Df2YJ��Вk��I�5Y�����2>MefA���EM��m�',l��ss�K�՟=��~�,C�aܠ��02�BiN���#�5��Ql�k���G��vtkS��6�鹊.�>���D�:y����a��6��v(��[:���էxX��ȍ]qţÌ�7H(b"��4ԕSD������J�6�����b�:�� m=*t7�܂�vU,bMa�oU�ani�w�����*���$C<�Zۿd*��"M����w�*a|��~�t�!t�Q0�L��؟M)�������iX���;?���Q�.��|]�#k3i�5u+%B�,����k�b��:��"�f�8�i��i�H+�:�����}�<.�m1�F4AF8��9]�n��)gO���s\���ʇ���ܞ���N���P�`2�Ғ�EW��U8��-	CⲤ�e5?@���s����1X�~pĕӹ�tz'c��/?K�0��~���]Ԗ�F��������[b�n3����2
b����	���NF�Q+�X��w��٠�Z�A~W�_dU���S���6mF�߮�>ߠ��Ŝ�=2����o��
y@�L�WmX�22��?ԁB>GE�����&�_eC�m�L�tx]TE��uҲ@G:��L�h˙���؄iH![�+�(�T��\����߲#�B���q��	9!���f�`4�Y��r�������$ �B9P���O�i���:?d����p����ȸM_����]�)t8epr-	ڸ��A��CGXb�U7C�r*�n?��L�$�;�{�q�&�i0�@�b��%ǭ��t�h�wU���*x�څ��l�|P�o��@�(��e�J�u޼.��a	��N�C-!���-w�������Σ�[y`[�
D=c��d��A�ɤ��a6(w��G��UpF���tc���AT��Dt�2:=��V~ˀ4pT�����a�.��a0q�}��=L@�צ~��~�x�*�]��)�/f1�܇��{���$TMHE�TZ=c��'�i�J@�Us��E����$֝�ɝ�����~�oZ�~��g�/�i�D\�6�Ay��gB��˪����#f~�Vcp�����j.ؽ��y[#��HP`A�1+��>�&C���vسb�1k�j����ť25�4�ҥ��>jѪwZ+�vkm9�� L�2�:��quD�����՘��������������E�Of�Yc<j�%���R*1�mD���-���(��G(�YJ�ޞ�5�+"�s��3$y�4����L�*��{����~�@�u,�/��3E�_���T�!.�D�Ư��~N`�_@�#e��[�5�1W��x]�{ni�WU�;6��$�޳z��j�;h�AÚ�V�&-�bؔK���"3dě���?��$19Y�x�*��ʂ��(�t]m�i�E�e\�N$� ��b%��+�� ��w>���^�B���AN0l�3=O�`?]����1�It� �f �� ����i.uA�ѶR���Խ��p:�3P�=��,�2�R�u��:��G92�F�M*O-J�x+���g/��xP��3^\2��}`�]O��HT��T�����ע)����s[\l]��g�������^�i��)���nMC��V�;z�,g��*v�����_'�������Y�(��X5�[=8U(��=�����ur�T5��������jO �Kg#�!»�`c,���~�L�ӷ48�ij�"�ϧ֓|�����ı�W��Z���ż�_t	Ё�H7��[�tR������iO��V��5	B�k���3@�� r�O��c�mH����k0� l [HG6.\^0J�O��fx��M�[k	���9F��3\|��XE�>��?'x��:����
��LiZ|a��-g�GUE/�)
EV��A����j�e���2�7�D����ƃ�o,���M�}��$sD�q3�����8�[�:_�,����о���^��곆�a�i�����>®a�e�]J�.��i%�Ԇ/2�z��k�������P�W��(��8N�*�@X��R%�n�98���e���x�� 	&@��r���ѐ��:�>��	��[grE.KOw~��Ї�6��e	:�a�荋LXq���p�� �k����"W�y�3�uH��a�2�"5���]�9Hyq&��fv���q'BO�r�a�;����3�2���Yn;�<]��v�ޖ� ����H��]��M;����F;�zdL2�Z�ՁV|��H ��i%�-.1�R��ŔV8]����.��G���:�8Q��rN��'%v���[`I��Ǜ����.3-q����r*�H��C�ԻH��q��އ��МY�9�nb�W��&�*�%>۝\unb�}5o�b�n���w������*�яJ��<�s�eǽ�\�L�ς�w�S,|�,����Z�T-Q��-x�>]�)b���?�{���5�c?Ԏ�Qu�"L#��Ƣ[�+wf,S�=�������:��8�2�ُ�+��0�,H}<TKg�&Fڻ
8<��]��;��Q|)d|���s����-�-H/�Bt���"߹S`�k���]���z��m��C��e���,�]���9䥹n1�p��s�jzͯ�� m�V�	~��]zƯF�~��^��1]�����:
�e��<��92�F��*+1^�X�JswcuR�HwA��h�E����幽x�\Im,����]a�K������2w�ő�p��p���r��m�f2�7?:{�>�eG+���v\R�hb�_��S�u�#�T���u���G ��L,���7ت��!A4��G�T]���
B,�ũz��E�<���^2!p��fw��󿬐r$��cu��>*�������F�O8�߭e�ީ(Ĩ�V��9(}M�U���hձc[�6�ˇ-/�K�pʍ���bd�0C�O�T�]����Ȧ<�@�30�,�bD4n��-t�z��ۼ�M&�4j���'1�"�N���@�[��~��J2
"��ǎa/`Nw#)-�f��ew�ۉ��v�I`M[ߏ��0`'c���dVz#<<��� ~(]_Gh�p�2��2c�����W�@{Dt��I=��V~q�9p�L��A�ڈ2a�x��Ǯ�����=2�}S;y�k�^^��|qʏs�/�BS�m��{��.$���E��#����i�٨{J��+����"�$<�Y�ï����K�v;~_��U���*�S6����n�}B�ڲːV�̌�w~?��c2���_��/��#H y��1��P�P��,�3�h#��f�A�w��W�Uj���Ɇ��2�J����Ϊjw��w��bv5}*JP ��a2K��v�vcZZ��p�����8`],˒"���/{k<.G�?7h��Q��i4O�����}���%D܆�eG�7M�<�eԉ:K'��f�-�
U�D~m��Iz����ص��k�Uu���|���3V*���*(bSY������:F�������w��T�t�P�}��J�G� �S�Kp���=�����LŦ4�b&���i >�%�]��tL�RM_3ڇG�9�c�u�ۗ���;�=���   �R�����d}������S��#*��������.�Q�0�Y�yC�5:���UG�Q�E>4��"R����g��fyJ�g��_[K�y����S4��T����t��n!f7��7`Mvܜ�Su���"��م�dt^-<��n���`Kڙ�����f�CQ�_1�P{3�JB�-�?����������^ˈ�?��]#���lk��y+��5p�F�-G�<%Yq���xgᐞ,�������B'Ŧ�50�ɬn\�̙��J�&�F���2���-�w��n��S��Q��I�u���dW�i�^�4^@�et��lթ�A���V.�JpI��oZ��0�Q��"�R�+&���Z:v[g�c�ft�o<i?��4"d���ù4�g��$3;|��w�,�woٖ�t
�i���i ��IN�@
�e|T1!��L'f��n�և(7e�2I%���ц_�:��G#�b $�֛m�~j�g��10�?�T�9#*����u`�4�����>y��0��eU�����!ht���'ek{y� ��D})�8Lθ�~��)X��j�/���#����%;2O�9�Y_�ג����Po)h�h���{ar�c��{UD��a�v��yU=�(>#c�m$F�:)6����n�/�(���c1�t0f>�W#
�FP���oZ�Y��`99S��y1���t�˙Ҝ���e����ǘ����|�*#=E��b�����;6�e�t*�k�7 
6m�?OI��s�jSW����£y��L�m��?�M�DGbh���:�c�
�;���LE�D������{*æ.������f^�:��Aj���y�^���;�\݋j;���n�t�� K{e��A�Z��x��E�������^��@ �R%b���i��FZ�I9;l�j�#��.�7=ў��n� �(�m�Z��䃈l�&_Lֹ�����+�U�Ӭ�G�+8dc��&�?B�G��UYt*�F[��%*_t�j�o����-[�hA�Sݔ���[���\1B�v���:Kt ���?�˴h"r$	R�[��H�:�_���"l�g�5���v�Wh��������%.�YK����(�L5����+߅a&"�F�	�1Be'm��m��s���S�=~#_
D��a"B|��Zz�ۛ����@�سQ�LUN�Hӎv�b?�&4���.{��<�W::@�üm��7��vI@�[{�:�B�U���~�i>4q�h��m�|H)[��D�֐W����bl"��o����b�� �!ד*���q����b��<o���n*�w����{*���e�K<sU��@�΄���j6�w�z�|�2Cɕ�o�]�Q�:>���y��)��������&%��'�?Q�W�����#9	��.�+4B,��ތ���+����Rd�8!���*�c+�}���s}م�<o���F�x8wK]a2����)h{��	�s��=e�����}�!֞��ߴ5�`3I��������~Cc����Ǽ���̲� �1y(cp>���z�m��ЙM��0�~u�]��	F�Z�'�5k���.��K32
#q������F@p+L�kX-ϩw>�Y�H�`A?��@<3V!��tr��w��m�j�w@��"o�]�K2r��%��+�ۍ1Cmb��2��h?u ?>��G&����;��#-_�.��)(��7�T�\�u�V�G��L� ���7����!����"��T�t���dc����C�Ϯ����V!�5fR���r	r�����8��U�c�4�ܼ���~	߈,���j�ü��Q�򀔳DM�L��@�,�,���d~-�AC�k�q�D�b2fC��4�ϧ����G����׮C���0��b�@{���t#���ü5@�ϣA�䔡�}����$@��*��o^J�4����aʻ*Nr[H-"�����w��L���$�[����o�c��Rd�ܬ��s�܅�(�g�GC7cp�E��_�c���B����=t�j=")�~L��p�j���&��! a�0zʂr���m=��<X���e�=}Y��^_f�J�]/�h�裡{j�K$�ȠE|D�K6��iî���[+��l�g�$w*��^�9���:�p�	~���p����6g/qéB]BHl{ˋ����~��3cM���U*]�mIx�^�Wy�S����PaVh�H9�0:إ����^�r�T����j�#V��m�2VPt����.	jRk'w���v�O�p� MЦ2Q����.D���L��$�ŭ�؀�bǄ���fV���Y��2���E�1cT;%l�.�b�I�GiҶY�����G+��4<_3�4�f��m�:�-���Bfn�@F����/�3&���?�B��D���]YN��@$Ie��2��FR1X���k{�;��(�Ҽ�l߲Z��t��KZ�h� ��1��g�����oK����Jv% H��{s� U�9zx'_�Qj��l}��J��ՙ�&��e]pgNE�+��G�� ��<:l����d��ʜ��%NQ�3~��`�������fI5�D��� �vs�{��1�-u������c`o���S:�+��>vnMd��J�u��:��XG��=F�~mO�u��y�j��gpM��!�a1�\Ӄi}![�Oj6T�`8���
�2�)O�0�bL\���xE��_j������%)%n�"����kz]�UH��+.ȶ�j��>�m����We�+�鍨9��\f�UIX)�5��W�6_��I5x�y��qw���jp�!K`�e݂�A��o�q��ی��b�8��j؍b�襬|^���n�R�卉ڷc2W���5	�}�Hx��E�R1ZF�t=ic�Vy�5
/~�6�di�[z���"�cG����kPl!�[hT�o>�0�2�Ow\x�M��k�Z�:����#|�E}�����x2����Bo
t�i[�J�nx�`��E�n�
���yw�;�����fNn�S�crP�;�(�o�y#�4mCz�p����{k~I�]�q�F�1���t��^6������A
�H���1��rjF�=�+�KdX��wH`����iA�ޣ�
/K`m��?���mq��]Q�Є���{�2<��(� �uf���Gm,Le2�.?�,�>��G��7��[<�mN�_0yU��ʫ�L�T0�u��G�jL������O:�!���,XT����/�V抺��M�C�A�Zu`!���f\���D}irI���i����Y��œf�_���ߒg*�-�M����3��{�M��z�q��8|��P­-Ti^�5���N՞bi�OCx�Lՙ��%ɧ&��a������0��bI^ �x�$t�9{LX��7�Y�>��>�����K�@����1�JǦ�!�aT�N<��-,v��wr�Չڙ��.2[d���U?�cLP3d���A��f
�(�}hGM�p1��B,c����L)*�Ey5tbvZ=�h~V�tp?�<�0���6Ma��i���{�Hx =w�:bd���&˽#VM�hw ʔ�:/1��ܲ7*{t�$?w�E�T��ir�� ���p�	�q]H$����7h�][5�z�V~1 ����o6q	��D�Bҷ��U�\��? ~D�3c׺��<��w�=بI�y�ۗˎǾPk�1
Yܺ$�Q���h�/؞-L�|>�jx4���T2�����}�ĔZj\��wE�vZY2�S Wd�2Pf)�Y�ND�^��V(�nA �"���U��Ѱ�1�(Y��<�t�ؙ71�1#�O�8(��U�G�dYuz��#&�+�Q���3ϡ�4�8��˷v_�t�@�2�z�3�����煌h�D�Nm'E�N�F�@n��e9f���Sq1b����{9�������7��Vr��
3��jh�Ś{�����ެ�O~K����V�o=���
��9��
x���� "�v�n�_j�a/���A�egT-N���[Vw�꘍F9�b�!�˛�L��@lN��3�`j�G��P!I��S���� �.�W4P����ul15�ݻ㨭���e�T:{4��H���\�Y�u�y�:�tG$ǻF��O���Ѓ�$�g�z����k�\&X}�FeO4�9T�Vd�GU����)Mf� M8\WhmF��a�2������4#�)� �n�w�A�Yz�y+5����u-�Ȑ��7�,疫<�D��s7���f�wU�1d���!G�@��]_5P8��v��j�9K����L���t���Ϯ�XC�ȑ�8�'j"�/�r�|(<��3Ĝ�z��ҷ-�\��M�	;1vH-�����R;��ľ_Xi��\VCn�5]֓�|ko�%R����c����#k���l+�2�[��.�0u4�O���x����qk�1��DŔ�>��||��EG&0�L=x|E�RS
>��ie�p�M�a��O�EZ�8
��I�gE�4hJ�D�p��ҝ�p7[�{���@2,���M���d�$~T�q�
԰�2��c���|,���^|+��.a�����!�m�4�+��,�>M'��P7�J��V��ԑ�����k�X��"�&�۪n��,�,h����X�On%Zh��HA��n@�T�V�	W��0rG�ћ\q:Qs[=ޭ�_�rз�:�r~�C�;X����:��F���L�p��RU\��%��@@j�p�݌�
��q��;a�,�"�Дݎ�9���&V����z��ըO]��a 1u�/�3�P����;�F�<h{��_Dө�� @�����H�`��0�F;g�L�Q�֍�)xL�:���0V:QH�mw����29BR����;6B�t��jj;�!�n��v��u�p�\���|:)�X�SՏb�����$��;9��YA�5A�����n�k�*J�����76�#�m�h)V�,��h����B�4����y#;�׸u��05V��;*��h͹v���ð,�Q��x�h��(�a��xG�ei�}W��)��z�/��B��c�XWS
�h���)}"��Bud�OyN	�Wn����
�)o����yȻǁMd��Ӆ)]XWsy�\�w�h���L1�˳��5d��	Lh��(�Rխq���_��a1�5�vDN�/=��u�5a��e�$���Z�������$iҹ��'ڲP�k_]L�>s��<�&��4Z��=����W�	�Zr��qSLʯ��Ԫ�E^�@*�F��D�@�7�r�
�\�V�Sl�#*��̩V��ň¿�?�7���1Pt|�91ZO��S�q��+^:�q=�y#&��h�v���`vV�v�k�����sZ!^t��*&R�{�88G�W�Q��}G!ދ?s�~\�,���'?A����M�/���~"��͝���O�q��ھ0��|��M-̮ڮ�x�\�h'a6Q�h_�ږ÷?u���x(���4ɱsU�G�'6�f,�<6yĸt;�G���	6�4[nL�Ė�ƻ�륚!Ԏ*{.�^=V`�F�ӝ�R�����W��!�y�v��sK4,��x�/;�b�H��j���`�z�-s���>���W��0/��h���vWzn�;B��#���z4?ǇLu�v����Y����B�4{��'�TN��>��X�w�N:r�?��4�|�"�� �e�i�HQ*4�����A)ӽ.�^>���FWW�eHi����+h�;����
�C��D(`�Iܻۋ�/c:�'*[+P��l��CΪ�șa��.� Tg����B^7�P��Vu� !�;A�d��nˋ-�A�ڠ�����6��z7�N�xum�=�{�W�}w[���X�Q%; ���~X�ڲ`I�4=�śYѱ:c�����\��Rؖ٨uG�9^q�I�	�ѐ�z�ɣ�;�"ǉ����w��b}^�-UC<<�p � ����a{
Y{Db��J�0���Y-_�����2s��e6��7z��1wJ�
!�X8��i���J����J9V�W�C�V_��࣓A9�w^Ç$�UF�ۆl�c8��9M_��d��yyq�}9F���dMlw%B���ߤ)�E��<�,'���9�V6~������~���~�TW�@\m�\A�M���n�g �%8��3E����e��$`��G��.(ͩ G�E.o�R{8��z,"K[�ķ��۲�N���׾ӪIǆ+UHB�z����6
9�nw +�9�Ԧ�"�c�}���Y�wf��[�X֩���
�bS�4�ؤ�y��f!bE�z�.x��`CΡ�&��U�s���g){�,|���.d��q�@��8_�gɈ ��)�e{��A r� �z���CUͤ��Z����}K����L-�y5���8����"U�/����'w&(	�/hT��P>Y��G�4�Â�����<���]���/���4ngw��{*���	)��=��<H,����Ұ(�����#��x�	���N�}�ړ�Z���b}�䡆�����{�m���Q;�se�':^��-�3�h���5|�d�h8u��k���@H��{w+���˫hJ�KT+��ͩԂ�@b��wp��J����t�J��"�7�u\���݉�����L����_��WK��x|(�e�q�@�2���� �I�t�6�0d�#`�>�:_�qF�D�h�Cj�H���Kl�L����X��]��v�5/�j`X��C�l��K%��ћ�g<�\���%(|�f^X��}��a��bI�[3�V�t��%����x�;�Z� '�z:߀��β�5�`C�ľ�Dc�aU���-i!����(��9Qg�:��4���˚b�R�nϱ������0}���f��a��W��K���*�i�O*�����~��fn=�K>Hgxcv�8[��$�aA!���n8`_A�q3ĉ~��u�Α����[R�5�R�#�H[���������i R�_�e�^���g�7D����Dp�7q,d]^�Oޟt��q����g��^l�5�z���7ϳAr��ǇtV2�(�*�EL���J��Jz/b �A��w��X`ٜ1�a�Ͼ��r�Q���f���^��B�(ޙ%Ʌ2�X�2�^��m��,�z��B�B6�~�($�%M��ֺ�z/J0�M�c������M��-�٤�Mf�P�7�M�T� (�yN�3��ܓZ ��	4�J��ԧ�!���`(�I�o�ZjG��M�Á�9n�6Ml-o61+�:�����/�~4{����-��(ф��6��YOЅH� g��;���1:�s���U��Ļ�j2�]��ƞ�����uG�H�."�\Ɓ���p���pJ�]��"aN/���.^�k7_f��(���X�Oy� ��HݛD=�DZe^�7D�L<��މ�Ȉ�k�ݾ�a��D�9-�`���ٟ,�zo6������3�j�V�'��> bjӝ��f.���h[��%����ϧIg�ܤ&�^��J��p�&�=u"��EX�7��"��
�U�g�T�&�KvsRf�3q��Űh����Η�{p�R����ׄ �0(R��Y�az�d���_��U�:@����d�1�TD60Y�ty�4�:�(ά���Q%̎>+w.�0sXv�g;��y�ܥ���YK�6Z��S+��Tx������y�~7��`�z�'{Sl����w���2dT-��"n�Ί`�%��2�]�yQ��%�����'-.����]P�0C"��}��Zƈ��������Y��k���b_	5��=�0k��Y(�6���~�E*��B{��YN��?����nu��ct���w�&����t�23�m���N,n?�S0�~��%ț�i����KS@�(�f �������֭��ȁe��riZ��]�(��"{���-�GZ���g�f�wo3�����5"���:�4/�4�{�@|1A,�Cļo�Àtᚑ�k� J�dIŮ�
Q�|��t!��	��E�W�>!$7���I����(���d��m#��$��o�RB������#F��40#��k�#�k8��H>u��4l���-wg>й^0�jaU&���2!?��^��k3u�xG� �o2��TB�cX�Ί�ٻ�s/�t�;n��p�4p3�׉��ǆ�)��hj����r+�%���]�v�%�U�d>�џ��������]��A��J��w��K4�>�4�#�,2P!�=o��p��Z9P���p�9��e݂���D�reS��bP���}���0*��Ň ����eF��*Q577��6���?F�{��q��!'�Wch�*�����hL �Ym��?��RD��Bl�������u=hLJc��) �Ђ˽R�����}��7��^&.�$�j(�P�p4D�qӦɄb�{������w �'.��t��Q��x��=E^ ���V�h	e�4  F�%#g��q���Zu �;l�̓cВ 1՟nwA��9����(ϐ�Z�!��{�xlO�U����?G���§L�?��(��o8�>��D�B05��QR�Y���FRQ1%P�av�oe��,Hƿ�@S����[ځ�\�-����t� l5�?V��hY��	i0�[��J�������lE8�5.g�vש.h�[/��4��?Y"m�¨7���'515D�Z8�j�=�sϹ����i�'���us�۠�~�=���V�l'a�0�k ��TªZ4�6���lƮC1Z�.vL�׽~����.���s�:Q óP����v �F[���"��PN�Р>Nq�o�d�H �e*B�mK��c�|޹(!��q����b�م���*L�i�ү�N��b%�o-�nA,!w���ی�*t�����<�p�ۗbф��ӥ��Ww�yy|���LO�L)Q� ��D���)�#z����ާ��?�ٟQg�ƖT�#C�6��+�@U,���C�������vi��l$8X*��Aҕ+��{�^!�}�sp<��	!bF��8���]xJe�߿�)?��_�
s4�j�D��_=T״�ֵ�Y߫Wk`
�ޒob��dĤ_�C����=���"߸����	;10kbp��%�e�z����`���~v��]�(Fsd5��O깬�_�F�O��@
:%���,�k��F��s+��X���w���+�AV�I�7z�-<�+
��$�m�7�ά9�����t��2iG�����M�$g3m���2
{<?��>�,HG�#Ȩ���R�_=�E�_�L��T��u���G�jL^����$��\��!3���y��T�������y���>��N�g��!b%�f�.�1*�r�D������_�nn�s�4�A���߿����ځ��H4��k�M7���)Qգ�L��=��-�-|�b���?b�:C���F�M�$`���o���֯�%�0�B2b��ǅ�`t�;7O���l����e��M�T��G�@�X|�p��Jd�����a�Ni��-��RZ�|w"��U��{cr[Q������cy�d�ƚ��sA�(O��G�4Pp�,��c�_`��d����tojk=�ޮ~��p,Z ���#̺ia���9%ʫU)=$�'���H�:�P���5�L�</>�_g�{�'�$,F�E�h����iz�ר-�K�?����$����u!Z��vd�Gi~u�b�����6�/���M�B_��˂�V̾=9~�l�c�_�̂$�İ*ؕ�Vy3?=˻�P8���t�ǆ����-浢�؋p��	߬j��ɸ�a2�i����q��j���w2�v�6?:� $ً2�t2�fiyD��l�#z�[�����4�3�����A�>9�Y;���˗�ų�1z�K߂��T� ��G �yY"�ܞp3g+���K�3��+4e$��$(}�ĉ���1_��@}�U��3���K���)D���WN8NB@[��e�t���3�1/�ҚPr�{F0/�^�<.���ދV��BNOh�sA��Z�����:ۧK���<�]��vH�׮O91�x��������~��L����U���e4��N��s�h���ު���O�����堌�{)N�w3_l`h�i?��R�IL
���^ Ņ0��d���iu1z�*�Ȩ�M
��]L:�B��l�@�fKu\��:���G2F�9�O���Pm����g��Pc!����\
�}8=�Oa[�T�$��W�G�)�c��m9�\Dޯ�����
��g�,AU�)}t�n%aC�.�uzt�?�����[7Û�"��8������ �Q0���3��U ��q@���t��k\JT5�:��Ѳ�l�j'5�K�6S����8�����F�$�����]8�fj�����!|��'�c�ĉ��U�Z���	�	�f�Hё38�R���ī�7i'V VpA�5�C�C�M�����'˖c~V6��vkw,l����e�0"3�O�k+x�o%�Xkᾠ����� �|�
�E􁧆_�xi@ϝ���
k$ki2�EҺr̳�&cE}�
�z[����&w3֠=���
^p7h|t��/ʃ���,y�M��Ĉ�$K�oq�5�߃i�&p�E},�^Q��u��/�_������A������>���=�_J]B��A���^��R<&k�#�Ͼp�(m��z8�������QX`p�%ǢT��^����f�����N�rt7-�h�I:�m_h�U��F1rtR'g~}���hͭ\�o:�9����UL0���#��[�̀ć���Q�z��� C�a^�+"֭���9 E&��NԴ�I�%Ojj�a�.צ|e�3m;(�y}�;�R+<5���*�Ӷ�� ����5�H�[���;�x���2�RVL
1��x*VT�H�H�m�+��j9�1�1�C�H��r��ڷ7����Q�O��#�츆2c6�n��S! '��_1�k3����w\������q#�p���8�Xc�����~�ۋU��-�;ϸ�����t��Jmwܨs]) �h�ǉ�3ߘr�"��3댉��"v��>U��>���%i��(��K�s�&T�]��8��,��>ןv#��BPbho������9���1�{f��݃�;�e )eT3����Q����q
*�����m������ae��*w
�7��6%K/?�������"�;W��kݓ�1_�L�km�<�?tI�D��ёC���؛���֘�L�*t�7��ޑ.��3�����;�x&�^~R���jɱL�1��R��ʕ��"����V�,� ��EN����xt��E_����ͩN�P ���%�Q�������Zv��;$���T�a�ϟ���I5���(��Z΅����l�V9�ٴ���չ��'/��e��D_8����]JB�v��ҿ�Y,�F#�%�YLb��o��m�m�M� ��S��ҥ)W[��\�tk.���� ��V?���h��	
pW[d�p��Q����lf`c5o��v8^`h`���p����Y�Yj{©о��B�5r�������M��v�d)��\^��sU'%N��%9LsF2IP�E=6(�r�ſaګ~�����[�ߪ�[�JJQ���r�)�� �vM����ҽ].3�����:���ty���}vI[3�d������p�!4Iq>x�%4�H�ef��Ԏ���14���Џ�F���b�d.���p*M+`��m���Wb�rDo��n��+wk������*uO?��!<+%�����O��"�|w�f9|��^�Mp�mN[QIB�V��1j�)e:f�A����ިB?���Q��n���9#�F=���[+���,f���D�R��M��0x�8��M���+W�?��}��<'�\J��Fm�8/��]g�ʠpO) Y��`��sUl�n����0�5��V��l9g`��V�p�Z��#�����C���l�aj�y��t112Pp�L̹�
,z`��숿����~7�]��#Ft�v�߇R����������C
ۅ+�wgr�L��F���+pX�hw�G� m�A�i���|��,$�/~�m_j�/'�>�4�U�2*��ַ���؂�ER�m�2k�V?-&�>;��G��[ȉ���NN_^���竭�PT��:uKK�G�+�L?附���}�7!t� ��wTP��]�*�x�B��&��,���!���f
�6� �rwR���i������������A�@;����{Y	�	 `�L^XM8N*�����D�b>����-�ʚ#�����b�k�C�CՇ/��}y��To���ϯ�S�0�(Pb���Ǧf�t�aB�q���h݇芯�p�5�yH.|@��w��gGJź<����a�8�N*o�-�([j5w����x���[ҕ�ڃ$�c:۴di�X����֐(��qG��!p�{*pL�c�Q����ٵ��t���=���~A\p���^K��2a�c�:�f�v�N=efV�l�ST�@*��s��/_a!ܠ�{"��$���E4ْ�v��@i{��N�'�^<�%�$/@���϶K,��(�E~v���(t�]�6��a�FB q��C�2̟��~��c[���'�%���#�y���|�CP��������?�������v���Ajf/:ə��2*���ץ�V�j
�w��6v���ҳ� ��2�b����D�.j��%��ķ�P�����rp��7_x�Y|���V��F�:1q�ݺ\���i�n}G!�3YcfОя�+a�M��y3�ԁ4F���%i������mR�@�_�ᨼ@3�ȃ��A����cD�MM�N�Lw@�V�eg�ү��1�1�Q�A{g�|p�;�t��j�o�,�����hc�����))�{sKW��{��4��G�츗�92�x�/ �	R܂$�n��kx��B~�޺e�N�s-��P���ؙ�P͓Е=I$f��� �\�#N	��36&5`X��R�U��I�y��.� �at�żƬ�)uZ�o���i���͓޷:i�y���*�S���u��:O�WG�dFA�O�Y��1���g(6T�!��(;\�Qv}��HO"R�To󒡵����R)Ӿ�ΐ�\�!�t���O�ͳ*��h��b� )��Jn������z� T��0��\����C�%r�D��+����񅙈��U���������5��j_50!E��m�M�j(�GK�D�:� ��$�)����w��r8p��j���Ϡ��|�^LЯ�
 ��E^��������	���H0���t�<R����,m�i�o�V1��5�I'D���đ:qֈِc�0r�Q%.k���l�� �'�0c*O/KzxTי��k�n���2���L|�.[E5*���̈́x��I�<��
,�i�һ�c���EH֣
T�1���'�8E��I���7����:\��OY,�sYM"P����$,�wq�0� [��Q��sh�,�ь8�����@�i��}�bE(��h\>���˾&�J����Y��?ւ�S	k�$��m��2����[�ZF��È-XA��%��|�2Z����q����y>� �r5>��I�<:�(���{���r~�k�q�~{ч)�=�:�e��qLq�g� GڔYM��nU+�^z��2#��߯�A��a���"n�C�KD�9�*L&D��/��J�-O�8�a���?k3�a��t;;��<0����=��E� .'T��H2G�^�5;Ut��[��S�L+!��l�V�c:HyQ�m���ڮ�V9𢣢2'�ij��.T�b��������vLpˤ�R�����FxS�U��(,+��J�����A#�؀�e�\���ݰ���em�u@m�#DVv���#�~ɳ�z0�ϛ�������㹤\��V
\;X:%h������]���Q�_]�V�4(.Y��N�x��#}E�=�ס���S��.�B�L�|D
#����}��B#0�O�Z9N7��W\9���Q
r�o�\����u�dh�&�WWa��\��G�֝�-P1��+��d*�>	zs�	��[ A�27,�%1�mv�q�(h���OK����Z�H��и	�8=�⵹��z�?��̕�]�u�lv�*U&jW�Ȼ�=Αe����	�ri�(Sz�H��숪�垷��A��￝�@8��rY<h׊$h�A�2#�8�za����������� �P��ٙ'��Z�������q��_^(�!=���&����ؙN�$�sk���LsH�Bt9ک&���8&�bWS�4��J�!xs�_��ڱ(ŕ��ZM�מ�l$��)�
�/���q�ܾ�,�p��U�M�!�"J�T�]'O3����B?����f쉋�M=47)�U �j'$��,��\y������5��·EA4�s���I<Ʃ���HXw���8��QD@�Fǥ����R��y۱~��ϱ���b�syΠ�W������蚉�_ ���7`YM*-�:�l��E�C�ި���;	�)z���飽B`GH#K�Y���z↑��������p��eU�B y��+�T�e8������]�|s�-Z�����ᐿ� ��i�n|*��@U�AWZ�.��Fg����.W��i�Ǳ���;k{�8�C��D�8���k۹~�Q|S'��8P\*�<~C�3q�G���7WT���{
^��UP�1u�q\�ҰA��@�y6�[��8�⬲��.��ׯ��x#����+�$���[�ݟƷq%i���1���üI[���џ�d�|�(̣�+�����u��:^ߒf��KA�~8�\�U�:w�"�2U�ԷѬL^�o^Cj�$p���BV���D�Y�;��'�0�������-�؅ ��X˸��a�_c�J����;ȁ��'Ås�SJ�E�W,)nV#�_���Q�!�k�w�=�$w�����l5�w��{_��	d��?�����CE�9����lx�p��͹j���7ƪ�'���9�2�~N�2zV�!����D3��Ʈ�G���>�;}���~ �B4�����M��t\�ec�$6��5�.� ��PE\�[�@��=�.�[pG�>�[�"(�w/�q..�vr7�{��>O��.��O�2�TS�Z,D�I�e��67��><�i���%�:U3���w�/D��K�����/�ǵ��1��3;��R'V�n���gHb 8��G^�'��>�؃��!��ϽF���Dn��7?렭Qp��=K�=�;k�sĨϯ��� +떇���@�a��R�v�3�����D*��9���ϟ6�� �4�R�I���ۑdJ���~y�؄��|x����z��*A�0�:7y��:���b5`Q�>_>�<�*.�Tg�k�y]s�	]�K�$�ʬ�#S�HkT���rޞ�	s�f�7]`Z����S�N��ȥf,�d���-	h"n�w`X���gG�ZcQ��D��^��w�-��=����}�Lȥ(�4�Zܺ��P��̯2lk]h8%J5)��ç���Y�Rr�/�2�]�Y��[��RK����B�4���Cn髒�����L�,&좼��&2��q�*���dv�n��S�Y���X����q-qi�8��S��@�H���̙{��~��I�W��S�oZ-\/�>��"Q�}X�:�qm�Z�x�g�f!�o���^\"��$�4��kӑR[|˛�وo&�t��5�A�� �!I�/
gA0|a�c!���t��[����7��I���>�Fl�U��#D�l$�f�(�i�Fu��yDm��0����n�#U����_u�r4����k�>�8 0��RU�¤�?!U���4��k�*����+±-��E
��e'&�Z:�X������8�P�F����;��t�F�<V��3I��h)��/h ���H�erAN+䈍�����v7�U*��>��ԟ�lx�w�� �؃{{�R�ڋ���a&+>�i�#7� Pw�oǬQ��k]9�F�ƚ��P��X�Üک�ei֦x՟���Ž|�}*p�����'����h\e�9
*,�I76I6��?�uu��,����W����?ڣ��L��nm��K?	��D4�a�yaАp横ڋ"L �7�,�-�&X��h1J���fy?�Z^3�����j��������U���}s���۸���X� X��:c��A�x�ӏE4oP#*�;�/{�* �/�%����9)���$ZK��;��W��Հ�D�מ>�H�MB1(��aZ�|ʿnl�V&��f�ծɧ�)�����@�8�*q��lBF^	�'�`Y!�lF���%�7�6o����W�դ]S�e�Қ�Z[0�\����g�" �B?lLh/ �	�b�[�9(�'�'���l��v5��%v���h�	m�e��rp�Y8S$�~���9M)5�k~�p9D썑�9o@3�3��¾�D'����:�Ss��D��=+�X�F�1y6a��ˠP��pvڪp�1�F���w����Ǎ56/v"#��S�x����.��ջI#\:�`V�	���$�v�=�[�U�1�f'��v:Yq3�ú#�H��;!s�M����   N   Ĵ���	��Z��wI�+ʜ�cd�<��k٥���qe�H�4͔6Z"<ɑ�i�6�3{�\2V��<d���fJ>@,o�$�M3P�i����d��f���{�9ݖ<Z"��5�����@�MC7����O�5��4_@�,F�@�x�cB�c���'��l�������.O8kq��8 �"/O�!�k޿q��	QǊ o"��>�P�޴4.��O,�Ӧb���u%MHy�A�{<:1aO�)1[�A�΀�H��(]��'�n�	B+�C�'K���=�XUs���X%�h u�c��'���ቨr_�'|P
�g�=-T�8�F�.��Dڝ'�!Dx�_�'k<|ku�ʣ,6��À��+;��@a�5f(�"<���>�1���"�D g.m� i�d�i��Ѡ�O�8�{2`S�`z
��1EDx��9�M��0�2^|"<�G&��\ᔰU䄎׸-�iγ
m�I�>a�L=�2�`�F;� ����*}�H��ӭ-XU�'U�]Dx2�JA�`��9�e�QJg�%�=�.!�?<"<��O���`��3+�����_�* �)��@�O �L<Y1N��=LdY����`�e�ÉMd?�%+=�B���<�1��UVU���'HD�8#��ʟt�O������*1�n�q���y��5jb�
ED^'�U
D*��d?h@$,Pi����$��xr�x�ݠp_�Xh 6'V�h˃�&����$���u� ��G"�E�P�-�W����u厭-��P��̜��y� @� d  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �    �  �  �    _!  �'  �(   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒��'��h�]���G��1y"Y;��=m����"D���)մn�%����;H���o#�	#&���ٔ�G�OaЭ�G��?7t-���Y����'D�8K�-
�8�n��K�E@�����Y����FPy2`����I�w���Q,3dq�� 2)̀jΈB�	�R	DP�`%�'a�E�plȠ%n(�(�HL��\rID����S$U$�r|�Pb�,=�<A�F1,O�����Զ�x�������2�BE�¼A���Y�7�l����b�<A��~�4)��k�O�D��~��v����$��9<��!�'�F�O8h�H4�F�?�2�r&ʘj�P�'?D���ȶ�^��S�O�x�^���KD�o��mId�՞|��E����
���K�ҡ��	0 r�|�5����i�}Y�)\(���!���26LP FƷu>@���*,[2�9�$k3LO�As��iluC���!a�\����']�Ma7��$W��BD�U���� 69xVkÇjl�DB3�\W݆��"`#4�h3�#	]`h)q��wr~���1���7�~����S��Q���q�' sV�a�/�!gyr8a�Aw�^���4�lR�k�3j�j$��x�6A7	�e8��4�Ə���s����-*�h�k�B�44:�ԑa94�� �
o����LLC��
Or�����^�>Y#�����<Y�P(xf ��OF:y@`�u��E��q4Ѝ<����
Ӎ�.��P �M�.�aGv-������`���Ɠ6�I��a�+J�����±x�Z%�O>���I�#qh�H2Ȗ)u:-{��i�{���
0�t���c�+!�؊4����d�;Z8�1�f�֜"��Jwb�;~�V���K�.6h�k%��|Bm��]���`1�Ksڄ��/ΐx�l�$o�~h"��#V��|�0���l�M��B!�=`1܇N��z2�!�cCD��W���靣�<�Î�.e/*`�cI�K�a�%AV��X�JE���� O/!��/J�<�+d� ?~��u�
�1O~��q�3JEn��3�'mO&A�Պ_0'@p�a���vy�ȓ`o�Y��!K3+&�:��[�r�<�����52/O�6m(�g~�b˗��5�WI�I�$��*��y���/?L݀�͕�@�<H@ĢA$�M��헉[P����x2j�!rHW2t�����:)(&���I�/X�H�'m�h��ܑ;���c(W�9:�'x�Lq�o�4ow��Ue+����'!.�8WΟ��<8��V�4�>IA�'��0�Wm��a@��Y�(�
ni��'�r��DLǒ#d�H�F�7��'���ӡK�R�b�*��+)֌��'wLD�g�\1'��#`ŭ*(��'66�f�	2ʱ�h�?MDIy�'� ���ݤ���PAGτab�'->X�FH��p\j���)U+ul�	�'~��+���\�tq��K�6l0J	�'F^M�2-��=�&ę���fp9	�'&�z��z�@���z|��'���[�M���D3cĜ�>��Yh�'���g'�%p(�T�A�>Sp�	�'[�y�5 ��:?�T�%!�>�v��'��5� �#�D�85nN<�9��'n��zB�wxE��I�Bl��"ODU4�/:�9H���+R���"O�r���r��d ,Q�ب�"O����.ف
�v@���N-)�yz�"O�h{�Nՠbǖ%�!�Kq��"O8|P�,�&@_�U� ��"�иB�"O��q�d���Lpz*�){���g"O�0����@�Q#�!�H8��"O��C��+E2Tbc��S���!�"O�����O�f�l��*��@Pa�$"O@d@�c�2HZ��҂C�A�f"OB��E�@�F�+�.چ&`�5�"O�d�P�NKȀhE��OFz�"OZM�a�
?d4�b!E��;cj��e"O��p�O׍Hn]2be�$nV�Ȣ"O<�K�@V'*�&%���I�aH}��"O�`@ M�d�Y��ɛ,4�Fl�"Ol��L�(T݈ԛ�Ԇa���"O�0bR� ?' Epg�V��썓�"O�0�Df��qEjB����DԊ�('"O �:bN$�H��BRҖ�a@"Oĩ�D��Z$��
��i3�2"O@�c�B�(���8vϔ2N�Q�E"O�( &�T�o�Tc���K�9J�"O�c狎+�X$3T�b�΄0�"Ox���cS�p���%�X�fx"�"O� *d�'��0oj��W$D=e�t���"O�r劝�1���Y���LƐ�@"Ox8�Q �kv2��'&�.b�b�R�"O<�CֿHN��EܕZ�>��u"O�i��	���(4�Ɂ\B�"O��Ai�1�^LI��Z�yZ��0"O�
��?f���i�7%Th�S"O^h�E�?��cqoر]��R"OV3e��-v����fj��U�Qf� s��cU�BoX�`�m${G�,������=��B+D����8C��4������t���(D�d���/ l�&��b&D�D�F�/Kx-����6�p\�p!0D��J�(J��HA��H��9/D��33D��)���$@���B�5{���0D�,xP�x�DY�զ�/���y%�-D�,��oU�^�bEqr�)94�ٱ�,D��SGK�Z���!a�O� Q��i+D�t	���/��$�c���,\� �)+D�����T/Ԡ�6bW8%_�q)*D�\q�牤+�ĉ��Y3S���q`'D�D�G'�0e��.�Jv��� �#D��(���)tDɠ�"j��1�N D�t��G��^�$ ������?D�<�ALW�}*Q;,�>c�E��"?D�� �i�&�6QZ%�Af���d�=D�P��m� Q`C���+D�(8R�g;D����8x�̜ґ�L4/���S`�5D�T�H s�,�q�H��'�N� wN9D��R�͂L�����K�j�� �`8D��k��3R����P�^�'��D`�m7D��O��Vm�
d;0���6D��c!��[� !p��)� P��1D�(�@��=:�DX���F�횁S��/D�@hČ�9n�A3�G�?9=�1Q��-D�d�M&>�RLR���2�b�`�>D��XF��f���z��!��9�L<D�4�e��/ژ�ɃǶ�,\�f�?D��	��[�2ج({k@�Mح�ץ<D�LQCN�!�X��1k]�WcjyF�?D�4�իQ�`�����Y�`6f�qh>D��!R+J�8�iGk�*�81�%K;D���d M�ZXy�jW�*�ň8D�X���J�0��)T'��!8D��!�����؈�0��3]ޜ���5D����R�N�(�D�Q���%J3D�TK0� 'h��(�M�&u�x �@E7D�����)fH��j$ޘE74���o3D�p�&���_��X��ڞ^m0�P4�3D�@bp��?�X��G�Y"Ѻ����2D���amʣ̚�
'g�#M�IV�2D�x�iٖzE&q��Wk<v�1!�.D��)�-��p|��t��b�M�&j7D���.)�(T�r,��s)D��bF�?&M~�����iS��:2�'D� �f@K�
Q���3톃RZT<aC�%D��3�/�.�ȔXK��:��!�&D��Y[y�8���(p#@=1��F��yb��kFMi��N������y��j6�,��H�&��������yn�,jz�2'N�4w �$b��yR��O����iWuh��ՋD�y*�!L�~	K��8U0$4[�����y��M����#'� F���s���y
� �,0f PI>vd���>� �"�"O�<�B��}~l2��^) D!"O�� ��{��r�\�#���"O���3$�
M'LTT*E�U�-[�"O�$�@��.���s��3���['"O�#��I<ے`��lĭQ�"O�$!H�p@�)ѠK�=�Zᚡ"OL�;`�>NVX���
�3�"OB���#$�1�f �`y�3�"OP �0�#Y h��`��!3`nQ�B"O��Oǯ}�h�r����^2,�c�"O(u��h����"��Rp}Z�"O><�)r�p��Z$���À"O~�x�-
	l��xa6d:mРc�"O ˂Û?Fp9�q�
*�����"O6���F]A���*�OQ�4_�y�"O�]�� �9.Ș���
�|\��4"O:�&��8^�)��QN�^��u"O6������n�m
���/7&�"O�,��EHҁ��/�N�k�"Oȝ��E�yXj� �j�	l��X�r"O�`��h� �4�#�&F{� Rt"O��â��ZӨݲ���
S���3"O24)�,��fLjP: ���Tʠ�@w"OjtCsI�kp�IU�T2s�|�7"Ob=�MߟQ���{r��2R�� su"O2DA�2e�dP!�
�S��9�a"O2؂�F�Z����b�T �~,�`"O<)��K�1�`jc� ( �Z8�"O*�CE����:���͂�v"O���SC�+C����J5F���b"O
�Q��7������!X��k�"O,X�S��?���1�jA�%��"O��8%HM
7"UzT�O=-�i"�"OJq���ѓ,�JZM��iD/װ�!�I0vL�� �N.��a�K5*]!�ʹk�nh���R-r\h�k۷3�!�d�z��(Q��vU�*��=�!��/Ws�=Q�A���P �]cW!��ʞ,��?g�NM�5�U'@<!���ⵒ�n� {�@&�`�v"O�A��ҕ0FrĀ�	�PV�"O��+D*7B5�i���oc����'D��s���?q(�c�G�A��y��(D�\b��9{\��$G9 0����'%D�pk���8��틵�[�و�#D��a�@��	�T�Qs ��Iq��B�.<D����ܦ{}�TCr��ELА�ǥ4D��+�S�4����ĕ�Tu�(h��1D�4��_�VXp�ⱭΆj��h��);D�t�Q�Z!V�2�r�KpD�8	�:D��+d��!n'��SG�F�#�8D��B�!V1���G(D�1>.���"D�x���VE���3��G�ZM¤���?D� (tn �7���c���&O��P���;D��;@�J!�>��e� ��BR�;D�l� a�j+&@�Ţ&[�h|"�<D� a�!]�[��	o��Y�4�Ӆ	:D��Xs�C�M�@MSD�2<��ҡ8D�l�D@�-���Ƣ��D�@C3�5D��x�f����`���M�g��l(2N3D�d���P(xd"��H��4m;D�Y5 �%����bo��F7v�T.D�ӡ�@�V��c!�&����*D�� 1#����p�F�C�T�J��%��"Oj��d!��Z���2�e��]�8x��"Ol��d�\�,�ƽp���xF.�$"O�(�n��j�@�p��L��!sq"O z 朅=���0-�d,�d�"O�m��j,��cv�ёq�QK�'R<�2�1Q@0vk�8^�U�
�'.��c*��M�hW���p"O�t��͜>l)��5xo��R"O|�"�S��p���(Q"̛ "O��*6.�
*�����ZQClA)S"O�a�Ł]'f���#̧�ڄ��"O~�gɗ���P�B@�z�>���"O��҇59T5p���4@ �&"O|�̅�'}ؠ�C �t��r�"O����C:B�(X���J�Xelq"O��jԇM�ɦ�]-|A\DC"O��k�n	G���T�>�p�$"O�	���|�X�S����i+
��"OX��S��1�$q����Ė)�"O��X�MD��a�#�|Z8�h&"O.���i��}��8���@ވ��"O̴�~I��L۝2\�MX�BJ�<�Ā��7����
�N�į�{�<1WgBUq�@F�f� R }��	��<c��̥a�޵�dJ�6K����ȓ%�vⶄ�A�½rM��(�n���S����w�A�kJH�ր�,�>�ȓ}��P	R�s���f�lА��ȓS0��#h�h�p��$�BR��}��J�� 9WmE�"= �������,\��"O� 1wF( ���1�hD�M��ͅ�hT��,M���釿*�����AL8Гhˣ"2de� �7�P�ȓG㚔����|���G�[�
�����`�T�\�<t� A�_�|݆�~����$N�6�B�2�阭E�b�ȓ	�	 '��L��CR�L�s}N��������2���)�?
Ը�ȓ_�8�v��P."���B��6��T�4�[�
/,`���.X*s˰�������a�js�m\�4}��J���d"�J�qq�,�cDi�ȓN
�xb�),i`��lÊI�|��ȓ ����5̘9	�]�䧎�-�P��CP�-I�fK��̑�Я��u��k&�E����??���Y�ゝ+:��ȓ]������2m̕��m�}[�1�ȓ7�2�P4�Ȋxf���+�4�i��n9����W�`��aG�)�6��ȓUyM��>U&�� ��HMnx��>}:����G#XZ>��j�	vن�)aT`��K֒鮙S6%v�$@�ȓ=U0��a�D��<�cQ�	�F�ȓ��A�Q��P����k�8���^�R��CR�%K�lM�(�N�ȓ�
\��_cZ��B�읳.�d��v��d�sn��W��LC����t��:�$9j��f�-S��496�Ʉ�o� ��k_.H��ڃ�ծF:��ȓlF�m��P�,����C�X1��\�ȓd<����vê���#�<X$!��G�e�1AXe����+��U�捆�=j1���'*X1��C��&�Ry��S�? t�th�ii8��g���j��!"O�mpS%R�B52в!���)���˃"O$�rժ6�ʡ[�-͓A6�z7"O6H�D��E���I;8 ��'&V��#hڌ>�dK�b
�e
�1�'@�	��S�-��P �W�	��q
�'����
X?rAf)���� i���'e�!h�O�7h��۶d�&	�8 {�'��1��!H�kT�����FP��'���Ȳ $�±�cbP������'z����@�����Sy��'��e�QN�!��IR��}�*hB
�'�j�0I��S%�#W��l��ȡ�'��9@ ���   �  <  |  v  �)  5  Q@  -K  �V  �a  Pm  Jv  �}  v�  ��  ��  H�  ��  Ф  �  Z�  ��  �  c�  ��  =�  ��  1�  s�  ��  �  ��  k�  � �  X �% #- �3 :: |@ �D  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�Y�G{���˾R5$�Qb+�jBƅ�7��Oi!���l8��Ӄ]*W>�\����]O!�ė��ތ F�8#"J��7Lb!���P~��#���(%l�(.ԜoI!�d�0c>��=`�r$,�
�!��LP!���6HٮsX~��!ݺ�!�Ĕ�m��G꟯i�̥sQ �W�!򤃛]Q���D�o��Z`A03�!��R�6j�l��B�^ ū@��;Ol!�P9��$`b��e&Ī���c@!򄊡jX�QTυ#i��A(PhˢF"!�D/2��`pB�]�6�`�6��9!�dEE����BݙB~�tK�`I�W�!�DV�=�i�H�!(^n8�䏔$g�!�$��mMX���9OT���n��O�!���-
l��WoР>J���NE�ni!��K�4�VYP�ɑ����+L�xT!�$�4<{��J��! �PhX6*ʨI�!�Ff^��PR*C�lʹ����F!�ͪ&�����'�4j�\���(�8\!��/�:��������bN	i!�$�<PⱫ��53���{J!��@�S�vL���?ʀ4sW��*t!�DT��`Iȧf yƬ`�c�]�#�!�D�p�,l G�.x��ᲆ�T<@Q!�@7_�����=�"|p0��-N!�"F^�cbI��i��,�g�:'�!�0�@1g�żm]�,�Ҭ�
3�!�d����(�qKrأR+�<q�!�ںO`�i�눏`�p�5mܒ<�!�d?B�>�1f��~�>�#���0b)!�$C6h���@焐K�и��)4!�� 4IAI�R@`�g� @K�C'"O�ِ��3|�V9Y%hS?<v��"O�y���<9�t��'��X=�"O�a��Q�/k ����$�Lu��"O08DF��D��6.M02㼠���5D��")U+e$l�ȶcX�6���Hu*8D�T�N�,N�n��4h>~��ǈ+D��@� Aƒ���eT�VD4��%D���q'�
1��Z&�Q�9h� 6D� ��a��1k��T% ���J)D��(�f�4��US L��1�z]���4D�p�3ϐ�ѡ��R/BI���&2D��I��.��s���p�� -Y����@�Ta��ցE��1 �oÓ�y��SZh&/\�SIRݲ2��y���(@��Sʀ�9̸3�j#�yB�ZM�z��?~�t�>�y�NÙ[8,�kWG!hQ�\�C��+�y��/����C�úkl�Y�-�yҎE G���롃�f�P}��eɱ�yBbӣ6OI��G�s�@�a�NI�y���(�=�"#�1lu�l�7' �y���8l<v1C�G͌eI^yD犠�yHг w�Ժ�=S]��������y�c�'�8*QE�K߾ț ���y�]*�������9,�ٸ o�#�y��M�j��D�2|¤{�G��y"#̽���h�A�a�Z��1Ů�y�)�s�0	���\Z�����yr�	z�H���+1��	Pj�3�y��XZXt�-�%`��ʤ`%�yR�IJ�P�����XWI /�y2���U?E���Ԍ|�j�!���y�c'�V��p�P��Bh7�J�y�:v% �𥑮r?l�i��y���T[�)Qg��}�`P1���%�yR���.���8�C["#�v��AOV��yBn�b=�A�X<� ����M�y�eD�_"J���t2a�5�̂�y�*��X`Ht���:�xED���y���1�J�Bc�"��,zu"OH5�5����\�B�ʄA��=��"O| [A�Ȯg��c/,�,��"OBy�hP3&>(��AI*�H�s"O��Ru���d�B�@(�&���"O�j�"�	�S �W�0�P"O������n[�}���>K�Ь�G"O���#��q�)ڒ@#Gt���"O��S��CT'��kR�Q�11��)@"O60�«�j_���hٶ4#�"O|P�d�I�j@@�2���4�,"O�@S��W���@�����TwB�(C"O��C�C׫Ix�Qi2���H�X�6"O�ɱ�dZ�{��ͫ�/��	l����"OY�!/\  ZR��BHW)+pD�ٗ"O�q�@C�lx�#cgިk���P�"O�lK�&T<T�����o�t�2�� "O|iA�,���٧��#&�YzU"O\ȲX*��9[V�C��|@r"O�-�Q�j ��	���`V�lA"Ox�ۡ,�:m�d��qJ�i��h"OD8bC ��\��c'/0f���)V"O� �/<]���z���F:z!�E"O^���'�����+�"ԋ$(�S"O� �x{U�jHXAY�̓v�x2�"Oࡓ�O�B"؈ �Z�6�1�"O�Y$�ِ$���RS���>-vd��"O�����?Kr�HA���X�=��"O4A$!8<���M��L�`��'z��'��'7��'��'��'tj�1���<w���G�B���'\��'cr�'?��'a��'"�'R.@q��y�|$�QՁx�ځ g�'��'~��'��'�2�'���'6�0�M��
���U��1�� p�'�r�'n��'R�'2�'���'�Dq���+K>��`�3������ş�������џp��ݟ�����4qlڌ^Q�<��W P�t�ǂ������ԟ(�	���Iʟd����\�I������Ԫ�^�h�c�I���3��P�	�����ޟ<�I�,�I̟����h�7ɘ�!���4&��W�����JΟ$�	ڟ������	��	�$��̟{�f\�`��<h�c�� �x|��iP�������$��ƟX��ٟ��	џT�����I�Ε�!�����P��
V����D��ޟ����@�	���Iʟ��I��|�&��D�d�r���>�D�$������ ���0����d�Iß��I��$��6&��,H��[�e�6!W/_���ş��	џ��	�t��ȟ,���,۲�%M	����[�ТZ��Y�������h������	����7�M;��?Y�R��"��8a �i`��0k�	۟8�����
殮�PHE����1@�x�Lj��@i�V�R���4��$�O��ۛ}`��0��F|r| o�O���\.;�6�9?	�O&:��1�4�ƆX��@�3ϔRk�,�c�U!�'jr^��F�4���Mx:��n�2
�1�	]yB6]�r<1O��?mC�����Q�_�R����k=���^.�?����y�S�b>i9���٦%̓UF��,�= ����q�eΓ�y2,�Oܱ���4�T��͠^Ԡr䖌ײ#� �+
��d�<�J>�B�i'��yR#\$o����T�^�4	0iR4�O���'/�'��>!B	 [,�"Ǌ'>�J�b�%�M~��'�rH�D*�ØO�pL�I�C�cj��I��ԕE,��S�#ξ?;��{y�󧈟󄊡8���ł�	J}�4�� �����W$#?	$�i6�O��@
u��m�⨕ptV�CՂ�l�D�O����O�s��a�����&�����Tn�x�ҥ�����fD�DbY��䓜�4�F��O����O��D� ��;amߔ{�ta˄0V#&ʓ`��H��X%B�'���T�'EV�/�8PI�����|Xƌë�^ꓟ?����S�'.ݶhj�[�RjhEI�{.d,�!�Ϥ�M��O���Ǩ�~B�|�S�Ȫ5��'Yn8�g��[0�٢�����џ�	����`y�cs��̪*�O^e��&��Z��ոal�
X0&�92��O.�n�x�a���ҟL�I��0�h��Q�պAV6L`��]���m�Y~"�H, F�T�w����!Γ{N�DHtN�
>�ā�'��'���'���'�����V�\SR-�sř�"�;@#�<)�~Z��,���D�'|�6�>�Ęw��� NĩeZ�a+~'��O��d�O�)C�P�\6M=?!f�W>V��"Z��d���Ed!��	A��O��I>)O��O���ON	 ��(~ M��DOw���f�O���<q��io�x��P����|��3�<p��6lWd k'�����H}"�'ҟ|ʟ8\ S�	O32 q�	R.L�)c&��'�\���b�P��|1h��D&�L{��N�X�`�0o
*&$�DIH��<��Ο���ܟb>�'�F7-��6����I&R���H �
3�Q�3�O����Ϧ��?��S��I��ˣ�5o>���![�z�~�������B_릥�'�����[Eܧ?\�z�J-)��Ժ'��U(�Uϓ����O(��O����O����|��C�/vqQ��«'Yl!�D-w�^�?Q���?�N~Z�4䛞w$��0(g�-�5���~�P��D�'�b�|���ʘ���2O>�[�ڪD�𙑉 �>�I 3O����KC�?Q��3�d�<ͧ�?Yv!�`���Gx����d>�?y��?���Ӧy�@ F���޴�?�a"�4{�j���)8 �8��R���'���?i����]���
�5` L� �A���'�  ���/�����V��~��'���Q��A� DM��8��!��'dR�'��'��>��ɗ#�PL�t�Ug���3���_�M�	�M+�+��?)�EC���4����NZ�Q�.|��L־,�`��a>Od���O`�d�7�6�+?��/�;R�h��i�y0�.�-�f��G����$���'3��'���'L2�'L�� G�i�ʵ{���N;j̩�P��K�4JZ0t����?9����'�?���ɤqs$�x� ���БW���ß��	^�)��NI�4�/��nh{2��i	�d��F��E�'e�����Z?iO>�(OH����$2� H��'
JcR����On�$�O��O�<�A�i0�5Cs�'�@�ӽV�� M�2|�d9�ɕh�4��'��ꓼ?���?a��XDE�}�᎜i�$ ��M�����ܴ��$�>,�Ƹ�'�Oh� �m0rD��+\�聀��N� @9O����OR���O��D�Of�?�'�:W�v ��*�|�b��蟬��ß���4	�Ґ�'�?��iz�'b��Abд^'�����3 ��p3�|��'��O��	�7�i%�iݙ@
ޚbHP!(����O�hpRa(�����BE�'��	џ���ӟ$�I,1��%,������$>��x�Iܟ��'��6MW�!��ʓ�?�,��,��K]�<%T���D�=�����9�O��;�)�$�X�YQ�� J^b$�pIIR���E�5
�.O�	���?@�2�$@4R�F]z�ķf���w���D=T���O��O0���<�ѿivj���g��g^T�!��
� L�A!	����'�6(�����D�OXͻ�D@z��I �J�g��@����O ��L�R��6�'?�;W��A��b�B�X������Ee;}��&O�.4�ϓ����O����O���O �$�|2� Ҽc\��VJ3BP�e�7�]&^"�֫ t�����0&?�I��M�;	��:C��7d�DX
��W*Qp���?N>�|�����MÚ'R�6�K�=(�##�� >. `�'���S��x?�I>�(O��O��t��- ���%���(�C��O��D�O��D�<�ưi��l���'��'�x̋��SAZ����$�oR tz7��E}��'�R�|�j�	��4R��&	�pxTg������Vr�H��8V	1�`�h�S	R����s�5I���!`���8W�0���d�Od���OF��.ڧ�?1����ȝ�e֦Z \�RN%�?��iC�y�d�'Q2�q�>��]�`�p��A\�t@���3����۟(�	�����oǦ!�'�F�����?5�a��89��E`�D�8]:>��g�N�/'�'?�i>!�I��8����\�	�ppD�q�m��O�Z}��ܗn�й�'Tf7학,����O���,�9O�	A�M�"��p#���6�xq́Q}��'��|��d	Řz�d��6*ܐz�zt��-�d�u�%�id��lјu��,���&���'u��*�d�2L���8 \T9��'"�'b��tU�Y�4g�����8 �׃kZAB�M�D��T�9�6��^O}��')��'�T�e��='l ��K%S���1v�BM͛柟ؓ��X�U�������L��6A�V��P��CL-V�A�:O��O��$�O"���O��?]���#I�M)ǥy,���S��ğ ��ן���4S
�ظ(O�o�Z��z�س'�E�2���b7+��$���	�擙2���mZj~₅6�,���,sӚՀ�N	$7$R��C��|?�L>-O6�$�O��d�O���e�\3*ۨ���n�/V�0���O��ı<i�i=n��'���'_�S�Mn��Ё�#��PȐC�?k���aB��ߟt��[�)�o�9������=z�hj��P`��ů�.!*O�)�?�?�t�!���8C�� B�l�,!jD�P�)D����O����OH��<9�i%\��`S YA��P*�G��a�gN!�'|�7�#�I�����O\�Khْ̖,�߀,�.<�dm�˟<�I�gZ6(l�i~�l�f_��Sf�I?1����%��e�h�e�4�<���?����?����?*�Z 8`L�t��͛V함lNp)��˦ɑӊ�����ʟ������y7�P6H��u
��[�T�a�dR#sb�'�ɧ�O6m�P�i���8̔4#�>��x���)��dI3B�����'��'��	����	�[��̀��>��� ��O"��	4�IƟd�'2�6���P�4���Ol�$�9_,qB6E�%vl0{1D��Y���<ЩO��D�O �O�1;�������f��|��c����1�/5U��o:�S�U��d�O��1D��H����FbV�񃀋�O����O��O��}R�ZU�Di�������Cy�Z����ԛ6��uZ�'a�6�&�i�aR��?�B-�-�r�(T�rcs����ڟ�������mZG~"�<
����ӗV,DF��
O�r����R0�(X4�|U����������	П8(v@�?%R�pN[�*p*�Xg��Sy�+g�R�pAI�O����O�����G�K������;��y� i�?�ҥ�'b�'�ɧ�O[v���(H8Jd
*�u�\�IGoZw���|s�%�?i>�$'�d�<�E/{���:���7Ҕ��J�5�?����?)��?�'����ͦ��v����KPkډ�,ɺC#���u �As��/�h㟬��O(���O��ę/昑�����ոgm	:g�δ��}�>�%�!ҶF�?�%?-��-��i��A���mM�G3��	ܟ`��Ɵ(��ܟV|���?���\�M�z��R�R\���3E��ПP�I͟ ��4,��t:*O�um�Q��22*2����;�\��k�%'��	؟�S�E�c�<�ed�d2�[�"�n����J$�Q;�̞)r��Io�Uy��'�B�'s���I��Y�D��	���
B����'�%�M��̈́��?���?q-��11w��v��C@*�©���t��O���OޓO���J  XD@|�\,t*�r$� �R$�T|u�}����
Q՟��g�|2$�x�ґ�D�8(UTm��·/jp��'G��'���V��iٴ%����JV,J:��P��,����?��yěf��p}��'��:�(�4e~�aZ��g����'��! q������"ej�}���g��)� ����A�%�f�z�"�, �6On˓�?����?���?������-��!�0�C\M�hPė+A5
in�>[�l�	ٟ���m�؟�Q���K3��B�]��ǆ)k�2�p$m���?)����Ş ���I�4�y�-��T2h!E۸!В �Pmn9͓��� ��p&��'�B�'�f���¸/�~��F���~�zH:�'���'�]���ٴ>6�Y[��?a��JX�`tN�2K(��I�7	�xu��r��>a��?QK>ң�f�^ᓳ�V"��033�O~2g�(��#�d�0ǘO���	2GA"��A��%�Q��.s�'8.�"�'���'C��S����'#��[[,�`�F2#P}��S؟��ܴMn�� ���?�ſid�O�]�	������1	 �H�B
\2S����O��D�O���֪xӪ�=�0���L�?����D$kH������A�y���z�cy��'�b�'�B�'�r�V��*�/�K��s�NWS��ɰ�Mq�Գ�?q��?�O~j�0�5z�A$�qRPؑr�T�����Oh��.��i�Y`2����P3,ݞ���N`�Cd�-
��˓;u�|����O<�2L>�(O�X2��]�&���KB'f:�};�C�O��D�Oz�D�O�<9�i�����'��|8an�
P�`�JF-*G��'8�6-+�I����ON�7�[��Ȇ@�R|�ҥ��t����u��?�M[�OЉ[��-�
�!9���������3�T��Ȅ]@�D#S>O����O����O��$�O8�?�"�9��}��O��v�X��П��	şL޴^��5ϧ�?Qf�i��'{��T'���`ǼKԲ��4�|�'��OͶ��i��I*IR�G5��ݳC!
�G��b���;��>���<�'�?���?!��k5��[�E���Q-��?�������9��,�䟠��Ο�O�x����˔H҉	d��?7$xȨ�O���'���'fɧ���=w��F�:U��Qc�$O a[���g�>7.?�'�@�	~�I �d|@�XoW5ތ��L�Οh��؟0�Iɟb>=�';06m	�+Pxy�d��.h�v�ÜsIv� �B�Od�ęǦu�?٠Q�l�	�p�!q�n�F Ad�D  �A�	ӟ����٦Q�'N�j����?1���ko�>),��u!�/z0+S6Od��?����?����?����[aP~\a,�*	�$�;�!	3Q��ul�2����ş�Iv�şpB���#��C#@��%�����O�
0�/� �?����S�'i��Hڴ�y��P+X5B���,Hh���L�y���($^�����4�&�Ԋ<ȉ÷�\�;���ud�&�����Ob���O�JΛi�/b�'�Rl1Y��gY a���H^�x��O���'���'c�'3�x�ҋK|N0p�Q��+ �(+�O�`0�� �]Vm/�	��?QVM�O��@�k�/�6��r�-_��a�u��OD�D�O��D�O�}��+���KA�۬(P��� �ČT�vl������(
>��'�`7m"�iޭ 
��B��jb��(�B���d�(�	Qy��N�#����4��,D8d�T��ERP"P&q�N��JT/T0hhZ0�|RZ��	ğL�	����퟼�al��Nڴy���%t.��@�jyreh��a��OV�d�OҒ�P�Np�Ѕ��Q�@�%;X��0BP*�>A���?M>�|���B,o/���Ă�7^L�h�d (�`�BX#���Œ4 V���d�&�OP��@iÏ�6S�iC"�C��8b��?����?���|)O2 l�a6��	0u�53���G݈<�V�]X�2���M��b̠>y����H09!�ݩ�V�D0�L�ߝ�d)�D&}�|�|w4z2��`8�O~
�;$�t�S� =i�(`b)1� EΓ�?����?����?)����O���˝>>3��a�쓂_C$Kd�'���'�f7mn��'sW�6�|�ņ�j�>�Ae�>.�^�p�$��K>���?�'<�-�4����hT;��
8`��4HSb�,���l��D�	�䓙�d�O����O\��ҝFb�Ix��J"3�%rH�3���O,�`��´1��'�_>���ٖp�^P��vN e`ud%?	�S�d��؟L%��'g��q�WFF���'�D�><�x6��0�ݴ��4�v�
�'��'���QjK�-�z��5y�ܣ��'��'�����O��I5�M����Pv,R��C(v6�<H��	<�:�!���?�!�iJ�O���'�$M�e=�p)G W���B�)Z�"��	!�ZYon~�c��rv4��+��	,K�fL��e߸o�F	s��6�j�	Dy2�'�r�'XB�'��X>��wl�_�����L䀜:Ҭ%�MS���?1��?QM~:�9C��w2�Px�Y�]��YjB��FƠD�!�'��O1�N��(~� �I(�l�I��ɻIe���`KM;97B扜tn����'�Ԑ&���'��'N��@v�j5@sH�4�) Q�'4��'��U�8`ߴ^x�����?A�'H��s���� d��ԎVlh����>q���?�J>��-�.ܻE��D���(��X~R�;5���i��O$����i��DP0E�A+��)��"�I�3
b�'#��'�b��ҟ|��&[�)���SD&(Ѳ}j��ğT��4��D�,O�in�d�Ӽ�$E
��*���݉8p���,��<)���?��?�p�4��D��N5��π "1�����o��c���35��b;��<����?)��?���?��㝭wQ�|"fd�SA��q&%����ğڦ�;aN��	��8�����|6�\/U�2Q��l	i�IП��Io�)擉���8t(�2(2^�*��7Bf�k3O�Ʀ�'ܰ��|?YN>�/Oћ.�?K.�`��N��2�2�+V#�O����O���O��<��iP&m���'H�Eb@!��"�7mR%%���'�6-6�ɇ��d�OJ�$�O�!(�K��K�(UQ��R� @��D�G�B6-!?� �>c	��|b�;ʼTː���^�^��C;.Ql���?���?����?����O�=�$��PQB��V+gPl�7�'1"�'�67Do�,ʓ��&�|�dυ>�ԥ�4ᙝW�(E!���jM�'�����ꜳZ/����8�s��&�I�b!��d�h��0 _,G"|�� �O^�OV��?1��?���ܠ�JaJ_�*����u�P{� (����?�(O��np��IƟ������a t[�HS���X�����$�g}��'0R�|ʟ��2d+[�p���)>ԑ�U-({A��3$� 
I�i>��7�'"�D$��X�#ف:E�T	T#�^�9���Wşt��؟t�	��b>�'7-�4�($� !��"�p���V?��E�!��O&�������?��^���I�O*��K��LD ��*E'���	��@����e�'�R�q�#�Qܧ
NDR7�Z�D� �s�g����$�O�$�O����O��D�|
!$Q�!p�)���U#2L��hS�n��������'������'7=歷��F��k5�墎�\��͉�e�O��1��ɏ \մ7�}�@)C���X�s���K�6�D'i��i��ź'�lS`�zy�OGr!�-[N�!Y���<|XႧ�"?��'"�'S�ɘ�M{7�
��?���?����N_Tqp�kX"v�}��͵��'���?q���S-�Xc4ޓ4���G� ���,�'h��A�؜4q���)�1�~b�'�n��q�+oU&؛QE��0�@�u�'i��'KB\�"|r��,�qH�㐃4a�x@0M�*7Zժ���W�
R�'�*6m"�i�a�Cmɡs 8d�S��2	����j���Iޟ��ɢ��dl�~~��L�%�,P�s�AN�Tpν��ڃqq�� bj�����4�&�$�O����O�_%�$u��	�E|�S�6q(B�IO�fN��'����4�'�����޴v��<�B����[p��>y�����O嘼�妛���4Ȓ�;R����!��� ,�=�U_��B2�G����o�	By�aU< 5�pbB 9Ό�q�3r%r�'|"�'|�O�	��M#�)Q9�?����"$�`��ŲSX,h��I�<�T�i�O���'�2�'2�Ѓ�٢�ˌVn&��*��{tP�SB�i$�	�$��3�П������&_6��0���P�����
�����O��D�O����O��$$�S.b�$�0j�j�L�[Q_���'(�|�
���7�����e'�LK��#0�{f�0 ��b,����'>�<�i����D� |ړF-ư�� L�T�1��<�2�r�Iey��'"�'���"~����O2p�����P���'��I��M#s�Z��?y��?1(���-6�b�L�/��)�������$�Ov�d"��?��SM	�@��+��
U���2g�(?���h�������ă�Z?QI>`j�: ����/ND���ℙ�?���?a���?�|�+Or(nZ#Nl�i�7�ߙql�$J��
�L~�D��c�ן��ɕ�M��"(�>��t��A�X�����E�ϙ?c�@A(O�	j��~Ӯ�D�u8�����)O�H[�`7~��I1��F�@Т5O���?)��?����?Y����)O���O'j���p�&_�L�1m�!dr����ӟ���~�Sӟ�(���3�d�&+�����ќ
�DA��#2�?�����S�'Rh���4�y"*N��=(V���16��@�.�7�yr	ړb�:	�����$�O2�D@�m���U��,fr�X���'zC����O����O��"���М�?1���?�׀Z�"���b�)K���9��͍��'D���?a����-�x�Q���>� �`ҡZ=��'(�=�!�H�z��4��şة��'Rn|��Mn�X��,�#;���'c��'���'�>�7�X���ɜkr���F6���)�M�7���?���Zj���4�F��C\�p(f�s!憒bJ>�2OD�d�Oj��/~�6�1?�����E����M��iZ�!�)/]xSA��W:�$�|�',R�'��'H2�'���a%͉k*�p��(�^�1�_���ٴ�A	/O��$#���Od����:)$T�`7́0%9�`�V��n}��'n|��T(ǟ>,��+��b�2\j�M��qe�iU��4#4���O`�Ov˓K���#F��F@�6� �>d���?���?���|
/O�=l�<T0U���,� j0�
u|<J2� �)����I��M�¨�>y��?���d�(��~o�h�&�Y$8��l�T���M��O��˰�Ç�2����w�Ќ�����b�� ���.@��(�'I��'�'���'��⬀񊁯
���b�<~SN�IM�O���O��ȔC�E�'�?��i��'2�K�!Ss_����C)ܱͨe�|��'M�Oo(,*6�iA�ɃL��� *9�i�#�B<	���)$�v�� �Ӄ�~�|�Y��ʟD�	��Rqc�n�JP�+Q��=����IjyR�uӖ��#G�OZ�$�O��';�X����
沜�0G[�}�u�'��듶?����S�.T ��%Pv$�<^��:¬
�B�f�5o
��eQ���@�"��W��#	\B�kǂ��;-f��/�o	����	՟��)�SCyR�gӄ\��T Q�M�S���f(bq�M�1�H���O��ln��.��֟Ȼ�bQ�aY%jH'&>8X���LyLZ ӛƚ���̐�T�����gyR�@��y)�΄�)|#�	3�yRZ����������Ο,�O��Co�7[��V�0����ᅵ�M#T�ҭ�?)���?yO~"�p���w��w.��x��89��+`P�� �'���|���EO/��:OP	�1�P C5�Y0�aʷT���f1O�V�؅�?��*��<ͧ�?I7ΞC��JŢ҃o@�I��
�&�?9��?�����hQ́fy�'�$ؙ��ڟ(��щw,�}�8����Q}��'K�O���$FL�=��d�5N�#�:������h���u9$�f��r���HS����p%����۱,Ш�+�I
���	��,�I�xF��'�je@EH�.�pQ��*YQ��Q��'�7M��^���O
�n�o�Ӽ�W� V X ��U�l*����<A���?��X��4���F�(��x���Y���!g� �aB�x��b�:��<ͧ�?i��?���?1�@�z�ޘ�E.n���dg\���զ��p��fy��'=�Oҧ��/² ������A�S�(�ꓮ?����S�'De�P� 
�@A��9v��b(H���*�M�_yB�i�,�������;)3��H"K�
�����)�2K{���Ol���O��4�8˓�V��4=��	s���H)r��Q��Cy��n��4��O����O�N�K�f�qv�&Q�̩ ��W,X�:%�|�N�^��%2Wo�?�'?���5sL�[�����`����#4�����������	����Q������d�
��y�A	*{�J�����?��g7�f������'�x7�8���1ξ8�����|h��Z�l���O|���O�Q_ 6�"?I�����0�Ǥ87��@
Pc��R��9����ON�{K>�(O�i�O<�D�Ox|[Ǧ��:�9ɧ�	4�t����O���<��i���j3�'�r�'�3�<<���՘|�D���Jy��[���쟰�?�O~�HGw���6��MQ�0Cc�ǣJ{`��7�L�4[�i>͑!�'D�H$�0�%'�Z�Y� �ɧ#W1�ӊ��8�Iğd�Ißb>m�'�87�H�#P�h���+]B�aGǭ9��c�O�������?iuP�4�� g�� )wF�.df���S��/=�<�	ӟ 8�ˆɦu�'N���*��?}���X㑗U��Aj���d�N 2�3O˓�?!��?q���?q���
'�����G�;DL<��&^�:�PlڞNz���	ȟ��	T�Sȟ������&E	�4+�)�F��vA�!���?I���ŞD&2�	�4�y�"�A�F�K�0 
���I��yri��D��ɚo��'��)*3C�#-5��到&�������Q���ش/C���?I��*����W5�Q��K�UI�����>���?�O>�n�s�̭���'%X �%�|~b�54�p\�'�i@����'�"��;t���C�H�-��)���y"��7�DbѮ��#��`VfA#j/�eӺ!Qe�O������?�;oa��`g�a|lI��,�i�ց��?���?�����MK�O�n�c����M>b��E��5m8(���<���jL>�/O�?р���q�0\X�����*e�"Ml~�n�~e����O0���O��?��A�Y�p>�1Q*ۈg�Έ�w��+��D�OF�$��)X:�&� �
!b��(E�߬IH�l�*yӄu�'�fMC�D�O?�J>Y*O>���9D;",K2n��S!�-�0�'9�7��+�6��3f�b`3��+m�
H��F��$����?�]����̟��I�$�@=��(�1�M�uKY�+���d�Ŧ��'��Ț�k	�?ʤ����wr�11V���I�а1� T	]��裝'd�bj
�&�f]Z`(X4n"�8�Ɓ�"��'���w���F�?M)޴��r��<@���=ɪ�f��"6��1O>���?�'E���s۴����>�=�!�,�r+��lyĨv͚��~"�|"]���?1�C�,�h�A��ޡx!$ �3��K�'F~6͖9,��$�O���|��d��#�\�4��*�z�TG�E~��>���?)J>�O�j�0@�� ���IAa��|%���Ɩz�h8�N�L\�i>����'g2U$��i�Δlnd��b��^������2�$	ٴ|�>�S7�N�A����X���K���?a��xh����[}�'c��I�$v�a(��F�cZv��4�'����4��v��x��x�I�<ITG�D�@Ai��K#��OQ�<a,OB��$(�P��ʇ�Urܔ�$K���1n�i�P��	۟8�Ix��ě�w�� �2h�>?�F	#���SQZ��'�R�|��4GؽL�&3O� ��c��\�����W�E1"�9�1O�Ū��]��~��|�^� �	ğ���P�9#��J�Ɔ�M���l���X�	���jy��k���[q��O\���O^11],fͺ���A	B�E���4�Ʉ����O:�)��?���inƌd
��F�Rk�������c�¦m�K~�QI����	�w���!�K� �F���J�0P��	֟|�	ҟ���q�O��"�!���[��;Kh,;Ǒ#M!��yӼTYu��O��_ŦQ�?ͻL�&�Q�Fˀr6��jB&^('W�`��?)���?��g�+�M+�O���J���t �9|[T���-L�h�A��LN�'���ӟt������$���l"#�U�6VP�h�CɆ����'7�6-Y.=K<�$�O��!���OR�16��WЈ\���
+S5X�Br��Z}B�'��|���W"4�$�� ��[2�,KV����TBf�i���
n�|��&��8$�p�'h(�!���K5L�bn���pyZ6�'�B�'������Z�@:�4u�)c��.w$L�	{�R,J���=R���̛���r}��'�w��cCP�NAvt@@�qx��/2U�֒�Sd䕣���SB���5AD�H�!��s�%E_ �-���y�@���L�I�����ן|��U�I4*`B (B�N�;���?���?���i7�*�O_2p�>�O�i��H�?(��I�۰&��b�<���O��4�~$JB�u�<�Ӻ[�����2��N :�,Ms�X>J`|H��f�x�Otʓ�?���?����puCA�XG�joA�R�UY��?�,O
�mڎ����	矀�	N�T��X_v03�P�B����aV��yB�'���?)���S���C?v�B�;�`��l��+�JB��:�bW�ñ<m60KcY����b,�w�I,��B&K�t~��)T��h,t�	�X������)�SKyr�n���P�.тp����F�:8&���%��g���O��l�e�����ȩO"�d���^A��R�Cd�ɥA ^�f���O��!ҁb�T�V��`Dk�?)�'��Q(��I'����r/ҝ� �1�'^�������@�I���	v�T�ҡc���&��i2e"?v7��`
���OV�D ���O�imz����G8��p'4�Ё� ,�ϟd�	p�)�ӛ�>lZ�<�I�io~풓����҃�[�<����.1;`��������D�O&��H)?�H@�nW6o$��W������D�O���O��h,�D�S�?���?I���n�"�#�H�"`��n�8���?��^���	�`&������"D����p�h$+-?1֍�#��9��W���+���DV6�?ـ�Ó$4��r3
 &d�=��n2�?����?����?Y��9ﺸ�+D[��Y�Fdݵ5�Z�91�O8�m��-����	ɟlRݴ�䓗?�;^h:�D�۹ �$`#W�`3����?	��?��K��MC�O�j1����CO����I<55~(K��6�FIqN>a*O��d�O����O����OZ�:ud߂�$9Be:'�>�i���<AŶi�8-@��'�r�'��O���BsxT�	é�5����� T�&��?�����S�'N�܁����
.�1z$ʟ�w�r)Р�̏�M�DU��;�O��Ua��#�ġ<�Í�&�v��I�'C�Nq�PC�r��޴��,#��,5� ��4�n��c(��K�0-��Lt�&��	\}��'W��'���Z���&��ap�nc!&́P��m
�i��ɘ4]BjB�Oz� &?]��9�6� a��i-$��vj��P^*�H����b!&D.,BP�NR��8����d��� @�4ʖU�O^6m �d�*n����H����0P��O?b�O��O�i�%�T6� ?��n�����¡V�X��)W7:��q�ș�?9�i)��<Q��i�%(�cE2���2�� �OD�lZ��v4��̟p�	d�T�E�/<��3$�n�[�o	��� Y}��'��|ʟz��bㆄ<� 9#�^+Q/r�󕉗6|\�rEd�$������ZV?�O>�тϳU�� i$LY�cba���x<!�i
,3�O�"5>.!���%�5�F)��c���'3�7�6��9����O�HS�\�Kh(@K���z ��s`��O����$� 66?9W� ���ky�A
�.P;�"ŭYkR�Ҵ�yZ���	Ɵ�I��{ӄ�Į|2pD	#IL�����F/�X�c�k�f�	�bW��'~2����'�D6=�c�F�<躤`WC#a�X����O��b>9�cE���$�V,�u�[숅(&7[���^"���W_�h!��R��욖��k�P%E
�"9u�0��%?��5r�P�g��qy�7,�L\$o(����-��X�DM���U�ҢZ
N�41 �M��+}��ɋ�"���#F�}z�􁍵/K�ʓ���@2ߪ �""�� ��(A�]���,<Z�����&0 �Dq��Ʃe&t%@��W�r &�C�KA3�,�%�Y:��e�D��<X`��t�ɷQN���Z�^X�|c�dQ�s�Z=r �æD�Z$ �D�(_P.��)51O��'�9HQ3����G�q�dA�M���?���]�O��<�4�υM�T�����%����'��'K��'$9�2�'��qTl=�� �)0}4-�b�&y��oZ�d��fy���*^���?�������w��@zDeP+t3�I�C�E�3։'��'�&�����?)h���z��D��&��p�@dv�:ʓz؂�X�i��'���O����#���10V�x�"�	�F0�릝���:���ʟL$���}� �P���H�h;�$�4�\����3�i1�y��g�Z�d�O��$韮��'6�	2�R�(�%E	����$L�]bܴ�z0�������O���ثV��ʅꈖ�1��,�G�B6��OX�d�On�y�h�H}�Z���	\?9�*7�x��r�S�c ܙJ��Y˦�'��	���'�?���?q�*��g ea���!�� 	UŞ��f�'��9	���>1(O*�5���H�AanQ�G6�XI�ۍi�t ��_���b��k�	Ɵ ���H�'�,l[B݂w�๰ ��
3���2f.� �������O��O����O2�1�	1~Q�fOdQI@iX8���D�<����?�����䎘,�V�ϧ[; ���"��@��X�~P�o�Byr�'��'b�'LҽR�O�X��ȿq"���cف("��pfQ���	Ɵ���sy2.2�r��?Q��$x��r�hS�E5:p�OX33o��'M�'g�'�Vp2��d%�D���hk"�QyC.*n��'Cr]���"�(��i�O����Ԕ#V����h�bf�Sf���j�R�ҟ ��-*����?�O�j��� Ŕn��-3���ٴ��Č
D`ԕm�����ԟx�������,iL� 4�E��
P<�D�Р�iL��'}8��D&z"��.'-b�	�G��M�26�*,��hnZ�������`������|��@fJ���6��B�n���q	���'���'�ɧ�9O��d��	����-�Ȫ!A� ��g�T�o�� �	�� +j�����|B���~r�c3B	qw����!AY��M�����x��3?9���~ǤKJL�鵁C'x�� '�M��3?�t�*OL0�O'�O$]��S�WT ��HA�R����C�I=�Z��?A��?1,O88P�W�J�(H�F)�wϤQ��	QB<��'�L�	�L%�H��uG�*�p��1� �_����^��M3��䓅?�-O���YN�h�S@�h�a%�VV��@7-�O���*��ПT�'�����4_�\A��4�2�"�?t����'ob�'��V��K�T��'W���e��K.y�#��4���R`�i�R�|�P��֟줟\�֊[�68f��u��>M����a�i��U�l�IZ��q�O��I�?ט�L҈u��k/Hk���Ë�<0O����<i�Cs��u/@�0Ճ�̿l���ؗ����On�ʑd�O��d�O������Ӻ+D4���kW�J��h[�(ӛ�'��;$#<%>�h7�QwvT�ԅW1'
up�gu��1���O���<�����?�r��'�`Jwo��[���(�BA>��$���b>��ɥ'uf�ET>A& 9Ҥ��0�$�ش�?���?�����p���d�'���X22�L�Rd9�ԴK�cF�F���'\�'�2�g~�'��$ߐM�)h]%N|22�V!��n�㟔���Iy"I�~"��	�e6�Is-.W�ܰ�r�����O�D�B�d�O���?��t�B�/:}Tl'��TY�yH/O����O�㟐�Iz?�@*#�!���=#C�Ϧ=ڴ�;?����?Y����$�3���' 줄�j޳#��h���'�fD�'���'6�'��i>u�ɟ0^*��P ݩEt�d1[�nmV�K�OJ���OJ���<9KC�X%�O &h����B���b�A��E��Ix��c���3�d�<ͧ�?�N?�y��� �ҠbË��?��E�`Ӵ�D�<��.�D8[/�L�$�O���ƚ��5�xX"�(��T�mx��xB�'�	ׂ#<�;/�P��S�U�w�챑�n�
p���oZjyB�
?u�R6� {���'��$G%?�S�ӵ2�����<)�=P�B�ݦy�'\�'�������f˖*#����GcZ/u�tI	�Ӷ�M[ч9z����'S��'��ġ?�4�Va�^�_f,����D��hl5�Rަ���Ο4�IM�)�'ÚP�	�0�Y���?|���#pӈ�D�O����z�S�d�>�ǂ�Hv��*�,&��|P+%���YK|��?���z��b.	~�~�BF�<�А�U�iBB�_0�����OFʓ�?�1y(t)ʵ'�; ��@k�� yM�}mZ��\��r�<�	�����P��Cy"�h��8��&L��)������p��a?!*O|�ħ<)��?��R��Dd��nx���`����P��4	��?a���?����"%_vD�'a���AО<��5�w��, ʅ�i���韘�'�2�'�R-V�y���[��a�ňY$��j���P}�6��O��$�O����<���,f��ݟ�cW�A+DaC��	�]��L�#�"�Mc����D�O���O��K7O6��O*���AS#��y��*�T ��*�Ԧ�	����'���SΫ~j���?��]i�@�J^{Рi�Zr���S����Ɵ���7xİ�	n�It��U�:d��LI]�&�SĦ��'_�D��hӤ�D�O8��矲էug�>d^��x��U&{����qN�*�M����?����<AM>ь��"��@���B�Kc�� 렂֜�M��&X��'�"�';�Dk�>A.O�,�0-> �8�
�Ja^�ഢ�禅���l�p�'T"���O��0b@ɀ�f�r���+\�u�`�����	Ο��	!P�*�Ofʓ�?��'=��B����8eKVO�r��۴��2�Z�S�t�'z��'~�� j��˅7t�ăg�=K����6�iX��	x*���$�O6ʓ�?�������-}�MRI4��I�' V<��'q�I��x�	����'��zV�֡"�~�P��Ή4�|�)Q�>g]h����O�ʓ�?����?��-� me�MSc�V�4�4]���� J��̓�?A��?����?A+O���%�O�|�%�Uk1�q�R*խ�T�Do�ަ��'��Q������$�ɖ?�l�	�����L��%������y�b9K�OF�d�O���<�m5�����փ�.^��4�j��X��\'��M������O��d�O��X�0O��'��3�Ě><0��R[{8�(�4�?������e����O��'f��jL�3&(�v��+V$���գrf��?���?��mV~RU�L��T�v�0�Ι6,x ��N�$A�,�n�ny�Mu� 7�Od���O��i�d}Zw��<���ۅN $�(��@W�*�4�?���9%n%��?a(Oj�>�bv#w��čv���8c�]��4k+�A�"�i���'���O��ꓪ��A.Ly<����X�k�!�fo	��Z�lZ	$*P��3���2��'U�p���j�:�2Q`3���M���?��V��x�fW���'���OЍ���F�Z�v4#�#�3k�� ��i3r[�0�G�e��?���?����#0o����M�'��q�TK��S���'Nv��v��>y-O^���<q���^�Em�p 3#��	;zt�&��i}r�I��y��'W��'^S>牋?���Z#L��s�� ��Č3��5��N��ħ<a�����Od���O�8�ukH"B|e���R/V�bh9$��%��d�O*�d�O��D�Ot˓H �2�����Hp�����Th��b�i�I��X�'�'�R����I��LW&x��ˌN8I箒u����'�B�'��^��P6AF���i�Ok��' D9�+��U��J7�ǬV����'t�	�����˟�q <?q�',�dz���M� !�DcC�d�Z���4�?����䎗k�0&>����?%z�D.XeSgJK�HL&����?��SJ���������E$t��HS��¯-Y�1�����M�,OTt�s.�X����D�����'�����D� '���0",WK�=��4�?�l�E�����O{�({�>`�r�
���S0��۴/	L1�i���'���OۀO ��ٓw�L���JY�2�ƀ&S��tm�"�lM�?9��4�'��b�	"A/�hZ�d��K�+Ӧu��˟<�	�B�pExJ<Q���?�'<���c>`8�p��Ï�&���޴������S���'ER�'/~%֋�)O ��m=/�ܔPU�|�x���r�L��>�������Ӡ̈}�r�+��U�aPE�JO{}�Ȋ�y�X�����&?�ʣ�^�LY�|��A&����҆{��Uӌ}��'��'y��'�Q�EË����Ć,�<$jޢXR_��������	}y�/@@J��s����2���<H��^�1�p��?���䓃?��Y���͓\�����"c�
�)X�LQ��R���	ٟ���]y.ǧT�8���4�V.,ydb�9:��U*BU��U��A���P�����Iz��F�u�����3��	�	�"ɛF�'�rV�H��ƀ��'�?��}�P�3�I2��v_���
�x"�'(�KE�p$b�|ҟ IY��� �T幦l̪؅L���P�@��BU�MK�Q?�	�?u
�O)�v)O>�Rm�U2��5
b�i���'#�I�f�'B�'q�,m�#�M�[����ާ�̉#2�i��`fc�Z���O����0a�>�#�[
21e�]�W���[���*���&�y��|����O� 0��d�.4#ǋ�-w� E��l�ڦQ��ğ�b휅�IşX�O��O�$ �EO7_�j�/X�+�
l��L�}�'�h�"�D�OJ�$P.�\5���^9C�ր�E�F&	��m�런!��ۨ����]���'�B�>�A��?Cy4)��@Y�Nxi�`�@�	q�	��p�I������Y�a��1[� ��}���^���!���6�?I���?����?�K>���~�DGӆ�#&�U'\�z��S�M��o~R�'F�]�p���	�8-�ɼ8�, ��I\�w������B2�J��ش�?���?iH>	���dӸ	集jE�r��5�B%vk44��X���$�O��D�Oʓ"%P,������?��a�0`U��Z��@C�9T6-�O&�O�<�5�$8��+�>>�y�Ys�lZן��sy�L�G�����$�81�	L�(�N\��jԥU:P�jYC��p�	h��#<A�OM�u���1U>e�p�T	T�)X�4��d\j�Эn�ӟ\�I������4�i���ڜx0��X�x�t�iLb�'�حK�'�N��<a��$��F[���ȏ�;p.(���K��Mc&7A���'B�'��dI�>Q(O�5�b =N�����%�m���D ���k��8��O�B��(q�t��L� s�]���ݘE�7��O��D�O�����x}�\�p��y?�a۫l�������3.I��T��u�Ity�ᔋ�yʟ���O��D۫%����
�"g��@�1��;�^�oZܟ ��Q����<	�����Ok�p���T㜐�p�:$�5כV�'צ�ښ'n������ٟ��'�l5�f�F%q1�=�Q�ͣ!4jpXr��j�h�����O�˓�?����?��
�V�B��s�9M^؝�5E�
8�l̓�?���?���?�+O���S�|� `볂N<i���Y�k2Z�	[�iu��4�'t2�'�rB�=�y"g�/fǂ���
�*_��deT���6��O�D�O"�ľ<9#l�[[������>�(���#ԹnA��SP�FM�6-�OR��?a��?���<a+O�Q�4��C�0	�D�-��i�٦	�Iȟ,�'�vX��~��?�'Z�*]��N	�A&�����9Nx�t�Z��	��t�I����h������#��=0`G�dX ��*]�[#@m�sy�ڤV&�6��O��d�O���[\}Zwn�X����[G��S�m
�2���Cٴ�?Y�$�j���?����?���T�S����¦c	u�^5�g-��?y���s���R�H�Z�~,ۅFܷ0=ƙ(3M!D�T+�jE�2�B�JQPD-��U�α��n	&I:\Q(�"_�ɻhQ����eA�=:��/��A���V�M��z���mH�@Y# dQ�q���].�Q�G�	�/6�q���e��$��qp���"py�=��@�sf�u���@�:x��'�%;^u�	^ß�	۟�I��u��'�0��P�VM\;k�v���Q�t�b��.�������ޥt͚�z9�YG~ҍ� 0W�\�o�I���e$��xr�,`C������W�A�j!�)$���82"=���N� ��ie��$H����F;d�E��ԟ�F{��P�IQ����#�9b3�8�!򤑒4E��Y�ƛ ���� D51O�D�'��;Y|ى�O��d��
��̺���	R�~���&�(Z�d�O��ʂ��O���y>������� � ��~��h���"�h��@��ZE��� %��t��<#���Z�T)�FI�9Y��J�n	?~ؼ��ɛ$Ũ�d�O�˓o�Yڀ�ҽ)M*As蓂3X>5�<qߓ-B:�2�F7a�R!X�JΕ�����R��f�U�3�\���G����ٰ����y�]��Iw��*����OXʧ�ꥱ�r�| �Q��'(���+�I�>$C:|����?I�%6�(l3Q�ǅHΤ��!���)�|���)p�:��hk�^�{VT��=�aj,�Dx��0ҧ |ҡ�T��?�"�R4`��pd�q�O.I¥�'�2�П(�s�� H�H�`��A�q�|�c�=D��2���"�2�e��7���B��(O��Gz��\�GD�u�R.�1!�4��LM!��6-�On�D�O�h�R��=n����O����O�8G��Zԋ��Tl�w�U
+*x�OVd1D�X�XaxRB؀%�L[ӏ
}�F��a�^0FR�1s����e�ASq��'��9��+\bp��&E��"��i�'���
E����'���'>L�1杭Bq�]��V8!����|R�'��ѱ�# &�	��\����O@�m��x%���ĉ0X�Rp���-�~!�a��+m ��j4-R�Fd��ON���O���O��h>�+�kޕ�TՊ�.޿\��)#�U�sv�8���px��y2-έ@��g���$�ڑEoLl�� `Sx�� �֧0<�y[���><|�e@�狤e���$�O��d�O�ʓ�?a���9\Sj�r���=ۚ���l���y�j"<#�*[5�i�L���'E�6-�O\��'p��%aN�_�(Ze�S�!<|1�ȓPQF5���x�X@rt��
m$�$�ȓT*F����|U(��e�b��ȓ(���_T�k�,�P��H��<�q��t��T-Ӵi�NŅ�sa�1Ȣm		�f�33f�Xo�������b�6(�f����L)zOp=��qq��5怰sjD��/���4݄�1���I=8ƴ��g^�G�ܡ�ȓN��98���N�4� ��M�0\��e�fZU�L�P�����3�|��ȓt."u�� ��8H�6b�$���ȓ5��=�!%ЎcT�ɻD��I�8��ȓ"��,��(��[f��+G��� ]���ȓ8��6+A0Y�,ÇB�{|-��9%���h]ኌ!2�N�]T��ȓvXn��,�����6�U3F�:���
HY�Ι:s�T�!-���t$�ȓT���Y��ȥu	j`��h�q�ȓ
�TH�v$d�RA���d�i�<�U�_�2k~��l�Zo�T���~�<�2�0خ���"89"��� �w�<�U�@!4��J��ہ�"H��}�<a`�H�6t,�#CH#���%�P�<� ��i�W
�b{��ɪFh��S"Oh# $Nތ�Fۼ��E	�"O���@�ʘtd��AТM�T�l�P"Of�Ə��x��ǜᰐz"O��'c�3UW>�ȓc�}j�
�"O�IJ�]���=�7��JJj�2"O �Ѥb�|",��SO��,7V���"OHe��-�#@s
�@��!�hLy�"O�h��ܘ*d�87M�� ��q�"O�́ԭԁ!q���+��z}8P"O(10R���I����ʈ�-�v�{�'��"���^��(R4���6`:�i�'�( w ¹B�Pm@G�D?�T}��'c��Gi\hUj q7Iʱ_��H�'Z��3j^\��X4o�0 J�k�'^�0d �4Z����S��3 �a��'�H���&��4���0���2���')P�z.M8
��2��F'%��P9�'�� �L	;{��'�ِ"��-k�'5�<�gl�f,Ñ5���'v<:Fn�c�tqҥ�n����'N��I�*��i�ĪZ�"ԋ�'�ܕs�6!.�Ai�4��D��'��y�q�ܻl��`(�/Z�p����'�"А.��a��Ɖ�l����
�'��@�n�,�v!��lW�i�T5
�'+z��&ȇ`P�=���c���'2��) %�4&���v��U�Nx�'=!�^�ڜ��&�5N��E)�'":M��+�
fBD�i�e�K�v��'�*D�'\>h�kF �HB*5	�'%�i���٦a�~tk々���'�|����¡8�()�.ȕ
���A	�'�^�2���1+nhǆ����'3�1c�۷3$.��g$X�I>H��&�ZX{�e�	n�|IR���{
ZE�ȓA���X��[
(p���Aẅ��M�:}��
�|�ε	���R���ȓ1�
�r�h�F�V`�Eɤ	��T�ȓ.���%(�w�PI$����@�ȓ3cp��(L^XX+�'�`�L�ȓ�BH�d�U�3���PI�A>���ȓ>��(3�F+6I�p�kI�J��-��k�� �EG_�$�x���Y�Z5��T*x䫴��k%@�@Q�\�0ж܅�ô�xo��Q�t�`6Cq��]�ȓ?�hPᩈ�\���I1(��/Sv��ȓ�����R�VX9�߸�R�ȓ�p���E��>a!��9!�Z��?y�]�s'�?����ѻEӚ%��E���c%�?D�����:Ψ(�@���$���� I��N���4!�5�O$�g�'Jj]P�"e�
I�����g��	�7Ř��(Ɲ$�J.H���b'�(�JT��E*���4�'�~YB�fB,�!b!	�-�H��A�R�m�T<X���/��M
��D�0d��A�|R��cPz�����)�
E��v�<�F�M&	������*���'�S�,T�e�6��Oܬ	�I�;8��ƍL$��B���j����߅+��0�4�(2AA&�2	0�)��)Q)a{F0��L� 4Ψu�%�c��P2o-$A�B[�2I#7Z�Hq�i	(*����zR��&M�V�A�A�h�U�d�&O6h�0�-^�DС����<��o�1�v$�C��[�6���HK�@X�O���7iǝCR�@
Ó]�X	Ӆ�)}7�u��m�a���'znE��cʒY���G�C�:�0��^D��KϚY�H=)�3H�$�Z�֯`x(E8�P�F� ���@aE���pX$�s��{)D0�&1Ԍ�;�]"��!�jY6�PAQ����xH�wƢ>���2�Ft �)L>^�2��O��~g�C���r6V� RhI�&�;^HѲ����Հ�&��@��9�e�]#I#�a��&C=��Đ-O�
iZaZ���$P�@�@`u��6#(�O�cbax��S0�E�.ږ�I�\���-�*z����Qi߿r���U��zyB"�<��3w,\�u��b�� #�3h���'E8ZIV'�\0dꖵ+}� U�O�O����E!�:DO�ā��V1fCn�	�'�"2$%ےz�t�C �Ǆ���kE R#�2,�!C_JyB�%�	��^�j��O&i��� wb�X�	� A�l����'�LЄ��qQ�t�"�)S��Ĩ��O�[�6-Z�n�d� cfΨx�����h��b��\Ae�P�Ut�]y)�$S�� �"%�f
YA�˵"lC6Y(r�R]���G�p	�`��2:��p �H1g�8�xP��˰?	���%I-VY�w��%�(���FByb�-r������W�[�B,)vAB����O�X6���J3.`n9yA�[	�yHܗM7jрp�U�`��9�go�.%�|�p�-H'Z�'�t('?QƑ����z�H F��]FҘ�U@V)���[f�ȓ5�ʍv�ܽ��B��7�Hd����j��+��9{��� �џH K!A�6m��$I {�m���=<O6l�,Y ;��l��ˍ$ 0�0sI'F�YF�.<.����&	W��DC��B�鄦Z��2�⅂U�hqO\�@�"�+t����\tU
��}
��eNH=H��#aXt8���R�<�T#T5�̠Q����>��틄�B�S7�:(x���O$�}�՛2���^+8t��t�h��'�t�:��޺c���KT ��V%<������9"`����iQ�3,O2�Z&��+T����O��+t%�@�'Z�Mґ��4�ȩH�4>��l�B��p�(�i�d�h�<��$!*?�hPi�8MR�� ��h�'"�1�D��o�O������#"�-C���0]zư��'���Y�jܘ&�6��Αl��|q�'8�x4 Iw\
�x���)k:����b�м�3�^�z\Pw�Ѝ��q���ĺ��N�ۮh�ϓoiv�ȓv�: a�)��d#�(1��A<����6QԑҴ�\ #��@AP��O��ȓd�&}�w��'���ȓ�D�X�Ą�4�|�ش��%u+ve�aֺXm41��Y5<�1�'�X-�t�ˈ"|Ⱥg�݆���sfT��f{�(E^�2�҆+ߜ*���#'�!�DB�I�H��1
R���a[�ᅔ�Q�h��IC�M�?]S� @�݊�)���Ƽ�i��/D���I4W�|�Gg"5�n��GB��`3e�)�)��4�7ɍ�
�%��#���28���?D�lG��J�6�p�J-�6���C�>�7�Q�O_a|"a�hQf�cU�ܣ!��`����y�ٮ/s�8B!�Xqc�ͩ�y2��";�O�D@�lX�	Ɯ�y��ޕj'.��$n�>?�:��×�y���(,be�`Õ�>�Ρ�@.ơ�y2��K�N��f�>�豷�C��yR��u�=sf�O,<���U�y�Oą(�$�:�%\��B��#*H��y�mĆ.54��!*��
����y��
�
B�か�[����)ƫ�y�ʟj��X��Ϋ#�jiX��U�y�냭Xk�x�#Q�� �e��y���=^�H(x�(�#����jƟ�yr�� |CΝ���[�K:a�b��yBb�]���B6�}-��;Bᐐ�y�Ϡ-ADx���?�<-:3n[��y�O�"lwX 7�*%����7�K��Py�-1�HypĬ��4h��3�mh�<���&z�Pc.)~\���e�<a�Ƀ�/� @DG��
���LEV�<� [	!`p��G��2o� !buM�m�<�����Q�d�0&I� 2�Lj�<��"��;W|l{�.3*�����m�<� �@��G9b$��
�ZX���"O��1��D�'�t&�WJ�"O���I�@v-���@�X��x��"OnX���F�YH��K��ê+����"O"<H"鋵hMl4�@�əY2��"O=���7P�ʌ+uh]�<;��"O9q��'	2bvZ,�\�"O����VN�m�嫙��d0�"O~�;��A���'��P<q�c"O���s+�#�r�*�(÷;(�S4"O�e��/\����طh�F���"O� ��f)m�X��^i��c�"O� �ѪE�Y����6o�"m����"O���e^()�ȝ��(�v5��"Oܕpb����jS���1:)��"O.���ĕ�-�^�Cw�[�O뀔��"OV鐡L/n9R��EJ�J�(,��"O��p��)~��a�5QZ|��ce"OH@�6�O�@*�	DExa�p�"OV9�`�T�c�l��@zaH�yb"O�@�e�����.pR��"O����!�Y���3�ń	wT q��"Or�Xw��mܦ�WD� �TI��"O����υqf�D1ҡ�/%(����"OZ����]Xf18��"0ܓ�"O,�*q'�8�H��%P�z0dzf"O��XQ�7[��9���p�V"Oz���7G��TЁ�K	�VI��"O�a�W:W��Pvc@��Ƹ(�"OF����1N�BB%�H���Q"OVL#�B�5����	��e~� s"O���G��O��]���K�Wk0lK�"OH���"�*:��X�%@Hcf Ч"O*<ѕ���g)���E�k�l�"O�=3��>¼��%P�@R��"O�h���"KQ�|X�F#q<ּ�3"O��#��)@R�UgF%M�"ON=f� �8-
<��e�|��#"O�0Z0�k�z��@��޸�k[��ybkD�!`�$	�쌳b�謣2��=�y����ڐ�gC�?a|%�b�$�yBGӗ{����F��J�[B�C;�yҎ��{��	/$�Xr7hLrHX�	�'ڜȂ�X�a`X�B�Z2,q�'H�@R������{ ����k�'��|j�&/�&�*�+���R, �'rR����_�d�L1�H��		Te��'}����Ǎq��#��?J���'���h!�	;A&��2�˞S��$�
�',���!�X�7�Fx{���#GHP�ȓa",��厢kS�X��Ǐ�F�����s��%��"K+7���1�݊V⭅ȓ �dT($'�*�^|b�oԮ&Y��:���c�
�'&v�zVcP+A<0��'��度셗N)Zq`�'g��ȓ1���&%P )&�1"G�*�%����{��ԫ[g@Xa�@"���ȓ,̺��D)|�nQS�C2[�l���@0p�[\����C�"�ĭ�ȓ?qP|Ӄ�R!�bՓE
ʄc[��ȓ�zX9�$�$Ϙ�À�87L�ȓm�|H`WA��^zDy;�k�h0p���Z��9��� x�Z�I�HU=��b�<1`Ο��Q����r�HB�BCC�<� ���� K�4����4�4��"O	��)�=q��XJ�(��;�lU�r"O�B���^p���ѐpy4�R�"OT����?E������Co�c�"O�ٓE+(6�.�󵫇�G^�%"O&���#e���c�뙶WE��Y�"O,�᷂T*Z��CQ��}TC"O�!�� �1�n� ���,Lm��"O�X��jE�f���pPş2%Cn��"O�51��o�HX���2nN��2u"O>e����2A������]��X1�'�:XY��S�	9I.tW<���'��@#�e�5h^�Bć��_?���'/��	F�P�i��%�ˌS�`���'E��B4�յG F�Eh�;�HI�'��4�U�9lذ�4	�!w���
�'� v�B"z78y����� _n̡�'� �f!�+l6l��c�ʎ"�nx{�'��8�jQ}��mH̃!䢔

�'^�RJ d�$!�.�On�Y�
�'��9�C���:�,�X�B��N�	
�'O����X�B-�XB`_�C��ԣ	�'n�`���ϋk� ���X90G:�s	�'��{`�%fPݡ4�ȰUE��H
�'xբ�̋�9ذx�k�T �8
�'hC�кj8��3n��Dy8`
�'��pk�!p6�� �Ͷ8=:4

�'X��3��65QΌ8��U5+gR a	�'���V�M�#�fx�d�J�'����'�Y�5D�>P�쬳���/�.���'�bA��V݄��ML�x6>���'r(q�cR�J �|��G"n2���'�T`Pt%9!�~p�A��m%;�'�z\��Gԗw9� ���x��Ua	�'�F���ʑ?�����D�6k�$4��'V� ��Q�|`RfK�]��B�'�s�[`����f���S��*�'��P�Af���d�����z���X�'��� S?J��x9�CT�;�0Z�'���	LS�l�`�-�%�m�	�':(��Iٻl���l]�5�1x�'5R<���ޑ1�<E�+J.H0Ś�'�@��� ��1�3{8���'����K��P�7@V�//^�2�'6�fkΞ_� Q���~��=��'~��%м�z��u�"�'�@��$gH���r�gI��	�'��5�cA�y�
8�랛j� -;�'����u��$(�m�q�N[��l!�'����� O#s���
��ԖDjN�s�'�5�
J� 9ys�jR:B4,iJ�'ܴ��R��]��홤.�9A�I��'�p-�1��4?Q�(�éN}U�4��'�P��p�ґ��"�	�t��D��'�JE1�	��w	�,�Wk�~���';� 0rEņb�� �b@D^�Q�'�8d(��A H�b�GN�ZG^�' �J� G!R;�a_�S�L���'F*�;S���g� uA_2vhd��'G�e��Ζ8������ o���"�'�v��eg��8����	oږ���'�V��e�ǉ��*� �jf��'� h2��cr�(F��9ʮpB�'��	�j�I�@L@wf�*�L�xM<q�S�? H��#f[�%��1�		=а�t"O
i�e�աfb:	FR&^<q�"O�貆���Tx��0%Or.���"O\T����%n�T�����$�a"O*d�b,`�ѱ`NbѨX@D�i,���=	�ԓE�[�� H�@�γJ%!�T#5H�Ѧ��6��AH���7Ng!�$�1ҭ镄T�+�H��o��_!�䖔G��bs\�)�.��m�!��f4����u*����<[�!�DЊ-1bh�� 	뷦�)�!�dr�Xp[CG�(Г��Ȯ/!���(00�C�	e�C�xd�"O��*�Ę�H�������c��t@"OT,jt��3n���"��	6:��c"O�0ۓ���!�.|z��q����y�HɄ�~�j�π�0�<PnL�y"HO�(5�$�bm9%�<,�
ޣ�yb$�6KMZ��R�  Et�qV"K��yR�Λ_�B ��+L��	����Py�H:��f&Íi���2��~�<�C�L��ܡ���NYҥ�E��V�<!��Ńx��)so�4�t���+H�<1U�Ǡk�Nl�F r��_D�<�$*���l#��ofn���Ug�<���&X��'KFEMR�Rf�<��- wK<���V�i0�F]�<��!G>\�HT��i ��G��V�<Y�*A�%�@X	
Q\�`�Ā�Q�<y3�NZN�IqO	�,X��{��w�<��)���J�</>ХB�O�(�y.�$}��R�H�&5(\���!�yK]'_3Fd�GO�pެE�%P��y�;��$���5a��3��/�yB�Uj�h��b��W �}���6�y��())d	��o ?��ؙ�D��yr��$��m��X?:��l���ߪ�y��
���Q�P$�mjT��FF�y�o_�v��ib(�(v��$e�&�y"`[�h��Z�'	���cT���y"&@*g��@A�W�0)6��ƈS��y"��,]��B� �-{�$@�D��y"W��0��%�%+J���]��yb`Dw�"��@��'�E�W.ˊ�y�f������E�&j;D�  ��ybƀ�l65���۬-zȨcF�Y>�yR�'nvp���Jyz
��`BM��y�@L�_����%��j(�P@b��y��U%x5��M�@�����y��~&`�����,L�x[�e��y�˝ ��4� G��U=�|b�"�.�y2�^�}�"��	NZT��#�;�yA�L�l*�
/y
�Xc'�X6�y�ƚ8r �R�L=W��G�Z��O���D�z¼I�T���Ro����N�<!�D�e?�1� e^2$��*�̏ !���  ����Ǆ��DZ��ѕ�.E!�D�h�*�����4|ђ�&�
j!�đlݰ �pƆ>V��З$�5a!��3E�%I�E��}Y*�*4��raxb�	%Aޱ�����΀X��J�x@�� R*�CWRL��	�% ��LH��m��[��S��\Lb0��Vx���.o,�[���8��s��$$ۜ)��S�? d�8��%W�����DV1ru�!�F"O�ej槏�|YL���(=L���"O^�)g���oah�B�Q�I�"O$��c���.���t@�<��L��"O�1��^ff}����Z�x5ib"O`)��Η�/>��⋄��\��"O,t(r�I/���+ĐM�z��S"OX!�`��;J��*�iF�\S���"O��C���Hi�!�E�E�z�)"O��*nI�G��b�$U�|	�s"O�}��H�v\�w�]
���"Ol$iC�V��1�B�Ӣ]�j�б"O$tx�B+Xṷ�����j'�h:�"O�|���A�L~�rT���'nnu�@"O6�i¡p䈠҇�=h@�v"OR�˧��z֬�bGO��M+T"OX�i��PҮ%#�&�T�H4 "O<��b˞�C2p��@ȸ��j�"O�G��^ �%�`bC<[@�!
�"O����Ì,J�q���;�.5�"O��3G_�z�P�x�j���r,�F"O�S���'|�Z��� ~���ۡ"Ot���ߞQ�$���R�Z��1x�"O��ʲ-'$r��ٲ2�*�&"O�iQ�P�_w��� �H����;�"O���4H՜U�J��K�-�4��"Od��p̘�$s�%�֬��>Ƹ\c�"OB��_����W �q"O�� ���^���ЧسBh�3"OH̺���1� ���U�K�8""O,����V��@��	:���"OVk�M�ZfH�f�4,l�T"O0��P�%C�|iC�P�BP��"O�E�RJ; �⤲���.h5F��c"O�e�w��$lPjq �@ѝZ�e��"OBMp'�P	
V@@a��,b��"O�`�R�M(Y��y�B��2*�M`�"O�Y�ÊG #���3�gO�	�8Xw"O�꠯T5|�\�����*D��}��"O���*ɲ��tY��Ϻ!ό8�3"O��)�嘄=��Kq�B�r�!��"O�0{��{�ޱ�Q��D$,r"OHl�N�B�tQ��΋%0h[#"O�͈֫�9y�Q��K��8�"O�� 'D�(IdBX.:,��"OZ<)Wa�&�b�^�s���r"O�p1$�Z9j�����i� M�Up�"O�`p`욉�v�����a��E#�"O�P�׍�%��t�4N�py��"Oh�S"� k>��`H4	�2-QD"O|��D9Ωa��\7^�^�e"Ox����9?0��j�F��̙R�"O�5He��PaM�V!F,(�"OLQ���Ӣs�����.
�S���5"O����j�Hb���1�\�y�B9�%"O�H#v
�k^&Da�m�8N��t�6"O~a@�-D� A��Ƣb��:�"O�1��¿�rU�6'Y��:ȣ$"O�X���v���ac�Y!�J8��"O�I��^�Pv�`w�֦	8��sr"O�x��)�<�v�@�Q�T@"O�����υh`�(�)Zz�b�0�"OLa����?����Hńo�.�
E"O���V��G�ac���7m�\���"O� �٢U G�q|��0��{���ä"O������,�����!;����"O���� .���Yp0���"O���a��92Lf����2j,`��"O,��6�Q� �4	�%�[�DT�}��"ON�p��K�&�Z�#��ϙ@>z0q�"O�X��I=s3܍gP�� 9kR"O@d�W�Ȍ@C�Q{�Ԏ
zP]��"O���K܂X¦�U�����˧"O�	jqƄ�Xȸ� �͐-����"Ov\�R�. p�S�/�~��0�"Ox�R5H�Ry�.[
O��]a�"O�9Rp鋃���S�ʂ�0H@"O�|�`� �X��y�NܓA�x���"O�q�wJ�"I�fE`4kZ�H��5("O~�R&���B���j_�O�$`"OX�r3�H{��1T+�d��M�$"O�ȩv��3Nt�5)���`"OPy�@AQ�$=V�s$�T�L�j��2"O�EP��
3��Q�2�A�;�����"O���p/I(VH�E�n�8�y�"O��{�1C�R��B�_�"�C�"O��Z�e��Qe48YF��K�J$�"O��˄�؛6��� ��>C�hE�e"Oh�9�	E\�=�cڧ#���Є"O���A���S@�[� ���q"O"�95	�g��K��O}�R��A"OB��&��-�"��J�?��H"O������#@ND
ō��f���`"O�]�"@S�+V�i��/�Z`��"O�A��`��l�ʰҲ��#2�f�jt"O�Qkw,�T�"qуO�i��e9�"O�t�ǉ� �ZM���]'�hDrC"O^��p"�ꪑ��h8q
�"ON8����x�������DP"O���􁍱�\��t�L$e�8�"O8ͳpJ͕#�q{�-��[6x�"O�]Ӏ��;e\r��فM���@q"O���f�>`�����훢N�BU��"Oй�p�ځ[	L�P6l�)*J%��"Ok�(K�.D�y�K3�L���"O|��j���ф�S�B����"O����87��)P�چT�$�S"O8| �$�n��M���R�b1�,qF"O<	�t�\h�l��aF
�,,h�&"O���C��F�~�2vD��'qp[�"OE�f�)x��a�`��W��E"O��K�+C��T���h@�'LRX��"O��Z�kX��2y�&�L�:h�"O�@��	��*�Ӂ��?B6��"O�+��T��ܸ�Ɛ�o׀�F"OڽJF����ڦ'�6M���!"O��WCT4/�8]�T͛�~��\��"Ot��bϋ`0԰���ݙe��d�"O$�c�J=ohbzB �7Z\,��"O�4��Ə\� ���8<T�taW"O�,�2�Øq��<�c-U! It��$"O`݂S�ӽ{Њ%�4�!w@�X
"OX�8eĹ䴨8bm��E2|]�"O�mw着oB��)ǋ��?2�5�p"O�Yt�VkD��
������"O�с�@Y�?vm�r	W$�ę��"O�l� *�)��;���*ڴcD"Oz��5��c&�
�$��j��+7"O� �I��~H�I�E��wQ���"OP�(��n�lR��ՂW0�ēf"O����+'\Tm���I2~%�@�"O1hE  �u��Ra�&<���#"O���a�^�a��ѩ�L3e;�ma�"O�����́9���K��P@J̚�"Of��!�S�$����s��>9���B"OE�a%Lg*R@b��cbQʧ"O�HŠ�xV����a0-d��C"O��PLT�yT�X{qK���$��"OH sb�5�4d��IG�'1��(s"O*��,�V�
(�d� 9���$"O|� �m *S?��D�_>�@�� "Ol�   #&,��k7&Z1ఱ�"OB�c2�Ym7�(�%2D�,S"O�e��ߗ��%��d�/��TIa"O��%.�̵�D�
�V�^�I�"O�P[B�A�V��I&%�7|b����"O�!!�/�?1{�m�s�N�&^��;D"O�\{�/A=3r\A��J]�IM�l� "Oiʃ�׊G�ʼؤI��I��0"O^A��ؼ~X@�Rt	���2&"O�ȳD�	&9v`�	�+=`���"O:�prj��J$>u*�(�#bJ,�"O�\����=Zph���L�>�@Y�'"Of:�R��8+d㔰1�PQ�"O4�y���H�ݨ��C#@�)jF"ON�H@�ЦL�9��ϱG�f]��"O��OŸa:1:#�^ �\<Q�"OZ�s%��'D�KC��$^e����"O�p��c�)����^H��8�"Oz�Q�������&�R�h�p�"O w�L�>hFDZ�vm��"O�8����:Ҝ�d�@t��<��"O����n�: ��W��?o���$"O�(1A"Edrt`�@��p�&�+v"O�M�pH��/݈�� `S"h�=�"O6�	�I#*]���P����v��0"Oh�B�� W��t2g�,[xlL"�"O~�@�(ߗ_x�@Ӭ�G���"O����B!�Y����=*fD�Xa"Od��a�Z�[ �y�($,��*"O��D�U���l��@3t�PU��"O,PB3�Љf��@/��7�^��5"O$qSA��"��� N��#�����"O�y���h<2���gĶ�b"O�L�.ß>v�e����lq^-(6"Oh1�/��V��a�f%P�h\v�� "O��#$ƞ&�-a��% S(9q"O� ��/@�/�d)IF�h*�*�"O�E:�×�p�r7�����*�"O�u@��QBJu#`��
�6S3"O9r�AZ+m��kADXFZ��32"O,q�2h��4�A���Q��)"O<q�f$�,L�� K��� G>䒡"O4�p���5�b�'Lڞ=0$��"O���
7E4	�k],=2�S"O�h�lߦA��zӠ;(��3"O�+⣑5)f��J��?z=�"O�]Y��&�"M�(W;o�.9�a"Ot$�aԔCB��(Щ��Y�"O0�0�,]�Y�v	�iЋ�+���:O���Ī��g`����//,�. �7"O>4�D�Q ?"�Sf�#��ȳ "O� �i��L�� ]Z����4�o"O�L��!� h�QU(	9x*��A"O��2vLDʝ�n�,����"OT�8 �B�K�|�yR͎�F���{�"O�x��hZY���bT�8��=�G*O����%2!>XB���64 �5R�'���fA�L��aCR(��Zc�L)�'GU�A�v��)h�"_.)����'Q���2��y|^���_���@��'���3�ݶ4垙J��5?����'/����/A%�t1���s��:�'��ˠjǲ,����	�}T��k�'�`���hܬ b|��u)�+�tЋ�'Hx
�$R�n>�{�N�F9��'9bU�2MS�Q��5�n�������'3���GI�,rR�X�V�����'��$:�ʏNn19�Im����
�''�x���9J���裏��l�Zu)
�'�(�9�`K�P��y�k��p|Q
�'e$cTHɮr9H`�w�"eŶ)�'�ZUv�Ѽ\܄�@�m��A��'W|�Z�/C�8��Q����9`$���'���3���==H�#�]�8�6�!�'��JĂĢxY�k���+����	�'Sv�y@�'p��`�u�(q�x��'+NY�B%�z&N�iV�G�L���H�'��Z�mב]��1�m�1<��j�'ľ�SSS.�\��A�%��k
�'m:��4���-o�!�����X
�'�$�X!9&�!��ȩ�A
�'B��"�G#%�JQ"��N T��	�'�2`��O[�<��x�V����R�	�'�<�&�>s���P���2]��'�J�C&j�;3��Q��銣�Y��'�����4?��!k�,���T��'Y��8��)"���#B{�N���'�q�Jԭ+�EA#��d����'HP�����Dȹro��X����'%�;2�ƶ\�Y*gN�z<���
�'ֲ-e�����-Yvl<x���`�'��`� U�&�Є����� {���'d�!�� �
�}J�	�,a�
L+�'�@��'�Q�p��U5�ڈ*�����'��4�"�ԙ"����S�T�ej�`�'�8�r��3;E���2(���'N����,J���)�nB�u� ���'��hY��Z��8�F教t�R�c�'7��p'm�8i"=	�,P�tvF���'�6)i��u'��6.�|E�-+�'���8�P�?�Jab6G���q�'��e�]l�j�	��֠���'����쉲b<��J�.�� f=��'_f��PP���Р�x:��3�'����)�C��=b𡖂C�J��'Ƒhf툎pg�u2q�S�4"0!z�''b�!��M�Yy�m�P!��uK��B�'�엺K�0�у�R /jP3&e@v�<�L�; �xy!K���}XՃo�<1�$ۢ_0��[(x4����n�u�<����@q�͸�
G�(�@�ox��'a�Q�1�"k�@�y0K�񆁈�'����������BLݜbxa��'���c+�:e��Q��N�@��
�'�D�#F�ͤVi yӢ�(`T�
��� �q��� �0P��C(3��Ȳ�"Oԑ2e'�d�*Y8B`�n��P�0"O���R�%��R�_'��&"Op`kpK�#;�T9D�_"��<�u��b�ORe@WÃ1i$iz�bZ�h�.�'P�(A��K8��E���e?\E��'Ĭ�IFLOh�ȼJ�B �dn>�:
�'G6hQ�'�΋p4�@�fχ�y�9F�DL1��F�l!M"FK� �y���1a�p���d(  �d��y�C�F�#�#��ؠ����y"��<.I����d}At. �y��߻��8��	
�J]�uB�J��y���][^��$���%qGĴ�yBJ��J%��F �]�CbE/�yr�WeL�Ih� ��h!���y��C<GnL��mS�7�}@��I��>��O0�k���4f��W�<)d
��"O�t�KW�`)���F$��"Of� �!
88l�3�����ɐ"Od�	D�|S0Q!�<K�`�"OR��q�ǧ��[��1_D��q"O@�2��ώ�lH����#��]zR"O~0aE�L\6�[  ��"5�'��7O� R1億LS�I��!Q��]j�"OP�c��X�dm"QFW�]�*0��"O�ų�듐x���ڱ�:;u�@��"O�V�Gala�c
y�tX(e"OB�R��A��&��$+d"Od`�dg$l4=B��)%QP-��"Ol]Ò��
��Щ�H8��"O�h5��-"���`&�0B"O���Q�FA�9��̄3ʴ�g"O���O��n�+E�$"�
 �+\�<q��t�<�R�)Km���s�o�<��D�K�āmA�9ܔ�׌A�<�`�>��P��X�Q�Xz&$�x�<)!ϫ^��S � �@I4��n�<�oC�Hh�x� ��Ff��u�<�gA�	cj�J��Z�e����q�<G&�""~� �7��|)� j�Nt�<	4e��p^��9���:�2m�T%m�<5H�+~&=���od�ȂJ�i�<�d��'T9
У���`-0�+Yh�<� L�vruIG,{4�:q�g�<A�FM`��ĥ�;d� �O㟐��[��u�W�
2�ri		��L���0�l˵/z2|abG�y�A�ȓz���ec�b�u�u�MS�t����$)��H#���2��:(��������*���x����H&��ȓ��U�_x�פ���J������Rk�زt�w+��eY-��p�����N3q�!�eo^�#y�x�ȓw܋7+�,\{G�Aw�x��ȓP�	#`ɜGĐ	;g�k��ȓX�Ɛ{���3Ҙ|���ev�q��e�2ա����"�x��djO 9�t��ȓhq��׊A�__~���������ȓ�
�+ŋ	Z��%@��S8�!��QZ� g�H�O�|�[��_�a�نȓt,M�dD�>�������.v��ІȓrKV���2/DV�8��O�3E���ȓ%�:@c4�2�|��.�bS���S�? ZAH#O3,Ty9�HG�lx&a��"OD*�)b�p�)�iK��j�"On5A�>���P���/J-�%��"O0ě����p�	 �_�>�Vx2r"O`XaU�����L�a�qs�"O�`���2|��s�Q��~h��"Oʱ�p���G�<)	r�� +����"OD�͞�l�!%lR�4��I+q"O����Q !(d9�M=�]�'"O�d���clBl��h��Y��١���2LOU�� u���ԅ�60�v���"O��Em �$��5�Y%J���q�<Y�T%wL�IDj7
/���S�<1�,�Y�|�V��6mN̠��G]X�<�`ぽZ�TpC�M����aI�'P�<����
]�l�y���Nc�i	4��O�<��h�?��s�c��<�䙻���L�<q7�H*�$��E�䴙�L�<��,Y#`f�Yt#�`�*����K�<I��>��p�����"}(�cUn�<��e�P�:�P���5~V�a�f�<yVV
U�1r�Բ00��6�d�<�W��:�6�w�y�p�qf�^�<	�J,/��j�J\bZ=(c(Qa�IB����ʹ=�Z��e��.,ʭӢB/D���@+�v�yB�D&F�����.4��PԎ�7n�$xa��'A\�рX�p�D����h�Hps�וN�ج�W!6D���B˛�<��8kW!	�0&��Y�5D���R/�(@�kZ���9	�`5D�$+�I԰i>��ƌ�
f�ۧ� D�(���I��xI�M����R"� D����EV�'v"ĪQ�`���!m=D���W�D�S>���a��B��!�K;��.�Od�ʱDC�Bu�����I�(�p�y�"O�QRQ��:t��|(v�k�dZ`"O6|P�Q���+�P�"O�E �F5v���*�)�(m���"O�����I~�a�G�W��"O��Ôb�\j��dˢ��s!"O�E l��Y]��@a@ ]� 3*Or`��4Gy@��>y3p��'�l�9u�+��i�T�B�< �'/"��o��$��;�	�	��AQ�'?`u��8�D���NQ�A����hO?A8�>B��	j�e��<�jukCF\E�<�Sm֢S����(I�J�ȑ�D�<aP�I�LRd�#�KU.6��UP�O�X�<y@!��>e��ʈ�V�BP@FVT�<���ʪ/N�pjJ�[{x��R�<�u�Ϻ2�NŘ��̀G���
S�<y�	�D���b"ҹS�d���J�<�e �^5��@�ضYJ!�ч[F�<�ԡ��hjb�ȶ �,M)R,�E�<I�^�$BnE9��^�k�L�p���g�'��'�q��,�$�%[7~����!�6���'J�����#w����@O�/���b�'�,���䂽*	a@�)�Ց�'8(��	'wޞ	8�@�&=~��'����g�Ǽ �*z�<���h�'%dE!P�$c���E >yq��Z�'�.�{!�X%69^,re$ȐjK�͊���)�q$�5rp.Q��̙f�<}�D���s���c��C�0���|��ц�S�? �5�GF� 	���4rK6�;p"OڥPqgڪ7?�a`���������d5LO��ȐEۖ(��yG�ɨ]�B���"O����4�Ha����u�"O�}@�@'���ʑ0p���Iڟ��Iş���3LG�X����g��3y���ȓ&cpP��
�3�t=趩�g�4݄�Jn�E�ց�.~H�����_�3߀���K������d\��B��7k�f �� d�����2w�<ٸ��2��u�ȓ�&�u�Pya����k ̤��\W�E����ۃ�Î$���"W&�d(�Sܧ��\�#�c��T�լ�W��؄�D^�2юN�[ydl d��_�2�ȓUV�aه�6SSl�'��0�KE�<�F&�7	uTi[Td�"����eX�<AФRX1^�y��yEF\S�<Q a�=~��$�5䏓J�DA��g�<� �Ol�J��O7L���z�
BN�<iV�ƭ-.I�f\� �,����J�<�G�7�N=�$���$��E�<��E�?��$�&N�.M`H�&C@�<�v��	X*�1W�Nq	���[�!�$�M�<s3�c���HÇѸ^�!�$ �"�t%�"�Щo>�3�LP�,�!���$T�U�.S�h �m"�� �R!��
;,��a#��K70�鴠�6O!�˺fh������4%^�ڢ`��M3!���_~��K�F����Y'!���!^��b�W"I^���wo��rў����oa�H��fC�#��<'�Rn��B�I"
��D���]�Q6�Ց��g�B䉈;l@���#. ���{��S��C�	�l�vMӃ�>N��qRG䟳1j�C�I�.����a ������ע�C�	�NU|q����@F���cVf�jC�	6�r�
0G��J�A�+%
DC�d��@&Lٽ0mn�"X1a�&C�	�0bd(!f͑d�(9y�i���B�I9:h`��E%I�-�"]���GҚ�?���I��A�l��D�r������g�!���u$Z���Wo��0��Ϣ ,!��~�Ҕ؀/ �y��i��!�$�S�.�{��,s\@�k�"�Y!�$́+�v��G��<9��U�>�!�d��9�:�V�z*D�zsa��7w!�d5J��N-mr�j�m�ym!�$�;'�����7LZV���,�+.q!򄕘�,t�R�UJ4���ϣw\!�D�Ip�8�t%\�t+v���G:!���'C�&��奛�e��٥JL�N6�y�ቇ:9T��5f�WPj5ku��7� C䉹�����fÃq�T��	���B�	�sf٫���9i�*EKN��l��B�ɷ��zpb\�;�
qs`	S1vJ�B�	^��%`��V�*L�4�qm˦>��B�	:7a�4 ���>�0	��H�c>VC�Y�
���d+�m�F���l,�C�IyƄ15��Ey\$ڴ�J.!��B䉤eLHSd曟Dcb`�lt��B�6[G��r�׷6F8�bƟMC�B�	�H�J�8��J��$�q�����4C�	\�Tx#0���R��	{��N{L8C�I#R��-�4*���)��X<v:C�)� j�X�,�<@=���O
��=��V��D{��i�Bq�ꊱVC��#�V4T!�	�2�P%N!G/&A�W���k�!��;X�z��@�,n�,����67�!�d�^/p�"A�+ZN|P�"!8�!�S]��;��W7X"��8��;�!��9;���a�Ҡ"wJp�n��x!�Y	��[�H'
]F1b�� m�B6O��`	�$���b����� c"O�d��*��ou�\���0��T��"O�A!'��&�� c�#
_ ��B�'?O.�pነ	kȘ���
�	i�}�P"O�Skܬlg"|觯ɰV^�D""O�Ap�
���A��k����p["O��9c�@3_ p䛃�+fr����'1�Ƀ:浸�c�<*D:D��ƞ��!�5�&$1&���(ȪL�l�N�!�dS�&�ܛ�'�Q�ɩiF)I�џ D��d�*(�p�R�ڡ"����.F��yBƍ..z¥Gٙ��(�F��y���x�\Y����
V���8�y�#�Υ�QAX�v5������y"�}z���#�-��P[i��䓥hOq����A�%���a$�z2��ؔ"Oݑ!	�v`V�ː,��+`��' �Y�HfD��H�&h&r�ӗ�A�P�!��"~��q�g �wB�x�.�B�!�D��[Ê4�F(���D��%;�!�DA&Vt\�4�)T*�����fi!��ţN��@q��ȫlJpXæN��!��B�i:�%��t��H�%O�{�!�d�$�L�� �Xo
 3�ډ
�!�?�p�f�ʍ8�h���!�䈿g]�b�bC�M�0�aF��!��<-ҐtP0I��N����6�!�Қy�.�ڳ��"	��jB⌲�!�d��Yi�dy��L���X1B��r�!򄊇T�lD�Ŧ9tV�-����>
�!�ƏP�μ��D;h(��SH�!��0W��)� ��a��-H2HZ�WX!��3HI�l�@=b����^%fH!�D�gz���s�"*����a�~-!��	n|�bL7m�����_�OB��<�v���I�i �CZ�'Q ��,�D�<��AT��E�Jg�	u��Fh<i�h�[������*p������#�y2���VQ��R%��l�~�+��8�yb��l�`���I�8e&Sk�?�y���*�V��r`Јc��5�m��y�����	6#2%����.��=I�y�G�:qF\�Ӱ�@�'a�-�dHM��yb �74z@�T�	��n��s@���y���h.i����gR�P��y2G8t1�]Ӈ@�#u��d���ť�y�U���ab�b�(g&�a��c���y�� 8�(��t��Qx9�����yB��I*�M�HX  ��]#�L�'�yb
k4E��)�~�rS���y��3 �@�ǌZ�ݒ�.��=y�y"h��C}����>:Md�=��'2ў��'�H cf �����Ɗrެi�'Dƨs����4����k	�Z�@l��'���ȇ��0e~���O
5ZېQ�'��$�&�ҘNp�2�+��J#�p3��� :�0��4`�>�
@?*4��G"OR�Z��ڝp=T�@�"K4L+�m�V"O�(��J�n۔8�#.���|���|��'���B�LC��r�Z< Y0Ma�*ݢS}!�B"-m\)D�bX�E�FiL!�Ē�f�T0�A�6;H��P��̸F!�$�>iy�`�Q\(Ɲ����/�!�-{��uc&"F�L���3q#��N���<O������(/͂������Z�ӕ"O&)�p��t`�@p�OD4��}�q"O�zp!��+�T��UOO8��p�"OD����9G�:8�4%�"O�L�R�X:��D�U��4!�5"O�e#V�Ֆw�}#���"�
�s�"O�ݺ��Ԇ]oݻ�� �/���v"O��MT�xv� ��"��ԁ�"O� y�jM+Y�8TB�Kgl�8�"Ol}���	 ^:�`�;6|\�"Of�"%��6G���!�/L�q���b"O�x��._;�6�cũ��`� �)�"O�ɻ��^�[�ЬpW�Ē(�8is#�D>YSHLzFYw�T�=X��G"D�������}%4p� �$#�=�$�O^��>�8v�0�~���T/}��[�)D��c���f���'E�2iɔ��`H'D�,�&Y&*%`Q��R i@�a6�)D�h*SdV�X6 0)*�O)N,�1f*D� � j�#g���៵8�j�z��&D�XHЫݮ� �q����-�8�H�l(ړ�0<��b8Z�!��4O(ȡ3v�P�'Fa����?��HPF�&_Wΰ
7E���y�HW�
�rl�"���B�'Ȧ�y��ԍ ��M�a �8�&��V�[��y2GǇaf��B6$�3Č����yrC�)��E��-��q��A��y2!? ����R� ��Q�@ �hO���D>I`2�a���3�V�H�!Ǯ6�	I���r�RT5��
�L]�'���	&�Oj�9�I u��b

�r�D2a4B�ɧ!��sTE!D�l��"\73��B�	!F�@�薩�<F�+����dC�� И���V}���U��Jb�C��</R�q���&R� ���A1ZC�Ʉ ��h��ȏ�`������+���=���^�4)ˎB7�$cĂ#Z�<؇ȓ-�@�͍�+�Ό W���7�
-�ȓuܽh X�2�>�������:t��%>�aa˂����@	3:d��u��0�ȍ��Z��K	;;�e��o� 5�$�R�V��hF0 |8�"�'�����-�� ~<��A����'��mBB@�0������}Y0 3�'&�`A��#��K��ٶx��y:�'�d�e�XU$$[�ʜ����',bU�
I$u<( HY���g��V�<�ӆ��$8@�=ƦqKv(�P�'?��v�@�wE؀+�'ΜL�֭B�'D�(+%�߂]��d �$��wr�u�&D�<��+,�d8����#k#D��� �&W����@�F�~�i�i5D�,ڷ
�q�x��e�����{O1D����'j�,E�W�ǔ��$�XHB�I�$&Ȩ�5'��[����`�ϒ(��B�5rZH�f���� �ϵn��B�)� x�b��A�
�u�G"O�p��-����Y�A�<�A��'?1OdY��F�R�e��i��Yr�"O��(� �9*)�jg�t�V@""O�l��晙C7,$X!#�/ eX1I�"OĈQ��4�H��#VoD�	��B�O2r�*P�J�E�$ݳ&�D�qR�'�ƥ�#d��f���s읈4|p��ϓ�Od}��LK�
϶h��,�)X�u9��|b�'��x�l�$��;��$SdN���'9����ꊼ'��Xr�H=\�1 �'�)#���B�
1b��ًY0�'R!�3�Hή��pF]!Ph�
�'��D�-
Qy��@�@�5\ ���$,�D&ZW��!A�<�򎁻!a^��W�}�I}�'�1O�d2� ��a�Z<KS[0Q��c�]��F��D,-���F�p"����	Cp}!�d�T�Qo�7��i�#I�s!�<C&jH[�W+&�]Aw�Gp!�<<�}���1��DQg��l!�$X�:�j@"���$P��Rh!��9#�jtjF��'+�8�@ٍ@O!��U�_ˤ��b�ݶg�,�VNҩ7k!�$����<�af��*j��n@�7!�$V�8��!dE���Kb�V�Z(!����p@�6t�(;��Cn!�X�u��5���-	x�F�PA��}2���RmI�j���:an'က!V
:D���PG��FD��q�ӂ
n���:D�0q�h��B���	��Դ+�DH7D��q&Ř�b�庁�ߤ#|��[��4D��*�bR����]\+��p!1D�� ��`�bI�/��;�d[��)D�T�[?t��"�^�6B@��:D����	�C��%�b��
ar���3D�P�6��Uh�T���֔|r22#�2D��c��҃�,��e��7
2�p;�,0D��:�cq��P32`�<X�\�9��-D���@C��f�Qf����B�*D���B:k�|��/_Q����(D� �cܟQj�pF�H]0b""%D����h(eb��ѐKE�G�\Ig"D�lh@C�$��X)�� ;�%0��O,�=E���Ϳg'|�Z���TR8a�� *��O����\�i$pB�-I��E30��(�!��
�w��93�F���Y0M�%�!�D�-r]:�x«
�>�Z�r��/k�!� �Z�1���͙^��z�l��*��'�ў�'�yb%���\ģ%��2Fs@�Su��%�y��þ���VMC=��ezeL���O�"~�D�@�=�=Z�i��Y@*8�'ɗp�<!r�ÏBk$u�����qE�R�<�_�ub Y[�
�&l��i�Re�t�<!�.�p� �p�� (�J��{�<��͊M�r��'"X�Fz  '��x�<p�ޖ��Ql�"	�g�t��Iq��|�qO����J�Y��Q@��#�OR�4h�"���@+ë���$�ȓ/�N`�ÌҟJ����B�1�a�ȓ]�}��y�̨�7�	�t��<BM��"ʰ����R�ZĄ�zb,8�U��-]��	�An�=_����b����?\m�)�u/]��X ��<�L��ve�**�����y��S�? ����P�r�y镈�4l�b"O6I30+>Ce���&�A D�yy�"O
���	p�Ѻ�̬dN����"OH|�Q%���Hg��lb��"O�y�$jںk�u�V�^te u:"O���%��|iָ��ʘ�f|V)P"OH0Ο
H҂d��ʕG]�)h�"O�%Ҳ�O	r2Rm;�fъP���"OI0皐~�Xc��>FnmY6"O�a ֡�~�ℊU���36 1D"O�e0��#/�~0#��8Ұe��"O0!`Gf�#&�b�֧e�@[�"Ov|���[�b!�� �"��@��"O��YEK�=��k�"�6O(ŋ��'kqO���)����QJ1 &	v�+)OD�=E����B����G���X�7�R4�y"�� ez]���,|��\i hU��yb�X�p&�S��l..u"pd��y����>BI�e�D dŐu�� �y��Zʜ� sˤ ��N�y"��?�"0A��7qs��a3�܍�?���.�?��6���r�I�@�25��a���$�<���d��@qf���&0@��dq!�!e��|�iV�&,T���4~<!򄋎F����02&.PJ���0&!�dȍm���o�Z;D��D��a!�$X�!�X�v-��-/B	 $!\�O�!��L� �!��/[-֝���I��'5ў�>�h�\Wʖ1�҅Nn(*�[�.D��Y��)&���$�Xl8u�h2D�\j#]�!C�|a�%O0�ᓈ.D�|�� &/������1y���a�'D�h;��.x�$D+q+ڑ{H�x�V*$D�<z���!�l@�@%�;o`�\�$$<O "<i��&w\)Z'%׮s��hgG�F�	~���Oe��c�;p L�5�����<�'ʠ�pՄTO������� �'�r���։f�{4k@� �T���'�B�8œ�Bh���C��'��Z�'8�u+F�<IJ.�Q�F�Q�FPs�'�n%A(بGNV(!W�y4)t�<�C�� r��BJ>n8x�Ĉ�s���0=�,�ؑB�!�&Q!q%�v�<�f�#{&�yk�kӅxHU�!�Yt�<a� R�.��1�ڂ&0
���o�<�b��?�^DX��Z?Nr�(#g�D�<�D�2�6���վQC��ҕ�YY�<�f��%�r��tAA��K�Jh<�X
G� ����;ls��w
*��$�<y��0|�߭-��BC�N
D�\U3S
�ix��Gxb&�<2�{!+�bL��Bv�\(�yi�6��J!�d����5�^��y⨞�q@�iY$E�NE��*�'��ykF�,�Ҁp���?��2�Γ�yR�*�#�%S�B_hxBÍY�yB��E���I�ś�A ����DJ��y��s���35�$�4����OP�=�'�^D����N�䚃�6�^���	
�T�E85�� ����g�L���O��\��F��t�H��Pi���X�ȓCdU�4�Y�s� p����*s(هȓv�u2箌�@6&�JDN�=���g�J� Q��54����j6���I@<Ѵ��$>��d�wI���4�0NEi�<� ��D�P"-�d�)��ע|>u"O���wkZ�:mE{fo�k vĻ�"O�*�IR�Z;�Z� G�+-�""O@躆o1�ԅ�&�U�*��p"OΈPM�}��h���R�'�v��"O�� ��܂z��]0��A?K߈�sF"O��[f�I�W�xc� ?m>���F"O�<�Z=]x�!6(2u)�P�E"O���f���B�)%ҥR�"OHD��zb�Q���0��}��"O��Ѝ�8qp
�󢦉j���1f"Oh"�O"i��a��=��I�1"O����%�:T+�x����w���� "Oq�\ rP���5a���P"O�2�.�y��l��/�������"O�}X�ED ��Ċ�.��@�(�@�"O��hGm@�R\J�M�-T�ʁ�"O��JR����"��n	���0r"O@���H1iRPM�,�#�"O %��X�5�8=�a��@$��"O��Q�sw| ���Z&5����"O��r"�S0J\rċ��n��5c"OfdR�F�)i�vi�5(��l��<�#"OZ�R(ټ?��mۤ�M!P��a2"O��Xg�(:߬y���4��в�"O�\;!��SE]��%2bآ��"O�uz�C��E!�Ȓ1�a�~K1"Oh�d/-unXr��0�X�P�"O�BG�*#.(#��>u�hx��"O�M�q��?J8�y�o�,����"O��Q+�.���n��5s2u�"O�!�.S����m�wD�!�d�+3~�H1K!�6h���?�!�dY�!fth�e�"��DY�.Y5c�!�d'��Q�$Mߎ�b����!�D%2zę�d��=�B�@���K_!�G�K��xˠ蒋}�4L�΋�,!��̥"^�:�H�;v�e�Tb^3!�$�%��@�X�NH��󇀞#�!��S?4
B�Q'����	�!�$U� .m���S�4;޹��'̾�!�d�F��E�ͦHX�A�P퇲i!�d�#���r�LU [S��#g�2�!�DBC\R�p�M-����%r!��� �X���-^�!I8h��x!�$^�r[�d�ӭ�{=(���K�
$j!�d�KI�09C�S�e"��yC��b�!�$�~��q��ſJ:ъC� R�!��ZԤ�ˢ�W�%��dX��M�|!�ă�u �S�T��P'!��%!�ц% 6�dZQ���Ѥ&�!�DSrSf ��oZV�,YP�f�79!�2���8�m�%2�Q�ƉJ:!� R�����!Rɺ,��e�#w-!��11-trƏ>SS������w!�V�E�4*�jQ���x#�H�'5D���s��<�@��޹"�N���6D�4j��ߺI���I�:��X:F�0D��;��K�-�h0*�����"�"D��t�0̰�"���' ļu�!D���GNC;2��y:�bO�jh�@A��=D����W�1t��i˼)�ވ�:D�|�@�9 e��r ŻAA�M@�%:D�P��mR2j���C�4�����8D�� ����G1%�`���@�f��Q�""O�}����D�����	�4o�L2�"O�=�Q�Z8D���Y�/�@��S"Ot �5�a�D��a�H;9w�	�"O�����)f���"P�DenT��"O�mh2�\;(�,J��)*]��"O�ݛ���	� ��"BjTHR!"O l�WkW/(L�T���.i^�ɥ"O���ԸQ��`�ƀzS��)�"O�|�$��=�H{��B;~��R"O��r�\
�I�T��6ǔ��"O��yE�^�l��:Ua�9���"ORQ��H�	��u����z�"O�A�턀f�`�ԑ`J�P"O�lK���3P"%�?7�@�2�"OJ� �� �EPE@ z�S�"Ol,�"��-�&�т	�>Yƙ��"O؝���[zO��#���k����"OdA�/D���	b�<.�z���"O�T�e��}K��׽W�|�ks"O���#�]"��ԍD�"x��"O���t)!I<(	�@P�N�N�Xa"OH1B�ks�r���-$THpH��"O�X("͇�%��$�Ɓ]tބ� "O���$B�D��O#�>���"O�B�O�;���9ǌ�<]�Lk�"O�<(Ѩ��\Sl��6�L�7y���`"ONH!E�]����Y�끹���!"O���M�
-��
Y�md����"Ocf	%X$�ʦJ�6l<P��"Or�;%�ݔR�y��n�	�`"O�GEC�.��V(H4SV$<I�"Oԍ��(��ialT
QS�q�t"O�5`C��0�< k̙P���C"O|QX����z|����O��9w"O�Ԣp�L�G���KƤ!K�4�"OZM �'�{1`��6#�l�j"O�m)DO�к ɍ�dc�Q:c"O�YҒ�E$kl�2�#hP@p�&"O�)���Nؖԁ7�_:@�]� "O$Xz�
�]�.�c�OU&;P(�"c"O/<H4͂��->@X�@�K��!�D�pP<ű@���	(�aq���!��Q�j�����>=8�8�/�(SS!�䙜5��۶��Y�Ƞ\�Y�!���%�[�,�,�9����B|�'9�� �L����Żlݰ�'8��KҬE���%ϏV� �
�'��$��C�N69*w@Ҡ!4"7"O U�2�Gp�BIPu�5/6�� "O�|;wmF�>T^���*D6'+8� "OPis	�.!���$'
IC�Q&"O6y��Gΐn\�����F�T%��y"O�p�aHM!h��ǣY�7�9�E"O-y0	�+��Iql�p�s"O0��c��s�~%�eN̈{+zMzt"OD`�u���j�����{�6"OQ��)|� 8dB]}�]k�"Ozr���8��
�JD�p_�M�a"O�\�CN(W����ٌqX<��"O��֍٫{#���C�	|(��W"Od��`�\(<�e��	�z��q"O�u!�h'����ED�$
�R&"Ot�X�!L �hXAc9 �|� "O� ��4)U2Wp��b �S�,E���$"O|�6c�'lN:�� �  *�,��"O�|I�e�-�T\u"V#��`G"O@m�U)�lR,��f�n�M[�"O��z�τ&�1�)>^4 H""OB���Jvd�����'_fӇ"O6���K��e+j@�9u?
�at"Ođ�U΂X�~��E�U0>q�6"O:��G��8W:�{��B6���"O������B��d��7F��Kc"O�ի�fȀ)�d+�$V]�� v"O�*�*��B��j�	�_��mH$"O�p��.N /�.I`'�.q�){w"O�$��ЩX�nͩ4��39�ֹ b"O(rԯP�dte�T���D�j�"O��ʲ�R�[b ����&�J��W"O�M6_^�
2#S�|�n�jS"O�
d׎uv^Lc�Dĝ.�0�B�"O���#k���f` �K2����@"O6�05hF;'R����#8��uC"O���eFG�Em�9��R/.�Д�$"O��*햨+��:F+�:X��c"O��C�b�;�Z9j�����,�T"OJ����-nЀU0�A�WItyb"O&tĆ0z�������f"O`�BV*�3�f��G�*tF�*�"O��; �.;��#�FƼVQ���"OAIA5Ba��Rǚ#$>>Ez�"O�m0�C?Zt@�O�]�h�*"O�)Gg-f^J��s,�!\@��"O������
�RԒ�)Z-e�$�!"O�a`�)�(�������(k�5K�"O�5P��~�y�7���|��e�b"O�Tcb���"Z���隍n�t�R�"O�����E>^v�(��E#,��,��"O�u�6�ҏenqX�$;J���{�"O�	����s!v�KP�3�(=�"O�X�4�ع nҹ��/vu�I�s"O���
Zg2a�1!�DD��"O���Db�Fel�{��06}�g"OH�bē��\B���$�&iB"O�D#�)+`-�!�=;�x�b"O8��E-ܐ�4<�� ��V����"O�����){��m��n� xa�9�C"Ov]i��;{�uZ�h��1j�"O�ɀC(!c6��#N�%U�.�z�"O�0r�M�)>FBH+T�N�a�$\y�"ODD�S�NSP�L�I�e�l�Y��x"�i��b?ik�V�`�$Z�!HN�.G!�$ѣEq�S"����Nl5�Oj��$B�i�t��1�M8�2�[��%?!�$	xj&��@�(-��-��+4!���2��Pa ��y�qSO��r!!�DBzwz�۾�:�y��!���W�HRU�N܎xۇMS��!��	���s��f�
�I�D64�!��;A���p�"[>n�3'����Wx�P�B���X�
����¶d>�O��m�ƅ�Յ��$��D��x9����G��h�i�'*�n��#�O�&6(��Lږi`gO�(ex��;@څn$BՆ�=rҙ��jX/d��b��q����ȓ�\1��2M�
�	�E��M�*=�ȓW�V Abfٵ9%�U��`��;-��S�? tHE�P�YJx�R@i��O(V�w"O��+![�-�:}9s至CB�(�"O�	3����"��8�X�V��Y�T"O�@Tj��"��-��^4L=�mk�"O������2�Zh)��̀x3Hl@�"O� p��8WMdDmտu���G"OdY9'�|H8�k	� ��a"O&5�҃�������q� ��E"O2��s.�
Θ��`�P�7�B\�IJ�Q��'6�X�dB�.�@�ċȄd8<�ȓo?數�C�lnle�e��VX.$�ȓo�Cw���"��Q��>T5��&O^�	�=�N��Ꞑ|��9�ȓ3i�����>#b@��g�]��%���B≬q#P٘����~xi�&wbC�ɶزe�uHװv�PA��,2���0 5�����@�=YU��g�T��a�'h���l��h����T����x9�'����7��h��RW%~���T\���'�>E��'xʠ��K@1����F�X�^���'J�~��yB���$���݄q��ls'�.�HO��S�� sqd�-��$s��xqȜ�r��B��*l@U�v`O<,hQ�'��2(g���	1��'Q�?��BK:.�X  ��=tq�+LO��h� �(Q�TZ�bU�$��s�C)�d{Ӳ#<Y�y�J��,�j��c�-��$� .�yB%B�8��L�F�R��w��
�y�	� ��j1)u�����0<9����Gq�e� �?U�hԳ���
S'!��ܐ9�\ñ�F�!��#�BL	!��jG�ɠ�� 
�|���8�!�[�RZ�	 ��2\M���ׁt�d�L	D�'��Ց��B�dJ���7�̋���<��'#1��@��d�n���+e+��@`�"O�p�0��D�^���IɲuV�����in�I�<IٴHO�?7�G�a���4�J3&����p#�L!�D��cW���D��Pّ�b׹y�Q�����<;��m��!O�Fpr5#��B�	1x���``$�=+:��6dߢa����2�S�O��0�σ|����Fa�<ݎ��6"O:�k�G�r�����ʌ�40n��Q"O��v�T�cL��D�u�|����O��	R�$3�L<ͧV,�5#�59M:��$!�&���	Y?�T��(8+���cE^7cl�}!*O�$�<�hOq��D�7�F�=�T��6��i|����'^�~�$}��J�
d�P	�%B�MbY�<�
ߓx�ԭ#��n��@��.�Lm�D}��S�y�"4;(� A�:(:4�H�,4�B�	�a 0��W�v'J��F�"�xB��;T_*��@�=]����� ҂C�IY�i�u$\<7��R�!�RvC�I���Il�>�qR�d��_:�B�	,d�@`SQ2"q���C�_�{�b�LE{��tI�k\x g�B*�pt:'"֟�y�L�<B8Ę�GC(��$�&'���'�A��	�4{�;3�
fOn�h�i%)��,�S�O��&�P��d"�/ʁ��0r��ĺ�yB�D�HG�I@�JD�Q�����~"�=�Od#=���F�2PB�@� ~��YG�U8���I�8��'j�X�Y�N߉;!���2g(�D6�S�y�81@-�-ct:D����0*��yFy��j>��!خ-����/��C�Za!�#<D�|����,����g���%�pQ	#�8D����Y��:��f-T'�$�d9D�� T)��̒kL�`�	?<�L`4"O�JCa�=' ���e�S!H��X�"O��Q��� f�p�T�
�It��x�'�`��NK�T�Y�)Մ�A���?a�'��y�����*N��P(���	�'��){�VNتa �ϩ;�.5���d&��?%nڮ"���a7�T1*i"��p���U��B�/c,Z�Hr�
�$�X�b����"?�Ӫ/ڧ#> Җ�Z�}V��3 ��/"�Єȓ%M�U�p���(&���D�s��<	��퓋}��i���G�O����
T8B�	�f��D�BC��$B���F ��O��C�d�\i�F��$y��Mr�S������"?��O>�q�� z-ԅ�#��w��ĉ%"O2�;�KG�������V��}3��h�H�>�I>YE��oHp#s-��>�~�(��V8��Dz� L"FW�0��F��T�x��J0�y��'p� 0��X�P�K���O�=�O�� ����,8(eِAԴA�'��d����a&ԚŤ��2�}��'�����͔�y��ec`��� u��'�R�ib/C�|�����}'�=���.O~�X�9C�D�AP�-[�H�"OXH��/	q��b�,G�{��ʤ�i��$�"�X�dgN=S����ʟ�5.!�$�1V�]�&R7x?�EѧFԊ!�3���8��C�r8��ʶ��8�!��2R6���*�L!j���cU<�!�ȥotz�!��;	�T�68!�
��}�U� ��� 	sB�-+-!�+#ZD�II�g.�p@��v{B�ɕ]4"�� +�"K��T
D�[�����9}BE:
k�pc�݋���!gT�<�!�$�1:�ʢ.N�@4��P��gɡ�dٟ<��q'���]J=R"���y$��b��H�E�m��$��5�y]y>��
g�XL�fș�D�:�y".Ȇc#� �W�Tv.�u�#�yb#�*s�)Ѡ�NG�`r�	ƃ�yBǃ(k�9S`�ěB��h�g��y�@,D�!Γ
7A��ZD� �ybd�(!���!eO�~o\�B�f� �y������k���.~)�؋�.Ł�yBD"x Fa�1�M>�HU0cL��ybmSbA��hSl9����ǒ�y2���J`DU6/��"(��yR��#v���./����1#��y��	?��9vAޣ;Qx����	�y�"��������-,a���y�\�-�j���MU�*�4xw#�<�y2hT�CD
܃�MYX��+����ye͕Nz���Æ�|bl���E�y�I�N�l9��	�j�����y�1 ����A'[$�Y©���y�훈Ҭ��c�<�|5���-�y�kP�ʨ�ؔF�(eYа&I���y2�lQj��aHҗavl�Q�MM��y��W4&x�лGF�9Hn%�$Dɇ�y҇��مA:&�8,��e�XvA��'oJ�$�49��׫ )���K�'�V�9u��;?ˌ�@��Q�8��x�'�Xc�ʺJDa�����xJ�'��E9W� 9����٠OgZ�(�'��XۅJP$pl1�G�$H�@��� �ӦΗ�A��c��-{�r�"O��GY�7 �D�F@ɣ$"O�a92eد;�<��j��8(z��"O�a�3�C X�:���
-��Qrs�'�D�y��@E�6�A�Z\d�{��zA��O�3r��(�'��X�6@4s���أ�ռ!�pH8�'d�8�� �<)���%�1����'&,t1�[�I@HÔ�Ŭo$L��'�ƵB1�R�i-��sG�\�,1
�'�����ΨP�0E�B��+Pݐ�j�'K�H�d�8���{��P��hb
�'�x���RT ȑ�,KC���	�'v����G"d~��:�qK�&L��'&��� # ��p3@�^1]�6�z�'�b����%��}w@�bv��
�'�����[�d�h��3_��e�	�'�&�� �	�/,���siX�S��
�'�2�"P�J�M�i;3̀$�n�8
�'�&Ԙv�E,.+�L��`X�I
�'��I�$$�6f"�C�D��:�	�	�'T���#���M!Q#F0@���	�'I�m�u�ٯ)�I� ��+:�r)9	�',����U�>H��B`��;`)�'�����X�zR�Mq!ǀ;$�ف�'�$D	��Vyil� 2nT���'��p��H�N��AZSh	2;�vآ�'3��e	�LY��zS��jځ��'T�d؁@ң? |=Q�V�y��Xz�'�&%1$#�C�P�����qƱ(
�'����3_upt����F	n%F(��'���X"�D�:j���#)C�ȹ�'JVT�L�X�Vd(�`�)��\��'�j��$@>+D�98U���F���'��Ɂ�8^�x�*7�z!ΐ+�'��	P1(��\�#�	� �de�'����#c��~, �g�6��t��'f�}�tJE=b��B�3��9�'����'�Z���c!D �._�D�'uLH�V�f�\t8 e�.$�P�@�'�nH;W@	1�X�c3�F����p�'�R5+��V�'�H��q�ǆz�lb
�'��;�� ,n4�C����y��@�
�'Y��8���(���)�J˼|�y�
�'Ɏɚ�M�b��Y�g*��E"
�',��HA�mKr�*W�4|-�pY
�'V����_7�䉰�l��kV� H�'��@I�F�e�KFA�k�̤��'�$a�5.Tmv��e��/bA~���'?��íؒw:q��R4"4�h
�'z�D�')h��GP��!*�'	D�y�k�*qC�+�/WzސK�'	�a���˒� ��p�.m`�I�'M�8�H�q:F�{W�Ҥe�܁�'�TȠ�*R^0��ݗe���[�'В8s%"�7������?x��Z�'7r�j,\(�R����Ă2(t�'�6P�� �z�l�`��ŀ 4� �'��PסU�����EI	���c�'�<���Y�g,j`�@$�Jp u�'�[0�b�0	�MS�Fk����'����t���/�l�����A+�0A�'"��QgG����xԀAo�	�'�8� ���g�ܹc����6$ܻ�'�$`# .ɕZ��#!�JRr��
��� �����VT�a{��ؒ �ʤ@0U�T����cJa{b+ĳ[�>�� ��lPY���͊�p>IE��6(���̖.�	y����k�b9X��GM�`B䉂EU	�)��Z�V�#��<�B�\��B���"�ӌ#���zg����O50��'䖌s*P� �\��Y0	�'_��*bC�z��`��q[�3��	+p%<P����wY� 1�E�� [����G0﮽+�D�EU.��#j]�e�0D�"Od��ꌔ'�8Ab�	��!~��n�K��LA�MӥE��2��+L��.R�1V�tGxRB��7�Jxy�AL�F��xV'��p=s��>.���7�U�8�k�H!K�4���-�Tm��@бe�@9��A��(��䕺i��xb
�#Lb(#C	�ArqO���ԉC!=��eK�'P]I��L�:��O:0�N�R�ք�wk�"�'t*,"M�?^^�G�=Z�$G v��ԻE%�Y|��Å  �D~$82��t����y�)W�3rv�v�Q;W��,i5����y���\c�JL HB� �0�� 2��6��<���4�a�#�x3Q�M#NI�$�O��R6ON~�0�hg�K\�I�G�'�f��CQ�+�>����} ����S@ʁ�sN!�nYu��.I8h�d�<�L�Qn��0<ٴ��d�5XebD�1��m�L�1��y��L܎K���
��XV#J(#3��N������N�#>ic��a�f��Ђ�=I��Y�QB���?�E�z4`Ѓ�J4f��3�],z�ǀB;��d[�a�?;%�q�e�y	 H�
J5��B^Ƽ�+��z�d���΅66���t��B�<��Ë�6��p*�}Y֝�RI�X8�H;���f���/K9uR �0K�heT}���U��{U�и�̗*�V��(�GƼ9�D�>LO� kd-� e҈pz�χ?`��%2�-�.�6�;��V�f��3��R߰�I�6���Fh^�$�џ�h��> g��H�Jȯ95&u��!#�I�.�PAű@j�)i��ǫT@�S'�b�gM�\�~��	@BX�D�ܧHq�8��'���ë�D�d�s�O
+o��j'
�9��P���?q���Ҧ�)�u�B��>���UO�)B���� �pZ� w��#�yItg_<� dҝ�d@�]"w�B�ɖ��)T�H����d�׼i��QI5�T���D� s�L��V.�*��d lt���dXI[f���*#+nџԩ&N�b*(y�U�Ϊg���I�� 6^x�2H�"u��<����.y��PCWy⤆�0b��92�'b&����n~�[��]�43�3(O�=�.P4su���l��K#�ݓ��ڀ��1�J�Rɇ�"��t2�O�,B�`���6*�~B��
s�Crf]3";�ӓ��U�ֵ'�Ѱ&b�Cr�2=��@9Ջ=�i�>���BR�ڄL��`&"��M�bq�����@	F��u��o�̋qM��¢�ٖ+�[~4�fJ@�ў���K�h�x���	H��,q��c�n�����8�"�?I��D� J�A���٨\h촲��ө#���;u�H�E��z6$V&!�t�z1�ν�x�g�8����
An��[�E���$>+p�����WV̡w�D(on�ѳ�0��3?j:�y���'h]N��#Gu�B�	�6ކ�p�E�B�py3�^�S<�
#�وD�R�t� �7W�I�Q%3�i�5U��b.-8��� M�pQI�k#2����`&9�@��+6|�Y��큨9t�*���"c��n��B���`�j��$*o��d�G��,�����_�"�x�-�1y���#FSx�F�p�	���� 4z
�Q/�D�1(�C�I�!�%��ዺc�m5nպ%��b��K�ɽ-�f�P7 ˄,�c?�kB�%~�4E�P�N�y}D�B�F+D�@3ի�k�@�f��풝��Tu+ÏAm��i4��1�~2�K�ʃ�|��a�ᘍ*�(D���f
S�)������7N��r�A�O4��2�(4�A�(�-�<r�քp�UHb�Y- jxÌO���Q`F�3�<�p��C�z�ôč�l6l�YP�E\2H��OJ��&*�'"JX@rSƉ�=����I0?�b#հJL�������*��4aw�I�"�l�;����y�-��F�ZrR�+G+�r/��R�޿jӢ��<E���X��0	�	�	�>����=
/r0�ȓ�^�(���-	;ą8��&|MJI�'r�#!�W>M��y����%9"�{�'C/~�&` �5�p?	e�R�vt��+TGȴ,L4��6"ܪ5�>���-D� 
�b2"�`����Gy��+D���� "���LŨXƬ J�)D�\W%^
� Yh�B��0/'D�4�5.�q��9S�Ɣ�ij2Pa� .D�0�'땼;�4C�'����=Ҋ(D�� ��i䋐1f�<��*QMD�9�"O���U�ͧO�T���(�zB䰡�"O80�S ��~;P)���OU9�(� "OT��Ƭ�I�\+%��#P���"Oڵ�����-�fA�'���$�P�$��xpm�Óo�HU���	��L�&��'{����m�@�+U4DP�X�dP�>l7���|����'Sp������A�e[�0qNpi��dǫIn�eR4����'EҲ�H��. 	J�x�H\ݬ��ȓ0
]8���.7QV��ƕ 7Dj�'��\#]S��OQ>-��O�RAlT��#rJ�QPL-D������8\h����%����Te�9��II !{��m�3�/m�`�z�Iٻ���J����d��n�x�y�.�]���aa"|®ك��Q����$��B,)��S��B	J)2D��5��  ��Qj����0�!(1֭�RB�BV�B�	�!h�}�e Q����JW5h��8Hy��+B*^Y�ҧ(�,�R%�z7r� H0Aǒ�@P"O���6n ��W)�`�`����~��Ҕ3�D�8�/%��䈤�Te�1E�=RN8r��&0�!�����]x���0���� ��!����W���E8�����hX\��[2x�d��!N�%��xbM�o���<yF�Z� x�P��[�u�:P{�jPt�<13Ğ�5�&��1��]c�D�p�<�#L�&66����ɡ��@v��m�<釯׫}V��T'^�U�������m�}���xC�6O�Q �z���咍O��a�O�qSA���ussc�?�)�D�9T�^eʀ?�O"$q���]�hI��g^r���I2+x5�U�:�O7�]Z�O�3����a藲Q�dY�'��H`2 b�0a蘿Ue���,O����f�Z��O��|AhA�;b<��	�O�<��@\�<-�^l�lD���1�c��@�z`���>�3NG0����J~�=yG.�R�j���靝7��-��M���P7n�"��<�g-��x{����a�1V�8�Xr��}�ab�S�(ݢ�[y޴a�&�Х��O\���i{�m�N|꧆�B����`ƺ_�r9gk�N�<�����\2��I��\JyRI���2� ��X����5�މ�T��FL�9wb��p"OZ�2��0���'J�t��C�Z�d�'�8�#'2��D��L�vU����a��ۗ�7A�!�d�N��C�Ζ�i�V�;P��0�Q=�n���8�x��V�϶kL$��P�G�e=�xN�	?٪5�<�O�!8��aB4������b�<1�A��9�����όDL��@���_�<Y�V�R�ƈ��]	8�� ���[�<�aM��h�+��Af@ (f!NH�<����"��]�b�Q��8�AF�<��*����貂G��0����|�<YaLT\��D�d��O
v�#/�r�<�e���L�!і{����b�XK�<�2'ԁO�.�!tJS�@���F��H�<!%��$w���Pp*��[��Lْ�DR�<yd��Q*p��c\�s���J�<)��5!�]!c��P�1���J�<i6�4y^8�bE^�
/�}h%��D�<irA˼�;gJ@��I���B�<���֛�1���g�
��q�<Q��$�PAJ�L�:��e]r�<�d��;z �S�AݙlHQRja�<i4�݂_�����@��s���C�]�<��k�(h#<����ÈpM��ehWT�<��ƐF��]'�J�!��ɠE�^[�<!�f
ވlbtƓ��U��
�R�<� ڝ�&/�r��J�EJ?&}10"O@�^-ٴݘ c�u�~ap"On�T��
yvdM�p�0�l�Q"O��x¨D�?.��S�Ȉ"? d*�"O�<�$�SS.:�k�`�/S,6���"O���u�D�Xe�2�\�B����"O^ej6���`9r)�Q������i�"O�e�ł�^~`��P��`yj0"O- ��<xSX�oH�j�UAI7D��ɳ�S�z�^,�Q�_�e�^�`��!D��[alI�MRt��g	l�vi��=D��91K�?m㪈�5ņ�if^��`�?D���#��=��\$%�,�p�c?D�HH�]9 Z√�![�o�x�Jq6D� �_�e���u+�"�`�Hf�:D� �D�N� ff4Z0��>e��(׆;D��ct�=%Y2E��1f�%D�X��	��(��yb�j�v�6+S�6D�t�'�&*h�(BN�bV�� RE4D��!�`X�`؈F�--h����?D��:#�ũО��qC�+�0�H2F8T�<+�@��:��BX�}QP�I�"O�X'�	;Ah���6��/�|���"O(X�4�آ>R`����&_�ܒ�"OSZMߞ5��Q�0�N�в"OR���"g��3�*��
��	��"O���@Y���Q(��.����U"OY�u��X�AYUf��]���"O�����(�T���R&C��A�"O �E�6$��@&c].O��j"OZp@ [�3�0��0�˽&l�:'"O����D�b)f�h���)5H�c4"O����F�,��+��#"�af"O���3,]~��Ǐ�6-ɒ"Oy5I.(��C0F�W뾹��"O��d��`I�1�vb���T"O
�2M�<{�v ���AQԍ�e"O�k*�*P��X"����#g,�q"O�z�c^�������#A�Q%"O�|�GW.n�f(�&�M�P�My""OB�{�E=
��
Q���"[�	s�"On�!�L7(,��A�s�iY�"OD�pQ���+=�qȰ��X��"O�I2.�>+�<��膴'.�pp�"O��
���tr�t
6�ۗ2��Zb"O� �J�8�>�b�!��p*�"O��i�AD&9uV�!��T���)�"O\8J��+�xxX%BI��ĭ�r"OZ)�T�; 0�@	h&�:�"OH��j�0}���W�k.��b�"O�H���́�;�O�s�"O���ֶLL��;���#ft�Q"O�W_�j��E����!�L�u�<����3���0��,�l��5-�l�<!4 Q�_�f�B��.Y�h$b��Hn�<Y����y2@S�/Ҡ���oIq�<	f,���}"�KJ��9�$�y��O��D���v�XqC��C�y2)�l�Љ9&�20�fā���y�Dԗ$IF��'��.��4��y���-/���I
�R�te�2L��y��*�t3�X�Y?��0����y��D���qJD@\�]�J٫%R(�y2���v����`+K�:ݸ�A%@��y
� 8<�sO� gֱS��=N���"O�ey���;��t+�
�j��e�"O�a#��Y�+�H���fV+Cc�x�"O؈bE�;���iR�A�)�h�`"OV�V��$w��X$�3G�lݹ�"O&��Uo�<�`���ƽ �F]P"O�us�mG�5&ؑ�F�W�h�jpH�"OZ@2���6��aDCQ�"�0�'E�@t�H'��		�P�˥盿>�\ 3 �Z�j��B�Ɂg�z��b	�;,��lث#�rb��̘*!�xhF�Ӥ;����`�m�D-�[\B�I�v&�����Z�ڸ�0�L�{�48Q��9Ol�˓2��	��L����\�h�M��抍4��P�?4�����:&��U@��`\L��`�5{�^�3ª�pV���	`�)�$K�Q�v��4܎b����dR�n���]a����z��Ǎ	S��)r��9����'�>Q���*=~�4��g+'�t�N>����)!�H��C���T�˵�k�L���*OB��"OƉ(��]V�0�så,\����ꝋt���H%+C9�4T��E�-
���&:��%JtV���J�7!���I�8ͬlh�OZqC@A�"��&XlH�)K$O̲.F�9��
�	K����3F��<�r�'C�XS��8�Q�Ac�h�S�}�D�9(Ǟ�g0O��&%�rM����~ �pIa�,�0��u��:nd����iӖcɆ��;;�Xa� [�G4��qq	V�BF������hdcX�j!zPd�::�@!0@ڃC2���'@L�]�{���0���sC�-)d)� WwPB�ɝ`2t���5n̄j�P�Gl�	F�8*(p�1cM*A� �k���a6x�����6jȔB��Pxy��
r�ꬡbO��,��DY�̺�p=���K;9]N��N
�-��;��� -0\H�!I
eTB��b�=q=H�L\ ��ߚ����6_pe�A�6fŀ�)���'�h܋T��D���� k
�D4���-jfM�2 :�5�#�ihd���
S���s������U��FpC��>Ϧ=Rga߫�F��ጄ5�v�#�lZ#t�ם�U�fKa��Y�F4��OkB�u�m����'�"�j6&�pv!�$w�B�)�kG$9R���YQ
��d���P�y)��#T����(IT�	!��RE�.�剰��X��J�<&��@�	�0e���?A��(������SŞ�났��Bh�ayՃ�~>V��V�"%�"�X�����
J���r$(O�Phc� � er2����J�R�0����  [BRX���� )K�a��$6�b�&|�d���B�"DAK13�H A�7��q��^6I��I��.P�&��A�F����}��
�9j�@YBeړ�R� 9?��F@Ag�Ҷ���C�`���u��PðA�:P�m��I�VɕI�,h�a� a�"Pp�Q%lɎlɤlv���ŝ��隕-Η=���
sI4�vOr$g��4;U�`�ˌ�R�>P��6,b4�[f�@d�6A�q�(XW�u�
�'�����6P�%� Gf\8@,OpPI���`��Ш��$9�Dlc>I��@Gen��qf�V�{08��1D�Dq�Yq*�e�T�)�,!$)���)�"Q!Z!FŘ�) �A�\��Hݰ�	 ?9#� 0i9�BիqZ���C<1��!:��1�ln�Ќ���S�D�(�SK�2,����L	z�4�h�� OԱ�t)��mH��)�Q)�tˑ�'o�)iW�H.G�X\m��v�6I*�*4��a �H�=�~@q��ĭc�!�\.FZ��FR ,\�-��E\0&��O�}9g�H�w�091��K���n$�����V� F�ԃb2R-�"O��;A�-y��u�5�Y�!���Ύ�v����l]$Xt����h���S	�Qw+��@h�i2�ܣc�!��-�44�Ǉ�w_�l���+���zv<� 7ϕ.�t�剾>�� �,�&c�fpkCX	����D�7d7��!*��8��h����.Cl���DŲ7�Z(q��7ːx2(����)���z(�|�!��<�O���w��;&;89�3L[M�KTY�4xes�cF�1{T���U��sC%��0��(�Q�	-�4	QE��86Q>T0��ͳ��)�矘�c�ܖnԴ�
e�C�T�j}y�+8D��3����)�txrp��#&D�a�"?��`ƦTBD�
ϓd��tZsj
4O�f�����	*���	����K�	�<�D;R&雃g�;�!�Ē	��Å�@�dJ�98����	?!�� >�)�숪z��$��KJ�(6"O(�[QH�4EecQ�)f�� Q"O\̃f��&ʹXg�,C��h�"Or���ㄿKf��3�G�sB>��&"O���$O/�Q�AcV6i5t�ѧ"O�)j1�ѨQ%!Z#!�IL�)Y�"O� �&�w*��!f܏z,f�: "O�T�Qޡ{@��Q&תI�� �#"O�M��lޓ!�DX��T
C,$���� hy	�S�X�U �&O�ր�Uo�u괉���S�P�²a�< �-�0���Cj0�beEF�.~�����3�#�:�*dXԫG�K[�GR��_�؛�!o�S�q�4`0M�*��)�G!��J�fC�I�l��} Ԁ�����c��%Ѻ�~n4�gϏ��`ҧ(���q�`V�:�`HГ.ǸRɑ4"O:h+`G�c#(�&��!㞼�v��@���&��РH=БѳN�b��i���8)D�b��M1�Ġ�'��l�,,�$I_���
V#I_~�Ї�	32��=IEj՛I��d�#T.%Ot�?1�ĕ�Sc>�z�$�I�4X�J�yr�R(d1�uxCL;!�H�����#%\p���E�F�Rn�� a�Z�/�S�O
��c֮��`��"J�'4��'��2t��OD���'D2�v9�.}r��g��"���{2�$
���rs�ƫ��� gY0�x"��L��B��}b�����Ýh��`[����+�������&��"�Z����X��p<����Ct�b�'mW�R�2��dJ��s��TZ�!>D��b�M!.O 5XEļ5�xpؠK?D�4{$��>�l�AA��7MU2|p��<D�p	aτ)Į���-��&e8�[��;�	�3�%���'�x��aآ�<�[wO0I�H� �'�h�1��WI"PX B�(_=>�ɡFM9A��`��'c8�z0�٦~���P�l�-,�x����A e��9��3��'w|��򤖺N����Vj��m����eNx5���u����e�&Ֆ'��QP��Ǯ^Q�u�OQ>E�R)O�Rۮ�b��E��h�f�1D���ԡP'8�0���@�=+8�7@+��	�yB@h�/A_�3�ɏ7\P�2��1'�6=���?���đ4VH��B^m$B͓%�R�w��K�w'���	���!�"GQ�����BaDb'��O�u���\�S�*���RjM2cV��dGL
�B�I����d��1n���H	&��ʓH>ʘ)��� N �ҧ(����e���s7�чM�$*�8�"O�H�B�Q9)%��*���)�{���d��%1T�)��'���U�7��F`�1L��lx&�*!��՞2vABaj߯U��S���QJ�Z�W%����$�Ͷ�s�F�7�8�h����1��xb�8�hx�<y��P.)=ʭ�ŉ��6kxy�Q!�p�<�(S�3�hu��,߸U�� Lr�<y'��/N0 K�A��.��aaw�<G+_+|�(�Ae��7CR�5��[�<��*/{X�U�G�?������P�<)g�`���������ܛ��x�<�Q��B�=����B��a�<�jJ��y�Ӥс\��=�ΜG�<�VkA��V�P��֡ ��ĂB�<�#mïƱ��c$�c�$	W�<�Ggαk{�����(r���H	h�<)&㉘/� `�IJ%�lA҂Ze�<�t"��vv���G��,B��@h�<���7N�8!���U�PD�k�<�D��ZB���(�Bb�����]z�<ɆGT<U�\�06)�>���W [p�<���F*|�!ag$�0)R5��x�<� ��B��Z؀ѫ�S� ��"O�R�Η?;*���G	�xg�AB"O�KG�F�'�4R���g6~v"O$�Sr�>K�ܘ��	��!s ɂ"O*Ls��;;��%�ǡ��;Qa� "O���@"��d;JAaРV�-e�y�r"O��b��<i� I��5+�H�<9rJ��ˀ1�+Y�T��Z�/JA�<IV,��.+�ZG�M8P �G�B}�<a���:���0��
�e�GM�q�<q��;0L��:��	�c��Z�+^d�<��. �izB&ޥiS&-Y� [Z�� Y�7.��+p��s�n��(�-���i"'�3S�D*)D�X{�*Z/"h%c�N��˰�mY�<�aξM]��	Ţ�J��I�w�*D�KC&�T]�	G�<��Q3'K(D��i���3�*]q��I�v���&D�pH4ˊ!a�l��/�?�8�pB!D����W�&t@L���]���7�>T�P��:�ZaSƋV4`�lB��I�HO��Ivx�G�_4cZ�hc�ȸ9��ɽz����J�3G��S�'���O��Q���D!�6h��^�0�	\�YL�I�@y��	�1v��DJ��7"ql���ƭJd�k�$D(�t�'�(��ᓶz^�}�!ٍ{�t2P�O�!��l��E��1��BH	�e�3�	V70u�q�f�i���G�@<bq�O��@����<���	ç������ͥ��Ѭ���F��'n,�����f���$�>%>�.~���.B@,2� �����v
�@�Q�S�O ���*�*�䪚����p��O���P�'��좐&� �0�+�M.EsP�8
�'Q�tqAA�6�b\o9E��x�%"O����M�,���"C>0�HxE"O�1�cPj�a�A��0ި��"O���4�Vwδɔ��Ŵ�u"O��K& ��� ���ۗ7��C"O0L"bx�z��R�(MjD��"O�!�df�.����ǜ#1�[�"O�x�)	�"pUZ2)N$\�2���"O�����Ox�UJ'h����"O�D3&D��(�A�C/9�0#�"Op ��KL�����O�*#���j!"O"����ό<�r���NҢ0��ٳ"O�}��)�+��+ .ߦ-�t�"O�\q&ݨ�2�a���p��˶"O怘������k܊D��@"OX�����wڬ�� ]��R&"O�P 2�^y�pq�*�?+t���A"O�YѶi5_�>$�뇕o����"OEr�o<��Znb ���"Oz���ѹ&܁R����:htIKT"OtŨi��,�Ƅ�d�G&h��"O���+݀`e�p���3y��"OX���-SCJ@��e٬1��4��"O����퐷J�z�b��<y��5��"Oz@Q gݝX�ej��K$iD^Dh�"Oj$X4n��o4�2���?H2D	ar"O��G�Q�1�"mɏs0(��"OT}���O�]�4Y$�ؑ`;(���"O<`q
A�%@����.!(�"O&��g�^�sR���&.Ѽ#�"O4�aS��"tò�j«^j�A�S"OZH
%+L�%z`5@�ꈉ�͸"OD���<z�(�	�##�:=��"O�=��I� G�~��v�˛�.���"O@A�a�� :�(!2F�R��7"O� ����*R,+�4h:���27�TE2�"O��)�*�_�Ɓ˰EʬH^r�`�'"��ӦP�#��X"�",�d[�'�֭�v�Z`�����\$!�-*�'�h�dc�4@�P :)����*
�'�>T����A>�X�ЬW,���H�'6���g����!BŌ�Z�!�'&޸S����yJ]�.�~��pA�'D��"Mɲl�\1
��Ջ!�Hq�'�N|� �06���䍸O A(	�'���BC�G�1���(�b�HN ���'�����^�������;"���'��,jW�\�N���).k�i��'�Rt�P�V��r��u�F�#����'n�4�pD@�D�H�U��6H�|��'v�Y�Ү��?��h��L�t�z�'f�Qt�E�*ŀ�W&�	)�'qRH���2\؈��+ #R�*�{�'��Y��I /u���s��K0!�'L��*Ձ�P��vk�F�`	�':�m��K1 a��b1O�/:ƼI(	�'���ZC�&P�H�U�θ=�\9��'������pL�Ӿ���'�Ĕ��Ƭ|�r����u�t@�'����8��!�p	6u�8��'Fv��nלz.j�����q�'��P)���+\�֐����H�	��'J�%�`�2% �=��Z/B�X�q�'!�Q d��FERdTȲGW$��'	�hP�b��-�&��S&�G��q�'*�d�4N��1�đ���2g�v���'q:����B�y�D��QGڂ�%K
�'�tZCE�t���Ɇ��))��C
�'�T�*���>r���ǘ5"hpi�	�'���CͲ)�Hh-��/�jqS	�'}��Z֪S**�<ӡ.�#:B��'��j��M�N@d ��o�'`}`k�'&&�`5��F�зïTGL�
�'�^���Լ&�l�ׄ�Q���
�'K(��fR%^�
�FD+z��A	�'�*�86�H4I�je"&F��b� ���'e.�(�fݐr�Ր.�,UD$ ��'[>P4+ϓJo�]a˘=Q�y��'���9����JFhӡ.,H4���'e�Q�c�����b�_�;n���'�+A �ِ-���5�m�'Œ�AP+��
]a�� ���'�<�2�f2M�*��G�E6ABZ
�'d��c$�8W��E�M�33���	�'6�����1:�R@�3�Y|�����'���; #x�^��BJ�@\�,2
�'�<���C�x�"�R�	ǁ?�ب	�'8�p�!h˒s�x9�� \�A(	�'�.b��'mr��WJA�o.�ٲ�'	L��gmX(bՋ6 ��T���'�@ �!��L�,����2E��1��'/B@���p��h+���@���'�DA�W-H�:����z�  X�'7�hqE�FJ�ȕ��$zf�i��']J���d�:cg:a�]��j4B��y2D�4d�d��Ү՜|d���y�L�9p�jw��x0�Ӄ�N��yR�C�V�A�e-V%���c�H�yr�2b�={Q搃#�H���y
� �q��))z5>#�X Y���V"O�%h�BF0k	ڥ(��!��-c�"O-�d ��B�{�b@^d1��"Of� �o�`�I%��*=Qz=�3"O�}B5�L0?jt���;@;̄�""O�1p� �l��W����U��"O�m�"��.Y�j��� �(�$�"O���p,B�~�%�V���dV���'��t��T:��y�#�S�vK��P�'�$�b0�W�*LKS�вqH���
�'IJ�"��h��xE��h��P�'::ɱĪ*��D�I�S��;�'j~�#j�jG�]�7`�R�B-��'����U�ɟ��(�;�n�a��r�<Y � 4����i�9gO�����j�<QR�ĵz��P��ѮS�həF%�]�<aVo��&��x��M�#��ɗI]Q�<���̽)�	3�`B`|��-EF�<�`fʦ{�,�w`�x�N��K�<�E�Ӄ|� �d��'蜣�b1D����eU(���b� y�=D�x BL�O�Tlb�(6ڢ,z��;D��[#�
]�`����>/�H���M;D�t��a���5�Qb��Kl
( �;D��" G��n�b4�ȃ�u�Ľ��$D�ĩSD�3K�\\أ傉;�Z@�k#D��"`ü{�����.�)[�N)5D�xjs���9���R��J�nOv� 0�&D�������K���:�cGa���8D��Y�D�
�� h$�� 
)��5D�L�Q$W>vS<����Z�2����Dm)D�hr�EњPJIiF�I9ΐi&�&D��
�W���e����9�p��$?D��T�M5�v�bB�oSH<D�ܱ��OK�h9�Q"����Q�U�:D���
�f�z@����`��PH`�*D��3��M}��="��E+;�޴�1m=D�$�t��,@�
z��c�,���6D��CqJX�3~�e�Í�"2A)�K:D�8�צ�w}Te �П)]Ν;ԁ7D��A��D��(�GS�H����g4D�� �L�,O*^1$E t�0�2�M(D��Q���A̬���ٶ7��!�$(D���`�\-i�9`�%z@(C�%D�p��A�lz0���fPjb7D�4i�(�?_0��&Q�,�Pm!D�X��C�n.�*��9�	���=D��A�G�J�����	�Y���JF�6D��Z�ώ�u#��t-�	+�+��.D��+����[����LƓP�b+-D��9qO�XAH	���8�p�8�K+D��z�E1u?��$�)�,X(�G<D�術ʶ$�ܑ�v�]�*H٪�?D�`�7��0ut�:��Z�w���9D��X��"�D컐�D9$��+"�,D�H�dC�U�uH���,�!�#6D�P��c��������1yw:�C�$4D�ЀeT,
�R\���U2`CR8�E�3D���`�,[���U��yxÕ�,D�X�6EJ�x����BN�S��aS7�0D���!�Rs"�P Ά31�=�TK#D�`WFO�{80{i�e��9��.D�\q�@�7�B��gJ���, �i(D�( � ^EgL�AR �1�|��!D�� �-�Ȅ6/�^���H�~.@�"OP�+U˞;y�l��1ᘈ�~���"O�M��&���!�&K�R�D�s"OZ�w��Rd:%! , �Z8�"OҌ�G�R�y��@�aal�-H"OVȠd
ȴn �|K�ɮs��M�6"O2d VC](Os���I�!��Q�V"O�Œ'��v��DHR1SzΌ��"O����?JHa�fݚ2]ht!�"O8�Y��(�2]�Ě�EGF s"O8u� �tabxZ7��9�@"O��C��5�! Ū�)����W"O�2�lR�8���"�̪��R"O.��B.��F6���s���ڥ"O����OB�V�j�KE�J�~d( "O���w�͜w���a�W�<�jQ"O(���-KE�P�ǉD�t�L��"O�L3�.�$���JǸ_l93"O~����B���ЀIO�4nc"O���H��7��m���m3��A"OHh�ª����XRf��X
���"O�s0��"}l$P1G%�
l�0*�"O�<�A�_��5��H4av
p@�"O�2�9 ����e:9p0re"O �����V��j4��>BA�$`"OΈr�+F";@���c,)G��"O�4KW�[�_��z&#�
�v�r`"O�q����v�<���hҡ���B"O�ht�+���jL-
��\c�"O:�:1�[�W�p9#�E@�����"O�@��)�LH	u%M�J�2�"O���Anji�����$�Y�����y2�';�&�y����`I
7��y�M�;t�(�5��m#��O��y��%T
�j3'���J2���yR�P^t�6��	F	���
�yr���J�H��AN����
Q���y2��8X�6A����~�V��SbE��y�ʅ�.��$"I&'�a�&� �y�!3>d�	r�[&le�4à�D&�y�j5_9���G�gǔ����� �y����. `  �    �  �  �    _!  �'  �(   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒��'��h�]���G��1y"Y;��=m����"D���)մn�%����;H���o#�	#&���ٔ�G�OaЭ�G��?7t-���Y����'D�8K�-
�8�n��K�E@�����Y����FPy2`����I�w���Q,3dq�� 2)̀jΈB�	�R	DP�`%�'a�E�plȠ%n(�(�HL��\rID����S$U$�r|�Pb�,=�<A�F1,O�����Զ�x�������2�BE�¼A���Y�7�l����b�<A��~�4)��k�O�D��~��v����$��9<��!�'�F�O8h�H4�F�?�2�r&ʘj�P�'?D���ȶ�^��S�O�x�^���KD�o��mId�՞|��E����
���K�ҡ��	0 r�|�5����i�}Y�)\(���!���26LP FƷu>@���*,[2�9�$k3LO�As��iluC���!a�\����']�Ma7��$W��BD�U���� 69xVkÇjl�DB3�\W݆��"`#4�h3�#	]`h)q��wr~���1���7�~����S��Q���q�' sV�a�/�!gyr8a�Aw�^���4�lR�k�3j�j$��x�6A7	�e8��4�Ə���s����-*�h�k�B�44:�ԑa94�� �
o����LLC��
Or�����^�>Y#�����<Y�P(xf ��OF:y@`�u��E��q4Ѝ<����
Ӎ�.��P �M�.�aGv-������`���Ɠ6�I��a�+J�����±x�Z%�O>���I�#qh�H2Ȗ)u:-{��i�{���
0�t���c�+!�؊4����d�;Z8�1�f�֜"��Jwb�;~�V���K�.6h�k%��|Bm��]���`1�Ksڄ��/ΐx�l�$o�~h"��#V��|�0���l�M��B!�=`1܇N��z2�!�cCD��W���靣�<�Î�.e/*`�cI�K�a�%AV��X�JE���� O/!��/J�<�+d� ?~��u�
�1O~��q�3JEn��3�'mO&A�Պ_0'@p�a���vy�ȓ`o�Y��!K3+&�:��[�r�<�����52/O�6m(�g~�b˗��5�WI�I�$��*��y���/?L݀�͕�@�<H@ĢA$�M��헉[P����x2j�!rHW2t�����:)(&���I�/X�H�'m�h��ܑ;���c(W�9:�'x�Lq�o�4ow��Ue+����'!.�8WΟ��<8��V�4�>IA�'��0�Wm��a@��Y�(�
ni��'�r��DLǒ#d�H�F�7��'���ӡK�R�b�*��+)֌��'wLD�g�\1'��#`ŭ*(��'66�f�	2ʱ�h�?MDIy�'� ���ݤ���PAGτab�'->X�FH��p\j���)U+ul�	�'~��+���\�tq��K�6l0J	�'F^M�2-��=�&ę���fp9	�'&�z��z�@���z|��'���[�M���D3cĜ�>��Yh�'���g'�%p(�T�A�>Sp�	�'[�y�5 ��:?�T�%!�>�v��'��5� �#�D�85nN<�9��'n��zB�wxE��I�Bl��"ODU4�/:�9H���+R���"O�r���r��d ,Q�ب�"O����.ف
�v@���N-)�yz�"O�h{�Nՠbǖ%�!�Kq��"O8|P�,�&@_�U� ��"�иB�"O��q�d���Lpz*�){���g"O�0����@�Q#�!�H8��"O��C��+E2Tbc��S���!�"O�����O�f�l��*��@Pa�$"O@d@�c�2HZ��҂C�A�f"OB��E�@�F�+�.چ&`�5�"O�d�P�NKȀhE��OFz�"OZM�a�
?d4�b!E��;cj��e"O��p�O׍Hn]2be�$nV�Ȣ"O<�K�@V'*�&%���I�aH}��"O�`@ M�d�Y��ɛ,4�Fl�"Ol��L�(T݈ԛ�Ԇa���"O�0bR� ?' Epg�V��썓�"O�0�Df��qEjB����DԊ�('"O �:bN$�H��BRҖ�a@"Oĩ�D��Z$��
��i3�2"O@�c�B�(���8vϔ2N�Q�E"O�( &�T�o�Tc���K�9J�"O�c狎+�X$3T�b�΄0�"Ox���cS�p���%�X�fx"�"O� *d�'��0oj��W$D=e�t���"O�r劝�1���Y���LƐ�@"Ox8�Q �kv2��'&�.b�b�R�"O<�CֿHN��EܕZ�>��u"O�i��	���(4�Ɂ\B�"O��Ai�1�^LI��Z�yZ��0"O�
��?f���i�7%Th�S"O^h�E�?��cqoر]��R"OV3e��-v����fj��U�Qf� s��cU�BoX�`�m${G�,������=��B+D����8C��4������t���(D�d���/ l�&��b&D�D�F�/Kx-����6�p\�p!0D��J�(J��HA��H��9/D��33D��)���$@���B�5{���0D�,xP�x�DY�զ�/���y%�-D�,��oU�^�bEqr�)94�ٱ�,D��SGK�Z���!a�O� Q��i+D�t	���/��$�c���,\� �)+D�����T/Ԡ�6bW8%_�q)*D�\q�牤+�ĉ��Y3S���q`'D�D�G'�0e��.�Jv��� �#D��(���)tDɠ�"j��1�N D�t��G��^�$ ������?D�<�ALW�}*Q;,�>c�E��"?D�� �i�&�6QZ%�Af���d�=D�P��m� Q`C���+D�(8R�g;D����8x�̜ґ�L4/���S`�5D�T�H s�,�q�H��'�N� wN9D��R�͂L�����K�j�� �`8D��k��3R����P�^�'��D`�m7D��O��Vm�
d;0���6D��c!��[� !p��)� P��1D�(�@��=:�DX���F�횁S��/D�@hČ�9n�A3�G�?9=�1Q��-D�d�M&>�RLR���2�b�`�>D��XF��f���z��!��9�L<D�4�e��/ژ�ɃǶ�,\�f�?D��	��[�2ج({k@�Mح�ץ<D�LQCN�!�X��1k]�WcjyF�?D�4�իQ�`�����Y�`6f�qh>D��!R+J�8�iGk�*�81�%K;D���d M�ZXy�jW�*�ň8D�X���J�0��)T'��!8D��!�����؈�0��3]ޜ���5D����R�N�(�D�Q���%J3D�TK0� 'h��(�M�&u�x �@E7D�����)fH��j$ޘE74���o3D�p�&���_��X��ڞ^m0�P4�3D�@bp��?�X��G�Y"Ѻ����2D���amʣ̚�
'g�#M�IV�2D�x�iٖzE&q��Wk<v�1!�.D��)�-��p|��t��b�M�&j7D���.)�(T�r,��s)D��bF�?&M~�����iS��:2�'D� �f@K�
Q���3톃RZT<aC�%D��3�/�.�ȔXK��:��!�&D��Y[y�8���(p#@=1��F��yb��kFMi��N������y��j6�,��H�&��������yn�,jz�2'N�4w �$b��yR��O����iWuh��ՋD�y*�!L�~	K��8U0$4[�����y��M����#'� F���s���y
� �,0f PI>vd���>� �"�"O�<�B��}~l2��^) D!"O�� ��{��r�\�#���"O���3$�
M'LTT*E�U�-[�"O�$�@��.���s��3���['"O�#��I<ے`��lĭQ�"O�$!H�p@�)ѠK�=�Zᚡ"OL�;`�>NVX���
�3�"OB���#$�1�f �`y�3�"OP �0�#Y h��`��!3`nQ�B"O��Oǯ}�h�r����^2,�c�"O(u��h����"��Rp}Z�"O><�)r�p��Z$���À"O~�x�-
	l��xa6d:mРc�"O ˂Û?Fp9�q�
*�����"O6���F]A���*�OQ�4_�y�"O�]�� �9.Ș���
�|\��4"O:�&��8^�)��QN�^��u"O6������n�m
���/7&�"O�,��EHҁ��/�N�k�"Oȝ��E�yXj� �j�	l��X�r"O�`��h� �4�#�&F{� Rt"O��â��ZӨݲ���
S���3"O24)�,��fLjP: ���Tʠ�@w"OjtCsI�kp�IU�T2s�|�7"Ob=�MߟQ���{r��2R�� su"O2DA�2e�dP!�
�S��9�a"O2؂�F�Z����b�T �~,�`"O<)��K�1�`jc� ( �Z8�"O*�CE����:���͂�v"O���SC�+C����J5F���b"O
�Q��7������!X��k�"O,X�S��?���1�jA�%��"O��8%HM
7"UzT�O=-�i"�"OJq���ѓ,�JZM��iD/װ�!�I0vL�� �N.��a�K5*]!�ʹk�nh���R-r\h�k۷3�!�d�z��(Q��vU�*��=�!��/Ws�=Q�A���P �]cW!��ʞ,��?g�NM�5�U'@<!���ⵒ�n� {�@&�`�v"O�A��ҕ0FrĀ�	�PV�"O��+D*7B5�i���oc����'D��s���?q(�c�G�A��y��(D�\b��9{\��$G9 0����'%D�pk���8��틵�[�و�#D��a�@��	�T�Qs ��Iq��B�.<D����ܦ{}�TCr��ELА�ǥ4D��+�S�4����ĕ�Tu�(h��1D�4��_�VXp�ⱭΆj��h��);D�t�Q�Z!V�2�r�KpD�8	�:D��+d��!n'��SG�F�#�8D��B�!V1���G(D�1>.���"D�x���VE���3��G�ZM¤���?D� (tn �7���c���&O��P���;D��;@�J!�>��e� ��BR�;D�l� a�j+&@�Ţ&[�h|"�<D� a�!]�[��	o��Y�4�Ӆ	:D��Xs�C�M�@MSD�2<��ҡ8D�l�D@�-���Ƣ��D�@C3�5D��x�f����`���M�g��l(2N3D�d���P(xd"��H��4m;D�Y5 �%����bo��F7v�T.D�ӡ�@�V��c!�&����*D�� 1#����p�F�C�T�J��%��"Oj��d!��Z���2�e��]�8x��"Ol��d�\�,�ƽp���xF.�$"O�(�n��j�@�p��L��!sq"O z 朅=���0-�d,�d�"O�m��j,��cv�ёq�QK�'R<�2�1Q@0vk�8^�U�
�'.��c*��M�hW���p"O�t��͜>l)��5xo��R"O|�"�S��p���(Q"̛ "O��*6.�
*�����ZQClA)S"O�a�Ł]'f���#̧�ڄ��"O~�gɗ���P�B@�z�>���"O��҇59T5p���4@ �&"O|�̅�'}ؠ�C �t��r�"O����C:B�(X���J�Xelq"O��jԇM�ɦ�]-|A\DC"O��k�n	G���T�>�p�$"O�	���|�X�S����i+
��"OX��S��1�$q����Ė)�"O��X�MD��a�#�|Z8�h&"O.���i��}��8���@ވ��"O̴�~I��L۝2\�MX�BJ�<�Ā��7����
�N�į�{�<1WgBUq�@F�f� R }��	��<c��̥a�޵�dJ�6K����ȓ%�vⶄ�A�½rM��(�n���S����w�A�kJH�ր�,�>�ȓ}��P	R�s���f�lА��ȓS0��#h�h�p��$�BR��}��J�� 9WmE�"= �������,\��"O� 1wF( ���1�hD�M��ͅ�hT��,M���釿*�����AL8Гhˣ"2de� �7�P�ȓG㚔����|���G�[�
�����`�T�\�<t� A�_�|݆�~����$N�6�B�2�阭E�b�ȓ	�	 '��L��CR�L�s}N��������2���)�?
Ը�ȓ_�8�v��P."���B��6��T�4�[�
/,`���.X*s˰�������a�js�m\�4}��J���d"�J�qq�,�cDi�ȓN
�xb�),i`��lÊI�|��ȓ ����5̘9	�]�䧎�-�P��CP�-I�fK��̑�Я��u��k&�E����??���Y�ゝ+:��ȓ]������2m̕��m�}[�1�ȓ7�2�P4�Ȋxf���+�4�i��n9����W�`��aG�)�6��ȓUyM��>U&�� ��HMnx��>}:����G#XZ>��j�	vن�)aT`��K֒鮙S6%v�$@�ȓ=U0��a�D��<�cQ�	�F�ȓ��A�Q��P����k�8���^�R��CR�%K�lM�(�N�ȓ�
\��_cZ��B�읳.�d��v��d�sn��W��LC����t��:�$9j��f�-S��496�Ʉ�o� ��k_.H��ڃ�ծF:��ȓlF�m��P�,����C�X1��\�ȓd<����vê���#�<X$!��G�e�1AXe����+��U�捆�=j1���'*X1��C��&�Ry��S�? t�th�ii8��g���j��!"O�mpS%R�B52в!���)���˃"O$�rժ6�ʡ[�-͓A6�z7"O6H�D��E���I;8 ��'&V��#hڌ>�dK�b
�e
�1�'@�	��S�-��P �W�	��q
�'����
X?rAf)���� i���'e�!h�O�7h��۶d�&	�8 {�'��1��!H�kT�����FP��'���Ȳ $�±�cbP������'z����@�����Sy��'��e�QN�!��IR��}�*hB
�'�j�0I��S%�#W��l��ȡ�'��9@ ��P   $
    �  )  �'  �0  �6  '=  |C  �I  �P  �W  ^  \d  �j  �p  &w  g}  ��   `� u�	����Zv)C�'ll\�0"Ez+�'N�Dl��T�1;OV��g�'D<y�g�4gfD� .��ږ}����'?���2�O�Ey���l܄@��"4C}ݑ�+��?e�'�W�?��F�8?�X����k�&����	uV���%�}a
U�l��KV ��u!?��4�'�*��&I:M꺍1���"OZ��C)B?|��pL�O�4��]�Fk�	8�ΦuᔣRT�I����ş��N"o�@��`j�~��2�џ �	��M�3�ƞ���O �{�����O���L�;^DR�$�@�H{��[���O�$�<���?��#G�4�'���)����D�ř#�Xݻ6�_*%&!��h>\�xw�!��q��������<�M>��'*����^T�d��m� �
� �T�r�QaB>�?���?����?a����6�I;G���P���^l�}
�@�N*�d�����ش���z���� ��i��4N��� |�\��G��I���2<��a��՟
Ez���O�Ou��"C�F;�X��f��H�*j�XD Ԭ˅��|�ӿi7���a�S�?��S г�VQ�F��0�d��%��D��1CN��M�6��,dǈ�`J�?zO�ɐ��A����5)�=���iӔ�oڵ�
�A2.�WQ�	��D1i{xi�4� x���0d���Mk1�i�27�N�U���<��(��/=El`W���5�*;��ē�f��e�^?�	Yb��C\<ɢ�i%�6���8%��3��Z�jO�j��苣HȺc����#�-���3B^�F�4 �4`�T���ޠH-d��ߑ8�D8���'�v�Xgk��11.�z�i��'�
��'6�O����O�MP���ݦ��I؟���D�R�J�p+
�2�2-��d���$�	�\A��������'sƪq�6#J7 �2��'BS�
��a7n[+=o6,)s�*C�ĜA����p�f	�j�>Ā��^L:�k�*J�  6����Ż�C��]ʰ�w��HO���V�'�R���a�i��[)~ ��I�)5*��Њ�Or��O��"}:�J�Aq�}�%'��{��y�'�O���ɟGw
m��J�f �����9A ��6��;@p#|��wE���i3I-��1��9xd�S�'����g�
�IБ�*3�T���'��H�G�BNP��i �9a|@�']f�2p��	!��܎,UV���'�Ą"T��$7x������� �'T�CM�p�����ے	��	��k/��Fx��	E/k|�ٚd,�p��{dOM�	#�B�	�lL.�b�s�H�*A���B��u�q��W�
�a�V�F�fC䉄K�*8�f�ky���4&Ƴ1+�B��;%	J�I%6m� � A�.|6C䉩<�6%��aC9P_L�H�F�&5��r����	f�,��MF�35a���Z�}�B�əl\HS)Ż 7�ܹ�c؉�B�	:	��i���S�\�a�TP��C䉸���
�w*P�"B��zC�Iz�����/H�h�8�"p��d�-�d�l�Y~BD���GK]:B�{�J�7�?�(Ol���O ��@�P�E���1�r�����ȟ����J9�bq`C�6��Zs�?O ���	�hڽ�ea��#���$ڊaR�HZ���!]�HZ'$ժ:�ax�f��?!�iP7M�O�(��ʦo�8���Y��N�<y����(�Ա�0KF�|��]BgO�jon�:1�',*�$����B���u������|�X�i�+���'��.�N+D
ÆH�)�8�����Qe!�[7u��q��j��C�́dMA:KM!�K�7B��r������c$ �	.!�dב!Ɛ�GI�1s&�ش-SB!��$�@��wKɗ�H�Qn.w!�_pf��`mL�Ey����M%Pb6��O��d�O�!r��/|�����O2���O��.N���MIA� � ��9�����5F��;R!RtRs%��Y�$�� 3��O6O��b2/K8@��`�Ӊ5�A��  ��V�K����?u��P �\�f(1��	QPFQm}r���|(����`^oɆe�eÕL&�V-�<Q,Ο��|�I͟\����<9Da�&��\�`)\�"�ji�ȓp��@ �\�M��sB���H�U�'��"=�'�?�/O��a�O.Z2���ǔ:U�ʉ��Ok��!�Ot|9�!�#O��a���%�X���-��s`!��8y�l<���T ��y�"ʓ>�6ȃ4Ob,��U�E5�|3�C�/�摺vN<6�@.�OH����0:H��;�� ���c"O��z2I�6I;�q��L<_��,#�|2�n�^�O��S�Fܦ������
b���5�ƌ� d
��ߟ �I� Un��I�|̧CvH#s�!� �)S�|���� ��c U9@�桩"oC Mqv�;�e�'���fIC�O~�h2�K�3:�(�s���<8�b�Ƌs�"́��ݬFi�/�*zd��	����'�.��m����B�cA�:�jx��?������(���b7ͨc�L���/`�T��'�V��߉T6"Шa�^�L$fJbP�(X%��1�Mc���?�+��d2�l�OL4�s���sJJt���חr�"��O����@q�KGբ̐�I7�����E�W�͟n��GoФi6H�.��0��D�!kлd��5�ƍwS�l�Ҋ�4�̙�N|J�d̆6|8��P�J3)�T�g��b~���?�����O��e�k����Bθ	h��K>���0=	F��M�Ve#�5t���`�'�ʢ}�'R�
`
�sBKX�������с�M#��?Y��'��
e�P$�?���?����y�����������H�z�	��7�h����X
�o����QrP>yϧ��9h��C���d�N�3dw��t����d��1yݴA�*գ�����O՛i�t}lҊL�������)q�\|�s�X2�?Y�OԵ�F�'>��'�O2qJ6��q��\+yZ� I��%D����׌ b8I ��#��}�e��<��i>��	ly�hZ�z�4�q�]�c�̲u�X��u$!7���'U"�'���'8R3�^�戉j搨��N�s�����3�F���ȅ�D;.�ҡ ��?���+ 2d�#G��CTz�����E�Pݢ� �=R�2���;��9�4i8�"=��&��	f4mkB+T�{K60�uA�##�p��I���D{2�	���ub4c��xI�)Jd�U4C��Ԝ��.�'FŚp��*��
D6�Od�n���?�B�nҤ�5xW����\+$���*�SX�<V��H��$�fa�$kT��r��BV�<ц�ïA�썁�ǝ1�N�b�`j�<A$ 9��A��i�4nʥ��d�d�<aƢ��*�<Q��+��U���"��H]�<�@.��6O�L	�:,�Lx�CGX�'��m���ID8C��B�OM�C���o�OI!�$J�t:�F�Է�P �$eA�cE!�d�U+���u)@`˼��a���k9!��$�B���J+=MH� EO�w$!��;^�t����.]�d�B�<!�$+#qd�qe�D"-�=���⨉��O?����ً<r��`u��o��`8q�i�<�P�U2�qa�k�A��y���L[�<�)L#a�h����I�5B��A�<�3�j�A�7�]�&B4"�/}�<i"�A�i���W&t8�¥�|�<Y0��=f�k���=#yb�-�uy�C���p>���֡��P���ôP��a�dK�Z�<���X��Dݚ`Z�!��P�Q#�S�<D�Z7��h"A]� (�*�*FT�<I��!}xe ���9ju�S��K�<ɑ	��B`�HsgҬ�ڔ��Ex�h�Pk��l ��@�s�03�O�@]~AC�%D�X)!@�^�.IC��}��fi"D�,�@��$a�X%�u���~��$��d?D��Z���#AX�r���M\��)2D��V�I5c��4Xeǘh"����-D����L���I�E,�,/|���"�I�H	>�~r!�U��N�q����P���ˆR�<�� R�G�x	6L�{�*a���IR�<(�,��Yؐ+Һ4�PLA�/�T�<��h
� ��Q����{̥��
e�<aEε���-��G��]IӃ�d�<A�A�._q
��r,��Eu�ɕ�A�	�H?�S�O�Z�3�A�.Y���r�BՌu1@��b"Od�[a/��M��0��`��m}���C"O�����.0d� �0/(}�Xc"Or�j��-3���:����\�&�t"O�����J�r�o�=�hu�""Oh�A��K�i��g��qAgU���P�=�O�H2#�`�["�B�Z�l��v"O� ��A!�|K�P'��j�z�B"O$`�6�F� (����JR���"O�H����3R���s��@`X"OQ92���]c@l� 1.��a�'��}i�'ش\��n_
���
��f$�A	�'��p���ֹt�qc�ЍX���0�'v���nK�w�>L��%ٔIf�Z
�'�^I�惖�>��(�暖FD�`(�'�\p`�˧i�p][b�B*HN�š	�'t�Jd]�9�ND��a7k�蓈���"|Q?���WGn�����d�Z��c*D���V퀴p�4C�	��(a��1�(D�|Kf��l9~!��O v�2@&D��j�($u��՘�ψ�^�@��4�(D�	!�O�;�>p�íŤd�(ږ�&D���%n���ѻ�`��m�<��l�O����)�]KFH��g�hE� ���CQ%�8h�'��̈�nґQ�:�D];BֈE�	�'�`��/�^(��l��<Z��k	�' *i��bO%v�DXZ�GU0��U��'������Y�=�fS�%��K  Z�'\x0��
5B�C���J���-O*�Z0�'���b�+{R� @d*ǔD~�Z�'��0N�'Z��'�/Xp�=��' ��Ȳ!P�Do��XP`Z�a\,��'˲����8~&���CG%]R��'^���͒�u&5�pnZ�%.��Z��h�I@~��
,Y��00�
�����9]�ɩ��*;(�H��LI�9���ȓ����I�4SSG�*`��ȓ�ٲ&#ՏI��s�%
	vR��ȓ,�֙���I��r�z�̩��y�`w ]-5*��Lž�G{R�A:������2Hˎ/��as�+��y��!"O�� ��Q~hD��&�[w��`u"O^]��&ކZ����dH<_ �"O2	�B��>��Pi�
L©;"O�Ui`Q�08`25o�"t�n��"OFu�'+
*%����(�M�FI`v�'M\]����,_U�����+L@f��6��Q��@�ȓƅ�'��Sw�
�IB&h��q�<�'����A�43������i�<!��K2lD��WC�1#��]�SeVO�<�\ڨ���� "�Z�����E!!�V}V9�����6���ۓl@< ���9E9$����/gT,��.X�H�jR'j˂]�!��ԣAUԙ�Sꘁ ���h׈ȷO�!�D�B�����K@����܃Kn!�$��S��q�b�+8����|��	�'9@��0-��g�ФX��S=0^(�	�O����t�#@T�@ 8�A�G��m�ȓlH��%��vz�t��ɎN������8�0��>9�=gj�p~����p+��sn�5z���ÇO�$��[�^���^z��ܳVbS��	��T�&Ѐd�1rԱ����]��F{������B��h�B����m�V^=	�"OV�8��L�{��C�J�?�b�YF*OX�C��h�z�$�#�X��'(P�z�l��|0z�xU�4l���S�'~�S�&]�j�L�� vI}�'�8���}\��;�'Gz����LU0\Gx���.sV��b]8��K���,q9�C�ɿ�N�����G�z���l�+���� ����MR�i�(�faTO'��r"O��V���o��� �����U"Od�����t�&�_��yD"OlD����}D���CdvxфR��"p <�OF�!�	j����U�4<T���"OЙ�M��n]r9B��/3@�R"O��&���n�b+��J���1"O:xxL
wȽ����;J=��3�"Op�Jl�;a�}�a�ZC��� ��'y&9��'�f,B��<.��7k�<!2�R�"O�-5F>�
�Ã�\.�ZyY�"O��{��D�X.�YS,�����"O49�S��9Y�N=9�`ߋ6��i�D"O��֡˚;td���  5R�6�Q"O� "U	ǥ{�H��v��r�P,��� Uw��~��AW��Hw��P ���5�Tp�<2 �TW��(��g ��J�K�j�<�"�(4*X���nL�� L���e�<�7M�"T^� v�W!3&` ����a�<ٴ��w �hF�3$�@��C�<��D�KJe��m70;> �ЃZ����FK+�S�O*�y����met��],��"O@�2�����⤜<N�V���"OT�[�J��a0�}�VJ�5z>9""O��i�?��3gÞ�8y1�"O�����^�趧W�qe>��v"OJ
�	�$.1i��8d��\PZ�D�3K.�O�xH���,&�J�A��o���%"O y:�D�2�B}��C1�¹B"O:L�陌|�
h���|\�"O�@YE�U�z�b��@-� fI��"&"O��wh f|	���7"=�8���'�j�8�'&��ĥY��YS˖��
�'FEt���z��!"�������'z"��F� ^C��Ϗ )Y�z
�'l���� !^���`��(�J��	�'g޼�N �$�Y�"-S�q(	�'g���p&^{���0�Cܲx� (S����TQ?�7Ə'u,I�KD������$D��1aH��d���¡;�P��5&>D�䪧FBSs� E��tR�f�;D�4�g�̊)+u��A5�`;�=D�0/��Ow.5��Hݨ'�褰a�9D��*"�G� h��R	"�r�S�K�O��p��)��\i�D[2��M��@�Q�����'y�٘0�Z�#�,bU,D,�1�'Tp���C?=�=y���8T����'�ޥ�G�\80 ��@��/�x)�'-�}����	d�Y��)VEڡq�'���#B�O�O�~����9�̽�+O����'�|�F�_�T.��A'�*W�pY�'ݬ�r�.=ơ���#�LC�'�`s�EY~�����Ġ��'(̰Ad��\�DqV����X�'�x�SD�,.�v!,�L��;�y�:��0Q��"]\X>����T]tf���Z�ň]X8(�(�h�`(� ��m�<9�H؎G����[�g�̵X�Og�<��jD��.Њ�Ƅ;>f�H2C�e�<�i�N��q�1�9 h\2�_�<�6%�>G�9�@h���d����^�'�N����	����]���`!cG�!��:䁻��Hp�|�`��[X�!��0�:M2dGW��ؘ*f_!�� ��`�灝H֘�y�JRU"O8���%o�1��&݊ �
-H�"O�1s,�Jr2͈���0-�XEz��'8\�[����1(����OƘ�j� \XQ\��UI6��B�LL�Y2@l
��ЇȓM�)������H����	(���"$5��I�(6c�T�'ۈ�|͆ȓ`��AI��Z�rbЍ��Na(X=����Y��@��D;L��dμE�.��'����k>d�Vk��LnY	ci�;.=�܆�چ}�Qh�8X�4��o_�C��ȓp��)�ɜ�k�lyfMG[����l}H�bҡÃ ��P� DJ�̈́0��6��0a7,��/�R� ��J�LC�����03� �I�6&@yPb�CM�b��P	D�o�bB�I�0Ƕ��$�E!e%XL+��N~>B�	�(��=`��2% r���H��#�B�ɗ��4�3��i���v�	9@�@B�I5D|�c�[�lk�Y���}^C�	�s�I��H�8�g��]4�=�wc�O㶸����+PwL��3��,T�|��/fb1*  ��`y�CL*B$��ȓg&P����
>M�
��� �$b����J� $	�5M6��i�J�+b�� �YZuH�=�r��o�$k��0�ȓTՔ����B,~�6��Q
rp&��	��#<E����}I�Tg��BLa��R �!�5	���Cn�&P�qV;h�!���W�С���E�F �!xVcJ�6�!��;X\��KԏZ�����еQ�!�ğ�&М���#�y(a�?@����D��=���N�X���8i�s2.��O�����|�����������x�aA��8 ��P��?)Ô��?���?9��!v_��)G��>�l�Q��Pcb���@�h�t��/�,�(�g�֎׈O^���K�^2��Ӧ	�1�b�z�lr�ђ�噩&8�ɠ�Ci#����a,o<��d����O���&�ӐD���b�ˍ�������2G.˓�0?� �M(�����ƎN��AP�Kcx���dZ).�%�,A6�[�%�mm�I�bn���֟h�	_�T�UKR�'N:9��{iyQk��ia�Y��L��?��HR#����u`�'�ܽ����=,���t�'@⁓��ӂT�]��lZ� �q�ԉ��"�
�e���s
�^wn���~-@�^l/Q�Եo�X���r��'��������ӂV`��RC��&ᾼ3K s�<�A�E�c�*�p���i60��6HW�'��#b����bQ@2�쎽P��Ƥ���?���?�V�8�y����?1���?�ƶ���;|�Q�-R:��0�'@�Ş4��'�Ʀ�3ra�4���Yv���?��'��'
`�x���Xj��a��#wx�*��K� ����&�`1p�ød �SΦ↖x�+��r0�]�D���41R����d�=#B�'�r�D}>������P$I���!%l��Պ/D��
"��S�H�0(ʁn�l5B�@�O2�Ez�O%bP�@��ԹI�]sbm���
h�c� u��2ش�?���?�,O1��
�[��pa�5��%O���D��� (a'�M������Bx�`Q" [z�&%a��T!���`[13�jh$�fP��@�Sx�p$��O�-�֪ټHJ�R�k��q�\�e�O�=����&
n��3�E�!i��5:��X�P!��^_$P�� �'~zU�ڇ��I<�M����G�Z���~�MO�
�8�2��8�B�ꐯK�����O����O2-�Ѝ6y��d��/=`�&x�i>�[��+�#��
hޠ`0�=�]�<	fE܈L��q+�A���)�	=�<aA ��-�B��g�7�x)���O���3�S.o9��c���:���D�7L<��0?��	�I��,��׸�x��u�Dx�4+*O>p�'�&/�iRw�
d�fI2�]��xr(�����ey�R>����ȑ��ʏ3;��"��/T�8 �ȟ��A�����As�)J&��8��S�OF�$�$�=#l�ms#O	l\˛'r$z1 վpW�`s�ʵ!�?ճ��"3�.k� %w�!���a�4*#�Od�D<?%?Y秀 ^����1J�%�ߜw�v��"O�XHb���L	V�y6�Z:���`v�	
�ȟ�]��A1�f���!ˠ��a��Op�$�Ov	��ʎgVz���O��d�O����O.<��(D�/^@�(ݙW�tq���+�H��"�%e!���g� �'��'�iz�NG�+s�$�'��9��=�D�Լ �tD��$C�z���o�!��id� ��I<�%
C*��pScwΠ�"dKb~����?���hOv��f�n�% ]c!�ㄔ�e@BC��*YA��XҊ�6`��e݁ b��r�����'��	�;��D���]��64����L�&1���Sş��	ӟP�Iwy���̀�u|<xf�@�E�	Iin���G�W��+�jʒ{%��t *<O���G�kJ*��u�J3r��{�d�7����i2|v�"��$<O�����'$�����ǭ/���#U3C�v�V�'�ў`F|�k2#�:���A�	�̉!�y���7p<8Rk8/t\���0���Ҧ��	[y��Ί��6��O���|>���
L84���v�rp�Qc��O�i��On���O,����v��u�D��#�� �ug��a7صӧ�ө&Xz�IA��OJ� L��v���)+&���O�+�T�95&��VC`3��¤z�$HѽZ#=Y�ȓ�����G��+��C�Et6\��^"6����	��?E�t�$h���G?a�.�YrH�A� �@�>H�I�.�hy���M1�@T�`J�20�$��?)��?��4���ӥ�D���Z0�� Ҕ5�ׁ$OУ=!Gg��|(0hr��iR��pDRC��w��%���~ڑD��A�~���Gn�D-��hS}~r������,}*��$^$m���e��	]��ԁ$]�Z�&'=?94�>	G�WR�d�K�S}�|á$Ó��I�%Z��b�Q�}��L�0��<�r�[�\QԘȶN��+���	Ҹ9�O Y�Ov]Q��>q[?-�6�]/`�E �/Ӭ1����+�O��
F�>)],"�zW�mh�(�Y
q��Ţ5���?��u�dt��d��F̛vIƮI$��ӗp�R���j���D�O��Nj�?�Ĥ6#N2g��!`�t��n#�~BH�����|�k����'�J�!�c�9'dFrî��8>	p�#b8�; ��l�	���p�i���|��Y�J̍b�`�L�U;���ɟL۴�OjX����<ц�QE?釈&@��C�f��OQƐ��K��r�'=�l�����@�B���/�.m���'�t��U�ZG@�E��'`����ߴ�?�)O4��|�S�l�I˟�х��.J�X)�v�*N���
�N�����O^��hO�S�K�$)�4�I�&�Hk�I�W��C�	�]���7b�2Ŋd@�&��C䉖jq��P�ܔSI����L�#��C䉪�=�aƍO�:ٔK�nC䉲z��@Rb�˃v��요�C) (jC�I-5�:��$͐%.~�Q�k �w>C�I[�|���u�\���;Z��B�	�aRDl�QF](C�*5�PJ�K�B�	*!wN �6�R[X�0թظ+�B�I�F��i�EQ
~$R�0�ɷ�lB�I�d��H���'H@(G�GJʖC��qt5ض��w�`H6 �7`�dC�	3��b�Ď%��Q�q`I�4(pb��QrJ�r��R�茰5�xCgL�/���ᦏ*z
<�����b��V�J�Y��t�`%�a�0hȖ�Rg�D�/A
0"���5���V�����E�e�:���#�U����S�V�r�Tl@W�|x�):3�ޯ7BE���#K���4'�>� -�p&]�v�[�&Z4J
!poq�ZLխn��P�J"h�����Uҟ\��/)dd���h�S�,O��PS����	a�V� ��!r��x��5�O���3Bڮv/�tw���1*%Y��x2�L5�?a����'�ħr��1eJ̾n���9�
�=(3*=�=Y����<�T/�v>"���@���Uؗ��U8�s���5U�J	��#tWr�#�/P���d�Or��D_�٘��~*|k0��"�!���<��!�S�L�)&�W�!��ݏVC����̀+WҮ��7���m!�$���Ԫ��0 �ݢ]!�Ӻ�ࠚq�C�z��+��Ͱ�!��#ж�H�-�r�L���
9!�䋌ac�5Rc���.Sԁj�-C�S1!�� 0�`�DAz>�j���jל]�"O:i�0&�6X��C�W�4�&���"ORaf^tռ���.h��aS"Oыp�72���	"�����1�q"O��I6��	z��3��2"O�-)aj �[s$7�:m��0"O\%�u�H��ZH���Ƨl�V��"O��j�?dM����H@����1"OB :��F�2P�1'L<�V`�t"Of���-r��j��J2U��rb"Ob$��A��7�v$��g�^�=)�"O���8 p�$�]�*�S�"O��S�>⸴(F��l<��"OJ̚���]P�@��A�'���"OH�ؠiٝ۠k�	�,-��XQ�"O�4J��:�J| ��\�����"O�I	� ^t���%�V�8�qJ�"O���Ċ o6��C�v�f0�"O� 0�鞖U����"�Y�J<�b"O��[��߁g�L�!�
}��"O�$�eo�E��%h��ݨ�ąsr"OޘQS���>��Hr��!3@`2S"O�\���	#8��X�=A��@�"O�}b�C�)p�br�5P.JYV"O�)��@�]�L�	 �ۤ5�����"O��r"�J�<���Ԣ8�� �@"O,�PgF49�=�$m�������"O�-��8P|���잽��Ի�"O��&EM5?l>��lǴA�00"Of�C&Mx� @*�
E�VT�U"O�1y��8y�n�ÇI\�b,�5"O�y`*ܲx($�0�n����	�"O�ԑ+�:b�$m���"�s""O^2��6G"�@�G��	�@"O^y�'/��J��0J�D���"O��t�/S����Hӎ>�8��"O>%�'���~�����͡F�2F"O��!vҎjN���cm
B%�a�Q"Oj���L�ț�!���Tq� "O>���>
�����P$	%�"OV ��E�*;���dL�a��d�`"O\�Q�Zv�>􀕢y[�	��"OB�����*R�E	��E��|I�"O�Й� �������� "\�$��"O�0�D.��-n$�2 �zYі"O�q#bD*j�X����$�>��"O����a�.'����S ^�S��]�V"OpS�E�$�� чB�py�Q"OJmx$��D1:�.էC���"O*�z�U%�f��q�	�+V�ɛ0"O$1�s�r�֤k�Kn���"O|u���3�L`� ǒ�q;���"O���兤��!���+V3���P"O(t[�� m�����}.H��"O|��'L)~a7�H�Z��a"O�qg��࣏#tt�6d�9�y��>��c�l��9PMr�����y�ʏR� ���˞�.ʹ؃�h#�y������D�,�6]a�J�5�y�,�gt�27!Z� ��p�Ö�y"��u<$+2�G�����3��y�Kмm2l�(E.n<�A���yB�#s���3V�'~+8�ZV���yh�V�t(��I�y)HH������y
� �qR�KT-� 	�Ǉ��v. �"Ova�r�@?Vb<�4-ӯ	8��6"O|9�$@)zj`A��K��L}j���"O$ ��ڢR��L�3���Rd�m��"O]1w������]2��8T"O$9k$H�@E�sdFγ\uh� S"O�y;e��0Oov#���N�H�"O�%ʀ�$@V�;&��88=
c"O�yX����L���շ8�}!�$�b����k͇_S����:-W!�D�9x��1 �K><��[�J�~M!�=wPف	�~3�da$e �}�!��M�FJ�UZ���')�فtd]:�!�$�<a'�0�e��w�`���{8!�ā
b��1�f�94 m��-3�!�D�*H� �q�R;\Ձ�BT�4�!�D�3+nH�8P�ڼ`�N�X5/M�_�!�ރH^���*$?��,`WNM$P�!�Dg�nܻ0���:hl!HH�P�!�Ğ�w�.��'&>²P:Vh��u�!�$:>��u�T*�Ҁ��-Y�!�$ݺU{��CBI�}
ޭ��G���!�4��Y�GM��R�L`���6�!�Ĉ"Q�r����X�0Ly6�յ"�!�W86[Bȣwf}����[�)�!���/2�p��,�$r�=M˷3�!�?l	8��R����Te�|�!��.H�B\��ҝ2�B�9�CǗ|�!��V��J�I�&�3$l۶�ҫ4f!�d�;S����҉��V��[3,��b!�dā5�:IP2�Jl���ٜ/�!�$�#yn�#�mَ4��0 �i�x���d�P���H���9SQ��#��	:�y�j@�3���#g�"���Em��yr����ǫ ln|�6��,�y2��3��!�&��L2S
���y�j_���I�o�� @&�УG-�y�"I��*� �u�.%��+/�y�Ūv���`G+�l%��ʢ���yR��2
_ځZFҏi��Ű��[�<�!KK'UnlP��M��!�8�kz�<91�D�	�:}����*J�uL�p�<9$,�J#�%B��éB%<��n�r�<��g� 56�����(\����w�r�<у��'�`�nJ�f�m#�d��y�+�����0A=]*��t���y��ʅ
�(w�R�8 |z��Ť�yb�ɣ5��@p�J�|��]`��@��y
��̓FZ<oH�T
��y҅�[�݂�J��N^ز�׮�yb�-d7*�zf�M$P-�r�R'�Py⤇,G��%��-%p5��S`�<QBoy�|U񤨃s��jT�ET�<1���2�ro�
<q�KP�<Ad��[�H�C�����`��]G�<Q3�S/s�`3f�K*�n�c���M�<��Ӕb�ؤJb��K����寁K�<����J".Ti���B�@�c�bJE�<�g� 37a�=&�R>�hiC`gx�<�V)Ã7��r���^�F5⩔L�<!��Heb����fz"A %�H�<�Ό;~g��H�b��~�!H���C�<���X�bO"�P�m]0R�:�ȄCIX�<I,�e�n0�')�+1}�iȐ��z�<� �@11jΝO��Hӊbz�y�"O,dbŠ��7�h���F^T^��"Or9��G�x �4����B^LAT"OdX4��(e��PTfţ���"O8Ipք���2f�'D�2�b�"O�E�eM(U+|t�ʂ�&��U��"OTpa�J\���%[ 	����"O�l�gF�'���a[�B���S"O,DAqGϹ3S�ȫ���.m�Req�"O�����E",1�u&��-�멋q�<�&��=F7<DJ�.�V�(��w�Bw�<��CO�O#�I(�a�|Ą�H�>m���һ?P^�y�3?��ȓP��Jui�5�Ĥ��*ߕg�84��yD���eO*O�$��C�D��ȓ>�<�� ^|AJ�.��R8�p�ȓ����c�"B����	�P���ȓ$LpP�@���؁�k"Y���ȓN���`uk��Fy�4�����9�a��Hq:��d�ƞS�� �ȓN��ŨB#�CL\p���Ʋ|�0�ȓ��yec�9+����!�
�xc�=��*��H�c)�:�|���D�Ǯ��ȓO�����@jΰ�A ��DS�d�ȓbX���僕Y7�5	1nO
/����xLM#hK��Q��(�\.�\��E��A�& F�b�da�g�L���ȓ�f�ba�
�gg��T��-� �ȓ;�֠9�.W���܀@K_�^�jU��-"�\�/�;0S�t���% n 5��5t��h��I�_�N�iU�5%�q�ȓJ�YP1m�#Vr�A����3\�ҩ����tcd@�'�Hp9&d�3;;�H�ȓT�����D�R���F-a��\��)���br��;3 i�ŊX,$�Ȇȓ!���d'I�^�d؀�E�IV�ȓl ]��'�<����ɜ�>���P��q��jd����N �D�ȓt0�]+�I�6`;�c��8<�ȓ9z|�R�L�U����iœw�����[(���5`G6k�L�r���g ؉�ȓ4�x՘��3>�Z�S�F��?����t��E��#�Su�A�o�>G�Ե�ȓ"�{�f�*�|
c@Y=1��L$������e��dR�7 )�ȓkI�]5g!x��Y�h�%�d��ȓ;	`�X�Ι)�<���P
o{z���{�t$��V�+n��g
BU�B��`J��W%��U�h	<:(����d�zC$Z�^�zbκp�:�ȓJ�\-p��6E��NI�s����ȓ_LX*��ڊ+odБ#e�2H��X�ȓ<�B�0v�)ՠMAb
2jv-�ȓt����*ӭ5M,0Q��M,Z���ȓ�`�f� �h�ꌫ1��i��@ж%?m�iK�iQ"8*p���$}��������"KU.x��LW����'΄	bJPAB��+�Hą�B�`��T�U&R�d}��E y~hp�ȓ	8����kz \8�d��\���B� W��h��<����?�&��K`�LI�N�r�$ȓe?{���ȓ&Y���)cK��¢5w���[�e�58���3��ƙl*Qr�����'C
l(�M)�C#s�$���S�? ��i��p��`ӺO�L�P�"OR�
a�Ңwȼl�����"O=�ɇ�J>�M�q��j����"O�Hq&h�q�$��r1�`ZS"OB\�c�(5~ܑ��[?e�HPa�"O�X���L/0�a�h�\%��e"O�л�f�_4\�s���u�q�D"O1��,�#a �P��$���1�"Ob��S*��%3ء0OʱP��0ʇ"O0a�G��e��<
�o�S���f"O�A��LG&Dl,���.Ǎ7�2�p�"O��c�d��G@�! "�Ȥ��T�4"O^	x���z�A�BZz�z$"O�ڀ*��L���rD�UI�"O:�BU�	�Z��`�ʔ�&KV�St"O��Ӵ�{��ͩ0)M�(�U�"O�q�.C
EƐa҆�"a{�� "O&Y�cFȂd{���1�J;z���"O�(����')'�	��>O�M��"Or!����� � ��I�+mY40��"O�m�T.ˎWю��u�]�pP�D"O�Ux�%��h ���ϻ5T�M+R"O����ˎu�� j-E�D�T���"O��K���{�j��Ti.I�H��"OxTR3�¹!����v�� *��]Jf"O�1��)�)Ja���%�~�f"O���&m�DoTu���"}O����"O���S�M�'��9�V��"q"OB ��QV.r��Ph�x-�K�"O��vG��n����,,�H�#F"O�	��I�*KT"�2�eL�(�^�2"O�ٺ�˸H?x��E%T�'��8�"O��H7�ݜ6>M+��dV�,�"Od���E�"+�V	b��Z9M��Y��"O4�2ရF�~�Z �ɀZ��A��"O���FNd`�!�՜o�0��"OT��o]7lA�xXv�6O¨�!"O^��e4+봔���T Fl�@�"O(�֌�4?��2ᆀ�hk��8c"O��b�n�:l|�}��L$�\��F"O"L��@l"�Kg��e�"O�!�+�1FTz�kt��/zbT��"O"}�D�&r�Niڣ��3[��	�"O�0*�����*���O(<��"O���g(��.�.�p��3d�ؔk�"O�X��w�YtO�)P5iQ�"O�|ti;[)�ŻA�C�v�,#E"O����a��[X��F�-��	�"O�B��d�`�<莀a�"Oԭ��oD�x�bUXq�X Qz�i�%"On���9s��0�5�H5s��*�"O���G�Ȼo��l��D ;���s"O� !���c�E��E�Q���Sw"O�P���zŀd��"&���"O���A�N(n�4��B�&)u��"O���R�� K�6a��}`�CF"O��d�[pptE�dΊ.6_�X@ "O2�8'��=i��%�N&m���cb"O2�9W���0�Ь!#Y�ҽy#"O&�`���Iq�����:ۤ��"O��C�놓Rɪq8F
�/4�:��"O\Rp��;l;,uiU�	?��s�"OUrM\:<��C�" 	�"OƐ�#&\h�Q�77���"O� ��c +���80��:4"O�l���m�����
�+֤��"O��S�7Ξ�!�h�@�!�"O�"�BF=>Dp������D���"O"@x��C?3�Y�QN��%�0�y�o��s��� ��r$�p2M�'�y��Du���u�ՙx�����CT��yr$���,����BX1�i��y�Ac�"�Y�I�	݄�h�A]��y"��#S|�����Q�\Jŋ�y̕{ʬ!E�Q'~�� �E�yr@�&i�1�CEZ�}+9p%.W��y"H��.y��ʅ�Vq�Z��4�%�yBK��h1@#E{�`\R�g���yRJ^$#v���g��	�	=c�B�9BFʕ�D��Y���2Słe�^B�*f�ਃ#	I� ���Q��>N�4B�Ʉ!�r]���C��#��){�C�/7�cwg�rl0�#i�_h�C�ɝEKj�A�� ��q"�ʇU0�C�ɡ"�J�#�JՔQ�eS5�I�r	|B�ɀ@����p�D�6�� '�� p�pB��:s�1S�'Q�j��p�NN�4"8B�I7�rdIUƒ��%"AO�H_�C�IDyx�����,P�珟;C�C�ɟ.�~�26KC���L0G)M	?̐C�1dE"�@]l���$�$r�bB�ɂW�6�h�f٪R̀���ٌ�yr���Vz*�)��X�z	��ڦ�y�iϨV�ZuJD�0Qt^,c���y�C��2�;s��u#�tJ�_'�y��W�|��裮T�f�̑�#F>�y��@.$����G8c[��"��7�y�̊%S�9�'n,n����*�-�yr�ս8`��+
�b�J�S��yRƬc���`ee�t#�Z��ybI@�tĝ��
E00�.-��oN��yrL���Df (\�a�@���y2@^�w���'<��ɡH¾�y��#by�-P5�Y� 9���4�y���*b�
��YtD���G�BC�	<&cr�#�Q/��#i�{�fB�ɕe�>�i��+z�y#�G �C�IE{��1u�9�t��g̨e�X���U(��ٕ-�R��-� �H�Is�4�W�7D��P�#ML� `���"�8�eN#�E����.��O�P�Y��S�U:�� ΍��=�
�'nK���H s���=H��bȟX��w��؁0Qy���Z�|ie����K�6>.pB�	�E���qa]���	���J�9�N˓5�vM #H�k���9	ÓoJr��Fʪx;�����3_X����+GN�}c�㋲�=b�!��$�&)��[+-J0a�F�(��I�r��㗀GMk�bEˑ=H�<YԋT�2� ᓈW$��`I|z*Y�3���%ڛ<
�(A�h�L�<A
!1��8c"��I��L�'d ��E�f��� �؄8B`�D��'�:Mۗ�'xg�-���W�}.4�3	�'���+��_��V�����2���Y��˟B:�d��eU�[�p8)�"K������/gآ�uDF�;����G�(vp�{�'ʞ�Ԉ`�'Xz��֥V���ڽy[l҂�׈-�j�'� �I�l��a�l���)O=xɑ��D�<8 ޥq����X���G����v"��"O�|�
ق4"�2�y��Ҧ.c�<�4k�y��I�q����Ìq��D	#	�%:\����^	�f�����
SX0Hl�;?:!��ע"rś�*̉a� e"&J�%X�~,(&�iR�;5D�DD(� c�~Fz
�  �3���#��{��N3$�s�'+�52GI��pw �1���un��� ���N� ��g�'ߺ�X�.LO�a~r�;,h� @S�i�^��B�	��O=#6�J;6��q�.�tS��@I?�k���&TS��7a݂<9$1D�@�v���R��|{']#����4-W
�(��ޗ7r�TR4J˸)[ #~��i�*� k��A;3i��C~Q�ȓ1l� �0,
�0Є�
$�Vdq����'C��
E� rh�C�{F{��2�j��pʑ�}BW�_��p>q�M�>�h��DX�b��:7u6�8%��Ґd�B�X���\D���U눼y�ʌ����	[x�D{�+1*�~�8&g��r#1��qaeɨi���y�(E��ȼѧ"O$Q�B��y��)���/ .>%@6�'��6�J%3���ȵ<E�D`C*��0cu
Y!J����`?	^!򤈻3�@�*ܕ>0ī��KZS�k�`9�S����<1f�U�M���*P��h"��T��L3b�����0��#%�t�z`J1@�ІȓH�P���aH��<�C���^�p��K��؇��h�CF�VKz���yk �6j7��"s$[�'����ȓq�މ���ˇ%��!�����<��h꽲�
�6~�yJ0jX=<\`���w6�t2È��Ť͒�CY�hq$u�ȓ36
�#�̩H��dڄ
ev�������c	��L�w��W��d��D?�H:d-C,��)x��P�q����+��ɺ�'��VA*�a@oM;Ģ���H��q酤R Dh�p5����ȓ�����ڳI����El��+J���ȓ��0�F��-D �@���J�l�<ya�O>��i�JÁ
�Д��k�<����Uk&h1�$�+�0!����k�<���_�D͌Mk�؄X���%?T���7�It��řS�A-#	ı 4D���D_%!.�`�&d��1܂�KA!7D�Ta�C�g���P�$./~$�f5D��R�B�(�� i��N2�
����5D�b��2 L��`M>x���$O3D�h`+0eXx9P%�������-D�@���ʠz����ǐEnm�Ԅ,D��i��޺Yr/F��>��L=D�@Y2�7S��H�oE�-_���<D�DhեX�Z5ʩ� ʁ�*��K��:D�� $O�F���D��q���W�,D��3V��Sm�u�kN.L�̉��%+D�쁂�H��	��]����ժ-D����@�F���ڡӆ��B *D�,ې�ޫTT�Se͟�R���,D��#Įώ4��ACKM�>�$l5D��ӈD6�\���a�<9 �N3D�hh�3V2����
?k�8�Z�!�D�5T4ҏZ�Z�<���O�s�!�d�#��PI^()��q��.0�!�$,�tb���g�N�����(Q=!��P�ϸ[��	<5f�ӳ��&9!�ՐC����*%�h�a�QE!�$�K�Irץʛ1(�'�!�^�BB̹�s��!���q���{�!�Ăv2p�u�� 
l"��U.ߒQ�!�d�$P ���Ǭ͞e�@A�'Ch�!�D����vΜ m�L���`΅u�!�DZA���*ߟDäA6�ҥ3�!�DS:?9c���&87<���!	�!�dS�&	���D�F���E�����H�!�Dє,t}0��!E�8\���R<I�!�� ��;b�˭?wiA0�_E6�P��"O
4(ЉW�Ov�4�Q�L41+�"O�Ր��MLE9#Ȟ�jT9a`W)xZD!�`Y��l9�dE=<OBab���5"fH��L؋^H�Ÿ&"Oڜ���%�0�`�h�Y���"O�|�P�
)���K�%}R�|�"Or=�G���J�F�ށ�"kU"OHi�%�Ñ;��Mj��E3��8p"O�a�C N-\NA��C�)�%"Ona!�?<�|$	�엿
��Y��"O����	�i�a�L �~(9@�"O�� K�;l����EG�s����"O,�"��M��Bݘ�5��L�g"O<�3e�[-W���� L�
�h4#�"OE#�cE�:r�;A�үU��JA"O�A��
t��m�7�ϳˤ@K'"O�Q����x�j\"��vY��+5"Ov��e��O��Y+��˘U�u"O�����M"gE�M
@LM�HB@�"O�T;D��&n� TQ3�
2-B����"O@x�@A;9�R�%Ǜ2k8xP!�"Oj���G��x��j�%Τ9��(r�"O���Q K�,%ہC�W�2"O��a�C֙#|�0��L*�"O+�g�<�=�Զ�+$lzC��  p����2~�!Ѕ�[�B� J�Z�Cf`B13H��� �IS`C�ɁDP>���X���v㟵4�B䉦*>�=:sB7s|���s'�a�B�	�0 yA��8WgxU���Q/�B�IX�t���C$�
8�tfPvs"B�	�Az�$�V��C����v? dB䉋fb��T�71�������Y�C䉜nJ��Ё7��XG㜈|�tC�ɥ0�b��b����(�f4p��C��$h&�9u�B�J
 )���I�MK�C�ɻ]K���H�A��ș�뇄nd�C�I73>�}ʠ�J�x�ZLK ,��>:TC䉁#�.蘲"�[v��q�BzgfB�	2+�@ZA�̯n�%�$�<,iLB䉹R7F]� ᪝�g�N.�C�I�yH��Xb��50�x�;Ң� �C�	"�X��A-G�@�X����DW�C�	�x.��FiA�'����W<j��C�	%g�rBe��{1�	�?}O�C�	OE@Hb��`���r�"�C�	6C+���	�L��@���ç{��B�	�<#Ԉ+`g��|��@��땑1�B��+���q��;~�б��Fo��B�	)�NP�S���yṳ0�	��x�B䉯Qj��9%,�4aɆm+�gˮm��C�*�,ak�Y��R��c�Ȃ��C�I�/"���I��&D��F.��]�C�I�e0�Cq뚺O(Q#��F�n�C�I�kf�}ْh	�vLmiE�H?C��2;=�	Z#o��VJlTp'�ō(�B�/J
h���"J�N�R �,F&�C�ɦU��A��� X�8��#�ߠb��C�	&Q5r�"­�9�p���L?e�C�ɬoAj��d!הh����)A��C�I0ς�т�ã�,�JT��	��C�I5Lʀ�׭ԪJX1��^"#6B�	NiÀ�ʕ[J%1GJ��J��C��I��,['&��?��ئh%�rC�)� ��jO
&��j3h�m��H�"O���ւ�2: IG'��e��L9�"O$=��L��v�P��,7b�XC"O(�`�\?���&��_�� �5"O(="E
P�� Jޅb�<ٳ�"O|���NҴ=��H
'�Ź=�k�"Ot� �))wUh�Ȑy�$<CQ"Oи�����L���B
����
"OXp��c\�`��0�N��z��l҃"O:Qx!/:/���RN��`;�x�G"Onx�`�X�t�kq�4o d �"O�5�5�G�j�n��f�\�<�T�w"O��"�,E:Un�tq2J�&K	ri�"O�Q�%�W�J��!i��[<L� u�"Oֈ��.!������%:$4���"OF �
�R�Uѕ-:�$��"OJ��T�0f�#�Thpt"O� X@CQ�~~Xy���\��K"OZ���덢B�^�Q!�)_? �yS"OD`��,�
G.�Y�	c n��B"OXL��I0*���ƀ���i��"O�PJ�E��n�Ջ�+С��I�"O�L�وu���:���!���g"O8,Jg���L���� hȖ ��:G"O���Ϟ(�DqWlA,�F���"O(X1�'T�<؁g-��.Ę�"O�����q(>ay�J:p�\��r"O޽�r/V�*�L��v�J�[0Jt�e"O*THf��f���B���62�az"OЁy��0J��b�ɱb��"O"-H��l�����ą/��8� "O�9�C&܊`� $	��Q"<��q"O�����%;Y	� Q<v&<c�"O)���˅c@=�g`�4\:�L�"O�e�gA�<��XRr
~'�u"On$ �H��ph�ٵ���nF֨z`"O^0��FC�$����7�L9���3�"O�=P�ƍ��Ҩ��m@�~�>LY`"O�$���+'�j�h��{��TYb"Ot��(M�o��E{�;`�:�{�"Of��g*N�f�0�!5��D�0��"Oҵ��%;r)���.|�I�"O0G�֛ d��q&_�Ch���"Ob������Y&�娧%�`���V"O�3�܄�H|3u��Km�X��"Oԩ�r�["!X����-qe���f"O��S���w�x��UۘOVX�1T"O��J/EZ��QP�K1GvJ1��"O����3f�DdI6NǶx�N5�"O��s�Ҭd0�҇l�Yg���"O��X"n�~�DD,��k\,kp"O�,�I�odȲ�H(]pށ�"OT��ai�c��F�m�Ƹ*d�$D���S���n�Ҳ	��*��k!D�XZt � ֌�"��Z�v��t˳+$D�{�)َ{a�A�%%�حr��!D�l0��#fB�)w��4A���2c�1D��削^[�	(vE�>�X�{!�=D�4r��=�\@b6b 7M 4��(D�tI��%E&��J��^����%D��"��9-���+B���j�ܡ�3�&D���,:*L;1�ځD@y��(D��y"O,1J�=����j(��O*D��P�/f9<9Tpʁ�2Cax��)� �T�D���f�d$��i����$�"O�L�C�"��s���7dJ���"O@�H��9*�5*�/��$�3�y��4s� �u��i4�}"�A��y��S�coT1�gȝk����ȃ�yRn:^�ā�VL�pEd� 1���y2d��i]�8�ܻ27 ]��K��y�.�x~����
�.�^��WO#�yi�;c�M�����
~@hb���y⍈�_�֜kJO�nR0�(��yr��!�lס�"RQPR��yr.R)��yh�
�}bt��+�y�o3wE�T����m�4 �A�y��Θ"��M@�Ԅ65���,��yr�Y[��<c��ǎ,����^�y��q��0Gˇ)Wy��80�E��y�V'p�ܫ6���R'. �bH���y"������;�ֈ���[���'O0����t��D	H�	�X�'�`7$P�%N:l��C�d�ț�'��1A�#���J �Nrɘ�a�'T� KQ"A#R�չ��FB

�
�'C�%S�!� �xذ���r���b	�'��Dsn�8b�X\���6W�f�#	�'�LYۖ�:ix��;� S�S���'*\��G!�wi,ջ��6PC(�Z�'�*<�˛�Z��x{��ݞ��0x�'�$�Q��L	E��vOE����R�'/�y�BAX�z���*�@��;�1K�'`x��T,�|qZu�ʿ!BP-[�'%|廅/��0i<�����FTh�'*�%�S&	��+��K��n��'M��i߾<f��e�8;��ܠ�'�&�K�$�e�.�9��Z� �U��'Z�Ũq�ī n�*�d�T���'���QN�w�ĭs��H!Rݑ�'Į��v�Nu7�1��l�H�'!j�Y�	�w�`I�����&gj��'�x�
��D�1�2Y�'˖n���
�'�2�hď�!,>X8rm�EI�#
�'~���f��9^xq��hD1@��
�'A��4���U�3�|ܫ�'�8Iؗiʋ#� ��m��Yt��R�'5f�ȗ�W�'�� 	s&ĘS"�}2�'�p�aqK7i��y�N�7Şp��'/��P���)�\ݡ���0+[���'*>,���[�Bg�x
�I�7w����'(*i��'�;K r�0`�^�.�x�q�'� X�/ްf��qV-4��'��"q�,3.�,�%��-��R�'4�	k�g;)f<y��0#bt�i�'�����$���S��Z�1�'H�����#_�Z#e�@�����'��xtϑ&k#�kRmҌf�5��'X�iä�Drp�YJ̷K7�
�'�Zm�RK�'?N��PQ�H�Ze
	�'~b�YW�X4t�X�b�:BT���'�l�j��K�AGp ����:1
D9
�'��A�W��%Wڐ#%�V�0$V���'OL���
|���ȓDۍ5����'�:I�!�����F�|��\�'��]:LˤH�y�Ӏҟa�0�
�'!: �E�'hf0U8#a
uk(PI
�'c}"�8�8�y�J�rF��	��� .L�!��]A䀠LX�~ό��"OL��peFb%4�ru�7.�ֱI�"OΈ�BFHZ����J�HV��kC"O�,� ⋌'jh��I�r�d�%"O~�A�Ǟ�9(]��һab4���"O�e��!_��s���\m��IW"O�pŦĆW���cq�Y8{[�0��"O>娲�֦0�yf�=절�s"O(��E����2��Է=�9���ݎc��{��(%��P�Ĉ��y2���_��)T@F�NPE��D���y��D�0g�ATA#�Z\��̎�y�O 8\*�XAꙪ"�z�O��y�h�9*"�# ��2`�NԨ ɩ�y�%É`B��2i��qх(��yb.�?i'F���� c�N`i�e�	�y�cԴ������A�XH�1!�BC��yR�Ȧq���C�~��ڣ�F=�yRGE�3sݢѥEJӞ5SA���y��|P�����?�Z�c�'��y�BA�<��Aˀ"��>tZ����M��y�
B��a%kҨj�F=3�L���y��uz�	y�GYS�r�JR�Y��y�B�2d��! �[�Fq����%�y���l�r(���!f2��Qd�?�y�eD�(��E��@.08}�#-Խ�yr�C0/J@�C#N�20�Re@�y���j��l�$�åx�F�*q���yb��,�h�i"s��J%���y*ߤ�4�妀�d"<���̧�yB���oxTD ��=S<�Z�+��y���0S<�CV��x���O@��y����HX`�L�n�n9I왗�yV;N���PbG�;4�������y2��w�|��X�d��E�Teϰ�yR� }?|�2��(f�<��,�y���0Q�6l�$A#3&����y#��v�Řd�(t�[����y2�B3G�Н(�8~�&�����8�y���1��<�S
M� ڢR왪�y"��V�h���b״$1��dZ)�yAR�U"�ȋr�˙o�@�(ˋ=�y)O�DI|����T�p�"\�����y�%��*(r�I��3��2�����y�Ƙ �F�	�ɇ8w֔"��4�yb�=X9�wGE,8�F�h�Ο�y�%�&�A���@��t�0�n8�y�͙�<6�����- ��-�E�%�y��5L����T�V��JU��y�hĸ+ �As�ñx��0���T$�yBdܐH��	.��w9� �w�׃�y���$a`ѱ��ܱӰ�27C!�y�H/]<���D�l>�#W�V�y �l�G��y���x�I���y�.��<d��8\��قuk��yb��l8PÐ� 2��W��y�fF�}��Bé�.����B����y�-Q�<!��`	N�j�q�a��y�ER.a�%��/@6vJe�a ۀ�yR��;L-z|p���3��!5�y���
/޶�ꡡ�W7b��`/��y	ZB ��IIF�1J�	Q�yҬ�Q��A�����v��` )P��y�.��SR���$�ߌp���2$f�:�y
� ���ECmR``�0�>/a��"OZ��,M�T8z�E�%�B�
P"ObE���	v{��x�F��B�yȐ"O6`��/� 4����\@�"O
��t �YgT<(�* �p�Q"OT]bqM[�l����x��0�B"Onٙ�ܢx�P���D�>}��Ő"O�01�O1G��[&��In�I��"O T����1B0)�%�S�X:EC�"O�����8c�C��{*�1�"O��ZG��|�,1)f��5*��j�"Ot:��	g��,@��Q)8��2"O�D�'��ؤљ%�_22���t"O����<}����0m�'yR���"O��@�L_ Um�Bc�5c\v9k�"O� �4�܋f
�E��f�،��"O��F��L��SG�K"0��D��"O������g��%���:G��8��"Ob�PA��N��b/�[ɂTqD"O��􈈵�젃�m]����a"OZ�r��-^�d��b���v��c"O����A�1��{��?�P0u"O�hP��	{�9�@B�W@ޠYU"O>|9f��� i4��#6� :C"O ��Lh��y���#|��� 7"O������NϜ$�D.ޗN�ĥ�V"O�u�4"�6��-��,�)�ƴb�"O��⧎�(��e�f�Zs�@�"O�T�c�#}��(���6���@""OT�"΁ ;�M��jɛ�X�)�"O*@�G��<b'( �S�6�iD"O�Qiu��(x�"���_	(���"O���%���f�,Qd�U��q"OfA��3	F��s�aL� ��8:"Oؐ�K��F9×m͚[ङ�"O�!�%��9uZ�`��iQ��v"O6�� �.1ȁ��*���"O�b��m��Ð&� ?�VD�R"O�1֍Q.��Yh�$C6:
�q+�"O��`V���c�E�6�x���"O��27B��Lг���j��5��"O~X*$j�e�*=�׭��L����"Oeʢ��3c�\���8"�����'�N�� b�KsPt�U�r�D���'�V�ɁHʮ|-t<��Z(5 ����'�0�o :
zdt���E�+���'g*�J�΍%)pڙ*��Ml���'�FXQ�J'8���2V�F�dN�=k
�'�v��.��D�&�K�x� 
�'�`H�B�;XU\QІ�Ov��i�
�'R���Alͷa:n��@b\�g3@;�'�j����Ԣ<G|�	p�ϴ`.P��'Qޝ	`���B�
��GL�_�V���'4<�l�[@ҍ�ck��m����'9(�"�G��:���"�z�(�	�'IZ娷�܁y:PI�Í.(|ʈ� <O ����V���胄�%�}(A"O�����9D:����G>%��zw"O�1z��?B6d8p��b��-�4"O6��@��%rʶX�t�� UvZ�ZD"O��E��2K�B�iR�q��"O|���_�t4�e�6TLE`�'g:0��JO����0����p��',҅��NG��^0�!����Y��� V̱�L�N�f��"c�������"O���¸^*d���J1 �����"OڹK���$m8�bK0x��᪡"O�T� �'�<�aKW=[َ帀"O �kb�̒q%v)Hd�W�쌴Q"O�m�����A��[%	�l��v"O`4��\�LTd� ���ZD�"O��@ִׄ �9P������B�M�<��³&"��W�w� ��¦G�<��U<#|�)4�U�F�@Y@#�YA�<I�d�%0QI���x�$��2J@�<�5Ł�<��qJQ*m��p1��z�<)tM�7��\0��&>\�x���_�<1��+^I��2�F!8K`���e�\�<9���xUʵn�6�^����M�<�׬-�|0�%fX����eJ�<1r'- fb�UnQ̅!�.�^�<�`�ְ+u&��UD� ��t�)�X�<��2E�����ʛ4Q��:�`EK�<9�CH2���h���n�t�rLP�<y���:�Ȧ	$U�x���g�<��C=�:Xy�+\p� f��b�<AqIɻ~|���Η�<�^͐�VW�<��	M�Y~�J��L�\ًF�I�<�u�Y33>�@�G�B�6j~�0�JQ{�<�%i�YO"�ѓ��I>��`_�<a��܆Q��0҂ ��.X�ЄK]�<Ib�Z�X=� �0&K;jG={���\�<J	0��!u�41�0d�d��d�<�5.�5; ѶE��z	�p��A�c�<�Bj�}����-��y�2%"֋�W�<!b.Խ ~�8h���A\����V�<Q�Ȍ ҜP�&$�P�YP��~�<Y7Y2���ba�+}���q��C�<1��ɪ�vm�pDīL��0���}�<qQ��
���£.�9)M�@I�v�<�&�I���)Ce��{6��"�Hr�<��=$����#�m3���Y�<��.�%$�<8���5&\�D�3�U�<I���R X�K�杜V�l�G�O�<aǅ�	#`<���F� �h��JOG�<q��7(�dy��Ww�4q3�d
h�<96�шY�^ ����4Q���#SF�b�<�	[9(��8;�◇Ec����A5D����H��G�$4�'Z�0����0D�d��J����6|'B}C@M.D�<�`i�YN���O�&	1s�*D�\�7�B-���V@��+%�<���%D���"m��e!(���*L2Z0�d+��/D�h"�i���T�,�,ʑ&0D�����Iu9��ÇBіi�s((D��u#�Au2Il�<BA�}5&t�<!�ĉ	 ��3�6��$�D�ȓ���R���@��k�"Ǝx��܆ȓ0����#R��̕�֢��d&��ȓ*L(��C��)C�4e�&Q)�=�ȓ5�Zez#�P(;�"T8��G���p�ȓK5ڕ���ÞBS��B�� gBR��@�3C�V�lJ>�4��eo�X��lV�%`�8O��q���;�͇� �z�� L��9��I��ȓ@��XA��P:J)bQ�\�D�2x��qha2rg�#��R��ǊM��>�n�@�e�7��,���P ��х�S�? R�xu��?0ܐY�i��X ttj"OV�qw�F?u�t<�T�޸y8���"O<ɓ�Ξ�J�25��ņ�'� 7"O4A�#��SDb����(p���$"Oi��D���De'~���ӳ"O��uH�r�����f�%7����"O4@e��2IfX�!Š�>�:=R�"O ���jN?hl�@XC������"OlHb"�]/c�V�3�G�,?��a�"O�8)�͠q r�P�K3.R]1"ODdC��ڠ�=�c�MM��;���O��B`�M��O?�IT��!��[�'��`҇�a^H�*Q�k�`)y#�A>D��8�b�E�`��>����ްh5��)E�
݈q�G���D�i��衦�ظBF1�	L?B��p�ҪOa�c?�؜&ٶ�Q�őF5�U2ԯˏ�b6M[�6���'����?�D�ܴ�]:��J}Q�U�7CA�
��?����	3oX�ip�(ˤ})F�Y$�F�<�5�i��6�!�����m\7(t�i� <W�ƽjTD�!��IZ��Z�4��<Qǫ� _@ce�[�Ȑ�R��Aӄ��q��2a�r�������ޱS��O^��Fx��˨C96�����r���`'���R(�Ls�%]62c&�:ǎD��8X��t5h@/�`�:�zuj%�^!(�ZT��jzha�c�'U6��u�'��7/��Y���	T}H5A��Y��ƯE�**��(�y�&~�H�*�씂-�����G��! �n3�M#-O�d�o�J���<�PE��u���2���4��<��b��B�$�20�ϭ��<��B��$�s�K=E(�,���GޮP� IՂr\�T���R��p�9+'�h������&�bQ�*�=F;X��3Aށ~#le;c U��d����=}䉉t��$#�^�dӄ}�QL�*t&tS0��	�,�`IX��MS����$�O��ʧd{h�āމi���:�`��6P�T��3>̒&��7��RW�
�]�����N���mj�Z˓b#d�T�i���'��ӡ�^EHQ�иo�
!Q�ힹ"�:�'K�?y���?��l9�M�aeԩU�ޥA.�=I<ڱ�'h�d؈႖�P�����n�vFz�F].LW,�yrmL�uj��c
*]T�AK�E
"�@��F(["ym^ͩS��f��"=�w�̟L�	�M�����鉿Ж��d&)� ԰��,X�x�	`�S��?9��2Zz���7,cH�QK�#�ў�&���42[��C
;����K6{Ո�{嵭gG<��435��`�_�ԕ'����O�'#�t�K vʼP���%FI�1���q���r��_�h�9�\=Wh�r����Ͽ�tON noȄ�7�����`�˙񦅰3��@�j�iEF&̤�2�n��7� (��\c�"$lG2RSś�,R	]��5޴C����IП�4�?Q���i���	��z���T'�,� ���',��d%ғD�Dpӆ	k�� ϐ���Fy2&hӘ�l�~��")�ծ;Q<�l�,Ghh��aPZs��'�rOQ[�����'5��'��a�~*�47�Ą9Ў�V�̌��Y�@'"M; �@�9��mx�n�y�\%I&�/7����Q]�'����kӍ�D�Rѫ�:.���8�JvӒ�[ /_Zn�m[�Z')��O��`S�y�>p�B��ă4:~���lP�T�H�$E�;@����O�0J���	�'�����A�	���J	��QÌ�8,O�����";�K����-�P�1�h��Mc%�i��'����O��'��&�O |  ���ݨ���ƎIznT�ǎ�;@h�[a���i�w�2�8��"��]�t�8�8��B�'���a��F�p��da��K�����A8Yg��YD�W(O�~�.�s�K�,q� k�Gf�<�<y���g�>S���Q���"G� �}&�π ��r]x�� 1�Z#i��d��"O~��֊J�6�h ��dػ��	n�����&�8t!��F�ZQ?���Bo��8��T��)I��[@�!�q` �Ʌ�ȴFa4,"��Q�"� 'P]܆TS�fB Li(%۟ўܩ�)P�Q�%
l,��rn6�O:h�0aD�w��x��ŢZxS���K6���`�( 	D�QaŶt����DN;�����8�>��a��$��t�D������$�t9�e�ѣ@G��bӵ3����f�Ƌa2쑡�!T��y�dD�H��P���f�,I��؍uK@���d�p=Bq ��A� |��@��s������-���zc֖H��!�B:D��yqE"�QY���O�@���K�Sr �Q�۔a�H1�������Sb�'v����'U7(�������'���*O���sj�'븧�ĉڂ%���H�g�(��pMZ��|HJ��Ï/(гFB]2Ю�� �'�l�V雬�(��# +ۂ%�M<���S�cd��)�<M��B�v�P�C�O��(#"[�����+@819��NND��B�)����'E�)1/
ͳ�O,g'�)��zZ��JC�Q�/���ZF��?+���?5��U%P�SE�1v��Q���C *{�UE}r�U<Q>�4#�ɟȨ`��YXP���!w(P���i1F�[�S��0	�u��r��?Qx���P	/��8U�M�G����*9��D�(qgr H�����~�HF�!�N�Ԩ�����aH�ֲiK�A̦�>��c�N;��Q�'�V�y�NW������:��T�J��I�o r*$Q�f�	?(z��*ܺCp�݋IS�iͧV�(xA&�:���'�W��Ԅ�ɲ92N9� %�]�^eY6NK�d�&0�ࡑ_���5lT�`��a��B��UP�_�����,0:pEp�) �2N ux��*��>��W2���D2�ӛ5��-����|�p�	���$%��a�hY�b���7�ǟr�)Qb�韜=G{bמ���D���Ls���~��U'q��� &X�T?�� ��B |��Z��0wKR�0E�U&Qi�i��k �r�"=��	6/F��իɧd��R�=A�rO� ��F�x����6aE�V�x1�S���ߟ��)�@G�7-@�:B����X�W�'t��9���o�`13�'��n��!B�D�����L�3RqOf�}�I���K@���h"Ltɢ�4�<C�ɆL�z��Fl�/,���C�<EC��3j�^�ȓ̖O��%�B���O�-�����4���I�]��i
F�V�"b�6 !�$�s���Z��`��\s��2�F#q���*Opűh�i�g�I�j���xT̘63/ޘ��˲dvPC�	5R�d�aǛ�]td,�����`��O4������94��Q
�I�����长Z�u��>�*A�㉧U�z��`U7�,Ċ$1O,������4�̇n��YAR"O�@��m0�z�h$Ď>�*�Sv�>���Ȋqn}�glӝkT�#~bw	]:F6jt:5"��P�Ԩ\H�<�'-?(e,��a�<k��������}�l��"f�y��I�By�}&�l����@�PCê7s��q� ���+Җ�<h�6����b,��(6]I1��%l/x�ذh؞@y��ZvA�Yz��ߋ2-��kd�%O�a��z'ޜ`�TZ6��T�}W�U:!�0Y�qK��5�Od�r�?O�1�rȂ�Ll�	��|�p5P�>93����x�R� �8`V M ���,�Tp|��HJ44s+�v�@<r%�GW<���؋h+��;�A�8������1=���vB\?��
k���X�i(��c@�FGy<����ǐ'bX��&/U�X�u q�'Xf��A���ã�8�rWdуW��d P9>�!+ҨsN(�ϐK}��Ȉ[�L�K�*���i!6ɻ�PGu��I�ƥ�j�0��dޭcHx�W�>YPjƧ	�~� S"s�չa�9�� v�:�>�K��>	D�����W�ߘu�ax�$��I��p��.�@�����L`�tˏ�+2������}Hb �%Yx�|:�@DA$L����
�4B����w#
Y0 (��x�hnĄ��ԝ2�vx"�L� ��0��&L+k�Z�c.g�Z��́laֈ���U_yZ���Vk���W%
9
v���뙽��=��G�Y���� �kӖHc�E35)e��G�x���Rӽi�t96&� ��\��O��͊D��%>7-S3hP#sL��uY�a"r����O��7b��.hİ��Z�T��V#�,��'��!D���n���g��!��<��bE/��l�Q]'S_���A'CM.Bd����铻�`��@�SW A�@M�#��=��Jb$L�"O�u�1�/L#��Ha��/X�X1��'Q8���b
�`���ɻn=Ҡ1&�P4(y|ܑ��2�����G�wp=��Z;�M� ��Pu�K,�BZA���V"Or���T(��aQ@��y� ,���I��M��k���h��q��80]4(#�U�h-�E�s"O�0�gޅk�Z�8��]x`��"z�U�����Ol��gH�
EV���M�3k�`�"OaZ��Ϳ-� ����-AQP)s"OV�+�NS�1��$j6��,@0����"O^�u&$4����ĥ­(Z�iU"O��Q�)�5��:��ýDp=��"O�仧��>r�\���e�=��"O�x�l��iT�9bN^?Y�� *"O�y�Q���M�	����'M2@E�1r<�h	$����'ܬ��-�0#%��*Х.I���	�'_�d1ǭ_� "p�g�ς�&H
�'#�`�N�&R:�Ȇ�.:���	�'�����JX�D��I/��%�L���'� 8���6Zyڠ��$3n���'Q�%�ޑ$��0���`�' b���,öo��HЪ�~)���'��:�酞	���!�AAp#,�1�'�p=�D�0_>1� S��n�x�',X�9��M�d%B)���η���(�'�V�;q���n���!շTX�;�'�����^�/7�*3e{x� 9�'e Ъ"�
M��m(� ��k&}*
�'Vj��を,	p�|�a PfG���	�'��Xxp�,}D�ԠӄE�^Df0�'����K�d�C�U2Uòл�'&z��P��XJ�R)H�h% �'��
5��T����#� L�rT��'
VĚ��@�v ��CոB��ܨ�'�Ρ�d�S1E,U��EP�8.*|��'��0�u�ՇJ��-���><\�
�'k�u����h(� "%z=dB
�'�*$R��	�-��M`M6M��] �'�lU���ՋG��8àE0�Ҩs�'�1�	�3Q�����운2��(+
�'C&@��܂o��䨆���!hf%S
�'������b�f�c�G�$��	�'�q�C�-5�pb�B݁�h��'Cܫ�*�+4���'9 �<�a
�',����lRLi�Q��'x���A�'�0�1��k$���%�x��ܱ�'�EP% �.&�ġ!�1�b�k�'�Va��%KK��uK�
ʅy�"��',0pIL�0�D� ���%p�
�'˨} ��$X����ت>M�̓�'.�9�&P2i���a�HA�>f��'t�����$<�x�tmX�*o�9�
�'ሜ���O�E�8���Y$plt
�'�|����	 Э
������i
�'��C���b|����{O�H�	�'Z�S�ə�����~���q�'�n�H�/�S���Ibd�6dcLJ�'�zؚv�°
�H��Q��Y�T)Q�'�2Ub�*�0h�`���!��a��'��\�e%��B����%3�	�yR�C�U�l�4b���誑�Z,�y�M2G�X�Bl�!	t������y"Ņ=�V=+���5#�`9@���y��MH)\����R~�y���yBLT�DLѷę9 �`q���ˠ�y�P��bͫE���M��}Ƞ��y
� �(�Ӯ� X��ǆ�_�>��"O\@2q�V ]��i�(@3x�١�O  ��M�#F����)'���k��"ȉE�>}a|N�*��}�ÃTϦ!C��>]�ȥ���V/@V���"O�{ �K�*�,����.�"�1a��ߤ3 �!���0W#|JR�ݮd�Q��҈嬭㖎@z�<�PcP�`��[f��c��3M���a 4�'`�>�	 e��z�iF�I�(����Y1I��B�I��8���\�(ሐo����S!���HE�S���Dx���Cg�$Zjv<ꃮ���{���;�AP�ؙz�����$�1�п��dQQ"O&yq �	�-��T��ŕ7f(���DžA��}�"�ёc^z#|�T�H�|�r�@�(ƶ����v�<��
���ҭ��h̹S��ʭh:t� (� �'��>��Zw,��:��d�:a��C�	�8��m�s�Q='���b�fݦG��Z�8��K�KK�i���d�PꮸR1��U�ʁm��Q�a|hT�n��u#D(u~��5�J=m�(����L�I�Y0�';�,z��۝L���!rf߿O�>]3���S529�$j��;ҧTh���κ:����y�؇���)Ado�R����BI�
���a�f-�͒2��"&C��Z��ȓ�1IGC��>i���'�B*8Bб��?��54
� W�~���T+*[B��ȓV�X��7ą�
�b��oO _�2��c�RA�C��N2��u�Y�E�L��ȓbf�3`a*S�T3o���"O�T(֔E5�@�@�-�jS"OL���NP�?�����J�#�P���"OD���C�� �� �u�3{�� Z"O��X��ރ`��l�O�4-���S�"O^\&�Իe��$Z�!��$���W"O�X�-tRY:ԀP�M���[ "O��d��dF�1(��ߧY>:y��"O��b�N��`¬�'D2\#�"O�=�4��c������ֻQ0j�A'"O��Ŋ��8���� O >+�8��"O��YP鐂C�^3 �R4�q""O*���M�o��Mn��7"O���+DQ9 ��Mч_�� �"OD0�rN��?�5����L���!�"O`�+�
��(Pl7�֕L��q�"O��1�#�N���.�2�ڠ[�"O���g��?c�hF.N�0�YZS"O���G�U6=Z�Vm�ȓ�"O��ɖ�[9�0�2��9�4��"OH�2��+8��bkL2D.-i0"O�<K҈Q�4il�TiD	�9��
O�-yT������⊼G�vx���YW�ɩO�5J�������O3"���ﶪ5�`%9D ����&v٠-Ʉ���`�5�.3Ф��'H%��*�|�gH� ���}&�L�բ�>&ܑ��Fϑ'e�aRͬ<yg�֚>@���i)}��$��y:1(P/�a�*`�\B��!@ӂ�&D���$(��H���'N	$�҆�*v��]�J�8h���P�~��'H�2�di��]��'�ɳe�ߘ`2|YS���3��"�s����e	�g�:@�F��v@�%���"R��A6�c�L��a�	�"�L��J�"|R c�W��X6f��eHte�q�d�'�T9;4�؛ٜ)%>��ΪoJ��0��f��ճd�T��o�˗I�k�g�!��ȱ^<X�z�S�n��hN�M�'�j�Q�T�TŨ1�Oq���S���.J�@��V����c�U�D���¤KA5�p?��5��9��BK�:��Y��؟(2�?qx-{@N����&�3b�DX�c'Wr��.��|�sa�"aR�k��ͪ��X/���AL� |� bR��x����� � nZ�BK~�bѯ���S�O"�q�d�� �ȉ�@�!�.��Ó+�5 �̄��S�? R1c��O2�0L��ɣ>�	R��2��ɓElpC6�3�I)Y������
}ֶqy E!�f�'��e��J@J�S�)X��P�-��]z2��`�{�D��w�Ȉf�.Lȵ�'J\9�&o�p����ǤV[(X��e��������g"� #T�Ϋ|�\Y�b�.R0�����n�:%�3���ۆ����X�$��s�M�	d2qO���lX+�S�D!� ��p��jB"O�ԩ"H�e��M�Y���Y�"O��j��_溈B5�<�4QP�"Ov�餪�4����'���$��"O=I�Î)	�����=tr�S"O��C` ��~���w"�?ξ�E"O2�a���r]*���BJ%`��|Ё"O�XX��1��R�B��q�U"O|a(�HN1|�!!M��j8ٵ"O2��RO��n/��"�Rw��y83W���"�KqO�v��q(#7O�!UH�{�j`YF"�<��qæ"OBU�*��Q�`�Ѕ+ǲ/��]yПx�KWgZ:U�� )hXT$�P��П�� �LR#9+�� _*!|��i4�'c��c�3kB�X1�i�mB���+J�^Ě@�&��0��e�6�>������~�e-=�l��B��E_��*�kԼ�OB�Ⳉ�E"hiJ��d�M�'l5`�lþ5؁�3HL��?i� VC�"�K�=lO��B�c��\���`P)��m�Z�c�O�B���L�2x�O��K�2D�ꝙSzb7m�!-�^��b�</&x�wt!�ͥ��p��um��{�B=��O��L1�܇z���Ta���I9��ϧ%S�y "�2bA�� ͍��م�ɰoq�|'�ħ�x�!*� 6c�1%�]�uV|� 	.�� �O>��D�3����!���xJ.�0�i�c]D�af�:�sO���0��b>��#(��Vs�R�#Q��a"��OY�(1���y��`��O!������*X����e2ь�j��ҧ�I�j����4a<�M3Wo��vf\�j�NO2U���"�|�<��A��
�+@�
�c�2�x��7)� Be��s&<,�|R%�a�K<]���R��:P	�h1�]��܁%�< YfBR�� MH3������%�!%wN��=����'̱Y�z�8XfFI	5V�C�' �U�)~�&��%

p��D��'��
�;�8��a�yu2�N>�&!��xw6�V�1�}�N�cdʖ�x�Ip���J��ȓY�z���
�j���TC�
 4̸�W(b�ʓI| �`��xR��h��x����%D�pxӎŷ�Pxr��(�d���M�w$�|�I�/U,�R��(8�Hb�w���C��� hҡ��#�>nw`�Cf6O�yBǌu���eϙ4�y��<��C@�/v�P<�`�J�y�.�!���7ëjB��@�i�4��IҐ��A"ҁo�ȹ��P���;#LB�G(�0&G��k\�B�I4DvP�W$�!*�&A���t@�m#4ᆧ~@Γy���!��<�3�d}w�r�K߿\T��e��z���D�?8�V�S�
�R�a �I�g����T;3���I� �`����&` s�L�]�(3��Z2
J�x�L�2uRb�c �͔o�80�b�i� �O�1���v"�{(@�	�'K>�0�E/`I�eQ���aI���,#'$5S��$,�D��U
7�� �@k��Wrv�:��Z��y2�U�R�|��dC!?u�$S��A�~�VmI� L
H2�	2D� ���S�l��d#}�?�rԳ������%Pr̍*8xV����'���Ie���,XCFva�'�*7��� J�7fR|HcF�$dXM�£;����Ub�m��$�H���$3����(����1k S<n�@�ϗ����)���������u�)�
sA>q��K��K2�\��雟����%Xi�@���N�ay�A0,�����5Fyx��\N�8���\�� I���P�Gc��>B���Ip!Ս5��=���֦27x%�K�.FB�C8o�!��T^n�S�Ԫb�(p��L�P��i`�ņ6�^�jV��<��݄SWp�S/�h~Z����ˌ^�:\k$���QZ֝����=	��]V7��iU�k�4 n+'�������7;@�¹iΑ8uĐ>zYZM��O�Ԋ	#x���&>7�� �l�A��m�����D!<��O�$�Д! N�Ɋ��;Q�6�{���X��-)�a)@�\n!j�DH���<� ��b�Z�%H����!N'y�<���?/����$�|�d<�'!�d�[��
�v��w��*��L[#�T]ӴE���My��]�0����!�M�2��I�E�m[s���>a{�f�#KЎ��2l��[�FAST`X���=�uʔ�F�� �F~�L���0!�(�3pL�� 0)ɥ"Ot)��)i'8��ae�4I�h�E����zDfDg�Os�2��^N)K��m|9��'F|5��oA�>�a◈K�~ �g�׳[����{���'g��C���R��S�P��as�'A�qz���?˂%�џ���'n�\J�gZ�"0�x�a�(
�.�P�'�`�zCk�,=��{�=���'q�D�\�Z"��Ap�������'��� �D�����@�����'��"F�͞�c���6!,uY�'A�,���T�W��\rr��	"X���'��!Ɨ��x�aFב&�p�:�'�d=�`.�*= �Z�j�er�'�EXŦ����{ K��I$��*
�'r�ԍ��I4�a�N]�=����"O��p��51��m;
��H�ԝ�"O�E8�L#z|�
' ��(�q�"O�p{��֜Z7�MqщQ�h]�@�"OȰ��Q�@��z�G�*!HR,p�"O��q��S�%-������PƄ��E"O� he�+6]А�0G��$�� �"O�=��HR�f�`�&P�#��p!"Od�$d֜%���3���;M�~��r"O���$�]�$�i��� .B���"O��*�n�-S�-�'�X�\�n$9�"O��xq��U�p��c�<��)�"O�ٸB�WZ$�V`�|h��""O��d�P*k�DMc�U 1�:@H�"O��!lF�^)�,@Nq��@�"OB�K&��9B깉��ܟm��hi�"O$H�",}�$�C!c�f��*�"Of��l��p�ՠ!� p��9�d�<�c��`�rʞ�&�����Z�<�%,���K��>��x8�i�[�<�#Cw��D���Y�i�D�R��T�<�e@r����c��-C��QWoP�<�V�K&��%�Ţ_���qC��O�<qe)I���]��G*��لD�B�<��-�s�4���j�������<AG���Gp�0��+I;_U�|���n�' �L"G [�VN1{�ei5����'欱r��ͅA�%	��.Qr�
�'Uڍ8���0q	@��n�X���Y�'���`sˊ��
]�0$ݍV�Nx�
�'t��jU�g��b1�Ի]��z�'8� j�n[`<��`�B��,�
�'��Tj$�J.t*ԣ��SG$�i�
�'��1`%�^2!ll�`�L+���2
�'���s����zp��˝�v �
�'V�A�"e�6)+�J[�l�
���'S\��5�ֆ}zL��)�!m��H�'%6	�DUT\�P�Z�Rz���'��Fy��.pP��<�d���+�`p�P�$]�T�ÁM��M��,F$�M�O�?ip�a5��1���{��DB3�ކ7�������$�0�0|����U90)�f�Y�""t)����<Q�#�>9 ��d�ʧ���Q�AH�5\x���d+<Y��ũY���_�%�Z�S>}��X%Ԫ�k�(s�2� U���,�F���~�=J��ʧ��O�TQ��<��BSwH���� �%��I�MX�%)�S�O용�E�=�J
��+<t�M�׎�>yG�0vn\��O>9�牡l����@7z��<�E�~��N�`�p�wo����3� (�"Fõ�%:�a�+Qp8<��ҬBa6X��"#Լ��Oq:ʧ(�`i�'�ԇy�!p�ǃ������/�6{Hy�W�Q�'z��ղ��O��:LF�0Ԏb;R�Ç^�&φM��D�C�:�)�#ſ|��1a�l�T�s��s��(bAZ����Z9U��H�X;"���?O��[�O���	�ra���e�S�JA#�A�	kL!��#(�N�Zү�4����@�1(!�$�94���hPʑ� ��Q��o�%!�䋥zW��2���u����[��Py"KC�nE�C�b0=�`�)�yk�1N�BTۄDX�H��AP*Q��yr臱n�4D��?�Z� !O�y�&��j-�(xtӷ?:��B�Õ?�y����K�\�����!F�Z����X8�ybn\91��̡W`B�;﮴y���y�Z�)�=`OP�0�%�#��5�yB�;	���c�.���s�O�1�y��O5-uL�I�b�j��3O_��y�`�+���[�C�,G�t���.� �yB*N�9l����6FR�x;E(�yrE�r(���%C�R�)�t���y�M�;jጹ�c.Bh�����y�$�/�:`j�� ,{i|�Y#ɫ�yᚂ��{5�AR(��KD�y���T�8��Ʌ�@r�����y�ܓo�dlÃ�M�E��q*�h���y�`ϸ4�PK1�X)P�1Y�j�&�y҄��
\f�b�
^=R)�lqu�H0�y����Eh���	C�teA��6�yb�2b���Yb��A��Z�O��yR�B%����T�+<0J��ќ�y2"_'�`�h�T)&{�����Z>�y��T��Y����5�`آq,U��y�枏O(��"R��'��5��i��y"�@�wvi�3�@�{=��1� �y���<���q�������n��y"�C�c��2��W�rڎ)4"�'�yr�̵hB�tc2��n��= $���y��� �l)c@��^�֍˓�̓�y���,�҉I�&��Uz���&��y2!Q�r��}�Kճ��%!���yBI��h�0�LZ�
��Ĳ�yB�l\��w�U� AУ���yr�N1H:�}8�ˌ�L<]2�G��y�kƦ����׊���=��f$D���)O0N����&�'>�eK�-6D����K�2� ��1�����3D��:sJ�-s`E��\� y�L�,D�8�C�6*��;a�Y� ��X*r�-D�L��t��M���ˀ Ѡ�9D�v�]5�\��b[�CF��&6D��`DO�o�"�1V��v�&t(4D�X;�(]Z���K�=1^xn0D����F�y�q0͘�1�1�-D�\;���:`��욼i����� +D�@k%o�e0���j�J���(D��K�Η5<�~`X�ⓧ=���z��:D�H;�M� {F�
p����j`e=D�<���(%^eA�AΖ���*�<D��æD�+/_���9�l�#l:D���"@D=X�C0	B�D��S�,D�djSW�1NBWAϟ<�����)D�h��'��G�"l�g!=O+(��F)D��CA�L��p(��7��1yB�9D�D0W�ɠg�D�r�ݷ~
��ِ�6D�� (��t��!V~f�ђ���8)��"O`XC`��(�x�y3���8n��S"O�����'�	r�I�1�"O�\J��I�_ۂ��am��.� ��"O찐T��?-zT���	N��5QG"O6Xro &��8��������"Oܹ�T)3�X�j#�9����"OF�A�뜭�8�$i�;�"O@IK���(IR��Q�v�V"OlոL	�T4���< �T���"O��P��O�,	��	�*0Dt.��U"O���S�l[��0��Ccδk�"O�Z `ÐB�({���+\��A"O�H���P�I��Ϟ�"B�ȡf"OBq�U g����A��Ch,�u"O]�Ѩ�XI�����-k.���W"Ork4�� 9J��wk��H)0�R�"Ov���L@$0.�%ᱤD*��S�"O0Y��%�t�g�g&P�`�"O�]��e��X�Rڶ_�q�3"O��z�o�� �󖁈 C���@s"O�\�r�΢����z���g"O���R��h��kԉws^��"OB�S�K.	���/�`Ib=��"Or�b&@��g�R]�O��=��"O&0�W�A�q�����g�8  "�:�"O�dfL���i���M)Q��K�"O4	 ��c��*�Ԯ���3�"O�hP�@
g�F�sb"V)^@�JC"O�a��)��<(J� 5!�Tx�"O�u�H�
ZbX��	�d*�:!"OtQ��� ڪ|"�M�Ch2L��"O�����iq*  ��Z%/K4%J"O���D[�l$:x�Fƞ�8b����"OHe�g�\����P��zI�"OZ$AQ"ЎN��Ax�#D:�(��"Ob|��'X�%�V0  G�p�'"O ( �FF�)Ƣ��` ]!��Ab�"O���RbM�!�Ia���Yq��� "Ov�V	�/9*�a���POdh��"O��coםZ�$����O��6"O��8���]�3w��/W,!s�"OL@2Z�=d|�В�?m�)��"Ot�T��&}�.����%�5{v"O$���- ���KA"K���"OL��$J�3��Y�d��.ג	"Oxai�[0��GCL�@�DI��"O�q35I����bs�O&A�D,�v"Or����C#*>�Q ��Ӂ( ��"O ���d�!B��-�����HQk�"O��ET�j��Ӏ�>0$%Z�"O���U-Z2�i["����ٲ"O��� �|S��DM43�J�
u"O�}��.\2"c�7D�lY20"O�颵'�3-���Uh�9E���i"O�$$^�R4>q��'�3�`s�"O� �m�
y��T�7���x��h�r"O�]�C��
&�p��X�h����"O�A�C61��2Ρ~{R5�0"O�D	����h���� 7c"��D"O�qJĮ֮Dp��Zt�J�mP���!"O�i0��3(����+�'�x8h�"O*�0�ǡ<`�H!� �xB ��"O\E�V�8��a�!��Cj�M��"O� (%�e��C��	�C�;8��S"O����F��~y3!��U��M�D"OB�(c�ά.�bP��O_�X�i""O��s"	�8r�#��L�iXa"OH�I��(%Mf4bU�/bZH��"OЭb4�
�Z��\є�M�n��S"O*�q���
#��{�B##܈!b"O�4 (T%FŢ!�1M�$�����"O�h�C�ىZ�h�p,�*xŐ ��"Ov�� �$�'�I
F�4@C�"O��r��?Iih��c�2.:�	2"OdY3쑔%N�(!�I�X%�ͪ�"O�M;UKLj-�Q�;:��`1�"O�̓@��&�.��$Z35��x��"O��2���@}H iN��x�T"Ohi���Bo<}��hS.VmQ"OB����Grt���pY�"O���#oQɴ�I�b4��]ru"OԀ8�fݮ���ʣ$�
Ύ��"O(|Hi^�{�8KUH����a"O8x�F-`h�c�̦x�P���y�Ā,�x����ɬ	d��؄����y��̟`�ei��
< Z�̵�yb(�9!z`Q��"��s/��y�J/s��I�P$R<�̹;�%�y���@Xx`�:e
$E�U�ƛ�yI�&<�1 �lN�Yu��@��?�y�e�7	���q�C8%��Uhs@0�y�.�lA����45�x2sk��yBD�4�n�X�/֣��#�����y�h��qC.��+�-
ӄ��y��"\��1;f��5�%CG���y���+| =aǀ��QY %��HԎ�y��9^��8!
N�=f��+����y⩀���̱��2�PbdmL2�yR)�
)������6;�&ɸ�+���y��@ ����W����"`��ybɚ�)0Te����5|FL�@�	���yb�	'�zi���v�^�:����yb�P51�̈�- m��p�͈;�y�ș4� ��'N:�U1J���y����i ��U��,0,�ɔ֩�ybɛ�F�@Ż�aE�*�����
�y��)��Lp��W>(,:�����yr'7��z�.ݻ��Ab����y�lW�R��=��'>i=fyr�$+�y2*�^@T�bA�w��!-_�@��mG�di�X6vE;�CQ�+�虇ȓGa����և]�j\��Ɉ/=7j���y��#� �����gY]�v��ȓ�x����ܬy�B�1���j3�i��M��i�gͪ.Qd8Jc �3�d���h�=ۥ��U�DZ�\� �d�{�<�!`C�8��$(�MZW2N`�w�%D��"� \j��T*�g� �"v�%D��	LW7G2�Q��Lj`��j#D��b�N�A8���C
F�Y��d��"D�D)�m�tD�a�E���<+�+"D��:c�Js�@��ʎ��h���h#D�XZŪ@|�d,k�hH�LbF4BEK$T����'��td��	�T���u"O�2�!dI�4@a�Z 7�Π�p"O���T��� i׀G�1� �H�"O�<8�-�=�hĲv� ibN���"O� 9�� Y�y�R�]�d��ɘf"O֍a�'L�zDD�t��I�8 k�"O��GG�7S ����e��F���"O���#�N2VHifD
M� �"O�L���ыmc�Y{���ZF� k�"O���℉�cϒУ�ʚ]�<Y;�"O�����BS�ca+Y�?-Z hq"O�`i�
�"(��1#e�Q/"�5(F"O���^27x������)z �"O\   ��   �  /  �  �  �)  !5  k@  �K  �T  [  �e  ul  �r  y  G  ��  ۋ  G�  ��  ��  N�  ��  �  ;�  ��  ��  	�  ]�  
�  ��  ��  &�  ��  ��  � 9 � � 6 �"  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�9�x8�� |e�o2+̒Ѡ���vaz���O��8�[&&$)�ޭiJ�:ǎ~���	Cx����ԊE ԁ�)�p8�k�>�����$ʌ{B��/���2e-P�n��%g��y�B�v��`���<��tρ�yR���,�wI6d���1o��y�FD? Xp��T�ԥ�1n��(O���D� "� Q����
7�<@��A�<zQ!�	5t����W���<&�-b�@�;�B�ɞ�H̻�kB�9d���_�Jؼ��$�O�c�4�C�
(�<��쓧aɈ���8D���K�&6t^��Un>{Mn�yRd1�d<�S���\��@��e}P�2.�=�v���6����I2cS,��&��:z����y� �+X�$"s���m��	iܓ)���F��#^�.J�e�u�nԄ�k���E4s�D�6fٓ����'2ўD+�"�٨Z��\q"��*o68H��y2��'"��
�(|B�FJ���'��{�Չ8༫��V������
��?�ԊaӌyZ���k-�\�dG�MJ5��"O2T"��Σ.�B�C5�6x4`��D�'Pў��"��12�Hҷ#�ui|x�t�$D�0���� �BMK�EVNfHqȡ��F{��iC��FhZe,Vu�]BD-I,!�Ą�4y�FR�\?����S�?�qO0�=%?��@�e6p�i��7e����4�|��!8�0sf�O�,}K$~*C�49i\��ה1��Ɋ�n
�<^�x"�I�]'$��iغ]��=H��ʟ {B�	3YPI�"��F�di�&	�Z�C�	FYrUh�ڵ|(0q
H-�C�IpE���ӭ�0p�N��`���HB�66d�{q#Bh�|c�J��d9B�	jNm�#bN
�����"9�C�	�r#��0�����5� �>@�C�I�b֬�bM�:ƌx�rm_ >b�C�	:P�4b�^�3�|��ӨɊ(��B�	�*}(�JJ��N���(b��B�	uA�b����X؀⅘ � B�I�l"��P�V@z
4���5DüB�&j��kT"D�iP��1��%�B��.�ҍ��J��i��-
`��=�B�I�Fv˷�[/>�A)�%�5D��C�ɜY�&�8u
�%w�HeB�K��5;�C�I&
����T<Hi9+^�y�FC�	<p��4O35�@1�h]�ZC�ɒoP6<q��Т=�f�a�]#^ЄC�ɢ ^���.��37(�(��|yVC�	�Oˆ�)�,�+��kTU�8I"C䉕*�����d^p�s�nS7;�C�	�?�(AD�ȿ;T�@TL��C�ɤ8�P�A@�#kU��B�Q;�C�		gN��Z��Hx��L�ƏA�,�C�I0U�d����'��5#ȟ�:PC�I�>ъ�!��M5%iL����P *�:C�	QNu95��	��m�D�ɪ|�XB�ɐ|�,x�@X�{�u26cC�B�NB�	�}H��J�Wr�TAD� �"�XB䉩ߠu*Tf�;O8����H��CB�Ɋa���󢌂�qtb��O��C��^it�r��u�(�OM� C�6h}����,��P{���C��B�& ���23o�����%�FH�C�)� �qR��ToJ#W�����"O~��GV[rD�$f��xA�Pz�"O�a҂d�)Y�	�gK�Y"a��"O���'^~��R��I���!"O����O�z�{�d�/V9�"�'��I͟@�I����՟��Iɟ��	2S6�T��A��$lR�΅�<*���	�d�	��<��۟<�I��H�	�����3���CU>�`�(�#��I��� �I͟T�I�X��ПP���`�I�Ȥ��,��9����5O\�'��e������ן$��矔���L�I�t�ɸ/�4P��n�h ��/�������O��d�O���OD���O*���O��$�O����ۘGo�s���:�r���O���O����O
���O��d�O���OXu4��Pg�1��
�R>��3 ��O���O����O����O��$�O����O�p0"��	��]�C�Nr��Z�m�Ol�d�O��$�O��d�O����O��$�Op�S���7�"��kO�[�P�ª�O���O ���O���O����OD���O��f�ʯ��񋏫"=�����O����O����O����O��D�O����O���!+X�-ڂ�X�cU�݅�	5�����O���O����O����O:��O���[�Pe�e_�"�x�{���������O����O����Od���OT���O�.�ddX�� ��6�:��1bV#w ����O����Ol���O����OD�m�ܟ��ɣ:7lxȷJ��8�X�`�- v��+O��D�<�|�'3�6M�<& �d3&
�q9� ����L����܃ڴ�����'"B�_�,��)���]�bY�� )ǘ0�"�'�t�
d�i:���|j�O �x�R�0ŋ;��H���L��:,�<�����"�'`V�4,��xm|�`��D�h.�y2d�iC�t؈y��Ϧ�]$^ �y0� *HЃ'C�2-��E�	͟T�����g��7�g��
	"U�6L���@�k��K�iy�Γ
J�H�z����'�dC�D��d.��yǣT�w��ѝ'K�IO�I�M�w�{���t� �H�����o�i�AI��*�>���?1�'{���y��Y��M�f�%��l���\��?�&kډM)2��|�6K�O0�[�`4�eB��a�
�Kt�Vq�BP.O�˓�?E��'�Dyˢj��\ъDHVOG�MJI1�'�B6-����	 �Mc��O�l�"���1e��R��&vrx��':R�'X��Ƕ�����Pͧ_���DO\r�@E\�&��J�
XӾ�%�������'H��']"�'ވHh�E�{�Ƒ�e����� �\�
�4ubX�����?�����?i���
t��Tȇ�
' �`L���\�i
�Iޟ �	]�)�o���H��T�*������t5��C��UҦ�*O����m]��~|�^��K�Mѫ5��ل�� �\U��N�����ןl�����my�n�N! 5�O����E_a3��!IN��r!�O��m�b�vd����I�����$͹�P��V�P�^l�@�恉]��$n�}~��.<)�vܧ��� a](�zR������@��<����?���?���?����9:��-�S!�>R^�3b'�u�2�'�}�l81��?-��4��p�v��̆+_�aHs�7@pIKO>I��?�'-�H}�4����0�JWUF��X�iN�n����ƦJ�?eD?�Ī<�'�?����?��lI�B�(q�ō�A3�)�G�>�?�����$�զa`��쟌�I�ؗOи�Xa	�%F�
�Zp�L6d�%y�O�T�'�'�ɧ�I�^)��C�ҎG��&�#t�f���"G,<D@7�9?�'����w�Pe�T�"c�-}"�􆐥ehv��I�`���X�)�xyo|Ӻ@�񏟚Zv,y���a�ԥ�]������O��m{�fo�I����lG�	JeNZ}b8���hݟ����u,�ql�p~2���P�����$ݔD�(��܀G�4麃`׸ ��<����?����?����?A,�ʉ:�B�JDF�J�'?�V�8���	B���t�	蟌'?}�I�M�;4d�Y'�oE��t'G�Iټɓ�O�b>���cS���3@&N4S'<L�3�i�a��@SUb�O*=;K>a-O����Op�a��O�q��j��D�x�E����O~�D�O���<�s�i�ƄAb�'�2�'���{�*@4���C�l�h�`��SP}��'tR�|raZ�z'P�郋�k܍�H���$2<H���-�1�.h��(�,����}��)��N���Hh�,��0����O^���O��&�'�?�wB��_a�m�b\9������.�?�7�i-��"��'��f�����7<��h5B�4��*�c�(�������I���rG����'��!�����?���a�\����`��S��U�"�'��i>���֟���ޟ��I��1��âBy:A� �ǣ�,d�'͎7�<W<���O��0�9O)��Ĉ� v��k1��4w���ْ��F}��'�b�|����sJ�"�3��y�cė 9�$m��Ē���/[r�M��� GB�O�˓#�����X�sn�XAG�>{�^�����?���?i��|�.O<�nZ�/���I�1gn��b��$]��1[=�h���M�J�>���?���"ŤgFH�D���o;r|� s#^�M[�O�=PDB	1�B��d��� ���`(z�l�:4c݃_�bcu0O����O��d�O��d�O�?�і�B>>���k�vXx�e$�ݟ$�I�0xݴk��`�'�?Q�i
�'nlb���T�l�k$,�8h��A�`�|"�'��ON�|�iS���EJ0�U�;�$�BDlL�9�p���LF'`��7�ĳ<ͧ�?	��?�FL�h��yelN�A � �/N�?�����D��Ǫ����	��O�R�2vK��W8 ���aȗY�U��OLA�'�2�'�ɧ�I�9d"bu+�mM�|��
���
���3'"B;J��6�'?ͧ�.�IB�ɥ u �T�޹��0j�����ğ �I�l�)��kym`�,A���	�����r Y��8i��G��I�ʓ.i�v�dX^}"�'��30@��v��8�߷X)r ���'rF�,(G����(PA�#&Mq�>�0aY�-{�
cFY'8�� �0<O�˓�?����?��?���)W>G�XkE�V�My�XB������nZ
x�����՟���n�s��2�����Va�f�cC+ݢ��ԘD$�?���S�'J�$̘ش�y�j����T����LC�����\�y�hˮ/3hm��䓛�4�&�Ā��6t[���F�̘S�ӎX�\�d�O*���Oj˓2���&UZB�'#�܀Ch8�(WJ��Ѕ<uz�O���'���'��'G"�i���T5��FF�t�b�On��r��8"8�8%�!�I�.�?i%��O��ZS�5��6���ޜ�ӆ�O��d�O��d�O��}Z�jB<"$đ;td��=x�J���` ��O-"��+�M��w����48�n�Pq�Q�o#�LЛ'_2�'b� :��&��P`T�ۍ?��=|�nis-�GA\�Q��rpȓO^ʓ�?Q���?����?��J��1	�Nϑ�BD�V���|�:�-O�8n�,V�'�"���)�&8ʖn/J��=�m��[�V��'2�'ɧ�O	���΄&�ԅ�`�N6�d�E�["P�L@R�Oh|I�K
7�?Ѥn5��<iw��=��bF�@��Q�����?���?����?ͧ����=�g&��W��77�z%eN�� �D�o�0�ش��'���?���?��U�(M`��mE���aB��{(�̫�4���	�g��}`�Oq�O���,j��9)r�ϗ(�t��eߓ�y��'�2�'Cb�'����B2%��E9���\C $�V� �V�$�d�ON���Ҧ�z�q>E��,�M3J>�rO�$K�&t�'��	=��DC��A]��?A*O�1/q���*��MRƟ�Q�:�8C �qNA+�ϛ�$g���������O����O���eN*m�G$��0�y#c&ِ[�f���O�ʓG�6!�'�2�'��\>�y0*�Ed��(4��:��@rD�:?1UY�@����@&��'$x�9c�����cG�6�|qJ�'�Y�T�۴��4�v1B�'~�'�K�<�����8~L����\��?���?a��?�|/O9n5]�X+ĆC�{��ٱ�[�rXP*#�HuyB�x�L�豮O��$E�I�"���\�dP!�Q<0���$�O�m�i��z��:u���@�O�b�0$���F� LYriS�[3D�k�'���x����8�	���	X��ˈ1숩(Gˈ�/'�Yr����6�Z��l���O
��6�9O.]lzޑ�#�Q�Ov��2u��:����m����Ih�)擟u�fmZ�<�!
�r�8Pr��7��LɐØ�<9�	�L�t�������4����O	%�Ȫ�D:d�F�Ծ�����OP�$�O:˓�F陳Q:��'M�
_g� ����:Gc��P���,�O61�''��'k�'��5jТ_�<rNh�i�vF�J�O朠�I�5{�6�&��k����O5�SD�h�{���*���7E�Ob���O�$�OF�}Z��LFN�9�KT�v�RX*ၒ�,	Nݨ��b��V E�K&��'�6-8�i�	{Q� �s��m������f�
��e�0���H���`� nv~2-ǳY�����G�ո��o�}#�	�P<V0R`�|�Y�b>c��*�AQ� ������Ոn�eh5&,?�ŵiC��j��'��'���
 ���.� �رgT7�d�Z�Ne}�u�4��Ş����"mN%ȰH��I�t�D0�M�$P�,�%�ӌ$�d)�Ħ<�`�	�y�z����VӾr��ǭ�?���?����?ͧ���J�m����ǟxr���=��@A�A� ���w��Z�4��'8���?),O�H���cjɢ�A� =qƝȁ�ɝx�"7�6?w��2�L�I��䧶��B	�1蘨xЍ�����QCÍ�<���?����?���?��T�Z���Lj!̎"ܚMp"ۍ_ ��'���q�~Ek૤<�b�i��'eH�;SS:�i��Q6|ݢ! u�|��'��O��hr�i��	� F���q"�l�����[OȐ!�
#��5�D�<y��eE'z.a�2!��Ths ���O��nZ���i��şH�IF�d@�&]�Z]��,��:\h�0C���$JJ}2�'��|ʟ� ��Ć���9�Ҥul���YL.IC��oӨ`���thc?�L>�1�
AH�C�䈑8�~$�⇖��?���?A���?�|z*O�Dn�C��*FgI�j�Hph4�k��� �\��ɣ�M���>��U��@*���Z\4��S��ZX�P���?Yw)^�Mc�O��P^:�ɔ��� �}P��ЛI$
�F,h���v3O˓�?Y��?q���?������0q"�"��5q�r�R�ʅFK@nZ�
Ƕ՗'YB�i����]!J @��7L7BňP��F+x��I��h'�b>A���٦�ϓX%S��KpV�4�Bk�@�T�����O�"L>,O���OB�J���^l�s婜2�>9)5��O��d�O��D�<)��iS�����'���'�\IR�9,<a��';U�����dYw}R�'�B�|�� vFҁ;��<e6�+���=��$#y^E%'e��b>���O �4�֐����Gg`tA��D[,��O�d�O�d=�缃צl��tD��?�>@�2�^�?��i� Y��'\�o�<���-{�
@Z��1 ޝ:Ӈ&���	ğ8�iyo/)��o�v~B�L0L����#��U P���l�� ���,pH>�/O�d�O����O����O�7�ڂN�Q�VM	 c4���O�<Yd�iB���'=��'��O9�ȉ  y��I�
D*[3��ɂ@R>h���?����Ş��(��P
=JR�3��	݄�@��	*�M�'S�H�& ��4H�d/���<)��=��Й�*�-W�:-��m�?�?I���?���?ͧ��X����P�����] �Ճ���u5p�"���� Zݴ��'v��?��ӼV� tt�9LE#��e�='�0]��4������Qa�O/�O���G�/7�Ukg
u&R���L�$�yb�'���'�r�'��	S8!$>�J���4p�Z	k˖_i8��O���Ʌ
m>m�	��M[O>�� �clQI���+r&�г7������?���|�P�Q�M��O�n�,I$)�E(3=�l��⑸�T|H���O�1�I>i*Od���OB�D�O(�ˣ�9���[�J�Hd9�@�O���<��i��Y��'{R�'"�ә!���i�֝�s�Ք}��U��������R�)rV�P�Z�b�y�F��PT<�K�f��� �� �LiP@[*O�I��?M ��+�����^�\���:|@&�d�O����O���I�<�Ǿi�P�
�F���Bl�E�\)��
��|�2�'V�7M=�	�����O� "VaR�F�	�OXts�!U�O"�$��`�*7�5?�T�Y�Oè�Sqy���^݀���ԑn�pq�R��y�]�d������������ �OU�8���ŠHQRay����2�gӪMi�O&�d�O����$R���ݛG�z�{���7',�Qcn�!+����ܟl'�b>ai�+�̦)�x>�M��)(;��r��Q�G��h͓l��B�C�O�qL>Q)O���O�������l��H�J�-��i�#�Ov��O��d�<�ǱihdLB��'���'3��PW��	�ư�4�?M+�$����^}R�'��|e�$N��SbQH�\8�����Ģ>���Iv�~�l`$?Qs��O����j���s�Q�if��+�Ȁ%"��D�OB���OP��.����N�|�H�X�!f�z�qfEK�?�ſi눵I�\���ٴ���yW3:�����k_�%�L��G���y��'B�'9��R�i��I!S��m���O��|f��Md��`�Ig�����w�Gy�Oh��'!��'����f+���EjE�ؘ:p���X�剸�M�����OL�����^-�~�!��n��� aD��Д�'�R�'+ɧ�O��q�%II�V85`�^�:�IQG@�rɛ6����%����!�D�<�H؁eE�CD�D�I������f6m�O$�$�O�4��˓w��7����,HR�L(��U5F��+���y�j�z�x9�O����Of�$Z�4B�< ���l�>1�e�`��$!w�fӼ����ƣ��>M�]�x� ��S�$1#� h���c0��͟���˟���ߟT��o��B'0�;ä��C��� �\Q�����?�-��&n�7a��I��M�J>��.��k@�\B�	5�ʠ`GlW����?a��|"oى�MS�O$��oN�? �����6#zT�4&|v����'��'g�	�|����	o���Ж!
�B�<$�B|ī���?��������̝Ɵ��I�|�O��ɨǇ� &��q��bI�p�\e��O ��'���'tɧ�ɘ!6�`dʈ�i��Kg��(ߎi�c�ߐt�p�˦���S=!�2M�C�ɪH����� ����CZD`I�I�����ɟ��)�Ny�nz�F@Q�!^�~��S��AR�d�g��$�O��la�3�����5GT(:�Bth��K{�M1CFGvyҭ��;�������-ąI����FyBn0f���"`�Yh�/�yB^���	���I���	ȟ��OK������L��3�t�� s�����"�O����O��?�Q���3@�e�zЁ��a@X�MQ*�?Q���Ş-�R)X۴�y�8���˙?zJ�<RQDE+�y��*!����I!�'��Iß���*9��@ Ѩ�T��Pv���!}V���̟\�	Ɵl�'u�6�X�!�8���O��dZ�,��J�e.�X�"̄=]���2�O"�d�O\�O$���0qRJǢu ���,O;~�	�E�����*|@i%?��t�'v@M�I|�aU,�,XP���Am�<=t��Iܟ�����	Z�Op�ͭ��
�n������St�Ҭf�����O*��Cߦ)�?ͻ5]2�bq̖4?J=XDl՛�>l��?����?�â�0�M��O[�惴��� ��)'�H�l)$�3:��
��"���<���?���?���?A�l̫�$4s�F�3|���D�4��˦�
������I˟%?�	��h��Oq�R�:��M��O
���O �O1��}zS� h�s� �)=�n�Ȗ�X�$���Y`�����(I4JL��A��ty���m^�Z5��#B((kT���0>�b�ix�h��'yLd���E	J������H2sl����'_~64�I���d�OX���O��KF΄t�Ʊ�b�$��I�Þ
4��7-+?q@'U$���j����:¦Q�ժ5���M�iJ=�A�p�P�	۟�����|�Iݟ���0��d�R=���V�T��댜�?i���?�B�i����SQ����4��[ڦ��ׅW�r���+߾0��Mm�	0�i>�YV�A¦�u��W<!REY��è2��g	�"V4�ca�'!8�'���'��O��Kd���˨�B��9Gʨy5���M��n�-�?���?q+���� 
�������1"邃���S�O����O��O���DW~лF����zfCA��lIt�#_�d4lژ��4�:���'��'�<�ꂉƭJU��Q�ꉁN;��a�'�B�'���O��ilZ�9n  $f�:�l0@!��x	��ɡ�����I&�M��r �>���d��hX�-��qHn1�a�ߧz(\K)O��Qիjӂ��꘠tJd�Iߧ��DP�lM8�rTo�w�,��VB��ģ<����?����?!��?9/����	ծ/ �}9r�ĸd���)4D�ͦ!�U& �������
r��y��*X��P��G�3U�I5O��d���'�ɧ�O:~-1��i�$�}H�L �ǖ�C�-"TR7Ee�D�rH�
�'��'��	�����^R$x�dػm;fHBu�8mN�`�	����	�ė'��7-Ǝ;2^���O(�� -�1
�Ĕ20H��ℭh��2�O���OX�O���<"p�Є��wr��F���b�
C5I�d�ZM)擶vԜ�0J��.I6�QY��Y�''����ѭF�(?��M�ev��c���2�3���ϼ���f���x����#_`�s��S4֘�T�D,�m;�
��{�*Z6B�����˂.V8�A���Z51�fa�P�ș`��Q
�^�������L�Wi�&�ȡAu�_?%�6��шÏL�.1�j�tM	a��*lTAP�ǄJ�Z-L��4
D(�Xت��D�z��hb$hM?�x�!"G�e��+�4|�:�1 B�$T��R�E}��JC�ڍ�M��'�Z�h�_�Ȕ'��|Zc�Y�FP_��ic� ��-H�O ��n;���Op�$�O��KzD�
�� !R%�	y��u�&�ք}��Qy��'*�'���'������wX�x���YQT`G	0H2R�p�	̟L��Hy�7D�p�S.��l��� �d�I�⊫u)|6M�<����?�=j&[�'���w�[*��I�͢5㢽өO2��Or�Ľ<IQ��C
��������m��}���k����f�0�M;����?1�M0�T��{��0�U�&j�p��B�Ǜ�M��?�*O�!�a�G�T�'?��O�8l1"�H�:8���Q#�pXZ�Q�I-��O��d��JL��h��z�xɡ'�'	o�-i�)�1x���mTy�GP�NT�7-�O��f����q}Zc,�py��ӾY8���$ГW�H��۴�?��WJES����Ƣ`d�5莦s���"���	D�*�# 7��O �db��)�`}RP�� ��V��P���&��A�:��pcY+�MkC�%��'��:�$V�
�މ� �Hr6��&�\��l������<���1��Ĩ<I���~"P!$���' 3�8� �����'�T��|B�'���'���P�$�2���$㌲Jc<͉�kӐ�	(����'���ğd'���&�5�BꅦIP�R$+�y���g88�zH>���?	����DL0���PB�0=
"�����m>x�B�	N}BY����J�	���I�v�������DV�A�,�<�.!��c�Z�ӟ��Iɟ��'�bE��r>@&mПZ�>�[d�	�L ��dӮ˓�?�I>���?)0�� �~2����S�42��V˖����O��d�O��@����R?]�I�A�!Y��D�N�,{�\��@h�ߴ�?�O>���?�'�DB��X�+���w�����hif0l�ڟ��	`y2�*\���'�?ᚧb���$�l:��"�&�B\�e�'E2�'�-����?����^�ԑ� ��J00�ǯ�>a��Yi�]J��?	���?Y�'��� ��s#�R�({��	G��CG�i|RZ����K'�S��'G���5	̛]��e#t�R��6�_�S�@��O��D�O�)�<�OF���+Jo�-Jߐ��#�y��,l��Ex���Q~!V����-���
@O t�$�o�����ԟ�A�G�dyʟF�'�Sg0����!댝)^0H���"V˱������� @s��1җo1nd��v�L�D����˓I���N� �5L��K�T0�%B�}���t�x�͔;��'�r^�D�	� I������?a\k�f�15D����oy��'V����O��I�z���z���m�ܙTi�$i�7I�"����(��ӟ(�'=��@�x>���Lm���7�A7�`m�0��>����?�L>�(O��O����	M@��mG�`/�=����l}"�'j�'��	�]��M�N|be� �س�*Ʊ��(R�l� B}$c�i���'��I˟ؗO��Z>�cU�ӳF�4(���X�p��Ǭ�M�����O���ɹ|����?����qcR�jd���ͥA�"��H�b��۟@�'�m���f��ūF�6/r���9zbX�Q�i��Ɏy��`��43���۟L����Y�����5�I$v�m��!�^ۛ&�'���'�bi�~�-O��禅�fE9y�q#"��a�B}9�Hn��)���O����O���^�S�tE�)��j�DDJ�,ec8��YN�Ex����'��5���$������2�h`Ӵdi�|�D�O��d֋o�f!�'�������9��ň_�#�~���.�K]8oԟ��'�*|Y�����O��D�O�� UG�Y��%���)�� �B�M�	�z��u�O<ʓ�?q.O>����{�,q=�)3F@�]!��a[� �aq��'V��'�1�vUBņЭ��$�㞈Vؠ�5���T����D�O˓�?����?�%bXV�֔����3��k�es�i͓�?Q��?i��?�.OmёD�|���v�T1+D��6L�YrcZԦ��'��^�����\�I��(�i��0�GX~hx� �C���@�>9���?�����S�2y�O��Gع[:̬cd���lW�kP��<t�,6m�O���?���?����<�N�T+�IN>���J��H�gӶ��O^˓$��W?�������#9ʆ��D�H9 �l�aAH9c�6h�O����O��K���<�$�?ݻb/�(��I8�hQ�j�Z�HF�l��˓X��Q��i���'��O�Z�Ӻ�U�7\���.���9�d�Ϧu���PЍy�X��5",�9`w�D�7'�D�'BKF|7�»�P�lڟ��Iߟ��4��D�<�@���K昗�l�d4�)P�$p�m3�4/����?�)O(�?��	4s&dd��A4_�8y�3W:J��ش�?����?IT�ɕ
�Ity��'����[a|RQ��.`m��h��A��f�'(�	Y0��)���?�O�NzBlY�lR�9�b�> ��4�?�"��9[��IkyB�'��	�֘1�>��aH�M��Ai`�,gOr�������D�O����Oj�'H�S��H{ڀ�X�يrx\�񄏎���<�����$�OT�$�O�G�M4 -��R*Zg��9�K��l��$�O(�D�O��d�|Γ!~@���>��ey�2i��J��kX��&�iG�	���'F��'�2�'�yZc���� Ozi�Љ�5)��UH�O��$�O<���<qS�O!�ǟ�ׅ=܌
Uʞq{���d��.�M�����Ot���O
�g2O����@x���k�N5��Y!/$�)3�~Ӏ���O��E�.8��\?��Iɟ��ӂg�Xp p-��O jH��΃-�U��O&�d�Ov�d���D�O����O,�S�F4��2��X�@�!����}��7��<��L.���'>��'�D��>�;m�n�hp��7X�I�c�29 �n��|�ɀA���	���9O^�>EZ�L�l�����@X�U@��MK��ʁ5��'���'���ͦ>�,OP����v��s&@Z8��hj��ڦBt�o�L'�����.X�8�m@8j`��#��֘) 9�Ƶi%��'�rDƥg"������Ob�	�9DizE��L5�Rq�H!:��b��b�'�	ß�����%-�{��Y�P�&W� �Lݟ�M��84��T�ܕ'W�^���i�� ��� D���-L�,����>���D�<y���?����?�����66�#+Ԏ9P"��$(�0��s�a}�Y���	[y��'0��'�r%�r��K�DTۑ��F���	�E�y��'+�']R�'��	�vu�%z�O��,�aJ���)�z)XmZ޴���OR��?a���?��OW�<)��_�{�P�D�--4���]�?��f�'��'��W�(�R�=����Ok̄�z��JǬ۸\��л��C�{�F�'����I����cp�ԦOԬ�#A�"g̈�n	�B�)�U�iA��'T��"eT|�H|
���:#ɓ���c��C�=Ӝ(�$�]c��'z��'�E�!�'��'��IJ�!d�y�Ӫ�,���b����&T��X�gV6�MS�Y?����?�x�O���f�)��s��Т� ��i���'�d�Y��'��'/q�HI@C��/.f�h�dXJ�y+t�iUN �%�o�\���O������>aCI�[�T�s���9L@��\�|���?M�|r���O�s�	-Xhh�4�Z�jTaL�}�I˟��I��(l�}B�'��dF"fP�y�E:p�R��"l�.x���|�� �.�����OL��1u^}P` �R,�U�!�"���m�꟠I�����?I�����+�jJ�'1�m��A�)C?����A}bKO�yX�X�I柨�I`y�Ɓ�Պ��ԫA'K_Vpy����a����(��ݟ�$�`��ݟ4pdB|0|8���=8ѳt�ʱnV���	cy�'�b�'��	�����O^:eK�h�^s�51 �54��1��O����O��O����O��x���O��+�fA�u�.jԪ-����=v����?i���?,O^MbT��uⓂ,�$�Ħ�)8R(ak����# y޴�?�M>	��?9F
(�?IN���b��e��тFmT�@<�T)�/s�����O�˓@N�\�e����'��d�\:
�\ihg ��	�����C	Oz���O^ �g�O
�O�S���R�����`I�-��6��<Ag��������O���PD~
� n��QI�~�t����W
@��i2��'� Ii��'�ɧ�Od��(�B�	7G6���S?Fhi�ڴ#�>�׶i���'��O�b��(����h����e�]4L�Q���Ĭ�M3�)ȧ�?YH>��T�'ܢ�+(^Hz�Ĉ>S�
A�Um��E/�&�'N"�'�|Y4�%���O��D���J��J� �2H��7XW�y1#�'�	��@'�8��䟀��?+讴j����NȞ�PP�U�}0�ڴ�?Q�B�e	�'���'�ɧ5��S�`�CR΋.��dⱧ�!�� �e\:�d�<����?1���&\���m�&�ެ�U@ůkH��%�q��˟�IG�˟��<"��ě*��-���J�K�Hc���'f��':�OiN �"|>集�,��1�僉2hu��2��>����?!K>���?	�B�<a�D�L��l��/LElyv�C%K)����\����\�'L��(�iS!)>-�3�$W��(�i��xDn\l�w�'��I쟔�����`6x����PO�$����<rԜ�=9���OjU�D�6�8�(4�D�G!XȈ�"O�1Q�$۸s�(�	�!���q�O��sW�V<iX��Sc�Q�1E�?}��C��-V���g��q�i@�h���(�O$P�e�D ��kE/�j�����$PR`t0oM�\�
��YP��犓)$+T�2OVi����%`��Y�����u%"�jG��L��KD��R7�@�d���?���?��u��ΆD(8��k���@V��"3�AE�CP0ٳ/W�d��,X1�&擝���|ɲx�'�0k��t���$���/Mڸ�E	@�|��q����''�L8gt��a�[��4����]�@ ��\ӟ��'0�@���|Z����y��a��E&'B�H
���y!򄁓�\��"Ɉ�h���QQ�P1	s�I��HO�Sgy�*�2C��H D��[JD�3IT;:�:��d��P�'���'B��]П����|j��NL��9SP��'X�JX���+�a���[(6����'�H��eӫ0���ZCΜ vI�O 5
5�=r@�<���D��G,��ba�C,?tD�� .��:��=P��'��Q�]�$���F�lE(�˕�"Nk�}�ȓ<����"�
�0aя	�<,��<�&P���'<�M� M�>q�^�bъ�9��aŊ�4|H%���?f��?������o3UܝÎ���t�i�.a��a��2`��*5pPI
Ǔ/Kn�!�H�v�:@ɂD6�M��
R����Ao�������Q8����c�Oz��<��b�)vW������
/�FظRD�r̓��=��*c���BSe��fH�(s
�k<y%�i���Oӿsa$��"f[��]ɜ'�ў"~�d)�)�E�1E��i�h����]�<Q���!YG:������xl���GNY�<qd�)K\���Ld��@��~�<�#k�jg4���%=;%���1��y�<�O�\�L�"�H7A�����s�<9�A�2��(a�2 ��Rx�<!V�޼�nl[Q�oő�P�E�!��ܙa��`S��I�k��ٚ_S�!�d&+؆�JT��:��(
��
u�!�DC6$� ��4�-GE��� Ρd�!�DY	m6�+g�%\%�}[��̸w�!��/o�U��[/L����P�r�!�C�t�=��ˊ�[,�
S0O�!�D��`����A�R;P�؄!�q�!��,7�¹��NR5h@nh*��/q!�P�|��$�@����y���2c!�ҧu�>p;w�T�Fy��`��kL!�$��0�A���];c,�%qc-��!�$!"G0���6+�9cU׭]�!�!l+^bD�=�H��dᆸ1�!򄌨q��m@�.��hip��A�!��]��y�ώ�F����e���qH!�dM��X��W	S�P��@�>o>!�$�H,B()C�d8�EH�?i�!�D̻!.� zF�'h��"��;g!��A)n���
[�)t(����5!�$�,Ͼ!��mR�nt��zP��2#!�$J`�j,�Q��:��:�i3!��3aYF���✢%D:��pIݺ!�d��I'��i7j�W�M*�N)]!!�� �iB�8l��6	�0�,��s"OYh�'��2����j��HTٚ�"O<��Bt�����ɒ!P2� ��"Oje��e�*/Q�i�Ɖ@�6�x�"O��iD�LVl�͒c(�R�!�"O��S�B߁.�̨�w@�>:	�d9�"O<,��ǴC�ҁ0f��6|���"O4�����rh�x&%ǫye��1�"O"c�e���	¡�_V|)�'>�AB��!��X0�B>l��x�'GDՃ��W��DA3�J k����' ����fU?4P�+��J�e��Q�'�@Hq��%<�n!3�a�OX����'!hI��!,�Du�d��>��|��'Ĝ]iħաB��@��NǠ-l6A��'�U�`�ڲ8��y�C�����ٱ�'��x��[��F��BeN3uP%z�'�:p �MF�}�8L��f�}�����'� y�veWZ+��8`�,#
�'���ꃦ��e����]�2�'���ƫE9	ݔ�(ԕZ����'�\BզV� Y�qkS�ߣ~�zDZ
�'Id�s4��J&/�#yM�X�'T�Tr�ի"�BőFآz� �R�'���Ӄ��!�4�[v��1y� �'7��
S�K�pI��+��@0y�:�0
�'�d��U	��7��\B���q.Pݐ	�'�d�RF
�_�C�ٻez� ��'6h�hw�F�o�@���
�aG���	�'��]�"aR	5�:�ɴ�K#n-H��	�'P:��i���01K��q�n	�'y�]�%_��8�ۄ�Y T�@���'A�}�N�:	�j�CÊA���
�'~b0�G�7�ޘY��9/6A	�'W�EӵJ�,I8[�+�1��%��'�,�)��/bkxZe�ǥ��P�'�^�B��yZ~Ш�iR{кŪ�'>Iz��KZ�.����v���'�E�V"1�,�3�'|�Fɛ�'mh�h���&�(ab4�_�b����'����R �8�@p+�o�$R�TE��'-N��D>�����4	�'_��a�*Np�P���W�B���'t��
c�W�X��$�6g�1��4��'�B09�/�t��)��Y �R��'"J�K��՜^&[�HZ1#0vŰ�'ޒh�b܂#tx���3 ��P�'ʸ}Q���+N���1��9<���'�pB5퉤����ٝ	꾄��'Ǌ�ybf�^_,m*�F����')BlQ4BE�!�*�@WkΧ�f�[�'�Qk�^9XU���6�ְyR���'��@ZuhY�
"�,�S��$o)�P�'Ru��+��� ��-a���!�'�f�1�nRg�!H6)�
XjH��,-$!b1�V.HK��Ҍi��B�	�A�`YB3�I�I���a\55lB�-}|9�l�+DXE���$Y6C�I�0Aɉ��A�{�4����P��B�I�DL����כ����-��`��d���v	��~����;U i�O��0}8���Bq�<�7 W���A ��F�P(xn�;�p�ũ:��Dѫ0|�?�'8)ٲ�ۛ{^��T�DMS�'�m�4cL�U4��F�*>�� *d#���ƅZA�_a脭�W�9\O� �<y�,@*�M"��{k~t���'�R��$ePU��Y���/Ӟ=h�gՁ$���hG�I�&@!��P�y��?-0�<Ӗ�
�wt��@C��$�5 o�C��~L �����'Z��?5���-KqvX��.QV0�GN;D��[�a�*[<
d���Zo�*a��
�U�f����P�Z��6�@lqP �|
�x��G�6�2�A�E��!.>�p׎4��╢��y��\7
�^�:Q�p.Ϳ? �����0#@<��Ig�����'�J�J�/f����Z�pޑ	ÓXT@y3��H%$U��Y��(2�`$��OU3]g�Ts�@'8�t� M�zTB�07��b�%9).��s
�:e+��
�R]��5JVA⎀=!��t�)�=}�[K�<Xb���O�V'�C�	S��X8T��s�8	U�A0��p2a����
�3��O�B#:�e�kv� !�!!O������y�|���+��!ӓ���F��(�
��$)cw/�!y��9�d
�b,P0�EF�6w�����6j^dлu��a��Ĩ�ax"�΍g��*��U�F��co.�bJW/b�BH�1��!1�!��O(<iS��C�n\Qk
-w� m�'ŁC~�,�4f�`�G�#G�
Y�s�ȭ�?�}B��.A&�t@�Q�d�;�bS[�<Yq/�E{��ɗ�Kjِ��ܱUw�,S�o
|X��/J�I~�P��/B�<ͻo<�֫�/�����j3.�����F�<�g��Np�8G,4�E����9N������3Db�D�N�oX��c��=�hO���B�a����IԊ)s8���'����������/�+&�*�B)�&N���ɗ�D,U^��yb��h���D�8�Hń�I6f��r����i�K�o�c��k�[�/��da�aNH��Q�r�,��`G�?Mq0Kĳ/�2x���]�p*p)Q�/"D�̈�� V���*%��0��@�LѬh(�baaK�B�p��틄�p�.I�]$��pc'�/u�s��@��B�	:A��CƎч����<m�����)D��}���Ly}�K�A�g��&����#h�$2�t�Pq��0,�*���	9
�h��PM�6�Z5��X���
��G�bEx��f����ы���@��D(P��-v�0Jt�hݥ��' ��O�xP��..���� �ۃf�U��k�ႀ��RP=*Dd��h���YH��)�}�(�XT�E�������D�`��� pZU�P)m������$4��h����=j�E��dM�{L�L@�`��a�,9اJkVd����TMfi,O,��ߝ��E���AR���u�����"����j��v�ʄQ�	�u��d���҃j�6�i5�DE���'�:�S8%p|Rs�Y&k,<��a��6S����&S̄4pS�S��6��D�'L0��]�	r���g	a�>E�g�\�nᆸ[W#$���AN ߟ��j��U�RA1F��_d��c�L�!�X��-ǐ]�"	�3n�"j:>P�IY;��Tt}�F��6�����KA��lSBA�7J�(h�'v�Z�MڛJV�2R��9ċ�iG�eZ����i�
c%�{�_������a\:H(�4�T3@ ��ȕGZ�Ƥ���r�F�k(�i>��/�h�qq� 9rԡ� +��y�.C�I���)��Qx5�%
��Э1�p��Dϻby�Op��'���� �7��'�r ��"&�p�Gߖg8�X1
�b��q�O϶'��Y3��@ G[�
sm�=Bn�7�ӷ|7���ck�l�C��{D8|�s+�.6��?6ņ9�l�C$��|����)�s�	�U�����!� �l�q�2^➔�`/^5N�5�aϘ+M�Q�e VOv�T��	p�ʡ��I<C�R�Ћ�5����
A��1 !�A=Q����1uf�杠ti���.X��@ �C�L �B�I:+������'�L��K�#y�mq�B+ߙm�~��Y�E�ؘ��!����<.0�#ף�)�@��R;���W;�4$�2臅p�>�х�iF��Rֆ��s�Rd�Aw]�5�blX%�8�:s!U&��r��-OXT�c�K7+B�Zt�ǤL�pܹ2�x��B�	x�wm�
��p�bM���'Q���po�;/e,Y�$��UZ��kMHX(<�5'��W1f���n�5&�j��f��B)ykF9l�Yaf��j��n���{��H�zN�sqf�3L�v���̎xH<!� ]!An�PQiR�h2�q�	�7V�O2 ���Z��壦 dQdu�4�>�q/[0$@6dYQ��:P  "'QwX�lʶ�Ra��%L^�.��d	rʇaޞ$z���]����C�2!��}��Y�자ر�ߘzd ÓqR��\�r�@��H�C�ƹ&�@���0aR�qQ(^�b�6��W�,��.V@P�P�*NP����I%n4�`�	U��8�!�گ^>��Pl�H�|�%���\���蓪JE6)���Rx���w���B� H@�M2��[B	����'蒄�JͷO���
��� _�ҷ &Y�(�}%��)O>�l)L
&�|�I+O.Y���ȂeT� z$h�*MS��#G�'Բ!x `�
Ӵ�!C�5�� ���C'X59:B����N
8bhY2�i���d�{����a�\���O��㉕-I�R%�V�5(l ��F�u�l!��P?yXؐ�#E2��Y��p��,~`P�@��AHԚu�I*�N ��I#�| v⃑\��H0�@�� �4�$�! �>�g�$c�h������|�'���RE&l�v0�Ńց! �-�"O����bR�m�,ts�H=v~6�+���\�&4؂�R��a�oß�p<!�f�'.Dr��Z�(�4�!�\[؞X�����D�iGn�:\ ��ġ����s�f�'V.��� $�(�Y|����I֡;���q�-D�̠0!��e��r()��Ď��B��'�<�bg�a��H�Q�K<m��C�	����� ҅(�,���
mپC��uY(@BwG\�O�¼2P�X {��C��.L�����N�`���k �7ffB�Iy� ��R�@�/L��iŀ�Ki�C�ɡڮh*w�ּ�r�8�@�F�>C�	�c�|5�5�4�P�����;R_<C䉒�(��V�21xV�i�
_��C�I�UCh�`FL�#[P�1�Ȁ4'�C�ɚ~x!cTCRY��!a�:��C䉓1����I�*u�t̃�I0��C�	�?�T��ɐ0�|�T킁lfC�I�M�l4Y�+��0��'�
�NC��D�@���f&�f��6BC�*�<C䉄Qq�t��D3j�=���"BC�Ɇ|84M�CA��[���N0B䉂Z��Q�#�[�@�nAp�n��|�nC�I�G`�Ͳ�`؞
�������U�6C䉾o��(0�E>����B�k��C䉱;�~Q�J[�}�N1Sbo�q��C���F�ǣM�T�����0HI�C�I�EvTomR2���:$`�(b�C�I!�B�B7I&7��˛�t��C��0��z���'qJ��H �	5��B��pN��	�`�-6�x���Y�S�B�5*�䴠vG��{�XUS��Ӭd�B�	!���B6jL%�-
�,W�f	B�	�R0��{#��;gf�1��԰c�C�0e&�Q��*y$y4�M)�C�Ʉ[L��e��z�<8�V߷��B�ɤY��t`5��,�2�Q�\:،B�ɔ�<"A����bw#ٗ4-B�I�b� Roأc$8,�w�֣)�C�ɾ:f\�cW�ĤyG���'T��C�	�{,�U�T&C�Lٴ%���Me�C�	�.�F�8b�:q�jr!��2lI�B�	a=�ܑcF��	�JM{�EH|TC䉉7��r���M�D��GA�6C�	�]fઔ'�-J<Ĩ�C�\B�Ƀ*P T��5�����EJ1IHB�I9IV��R�F�,MOօ�2�	�3�DB�I�O�4�s#�,/����Ʈ��3�PC��3hi�q�ɗ�\N�}� A��B�	�~�9��.ЃH��4�M� 1�B�I0o�0"EȩB���7o 3vB�ɗ0�d\�T.��f��Д;�B䉑A�h{����8c�-͊;XB�I)6LRn��W����R��g�dB�I6����AC� N���A�oX�`��C�	&Q��q�'�RU�	�CӚEz�C��Ĉy�
�&^�9� �-�B��2h9�<�� @�
Uf��MʞYzB�ɘE�)����!L�p��'hTB�	�)�l��2�QH`�ăÃ	K?"B�)� ���q��:gHUQ��Ǣ��a"O���%�ضY��У�<i�Nq�"O��ї�^ RȰ����M�z�d�*�"ObD�ȊYmn�!��`�p�"O�Eh��E L]2p�<^���Iu"O��R&p����lКg�� ��"O9���h��e��Ƕc���P�"O�U⢩�yb����Ɖ7� "O.��EIa��y���oZ��E"O� B!�A�p���(q�#G����"O�Taˊ��k����0;�"O���S�UB�Jm�FϷ8z�x#"O�x��F�K6^`�P�K�B�P 0"O�<��n��a iF�_�k��}�"O���2B�Y�8$�t��!V�4��"O� ` G�B��Q��"�p%�"O����M˔y��E#��O;�V=JC"O�dH�a�!��I�w+C�Fv����"OL�P�U1}m2��kQ�q�1�"O�m%
\�,&m2e��0m;�"O5[&X�rg�}3鐶o\P���"OX9S�� >�8�&� �%FF��"O>����:$�l���׆R���E"OjC�EېLS��Z�F�`��i�&"O1 �7P�5�޷'�m81"O�A{�+42��T �����`"O���GM� g�h"eG�B��,Ib"Oj5ug�:�Šw$��d�\%1�"ODI��耲-�i�!c ??�tx�c"O|y��F�%XNyJ��� ��"Oj�ᔃV{2N�kE�"�<��"O�`k��
��E�B�<{�F�c�"OL9p7�?H�,���I�[�.)	�"OP�H���ltY"�Ő![�,1""O�(�7K� �����'��{�"O`�4�܉M���¢LIU4uR"O��+fm�V���A�K�o&��"O݉��X�6�sb$C�L��`��"O�����݈k
 �B7�ڎI�x�t"O�t��K�o�;�ț0��Q"O�u�/��T X���#��A�"OFh� ^�[�2-�S�{��`��"O�I�d͙������&�"Oz`:v�U!1�px��c��İ�"O� k��v,i3SE��3�浣�"Ozc��@l��K�d�/z����"Oԝ1��6��Ms5�V�{r�cD"O��BA%Lp�.��"��Y 3"O��R��V)<M����S�	,�"O�I�TiK b� �p
P��s"O\A8E%@; �H�)���!r�$k"O E�rDŻw
1��!W��t"O~]�Ql�"�����L�l����"O&��p�_=T.��@+�,l��9�3"O*¡eE�eudD�0�h�2"O�!����4�ʭ��pV���"OV��tE.��S7[	+H��""OxA�²<��1jQ
�-	(a�Q"O ���햗r�j�)��P�*��"O~x�r�-O.��F�H�Z�~��"O�A�S��
Jzfy�a-;_�lHr"O��j�:+Ya��W/ ci��"O$�ГF��:Z�k���O\�Dx�"Ova@c�'Y��ah��PFU��"O� �U��S?P#`h#qҠL*�"O������i�v	�$.-L���"O|�` ��Vy:� G5&�RD�'Q�صM��/���1M 9��J�*(D� SD�B�F�*w�\'d�$��g%D�ĳ&��o (5�B'=R �-�f8D�,
�I�!!h-���<С��3D�����O�v|>�K$��Jvtu�R�+D�$H���d�d�SÅї$�j���<i���ӆ:3��i��5����K߅kt�B�	����	�
���{���BfB�/A��`y�Ȕ<#��8��S�i*B�	9O���g^�g�,�e��0QB��pK�)��N$��`�Ϙ*f��C�I
J�H���l��!�X�����e��C䉙�N|�QK,��aT�8FtC�I�* �	E�Ɓ�A�c/RG�B�	�_�vM��n�:�A�ʽF,�B�I�;A1A`�>w7���"L�:��C�I1@������:D^��J$@��h�B�	.?�zY
Wd�r��L�� �,��C䉱|���p�S�z\!��.-�C�Iq�&�8�d˘_fhp²��4��B�I������,r8r%"��}�B�4I���C��`D�t�3ԑP�C�Ɏ%�|��"K�?..lLR�k����B�i!b�Ӣ�M�L�\(�Rˈ2U"�B��`a\Yj�钂&��$��fJ��B�	� sf�ɤj�&��H��I7��B�ɋ(_���O�0�-�CF�hn�B�	�*	J�Z��D佀�#�vB�3UR���دf�h+"�Q�hB䉋Y����b]�9�hx��͉{�TB�Ik��) �A}^D�p�ϝ1�B�	o@�D%)��#��K���C�	&�.%��*��Rc'5|�C䉬2�l�iB��
b��MS� �H.�C�I�Z�#B#�r�J�9��C䉆�d���\�!g�Ѝ�C�I
��x��'Ȯ�h��M�opDC�	�X�ɀ�}T�If��B�hC�*���0�c�	U�*�*V�L�
C��"`�Y�Q��>ʼ`b�!��._�B�	*;�}�Qj��F���Y�DH ^ɚC䉺b�H��uM'~ɐ�i�)F8�DC�.]���)�#ڥv-:Y���7??C�	7` b��!@���`u� �+��C�I6k��<��.׆F�&<���{�C� y>
���Ar�JE�̞98��=q�'c$8��FꞲ*���qW'
�o%@%�ȓ;b��pM�%��#�բa��@��PpR���!��M`1,F��!��UHv`��I�2\��+Tb��0#�E��P�)��F�2x�>E��b�:Ї���!��4`�$��+?x�I��
��tXtǒ,7R��1�n��8�ȓ
�:ݘ�)��Dk�͑�9T����ȓ#Ϧ��EL��";(�q �V+�����Gul�3� 'I����(<���ȓ;'���Ӏ��<�$�Q�W<`O�	�ȓsZ��1��y�,� ̑H�V̅ȓ(�*uXT��2��U�!���6��Ԅȓ_3�	!+�c��A��AH��X1��eU$��� �'����	X1C�T���S�? �-9ԅ�*|�*<A�ӛ&�ȕp"On��F�ۧG$�{#g@�)�F�)�"O��Q�G���l]�x� t�V"OD`��JK���B��	�N��f"O��y����?�H1�%ȇ4?4��v"O�����
@��d"��Y<�5q"O`�P$	%i7XP�[��2�"O�;[r�9�o�%Q�d�i�D�?�y�F�}���"	�FӞq�l��y��M�N\�rIS��Fk� ��'���-ȓi��-����;?-��'i���da�(~پ���E�
B�u�<!��N`Dܺt"��e��0��[�<�Ř�Mj�]+6�<��%v�W�<ф�8�NQ��V����T�<aQB���c���]��j�Qh�<��:���oY$oL�AB��\�<6�	�~S"eY��Fb׬MQ���~�<٣�]�cQ�!�q��{Bi� f]x�<�p�@�U�Y�!؇+���`���o�<y��\�3#���C�8�v�2��V�<�e �&O�511�le#VaO�<�5.MY�R홲��2`t�@M\K�<�&m���`�� 0q+�QL `�<!uDM�5.���� m��*�.�X�<y�d�wS4��0�ƒ8܄H�!C�X�<	T��Ymh�8�A\�d���ԏ_�<a�J���,8�EJ�	�́u�t�<	%`4")��괯��H�yejn�<9eA iؼk�`B�3�:�ˌh�<�Qg@�Y���	�~�� ��dHh�<q�AP�X`���(�mA���l�_�<�2�A	>ۚ���	ه*\Qa�"�X�<ACO\�6�����ʅ �ؼ�Q��R�<IT�ݨr=8��%�_�ɘ%i�
KM�<#��� ��:�%��*6��F�<Q�U^kj087��g�F�I'�>D���8�Z�kV�� ���l(D�({�
R�¹RA��? t�*D�(:�GE�{a��EC�g��D*D�I��7g�j��^,z>����)D����.ܘ� q��$:>T����)D�t�g�L,~.���O[�Y�*� �d,D�<3!VZD?v0AQ�<D���c�w�0ك �>T�`B%0D���p��5g��"��4"І"D���Uo�Eh4K�,[�Ҙ�!h"D�dP�L�4r:��IUFʷ=��hs�c;D����MD�?1�y����%�p��%),D�4*T��<' ��FCZD��u�&D��g'�Ui@ܸl��-�<�hR�&D�(X�B4{��` b@h��*W�%D��GI��w�А�RD�a:c?T��/�������sr�"O.	����"�@���'!2a`"O"@�����Is��&��e"O
����*pZ��͓�e��(F"O�d�`��Q�d����DȆ��4"O�$8c,�2k�je���&k�`�A"O��vl�0+ݢ-�Ś�ʼ�W"Ob�p-��v�:$���ה{��Q'"O�au�G#N3p�U���7�|dK"O�(2��]; b�䳐��	j��6"O�q���90z��(ƍɺm�F��"O� P���d�!�n�!J��9� "ODb���ݳG獲ak̜{�"O6���f;(*(��ǉ1�1Xf"O�I��W*H��Ȁ3Y��1�"O؉�G�ȧ0*4@$L4yW���3"OD�صdF$�L�3󃃙?��"O�cU�_/P:\[���E4�89�"Ox�����p�D(�w���YL�
�"O�t�S�0�h=� '[��F"O��hn&=Xd !��IK��;�"O�D�B=]��$Ic��Gv!�"O�͛f�S�K�r%����N���"O��O"�A��Բ5��]��"O�D{7Ɖ���)91�ҳh0�0�"Op��G�m��l�H�(�����"O�ъ��ԙY����pgB�s���)�"Oh,˃�� �Q�����܆Lc"O�$S�ꃬ*Ʊ�į��(6�q��"OVb����;�̛Ԏ�>a+��f"O�P�L�"
��y�k>+x���"O�J�fV�)� @s���7%}�#�"Ol +�8��@�wȋ ����"O>�p ���2D<`�c��8�:�"O�0 ��í'e�e�Ɯ���a"O�������,�,�f�\�N�R%��*O:��H�$("\��bL RL�!j�'44P��#U�q����璻EQd��'����3�X)=D�"���<��
�'�n�A�Xm줘���%���	�'��Q�
�f�lI��� ��-r	�'7%9�G�*w�$�˱#�1j��] 	�'�4d��̗-�L����L`E���'+���`��51�����ZbLH	�'�F���$܂<���@��!R���'��]�JW�H[�\Jf�ޡҌ���'�z���/��3�	�ϗ�<L��'i�-)�Ϭ"�����]���)	
�'���S���_h�7g�?�����'��miC,�RB�	KKujR���'vP:�!O��E��N��g�I��'ZF���
V��"P'@Y�x�Ҙ��'����0��<��p�Ct��Ը�'�,��FjZ�g�zp�Q	v�����'w�m! e�=;b�@2Dq��MR�'�	��$ap��O�
W|ވ�
�'���($kO<�Ĺ�p��#S�.��
�'2D[4Ɲ�*�i��	�w�X���'b:t�Qo�q���Ǥ?n�BP)�'Wz(�RI�o��=ۧ�B�s` �'���"4 �(�*U��	F�d;�r�'�ڰ��L��PE�1c�z���'L�� ׃.)Q(�`��Q��(j�'��,(Ԧ�aG����E���C�'r�X�&�;l%WK[�r*����'\<`a��0���`�iE54�*�C�'�PY	���Ea0L�C�0[��i��'E���aDź43��� ��c�Ly�'�A�@�P�]TZ��'n[�i��Ui�'+�uI!�B�@�y�.į_#Z�C�'��q�m$��7N&(�
�'tt@��iɺ�^'x����'�H�O�0b�&���� vG�Yc�'�V�[jҝ/{.4�f�gc2��'�ق'��-[�n�k脘n�*���� r���
cnR�@��^�&�<JG"O����X9����Oqܩ�""O \:B��1!��*7�+��us"O�+*W&8���S7�O�J�H]Ӆ"O�A MJ$��p�e'�R��"O ��r�X�}���+:LHi�"On���-Y�"�y���â�bb"O6,��
&4��`�ЬL�<�r�"O�@��*+,��J�
�6��"Ox�s%]�ڈ2�%� �"��q"O�L�����*�H�(0�X�/�B���"O����f̔n�>�(�Q�<�|�["O��cgnYQ� ���+E��HX�"O�D+PnËy&\m��mO
�&�JF"O*p�ԣ��jk�,DV�ԓe"O� `GЩ����pM�6o����"OF���*Z�p8�(RBք��y��"O�H�0�74���ʟ!�� E"O�4��f �x!�,�3��$�"O@(���1@x�P�b��v�	�"O��;W�˺j�A���x����"O���rث��D�ъU���"O���5��_M���KU�uۮeY�"O.�8t@��=��@�\ժ�"O���"@
;o^|1Vɜ�J]����"O��� K�3�xPK��_<��U�T"O�y`��Lt�E��T�Ѷ��"O�DYg�C�m[��c5��\��%"O؍� BP5����K���YkP"O��ѢCo��q� �$�Z���"O�D0P!_�l*ZY٢�վl�y��"OJ�S�f˨;�D3d�,�.��g"O>�A��l
��5�(J�T,ã"O��p���a| �GB�����"OZ����,�LU��jֿi�2�;�"O���fP�[�TwK�v?20{�"O؄�6�2<o���oU5(��a"O�,�F�3.8Š%O
w@�!��"OX�8u�&&�
�Y�.O�.0�:�"O��r1ކf1������u���X�"O��[���F(�h��Ŗ`�t��7"O��5m�-C]H��� L}��!b"O��֤-Ql@���Ln�uw"O��������Y0�EܖNj��&�|�)�ӯ:5��ōB�k��D�d�̭I�BB�	�~v�5��H�3$�v�%L�jI6B�I��Hh3��ӏl�z�2 ����C�-RZ�c�@�n|��J���C�I;W�P1�E�ϥW�b�[KԤNƨC�	'V��pA%��>j�P���b�l�Or�=�}Jf��?Fp�� L�����KDA�<qa� �(�_�!h�]ZC�DX�<yq攋}BS��٪ir�{��	@�<�u/Z�b̹0��g	b$�P�T�<��սD�E�&�&u����`8T���g{y�I*D��>G8�"�,D���1�ֿ�,a�E]�`-0A��5D��qaNW�7�.P�BbF2m��(S�4D��+�*[&iDV���+��� �.D�$c�M�5��%��"�8�¸�tF.D�dS��� x0)&��e֜p�h*D��V+�=$ ���_�^��c��'D���'��0�<qA���:B깲`�%D�\Y���C��-x��#aXq�	}���O� ��a޶	�0J=H8�Q"O���Ti��B�4�f) �0��I�A"ONA�e�-y�Y��ӞG�f���"O~�悒2.�]�f+]!��Ev�<�0k�Q�h�+s�z	K�m�<񧀆,2/�Q��mM�]Ul�Z�c�R�<�G"^J|�F&N�2=��ǒRx��'fTq�I*S̬�;���*s�x�,O�=E�D�ެ���`)
9;���F*��y���$	 ���KV|�E�	)�yroT J�D���^�I�)c�H���y`H�fs�(�ET�GXvmBd�B��y2�G��x@��(G��t���yB�<Ҏ	A僒>US��:���=�yb�˛n��y��Dw �I1��I�hO����оL-�Iز�U	5�9�o��q!��К0�x��A7�&q�7�B6>i!�dA7z�|�笖$��1��O�	�!�R3EL�8gצLaĈ��H� Q�!���+$K����!LY��ْ4E�4�!�d�&X ��5��>�ʽ��� ����A�'��R�N��xx(�0��)z.P8b`"Obؒ�_�E����	�B��z�"O�Y̊�#u��)Ԉ4r�M�6"O����D1c˖mTBJ�i�4�"Ol�)�	.H*�qG��xN4�1#"O@�psd��4���ꀏ?�Ʃ�"O%�@��-3��8jS�E:$�&����2�S���B�L�)���}�>�J#���=!�d�����+�dW'pvN�Sa^w!�DP B8��Q���Z,i���=I!�d@�h��Ip$�KOzR�+~ !�$Z�e.\�0�PZY�Q�7*!�DH�{���G�x \��X�'!�A&����#v^ଐq�� !���_����Q5mtD����	=�'Ua|�b�?e�@�WI���\�2��-�y�j	�)�nl��'�H�jf�گ�y���~ ����b6ų  X�y�hܵ �0KB����ۇ��y��L��R�Z�.�I^^�9'͛��yҥ<E�Ȉ�ĉ<Vvd����<��'�ў�O��̺p��[����D�׫Z�dU��'D��炄�[�� ̶Y��S�'�T���B�{�<��Q�۬W1`���'ĸ�1��A>}��i�	�
=�Vx��'�|}{����@)����-JT�x�'��E"�0�& ��/�-D�H�'�"d���TQ<�����-���0�'p�RI_<f+��6ʼ��ay�'B(�٠$	)Y���Y�Ǖ)Kh�y2�W�gE��ђ�IQ��+��y�%�j4B�j��]�SrP+�+��y�%�\��X���TQ~Z8�v�%�y�lS@����d��s�ҡ�����y�[�%qޱÕ�Ԑ5�`"f��y��U��2	��{zla�r◻��=�$3�S��݇0����Y#Y���WC�o�<Y�2z�,����
�< �u�<��υ
����T���a�'��t�<�6k���|j�'��Q��5�ƏPl�<)��p���OP6٢%� i�@�<y��
.�H�ǁ�9h���Λ��8D{��	�x�ҝA%kP�`/Z���Ɇ�V��C�)� ��񤫖�+M����F�A� ��"Otu���Y�&�48��)��b"O`L���і%�����"�!as"O ��7#ܩc�lĺ�C[�i2���"O~Q��
���f�6��i��=	a"Odx(7o"CH�����e��ѣ�"O�����2
����7��:��Q)�"O2� ���$���9�#��C_�#F"OȤ�t���Z>,U�h�R���#�"O���Qㆠ3:��G�)	n�4"O��a�ܕU��-Iq �!/ ����"O�����h=�� �8� �T"O`�� ��:n�p�f�[�#T��*q"O������9��|�c�H3Q�u��"O8�pV�H��|f�C;�E�"Of칑�ٚ��)���r.p�Z4"Oв��T����͈-4M�*�"O\��2:2�^�[6�*#Zi;W"Op��@R5Ȕ#����:�x�"O�i����m�x}u��i	���T��G{��	�J ��QH��N ���2!��#^��ۥ�פ4����S-B�">!��U=ˮ\�"oHyͺ��ҭ¸p+!���8�~9yd�_�M��Ku�M!�D���R���ְW2pSg��!�L;
�֔p��B���<I!�dʃ.���I�%�
d	�o̽xGў���ӷu�0�0���RFy
�ɞ#{�DC䉥v���I�i�j�2��%eX��&C��H��m���Fb��s�*�M��C�	,G�r� ⪜�}���qlU�>U�C䉊DRpT2��X Lt��Q�V�MkNC�	&z���7M�Qt�dP' �
WlC�I�!���6,Q�>j�@8b� 8$B�ɷ�.����ð�*���O6�6�OT���] H�AĨ��4��< c�*j!�DVqq��I�XW�rT#��{!�dƌt���@�B; �q'�4B!�dH�D>����	Z5�)3�B�(p�!�DUJ���bvJ2x���]�n}!��F%�iXs�m�Xh��(�"Zu!�D�lij�q$�g���{����*�!�_��v�#�r�+"@�!�$�14���Z7�[=(���*��lj!򄃌=(L=T���B��A./]Z!��	1�I�ЪXo�����&R!�D�Z�	����W�"3!�M� E�Æ�:$������c�!�D�j��J�46|�̗�$q�O���$3B���%&C#%�`z�-�<0c!�d����	W��E��^�P<��@�8��h�����z�$�X��фȓo�0	Z�ʇ�7%�  �j��:Y���MZ��$��޹Ӂ�͐I�^���<�����N
�$��6(Y�rH���O��2F(Z:�N8��U�v�j8 �'����_<4)�H+8e(�'qLP�%��$�5�n�%@Ȟ�
�'� "��pTî�$2��z�'ܚ;ɕ�2w������-��P�'���	 ���y� ˛)�H��'��M�W��PCp�2MB�7ʤ4��'P����NK��l�Հ�+{gDQb�'�K�\$��a�(��#�(	�E �{�<� X�[TB=8�`9��ހg�&��"OZ��ƣ��y9AR�\�F40�"O�����)V��-�4�ݨZ��M��"O.��I4Cpݙcd�P�� ��"O�����^�&��rt��4V�T� q"O�M�$j�_u�=H�RD�����'�!���K�\Q�#B�=
�y��(�F�!��^���FP3~�t��1G[�x!�[�4M�� �Q5p�*��LV+�!�(Mr�,s��H�(d�b�
�J�!�]2]����#@S3� ܐ�h��6!��5Y3�@�eA��"rFLI��_�a!��6%��x e�K�pa&�k���i&!���A�����,5�T)ɲ)͓�!��k�D:p�I� �$L�gi�v�!�C�I.��r[u�t)�@��u&!�d��q$�j�j�R��@%�ʟi!�Q'���Ĩ 	$�ز'*��d!�dȮ�a;�E&��<3��X�E�!�9L���3!��T�Z�
��E!�$_+��U���J<��A�V�A	n�!�30�a�	�L�:��v�
On!�J�^�􄠥`S,�Ճ��ւ�!��;I~)(���%uh��wgN>�!򤕫^�0Es���L9.���E�:�ў��I�)pF ���%m�Px���!^��C�������	"�>���%C���O���
T#l�P0��8l,��F�ad!��(3e+���Zn䱅�Q�TN!��V9�(x�5�Ї?�M�CWD!�d�)Sn���Âr�遐M�,4!��/���'h� �܈6k=A�s�	N>ł�hG�O�A��U S ��3D��ӇJ��@�=�Ǚ`� *�"�O
�=E�$�Q|��j7� R��Ã)͸e�!��D�@3�-ÀFKxdʆK��!�ߕg���g��)O$#ꀚ-�!�d�'S\�!R��5v6�4(�1?r!��èRV���F #��wHĊWD��F��|ztÝ
d]*�jSAC:M�!0�+D��q`�J��D=tH_�g4n��3�%D�|�I��KJ��������S�9D���#�]���AaG�,��� �8D�L+ E  "�y@7B] c�ظ#� D�<��Ô
a���	C�����>D�P0��êo��l2U�V��8KC;<O*"<�V���?��5�# .4fT(�Vu�<9��>Hk"����ϩN\$P�c�o�<�FB�xy�*�#[��4��Vi�<��R	DA��!4/)O���Kej�^�<�D��B4HD�
D���$�Tp�<I�`U�d}t��m� ��1��Mh�<і�K�k�,u�£��^�u�' �f�<���-Ks�	�^$[J]څ*�d�<�r�1�t#��W�@I2���^�<�`b9}�`C.L]&<�H$`P[�<�`3Ӑ�Q��T�M{*�	҅�^�<���ÓE����	$��1
X�<���/7��	ad�mE�<q��Y�<9�m![\��b��(��)��@�<#M�M�x��D/�/5�@�H�{�<��۠a��[d��<U�e��R�<9rl�m�ε�!Ѕ�x���K�<�b��P{<�E�B��P�&�r�<� �L�틶}H�"����:l�#"O�]�+�&ݫ�EG�׎��"OFhs-4������R�P��R�"O�@�ÀA�xޙ�S���d����4"O шT&־�:`xr��~lv�(�"OL1
�cG?c`5ia��":�R���"OH�ׯJ&6�\|�T�L�@�0�W"O�����f�@�
3jؔ~����"O.U�`%��z���#*G�/�؍�&"O����Xa�J�Ǝ�E蹢TV��D{�ɔQ��$���L�3�HB�=�B䉥yd5+B�J4c}��d��:�<B�	7��zB��Ij��yDi��XK
B�Tm��а!E�P��S��:sC�ɞf;�
�T�k$� ���~�B�IW&p���60c>x(�C�&�B��:�v���X�z:d��-��84��D-�9�`!�>Պ0��;��U���;D�`��F�Y�0����5:V ���8D�4J%"����]��JR8!"�ba6D�L���y����3Fb��c5D�,��(�	~�.��C(�8��q�=D�af]*S� �s�E]Iw��;D�PH��z�������$������O�=E�D��e�8� �n�/(��]˃m��~!��Q�myd�&��%l�X�ӫ!+�!�DLgIt���KXXj�h�D�D>!�"Z�8`d�!s`"�H���'�!򤃭 ��q����G�L۔�Y�O�!�d�5M���� 2�86���N8�B�	�y���Yq˗Y�8-�sk�"^ƒO��=�}FI$w&��򦀠e[��(��U�<A Ό�!<�pw�M"^"��ReR�<��%�[Y�Ts@��($��u�K�<A��&L`9
"M�����ME�<QsZ!M0�耏�)�2�)��y�<i�(]�x�A���'�h!$�y�<�C)ҀAh2%:Ҥ��Mh��u�<�Ye����'_�\�J�E��)@�!�Ă��A�!NG�1����Oߠ p!�	�`��Gը:�P�yaB8Hx!��T ���`e��3�x��B]q!�DZ@�fDᄠ�1�`b�bh!�$Y�s6�T+ƀR�C��YuYGP!���?�ЈR�Q,^]��*3`!��T$��рK"k��}��Ǖ�eK!�Ę��@�sM�.��"%�4�!���/'D@�k�D)B���Q�}3!�-���Ps�Whp`��[!��-'�8=p���=z�hP&$1!�E�M��T�Ɵ�F0���"��6	�!�d�=Ů}�%g� .Z�5Aٔut�	N���B!��:�̐�V;D�H��
!D��ȱ�?X�D�U���s�tKB&3D��z����}q�ɪTe�+\'`��L/D�,�0 �&j��`S�A�rGnt�� 2D�� H�B�ęq l�NP!��<D�X�ӊWw�����
9o�v��%+-D�@��o�[Ԣ��w��L:���'D��!6�8�� �a��ޅX�@B��k�ޠxf��<7�zqk@���PMdB��?���e��(~)Q��M&��B�	�p/X�� 7�NspeI?C�	�fn��4���]o 9�1��U3�B�)� ��X�ʚ�@$���(��ި�B"O(E�dc���:-��{8�u��|��'�p\�v��B��"7��i	�'\�0�L�\�@L�%�"Q�����'G^�:1��DM(Q{���FnΥ;�'B�[���o$YҶ�=�x��'�
���:��%;�#�0d޾!k�'٢�xCɕS�"��v��9`.���	�'�����Nc����v��;.���x�'|��+g��yg��A\@a��'�)�AO9z�
�:���J}x��
�'dم`��jY)�J�E�L�s
�'�R`�c�B�(&�]��&q�	�'� Y��T�.ܹ������'=z� �-:BHi9F�ݧL��]��'����/��F�BE�B.K:�l��'nx��$��x��$Z�	�(I�J���'�@ه��<"����0nV�n^4���'
f	�5�R?=Q� AE�Q2�'6�i��o!}�|*����+
�'��� aL8/�vL�n|�6��
�'۶(�#��u���g�'���'��{�M	�}�n��K(:x���'�`�bዉo�̌�&	��i�.���'�|��( ���Z��{�D���"O�(�_(xfO:	�T��K�0[}!��<�"th#����i�4��!�$�'���劄6�����/DGH!�D͋l)�Z�K�3CΉ0e>!�ĝ;0�2 �q�k(,�I�-�,lU!�D|$����CZ�P��a-D�E!�$	�\ �Aa���Ѓǎ4&A!��>[��l�1��%�&��p�.0=!�+d?L4	�/��z���?~E!����bt�UlV�.��q�Ƃ���Pyr�3L6���7���Ls��pm@5�yBK��*n68r��:H�`��tnP���O�"~��T�x�Դ����O�x�!FW�<I���4|�|@3N@4��T���k�<��C�w�uZR�H L�Rt�s`o�<��n�_���� "Z�Ȱ��k�<��I@7'�
	*���WT`pS.Ne�<��eޓa�����>Xi��[d�K�<�&��+�{�)�0�R,9�ƂH��0=р"�-w���kĠ8����J�<��e]�`'xI�����Z�C�B]�<�BC Z�Dp����c�� �`��W�<it셷o_(<['I��&(�x�I�P�<C"��Y�����I=3���J�P�<ye���cR2�)r�f��	Tc�Z!�ď�,jh���B �L���"��rW��DƔ?�Ra�A�"y0-��G�_#|B�I/c6�0�oW:	��Z�"؆XvHB�ɬ9}�P)f�� ��8�E��i�TB�1O���.	��P��jE.Ecw"O��:��J<�Q$�3�6� �"OI�Ǉ�@5�1���O8`Y0qZT"O��q��1
��ț�j.	�L���*LO�i�SK�`�%JԼ(�>��7"O
��FCҐBT$`�����)!3"O�}�MI( �����g����"O�8#���T"��@��zk�"O��w�
*BL	"פp�t$�a"ORTj2"7��:���)���p�"O� �U���CD��#��d��9c�'w���V6vpI�ӣVy�T35D��!��0Kzu1"n�4a&�d)7�1D��f	(>��L���m�A�R���y��Êj��[5��X6�25��y�
�Evc���*Wd�q�.� �y�ɑ� ƙ�����  ��'��>�y�i�S$7˒"J,"�Ss`@�!�Ă.#���f璥Y�z �@�K�Y�!��4j���c ���|`����$��!�F�pE�AxQh����b%*G!�0.�!��*1챀"!�!�!�d�+n�T�W.Q8Zc��CC*�!��D�^l��G<1��EF�0]�!��H��ҥ�)bJ(t9��H�!�=+_�IHE���$�0r�m��!򄟸6֜so��Wk�})��-(!�DK�:L� ֫�#
�I1�K!"!�$?h2�: I�`�s�蘼�!�_�c�aaD`�'\~�2'@�*�!�%!�ִ�7���u���S(.!�$�#HΦ�1rK<�n-�@HO)!�$�;IX��`f�����qU��Lm!�¥	��u"����-�� �V�vS!��O0\�.�a`�:gs(i�#
ʟT]!��'LT��%�B�CT��ZpJV�{!򤗲^ ���t)�l;|�H5/�m�!��O�C�v8(4��f���9cJ9H�!�$��2����&ߵ*�f�i�LT�
�!�/Y>tG�+��!��.;�!��\061j$�ҔV�$\YG�Y�}�!���w�,�K �Q
i�P�3t�� t{!���&��Q���@�	~t�¡�)r!�їB]n�!B�;m�(���LLC!�D��n��Qr#��H�b�a̮�!�䟽T!z�s��9����!��N���$�:]�P��EC�Fzơy�G��y2"�4 ��x:bD�>ꀡДƓ��y��y<ȕ� � ܺ�h�7�y���J�س����3�^��yb��vu���tCR��`c���yBF�9k�} �kL�	Q��y��_�c��7Ɠ�gx�E�gIޅ�y�BU<uH�R��A!w�8�xoO��y�/��F�.��eɆs�E�Z��y�M�%8��+��� q��t#�)���y"�C.[2`<`0�DiƖ-RT��y�� H�8�P!�Iw��,h���y�N�Μ��$KѲp��&�y��0Y�d���,)����ޜ�yRe΄t"��f-���4R�y� a��9��҆�����yb�ݶ0��%C��÷9���k��ݩ�y"aL�X���D��0)L,#ֈՌ�yR����9�U(ۓ&�z �_��y��1L &���f��2L)�l���yRȂ
pd�����J-���K����O`#~�`�D(��\�-�VA�q*����0���t��:kD��V�B� 4�ȓ
 �ԋĆ�:Y�XԯC0m���C���i0���0\���B�"n8�I���
�p�FL�a+�ܫwO܈3���ȓ��Uy$�*GE�Pʢ� <$ �ȓR��$J��aN�@ڴ�4$$��S�? ��Yg�ғK�U��j+.��y�"Obb���* �ݫ��&|��"O����g���ȹs�E�����"OdQg�ԷY9�S1��k�����"ON3D��h^Q8��XѲ�"OƤ��b^vu���Ԩ�?>(��q4"O�Yv�֙��1�^�R<�hR"O~�S�O>G���Ғ�]9Ү��"O$��I �.�W��`�&��F"O�a0���YoA��C"��"O�8H�3%��A�-� +ti{�"O� uI�6/ �	���>-	�L B"Ob�ȧ�]xZB��U�.�S�"O���B���~�ƪ�+NF�{�"OL�d�0l"�D� ��5q���["O���	�Zu��!��8��b"O,Q�H!U�:əQ%��9�tt�"OHH�y���g�\~*��g"O�E)�-�� ǂۂ`_�7xp5`�"O�р*ֹA�.�xdO�=� ��d"O|$�se���%s��#K����4"O�t�PBA�t��rge$w� %G�Io���&JPK��I톛0Z��j��6D���S����0l"�,��l3D���d��rȬTs�&p�ȹ�'�1D��W��O���ϙ6��K��-D��%�N�sp�&�/
x�T�/D��ٲ��]$�-�F睞Lv�C��'��O��S�]vb`�Ɉ�s���X�D�^6���0?�!+7�. �*�@m���$�l�<��ʉ�9?�9�D�!-�\�C�E[R�<)%n�i9����)Ƞz;�D��O�<�b���� D�&+���IlMJ�<�* 	~~�@�Kؔ$�n����D�<�S��L�JI:�O	5�����C�<	rɝ�'j^(�0�����V,�T�<����#Ҹ�ҁ▰ Ű�£��i�<���;b�ň�� �5`�Am�<	��ֶ5�bl1���>RDڥ���S_�<�7�4<,L�:O�j��A�<��e޲t�0��g�՟lQ�(B�Q�<�Gn�-�*��K�U�Ft(���K�<Y��'~��}SQ-Y	I��@���l�<� �<���� M|��X�
d�<YE��L��c��Z֍�#�c�<�d,����&#Q�?�`�A��H�<��ɇ�,���N��.��`A� B�<��g�L��ك��/{tZ1�b�Xg�<�r�X�LO����`�)I�~�B`�<)3o��0S&'R�h���4FM֟<F{��	��M�>]��儚+�`�k�⁻lnB�	29o�)�f�
/��X�e^�f�B�ɘd��P`"��$�n��(�ec�C��R��p�Y�3"0t�"P:��C�	�0���#G��6A�Y��IκB�hC��/��y'jJ�P/8�(̸C�TC�I0r�����fܗ@� 9���S�l�$:��jc�
/|Z�ۇ��ظë!D�tR`�ۤy�Y��͑)E� �T�?D�9�e��'4�TS�0v;v����:D��
R'��H4r�
0�h�zs"8D��Fx04�t����.�`C�	Ihu��nǚu-�MBr�םb��C�ɄQ���`��8��\��(ʢkZ�C�)� ��q'*K������df�v���"O�]���{.�����)l��|p	�'b�e�����P"j�3����MZ���'�	#u/�yezD�B�<���'�j��N=|Luk��	� ���'�R!�ěBbdxCƍ"��!�'�hC0oJ,NXv���.#9P �
�'�ލ0�*D`xNh�b@A8�`�'��ڱ/�;=� ;�)�d���'h���oLC�쀐)%6���'<1灼;vfp��b�� �����'U�Q���8�9�@�$>���'uҭAЭH�F���2ä��?�rp��R�'�B����4IL�4�3���(���-O�q3F�R+�xe�_n9`�"O���h]6*���Z&&�BI��"O2 ��GǙL�����*�x6"O�4y5EB\0lk�`0c���"O0ScgP�H�%A�^
)U"O���f�^�����9"d"��"Oh����ԓB�� �Њ{�v���"O�0����v�^r�� �*(!���7v�$	3)f8|!81��5-	!򤃿'8�d�ΐP0�ɖ�R�i�!�11���8d�ޭv0f@�Ō���!��Eg�R���f��c?���qe�R_!��A�-�*�+��T�!�E�S@;!�ϵ����)Y����QbD��I1!��sņ�(P(+,
%��#T;B!�5}�F�q(�w��(�PV�!��I�:�;S�[�~al��b5b�!�$��<X���D�k`z=�w@�'t!��D;N3��y0i@fV�rE�R�t�!�d�G9z��@`^���Wǟ(�!��\8��)���\�ЕŚv�!�\#g���R6�
l�d����:�!�	��(�ʂ/4PȤe�PǀBw!�D���^�	o������!򄜍M�2]�#����L�0�%_�!�^�0
�m�Ã��q��a�U��6p!��b����0(@�M�>�{7��}���9OZ�9��o��Ԣ���4L���"O�1�|�xf�e9j�@"O�\*�i���xp��cū$�xS�"O�� F�>7b��CǸS����"O\�xv-�fi,H�ȇ�,��qؔ"O�@#���:�L;A������"O:Ԁr�B�6�@@'��0B��t�"O*IYvf	�`��)FA�jP
 "O�h ���\���с��6 ���0�"O� x� l8UA���c��-j�"O4XDl�A{�Q`&Ke�:�"Od�L� Z���#��s�ۦ"O (c��	[ۢ5`�M�LF��b�"OTuSpo��h��E;dK[�<��"OԨj'g�*
qN����6�$\[a"O~x؇�	�R��y�@�v"O�!6&ܥ���u�\3����"O���T�I��M9����"O��C�6/n�ģ�,�#t��ae"OvP��? ��h(���>!+6���"O�kr�+���(�B�'@G ��"Or�[�a$�tcT���>��3�"O�@T'�FcRMr��ד[�: �"O� �4�!���eK���!�*��8�"O$LYqk+7T�w+Y�8L���"O=���!<0&m�'F��"O���1�E������ŷJ(PD��"O�	���p���A�
�S��q�"O $YE�L
��04�R��ެa`"O���Ռ��L��x��ܚw�4�"O5�B�=0
�!E玷m��;�"O���$��	��@�B��s"O\,��,K�'�5�I�0J��ݙ"O`d�Q�Њ#������/N�n��`"O���c�30�0��Gb���"O
�@Fd�u��Z.D�)E��7"OP���:d�$[�4Ԝ�`d"O����5X"�\ڵ���.Ѱ�2g"On�2į!%�9�����hx7"O��,�$+��Ȕ&�zS�"O���k�Ր�rD�NA���"O~���o�JD� c% �q�"O��2��/��Tk��\+�r)r"Ob���#UG\�/��x�"O��Go�$J�@Wh����"O!�V�V�u:6Hq���7����NK�<��ˁ�����ƙ'�4�apa�H�<i��J oPlڃ��>�0�eC�K�<)�Cn��}�!B���<�Z�-OH�<i�E�
�@U*t�QY�i@�N��y"�@��^�Z��k�,�c���yB ןq���U��z��}pC����yR�o�����fM�@����G$��yr
K7!�8��`OB�6�&Ĺr���y"�^�9C�i��C_�-�<�"�DP�y���.+^���B� �섛 �8�y`�G'"��&�#W����t��}�ȓ'YyrR��3<��{�"č'}>܄�}�����c˰re�� �@�#A���G��ۀڋA�	�兗,W�h�ȓL�r�(2�'�,��.�.+M����.˔h+f�%c�Ƞ�q.�?�>}�ȓ��0��`�Qb�а@ F?+��4��Ғy�c〓]�P��� ������ȓ� ;�LDc�Mp�J9FȮ��ȓF��Q��<+|r����4Q��P��75�D �̓�2W�S� �	U�<��\�y�	
E�d�97�B������\���EW�-���
��N�fą�Oc����)P����3ʤ>6b	�ȓ5����5Z 
D���/&����\�s��Ug�H�m��/��Ąȓ���Q7��� ��t/ΔZ�Ԅ�{��Q/N3�"�x��
>1��J��x[� &"Z1�iʏ~z:h�ȓo�j���- �5`ׄ�	}�ȓ'�Xr�Dj��;r�ٔ,��A��i%\�t����bqΈ7|����f�3��*{�f�!Q$2�����w�S��;J$a*wL�~��D��`��A�١'� ���\?�ڼ�ȓ��g�*>V}��	.����q�p�w���'
�a��q:D�D�D�ɩ�����1�9@E#D���#(�"/�4�9cV�}F1�p$&D��Pg�Ǎv����S�S75=ڌ��(D�<���_)}|p�p�\=(�a�9D�� |��E$�\~m��@73��HD"O�=�46�ơA�/ըi�~��"OHE��I��R�n��¤S7]��W"O��X n6Hk���:R�BYc3"O��$a����A� �W� `Z"O�����S���AcB �3�"O�$"�ˍ�� ɍ�j��t#t"Ovd��g�5E����
 V��PY"O����B[�*�0Y��D�K� (�"O��+M�w3�taE���
!Ó"Oz Ȑ@۫|� 1�����=ِ"OLhPTE��\�
=�� �:#�|@A"O���-Y	^�� ��\��`b%"O�5 ��Q�(���3fE�����"O���D/y���fA�A��Ma�"O�)�%K�(�p��B�"Op���*]�_ih��eb�3��8)�"O^;��ÒA�\XsK�*+��8��"O��pr�C@�}� �-،�Q"Oi�_�j�T�CY(	ʞ�@�"O.mk��C�-{���	O�ڴ!�"O�y���1Dk���(��V���q"O:�3��T��4��'Gq<3�"Op@ɠj4!Ӑ��GHY	|>�<��"O�i��j��������#Tݮ�"g*O���`ʂ���c������T)�'� �K���?pԜ+�E 8i����'\@'���E ����GE;h�P��'���D�̍X�b-�AF���(�'XPbWe��Nj���ₙm��h�'���!�E�,BC�10��/c���Y�'A�jr�K$uڤ���ÝWl� �'.��(�m
�1��rg�Xb�B��'�.ґk0N�	[Ġ��a�\��'Wp�y��6x�"��B��&6P�
�'&z��$��8eg���I�,����'R�`�Ί!�����K��|����'_(S��[� ����J�]�z@y�'�xa24�"|6X��[�[��H�'X��s�HG�!�t�Br'�IL���'��Ey�f�k���!�M��(S	�'L�]�4���Vz���D����'����?Wg�*"��;UR��'+\�я�_"@�Ɂf��7͒�i�'Z�܂"gX�$*=B�'�5^]�J	�'?�yX���J/�ܑתӘP�|�Z�'Ğ}�e�U�\9�P	7^A܄p2�'�d"��37L):��_2D�:T��'������MW0�	@�ȗ2T`Y�'	�``��V��
m��%�TTXY��'=U[����`D��Ms�r!���V�I�������6�Ȯ<�!��;S��H�"�J$I��@��� �!��Ǿ9v���h�ot�bt�Ѩ>�!�d;3�3!�M�7�h�%D�>(�!�d�#e"���B�A'g�H�`�Aw�!����I��=C�l�`V�U�6a!�+@���� �\܀�0h��8a!�J�-Aba6Ȋ}�T&Ñc�!��PA赑B�W%���EHR	:t!�$��yYh�[��O�k��qa�[�V!�$� �*@�C�J�9V�
(l!�Dބ��1�mLYE4-���Y�N!�DP5S� �")�}�d��6!�� �I�"Y5]@����)̱��"O�tS��L>@�����7z��0c"O8p����/|��d�h�=�~�b�"O�h�v�\�dv�U�'�1��F"O�ء7�Ӯ=R��3��d�6"O����0 2%�C#@�'c6���"O(	)V��8���Q��/@����w"O��EOV�S2Zݨ��C:F�P٩0"OrEK"U�#�!�rm�0�@���"OԐӥhL�.>pr��,S̸I�"O������i���V���f�P1S"Op��C��+U����4m&T���"Ojѣ7Dζ�`���KO�9D�y"O����ß%0��r�d?s3@qt"O��)��k���2�=a�\K3"O���!A5!���	ƞ�#q"O�XY���[���S�mW�:�:p"O�=��BpJ8P���& @�"O6��ra˃�H�ǟBk`"OX�p5���>�T����C����"O��	�/��nBI��)66� w"O d��˔8t� �b�F�8����p"O@D"���7p��ūA��>a�6"Od��3h[�iA`h�Ӻ�4y�W"O���S�>V\��`R�fX P"Oh\�F��U���v�"~=~��w"O���P�յ5�:���>`%,)�"O�`��.��|�f�3�ܽ�R�3p"Od̛t� �b]�U�6<.m[`"OH��%Ϟj��#�I�]*X��r"O25P�&@����jEH 2"O4�Y�%�>�,h�"[c�DC�"OP�L�H��r� ��Y��"Oz����2#`p��֦Fe��J�"O~`pF98��Ї��j@��"O� @IA�m���e���Y{JX��"Od(�5L+��YU�O�'_&Г$"O �x&���|�k3c�:A��YD"OXͨ�Ϸ���)aT�%0#"OԥAc�G�E�r����}�:���p>yO<��c�7>|r��r�27\�`����t�<��!��^�z-��ҭ+HA�"�s��+P��<���9pHk�  �Ҡm=���Ng�<�Ҏ�&d��B��0�`1�bNW�<Ɇo�EB�ҡ�IW\Q�<iu@ �oʮh�qʙx/�(:S$�N�<�tM�	�H%���242����B�<I�KR�=����d�P�X��<�JA�<9p�.�%c���Ȕb�ŝ�U2�C�	����j��BR_��ۧonvB�	"9�AjE+\�  {����'�B�	�E6�C����F��mܲ%�6C�	'5[��ˀ�߂'�l�p5~�w��!|O���,�S�
%.M�**�0PE�'ݰ�l0�t1�q��Dz�����,B��-12����#PA���㴅8V����D4ړ1i���ӥ�Mzn�"W��lÊ܆ȓ"y~�9��^0Bi�?Dl|��u^T�B-��y����#+�9l	Lm��t8, �1��$8�9z���7`�Ԇ�}���e�O� xٱ��5,��%��%�@�j�h]�OPy��Aa���ȓ'��y�hY�x;@9 �iH⼄�S<���a�G�`:掞*����S�? |i��*'�z���M�$�04ٴ�i���.�)��}⤯�	4�:�A�I��r��h�8D� ��7��]Z"�^��F7D��
@�/유���џA��YQ£3D��*�"U

ZH�L��#��1?D�H�G$5�Є(� �2iǌ��g)D�\p���'MZ�@�L�m�r��:D��(G�ٙ:lXp���#0�h@�.D�p醉����A�m���\9��*D����U�=gČ�櫓0/����5D�󪂂n��9���B*D (��3�O��D�:��CS�k�H�e#��j@tȄ�RU
ݚ���2a���1�K\�z�Ȅ�6���0
ft���w�Du��Q��Ih?�(^�6�{�H�WβX�����'��I3�H��Ic���#��?<� �O#�zB�	�:jPM1r"�P�����b D�48�?iӓ\����Q�C�D�<����p
\��	B�'��]���/&��mʷ��<�Ǹ�yr'X�C�`I@�)o�’�I�yB��e���"��&7��<�DOI�y�H�>L��� ��:${������?�y��2\�Da��/��@�z��5�y2����]A���7�6��5����y�K�>l'Q�U�����t�E��yb��8c
����1�4($�؄�y�ĉ@��@���I��Hã�	���'#ў����{�Ç%��  �ư-T�p��"Ox��s(�2a���Ri\;Dq~���i�D������ēp���舣~����/�2|���ē[��D�T���A"�Q�R�
�ѳ�$#|O��� �,\�`6D����p��O���@[~
,y@��=⩛��6D���$��7�Ƹ�����{[�,1e"'D�@�����/f0���x��А��%D����P/H}�s��}���Ԥ"�`���OD�XP��\2:�	
�bU�-��a��'��ECP!�"N>hHk�k�8T&&����D+<O��(�#7?�ة������E��O���1�MyȨ��lԶ$ɤ�����]�<����."xu��F�5����ЩZ�<��a80����@]).�"1y�i�U�<�W���m:���'~I����T�<��E+^C,�b�%N�{	^��-j�<Q����@��Z��ވd���l)E�!��E���a�%�[� �)c�]�2+a~2Z������j����ɛ�FO� �&>D��b��?(�2�¶�Z�V5��b�g<�	�<I�}J~�gu|M�",q���&��t�<�`'�$όMQ��`,�`("LR�����y�^���ƻ4%l����P;���	L�-0GĄ�Nޞ`�ِ~���ȓ4�Ɖ� ��<I��[0�
�j����ȓ3��`�+ߙ|T"hq㬅%2B:<��BZ�1��iK�|�d� ��|��	l�	�-�@@p,��K�\]��-"�C�I)�ȱ�/0^G�HP�=���<����*牝'T9p�F�#7�b����C�ɭW=fiq���8�X;c�8;�2"?9��S-||�!�5�'B��H�Y�pC�Iߦ����j�(�����Nh�Q7
�<����	Q����$صU��U �a�4M���9ғ!�fEK6�T;�$|�O��s����ȓ��=�VD���Qk���6���I��O� �$�E��/��p�.ݱ6�ś��'��M~b!Fw44�
c�5|R�l{�e	��IVX��0"�8w y��/�<��y$ړ�ȟT��d ۓ�X���!�1d���a�C�<����Dj��r��/D̈ek�XX�\�'��	�n���Pe�Z���q�����B�	�O�d`��/\r��h�wd�0l�*��D7�T?8 �t�t�K`��$������/D�p��EQ��XI���A"��Y��$�O�c����Y��S��؋x0R�t��I��*D��ztC��nu���l�5�!�'�,D���R)��P��p�B��K�NY�t 8|O�b��C� ��w9��@��	�%�IS� D�p�Q
�4t��k3mǤ!�"Y�R�;��Ʀ9��%=�)�S4������8{]P��FєW�^B�I�^*�i� �:��M�7���u4������O>�w�  �&%��;2l2�Ň�5Y�"m��z�����D�D������d6LO���@��}a� B7l�2_�$���'Xў"~B�-�=Q��|zP�`�d�K��'�y�
eB|��!Qz�{D%	�䓯hOq�|9#Y�X�4�tP��" �a~�T�����e��!vV���4D�h	QK��$e�u��=Q$)%3}xR�ǟ�(���c+|	P�U"o�]��,0D�d3AIŦW���G�rN�ف�!D��rmT�rWp� U�L�=������ D�p�6��hD.���/́Y����f:D����Y�}"�X�k�(�"ȣg�%D�\
�
��.�F���/FGеh& %D� �0d��r7E�z�t�%D���%E
�y�0)@�遾/L`eP2 D� p�Ƒ�ZT�\AQd�&�I&�?D���"����L1{�k�f?D���'ߠ���D����%��y�!�D���8����"U��rET�!��̹)�`]��l�;���C�a�!�ē�t���Uj��G���*��ZS!�$�-�����/Y5��4��P3<!�D^̩q�J�#xD��Ϲ$6!��S��E��-�5e��@_=S/!򄚍E��i �N<<�
�jՏ�G!��A�}�(j�T�~n�Y�$��!��-�
ʵ�N�p�<M�Uȗ3!�|m�l��/N� �y�a 1!�j�h��	4;԰("�K�!��4��8�J�'9�Z �cnӣL�!��76"с�
��^�$�p���Y�!�Ē:a	
�S!!s�X���L�\�!���?/9�+� �%pn���+4u!�%ab~��&�T6:d*]AԎ®#�!��:M��S�
�S$��q3FD�!�d�=b��X2d�$�Tc��A�u!�	�@j��:$F�1���Ȇ�ɗ?�!�$ bJQ����:�� [`�^��!�d�B�&��P� ���P4f�-+|!���vڀU2��L9t���e�${!򄌅D���i��֏\	��qt��==�!��!E�^U�eC�`X#m5!�$�*Q�ԥH�oI(�%
G*�3r~!�$\̮��p� 1�D�"w�єy!��=%�N�2`�X�6���J�v1O(��V�� y.�+2���\���$:%qJQ��dɆ-�^�S&�^	~l!򤆃{6�Y؂ƤX ^��� D�]�!�� 8äN۟ i�Vo�'��8��"OZ$HiA8�"���)�y�T\a"O$�*D�D2vq:%����@6j�c�"O6�����%z� v�O�`)����"OL��a�4"z��b�	/p���"O�(Y�"
���`&��D�l�"OȠ�fK�g�E��n�^�^��"OK�{eR!��eX&Xt����5�y�*�N_R<9�oϏ_2^!ɰF �yR�N�~��abS΄�O}����%���y2L�4.�#�NY�;�Zp�h�&�y�c_�^�@JAnT=-�);����y� |`-`R-]�$O�A"�׊�yBB%"jX��C
-���33�8�y�M�)+s�Y�q�,B��e�2l��y⇀ n�*m�m�GM:@��ϝ�y��IF��#7j�:Ef�+�a��y��ۋ�b���Z�!(�eH�B���y2F'pv�}W%�,�%�`	��y2���T�lUl��},z�!��!�D���rt��^eP S�ٔ!�Uq{ؘa�gS�Ig�� ���M!�	0#/2]�n�5Z�^%��a�4!�'C^��2C��e�hŲ��O
!�D�|8�p���˨>�hP��1^@!��<@���8Ș!�N�Ũ�k!��){�D�����+�����Ş<�!�9P0�=qp' ��Z��Y�H9!��		-�\�"�۱����c��6",!򄀳�6#�"� B���L�/!�$�S��r�Gk�LP�!R�U!�$�$=���SĜ���%q���[!�ݒ5�D���6����o��!��6�ZXy0f�c3��8&�V@�!�$�O�6a�g͑�E'�a��#X�!��i��æ̖ ��l��a�!�Ԡ%�P�zpa �>����UƄ.+!�d\���#��6ov͊E�&!�d+dWb��g⑼*X�೰���!���O���	i3�u�b.A!�D^�i)�!"�]3:�3F�'`!�AB�=vR\n��"�D5*�!��D#lے��]�|%��7Β�']!�$��<SB$�BR94�i('*�6Z(!�ب`�
`�V�V|��w*��?!�a��y�`DR��A�#L!�DA/��!	rK,O�t�2��.�!���I;B�q��f��H��V0�!�D7m�N�C�Җa$���4�!��EJ������xS1A�$a!򄚕~�"���N�i�~a��
?n!��9\�l�qq�!}.ČK�hZ%(Y!� �G�D����[�����7!�d�&`���<@I /�q_!�Ҁ��m��Ɏ�K�F��#a�3|�!�D�'d�n1���Xt������R'!��"@���`�k����OڟB7!�D�H%���m#w @�S!5^!�$:,���(E�S)aH��"f�ĨJ!���P������y$�8����F�!�d2l��X�`	�B^ �� .�!�\v��#E�1��QSd荴+�!�dW
k��,��5�tl*�"q�!�D�3kT4�g�W��\��	�gp!�� \��DN��Hvv��r�^�%)���"OJ�{gA<q�q�[���9�"OR��`kԚL��ݐbQ[�@d��"O���%f���݁�Q _d�Q��"O�PYr��-u0�2a.m�qT"O�X�3K���}36"M�\R� i�"O�����F�� ����
Nh1 7�O�<:�F�4�0>��
��z� �*�/ 2;2	���C|����阼.�y��(Ƹbc��0�ĺaGB20�C䉐?��!ÓE[�K
(X��͗ �O H��M����H�v�w��	Ǽ�J�b�<AC��!7"Or�c�I�0/0N‚<b�@�W8r�P �bc��<Yᣆ�6����'�]Ę_����w*K�g�s
�'�*����[�H��"d
Us� -�O{}�	��JO#D�D)7�'�d��W�P�}���')6���Ǔ_V`AW%&���8����M뇎�*'�ͪ�D0490ks�<�V�DOY�"�hZ�w�i���Y� �b�oU,b��Ĩ)�'1Dt�'ܻ|���wf�2q��,"u �P�Xs8��7i�8F�ȓ�"PuB-��'����d��g�I,+p�� ��	xB�|��C�	�:�Q�܋4�)Ѷ�Muκ9ag�2Yލ(�`_n�ܰ��I�9���+�)��B��%KB�H�q������ZQZl��'Q�Q��'�Hxs%!�5������2m�PD�	�'\������,mwJ��@"��"OO���9~aJ$��Z�������v�v�+1���?ӢQ�g&�>(!�ɠC�,�`�KH��P���N���tI���$S�8�p��~&���f�Պk�@E(��Jx�8��l24��"M��p���a�Ԗ�	�D SӠ��pgK¤��7G�~  �	xcX� �G�V��D�:�ŐQmÅ�y��]�7��@�E�$F�j�mW2�y�O�1���[��ت��1Ѹ'sf�#��y儑D�T��	s���4�B�k<��BA8�yr��d]��]g�� �T)��C !v�A���%)�8��4�་�)�72�quBK(5��:��A`�<y �x_FMӅ$�(	��5 5�7�y���7XO��� ��Q2�u{ �[}S^}GxBa)(F\�	�A<H�H�XwG��p=yPϒ-W6½�#��@���	@Wb�K%A�6|���3e� %+�� !4�>U m��?���Q�H<+]D�i%㖹wJ���=�Qk\�&�R����W@�A�bJ��Ʃ{B�E[t���b��,��H�a}"T* D�c�k��6��M��\!N�P�m���Hy3iچ�5򱤎b��	S��7��O���]�uv�C�nM�0�i�P��	ўB�Ir��$�0	M2s�v�p*��jx4`��ϰ
��<;W���
���f��,�I�2r�xc�����աZw��*�I;4��9���;�O�h�f�$PDD�Ȧ���D��RQI_�a�Ԋh����D. ����څر��  �R �1LM�e�ĕG}"��W�=R�+D���(
vN�8|܍���S ?�L������4��*��7��xªU\4���-��rU�I)��ێ�~lLl����ro˫+�nd9u
	,��`�����1h��`��Δ�8�H�ل�4�y��ڄ_�օA�NS�nǐ=�D�P[��u�u�@�<���2O�M�M?m�-8��(���� ��"�䊂�u�a�.V�4;ZLmƵ1f�1�D̫4t	��A%U�plk��FEԠbC!�`x���"�<s��qq�o8Kz�  �@�����=0�)ԈT�����UE�d���n��)tx{�V6���dM4�d0��K@,<ђ.�2��I�}��@82e��h��ٶb���d�Rg��;��p��,�*���n��<q%퇐5�vXp�	�+|�Y��h�R�h$	3lFD����ؔ*�v��|�J>�G�V!ug�%�BUt�yل)[B(<1w+�
PqR2A�"<�䪐`����T%  ��C�
"��ٚU��m��k�8"�NE��ժ"z�x����愈{�[�R���a�&ի{��y�#e		�1�#"ś�L����E�%JEr���'H�'�u�?�0F@^�
�B�D��[0x��ջ%	�,a���Vi���yr��(��i���v!v���`�% 5�"*��Qm����;]��x��L<��&�%t$D���W�4��A���Oh<�� rM�Cf�@�N����>�����W�8g.I!�m8P���퉗&�h��V�*Q,}�b�N�Z�N��dJ\�����V1S\�زa��u�Ub��_6Dkt$�r$~C�I%.21�' 4��tH��&=�㟸�ф�1J;^lBd�@jN�>�C�.�D�G,�)Pn*5aӋ;D��Q�����V
�4U�x�&F����p�X5Q<��R�>E���L�b�J<��"1pi� �"	��y�P"�YS�Qz<N�Վ\��I�8�h�b䫜�6ax���u_�!��ϘGP֐�MC �p?�@`� @z̭ �$ا6z1���E�X�P��G�cL�C�	�{s��g�r9���V�P�@���>�g�A�{9���C,��\��Qu��!	#����ő�.k�C�1[�f�	ڂ�x�E���I�5TZ���Ć
;-�����	�s^�#\��Q�D���9!���J�.����%SC��ˣ�D
E�4��H��cf��w�\�.J��'hTs�Fֿ�̈́�	�S
�,���şQ=��������>1��N�K�V�1�C���(���u�A�!��Y�:����c ���^l�a��� Hp)�F<$xX=�Q�.Y��U�4���c�ȏ)	t�^��yV���ָO�����dV�:T#�n.N�f���'��H��߼L�e��Q'x1�|�-O09{䁂�B����6�Ԉ�j��'�nU����f@�D��jօiP���(��ڥ�_��P�R �\�C� � փ^۪-c�N5�p&'� �ք�enA	;����#9�fw��`0��:^�b>�	��i+ȍ�wÞ/��!:��=D�\B�'�7 ����!)l�˷����y`�]�c�Q	@�>E��I_*m�p���aK���ꗐ�yb�8IJ��"J�j¨N$��I�@�p	�D�I�ax	��+;t�#�LP�%(��p��4Ͱ?���R�R~�y 憧	����q>p�Z�nW�Pxr�G^D���X�u�ԍR��Oqek7��O�����߽* ����ӠD,��9�'R��c��F�(��7 ��aM� ��'�P��B� @��i9�Ċ_ZX��'[֩����i���Hg
�N�=��'6T� o�8��+��FV���'u����@�H5@-���DK�l�
�'00a�����o�ԁk�.��v�	�'�Ę��'�b���`֥d��Q��'H$��3萎4�2	�g�d�$�:	�')H��M_Z�A�C)��������AI�>�@�<:wp$�Q��|�<1'F��mz$�9s��sd�W��t�<��EN:�@=R����R~P���EM�<���V�8Z0�1���~��U	��P�<1�^#oe(Pr4 �+R�1��!�{�<I�j٨]�^ձҩ�F6Ld)�N�z�<�"$Acn�1+���X�D�9R�[t�<3N�9|��ab�O��`iQBXy�<a��F/���� ���Q�@p�<��!ԣ��;u�@��Z,z��l�<�q�JI2`RD"ӓD����k�<�杧G���6A��d1�ree�<�FbҵL>�S	����;��a�<�3��%�|����G8+�zmS Oz�<�2��+ t�3v�W������p�<�1�_K�� h �>~��r�y�<���ڿb�ޥȱF�M�.� dB�N�<GG�fA�	�s�M YP ��l�<�r"��~�ps֪�(����c�Do�<9�G�G��I!�M�����R�}�<��RB�.�c���&7�>���ALy�<9��ƬEV�s`���3�Nh0��I�<�#�ȵ,��6
_�m�AϏG�<1 "����Š���h��|�<� v��ƃ�#Fܘ��͓9�$�A"O⁣Q�@�) l��1�.��e"O��A��`s�)�ad��p�"O�T���\�ٙ�KK���S0"Ox�ʲ�Fp�-�E�ȱ��\P�"Ov�WI��9%@	���R`���"OyrCӥh�^<I��,l�T�a"Odj�o�2ف��f��D  "OB��e�cuZ�1ƀ� ej`�1"O���fꀚRe�Q�� D3;��v"O��
b
��6�^I�C>��E*"O���s+̲%�A�A�Ɋw� љ�"OX�/�.� �)_���	���z�!�D�Z(lȕO5f�4��F/�@�!���v&��Z�铑xV�ݡ1lܤw!�ߚ<~��F%L�=�4ˆ'<C!�d�Y�$=���<+�����)Yk!��5q�h����Ѷ/�B5Ȅ"L�!��h���.=W���% �
[�!�@s8��J#����	� !�d�$4���H���]��R	4x!��JVW��9�i&Y���aaL F�!�$̞P��]�Gi�@M0&*�=�!�	�5��8�d�ɐb�`�q��D�Y�!�d(v'\�:@/B�$���R�J�!��6j��4ӱ
�+o�*����03^!��Z���I=J���+X�:C!�D��04A���/�����@4\!���/%$Ē�mQ-{�ŁW�{m!�)3 i��*/gr�1 ⟊6,!��:L��T��=o�ذ�q��,y!�� o5�=X�IR6 ���2 �Z e!���=u��x����'��t��g�FX!�䞑U-�y�҇�f3��qѐTA!��\)�������(2�|(�'K�yS!�$Q4|��d�T�Y1�|j�\�~H!�dЕgC��	�G.p���4!����ܪ`j�R�0a�+O=/!򄏃�<1 �*G�d$T@���3I�!���S�E�� A0V�'U�^�!�DN.j0�Ycg�e�t����U�!�D��
$R�&�7<>���ݪO�!��F9J:���»Z���A�gT�4�!��"�f!��*'�ҨI�� 4V�!�R*�(s�Q�'��e#䈳0s!�ć�n2dd�7.M�[R�#b�_S!�$�L��'(I
hZ��B!OI!�Dx�bcϧ|�F��E�Ι _!��F�5EjU���r�"�ҧ��"do!�d!H��OW={8�����7nT!�Ė;0��u �&	&^0T��1n��t@!�ʵ2t|��B�>6t�T��� �!��*"�fB�<c��J�͹Q�!�ě�r�N�s�>�E#�`�6�!�<���ۓ�=Pg�К�A�:{!�@�k�& ��90�X���"Z!��K�
]�Ʀ
mr����P��!�d	�8X�J�:(o��c�@�-(�!�dY�o���DA8���Q���!�V:�$c��C:GXA{�%T�3�!�d�\�P1���X9�p�dJ�U�!��q�
0��X )n��u��/e|!�$F�f,*��,�y�.P�5
	�T!�$��l"�1*�B�$U�����;�!�� b��U��$g � +EbL����@"ON�;���PA�|Zbπ�ռ@��"O�1ڇ-��cZ\
���2����"O��9p.��R�B���h@��P�X�"O�Z#�!i'�] 5FΒj�
�!r"OZ��G��lY`�98�x$Q�"OB����7D �B�^�"�;�"OR����A�!߶tS ���$���3"O1�g/H�1��B���^��C�"OЭ)�ȇ5!n��q�6�����"O�Т,�2Ղ��IN���d�O� x���0>�UOM*p}�UA	6U��eZV��U��Z$��3xѨ��I�R�|���)�J����œ!�B�I�;et"P��������$@&�O���M3&F(��3�G��H��H�'�9E5��a�b�P=��"O(�5�
Y�RMC�KZZ芥��N [9�h�ծU�<��.J걟�'"D`ұcZ���J&h��zHV��'#4���EV�3R
D,��1%��bN������0Ut����Qa{B�_�(�c N�=5�	�����p<	�N�:0�d���(4 .��ߴy�����W�xz��a6�X�ȓ<��5!�����E+g��:��ȧO-��NU�s$���WG\:E'�"}�aFL�aE 9ƍ
F�Bt�J~�<Yw];m��!� �?_��u���p�΅��H� "	�8�n��}&�0#r;ug�K�O�r���ï?����H�@tȳ$A�h!�Q6b��.w���OE�:GX�FP\؞����͆Q��9G���4H��)OB!rgH��J���i%ir�ѬA=�8K��ܮ5�b�K���ya�p���8êU0 /����6��	�aRL	a�n�.��S%��=��e�@+\!�/)<C�I�b�T(N�q~8!rKٍn�$DfA�C��-d3�����L<�r���Ԍ��/Ƭe220QAGh<��=F����̊d{FaL�{I��KT�#j9� NlS5n!x�V%�X���'z�  �.3t̓C@���I�2uf|�t(\6�0H�ȓr��{��G0p0qp�³ʾ��=�#YcSj�S�e=�'z�*ᚥ� ��3G�+JV4��Ht��R�� ��1aB9l�фg�$&��O <x��Y�Z�b 2G��T2��.V���:q�(D����r�@�2�$ =@�I��6%��t�A�/��\�CT�%����C�U�m��۽R(� b��zR�7�p,+.�e�� ��2 Q�D3.�XK�@,c�Ṟ!
O�Е-%\�iОkkX,_1:%�=q@a]����P�ˈTo�)��:�Ӕ!(�<8d�r�j���\%)�B�ɪ1s,�����cfJ�Y��[8{��2cgR�@/։h��U�&��7M_�����l.u16�ъ}� ����xZ!��iϔ��(M3c�M�e��O�	+n��<�@Fۇk]�U���'�\``D��P}0�M��$q��8	��>7@�qX�>a����$mPD�'�/@d�M��3�b�U X�r�����T�)� 3R-�p��("
b>ћ���^��걌�?�Դ�"�:D�d��hQ-E��$8b,�W[J kq-�� �$@f3~��r�>E�t�]p�Ȉ(���$�b��a��6�y�Ĥr"d� �+��-فJ��	CR4Uc��_�?[ax�Mr�`���*JJ<�QT�	x�vl����,�.���K�&�Rxb,��#v��k���3#� �HztB'�D�=`R�0�N��*V��D�I����~Z�����~�Y���2D��Ke�E_�<1Â
�XF h�/��9���X��n�<�4ď���쩱`I��2�$I�g�<�3��ZiH�A�.oBD�hW&=D��v$^�̽�uM1#�BQj�A.D���c넶e�0�A�i#V�B��E�,D�̰��ٹ\�P����WYL��r�'D��`��Ÿ5G�Uyw�[A�`*A�$D��  ��b7�<]�6���H�6Ȱ4"ON jm�MY�3�,	4A��	�"O��Ā�H�z���y.���"O*����2�
��� �H�J�s@"O�EK&E� +����!6&-C�"O�E�)C��H���5\Α���'��M��D�S��1A֢H(=���N�0�N���v<���W+���G�2'72�F~�	!D�pH)@�ɏ�CL �ZF�����O !�$ҳd:��kg��<��x�j��ܻ:���7mF���)�'�� z�N@�AZR��懪tf�u��b"�:A�ɻV@Tir��H�ht�O���R��7M�:��Ó����D�:4��z����2�����I�?bfx2c��l<�7�7X��aQ�A8X�"��aO�DN�F�>��"&V�:o�E����B��y��?/`1��8���{x�(�do�m@�l��"O�,��P��tmqQ��,?@���OV� �Dl��D�<�O�:��#����@��9`����]�P��"'�O��8����(�����\2+�6��C�0�t��ү�>q���6�Y�%O���U�ێ�0,A���(WW�b����Z ��`�ʃU^��3�P�q(�
V�`��f�TF�r� 4��I��x��V�z|0"�����I���O��~�cm����͚u}��!�X{��I�z�xc#Do�,^#PR	�'�V��a�Q�[p!��f���z)OL!w��^��5zs�%�d����'V�Õ��<����R�O�a���A�oh,8���e�:�G�܁+�������i��#�	s�R�Q�\4��
L'ujN5��a2�1� �{%H�!��b>=r5���S%�̡�%L�v��0�Si1D���%$7WݾxA�NT���6����ʖŊsl��>E��D٨`<QG�E�p� EX��ߖ�yb�_�2�����Ip�9×k����1�J��;vFax�����8%I�����Ib����?I��G3?�H�b�/=/��+��p,�6�
�Px�AD;/k8ehGF�3�~c��R��O���᝙��O<����Ď�7F��:��!|��x�	�'�l}�f�K�a����;q麄i
�'G�-��n�[�f����(_��9�'ɪs�j�9u����a�Ĳ{�0���'dH�������0���Od, ��'����
/�챨sk�<h�	�'_0`A�d�1��P֏�(%�j���'8mC!LP�Ԡp6D�:ʶ�h�'�)����_�4�+���>{�d���'��e�T���@�p���$�8��'�`�)0n����Z��H�(���'�ܬQ�^����aS�@��I�	�'p(�)Cƚ�!d�22��<&�b�[	�'`�t�P��={����A�;�h��'��#�0j���!C�����'1�pw �[��Q "o@�Nv���'���@�K96e� ��P;r4	��'o�,S�G,��!�ш��ҬS�'�8����!��괊����2�'������-O0���H�qbd��'k�c,y�¼QÍ��s�H��'l����IO� �BXB��Py���8�'ubݙEk�')��*����T��
�'��؉�GѪw�yj'�֛i�yb
�'�RE��Y�0�=��1?���'GB�[��	�X
��
2L��4#fM{�'H1"�l�n5d3R��0�����'L-��Έ%KO��:�ݭ?�.`�'{��r"HH�Py�`(���r�	�'*���H�)��"Q��"s�zts��� 4�g@��N$��$��R1`Y�"OjT�ɓ�R��1w@�e(p���"O0H3��0H���ԠS�Hq�"OXH���YA�}X�I:r�8��Q"O\����!B����DO���QY�"O�`ڦ��|rpȢ��00�~D���d�7�`x���%j%t��0��+1O�ͩ�̌�z�	8pI,�`��"O:1�CL S����s�S���F"O���զ"L�8��@� 	��@ "O�-�u.�SS� "E�	C�j��7"Ox@�Ԋ�>g|�u� %K��f�j�"O܄1���'9�4�9�m�q�y�B"O\mR���-y61�c솣ng��A�"O��rA��m���rk�?\>j�"O4�ρ(hI2�5@FX�Q"O��QA%&B�"�q��&�|1	2"O %�P�Ň;v����Ǜ�T�Q�O<С�.�)�'DH\Q���  �uP�d�b@�u�4��%<��;}�INZ���)�2t{�fQ;Az�i)G!�%�p� 0� wy��\����S�
�䨛���8B"}�2NB�.O��(O���E��	 �8�ç/L*��a+�!j�����%.*,}�'�UӰ��&>.uYq�;�'/M(�C��~��L��/��S�����Tӛ��I�IF$T�m��Xa����0|j׃Tl��|�f��<;�,�Sr	�ɖ썇kǜɻ�����ӊ�\@�P�>^�չE/�#O
R������ �a��]}���6��CWA[`�R4 㮼�d�M(|�>py�!Q4w,A�'w܀ʧ�O��1Z�.�DGt�eD��8�f7u�)r��J"#;�Ͳ"�x�s#�;�
�k��(gӴ���ʄ�7Ϛ4+S��8&!Ȍz&m۟Y�NLp�	32��)�~�v��p�)^���X�,T����N�.Δ�e*��@A���Pp>�D��I���PI�5h��|c��P�nAv̓�	Ϙ�fX�vI��V�����	u]
�h��
�X/4��D���q�j�l��>X���&v��:$�1�f���"pl=���)�����>qVkE�>S���˓pJ�US'̷e�^@X���t���@��fʆ�y��j�'�hX��m����DR!�:���ŠM�5��{H��˳�=AL�-�1f�_�����zg�T)0�DE�A֕OQ�ȓF�����|l�<�3#;� �ȓ�(�e����D�(7�D�g���ȓ��-��F^�;~���O[,C�24��N��uO%h� y�w鏱8���ȓ��0����-l�Ĝ�w�A�~)�%��px|�t�[�L�Qς X퐔��t�J�P���lOJd����%6l�ȓ*�a�T�Ԝ
0娃��"(T�u�ȓS3.�Zś".�\�xAh'XT���ȓJf��0ЎN/*G��zBgA���ȓl�zr/Q�%����� JV�nq�ȓqZ���D#� E�Fn�,E�  �ȓ���1����X`E�M�Z��ȓ���&H��9�@!�M�.$wz݆�ɮq���S���A�c�ʴp�-�ȓɂ�!�"&I^��D̰y�zɄȓR���S�U-"�8���Ù�1G��fQ�d����gG ��� �sG�Q��^��y����w�x�#�"aAj��ȓ����dւ�  �1Ɯ�K5�Y�ȓdB��fb .]1+�@^!R�TH��(���[P�
�X��,V�&:�`��ȓq��I�
_��#��G�^���me&�X�.��S:���P��P��a��7h��K� ���.Tb�ރ!�Ňȓb�H�)�	�I��t��j
⑇�}i�r �6��(`��"��ȓhX !Y��$!Xt� B�}�$���S�? �EK��ќA�8��s�6���"Oz��6Μi7nI�`딬xϬ�s�"O�I�A�/!Z�@��j̔l�HM�"OT*�!ܚ٤�ǚ3ѐ��"O��Z�Z�o.5��сV`@dpS"O���vIF��u��:E|nA�3"On����E�\�`�I5���D՚���"O�X����'���䈊lZ�PB�"O�	RQ

�7��J���Wd ,@"O�DbkH�st pCFlg`��X`"O���vϗ�5�H�!k�i�0�"O��"�DU�H�\q�����,�"O�pJ�@�ut�1��D�#�ޤ�"Oz�� *U�X��q�敛z�~��"O�u�kE<��)���I}��Z�"Od%"��"
4�"ΩN����"O��x�Ʉ j7R��aش5�X�j�"O@\	R�ғ!�6��Q U, �,Ղ"O��ؗe��+��Y�4��"O�����D��1�5��|@3�"O�I��I��hU�1KF�+lf�h`"Oҹ�鄁7d��1'F�]p�"O��#Q���m�`����=�$ݳ�"O�m���<M+t0��-�hq��a�"Ob��"�V���#�ZϲA�"O�J������x���h8�ȓ\r��ϹAJ��aC԰~V�%�ȓ�|��� �(+wXÆ�+�:@��x:�yŉ:`�h�rrlV>h� �ȓ�P��I���"7`�\���kL�1���1=�@���Փw���h�n�@�� �g�2vlB�"O�T�e��6|�vI��Y���ɤ"O�}9�+�'�}�BG�&�T帢"O��� -�	V�\P1'�A�-Su"OZxz��X���C�&�<Z�I��"O���e�2{"e� Fܒ,k�-I"Op�6'H����9D�ùr�H,0�"O
 kc��'%E���m՝[���H�"O�9B��1���4KL�Pc��Z7"O��(�K�:P�f�!�)S,$�R0��"O��U�o�@�{��؀/�z�Q"O����H�P�HH@�бD��8�Q"Ot����$q��0zu�$G�q)�"O�a5AM-\�@}�d�1~���"O�@n�v[�2��ٔ*��y��"On%�����A�$Q���O�����"OH4�g�	�8�4���X�,{��S�"O.�a`@U07��a�g�Ǎn\��"O~y	0�B�?FDR��#$��=j�"O��*�f�2CD��UNT:��]�!"O�Q&�M'D�|$#�� w ��p"Ox��,!�XEi!�d_R��"O2tt;ӎ�q�k�nYne�1"O
|��eJ"Z�l[F�K�_;�A�V"O��7���<��c�j
D3��1�"O�5F��BD�s��*F4<+�"O ��� �&W�` ����+n#��p"O4U��Ć<���"��)wЩy�"O������:������'sD�"O.���} 5ʄM��SHZ��"O��a����#��
�O1��1�"O6�1 Z�`���D��v�XI��"O�u��c�k� 9Qd�J2�Bq�S"O� DL�`�H��n��ՁP�����"O@��Ek_�9Kh��U.ʦIx4��"O�(��G��@Z���� !e"O��7��;�֐0�!�)e���"O��K,L6c�`5��� D�"O�(Q���y����]'9��"O
a��.�N9�����X��\�B"O���D`L�A�� ��mX5N�rQIV"O&E���҇O�q@�ݶ2}��Q"O`�� h8_MȬڤÒ/�n�a�"O�	�Ԩ_�sF�i�GCL�n���H#"O4�B$�5<�1Q�L�6�r��"OZ�٢���!V���!Gb�UjG"OH����64���a1 \R�8�"O"�1�b�Y`����e��"O��7e&c
N�k�'�C�>4S"O�!�-��i>�}��G�")Er��c"OuH�H�A� �16�S V?@���"O���3��t+��I��\���"Oj��ѝx���s�#�,Rj���'.�B��sB]*�#�.�|�K�'����CF��lo%C#�3{���'���c�g��%�@#J�k^y�	�'��)A� �L�����	�'��1'8��h &	Du:;	�'+���b��X;��7;��d��'��9A�i��.�A��?A�m��'� ���
�=2B,1!�@�0�c�'�U��NF0f�`e���+$���'S�=Q���&e�jc�˴y��p{�'|�|#����J��2cݳmD�� �'�&$��Cн}	&qS���dv�U@�'�L���I�^v-��Q־Ѹ�'ي��6Ĳ�ѱ����$�0�'�f@�}-z}�!�ޝ#�6�"	�'��D2gN�$ת���æD����'ZDP�.ZXG��1E��q�'R�h�S�b���S�d����j
�'��g.��g=�LC��ԥJ��	�'��� S$�=zЂ�C�مH�R�	�'��0����-2��r/�?�:�8	�'
��cE �6��X�
\�8q����'M�q�d����J�$65�i�	�'�vH `+׺;-
���4���"�'�������"T:�c���b�J���'ۦla���4<`���T6Ĥ`	�'����m���`�@��bk����'M��J�H�-�@끅����'�U�u�M�PG���nYְ��Ib�<��L��*���e�D�w��w�<i�L,���rh�	��52T'\I�<�dC�x���N)3��9����[�<����0 Q�ʁ�)�4C$�Z\�<A'X�U��(��4�vp�7m	Z�<�0H"c]���B�QZbе�Q�<�ԉPS� TP#A�*tT���J�<I�狺�jA��Ά�+��l9�]M�<�O��$�[&[�^i)ӌI�<����2�4��6C�q�D<)��\�<IףE2k��*�,Շ��i�AAX�<i�L�/��I4�C�8�h���QM�<Q�ɟ�\iC���v$�&��}�<)��\"�d0J>z)����u�<�U��"�t����� �4�	�)�r�<� x��2 Q�s߄�;5!]�hL�l��"O�$�W!!R�б:�`�^�T-�4"O�15ǜ4!�0ා��1'���"OL�0�ŝ�j��p�t��8W%�""O�˰BÈK n�i�P�H�@�"Ola��'�	��:Æ�P��Q��"O�\�0�K�`F��`1�̍z��Q�"O���4�I�8Ȕ�ƈ7`�V"O(�;��/Sm����FQnKء9`"O�`���^[q$F�[9�U"O��B�/^ R���iZO��b"O��G��_ޜ!�R�Qu�*O�$�e�:&.� s%U�nq�a��"OrA!�N�VZ�z��6g��kW"O��Z� ߈O��T�n�&�Q&"O��R`a��`}ޱ3&DP�z�"O>�hG��]��I���6Q�	"�"Oj\���l��,�E-�	s�8��"O��₇ :�ݺ���/m�J=�D"O����+f�����\�N���"O4�J"�R�B���6FI�q��a�Q"O���CY*P��ׅEn��"O�A�aO�3A�^}���Ͽ4u����"O�}"R�L�>4�[RNӲB�)8r"O��g
S�`զ�m�+K�S�"O4d��F�Mf5��̍l�j �'"O� ����;0-|a�񋌍w��-�$"Oh�4�
"p�9�)�'E���Y�"O��ɳf«%¬D�`I�&#�29��"O��x�N��*�����<3����G"O�p)G��(u��V��Qv"O�كEY�P�@Ę1k �E�:	�b"O��  �Xh�Q��J=s�ĕ�5"O`�`ǃM4~�����Y�tX�"ON��E�?�4�k�F�a��q{C"O�m��   �P   S	  �  `  �  y&  4/  v5  �;  B  TH  �N  �T  /[  ta  �g  �m  ;t  |z  T�   `� u�	����Zv)C�'ll\�0Dz+⟈m�Oh��5G��DB� �8��GPz�إ�7&=Ĩ��(C����AL �$�e��I�{),Ȯ;\����'{��@��'�tp�g/;�ԩ�aIg=ZaRFT>*��m@�I�5iR^�i�7�Ͱ����LsA�럒�D��.P]!4Dљt�rh�bO<[V��X�̈́�JZQ�	>�I�
0
!���ٴ5x���?���?I�'�2ubAC���V�Z3m�j����?)�%�>K�R��,O����"o*�)�O�牵s�v4HP.F%P��l���ԔZ��$�OJX�'���'[�M͗���z�t�jBzLF�H�*.h�89�r$9D��K�V�N����,�� L�O���g0�A����Į��u�㙖/E�ٗ'�<�ӣ(tI�D�	�
�ry*��'�2�'���'���' X>���'%���	$��h�
�g��{i�@�I��M1�i\^6M���	��M{°i~P6��A��5s��(�O��ɩ����zp9����9�ȟ<̻�	Γb���*�P�b��%�ƚ
c�\;��ڏǤ)uiv��lڊ�M������c�-Q��T���mx$��2Of�⡃����?��-A(/b�=`T�:@%���#k�q�(�r��OZv���d���nڥ!x4j�n�0��+�+�|Dۦ-@�*O"uK�+^�M�v�i��7���*�c7/ȝt�6H��#ާD����~#�\ &�3݂�� ^�}k,�7bH�db�$lZ�M�$�i^�51HY1��x�;O�4�%*��[j�Pye`O�\ѥl�>-��D����Ȫ������3H˲��	W�:L|a�%
B\Xa���%;@aB���'�|�藝���%�XM�0"g��(htd����$�y�B��hb�@Z�!�� � -�y�@�?G���8�瘁E$� ��y"�@�Q�ƑSU�L�	���3e�y�+L/t�0�!�W=s�F0�'����yҭĤ[��p��ĥh��9�EQ�hO҉����\CZM(�������A�4�B��6f�Lбb��9���&N�:b��C�I�A0}��/C�!
�帧, @�C�I�(G8}땨�>Q�1@+�(`�:B��"Ze�0�=o=l�F��"WB�	�NP����
<��ȡ?���?!��"~BQHN��ʔ[Dj�X/�li��-�yҡ��`��T:��HJ�̝��D�y@�	�����j:>��0 �)�yRe�C�$\�Q�2߶U�M���y���+�`�'D7W��t`���y2O�k�}RSA]Y|�9��lǉ�򤒺
��|R� �5VY1�M�WYr	�e]<�y����}��MF�:W`y_��y�+2u�bj'�r蛢���y2i[�h�t���ʎ�d9����ybؕ_ Ȩ�QI��\���Њ���<�a!X�X���'���
k��,A��K�4�|���!K�o��'�b�Z��'�0�X�0@�Z5&�<���'jp�EHW?@���8����:�̹F��#��MF~�HI?� H�g���?�ܼz��4�ɳqq�
snt�L�7f�/
X�D�A�P���|���m���C�ウzhݹ#�/��=HDC}y��'��OQ>�ZŦ^�~�|Ѹ7�ʿ,$��g�'�O�i��A{0ժ֧ (+R��A� 4%��d"�d�4���C�9O杣>cV];aϖ4�� ��^�c��C��%�����ꂍ,���3̗*9�C䉞g&�[,��up|j�!��y��C�I67Q�B4]���!+U��LB�ɵd"���%|<0P���9�nC�	u�4P05�7S�8�����E����ܺ,��"~Ұ�<vI��F��#8\����y�&�'�f`���#|���-�y�fC"��!2���%B�yEK»�y��/���:ŁR�|֔� ࢙�y��E�gqF	rE��w#\��Ƃ���xbe�6&�����! 21�T ���d�ze��'a|��VN��9P��B�rV�!��߰kdx��'�&�q�V�W;���'+uQ�F⒫�xrGV�U�|���6	`�(b�%"n��HA���2d�y��)��]u��#���y�,[�M*��8 ��1��r3��n웖�|R�B��y���$K%���+�w���X|I�?O�� 3�ٰ:���O� ¤�tMěc3��#$k\�0Z�&�'q�
b���n��'̒���+5 o�M�hS�|�
Ó_x���	��	П䚂��B��!θ	�SDPMy��'��OQ>9{gB��6����'��&Q�m���$�O���	*I��)XD�&B���u�=3r�$�<�AK��?����?i+��a�� �O�Ms�퍭d(b��z��<s�e�O���1�R<��B*W\�b+L�dg��O�S
��K�H�K�h��I�H�6a5QtLx��#��8n�Z`��_�E��=�O�v�
�J=(������%m�D��Oũ�'x���<	�㜉/7j Jgkʍi���J"�`�<1��	E�R�-�$ ʈ�+]�'ۖ�}�bӼM<Ctk�* n�kĠ��D�O��$ g5>59���O��d�O���l�a�e�)G8 �;ԪQ�M- qiՁ��	��M�1R��z�O��l��/��v48�Z��Gˎa��1Kh��bC���`|b>c���PN�|'��b5EZf,i!���OMm��h��L@��x�|�'ra�+o���d�+m����U
��;^�{�����p��:ڊ� �(��Fb�,�M������������b��9 l�j1
�	�Ŗs���jcT��$��/HEc�%D47}���F[�"�!�H	fl*����/`L���$��!�$@7CE�X�2IǶbJ��5c�1�!�d?:��u)��d/u��Y�1�!�DZ*S�Z���
4N���r���*��}�GL1�~����x*���1�l�r6G/�y��٧j��)1� �w����6e��y�!I kH�f�Tl��LBW����y�m��z��D�i���uaĔ�yR	2,]�ѓ���2C6���ޔ�y҂�HO�����G2@X� �$���hO�H[��ӱ�Z���$^3K�KG��9Kq�C�I!j�`����<��! P�C�	-Ga"�0�ވD�b���p5�C�ɨN�Cd`�.#jk�eXbZ�C�	!�n%	��X-t�� �-�0Q��C䉕)��ذ���5,�U���
� ��Q�t"�"~���Ŗ��bRO��Q�m���y2� �6=I0�
2�mZV,5�ygԝE�,a�֏z<x��Q�y�AC�VN*��k�̨���T��yrbU�]F$y�rmƸ_:5hd�Y��y �<�"�͡.�Ͳc���DUIx�|��g�t1����c�湰�œ,�y�F�C��� qȑ�hs&�iRΑ�y�*>F �Sk �(��I3�yr��@�u��̝bTн�m��yBbC�O��M(���0W��)��G���>�c/�^?�l
6Q������<$r�Ec��o�<	go�75�p��	�l�MAҌ�h�<I�4��Cυ�y��Pd/�f�<I����q�P3o@�Q"}(V�Qn�<�e�\[4����oڄ}�l�l�<ٓe"�dupц� 5~$M)��p�'=����i�2cdc$I8�^�3�#�)�!��+>Wr ��ȁ�Y����'�Q$+�!�R�_�<���O������b·s+!�Ĉ+�NQ�1j�<?v ���AB�R
!��<n$�fEܷd��"b�3r�!����rH��4�K2T�u:v ��r���O?! KG(h��5��cR5e< 	���P�<Ir�C
0ӈy���΅2�֙"�O�<)�*Ǣ	�l�3�H��@d�g�BL�<��B<g�b��be�;g�5 U�SC�<��I�݃��CZ��е��i�<��&З�B�p�G2{��<JM�dy��p>�1���|X���E�	�ܪ�B��y
� V��������3B# gY��i0"O(���U�.��Mar�<7bdȣ"O�ݹ#M�	�����H ^���"OX��e=1����u�/?F:t�'�����'���R7a�?���*_�q��'F�ٚp卹& h�3�T)���'�L}��i�-v�s�i��c��"
�'ւx!�� {�T	���>#��D
�'���x#�R���Z�ߊ1�(	�'+v��v�Ɩ[ԡaӤ_"�����D5b�Q?i¢a�:F����F'L�]�0�8� D��b��M�� �c�]�K�,=	h2D���1R������ꂪ,D�̓�l�5E���E���g��m���(D�t��`V=C��:�M^)irFlj��+D��藪V�P)@�g�\�Yn&`Q��O���b�)�ZL�a{�̃�)�dI��%�3 �>$��'\�!�P�[
�U����t��%8
�'�(D��o�;cEŃ�G�Ԡ3
�'Y�q��� �#���g�<Y	�'w����C� ��6"�*�Y��'X�P5F�2���Sa$��� x�*O6)I`�'戱��@��Te��m��}W@�
�'X�L�wk�w脅��eX!,��Z
�'a�� �&l=�pчI&�
�'�@4��,O�$�"�����i	�'�1�O��;�9��Da/�����U�#z�z�E�o:��A��-L��Y��O]D�s�*Y7D��(g��)M�9��o�tL6 �V���h��k���ȓ=>x�*�˓�p�j�92�,��(�ȓ^\`��6�)�d���愃u4	�ȓc'�u� ��Fy���(�<x�5F{"6���"��.�*���.Vu����"O<t��f@c=�t�Gc&�d�Bs"O<�if���.#�d"bl��denL�"Oz��A>��P�ԫ��{��\i�"O�m�TĎ�����P#�d]QV"OVɑ"��T�l����D� 	���'�f���� �@Q5ק"$j% ��L��ȓ,���[��>�7!M�Y��ȓ��T�a#��xdH"狛�z��ȓ%�x*"���Lx�`��;@h��L-8,k���!Ec��B	Y[b����s{��P �;�0B�*ȩI��'��8�8�b��틊P�a����1ĠH�ȓo��2g�A\��q���"Zi蘆�_U&�Z�_`���C�ڢtB ��ȓ:�D�	�ad�\�0��T�@����A\:�����z�\a0J�5:J�-��I�E�L�	�c��CU�E,$�lDr���-]ڀC�J`V��nJ/oBL����#7RC��
V�����U�e'4���#z�^C�ɴ<_�q�6��`g�U��JF�%�(C䉔~��Q����'[��P![��B�I�]+�Oq�~0ȤA38��=q$�x�Oh��cO<]���Z�(��(�� �
�'� ܉�μk��S%��� >A�	�';�Y�wٮ�p����g���y�	�(�8���BR>y9J�	6���y�ĖhhR���"j�������y�fC�\W�����U�9�z�PA���?1�*�a����r@��q��X��%1	(h�C>D��rĥP�W�B��'P�\����M;D�� fH;1��X��4��%�u��X�"O�e)�@� ���p��P�� ��T"O�@r`N�s F@�vc�!�J�h"ObI ����kz@���a��;�`�T��2 8�O��3�j@�`�����D�z&�"O&���G��Qт^�4ܔ��"O�����L�n����9��!e"O���E	�/~Ֆ������&��G"O(���#��a� ]#D�	��'A���'��d�VHˋ\Ɩ��7BK�[���'`P3%#ZG�d�Wd?*�"b�'>�5*�%G=O5 �d�%|�y	�'��mP��^0����!,�tw<`b
�'g�����P{���7�:p-�)�	�'�
�1��~�(�G%½��mӉ���}
Q?u���
$�d���\��`�! �$D� �uˀ�W��`�\=n�^�i&�$D��pe^�b/>,!TJ�fKX��b�!D�Ī��@�U�����o�cĊ��$�=D��Z����\ٚ���=K���d�=D�, t狵<�t�6�W<b��&N�O@�0d�)�/2��@��A�'U@��u#J8V���'��4��'ж1Mu"���X�J�'$��e�A�v^�t���P4&��'�&ip�8	��f��5$��X	�'N��۶��
������;*�9�'b@�`�	�e�<�aE˖�<`{)Oh�	7�'�j;�@��/kU�Ȥ�t���'\|+fͥc�:�e�6Ɔ���''��ۑ�S	4!����Ϝ�H�`M��9d�!��+0�B�H'��"4��ȓ��Q+���U��@��Y��Մ��� Y6�I�$ i�t�?f����Kz^dB��#=N<�"�dS\��j��͚,`B�I�
�"0�k�]Cd����.B�I�����,�f�[F�
e\C䉌7lE�7e1%�TՑ�	�3�C�I�%��c���h����-C��P�=�f�X�O���)������C�/�ձ�'S�4�*#pN��/ӳs�Z�	�'b����IW�5�}�!�-n-�p��'I@�yŢ��T$`����O�r�	�'��,��+Nzx�45T�qB	�'�N�B���.|��� �
� �p��KҀGx��	M�7R(!�!Ł&/$��C�3r͔B䉿t���"��+^��'X�$z:B�I�;�ht����o��C���}��C�I��)t��+4�q����%��C䉃A�V�Q�˭w(��"*�:r0�C�	�+$�i`F��S7����C�_f,˓I�� ��I�O�Tak�,�B��b-�9�C�	�w��h{�!� �2��N�8RB��=k1��RC��]��آ@ML�QcLB�I�=�1�����-VB�ɪ/�Xl�� ����dT��$����5yz���/���ڧN����0`!�&4W���@C5;��i!�W/Y2!�$�7��X`� ���B��q�.>!�$]~:D���'�?��	Z�� '!�d_�w��$ �E�M�2�*�
Pn!��/#����-Ŕ,�tiȱ.˷\ў�[$7�_�v�jwi!1X�1�V�Q�����+�NĻ�:0������E
����(��(�d�/#ޘk��%6�,��S�? ���į��#m�L
uk�((���*O��xA�\|<m+�"9	�����'V��g%[]ny)È�p��(��4�ȬEx���Ҕ+Vb�j�FP�2 �,�4C�I�������T�ڹx���3htB�	�"TJ�"�!u���_�3�jB䉏h��IH#$��5��a�h�/_h�C�I�N�4)�ՅR'	:n]k�*�
`eC��.hZH@�ʫ�PqI��@��ʓWP����	'm;�P����-U�JY�jޱ��C�IqH�
\�N�t���� 0H~C䉩9�2���$R�O���9#J�s�C�I�l��B�oT��v-"܊b�'�nI��	�V���b���~)�n<����]��XBWi��' U��f�H��ԅȓ5���-�C4��!���h��u�ȓ4�Hx���S�cp(a%��&��Շȓ]�h	�hɱ��t��/ ��ap��] F#䀑��Z:/�����s��iɦ#�y�r�*d�C6_zZ�F{�%�������ӊ$0��yp��;q���"O��V.b�D�F��;CeZI�u"OtH{%ƃ�B=y��ͯW:\�3T"Oȼ�S �:
#�hja��$�8�T"O�᫡�bht GL4k��mµ"O`��f��-,��K�?p�(�bQ�'Yd 	���D2�<����8I<��o���x4�ȓn�F�G��{0^R@N�5s"n���`e�pS�Þ? %�QR,�-k��!��!�$ɳ�SmP�m�2R�$�<ćȓD)��+�〄��$�D(�Ɠd�:W�\���a��C;-�̨;����	8���u����'�&���d�%�	7+�HA��c�TLZ[�şP���T��(���(�G�j0���aܛd �5cDm��N2{f��ؒL�����;	��9�E�Bݎ�Z�'�(جAc��^S(<��BE�$���D��)!F�:5�]!EJ�#<�H���	F�'m��I �D�2&���s��;y6��'�a~�(��\���2�*�@7Ȁ)�`���>�q_��T��.t�V͂P�0pE ]sԨ�<U�]0�?���?�)���As$�O�ir\A�F��n�1@�u�g�B�8+��i����O�����S�t�)R�e�6��NN�L ��p�dZ;Y�d	d�:���Dc,d�s�>�'Q^�(�g6�`0$�S	m���̓}r����ʟ\��'����_<d��/�|rUS�!E*�!򤁚TFV]����&hN�9jd�۹=�ўD����ȫo�U �)����@�� �L��O��d��P�����O��$�O�����N���{X�h��eY�K|���@������D�]0��d暷8+:ˀ�3J��䕝F᰼s���7�Zܸ�EZ=}��i ���;Q�0����EkXhU���?ݻ�a��,�h�oO�KL&M�8tp��z֜��'��q����?)���p��AW	�1�kP�5l��A#+D��c&ײ8h�xB��1~��n�O��Dz�OJ�U��cЅ�$�B���%Ճ]���T(^)_�
M#UgD��8�Iԟ���6�u�'^3�ܥ�'�D� ��낭�-&<ɃBCA�:l�S�8��t��I  sÚ�:��(�F��&D0�P� ��+�ذ=fJٟ� h�#݊a{�	54m�LП�E{��Io6�p���{����L��MvPB��
u�Zu���_��i�THÑ&ʓS�V�'U�3�����$h>�A�ӫU����T"� K���O(����O����O��8���+/�!��d"Ҝ�i>�R"�̌<��Å�\�0ZD(�%L9�r���O�*XА͒=���V�g��x�g4p��	!ٌ@>�Ē���O��D(��
p��p�Հ0�d��vFΝk���0?�`FPD����A�	UD�R#�Ax��C-O�	�uE�vW� ���!S��q�Z�tQցIҟ���� �O@VY ��'�r�S�6>
!r	�K>԰�Ʈ 2���
��@���N�6�է��'�SK��ъ�#�R�H�	�8BN��I+ٺ�K�ˈ�4�r5*�O?�sv��3g��'�fպ1[�jy�$Kp��O.��=?%?m秀 r�FK�.F�ш�� l�)q"O�a;�Z�{���1�I��b��I��ȟܙ�I�l�^9 �ҍQ�,�Y0��O�D�OF�s���L!��d�O��d�O ���O&Hr2����\��+��:��bk�<����Q�
� ��P��8;���#V�O`���"B�u�tC%+Cx�+��=}p�A!�'wk2<� D۶F�� y���g�%?�#���@�!�ޫf��`Xu�J~�#���?Q���hO4��r���@ʇG����B�#�B�	2F�X!���<��ęG`]*)���d^p�����'h�?
Z�4@q����e`�9�܅stI�8bu������I����S̟��	�|��Ӡ#�X|I��1x6��:6�LWH%c��]�����t�'�&l���<e�<�qV+
�hV���0OB]�"�Y%�׋W�`��$�0�҉���F�J#
b,(�K�G�"F�B�t�'r�@����^Z�����^�� T��'-b0��Kf:��8c��n�~��(Ofo�ٟ�'��,SP��~�����J�R1N����5��� �Ҫ{����ޟ���(/9r�����m�ty�d��47؈
���p��g�L��|�u%KY�v�	��^-�Ta���D$�פD;K�]Q�o���<�)�n�s��A�)�'Z8q��ğ�|j��^�-���sU	��Y��kyr�'�Dl�#bb��s2�όORbl��0��	 2%J4jU��ʀ��d�T;SG���?)���?���L��AŗS�n�ڗ�)Zf	ZS�5O��=a��Wi�5��Ig艺�j�e��S�Z�%���~��MY�z s���"������x~򆧟���0}*���\�m5�z���s��X	Ș���??��>���[��i��]~�<��E� �(\����>	��O��}Γ:PŚ5$Hj�&�7I_�p��sV%�S���x�$V� ��5�SG T�Z'��#1��v��x�R��U/u�����D��*Ć8��Hv��>8r��)�i��P��I���,'�'(�7͐�-X�D�4cwϔ��&��E�I�8y"�'�"�$�*�� �c��-9�ً����O�������S��'��X�O,"fW�*Y��[���r�ȑ!br�#Y�y����?�ED�<)��ī�{,ر��;��0�k�?qQ���d�qo&?��y�f���~B/�V���6��܃H�?ɑE/�O�a��G�/`2h�6�"/30�V"Or��S��5#GPM����`#N���i}r�|r�'p��N=O�R�r���x��*�O��BPn��$�����1O�ip|��.�*?;��I�|��E�M<���)��u4�a�b�$C(1��S�!�Lb(�0"�&(�E3#��]�!򄊄df����S12��� Oż/�!�d\)K�N���DA&�( ��Ň!�D*'�,�Q*�:�F��!�6
!�d�43` X�P��W0�3f��!�(R��u���(BT&��u�X�=�!�=L�b��0yL���* �N�!��t6�[�m0oB�1`��5!�S;	HB�"���,
�CR�G!�I�rfp�Ui]�b��{@���!�䆘��m��T���h���72��O���^�27HY��^*}?ƑI�NC�e|ҵ�3��z�LT�Q�϶�Q��%Y�t���HF0���a���a��~�����^f��k��|�)'�R�rZ�P��+ƙ7�>I��D�G_ ����J̙iך��h�?��={��N�)��w"�,��Lr��꤃�R�n�:U�ߞ)�T���Ij�)+�r`��l5ze��釛X�i�ȓ]i@��"ؓq,�(/��) � D�8s��VB�|�;tlW�ˆ!��#D�� �t$��c�<�j`!��6D���O6N�&+BO�+|���!s�4D�P�
�;��!�!��=3�d��ԅ/D�xJ2�W��D��Y�8�� lŃ�y�m^�s�
�o�y_����¼�yRNG�l���D�E]gK�y�	�g�ll��B��8��\��y��F�N�StJ 	t�F�۷�y�)f����쑯}�xĘ6���y
� >�k��ˍf{�1Y.�$z1A"Oa��eP*)�>�`�MJ�g��`�"O$a��13�68���� O
츁"Oh���版�2���_*��U"O8h�Ԯ�(�x8��ԍd�1"Ot��E�P{I$\"�����"O���C��f$����!�R��"O�|�v�(�ABC��	�$*"O���2�̕|}�yPb�)7�0ՙ�"Oh|c����7HdJ֏�8V�D�0C"Ov}��C2S��X{�/Ծ+�$)"O��j���zb���s�1D4@�Xa"O0��垸�t`����#'d��u"OH�D$-����'�e#�7�,D��#S��Y�|� ���,c�H,Y��+D��1�+o
�pI$#_/##�xѕd<D�|J���&bɈAb�o\�5��D��;D�0F�&Kr5���Z�(֔I��7D��Is�S3m��Ih��Z��y��n)D�4I׌^�B�`b�$E]68��q�(D�8�ݗZv�����N* �j#D�d!1*�*^Fh��m�17�y�B>D��K�%�6���Q6�;V+����:D��#�-�7����p�[%}8�0A�%D���C�/���4��'d-x��!D�\�um�[u@ ru"V+(e�l��H?D����?f���4`_0&E.Փ�1D�P�b��i����(�1e�FPG 0D�����!z#��@#	�?�~�a�-#D� \��O�5ز�;��G< :C��E��E�+x��U!$�t�C�	�V�l�E�4Sގ)ۧAB�P��B�I�v\�a���$f�i�e�
=_�fC䉇C�XjBK�)�^ՊW�M�2C�Ɍ �jaf&p�Nu���؂bR�B䉻!O����t�v�RH�?~��C�I�qt< ���R�:�HÌ=A6�C�I�������
QT�
��#�VC�ɝ�褺��|��IT�H_�<C�	W�l�O��!�J`��ƌ�TC�I��6mJ�@88lSS� p�:C�	._�h�� �/M��y �k]�C�	;S��JW>2���J�JAFB䉬p��<�N,��s����B�9f��l.�9%�}pd�D�b�B�	�(d�����H+b�\Ԓ��׈c<�B��?K����!�A�`�J�h��:c�|B䉯S��{A��=O2L���"cM
B�	.���"���.w~ P��(L5�B�	(+��t����8p���`B��C䉌k8z��t$��l��ɚ�J�6B B�	�cM ���ʁ73�yB��N9�C�I��r��M%+q<�P�)B���C�#����ã[�$0P���,��B���
p��*M�6�M�♊�rB�	*.��XZ�2��<cB�s�PB�I�*�8 I�gE����i����XC�I�W*�����E��I��mO��lB�ɐf[��ö���/�
;��B�8NB�	&FXyтD�/�1�QS�S�xB�I�;<r&k�������lC$ �C�I�p/� �Ĭ�7P��)h���\=�B�IfH�H�u��q3�KW3*!�DҹW�I)C˫�<6�U�!�� SQ��&k�y�$_�H���!"O�r4�,S��a��"m5$� �"OnM��"�5�{�(&*��9c"O��y$�Ɛ��A`%�^�2�(E"O��"�S�7�.| �o:�"q"O���,R0i`�!�d�7��<��"O@U	J�3���j���!�z�2`"O���I�!d��X�C������"OmЁ�Ɏ�\ Ȁ�-��M��"OD)��b<
�h��AF�.�xC�"O�93��ts�jqe9\�~���"O�=I`)��b�<2�c١��H�"O�9��N�H�t9�C�s�,@"O�LY4b'q8��-�"T;@  �"O
�@�K�*�\4�U&;C>���"O
 QU�=	�q�4�w[�.)�"O�\:VLQ�t�ĀP�Vw�I�"OxqVb�R�)��^�H�� ��"O�d�q��:[|����
�x��"O^d��FV5�j�$��h��:�"Ox��Ҫ�*Cy�i���)5jޠ�"O��E�`W���RE�`2���"O*�'�Y`�,��6E],�p;�"Ov �2�>e:>���%�~v���"O�H􁘟~i1ˠÃ����"O�U��f��d�\SG)��@��(��"O0�xW��o�FH��%��0��Y`"O��[b�Z2�|�y�O+��b"O�K榈�u*�!6O��g"O~��C�K*ƔH��D?�Z��R"O���Fכ0[bq���d�Tx1"O�!q�O-'bp����L��$"Oh ��NS.G�|�� gRC�sa"O� Q#�ӃYcZ1�e���|9�S"O�8q&�J$��,��C�Z�*Ń�"OP�#���  e�@j#i
/7���H�"O�9�'��F]��6�	a�f,)v"O`1sU��'X�~ApB��&jzj4�F"Oh ��oƻ)J�zw��8E�cD"ONd�g�S�y�8}J�Ò+r��8s�"O0ň�B��\���%x4r �%"O ���hG�L�D� ��+%n�� "O�a��ȇ�(|xr�\h�9*u"OP�b�#Ϻi���©�
j�1*ORԡ�.�|������y�����'p�$Y�/[�"1NM3J�rR|�P�'+��z���@<�"bK�`NZ�'����疙QbiT@���'o|Z4� �;�=��x��j�"O@k�#ƹuhܜ�Ca��~3"O������T�`g�78�&�k"O��;� �($HѶ��E��E�@"O�9Te�Na�e�F쇸 �h5c�"O���6�B	���ZW�J�0*�)�"Ol������T�f��N4Dm"O,�!���?b�Ehef��1�1j�"O�-�g�
4d��Q�B�$n�(�"O�y� 	�%V��(���0.�Y�"O.}���0V�-�T��#bX�"Oh�A���87��lQ���(r�0�"O:\x��	)��rR˄�|
�@4"O<�KWH�M��(s�6\gvh�"OȰ��L��0)���"Pd��c"O�����BH���3�
N_�� -D�� f�Zv�u�ڝ����K��0��"OZa��͌��<�:7o��|��I�"O��8�$Bj1�l�EP�b�d���"O>u��oɋxb�@��ҔZ��dB�"O��wI�
0�� +���=j�"O���gT?p �PQs�.*�p�"Oղ��HAt�V�F�[�$x�&"O�qa��g%��P��šp禌��"O�L�tEٮBl�\�׋Z�R��+ "Ox�����4wTdX3J����(�"O��kg+���H%��ꎲNT�{b"O��:7팴,�� �eK�!Q��I�"Odh �Ds��M+��Hb"O|��kJ�7���ܦS�`x��"O |f�.9��pVcT�i��;�"O��@�kL:0���'c@�g"O"U q#�,%x �r�P�w�`�ґ"O꡻w�ӆG��q�(Қd��M{"OČ�!�{�d��6c����?;�!�ĉ�Lf`X�J�p���a��!�q̆%p�I��?���"� [#t�!�Ă�`��e�ҟ�.l��@-mx!�dWUp٪������@?!�$�$k�d���EJ����
�u'!�D��da�M�&R$P����M!�DN�N�i���@C� ��!���!���fG6}�D�K4�Ȋ��~Ih�'��{���P�l2��Qc|�!�'��qhӁ:}ȉ!1�7;	��'�$�ʤʞ�h��x��M!Dʦ�*�'M\����v)���%E�%�	�'��:���Q����H$4;�$��'����U
6a�\&1��ɩ�'��)#�:q��)fQ�,�x��'�n}�@Y#��ʦ���P,a��'^�y[R,�����-@T��'ԚĀG	�����@� �yS�'PF;��@�嚰�Anنv��H
�'�TH�����:l��S��]"[��و	�':�4	'�[�:�j`+&m_1b9��P	�'��5�؈itY�vJ�%Cà}Y�"OF�ct"�uFZQ�V��3s��@�"O��t�N,E��rS�E+[�Y�"O�P��	w�i�0�Q����H�"O`E�2�^%K� ��zH�"O��@0�-�ТSe�#�^�#7"O�a�E�)F~�0�7�G����ʗ"O��P1k�
'j6lY��ǜ0�� ��"O����ҼZ�t�"��>F&n���"O��jՌM���Q ��l�l�"O^ps$o�3)�JBh߸O��-1�"Ox@i�NH�Q4]�r�	-d����"O@�8��+,�hQ�!�ZlP�  "O�=��	P&hr*T� B�']�Tu��"O��Ce��*at��r�׊�V�Q�"Oj=�Ќ��a�����	��^�r�"O���G^�
G1���_B��Zv��?<�-:b�H��:�9b�F�;H>��� cVH�7@� ���)ֆ�o�<9uAލ\�T$���=���F��i�<qPN�:?� ,Q��fV	��Ug�<��n�ssJ)��i9��(ϕ{�<R�^��HlZA`�9c@=� �b�<�͞�|s����RU�m���b�<�a.�&ʔ0p�I�C��k���S�<� ށ��*�=K�N@`�C���M
b"O,�t�S�s��|2��A�,�k�"O�(dł_��x;G'MTf��"OJ���6^��ؘE���9}�Q�"O��al�)4�����kFl��D"O X��O([���A�rڂ@�s"O0y�*��w)�M����xȸ!��"Ot0ر�F�"���
��U����"O6�h��^�Y-z#�ED���0�"O�5�f���?{x:U�O-��u"O�鳫C��4���6W,δx5"OZ�sm	E{�KA	ɅT*��" "Oȵ��K�W�(�	2(ZU�"O�4²Ƒ�."�C�	Z7鴴[V"O��k���V�$�G-%�z�s"O�	��D@C����q�Υ[��0g"O�$K�K/"pS����T�C"OZ5#��ܲ$�:mҷ�F�"��=:D"O(Ȣ3�Ȗ;tԈ��N߱}� �Ӵ"O����B4a������͚A���	�"O�@y�mT�b,����Oz$Z�"O��RA�	� Q���M	�Zh���f"OVY(`G
S:<���%ǱjV���3"O����F�Ĕx$fK�_����F"O���$�>pZ
E��T��t��"Oft��CΞ-,]�1��:!C*���"O`Lq���;G2�2�iH1�D��"O�a�p���^5�{�c�YbN�y�"O� *���B墍;X:H�"O)Iu�M�Ԧ b2N��q"O� j"/Ev�1p��9=�`$�g"O��bf�F�"0{���	k��Y"O����)6sȱtNWG��`j7"O�\�dD8+�4��ˋ�#*,T��"OP��F�K�.M�!	@,6���W"Ox�tB�xS�I�g��?bnH��3"OlXڶ�ѐgŪt�%�̌��mS�"O��2�,��}����JZ)�t"O�@� �x/�1��Q�&��#�B�	�V	�g�A[����h׉/�B䉳L@:�g	�Uq2�S#E;6B�	���)���"�p�[�ᕌ$B�ɰO�Z5�����<��2��p0b�-D�xh�Krϒ�Cv��E��M,D�8�:r�LEfF�l��:�7D����fF�~�أŊ�4&|�K4�3D�D����UӒM{UjAt����&D�;�W���I�O:Xͱ��&D�0+b���� �f�Tی��J%D��ɃE��)!�q���G�[n��*#D����8&�� ���mD%pD%D��C��-(aĸ�QaǄP�@��j>D�� /�#W��}��H�N�<]���<D��+g`�!�L�J��/Q�	��6D���V�@?5 ���+B>r�uP�N D��Y6�>05� ��!���Uo8D�xJ�L��mDj�td��%OdH�D<D�삁��>�j��ړz��(�/9D�LA�v.�z���<+���:��'D�����Λkid��q�у5�0u���7D��œ"jD)�)�91��X�(D�Ȱ�oS o�
�ˀOZ$3�Y
`#(D���f#HG�e��I�+�֩��7D�h0�N�B�q[0�	�6Ð�au�8D�� �Qd��c�C)��^�	�"O",����PJS.L>V�b�"O��b�/�n���:8���c "O�p9b2��ȇ.��T_4}�6"O�%�C��`�����:T�)�U"O,a�RA?)��`��#ٜ��"O��BN��t�>�1�%�0���"O�\��&|<ā���6y&�"O�2`S��4c@.S xr�X"O�ՈQ���0EDA�`��"O
,AA�����;�#�I�D��"O��+�8P��<�A�<e��m��"O0E��΍A�%���?KK����"O�й�*]�1�$�+ d��Ht�[�"O�U�KǽG��\(��^��9p�"O�i��ўElݳ��_�<��\��"O�jg��3P�\0ti�1��"O|����	3$T:@�AR�b!"O[!�l�f���
l��M�"O*4� +O��ʕʊ�
.>��"O6u�=6B���޹c��`"O��	��G�g�,���$� ��R"O���d�?��hB�f>�ͩ1"Od0��E6,Nx�tb�b)h��"ORm�R��#2`���@98!�H"ON�'N��0f��H ]�Ǩ"D��xG��@��P �m_�u7�q��'���*4*Q��ÉPf��Ta�'����)׮&��a�c���c�l���Bv�Ը�F�~��eE^�����j6Ƞ
A�I�=�� '��ʙ��S��A��ȚA�`�Ѐ��"G}d%�ȓ~���R��=n�%�
3�Ą��h��6��`z����)���̈́ȓ"�`Y�f��3�!T"A'��ĄȓQ<U�@�	�>�Pm�2��-TXF�ȓ#��G%�tt٩!�3#x��ȓ=��m0�KF� W�y�C�RdPp���t�#��ʙ?�ָz�A5��Ņ����D�M�hBD�
P��]���M�8�����G��fa�Wm݄�c��*�ˆ(x��$��@�2�!�ȓRC����L�
��A�&S�]�ȓ)���ގ$�VS�	^� ���
!�����qw�I*�Ý�M����ȓ^Y��z�Β�lx9�c�<elĆ�N��y$�ԃRg<E�e_�>u�i�ȓQ����@_�[���D�FbC>�ȓF	� �H�n!P��H ��]��T@u�P��#oD	�`,�z���ȓ6��m��ͦ~��d!�E��W�⩄ȓW9�XPf.���U��ʃ0���ȓ9��<���t
�F@��]��nP�Q�S�X��$X�SF����ȓ�ș��ԯyj���H�
1i��N�"͓��Xjl�p�$��;&��Q�ȓ3� p�;�Nc�hWX���v���e�7)�0���/M�݆ȓp�̴!��N9p���P�R}��6I�iB�B^�9��Ÿ5��
6�����	<,�PA��7z�d�����T@$Y��}���#�;f�Hȵ-�%]b��!>^`a�gĒ)��`��K�#�z���h�b$� l�j ��镺,t^���S�? � �� s��i��g[�_�E)0"O��2�o�+��Xp�ِAz��"O�܁��?<�X���W�c]����"O���dA	W��a���S�j���"O\�@g��-d_�-�de�G5|���"O��З�\o�U*�ŏ�S�ܴz�"O�x�S�	�$	.q����/$"�
5"Oܼ� 	WCj`
 K0 �w"O04��	K�N�0��˚f4+"O���&�H�w��
�Q@�"O4�r�8%+|�4�G�Xfᓑ"Op`���� �T����="bc"Ot2A [
��$YsT)B�q�"O���T��(m�
G�=S؜9�"O���Ą�B���S�#mjj "O�@ �M\�c�����Vl�A�0"O�a�Bf�AK<]B"�:7\4L8w"O�(ĖE<��Sҫ��8�.���"O�Ͳ�,�"��4�v��;���"O���q�
�r#i�Uk�s�T铦"O�1�h�J^���
\�\>pe�D"O�4��L_/���MN�t�u"O ��"�	^����X�M�(��"O�-�&�������n>ـT��"OVeJ�%��n�Xd��lU�H"$ pA"O|�{5�G�M��Ac���fE�a"O�=���$�2��D��AD@�"O���ț $��Q'@��^ ���"O�����*���2dݖ"L
��"O&��%��*h���ćWFbm�4"O��� O/>�y%�ɟ$��*�"O�Q8���3B�������J��b"O֧�i@0t[�'@,ҰI�"O�qX�*Xrv���W�+'9|]�a"Op}90a5C֚�rŃӬ!v��#"O�}�"�ώ�(8Z�B��1r�X�V"Ot�#��&��8�O�a{�U� "O �[1O+]LX�ȉ�/{!��"O�\���D����O�(,z\@y�"O�X�c� �^A��Cyb�C"O(@�i�D�����#�-kܼ��"O������W�x��ɛqeyf"O>���G�<aMf�42���"OV1Y��؀T��� D�A�$a�"O���Ŧ�v,�8�ce���A"O
�sg����a��IS�0(��"O���#��?S���)2s��KS"O��k��S�IUs�hʨU�d-��"Oy饍U;y����U�ӕp��|��"O&1�fe@�8?LY�%!,cSv]:�"Od Jt�Y�O0�k��Ǩ=jޕ��"OJ�!G,Z�SX�
2ȗ�1��"Ob`���y���"��*��:�"O*����������هD���"O괻q�L�Q�M!�Ѥu�L�"O\��W�6�༡�eZ6���8"O��3�͐�Yo^�c �,ծ��%"O�M�D��w��9�4�,+�9ؕ"Oj��ac��MA`Hu#HY���"O���2��;��ل�a�y��"O�y��>F�zE��'�%CFz��"�Ě1}`mW��p�p1��/����'�Z|C"¸6TV����.�(��',zmx�	��Si|m�󄚏x28tR�'�+G�i�y�w%3��Y�8D�� �\��h�3��eFḚhӢ�i!"O�q�B�O�7��� ��1���0"O�uqq�Js���T��Eł�R"O�A����rOZl8GJ�)�jp�"O�yѶgP�S4���
ɝI�|(R1"O��Q�L -��q+%kQ<;/��7"OF!3�!�:��2j�:�C�"O u�pj\�Ct�k�J�8]�4�"O��� �D.E;F=i"L/;>�X��"OZ�"��J]�2��e��"OV�*A+^�_p:��ǩD!$�m)�"O��a��� /�Qza�ߕ
�8�̓rРh�p�K�Wt遵��Nz�͆�U�$�hT�� Ia.�I ��ɆȓetX)P�Ғwը��WF�Z����ȓyqԠzu� �<^���C� >Z��ȓr��T��'��+�*Mq�̕A$��ȓ*o�����r&|�`MD�8~�0��dy0���@�S݂9CF'�A���ȓ�
ak�kߤ�ȱ��H��Gu �ȓ7䈽jT�ف9Ł��-7��t�ȓ`�.d���^�rz��Jt�][�l���� ��#ت�5�*tִ���(���"�#)������Ȟ����:}��6O�)t0��A,N�u�Յ�Z�*SwY�&��Əǲtj �ȓ7�ԡQ'	�B�pP1$�&z����w�z��IբP�be g(�mtlC�ɂ]�.Q��N�>K�����7 ��B��,e=�u�R�]�:�й� �"TRvC�ɩ&�P��B�rEj��B	1�pC�I�Bi ���T���V�8C�w�bpt��e�BU�8IG�C�I�5� ;E�ь:��mRDO��DmC�I3:���x��͒�va��,�/n�0B�ɋa��y'��&� �i3�
�9c�C�IN�tUk��>����qǺ��B�	���� Τ��Y�tm)�<B�I�eX�Aj�@�)�k�-#�0B�I8>��T���=��J�m^� �jC�Xlj+	�6��Q,G�DC�@��1�OY9@ђ��j�r�C�I�`�P�DgQ�O���pG"�1��B�I�&��`��aL�Q���B��;&�B�IJ;с�@}~�)�(���B�I(]9���č���DG�]��B�x<v4x����jҊ��Ƣܵc�LC䉗X�R�"O?�L1X�왚�.C�	 H�q��&� �hSL�:^C� `�&a�% ¼K�P��A�FB�+�pzfC�g��$���T!0B䉯lM���G*�g�VDJ:��C�ɒ3����F-X�k��#�iS��G"Of�S��_]G`@�{&8�
"OZ C�"�$[�����LT#[��"O������3S�02�i��5-�e"O�y��l!9b�$�W��<$=��"O�x���Ģ)1h�a�N�~�B"O(mȷ��L0 @��F�0c��tK#"O�1���48h��3�K� �i�A"OPL�%��L쩐J���H��"O �+Q����z��9�(p5"Ox�a�]��U�w�ŷm�ŋ�"O�DIu-V�&Mj�`�%%���)"O� @���D�T�X�sM��h�j	(T"O`��f���8�M �h�&L��"Oց0��S�kƭ�񋚺'�b0Z6"O�����
a  �M��$��"O� cI����i�ҎD,q�F��"OL ��e>C�D�{S ��%�%"O�4 �,¹~w��@v�͜tL͘S"Ob�)�Z�(B&8ŝ�:0 "O���KT��Qk���+�� �"O�E���h����O!T��M�0"O�]{'%C�w�R�T+g�lMS�"O��H&A��8Iؒ�U�b���E"OthB�D�+2��@��&R�a��F"Ox� T�k~ܣ��m�R�B�"O�x3$�<'�h�Zsŋh^��"O���%��)<����'*g�y��"O`���R�c<��˷�XZ��m;"O��c6�@?J���4kKz�{ "O�� U�]�5�<��a�;Ht�s�"O����>-qx� Ǎ]��8�v"O�r�o�;wIN��f���6"O���D�D3 �܂#�T>7�l�ٷ"Oq����7�� �֬�(2�J���"OrX�I5�`ڔ!	��X�"O���2AV�};�=qc'��
H<�zu"O��0'�ح��l��Y�DL���"O.	92dۡ���x�$��{�]p�"OXmp��˚=�V�sBM�gJ�ذ"OV0�c)�?o؍�U�qd>�*"O�Z#��+��H���U5%F �v"O���j�4��͚rl�UL `�r"O�1�$h�J�N00�i�0BXT�(V"O@d�4hT<r��`	Th�*@�Q�"O�X�qa�,޺�D�"��R�"O��Q�d�u����0�N�p7"O  �&��x����3��
X�M)�"O`��&�۰|
և��Pe <Ra"O��;G�ь,�[Ռ�5��Q�"OdUc��^�.�:F��>ݚ$�c"OH6��b�����,�X���"O �{c(H����!N��$��x�u"O������vP�qq4�Sk���#�"O��@!���6V(q20�Z%P��9"O�BwC�Zafٙ�p�X�"OJ�J  i+�8a�q� :U �*�"O����j�y� �qOTn�]"O@h®�4�!-�f���/�9S�!�d�i�[�0�L��NHw�!��92�3PBL�
E`U[��F#9�!�_ Ft�wB�3{�|h@��`|BO|�g��"� ����-��+�"O���%�i�tP�wo
�z�0��"O:���i��@��8n��L���!"O�$ըR�7+����Ύ�1�!���X3F��%�!>����)a!�Ȓq�vH���Қ}��-�Wb�.�!�ğ2P���w�N�x̺�e�!���_��$3�+��S�)3S��2!�� 7Z�Q��M'W�v�`�_�2"!�V:2/~�A�&ƛ6�ti��O!�?dxb��H2/�hq���I��!�dN�X�F��V���\�P�O�Z�!�����37ܺ����!-r!�ӢA��iq�H*�6�8&F�]!�� �i����/^���êFhS�ȓ"O�1��8&�}��n<s��0�"O]K���Z~|ipm
5MN~�9"O��'΂�^3�qط��)[dY��"O��`WL͌'�� ���t(�(3�"O�� ,M�|���cɇ��6"O����?Q� ���.s��S�"OBs���p�e�Vkr�DX�f"O^��w��#*�8q�B�P̠�Sb"ON�����,���Bt��#��-�y"+[,H���ȱ$[�G���`/K�yҩ<O׺lZ󋉫h��u#����y��S�_��xjtM8� ����F/�yb'�4z������#(�,5���P��yR,	j
�%a�"%$A\��� ��yb���oi�Z�ˆ�G�Zݠ��yꇱ@bZY2�#�3]t� �Z�yB뛴(Y>i���:2E6���.��y*�b&��F�TKlI�n���y"�ċJ[&A�d@A�x���	�	ܟ�yr�,7�v�
#gƟo�lRvFF��y�mכO�x0�3'I�1cB!�E�F#�y�j������M"r���<�y�i�.|+#A�V�m䊅`�,��yB%��>�4p�,՝c�Uɂ��3�y"/�	Gh����4�#�K���y"�%��|)�vJ���+^#�yB��Y~B(;�".=7�4���3�y2�ߐD`���H�9�*�-��y"�ÿf��E�+h>��"#!� �yB�P6i̺Ӄh�<W�p� ���yb!Sh�5�fF�0K܀�s�@���yrNU�d0�erb�=q�E�A␅�y���Y�PÔ�X!:��y��j��y�G(4{n��Do�#���A�M
��yBa��8<�*%A�������yb�HYn��섃bq����
��y"���K���&Y*�Y��lȅ�y��ڋ;�*��EK�O>���C��y$����{G��I 6������yR���~!!A@
?��8����yr"�'VX�h��2` X�G���y�!�#E ��ޫ9	q�фN�yBE�0ER� E-�,���i-�y�_9b�����7�B�(a��$�y�=����\�l�f=���2�y""[7ip0c��a� �ё�F�yrO��'4�-�ͅ3Q�8Xr��T��yr��	��&E��R[*3��@>�y��ߵ8�ڜ�S��3Q��x�A�8�y"�]�
#��f%�-y��m���y�Õ��"S�� �Ta�鍕�y��ҌVC����'�<�8��e��yf�LH�X*'bO@/�9J�-\��y2
�e�.��@���k�zrBƏ�y����.����֯0`����yBAVQ@<��[�Z���֥��y�	g1�Dr�� gY���(�8�y��:]��lX'�M�b���{���3�yRe�eޮTrDU'�b	������yr��_cȐK�E 
YP��ץ��y�/\4������~΢������yb�D�j:��7�Ίm6԰`F���yf#f ��ږL_��䫤�D�y
� �1 �l�p�'ʧ#4$q�"O���cӃ�6�����)�4��"Opp�Uς�O�FDS�яO�(�"O�D��.v$�UK�� (0�"Tyb"OJ�`�W�$��н�v�"Oa����3]�1rV��$�V��"O�(s�ǋ9hH��	8x,�<�"O�(��V�L�v���2b�E)�"Oj=@�H@�D>�x�� �J��xb"O�\��I��-/j���*ӕCJ�Ru"O`PiUZj�	 ��-<�l�0"O��a��K���c"��Z���f"O`�3���#1��C�͍�x�"T"O�Ac��+�4L��N���UR�"OD�3jWqy
]0 RS�Fqm&D��e�U�a�(���j�~q��8D�4��ۛS��x,M�,p�q�))D�+��ȘhR�����8s�2Mҳ�)D�h��eW:9�^hz1�N;�*I�F-D���R��W�h����%Mܰ��#�*D���祆����RWd�_d�!��#D��J�n��&0�t��/%�v�AI/D�<��� W!~�6(̓I�����,D� h���f���R��"Z��,3І)D��yf�\.*t������	�*drs#*D���E�#�*eht�Q20$(c'D���&D@İ(q&δ��05*O�a+wK�.2ذ�0�/	:�x�@"O��c��ĊbE^tp$lF�9�t04"O�0�Ağ�6�6Y�ӿ\��d"O��s�o�/2�<���#��B��4�!���s[�X���ݐkW\4pi�3�!�$��[r~EbG۳MQ�9*W.��%m!�dōp�@��y=�p�P��	!�$�����'�
6����>_!���q��F �$��B4�!򄖽X�$,��W�<�����*�y�!�$M0����Ŧ/��(JQ(Y��!��
�f��OӐ0vJA�A"G�H!��G�;����$�"Xb��bW�6!�Z3z��*��!1��1"Z�zD!�Dك��R����E> l �����!�$ )�@���nwl=�)\��!�$�T�उwɗ#>.��Eϔya!�$�5|Q�0�$s,JےZ�=c!�Ğ8�Z$�V�۸#P|��֘R!�d̿8ϐH�B'ŝyz�H�q2!�$ۢr��c�,����M��!�Q�DĤ�j�-�l�j���J�@�!�_&%�-����g�0)r��<9!�$ߑI�ik�H}��Yj�I�!� W���sEĆ�B������("!��> ݻ�B֫O����'K6JF!�ą�H�D��J3a��1Ȳ�K;p6!�DX��������e��Ǔ� !��-���ڒG�ֱAf�Z9i!򤊃�t�0��LD��|sC�&M�!��)7���ej�i�B��p�O�Py��w�T��# 17zD�P��Y��y���^Ol]��nF�#2�TҔ��y��@�fF�0@���lv��S�D[��y��F�,��x��G��K���P�B��'�>maTR�V�(B���3��B�	�`��Ŋ6� �SN65bP.�,
�4C�)�  ����.:�Z�& g�"���"O�98b�LXD\�Ԣ��B�@��"O���sÁ1-�Tx��L<ai���"O$�Ig�G2�����'p,b�"Or���"a
$r`@�p(�;�"O�B����p�K��&4C$���"OL8H�]%1��	���7)$4l)�"O�h�6j�(����(��&��V"O^����=��4�bgK�"O��6O�7U�1Xc$I%f��$ �"O<X�+��Ŝ�	SJѫ1�b|�"Oܽ�e��/4�H �9N���q"Od4
s �g�Tz�HO�	jl��"OlH�P��QZ��I��U2�����"O�C�y�J���K�ka��)�"OnRC'�0���z6 ��uN d;�"O@Ek�ʏV��=ځ΀#�%%�ybi
�)�F(����^� A���y�V	[�Dx&IA�X�0�Kaܑ�y«�	��	yc͹O�1�P��yrmM���1He-�p���2'��y�m&R�|�h��ATʍ�k�y�
T�e�P����Q������yr
� �X<�lF$�����F?�y2��g���!O�vV|�ɢ���y�8Y��X`��Zm�hP����y��6.^����@;L\�����y"�N�[D8������J�n!�"����y҄A�Z >��bDo��r���y�b���b���)^�:X��#�)ح�yb�Mv��aW;+��Eq���y!�1�H���a��V��C$��y�.��i;����O
%��tRCV��yB�\�2{v�vh��lV�+C���y2#�@�=��΀bAD(D�"�y���!*�xP�s��8`�fa�s�
��y���	���[�ݴ]B-y�ŝ��ydE<#�8!NWjD��u��'�yri�	Y��S%+�0d��)i�D5�yb���(`	��d���S ��y��K�BPȌ��F��f�(�!��ޤ�y�W�1f��KF�F����"«�y�O�f�������dy8��H��y�
ؿ RH�×n�Z�n<*�ˊ"�y�E�+��h"��{�61�#+���y"IɇW���z��z��ܳ6b-�y�
��mav�A"n�>�8&�	�yG�#���X���^����E����y�&	5<M kr��Tr�]p���y�#ڽ]���eo��yׇ�\�<��oL���U����7[&D�e��]�<q���X5�E:�"�y�>P��f�d�<A�e	7b���E F	*�(�C��\�<I%�H�
t:H��F��+���� �Q�<��kڞ3��u C�5�ŒTLJ�<�gS�JSB�Х0��
�B�<���Ճ7����m�>;�2��P.�{�<Q�"@3QX!�����)՞�q�C�p�<�֦Տ�ؔ���	�zB1�5Sk�<��d׊e�6\�bM�oc���Uf�<i��L-����t$�n�\EyVF�_�<�wa;|{���P.J��Q��UX�<Q���ݪt��/�K ��s1+J�<QOQ"}���S#U\��D'I�<� J�
!��)���sGC�$M�ذ3T"OR����)PI�ai��D#C�F���"O��1m�7t�01;f�Qը� �"O� r�d��0�c�CJ��r���"O���A��-��jvd�H����"OF����&Y[�u�e�O�s�*��r"O��{���Y~Et�N����"Obq��ĔnZ�[�ϑ00:E��"O�����C�~�P<���H �$��"O^ؚ1ϝ3U,����{ bHf"O�⑆�	����c��B�ؚD6!��Y�on Ad�\9�����#�6�!� �/Ծ����<;J����[OL!�䝍(!���	C�t�"�H�\G�!��y��\�T&̮0f�pʐr�!�d�($ZAH YS��(	��e}!�ĉ�"~�xPL��&�ɰ�ӟ	�!�&7�6�!2���D�z�tNR�$�!��ԨH��E:�N�7{d��,��!�D�g�ĵn�%a�����	�!�! �V- ��(��}��͕�!�D��u��Ѐ5��b��m8���!�ė1Z�b% CY0���@���:s!���B�b�2��z�:T��v�!�� vz(r��mv���DKp!�VY���X� �9)�)A4�H�K`!�$��|�`��EJ���$�!�I,%L!�D�Hξ '�T�D�V���C%!�$�|#ЄSg�̾ay�q���'5!�� <9%���`.9>\��G�Ѡ"!��(q/2�)򎅘vP���s� 
!�ǈ:*����D�4��)����!��Sߺ�YU��D�P��wE��P�!�$�����Kcc���,SV�ar!�$	�}��lXD$Ɵ|�6(d�
2X!��צ$.�YSp`�9S�ک[aϑ�}T!�䙺iWd����E�� S1E٬S!�S&J���&	�MrP ��e��"O�a��L1=���GF��(;�`��*O�9��MQ�
Oj�r&AMw�h8�'B�9P୘�P���� ?Eb���'���r��̧m��d�)I�7��0�'���I��
�tkpT�1�4-�Ό:�'��а#&N��ٛ�N��8�'�0��ԮN�MWP(r��О����'פ�H�\�<��r� ].-�
�'�D�XwC K���!�᜴��X
�'jZ4�1� ��aQN���>��	�'B��r�mP4c6�aeBù(e�'*�P�U����ǞI���9�'�x��e��'MҾ����<ȅi
�'a����ϛ�` ����)/\��'�F�����'�`xC��Z ,���'��X Ś�6��p���C'Rq*�'��L�w��,`��.5��̚�'m��Г�#^�� �.�R��	�'����+Ē]3�#�c8�X�0�'˨���Å�R@�B�:��p��q�<1E
$�8�(ЩU�z�![���q�<q��
n0���aY#`ܪQV�<���G=+j�1�) gj2��rj�T�<�V��?��A��Sg�y�]N�<iA��>"������N�p�)G�<q6�1Q`��`�J��҄H�W�<� p��t"�'R����C|x��d"O&D��HW�}��!��ms*��T"O��ط���J��R�o4vgXc�"O"-&e���M�@�6�lZW"O�%�A@���k1�� /�=�D�I��؃i��*�6�	�:e$��M�U�>݀��(C�qOl�$�ho2)�#I�|h� s�N�'6����O�����w'��r��k�D�����&z6E�hȻ*���p4FB�U"�}Ҥ@����=p�Ǝ#o�[V�X�E�����3���{a���O8��7\�Fde�k��?����������w�ڟ"~��k�<#펟>z8�醈rX���$�٦e�	���ӰO*�[�g�ds:$a�&��4�W
U��M{���?y)��T
d�O��DoӒ 3G$�4�,�`�l�2.I�R%�!@)O;@-���ݱ �z�J�ҟ˧��^c]�A�?Nn�}caǔ8��޴"Q������"]M4HsacɚH�\�y�D�G�<�|�1U`�0�'eT,#��4 � 5�8)o�g����O���?AE��&~�	t�S25�F 1��  �\��㟔����܁A�B�X��p�,%V"��&�b̓)�6�'2�7M�!l|��qɛ���<�N�fS�|Q����MS˓`��A��O&[J�� �1r'^`�u�R�3�n]���_�
�ґ�%�H�`���[~�'���IƇD�lu�*����}����`���V�8�3K4�ٶlE��i�J�[�� }Zȵ��K�2Huc��J�9�fh��O�I���'S�|��'Zb^���4M�(m*D��"�!C�a������L�Mɇj�3��`Y��]�t*rY�i��'O������'5�S+m��l�nߺt3$�C���`Ęa��L�'����	��<�	�4�ԟ����O��	��ݲ��� ��|a���%�١j���rfCM�"��`F_�L�ۍ���,�\A&Ć>^�*,��*��r�x�M:��}pF��*��,Qc�%���9`�	�2P��a�T�'�D�P�Z��D�^'WY2��A@���M����D��˓����|�ɭA�Vlj�O�Q��\����}�<�!%Ǎ?!�){���$I�8e�ck�%P�x�v�$�O̰mځ[��`޴�?a���?�]f&��
��A��Xy�)� 嬡z� �D�O�d��pIB)�dퟻ[t�=[�#�xT�Xs�O'���!���XL�� �H� }��k���+�p!�N����wB%r�T�: �<c����9
�F�2�՞zY�����I�2�d�OB�$>9l��)��-	�뉫�
��q)J�QR2����������\�,�Z\ ���-�D��1�"Ọ=�|�°iy�,r�L����$ez�GŻ!WV��>�=��O��$�|6�� �?)��M3�SfGr� ��w�| B�P+ntV��&��_ Д�Ĥͪ$���ן˧�b]cLf Z���92�,tB�����F݊۴oc�D��}��y��ڠf~A�M�Kd���|��[�"���2
`�B�� π�m$Q�����O��i�R�sӠI�P#U�#+��ag�"r�|�S%�O���<�O>���Ԉ�
S��a���;+�
^A����Q��B�4�?q��i��Sͺ��ꏇ29
-IR.SX����$H��`'��퉍wBf p   ��   �  <  |  s  �)  5  H@  K  �V  �a  Dm  =v  �}  `�  ��  �  5�  y�  ��  �  H�  ��  ��  P�  ��  '�  ��  �  Z�  ��  ��  ��  R�  � � � A �% - �3 $: g@ uD  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�Y�G{���˾R5$�Qb+�jBƅ�7��Oi!���l8��Ӄ]*W>�\����]O!�ė��ތ F�8#"J��7Lb!���P~��#���(%l�(.ԜoI!�d�0c>��=`�r$,�
�!��LP!���6HٮsX~��!ݺ�!�Ĕ�m��G꟯i�̥sQ �W�!򤃛]Q���D�o��Z`A03�!��R�6j�l��B�^ ū@��;Ol!�P9��$`b��e&Ī���c@!򄊡jX�QTυ#i��A(PhˢF"!�D/2��`pB�]�6�`�6��9!�dEE����BݙB~�tK�`I�W�!�DV�=�i�H�!(^n8�䏔$g�!�$��mMX���9OT���n��O�!���-
l��WoР>J���NE�ni!��K�4�VYP�ɑ����+L�xT!�$�4<{��J��! �PhX6*ʨI�!�Ff^��PR*C�lʹ����F!�ͪ&�����'�4j�\���(�8\!��/�:��������bN	i!�$�<PⱫ��53���{J!��@�S�vL���?ʀ4sW��*t!�DT��`Iȧf yƬ`�c�]�#�!�D�p�,l G�.x��ᲆ�T<@Q!�@7_�����=�"|p0��-N!�"F^�cbI��i��,�g�:'�!�0�@1g�żm]�,�Ҭ�
3�!�d����(�qKrأR+�<q�!�ںO`�i�눏`�p�5mܒ<�!�d?B�>�1f��~�>�#���0b)!�$C6h���@焐K�и��)4!�� 4IAI�R@`�g� @K�C'"O�ِ��3|�V9Y%hS?<v��"O�y���<9�t��'��X=�"O�a��Q�/k ����$�Lu��"O08DF��D��6.M02㼠���5D��")U+e$l�ȶcX�6���Hu*8D�T�N�,N�n��4h>~��ǈ+D��@� Aƒ���eT�VD4��%D���q'�
1��Z&�Q�9h� 6D� ��a��1k��T% ���J)D��(�f�4��US L��1�z]���4D�p�3ϐ�ѡ��R/BI���&2D��I��.��s���p�� -Y����@�Ta��ցE��1 �oÓ�y��SZh&/\�SIRݲ2��y���(@��Sʀ�9̸3�j#�yB�ZM�z��?~�t�>�y�NÙ[8,�kWG!hQ�\�C��+�y��/����C�úkl�Y�-�yҎE G���롃�f�P}��eɱ�yBbӣ6OI��G�s�@�a�NI�y���(�=�"#�1lu�l�7' �y���8l<v1C�G͌eI^yD犠�yHг w�Ժ�=S]��������y�c�'�8*QE�K߾ț ���y�]*�������9,�ٸ o�#�y��M�j��D�2|¤{�G��y"#̽���h�A�a�Z��1Ů�y�)�s�0	���\Z�����yr�	z�H���+1��	Pj�3�y��XZXt�-�%`��ʤ`%�yR�IJ�P�����XWI /�y2���U?E���Ԍ|�j�!���y�c'�V��p�P��Bh7�J�y�:v% �𥑮r?l�i��y���T[�)Qg��}�`P1���%�yR���.���8�C["#�v��AOV��yBn�b=�A�X<� ����M�y�eD�_"J���t2a�5�̂�y�*��X`Ht���:�xED���y���1�J�Bc�"��,zu"OH5�5����\�B�ʄA��=��"O| [A�Ȯg��c/,�,��"OBy�hP3&>(��AI*�H�s"O��Ru���d�B�@(�&���"O�j�"�	�S �W�0�P"O������n[�}���>K�Ь�G"O���#��q�)ڒ@#Gt���"O��S��CT'��kR�Q�11��)@"O60�«�j_���hٶ4#�"O|P�d�I�j@@�2���4�,"O�@S��W���@�����TwB�(C"O��C�C׫Ix�Qi2���H�X�6"O�ɱ�dZ�{��ͫ�/��	l����"OY�!/\  ZR��BHW)+pD�ٗ"O�q�@C�lx�#cgިk���P�"O�lK�&T<T�����o�t�2�� "O|iA�,���٧��#&�YzU"O\ȲX*��9[V�C��|@r"O�-�Q�j ��	���`V�lA"Ox�ۡ,�:m�d��qJ�i��h"OD8bC ��\��c'/0f���)V"O� �/<]���z���F:z!�E"O^���'�����+�"ԋ$(�S"O� �x{U�jHXAY�̓v�x2�"Oࡓ�O�B"؈ �Z�6�1�"O�Y$�ِ$���RS���>-vd��"O�����?Kr�HA���X�=��"O4A$!8<���M��L�`��'z��'��'7��'��'��'tj�1���<w���G�B���'\��'cr�'?��'a��'"�'R.@q��y�|$�QՁx�ځ g�'��'~��'��'�2�'���'6�0�M��
���U��1�� p�'�r�'n��'R�'2�'���'�Dq���+K>��`�3������ş�������џp��ݟ�����4qlڌ^Q�<��W P�t�ǂ������ԟ(�	���Iʟd����\�I������Ԫ�^�h�c�I���3��P�	�����ޟ<�I�,�I̟����h�7ɘ�!���4&��W�����JΟ$�	ڟ������	��	�$��̟{�f\�`��<h�c�� �x|��iP�������$��ƟX��ٟ��	џT�����I�Ε�!�����P��
V����D��ޟ����@�	���Iʟ��I��|�&��D�d�r���>�D�$������ ���0����d�Iß��I��$��6&��,H��[�e�6!W/_���ş��	џ��	�t��ȟ,���,۲�%M	����[�ТZ��Y�������h������	����7�M;��?Y�R��"��8a �i`��0k�	۟8�����
殮!KE����1@�x�Lj��@i�V�6��4��$�O�T�'�A�N���k��1Bj�O4�DZ~�,7�"?��O���i#��fZ�P��|�a,�!W4�}�'+ϝ��'52[� F��$�p=�j�C��L �S'�܉utj7�c�1O��?�#����/��AH �ʒ�
b��h3�k���?��yX�b>%�#E����%*�1�%��:s2� r�� ����y"�OR� ��4���d�2��1q���P	��TÄ�4c�D�<aL>�ҵi�� C�y��
�iܸ	�c#M
���@�#]�O*�'�b�'�d�>Q��^nX�3��E>�`%�B l~��'�@�g�B�ژO�B�	�Z���W�j�v�0��?Ѹl�թ�J<�	Xy������N�tµ$м²u*��2-'�L�E`e8?I1�ia�O��zϠ�٣`��_��A�N��"t��O����O�ԘD�lӔ��������ݺ ����diF�B�d;F_zf"�O���|z��?����?���(�����{��\�$FϏn.�	�+O�o-;|x�	ޟ��	�ޟ��� �/l��1	QAUF�P��̑�����O���3���MT����!����h���B�Y�"qmx���A:��tL���'�x�'�Z�9��@�Y�1���JWl�S6�'���'��t[���ش"0-k�f�����>(L���A�6PP��U�f��VD}��'-B�'��롮ֆ2�Y�r��8d6����4ț&�����(!y�Q>%�蒷�&mp���e$Ν"��:�:ON���O|��O����O`�?�3Aʻe��Y��=̼Ȫ��@y"�'%�6M������O� nZH�+(���c�/- ���oK#��%� �I���S�E(�}nZ~�
,7��[��O�N�ֹ����=%`,�#���|褚|2R��ɟ��	ǟ4��
K:u�P��C���wC�t2�N��X�I_yr�m�J����O����O<�'�~��gbڻn��p��:���'�&��?�����S�T!́yB���D�P(��|9�S)!¤�G�M�V��擖;k��?���a&~�R$NX�lG>8�DcʘB=����O����O���i�<��i��d�Vɘ�l:���C����є	O-k���'*6�1����$�O���	0���R�>q7�(zr��OP����1Pt7M&?IA��9���>�3�j4V�7�(d�4�JG;��my��'��'���'f�V>�q⦉j�Х�r��([���UnD�M3 �W��?1���?�K~:����wi��qC�OK���"�lK��'T��|��4�U2ۛ�:O�8�� �N-�X�6�̌.��:�9O}a����?���/�Ĭ<�'�?Yv���*�PFF��) ��R+�?i���?������F�-��N̟�I��l�$&�]�,YR��
�^ӴժCdHW�Tv�	͟X�	d�n���qF#��H"Z�`���sx����-ʆ�M�}R�M�����+�palQ#M4R��p�L��>h�I���I͟���L�Od���>X����W�ASԼ�����|`�l��5�t*�O:�$NǦ9�?ͻe�0�q� �\�Y�G ]�G����?���?!ìʸ�M��O�@�c�6����Tt
h���,��$i1��.3��'��I��P�IğX��ܟ$�	1\�8-�1j�$6d%��)���'F�6�-_	����O���.���O>���o])�li����&��ON}��'|��|��$L�J�~�1���YO����%��_��!���i���| ~i2��OڒO8�H�*Lp�m���zɣA!ܣ
�B���?����?���|�.O�����X�&�$_3���K� U�A�-W��$��I�?!�_��I����8V|$��I�$�ܡIW!�n��Ť���5�'cl�ծ�?��}2�{�? 00��$o
�Y��G'S��)�:O����OB���O
���O0�?��̏]��T"\�^p�A������I؟Ȋܴ0�}Χ�?�ӹi��'L���''�68B�h��+>8^�B�|��'X�O̶(�2�i(�i���g1+\Q���Ǆ݁ޖAd���h��'B�	�����ڟ���� ��e"�� \ �+�Bʼu�,�	韨�'Ɏ7��S�@��?�/��!���%#�ڰ�u	V�hLZp22���y�OZ�D)�)���^)'�[�ݘ[ͶA�c��*:���J�@ԙ�/O�(�?yg�6��7}y����Hi,�Z��T�,����O��$�O4��ɧ<�&�i��2G$ĕ|kh���-�C�>�oB�s@��'�7�2�������O�YA$k_\N�`�*}i�d��O��Į��7�-?�;r\f�)�'��_�����4`r�o$7���Rgp�ܗ'���'J��'���'	��R�~e�]D>�dK����*	�+u�� �I��%?��$�M�;�����d�}��D1:�(����?	N>�|J���+�M�';Z� �3LMC�A<l:Q;�'��y:��t?H>�(O�)�O"�����G�6��-�M�bH�Q�O��D�Ov��<��i�:�ˆ�'
B�'<�q�eE��͂F��lu������|}b�'|��[K*�$퀈Y�v�jfT���d��p��1�ɨM�1�b����H���%\`a���^������z��O@�d�OB�$�'�?��L�6�����%~T9�!Z�?�r�i9l��R��{�4���yg�]���Ź�K�5FC�l��eȌ�y��'���'Y�M!e�i6���1�|Mr�O7f�U��6
Б� �<J��
L�Iqy�OV��'�"�' Bm
 a�F	��,A
(�٫� =��ɼ�M�a��?����?yN~ΓG��)�qAރ����"��P�e��Z�|��̟�&�b>)8&��;�Ȑ�U�5���CP=A+��nZ��$8��z�'��'��	23�f�`�B]���Z�Ɏ�!d�Y�	ޟ��I��i>Ŕ'����=t��
�/R�9�u �
:����GW�q�2�{�
�x�O4���O@�D[�_0��C�`,[��؛57.D�uFe���bo�ܨ�����>}�ݭ��!��\�`�챳/��p�Ih�	ӟ��	��X��|�'65�}0�@� !���M�غ�J���?1��7�f�<�b+On�l�Z�;��aKW�
�4����烖)�lq$����Ɵ��oZ~��N�wl�r�ٖ"���xw�71/ڸX�G�p?�O>�+O����O��d�O܁��e�%1讠#!��+`W��T��O ���<��i����B�'�'b��P�t<{'�*^�
DJ3���[�Iӟ��Is�)B$�'cլ��U'ɦQ/JI�PgK2E"yꒉW�Gu�xZ/O�iɦ�?I�I4�
.SƜ��,�.e$$����8t_����O�d�O���I�<QC�ie��� \�:t�,�zs��� ���';b$n���l��O�d�
j���f�^9^��ز��_Hv���O<����lӜ�;`
G.����d���Jb���
 4���'��I����	ʟL��ϟ��	Z�t��,tsF�I .��\���26*�=H=�7mCu����O^� ��/�M�;L�;�B�1�ƭb�%	�H�R���?	K>�|jw�
)�M{�'r��T��?"(��;�)�'䊠x��s?9M>Y)OL���O�m�婍�<Xb��A�Ԙ�+��O��d�Oj���<ac�i�
�c�'���'��]K�b�.%����S-�[�p�J��D�N}��'�ҝ|bjM# �RQ���.�2���J������9 ]$Y�	s�pc>@��ON�$�1���ャJ���7Ȅ��b���O~�D�O��5ڧ�?IՃ�.J �`ƨыfA���3��?c�id�up�\����4���yG���NA�Tju������!�y�'�B�'ꂔ�Ƶi��I1p��H� �OP:��Я�J@����ŁXF��i7��h��Ky�O&Z�M����?��2������5uĹ�㍑�B	.()O�dmڼf���	ɟ��IZ�ɟ�D -T��3�g��qWS���d�O��*��i�{���Q�nJf� qp	\Y�����x���p8�*'̾�H%���'�(賷#E6��J� ]K$�B <�"�'���'��O%�1�Mbm@�?��̆x�8�@�.VMn|�qgʜ�<7�iJ�O��'���'\�Ӄ'K4գFظ���:C`��6�0�i��I�qJh�ПR���n'�,ٱ�&c��H
�f�/k���O���Oh���O ��:�O��qC��	;-�U[�G�!x���	ڟ��	��M;�L5��dGݦ�'����d�JP8!�������se�JO�	���i>ywa�ܦ��'>�=��hX�.@��9g EV��j',Q/S����������Ot�$�O~��=)v�ʵIŇ�Z�Ȇ�@����O�����!����' �S>i)�`�<'G�����1A@���;?�2W����Ο�'��'[��!�j��0��D���D<�E�5! �H�
-�"+��4����5T>�Ot誐���U�0��#A�0�`ub,�O��d�O��d�O1�z� ��fo,8��L��%��t!��d�zЊ��'Ol�v�t�O������J�G�5`�@�HN����$�O����Cz��Ӻ���V���H�<� ���YT��xÀc�zPI9O�˓�?���?9���?����ɍ-"nά1�R!x�aI�7-�hn�T��@������Z������;V��\Kj�Z`c�o6F�I��	��?�����S�'�ܴ�y2D-Bf�T���H$�b�a�_��yrM%iʈT�����d�O���[<M��p��LȞn�B��o�=+�2�D�O���Op�4p���D�b��'�RM'fd+&c�
X�m:�B+Y��Oj��'�"�'�'!�K�lr<�"��G�Z��c�Oz<�D��b���#��^��?q��O���
�������%��I�@�O���O.�D�Op�}���e��Y��ec��isVMK3}��4;�3s�f#��m���'�r7�-�i޽�
�?Ed�����D�y�-r�x��֟�I� �:�nZQ~R��j\y��T��!��&z��Yr��$��J>!*O����O����O8���O��ؠhG.5��3��Ol���� �<�i�ljC�'�b�'��O���>q`�z��?J��8��{&���?����S�'8Ո@� ��>J��Qg��nٸ݀�EF�`�m�)O�e3t�P��?���/���<���N�|TX|���^4d�>��F��?y��?9���?�'���-��͟� �*Y>H��T��Ok ���bvs��de;��O���'��U��C��J8|L�<�p�҈r
e��cӏ$֞�nZV~��ӃM�T��S.G�O�����u��"X�"�E�f��D��?����?����?����O���&/ʪ9����CJ1>Q&�*�'��'�6���ad�˓s���|rh�C����ψ�YLH-���D(��'����b����f��ZW��)JNBm�A��I���ͣt}4����O�OP��|����?q��R�x�*p�ż-�>��3ϝ�
V��8���?�(O^�mڳXPr��Ɵ���D�$�W6s�\�sh�'����,G
��DX}��'Br�|ʟ�y2F׸]�0��p�`��x�D��0c��{�d��|���X'�$���{��hŀҨ��$�d����Iǟt�	ӟb>y�'��7- QA�1��G���lP	���5F�!$�O����զ��?�AU�$�	�l��I�$OPL� ���G�B:.@��՟c��L����'TrD�$T�?���|��6L
'qf����JDL�v��"7O�ʓ�?����?���?!���IJ�z�ܜ��d���䱐־)aЄl�+��`�	����IV��������K��N�������^�J���?i���S�'x��z޴�y���+^�$��gU�0~��1T逶�y��	NuT���䓸�4� �DU+xDhd�R*�&R]��TaП 9����O.���O��"��v�(.�b�'���d�Ę�g�͌8?x�	ce��g��O���'tb�'=�'ː�8DB�p���Q�����O��(!�DbX����k0�IƘ�?��K�O�[��� �{��M0n��c'I�Oj�$�O����OT�}J�a��|��3
F��ϑ;1n�aJ��Û�m��b��'� 7m#�iޡ�Ŏ�z}pp��!&����e���wy�n��&��6��������;� ��7�n����e�#G,��p�|�U��������	ڟ����lZ���tT�Q�	:6�T��E�wy�
b������O��$�O<����$A�k�
S 6��"7��: (�'��'�ɧ�OĐ��eD�.-�65!#��^4uȲ�U^����_�p�t$�V6��l��Wy2��t�^�g"@�h����/ U�r�'�'��O��ɶ�M�/���?)�-G�H�ȴ�P2%��c�d)�?9Աi��O4y�'��Z�pЕ�\7J��	�E���eb�Ǻx�B]nx~���5p����r��O�ɗ�E�F��4%�Wѐ���l��y��'B�'���'�b��"d[>dh��ޣ/��Ĉ�H�������O���LǦ��� :ZǸim�'(}�A��(qf�#�/_�Dd\�q5�|��'�O�:H���i!�i��A+Ǆ >���1'� �LPp�@�0V�vP��:�'���Οl��ӟ��I�G(�� $Ċze*�߰}"&Q��̟��'��7ق`���O����|��ל[�%�C#�=)�*����_~��>����?�M>�O���AD�4_��=�����L�Ȥ
������i=�i>r&�Ot�Ot �!
� Q�"��R%\"i�`��3��OX���O����O1��� l�6�Ή!���T�*l.4�!۹Bl��'O��b�<⟜��O>�$	-qC�a����+Hvqy�M�$R˓J�-�ߴ��d�+>���'e�@�	�<��0�]�D[(I�sH8 ^p$̓��d�O����O����Ov��|*"!��1��<l ބ� ]�?>��fڢ3B��'r����'d6=�(���&�*H���}h3���O�b>!
��ަq�7��$�Ы��&�L@��I�P�ϓ���Bn�O�T�J>9*O����O�Ȳ&$ڦI\���%��jY6Dzs#�O���O��<�u�i�z��R�'R��'���X��H$<�~P�Y����D`}��'��|�� HM󡪞8�"i	�=��U=\6B�V��;~+`��{+|��]S�F%;�ሳo�&�"s��!=Z���O���O��$:�'�?	��N/~ϒ��BL�S���gi��?!6�i�ց�%Z����4���y��
�"����ZE��R@��y2�'1r�'�J���i�����D	PП� Ԙ�j�x��/V�M���ge$��<��?)���?���?��k\�!)ބ0��8~�.DYT+����1��
⟀�	ҟ��ґ��h���x�m^���!�e�����ß��Io�)��]��L��nV�L��m�P�گ:�L	�����'���2�h S?�L>i,O�";�Y��O=K�r��EZ���Ox�$�O��4�2ʓ!��$��-���R<`7��&O�n�#.ͯ �b@eӢ�lH�O�D�O����+ �����aiՠ�ǂ&��R��c�H�:�P�j(�'��[R��U��L����l�$!C���<Q���?���?1��?��t+v�T,���;=��al]�R�B�'L� dӬ�C�<�B�i�'��@r��g�~��5$^7��z��|2�'��O��\׺i��I� М�Q�>&�3���4�V����%A��4�Ĳ<)��?��?����.W�0}IEC�T�.��$.��?������p6A���I�h�O������z64�*/�R�e��OVd�'�r�'�ɧ�鞑)�Щ ����M��@�Աs�����X밈�����=��)�W�`L|i𓈆�-�X�-ul��	П������)�iy��}Ӻ����ɭi�����)B�T��a�*��~�ʓV���DCU}�'��<��F
�%
�����=F�إ��'d�bJ�*�������iI(oq�ȵ9�
! ��p"��,�`�1O�ʓ�?���?���?���)�?d���gċ3\�m�����U��Mo�T����I���u���i����ck��	��Ǧ���>�[7螭�?����S�'�<�ݴ�y��J� �P���Y�[|X��*5�yRU/!y�����a��'x�i>}���(��}{db]��hIܟB�`��	����̟P�'�F7��
Z `���Oj��:���$����m���{ �$�p}�'�2�|O��^%&�a���#^����ߤ���n+4��
i� b>]h�O���3P��m��
�F��t��C���$�O����O��S�OrLB$d���Њ$G����ɤ��~�*��(�O��D[Ħy�?�;��2����Z���	2��HzP���?����?QŘ�M��O�L3�О��KAk�qjD�S�w�L�i��X$�OJ��|2���?���?A�%��X`r��{W�躱� A���(O��m�#M����ğ�	}�Sğ��d�M���4j�/ю �"�n����O��b>IZ�(L*R:r��'� &Й�F��	N��#��[yrN�($,��%�'-�$?��,��̑8�~�j	&D���	˟p�I��i>ŕ'��6m�6cY.�D�W^.Lۀ��i-M�p]�� ����?�0]�l�Iʟ`��-}0åmP)g@&L�ᝍ^y����(Z��'7z�2�G^jO~���
�`AKV�*r�0���":6!��?����?���?����O�`���Ҷ�rzg�P8!�)S\�h�	��M�4l�|z�f:�Ɵ|�Śj<��gcc:�xDA�.՘'�B]�� �͔���'=Pt�Ƨ�,eZց���҉W�̹3U/��Sw���I	-T�'v�I՟����<�ɆY�X��B�	d�$m{��,	�0��֟��'�6��)J�����O��D�|Z�씪{�Bt�CLؔ%I�a5�f~"�>a���?�O>�O�\��0�I� �
=b��1U�ct���F��a�iI�i>��O4�Oj��e�O�T@��ǅ���i�1��OP�$�OT�d�O1��ʓGK�Fk�; I��ɐ�|�n4j@��&_b8���'��f�`�L��O���C)m�a���j����#^���9e0��ڴ��d{�(9��'.�t��ʁ�T��*X{�d���+5Ox��?A���?���?Y���IT�kl��P���"`������M�0�mڶt�$�	؟��Ij��؟�������"PSb"�/Ѭ2��)0���?1���S�'j��@�ڴ�y��h@�i�F,D�=���B���y��o�@D�������O���`=��r��Up���/X6V�����O����O8˓z���_�8���'����)L2.�;3�D�*]a	ǅ��v��O���'�2�'Y�'\B|�Ǎ'c@����l
)^y�`��O�������L����A�?�ĭ�Oҩ�%(B:G� �br��0���y�b�O��D�OL���OT�}�;c1L��'	�$Af��Ɗ!��Q�W�bP�;���'�d6�$�i�]y3��hy�T�da_X��D��Fz���Iş|�����l�N~�֬9�����s<�2ekE" 9
ճׄS�g���rM>�/O^�$�O.��O0��O�p"�fсV�&ਦ ܤ6P�I4��<IA�i� ��'�'�Ob�	g�ȉ�����h�@�OBQk���?A����ŞiX8y�V�"VL �l΃cV�Hg���M�O�Y#�݅�~B�|�^���V��>�6��R�K�8 cB�L�Iϟ��	ן�Ay�iw�ȑ0��O$W�.�Ըؕ�{3�Ab#R��?a"�i��O��'v��'���	m�.!Q����@p�H[�6L��i��	#mx�	0�OBq����J.v$ �p0ج��.�.�D�O����O0���O��D'�"b+�BuNˊ|N��4Kɫ�-�I蟀�	�M{#�>��Ć��Q%�$PW��(�����ހ.�"娦�P@������i>��6\���'ԭp
� Bd���F81�ָ�wK�fa�t�`M6�~��|�R��˟�	Ο��T,�v/��Y�T�"��8J@l����ITyB�dӬ��O����O˧�@�AeF"`�BM�u���'�<��?���S�$
\Mx�08Ǝ�a��G.S6J�����Ŵi�(��R��*��KX�ɬn򈠙 ��:<�
(3rGȭ0(����̟�������)��ay�(~�d\�PD�'t��Yn�>W�AO��D��d�OZ�mZ~�k��ҟ|�6m]7tN��Pe;oW�`��d�gy�=v�����pC�GZ�P�$�	ty"E�<�`���A	B�`�9�!�)�yr]���ȟ �I��0�	��<�Om�����H�S_~!I�jh{����r�{�:	b��OZ��O̒�X�$�Ԧ�݅t�B)�c�%1�Ą��T{�����ʟH&�b>A�	�̦=�?��8�҇�	9/r���*��dV��̓(}(�(��O��@N>1+O���O4H(D�M�k��q$���;��0"�OZ���O>�$�<�бi�r=��Y��I&J8d2�jc�V�)E�S�t�?�@Z�d�	k��<��9�%ܻL�\IHF���'���'�
a��枔(����T��՟��'���Ctm\6C�-*P�D� R���'�R�'yB�'��>�I^o"�����B��}ѐ�=(���I��MS�M�>������?ͻxs��#��l���"��b�lϓ�?���?�U�Ǭ�Ms�O&���L�8����"QzQ��I3J�*x�k
�T�2�O ��|"���?I��?	��GX��QOʤq�<���	��8(O��n��z�'7���D�'z�6ʻIb��ѕ#��X��q�tF�>���?�N>�|:b�S�(�>��M��y� h��G|��i��4^��Ɏ ~��Ӕ�Ob�O�˓pf���^��Z��TEc�)��?���?���|�/Oܥm�<"����ɯ!Ƶ��iy���Vn�*v*��	��M���>����?�;AX0��U&w�I�C!��Z��£��M��OP`ks���d��D�w���R7�ˡ�	���!z�	i�'�2�'���'��'=��˰�PaG�L�q�H�S�Z���O��d����C@�Uy�Ga�j�Op����P��t����B1�:�&���O��4����(j����^<	a�A�S�T}pr��T^�X�@�N�'�ԇ����4����O�$1I�u��_*:�|U�U )�T���O�˓K��&B�$�"�'rZ>�Ø
>��u:E	�X�� �&�.?DZ���IR�S�t�J1�A%��R�\<ï߃,��l��M�YNhE�Y��<6tB	Tu�	4 ��`{�(ǻ"��G9��\�I柠���)�y��e�R����>	����U�K3�Xc� ��iHL���O~�m�S�Qi�I̟���ԴL�J��zkH����f�p���O�h�#y�6�j���"���"�O:ܱsFħ4}D�R�	X.�؊�'e�	��4��͟�	͟L��Y�4/V�!�ũSh8:����4��i�:7m��+t�D�O^��?�i�O|�oz�)Q�I<8L&��b�K7�N���F���@�II�)�:[4<n��<!1�VV���JA�]�\p���<q�dr��' .<$�Ж���Łxb:I�,T?	7���t/�>3�axr�wӒ��d��O��$�O�5�bgh8$��C���&Nn��O���'k��'��'��xa�Ϊa�\�C� н����O|�P�BZ'FG�7�C`�0N���O��s5�G�p�ԍ�QæG��e"O.=��gF;j_��ZU��Z0(�9A�Oo��(��I�(bڴ���yǊ:fԜ:%�OvA���<�yb�'���'�8����iq�i�)Ƞ���?��IȨ4F��Ñj>؀�.�s��';�Iv�'��T�.�%�\��T�ƅ	~~B�bӢ��G!�O��$�O��?��̓%ٔ�	AJ ���%]���$�OX�$%��郊,{�9�Uꌿa�~�3��.y���cv�@��'t�J���]?1K>Y.O��l�7) �����y�fXB��'Z\6m� &���I��йj/A���A-U!�����ݦY�?�CW���I,���I\��XT!>��jEAZ�R�R� R"ҦQ�'GJ�J�*��?}�D����w�hp��D$���c�/Ǭm�RLJ�'��"�C<n0u��ؔO�����K�"�'�"{ӄ��w�?M0޴��+����j�6��·�2eP84�J>���?ͧ8��e+�4���ʷ%�tIipD��9���D�z�AՔ�~|�Z�t�?�'fS	?r��)��I"t���Iw�'�,7���O$����O>��|�q`EQz�hp�ߐN�d���x~��>���?AL>�O��Ɂ�ڛfn� �f�U��8�؉6�{!�V�$�i>A���'7J�%���h�c�\�����~v��@�3�<bڴ�`�kcѩ*<����,ٿ(�����E�8�?���@ʛV��Sr}r�'&h��5瞹8��� Rkđz�f��O���A'(�7>?�s�T�pq`��py�9Z�`�c,�
~��vH��y�U�,��I�n�����I�`ٓ%��<���شt���)��?�����O�6=��}��킟>�hq�
	�.�1Å�O���6��I�; 7-k�� ��b�b�/Z�|j0LB�0��X�?O��������~�|�U�����@a3̚2���+e���_:����ޟ�����4��eyri�,�!A�O&���O�]�¢P*_�x��֦{� ��f�:�I#����O���.�]�.o���6Cdd���çI��I$l��(� �ۦ!M~������ɛ��|�ï�U�Ӂ蔕 -h��Iퟘ�	��@�IQ�Oj�L2|&�����Y��F�T�2�gӀ<���O��DZ��?�;/\Bq�L-��=�-!SӐ�̓�?����?ٔ� �M��Oq�DH�4��T㒷Gͨ<�T̡�(�A��ƌ|�'��Iߟ,����p�	ݟ��	4F�ݘªнi*.�
��K#1Z�'��7m͠_���Ov��?�i�OT��j�� ̎��&O%)"�49���E}r�'���|��D�X<o�P��6m?��I�F��
7� �ӷiOd�4��T8ᇹ��%���'�j��`�E�.)ʌkpNN1|��=+c�'���'������\�X��4\w��I��6UF0��M�V*����$+��{�!ڛ���Kv}2�'��w��l���Cb^i�F�Cà��&��	g0�&�����۩/����J�������9@a����ПI�ଈ�Ev�����D�IٟD�I��"�� AuB]�̊�3�8���mQ&�?���?�r�i��<O�bGxӺ�O�Ek�M&�a��@)e�
*�e9���O
�4�<]��bӞ�Ӻ���0�t�PGeZ� #����"� t 00�pT4�Oʓ�?����?Y�����R ˽a{�l�W�����%J���?i/O@oZ�hz������	N��:[�1b`!��laa���y��'���?y���S��.)$@՘�Y"�	�EN�/���CR!�f�
aU����(�G�ɦR��Q�md<x�G�:r��,��ҟ�Iܟ�)��Wy*qӸ8�s�3���!W0g�� �R�z� �$�Ov	oZZ����
�O��D��	��I��  ~�sэ�5d����O,4vGhӰ�;hҨ�3��?Q�'ܔt.T��;�
I�5�z��R��y�Q���	����I՟�	���OZ٪bg��Lب �LJ&g$u!�#pӬ�s���O��$�O ����DE���E����H_�]y8t��V�2?BM��Ο�&�b>���F��4q�ؠ����s W-<�ϓ�Ĭ�Ai�OdՙH>�)O$���O>��G�:ਤP�^8j��hC��OF���Op�$�<� �i�z9���'�"�'L ɒu��w�D� ��B�=��a�Ք|B�'����?1���e9N��b36vW�� g���	.߅hb�$(�n�`�ӁieBn��427��w�@uKR�� D���"g�������I̟�F��w0J��QA��r}hS�׈�1��'.�6�E�l����O|�n�K�I�����!Ϟ��C�	���y*����x����O����O�u3!�rӔ�Ӻ��BC�J�L֜6�lp�" Q���\��O���?1���?i���?Q�.֩�q%�\k��R�(Z�1!
}b+Om� %Sș��۟��In��ٟ��d�� 4�:R�5�΄:����O��!��	��"���`��Y�r�&���ɑE��|Y�&n���'��(+&��C?qN>�+O�(�j�'���<��cKJ�a|B"h��u�a��O^-��iǷZ����/D�l�2C��OVpo�_���	ן��	�$kg�)>��p�!O�=���&���1��lS~���j����ӯ$�O�w��e�$�q0a�J;(���y��'z)Qb �8��L�P�H:� 6��O���O��m�B���ZC���|R�ǸU����'%�$P��r��C_g�'�����f_ћ���]�U�p!
e�� �>�{7� (hBT�O�㟸	p�|B_���?��Ə�	N��GڻI����c)Q~�'At7K*~�x�d�O>��|���I�yN !{d(�0,ѩG	�~"��>����?�O>�O��g�#7����O]�@�İ��X�q�D�B��i�h��|r4ʵ��'�DY"위�ʜX���3��xrU�:��9�4<k, �v�6(P��v�D�#�4���R"�?!�dԛ6���u}�'i�P#I�HiM��,�.<� �(��'7�H��{K�֗��HR'RFW�)�<)��ޞN��҄-5)�ѕbK�<�,O�D�O����O��$�O��'d�E�c+F&p���3�N��TR��i����D�'t�'5�Owb w��t��Зh^���(u!�?3n��$%�)�S�`1��n��<�Qɍ+?8u�C 5�(lX�<��CU'/��􉠨�N�l�9r�Q�ū��N��ҸA4JT�5�f�� aI�%�a�f�W*&|�D��_� �T�R@_ڢÁ�F	T��3�DBG1	D�]�2t�D�����̉l����0G��a�FE�<�"�B`t8i�OA�ccY�=���E�y��-Q0�!TĈ����:B�|9� C��hɄ4@��o3v$��Θ4Qd�8sת��8\x(P&�J�I����G�4y�B�(�	s�ֵ��GO�U�H�q�E\�!P��^,�G+x���s�ːN����C�Ѳ
&L�WA�\d���'xB��g'���CO�0I��[��U�Ti 6��O��O����O���O��'t<ۦ��k>��H#ᑆx~��I�4�?������O�N`�O+��'���n34B�,p���nG�	` ��:�O��$�OX9�7�(�IG���1Z�| Ӱ+Ɇy���9�k즑�'AN��$�l����O~�$��Ԑէ5�l�.[��Rũ�&X`�2���M���?y)���?K>���� 4j�M�}9�<*E,��N�*��iE���PCg�:�$�OH�������'��	�h�L�UJ�*_�M�5�ظ��Z�4C���[������O�	�%Z��Mq�ǔ�,B��2@��7��O���OJ-��v}�W����^?�M�B�(�j��*~P(�`�k���$��W�
��'�?���?Ie��, U͍%�q�1d��a͛��'���!�>1.O:�$4���`xǉ����4�Q�� 3�IWQ�x
G��L������� �'�@�¤�,<e�𪉣c�|�F-��L&����Ob�O<���O�-�T�כ`VPb�UY� 8Ej�Xn���<���?�����.z��!ͧK�J�	��Ǳ��p�kN�v-h�lhyb�'P�'?r�'�j���OTT�g��#W̵K�F]�VS��#�R�x�Iڟ|�IQyb�W-v��ꧠ?�g�FL�ҳ��`>\�
����.
�l�ɟ&�$��ɟ��w,�Jܓ��$p� �ᐩ���ؔ32X`lZן��IryB��E����?!��:�l?�@䱃+7;B�zs�6w��'w��'މ�����?�XSO��`��}*&8!�n hvjz��˓4�f�C�i��'��O�n��;�"X7Y@���=R0t�c��Iȟ����G�׸O���`,�7[�<�Zd"�o��h��4��`�S�i��'X��O�lO��W�rX\��ޤ5*4��ʆ��nem�˟x��͟�$���<���W$i��8yG
�s�:yb���i_2�'�RJ�A\�O��O��Ƀts̚��
!�|x"�Mׯ/s�6�OޓO�������O��	�A
I�b�2G���!�҉#��6��O�����<I�W?}�?�P�/A��Y�Jښ
.���Q(��V�'��B�O�D�O���<��b\�K�&�U*�h���[q������#�x��'_|�R��]����1����4� a���RY�7��OJ�O��Ļ<i�g���Odx�:v���E?؈��&�
޴�?�����'0"^���ih�ri!����w�I)w��x-F=cpT������ICy�R�)���,9�X}�B˃�!�� j�[9(6m�On�Op��|z����ӡ"����������	C�0�6��O�ʓ�?������i�O>���k�\�W:�`A�[���|�S`�M�'4�W�`C%f8�Ӻ�0%�#��@C�"�9A�ԣ�P}��'�`��'�2�'V��Oq�i���뀣X`>� Y�/�% 7Hj�|�$�<���G��ħT���!��'}[�1#��\�knD!m� yF��	����	�,�S^yʟ���T��(ujr9jB/ۨB�Ea�N�D}b$���O1� �D��S��a�g#����3O�<@ڊ�mZ���I��(J`[���|R��~�M�E�v!��ݛAr>����*�M�����C��3?���~�M�9%���(��.)��� ��M������-O\��Op�O�)�Ϛdy�)����(8%���f�Ɉ.��c�D�IGy��'5x��B�H>d҅�%g�kl�5�	/5�	ڟ���h���?�'Ū�*��?=�R܀�f®4�	ٴ,Z���'�b�'�_�� DiS&��d�ֿ.f���3�-�l9�/�>���Oh�+�$�<ͧ�?���H�4ʬ��u�^I���OJ�L��I���	��`�'+���AE)�i��^�v�B�дo�~�P�CC�Z\tn�ޟ&������'7�'Z\�	S�	ZI�\�P���b)��oZ��x�'	�KT�.��͟`�I�?��,#I�T$B
P��p0��	:g�O��ĳ<��J�_��uwꘌ_U1�t-[�5 �	�E���M�)O������1�����d�x�'��b���%���P$/O�!�l��4���O���x�H�s�p��M#ٔ ۀ�'nR��@ǽi��H{Ӑ���O������d'���wCv�����y>|�����91(ȑ�޴�?���?1O>�����"�yIC�6��X��
�
���n�����ܟ 
Є�Zyʟ��'֒X��P�>��9b�/뮴��6�	��O�B�'Pr-DL�.�r5$��b�)
q냁�~7��OV��F�a}"_�(�ISy2��5v��j�r���۱&Ϝ��e`���M���J���?y���?)��?9/O����J74	�T��\�wj�"`陘~�}�'���D�'�B�'��@֔�8�@CBטt��"G
��Gĸ`��O����O���OJ�9P9b�5���0�� +[�@s,�G�d��iN��ӟt�'Or�'N�FG�y��%k�=AbHI>�˴��]��6m�O:���O��$�<a%�πP��S��Hc�Z3D���@�-ؙ�@�ΰ�ֳi��R� ������Ɏkj�I�T�I=D�N���m,
iS�F��0ܴ�?	���Ǭy&2��O���'����&X�q��QY��[Cnʓ � ��?����?��m�<�M>��O��i�qp�
�N��h���4���إbt�l퟼��ӟ�������PD���-R��w'[yx���#�i���'|����'}�'�q��0ڲ%S b��)�EZ,"s(}�6�i��|�u�"���O��D��0��'D�ɘ-b��a���9&�r���?�i��4k>dΓ��d�O��?��IV�t�K�ҟ. �٢�	d����ٴ�?���?���A�B8��_yr�'��Ğ9a�@|�A�ȜA@v��4)7:��|"*��yʟt���O��dXd�? 8`׎�>z�t�rf�Ԉ�^<��i����^6�����OJ��?���f5pBR�;��S�� *�H��'7@�@�'��⟤��ğ��';x|��m�~3�X���I��ٰ�(K�8'����$�Ohʓ�?���?	 ��X����޽<�pY��55$H��?���?Y���?	-O"��PM�|:"��LY�&�#,�,9��Yʦy�'�RX�|��ɟ��	1RG��	6��a!bh
6&�$�S�U�o65�O���O����<��'݄���d!2k�5<$1[�& 
u&��A���M�����d�O����O� �5O��'�4�cE�	y�ua&U�X���4�?y���$�2i"��OT��'y����"}/����	�af��H�	Uf�"듯?9��?��Lq~RV����%WZL2�� $(��H�Æ�IR~�lKy�N����7-�OH���O��p}Zw)�$�
lc<,���l]Ȧ!�I̟\�Ut����ry��W.�.�8�#D�s�Xp �h��iTG|6��O��֛6�O�z���D�$S��RG�]	�b!2���
<rl�9K�*����+�������B��ar�~��K9�MK��?I�""n��0_��'%��O�M��X2oڈ� ��.1p�ǽi[�]��;��|��'�?���?��i�c��e�3H�L^\	t �uܛf�'�d����>/O��d�<�����c0Jl�G�[�T�3w�[v}bcY�y��'�R�'�^>�	�F���jwcG�R} �D��{�$Q)�/X���<������O���O� �A_�b.�M��ۍ9�%��
05��O��d�O��d�O�˓hL��5<��1ˇ���`=X4HT"��S;qS�i��	��Ж'��'�rb���i�#$��� ���""�=r��=����'}��'^�P�0�'A���i�Ok�^ �d%˒���\��$�g7@{�V�'J��՟�	՟,�A�'?�'�B�;��٪��ݐf�[�-�1�޴�?����$Z�{ (�$>��I�?�;�/s9�Iq��!7��S�����?���k<���������I%Q��t�d;�P��ďǓ�M�,OF)��
R�uX��2�d��h�'�噓c�"u��C��Zΰ��4�?i�Y[��Γ��޸O������)X��DD]�O��ժ�4zB��3�i���'���O�`Oh��Տa3�0�1���G�L�c���5�dmZ,q�u�?	����'T�!H1������%�:���}�0�D�Oz��E��'���I�L��i�uc�#
9b&�jG��*f"ao�|�Ɉ6�.�)���?���z����o�3%�vyЧ)7	n��c�i"�2c�L��D�i��y�'Ӷw��)@�����9"�!�>�%�Q�<A-O��$�O.��\�k��U�s�t�E�%�\�	��L����>�����?��C����שP�X�8�HD�����w|��D�<����?A����$	�@o:\�'OPhȹs
]�Q���A(��2`)�'���'��'���'�$��'6�DB� O�5W& �󪄨�T�9�ϲ>���?�����*{��$>%���^�HJ)��_P��0�#�M�����?	��=�:!͓��ɬ�h���X!j�pY�c�A3ha���'���- �d��I|����2F�<.�j�����c� ����C�=@�'�b�'�V5R��'��'z�I�+Y5�	Q�D�/-m ��!�,$�6[��9�,ͺ�McCR?��I�?M��O�`"��Ѓ)V�x�3	�k�BQI�i�"�'E`�!U�'
�'yq�R��<[���ɑ��cf�A�2�i��0ћ&�'�R�'���I:�	1lƙȲ��Z~�y�a�V��lCش8�� ��䓓�O�2&�+ߺ���$&�X��ф�|�67��O����O
�k�/�O���|"���~���Dp �c$��a˄��Ջ��
��	;��'�?y���?��Ȝ�Kq ���䌞dޠ)I&C�f�'������>92T?���ȟ��OԵ���E� gj�Yq��+RL��xR�|��'��'-�'�-YW!1j�"��R�K�W����Zp(Qw�'��'���'�'���O�@�cǻ>�ČJdgAO��=�iW���O:�$�O���?�uf�#�?��=s��4ah` ��}q�F�'�2�'q�'�"Z�p��l��$ٗ�Ӕ\DA�-I��I�V���	����y�,ò((�����싵]��8���'^��B��˦��IZ�I؟�D}�ɣV��H��O��@w^%H�M���?y)O����k�S��ӧV�PИ�AV�!r��q &K�.�~xIH<���?)F�NS�']��M�ꈹF�J�(�x8�҃��<���Q�찄�Y$�M���?����J�S���8'�X�S�:~�� vA*CB7��O���CW��Hh��'�q���2����nP.�����g�A��i���[4aj�����O������A�'��I7d�y��eS�q'���]�3��jݴ^��Gx����O���v�\��`��NG B�`|@�-�æ��	П��	�l�Eb�O�ʓ�?�'L{�ꏌ(�0´��#+$"�4�?�)O����=O�S�P���{��{�l|z�K��I��,+c���M���;�|-�Y��'�T���i����$C�$c�8iR�ε<��Q� f�^���
	T��<���?�����DËU%Bm��&� p� Io����xA"f}�X����Ry��'��'�x�e��!iH�#S*�
~ �Ң),�y��'�r�'��'k剽����π  e)u�$)�Z��PgP �L��i��	ߟ�'�2�'}2A���y��>�=#��U�E��˛�u�7M�Ov��O����<Qd��&�����X-1}r�#�́�qv�\�uǌ�Rh�6��O���?I���?I��<�+O��:P��H1��!���e�v�9�٦	�I�4�'�"�$�~2��?��'Z2B��w�E]-.��*vGA�����O��d�OP�D=O����O��D�?��V�O�N�	���N��FJ~���V~�4�F�i���'B�O,N�Ӻ��N�=�� 
sC�7Y��!��-�IП���ep���I��If�'}�M��Ĩwނ��j�z|
��I`g����K�]>�����U�~ 
�C�Z!�4+���)Q���6���>!�<�r(Șɠ��q�Q�'=@8�SL� ?��\iЏ�
�Fuڒ��45�lYR�j��.�*�@R���1Z�F�&e>�K�)	*��|p �SB��e��:�zA ���+�њeE�2MnS+��H�x��S�ciÄ!]<b�������|���O���OJ��;�?A�����"_�<0`$ֈ�@[3�V7�M�f^�4 "����@�`�#��0�[���3�)±n������5�c�D�b�b��e��+�NY(R�_:�JJ%鉫x1X]R��{�Yj&J��cP$����O�D?ړ��'n�р�Ë�7��13tLA�"h�p�'	ta���9
\Jpġļà��y2N�>�(O����M�V}��'�\ �Ƣ?kr����\<Y4�Y��'<"� /	X��'���$Q�H�acP�-(�U�(�Tp�۲�BD�F��R�,��I�X��{×�c����'��`����?X\%m׭qƐa�L���	����'�p�!Cޭ**T1��U�k.	a�y��'-ΙS!K޷b���`@Ô]��|
�'�06�ǉbQΙ0�&�'�Ήʠ����Ŀ<� I@�RL����L�O���'��Kd���a����F�7B�Q`��'��(Q*�"e�by �l�O�Sz��j^�(�l�J�bK;;�=�îY����Az��
�eЪْI
�_T�O�$=�g��6r|R���$9�eHL��ऀ�O���5ڧ�?��m-sV>��/ϼOC���U�<�W��k�V�2��ϵK4 ��
QI��8����Z���(���t:�M�$�(nZß,�I՟`��E�M��	�h�	ҟ��0{@>�S埌Q$rPIۀ��'� b.�9����,��t�cJ�#�d�v'W�q��U���"?��+����>�O཈c�D��� �+ܨ�z��O\�	T��)��O���O����*�
�d�R ��G�hHbb�)��!|O�#���su�A��G�����u���{�4�?AH>�OM�I�[R#���H�
uXVѺMN*�qc���>���ȟ���ٟ�Sß��I�|��@ͱR���R��6(��Z�KN�/�Ԋ������>4l�+lV�s�7+���׍K�(/���$M*��>	�$�
�l$�J$KH�����[�"
����ϟ��I���'%����==^(�"�D�9���Y�n)\�!��-8��t���t��M��͚�1O\�l�۟��?�O�x�dH� O@ ��a&��0�'�(Tr��"��	���"s�	��'�VPĪC�'v���cRh4Li��'>����ה�-뒠	%*�ҩ�
�'P�HDt�d}��F�ObJ��	�'�TY��H�m7>�����#]ֆ��	�'�0�SN�2v	�cM-W�|�[	�'�P�����S��T����R�~M��'�-�VC
�^�Č�G>��+�'��Ƨɰp�"�Ɣ?gZt�
�'��l���I'@.�lK���KP(J
�'7I�E�.�>�@���C�\X��'����<�Ty��/�`�1�'�j���(H�Ҋѳ6'Z�+���;�'הaЂ����Y���� ���'qF���̌"@}�9������͊�'��ŐQG#im�`�$b��ꜝ��'6�����������I��)�'`������6Gf|L(wdL=Q�T��'�����ƨ&�r�/�V��yC�'�65`�%/�J�	3B5� j�'o����
B�]��s¬�wyFdc�'�,L�w�Т&��%ÒǚtrDt��'{.q)�B�����ܞd�4���� ��RD8���ٳ�R�B�<��"OX(I@��(����˟ :��8�"OL5�h�%����׻0��!�E"O֨A��8��Z��J$��"O%��D�r8r�@K�6�Dx�"O���{���6j:Fe�a�%M��yRf ���9)�B
-��LCe����y�_'VR�9yf�M�+�H���G �y��];<�]�%�n�Kq�ײ�yr�e�H�'Ć�oC5�`L�&�yb^::�t��iǈXb�"��'�y""ӘY���$�B�dZ�
�a�y�GU࠼�c��rî�
�y�ߠ(����˫?���`��B�y� [�>��b���;�b-dF�1�y"l��+e<pXT��==:�	u�2�Py�E��8"|�X2	�%��Cu��s�<���T)����h��66�3�E�G�<y�ɏ����7h��I�8I['��l�<a#�ʨҷjz�4m�G�
j�<i�NĎc�� nI�����rTd�<A�^9��g��_�����BV�<�2�����2D�i��08�.j�<	f�1kбp��݇`~\i�&�P�<��
tp�r��P���Bd�<a��H�wy���fC"��k@z�<��C�\��i�"���JA�]�<� @� J���J4�U�f�����/�[�<�g�U�_:ְ���ү��%藯�Y�<�)Y(H���F����+�$AY�<��� "*	�e�vK�<;��)q��V�<9*��xpe�RK�*�<m(p+�R�<Q	��yԁk��-��z��N�<�&OM29�a*�iצ{�b�Z�DQB�<ف�[�#X"C�  �1rQ��f�<1�G�HJ�T���<�0�Rf	a�<����b9��i S�r5��&Q_�<�3mˤ+�T�Ƅ��o�t;�Pw�<����ybR��g�*��'�Wh�<�T.R��Ĩ��]H�*�	�e�<)Ǯ��%�0�� GQY-���y"X.Wz�Ap�ÛG٤q���yr�� _���L�k�:=��G�y��E�?Ȥ�"o�'^�6(��(��yB&�3�Ĉ�t�C��l��c��y���!O�*|�*���T���$� �y�� 8{��uH"�
h���p���y"O'<�N���`�4u����y�W��B�a�&���L	d�_(��'���K�$*�'��$�A冷9tB`�E�.	XM�ȓW�RupW��	\a���Ub
�Rc�u9�,Ts��+M{��IU�����e7�a˃�ɧW�l��	<a~���'z��Mв.�t��dJ�8�����T��?��I(E@����-�,���D|�WM� ��'���"� �<�@���C�E��rtk���/���B�-��(�$ r�FY�"O��×B+ d�S�=65�$H�
,H�]j2[�Y�R+Y�d����F#0D�S����w��87$Q�F���F	��P`�H�'�z��]�kEFi�`L.*&i�SR^R��Rl��i$��m�$Yu���'#�ls�'jS4��'�b��/�[ǆl
�$V���Ó8	�x�lBDa�9#� �3���Zᚖ\Y�Yjf��6�ځ*�FI��.�4��yUU�1B��$�U�N��ТΎx^��L����I�]q�b�$!�\x�FŹ2����S?)j`.�Q�����]����cR�c%Ժ#�!��C�X\@�ģ¡!-\ ��]۸ŉ�	�- ���n�5,�j�3�C�\TP�AD�ã%%]��Og�@�^�8�C�@��������xb�P��� ��(��؅2���fғ&��q)�^�f�|kebh��*D�����Z)�`5�Q#���U�� S��7�@�{���g�ax��rߖ�� ĻFv�<�ӦH1�&�x��I��J�$��&`��[�e�oy�*�<Ó	�t��Lm������Cl�'Z44 ��`GX9!2m��<r�J��O�O���Zh�J�$�(A�kн�y"aKMT���4G�`��<�S�]�_���Bi.�� �'=~���x�^�����!�2tIW�Z۰��Anƈ1�a2�Olâ�A�?ʚQ����4tz`mR7�a�h9�KIJ�tT��F�j�0:���G�j9`�	��2�u��ι2�
�>q���#�X%+H�]�)ץ����v.��~�<%���P�c^�qf�T!g����#BH`E"#^��p��+s���'x(q @ӵZ<���w�ӨP�X�J�O�O�r�c�
\��|mmk���
�'6b�V̇Q��zP@��4��$:f+��-E|�q�OL}�,�Q�ӣB
��)O���PM�i�����h��R�@�ʴ
O�@�ү�-	LT��o�L��0�KQ�}jҖ�T;x&��0aZ s=���Qh ��G���1B�I�����	?��3F�Y�?i����0�IC4����]���EzҌZ�+����L=5%�-�&�D1dIjg�<�I,��*�J_�suԕz� �Hܧ
mh�3�}�����P� �%��%� ����sd�
���%~x�(PFP0l��;CnM� ��D1�g?�@�4}di��֝��%Zӎ�^�<9&�Z*c��]�D%�J�l��]�<1b����=��f���<�R��|K�����T��J�QX�4�� c�
���M�R��,	��
2�
�qb��y�Y�\D��T\�.q�a��k�9ÈO|0��3�'h�i���CR�A��GJd,�ȓ2|���6휕4�5��	D�\�ȓm5��f�lV��	�u4y�ȓ6.$d�#K"	xL�#~:����o�i�I?<n��Cq��=[�H0�ȓ8q*s7���A.
����@vC��ȓ&�:,�s˗2Q����P�͎C�#��i(&fz���bg��"A�jC䉉AB9�6DG�-$^��U��-�J���%2�La	�҈ ����(D$ވ!��܇�	�|+�\��?OV�3i���e���!L�$$�'"OZ0
K�$W�Y����O}�����I�~3JJ��5N�3&V���Ⱥ���4@��B�I/E��2M
 )R�J�Э5����Ě�%۴�"~�ɸ/
^(��	�h��"M/RbB�	�Tu �	�M�	iL�a,�3	��j�^h���'�̽���϶$��ٶmo^�"�'T� G�����)Ua�)�����'-r�smM�dm6�u�!��1�
�'H������m�hX+e���: �ĩ�'��|;C���	~�|��@�9[�1@	�'�����"����-���?~P]3	�'� O�-���IFj]"!��'h����?E�H��0NLR��i�
�'*�9p��
�QF���J�L��	�'����["J�UgPt���1ZC��<�ڑ�Ԍ�YO|�˝E�B�I�� �A��.�,��0ilC�I?���`��P��%�sK >u$B�ɨ(3�z�E	h�昪6BIFFB�I�+�¨����?zM����dW~BB�Ɏ"'F�q��9h<ڀ-�g�BB�	�D���������. �C��~�XB��B� ��mR�;d��B�kc|B䉩t�*���)�=��b�#�ZB䉼��0��I�[�����NNq��B�I�eÈĺ@i^r^Z}��-�_�C�ɛ"#p�	"�Z�%�Fej�Fŀm��C�I�Ys�Y"�J{���s!�@t|B�)� (�����3�"��B�6!�
�K�"O���`�e���[��O�� Q"O�|��'��nҎ%H7�Xg�2�"O�Q�-w��3�/ן,f���"O��M�Pl�e*);D�@ 9"O�y�Poف6�&���AG�:�@!�"O�y�V�T+F�v��p��]���w"O.L��&I��5p0�����"ObxRC�\�J��)X�Þ-p�0��"O��J3�9�*4c��h��"O�e:��F2v8�a�<Y^�Qq"Otu�֠l&y���oF�"Of��AG!ތ�(��̸O�$���"O���W/�K�f@�/��(��qq�"O؍Ru�dx��P�F�#�p��'L��"@D��	�ȟd��t��'��Ǎ�wک� �ӷ[�t\��'Z0�*栃�0j�x�ɐU{~t��'F)��癡,Z T�b-ɓ�L]��'E�*ZU��@e#Q��I
�'Y���6��o�شBM�EX
�'nd��CӡSjTI�GJv$e��'K����Կ4�mtI�zV���'d�yґ��E-��8D�	t�
���'"��]�+�� #d��8���j�'Xn9��CM:eZC�^�6�����'�81��+G5XD�A�'-����'��;��|��))%ϖ�'��9�'�`up��J'����1iU�"�0�'�x�:��
*qHޤ�⍺"�PE+
�'NT=�3eݮ�ڨ��A#%-�
�':Lupa��(\�>yy`E�#NJ�8�
�'+bq��3l�ܒ7Ȇz�2D"
�'WppS��*v�
TK�%�u`
�'lƱqǡ�lO��٣� ���	�'T���͂�e�,S"��~����'+���"�ŠP�uH�&&uA��	�'��z�q#bݠ��Ԙp3~���"OHɥ� f�&���Ē����ʏN�<�ucٕMN�l�e&��o�8͸�̉K�<����U@�m¢�Ӡ�~�� �FL�<���1��(����%.������Q�<IG�T.f��ի%;!��HB�~�<q A2_���RA��AG�����Ev�<i�,F�R�\ic�H�b! ��u�<q��Y��H���B�'��H�"s�<i��(x���,-�JQH�Lp�<)N��H��7߲"��1s��s�<��(��F��| 6�8�]�(�U�<ѧ,j28���/H�J 0aI�Q�<!�-����z�ō�;̺�S�&�M�<��(��v8�a
�H�")LЫ�̞F�<���E������6�d���d�}�<���.�U���b�6}��
Nx�<����V���F�� T�u�<q�jۛD+�e�%�u�)��ϢT=hB䉭-s��$�O�b8%��$0C�	�qv�Xv�D�{����j~�B�	)~�{fk�& 	��	�g��B�N��$�]?y�d)(ԁE�c��U��DeB�+��ϊ�*�֧��2��t��P{�0q2�5��p3f�; w�t�ȓY����E�1�P��G&����ȓ(������tbѢ��hu��S�? J�0�$��kY�d�i�)�6�P"O��6"8�t�2�ߩQ=j !"O�$���HX1P3A�.n�U"O%Q�V.l�����@�a+~]�b"OP����ȍ"ֈ3���]%T��"O����gn��A`L߅O� �6"O2,��	�*~���?)f8�v"O�9��xj\���E;	diz�"O�Y�$��8��,X@K��Y�JY!g"O�%�Ō�-���v�]2RK��y�"O��Xw��7?#�����0�y*"O:pr)�����S�H�y�A2b"O`YP��KQH����n�q�f"O��Y3%�O5�!pc(�o̘|j�"O\	9#ҙ_�bm��F�P��&"O޹"��[�G!�]��g�,����"O@�����_!rx�@��P����"Ohd��#�e�P�F*^9E�`���"O�l��I�Cu�GJϖi�V�B"O��be�q�zd�B�D���x�'"O4�@�,b��&i
-~��a&"O��1�-CWxb��z.%h"O��R ��U_`	"�Q�/_0H� "O���D�8%��:ck�sG��qb"OT-ň'5R��ak�+��a��"O`u9��%R��tj�2]<=�"O��b�MG�u2q��^�"m{S"O��HC&]����'�ǭ
�!��"O���`�V
T���4&�7D����"O�[��ĿE~�{ &A�4��H��"O [��$�r�j"�
 ��2"OL|���*x�LPA�M��*��XP"O$�K#"И�h(�&��]+h�"O2��c�ַ*le�u�l��"O�Uh#�ρQ�t�˴c���"O$�s$����@�I�8�R"O���#�1f�*I#���ٱ"O�5�`/](&P:�
"`CF"O^�P���?'-Ґ��hۨe��X�"ON���Ɇ�� U�
�p��@w"O��V�R�T%��Be�ɅF����F"O���ύ�q���#w�՘,
F=P�"O�����P%J�X�ѣ�{�rL#�"O6Pz�ꄰP�zd�N�g�0E"O�و%�A�9�9�H�C�T�@�"O�9@�Ό|�*�W�݇�6Aiu"O������P��!(A��	�ڝK�"O8�diW#0(\X
f�߁0�Ѻ�"Ot|�0C[������$���T"One��b���B�I�%b�qX'"O �J�c�at	�I�!�D �7"Od��᧟�9ѦR��j��Mh1!�dN�V���3�;`�� �3���-!�C!�^łGJ�(tx�9ssA�!!��T�!Z�@&XZ0	�aBA�i!�$K�x4d��Ł���
uZb�G�w�!�]�"&%��Λ����R 
�F�!��"����E�"T�z�KqMMv!��C /�ĠP��$ߢ�Y����W�!�ą�t22\Z�M�*{�t$��� /�!�$��!�� ���O�&�>��!$�!�ĉ�(1�����O�J������8;u!�DU�Sx��5�Z�N���ڣ�D3zu!�$.��qH��L�^�����%h�'��|
� Pm`q�S�5�z�+�HI����"O~8����$��9��h��l���E"O���@D$Ҭ2��҇^����"O��"S�T4��)��H.?p���"O�����ݲ�g�1v��i��d_Q�L��i�$`i�Fb�jA!�S*���S͔ Kr\r�!]�],!�T�cz*����G<�a!y7!�Ube�d��ůEz�ɀ�]��!�ēA.� �^��3�9E!�d��j��s�Ʒ'H0|�c-�+/�!�$
_�R�����]d-����2Ex!��^@ሠ34�&>T�艥�)iX!򄑩	$�
�*PM�c�N!�D��&�;�#ڍ2�UP� �3;!�$K�$i�6ɯ?䨨ȣa�!���	�\��*�!E����	i�!�Q eWF��F�R��X���!�$�=~h�)�*¦K��	�Y$Q�!򤝻0
�4K��\�?����&d 9/�!�DS1� a0Wş'��4,�1�!�ڼel�h�Պ٪k58z��]-b!��(�T�+$�SO%ڄȁKB�?Q!�}OXEၥ�j$y�
["J�!��L�y/z�g@�3΀�$R�ZA!�βL&�L����o����4:!�8S�}S0XJ�Xl�7 K7dL!�d�#$��暘ksd)x$�Z��!�ta��H&v���h�<n4���'����0-@>���۲ ���$a�'���P�n�#_���Se�}���'q�L+��S�>D�Ód��^>��a�'�HE��*Gu@�a�K�Pa�tz
�'F(<q�-Z���*W�P9Hn&I�	�'��LhuJ� �6p
�I�
@"v8�'l8�IRNH�(R��6�S8I��U)
�'�v�� ˭>Z�l�V��A޴�{�'�f�w+10RtS���
D�c�'���p�@n�I���s�Y"�'߮M��b_-b)��:����M�F�Q
�'�PA#�Z$��dI'%U$F�"-
�'!��"���� �̏�E�ġ��'�|-����P�Q%Q!��l��'��!
@�N�3ҡJ���'�� �E�"�#����Lp��'vd�b��?;Tℑ�/	
G�T��'7P�e͑7d)�q�V�MR���'|6�����$ ��3}4�a��'���Z�
Ja�LF�y�4�
�'�q�����]��� ��jx`	�'y��1��hWfI����&[�z�'�*�"F�'@,����LG�&�<�@�'�}��FKF�A����U�
�'7�x�ĝ�q�h��a
'<L9��+<O�e���S�4��T�@ 9�t�A"Od��F� /��l
��:�b�B"OI9��P�k:�Ɔ�+/;�t��"O\��6H��n�;1�]�}2�	b"O����-O/k8&�Bs�C n~���"O�h���/}�P�ԫT�L1���'9��ps���R¬���F/~Qp���D�s�<�!�:'�~��6玟?.$�C�q�<!�iUv|y�2/��Ey��q��k�<�R��%��L��$UD@�
及k�<� ~�1ǋ>XA�8"�%�!�ހ# "O���(��,�DF�!r��q*C"O�
��2T�E�S+������"Or0YS�Y�s� qDA$8�� "O��gMK�l/�b�b���rl��"O��AB�Z�PT���lI�-��| "Ol�8%��{��2G�i� ��"O�ڢ�ץ@������#cv��q�"OFt��k{�Z�!!� {tΠ2�"OBE���S\U*�A�o����"O������9���ᄉ�%li,#B"O�qģ� � 8B��K�7T��!�"O�x��q��@���!�R���"O̜S�f��Vq��˟��u	�"O�(�(��7����-��I��"O|�����[�|�%�߄��`6"O�U/��q! `Sqb�%��S0"O"0b�d�!m��� �9^��h��"O��JV!*��U`2��".�����"On��vfJ�M��9y�fB�i��1"�"O�,3.%
��e�% �t�h�"On����|1J�d8g�v�9�"O��03�S���lQ�H�E�5�v"O��(+��rO�`�\N�^��"O�L:!싮{�r!)�٦�+&D�2dG�uB�ɵ�\���Y��h'D�l�A≽E�ꈁ�ޖCd�P��&D������2T'$}�0i���ĩ2�-?D�����/�Fq����4W��1ȅ�2D�(:���:Wo�����E�kŭ5D��XW&�lF.(q�B��j}f�-D���uBY44n�L3E��/;��@�H,D� *`/�!}=�5�ٛ'��=��*D��������A;w1f���#'D������)�8Lz�iϩ(�F��$D�0�&�0H��刢 �*���"D��2� }^bXz���h��ബ"D���TL�f��:$�Ǿ*��"4A D�����#�9x��ڟfg()k��"D���v凄W��I����[^D<p�#<D����.�G��T�7ED�Fw�p��%D��kē��>i��`B�
d����o D�\�f��'�Z��q/�f�Ny�b�9D�Dzq��?BiD����&:�BR�5D�hA�#���	�)�'�ƍ�Ud5D���/Ґ<Ւh@b�9u��	 �$4D�0QPC�v�8�*f�F�C��mz�M0D�Xb���NC�H��!L���8D�:D�����C;��d��E�+n��J'L+D�PI�a\<lܨ�B� v_p����'D��s�ȅb*b�ps&2'�J���#D�L	b��7&���Z
'D,��6J>D�@��l��s�a�#<����<D�`�I�s$��`�c�(Kc�<�'D���`	��mPX�����(�Z�a֌*D�8���ȕ9�H#�F��:V�<D����^�RQ�C K7�̡�=D�$��`��b�mIcd�5۞Ѫ�#/D�+��,n��k�GE>�b�	1D�,`Q�2A��:u��)(K|]c-D���eG'b�0땏QrB)��C/D� t�.^�H�2���J�6�+D��[��T-��II��~��9)�%+D��R�H�	�vm����d����(D�� :1���L�����J-]���j�"O���4gJ�g����F)f�H0��"O�䀄%�	N�"����%!��b�"O 9�P��J6�Ԡ�9� h�"O�͐���?Q4���i���:��"O�\��⓹r,@	<IAP �0"O.��FhڨV^u�@��w�L%��"O�t;䊖%���[���1c�����"O���/��P�H���I#��hw"O��`���L��_�f!��C"O$�lG#6%@̚�ƒ�Ru0}S�"OX�c���t���!��Qmd�r"O@Ź$��j�b@zĕt3T{2"ONp���*��8��%^up]��"OX$rSϚ&U ���� �u�ɪ"O��h�HÆ	�ݨ��]�Cd�%��"O2��J �6��X� �حj9J��"O�b#
_t�d�+J�n(jU"O%:%H �v^���/A�~gFQ!P"O�x�g�5����ͲPR� #"O�$��%�A=ՓSb�!M-.�bc"O������+���v!��#(�lx3"O���EX�<(T���F6uPM+�"O=ꒀإXr�`1SI]��{�"O�IR���4�����ʬ	����`"Oʘ{d�E�����U�H ��"OҔp!��" ����֟,7|j�"OV%@�B�5	�H(�Rl�7�@�"Oز��zZ����jF�E
l�b"O�p3���zM�1!��6|�Y&"O�h��T�Gez8�7e�g��5"O�iC�
>ʀ�C��$�DM�"O(LJV#�-I�:u��G�x�aw"O���8��X��Fr�����"Op4򇎛�6��Aˏ����"O,�y��S8V=���!D��P���"O�Q��A�3~�T}���1Gt�x(�"O U�UME��� �Q4��
�"O����׃up� �c�]��l���"O�쩕(H�i�z��E�ة�Q"O�P� T��#�D�ح��"O���R�9p7�a�TX�w�H��"O&m�gO�n��8��̡k���"Oб�&h��] �Ӣ�� ��D��"O����U!'��:��l�K�"O]��a�}�޽��@�"�(�S'"O}5�q@@�*`*ԅ�T�"O(�)B'��I�(� )�
�a�"O׏��Xu��C�-Ţ�I�"O�L �kJ_x=i6���Z
P�q�"OTLx�)S�(p3�,�ZT�"O��z�hJ9��H�*ǍL��0�"O����\�>�(�)[�t�P�"O�I��7u���8�Ɂ�i��%!�"O�͒cĈr�
]�w'E8g��Q�a"OL���C�sk�����	�����"O\���"V�T�UhY%�����"O2�F��BY��aW\��0+�"O�x;��_��p����itn�@w"O�p@D`��s�fpi6O1up� PG"O��r��O����ɉ�fU`�y0"O�)���'WN���$��O��D"O��:Uĉ�7��{3IǕG:n���"O�Y�a���@���?(���"O� L9�!L�-J X�g���Ta"O��ycN�FN�a󐄔�VJڍ�"O�l�o�mp|�0&��+\�@�"O�8�7Ƙ�L��*�b�.����"O`@wH�� �x�rp�Ɯ��"O�l��Oϯg]hKQ���e"OfM�#΍�AdX�0!g� ZG��4"O��0���Tm`yJD��"~M��"O\���.Qژ��$�(��ݙ�"O�M�2gM�.A&� %����U{ "Oj)��e�6v�|Cv�Ĩ֞�B"O$ds��+W-�P��@��f͙C"OhX�
ȟ_{r`p�@���2�!"O2���� L��ܨ�e�/a�V��"O��+D�sP�ٺw��i_��"OԜ�j��Uz
F��}ґ��#?!��ձ,{�qa%O�&���j�/¿�!��/&���:b�h)8�8#���!򄗎8D��*�Lׇ�9@T�F:C�!�dY��J$!�B�,j�]�K�ws!�DC,���s@cZ�+���� m'yc!�Ý6���׆��ы�(_!��bŚx���/���k\�0/!򄐖|ڜ͑��ޅP%�T��j�$m�!�A���9�2Ʉ4")��I0�!���D^ d�(>zdhX�刀�{!���I|*9�I�,bc�eb�NX~e!�$��� X���ґO!�+C�^!��C:lª`s�"=5�ѩI�?Y!��8PM*"�o$FYH�ʉ

�!�d�@tzu+"��#y!z���iȋi7!�䂣�Fȳ����=�E��8!�$îg���A��[�z�!�@j�&R%!򄎗MFd���Kצ�
��f�y#!�$k���a7*  ���խ"!�؄{���Z��U��ڵ�n!�����izEiۂ� x "ο*�!�$lh=�d���(��1��T!�	{B�cBK�G�>9�5��u�!�d;_�t"�J����,�		m�!�B��t�Ӄ\�'؆�вg��!�$@;J���Sf������4�!��zV��U�H)U�<�x d�%f�!��ߥ� �BcYg�dE*b��3K�!�$�-6*9�����E�^mJ���8�!�	�o/�����Z%Ɣ�be �"�!�̘�^��w�;2�p���o��l�!�d;��8rqL�4�j�a���0I!��L�h�y�)@��L�Տ(:Y!�dr��0��1+�:!X#��?!�:����w�̰�J ���Ĭn"!�[tݮdB&Nэ-@�pC�G�5!�ӶtT�!a�k�=�-�#Q�!�d��3>v��U�̸i�깃��� �!�D\�SP�
4�ʆX��p��a4�!��9I�@�׵9ΦqQo<�!�$����O&Ǆ�xnթR�!�D���N8��MR.%΀J� ��W"O���`��XxL1D�3�i��"O�I�te���D�B��$\����"Of1�f�"lNH�06��.�����"O�qR5ԢM�q#�O6�:��4�'	�ہOT=R����7	�;!�D#VyzP��%��LA+%(Y]�!�� ���b�UѴ1�ffȴV� �{w"O��J$�I:g?}S�/v%��""O`Z��̊W�~�Pt���PM`�"O�q{bo��"��Q�W�	:La�"O&���Ŋ3.t�с��hT���6"O�u*B��MrV ɠl(UI"Oz ��l a�ڔ.:�X[F"O|쑤�� |j��
�c��)�p�"O�ٳr��$�*�1���:^Pb"O�-���Z֚	�Ń��|ؑ�"O4t�L	{P��`���)�v1�"O��ÆO ��p��B�
�$��lp�"Oz�j��
\�P��DKՂRxD���"O"�ag�{��9��I�vu�hx"Of� �Y��(�*BH�"��0�"O��@��Y'D��=�����	"O���7�k�/�3jV� "O������V���Y�¿G����"OJ�8q�IG,iZ��Ɏ*N����"O��+Ҧ&^[|�8T�ҥ+�V��"O\���.si̤�4� !��<xV"OH5b�!��A�r�JP8�S"O(��,T=���K�"��"O�$Ka�9sp`�)���)S�@-a�"O�ةC+YQ����ON�V	JH%"OTx� NX_��@�r�t)"O����´{�-*r�	�Eb��q�"O@��e�<,4U�X(%!`G3G�!����e`�-aAC��`�!��^:l��R�6@���"�O�!�$��by
=@�����kM�c�!��K�����%�Z��3!�
!���?%k4H�� �˚�'yx&]��3�x��$�ʄ0T�{B� �t����R ��Ɉ�c���p"�m�d���J�
DH���n��͓�H"4��:O�%Q"T�H�*m��c�)�N5�ȓ*�tD�"F({� �� �
���ȓc�bH����R.詗��C�F@��ly���Ѯ�).�ppɂb�c����`�2hu���T�4PYP��'li��a%��e�R���h[V!� ^�H���2i���`�.; �[�D=St��ȓ#�,�V�]�x�t�$���RB�	�2��E�&GR|Q(��V툏?�B�ɪ+��Pf�{ب(��0��C��5B  �C#;�`��EV�4�:B�I�����S �dpD�TN�^C䉿1����mT�Xt`��s��
C�I�A#X���V�I�:h�jM�]��B�I�yz���WAзIj�H��g���B�I�&�}�M	���VJ��*LhB䉻!قƠ��m�r�r�~B�I�4�4�(��7�6���]h�C�(o㢩y�F X4P��3�+-U�C�I+Q�);�D�4 �ny���-��C�� �|y�D�� Y+G��7Cy&B䉳|´��׮]�w���ȓ{*LB�	�&D����nO�?>v�HuE��Hp�B�	�Zkb̂ S�F�*�I�4�����,?!��҅SPe1�n�o���@c�]�<�TB�5� 	��ι�x�⪌V�<	�h9x��E��2)B>0Ic&�M�<�GG�-�������/$O24�+�M�<� �2���nް`r�� ����"OF�2�_�D�ʳIW.N�f\	�"O���&#�%�Ve�$���;��IF"OH� pBO\0\�[�,S�$��D��F�O�rq)�.�/v�Jdc�H"�'�1H�W�)��(�`�W�
��!�'-���� �*&4TTk��̸ �ݨ�'�$��,ٽ\�T���	ue>�R
�'��y04č%�L��7�ž~,P(�	�'h��D�*F�R�`f� ���k
�'�z0�'��2i>(�E��H ��'�!��O7\�"���@'`	�'� ��DF�6'���Pc[y�P��'%\�'�@'RuP�v��h��'(�[wD�c����8T�Z!�@$D�k����*�aB�N�F�Z�"D�L�V�/f�"-SvE�_`��q,"�OR�b�J%���K� ��Z寙(Q��C�l��E7"L����%Rg )�ȓ\����aE8d�
�r3�
��m��$����Z�\N��� �T�GO����֭��f��@�R҆{Q���!Ir�s	4C������X�^݇ȓzy(Iy I�F��M�W��@&ft��	ӟXϓ*���&ѻp_��4�֮c��� �:��R*¯]ܪ�L�$nLXX��X��9�d-(3H��$� }<4�ȓQWEzkP�4t�]#�T�7*�I��G:fI�F��]�6Y���Ϳ#��d�ȓY[f�����./��{�Π~N��ȓؐ1��5q;&�8��%��3�� �!�M�:[�D7RV��ȓ=��s2��33�*����q-�ԅȓN�b��o|aQj o��t�$�\�<��Ӎ�� x1�g.���M�<�厓.���Y(W����fM�<��ǉf�P �rD�0:�x!�F�T�<є
�1I0�rXQ�İ�o�v�!�ę�p�f�éUfVk���+5�!�$D�$W��k���(X��c��o�!�L�9�<M(��Si�L��D3u�!�D��X�Z���坔e=\QH�'
0V�!��	��0���UV+���5G�!k�!��R>����%FƦu���Ȑ�1!�$��kV�d�	���iG�N� !�DX�:���(gKX>t�����A��OH��ڼĢ�RS�G�||ĥ!�"O<�����N�V�{GL�-7q~U �"O`���|�I���<j �:�"OzD�џi��P@%.R�<aT"O^�0�L@����!	�:�)Cw"O��
5�@' Lv�9�ə4��1�"O�%9,O�>S�Xs!(�>^�V-B"O��!���T�
�c�e��#zѡ"O2IY�VL�*���$<�,,R"O�	���^�$��ϊ%lJ�8�"O�P�7��9h��5+��F6m��C"Ov�����k��@�f[��<��$"Oޥ�LN�i><ey���� B�mk�"O��ɤDZ	5�0Fd��4
(�
"O���i�������W�μ&e6���Z�D���	&,�L8�sjH6hz�p�ȓF؜���	C�F�c`L2	ul�����k#LV�[2,�+n�
���S�? &0��M$&)>�3팇%�TLa�"On���A��n"(�#��|�P0"O�����Pj6q�!�#aĜ�Ч"O���pdË\;v �v�\�>��@�a"O��S�"]�Sh,�Y3/�@�f݀"O|����;��S�_�Zզ\��"OJ��*-���#%��X"O����S�R��S˘-eT�Q"O�X����89d��V� �b"O�	��!ߨ	B�ma���a�e���&LO�	��H�b�>$0Fנf�#�"O8�1��[�MU�6�φ@��CQ"O$��ʏ�?.D�&��H�DS�"OB�`.���`���"�<�*O�9tK��?��A &j���'�,���&4G �*�a��X�'���3��ەkZE Δ�Z xz�'IheQ���%f$Щ�&Kb�d�'6�IH�-�O}R�C7BG�I{�D�
�'�f�Q㊁�d�d�I�!k{ll�	�'��XAd�W�J����dy2��	�'�p)�1�1r�\�����3�l��
�'�n��B\�v�L�$��c���k	�'rLA
0��*s����d�d�E!I>��k j$gM��M���Y��r����������h�%kN
_����H74�t@�O��8W���@F%{�zрu�Ir���Z=5�����%�V�K3�2D����� ژi2��˿�6P�R�.D�T*a̘��D���.h����U�-D�$9��F� c�г�� P����l+D���Ŧ$;��-��\�u��ra�*D�XI�ˑV�|y'�Q{��;� ;D�X�C��ਭ��W��5%'�$<�Ox���K�1+���a#'L� 8�"Op�a@��:\����q�5	�v��r"O�x[U��h7А�EH��¡�V"O�Q�b�]2��S���K�2�"OP\�$�Īg�պ'�S�x��P��"O^��gd0V3�5k�oχP��x�"Ol=1��[bp���مM~R� d"O�$�Ь��(M1 #Ýy���"Oh���L�; ص��c��PX���3"O
�("��	q>�j���l6�鲣"O�sTcC�~G�q�����_6�]�V�'xў"~�K�5b�$]��G/}pHM�҃���y���b�)y�n�u#n���>�y2�_:xx�Д 	�!�du�  ��ybe��nБ���߶/�D�g�ò�yR�M�+����'R!��)�&�D��y�$J�=����Ҭ� I���yҠ���X
�B��B��ð���yB.��L6�����:��4�Wh��y_*~S
����T�e��@�X-�y��ѥ	����6���^VD�h&�ȓ��O��D�O�c>�+��C�Uw0H;�j	�
�D��)D�t�ذ�Bp��ɇ?n��E��i'D�,0�N�#�&][���p9��*D�9�.ݺW��܊D�P���,R#*D��f�U	pSh��͹`�nd��:D��ѡ�Q�@M�%�?:��l��`<D��+�+Y�-ຘ1�!��V�%��Ո���k��=fK^��Q�;~-��8f"O�y	�j��Sߤ1�͖>/�N���"O� 6�����@���2�ýs�M:�"O�D eW����b��C��@��*LO @���5>Ҿ��P��W$�s"O�P�o�j�H��� �q`"O��ak�|�>Is�&��@n@���I��D��C�'v�4�*�DÐj؀��ƺ4�v���,E�My�*ĉHy<A0g^�U�d��Fخ�s3M����)�^D�Ņ�!vt\[ΉB��U)#�W�Y��p����E�)2^*��7 =;h؆ȓ#���l��N�Dc���teZ��ȓfoD��F�q�3�Dџ�l%�tF{����K
��ؓt-�^] 5"����yc��t�P�𠕾j��D� Ǹ�yr�	bzec�E�t6e�B��y��H��2�j�E˦O�t�s,@��y�(̀=�@tI�h�(E|�{����y��ԥm`N�@,��A�|iȢ�3�y���$�q�U*�33
��Q�Hֆ�ybeS).R��P�Ç/L<��g��y�Q�	pDK��ֱ!����b���y�ؾK}`���k_�D�`��$M��y�Ñ�q��萅�7a�fpK���y�k>@<\�� VS���K��y��"r'�1:W%OHF�������ybD#�V�h�ֱ>� ċ��н�y"���@���a��f��nW�X��'�䄣��춹�")�.m��h�'�C�.Ǣ6J�U�*�&g�D�!�'.�|����

2���>Vq�	b��$;��=���%;���y4"N<���X�"O��ɂ-۞	��
GN
k� �"O4	��œDf���;a��Pz@"O����`�{ኍ!�(�0o�N���"O0�`O_Xь�
��Y1Qоi"�"O�EytF��[h�-H��
>,^P:$"O�x�[�P�Ia�ؠ��:�"O2�I�]��]�4f�ָb"O4�XA���l�ZA�ߛ�n �2"O�X�Am�J�p`˓~�<S���~�O�rh�Fa�,$}�,;�LV�e*��	�'y�)��H�A�Z�P���
�Ό{�'}���"�H�%�t�Z�x�
�'���������ag����
�'0h��TJ�r�p8vdϜ{vtA	�'�8R����� ��",���'�Yg�O.hr�; ��e��' �D��L�hL�w�E�@̈Ő�'���
cbҟ7�v̂g@�K3rd[�'E
�JGV�!�������&x�~M��'P0YPP-;�1��;w�v�Cϓ�OT��$�"e��e��o	�̛�"OP%QQ�0J˪hB�ހn�Z}[�"OhM�B�M#��o�<X�R"O5���*`o�I��i'~��c"O����g��A�6}�◿/���`�"O�P�Ԋ\=oS�xg�Ɂ��� d"ON��)�Qk2+\�C@d#�"O�uP�a����tE�uqg"ON��AǃP)���k�`Xbm��"O�lkҠԵ��� GսvDb)�T"O�Ր�[�%�a�`f\:M~U��"Ov�a ��3 �A��F����B"O�����T�#yA���9�L�p�"O� ���g吅��\b�cޞ:��Y��G{���9T�k`�'�.��U�b!�1�������M���q,T�K�!�$�|�r)��	�dPm{�@G5!�K�#�Z�P��O�W��3KĊ�ȓtLRԚ`K�h���C��vV��ȓ+�
��d
нZ�nLp���&W�J�ȓ.��E�U��"�H�QSO(X�Ň�	�<	6�ݚ|���D��%΁�p͎}�<A�;Xc�(iD�L"�<Y�#�x�<�hJ�[2�H�R"<�HQ�2fx�L�I�<9a@�+$(J�cC#_�j!P bGx�<%��c2|p�㜊�l�)�Ŕo�<Y ��6�DT���?j�N���BZT�<q��-$mp�2i�E�Ѳ�U\���̓+8�As`LR//׀yѬӏEʮ��D�Mw�'U��ڄFͣ&�t�ȓ����դ��0����X�v9d|E��S�c&|9��A5GI��g�M�S*�B�ɑ�̴��'K?�>�X-Q�:}�B��z=�0)�Y�m.H��KDnNrB�ɉq{tDx�o͵'���` }�B䉲�<0@GF�G#����O3^%2�Oʢ=�}�b��6�ժ@��zd.��kHF�<��LP'n���RBB�� �d��~���Γ=Z���3�P�^�Tӣ���pY�i�ȓ1�ђ���:ʂ�����"8��ȓ
�x讬4~���+��i|\���"Oj��N�!�j�ҁ�V*mh���"O YqԣG���X9@�������"Ob��,%S1�\#è�~L~�0 "O����
��1? �9V��R;P�j "O�|J5� {��Rn��H2��8�"O.�)�-ƾ/�)k�M�
$�!ж"O��yW$<\�p�%lR�c!4�$"O���ZEc��j��94��ZS"O�tB�#,d\���@��$�i��"O�\{�E�)3�E�A����*\X�"O����-c̘)��
�u�4P#r"O�X��p;�U*w)�/ �����"O��eD�TUl[�B�c/.���"O��I0'� Q�
��v�^ Z���"O��:���E���Q��Nr��Kf��-�	L̓}��h�6 ��[�d0�u��xE�ȓ*��\��"��S2���KT��@��Ɠq+8p�U��KG�8�cMc+>��
�'�h��g+�P��|:5O
�2j���'e�xp��M�� *�-c�R�'4f{w!�-e����G<1�1�	�'�t��bBg���I",E:-|Ѝ9���'\4�B��MS��9���#4D��'6�81EK(:¸�w���Q����'�����B�%��#'�OJX��'R�!zB�Ќf�<{�͕�3�:�	�'Eva����7a������F�1����''h� �S),R�9��%ƺ���'W4p���נ!���4-֡K	�'�97�J.�6؁p�IY����'��ӷ��q�.LrWņ�	b�3	��'�`R慼5��MP�ڥ+�H�҈b�	B~B�4C�XŒd���A���IX��yB�3�� ��4>�Q% ��y��AO�b�c��[�&�f�3���-�yLJΘ�����lbJ���y
� ����������b!8��m�U"Oj�!1�b��tJ�ËI{�(�T"O�!��Z%�^�
pi�2�.$@�|��'���< 4I����~\�h!'�2!�d�Z� <��(�;eV4�@����c�!�Õ�t�i���`�D�B0�>C�!�d0N�d@��c�cM($	6H\�F{!��V�;nQ[�!�65�4ȥ	-c�r2O�A�':ȲR��9b�h-kf"O$�����9���A�Mĩ/�8���"O�4A%��k���Fky�q"Ǒ+W�דLof�0�f3	` �5"O�L�&�B�e_ȉ ��?`�����"O�m��BV.��EB�D�L���q"O�-9� M��$�I�1/���`"O���A:M=$Y�&�L(v���"O(�S����Q�>�8�F��.�T�3�"O���Ğ�V��Eb�B�.T��b"O���$�^&D�m01�C�-�l(�"OrIk�\3^����F�6T��}:q"Ov�Z�J�7-"�M�&���Y��	F>�8�Fy���"�L**��]:Q�&D�� /¹R@J���ρ%e�Y��D$���O���>�r�n�	r�$����6埶�yrE�1>u%�Xw��ȉ"�J��y�JI(_�2��e+Q4�@�Ao���y��,}YhͰ��X�Z��4���y�kEF���X��ם���3o�4�yG�6Jwč���y��������hO���$�-f�b�q&�ڎ~�V�{'�	3�ў���65�6D���
�+�-�PF	�%zC䉣G3�D�r�24�`a��F�Q�(C�	o-l����1m�2�B�׳"LB�	�w� �HZ�_�B�*�aՐ] C�I�O�8���T�!�:�g�(4�B�ɭ��,�(�\�*��5�OUp�=�
Ó���,t2��M�J�� iU CMyr�'�(���|�հ㬚5g�8����yb��5�<
gDM�7����O7�yb��vh�����X�� ����y�DȄAѪ�V$6N�R��G���y��׃ �X�uM�'x���6�̥�y����VyX��t�͂�MF�yb�w�UF�4"B֜�T��;{�=Y�ZP�9rS.&�aS�-W80���
B4-����ôA��I^"y��ȓ�dI9�d��@ܦY�pdC��3$��ہC�S���)�#�C�IP4ܔɃo����!2�_�<o�C�	1�z�PԀT�%@���	3(8e��L](�Rj�*�,��2
��cz�ȓU��W�f�*���E 
����Sq̠ �'T�V�h��]`�Ȇȓ������\�@X9�m��bp�ȓW��0�ă�J��� ȉn�T���:�Nћ�OM	PẂ�n�,hxG"��6Va��a�!*�r��3�^�)�vB�	�������)�$��@�w��C�	G�����HX��T�6n�/�BB�	���d)�O�xH�KIiB�	-gkt�#藤Iy.�����?�B�	�C�P�mJ�=�q��.^�#�B�Ia�	�J��9��1��]�czNB�	�l��qcĝ8���1�[34NB�)� .�`FN� �ҕ���
�����"O�=k��*���*����8`��'�1Od0a�m�+:�$��w��>^�8��2"Oh��Dƚ,�R�s��+x�|@W"O|L{�^"|О]��՞[>I�"O�ևV�]��	�% ₌�G��[�O>�����H�6���P��!?�����'���Ab��x�T�K�:L��e�
ϓ�O��ӥ
4>vI��˕�:�&�
��|r�'!N�P��)Pa0�*8]�2�S�'V��C@.W����c�XH��9�'H��n���|±E��9����w"O�TN�5M�����37��D6"O���Ά�bm� 2&�lp����p��y�d��,ZLl̲��sSx�Y�����hO�c���Où�5��-��T��I棧<9��$;打LNdc�͖2|Ȭ)#�<B�/����H�3-�R��󨜝;.B� �x�hr��&6�����Z�c,C�I 1�� J�&V)%Q�!i���	e7C�I�[�H����[$	/�ȓ��+�B�+���´לn�IBP&�(�B�J��Aר\�4��M���5`B�	9>Q�����#	��"�Ŏ�z�B�b@�q��H)z�ђ" 
4B�I�z6^hA����Y�2��'Q{8B�I.��D�0]��{O�,P$���$?��Ip�â�;(�2 !d_E�<�t�G)BHr4(��m��� L:T�f����I!aP;Y:�,��@9D��(��X�g@���LM�|��R�6D�8	R�o�
��	�	D0���5D�t9��D,v��X���|8��d3D�0�E/�L1�1hvA�5`�j��1D���v�\:�(s�LR�:X174D���0M��'��["br[D5�Ç1D��F���0�6�C��7d*4%A�*D��)�i»���2��D���b�*D�ā��L�jpxXd�D	ۼ��1�&D��P�X�e��(����t�vE�l8D��Yv�\��Ҥñ#�4����"D��K��4u=�4C�*��-�'!D�ȢU+Y w.U#+A2l�^�X l�O��=E��lЩX��0 %��>�Z��t(�&�OZ��dU96�������b��F��8�!���9��ċ	+��'/��!�d�==BY2�֎E�ZQ�$��!�Ғ80H}�V�Cn���3� CE�'�ў�y҄@	va:�
�S�r&ZxZk���y�M�V%)#��	u��� %�F��O�#~�#��aXf%�EI�@=�a��@Bb�<���.c�����x$�]B��Rs�<q�-Z*v��<�b�\)���R���m�<�RN�/`�@�B��ɤL�����e�<���J?�0��e&�ؼ�$\j�<y�ٞV��!ǅ�W�bub��[fy�'�V��CFQ7& �S�̵�v����C�(#��[��M�(���,,�!��V.�(;�T+(�5X��.i!�\29#�"�$�H<FDr�(��g�!�D;"�$���	OS�� �@.pI!�D�3oW����� .���SUJE�,6!�Ā<��a-�4N1h��¦�~!�dE^-�6aI14��&O�A!�� x['Q�P��u�`����a�6"Ozuh%��1:VQh���� F�)�r"Ot,�aJ�	xy:9P��;� B�"Or�#W�KF��ȐMϔk4�2"Oz|�fҖJ�z�	;_�@J$"O�}��X0hP�)�O]5'Id�Q"OJ���:V���`��\�o)~<Pe"O4!�1_m����?�����"O���珁-��TA&h����A"OV���܍W�j��7l�9YH$�"O@|brf�]ò|C+�lA*�Z�"O�3��
qo>��i[`�X�"Oz=Q�N�I#<�1����0�lp�"O���2c����@WHI���m�f�'�1ObA(E�٤ye�s�,G�q�XP�R�8E{���ό`9�Ċ[�䍁��"h�!���6�"C�;� �v�Z�}!�DP�|5��yPO�*�F��D�� |!��A�6���!Y��5��ER�.k!�d��&6��e�
4��37DO	!���l0�ĦR,peƥ�cb��'[B�C�'TQ
C��Y�U+E%�$֨H��	Vy��ɼCu��S�N�xNjT㱁�7�C�Ih=jh�'ޖf��5��U��C�	�M�1j��LBSV\�3g�O�xC�I�HUZ�YAU�D76�±'��	�B�5dl8��F�.f�1S�B�$ٜB�ɤ����C��,i���©^��O�=�}�u�_O�JM��B\��) 0��z�<����	A"���k��KS�s�<Q0�]#\Y�-	\J�l���Kq�<�u�	�HdKw�@+O������p�<��`Z�A����c�� -Q"�k�<�&3��Y�R�J	.J���aTSx��Dx"��9F�����6Q�P�ʊ���hOq���y��ڀ
���Sg�R���5K"O٘��ک �Ls�M��b�N葀"ObAj��W$pj�9�Ӄ`�i�V"O���CAM�BCXlҀR
$�̨j�"Ol����G�Qjl ����`�Ȓ"O�]�7�ϗ/�-;�D�d*謠s"Od�� �	�b�$`D$7b����!LO���&�W+���K��9~� "O���%���U�Hcd�Dz�"O�Б6H%I ����%]���P"Oļ�a��:r����өf=�ԛ�'����R�=]]lUeI֓���'���r���gu&�$�؂��@�'�P�kEM�r���V���l���Q�T��'���O5f��,ÑPRQ�˄m����O ����+���K�H1f�"�h�"O�׉�w������"T�"O�u��'��MP�����2L�b��w"O��g��sS���r�×�\�Q�"O�P#�Ģm)�H��oX8ڴ��"O��Z��8�p��T	X�Hx�f"O\���,K Z�r�Lɸ.���c����hD��-�M��ih"B�Y�l��5@�	�y��N�W�:�9��=_�I�D���y��[�zN�[F)�X,��!(��y�G�1B(�\�֡��S�8$�d�O��y�lY��T(�	�`�����&��y�FF3'CR�s��*Zl&��Fʉ1�?I�'?�E2#X'?g�ɫ��j �p���� -��i<9%f<�b��\;�"OF�����8�Τ�'�Z�j�)e"O��zU�C$Jh�"JL"Rt��"Ov9��N-
�<P�����g/z�su"O�u�fnЯ'3�m�F�G�\=nP�2"OD8q�ހ`;�U���Y/Y���W"O����Ǐ��4i �<U��"OZ��6mC�-]%�Ӏ�J� ���"O~��A�-�v��N}z=i�"O��ڃ��Fj8�K�0 �a��"O�E�aK fhx��A/�L�*LY�"O|M��ɩq�H�`'�}�<�"O0�R�ґW���@bm]�C($��A"O�4��'��v�|�,��%�eP�"OlY@�h@/~]�y���I�f����"O<�s��	*U���  ���w�^�`�"O�dAm�;���
Qb�$3n�Y��"O��y���>�:6�S,��݇ȓCל�����G�����C#~���}G�`�6A�=;�hْ�i1yN��Y�h�vDP,rـ�z7�U)���ȓGW 1&g��� k@TD�����L�bgT-��$P7��N�ȓl�LT��ʹkT�p�Ղ M`��ʓu����L�P�x��B$N�D8bB�I=(eȘ��gI%:4�X3j��ȀC�T͸XA'�?	�H����M�Z�C�I�zQ�}��͞r�D�W.H,��B�$N7��5��J��K�H��.��B�I�t��<��M6&��S�J	l~B䉸p���j�!��
U�� a߻J�C�I�&�@��LF��֐#  �7�0C�	5"C���� �/�Ҍ� c�FC�ɱix( ���1O;��؂���"��B�I�r����F�
]&Z�c��V�{RXC䉿f��	� d��i}�mC�_�N��B�ɠL�"�y!  �E�s��	��B�;Q��t�Ѡ:.�%xg�̩�C��s� �$�Ыh�r�KBK�-��B�	�x���kP'¬�b%pq�a��B��g�uQ�͚��P�@�.�lB��8.a<�Cp$�=M�К�	V�`<:B�I1bd�-P�VYfq��`�7+�C�ɭ!�z��n�#9lz�2a�Ň<�C�	�Wv�D�힛EzP��E�s��B�I�@�i�U(M$q</sa�*T�����Їp��isƕ�H���"Ol�ٕ��Q7\t���I�Kn�X#�"Ox���ܟ}9��o�?��y��"O��-�"f�Z��T�4��(��"OB�0ī�)����1��xJ|�T"O*�0���o���cm�#"�8)F"OL�K�N�.�uf�k�n�c"Ox�(!��8̊<��Q�{n�܊�"O|`[FK��Gܬ��G��/$|d�U"O�m@���2O8\���/�4]ځ"O�4ٶ���s��<S����H{
"O�	�v��j|�q�E�NETi�0"O(b(L:g�
e�P R(7.\�qu"O���҇V(:�a�䮔r�Y6"O\��w��W��Q&DM���a�"OD�#-�+�h���f�:�"O�lH�h����J#�K�l�`�"O8���E*G4�18�j�3&5�;"O� P�	�����=��-F$��i�"O���MTgpd��(A�'��4�4"Oܩ��Hǻ
��Y
�HX��i"O �a���6�F�����..x�K�"O�y��O���
����rN�Q"ObA`�=��"K����)"OR#g��{|�pu@�&E�<dc#"Od]@��?:|��/ߠw���Hb"O0}��9�\!kD�I�b\��"OJ�9����� �	Ϡ]��T�"O�\��f\5z:h�Di_�Y�-�p"O�P/VFE���E��l2y�"O���nP�>� d�Ōh��G"Oh��5ǀ2x���J߳,�R���"Oꍙ4�����M���L?�!�"OXyZ%g\;��BQP����"O��y1Cݣ3"6��E��B�R"O^$A%a�D�@&τmf(�"O�4;�c��g�S4MQ�4�"O4��c�>-�u���#�thja"O��,u��j2hǎ%*��E@�yR�Ķ�>�p�E&��<h����y� �,�^�-� ��ʤ�y��Ƹ>2y�l)Nvf�Ҏ��y�<?ݢ�3��?A����nG�y�˖�]@����Ǭ!͢�cj��y�)��:��}i��}�(�gĝ�yB�U+I��p��0b�hD��&�6�y�c��P�j�&)�Pա�F��y�·�0IF�"t/��,��E��y���,�а�@
�8��M^�y�*	q�0�r#��)Z�n!� خ�y2BʔO�"�:�H��Kй�����yr�֪\b�beoȊm�Iх�8�yRʲm�[Ř�UsX	���
��yr_�5K�z4A�(z�> ��D!�y��p�R�z끿-�CK3�y�*�>��9"#�}x��qǉ��y�EF>,8�xU�V+e�9�Ԣ ��y��I�*�2̸��φ��ᄫA	�ybc�V�y��H�I&NTU�H��y�F�hJ�%
pbHq:��4&T��y�)���h�B=A���pS���y� M{X���팊<�� [��3�yrE��`��G� ���@�����y�8��D� o	I�����o��y�c̲Bm(8���=5'<���Ó�ybś�b���I�!-�&AA���yb�ˀ /F��a��+����+	��y"�>7*h�P�U[<|p�E�	�y��	f�D�A�iZ��zyA���yB�[�Z����QK�6^�������y�.] Nc�h"f��~U��ZU��y����!R��{�+�f��d���yB-�/E
U	M%)NْD�)�y�H�p�PcV���`gN>�yB�-rȵ#�ˊ}��(�u�L��y���8�Z�!.|z�r�%��y"&�=M����g�	�lʎ���Jߴ�y�+��+�K�D�:�,,q5@ϡ�y�(�9�Bq���X� �
,��+��y�͐,8���!����PDX��y��Z�\s)�F�̼bgF�4�yc�xA���+BXʨQ����y
� �%���D�pS1K#��@���4"O�� �"�!HӜ9`g�I6G�� �"Oz�%���q�1��D`��+W"O�|��)O	:Y>�)��ۉGIvQ��"O�u�R+�_x~��0�V<EF���"O��ZbF
F�T����S��.H!�"O<�;S�$U���nŝE��h�"O�i@Q�R�W�ⵀ�À�Z���"O�:�n&�*H��B�0�~X"OL� @���m��ڲl����A"O�}�aͳ4e�1����	A��"O�q3�D�fZ�hsf �$d�n���"ObUc�5;��-@��`�L�"�"O���4�FE��[�&�;�"OD)C���T���0�"��.��ų�"O�͈Q�ݏ R�[�X�{P�"O�y����M�c��M�a�j�"O>!�$KV��H��g��_���u"O�����GI���m�"%����"Ob�!�
%4��j^4Z5k�"O�\:���y�(�b�JdB�"O�$���,[g�d�TǊ�pԎ�!�"O�d!��?H���r#��{���1"Od����I�Vn1�u石1��#"O$���=O���P�o7��B�"O ���Z�3���iEU��%"O
��P ɢkq���'��q<:�e"O@z��[�Z:F� ��<�Fu1#"O�R�bۮjL,5��%T��E"O��ZBC �m,�XB^By� !B"O0�����Y���!�3(B\3�"O>p�Sj�e�u��H�)�uR"O$�
fG�'�r0�Ҩ��4�0yX�"O�j�KF]�Q����	0}à"O�̢UI�)L}��'�
�&"��"O��Jq�M6��p��%S�����"O����C��-~� ��˃p�ܵX�"O~�)���ir5G�/P�FR�"O���Iȟ{�`9�%2_{�=��"OF��"K�`Yud�t�,�p"O��)����z>�!� -v|�9p�"O.��t�͒%`
k�Ę4�b���"O=ѥ���(׊DrF�:2� Ԃ�"O ْ���8X��7��m{�-��"O,���7\���ʲ]�1"O E��N�!W�)B#��'"O���5p.�Ȓge �w;T��"OH�6G��MZ�2�Ğ�X�D�CG�x·iO�b?y��>$��|J��nY�yZr�6D����eH�B��۠�D,BBtc6�Ix���81��11Z�)�l�	ﾡ+�#3D�t���Q�]wL k��ۀn�J�:g�+D���V2!�����*Q�NAAt<D��q���'�  �#H�(��L;D��eD�3[��P���mcޭ�tG?D�(���N�S�����'���hUN>D����'3,GmCq�Q��	��<?�
�e���o�7r+�
���=ޠ���@y��C4N}��R:!&j�$ G��y��=��ڵJ�-�bT4@��y2�W�m��s��N�~NM��kR��y2�E�TB��X%�J<�.ؙ���9�yT�S� ���X�~�p������y���/lʼ��kQ ���B�IR��y
� ���`��au����0\Lr"O��AL8��Xv�Q.q#��p"OJҷ�6��E�T%� �"O~ي�#��P�V��c�/["&["O�HR��uڬ;IսY���q"OH ��N�l��xT�>��a"O:��vm�(`�a�dY.G�Dh�B"O�	s3�Ƿ~�F!q�j �("Ov�� ��W˄�{%J�	�T)��ቻSQ��S�D��a��| �GܲG3�X�ȓ4��Y��D��a�x��,:!���n]�T��ꆠ4�D���I&F��8�ȓ�����KՓZ�f��0G�%K�pM�ȓ�Fl:G�,E����!���Iu(����i�	�a�4����N-&�ּ�r�O$HPC�I�]S\ej��͚N�a���3S�L��*^����-�,t�h�Q���& p����L�'���/��9���h&�S�����	�'�����Aی�肄U3|��҃T��26�>E��'Y���0���yx�FJ�@Z~)�'��`�yR���a&���r0@O*'
�pEzR��,�ȟ���1��4�N<�e�"��Sc"O���g�hju���\2s�FmȰ�Ot��>���i��I�@ B8tڰL�@�7&4az���Ñ���Zu'z^�� �P��'
���^�qYY���#��ܹ�̖�n���ȓK��89�$ʛ*HaY�#�-����ȓ)�𤌁3��%�w�7D�hŅ�	v�'��$��P�uA :����f	b!*
�'\!�/�h�pv̟"�(
�'̮ #�P�Zn� :�"�:�'�L嘴��2$��a�����˗��L���<a�홿>�����b_�5���mB��HO�ʓ�y�)��	1�䚧���/���呔�!��
Z�m� �ȫHN��ѣ�c��VV�D��M[��s��9P�!ܚB��d�T��1�lU�"O&��l���r���C�T����IxX�4��n��[��Ĉ�j
/��9��/+D�`�eL#)J(QAe��<UZ���O��=E�$!�=I�.�j&m�y�j�B�L�.NC!��B	:�|s0BM�����+ʥp.!�D�a�$ɳ3��(3d8���(&�Du�d�OR����|�7�
 @Lf#"��'?�@�G؟`����EyC	b? �m V)D�O� ���I!�
=Z�{lt3�f��;a~⁹>�A-	���i�GՖt���B&	F̓��=Is��&13�d"DcْFL�A��F�'s�?��������SSg� �e��d+D��p�$�{q�pEɭ��(��)D��A�bK�N���X�F�-~h��j�2D��#e'ֻ5� �w���g���i3D������^	�]��tAɧ*O�U�D�5Q��`���̑�P�d"�Ş��8#�L�ta
�I��^)N�l��$��)C�DX�K�Q��Oƣ]�$��>��(;<O޽�G�7?\9���#4��&�'ў"}:ش<��Q�v��5e�&�� Ls\dц�[Uj�F�&��,��\�}D��/(�Ex��	&l~a2��C{�<�V��4�����C��Wg�j���F�PP���"�'Qўb?�)p�ɷG��i��n�Ή�D�:�T#���i�s:�	aehF%�~e� 
�!�D� �8�9Rm�']~��w�9�!��9mj�AF�����c0nQF�!�� 6X���(a�2�PA�� Y�x��C"O.鐐*\($?�)���ɕE�yI"O��yE�yɧ!�d�V�@��x��'�����L��:-��q�iJj����?��'�B]�f�N�8�k�I_�=�NU��'B֭��A3��Jǧ.�T�ٌ� ��?�nZ�L=�oO 	lIa��J�_��B��=���k+75 A�a��"?���5ڧ\[v|*���^��q��P%U@����j�j-�V�0�$T�P���`3�Ș�'sў�}Jd"I(W�z@qA E
l�� NJ�<�a�V�U<���$L?5h$Q1$�j�<��y'&k%�S�d6��!|����'R�	!T����5 ��[`�q���h�nC�	�sd*бW*�&q�t�A �%+}~c��̓��'F�'�h��B	�&
I�(��ɞ1Or��Y��HOj�a��޲a�}�EϧS2�,0"O�R��P��ȐE!Y)r!8t[��I^���	 (�<�D߬n����_!��&����כ.:F���L�_�C�ɧ*2���'D�^�Ѓ ΐ-A��C��!6�v���ǧ��т��,?��#=�
Ǔz	��
H�4Yۚ-Y����LчȓPޙ2��1�q �mF�J���o�{(<��枧Fj�,�V��7 ��s���O�<���R� /��#�U+��
��O�<1'&C��*�C�%0�>���Cu�<��A�*!��#ȶb*���h�<��D�a������3.����f�<Q�o�U���0�fe�g��`�<���4�j��� U�$�z���nM���x��e�p�ytQ낰�s��+�p>iH�8␡Z$i_�P��$�0! XK�<��IE���dc�B"9�CW�J�<�gHr���!�G�q��I�2�Jb�<�&��<BG��� ���b�nXy��B�0X���5�+Sm�Y0�*�Ho�B�I*�n���/�.7�fl#����t�B�ɪu��@r#�Tc�x��f�..٤B��9]�
�� ���D�L����B�	�(�ɱ
�H�p�x�L=-�B�ɪZvj�Cޥ�J!#c�7!��B�	3@x6��C
��(]��.M�~28C�	#b���b��=G��� �K-8&C��"M �ĥG�D;��J:G>B䉄T&Hբ�'.4�u�L_�C䉈S��B��g9��x�+�P��C䉲!�h*���0N-�pPu���-��C��)wt�A�o{����a��s�~C�	�;p�@� ���'��x�&C䉝E�0X+v�A�f"v�L�4UC�I����έv�j|{5�[�˨B�xr��pr���2L@�#�;�B䉆z�Z=S7��6A�> zAʋ��RC�	�S��͛�
b���6f��Q�C�ɓU��i΍E�!�wL�"Cr�B��J�͑7@��wK���E��'!
�	�nW�xjp�(g���<���'��t���:���f%¼�r�p�'?t�P��QV)J�(��T�sX���'�za���K�rwPݚ`,�=l�����'�hL���=AZ(8��٭kc���'�(��V�L�]XX���r=X���'�� �@�/C&���A��x[�h���� j0h������LY��ǳ	֬���"O��i�� �n��眒d���˷"O%:��Z�Sh�¶H�� �0v"Oz�"�O�����s��U���*#�'����"�)A�b�i!K�
{��Ư����y����*6��'~)�@�A:�nM�`遾-9���'9���s�	W[�LɆ+^�ar�'�(a���B�}5>ԪӇ�Qg�0��'�`����%]�P�T!R�E2 ��'@BQ�  V�IB�dгL]�3� ���'��ݓt��P
��*�7)U��'�J���\.~0J�
�gۍ�̬�	�']�DE홥�1��E� cN	��'�p�;���#�h�C������'�r�S"�Ez��ՇM�x;��	�'�(ܲ�љ9����cԺz����	�'f�]�;D�]��j�%��Ձ�'ג�ؓ.O�%���*F�23r��'�D��j�-Y�EXcd�t!8�
�'ch03D�^�=d,�Re�زº�	�'�ހ�'F�1 iU	���fl��'vM����:u�|�Q��"�����'��-�@c
�{n����H�r�F4��',�ѐ��*^qd!#�ĆsS����'����C�T&&�Nh2��Ȩ��
�'���k�X�'��;BCZ�[`�(�	�'����f�$e���`�V����:�'��}�%��I�A��0ۆ4��'3��S�iW�m�j	� g�z���'L�h�m^ 4�8;���v�z���'0A�Ыʲ|�Ʃ�ц�'nH����'��\���Ӌn|��{�Xj(��'KP�Cb��M�̩���ل&���R�'9���r�^�o�h;�eÌ+�D��'�0�u ��(�L�կъ
<��'�NH�"J��_2�[�

��'S����d� L��/��w����
�'�ثfɘS�L�A) &j�콡
�'�lH�&nIL��D�3bL�d��`a�'�r<�f矼�����-��u��'{���eQq2�X3�ʂ�i����']����Q�z�����m�L��'��Lh3�\B6�#GaQ>y����'�t C���Nb�;&+,=���'H&̹s�A$˄��#� ��\0�'��'��2,�v0�vXJ�@c�'����1�ޜ4��@&�S�y�	��'U�]�e�Ɍ��X��[�{ߤ��'����ӊT�z�4�Av�_OҘ�;�'��c �*dc��r��L�_�$D�e"O�X�f��C��଒+I(��x�"O0����9��ae$VM� "O �����[�悫r �@r"O戰DC2v�`�Ӱǚ�HN@� "O�,S�(�)P���kH�,2�"O����؟~�\�g��5����"O���n޿w���"��
��X$:d"O$y��/�-O�������Tp��"O $�`b�%j�V=����,{
}B"O��ЈV@����#��]�<x�!"O�И�H�8�
������0!��"O�yaI�1��I�o�l��d�""O�	,���wT1��e�b��1v#!�d\_��0��.�Z��K'kJ!�� 0����,|�P�1���b��8[%P��R�z�a{��Ⱥq��[#� $v:3��p>��$�l*�N���3��*�&ARbg�!fB䉔arp��" �:�V����"�� �+����ŀ,!�}2��z�S�a�`YģQ�[%x�OD@�B䉳�����¸���	7��z��4c!.]O*��a�O�q�t�GL�����ͻW�`�W��QH$��c�5���ȓv�Z��g-Cg�Ԅ�3��04Z�P'j�.�<x@���8� �c˺c��4�����3�L�`7�˘vX8�V� \Oڅ�r��O�uc@bCL�^��'L��T� ���"�K0,��zȀq5�
�0>Y#I�^�8B5�ju�(Hd�@ܓ;\0��C�L�b|��Q+B%�`�3���x= 擦ٚh�R��7�r�#j�
B�I�D�&�`��U�Nq�ԇ�b��}p�H����e��Hw0TP6��G�"b>i0�N|��V!� �Rx�����?_r��u&D�˃��� :LHŐĂ�3;�!I�Y3�t�C�ՍJ& 	��!���1s���?E�P�] 
�=6X��C�@:����I(�����Gm��2�)h��c�}U��Rg�I�$������;$|����-wÒ�i�o;O�僡��Ɓ��
͡]/��x��$�_*��(u�ؽ$xͨ��\�m�� �"]�Vޘ���ѱ�Ԡ�f�3G�x��� �$9�/����	<��\��D���%bW�L8b����aȈ&+@��ꑍ#t�+Ɗ�<��|�r������8`��.كdT�� ��i�����$c�!�$ζJ���ғøl�c�+v��h�4(	+9��mږ�n\P��l�-ig�":,�]��LFEy������%#�b��Q�ԉU��1�0=a�)Q���t�Y�\��ɂt^�А�#hL��5�K(�$@�'*]3�nV�$Y�HE��mℝ��H�vA�X��.�1��'X&�:W"��T@[���:F"��OĆt8��Z�cNNP��a_��}���D�k�D�e���`�MV�N"EcG�W�`�d��(�
P�|m�t �6pf�96N˦
�,�]7[�*ش���]w��êOwÏ2 @bTy��3{�ɘ��QG<�VC�3F�v �Sǆz=$;�c@4A��K�퇓?z��ǳijf$���W����~:8kS�A7��䍸�R�$��^�0�j�b�72�џ|[ŃR�`Dt9�Jɋ~�´+�.�4G�N�p�+	�
����&O�撁#�ITOyB��>�H�[�'8�)G�s��9@��M���.OʥsǤ�3cW8e���j��b�]9w@
�؜��/m��tX��0i*`��&�=XB�	%T��@+'��b��g��!Hz�J�5p'�ə�:|iIq  �i��l�j������~݂��3+�S�f}��I�h����'6,R,�o�&@�IQ$>��8�!B %Ø]��h�M���L�(U���l���vk�+=�>�?�A�
���C�cڮ�����R LH\��d��~IJ@��Ǩ}�8��#$���xb/�6i����A��X���w�<��_bnv�r�_�i�����Z�4	�E &f6�S2/x�x�I�F�u
�GѦ0��B�I�b�rب`�ݜQ�n��C� �J��	���!�+�>K4�X`�-���I6
�	��ђ���7%�"	[TBT�0�`����	��Œ�J��f�!d�O�
&�I�!S�[�����-�G���0�ڕ<0��$Ԝ
��e+V<IÛ4g��x���Q
(Xh�diވ2Eg�#z����,�o[�UXu���<j!�WO�Q��mV(���s�`N(xGE��$^F�t�Y�	��\'��"��������T�}ST9Z��;)i!��;^W8�5	��}E��eZ�hࡳ�RT��ى'�^?Q���O� bP.i��\*	�S
���"O�$��F[�\�����H�DX4�(��'l�튕ϐ�:��D��SNX��pdŕ�#��V`'&���ю=|O$yJ҉������%U�b!R��T�Sq_j5(��T|�9�'�V���/�R�ڥ��/�c�Ht���d��,�v�����j��~B��3;j,�Ǭ��k�L���`�<�%��m�L���K*Osb<�ŏ��a[����
�ʲ��'����O.�Rҡ�i�H9@��`�~@k�"O\ !��f�Q�ء~���E��,�s
0A��-��ɒ>?�az�>Cލ�0H� &�b���I�YI����L�.�6Q��
:U��E�ϗ�y��i�����J��'�Ɂ���y�ɜ~�"��"���UQ<���c�y��~��$�e)
�D����&
?�y�M�*-���A��߼�25��I��y2��(6�d�`Z$�psN�,�y
� �< ���<��JA�/6�ep!"O`k��JЩ���("�q`d"OhDj��Lʪ���3����"Ojm���~�-w���CAfi"O(	��Y���'�ޮm�j�9��DW6W7���(��%�ġ�pH�I���+P�ه��(��1;KђO��CYнpt��?1�%��8����`F_7����v,��L�>tGB#�~b�`�O�q��	nx��#_,]o2<Y�J��?�BB�I�D���S�۪p��jv���r��ʓn��Ac�اS�ӧ(�p�����FD*�� �V�m�8mc�"O�8�ɑ(N�5�W�TC��&O���(; � hu�,����(쨉��ߴ\��\S�#�^n��)������;6*�,)�!�NM9A�Z<´��ɴ5&�� �M�3n��c�`���?��� 5kԐq�/��H >�t@3����R�� �H�g�!�d 6[x�d-ЌO`}*�`�)W��	�B5N�U���{��S�O�J[<ԭ�Q��d���J�''�đ%痞vuA�u$ipl$ Rb.}"�?!���x���{��A3W� EK�J��\�L�3���xA�U��_&u�V����K��ج"c�l��ԛ0K��Hs���Ԑx�����/O Źv�ʀҘ'��@�D��\�Бë�yJ<��
�'�����cǊUAּ�S(7z����'8e�Q��;z�Hu�2��$�|�{�'{��+$H�*1u4��1�R��!=m�Ѐ��'5���l��U��*�/���ă�'4���'�ӻ����*�0Sz<��G*F76����'ɜ}������0�͚+:�(�����+58$�� O��ħ*B<���ѭP��u��'O2{��ȓq��h�g���$В.g���'Bd��3 ʸxF�]�OQ>�h���h$�L�w��i�r�!��+D���%'�(�����fso^�$���I� �ʌH&	�F�3�	�膅�`�0��[׎��X���$A➍ؐ��7���
�)Y0iv���� ��i��F$���U` %7N��C��-@dX�G�j�����Ӯ�F�ӆvS��b�G�6�h�6D��ZD�C�I�T�8+a��K+(u A�Ϣt��Y"��t��=��ӧ(����c��ppzM gӤV>�p"O�ÕN�6�����~@�P�j�p�$��`�(����5����4�j��S��>b�t����*f�!�č�6�����$��> A�1j��\&<e�W	O�-JP��D��%��D��k��l��=2�T�%�x�ׯ ��<ajP�{��X���Ҙu�����_A�<��S B�xpS���]r�Ix�<�%ș�K�0�!"��J�/{�<�D���X2��H�F�vf��KSp�<!2�D��hl �j^5X$d�Ir�<�-.x�DP��O� �,*���i�<�3�^�ufn�����q�l$p'��<���Z�N!�@L]�a�	!�Jx�<�7��H�����\� lRe	�`�<a��V�\5l�K���sH2 ��*^�<�DT�B�-)`C�!4��zw�G�<���l>@%brl|h]b��JB�<	!�-Q��[?�I����t�<�P�حd7(9[�'GkT�Z��J�<)��܋���1��b3����UK�<�EL��
��:gc�=&&�Q�[^�<A�L�?xxIݵu�\��FF�<��f�Awd���KB05�d5�D��B�<��h�)$����T�2���`KE�<����i�< q�����D�}�<1���,B��S��ʍ_��ͪ VU�<� �t�Ԧ-�ܘUlU)k��1�"O�q�C�ˇY܈QEHT�'� tZ"OTЬ�.Kڥҳ)	��Af�CW�<��+R~��Ȑ	�9����4a�o�<Q��ʖ(kx�bg�@W�A@B��d�<Iĩ�:' �� �)>fJ�arF�K�<��N+{ex��g�1�D�[E�NA�<	RGp��b·Df�+�M�C�<�#F�.-I�G�49)�&{�<q����F03uĚ(_j<@Y�L@}�<��Jصq����gS�S�t��6��\�<q���H�MF�#਄�3Gs�<q����L)���r$0�9'k�j�<��k	9Ĝ�R[Ph���b�`�<�b����җ�	䔐#	�^�<aG��,o`�ʳ�S�
���aCS[�<a� U5Js,D�b��@\�0"&�O�<	Q΍;yp9���12P�qV��E�<���@�S�4x�����ig�y��\}�<ys��$t4p0�H��<)��cT�<a� wP{�哫两�7���<�ga�#s��I�dǛ!h -	���x�<aR��1`).��3�@�s2`Yp���2s��A�{U����'�~hҤ�ȓD�t��չJ|,���4>���ȓ6_0E A��p#,�vN��+�ЅȓO��$g_�V� ��P�F�J�a�ȓbތ��a�<c�ʭ@T�J1渆�$Yz谐�۫<
��#�AɊU�H�����$��(�L$8��s�,��Xs<�u�L�?�}�T���N���z%����3^���(Կ
�4��ȓo0u��e13�����#!��ȓ7 �� B���p�A�'�0{V�؅ȓ7�Z�vĜ%:�p�ኆj�~��ȓe 6\�0ˋ �j<�ժ߇<(<�ȓ!����R$�)&C�d0@BY�u#��@�q��ж,;���!�֓1?�8�ȓ|�b��A����R�fݑ/�����)��h��N�FV ���ȓNV�{�'жL`x�&�� #�L(����31�Q��la��<D�LA��_�.lȂ\(y���ٖ�լm����Y�px�AHU!`� ���Z���9�ȓf��@�,	��)��͋{�8t��<,]:� 	44הQ11��m��M�F�8��K��fX!W��^���ȓ5�H����X��cJ3�ȓ^�f�i�Ǣd=�@o���,(�ȓu�~��'�O����HƾmT���La��	EF�<Ms���1�M�5�x �ȓ\"J4*�$�JĢFP�HH1��[Bq;d��x��Zb�ϳ�T�ȓ_؄�u@7sn�<)�M�*oz���I�,�yRA��᠔"!<�Ly��8��9Ѥn��H�An���ȓ,>%���C?U,���"J�f>1�ȓQ˰�B@Ī�*��ŏ�C�a�ȓE�0� w$O�:��iY�%]9�-�ȓG���$	�6-0Ե��iR�] ��ȓn�<nܰp�4���m�a��!�'B��x�� &@��%���5"T�A�'�^e�qǘn�A�N�~��5�	�'3�����8�|�"P�D�zV�<c	��� uZRdNT�P��`͈�����r"O�����#��)BÌ�����&"O�� ��Z� ��a�,��b"O��ȖK��@N�e@�a�B6��"O�K#��j���SE 4lՁ�"O~�R��ޣWw��J1��R���#�"O�����&� Tr,Y;JZ:��'"O��j�b�L�\>N��;#�'R*����t����,���Xa��/%Ƽ�`��J	��C䉗��X��+�6�x�KT%�d;�c��[���f>�i��2"�P�dބH~\q��F,%_�C�I'k8P� ��l�>Iq�N��8�ij�f��p˓)�T���L�$0�OC5{Q�	I>�x�����x���Ps���w�[��<q�O�?���@�^�~�}�p�'�0�;��]�Dfz�HE�X1$��<R
ϓEct�(�EY2"��(B�'�2���h�A���"ό��'%�L��'j\h���b�΄�M>�k�d�ָ����%���}�լr���@� �ĉ�3"O2e"ׄ
Jc(�ZE���:|�u�R%tA�\���TR�!��
^���0z����3�Е��͔)?��Ņ�	9o�H��3�O�l���}�0|*@�"U���q%�'Y�9�'H¥0~(r���1U ���Ш��,2�c�p���!#�7c�O|���d�A�l�I�0c�=jTG�O؄T
F�5��lڱ�^�%�}h蕁q�j	a�N&��?!��Ż�8zW���J"2) %�+AP�� ͣv�A��ӃR.���ź�*�A����4A����HҮ쳖�̵)FH�&��`�<�t��}�t���nK�0��JD�K@��'��	���F�	M�@�T@��y�\�ph��lN�$�,O����D����ȉ"4�3c�'�jex�"���L���d�x#�bF"!� �G.v�0i6 �w}2��U3l�����s�'z(Q��	�77P��GO��%;B�ȉ{f�-|Ԁ3)�H*���H�|�4�GO�p�y�(�B���;�4}��2����I:q�$��J�SƐ[vHO'�l�sgJ���zy��卻f���a�*fݡ��)X�bT9cNY!�����ЃcO�B7���e�2y��zO�أA��/�MBf��A�NH��^�HJl���Q�Ai�	4JՃQP�9�TP�Z3 �!R����_��Q��8m�ܽ�DE8�z�`�"<��JᾝK���WZ���"�sy�p�d�:����gE���Y� �%B|t�`(OF��S���*�
���F��������  �2%��6��uY�(��1z_Ѐ��#� $��0���@�t��C�:�R�ȯI�Z@aeJ^�f[�ij7��o(<�wj��T{0��D�[���!�7g�|�8T{�ӸIH�m��i��|'?]Ҁ�q~�_�n���g^�C�$��ubG��?QF@߆hV�P�O��3D?L<ux&�Ċ!�L�a.ڪ<I�͓a$��0<��� X+��j��Sjh2d��o�'j� �D�di*|�a�Q�y��1P� !�����`*�d�d�,�"hƆ#�!�X���X�E��PJ�Xh1Ɯ@�	?�RY¡v~�1yff�?:�@���R�'���"o�{:��e`��%;(t��K���3 �Q?Z́�^-&[\,�	�>��!��B`��Z�c�S�Ae���'�2��2�� m�����U�&���'�6��R�S\o2	Ӱ��Y�ĨĎ �Y2�uf2��X�e	H�$��I�s���! �<�6�FA�4��dÄ�����K(��/{�r�x���D�b|�a)�vX�AѠ'$�����-Ivl��r��&��,8�.:�ɽ;@����i�0���j*�Ӿ�v�����$�kf��O��C�	%5��ڕ/X.bѠѨE��@JfE�#�[��B��Z��~��s!$���
�`T�QxN8��*#D� �SfR#N&q���,Tj "�O"%�a$��[r�`�!���<��p�z)#nд��3�8|OEñ	>��zA�֫MT�p�%19��k�1?�$�
	�'	r9�'$N)x����Iu�8�Y�����?��2ɞV��1�~��bS%|��a
sO�7�����+�q�<a���1�Ȕ�&��>g��cE2F�8��K��n��c^�"~�I0U��j�F��L�����؛h�B�I*��$��(ߘ,�h����/�1[2�����'��<�B-G	J�F=�b��Y ��kS�v��i�͋�$D�1��]p
H@n��~*��[d"O�eW�L�0Zj8� ��X(J "O� $5�I�t��5�J*�i{g"Ol�k������R,T�|,��#�"O̠ZPF�FN8�a�k
h�a��"O�*�K�*S����t�U"O��/�'d��<�W�P� 
�h"O"���,�.�ޑBN��&t*�"O�l�Pb"n>�$N@^�0�x�"O����N� :z��R�Q�B��"O�HK�͓pE,�1p�I�H�ĈB��Τp`@�ZÓP������F����#A\�
ڱ��R��+V��\�kƅ�;WT����
`��X`�K�*�	�![I�i�7b��B�:PDbf�oR*���H�Ӝr�X��꘎EKz����]B�C�ɀ;� ��W�ut4��l�]L�˓^����J��^~pӧ(�T����])b�a��Ð^�����"O�$�EBE&<�ccS�u �@����B���'{����K'����L
5��c�:LQɓ[�Z��@@Z�h�#Hm��ճ�����@�s�j������<�C�$�/)�`ȺsD�>~>�?���M�:���q�.�IA���p�IY<���c��E�)!���4
���k=�����Y$"z�ɯC�D0Sہd��S�O� Qb%@W1���Z���"7$:�1�'R�I�p�LE+1B��4U��%>}B"�+*n�����{�Hݭ^Na�rlر|^�}2���x��,\�Z�	��q�Xݰ��k�)��Ŝa���i��~�� �d³Ir8� � �p<q B��$c������zL#"b!/'�U9Ջ D�x�v�ʹW<T���W 0��ݩ�C!D��a.�/?�����IG>�9�f?D���'��*Z,��ՋF���%ڃ�9�{��Q��'-��[ �I����D�ͱA*�|@�',��s`f���u{��P�:�6!*e��Wc|)���'}�y���<%���s��\��y�����i���o�8��'}IL!Z�'[�q,�8�C��tkء�ȓ���"��[�A��`c����';��'�n^`�OQ>i{wG��~[Ɣ�4*�w@&���9D�Ui�Qd���CQ�de@4��
���	"|�ް O�U�35U���ڐ%��(ڲ F�	ކ��$�"6�C�<b��! A@�bH@ʱl�=˾�3�����P�K�W� �:��	D�D΃�+�FUS0JHJⓥ �l��" Y��y�t��K�B�n���!�#dV���*�ؼʓ��y�Ҥ��?Dҧ(���9���'P*��Tz{�xP"O�47L��!��}��i� 6Uf��6,	S��S�j�����8���1j����e%� �(��#�ӳ9�!�ğ1h���b�(�2v�r��M)OD��a�,t� ���
���W�ĳ;ψ ��E�}��xR����8�<�'.E�:�b�)#��"i�x�<�����Y���QMn��4d�w�<yR��%w�e�)��y��%�k�p�<I1IY^ax�:�h�9/ּ`b�TW�<�S Ԃ%�ف:.j�Qs�RF�<Q�� �&}�l�RJR�T;>���`�}�<	�N#r�R��%��0S�x�#�y�<!c�V[|�D
w�C&jj�}I�D�y�<��F�x6D�K3eբz09�+�r�< g	����@Q�x �#m�<����+B�ܡ&Ù$ȴ#�g�o�<Q�:���(%�Q�/�f�b��e�<頪ˆ�ѐ޽A�1���Pe�<1Q�A3w�2��R	[2xW8��R��d�<�3.͝�m�uo�/8��}2�%SH�<a�	�"��l���_�Ӥ��s,�@�<�BN��4�>����ٹ,�
��^[�<�  �v�<f@�+DmQ���1 "O�Dف��<�rI�D�T�x��a@U"O�����d��h�����zt`�"O�]2��eJ^�0C��]!,�	�"O��À��G�����+"xtH "O00�ъݨ�~EF�=	4�LS�"O~��DѿЬ9i������"O��+�AS2�����F��'"O����ѤY3(`Yc��3z��Y�`"O�IUG=,4���#&�U�#�"OHX���d@=�$�1�P�W"O�T���Ks��hb� s����'L*����Q�e`5��E�hjp�BAB�RKr��׎��/<��)
�'��I�5�U�'�b������2m���'~:`���~`d1W�A�;�n 3�'О��V�R">��rs��, B���'�>|����){R��Y"JX�f%�' x�a�;/�`���K\�M;q��'�@���7_i��t�شE����'U�-qjr���q���S� ��� ^����CMk�H���nY�9����;��d�^�qÒ���=&�)�T}���/<������$�0 ֤F�x����J�{�B���<E�d�шa���
��_E�0ģ�U�r����O*@��˓T ���	�RR��B��6F~��8�.~Q!r$�>���!&�c>�%?M�%Ø�B���6�K,6>������]3�I6Y\`��1%ިT\a� E7[^�&�[�5'l�Ȱ,@:��@�A߈�1q�e ɧ�O����MI��J� �%@����O�Fꘘ���H��A�[@F�,ȶ�4E��h�=O���7|`��$�8z�Db�J�&�f1�ȓ�T�c�c�!`u�&H���̄�(��6aY:w㙈�.��ȓRd��.jv��2�̀G_���ȓ�<pZ�GJ��C#��4�9��VR����-�B�AV�6<z���6L�="�F�1MK�ـ�'в&P|�ȓR��t�cA�<܀I�0�JM-f��|p$�2W-Q�͡�� QT��ȓ_��Ď� �,1�E	��9�@�ȓuN �UJ��{�rA���Ŀs���ȓ=����VŦ�5�������B���fN�!M"f���I�J�X�ȓ4'����b�0*�;��*a!�ȓ6�JH ��}Vd���&�.P�ҡ��Uվ@2�`��a�XmKF��?9.<��ȓ���R��Ap�͘e I"� ŅȓT�#Wߡ%�`�8u)_�8��ȓp���H-'�b��,�-I���ȓ.@��G���:��SŃxW*��ȓX]k7�9�"��������3��"!�&h���k2n����P��}:hXHF�2ĉ�T6���ȓMT��go�+\lႵ��\��ȓ�	R�@@�\_�I�`�;sAd��ȓ6K�j��B?  ՂT�ݠd,
i�ȓ����ڡl��M[2�Cnb���ȓ+�h	�����3��]���ݴdغ��ȓME`�p���'������>[�	�ȓ"' @��],j���ڂd��A�����I�:�s�gE�*t���B�շ}+����m�\h�@�[Є�jq��U�pŅȓx�H�1IݡIE��3� B�g�"���'�D����B�[v]顦A�<�ЩW�jH �a��@A1F�@z�<A&�R1>x�QeI�*��  �FN�<� �񁖫��e�*C��A)b||P�"ON1 ���T��
���$��"O��"�C�38J� S�+M>L�4��"O��Z�
V�| �M��tD!�"O�8�R��Ty-T�i����"Oٙ2��']~I�K�82@���Q"O|��Bf|��
�(x)���"O��c�L"
�����ȓ*k �
�"OXhX�%��>:��B�E�p$"O|�b�O�bL( �`�=N`�"OB`��Ϗ
$3��ڲ-��k����"OZ4�5�
7��9*gF�:`���"O�Ȁ��E�0�B�#��,x~!b"OX����
H�ns5d_�V�X��"O���QJ�0��q0�@ "O�Ba���R�qcC� Ll�Ay�"O��[��b�D50��� `v (�&"OX�3�@�(�H�S#ܾ���@"O�Y��ܖ���[��ƽ:��� "O|�����L@$��0gj��T"O(�B��u��5FlI��u"O�qQ�䀆t*�H�J�~0\%��"O"li��É21�gݏ1���q"O�)S�&�+OP�e�G�ϛ@���"O`���"C3����2%��2V"O,��`�<o\,qe�<v4Js2"O���fҢJA@�9Ů�4q�d�K�"O�I�efa��Q�~:�iQfeΐd�!��7bu�2g˔a�B��Ę�9�!�d��l�D��� �DP����]!�E��l=��ھ/��AY� 3�!�$-��2Ϗ.�����Q"0�!�$I�(~(ת�602�"���>X�!�DQ69�j%�B�M*�fa���j!��,qL~�i�k�m�L kA�0f,!�G�S+�5���V0٬L!"ꂭW�!򤛩,M�=�f
�t�p]���!�
B��IX�˄�T�-����!�D�e<�a��� �P��߼1�!����(K�CAX蔩2�F��=�!���,��]D�d蒷�_�}�!�ď!c���D!��V�9#�v!�Ы|��y�b�3l��8�d���Cp!��	�Uir���nG�s��qzw+$QW!�Q���:t�O�w�XPq$ҁ!�!�dJ D��Y�����@#]�!�DUt TX��kZ3#2��!R
X9�!�ſ}آ�bd�ϰ@��}��ɡ)^!�$�%)s� {Ä��{{2*�h�6S!��Ԋ��` ��ޯjr���  Q!��L)
1�A=k楫��!A!�_>8Z|�	�!QH�I���a`!�K�./��� A�&�V��/�!�Ջ��Q�R�t���0b[�&u!�έn�8X�P/�4�(�H� �Pk!�$ۖJx�+.�d<����N!��b���3�x41����Sb!�d�G/�U(�lY;t&��#�O+cL!򄅕�İ�b�����_:>!�dT<u�mx�I�;:xTj�.2!�d
5d��+p�\~��X")�)�!��6k��`��fS<�uː�[�v~!�d��d�I���|(�AHH!���L�6���_��qt��<!�� �|��Z4V�� ��5b;l�Xc"O��p�#nBx�6�3k	��b�"Ov�[d��'������S�@	���c"O"��#,Z3+��CM���u �"O�u�Q�U55Ɖ�R���_���r�"O� £cU�(\!�c�	�9$l��"OM�ۆ'�@��`G�J�b���"O��������~�D`T"O
$���Z07�~܃��K�a}*��"O~�I$Ś7�p ��d=�p��"O�0�.�� �����W|x�6"O��ؠo�:��؈���^Q�]�"O@Y�'�y�v�ɐ$� R(��"O� * E��B#P2��ϛ"����t"O����'P� 4�gl�0�����"Ox�C@̈́,tu�q������ "O����-�)}����d�0r��	s"O����� [E��%O:wm���1"O�P�2A�I¨Di��ԋc\�:�"O�X��(<�\XrG��$Aʔ:"O��8�b����AD� '���"O�H�.(kjd�{���n�y+�"ObCNB�P��!�`҄�v"O4-2��(��4IY��J�"O�%���4���@OO�K�^��s"O���3�A�y�L��o��՘�"O
��'�p����_�w��!�"O}���:"���	�Q[r�Y�"O��ʚ3{�1�����B%	 "Or��U-�� �x*voZ�%�J�W"O���i�"�T��K).�|�v"O�$�îZ�����"a�IЌ���"O�E���)=�����Pђ�16"O�Q+@p�� �c�ˬ=о��"O��Sa��)Ϣ�e���=�ȵ�"Oz���I�EƲ����NE4� �"O������>@p^�����0A`%{s"OTY����i&
ݡu�)
)p�(�"O�h�`F^)��a	�^�l�""O��q&l�5K�X�8HB�I���Q6"O��R�^�4"�A�t���"OD�5̕�X�(�*��R1=p
i@�"O���o�7_��1��嚺PuAV"O<��q�Ga�}���Vr���"O��#Ӯ������L�9�)�t"O�ȳ%)�7+��1�fI�:���"O�`u��5L<0ѡ�
.���`�"O *��K" X�A��%"�,+$"OJ����#�h����2/P�(Z0"O���WA�
6�l#FHϸ1�ɗ"O��/K�#�h�1@���5SR"O�S�G�v���13�[83
  ��"O�2Q�U<+�a�8	��j�"O�eۂ[��F���N��9����"O�z-^�h���F�E�`��r"O����IuKx���G��-��;E"OV�gڷ^�zQSW��G����"O<���-�,-8q"E�Ȉx>i�2"O�q�C-�8=��m
�gJ�e����"OZ���$N�ll���'��1�*OȹbP�� DV<��B�3���9�'�����ҪMB�3"�&H xIB
�',�	D��*
?Q��C
�'Q�GO'�4`$,G8oY���� ���Ѡ~#z�q�����yxB"O����.x�9SӉƨ�RdzF"O�q�5n�<��É�%^}�$i�"O���]+?<�eF���G"O`P���KǄ���k��d��"OP�0��\J=�3吜nnY��"Oi�F�1u�r���c�&e��P�"OnͲ� �g�� y͔,H��a�"O줉r�N�X��f)��j��xK3"O�xP"�&}%�!�"�3���b"O�!���ߞLO|X�/��s�FU�S"O�-��A�
x5��O�}<d���"O�T�'+g%����*xڌ4nt�<��K�A��Sf�.�B�)�j�V�<�F�8�D��1aO �ڣK�T�<��d��ݓk*�hks$IM�<���q���]�2�P�b"��}�<9aJ)U�(s�W�0�:k��p�<���N�Dy`pi
PCH�Z0�Q�<�.[?2���Y���=�F����N�<Ic
A�S��`Q�ȯ0�xt��J�<����8H{J���³w����o�<rۧV��*2��D�2%C��Fn�<a6	��a�%+g�F��g�h�<Q�
��Kڬ��7�0_� �}�<I7 �SV�l���
�,\�m�s�|�<��J�`CbYhE��� ��;p)�{�<��	r��-�����u(��:3bc�<ѵ��|�t��V�Xm" �	c�<�6�G�FF�9��/a��(����H�<�'R�橘�@[�{��ic�{�<YSJ˔D}0�����7?PX!'�s�<	��"?����V&A3�g NI�<`AY9E_�	��Nşt�hH9F�<�ׅW�~��̳6�Փ|1�)�KAB�<I���&6�4i�F!E�e�j�z�<!3H�	! �`�fR�I��q�-L�<��$���(����j�0��w)NA�<ɱ�W���(9�.�m:z��ʆt�<A@��)���6lT:���0 l�o�<�`��:g�D�\�RYbу�(�d�<	U/�4 0  �P   G	  !  �  5  �&  [/  �5  �;  ;B  ~H  �N  U  ][  �a  �g  )n  lt  �z  h�   `� u�	����Zv)C�'ll\�0�Ez+⟈m��>���ɪ�l�D��'O�����o] �P4�ѠO����N��H'�tP�l��BY4��D��<L�;`f�K�'G�d��'TD
��a}��`��U�	Re��/LZ�ҷ��*=�p�!j%e��KǷ��a�"��Z��D�E�F"0� �ՑrǦl*��)U���,j��ɣV�:�3Q��#-z����4m���1��?���?��a� h�a��73��Y���4"�&���?i!�i��P���I3`�P�	ß��ɟVznX��ܔ +�)
7�Z��4�����OR���B�����/j3���?���=��a�5������T�!��ʲ��#�jO�+x�4��,���	s�'���Õ�Y�͟ ��k\:3b��`�j"��:T�'���'2�'��Y�d$?�j��k�d s�	��yz@yÁ�Rןh��4Td��%�|��'��7��Ѧ���4j���'�f0\M� ��B �#;.�B�'�f9"jU
�yY�a�`�J=Z}��h�	J���Q�����rT�˘�Mt�iȐ7�����-#N0�PZ(VU�"n�-d,e`'�32O��$^�и��A�a��$[-,T���5n�(,l��M��iE�\*�D�&� �pe��I��Y�W��!|��`2�͍W�6������4R�b0ْC�+R�M�j��:�� �ܷ$�>�	&��U\�0 �i�� �}K��B�@� �еi847-æɠ Oe�FÃ�������[2��*g�҉0-f�%�Kɒ��ٴr�Q:eO��S:�����2w��Y�����',��zP�%>*��iri]�W
0�9G�'��O���>���N���>m@#®��!�0G�L�+�!���]�XL�TmЦx��zW�ǂ"O��g�
-���ЀJ�K��Y�"O<-�AH�E����Pg��2p2�"O2(+'R~t(��Œ�!�Pl�"O8���C[y(����k�8!br�	�qW��~���
�,�F��GH�-p�I��
e�<q�K�&3���cE�>4�T�(_a�<���E`h���E��(�Hr�<A�G1v�V��B�b��HSl�<aug?bf���ȏ@P"���Vk�<y�*��olZ�9'ṇ�N�� a��$1I*�S�Ov�T{%o�Q&���/q��=#�"O���p��1)\M���:M��q�$"O�����0�J��D���q�F"O<Hc��H�0���P�R�t;�"O���g*H�VDÕi�f���!"O��ƬWt���g[i���Z��*��(�O|��o��.���aDۦ[�z���"O��&� �l��A��&�Ԃg"O�TY��K3spЄ��Ϊ��|�T"O�I��]v�X�ϐ)w����"O�9��j��o�8��V
�p� �'b���Mvӈ�d��YI�#B
$�2UÒ/Z� ���Qy��'���'WB<� ��/��ɇ��! �\���3����'  =�K�Ɋ6Qxax"%;}ԜpB��1tVv�� �'�����@�O�"��DKY�u�*�	Ó���ɱ�M�]����4x�3A�$@e(�QiOےE�/OJ�!�)�'��P���!3(5�-?;e�������?!VVT7�8�iC$%�D@:@����&�:4BO�:�b>����$j� ]����Ļ+��"��IJ�<��k��c� 3Bв&�l0�F_�<	'jE�|���!�/&! ����\�<� X9Q�r��k��F�N����@_�<qү̎Qt�Ub��4p��t��]�<Yg���1�c�`R7*��-��!F៴㔎/�S�O�]
`OcR��, �*&��S"O,tQ�Y���w�L�a��)"O����ɚ�C��YV��;.��!"O��p�-D� H���ǂ��.�Y�"O�h�G��c�6yF��<+����&O%�_�m�E�_ ��l�S%��\��>O�����As���^�_�.y�D<s��1�tOr<�GB_;1k�EІ�+�%�<A!�_:1m�AP���-���cAb	�5�0Չ!�'x����}�䍱T)�!oָ5Ό�y~!�$H�j�N���C���}�`!#f�X�ɰ�MKN>y��ەb��ӟpC��G% ༕k�Ă�0��ݸATҟ�I[�,���ɟ��'(�T���F��d	�� ّG���� D��PC�H(X�#���N9p%@�)���lH�q�V&̻/�P�Ո]4j�Q��g˿H	)C� �M��+0ғ_����I���'�|��H�^�Y������K>����QA�� ���N�4!��ɍ�?1B�T��yY�h�/",N�	��Y����'�Е)��'�"�'��7�!�I�0�"��)ɲ41�U�g5�T�I�@X_$҈Ct/U� ����"&1~�'��	��1.*m��9B�BP/�p��I�ETV�X�B�z�Z�Х ��-��Ŭ�:�� (A�N�KȜ���&FƬ��d���!a��O���>ڧ�y�-&��ѡ"�?�vH�g4�y��{^m���5��-���Q���O�F���V6vs�k7D�_�d�A�5�?i��?i����X�	H��?)���?	��yw�ɆyV�j�Q;T9]��"C� ��L����a*eJV �8
@�4r����|���J32�C2�ۋ*�M`S�2 �l�'�"d�m�b��0�:�{����i���'xȥFP8	�d�S���u�`������G��b�'�ў��
ۋHr�)�I����L�h�V�<��?���Їi�v(<mR_Vy¬ ��|R����ę�6s�$���ֲB����	�"*��#��P(J���O��d�O����O���c>�ZR$�� ����N31�j� a��;�Jdy�l�5$�rpmR* E�  /-��Aԋ�2]�FH���K�>�!׬O�s�X���Y�3^����i�BeDzbJC�c�T,hUCˬb4S�ME>?�E����?����>�~�d�₪)�d��C��u.��ȓ8��\[G�7�PY�����%���ڴ�?�2�ݓ���Y�W���7�
K�x� ���y�HP:|4�d!��B.e�g)�%�ybA�������ˤ4P��7��*�y��) �����19�k�"�-�ybb�v���[�1�v8iFޝ�y�B,��!��. ɡu"�!�hO�xR��S� ��$���'.�L�[�� 0C��0(��d�V�Ҩf�����B�I�+WlΧX+%��CX
�JT�V�<��bT�u@E��W�W��b��[U�<�#�P/s0LJ�� ��bG�
v�<9��(Y*Px&D�(i'�i��L���peJ=�S�OثD�M��a�Yj)<��Ŧ�v�<��펎;��+�W�7H8���g�<Q�(�%@�) K�!9:��ӰFn�<Qtkޙ��)�l��\��r�mj�<�Tg��J���.?�&t
#E�c�<�ꊥD�8 *ƥ�k� ���+�`y�G�(�p>���ΦSd���#�3GM��Kf�<�@C3A�h  -L�&���V�<�'ギQ2�=;���%���I�I�<���%^��t�d��K��IuB�A�<���؜g��)����*e��+F|x��bĹ�0T�Z�4h�Ałf�@R6�=D����?*7�eZ��AoM�d#Ŏ?D���ぎ7�� s��@��`�Pm>D�x��S�>�d��eޒ?Mn�H7D��#�셢Xp���T��˖�x#k6D�\�ʞ�;jV*ԊM$t������6�$��|E�o
	M��<P�@�-X��H�$A��y�A�/N��T�s��0[�ҕ)ٸ�y�@����L�P�A�@6P�*Ea�y�]cH�{Ĥ1H_|���[��y�6��D�ç��B�f�:�,W��y�_�E�@)��!˪'����B ���?���Km�����p��	7h�@�kM�IL�ȹ�?D�d�.��p!���>Ԏ�!��?D�T��EUP�P�V8n�8�i=D�����9�=!f��CPP���;D�ܫ2"�GNnE�e$�+V�z���<D���`R�W�v���J7\:T�j'�<!"�Ud8���A��V_H�R¬�6}�>�RB8D�� 1�G&I��(5
\-����"O�H������D0��N;~��u8"O�]0i !ܺ\A�K41p �#�"O8QK,s��q�@ ]Rpѷ�'���*�'�4���ʜP�J����F��!��'����A�'��p��-@��,�'L�a[W�ɰv��-��L�(,�
�'p�����RG�%(wh��L��ĸ	�'�D��Nd�p�RG(��x���'�R�@$�U(��5 ���h��D9{FQ?�� �>� ����m�84��F3T�LٲAZT��rV�e*�]3"O�3 ��%5�&���Ɲ
��|K1"O.�r�&<\�`���/��a�ʀK�"O��ⴊ��PY夊�6��91"O�m�gaѕ8�}Y��_�M�>�Yv�'��ҏ��;���S���VuT����#cȅ�'Rӥ�S�9�<̙�:)Z@��F�
-1�b�Y���@K>.�$��F�����e�qy8�0P��#|�����y��ԋ�L�PC�	�J ��ȓk�x1�B_� ����%n� �=�'��m��2y¦劗�~�Xs��L|�ȓk�F8�!ډ��p�W6COX��"�^A�Fܮ3���w��3D�̄ȓ
l¥�E
����e�"��K�vh��m���E� S�@�U�1��1��ɬNx8�G:P� �ʇ3f��0��%0L��B�	��x��P����*��G7HC䉇J����5�8v:e�4��8] $C�I��PֆH�&rތ	g��n�C�I�C=L�dcX�\�l
�.B�ɹ9Jtx0���]Q<�C��{;��=��Qm�O��ۖM��2O��� T'%@�+���� TJ'�єh00�ɒ׼y�!�$\�.�*������Y1��W�w�!��YHPH�OB�"���[7���!�Y;K�P԰��_�I+��$fR�zs!�dW�Q��x9`i��*u �%��7\r�U(�O?�*gmM�E� ��B�(5�����x�<a�(��;���ϟ$�4Ad�CK�<�c/�"�ɧH�+Qօ(��X{�<I��ыV�z�ys� f�>���u�<I�@�	�k�S>��ѐ�RG�<A�i���)�J�6@�҅Xg�Dy"H��p>a��@�@|�����Ը`j�����B�<�� &x�V��R���f�ja3�UB�<!�e�1	G�թ@�/PKB� ��A�<y��Iv�x%`ȧJ��p��t�<��JZ�m��,���Ԣ9r1*ƏZwx���1`����'�	s �Iӊ|��)sR�?D���	�c�F�P��˾RĞ��� D�l��D)v�hX�I�$������>D�d1£Ãv�n�����S ~�D>D��a�	����Z��� z��v�:D�4�"a�7w��u���-^��� �7ړ!2P�G�4��=���x�E��JfV�Cw��;�y"���G��X�W���ID%�f�R��y�F��z�ա�dE�4�Ձ���yB��
%�Hb�/�X��`���y�]�'^�52��PX̤qw� �y�!�#�������0V╺6�2�?�u��C�����hծI�,��h�H0lp[2�0D�lC�K�r�4���I�e�y���0D�� �<��IR
}r�@増�z�~	w"O๢��+�t��vK�9��i�"O�y��#�Mh<Lq�ʉ�m�` �0"O�����# �i��wph r\�p{W !�O8��An	N.
-��(�W]�8��"O�T���u�`���W��\�D"O��� 'D�aj9��m
7"O^��ra����eh�Y��d{$"O�v�/�����ą���˥�'Eld0�'�H�S�N�*��e���V���x�'��`���L,nd�1�f����k�'�� FE��T��2�.��yrF))������G�Q����DҬ�y�� v����GH�CJܼ�S��y (dTD]��f[�f� �22�P3�hO*�s��S#l��򡚍��Ѐ�^��C��.	1�(1C-٧\R��2)��O��C�I��C�\6���q��7i C䉾w�p��Ǘ���`��}lBB�:/6ѻn�	�~|8��=W�&B�I	�����H֓[ގ��@X�Hz��D�Cp�"~*�E��e`CE `^�l�M��yBB�b��a�0΀�Z3��34�_��y�+�l�pu��#�L$"�1#َ�yB��;@��Z.�>���8bݦ�Py��6~m0�I�`�#A�X�:��N�<���\��0�J�ƨ��Yr��HTy��֨�p>��E�pX��Ũy�4�
ǯ�R�<1"'��hR����J�!=��B���Q�<	��Yw�"�Sb��4��a�kQN�<A�ʚ�)|�=��L��hPP��~�<��k�1~�U�2��;|Ϫ%�B,Fux��"�ù���D��+����eÛ�f�4`��6D�� �W�2���Ӄ0ZDx�1D������^�",��lI6s�慺tE/D����-׌Ed��R�e�v��!"D�	�U�	��d���?+,Dr�5D�L���̍va���iøE`�P[�K1ړ:��E�t��:u��e��E�%�v�Xe�
�y2��,=�f`�3��k�|��bF�"�y"��bQ�젱�L�f�*4Q��R�yRKmɖY��<bg܅f��y�'^�N05�$/��)fɋ��yB,@0r��ҷ6V�@�H��?�� �T������q! v����0��=�m�,)D��c��~�8�@�&Q�#j�1�'�(D�d#񢄭vp1 ���"E�P��%�'D��B�o�I}x5�d�@8�1���'D�,�ť	Ԧ��Pe�#la�%CTD%D�\84�����D�]5�T����<�@��~8�x�s�՞"<eQsF�b��\Ӵ�!D�|�#��.3ژ�"
E/���W�5D�D@QOxe��1�%  �E�7�y⣂�;".���N�4��8�$��yr�^�xi,4*p�\�C�&4GS���>�è�Q?��D-�>i�F��X�N|�6k�a�<)��I�fq�͐~��騅�NV�<��#�/K�Z��v`�������X�<�5n�c��� ��w���a�JR�<���t�!bI^
����t�@M�<A��*L����Aۚi�	P�,ZB�'�.�����)<:��A�_*d��
�@իX�!��@+L��a?.���@��J)�Xɂ"Of@Qo4NH1��Z'ttq�1"O� �Ŋ�cMr���n�o�4���"O}ц�ޜm�� ���TM��"O��)�n+<�|�(�n�=5��Yh��'(L9���::W&������8J�H��Ċ]��ȓ�H	#"#�%OL�\����QE��ȓ�8���B��)5�Ms���<x� ��h
�h�� �Z�d�0���>v"�ȓ<ƹ��I:;��Ie���/��8��͆� �ٕin�aBԍ�1|�|�'�XD�J�~�JWG'p ��B�9o�dA�ȓ!N�8��Qe�� 8ӣL�92��bqx�z�.�;�\m9% ̔�v�ȓ<�f$� !�W 	���3����9D\�B�݁g;Hi�����Q��I�mLN�	*����"�:� �r����s�C�I�lX �N��P�2az��<7<C�I�~�e�0ꊝp�0��5Z:(C䉍;��`����F1�q��9��B�	!юm�QK�%��r��K�
C�=E\*�{�[x�u1i^�+�B�=��h�O؆-Y�,���ױ~�"�(	�'>����m^9J�TY� �&t�&�i�'��!Ȋ�;�r�x�"D?>:
� �'�h|��B�a
���μj�D���'E�l���Դ��3��-2^=�'�݂Wă|8ڝ)���4"���8�Gx��	޹(��۱8�ā�ႃ<��C��p��+J'J����.«I�~C�	�F��{�eIk�<���jA�t�.B䉣c]<�ȣ 
ua���A/o[B�	�1H�:#�C�LVƠ	򯄩T?�C�	�`֔)�oC��LA�_��ZP�=�O�<�bA�����O瓅vg�`�1��B@�0F�ȭ`����e"��ON�d�A^1 5��RG�Q� 	�`o���r�ƀsD�с.��%Zu�D+j�#>��ȗ�G�ȅ��+tǼ!QF��-�ug`�Nh!Ap��/��EGD�O��Ez�'�?)�ΘOϦ`UZ�N�4��'�1p�0�)Od���-� �j݃�֩:MѦ?,�}⢮<�㑕=�jjg@\#Wrt���fCByA�.`�R�'\P>��@HW͟��	�de�d�Ў��ufهȖ��I�dy�IQ��cG�1CJԥ:�����ן�b>�!�'�9�(��� C�Q0�"@z�����_�v�ɑ��kx �����؊�$�ϝb�!��텚2��a�W%E+�y�."�?�������$��p��f�
8d�)��5;��P�4D����@�U�)���95.ړG��?@�"Y�a�~�����*�N��G֟(�Iߟ�a3�P�t�!�I͟<�	ݟ�S֟��Be�s�N4A��!m�ƍ�Ч_�8�u	l
z�����n�=]j!�O��O.���Z׎�ؗK�X}v�����t��!fkߗGն܋$��".������1�x®S	��Ţ�'˪S���A��3��d��U���'�ў(ϓmҖp8f'�z����R�'9�8�ȓR#&�`C�h$�m��J�%��Sןh��4� �d�<�E��}*r�4$�!Y��P��KˈR <Y
��i�2�'0B[�b>��O"W2���تo���sU�p�hC�,	)������<�CC�gT���B��xQ���>b�ؚ��ؕ2;�%P'O���<���ܟ�Hӆ��V�P��˜3C�u�F���D{B�	'VZ\���P��ĺ1�R�y?�C��A�yynQ(yz�����.OA��:^�V�'��ɢ^�������C���y�+ʡRę�VQ'|1���L�Iោ@"+M/6 �qJ�FG��{��|J�DH�q Ԑ
��>�����F�'9Nؠ�ȉ�e���"5��S3*R��@���ױz�#>-lT8�	Ɵ��|���!0H�f!�2 ��q�q��xy�'�B��G�<BX�"�V�����)e��DpLd�t'��m�����J1ê<����?i�����|���?1"D�"% *MB5�Ʌ�tB#/ӡ�?�E߹`�B�0�M����T򧈟�����16��Cp�>.���(�=O>����'X`�p��"�|�z7؁2Ͳ0:䝊`� �^���gYV��O��S�q~
� 
Ii'��vt�&��!k�x��"O p��'/c"\�w-���퉏�ȟ��ᤫ�({�
����MS��?Y���?�o��j�D���?)��?��'�?!���v'D-�%N٩u���P�Rb���Dԏj�JM��C�"�j͟d�8�,��[  QIf�0Z֮ 2JޫW��e�E%c��e�0�.�'�M�J;�D",y  �sQ�@��c�J�	�8�����O��=��'k�}B`@�#���
��ԑs����'����RX���KT�}�$���F���S�4�'Il���#T�b��A�Q �ȶ��@LB�'K�'J�)������"D�=�â\�ᱬA�leJ}A��;I:��ϓD
��j��P�E�@-��o� �̤0��M�E��\k7������8�F����	�I0����E�rZ�z�nK���Ie�'���p�H�>��]����IpT ��:D��+���:N���ȲiN�vMX@8pi�<E�irRS�,��g����i�O8� 8qD�ق:�:a���"<Y��D�3(���OJ���� B����(G�*���<+����ǀ�>@�S�*����">���YS~>���!O�J#����F�?�R)Ɯz͐� �჎G�s�d(�P) ��I�Ms���$H��f���J*�6h��@0���O���� f���"P	���j�MF,)0�}R��<Yv�S�4`}+����+���&�Wy��'��ꓘ�Ϙ'�N���':� !�cE�UB �Ó�hO����3r*�U±,_�m���r�DB���'江n��'��%-���׊�:�D(����!�'�@�L���<aV�]9r�q��ʑv�le�%�ݫ� ��O|��O:Ł6�>�����S.�j��$P�T1V���D��F%:�Oj����h��䀁]�N<y�%� o,Hg���y���u�> �>)��]i�s���ȬZq�� 8F���&��%�?�eg�N���K��?�2Ĉ�9Xc�����ʝ]�T��_���	8\b �'��'�.1@M�<۴e\|��,�BE[Ĩ�F��vy�����ɋ�ȟ�t���ʘF�p�;QK�:��H��l?a6v�T>�-W��?݄����A >�x\�A�_�za��Km�����G�~x�$�O��C0Oxb>����Ob��(`��EE��0Z�D�O��x�'+�,��O�s��"���B�KղL�u�ed�.s\����O^s������G/�`@�i>C�r��ozRI�-��Q��!��!��R��l�'��	F�)Γ�?QuĒ�=d<�:s�(�����(�;|��I۟��'�ў�	:�S�/^�L�p��(���dy��'��0�C4o��[���?[�=�ȓh�0��c|V|<�C�v*��<N��c�C6c6X�FO�Q'~4��R7|1�t�8e�$�9�������ȓa:�,��'�D��k^�S6*	�ȓ	8��`$bӀ}�<aw�}�pC�	-zx ���Z�E7� ���X�O1�C�I>B��A�@b�h}B(yShj�RC�Y'�@�JCVy ��`UU�C�	�3,Z!��&ڬsE*|`p��'dlbC��7p��a�G�ۀ�]/66C䉽2�PuKa� >�!�ӯ^cW��ЛQl�<xbڅ�&B�*s��&�ў�c�'_-G��4P���G�4�� L�@թJ�$L�����CG�=a�)k�R�Q��̩so�	Z���<4�RV�G�4�%9�ߣ,��a�`ꄧt��*c[���M*���͖����B^�(Ҋ���DŉK>�w9Yu`�eM�{����E��v�<�&�M*w�"T��#k���$^�C�I�x<��C�K� Y�#+ʎ=ҘC�I�kd ��c��`�����oI�3�~C䉚B2���YcF\�xc�pQC�	�oװ�8Cl�1v@-�%h�Q��C�I�<�Hi�IǗq�h�P�"��I�C�ِL����$�:)�a� X|.B�I �d��ۿL�@�X��*�B�%J�&�Cu��f ���L۲e, B�	"97�s�]N� 0r���C�	�&�Ρ��k#Z3���r�ۊ'�zC������s=@$Z �)3`�C�)� �X�a/��@L��J[r��y�"O���2�R�(��������Ez,�r"OH)*q%4HX��V cb]��"OlŲ�)�8��@B��;ybz �f"OD�H4,R�H��+! ŗ%��m20"O���!�	?/�Ȱ��:
�F�T"O��k���d����g��A"O.�J#̔'�pP�ǥ/��r"OF��s,��;}nP1�&C�2���@�"O"�@`�D��[2f9�� �"Of�`��Çk�"��֨)�R��"O��T�K+!� ���<0��H+5"O�Ay���s�xY��@�e�
��@"O<C��S�o~:L��M�!��m��"O��j�Ə;~��(�aO�0H��1�"O�����Il��R�nȃp��0��"O��H���5�4Ⱥ��8?�+	Gi�<��ҏ4]P\[q�½�FB؇�!�$
�cx\C�	{�k�~s ���"On��O\q��`Q:����
�'� �2��3-���j�1B���'vŹpƐc���w�C70`�"
�'@
�����J�~�b�	 -):�E��'%&| �aI?vF�	R�HD�	X�
�'�Ȍ�G`��^�����Ĉ8n�4���'PXᐉ�-���� 'id�:�'zF�����#It��@�ޜZJ�]��'3\�ݤY)�E��&ܵK���'D Y�$�2ZH��! �$<�@5*�'r�	����,E��4�� 76��x�'��d�֫8p�֨��� +0��i�	�'(V��@�""���f�"�.!��'f}���	T�(��n݃�^X�	�'�x18���G�jE������p��'G�c&��p�:�Pi��"�%k�'�fd�`��Da�öE��	x�'J�\ �k������A\7n���[
�'J0Y��*&�<R�슫Z��	�	�'��%Q�n�)��${�n��Mx8�*	�'�f���
M�8,��I(L�
�'"f|��N�]՞l �k�o��lc
�'1��"��9G�����d��a�\��'�����P�|x��P�� W	�[�'�Ԛ�� }��=J K�� ���'ʎ�2ǭ�=������,<p�)�'$�X)Q��6��8;��V�X���'�Uj�&�[�(��c!79���

�'YL��$�>Jx|!#��*�5�	�'R��[D��C��<#�cN�$D���
�'�a��ٳ7Gv*��G"w�Z�'�)��';P��3������	�	�'ٮ����=�Z!b���
5���
�'�(UN�n�^H���>X
�Z�'ed��$A�$�&��2�ѶI�!i�'_�Q۵fǗH�*a�R��	Q��@�';��)�@θA�``��$>D@`��'�N��q�F�n�z-s��:c�h{�'I(�Z5���Id.�+�O�6h)�z�'�:{�lg^�2P�a3r��'l��s�ؚ7T��B@
Ͼ*��l�	�'=�}�A��p���喉��:�'��zv��V	J`�ƌĀ\��'q�5Q�l��Z�@&��Wh��';da0��8�T����T������ �26���fș�䓀I0�Q�u"O
���=:��p`Մ6,Z1YV"O~$+�B;.:55��&��z�"O��� �	�����U%I�M�%"O� �
�5��t׭�K|���"OE���
 �srN-�
ȹ�"O&�����m�j��@N��v��4�1"O��j԰�@%:ס/�"E�1�I�<)�A#6\�5A�ҶO���yU*}�<a)�08渀�K��P2*�aq�`�<!��@3&��A���P���3�^�<�Pn�t����3� 8�q�\�<��8�Q�n�I��x�%!T��Bc@ҟ��DI��
$,� 03J8D�Q�j��7f��a�ۇO�\�)Pk*D���mF��f+�/o�XԻ@&,D�����M	T�Z�O|dQCE.D�08E�����T��2xLF�L*D��Sw�GG�@A@��6T�ԯ<D���@�]-\�!G�X�+s��9�%9D� iQ&�a	�gV�%���S�f+D�`2�N�	NiF�T(�扸��&D�Dj�%�#\]�{��P&0���B��$D��Cq�8W��ӵ	ЕOi�lSF� D��a��*j��V-�`ec)D�������1�~��fM�R���4�,D�,�6�*-1�X1LM�__z�S�%D�<�׮R�&� ̓l[� :G�(D���D��E�X�{fl
';~6Ȉ�3D�� ���#�;&�j@r��4D���E�_��;��8,8,�ZQ	 D�����6a$��aW�A2���b�D?D�ZѠX�'p�qjR� =L�IpQ�<D���A-�:�Y�0�+|@��!ac9D��nN�A7���U%ُ�f�Ӊ)D�x
�͎�!3��3�Nn�!�w%D�4�ӊ
`P�|Y�j5D���3�r�k7̓�M4h��C�.D�zA�Q':�d5��fR�
B!q +.D��ZC��1a��D�#T]23"D���,ޣ
��R䊀mA���w�%D�8����X����w&Ho��$��l%D��� ���+3&C��t�1D��4�D^�4]s�AݱT�f�`�",D��j��3[�����""S�-@U�*D��`�m�&����O2`I�]"e�4D�(a�
��5�1*�/@�f����D�$D��(�"��(��B#j4~��W�!D�4�$�Ɇ=������(R�@rwM*D��QQ�@?��1uG�!�%Ӆo-D���`�\�'��-���K�L���d�)D��C7h��&-f������t�A��(D�\�U���S���	��C7Dn)�'D��:�C͘~(n�ڡ�L�68����(D��Bd��>�9Q��H�>>œ�+D�8���H>G��[����8њ�)D���f�܎IT�1�
R�H'D�ؘg�GF0�S2�
41����&D���D�y�jP�U�p�扉��0D���Hu��[eL��S���S2D���׆��-TS��0;^��J�+1D��yL�P��%+$D݀��u3��1D��r NAI�fx��.�whxIb �;D�X bb�!
����Q��W�2Cu@:D�� ���Ե�d��9t2��t"O 9���'J����O�BQX��"O�:�Ƅ�1�Z��Ɂ�zH~hR�"Oވ��ԅQ�����";B�r�"O�����\��U(�F�-)�ᨠ"O���b��n��s������д"OL�bmC*y��܃$X��v8�e"Ovi돎"�yҴ�4R��Ljv"OX���ݸT�|) ���,y8@a�"O�P���&9�t		0�_"1���"O�k��eo���⏌�5|�,��"O�x�NȔ[y��� �eh|%�Q"O�t#NA=%���G�~�^�q�"O�$������(�m�%����D"Ob�[��s���
2�d �C"O,�6*�3-�i�v�'m�ƭu"O�X{0�V<}ስ/�Z�r���"O���۞8�b]���%�(�"ODz��L 0b(�U۠%��s"O�1�`�$�}Cp��}�"�(�"O&��a$��q����F�U|���YF"O:ɺ�I=b}Mɕ�/��	j&"OH�����H�IL�p�X�P�"Oܤ	b��1T~܁�2oU2h�i�T"O�3���3�`�p&)�6�2!a�"O�)ңp���&Ǐ�xX�9�"OJ�K���46�-XtK��j��X�!"O��P�[!A0��dk,���"O�!�3C7E�B�C
H/�ֽ8�"O)v��PԦ������K5"O,!Z#뎯gizL0�I�L
Xɰ�"ON�
��>쁻	_�t��W"O8�cH"Q����&S�wTUiw"O�}��*U�8����ӫ �3�zYs�"O�r"oM� Gd$թ\d<n0��"O�0h�M%7�N��F�'f�4�yG"O���%!A�=d
�Qc��'G���S�"O���l[�D�Z�A��Y��"O<D� I�3�$��@��[����S"Opyq��:S��5*�/]*xpD�T"O4�s�K�3��\)7�(f�	@"O��F�[�w� ��BJ>,ZN��"OD���΍[>8�����8b���"O� S��e[r�Ca
J���aQ"O!ia�ש{�Ό�Aҋ���"O`쪳,�^�He��ΐ|wx({�"OE���6�+e��cN8��"O�嚁a�����&�./4�4J�"O �ВlIr�m[p�ǟ3$q��"O(18�
�=��U�dƞ� �"O�Q�c��Va�p��C�_���P"O�X7Ɂ�U��1f/�����"O\��B�S� $е�?Uߐ�T"O$A�$�5t+�xY���=���BP"O��Y�'F� �&�U� ��ոd"O���9ټmE��D�Yْ"O����m�\y� 3�PI[�x������3���t�T�N������	��'4ꝰ#�)�P%��'D>
E����'\��񣪃w�x�DS�l�J`��'��t��D�,?R-p ,C?Y�^,a�'�,dB���2>�!���N�z��'K�qz�&�@�0��"	-B7*u��'��Y���ӒmN#�ez��'�����ŝ;:�6d���L��vL���� �˴,Y�d���7K�K�2�23"O�jdK̲Y��-�����W�dy@�"O��9��;� �4fԲm�R���"O���dAM+@��U���q�L-��"Or��/B6j>X8GX���	{�"O�8�R��Y͘e��Vb�L�V"O:L���
^:nAzЪىLV�"O�RS�Q�H{�������"Ox�CNޕa���b�R���"O2��viٛ;E��y0 ݛ.a8��A"O�=��a�k���b$�,Pr��d"O0=2!c�(}��I�˖:9Ѝ*�"O�y�bC�=��8�"J�m��D�"O���ՃˊI-bL�S��N� H�"O��R��@|�8�#f��V}3�"O
�� �ŝ3%�h�T+�G�L@k�"Ot(�� :X�H#�ܹj�H|8�"O�M��"w���T��%D�̂�BA:�Tl�+��4 �#D�<)���r)ؙD,�;"�� �RD;D�l��eQ:<����H91l�蚣D9D�����^	bb��3��^��Sf!D�c��G>�����f޷QҪĠT#"D��s�ķ@��l�S��$�n�G�!D�\��mB$#�`q�A��m�Di
�  D���F�t�Y窀�Z�<Qs�m/D��`6�d������#_t�%P�/D����o?��f=I��сD�7D����
�V+"h��"�C�ֵ�t;D��{�&�/TD�DI���tв�Zeb&D�p�`痘{�,�9s�ˊ�z��'#D����O�wC(%��	7Kl�M���/D�����%M͖�C�)V 6b�@�g�,D����E
t��G��J�-R�'%D��v�Sfڸڤ������D!D���d��v��c��6V��p��@<D����&���q���}��S#(:D�h�DO@64
*�Ȕ�t���k�&D��bE�$ t���f�n�00D���$ ��8�� �b�X$�N=D�̹kS-1���;�'I6pA�L�`D;D�d���A��� ������N�!�L�8�
,SA�bLVL���Y
M�!򤚂o��@Ʉ.Q��L8�	�z:!�$�(*hh1�=�P�
�&!�Dݎ7�J��'(���T@ ��-el!��B;9J�d��%\�g]�����1!��W�YV�r��ȻK��R��Ө1h!�\�n��a�J�����$K 4!�d��o4�U1���Z���Je��V%!��͜g�2��E�A�tI�0R#�!�dH��� .F�*��)�ȇ �!���=��a �G�|�ʖm�y�!�TH�[��
�8�:��S	8!�	0b�HB��A���C�s#!�r�洺�Ē�0�④U�֚|!�]"l�~0ꓩN=KvLq
�nUQK!�D;�n��@�E��Qpr���I�!����B��wE͕o9�pȟ !�Ƣ%W�z����2 8j$��8!��@4.L�5��3⁳㭌!�ė�=f\ئ	ښmxn� g헥`w!�d�ڮ[�,U�}�� �A,t!�dA38<έ��㜄k>BX��!�g	!�� �(8Ō�� �5C]�m����"O�Q�mH=jsha 1Qv�d�`"O�YT$)�܁$�B(2fr��"O" ��CN��(b� q}�0""O����eE�7.΁����Yo���w"O���@���=9��Аj���6"O��cŌ�>���A kޫ��|�6"O�x��苵a�мc��� �8�"O~h�+�/g/�����ݙ:��1�'"OND�6d�_ �2��ۚ&�N��w"O�� g���&x������.:�3"O���qLA�xs8}HB��"�� �*O��0 םY�<u��
+���'�n3R@\3N�dYӻ4 �z�'%R�$�����Q#@�R�e��'��B׀�$|��-�H ,�c	�'<,yR󮄹q9�`�P�Òt��К�'"�Ss��r�a�&��eA���'W�Mb�����5Q�OP�����'��Rc��������Q.N�:�'l�=�` M8;�|��K�56�$�2�'������|�PcD�r��'��:ƪZ����Í'�vL*�'��s��ܱt�@���b�?g���	�'(��l)!�4u�皝.E"(B	�'����mY9xtP���0)�����'k����)6T�GmߊW���S�'�-�ׁ\�<J���7��]���Z�'ߨt{7�*U���c���3V��$a�'�JP�o� ZeJ��GP����'�����8D��!-LI�|��'u�xcQ	�,��l�v
�|�z���'����Җ tTI e��m�+�'+� k9Y}Z�A�O?̌0��')��@�[�u劉�đP�Z�'��� 4+�"XS�jN�<4T�@	�'��!�W�ɫ/	0��<0ZXC�'؅c��U
Ui��(�� �<�5�	�'��8��M@��y�'J	f,�J
�'���J�"�`5.	2
S��'�85�$J#;��q�[��(��'G�}�AF�3S�
��#ޥ8���[�'٨y��
=u�8y����/"2����'���S	9���#]Mɔ�C�'�p��E��boR��c��1Z�h	
�'�Q;�*A
eBL��dJ�Th@�i�'�*(x��=kI�N�Im�L��'��"v�m
�u��u JM(�'J�ڧ���8v@�td@/="�9��'M��!'�\&%4���#'5�c�'_��^�=vu�vҍ0�4%#�']�g�I�J褡�N^�/(.��
�'KT\��N��V9Ό�a�-�@�
�'J�LA�MH�L�j�hC�%JI
�'�����������CF 0rp��'�5��cذF������6`��c	�'��R���n��d�T���jl2	�'�iq5��?��P%��;c=���'�D����qZ�#��=-N!��'�¬#5 F�T?v8!5���4�����'t,3WlS�P%
��O�,�Z�P
�'��5��2��s`�4^|��'��0�ƅ'��x��W�O�I�'= �W
w���Bǋ��N`* ���� pM��c:	
r���-��n��B"Oz��F��4<zr��'���!����"O
�ф̊6sD���G�MӸ���"O<a��$1�h�rw��|WA`"O$���7��!'�!@VȰ"O�۳�V�'/F���f��j�����"O��娏v@ ڄ�Y�F� ��"O��Cb �2�Qz���<P�XX�"Ob�35�ƅG�������'"O�5�����Ru�, t�X�qy���S"Oj�s��?d�i�E��t�
�"O�ػi�Xܠ;`DF�^d�Y!5"ON��L�>s6�K0+�;Nl	�"O����L�%���b��#�0�"O�L���At��%(��K�����"Or�YU�W>&]
�2'&K�1��0�"OB������a{@���!W�jD�"O��wl��'�d`q�-_</�Nq�"O49sč�9r��h#oW�+����"O��Dgҟ0�L0��@�*2w|�	"O�Q�c��5 �)�	��z���8�"O����h��K%6��pjU�Z�1"O5@4_
���1�	[(:���	F"O\�Q/I� i�$!�$���"O�(b�%ū
�*�cDo�s���q5"O~�CD�# m�D���.,d)ʓ"Oȭ22&O�EirsFOW;85"O�li�$Y,g��qPc�#d�p�"O, �ǈ3; �j��B�u|�8�"O�@ka/P�Ie��S��p�X�G"Of4�4gVb���"�ޑ9��"O01�g�,�cB���"O� ��J�9aF+5��0C"Oέ���V�2����N8&he"OVT�c O$!���@8u|1�G"O<����Uؘ�(���A�\��#"O蜨�c��:��|)%��*����"O����D�:�p��ʀ>-p�$"OV�S��_�a�ޑ��J��F�<�z�"O|�d��Z�JdrG�� N�����"O*�𥅒�g�h�CרNU�RMh1"O܉2�@Zw�Àȇ1<)H���"On$"���7;|���L��!�w"O�0"ql$zx�#Cl��	�r��"O�4��l�s]S��5�>��"O�E��J�u�)���W�E����"OL��B RH'dI$�5o�ơ(c"O��H����x�T���H�	Cw6U��"O��I��-`2�߰U7.�I�"Op"d�W!;F�Ab2���d*�q2�"O��R!U/[��w͐�g^X�"Ot���l�h�*"��	(�"O�U���ZM�Z���ha��"O�u)���gt|�`��+f��R�"O@aՃp�H�ߎ����1"O���B�Ƕy{X���G��( �cw"O���Q)7A��˶hN&#h��"O�h�M�8��S�� ,�ܱ�"O�q#���)h����
M>;'0�"O��w'��-6,�0�	�4)�JEx"O��kb^�l�4
��
�dBr��*�!��U�0��d
�Y0U��'��v	֠I��qB�ޒq��Y�
�'�	�N��*�0!�%�4\��9
�'鲹�s W�(LD��TGτF�L��S�? p0�%.��k6�ܳ�'V/�ּZ$"O�Z!+��\��y�'ٔ+ҖD��"O�����>>�I5fۢFà} a"O��q� >Jl���e�
�����"O������B���2"V��y��	6��V�k�f$zb��n::C�	�)�H��aC�3�l��E� .ZC�I?�HDpϚ�Q��c���V��B�<0M���oU�6��K�͚I]pC�������X��e�F!6T_,B�I��`e���g�LC7C�7vLBC�I<E&Q
����xD�P�"a��g��C��� �f��<F�L5{DoD�jgB䉍8����tk,B�C�F��C�ɉe<� �F_�}I�Ր��PiJ$C�ɍX4��9g���yΘ����(>�.B䉏kD�ř�lD�`�87�c�C�I�}��\�F�ξ%(���FÇ5V�C�	��fx3Dl �>������%C�C�	��6x ���G)��.�z�hC�I�}[����ؑh��x{��XB	�B�ɨn����/��\t�ф��ҴC�	>xJ^Ac6�K����l�,	1x,�����sMU�)y��0j	+*������1� !݌$(lx�K�JX����nɮ9)�Q�8��(�M%W[���#k�	��k��0�֙��
�$�$��6Ժ�UF]*Nn��tEK�x��ȓ\4�����]�@��F�Q݅�$j��֧��khn�s���ZtL���4e���J�e!0��*]!t����ȓ�� �Ф��P)����aV�
�*��t�"x���R:��iS�d�=�����?� ��&q��� �c��фȓ9�4D+W���u2�=�uE��[3���ȓ\lY����d�T	Z0� �4P��s�W%�%��ѱ���W��%�� ��B0	�z���)ej�e�����-H�ZC��^AZ����	�c�.0�ȓF���k��?��Pi7E��`cD$�ȓu&*YXBAQ�բY�I�",y��;�.9�W��0)k�B��K����>����FJ�s�B�p0���,��Z�DaX���D<>����N�|p����6�F���"п=��٢L��<4�ԇȓk�!J�	��@��P�I��L�ȓ�F�t��7J�9(�B��䨇�c�>)���֢9�Dų1�
B0��ȓQ��9�`)H�s�Fu�"^��.l���P�yf��#X�:KoF�8��h���XX������5��]�؅ȓ ��,���IQиq�J���8��ȓ0R���g�5���ѩӢ$�6���~����E��/ΞHHd�AZ���ȓ�耦�
�����*:@��Pž��h@ S8,�)�nM�hMN-�ȓ&�������iԂ��D�!�(���i��ؓ�gղ]t�(�@��>S&ȇ�\�J��o��`���S��p-|���L㔘x�[.��J��Z�+h6��ȓKی�i`(�;yDN�"�B�?��لȓ�2�Zo�j���;#�	�N�\��]��8���7yR�BIK�P��L��1���T�+`|8�t��2>6�ԇ�S�? �s���4Tb5��V�r�!�"O��r�Rk]Zs��T��x��"O�(p*�*~t���Ih�"O����[},5�%%��2��;s"O̛��.�lL��c®�:c�"OX�a� ��=���r&b�n�N#�"O�iW�G��R���E�Nm�X�F"O����V�\�F���
�
5
���"O�b�@��%�d�Z��8Q"O>,�$�ׯx
.��A#`ج�"O2qI��*	�TD�d�ʷHp(��"OtT���C�G;*a��V�-c��[t"Oܨa5!�.^4j��u�B,-��R"O�y���S�
Xh��J�k:� ��"O^<B4��/m{lX�D��^:p�"O�eq����L�7�	�8�Y��"O�m���_%p�z�
p,6���"O8-�F���ۆ��E�܏]���W"O�������� #s)\$gQ�e"OЉ�t�ä��So�S}�q��"O���E�.��<Z�HLgL���"O$��#)�&~Ҙ;&(�`��h 2"OJy:�a�|� �9�Gϰ*崄�4"O�xW �FbԠ[�fG*;�di&"O$�⥉ē��\HW�����ˤ"O`�����#B�.AhS��25��u�4"O� ��ض-j����R�E�"OQ�wdM�[z1٦k����R"O2��tfz6�iT�
e�>ݹ�"OzmiLA�$��� t��%K�eZ�"O���@ݷ,��ŏ�)*Шx��"O��HG�Fe��s�o9�����"O�y ��	o=��H�B�6��"O|4�Q��-��'�� q�r"O���
ޅ vT|a"��㰴�&"O6a�E"PM88�dկ]����"O���r&µ�]�q��!6��aS"O05���k6*w��v�n�;�"O��yV��N�⧬W`�.�A�"Oʤ�@�L�&ox�`b��] (��&"O��rD�Ӱ, ����]�0�"O8�␌�B��u�@(@�uc�"O�1#��:Q\��hB@/%ŰQ��"O�r"(ֿC��pS�H
.��å"O�e+���$s&�%�R�Q�7�x��"O��a��"#�:݋#�֙�@�+g"O0e:sE	T!8���,�<14Z�"Ol�'L �J%�i�
�[F��7"OJ,2�:u����)�Q�dYb"O��掏&0��A��Q���"O�5bBi�hvܒ�N�@���a"OJpZ�d�,I��䭐%�Ե��"O�� #Ü�P^�Q��H�_���"OX�;�-��]����'^g�� "OmzAG�%w �5���QM����"O�s#EH�vu�)�r�>8A�]��"ON����@l)X��45����"Od��Ǎ n� 4!���4�I"O�r�φ�~�ZA�ŭĦ\pv@��"O����Z
)Ǧ$� �8]��Y���'(��D��١+�e:Ŏ�- ���D*-D��SW�@4zZ(�B'�,�t�p��,D���q[4\0-��*9������ D��QIԮ$/�\;t.[�U@�%���2D�� ,�:��ÁRn�9�˕�L�H8{�"O�Ur��	�u嚠I�
ƻ���X�"O.-0�D�D�:5c�DL���0�"O
=�`����0)K�Ã �P ۥ"O�R�#S%��T��1"�6Z�"O* ��]�Ȟ��Y�x�V"OT$���G�Jl[���J�$ə�"Oy�0R�QI\�cb� �PL.D!��4�t!)��S)%b����G�@�!��$sP���1�ݷo��}i�,�/$!�dY�w\L�KJ�$�|q5��	�!�$V�^���dP2�>1�JX�'E!�D�Z�y����bE�Bi[!���%�z�iQ�MR�K�(U#�!�dջT:ƍ��ʦW��U
�Z2:$!�Ĝ�<oV��B��iK���G!�ď+_M�H��
C�$~���e�	�!�䋈F�("T��Xh��ЄJ�
�!�D�)6�x����?l�l:��Ӕm�!�d�> 0i���E�P��5gR W_!�d�9e�JX�C	F�!Jh-a��A�!��#4p��!@"\- ��P+��=�!�$F-o�=���Q�xҎ��G ^!��3K�lY�bE=i[j�p��eN!�Ԡc:�: �_.w�lh#6gP�h�!��Y�mpPe� O�/�=�w��k�!�D��՚c��:XD�� �Ԍq`!��S3nH�dJE���iIV)��$�'*�!���4#V�0�JΆs<ZH���;�!�$F$`d4� w)ZbC>P,|�
�'�d����n��C��̯L;�x �'�!�an�|�x�tRi�|i�'���Tm�^rLa�@�H�zm:
�'�t��	Q�B�xXP�I:�v���'���#�'�9K��j����+�6%��'h����号a���k����2Lh�'
��"�ŝ�v5ȷ���S	�'��&�0ٲW�$�np���yr`�\�ZH;P�͟%�@��ʟ��yb�Z06��e���� �����yB�Z|�0"	�4Z�R�J��y��B@�d<�b��M�Z���y���S��T�D䀎�
$�1��%�y�AD�[��YQ�߶jFDA�yrBŮz�Rh�%nU�^_�ó�Q�yb��w�R��Ԫ�Yy�lRì�y���(��\[�(��>�ĳs	,�y"� �P��1ś2;Q�= cBז�y"G�5�*��A��9����F��y��V���P�gˍ2�P�B�F��yb�F.Y�x��E₣#�K�$�y�*)��; Ր ��,B�f��y"$@���P��^�A,��v�R��y(�&5�� �Bȸ0<��%ۺ�y��s� ���o�p��őƄҩ�y�-mD��qsl�<d}����+�7�y�l��3Ffh�4�ܑ&7�������y�^2�BP�5%+�8akg���y2��1�r��ā�K����˖�yr�اZ
�p�F <K��1���y�K%���0j�H�Q!�ϵ�yRD�����)jW*G��%��y��E�q��Is+�=���`f�Q��yB�Ӡ,-��)�!Y�e��1WI��y
�  ,0��ܹ~���t�8u�9��"OU���)_�`@ۭL����u"O�)H��A�(d`���f�l�;$"O��3uG�R)��٦!� �	P"O�����F|@{򏔕Q�>��"Oa��� <��M�4q�(D+��i�<q6B��FakG�)0]�a�<�I�O�6Yp��A�N�y��u�<�Ӌ���+Dנ��n$/�B�?I���@R��X.��b��5�B䉪a�h����!�VE�)edC�tְA��n� "��+�+C�.C�I5M%^�iצ �s�~��᠂<�C�	� a�Y����W�&����Ld4�B�ɺ&�9 �Tdb�L�u/���zB��"ؐ=Hql�L����ކ��B䉥��Y1L���$#�m�{��B䉨8.D�q������۲
�3ZL�C�ɣRqt|���2�������&B�ɰq�� U퐓P���bhX4Q!�ڎu$� ��	�}��h���!�d�U� W���t�����!�Ğ�AK��+��(P�'%6*�!�� �v�[�E�R�(A����!�G��ʐ�+G��U2g�[��!�d�)����o0E~`)(bc�>N�!��϶'��}����;m�Qr!���!��]�G�Jek�)S��[Ҋ�	 �!���0S��Rt�t�*uF]Nv��'~s�gC���k$�F6E%��(�'I�8��hċ �^�Q�GZ�B2�h+�'0���.�n�Ȫ��Ƕ3��h�	�'����٬n������[�@=P	�'(����%#z
��WQ�	�'�>�j��Qڀ{EI����Q�'߀��1ɑ�lHT�t�G�(�V�0�'� �T�P2y@us��.�&���'� ������	����/�>�J�'����K�\������5��!��'�بJ�OX��Ic�V�6����'�Z #���� �� y@n��.H���'q����V�)����w��Z���'=�=x��Y����z�阻)����
�'��0�aU��d1p�I��#zT�r�'m�t��T>\R`�����q�'���Dɚic@ ����	q&P�'�%�I�8�9��@��5�	�'���[��H1���j�MP܍��'�d�BN��^���ա�y�J��'�2@�@�	
^|���ʬrn4ua	�'�^@�w�]2"����:�A�	�'R.3S�Q�,Uuj	69բ���'z�eP�ބQ `��/ҳ-B�ݒ�'(v�1�G��`NJ�2E��&F�X:�'[��KG��0&ry��D�+7��A�'��!�3,2�ڨ��`	(y>�d��'�4�!�2���h#�W��4�p�'�NQ���0SF�#s�F;��ͪ�'���"H�h�Q�� '�����'��0-�\���	NMQz1j�'��dr��U�.\ 	�S&E
HP�Z�'(�YQ-�?e�	P �S�F5Ш��'�8M�Ǝ�|=<��JI�(��p��'�>��ᫍ�r�.]�vMB�p��J
��� �ĉ!(S+0���rTm�\���@R"OS�&�@gf���
�FJ�@�"OP�s$k>?�H��ugz�����"O�M#!�	>r�H�2A�N�X�*p"OFu�U�]�j)����K�>��٪�"Oh�"�(�$ {!*�h� �Ѵ"O�2��׼|H]YJ�@B<b�"Oʴ��EX!O�F=A� +x˨�8�"O���a锲{K`����=�H�Jr"OXL��΍y�ڤL�+d���83"OD�󷇈9^K�A ��&AT��"O��#hÑa耸cTj�>���"On�ӁA�O>�*0�ʅN&r'"OΑj�M�ET	�N��,k�}�"O$T�n �s����lѮP�(�w"O̹��8Dƨ]�#nѹSڌIx�"O.0k5`�h@�ӭ�x�l�$"O���VJO�=F�B�-�*&t�J�"Ov��7�ę1���!�?V��-j"O��!���6�����ys���"O���#H¦X�!`_�y�d%Y�"O�	S�ÉN8B�f+[�,��!�!"O��S�#�Vi4��#�ʫm��	�"OP�(Ԭ l�� ��H�p����$"O�{0{��|�r��e��X:�"O�d1�	�[�]"��T%y�����"O�P@���1醥"���`3p}��"O�����801��0��g�Pd9&"OnP����Ԑ��PW�:PIE"O��BMU�������x�'�ސ�R�hl���ǟ�+��Q��'4�}�G.y�F�
5X�(L [�'U�E�AL��V0y��A4�ʄ�'�>��S@�;Wl�R�EN4���p�'KN�QI�D�����DF?�d�#�'v<�X�d�<1�]�č@��R�(�'��Y�@J�.��s���tz6y��'怭@�O�=K�1r�h����'�pأ'W�Z���	�����,�'y�+��?�N�9&�C� �޽k�'f� !���7*�h���@~Bֵ�
�':�����;A���z6��a�䨲�'�2�xc��>
|���n�T�|��
�'����iʭzh���E&@�	�'�t-�G�I�I��%����,r�'��bq��/O�8��a٥p��Q	�''|!�R�Ǔf�vH@��L�y!"t��'C젉eK
�x�x�GG�w�&���'_J�Q�*� رH	�eb�J�'�ȡ���ɿ"�v\��c�91�N%c
�'~���&
"PH���! ��.��'��9C¥4w?v��PD�%*O���'dx����'����V��<O} 9�
�'wN��E�^�.���Xv�_�?UҸ�
�'W� ���	q���@6���1�t`��'�H�ђ�ם<���H�/���b�'�6����\�>Rd��F!4'�2չ�'���#��ǻQ�8%p7�y�'�ڡ�cTT&��g��$`J��	�'N)�PgW�=jD�:�`��R�x�p�'��{�A�>����q�W����'����=�htr�K_�U��C�'�h=��
De�M!�����y�'5���q���z�3s ������y
� "q��'ǣH���r�>OW�i'"O|<Å�߉�P���E�7c���Р"On�#� YM�P3�د9��`3"OrD�'�!{\Đtl�1x�Լ�1"O�I�Dg�]�B��bF��M1*O`�c���q��$Ȣȇ�*vLQ�'�8�x����ԙ�c��l���)	�'�
��S%���
�Jj%\��'ub�ۤ�N�,T�g�9t~,��'�`|k0� �q.lu��!MkkX !�'��Ygh2.8P��'
_[|iA�'�*���3}Q��ꁣ��%^���'kH��@0}�����$�L�'Ƥ�S�S�v�b����gJj�*�'nj����6�rL���d���k�'*A���C�yW~���ͅ�U��$!�'��%�fCJ�%E�pkA��N��!��'Z()Eˀu�*����^�J�C�'��ZDnQ%Qz8ba�A�I0$	��'DBl���ΪH7�-8�&�E��P�'�@m	F^���� #�/o�޵!
�'Ȱp@��3�,��֩e|$1x	�'�VIxqa�2D|�1�gNX���	�'f�9c7���Ż��
a��`r�'�tuRs��*D��ub�I&T�> �'���!� *kh��i�	��Gجuc�'�Br	��´�x3��qfщ	�'�vXcr��8L]d��5���$���'C.��҆B�T*n�+%j��<��'}"�"R$ҥ"�0���N�,��A�'�ayv�"@&�@�'@��x9��'C����A.*�.D9��P���X��'����(�)Q`T��KٍP\*`p�'؜�9R�а7���T6P�h���'�٪�L7e�������,=�����'��P#���H).�u�_�4�ua�'2� aA� !:���*���-��'L"��ׁ�-�4 @�i���D�y���*| ��#�}��:��2�y"Mϧ�P$[$cX-iZ��V�ط�y�H��1G�J�{�j�a��]�yR�	q@l�-�v"T2�k��y�H#PU�mq��Z�us(P��)���y�H�+b��*d`Ưs
ؽ��$Ћ�y2�΁��u���ä7��ԓFo�>�y2�W�N@0Zu,�73 ������y��Vo�@bl��+мDSu�ŭ�y��!]��T�2&��7���#�K��y�E�%<�k�9/���EQ��yR��fg���r/؇S���k�.Վ�y��� t���3R$�M�ꝫ&CH��yi_�6�~�D��/�ƍ�֍�yB�U�]�-#�c�#-MH5��'�y��
j^d\�wÀ��t@�1��yrkS�z��T�q�Z(e ��	��y�"J�M!2�!0cǂ
H�ʁ˚��y�.+F�jaH��-��Maŉ+�y�	�_� ���"T��������y"�ݓ��S�.Q��4 �M�y��4+.A��(�]׆%��?�yҤI�7�Ԡ"��^�Gzi��ׅ�ybc�`�|�y�%�7�@�5�@��y҃�: < S��N�/��xU䑠�y��G�"�`m��(�* k���y
� ���Հ�#������=0�2"O�5։�{�J%�CCW�]7���"O�I��9]{�<�sa��+��pf"O�B&m;z
��F|n,J"O�ES���k1�a�� �(t��Z���՟�[�EА8ߛ��I��Y3b���EW[NK�F~	qO��$�+4E*��b�ЫDI�����5n�L:�Oj��r'�W.r� ;��J7>�%���d�����I� %\��ף[I�DR����#1V0�� ������vnG���Gz�ݑ�?q��_Z�O4�FM�5/xl+��X�ʈ�P��1g�H�D'��i�Ͽ;0e9,��#�I����qS��e8�8i�4G���i��;6bXC�ɻ�0���p�'�~���O��ī<�O��'>�4c"��Ox����N2����CH�\��a�E�j�@���:JT�����Ͽk��M������2�>���צ�P��цo޸(a���6�Bٳ���6s����\c�8��!CX~n6���1%ut���44d��I��Müi���s��D� �yT`ve�F;�(��O�D%�Oz�a��҂V�x���H�������O
�m��MCH~r3�]��u�o�He(UX�!�u�8J�I˰6�Pʓ��E2`�iYay�g�%H�n;`�[�} `�uB�j�����[� �^E��ϛXĴ��G��lYz���$+s��s�i]�"kD,"f����{1gE#�8�2�F��Rt���Y?��ǩ����'Y��)�
�N�l�#�/�x$�I˕��O�����OZ�O���Y�D�	Q}r#_�7����v��7t��q�>�y�c��\\���5�
e�l��棉� ;xr\f�l}�i>q�_yb+_<�����cj.}*3��$��P�"N`�R�'a"�'B�X��'E�'�tԠq�iऍ;R�7V��{%��hW y�dg�,I������Wf����$�����ۅ9B��I�hԫT�q3��= 6��"S�2��B�,CD`HFzc��?)ߴY<�Q��M����UZ��ʸ�.�W���'��I�8�?�OB��a��,
��|���[�f�4���2�����`0�A�Ь_�Ki�H!���0�(����MCB�i��Ba�H )��O}U��n��?j��pm�?K�iS&~rqO��䚫�Y���Qz��91�V+q�~I�O}yy��	y�}
�kG�k�H�Њ�$N	�t�$���9����5��5^PD��3N�KӚ�i��Y�l�0��0�*1.�uFz����?���0���')�S�W���J[Ha��Y>N&�<p�oL��?������,L��_�&�FD3��׾SU(��R�'h7�ԦAo��6PT�q�%b�(a��|�����':%Pc�OF��|z��?����MK烝�=G�3o�
Z�Q�ܷt/~�PCà!��)�g�� }�tdb�/�"��e��r��%F�Ԉ�O�U�
I�@�{�pt��-7�� L_:)z�� )�����\c��ę�_��3���?~R�B�48R���ܟ r�4�?ы��i��9����[��1ipDU�-��!��'J��'�ў���R�K ��XE!���S��+Q�	�M�Ӵi��'��ĺ��F`��-�� �1B�~��L�I}؞+
   ����0d"̍�I���p�{1��(�O,��O����˺+���?)Eb��X�"��31���Qr?٢�4�Of�q�и1ȠH��ݝ?L�� �O@	��n
�#ڼ?�1�'Õt~�������	���$���	�t��ґb����H(��,s�vB�I�b�(�0$�,؄�@�΀kV(щ��?	�'a�`�s�xӜS����C��i�`(؜SV�䉴��Op���O��dI>3��D�O�d:^���O���,�"���p�\�ydd��'z8!�.O؈��Eb�p��S��:5�,�u�'�ܔ����?ab�A�{"}�� �^��SU�g�<�rl�%=�ac&��*�h�]|�<!�PN	2e���Y��-���<I��$�)QֽoZ�$��W�T,[DFhY���36^})v�u�C��'���'w�M8�'L1O�S4)����N�	-�l����T�j���<�DLTm�O�ڌ��b��_1��C�?O�l����$Ʃo�R�S�fpT����ƻ7�LD��P�rB�	��p��^�u��#JԓO�H���Xb�I:?��9���"*+��Mܤ6BB�b�jw	�*k�ؙ��o�>B�)� ��k���1Xk��J19���;W"O�Q�#�P)MG
%��NV
B���	C"Ob� ��UW���sd�&\��kG"O�� TH�2l��	�IfVa�R"OBEa�剩b���#Ѹ�~�	@"O�d@��D'ԠK�-�&]r�x'"O��'
�*���y��Rl2�s%"O|�Em�!
�L�@�YK�<pr�"O�\SR���{vN��S6y2�"O6L l�@QT�;CG��-�1"O�����Z#Xꐚ@g��3P�"O�%L5$6h)�b�D%a �ٳ"OZ�auf�ƙѤ'���z"Ofu#S���i:
����'?x�3P"O�:TL�/e�X��e	 5�9�1"O�Q`��	2V6�����*/(n�`�"O���(Z�!"df.s(��4"O�U(D3`���(���(�U1t"OB-� �E ���Y�F Zp��"O�x0�ڛC��1B�@��Θr�"OxD!��+v�&m�:'�ԁ�"O�m�$�@.#�%p�,���y�"O��%$��s^��d��P��d�"O4�����sV���2(����"OƩS�+E�/F�"��w�JpA�"O��j�ݾn���`W2�B�j�"Ox���]f�{�!p>e�d"O��@&G�&t�0��]��C"O�kA ��x�&Zs�T<V2���"O�4�E�@����RcS-1��R"O�f$Z�+f�����,<um�#"O��h3MLhަ�9�!H2CktU��"O4�'E�T���K@�܌%k49�"O6�2p�����
g�.U���;"Oh@�h44Ђ�o�,bc%"O�rW��C�0�[�.�4g�x {5"Oy�s��!`>�P�]9�i�!"ONR�-~GX�q�L�� 3�"O:8#�HA���'�<b�>�d"O�} 'M���R���*�>;�>�d"O� �lܷ_���B�HKO�iD"O(��d�J�lD��G�T�\б�"OB�{�O^�I��c��k��(;1"OT����� p�D�&D��0��I�"O2H�w!�l_|P��"H�0j@�"O8@H�Ő|��r2aH�2�꽱�"O0�����~�DS�D+Da�:A"O��@bm�;$vT˗�ޤo!�*R"O��!H��
���H��Đa"O�1�V<��`�w脺�!�Fyr��1H�c��|7���{�X �⌍��;5nX�<�DCPh*t�!tBw�Ra�Љ�T�	s�BA�ϓZ�Ab�)�?w����U��25�zP��	�{R�a"�(���L�e���4�k3��#��x�Ѻ	r��bu����������O6���_�'! ���!�	U�"4X�L�~K��!Q�����~ �U��f�<qb|��'D�0�m2�)ʧ��%���L+���:G��h�H��ȓ-�<C�(�Tr��J'Z�~e�H$��
�[���<���t�d�����K�
x<���$$����@a��:k|Zw���k-nHbO�	4�R�F���u�;�p`@�"O��pM�@�
Lc1$L���tq�"OyK�j��D?0��b�(�| c"O� ��XqKעUVtm9AL�P�p�"O&ř`J�%vZ�2C�H�j���"p"O�){s���x$�:@�����8�"O�]�IL�2V������
�F �"O��� B��u�ʝ�㧂�
Rr1�"O��;��L�Y8��Ɖ 	nu�4"O��� �����6� H���"O�mC�-�>)~��p3�@�Ҁ�R"OʁA$D�Z�<}���[�H�8��0"O`� ��-�9H��N�u�DT�� 
.<��ɀ8�� zVj�1rF�E G�[3m������{�O�,���A�"�(�/�(7:J�2u"O�eڀo�<-��-�.R�^ ����$Y-B�⟒��%�g�C�ބ�n�<_(Ӄ"O�"��c���]2G��n�k�Jʣ|�')�����[�d��b�^m��' ���0JמJ�]ڴ���M��U����d���"H�B!e۩[��i8��Veq!�$M�I4�R-�1P���FY�!��?8&� ��.�4�Ԁ��f݋�!�SG�������W�XP�CLٟ^�!�$Ӳ8��Ŋ6��y^��gj\�%!�$��y�I��a���)��1!�D�+(�jՂ5垈zF8�i`遧#!�L�0�l���wH��u�!�L���"~��9i'�}�!򄆓̜��3S��Y����z�!�d@�6��\��`"������!�<����5s���)�!�$L==��PG�B	}��;AO�!* !�d^��dy6c˩�����F�!�dЮFl-�����*��!�>�!򤐀~�U�ТƐNj(�ЁI�@|!�d�+c(^��4$Glr�5p2ϱWu!���, 
�I�Aˎ	�P�z᎜%	a!��Q�?�Fxv-7}�ZuI��ʶ"T!�ę�WZ�Y !L�#5����@@�O�!�ĉ�E����n?z�^�)�� �!��7XHI��,��m}hȣ�ǆ`!��\�n2j�XGl	� d:6ս7�!�˱U46�h���- N���%6�!�$\�h��|p��4m�����1&i!�d�p%�5�̀qߪ��ƀ�*y!�D;�b�ɥ�ӏ"/�`Q�l�~!�Ă�La��J���O$X�Z�՘#�!��:cȝ[0$��&���G7I��y�$��"��Sr�<q7�N�F��@�Ȃ:�4q���v�<���܈2\���ЦC�|f�"��u�I�tv�bs狷�蟊���'�q�L
���	��8K%"Of�K���#�Xp{��̠9&�q�hW�`��O\�P!0�3}��r� �4i�/Kg�)2�i���xҎ��qS��8yxX){���A(q�A)5�^��+G����tK� ki|4�&�e�y�K�"oal�&�<���	h\����J�3���k�{�<Y3@ /an�ۗD�;�Hʳkv��?�h�3k�����s�EV�b ��.,[F0�E"O<��QΙ���cs�H�Z��uʒ=�OЕ�'�5�3}¡V�L��M_�m��� �6��xB�.E�@�# �O����FmI ���$��;
b���I�|�(\k� }�����W�,"��ti7��%\��D�'d�JP��9h��R/ SU,�
�'���s��U��m�0��3Z�H:����){~L47�?�J*dOL��y�ΟW쀜G�Q�t��X�I���y
� phY�[YD9�&L<iJ�� ���(P�p������Tڢ�����>K�!� �_j�<�7	�#��(���B�G�\��!<�=`����?�	��G�DI�$�-��)�Pe*D�ě���qy��+&����*V�	�6Mn�=s�̀2�BĬ;�0�3���k|�ӈ�$lqK��̖$j6��!\�:�-��Mj�4�F�7��Yf�U�K�H��L? �D�zW���%ƛv��2��',��>}1`!�Z�vF?���!�<_�n��T�!Ky>�b�ʘ�s�ӧu���3���SB��	5M�ۅ˟ c�zp��0����p<�t��k����N\�xFDI3�C��~1�R!�k�tk�oT���`�Ʃ�T0�Ft*��'�p��$�§F�x)�ϜK�ؘRB J(<	掏�j�*�RlğD��xs
Ԭ��@�J-9���L�A�N���?et��D�R"L���!B�1�����G��|�ff�6ѫ�C��
!nm��n��X���g�G;`QT(��>�I)��	���&:ofX���ϙ0Fz��'��FM��#�k�-m�0ӎ{�Զvטhq4�X*r�}*�.���I��<��JJ\E�q�ʂ3��#�
�� ��r�MZ׬-:5+	-q"џH���/Vn���JQ�g0�w@��o|>��e�F*h(Dx����ҝt��(�� �18"���
��e �'<�v,�d�
�J�,����!��?y��N�V���n�%q�0iƈ�W�剪M�D� 32\�a�њ~�#�Y�8ט�66���ߒA�����ĨV�ƍ�	�?|@�h�ą]����d��x�£��R"4����%r6��#��<	#!J3
HX!�l�,]r�y�ƫНp��5��\�t��nԚM@0�ra�V�X�'�!�	�q<�Dg͈u�ax��*-��Dȳn4V���΅&fI�Iԧh�� ���GXPl]k�m��n[�|���l~E���d�Ie\u��	�Jx��"���}V����T���Y�VݒP�M�8�!��+Nb���'���,��t���;��@�����HH�YJ�2��;LQ��q���6c�f1��:�?�:sf�Lp�g3n�l� 2��[?1qc����'Lk��1��`gf!�&��ڼA��ZH��Ab�B4n�Y�&L�s���[e|�z���$#Ɓ�!a�>)�Gܳe��4W�X�QʟXy�@�(ly�	�P=�����(Ol�@���'�|�C�H�-hWR��W>:��A�� �+-�p)M �z�ף*k �&D��0<1E� 0H\�S��(��)3��C�݀� ��'&��i�����/<�%��._��l`���k�<���P�f푰��9/3n��s�Mp?�3c�����h�*�kD��YZ=�sGDj���Yd"O�ڣ`�w?<Q����!6��|�q"O����ɸX�H��T�M��A�"Oji�bI0�BmZ�	�V���B"OVT���U!P��i�(��$�d��"Od)�H�j�����I2�xt� "O6���dK�k�L���-����U�7"Ov40��9m��eClIt�l�Õ"O�X� �̆}�P��@E�Y�hQ �"O^4��%��XURЂ&F��D 8�"O���B��?pX�H�C#Ӱ;�a��"O� ���-(�Ƹ$3B�RA��"O�A�A�)3YR��C���L�"On�	�mD,Db"eg��*����b"O�`��,�� ��z!nJ�U+t��W"O@a�e�E����[#/E�H[V"O�p fNܒb�q*��O2*X�"O@`���G�vY����;>�`�h�"O*t�r�)u���s�Ĝ|��|S�"O��g �7	ty���LxP�xw"O�Dj�L��2/��7bY���d�D"O��éޮWG��C'��2`�~L�"O�h��J$X�Xeڑ-�(�B|�g"O� 㐊R�\EBtK�)E�4u7"O��$�(n�h�3,��S����1"OrP�B,)CN`@�7�L�)A"O�a�2 �fiJ2N��tȂ�"O���G�d���'��B�n7D�P�)
'DSHA�"�"kj$K�E8D��z�ѵ �*Q�����*4�5D���A��Q��5��ψp�Q�3D�� �ܱ�)сJ����e��T�b"OT�3U��/T�~��1�Ϧ|G��E"O�q�P�.߸I��Y%}��}��"OT�8@-8^|H9�i[q, �3"O���dj�))�0�q"@�gx�q�"O�z�L�&n��M�q�K2��4�v"O�D��%�J�I���S�]	�c@"Ob5����5g���&���5K"Ov�`P� �_M<4��A�T��``"OR���Y=m���BR�; ���@d"O"��,�4i����튮$y���#"O�THG��l�dS���(+Z��"O�zP�]�o��Fm�qF���"OfY2	��1^��,�/+Fj�"O����U�/��,KSZ�"Ol�)L�5(�M�ĀP6g���P"ONX� !f�bH�v�ť"��I@"O����'בU�ީ��m��~Ո]�"Op�1 �#18����C�;�� �"O"�(Q�(;*��1�&v���"O�������:%$��_�٫"O��5HJ�B���r�GբA"O�t�T�$��x��2�2��"O����A;[p�;fR���TÂ"O���ѧ޴b�G��T��"O�GI�]4P�%�ȚP.�"OƱ�! y�Ȉ%��ln�p8�"Oh�1�� t�ra !��)ZWl��c"OZ���n�Q�
���)�;k72p��"O�1��	߅���7#G�K���yr��z��]qK�: ��\���
�y�IGj5U��;'Ԏ�ٗl��yR���!�b���l6,�����y"�,3\|T#�X�G*)@!�S��y(�(jxy1%�x��0:Ʀ��y)��f�ap����<R��z��yb  ��̝#��A6<˖���e��yR$��oZR���agNڊtr�ͅ�IC}rd�B�~DQՊ���٠q�I��y�JUb�	Q�i��l�D��HH�y����\�Ҕ�3OL�8����4���y Ԡamf��OR�4���CT���y�b��e����Ɓ�	D�>�	�'̬T��#��k��|hFɋ�	�'��LY�%�:X���� �J�'$�3�18z�����Ӭ��	��'���e� �X�'O�E���'���{�CM.��yӠ�ݎ��L��'6p���E@�R>���k�<76�lJ
�'ϮZ4BN���5��\45l�As
�'y����<	��c"F��6i0�Y	�'�T-�b�����ҡZcd���'c��HV-#�޸�#dQ$�Z�"O��r��B���1��Q:AL@�"O>E���ɢ>��D"6h��W)`�g"O�,	�%D�J:�f߆1'�M��"O(jQ*��?c�4�F�g�d��"O�S0����xY�ӆ��.�x`��"O`���<��� ( �H� �"O
�Ge��&�\Kæ�u}��""OU����.)���[�A;��y�R"O�$��i�g��"vH��Hq�"O�m���&4�NKM��<�g"O���-sf )�#f�,��A�"O� �ö
��YR�l���Qܜ��"O�Ma��ηr��5Xgǉy�*%)R"O�<˳�\��T�� ��=�n!�g"O��w(ci,ɋ7bQ?�|���"O��)P��P�P�O�3Q�����"OJ 8dfV �b�S@������"O�ay�Aӫs;�y��6:�DH�"OTUP�FF'n�6�sF�Vլɻ"O��5"Н��$0��<�X��"O| �Uƙc� ��+�X���Q"O\�02MV�6)� :�`޶O��}��"O�����хP�4�CCnFW3(Y�"O"ɛ��U.ܮ��G��oB�@C"O�]�e�V�n5&}���%4�@k6"O�|�'�'��`hE��fZ 	*G"O�L+�ӢO�x��Î(!�(�"Oq�f�̊iu~M0�H��;�����"O�mcr�?S!���AǕ;��Q"O���"O�7�&� '���\�P�"OT����؄,�����e��2��%"O�M�"�X�'QJTړoX=H��	�"O����#nFJ��UEGф�;W"O\��A���1�e�<��PY�"O�hB����L>RQ�̞�M���t"OP�a�NثZ��|�G��tv��"O0X	"�W.�tL���N
-tb�"O8:) ���yyS�G�V]���E"O ��T�Q. w��r��$?�A�E"O�U:���� ,U�7#Z|W"O���,]�U���1'mT�"O`M� �_˒��1G;]Ա	f"OԤ`Q �6�l=��=V{�Ę"O"��rJ�	B�����R	fo�}�"O:	i�o��u�LLj��H0m�B���"O���R�u� ��t � �d��"O���#��^�pM�	�M�4Ғ�|B�'�bB�r�H	�6���y4��+�'�|t�5k��~���t
�_�<�A,�rL��R@ѩ,K^ ��N�<a˜S>�)� � #T~�+C�G�<�ϔ��Z�C��8}�ƽ �g}�<�eJ	�VP�gG�4���a�_P�<1DJ�"����<.�|)c�BN�<9sE�{�4D���L�IXШ��AGI�<�!�*I�*�C�[�d�Y�)HM�<�bU$o���2��g}Pui6dt�<a0��/�@��+D�d|z9�G�Z�<���B�[9	�fD�t�MXD���+�(X87���g��ɝ
0�dh�ȓ/7nF��w��m1�J�h���e�'�D��E̩Gc����ۮ^z���'KV����+k�4�6!ΎE��'���`�/�4BT�hJ�-O�%V<�i	�'u�+���42�.Cq�Q6m� ���'X�r
�:D������]:~�
�'�T�F�v\�k��O�O6���'�yz�ě)C�՚�M����� �'���昢We)G��)�Fz�'��M9��V�)k�3��7��}��':nqd�����Xsܨu�j}��'92�7-ͩd~ ���e�p��'��z����ڙ��+ζY�����'D���A��}�va���VN�	�'�����/#$VbB@�E��P���� ��@6m�&�2]�BDԟ2rZ,ڥ"O�i	B��uS�81� ²;U2��"Oh���>Z%�5�o�9
@d�{#"O0�A.G40LP�N��U=� E"Obh:D���T��a��_�:���"Oz��fIL4kr]˔7Bٚ�i"O�Q����!h&��#�O�`��a��"Op= �G�1z�89�IQN2�#�"O���[�-�蹛v	0�R��"OB�2¨�	T��&���Y"�"O.�*b����?�ܘZ��!4��P�Ν	P@)91J�Gb�5�b3<O�7�:��##Uvz�""2��`XBh^ed^B�	~L8��O�?����D�� C��=��S3�&���,��g[x�/�'L�\B�	�3^)(Rk�Hx�%��Ba*O6q���ՓW)l({�c��?�d���"O,80���=q�9�!��V��@p�"O6}j!��\U�q�C�Q�!����"O�	֌ưz�ZQC@�6��u�A"O��(�&
$&�J,j�AT*I�
͉�"O����p���j�^�^� �"O���qH������˂�`*4�G^������/_�1q��6@ExD Y8�C�	�HB@[����89{�,�y�dC�#zB`a�Q��}�+�Qm_�B䉞)�J�A��o���"�C�)"�B��R8�pC�=:IbMpᎍ�&����%�$O_����	6{���
&���cd!��p�6�P��X�X���p�J3X�!򤑟Z�peЦ`�T��T �7L!���Ns�T���%S��j��ؐ/�!��@
���y�
M?Ch�W�AU�!�d�hJ�M��a�����,��!��+F�LaIaL� �%j�!���Z��` �'��U�g��#�!�D�����1�Õ4}��M(���K!�	O�x T��aC�Di�۶-!��
��l�X�B"$d�mT!i-!򤆄�0œ%J�-�ȉ��)]�c!��)I��y$,�?{��mRU	C'i!�S�4��
b�S
�2�G�Q!�$R2�T����R"A�Ap�M�rY!�S�>�$a�/��y� ��R"K!��J=}�t4��D�J�Qx�E5rI!򤖜I����O_E t���$I/!�D�8`�Щ;�!�-�(�'m�Oy!�D�gY���b�C���=0�N�>5W!��^`��J  �m{���$�ŏ�!���8*���:v��nv S���~t!�ą3x�a{�l�l��A�A7i!���L�`�&"U�0=��'���P�!��ſi�E�
�T�8-�r�W?�!�[��j�O٪Zr�1윭*!���*\	ラH
/e�eR�h��5#!�U�J:��r���,hma%�#b!򄛱 DyJ�J^����DڪC!�d�3.N���D����S��B>%!�d}>|4�cq�����g�08!�DI�c�ŰT��+*�%bE��7,!�1Jj�D��nC�R�J��O1#!���f� �ie� �����^>e!��б$*ʡ���D�d�i���!�ݭ�<�aoɠ,G��g��{�!�� P���S�&e�l
�I�2&W�y�"O|���V n}�Qk�h�=)TA!F"O،i�F�;3�����g��w2��"OR������$h�H� $^�)�1�"O�U���P|�%Z�\�D���"O����M�{h��pPa��L=�"O����(#�@I�5A9��Aa�"O�|��iܬ 
J5�@@D"�*8H�"O��`�A o�����@�.F0�S�"O�#U"R;:]ۇ����E ""O=r����l4�PNڶ~R�ѓ"O� ��B�`�h)iDK�O�D�#"Oj8��F�,2�U�Eg�o�U��"O�U����(~����fR$m�(5b"Or!3��l��!���?vNP�"O°"&�נS�l�H�
�)8VU�V"O��#��t@���WK�W<�R�"O����Lf�=���U�4��s"O���g�&^[2�9F��a�}��"O�1 ��X�k�`KB���4�N8s�"O&Ixg�8�0p�Q/�.>r�[D"O��I���vp��2NA�3ؐQ�"O 	C���2�`I���@g��a�B"O�M:'E�i���ؕ�� ��"O�0!� mΌ($ �о�`�"O�k�"�9j�j�u	� K�P���"O���=eQ���&���h���"Od�C����ys�͗`�N��f"O����*�BO��9�3"O��K%�p\��K��\���"O�M�&愊? < QK[�#��i�"O�HR��pfv��J�<9s$Ha�"O0�3�ʐ��4̠�(D$]��"O8���o�:+u���#��BP�C�"O<�ɧ�
0��䐲e�� ��p�"OhT�c*:!о��#^% �쓃"O�@��\1)I�ȪvbZj�y�F"O�I GdN#MJ�8+g��}R���"O4u��ce���#G��|ȷ"OT��	B7x�����n�6̨݅4�!�d֩*_����/L�80� �.�!�d��"�.�)�!�"-�┲�1!򄅶T��%�C�ƄҚ���(&!�$�>5j�D��K�F�8�q��C��!��~���z�غ3��1'��"L!�$��]���7I[6W��p���RD!�X�"lz�qD���������8!�$ҋQخ�˴cB�B48�P��YZ!��߆O�&��c�M2}�5yկE;Z�!�dF�F�`�w�ҤrdD�1�E8tJ!�D��I؄�����;ZX�Pv���qG!�Ę�z��rE��;W�1��I��|-!��F�����ΗM:�0���S�!� �GؖmYcN� |=��� ƀ�!��d�&�i@���Q&�4{�瓕d�!�$ۄ^���Da!�.�n���"Op�ʖ�ݭ~��+f�A-P��<�w"O����N-�9J�d�g�93w"O��"�菙 �(P��"�ݘ"O�� 4�H���P��C�eex��"O�%bAO��	 � �n42\�E"O���'k�� q�^�>��`�"O�mc����� ��ȸ'w��"Op@�Ũ�/jր�1'�A ��Ě@"O� [W�*>u�"Ύ���*"O9�5��N|P}�u*E�
h����"OR���]�ol%�7�L.UCv"O�JuG�@����CHJ�#���"O98�!�$�^� H��g�}sG"O*tZ�m�&��[GɃ����a"O�)!�hR1?��8FC΀Aր�j�"O���Ŝ.'ZI�-W�J�J��"O
���A
�H�v �Ԇ��g&5�#"O�\��^�)׊�q�z��4Z"O���@Z�➠��CŤ0�6u��"O�` �@�%%;^�[��M�>D��sv"O�aP��)#;�i�a��(%0h#Q"O��Q@G�s��24eC;`7<-Jw"O�{�iV�/����X�W2�`�"O�X�E�ՍC��)���U"a'"Oص�@�E�B�v�A�ϛ�Q���"O��(��Q�t�3�G&.\�"O~jq;3,I��LR�'2��e"O.谳Oɢ*�T2��Sj��r�"O�u��"	uR��ʢ1���XA"O�`S�ͤ��Z��˨,�L�d"O�1���u�@�%M�+.3�r"Oơ�U(�77xc,Q�x�'"O��(���j�QL�X���"O�d(�`��^B.��a�3`ȴ�d"Oph�#ș	�58��7���V"O"���@�p*䰒���ڔ�%"O�Ԙ1��	o�
䩟�K�@<�3"O4�� R&f���B��L�ֱC�"O��@��@:�&���!�`�ib"O��9Q�̲f�x{�)D^�X9��"O ���B�1=8m��a�j߆�#7"O���$ۥ@#�;�Đk78��"O��!��b�16/϶k)`)xC"O �C���@� ����n1#"O���p	81:�[@�d��9��"ORM	A.@���P�V�1�n �"O(A��5 *���Ĉ)B�J���"O��x��
�v���8W���H�ZA"O��C�i�h�M�H0$"�"O:u�@��%�4qD.;��C�"Ov$b2,	���$2�*.�Ba�e"O��c"תyr�8���'�V��&"O��1� }z��&%]�"O�Ha�_��D�:bo��MK���&"OҼ24�\�O��\�!���m���"A"O��R%(Tw�e�S��w���"O�@��@�9^��T�����ő�"O�k��Ś>c��&]�k���J�"O��e�e��	�+W�C�2�SS"O���TO�xcZI��)B�����"O�5��'�/n��J�9>��=W"O���f�Fp#�T9����l}p���"O��å
R�s�¥�B]�2��$"OV]���@4�(��g��L��ْ�"Ol�C�(:Z:黳o>|����"O:-��
�n��}Г�
C��%9�"O�x�%N�
x��̚� Q).z��p"O�Ir
�dt20*w��6}Ѡ!"O�����3�h�з��1Z��"O@I ��vAfLs�T!�y�"O��[�茱��B��9[�ԡ�"OԀ ���l��(��_Ixxh�"O� �,'�^�=��MC'�:h�a"O���B�=!%T�P%�3s͔	"O4r�$qk����D�8�,8P�"O< ��8��X�'a��m��\z2"O�H�d��[�<I �@W�n�\�i "O$	�6&�"�\���o�h��Q"O��PR! "|�ɻ�-���"O��2
G�R�LT;�+Ȩl��E��"O��h��K�N�n��K�m�.a�"O���TK,]
�ʊN�>m��"O.� �"B2�e";� M{g"O�2%�+�e��Z�b��Q"O�ܺ%��0�ތ)%DҊnCLR�"Op����&ȼ��ă5l�4���	i�O\*�K��6��d�Q��0��MH�')��j�c�3��as�	��PL�9��'��p���� �֙��V* �����j�+R)�r��m�$-��JzY�ȓ5�Y��l�8&� V��n섇�d�\S�H�z_Ν��j�qu�u��c�4��! ��NT��Wf�"ar0'�����;E���qeOD/$L�4`W�
9D�vC�	e�Џ��\x ׶y0N���r����Xݜ(��0@���}7F��$ePd�'���Sj�l(�
r˸H�`�J8o�FC�I37z�1��^I���AΣ]�8C�I>P�Nк"���}�vc�o�C�I�jA�E�bN�f��D#U�˓�?Y	�����3��P�����.9�(Y�ȓl���3�.�@���mK�8N���,O���ĄV�Vp��n� zM6�E{�O"Qѯ�:]���qOё>�|��
�'�%����$/)�x�����	�)�	�'e�a�@GX0+�H��o��Yp$�
�'_�p�� �YPzDB� ʤz�=�
�'�;FL\�Z��p(�>y�
m)
�'��p�!����h4Hp
F`�&Ű	�'��Rsτ��T�8�)Z��и�'���ۤ�٭G����"-X,a�,��'m6�;�o�$gV�{�j�.t,����'�VuH7��e���b@��m��)�'����疗{0��ɾaj�x�
�'O�x��N^��4Z�(-�X�	�'��<���Ⱥ1͞X�i�B�9�'Uh`�&Yp�E��������'e�A���O@@����?ql�)�'�V�h7yST�g� �^a��'��̚�"2�U�f�E�'�����'�	���2��)���4-��Q�'����>S楩��S*4��'���xa�ƝR�ș	�ރ(T��a�'����� �XȐd�������'�ʤ2e퐣z�t��g�##N0 ��"O�U��D^n)�S��PM�\r�"O�8Â��;p��E�Fjk�"O�����^>�ZX	�E�h8����'%��'֕i�h�*�����G��ʌ��)����/LH���/L.e����)���y��R�0� �eΝ-L�H�F��'�y�L�ph�R�M&#�0Iم�M �y���'c�����6Ns�-��BJ�y"��u�pZ�F��C��0�B��y�+"���C0c�>Co��9$H���?���hOQ>I"�o�qنo�[��h�7�!��0|� V=��>F�0�����&R�L���D.�S��0X}��݄)��r����!��7�h͚���1�$��1�!�;�-��)�}����f����!�dق$b�*�˚?�����T$+�!�Ik��%��"Yv���X >��|��(���Ag%�,��[���/j��-�$��R�O4�`�N�&k�� �L��PZ�jN>������f`NȢ7@O0X���i��!�d��k
jyA�a�<!�Ԑ����7Y�!�؎D���u��j�z ꓈UW!�ě�G��e��I��-+��(�[/A�!�D�('�j�r�@S�5b}�!�ټb����5�g?�uz�K��=����G�^���hO�o�\]�cεf�F�B�+շ����/v����/Մz1ah��ԍ��e��h��3�U��Y98#�L��4 ���m+�!C"��:�x���^n(����(A����"LAa'ִ���P~򋙴c���C����
�� ������&��O���ac�&5�6(:�+�!~��R�|B�)�S��l*�FаȈ!��7}��B�I��٘�� +TɚX�""K,��C�	 $�n���rR�xI5e�)U3�H�
�'���񔄂�4��p��FQ��(x
�'�0Ч�^�6,�XP�o������'Z�����޷"��$36j��"�
�B�'��9PE�
Ō,ƍ�'"b ��'�dEI7��U����	�W��x�'W ړf��,�Ҡ"U�3:��Tx
�'�h*C ��/������0�LU
�'�-�Teϲ)�}s�`�8?�LA	�'����,�0.��Q���[� ��L;���+�p�h� �+�8 5���HE�6"O��ҧ�<S"@
A�;aH:���"O��p�� ��yd��C���`"O5�6��yh4��!�.b]+"O�|���M1c�	A �=K4U{�"Oz��׀ʛT�<��E10���"O>Ei,�/M4Naaf_)0"��j��'M�	Vy��Ӿxs�
��H��Q�0ˍ6�!�$ך�.!d���]�:L���� q!򄊯�$�*4N޳y��͢'茭$�'�ў�>�b�$H�3(��zh6D�����U�M$LP�N��d�@G4D���.Z��\ɉ���D�(#-'D�<S�.^?
�hq4� 4� i#|O�b�Xc�N+I^@�Q��M~��ɐ�3D���T@U�ʵA�ܻ#"����0D���U*��kp��0"�O��H+.D�T��)�+ÀM1DaM�ZD�Ф8D��A2'D~��*C��]W*��$`:D��j�Oӆ�<aඏ	*sb<�0,%D�@'��I��|��c՛Ng
@�#D������ ��;Db�"V����"&D��RU�\ւ���T�e<�R(.D�p� F0%6nU{��љK>��b��O�=E�cB?�4�''��6��([F�!�;%`,�!���'
j��Ǘ�r�!�$}HH��������t��a!�d.&����8�����Ы�!��Y�C<ؑ&�p��T��&G�i@�O:���#uG�=X@��<q�x�����3
��՚��� !��Aqx��Q���d+�S�π �ItlI�.�0h9��80*��Y"O����I�h*�A�"��%r)���7"O�M���1)xּ�f /z�0P"�"O�Ed��U�b���
+w��e�"O���fDn���3��M�B�{$"O@}��,�9	��Q0�G ^��|s�ONA��nT�	_fJ0$���	�0m4D�0��He`08�D�X�I(�)	6c2D���!�K��<J1jU5�P��/D�`pի��Q�(�aԸn�Ȣ�-D�̘�(X$U�Q3�%/&���I*D��ђ��;'�VU�E�8#4�ۃM"D�`��k���p %�k<���'i!�O��䃁D��*�p0�j�◵HB��5pr�M;eN
�G2�|��C� '2B�	7f�����b��*�>^S�C�ɦP��ӨܶsV�iU�O�w��C䉾4R�X��Ү ��iT�6Y�B�ɥa*K�[b�U�#DЬB^JeyV"O�42��� ��0Zcʄ#����"O��H"L\�"	��B�$��q�"O��9�
��m���QD���; d�!�"O�$�7��S���b�ذ��"Oݛ�!�b/��2v!��x�Z"O��S�*ܙ?R4��^����P"O�a��CT7��EM$�8i�V"O�4 �śq�F��W.�$V��h"O����^8`&�A���)－�W"O@�+�˄���٣�ʍ�8��'��9P���8(�f}�I2Xj����'�)3�_�Wؐ9�S�@cRq�')v�B0���IQ����!�(UʴJ�'�!ڱ��>jܐ��Y�!74�0
�'�n�f�B<x[��1�X�
�'�"�+�ȅ*A�� ��Ĵ@�X`�' N��@nS�Z���A$ŬJ�5!�'P(�1�C�a��d8�$P�P�T���'֪�� 1e�ՀU��-Ml�`�
�'�Qq̀eI��ۑ׻O�n�
�'s5Hՠ��@�M�PG��|:H�X�'��!���܀M<
	Y@K8t�����'����B�ec,�!�@�Yf�4��'����n��u�d�h��$#���'̮�u/Z�]��݉�fډ+n��{�'z1``��]Y�y���-�����'␽A�^-D�$�рI�L�襁�'?&X��GM�\KTt�ԁ�{����
�'��� A
4���#�V�l� `
�'��y*d�ƽ��S�n�yts	�'@���N����h�%��o�L���'�0Yx� �gs��qp
��7����'�H���dO$�.�2Aǈ�2D�J�'pv�S�F� 1����>���'���1��n�^z�O��7�T��'��y��\�VH*�1`.½x����'t�	�nS�G��U�$�r����'�&��G/8�mb�.R^Z`[�'�jgi� Q6*0#�
A��UB�'<$����նe��� D1)Ɯ �'������I� �"M�4-d��'jV�a�!�H��p����1*(�
�'����`���|}�s��2\8@j
�'H��5-F:%E���3Ōz�L��	�'Wn���j�x�5����zY�Q���� ��7�C�_�� ��,+�TMk"O,)j�.�$0jZm�VnBm�� �t"O�u�c��17`BA��i�eP6�'�1Ocd��	*�(�,D6O���"On��5��u�n�S�E��U[�"O~���-\;\���6%��ym�E§�|��)� ����uj '�<!s��o[|B��'0f�H�'�M�g�:9�AgβXZ8B�	S�j́ �ƞn���B���**B�	?9�(̘Cꇨ+��� 2��4b��C�`�l�A��� G=��]�Q4�C�I'�n� ��.N���yg�[�D�XB�%E��Х��I���J� Z�V,T�O��=�}�1'�ltH�1�=OJ��D�C�<1�᝙%V�ţ�ȁ�q�*e���G�<I��K�]Y��s0bƅ)�01��O�n�<9��G(EW&�����A~�qK��_�<)�Ꙟ\7 ��gET�N�(�«�t�<1� �{�|��!�#o)Pd�%%s�<Q�BH�%
�3�,�h����fyb�)ʧ+����eK٠zH�hY�Jˠ+ap|�ȓB�(����� ���~� m�ȓG�p��F�:> [�n�2U��(�ȓ����&`ťlm�@: e@�6�M�ȓ���1�I� {�ZK&������(�rΟ9w�^���hQ��܆�\�~ԠUJQ�^Gz�Վ�.'"P��{���{�b��iC4��'���@U��Y(�ԃ�Ӽz��,�S�ǊA���ȓ=�$)�ȿ��T㴀O��h܄ȓD��蔋�JV��2�@O���x��e+X���n��k��)"�%HD��g������%e�|@hƂU�#z����}<���N8�A�
� ���	��t�<)!���Zl��jS��j=2�o	j�<Y����&�ع8���/��H�b�f�<����~��d{V���?�~��0��}�<)�V22�5��o 62�x��M�R�<)ǓY���,�_"���K�<iͅ�X���L����e�fFğE{����2|������D6e�X�0��BB�	!h����I%n��
��ͅ%8B�	."<���H��Jl�a���k|�C�ɾ|r����%�� �T��&D��K\�C�	�T
�00��g�PL�� �w�B�	�:�l�
�.ķ�K���;�����,�x�R����ԞL�t[׍�'t+���y����X�x�� �3�H�@0����t��*(D��	�&^�> 8���
&�|8V<D��IM�E`Phڃ��ɥ�9D����IV�D���$�׀�v��& *D���S�֠
B)y&EX9%�&$��'D��
W�ˢ'ɚ5�W�U5U`�6'#D���\
�Jݡ�H�,e1�䰧�=D���� ��<��	Q�4��I�GG(D�8�w�[�$"HT�bA�-�V�Ȥ�%D�$��O��� K��W3l����6D����*��2sq��Рmi23�&D��F��-��<���� ��-87�$D�PH��¹�F����FX����#$D�\X��V�>�ɰ�3�M���-D�8�l�)7Ā�XG�
�;v��BD'(D�Xa���
�T�Ul�q�`�I�&D�x���fJ:��e�C�0,x�:Pf#D�� ��u��+t5� ���%���8�"O�U�C�U 4�|�A4��:yDT�w"OD��̌�SU�{᧞)/c��b��'(1OJdA3E��z>j�# �!pJ̤JP�|��'\�����@���
���"���'��M��h�(p���&�+�����'�<l� *C5e� ��.�2T�����'��x�A�NȾ�ʄd��di�
�'ޕb��=Lc����� $wR�	
�'880��W�� �9?/H�$"O��B��G<H�����BŕBUXT�p��!��џ��'�R��qE���}��Ȝ.r����'=��[�/[+R��y���xJZ)X�'`�1� �V�$	����l�R9�'#�Rb��2��Aу�F��'7�}�G�L1����#bCN�fY�'�� 25)�(5o�]rS�F�wX���';ĵ�'�C~(���I��n��)�(O��OV�?��'{�8�v�X$�ޅp��� 1�ֈK	��O�}���P:�`8�ZZX��`"O���sǗ:kr�])bb�0dy��"O
�@��Վ=��졡O��]G�|��"O��А. �7،�醏�\,L��"O���#�H�8'�Z5���wL�@E"O4Qؗ�J�j�
����n�H4���'�ў"|r�'���S�g�W��1����>IF����O�}�E`�
%;�$��	Z�l}�(*c"O(���_BŌ
�iЉr P�"O\8�dR�F��Xq`	�(9.<q"O�������5��-%KC|�"O� ;3E
�5�@��ˣh�����|��)�S�'��D8 �X�}�	� �P ���I'�T5 I�%�����eG-�\���	^̓n8��!���W"�!7��=m��l�ȓH�	�3�Z9�9�C��\��݅ȓ	�6	sh��*�LP*�V�0��d��q���S�|Bd:���9:��ȓ=:���G�ɍD�>$�t�J�0R�F���8�j�&a�e.�����Q�g��㟈�Ig�'���_3 �R��P)D�|X�B��&f������I`���'�p����w�lT�S�-<�D��'b9Q�� �g�j���K.t�	�'�tap�=$x�򭈒q@*��'�B����N�H��!�M	�@0�Z
�'�x�Q�L (����F���x����
�'l"�TgI�f]���eo�8^���C�b�'�:��@�O�譱�IφWqdp)O�O��}�A�����L�4����'[)�"Յȓ	�X����~�\�x��-`�"�� �q׆����(p7$'Tf�ȓ(�6��e����ĳ"���ۓ@ D�t"Ĥ�������D�R��d�� D��:\�12���Y>��g�?L\!�dȓ`�2E*d�c%�|��	ay"�'��O��?��{�
Y���7�:$X(��(\~9�B�i�� 7!�<U/Pa��3����B�N�N:�����N�H\�e�ȓi�N�#�
@�s�N>~Q0��ȓt"��Q���)������O��2���`N�c�#�T�{�@�9�v���y����IH�)>��#�JlJ�'���>\JB�S��|�`�BuI�/H�C�Ʌ$�)����T��Jv��{��y��v�z�"T�g4�"��V�Y]�y��S�? "�#��9j��(�a���]:06�'����D*��;�Z�Q�L�!oDp�e2D��a3��!S$�p7S(.|؉��0D��s��4�D��b�7/�F8�-D��p�j��D��BCJ�)�
@#��'��hO�	�a6����Dgs��J���4r��5�|��I�v���h�81hܼHj1D�t�t�ן�и��a 2f�Yw�/D�,03���c~�yZ2"K�z��P(��)��0<%��9ykN��ҍ-���@{�<��@P'�`�TKO�Bm�!��Py��'�O�#<�D[.A
��'��J=pLx��R�<Y�8X�p)W�ïm��#M�<�$�݈@���M��m���� Cn�<i%F��\���+_+>9[f�V^���hO�Wf�dP�J+l0 �Q�A�6۰M�ȓd(q�0�٥$�-�u�B�P��!�ȓ b@Q�#8ߖp2�
�HJf���ٟ��?E�D`�9y}`hs��j%��1R&K�|�Ig��x#Q�*-��˦�p��h��7D�,�fK�Z5��!��	ʆ��І9D��K�
�	�ԋ�����y��4D�(�2�B�?/�����NF׆0i�'3D��9Gh�����KZE,�Y7I6D�����.�x$����W�2k.D��8@�9xY���T)�`��Mh���O���S��}� ӊ\\*�K�:mr�B�T�<!�։;Tlp��7��R�R�<��D�A�V�����;G<e�a%Vf�<)Oۉ,�T1��1F�\"�_�<�� ?����"[*a�����q�<!��P�q�|uP$C�(Y�`�w��x�?!���Oݑ��kNC�ӒP=r��t"Oh���Z$%��@#�P�bV!F$!�Y�4�Ƚ�pܔ$��r�C�Q!�D�2@r@����N%쮥2��G!��"�4���Z�
M��L�pb!�W�=g<8���S�#��1KY;LN!�TsWk	�<<���۞/K�}r�'��� J.ҹ��G����a����&��)�'��H  @�i�� ��iS/l���p�'�VՁS��!LW|��7�EZl4��
�'���*!S�ց�D�?��%��'X>�kw��4G�b8:��̤DAf���'����@$�l%���$G4�ѻ�'麔���"
�Ͳ3�A}Zl�I�'����@a	��C��',0������d-�O����!o��)&
�\i�"Od=�UnL�E~��r��FU���"O���׃	 �M�ӆB�m����"O*�3f�Y+�zИ�ԗ2�pA	u"OD;ec:��u�
A�CXd�A"O(��%oѭ���Q "U^j�!�$˥,�*hi�'n�9��ҪOD!�D0܀A���S���Bf✝g4!�$��p���`b�@�y��`p�aA�|!�$I��h<#�$��8��D#A?4�!�D۽u/�U��H��]:�L&�2u�!�dʍ-Lqe�U�pw��2uϐ���'+a|b&�%��1� G����cf���y��P����큠.� ���O5�y"��4�h��b�����0.�yr��a�$�J .�{� ������y�Y4����G۷?��U`r�ȴ�y
� Rs`�:��ڀ��?{�T� t"O�Y ��-�(�QǧV�T�fW�X%���ቮj� t���@��M27�XDrB�	0*2��#CFB�pf�-CgD;lt�C�-���Ċe�z�r��C�I�%��c��\Q:f�k��B�,ל���b�#g]ty�T�U�"��B��%7Pd)��Y -�l�6BB�B�4 _���7fM�9V���T�m4~��!��=���y�l	m���J�
,�Ĺ֧��y�M�&p|0��!�N��`�6bT��y���o�F�铠I�%�X��sB���yb#H�%a0��!�Z����s�i��y��N-*�#LWZ�3F�.&�vE��'�.�C���.^�m�Sa�% ����'�e��H��e!Ҽx�M\�S0����?y�'�ҍ0��!
jd��Ɵ�I%����'⌅�v�X�I��,�u�RA�<*�'�.�Z	T�K]'<�d��z�<i���}ݮ@�*�0)d����Ys�<��$E)3���ITÚ+�\lF�c�<I��h?d��7	�q���&O`��C���Iw�J���Cc��zi
cc0�t�)�O��	8B���G�I�~�PS�й}��B�I t�b�`O�t�`��d���tB��;'�!)��M�U{B	G)֘C�	�-
� ���#���yB!�1��B䉢 ��uAQ�ĳG�hC4L��}��C�;m*<����0d�$������C�	�EI0D��Q�M>�C���:�C�I�M�x�=�$����p��B�Ƀx�������$ש�:p��C�Ʉ0����ѪM�`�� �&��r��C�	�v�Zȡ$a��1���7!�3Q�pB�I��=���&of11��� LҤB䉨%U��� �k��r��fZ�B䉣p�t���o�8yt)yu��O�\C�I�9p��Т���Acg��C�	�`Q�!���\.Uc�D�Z��B��.78P{a$p�ܪw�ФO�C�I�_���YB�' ��kƀ�TR�B�	UO���0�CY�.ț���H.�C�	4f�
����͂N*t�����_BC�I3~��Hcu
Cd6�9���64 @C䉑|Eȣ�˻X{�� �Λ@|B�		��@�"߲k��P�
L�vH�B�	p�����N(G��\��B�	�` .��DM��T�c��7hVB�ɛN�Y��U�(gJ�)C� �B�Ʉv��\1F�?g�tk��m��C�	�ej1�#��1;�Q�5�^�[q�C�+�>�s���
�Ԍ�$�'YcfC�I��X8�uA��܄�q�C (8C�� � ��$QT�m��D�z��B�I�ʀГP��JM�� 6iO;|2B䉡v����'�X�J�Q�̓�B�ɦ���ҡo�0(�iU
��B�	@�p��d�D	 �Q�4�bl�B���:��"�_�,l�q���8^��B��%��t��A�9y1�-*5m��i�^B�I�f����!���'��4B�I�M���SbP�B0��SVl� B^C䉺Av���XH�^H�C���B�	:S�Z�ŮA�,�7��=�|B�)� �L�7!��z��{�#/j���"ODX�o�7N@�H�#NE}���O��r �J]4��� R��BЁ�];!�\�&���S"�H/tZ��q� ��z1!��$1����
U<@X�jj�55.!�^#t d"3�)��o�~!�d��Q��ň�Ε��^!� k]�?�!�$���:�����L��8���y�!򤉛�4��!ٱ0��R���qsa~�-
�?aU�ݏu��0�$�f~����=�y"�L�r�C��!8I��s�K��yB�T�S����G��/�R\&�y�D� J��Y�6�G�)�x�i��F&�y�/A%P���#�B��h[s��'�y2Iͳ&��\(��־-��/
&�y���*�ڭ�X<��x�@h̐�0<y"�
ҟP$�|��#��w�E����=[�t P##V�<��^�|E����N 	�8i˷��N�<�nR6:�j�؆�	�9��(��C�<u+�?�|8��a�1D�p@H�}�<��HTkZ���E����\}�<	��n޽)�n)b����Vz�<��Y1^z�0P!�[&9��[1��x�<��K(f��x!��8+�ec���_�<y��V!��� ��	���rRl�]�<�V�U|~� /@�:,�j�A�A�<����'��y���e�1:�a�z�<A�G�2c������4BC0h@!�AR�<i�
����Ө�B�<���Di�<YÍD�
in-�	J�<Q��ƪf�<tbC&�d5�U G����M�}�<�P��O_b�C↜�Q���Q[S�<�� �"78d(�ڙP��H"`��R�<�A��2�\�'�À"2�ŀG�Q�<0����u�2����
�����N�<���/MAVQ@���@e��a/I�<�D6hd�I��{�2U�o�N�<yag��(Kz ��nY+䙴��A�<u�Ӡk,~��� 0k89C��z�<1.�d3�	:D
P�il�����p�<Tf ]�Q�rk�X��x�<Q�%C�*����3*�/���) Mu�<�@��T�s��W�tp�2�Yh�<q�B ��x�s�fЯ:ʎ,��o�o�<�2�]-@��u���@�H�~��k�e�<!D���ʅĂ/�� ;q�R�aD p�ȓ�X�)2�x�B���G���D��?��	j�ǔ���R���qN �ȓ� �:����\H� ��>��ȓ,�����&k���%�̭[P��� ��l�Va�qA�<;�	ȟD8,�ȓgb�h�$)�<[�S�F�T!��n0���`!	�e��5;���
Rj�Y��"dHԻB�!��`ju'L�++���6"~�9u�n�ʢ��y����D�9�wL�mxV��"�z�%��_��Y��%~����C�[ %�80��{��y�gR�,.���Ȓ4F�b���kЕ�⌘x,����(����y� ��5ij\i����-:�=�ȓ|���[t��̼\��������,>�8suC´x��4�C�R4Hrp���:ġ'GCWl�bbh�$	�8��T�4��"E�1�`N+r�����S�? *���O��Tm �&�0���
�"Of�[� %A�T�X���W~�]�"O^xPw���U��e!ƃM;;�d��"O�s�(�pXuB�oў9܄=�"O���I	D|i�u�d� X��"O����/ujȣm��T���04"O�x�%^-N(�4S��<� �p"O�,JP.Y�1��h���\$j�(&"O�0��薍i��IS)�&M�Ըg"O0���BEHk���A�k�<e"O|� ���.U�ؒ&)E(HD}x!"O2QX�5]��|P ]�3�V]��"O.A�	�
|;!fK
Œ��g"OV����Hk��wE�/Q��"O���k˃Bɨ��q�Xcp��"O:H�dI��艺N[#<R���"O,�@Ѯ�L/��MTJB^	�"O��8�IE V>�K��U�Z@���1"O���qJnB"e�P+P,H��"O�!�y���)�� �}��$Xp�!D�x"3���7I�]J�چB��D�%2D�D�&@	;h�p��ʙ ����E0D�������a��G6xC��S@�-D� �.
p8"0E�@ߌ��m*D��FB�50��|A�	sؒq9�`=D�·�ų[�`�gkQ�?�^a�B >D��Qb
�9#g
ѧ�.�-B�=D��5 �!͖�p�*K�E .� �:D��A�G�<� �v�ތJ�d4`��:D�B�h�(��u)�7Njd�Re�9D��gC�� �|�XFK���R��sB,D��)d-�	(��3O�;5E��T/5D�P"��ɺ�	�A�-V�ģs�.D�[���N��L#jۦ �
P��7D�kq	\>(�B'JY50����K2D�|{��ν�&��/�]�I¥�.D�<��"�D�R|s��,EB�Ƈ*D� �p\�*�z�GW6PI
���%D� �@�T.y�E�'��7պ��#D��S����O��C@����N�q�H"D�l��F��>��E��42RD+�?D��y��%f	B���؄3,8�!<D��5�e 혔�S�*_�P��/D�|���K0.2X�Q�o��@�V�*D�$Y�n�2��� �<TRG)#D��A�HV$�Z��v
hx���!J!D����,��]9�-�����!,D�`�@mJ;d�b䉗��	D��E���)D��:��\���x#�9���i�%D��k�Ã8L��W�&]����@O"D��!DF����2FO������;D��"G�J<���q4�))O��c7D�`����� Kɂ�K���(�E�5D���P��i��� ���-a��`kw'2D�<2�#��b$�R�-�v��	,D� *��7�����i�V��g�(D��xDd�6�f�
1Iݲu�T�P��$D�L�d��N�q{���a�~-9Aa!D��RхA7A�Mq�Æ9�h�B�=D���!�Ĝ`�b��Ʉ�8�R�=D�a4����25 ԱN�\��l%D�f�\�b� ��TW'b!��>D�˳b�'g9��W�Q�rx�bN?D���N�3��<��@�F�4�'(>D�� *�K�>*(��k���E�6�&"O��c3�҆aKR�{�\	(��`"O�dq�oʴ\�
���1uu���!"Oޜ�0���
x>�;��tb�m��"O���qgA� K��o�\4��"O�=��-�lJܢf��&Z�)H�"O,}Ƈ �X �ɐ�02�"O�]��dS�A���*E��-y��ԋ�"OZ�B�A�9 |2��e�VK�
�PV"O��{�&�)tw��$C� �@��`"O��P����Px0D˥�!����g"OL��W�H�!�@(�AL�s�tq�"O�!��K�`L�@ݹ_�h� "O�L���~m��x�l�dcN��P"O��щ�o���@�	�M��H��"O��B���.BŚ���J��
h�a"O؄�$��2*�.i(�	Lj\��ц"O~�{cȃ3z�,"w��'G�`#�"OT
�O��e��3��y/��bR"Ot؈�Q��E: �[�Q1pQ+�"On���/�
8KX�@�4@ؽɤ"O��@T�*D��(d�\�B0�`(�"O~�D8]�l��ԩ�R	�u�"O��ZqnT4t�Fi�ǩ�j��d
%"O��p�%I��^̚'��#v�8 T"O&� ��vw�0�� T� �`�"OyP0��T``@ɯ,�v 0�"O�qS�"�^�4��s.D�m��P"Oy���k�<���L)�0��f"Ob�"���C�z���MV�k�Ɖ1�"O	*�]~u`ɣ%M�;ͦ���"O�\2�)d�P��[��Bu!�"O0�S���#Y����j��Vb쳶"O�	07�^�R0Hp�7��. (Vr�"On �VnH.���;�OT�3#�-9�"O.h �A &�mїn�|��""ON���a�:i<;f�RP B�"O��SV�$2��D�Ŧ�#����"O�8�K�DP��Qr��d�5"O�9�"�Y l6��@��R|�kR"O����T�Q���3bO1"=K6"O��k�IJ'�x��':�(��"O��AҤRǤ��`�.I�2��"O��ҕ�Q,�:�,���"Ol�
@ᐼ�Wh�v�B�"O���W�GY���鋥p|Ը�"Old��� �@�b�Y���#R؈���"O@}9��P�B,�K&���X�9��"O��y ��6�(m�@���|�ࡳ�"OB��A�(,��d��[��Šb"O��h@(*vbpuY��:pv��9g"O��yя߷Qv��J�5D�X1"O�=xuo�
i� ��-qjq�"OT	��cx0��=9�Ġ�7"OtU��IQg6@낁��m}�Ӆ"O2i"4)݋��J͸����.D���sᑳO��,kQ�Ƒn�b`��)+D�|��f�d��r ���`p|	�qi&D�X2���q0��*e��.x��i(D�L0�k�&ZeA'%}�$�2D��Ig�$s{
���\ ch�	x�0D��1r���=%.h��V���+F�/D�X��+7v�TcB�ҝ)䍳��,D�k��� u$)��ϔv�A���-D�� �ѡ�і�x��2G�)`�tDy�"O\첵��N�x8������r�"O�I��bAZ8�P��'(t1��"O.y�%,��7���
���,��i!u"O�2�G�6t�ɪ-���k�"Oҽ�Bۈ7��M5C=Q��q�Q"O�҃/N!Ocv���X
/��s"O�5!5C�M�<X�a(�v�ے"O0-j��M���*�C�Rpa��"O���a�)�j Jϗ�Q
�r"OV-b%�V�E�$m�1�X��"O�5B���H���a�l��y����"O�``��ϬtTlJL�7� ��"O>h��E��7�A�:����2"Oƴ����-*��RB!}�%)�"OT�PErě��R#z@lh�"O�e��
5�>���eM�:O��x#"O�D�%���5��5� A���b�"O�r`*�����:u��p��"O`Q6lF�Y�f�I%�I�/�I("O�t
a�#;�6�<��r�a���yraN-���Tf]��lJ����y"�ٳ9�"��#/����R� ���y���G��Ƥ @dm*�����yRJ�3�,�x�"Xy�}	��yB+��u\$ȶ�����5�й�y����^=�LP�-E�����B���yr�7#�b|3PNV�N� �*���y"�i��hJ��9P��"'��y���0��HC�-٠K�Lܚ��H��y(��;xBuRp�>p������H��y��4�����J��*�y��
�ydQ�&����KD=�.��h���y"
B�"�Y�1	U�1m"�)�j��y5��7K���ٺ�%��y2&ɔ~��-�U�N W�ē�eL��ybm�������q�4�H��yb��9��)9��
��J$����yB�̻G?>FE�Ld�b��ɢ�y"�ˍx��ˢ��E����jN#�yB�O�݄X�/8U���4`��y��\�Z�	�fN�?���ȧ-��y�+�X�NШs�R(2x(DS0!��yB(6�,uxī��,l�B�e��y"�ǭjZ�|��a�8Q��������y�a!PL��	�I<�9c&L&�y"��[���q�[!,��JW.)�y��/����㌈;R��I4a��y$�5c���Y7bٹF�A�'��yrh�5�f�����;!h�*�g�y"�ǘM�J8��œ4/�)4`��yr��&I���ibDɷ&�4��Ƚ�yb ބ{1re�̎$�.�B�-��y4�L]¥O�(FP+ �3�y�aQ�Hl�\#�k�5��r�!��yrmW"#'pEb�H׸31L��#�y�-�30�4�jf%P�u/�=H��)�y�mܝ~�Z���
l��h��W��0?�-O�I�v"W�	�`)"���[�H<ST�`��������D,6&.�`2��~lB��`�pyWfER��D��i�
�Jb�\��ɣhY�aB�	�X��8;D�Ph">Y��i�>?栁�#��IJ�����T)!��H,��� ��L�����KO<��7�S�π � ��f��2� �*%�lZpO��v�V�G�
h�bZ�:j�}Z�GnyB�)�',���a�c��=�!�2��|Ɇ�II~B»$���3�F�n�|b���yR(�~�Ĵ��InU�P��+���y��=<��EAǡ�+m�؀ C?�y�^�z�$����a)��1�	�,�?ً��S�Y�ژ@�m�\%$Wp�����f/)ck�$RX�@���C�504`&�O�㞼D~���%-4ЅA�lɒ?�0�W��D��䓎��|%a��I� |z��[B<��*OJ�.T��!A��V=����j����D �S�Of���7�9~�8))�h�$����'U8ٲD��(Uށ�f�:~}X�������9�)�'K�*8���[qD�lV7H86��'+�x�U�S�=�f�z%��2B<Tq/O(��䉵b��@��%�$Y�*l#B�C�1O��=�O�rj]�Ns�t1�[',v)0a��y�˥v�2�zF��9NbL�+�8�0<9��d��D�@�3�c?�i6`��2V!���6S�d� F��46'��`�<�r�)�'k�~�pP��	��ܪ�ā3qL
�s	�'LJ�c�`��AC��bd�^>|�P���'E�\���8Um&8k3���+ X �'�^xa��N�TK��R�6��%��'΍���Քv���µ�K�j*� �'_���F-3||�c�F�(<��'������-&��Q(ǁU%;�>����'�!ۆ�9'X%�6
�:C
���'F������R	���6%<N�l�	�'�@���KQ��{̔�9�x��';n����?Q��UN>�z1��'ʦ,�&�>fO �a�gI�j���K�'�E��dU�[�5x0A��b�U	�'���1�&9A��Ф�9V�[Z�'�|Q��T�U�'���^�6y2	�'�g�Zd�v|���ݬF<@a�	�'*�!��*
��8t�Ա8+n��
�'$���[0`����*3<��p
�'�:=ʤ�)n�d��Q"wL�aK<9�]��Z�lݢq�<��5��4�� �ȓP |�8�B�-<8�%c�8]�T��'0a~��%�n���<qef��g��>��>Q���y�Z�z��bKчk{�0[��O�����O$$
דm^A�S�Z�p��D+����h�tD��I?H�6���'B18�Έ4�~X��'�Yפ��h��I���-��Ī�'��rg�b��E��癮'W��a�'����l�2t���0e��b8h+'o D�L�#Ҡ �L�B��S�xV.���+�O��O���I�-{��P�v�҅P�,8F�x��'L|8y�D�XӘ���iƀ[>����~��U�,�DS�i˜`p^�!�B�;�y�F� �bM@��*U$�� H���O�v� ���;@�]�������V~�'F2�� UdD�1E�>} Bdc���ybm�XD�����vľ0R����0<	���'�~5��J��sR��qMܬ5e�82	Ǔ�HO�t����'��A1�Q�?gb`I��	y.�>��d��'��ai���%����b#J@��y��L� "'�=�{�H9,�.�R��$}B�xb��	�E�q�J�/1�L�w�|8dm�n���m�3j{`eW��#c�~��r�VR
B��19`���רZ���X�S�;{����b��� lA��H6"��P�7�Q�k�|�c+<4���`NE�v����c��A�����3<Ov��}R琟BJ������O�̼Br�Ϳ�y�.ɒ1'~A�_4�8*"��èO,	qB&ҧh�j��s�!;x�p�Z�9Ҽ��q�$$lO��0f�E�\ �BP�2~H�>����	�)qZ��E�ғ��q�m�\!�$Z��8� �mX*�����M�qX!�DČ������O�:I~P:"
�J!��8j��y�|��)�A�P�Ie���fx06�
�6��
[�S��:�"O����~��傪k����#���{B�'(��%��Sgd��&�
����	��?ar�iFt�*����%{'�-D�R�'��:�"	���1�T�� 	Ǔ�HO���p��!��e��ϭK%T��"O�yꡎ���eӐ��O\�rW�>IT�)�S�~���w�,"��y�圊*d���d/ғu�>	���ˠ ��ۦ �B���ȓQRi�����1L���t��[�J!�'_�F�)��)t�Uj�7 ����f��N�JB�Ir�6�s�&A��\$��Gn��"<Q	�*XM�a� �ȁ]<~�5�ȓ5� x���d�\`WIN8��i��-�,��g��m2�KE%#�F�E}�;Ox�|d�.`��2�@�h������@�<I�fZ�H��y���v6c�@~�<�E�/UG��S�|�0�D�P�<��p�T@'n	q�HL3���N�<��@�u������X+  DH�<!g��	�2D�@MP�Ǥ�j�C�<!�'%|4�GƏ8��UJ��H�<��iA���j���'�0B�JDF�<I�Ɣ�_�ź���KW��3�Vw��hO�O����I�j�!��Ӓ*���0�'� ��5��&�d}Cf�!��u�-OO���@?վ�j� �^Ap���$�!��;� ���_bPa0�"L�t����>y�(2E��A᝝xxjpp�eqX��O�1�$e�w�2�0gW�a���"O�Q{ӌE�LR|�&ؒ
 ���"O�����O�yP%�]:��L�e"O~\��1�]���/氰jcR�8��	;�ѱ"��<�D��͚/@B䉤�����쌟n-����"�6=����M��h��P�l�#g:�9D N`�j�����V�'�󉉈b��Tr��Ҡ���M�|�!�d�<��uɄ�29�p��Sl�8ǆU�ӫZZ�S��?��b�.��T˅�^�ln(! ���l�<A�C�`Ā�(�w�R	��c}E�,��D,�S�d[*��cg��Ia�(X��>�#�� P3@<�.��׬A7*��;D��:#�R�LF����c�*>6�p(�D;D��R+آK�)�'�!߮<ST�8D��#���v;J�Ν�!�	p�	,D�<RN����2�H\b-����n=D��V�[�pZ�
%"�0z �Y�&.D��V�N�e�\���3m4a�.D���f�Ճ9��� ƿb�I �"*D��:���,���!D�	��ȋ��:D���M��c�ni�5.�#Zy�l�r�,D��y�kQ'|y����#!��;�*,D���ϭ}z��k�^��#$C(D��ƣ�|2�
#�P'?8�-���;D�� j����ճ)��%BE��41�A�"OH��A@\D�j0��<J�Τ�"O-#��ڞdVT�ˤ�ŕ��5��"O�]:F�\Bs���ԋ:sشh{�"O����*N5<���	��,�kD"O�(��]�i P\���Ԑ�2�"O��b4	���x���
I�6�"O@�D�E^�n��
C��"�+�"O�I�D��[y`���ǖ���1a�"O�`�WyQ�x� J��Qb�"OX���)7R�I#���/z��P"O��X�gC�	��E{1 ƈ ���ZW"OQ{@NʠWN�s�P�"{�LY�"O�����S�-T��p5-�ӈ5��"O����#�e끪:5�Xe�3"O����N�(~��&��[��(R�"Oz�bA7���ť["6��1r�"O�)�,Ӌsn̻&d���b�"Ovi*7%��{;�tI�o
�����r"O�% PF�(4Y��iۤh;��"O�D���B�:iI��(ڻ7�9��"O,��$�D��1I��
���t��"Od8J����2��2���!KZ4I�"O�Q V��4q�
���I	:XLQ�"O�\��b��p�
Lv+p���"O4���бN���d�U*�4�A�"O���%Os\$(䈍,d
h��0O\,��'�E���:V`׃=�����	M�I�jV�fi�qEɁ*�<B�	�`����P e�A���!&B�	<d��(H��߃�A�P �9Ee>C�Ɋ%�̥���4E��	���ޥ��B�g��嘶B
��ux!^��B�	�JO���!��iR��E�_pC��::w�<:�F[(A�Ċ�{,C�	�-�`5����Aft�F"
,;��C�	�;T8Z%��<P�*u@�
�bC�	גg��sv��`�V�?z$X�"OpPBt���q��5r2@��I2 �@�"O��b5o�$|��Q�@Ϫw�:P��"O�0�ፅ���aYЉ�p�"�q�"O"��*��{�@=�-�<@��4�D"O�lYT�E�e��EەW�h(�a�"O�M�c�0?�RH��� :ĭH""OFig#�R��@O�M��:�"Ob9#8B��`�/S�t��UJ�"O���ʟ�zp,%������y"�=
�X��1�I$=<�P(�'
Z@k�b�9f��s�8\e��'�*�Mt
�K��+0|��'�����ή{���5��j�j�'�x�1�мYs�8�'�K_�-��'�p�3r���B��N�A�mP�'�n�8V��.j:|��R�O-�]�'b���e�S8���h� ��K����	�'$��g��:�ph	���VѨ	�'� y�ϊ |^�X����2ZzB�'��Pq��%��B���@4T:�'��؀�\�s�\D�"���xۄ��'�`�ȶ!SRU`����$X� ��'(0��`�-,����4JˊQǂ���'���9B@
j~L#
�qR\x�
�'e�Q��%���&Ui������
�'�F,���K	p�р���t�HC	�'!0h�t���2\E�W��;c�H	���� �D�� ݞD"<8��J�dzB"O��`	J20�XI(A"�q[8���"OҌR�ȝ��A� ��0ۦ"Ont�3cX/^�Δڑ�E�a��X�"O�l ��9��-�&��-_tmJ�����#�ʚB�'���8�h
_J<�Jw�?9JR��ȓ����V�9�L�c ,��͓8dѰ�耥m3ҧ�����O�3:IX��hMR��yP1"OR)����vn�Y��������W���6���	X�B�.S_��)�
B�l��P�V&��$�7�O�4 !K��G�4p�tn�c�I!�GVm����4��N�C��^<��C�Ɨ&N]��U$R*��=a�a�|��X�QE	�ҘO
|�����D��f��YG
�
�'@H 8�KPad��%[2/�%���2�
���Ɨ�P�1�*O?��2/�N����,B��4���bg�<9��'y;r D&Ȓlv�$��by2�И%G�顳,Q@�ax"�v����/��0�8������>ѕ#�$��91���w�NpC'E���`1����8���a�'H���p��'C�D�3�#Gz�����+�4 ��)P�&�b>Ia)C.��|2��~W���$c!D���0]"0���V�P�T�1z�$�e�C��f���>E����,_=@�J�R2z,
��@,�y�H�%mK(�y�C�Oz��������ɰ"�����_MX��(p�PV����` 0�(R`%4D�h�B
�
P����}��-�0M3D�#�H#b�闢/# ���,D� *5�(e��"!�DR��j�l+D���p��$5���5#_9명�ei+D���g��1bb�p�뛭d0��v�7D�8�H\(k{`Ƞ!�V���F9D�L"�d�88�@������-�rO3D�<�R ��U��1�U�5��j�A3D�,���\->�E���hd��r�-"D��R(����B�-}{��A#D������K.���D%V��\���-D��!�C1hܨ:p.!M'�|JK*D���j�7:������̐m�Fh��@<D��PPGIl�2l1!M(]����:D���� c@��A��
��bޞ;��"&$ިvzӧ��BΘrZ~�Jp�J�S\���f���yrˍ�VZ6(�0�^K*�D������y�%���䅙��Km�y��*IMR!Sn�J1���R�R��=�4I�/�&m��IT�K�<�#�͎�N��IzA�Lupx�C��3$�h0�*7��큥��,!��v*)��4B�^���#d
��#�	�$:Ժt[����b�M�7!򤁴"*Up�J�*2Ꜥڤe�(T��"Sr�̙r�n�j?1���O0p�DOY(rZN`i� ?b@���-D����PYנ8y�ʎ�0B2�R3��OѨՍK����h���+��<�k �5�\�S񍛖v��J�$]��`A����BF��a+��h�Z�Ԧ"4�B�[mM�=_T4���Ao�$�=����'�B��2�,X�T>�v����P0�K$(T`,��~JS)}��S/T/���Q���<��G��<�J�jߓVv�a1�{ݞ�zRJSe7�4J1���&���-�&���1�	WP��4�&Q��Måύ!>!��B&��/d5j���cFB�<A�C��9�<K�H��7�q�#H���9�CN�A���R�!��>��6C��=�2��S����є)��0��/�$<����dN2X��|���R�����GR�@��K-p0�H`�Xފ�6F�=U��'��>�	><��Q�feE�b�$#qJ�
h�>��qq-߄{tXA��IO�i}���g�;k����0+��y�]���C�_����D�4ҚY��&��{+>���ELo��Q#�-�6Yiر�OT�ӳi�Ҹ[!�=?���B�շ�M�
�6g�&] ^�\0�0�b�<I� �<�N�x�׃'�����8����#-z	�ILhv�E �<ϛVDŭK6���3�D�e�2A��
K~�q�'���pdVR��oZ6��T"�.2C|�R�eL���Y��ύ�a�x�-O>`���F�j�1�1O� HT�t�$T��a�!h��6#Yr��$��H$���	F���O'$u�QhI6?!Fr0m�7y(M��bJ=��H��"���<�i��'��m^�8�r�͝{f]��i)f�~�ٵ.}2?��ٸc�"Z���S���J�������aҷ{k(8�@�(�!�[���z"I=A[ I�*QR�bܡ#���{�%A'�A0M<񧨋��'Y���y�o���@��uW���}b��1X���oء<`E2��Y�A� 1t"��^��c�()4BY����ē&�h9����d�rX�#��2�t`FxBf��NH6�b0�	B���0�ٴ86	
G�ˎh]DC�	^�B-q�&(c��᫕�P1�hT���"~�ɡ]P�s���X���k��R�`�XC�I�:?�<���P���CB�uK>C�I^;�TāW?v����g��lVB䉡p]n�{P聪i��U�Q��0��C�I�=$|��ѩ"���B�K�U-�C䉀{L8�y`B?rFD����>Z��#;g�����s�B)ӆJ����4�B�-'�)�S�p1�(4�/A�.�!�˳D��C�ɱr#��Ⲏ�6��!aRe��#$�'�$q��! �c>c��QdJ)Wܦ���Ł<H����6�Ob�31��]ZeZUMU�.8ءY�OH� v|Qx��&հ?q I cT�y����F�n�(�H�j�'I	��%JL?Z�JL�\Ĩ	��A�`,��P�H+%�Ơ�U�'^ZM����g���
��F��&�'��)#DEW�#:Ƹ��>i�,!Hh�Aɟ�m�E&��,���S�EF�-+�A��"O�إ �(�RT+�]��h@L?aP!�̘��'Ddʧ=Wf�#ꄿ��ݑ�V`c��׍QQ�h�S�	�
��$B=AM^�:�%�I��"ej�H	�tE�'PVE��ΐ��԰��!IR�m*5�Q�J�Fy�%�<�nUI�Y�ڵx�bĄ�O�ٻAm��b$�5�}�H���=�H�i�)��Q*�e���=�<�
6n�u�.L8Qł{8�Hs	�	��u �H%Z��؆� h5��nK>�� %�����4A�W�*0����On`��;����f��/���C�5�䪡"O�}��N��������J�� �5h���IH?��$��]��m�%ٟV\��ǧup��
�w���G�@zq)�F�d3&a�	@R���_��&!řk��0�W�$����ќcV�Y����0ij]"��̃}��Y��N�Y#
��j.���6"�b�V�E~b͛S�&Dc��O��{�0`���K�V�=����G�Xx�M�n��,R�E�"�J��DW.*����т��OJH��aGX9Rp�Bˈ,L���DX?��K�YC��0�jE�#(���S(��-
D>�ʶ����k�E��y2	�6P`�""�I(��!bb1�M�&�L ZD����<=JT@rf�Ro����J��O�H�íT5*V=h����"JL���UPxI�� ��;�ڽ	G%��	�=�e��+��p�rP4����2[�n<�P� �"�Z6�(�3$!i���1����'�� ã�MӺ��|�3�Jݠ� ��$#8��[�3�\��S
A�WB�|j"H�6�<��er%�e� =7����Xц�v�VXQ اO�)�,�.&��4�G&Y#S��]	b�Z�s�G,T&e� M��e�<W�Е{bǘ��y� ִ^}rͳ��ߡH�ȃ��yfY�u��?oR��4) >p�A���V5\wj��v%��ɘOC����/I1{@�A�!ʮEf�ѫ�#@^L�r��b���	�?�B�YPO]��0��*�"Aʱ�㍔����kC?c�\ґ�=���fW5(��<�VeY)Id��@(N�ٸ'0BA`��Q�0��I�~"��/hV���pM4c&`�镥ѥc�"pK[�	��ls��p>�2�ɗOZ��!�iC�%�]�zfy!�K�/���'�8خ;&]8e1'T�A��{����?�1-�P\ &��''��i�dj�4j�D��ȓK���C S�~; � �²
��o��uet��o��E�h8�������	�|9"�>��@U�8����,ef�Xf*6|O2��r&���$�{�8��ՠH�U��ya��/�Z,�(�\y��Y.��}&�8Ӧ�O1t�,�:�&�`�f"4��R���1�*�h�,"�0�@���j4��l�0�a}�B�Z�2Q4�]�S�B�i���"��<Y�'P�L�A�͢>�w�m�ލ��ޥ�e���DN�<��eR�N���B�$r-1g	B̓&z9#a牂������U� U�0�Hی�҉��"OR�U�50��j�(�p�2ā1jU YtqO����Y���5DO<�q�CMڡ�����1D��  �Q�:��,)A΍"��iZ@"OvxÐ�&K���DK�9%J��"OHd#$��"y�x��vй�"Of�k�E��+�h�ЪٳE���"ODq���Ch��F�@�8���"O����gT^	j'��j��"O2P��>�Ȉˑ,Q�1�&�"O�qb�oX/_0`e��썑b�vR�"O~h�O�?`g����-�`�"O������q���I�V y��m�$"O
,���4^|f��g��g��t�"O�Ѳ�d}�x�VE�;pT�"O��kf.E�N3�l�D,ԉo$�u��"Oȵb�K�(�*U�ݍQ��Bc"OAC!�NI���JأhW�f"O��CWa�`��Q���	TC�`�U"Oą���$�j9��) ,Un �c "O����M�y��Y���a^�=('"O&�� *L<"M�*�Gގ{�hM�*O� �a���.�KDL����$��'&���I&c:R1��N��!4٢�'�P��D@�%E��ls��ЙX�x��'�="��ݠ7b@���ͺi��`�'�p!��a��a�x��˝1-��'��|��eQ5_d�q� O l^.��
�'�Љ�U�SQ�J�`�	gv\��'��L�G�9�Bh�E-غB�����'�b��q��v�n�
�E�68�d��'�P<[�)�-g:�çn[,
���	�'G��0C�ϤQ_��#r&Y<yN����'7@�Ra�

`$����rSΠ��'U��U�oF�!��G�����'����e��6� ���af�Wv�<I�(ރTb�M�c��:��	'��T�<!�TA-�*�a�?BX�=B��H�<����3�t*q�^OR�H��@�<)d��^*AJ�Aվ2H�@��e�<q�n��}Â��!ǹ�b�@�N�t�<I����*���c��?tp�����}�<��L�/�|L���;BoXy���{�<i�.�?u<���kN�<������q�<AA�*s�i�tN^�V�>���$�Z�<!�C�F~z��C;6��R�[l�<	����s���b�ˏ�0�B��C�<�0A�'wNl0P1��^��\��Kd�<A�
C�d}R����TQS��}�<���3���k#^�i��xSKt�<�QǄ<@�
ɦ��d�1�TN�<���I��@t�L�t b�T��v�<�%ξ9bb�����S�f���_{�<���]�A$�d&΍nh|�@F
�t�<yw��LK�&�2D@��6������b�X5�(]�2x��R�"�F�ȓ!1�Q����1�
�6�>yN�܅ȓA�4�ᖃ?d�K�#�O���ȓd����\ke i�����`��� 8�ȶe��=��9��;y�P�ȓH��9���*R��%y���5}���ȓY��L���K8`޵����2%�q��X��X3�V��@��o�5P|,��!EI���<Vu0�g'7�l��ȓ~^*��G��3�NH����dS
�ȓO��=*v]�g�L9��T�=��r�j��eꀸ^I��p"��r�Й��S�?  �˲��5�4x�ыE�WZt �"O���"�ܼ�pפ�9/$<�#"O�`p��PQ�\@�"E�#c���"OBm�2e�ut X�V���a��,h�"OB�S�F.:���Q�D����|�"O�}�􊅝6 a0���y?.̩B"O^��E�^:�8�!H�P�r�"Oh�0��9�0xZ1ᑙ�����"O���,�3	&�@���x�c���.N��4�� R�L�x����L?B�*hj$�6E�����iB�Px�Nޏs��8���2&vZ�7������"CLҧ��2x u���[|�Җ�iZ�h�"O�h�)NE�����M�,E�icU�l�vbV�5�Y���U���(�%h89��5��]2vF5�O�M�3o��Tp��ąq,�Q�K�e�����Rd�HB��ZL��'L J��Lc��M�z�=�qa�sp�9s�dҢ��O]�|q�]?��Ec�.Ș!�d�J�'f]8�e�!"p��"���3�$���bYX4B�g[+$>�++O?3���>��ip��X�8t�g��n�<�ס�%G��P@��,T@�L����~y���0N�H1I���a�ax⭅�:>��#�I�KZ��x��Z���>i� Z�<�N���\u��1���!O_�8I"Nw�q��'��e��%N*+j.�r_�I,hͳ��䒥i_n}��*
I:�b>q���?[�V9��"G�Z�$|0��3D�զM�z4�5c��6Lqڙ#�r�����t�:|��>E���X7#L��mH-����F�S2�y"#�iXa�GT%�@�Х���ɨH��؁�oX���qF���|rӦWj"Y��1D�@k�ò`k�xҤ�F��I[W�2D�4�V�]�z	�5ڰ�޳q����#D7D�@����
╙�G�=�h��uC;D�$�����R�T�QQ+ܹh�t��<D���n��6��Lڶ[�w�,J�:D��QC�ϚN�41��׸!9:��1'9D�Li���;6������:c��*�A D��(���)y"�X"� Y�L����>D�xs��Z�C�,�p�a�#C�n�I=D�l��"�A8Ιhw
�\,��
$D�x��4Z� YkNF�Y�
.D�(��X�2� MY�^�&k���d(,D����
+��赍S�Y���1D��s#ٺ=E(h��]7���V�(D�8#�]0}��L� �Wl�����Rk��
H��~ӧ����ˌ����H�y��᠂��y���N�<�z��u b&V��y"��)Nt�8 �ҡ g�y�	D$)��=Z�*Ѯ`��q�ˇ��=f��`�d`��ĥ+��� �H/oƀ����	���Iӭ,$����#��l�Ǖ7U"���)��tqpI���0?�5����x�����O�2�(J�CБ]�!�d�g������J�,abS�[&%�,� v阨LŶ4��A�f?����O��q����-B�J��s�̡�"O�|�Va���l�񳅇�
v��?�`)ҍE��й2�\&g2��$��]]��j�a�)>G(AJa��yk�{R$ҥ�xh�w���XZ4%R#�%.� cC���G�ܑB��"4p
Y���d1��(�#�/,��G��%��AYgf!�	3*�� �G�7=*N@B��i��"*
 #T�
?�(��ի���2@����"|O�#��3M2č���)��y���0!J �T�M��8���'orP�T-��jv�7�K5Wd���G1
.R�Qv�T�!�DF�Zi��@S�^��7垏W��f�>$��u`P�~S��8u
ǚ^m��O�ؗOh�qQ�ޜ{�r���*U�@ߓ��1%��Gm�yYr�� ��Ik�	ȫwQ��D��O���aRn6e���'��>�I�V��P�T��$m��s�,�°�lZ� 5S�����:1�v�jR�
�*�`���0���2F*�('������"o������c����K�j�V=�2�L�2�R��FͿ+Y��O��{Z�l �+T~����Z*�M� 橁�#��wl����]*.�U"O\��W"G!A�h��Z�0*� cv�''z"���.㼑2B�0b-H��"G��`���'b�����!�Ɖ�+fԨ��2|m�8آL�`ܛ��@7E��[�B�4�-�ճ
�hk$�=*f7M�: T�*����#e���:\�t���,�O���@��A�8J���0tp#d8=����VJ�+����!ƵUJҜ�s�N?m��{)�L��Ay��8>e�b!R���h�4�t��'�_�+� �Iw�M�YA(Lz�0O�Xz�;1�6QH$F@D?��0`"OJ�x�/Q]WB�����O���*��'�-��eՊyx5�����ē��RH|z�fҸNn`zf�|��4�ť�t��T���_[v]k��i�dl�Q�Y�Z����Rf������&�	>�����L<1tm��miz���)\a�0�0b�u�'Bܚ6H�v��>����+��x#C�G6�؉�#�;D�PCFc�>a�ZPI&K�?5�hM��(�d6B���%�)����T$.T���"��&-�^E��A7D�D�����1�<���ϑ� }c�6D�t;���,?aB%�b%ʔc�*5D�h�ӈ�
m�"��V,L��j0�<D�py%M۾>B=1AW�^��V�4D�D��mW(Y<�=���`�j��u2D�����y����F��q�nA�0}(z����=��Ǎ[��x�JԮU���r'�j�<�!��3p�6�E
�*??��
�$���q �c>c�X0U����@Hqs4�9��,�O�P5 �{�q ���V�2�#�
[�q�G�����?a4.Ѵ$��A�Ù9p0�1r�]x�'���� L�ܑK|
4���$]�%�̗l.R	��O�<�D�I9pX���d�j����-Q?��D�$��e+4�F�����'����6A�Lu�EH���bäB��
h�����L�G�`iBA��e����.Oq�%%�W��Q�J?��w�K4�]��(3l<9kV�)�O�A[B��(�HX�!I�]\�`�!I?:�Z�������DSMv�\�"�ÇS�gG4h-Q���'ϖ.^.Tx��p��f�~5�f���$9�L���C��7?�Y+uH�7a�5I��
2zkv��)A�L�i�Q�՗�h���P
�4Y�!�	-}~�z�"O8ݠ5�8#�J�)�.�;`E�{4�3?�D] rʞ �(0��b'֦9�;���"43��S!��p?�c�[���Q1�?i[:�s�D��pi�RG͝�B��*j�R�(�'���1ʃ�q�R"?Y���F44� ����� �H���΁".�H1P���y"��Z>4�hcB�2��9C�J�R�>`��c6$��1c����F��'�p���TbM��@�6@X���'�"�x�g�z�µ�����)fe�ڴ�x�/�8�p>iљEg������4��8�/M���aW�Ō="B��V3O��Ag��|s܂�W�Uw�qC"O�]�шC�!��Ѳ�bllL˥�DK05>�͂s,Z�ǈ�qJ���

����P}K�Y�d"Ox��ՎF9,V2<��*�&N�lŠ1��]�|��B�>��(��l׫�<��'z5���%]c&�q�E����Y	�'��l��)Y���� �ƭj\@J0���hvh���͌�h���f��ɧ�O5|
`�C(B� ��'�@�~�	"���!S ��G����{��l�E
ȶ�����㙌W2�nM���3�x��O�|s�4�p��FL���rd���_\Zb$&���h���b�#M&8�|���X�nB*6�Lғ��6�>���ش�.%"��<���jބQ{a�r�����i��2�]�E �!���Ǿ&��D@E�J�t�l8R%�t�!��F�O�0e��G�|Y�lأ�W�G����'.w�鸆oq���R蒌��)[v��Wʕ���PJ$ʅB���$��uC�T �Ot���ePpL�@�&f*�h��F�y[إOP p�,�3}"k�ג�S��C5$|V���ϗ��xR�˾U}�c�BQ�[�@��P���A4��uǁ:r(݆�I`��X��E2[_��`�,O�k����ŲYY�Xм���'2����e���0a�OB��.��	��� L���,R�8�8�˛`�:���b�0�&�$��1kDD.�:Y�L�b��<=�ڨ��Na!Deۄ9�zHI�D89���4�Qr�\�|�'��@q�U	��+� v��Y��'IDex�Á��2�X�2̒�'߶|�0�� �24��dG [��z�'J6ʒ*K�i�����iΩQKԡ��'Q\|z��
]xjh+v ��S��=0�'P,�R�%�?w�t8��Ԣ����'����		�AŊ�de��<�q��'�r)���sw
U��a��ȇ��'Ć�3&���qD�5 M߀H��'�"� �!t2�*Gʔ+zah�'��`�#�G�H��j�ʬ/�,��'VXiK���=�X�nm^��'8���k�c8B��j��M�Z��'�@2�+�B���1t�^;)�E�'#J�
�H?'�,��0K<,.h��'�^��ƪZ�	� �*�/�XlUh�'�ZM� Ádqdb��!|���'|6����� k�Ⱥ���':���'��i��AlE%�aR��'D�l���-6�p�Də�J�կ:D����-�.��j�M���6D�TS3��Ϣ�� ꍌ)��e��8D���@�R6{;�����<8���J�)8D���ʝ'(8l����5�iK�h%D�$��L�t9��:�jڐ2y�����/D�(f�U,K�Tɋ�$�"�8k��!D� `��� ���GOԡd��8�a?D��3C��#>#����EYv��F?�y�A�X�� ɂ�Ҽ=��j���y� L	I�Y�S▋��8�3�
��y�C%lhL�YA)A��M�rH��yR��;y�){e�ͮ5XRu�n�*�yb'Z1P)��"sŔ�)�h�
����Ohe��f�<����ѥH�9O��E"O�PP�Еz+�q�S#B14J�"O�P�
ʪr�:����89-0� G"O"��*݂�H9*fb��h"� 9�"O|��T�X�&ؒ�o��%0"O��r�o܍e�uCP�H�$��4"O��cD�,!�p9���)zX��"O.Q:7d��j�eNYQJ�\ۆ"O�4ja���Y�4pCʡrQ��J�<�2� D��c���2ZB��(E`E�<�4 +)�^�q�2'�2 �D��}�<����5������^{�ux �D^�<�`+Y0G���C��L���f�c�<��%�\�,��rir�xp6��b�<a�%]	p�їN�"V�ؼ�R�g�<�Sd�2y�d��5��� �VCa�j�<����ڊ��c�� m嶸J�Ś@�<ibbƤM�L��̎�<�^8:��X�8�"S�@���M�'��7^f�ː"ԈF�A�'�F4�?�u��1(@�`��Y|�l@��#}�A��eKvf�1o�������� 6df���&/?E�.L�n�Z�˃0KԠ��6M��p Q��)u/�8�'��O`���ځh��#2���0�^�\��Њ]�<5*���>Y�j��0|�p)@?_i����9�)AgZ�� ���&J�O|��ْtW���~BN?E(ֆA�SЬ�*�eŨq���۵MblP3=OT�W�:�)�S�{֊�b�
�F$`P �><D�B�I�y�(J�Fٌ7�Le����0��B�	'I��b��M*^����0��(a��B�ɕv�"ȹ %�+P�<�U�d/�B�0o��D�Q#�.@4�Ġ�LrB�)� �d��ĴS��(�� 7/�I""O����
d�p�R�o�"�m�f"O�|��@.��|SE��"�����"O��E� (��:��oDR�:"O�h9���[�pd�ʙ��x��"O�� _�a�������)^.(x�"O^��Bͦ	R|s�b��*[(8K�"O�q+��Ϛ>��G�ΎUL>�!"O�	��D'R$�C�OkS>uȳ"O0���$s]JF�$x�!ӳ"O�{�b�8��-_?�a�R"Oeq�L�LVh�6��`�"O�t04��r��,��E�p���3�"O�l��`-�~����$sE��`"O�|�N�{�4���N58�5"Oa� ��;.���iCE�쭰�"O��a�i�@��]�eJ�T�� �"O��S�X�,����4k�:���X"O<aCdFO$
^ƱG���,0E�""OبqS�V p��P�Ń&D��!hf"O��W$ܩX�,P��0&5�"OZ�zg��:���5��`*�"O~�za�~�̸J��$S���"O��:7���5)��B��-!�$ǚ�h9�a\�^Ub0{�@��K�!�$A6=�smP8>Q���#@�:&�!��X�jtX���{<��f/�81�!�7Nt��f�-�u�o��!���i�]�5g "�[�Ȃ�n�!��G�p�fN2W���S�&�!�آgfڐё�4���\!�ĉ�nK��ţ �D�a`  D"!�� �^]\�m��JHġ�3IM�<!����L��''\�:B�A��
�?�!��L	g]B��SC��d-2�
>�!�
!�Z�§
,j�@�` ק8�!�)�pQ��I�3
y��dI�3p!���yg� �цV9{W�؊T��)e!�D	*2�楪��DML�	w�N�b�!�Մ澽��D��>��Q�n��g@!�D��<!��F�&9�#'(� #!򤅕�2��o���"(�?!�dڬ+=�\"B�'�D�s�V8!�W�v0L�q��݆:А5�Uk!��3GdF0�u���!p�C?X!�DȊOK���f�ؠ/�t@딾8B!��
D0��t� ��]��J�&)�!�d^:c�P���)��~�l��')Z�Y!��ˍf�@M8AE�/)����IA�#
!�O=b�&9�X;b�6�y��1\�!�$� 2a��ȥc3ڨa���G�!�DE��V����A�_A^�"��D��!��!��9�#C�K_�H+2���s�!�$Y}�0�4GD40R�I�Fې2�!�D�68�x�3�ŉ�o_Ve�G��l�!�#]�Ӆ��-/^����^=;�!�D���h`���i�X@F̛�Zߡ���.k+tJ$%��L�VI���yR$�U�$R"�+[Z{"Yb�'�����,R
>6�i��C�3U�V���'�f
'�!CpT�4�J,Br����'����T M0F����Ά�4xft0�'u6��۰9�x�&ؔ��e��'�H(�U��&�����JM"�t���� Ly��JV?Ő�8��K��4�1"Oڼ��J��j�~�#,�R��a�"O�8C�N�G Vh�� VC~ @�"O����!5NF�|���N1ffQkV"OB��Ο���� 1���"O�lA�vCPг� �c��6D��ia�&0v��I�(�8���5D��"&�I4l�� ��EIl'fș��8D���"Lf��X�2C�6.{�`y5�)D�l�VI�x�\(:�G%A��@s��(D�Y �˒ �x��.a��i{a@*D����L�-7��)R�7I�U�@,D������-�Zp�QϿ{��z�b<D������D
2��^JJE.D� ��`ՀUK��p���v�v�hDL,D�ܒf0�0�?	a4L���4D���E�ؕ'�Y��FX1 ,x�e�0D�Hz�Ie�&�k�DD9��,!D�t�Ы���T4���y��1�a D�(z@`�S���V.P�r��kF�<D���%_*P���������� �>D�܋Ԇ3+���	�
�H��Rv(/D�,��l��C{JT��M���"/D���-ŞH:V� @���I҆-,D���0�D�I�t��$�(Wy0��(D��	a,Q=u��50P�d�&/�*v�!�$�&-)���E�\e����Mۏi�!��� N "9je��>"�	�"�%%�!�d�4Rɴr�C�9nذ�[ ��,n�!� �"�0	�"���ۗ@O�a/!��̊i��q����3��\�So.�!�L�h��I���
�T��ar6�@�/!�O) ���,Y�]�Ƽ��.�$�!�$E�8^ɡ��9St�e���}�!�D�u��M�Am_|V���A�z�!��f5� DJ^?<]�z�'��Ux!��G�l�~p��O�pL p�DL�pr!�D�?s�:L;�I�i�w	c�!�dP�(EV�JF���^��т�@��!�d�X�0�(��A��fd�7��@|!��8/J���X5�dq��$�VB!��
	<�[tcM�Hu�{		(!�䟾F1x�ҠUh���D6,!�ڦ='� ����
������W'!�$�[�6�1�a-. x�hV퐾7A!� X���I�,ݦv��1�➙)6!�䂳$���"V06��=׏�"!�$OY�L���>d�|�1nҘt!���n�"8�'͘Y�@i�#��P`!�$M�=��2ajM+�j�X�	��|[!�D9al0�R�^N�]��&ư�!�$�4G�{�d�&[�|��d$�;{B!�)A��y2 I KȈ���LL4e@!�ė0(\���k��P�05x�œE�!��A�̠9��i��q�Z�F�!��ѓ=��H�!�Q�d��FiU�)�!��,HȔ;f��[r�-�U�ѽg�!�DT�@�&��eN�Wд�&��.!��W9{Y8��cUp�y�O��r�!�c�ԈhM&:��t���!�D�� ��*$'2��01D�ɟ�!�Df ��r��^@�"��`���e�!�d��#�3V
J2��-J�J+!�$ ҍ�Hw��!��Q�{!�� \���M�.� `�Ңr�&� "O��CA�F6�hy��!@ M肤�"OPq��.
��1��N]`�"O��j&N�L��t BnΥQ��zF"OU�r��Z�B�)1MH4bo� S�"O�xi�ȝN�uU�ϱsi���"O���h0F�+�ʗ	1[����"O��`7�ǃ��8H�iJ�}Fp�ђ"Ov{d�P)R�n1��.֋q@�$j�"O�(�G�B�+�rIr����~)���"O��d��'VLJ.@ٹ�"O�PۧDü/pNX�QP�[�"OrD�F�{M:m2gH�/BBlq�"O� b��#$����P��1<'��r5"O�`�"��eB��� �X*T�"O�Ы�j�&P�Q�`I�@Y(r"O\��5���p�er��53F��"O@-�߳G�5���7��#"O���Կ2��@ �O�0� ��u"O���僙�&��<���ʸ�I�"O�����$vd��pU���F��"O����<vbث����Ͱ�"O��%@Ыn��|��J�ˤl�"O��M��EX�eڐNb��)��"OX��gMġ\҉R��$��<�v"O*��bn0<:�C�����-�G"O*��` ��,ԐPM['mZ�]A�"O��r��rу��I��	�"OPX5iӃp� �S ���
prw"O��C�$�A=�1���!,k�"O"(r�'ĸ5a�x@�c�� �r-@G"Oh݃��U8��2Y�9=,��"O��[@M�	J��)�&ݏ>�x "OX���IU�3l��4T?F���"OȀ�3�F��B1���Ѣ���A"OD�K��V��)P�,E�~�	"On P2j4U�-��
�UE�!�yReZ�
DM�I��CN��y�M!�Q�G�7u�U�F��y"��5G��k�
K�F�p�h7�[<�y��b=
���7E��Xf`���y���(G����a$�<<�a�Pj�#�y2/�,�N�k������͉�y2�H�uV6��a�F������dL��yD�6e
�lxP��gf���uM��y�	����E�����Y/�y"����f�@v�	�Y�\�cO���y���xڠ���<�r*�yr!�SLx�KU����~���+��y���O�e�*�:5�a��J�y�e4�$��-��0��9 ��@�y�jJ�Kl�P����=�H�$����y�ǓJ�ݪ�dX78z����\�y"8}t ��d��8/q^uz3�Y��y� �sc*�Z��)�\�ђ)�%�yR@��1:�t:��%*E�& ��y�Q�S 0 �l��;A\Y�9�y��M/xq�OG�8x|�pE��y�"�<6E�boQ5v,1�X��y�G�K�p��̍='I��0U��y��;r��1��U�Q�d�Q��y�<9��1%F�TC��Sb���y�(�l�<sg�!�����C��yRaϚq�!�4��>$��W ~�Dȇ�S�?+�ş   �   �  <  |  s  �)  5  <@  K  �V  �a  ,m  'v  z}  `�  ��  �  4�  v�  ��  ��  B�  ��  �  L�  ��  "�  ��  �  R�  ��  ��  ��  K�  � �  H �% - �3 %: g@ uD  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�Y�G{���˾R5$�Qb+�jBƅ�7��Oi!���l8��Ӄ]*W>�\����]O!�ė��ތ F�8#"J��7Lb!���P~��#���(%l�(.ԜoI!�d�0c>��=`�r$,�
�!��LP!���6HٮsX~��!ݺ�!�Ĕ�m��G꟯i�̥sQ �W�!򤃛]Q���D�o��Z`A03�!��R�6j�l��B�^ ū@��;Ol!�P9��$`b��e&Ī���c@!򄊡jX�QTυ#i��A(PhˢF"!�D/2��`pB�]�6�`�6��9!�dEE����BݙB~�tK�`I�W�!�DV�=�i�H�!(^n8�䏔$g�!�$��mMX���9OT���n��O�!���-
l��WoР>J���NE�ni!��K�4�VYP�ɑ����+L�xT!�$�4<{��J��! �PhX6*ʨI�!�Ff^��PR*C�lʹ����F!�ͪ&�����'�4j�\���(�8\!��/�:��������bN	i!�$�<PⱫ��53���{J!��@�S�vL���?ʀ4sW��*t!�DT��`Iȧf yƬ`�c�]�#�!�D�p�,l G�.x��ᲆ�T<@Q!�@7_�����=�"|p0��-N!�"F^�cbI��i��,�g�:'�!�0�@1g�żm]�,�Ҭ�
3�!�d����(�qKrأR+�<q�!�ںO`�i�눏`�p�5mܒ<�!�d?B�>�1f��~�>�#���0b)!�$C6h���@焐K�и��)4!�� 4IAI�R@`�g� @K�C'"O�ِ��3|�V9Y%hS?<v��"O�y���<9�t��'��X=�"O�a��Q�/k ����$�Lu��"O08DF��D��6.M02㼠���5D��")U+e$l�ȶcX�6���Hu*8D�T�N�,N�n��4h>~��ǈ+D��@� Aƒ���eT�VD4��%D���q'�
1��Z&�Q�9h� 6D� ��a��1k��T% ���J)D��(�f�4��US L��1�z]���4D�p�3ϐ�ѡ��R/BI���&2D��I��.��s���p�� -Y����@�Ta��ցE��1 �oÓ�y��SZh&/\�SIRݲ2��y���(@��Sʀ�9̸3�j#�yB�ZM�z��?~�t�>�y�NÙ[8,�kWG!hQ�\�C��+�y��/����C�úkl�Y�-�yҎE G���롃�f�P}��eɱ�yBbӣ6OI��G�s�@�a�NI�y���(�=�"#�1lu�l�7' �y���8l<v1C�G͌eI^yD犠�yHг w�Ժ�=S]��������y�c�'�8*QE�K߾ț ���y�]*�������9,�ٸ o�#�y��M�j��D�2|¤{�G��y"#̽���h�A�a�Z��1Ů�y�)�s�0	���\Z�����yr�	z�H���+1��	Pj�3�y��XZXt�-�%`��ʤ`%�yR�IJ�P�����XWI /�y2���U?E���Ԍ|�j�!���y�c'�V��p�P��Bh7�J�y�:v% �𥑮r?l�i��y���T[�)Qg��}�`P1���%�yR���.���8�C["#�v��AOV��yBn�b=�A�X<� ����M�y�eD�_"J���t2a�5�̂�y�*��X`Ht���:�xED���y���1�J�Bc�"��,zu"OH5�5����\�B�ʄA��=��"O| [A�Ȯg��c/,�,��"OBy�hP3&>(��AI*�H�s"O��Ru���d�B�@(�&���"O�j�"�	�S �W�0�P"O������n[�}���>K�Ь�G"O���#��q�)ڒ@#Gt���"O��S��CT'��kR�Q�11��)@"O60�«�j_���hٶ4#�"O|P�d�I�j@@�2���4�,"O�@S��W���@�����TwB�(C"O��C�C׫Ix�Qi2���H�X�6"O�ɱ�dZ�{��ͫ�/��	l����"OY�!/\  ZR��BHW)+pD�ٗ"O�q�@C�lx�#cgިk���P�"O�lK�&T<T�����o�t�2�� "O|iA�,���٧��#&�YzU"O\ȲX*��9[V�C��|@r"O�-�Q�j ��	���`V�lA"Ox�ۡ,�:m�d��qJ�i��h"OD8bC ��\��c'/0f���)V"O� �/<]���z���F:z!�E"O^���'�����+�"ԋ$(�S"O� �x{U�jHXAY�̓v�x2�"Oࡓ�O�B"؈ �Z�6�1�"O�Y$�ِ$���RS���>-vd��"O�����?Kr�HA���X�=��"O4A$!8<���M��L�`��'z��'��'7��'��'��'tj�1���<w���G�B���'\��'cr�'?��'a��'"�'R.@q��y�|$�QՁx�ځ g�'��'~��'��'�2�'���'6�0�M��
���U��1�� p�'�r�'n��'R�'2�'���'�Dq���+K>��`�3������ş�������џp��ݟ�����4qlڌ^Q�<��W P�t�ǂ������ԟ(�	���Iʟd����\�I������Ԫ�^�h�c�I���3��P�	�����ޟ<�I�,�I̟����h�7ɘ�!���4&��W�����JΟ$�	ڟ������	��	�$��̟{�f\�`��<h�c�� �x|��iP�������$��ƟX��ٟ��	џT�����I�Ε�!�����P��
V����D��ޟ����@�	���Iʟ��I��|�&��D�d�r���>�D�$������ ���0����d�Iß��I��$��6&��,H��[�e�6!W/_���ş��	џ��	�t��ȟ,���,۲�%M	����[�ТZ��Y�������h������	����7�M;��?Y�R��"��8a �i`��0k�	۟8�����d�hG�N:`pLC¤׵����&K����_3�v�4���O>�&��O+
ͫV�� Wɐ�����O �$ڛl�07-+?a�O���5�$�<iZ�]z�)�=U)5/�)��'T"_�lE�DƷ�h �a��8P��u 6m�0�1O��?5�����@���b�h5��k �;gᕅ�?1��y"R�b>iѦ�S��Γ6!���֌��u&֝�$c�"~b���yrB�O$,��4����-Rg���J^�fL����]�)D�$�<AO>�i�Z�j�y����ة��V�U����b	��]�O���'���'��T>�05Ù���fѐ\��b#1?���bj ���FF̧bk��F�?I���gb2e"��F6�E�� ��<��S��y�,T��Sv�n^0P@�H��yB�|�!qӝ�@Rݴ�������y����\;]��Eh�D�,�y��'���'N��1��ic�	�|�#�O��)4n�!
6�%���w�=å�X��]y�O�r�'%��'3�i�3J^�<�W�Ւx��dC�B]�R��	!�M��V��?����?�M~��}�n���G��rS�4`�ǻ�Nu�$[�������$�b>yr�O��0f�X���
R`�3x���mZ|~�*Ȋ]����������;�
�j�#1�0��$�.;qf���O����O��4�|�
C��Ǖ8��-jN��	����!�3fc��t�*� 8�O��D�O��$��I_��ఫШ1뤔�'b�1\�Ĩ(%x�V�!�,�3s2ʧ��KT�S�U� �h- �c��0��<Q��?A���?1���?���o^�Jn�9�F�U�_c�hh@��8a���'���l��8)6�<a��iR�'�aI�� 3�@�x�ט~u\��P�|��'�O���h��i?�ɠDҨ�L�6]���"uIР��~]"��+~�O|��|����?	�N�
��S�l����"�C�Hb�����?�,O@�l�e�j�'R�Y>9���%�X��b�H��6�cw� ?y�U� ��۟�%��'6����'��ec�t1�O�p��k��Uq��,�޴��4��i��'g�'5�a(�F���|�cv��]�v�rv�'T��'o����OS�	�M��L,���b6�O�s�T���(1z�����?!��i�Oة�'t�d��8��H}�Z��V���'��Ġ��i;�	�f�:�����&�P�Ju&U�Ev4��b��fu�D�<i���?���?����?�*�2��GLؘh_̱�!�*q,�C� ��I;u��� ��Ɵl&?牟�M�;L�I�l���BǄ0u4��Ο`��z�)�(p40�m��<93Hڟ-����HE$P����<�"A�8"�^�DT��䓢�4����"X
�h�(�dZ]K0��/�O���O~���<���i��)��' "�'��|rp��:D֐yR��[��9ѥ�Du}r�'���|�\c�]�� 
���1ሂ��$U)vy{�`�^c>����O��d��G`���
�y�:��d��!���$�O���O��D!�'�?��!�~DŒ�O(:����?i�i*Z���'�c�X��]�h�=��J�ce$ٲpĚ5�x�����	�� ��Gצ!�'�,�&��eʀ)SF�iAL��lJ� C����$�O���Or�$�O��	�b��婒h̎$��PE��B��)�f*��R�r�'�R��d�'�`��gfG?IAn�#��[�~�Q�O�>	���?	M>�|B����L�jq�q�Ũqb C�_�CҌ��4��$]kM+�'1�'��	�$@hq[��ᐝ�g����D�	�$��ݟ��i>9�'G�7m�{����2F����� իmP�re�������?yZ�@���|��4ik�4��@S�(��(��#B���tB�����)�'�20��m��?�}��{�? ���2I\�*9l`���:rP"6O����O���O��D�O"�?u�� �-$1��@U*`e�!w�W֟��I�l�ߴ;q���*OPunf�	�2��	�@D2iM�[ �	%���	ʟ�/ƘmZB~Zw��Q[d��\��ϼSUXy��nٰD��L�g�	py��'�R�'���K�jz��׫A�9�@�@�pr�'��I�M��	��?1���?!(��� ��ׁl�|���_'-9�������O��$:�)rf���t#�&Y��N�X	�g�챂��_?|j�eX+O��C��?I�A$���(+t>2���(�Й��O.N���d�O����O���i�<93�i��E�b���Z���J��	�t4��N*��	2�M��J�>y��j�ё%��|���gR�R���?�3����M+�O���v��)S���B�8���2���8��U���ςrH��<Q���?����?a��?�)��pԬA�:Vn�b(ܚa��9�b�ͦUі�
myb�'s�O�R&m��n �k�l��ǂB�����47����O��O1�|�j&,u�6�ɨ;�*)� ��2n�RE[pH���c�,��۰n��d*���<ͧ�?�v �-��P���^O1R�I4��?	���?!����N���E��������,J'����p�ZԫƟqh���b�Mc��h[����l��]�'_� y�e�0lD8cG㍓���`����W�(��|���O���OD��3�֥BlR�i���/0�%���O
���O����O$�}"�MDd��5L|�Y�-=��I��G����/<���'�61�i޵C��ìZf��+t؛4,!�w��æ���ٟ4��mU�9�'fҨ�t ��?����5L��(�)����pJ� [��'��i>��I��<����4��"f�`);���5��v���)���'K�6�Ӕ~t��D�O���/���O��k�+�	�j�r��a.qKG��x}R�'�R�|��T���K?�4+�4P�`�`@�l�ݘ�i
�˓����n���&���'� 1��`QRq�䊶��
]lc�'_��'�r��dQ��;ݴ;4�Y�:�&� i�B��k��&Z٨��:��v���d}��'���'mژj"iF�Yd���e�^8� �*ڃ:��6�����ǆ6��t�	��Hɚ��5#;��jP����5O��D�Oh�d�O&���Ot�?E�-�;C��j5��ؾA���՟��I�P�4�n�ͧ�?���i�'h\��C.�!�%��$��\�uI!���?���|�#M���M�OҸ ��g�И��D�7FrF��al
 	x�Q�'��'���`���	.Q�*��H�D�ԣ� �UR���ϟ�'47�[t��?�)�z���)�0�VT v��%� �R����O����O6�O��;GM,��a
F�-H�q+&�V`�d�st�B�>LvD�"�ey�O��,�	�"��'�ҁ�`Ӝ�88�a���O Ɓ��' "�'��O��ɷ�M���O�T��s��X�(ڕb�,�0X-O��o�o��^��	��0`�ȷ{iJ4j�� *U<}9�oßl�ɹ�$�l�C~��^������W���\����a$x�a�i�)��$�<���?���?���?�+�5��ّP��5;���9��y!�	W��a��"��������8��ŵ�y�.4&�}H�7)�H3��6J��'Bɧ�OO|��űi�d�<"���*�c`���!	�zi�䎭b?��q�' �'��I��@���*T%��#����ƌ (N���ܟl�Iן��'C�7mVG����O���,��"OfaWc+�p��e=�	�����O��d3�d��s�>a��M�\�N��]��ɐ8D;F�P��|�f켟��I)#f8d�~2�t��@ʇ@�&�I̟\��ȟ���G�O'��O�*����	,�r�#��6U�Al�1�E�Of�$�ߦm�?ͻ�5B���)̳�nuɶXA�4Oz�D�OV����*6�$?Q�[2*WX�	-��zQ#��2ڜ�js+­e}`�xI>a+O��ON���O���O�=������P%���˓�R%QT�<ɔ�iӸD���'�b�'��O�"�?4�ai�h��zb( �f�2 J(듆?����S�'|F1�%��JCkT6d�N1r ��MC�O�JĈD��~��|R��	�n��zh"7A�Aj ��Dܟ�	���	ߟ�Suyblv�(I�v��O<8�v�Y�]i̝
��\�Y�3C�OV�n�y��a��Iោ�	Ɵ�j��@�" Y2
KH@�D�O E�J�mZ`~Bh�>���'��ֿC����L�+p�	Z�I(��<!��?���?����?щ��
ܟM�f��Կ�E�N� L3� �럌�I��iݴ��ͧ�?��i@�'Z%���*��T�'�Ŕa#�ͰՑ|"�'c�O�@�/�MK�O<�J���6a�*�	���-3|~0� ��2s�h3�'��'s���h�	ߟX�I���j�ƴI���PӯO6.% ��I��'��6M^.j�"��Ov�D�|��a��_l��V���V�6���ECR~2�>����?�M>�O����a��>��MQ(7�� C�N)�\	�#A #s��i>McU�'��y'�����X�!ؕXC�*.��d��K�ğ���ş����b>y�'V7�r�RT;Պ�<n$u)�#X�?���
G��<���i��O>u�'<bK�."�T���'N�M�d�P�:v�'���13�i�i�=ʦ���?e��^�� ���ʃ��u��MC�b���zC5O6ʓ�?)���?���?�����]�@������'�Щ���W2>e�m��Ti���'������'Ԗ7=�������K��A@��N(�Z�A��O���8��iT�z�7�j��s��A?"��K�SM|J ��-z� �#L:Dt�$0��<���?1Cb$�8��H(B��8H"K��?���?����d�Ԧ�kf��4��ڟز5M�.X����FP�{)�u�m��zy��Ο��Id�n�VY��D�m̺��W�ѡn��4��u9"��9TȀ�|j2)�O܀��_�N9���s��,ї��3(W�A3���?���?A��h�r�$�e� x�-�66܅yU��,���Φ��r������I��M���w R�cBFJ<
:<��ϿS@-8�'��'B��	�E�Ɲ�����P�iF�D�j��r���a6��$ �1{���O�ʓ�?9��?Q��?I�l��D8(�*9����҂�%V4�2/O��n�3\��=�	��(�	\���D�q���P%�Z#O�4O�aCu-H����O��D;���M�|l���7�y���Z	O� ���Ҁz+�M8,O8�S��X��?�7�9���<i�$�����l�9��y�b�>�?y���?���?�'���yQ�@_ʟ�P��͆A�������Q��l���{��	ܴ��'��?�-O>��Q�Z�X|��9t*H�y3<�ȗ�!'�7�=?���Y�
�h����'���c�KF*i+��:���H��Y�<i���?A���?Q���?�����(�\���%s�B� ��^�P�2�'��(b��+:�����!&�HY�hռ<�|ѳu-߷p�8d�2h�V���d�i>-��i���'S�Z�#[ x�2��c�{��-
 �E72�	���䓙�4�x��O��dμ,
.Q悈9�$������b�$�O ʓ~����\��r�'�\>Ȇ,��@�fyY$b$kH���??��X���	��%��' >mQ�E�<��,�!Wu8�[ "�$�D�k�4��4����'"�'o�� �M(��<�2,Ƌ;��E�F�'�r�'����O�剗�M���*1��D�3R���`��>u4�+O��l�]�3�I��ĸ�.Ϝ=�mۃ�se�cU���ɒK��m�d~Rg�5A��4��[�	�.�L0�/E�X����n+��<A��?���?����?�,�h�I���> ��
��3f�V(��@Ӧ�@������	ȟ�$?����M�;B�v�Q��=(�H����*gG#��?�J>�|�A�+�M��'�����)���;�N6R�R�'_�9���y?�O>q,O�	�O�e0���j��^���S!�O|���O��D�<y��iX��'�B�'��Ї%X�>;>��VD]�Q�����D�]}��'�r�|"�v���z�i�y�3#�Y����Ә2�(�C�Գ[�4��, ���^���$#,Dɐ!.��AGKN �d�O����O��&ڧ�?�EEݼ[�p�	���?E � ��ô�?94�i�\X{"�'ج6�0�i޵!�ʈ&h� �
�d�4r�xR`y�h��Zy"�X�TU�f��HsA�Њ& ����6�v�F��4��T	v5&�$�'���':��'k��'����_c�,�D�-�B�r�\�H��4*��i�,O���,���O���6!X�p�d����.{Z�tjդ�_}"�'�r�|��ԥ�4 Pr'+ѥuB呅14+P���'?��6l���P%�'���&���'z3F)6~,\��!�'/ ����'�r�'R����]��	۴5�hq[�N
Zd���9��h���G8�$���K��V��`}��'���@;��+ n�;Sΐ��Pc�/�R�ZV���'��J�E��?��r��4�w"@�DE,uo6��� _$A"��'L�'>��'"�'Z���xV�����S��#3U 	����O���O8�nK�6����|�P�~�b�n�"a����"��)��'�"������'ԛ&����Pd�2�c�<��a�̥(��Z�����|W�<�	ߟ��I۟�zd �Cj�R��X2Mh����4��iy"�c�vm���OB�d�O$ʧ/�`�Ӥx��Ya`E�;-v���'����?����S�4f�\������W���1f���vbF��� '��擟�����6�D� !��Y��-ήF�������l���O��d�Ot��<�4�i㼔��#Z;�
5Q�f��'&����9;剂�M+�"f�>y��P��:Aɖ j~�B��8$�|
*O �y�b���� 	Q�F��$�(O���2l��b�j��6�U���#2O�ʓ�?Q��?A��?)�����J�HZn0S�
�������Tn��~@�	���	U�s�p�����s�ې;��@����;yg������5�?����TOO�YK�v4O(�9��� ����9c�x���=O��/���?��>���<���?���F�?�X���&h�5���1�?y��?�����CȦ���LƟd�IƟ�8GF�1w��I!���,[��N��Q	�	ǟ`��E�=r��m�\3�bC�-��6X��	[PE�M~�3'�ODE���K�X}��������!�B�?��'�'���S�x:��>/�|	�#�q\đ��� #ش�bp���?�W�i��O�.C7�i�A&	�����c@O/.m�$�O�D�Onaʑ#k���qyzp��?� �����-��SLߵI��T	��$�d�<)��?���?!��?�0@�;80(���Y�EB�i�ɟ���Qʦ�1Є�˟���ޟ����Ży �X���@���a-_��I���L�)擉\I��ˠ#&�*�b�L� 4�Ȱ�Lꦥ�'�J8�dB?�L>9)O�i�A��8�pS^���D�Ь�?q���?!��?ͧ�����N���`�7Z�>�Z�&��1se�`�'�S��X��4��'>�ꓣ?����?�A�X�9�H�+)C��E�ఖ���M3�OB��cF��(�t��Ԁ�0;�$��^p���m\��OR�D�O��d�OH��4�S1C�-���N�J'��dK�@R� �	ӟ�����M��|B��N����|2l�#Nu�T�SHŅ���sa�-��'�b���tB�<*ƛV�����:D>������fq�!�g�œb&6�K��O��O�˓�?���?a��~g<�AC�ȲU�z"@�Zw�$���?/Om�Q8��������o���ȗ:��ōA&3�`��������C}��'Hr�|ʟ�H��Ř.�z���i�j�9�d��H*��h�(_�LI�i>1���'��&���(ð!�E�3�*
�����T�d��ɟ�	��b>a�'�\����6�RJ5��jU��J��A�Q�'�b�h��8(�O
��3O2��I�V9��Pw��h�&2��?I�Å��M��O�mSO�O�t�&�,T�\�ё��tMH�H�'��	⟼�I���I����IV��'�
L� �鐣ɴC��Q1NB�,N�6-�0*v���O��d.�9OAlz޽�׈Պ^� �-S:46�9���러�I@�)�847p!l��<y7�%�h9����y.AQ�<1���"[����1�䓢�4�����*3����ɝ�.���	X���O���O�˓p����̓���'W�w�$�p�A�hx��I���O�<�'�r�'��'�){�(B�pԊ0D�ˉ@�.��O��I�)��7�!�nP���O`a ��!J�5�FQ�Jx�w��O���O(�d�<E�t�'ᦘ����6��l(��5;o�ar��'f~7MB�D2˓DQ���4�0Š����1�$�!����~YV�QC=O��D�O�ZB�7�5?�U�_z�@?,ڑ,#j�Q��A�f:�X��K �$�<ͧ�?����?����?�����\�Nyc��_������������E�c��vy"�'m�O��i��Um��PP!�!D�0ohj꓊?������Q/o� ��6���}�:p���/�M#�	�!��I�w�Xt�g�'��'�`�'��t���]/j�* ³ ���P8r�'[r�'7����dP��شV�<���lo���VJ�>���`ac�Y0�����Y����d[i}��'���'�f��w%M�Y�(D�A�5ղ�`��&_�6��Pˢ��#Yi��?�	��p��^B�ur��Q%gOp�(0<O����O���O���Of�?1�s*�zo�Y�2�82���{���,�IןX�ڴ-.v1�'�?���i��'b���ڴTCV � e*3� 	�y"�'P�	v,��lb~2&�'AҺ9a��S�8�``�T+�`iP���ҟ40��|�]��������I���0Pcլɢ ��#]� u�u����۟(�Ity��dӎHȢ*�O��D�O,�'qxL}:��;����R�:(�8��'���?����S�d���O��(A��KWo�mr��?����t�7N֛擟�ӦK���-�ԮR3"S�ϒ��b��EQ�'���'����OV�I��M���$/z|�����tA�֍�l% �y#I�<Q4�i��O��'�Rb��h5�����5=V:-�E�V��剠$�llZJ~B�̓.d�H���\L�I�"8�����4���"�T"
����jy��'�B�'�R�'�B\>�H@�e�&X�̺-c*e�⛒�M��ŋ��?A���?�K~R��X���w��f�uT:�r�(k���'&b�|��dc�t�?O�J��)l�ȁ�ՅP��PP6Ol�L^�~��|_�$�	�������N�~<x���j�.���k@ٟl��՟ ��\y��uӌ�jPB�O��$�Of�;e��+ ����Ǜ�gcxJq�&������O��D;��Q�n��|S��!0lz��$�/Ft�	?B0ؼ#�Ŋ�_��c>�+��'��5�I;Vv�Aj �e��t`�I�<��������������Q��y����z���a���0��h���*A#"�y�2�Q��O�������?ͻH���Ŧ�9^�8)9�BR6K%^e͓�?����?��OF��MC�OȨ��M��������U��D�U��.�xb�'E��؟���(���ɯI�����m-T��Y���0�^zy�`}�6�`�<a����'�?��iR�$=�t B�*y�(Q&�9(��������`�)���H)ϐ$"{n(**�@#����@���Y�'? 5@bˋC?�L>�-O�hIq�R�N@u�$��`���M�O��D�Ox���O�)�<i@�i��i�&�'^F��GFE�*��D�q�I�w�Fl؟' P6-5�	����O��D�O��y���_��j�	��e��"��Z��7�9?���V"-���!������do�"ھd�AI�4�ޡq�fa�(�	��IΟ�������"�!mNT�`��vW���@a��?���?�v�i���O��hӸ�O"���2����EDY/5u�y��.#�D�O��4��qEoeӨ��|D� D��c�C+$˾q��Mע.V�A�b.�.�~�|�R���(��Οs�䈖W�y�%��%8زٱ� X��0�Ilyr�h�J�bb�Oh�D�O��'U|v=!��ʒ^�X�t�C�2*Z�'�4꓂?Q���S�DɎc���'�U�.��H# ����0��A)p�X]j�\�據�ҩYa�	/R���f��\Jb!p��>^������	ǟ��)�SQy҈r�Ƭy�/�8&�y�!UYxPsg�*G���d�O�n�B�����Ɵ䙇̔�;F���p+F8�T��S,Xny��?�������
���M�Hyr�T�t�=���O e��J�I���y�X���I�T�I����֟$�O����U,
Z�p��/C"�jU�nӊ�pP�O����OB���D	���CK��`���u$��K�cP�2����ԟ�&�b>s§�ئY��Z$��3��9�%U>(͓D�,��si�O�PZM>�+O��O�����;}�0<�q��^�8D�O��d�OX�$�<��i��0��'Z��'-�݋@"x�}S ^1:^T([���J}B�'b�Oʱ���Y�P�)*���G��Й�$R4	��i9�i)�Ak�h<�����ॡ�;'��#7��X��`�b�ڟ��I�0��ڟ�E���'n�4��ѝ0^�Z���7�%�'Kx7C�ʖ�d�O�mP�ӼC O� �*x������q�͇�<���?���j�n��4���F�t`Bm��'p2��a�,��~�<0ۣ)Q���Ó'?���<�'�?����?Q���?����/ZY�
�	nfJtd����D䦩����p�	Ο�'?y�	�c�ܭ���#@c����.�ʀ(�O��d�Op�O1� ��éOJp�i;�Ȕ>��]RԨ�A�i�Z�t���K�Ƶ��'���'�d\AN�.z��!%�sbvXC6�'�b�'����Z��H�4w��$C��oM���t ��]JL�t�Z�� ���&���A}"�'o��'Ά�G��h����8N��!��yN����rV��6ai�)*�	��Z����Ֆ ,T���~}L)CP9O^���O����O"���OT�?�"2��1!���P/C�'����L����۟t��4>�lϧ�?YP�i�'��9�˫��i(@(��sWj�pV�|B�'��O�M�¸i��	'e�����^ƀ	��)<hp�:(þq���`�	~y�O���'�2���)�ҍ&�̗�t]Jd텅x��'��ɹ�M��o���?���?�.��d��HeY慛��Nd`�r��l�OT��=�)�A��y��!6�8�h#� �L�&nݗJQ )O�8�?1D�-��E�L�T5C�HBm�  [�5(��d�O����O2��<��iL�аu#W�'�	���b4�H�Ci��[5�	��M����>��i����gB(�cOE0:�
Q����?�ӂ�(�M��O��3Bې�I?�Y���L�d0f&R?^
��yD}�8�'���',��'L��'5��_�صrB��F���C�B׺a�E{ܴ
��Y��?9����<��y��G%b�I��ׇ=|���U,ӈ#�R�'ɧ�O�j]���i��bQ,�B������t�r��3/��-<*h���*��Ob�S�jC.in\P�7(��a�&�r����0<��iS���'[��'79�'�#AW�	1��l�25�� V}"�'��|�z'iɃ,�18����2L.��$Y�:�B��	�MS4��d��R?���m��3��:��m�Rh�]�\��w�ma��;e����썅\̸L��8_�f-���!�M��w�pA( ͞9L*�r,@ 	��9!�'P��'����&J�V����	��%���F^�
��h8�B@�s2]��|\�8Dr&�g�!��J+6���nA��dU٦�;��������ڟx�*�/:]�� �G�+8�5���&��	ٟ\�	e�)�ӈZq����
�`�j�R�HP��5�����.O�0`E�K�~�|�U�ĳ��ݏ}.ĸ"�$��,�h)��%�O~�m��p�R��	!8��Y�LkE�x�R�לVǄ�ɂ�M�2f�>����?1��:ʭQ�Z�<o��P���>j~<ە���M+�O��)�l��V+&�I��<�qOL9��C�&C��0�;O�����d�D��7�D>?�%E��6�d�OV��]ަI!�5z��i��'�Q�s%��mOb%zᇎ
����|��'��Ou\��Ʋi��	�`�d��OϸP�l�ڒ�I+�A�r�A�Z���<���<1�B�
�Uu����O�t9DphG�J��OJ�m�a�Tŕ'4�Q>�ñ��9`�Jq�2�)k�	�N1?��U���ޟ�'�������N�<F�^�F�Y�I���PL�8&lUC��:��4�.����ꢓO^�2CJ�����$�+;)<���O<=n�%D��+�׎b�l@ڕBA�v�R��$�����	��M��i�>9����;Ԁ�6��`�>������?1��^�MS�O5 ����U����i;/Z.-�kɾ\��Ӈ+k���'��{�C��c R��f�w���Q��)|�6^�4�����Or��'�S7�Mϻ@Бa'"�% ���ZPbN;������?J>�|J����M뛧� H�@��L�BCV����W�w(�(&>O��*6D(�~ҝ|�[�p����0��.
�r�҅�`��/?�S�#���������	qyb�z�v<��'�<Q��:��$�shW1H�4Ja�6<<=����>���?YM>	u'̗�p����@�� ��Y~"l
;� <�p�i�ғ��EX�'�g$"v�1zN�7uЉ`@�n6��'w��'���Sݟ�P����w��e ���]�"LV̟��޴��0���?���i#�O������[�(�:_�V%����d�O��$�O6�Bd�x�~�T	��Qi�?��JĢ_�,�ĥM�] YyS��B�	Cy��'��'J��'M�Bʱ}��vhͷ<qΈ�b�]�j剭�M�aM��?��?qL~��e�yʲ(ٺH<���b�ܼ�rV�D����$�b>u��$�j���h �E��D��zP�o����dF "����'0�'r�I�m��p��bC!Z�@<J�n�8�9��ɟ��	�L�i>Q�'��6�Ъy����8
/r�Q�Z�7�P�/ �B�B��ݦi�?�eW���I蟌��b�f%H��S�D��� ���*v��ئ��'�NT:t��?����t�w�4�=WFR��p�V�t"ސ8�'B��'���'%��'h�2�97�J��*|[1n��i+6� ��O���OԸl�9���ן0��4��l�X�{łG!#4��X�L�b��=�N>Y���?�'e[�dk�4�����٣�Fݧ?�"E�jЖ�@'�"m���������O6���O��>��83+�2�����~\�d�O�ʓl6��@b�'^>����FC�Z}`2%]��n�`�u�8������O��)��?]����&���+�zV�����SJ�Z4ī��O��ᗧ��E���J�|b!I�Ga>�9��Y��b0[1d�F��')��'m��^��,�h�!!Ꮔ4�&��"�PT�@D��;W��$�Oȸm�j���`�O�G�k��S�daL���	�q����O��R�ai��w��U��?�'�ƙ�RŞ'a��q�`\�L�P8�'Q�IX�I�|�����M�t�[�h؆�S�w�Ms�u֮7�
��x���O���=���O(�oz޵������E�Qa ��LP��"[��l��D�)��&|â�mZ�<��P$mXi�w�W"�\����<����u�t��������O��d�$�i"%�ў_����Q;%��d�Ox�d�O~�U����ݮ���'R���!0�&�R2W�|�GC�)]�'\�M�>	��?�J>��	8N�6�S��W0�&TJ��t~�ٹ`���g"��!�O����	�!Z��F�qA�x��a�.V7�J��	�
��'Wr�'P��s�}�r�{�e`Qa4f��A�f�ԟ�8޴\�"H"��?1 �i!�'}�w��b˟�|}>���.ۘS�e��'��'���%��&���]�S�y��*!&~����ׁk2�,[0�לz*ԩ��|bX���Iߟ����h��ϟ0��O�\�4��&qT��
&�y��dӔ�����O��D�Ov����$·c.��0J�.�lׁ�1�T�C�Q������%�b>��%���D6�a���{�ɉ�="�nڢ��dN�l��1�'z�'v�IjC�]*�kϳ@�U"�	̣Y�����ݦ�8!�OϟD�U&R%���e��XJ��$�j��A�4��'���?����?��,� ;^<���&��8���P;xD�؛ٴ���n�!���`������J5���bL�f5�a���ޚ<��?�O����E'@����!�8�,� 	�<�> �fC������ަ�%�Ȣ� �B��}HgJ��$�� �Gl�ޟ��i>��a`ۦ��u����@ A&�A��IN���B��,��|�R���?�џr��ih�����4�x�'��6
~����Oj��|�֡E�(��}��J����;S��}~2ǵ>9���?�J>�OR-Cp��(c@<�L=}
Z���!�"nR��p�i���|��J��('��)T��u�T3���/��xRT
O��nڢl�d{է��a-�M t�#0}8mI�&��l���MS���>���
�T�d�۰=�n��Ɗ_�ح����?ٴǒ"�M��O<��4�M���d_�<��&��"�2a4�P��e�	rk�Idy��'��'�R�'�V>�J�]0?	����vE�1"pg���M+�A5�?����?M~��r��w��� ��U���kD�E���'@�O1��H��ff�T��5g�V$XC�>�Vl��N`���	�%v0<��
� }8�E�)^���)���
����&�Q�@ �D�'b��(y�%vPR�䐇<A2	�+���������=/8�)�#Z1O�t�B)�1''�1#`Y���y<�(F��'3�(p���/,��	�f��,.�n�5�9�X�`D�Dq.50�jT�PGґ�C�
����h�5IT��&W�yM�IP�����T�KT�%{C_�>�xX�Bo�+C1�d�� Z�M%�����:s�@5��c-%5ʬh�+��L�����Vf�e#����o��y7�#@����b�ݔ�,6�O��D�z���!w��o^��ͽ��<n���P&�������Pg����O ܸ��)y��9�F����ıi���'��	��l|X������OH�� "R��4�]6�L�)�eT�a�T0$�����`J"'�K����h��g���pD]�1G�Lk��3�M�(O��i&��æ	��Ɵ��I�?k�OkL�)O ��t��0�f$�S��J���'�B-��ub�|2�� 6�0��H�Jʠ� �ߍH�LEa�i&�1�%y�P���O@���&)�'���-tV�,"i�cZu{��V�r�J%Zشr��������O�"/�	6�@��_h(���X�J�7��O��$�O�PA�[x}W���	?Y,	91�N���F�s����#d�q$�ȳ�J�<��'�?���?AB�NX�F<��h�(�����$F����'8%�	�>�(O�d7��ƺ|�p��7$�Jȑ$��,/`�	�[���Ծ8�O\���OX��<qd@#W�l MFAt��J�12�\�l�'�R�|��'�r�J�Ph���T�RJ�@��G�@�%�G�'
��ӟ��Iɟ,�'�6�
T p>�Q�L� �Qs�*\��H[��qӖ˓�?IO>I��?	BPt}"�

ɴH!E�Z�@څ������D�O��d�O��a��Tk�S?9��

'8�hp��w�V0�@�ڹ|̖�Z۴�?O>���?�����'-R�*��IsF�PP#_�y��=rߴ�?������ſS����O!�'?�4���Q�X5�D�S:�]ʠ�2BOv�d�Oly���:�IPr6��>�0��6�Q�<ڶ�#����'-����j�@�d�O2�����ק5���#A*��b�`��&�i�F��Ms��?�®<��'q���c"b�7Q9� d�	f�Ř��i���	&Lj�r���O����TD%���(t��m i�&��E8��y������M�)��?�W�Q&�ӡ���W�A�����';��'�����4�4�\�������ƩZ� ��MM%9��,���rӈ�d+��e��Od������Gf+�xx�����. ��ye�q����ޚY6�~���m��2�! ����}�"ɱ@㍧EK�����x�n���$�Of��O�8#4ș�E��w����
56�U�5�Ϝ=^�'k"�'x�'j�i�U��԰3�
{�^ x�>l��{�F�$3�D�O"��?Q�D����t�(�V �T��)vb�X
 H���Ms��?1���'��Ix�7M޹P�����'�a�YY2�
J?��ܟ4�IޟT�'�DpҢ�/�iT�_}��j��S" @0��7p�Z�l�p&�����t�'�'=°��e�ԣ��P�`E�.�Pl��D�'*"`Ȉa��Sߟ����?�X�G�%8E�K�M���`�R']�.O@��<��V��u7���	(sL�e��������d�O�p�u��O����O��,�ӺK��o����KG+=O�T���ݦ��	Sy�I���O�OA̜	A.�F��颴��-���:شvz�8��?����?9�'��?�	�LC1`^L��A�-Hp�4�w�ϛ���J�w��b>��� `Ή�rG�&'��s���F�1��4�?���?�w��#׉��$�''���,.f2t֝6�rxb�l��~���'B�'�\�g~B�'��$�!I��[�,S�qvm+AlE�<��F�'#4c$R�������L��I��~u"��#�z�إ�A��ēL���<	�����O �S��iZ�AZ�j�(>��=�2�	?T�ʓ�?����'���O�(���7"��;�Ęm�*b�i�I��O��d�O���<Y�!R���ӊ,��:�iٔJ��Y��G	W��IٟT��u�	Yy�O�B�ݱ0�d�	M�0P|d� HN0[���?���?�*O�� WOⓌ"5j�Sc��N͚�a�=.�����4�?YM>+O�i�O��O�Z@�$g�&�� !���2>�Z�4�?�.OV�De,"�'�?�����N0�b��j�Z�1���=l�̐%���I_yҀˬ�O��9f������D����;hG��\�LSuDԵ�M�tT?���?�P�O��ʢ�U18ǌ��.ŵfJ-�M�*Ot�d�O@$>�&?7m�i� �'ة��<bR�R�k+�6b�� X�6��O����O&�	V\�i>MoڣT�F���#Y��X1���h���'���'1ɧ���h���цE�$`�L˺W3����
^.�M��?!��D���-O�Z���An�����t�z�C�>�f�Gx��(���O>���OE@%�ڞi�(ٱ��(�1:�
Ц]�	ߖ���O�ʓ�?q)O�����h�fN5I�B�z�ύ�Iv��+�i�B��y��'D2�'$��'�剔kG�U���mxx�Q�)Q�	�5��Y����<a����OH���O�͑�,$k�EC�/�<Y��#g��,e�	���	ޟ8�	y�d��k޾�S�p�@�SPmʵXGHP�Gϗ�|8�6��<1�����O����O(T(�>O���5F�q����@ʻ#���� � զ���П|�	Ο�'��H���~r����h��!ʍ0�(p�"��	��K��M�����O`��O�ԣ2O��D�O�(I_����
>�r( �)ǖ��7-�ON�D�<���Ԥ[Y����d�	�?=�Ł>|C��]7g�M���8����O��D�O�)�6O��O��S�B`�A:%��}>4 cf��47-�<ar�P�a����'j2�'d��c�>�;*Ϧ;b�Q&4�\�]�@�4,n���8���Y��	F�	]ܧ%�L�M�:= ��SOL���4}�zD���i���'"�O.����d�4-P�x��iC4\�ܰ���:�l��l���Yy��'e���k��3�@ ��tsU�N@���o�<��Пp�#����<����~b�=5�x�h&F5YB�-c1.��M�O>�g��<�O���'*Z� b�h5�U aT�8HwQM�aQ��i��������d�Oʓ�?�� @܁RFB��S�� ��#���*P�'�ᣞ'j����L��۟��'f"���
� �BI�f�2��X(�]
qG������O�ʓ�?���?	�#����}����"m����C�4�N���?���?A��?�(O:���(P�|b���+NP��a�9j @�IUƦ��'�2P���I�0���6���CL�))�g������
L3m��@�O���O��$�<�u�S7&��S֟,)G呲f��2�'�S�2�"�c߱�M[�����O��D�O"��4On�'2 ra�I"q}��Rg!�(SG�,)޴�?����D�д�O�2�'��E�Yﮁ����4� ��W'���?����?Ajc~�]���'H&��������=+�!ݚ5��Xlby��(�6��O ���O�	�Z}Zw�&b<��B�)̦e�l���B֊�M;���?�f
�<I����3��=�R`D�Ȼ`�r�Є凥@�H6 o�(m��@��ퟠ�;���<I�"BM0�
�dƻ:��H��Vw���h�����<���t�'�4�`�M0�� {`/3;�����sӒ�$�O��D	�|�0}�'���ʟ,�c��'AI<'�N!
Fj]�r�o�۟ �'��K�����O��$�O��Kv`��[����pc%��P������	lL[�O8˓�?.O:��Ƥy�E%��z�hY�����z�A�A\����Ee����Ο(������y���"0���BҢ(�|�sf��4VC�0
��>9,OD��<1���?�i��e ���RP���S!+�J��a���<���?a���?�����1�ͧLYP%�=3�L����<�>�l�hy��'���d�Iϟ��Ʊ~F��"L�h���C�'r@"�s��@æ��Iß��I��'��e�!��~j���7*ɜ)X����ۼY�A�W�릡��Oyr�'|��'>>��O��I�3���1'�-h���*Ǩ�"@7M�O��$�<)�͜��O���O��in�0=ѸA#t&�9t�.l�E�0���O���ٝ
����:���?���k�-7hp��9(�ݚ��l�~�=� ���i���'�?����I=P�68C��
*�94��yY5�i���'��r�'��'�q�$I���I�R X��"I6b�v�Bb�iN� �aӊ���O����-$�$�ɅM<P�����XP�d�#R�7��"ڴw��9������Ox2
ݝY�<XRhV�L��r��ئ���ǟ��ɮ+L� K<���?��'7��ЁP�/�f#�K�UT-�ڴ��g��|�S�$�'���'y� �Ǣ�DiٳCO ?j�� G|��Dӷz���>�����S7�,��lڷ!Α��L���v}be�y�V����Пx%?��ӭC;v.J��6�$3f�ԉ9�8���}b�'��'�r�':Zt�.ц ��!����Y������?��]�|�	ҟT��wy�(T�`��S�d��f��X���ø�,��P���	�t&���I��z-r��S��H�>��X� *�m�px�����Oj�$�O��Cj�A������O�={ڨx�$_D@ఊ��1?I�7M�O��O��d�Or��T?O�'�ШB����#�����'ܮl�ڴ�?Y���Q	bi�,'>e�I�?�B6Ӆ\b�|!���cΔ�����ē�?!��j�< �������K��dbe�
�]ZBiP���Mk+O&Ż �Y򦝡��0�d��l(�'r:�+�eѨu׎��R�nC��x�4�?���	,�?�I>��t��8�j��r.ԋr��iF�
��M��-}X�F�'h��'[�$`+���8Dt�2��ф41�5ka��3I,%`�4zg�Dϓ����O b�\�"�:庲�S�+o\	��dR���7-�Oʓj(���/O��?	�'r�����0[���蝫7�U��(��OF��'���n��hPS�+[$IQ@��:`�"7M�O�1�eeRd}"/�~���?�K�X V@Ǝ��	�jQ��X�1�d4���Ov�D�O���O�%��X�xU��F��1�Qg�4�>��?A��?yH>I���~�J�?V�F�ps�C��u�t�M0%	W~��'C�R���I1�"9��Z|ڨ0�m�o�p��ӆA��P�n�ٟ��I֟p$���	Vyr���M[��4Rt�q���z� A8� �|}b�'\��'�剢'ґ�H|
BB#d� pA�2!��C�!B�s�'>�'���Iof�<I#O�~��KO�z��7-�O���<�a��7Gm�O�2�Ovܔ��цg�![%��=�,Q���9�d�O��Ƅr����K�(٦�\�K. ���R�V8��m�SyR��WZ�6��O����O��ITZ}Zw���:�&˂E�2��!k�u��@ڴ�?Q�R�h�͓KB�s���}��C<j�F����S)�6���
Ӧ�aV\��M���?�����[�l�'#�����x�Zͳ�!.)��l�G�e����O��?y�I1p��y+B�H7j`h9��	i�r�!ܴ�?����?q���B��Iwy��'��՝*�.8�d�X�tt|i��ǣ>t�6�'���(x���)����?��*�Fm�Q�� ,��Sv�S���c�i0���7~2����$�OBʓ�?�10��xiFFQpӼey�b��;�Ɖl���Ky���'U�'�2R��#E��t�:p'ˊ8Pi8B흩�	S�O�˓�?�.O��d�O���A�d��|C$�8bU4�Z�m *8�8OF�d�O�d�O�D�<�գ[�>�� 
$*sb��s����c˫M�.�pS�im�	ܟ �'lb�'q"��*�y��ěs&8�PTm6	��Y����,��7��O����O�d�<�"�K�p����֘)B?����[�S0�����.��7��O^��?A���?�se��<�-Or�P�D\�xI�X0e�H�C�d���9�	ş�'I�Q"h�~z���?	�'<�>,��c�CX�Cpx��[���Iߟ��I-���	ȟ��	՟���A��b@h�uc�(@EJ"
ynZ^y�n��Rm6M�O��D�O��C}Zw������N��(i�R�h�Pܴ�?������?��?I���(ܭr�z!�^
tI�p�@�?ٔ���0g��
A����cH O1D��0�0D���r)?79�!@��)\��,Q���/�j��Sb�@d̢�,�^�)R�+5#�����'@ښ�!��%�:�V B�9��Z��#�@|
@@;b
�x#H�o��i����0|a��"G�-�Lp����-�0�J�B1v9Z@ �	�U����I.%ư0�2DT2_��e�D&�ܟ��ϟd�I��u'�'��5��K�EU���q{��	1͘M+R���83���1��S^�X0jմ<�AG~R�A��]�p+ڀI�`�˖FЍN���� ��=?��-�G�[�[IG�ę9� #=I7�޵1-j�z"ӵR���3(T*�b���⟘G{R���BA�����]�)\	(!�M���6�&"W���z�1OI�'��! G ��O@�$���.�蕞x%^%����%}
���O~�JP��OX��m>Mh�Ϛ�3���s�Y��~��?��� v�A�w���p �p<)��+1^`0�(�sy��L�]}��z�M�	����
�H.�x�Q��?I����	��t�JY�I�x�BQ���k�1Ot����6�V�ؒBݪ'R��J�Ka�!�D�I�s`P�g@&h��+	;f����|�@�'ӈ�� ί>����iH�f�����!�b@��%#�]P�b�6�j�$�O��r�B�%a"ʥ�~���|�-�D!.�LI���D>����>'�Kv*I( ���|���ɖ0:,δH�Ο*��tI&YP�<V �	ܟF�T�'}������zQtq��&� L`P@�	�'�Z`W�1iD��rV���	�ґ��;ҍ٧z��Y�G��f� 8���A.�M���?����Xe�3�?���?a�Ӽ;4�]!sAq� (T/H�r����Tm�%+�MF�p��/�1y4˲cҋbS��:��ϯ>����'�t�BvB�g�ɣ|�R虵 �3Iy��y�o��E�D��|~� ߌ�?�}�Iϟ �ɐ����fG�!M�L@$�8."M%� ��I�}/�uԂE�@�hٰ�fq3 �~���'ɧ�i�<�f
� GH�'�Z�޴�&L�"�J��Q�[��?����?���|
���?	�O���eg�0M�r g��%t�1���cv�7�'Q���䣐�0 �b�%<,�Pf�	rJJ1���'HH1	�_+Z�\EY��؊ D��5����?����?���D�O��X҃o�Gj�IP�c�f�)4g%D�LkF +�"�Y`/W�JJ	�!.�5�M;���������a�q�� �>�{���\!��?y-b�!g�:p��k6'A�!�$�@lHC���!0��I��S�T�!�$����� ㊰i�H��U	!�8-��@qN�-`j�:�M]�^�!��2H�fH��m ���&L4?!��Y�:�3��.U�,z�"��mT!��և��D�U;
qP"t��M�!�d�a"�r 2=�4ѫD1�!�D3Z�ȇ�N����7D��%�!���&$C��9&�P�tNP�CD
NG!��RO���p*��Ts�pW�A�`4!��9f갥�a!�)w�N 	�!ʏ+(!�䎂Xh��hp��P�/3y!�D�SK^��uƞ*&�2s��	,x!��a�L�t�P�l��ゟ��!��é6���4S�4���ǝ�$�!�Ę�[�8�R�A�L�\�� �A��!򤎷`n*T�& �Yk2!R�aԁ|�!�F+|M�d��:w^ P����%�!�$�;�d[b#N#2L*��*9l�!��D�uBr�q�	�#ScD�L�!򄅠M����G�U�N��	��M�!�ZnFT� &�hQ��!R�!�� �M2�K�Pk��i�o�c�^��C"O�t���ޢ�f0�g[�V���I�"O��: MZ�
�q�C�Bu�IB�"OR�6����Z�R�F$,V��d"O�d!��*ME
�J�7eENX�""O�+�ڧ'�]�%	�):l���"O�����0$���(7�̿�t�"O�ّ��ܰ�Y�" �P��چ"O.��4���ѭ�'A�  ��v�<a�CV?U��ZS+�Z��6�g�<�d[$p�tA�
��G$���	c�<��C���@}����3��93$Mu�<)3f�S���"� 	$r���%[r�<b���(�
A�ƀ�b3b!�tnk�<Q���:,�M��慔;Ŏ�Y��i�<�Ɋ.��kq��|&c��Wz�<��	-s��s�ÊR���q�s�<y���}�vf�1#�^�jbH�c�<��d1B�x��$ޫVQ���'�i�<i%�ۑ �걨d�N'���c�MZK�<A1��2W��h�U)L<]�����K�Q�<A�ܑW%��f��F	0�FS��yR��+=M�A�W�_8�|�ħ��y�HY�v�H���اb�j5yt�ٍ�y��)"��yw-NR�NL�ҥ�y�ƞ'1	�I�9*���+�y�KʅH��̑�%'B�"��O��yM�{�Ptkt!ЩHN@�5@+�y�e\��Mڵ�F��3�'P�y
T; �p�� �ǳrW�q��2�y"H� 330u�D�S;d����E��y�A2FҺ	rK�%WRЌ�e���y"��#j��l��IKo�`bi���y�I�4a����Ɯ��-�&EӢ�y�6,� ��f�`d	ֆ_��y"R�q�@f���尕(�	�y�-�%��1J���s�`��ȓh�xe�N�g�j�ضk];rЅ���$��N��ղ#f͑x����R-�F�B%�䙓t��<�� ��h�E�1
�b���:��5�ȓU4L��bƝJg*��@Ɋ-�P���0���i���F�����M�9F�Їȓ{ ����I�j֐����V�`��nD,)#hF51((�2��ʁ"^Q��h�p<�c`ʲp���14jT�kZ���c��Qg�҃)�r}1�׼5��ȓ����Ҍ`|�D)�e0���ȓ\lX�s�m�Y�P�д���t��?a�㓬��?M��i�N���q,�2�Z�
�#D���So�J�n��S!ٻ@�$=)"��8�ư�ܴVr:;�O��g�'K�ܙ��$�t50䮛�Aɢ ��`Y ��V#fD��E��=�$��PD�6����I�KW�����'tJ�q���S���A;3}�=�M�<0��
�z�x�WUF � uB�Cv0�"禮|�BA�'�e!�%�6])D� #.Pj�<��J
̠ !��_�y��JSI\�h�"�(V�����m���B�t	p���'0����Owk�0X@�;���^ۨi��MΨ�xrg� <tQ�Tf"P\@��s��9�V `��	�.��A�	,Y���d`}�	J�p�z���|�$��g@uc 㐔g_N�9�B'�0<9�1|O4�t��t���(�E�)N��P�RgMGRhEC���4Ӓ � g�>��+0?��9O��'Q�[r��BO�MT��C���z5�<u��	E�_t���+A��r�������h֚9'0;Q���j�h�WA:(,��3�B��xb��9X��8�ذm�����	�T�����º���2��T�c��;P��xgٲiC(�ԧ�[Wř�'<9qIR�_a����U<YQɁw�? �<:�-�f�adf�;5�6��Ց)���Fe�/"�V��`!���6.�n115�:��$=��`��MԬ*�>�	B.��(�ax��b�T��W 9�Er������P@f�ԥ1jrk �hz"�x�ey���<9Ó.�t��F��}�x�t�Y�|���'�z���R9�MHщ��a�	�R��8O��T����p��s����G��#�"O��7�M�O�|�1B�ǳD�m2�G֛�Z����G;c��<J6��6��O�=H2��V}R��m\�ٹ��Q0;F�)���?�$���G�e����jA
��MA�>��I"CTi�����0XuY��_�d�DdG~r�)Ҹ"Pc�xx�u�	�Q���&�Y*7�ꍲ��bn��U�뛴`��\���T'p�aY1�uN��
���%|�a�U�В�.�0!DE�3�G���Dފmք~5bD�`�W�a4d��"Da�o���M�{Y2�)vЄ&�C�	�`̀�)�$�r#���E�/*~l��ؾr�2"3�i����Gɗ]��:Z}���+OBA�d��~:8�1U�6vs>�2
O��	��@�5��#%U>�B���(���T���<PV�z��Ó3�����Y�{ڦ$��v���I�;Z�,��6��9�:�AXFoP/���`*R<�'g!�43c��|z�1:0&؎eL8	w'-�	3���K�Ĝ�SL��c���xܧH[Ε:ġ�(>�,5A�	V�t���ȓi��);V)�M�����Q�>Fd��2���#¡�d,>��D4�g?qQeB�Dq�4H2��O٢	)��N�<)��0���k�W[�U�Q��<�e��0ax�I���<9�A)=c�߿�rXQaK�gX�䲦ʆ<�:i�a���Ip��Kq*@�-Q��y��ހ��%y@g]9EP��aR&�"O���J$�'���;��H��� �PhC�v�p��
����K8p�YrFn̶V%��ȓaF�Xc��U0 �$<���/O���ȓ'�L����;C"���
ѵ�(Q��!�Np#r�D�\Aޜ�6MV�=��ȓ~8�pa4�ʺ+�&X�E�ŉlhL��H��y�Z�(�D�Ӡ�P�Z��E�~����?e `����b��]�ȓ/��1�´M���b�%�
D���|�M���'��ݐQ�V[
�ʤlW%�fu����y`�8�y�%�,H���lÉE�(�6�م�y�
ϤI%^���h_�7a̪�"��(O�P�A
Φ͈�$dX��Ɠ[�98t%Q�J���"O��$fߟ'mp���nY�N컇nX(Dj��9R���O��
b+�(rN����'Q2'�>x��"O(H{tiN<1���%`��@lZdR��᭏,�0>Ѡf�%�,)�em�= �`��$�G�<� �f��x3� �5�ّ��@�<���̟N��8�%�zi�Ap)�B�<����:;Knh��A�4G|�P�$�B�<��a��3��H2e*J� �#4b�@�<�@� ~8���2l��UR`�o	W�<���
%�d�t�� ���NT�<Y���;9&�|+Ď% i� ����M�<�`I�j)�I2qH�*�Z�Q) H�<�t(��!Ą�,b��L��G�<�I[�n��Pr� u5^��VC�~�<��!� �j��t��I/����b�<	���).�8��$Yp�Bԛ���[�<�v.N)cT�u#X]�FT;���S�<q��%�p�*O4.U�IӁ��f�<�����FM�% �~�� C5([^�<���Y����d5:� ���S�<yҩ�3��q��ذ,�`bg�Z�<�ƃ&|��&IvF�`�O�V�<aƭ��.�&XXt��S�H}J��X�<y�-�9c4��!"��=TV.�8#J�<���]�d$Yq�OO�g��M���DC�<u�0%�֡���zR��I����<� N���I,��z�E��b �2�"O��4eHs��`��%C�	y�"OT���(��ɱ�/׈ā9k�"O� ˀ'x� ��͕*�˵"OhȈ&�͑ \��P��9"OXMz�NX5
���Y�� )�b�x�"O}�&�/C-�I@k�%�|y�4"OvZ���lH�́S�C@���+�"O6�x �E&Xl�0�4H�<��]k�"O&ESF���Ib��g	�qFh�{!"On�1�F�$�\�Ȑ�ú:=���v"OԤCH
�Jv�T#%�9q"O�T	��(��	��'O�i��iqf"OB�ԽL�N�:���"�"B"Ol�%,��Nd���jA%}��"O��]2��1�A:���#�σ�y"-�3�*�I�ɕ1/�(Đd���y�ġ��JW/�qB�M�cA?�y���"Fx-kF�X� ,�g�4�y"bZ�T��#e���C`l�J��ǒ�y��ϴC�nwA�6S����G�
�yrO��8.2�C.KL���v���y�,N6,t�y�2i5o����'��'�y���-�0Z,��g	�˓��y�k�a�Q�&�N�w&�UV��]�ȓe7,��SQE�;��'s��?�*�Q�/�& +&�Z`K�H���ȓL�x�q��Ăx�!�2N�<]�ȓ�����B�H�ł4�ٮ��L��D�I���XA:�r�2^8a��-�Z����6jj�Z�) ,x��\�ȓ/�u�b��CI��l��[7��2t�eJw��f�~I[� �1�n]��Z�4]؆�ʓl/�Bv$_�#ŀ4�ȓ���"P4�آ��̗E���ȓTz$�1�"�"v(�Z��:=&ĄȓI�����ڧe�}:T�T$��I��V- A�˔;hI����F��\Q�M�ȓL����Zu�\R�!Ĵ)�d��ȓ.����1f�'0�j�h�&_��2`�ȓ^b��0���,��jѬK����/ �(���H�
�b���)Ѭt�Їȓr��	D匳i�h�h��\�V�X��HT�0��
m�Af \|�E��'�(����[9(MX�h�$0�
�ȓ  ��¢��6�|���Z�T��Ɇ�=0�Xe0T�z�*��ŔwHNԆ�,��3)V���	�$�Z
%d��� �p������nivp�,�%¤��	�t�0�jN��9�tC۠��H��A�	1"�,�@L3@I�e�d�ȓ:��[РH8v� �֯��	����k񎭻á kb��!@�D�Td1�ȓL�R͘D��1
�i�`��W����M�~(�	��BD�
EoV�)*���2�&,�l\V���n��4��dq��� Ied8�7�G�-2X)��i�D�r�bX�F]���`ߜE���Bc�E������>%�C��3��`��!�6љ��2R��8 �X�p�؍��=�$,BEȆ�[1�4�'*^�9�ʥ�ȓ%+&<��Ş3Ԑ�H1'�*n8<̇ȓ4	@A�UA�%^*tA`�n�* b�|��n�.�I013��3�!$-�\��S�? ��Z��_-�Ұ��ΐ#R��ݣ�"Od�{�CT�/d��2���'r�8��"O~)i���>-mE���%W�!�""O��k��L��!ȧ'�`=��pq"O�`�%�G��"̲T��%{��!�"O�0�pM0�2Y� mz�p�%"Of%@a�A�r+�ÑnrF1#�"OԍW��-|�� (��&n|ꩣ�"Ov|R�V�?�5�ś6Fn��q�"Of (w�٤m��C��<iF�W"Oj��`�q�ѡ"�T �@"Of�+SoF j��T!���<%[�"O��
��0z	�k��+32	��"O���4M��d�	�4u��t"O��
7M̿��He�'�@�"O,ň dU��XU��q��%��"O�����*{It��)����B7"O��We҉!�||[�H\	f��p�"O��p�#ߛ:���I曇�Rex�"O�d� UǊ=�&��p�Q`"O� ҧ�n�$TZ�W,,�]��"OL}��琉!���`*F8ڢ$3�"O�́��أo�E�p	X�N*��Ct"O��P�,�|��'D�>�`!"Ol!j��T�I%(��M�X��P�"O�`�ǆ*���B�T�u�kF"Oƽ�R��\i�QX��Ai�}�P"O�a�Ꮭ�bF�kh��aM��s�"OvDaG���2��Я�++����
`�<9���/��|#�/N1M� I �F�<7%'R�Z"E2[�h�Gc
F�<�§LA ���e�`~(B�@�<��-M�@DT0R��F,mH	
�f�x�<��E�1B0�e��Ą�v ���Z�<��`�46�,��U��1����7�N@�<i�*G=iNv=���U-H� ���f�<��%Y;=��!u���~ ##f^�<Y�jԒ.�@(�R��]��u[���\�<�G�ƃIy��� �� ORm�Ҥ�X�<92a\�%����r㞞�M��B���yR�P:���gF�.����HH��y�I��]�ՋY6"�$�Q���y����nT!�B����8� �fG��y"lY�eJ��c�����eHA��y�]���m�z�D�s�� �y2��68WJ�gOӀt�t������y�'�e`��� �W�d�FAY� Ӟ�y��
4mǲH� �۠����y"@Ň_���Tkβ�LiZ�C!�ybB�-�E��b�n��,�=�y��	�F�ZP���	�il��z����y�C�ii�Dx�OZv|�����y��ݍ}�|ZR���Q�D�yb��	)��`R
J[Q�-SC���y-�*<V�+�-�OՖ���L��y�b�4]{$,Y;s��,�ĪQ(�y"
 *����0dz�\�%I���y��,��(��j�(@,����ܛ�yM�3����F̾C(�f���y��T�c<Pr6k��eJշ�y""��u@L Ȅ��#���҃l���y2�R�.#F�Y���,6p9#����yRe�2<P��-��:84X8nT��y�oc���0�ݱ*5&R`�	���p>�  ��Ơ�(����Fݵ�m�"O����ݶ>!`��c�K
~
<��T"O�ahP�_I�� +�
�Z%��"OBE�t'��U�ء�OM�
�<H3�"O��B�ٌw�,в���	10h��i)���Z�9q>��@�}c�ူBV! �!��nW"�Ԯ��4U���䡊��!��R�Y��mz�Z@T�]���a!�D�)ô�@�f�18I,d�с�+p!��+�إ��a9�Pp��7DT!�D;P�0�A�_�^t�`��5:!�$��~���ZU�܄��A�یY!���*�
��E	�9�tt�%��o|!��Śc>�I�4��h��S2�=a_!�dO%�daE�)����c�7[!����Xe��&C�vt�a�\�1�!�dW�<UD\����EYʸБLW�]o!��:>m0�a�*�aM�1EL �f!�H�G.�+Ѝ,X~�QFŒ�:_!�$�2�m!� �".��QJ7!�!��'J�h�c0����XB��RA�!��oTę����&Vhͪ�Ə4e�!�d��0!�w �^��˷��!� �������L�V�%hϽk�!�O�xA�ݛU�^t~رs7��*�!�d�R��q��S=my�c�(�5E!��Âkb���g9N
�� �g}!��E8��	�ib ���u�!�d�TH!����)Abĝ+"�Ă�!�d_�5Y(�Y���DxT�x�݀,w!��S�@#��x��܉f�iP�-92�!�$��_����@eN�%���S�!򤚈�8M�W�=5Yr�#�0�!�䕧z��-���I {10}�#B��!�d	*`�*�ڱ�ȑ��*��ۧ^m!�$��2v%2�V,�l�QP�C8V�!�O>I�t|I.\�h¶NƼ�!�d���]:��D��6.F�:0m�[�<aנ�3^ؑ��m��^sX8iB�O�<����,���������I�T��I�<ߡ5<�����4S�����E�<�t�Ǽ#8D3��U�d��8�L�}�<)�L��:��1/�z�|��WI�x�<��S7	6�K1-FV����v�<�#�6Ux�"���9���Yg��B�	2(�Y 0l��EL����* �g�LB�I��[r)�^��zV%�w%B��)I�x�kA"�s��W�<0B䉇8հ|0w��9y���s�ȬB8�B�� u��qЯ�(z/� �'� {�B�I�{���ʔc���Q�A|9�C�I9fҀdBV���b(���
RB�v\�d��L�-1�!��/�)$]&B�I3R*�j�n�-(����sD�,V"<iϓ:�P�+�N������^�C��i��g�㤉V�Qt�P��gZ� 2>��ȓpU@@o�9�(���ړl?6܇ȓma���	�M��IZ;Ygt��C���	UӾ�b�0�A��kXX�ȓZr�)��kN�oRp���e�/ �*e��	k�'���a���:|��]���k�d��"Ol�����H��0�ʵi��Xxr"Odݚ�a�g�)r5dR<P�d�"O4 )��X{v���E�|с2"O� �M֋�?0@�9��Ц=�|�jC"Oh-ٶ�B�aFa�ᅼP�����"OH�ɕB��y/���f!�szP\�"O
���N�S3N�9AϯA!1"Oxa�f�y�ܔIt ��O�=��"O�{��� H��A��:%vej"O�Q�r���
���9Gϑ.r����"O�1S�	�+��;��XK���J�"O�p��G�]z,)���l�R���"O���Z >�ب�D C;M;=��"OBQ�S�߃~e� <*���"Ot�*�%I0:V<)�QČ(l��t"O<�; ]*E�AQCc�b�d� �"O�����^�~|b�@����`�4"Ob����7��m�'�v��Y �"O.yE��S�8��w��K��9C'"O�@"��ַ�ң"�-Y��4 �"OF8��-G�x�0M�p���1�ʍ`�"ON�Y2�ӿ:7�LzFb�n�6L{�"OR%����&v�xDcLQ#tJ���"O0<J��8Z��=Y���@h����"O�ɋ���.~����*��#nڬ�"O�M:�Q&yt��"'��Q 8 �"O�kSk�z�Z2-VcZ��#"O��2.H5.t��E�8I���q"OD�D%�e�D�aR���b<K4"Ot�"�� Vh9k$䅡v�ٚQ"O��c�T"M�4hu�����l3"ODj��S�*�X1�⓾5���V"O8��D�B�h���`}�.���"O8h�F�Ʃ5��AM��5@({'"Ol��G/�0N�T���N�E �40w"O��Q��w.��酨
�٨�"O�q��mR;J�8����4o�Ls"O D��QE��i�kP�[�m��"O��#�!����)I�O0X�ش"O�6#^���ޚ<NEҤÍ�3!�ĕ�@^��)G#�,,�	����'���aD'B�����	?aZH��'/*�@�l�l3�h��ٱ2g<t��'*�a3�,P$?"T�Ud�?10����'� �K�`Pþ<�QK�t���J�'�Ta30g��^3:���a���i�'������8�-��L:1%@�I	�'�|�c���0~��S�&S.Y0���'*��M��y.��auG�0�A��'�\�ł{ӒĚ5L�=}�c�'�*�I��B�5H&�z�� 4O}��
�'����*�?h&Y�s�Z�@*X�!
�' ։zQ��{�\�zC�ɇ0-���	�'�ᒻ�!��Ĥ(�p,k���yRàf�(|�3��N�SO���y2&�2��5&D�?�K�.���yҢS5v�j�K`n:Rra6 A��y��2��آ#�F��u'̎�yၣ5B{wM�1Q�B�n�6�y"#�s)��r#�D)���TƋ��yrFM�	��M����eɊ�y��"��� �`����yւ	�y�o��a�ð�L8�Τ{D�Q��y���Iup�+�	��6��9�F 	��y�K��	r�y�`(�(r 9�f���y�g��Mm���)תl�"���.�y,Xm!d؀NR$r/������y
� J�8I��Z�xE������k�"O
m"FL$[�L�B�ΉO|�\�!"O�:PDP%��� Ͽ�
���"O�$�%B�A@UC$"y��4"Oգ��E�x�z�{���=Vb,8("Oxt�i��D��Q�k�:|Qv�*�"O��G�e
��Zk��!Jn�Rp"O@��'�\�vyr9����04���"O���QM�$4�Y�&U�1��"O ����Y%BB���� �.$�P�"O���"���
�]" ��y�Zݳ�"O�]+��*��`��W�i����s"O*�k��ۋB�X���甛W�� �"O����Çz^
���E�u�^��"O2� �A�ȒH���8��!��"O<��⋘�a!n,��m�)�l�C"O��ĭB�:��$��b��4i�"O�U�T[]�-�o�-�m��"O���R!K<[x��sg.Q	�<
�"O�$XR�3tvx� 7+�8F�"�0'"O��NgU�����1&�܍h�"O*T{ ✀F-@�d�64@�1�"Ov�k��X��0���8Kf���"O�bjEsBm�%K���p�U"O��V��^�6��%���O�<LZ"O�u C�˞oa��/�,-ovсw"O*)0d"!2~z�#��"Qe�@��"Ob�2��L��D
>Y���E"O^D�Wk_�Z`P�;R%WRVf�H�"O��3c�P㖁��D(|1���"O��0��@�V���bX	:��C&"OVI����u�����!�Aװ�d"O���b�?8��E���Tʹ<��"O�hJ5��5. e�7 E�U���d"O�Dr�K+���-P3i���ӱ"O>	�uĞ(5a�K��s�z%��"O��1\&9�,p9���=o���e"O�4��$.]��U��DP�{���+�"O
q��l��P�ԀK��$OV�M�<i�'צ=t� YF`�X����L�<Ab��30t���-\�+��kp��m�<����J�N� �h�3j�؈��Fh�<)�-�<E-BH����Ch�ɻ��a�<��)�#��u�IZ�3� K#�E�<1D�A�,���4�p��\����<�1�Ӻ9��C�N��h�^��R�x�<Q���r̶Ɋc��vB����Lu�<1�I�u��"ʔ�� �Ik�<�2M�m>�l����,�XgO�<�p'�F�� P�3��Ñ,�K�<�'L�JZ��p�NS�!}B��1GIl�<Y��Y�L}>��a��",�j��!+V�<��_�>&�0�
�%S��kF�[~�<�2���*r�b���mh����I f�<w`�(o��9Rp��'� %��Lv�<I�cȶC��
�&M ���b�ğZ�<��h�92Nu�ፉ6<9�s��V�<q�ǈ�^�!'#D*?����3 �S�<y�b.s\f��`�ӻ#���Hd��L�<Y&H�E��s��9����FJ�<�3d�
%��I.�_���$ I�<��nW���a��T�EB�ı� G�<����0��	��@(c�Kn�}�<��M��Ar�Y�2mM�
|b0:��q�<� �<�1�E�20(p'�@�G[¬��"O����b^n��s��=K��3�"O���aK Q�v�J�b�i%f]�U"O��0���5 �F���Sw�pX�"O@+��Ќ?�$�0���ke��v"O���qm\�C�����/�[a��C�"O�d��Kηf<�bvn�;u<kt"O ����#ea�m	���b��8�S"OȄ��MZ,&X [a�U��A�"O ��� M�s`���	�?�ڍ��"O����
ё;��
�+׋�Z�bC"O��C����B��[�5��ڥ"O���񆘺a$��'�ǘ4�`%�"OЭR�M;�
�ң ��I���"OF@���J3�$�I���(s"O��c��RG ~��R胢� �v"O�X���<u����7��ʜ�� "O���Gە����GVS�H�+%"OB�x׏�5i���D�Q�@��E�$"OL,9�m0$5�a��]rG�)D��S��B1M���F�D)��.%D��H0bX$`i��c�T
��E->D����d��~���F:p��P)�7D����#�/��9��$ܣ��8#�8D���C��k|��	Y�,�X,1 8D���d&U9:�н�Ə��YD$pe�2D��@�(��/����(W�3x6X(&�=D�$k"�@�����)Ѽ�j�K�B<D��k��"fO�<�r�B�Vq�y��E:D�(�ŀ�6,����R��,R���2D�X�F* 9c���E�^�R�h1D� ��ʽ!X�%_�V_�=��)-D�К�h�:%ΚP�ٯ��Rb,D��s�!I�a:<ͳS�X	R� ��'D�X��BXX&�HC�W����� D� *�d�.�NY1�� �����-0D� А�7]��@	�n�I��m-D�H1��Τ{5�e��l��A�x}�q�,D�XJr �?b~Fx�� �-��-؀/8D�x/=+��#u�سv�
`5l�)|�!�ۛm���\�Y���:�^�2�!�$��}^,*l
)�Q�dX��!�"�D���+$�*�LV�W�!��%+,h-��N�+|"���� �!�d�%l=̱�F���d�!��&�!�$�-6���#���#H�h�F�e!�$B2K>@G�Y�d<Y���?�!���qx�TH�+ģ������I7݄��&�ї��Ⰵ�Ҡ�(]���b!��ZS�R,x�8���D�x4T���v��qs��5}P������ȓ�N1{
܂E�xyILu���ȓE��[�� "5�� 无���6%J�f-X�%�h| !,\���y�̱��J�Ml����&E3�x��W��=i��S�5NTh�"P�g�4�ȓ
jq�wFBku�E� %�*h�ȓ$�8�*$͞�wtΡ�R+�'��X��r�a*t�ʈry\ݨ%�T3����B�(sE[�[u\Y�.N���ȓr%��3OĄ>�ٸf�Ũ-�|�ȓ"z��a�5/Q�r&�*yT�@����<�#e��N�PN���(�EI ~�<�AX�?�MP��ͷ�`�Z�@Lx�<�  	��^�dr�x�/يL́�@"O4�C�!G�����@�
��"O)!�JtB:�y.2ޒ�D"O��"�
6XXd,`@.��$� �z"O��"�<h�dQ�퉶���w"O���8l�bI6�\!R�"Ĳw"O�"�mX!]ָYp�V:� �Hd"O�a� Ȼ3�ldnڻ�8�+r�9D���4-iBTZ4�S*̕��8D�Ӷ��q�H[pB1�� �5D��C$�·(����D�DԌ|J��?D���ˈh�4s5A5L�N�{��"D�Hi���vmN�2�G*"D�!�K�%w��z�"M:)Z����3D��K3+WU;h��A �UB��p$3D��cR��3(�LY��M�',���C%`0D��qo�/b0���.����j8D��Ќ��]�*���)ǫ4Z}�3c8D��7��5k^0�����(mJ�{s�5D�Li� �+`~^:E��K~�PT�4D�����/: �"e��H���y2�	�1@9  �:A��aW����y�	R6hW�!����i�hq�����y�H�jP�P�.��d�25"#ݴ�yҩA� ��a[�)�Z �$�%5�y��B:w�ƙ�`l �]� � 4F��y2`�W��M�Hζ'�.�	S���y�'��-���*6�%jZ�C�gT��y������!U�X$�NŹ�O��y�Q'i���q������y+ �y�C+`+��z�B9ιk@�J-�y�!h�f���Im��O��y���!�u�6�_�)�
���y"��v���'��/Ң�Rڻ�y�O�J,��ID�|��8�K�.�yBm�5�H���������9�ybO3,ܞ��"�V�ݲ������yB�֎G��s4�7}cNa���4�y��8-�\�1�N�q�j�sN7�y�΁/Uܴ�P�G��U�`z���y/֊2 ��DA
K+≻n�!�y���i���M�m�]@k���y�`C6-��ܯr_8<I���yү
({�lH�E2p[8�����yRE��o�V�R�g=v�D�d"ڝ�y�ś�v`��v!�*�t}DZ��yd�-y/����33����
��y«�;J̮,�t��+�޽ �A� �y��&�,rg��m��`ccCɸ�yr��,>�ƨáN�Y��[�L���y���,
OB|AGC�P��a`�
���y�)�=1NM�e�Ñ3�H�B��_��yr�Z}����f��&����A@���Pyb�X �Vd�w�r[��G�<��hV�L=��R
 �V�H!g�J�<i��K�� � 
�uZ���I��O֮:T$�� �K0,*��݇�9v����C�&e���7��,,X�����#�ڼD\� X��lB�ԇ�S%�A�K�3"�-{�D��J����I[~ҭ܋{R�'��2^��P[s���yb�~#0�̸j@Y�'���y�#B6����E��4�qAB
ѿ�y�@
/��k���pA;�I�!�y
� D�p$�=+D�ʀD_�O:M҆"Ob�Xdf�;"���'Ɣ_R|�"Oj�Цh���p�A�Z����D"O���SE�z�:aF��(
��d�IZ�O{l�X�
��N� ؚv]�v���'��@��o�.5�B5��N�Z`�<��'4����*EX0�v��Yf(Ⱥ�'2�ċC\ߚ��TC��S����'��p*Dvl�<�Ƒ�9�����'`���JI�dB�.F]i�H�'���2/D.��9P�F3�h�p�'���s�.��L��"E턽E��(	�'\�$�ɕ��ܲSI��<��)��'�� X�-��y�Q��ٝ<��u�
�'�l��*ښn��D;��?-����'EX�`ٻ+wvɻ��ѭ,= ���'Lҥ�#�/Fo����G'*����° -z��EBU6. J��d�c�!�D��	�i�@ӠY��eJ���7�!�däP�쬚��Df��Aےd�'�!�סJ.(t �ԏ���YT�\5�!��ɫQ"�u▉<n���䀔x!��U�f��l���6}�liפ�r!�&4����*�8T��{��bp�}��'{�\�$���.��^;������2i�!�ğ�\:<�hn��3��bS�X�J�!���3T����$�~0:|:��\�!�Č$)[�mJÛ�t����
Pl!���_jB�nÂ.r`�Bd���|6!��Fy���HTm��pL*�PF.��8!�ď:3�����D	��iR ��?�!��(��ᘰ�?/͌0c�.r�!�Ą�P,��U���A�
�!�d	pi���u���0�����@,�!�dӔ<�h��&�	�zt
���!�DY�>�yCT�";�*�۷jJ �!�	q�`�qƣQf��R��Y7!���9O�:���d}}n���(��!��[���ȀnZ
e�s0*�2!�(L�t�/��>L�q����!q�!���p�M�P�ǽDe:�"K�Y�!�
R^D�T+P�H]�� P�!�$��I?��Y�L�,),P�Fږ9�!��W�Ҥ�'�)t�<`����HG!򤂛H��9Ӄ��xbdD[��;B!��Пp��8wl���ɦ���9O�*WIC�6d����k��a`"O:X�� ��C��� c�?⸙��"O��T��8��g��d�F�/�y"���	�`4�a:�N�ԋ�/�yR�T`��h'��!7h �
��y2ϓ�Βxb�P�^`��m��y���	��ģ��=\J��1�A���y"DS���=����CHDC�	��y�F��C"�ZAf�??S�-� /�
�yo2`_��¥AI�v�� oҟ�y"�վ=�:�x2���>v�ZcnM6�y�k��@�ly`�# :����2A���y�ܝ1���P*N�/��S��*�y�L�
�(����'ҮeJ"� D�$���̦oJ� "Ç�Dm���uC<D�Ȅ)M�X�j�E���}�Ȓ�4D����A��e
�C!e��qBy��/D����`F?`�H ���!���$l!D�� X�CR��C�pX�1O���lhR"OfQ �N��80�MS�;��,�F"O(x�!�!X�ᙑ�^�<�V�9b"O�H���Z(~���,�]4�P"OL��VL�SԚ�:Dk�xްP�"O*��#V5_���au逤/j�2�"OrP��"�'��@��5v�j�"OZer�ëB�d�9�lĘE��(��"O��	C�M*N�Fd�kT�
��"O©�E�J��9��L�r7�D8LO�e9S.��^L��"o2rJ�%��"O�svi���j��v���:4T:�"O��	D�����Ù�G0Ҹ�"O�� �D�E�|�bA�jث�"O~��r%�:j#l�4��?>!Ne�Q"O�ث��_*N�bl�����"OPy�� ���*v��i%
iY@"O�[ �*��c�>+��I�"O�ux��ɐ*�8��f��A�6Iq�"O���)B8���r���Тq"O���E��`��9�pG�"��	�"O I�q/��O&�11����\bD�t"O2@k�Jվ4���Z'�<{M���"OZI�p'_�ywLy���L�:Q�HS��|r�'-�9�%���k�,`�EAߖ��Q[�'dZ�'��<>#�i �((�.=Q�'�JÒg��0����- �h;U($�|��'�ND����"G��^�H��'i(�)�8y�}�&g]+ ��hr�'Mv�r#OF�l�qG��Di$��'��t��I�
�90���C&����'�D
t���лc���7��]:�'@�U��,���1�I�)4�t��'���Jbl��<熡�d�4_Y�ExK>1�8X��coÏS��	�"�A�|u�ȓYk8e�0�����ȋ�C�5�ȓ4� �q�斬\��
�D�P��ȓF�|���-ÞV���2QOS�
���%��3�eԜ���@�+] ��ȓ(��eB/-�L�"@Ƞ �f݅ȓu"���K�>20rP��q�|���V)�4��-��$����-|� ��ȓ=]:��iT=R�*A���&d�V��ȓ+)�)��٤?�$���a *�����c�@�Z���2|h͂%卞J��1�	����bu��뗵H�H'.Ѩ �t�k�'.D���VŖ��'�= p�IA�&D���'��8ޢt�&��!)810m%D�̉��ĬqF��'n��z�%D��3��P:���S�F�
 �)��("D���
�	_�� ��$0ش(��>D���1$�<%N��B�8Yt8
�n<D��6�@�#��|8��j
dD�W�;D�����L<5����4'����4D��sb��|�� q�b�tc��6��?)���O֢�!� ����� ��PB�'��		�!��Q'�y�p�@�x!Y�'��ⵡJ�":��b�˰P@��P�'�X��J!����I�T,1�'�	0!$��\�ve��EG�>|v�p�'->Q����ep4�����BfT���'��yJ��o�j��oF�6�����d5�B��xCc��~�ĉ��N8�(��ȓh�� f��8i��QIW�B6E$���S�? z��adۛo��@�#�&��y"O�xGE�6:��Є��\���9LO&�����USBd��ճS����1"O�R���%�����=\���"O�䑁/��'����-	��Z�A�����o�')�H��D�۵qI�l�D��0E��ńȓ4��!PC��
	��#����X�m��er��'Z�}��p�p/S�B,��lz�x�#W�M)�b'��$P*�܇�O`���eL�30�CƩ�!CF�Ї�ybU0���$:���#bI l�}��@�4��T2�`Sc��C�ҭ$�F{��*�Р�pu_+^q��*��yr��>O�qPa�ٞRy\�`U�X
�yə	�:���
]�AV����E��y2��Zx
��p�(p=�(Q���y���F�ё�;MT���b	��y�$Э!=�������3�2�*j��y�lH�fH�R���=��5���y҉�.�0(jQF�2�vݪ@����y�Ɂ��D�3�^7.*�� ���y��PaEX4�� %�6l�b�܉�yB�� :r�S2�2�8!C�H��ybFX���B�c��flD�-�y2��8Du*a�F�ij���w��y�D_ND$8��I�S�j�kֈ@��y"�׵[�Eq���I~�-��̤�yl�%<�̄kB,�B��0(����'���t(N�����i�:#O���ȓ'�����Kfp04�@H̝A�0�E{��OcJ��$�6��0���F����	�'dB�3�O�/@�h�$��<����'�8��F�5Y�������~��a�'׶]S�@݇�nYa�ٯ�,���'3�@�3���lw(��F* 0Z��'Hi�޴G�U���$`>�8�'��ABBl��g4���r��g�� p
�'��pӮ�"m%�ib��d�J$��'�t�%OŊ�T!b�G.K�H���'\ ѩ�a�{�x-��Kβ=��ي�D3�[����˝>��2�(5�h���'�����N�L�=�t���p��ȓ�lUs�d��U��`����+i��ȓh,�����L!�X�`)��.��ȓBΝjg��D�l��e )�x��@��Bv�نs�U�D�D� �2m��<m����γ]�<����z &U��o�P�k�`������i_v �H��6�L���� v�S��ٙa+�0��1[а0�FS�]�c�oH�5��ԅȓV�
ؒ��ҥ1��9��ە-���	`�'���R#(�^zzuB�߹�x]B
�'�]�H���ZٙÑ�A�u�	�'�L�i�n@!T�&ea����Ի	�'3N];PE�P���QLB����	�'��
� (3�<Q豪V5{��l+	�'�x�H3لI^�A�ԇxNN���'Ѣ1�g+��{�мc�wH^<�	�'6���aT
H�a�(�{�&1I
�'8 %B��R�L82���q���	�'�|�+񢕂C�ay��_9V�y�	�'��A�*Y2g���C��O)S	�'(B��D� kdP��-�+�pR	�'~D�"�C��W1� P
0Ǯ�B	��� 4̓�G� ��!I���#%\�PE{��+'͢%�wH�� �"��t��z�!�T:N�"���#a늕1gʍ�3�!�Dطm��9p3éQn�	�v���\!�S{^@�fK\+0�i�c�\;9
!��Y�H�C�d��htC�6!���k�̀)t��4�h�c�D!��&qpvtjQ��N��#3��
9.�r2O���p�T�a���R����,u	`"O���7�גK�	�I���W"O�h���$Q��Qe�,�v�	�'�R5O�"�$C.��}�wƑA�0�s�"O=cC/�&i����OE�n���"OH��e^}�z|[�m�!�\9�5"O���2h�1Μ��%��Hƨ�Qc�'���|�X �Y�Z �;���{2!��
S����#�/>|х�V�!�d}2�$�2LM�  � �G倦y}џpD����2E� A� +Y�Lr#���yR@�4r�T�sf�8%�0�!DcV��y*PHmz��2(I+MPU3遡�ybgո_\<\2�
�f��1��O��yrˡrјr-S�	�Fi�Jʹ���hOq��y��	�/ḁ���F�j1n8{�"O 2��	"��P�fτ�F���'��8WE.�I���|�(�CkR�k�!�$��3� �↸^|l�F�Oe�!���2BΑʰ�V�j���	�^!�$��T4�W�Y�����hX�R!��(;R(�!Fz�.�Y���=!�d�&~����Ryм�z&]�!�
�z�0yhfȎ-�Q�9�!�L>J��a� ��NР�G��+,�!��X����Ŭ�.I:��4�!��8�4ݱ2E��OՌ S�$+x!�ݫfx��nOI�Δ�q)�	cr!򄆖T��Hʷυw0��rThFW!�DJJ%�$��Ïh&�R���TX!�L��I�`*$�p�"��Pyb�D�y���g+�,?x�]@�aD��y�ӷ'X`F��ڔ�`Ϥ�y⍖b��р�mQx�B�����y"�5�V��,�`��0�-
>��'�O�c�2��I�5�L ���f"�(77D�ʒ��hr��8$�H1�S�44��p�HG'z�R���W���Ԁ�p�<�0�/5aRC
O�D<����l�<�%�OH�����J[m�HY�I�N�<����1
ʘ`Y�Ɂ#��!���H�<���յw�z�i�R&8԰Xq#AI����<y�j<fH���ԐE��ŜY�<)U �t"�!���(N���HLX�<y��^4����@dHS���_�<1DD�^� 43�
�}ـ1K�ȟZ�<����C�2	6�0a�0[��+D�,���$J��R��[�4�Z�.D���Da�j>�3�M�7?�N�K� D��Z�H��8@���eԆ-<B"<D�TR��y��%�3)�$��Q�c9|O�b��&ȿ5��)Jb�ſ�x�+5��V�'U�ɥ�� ��j�cЀ�+�����DC�I���:7��"\a����!*\>C��2i��@�� RL��5�P�\��C�	z#��ҳ�_�[:Y��J���C�)� �r��G�Tu�VH{G��"O�p�v	G�v6,I�����q�θ�C"O�\��M+�: �
�~��sb�|��'��G{�\�Ҍ��f*�$i���6F�!��^9u�|�a�39�T� EM!��ݭ)��X�,O��<!#w䛈H^!�䂚p� ��e�]�x��UxF��!�$�Uf�d����'�ra #h��2O)��O�$�}hR(ӿ/H��!B"O�)�G�
|&�H
��
-�,�"O��v,��6hȔ�LG���k�"OB�R,�.�.a���8��}�s"On���G�"	u�5����3B@��t"O"�v��@�,US�f�q.�TKB"O�U�nݲ`q�q���� �"O~h�ħpfZ���. )��"O��$�W�j�Fui�Mǂ�f}��"O~@��
2Ak��Y3��"��Y�u"O�<�� &�2���̢y�H�"O"�h#�4�01�Aݛfmn���"Oj�C2#�8l�f�c�
T�g����IX>�cd���`�LX��A	���$D�`P�@&Nhji�iH�q,��rV!�D�O���>)�q�J3��ɵ�K51��? !�ĜP��X�o�Z�P���	Z$s�!�$��E1Z�
��'Ѳ�3�h�:5�!�(Cn��bB�� �L�%h̕9�!��ʖ&A�G�I�%� aȲ�Y��!��6d=�˔�>dG�ЉG��72ў��ቕYZ\b���p�`�����	"��=!
�',��Y�N�,(f/��p���}m
��!ϊ`���Dn��K����ȓ� U�w$�Ty��+�[�R��]��;2zX�K]���O!s���ȓE��A��X{�≺V�9O�Ňȓk߫�4{n�j!@��z��x�a�IC�s0Ă�A��0�o��S�Z����<Q�
g�����C�Phk@�;ݬm����<���)����b'U�DF���dC�I/ؒT�%�.&L`5��/A!bC�ɑ�؀��G�9+u2��/whB�ɋ�Ҡ@�z�\��f�P�7FB䉚t���w���V2��c�'v~B�4���cA�My� �C��|K��=��K]u3$T�6��&��|U�ȓk�V����(W.uA!(�(+$y�ȓ���Y'�;خq����OM셄ȓ�\�Q�-��p����$]�䕅ȓ<޴��N2L0����!1�<���*S��C�m�y�D!Yn��
�'�p�Zf���2�LD��Ė"mܚ	�'�	�1%8h���R�Z�hD���'pVl�FA�:r�d�q��J]��c�'�t}8s�½]���Iڀ0%��'��-G�\	��
<׎�'uN�2F��2M�a`r��"/�Db��:�'O�*�@��x��`�ͅ(0@8ͅ�?`�/�*p�2)+P�6���1Xv�����6I�L9*!�-QJ9�ȓ��̂�F���s��a>}��"O�x��G%舕����aL(��T"O  ���
�P�a��� eT��"O"0B�� ��m�o��Z�"O��p@�M�l�$@���M�Q{U"O� ��Q)��gL��pG�lE�`"O�<�"*F!1�]s�lH0QE�Y02�'�1O�li׮�<a�����˃�o*��ʰ"Oh9�eD�,F%ޑ��͘�(�=1"O�)��&��W^�a{��S*�s�"O��3� ��$E��ɒkΝN$����	G�Ob ��6H���TV0 �6�;
�'Nh��i�DTPɰ⨊3"��Y�	ϓ�O�4IF�C�"��i3��ר=�^-���|�'#``	�3Q�@|��.����'3$H��Ș�D�Ҥj� ��!�'��<�q��_(L�2�]Ya��'B�;���"13�D����%�N� 	�'��S1�K �^�� �="'�9x��!�$*j��n�!8��\|xt�#D{�ID�'=1Od|��i�2�~�I�oW8-J\EpT�FB��#�`��]2�B�!ƌ??$!�d���� ��j���D%�y!�dB�or��Q	�vL0[u��3!�dn�����&<o��a��ܵF!�$�E��y)�Y~mP��D��l�!��թg<��D��'^ UICn��N�!�$>O4�A�sOє�Ľ*�mT�8͡� 1E���$-���m	����y�����Hy�_u����`\�y�o�-$J�����ɵ�\��y2�5k"��4b��|#�U��F�.��>��O�aPm��&�����
�~�lY�"O��z��=[��=����h��b"OlLI�݅v���q#։OkN��"O�x����2@HT�5bU����"Od!͋�I>�Y"F�6���P�"O�E���rh�p��#T�2 Z�"OX(�炣==E��@B�yt��Ye"ODt:WO�y=�� �!	�@Xԉi@"O��Q7)����aΐ�d)�"O6t�t#φH6�p�՛6��X1�"O�p�ς�K�޽��D�a� l�3"Oj��1�I�iWZ�r!AI=`˺DaD"OI+�D,$��o�b�^=2�"Of욧o�)-��"�S,'�����"O`�Å�M%;
�}�wd�" �d�`"O\��f��pD�K��J�F���'�ў"~2�`_0yڜ��d*r(́� ���'�azrf��%�8��B�Ĕ~+���u�O��yRo��tx��3��o40��ӇO�y�'�8~��D-ŵd�.�j��j�	�'�X�Ȗ&JOE�aр�D82%jM>!���?��7v$��7���9�a�)oXI�ȓXY�Ԑ��x,j�Y�
R��F��_搅S'�Rz���pI��)�C䉆)���A�aܹCw-��$�B䉖s[��0�Z:O#�5(��	n0`C�I�U�
�3�Ԁ;�8�b�l�0��B�I�}��A��ȕ�JS4��odh��'e���H�D��z��P��N@�)OR����=���h�˗e���6bA�}��� q�	�@!qA@��]~nhI��6D����j�'G pHQJ�$7Zx�k/D��h�CI�O>��x4�H(��j�-D���뒌Yy��#�C3X5Н��J+D�d��k�(�R$� : �T����(D��9�Z3T�P�c!J�3�8I�"D�`�Ђ�Z�|�F�^�F��s�� D�� ,ѩddÄF3lQ*ao�y���d"O	�)Z6�9�v-SV��1�"O١�GjՒ�.8'����"O�<�3J	�$q�dB�G��p5J�"O��3%�Y�?���b�6�A�"O,���� >g���`��*y�Xkw"Oj���K��.�<�㄀�/U�`bb"OH��EN�f�L͙C�/-���"O�}��m�IK�+{��:����yr��.3!����X�x�}Q�+7�y��@�UԐ![b��� ��������y҂>Ċ<I��xi��K�%D��y".Ϯx�mcT�k���C$�р�yҀ׳O�<A��#p���o<��=��y �k�ɡ֢N(��-1�����?�S�Oa2�C�^�<��Q�G`ʃ�f�
�'X�葂K�
Xl�RתQ%�@
�'�@ $?�j�Ag!��v�ހH	�'�Fd�1�
p�9�6�o�J`
�'n��0Nۣk8�xx���s��܇ʓp�����I���"�؅���CC�'�ў�G{��3FE�@)WÇ�.A`�%��|�ў��'p�|���\�u�,�Y�íaA��3��6D����䛙9�0dS�KB�qfb���4D��r��˜���!f��v�p	�E2D�`H/ɤV����j!Jv��!$D��I&�ŨR�\�6�n~���n"D��C���H��	"���4#�Tq��/"��8�Sܧ��Iª��x�S��%U*^X��]�92�ʊ�"��S�@�}DX�ȓ�Z�9��2)I$0�`��L}�l�ȓ�N���ަ"�M	��֣9HƬ�ȓ��eǀ�@`	�"��9I�z��ȓ4���!#��H��� 'd�UP�-��u�'B��éߨvۊ�6��ZؒO�=�}J��6ux�y6����<�d��Z�<�P�.�&dȩ*�����Rn�<�r�϶A�X��գ<!0�ı��Ej�<YDo� ��14�V:�X�!ŀ~�<y��<;�5��15ܴ�zrMz�<��jI>�&Ah�Uhv�ʡ�MA�<�A�ՙ(�MKB�ͻ�#�w��0=���E3Z����
�@�A���p�<i�(�+I�!��F�	:�ĬQ�<�4��� m^8o~�ȑ�w�<�`HĹ|f|,��F��U��a$��I�<�r�0P�OD;�H�B�G�W�J�ȓ@�^��B=�V\�bE�gY�`��F�Y� �]U���`1��-8�P	/O.��?��'�rV΂?;F Pd�-L�Շ��m�'x̀هK�.+"*�j���TM��'i�!��b�~@�*��x�����'�>�I`��Ft�!'�Z! �b5��'���w�1#�~qŢU�wِ���'�=��	�8Q[Ĩ�$G>j���)�'W*�Z3��5OR��0�A�<<U�	�'�l8#Re
9�B� ��v�����D�O�"|�O�	�n11Bj	6�
@�q�<�u��7��m�Dڳ���� ��p�<Q�͖jт��*Y\rTbIj�<�҅ۃr�����@�*i"�m"�BNe�<�`��G�.=���B�.�Ѵ��a�<���C���4��6x��)�%蟨���Ywv��" !P�n!c�'�-�X%��S�? t�IȂ�2Z��V��<��q"O�u0��t8q���;XR��#"O�!���b�~1y��[����b"O<�3�oP]�<���+�̑$"O���R��u2Y1㊅@���C"O��U	F�~0�(p/�/�����"O��JX����3*�!f<��A"@��y�E�<e�D�?�-k�f�C��(M������ڷx>��)�ds�C�I�G�`�M��@S&9����7��C��]��Gh���d��R�� P�C䉀O"�9X��A�1:�3ER4ɜC�I=:�<i�Z�<H���A�6|.�B��O�p�5�Ƨ<mh��U?�B�	>h@��j�,�cP���@З�B�ɏEP�!��T�O�0c�g͇G��B�ɳi���A&���Q%T���	=[�dB�	�g�P�a��?�&��Q�4k�\B�	�:��䲖��Y�|���lA^B���0�@0Q�	��5��b��C�9_�4�@��Z�|���E����C�	�K��Ś�LN�1�p��	��C�	lL�R��N�+gDwF�1I�C�&hUx�;$O�[���gd���\C��G��f�Q�X�#7f�(V�<C�I>q*
�Rv��xQ4`K��S=	8C�ɂ&C�y�C�e��v�8'��B�I�h��x{
�n&�%
Q��B�ɷZ܌8�O�������^(C�I�P�<Aj0f�+%0e�+��B�I)U���X�c��0 ��Q�fU�C�ɱc[*q�WM)p�Xyr�̒M/dC�ɥ)x`i���$	Q��	G1�PC䉨)XT$�G�E�07<ە�P�C�I�k,`��N\�{ ��Rą�P��C�ɰ)�f)8�"��y]���%�^$0�C�ɚ6`j����$Tw�Q臣Жr�C�1&�8]�S파r4�[��P�sB�	g�Nq` "��+��#	���B�	8o.l}C*FZH���4�-�DB�#x:Ԩ���]	Z.nT���I��C�I�}��r��=��(C/@<$�B䉷K�\9SM,�d�X3�.l�C�	9O���:�h���dؠ��t0lC�ɼ2�b��gh��k��{b�B�a�jC�	>1EY����|r1�g�8�4C�I�R�H�����\90t'�u�C�I�S��ZTe�?2Hl�p'ȥp�B�	�'Z0���*ܔ�(w�G�Y�B䉧2h�4�@�O-^t0�4�"R��B�� 9r"�����Q�ت�hޠo��B䉲9/���ҍ�),��="DAݵh-|B�ɉS�� �]K�2�s&�۶A�~B�I� Ş|ˆ#�1=��r����+&B�ɵ@&�4(@�O�
��ܘW�xc\����D8���\�\���&6���3:!���=H�̺�T%l]T��lXu��ǔ�2�X�j�A�A�a���X�k�荒5$�3@�G��M�ȓ{hiۑ�P�mE�(h'̌5q> ��ȓw}��y��,�]�/~<����:E��N��w2�����o�H��ȓ!/L�[�̓E1�)C��!�݄���d
�O?:@r(sGn'Y��d��S�? Z �6 R����1Gˉ�0���I"O^�����gȊU�%�ۤ �Ա"OR���}4B5@�D����B"O�]�H؏a��䅼Z}��"O.iʤ'F"_���� (�3w<|{�"O�@8d!W�N��ɑ<\l81"O0m��� B�(MōZ�q����"O|�"s� r�(������"OR1(�"�+z|�e�F�z�:�+6"O`fkʟM���c`$�:d]��"O�����O0�����	H"Ox�*�
б5Uq��>pQ�1"OX�i�
W
��j#g�54"O���ǧz!��!Щeݐ�"O���LՕsQ�Q��(��PQ"OF��
V3q}�9	㢈&|���"O��ʅ�?�M(ӡI3s�&Tp�"O2|��N	�� ȵj3HJ��B"Oj�S`�!rVE{�LZ8+�9(�"O��@��Q�v��sU�Y�^),��T"O��c�"׭y�����!5��d"O��q�	
d��I�%W1�E�"O^TtǞj�0$�B�şsŐ� "OHM2�K��'v�$dг�N4b"O�S�L�� ��I{E� a�"Op�᳄P���H@+.���"O�A��hR�Aw�ݙ(G�!�A �"O
�ek�9X��-KeFI�-q�ԑ�"ONK���L�4$��#ҡ
�r!s�"O)��+A��L�b�QraHd"Ob\��I]	*�4MR� �vU��%"Oq2�-Z�0�؋Ձ��=N���R"O�ED��8hA[3.�1'"O�)! ��+}(��Fo���xX�"Of��S@K�$"np��J< �`E��"O0�7�$YׂyCMѫ#���s�"O8@�7}���s��S�����"O�̋�@��:���ť�A�"O=�F��h<@8Qc �`̲�Z�"O|�2��K<8ed
P��)oP��b�"O^�sqB�f�t���}Np�s�"O���Cַl����!��+����0"O�D@��=�`��R�
� �D`�C"O\�J/�,�
U{�.�2��,hq"O�,k�hU���#���:�
T "O��3�R��r��ìQl���"O���1�I1m�䤈�oɰ)Y��"OH�9N�LK��0vF�LZ�0"O��5(xP�P�5��Gh
m��"O�����Y{�|7�ҳS�j9�"O���O�s��Y�,T�U�L�G"O�Q#〉v&��aC�T�|�<E�"O�����s��� �I4�Q�T"O4���bɜ.�����ΚON@9	w"O��g���H�!�p�?c2`� �"Ov��nPyL���N�:`�B$"O�Eh�yY��I3�&1���2"O�L�$ɑ +�X@�X�N�HV"O�I�#��F���q+ֹ����"O� �Jʾn��`�R��4i�4W�V�<��� {Rj=A&�D�,��S�I�<�$@�hIF�6ȍ�xfA��G�|�<A�.2 `+� �Lz���-@�<a��8F����I�22B�:%��}�<� ����H�
�bA� %�4ŤlC2"O���Cђ?v�]�E h\ زS"O.�����l��Ł�d�Q0$�)"O��8��}�,��Bޝt���P"O��#4nˏz=�Q�k62��%��"O\Dؗ�Z��1y �V��<Ó"Ox��JS� 0!��T@l��"O��!6�
s�ޤK#�?%H���&"OZA�'�\�}��� Q��YU"O ��Pd�J5>�R�/SA$MBr"O8���8x�|
�-C:Q-�(
%"O�%b*��G葪&�[�q@d �"O4���!Ay|%"�KEo^B9�"O ��ǧ��Bn���/kR��aA"O�	�2囇^�$�8-�=E�6y�P"OR��u�6�ֹ�g�G�J�^X��"OZ��𮏠P��,�9�����"O.�[qT�)f��: ��b�ny�"O�8۰��9�.]���Sg��ԛ6"Oބ:�C��c�l�H&�@�6�)�"O`�*R)$lV�B
��R��0 "OVA�m�,^>H���I��Q�2	*D"O�T��l�'α��-Y�:A�r"OJ��W$)@Q\�鱌�-�a"�"O
��r�8dt���G!�j�z��"O����a��;���{�%��+t�ur�"O2K�m���E��D�2f<|ae"Oh<���@%RU�T�vP�5"O|<8�,�4Q���r �Hjj��"O��i©8qU:��p�C09i^��"O�)v��A�D��D#]7y���"Or̺3���1,쬓�,fX����"ON��2!�5�"fǇ\P���"O廦g�3X�B��՛
7�*1"O@z��P�QM@�A@��F8d�!�DʏR4T�&,��B��I1G��!�DΖy�9�A;R̸�I5�!����	�B��/�P���ͳ�!�� �:��4��X6��@`ۮ!�!����P�2�U����t�]�n�!��$n�E�a(B� �U���!�{������*� �U�!�!�ٯ{|���-�Nl��[�eO��!�E�X,�8�m�GV4������!�T�!f��:cIt�F��?
!�C+	�8Ma2��1B2�#a�p!�ə7u4�3�h�'ya|1�R��69T!����,�c����hc�tF�'|�V�)�:]jdY���.�8�vo�C�,C�$B�H�BԣL5�Xg,+�<㟨��I�(��$zw U¤�CSB8:C�I�*Z�Y��$�̙  T�4C�	�R�pa@��ՙ20����	�;YV C�Iy���*����>,�w(�4C�.5({�iݪ.�����NB䉶��l��Ji�f���lEG�DB�	�+~���`�M�C��&�����>�4%Z"52�}С�@$�ʓ�U{�� �'��`�1@�g�|袠J�Z�Q�'θx���6�E#��:�1��'A��C��s5z5B���?��3�'�
���E�B��s�\�9��ջ�'�~E��'N�4�<��!Đd)|Ez�'ʸٳ&�Y�z�B�	�*5^�x�r��� �=�ʍ/.$H�ҡ�>K��U�"O,A�"[�(�6����#V�ށ1�"O!�W��-�%ɟw��"O~4�I�#��Y9��B�MC$@�"OD��Dع��̋ ��%[&�ӣ"O�,;!���I�R���Oٍ&�Y��"O����������q��j�q[6"O��r��D�+����ѭ�A�*���"O���㎊�<'r�)q�![����	.~�Q��VA@�ȁ� �i0�pi�EA,?��9��i5��P��I?g6liF��݇�jcHtr��	���[�ꑮx�����mj�[�G�ͮqc`�N)3^<��K9 1:�bV
m�9s���%J�� ��I{�$g]��X#' ^Ӽꆎ�8, ZC�	�SOXXƤ+���6�2^�b��D<�V��e���K�@#�\�`k˒a+@ ��Iu�'d�e+L�-	�Ŗ��1Z
�'K�512C*<� Q�DK:E�>��P��$�>E��'��! jJ�[{�q�0��5�,���'���y��ڇ\��X����6� ��dڡ�HO���r���b��w�K#�̡3����B�Ҷ��(Q�1p�[�a�ц��	���'��?��e?�z� �3~X� �	*LO����ͬ@vH���]�1;a�;��`��"<��y"� Ô� 	�g�̕b�i���yR�Q��=c$��I\�9玀!�y�kC>C���q��ˑGs2�+Y��0<َ�d*&�U#�$p��8��e!��	�9;��\WI���W�%h!�D'*t|���:2J05�&�R7{g!��,O̊�P¯�-YB��B�G�Y`��c�'�̉��>��\C���	{��i����<�'�1��x&FC�&e�-+7�K	�PS�"O@�R�p,�h��c
N�!��i����<�۴��?7-^:��Eh׋Z�]���re�&88!�D��p�j�"@	�咴�@e�&0�Q�T��	,���{��Z8%����p�	 �C�	w��h��M,b8��3��z���$�S�OK(���B(I�� 1�Ԝ[ Ԝ�"O�`:uB���^$1��ӣf���"O�`SOڄ+��ʄL�~gY��O��	D��<�L<ͧ@F��2M�l���C�ئ���	i?Q�"�5RK.!:�å8�RT#N�P�d�hOq�,�ǧ�z&��\�\�����'�`�)�N��B�:T�xC�Ol���<Iߓ0����3?��᪀c�r�F}���E���A�e[��t	���${�C�ɴ�^� ��W/\�;3�Ɔ*��B䉅���J9j�B�S�@8o�B�%~ �Qg�T#$����b�OSBB�IRdTq���&-�YJDcD�K��C�I��i8�NM>sI�ģĬL�(z�c�HF{���ǅBN�!7 m�H�p�gI�yRѻT�
��m�(e��A����'!h���Ib���xp�O9)�q��ŕp���$&�S�O��V� xU1�l�T4Z�� ���y����l	�p�\H��9����~b����O,#=��F��{R��C*�Ds���-U}8�$J�4i2�+i�ġ���M�$�D���1��:�S�'oA�H#a�;�ģp.�/�ƸGy�
v>m��k�S�ʬ�E�)�@��?D�hsC��}�ڹ����8���d;D��K��U+Q��+�C�)��3�:D�� ~Xi�;R���z֡R=g���"OH�j�eK-�T��^�R�����"O�)a�H�m����� <�4R��xR�'�9�b�ͺ0�����
.=)�(���?��O�,�R/[�S��I��k�
��'@ܱ9�!��3y*p����+1^\@��$-��?�n3C@�p��!��P�B;3�DC�	'{wXi0Q�Ԑ]K*��5I
'V#?Y��(ڧ+w��IA@ȟ{���f@C�,���L����w G6���:�n�'[�`��'aў�}:s&�8fHe5(��p��M���XK�<ai��Y�t�㋜�P���21�WH�<��ő���u`VnʉJ�Z�!ԫVH��$�'��	.�9���=��e����=+,B��
N�����/ݒ���Jb��c�ϓ��'��'�J]!,^+_K�����04�L�Ǔ�HO<8(��!9����+Y�uf@��"O�x؁$Vf�~i��	�.X,�}��Io�����E������#w� )�׀G+y�!�$�
�)�-��1���A'�!�R��|!ˀ`�ot��C"�/@�!���MM��oμZFHM8E�L=l����I�\��(�N����s�&øB�	�n�аk�F�{~�3��C?F�v6�:�d��ݖ|i��p" �F���m!D���*\�,���$S��<Ѧ�*D� ɇ�ʔn��P�T��T���&*D����)��-�A����d��F&D�xh��)�����(�"4�׭.D�l#`�]�1����fQD��#d�!D��Qt�I�9�r��V��I�f��M�Dh<1a�ӻV(��/ȸ-^*�x#�p8�H�OT���.�7[�$�:����<<�"D�t*fB�$wh�!P�+\�zk�$D�Pɷ�{� ��j4��)��!D�Ăq!�4H7�|B�̓g�8�f*-D� �jͧjI�h���^G[z���I(D�T�r�O�W&���dK+YD�1�Q�#D����K.B�	[�kC<PLV��2+#D��[E�ށuN`�Vi�n.�i5D���$/��䐸��ߘp�^��w'4D��{���37���q��L�VY� �0D����a׬W����A�?��#��/D�,K�F��U�L�@r엽D0Hu�#8D��)��]M�����?�x![1K5D��!l4!���*#J�	u4!���.D�D��$�)#��m�L��,-+qO2D�XpV��6G�2���&W>�vm/D���p.����0@�F!j�h��d,D�T��Ǜ*� �C�y���*D��@���zfv�8�,@�3�H��*D���� �?s�X�����-Q�q��#D�4�B]�	��x�V ���5D��z)�/X��$��%�F�x��6D���gEz�#�ɖ6��I`J*D����0i�lX;Q�8>8s�I(D�P�@g�-����"���7�P���:D�<�@��1(S���t�3:��:��8D� �B��e�����:W���a�+D�+�b�:X���e��f����Ѧ(D� K�ÃU��Y��"��%����	�'��<STd�3ʜP��E0*Dp��'�!̗�6���f�%xD	�'���e�	H�J����ݖ�4���� 
q�0�[�q����iQ8�dR�"O�XC�F�3�4m��J�"��"O�����T�tB��`ߦn���"O�q��`Y�R5j<��i�:���h��':��ĩ\�Q�f� bl% VT$[p�:[���u�I�Rx�%q	�'Tf��5�� � 0A0oU�Uz�dH�'4�Qb@�oZ��G@3|���c�'�\-
��'��l�_|ذ���'Q:��6��S'ĩ�f���-���	�'r�A�R�Ak��B��U�
���'S 4�0cX�'�&1�L��E��'V��է�����V,�\�'0�q�S�D�l���@�Ў]��'{���6d jL� �_H,�l��'~0�� �<�\Q���Z�2��A�'F �)Ѐ�<ꖔz��R07_ĳ�'�R�Qgc�%E�ġ A��%�.� �'�*�� �!q���լ6�:�`�'�ށPM�;�|��������
�'��kek�XT����r���!
�'��]=-6�$y��I�y*���'�X��k &o�1G��5%@1��'��9�d�= ���P�Ϩ\�B�r�'���Ġ޿-�����l۸B1�Y�
�'+� *�N�}˨�z&�L�;�FmJ
�'~�)��,�%x �yq 
�*�nt��'uh�H��u�v�iP���Āqz�'P�I��h���w (c%��q�'��l��U�X����M�"�|P�
�'D�T����;��)�e݌�-X�'�dA��h�쑰��[:fHY�'�����Z�P�\� !�(UH�'������V6��z�#Qr44A�'HHt�Mۜ� !��l��C
�'�=���V��i�J^?[���'m4 ��� C0�����Fp����'��@�B�<4�^h�c�7
h�x��'; ��ǈ�5^��5�s!6 ��a��'�P�;�'�^���V9|[*���'��$0fJ��/>J,��mz�(9B�'���MO�x���V��/�f���'OȽ �&Inf�� �M2��*�'w��'M�#��Q�' �;��A��'�ʵ����<z���i͝4:���'�l���(ܵ|:��)6&�<7:���'w��P�G�pa�i�%�
��U�'g )�d��as���0g�xa��'<<p�[E���ؕjX\p$i��'b ,�	��ٔ�Hz���'=�IS3��<������#A�����'�F��!�хC����*�A*�T��'��� ��)"��Pࣦ��1ˠ�[
�'��E�b���Rt����<7e,	`�'��AR�DM�a�����A�u� H
�'�.��c���ҍ	�(H�]�� �	�'H2��M��Z������4��
�'(������_*m��B�K�4�
�'��A���ޙn" �\91R)�W�)D��{��Fg�*aD�85�TY�P�)D��!�`ί2�]i�c�5�"�9d'D�,�K%o"����.�JBj11'0D���#`�$.�84m�Y�$Z��5D�Tf�	�,���Ώ8��p�F	?D���dɀl?����/��B�8D�� |]�)�D��2ė�b���v"O��J�d@�r���2O$}=���"O�]Bfd�`�
 �&C�')���B"O���A�H�Rf� l+$,���'���H[
���?i��$����B��00']�B��Dz���F~�����GQ��b����g�S��,Q��S�M��]��GԻE
�8��X8xB��>f7�h%��z��B�jW9n�TH��\�U�2h�/O�Y{A)��pX�&>�'�t�z���!vz�Qq
_9?,|+�����M�R���JAhR�h/���S�՛[�Ơ�GaĲ�2��v�X)�0>y֎R ?�� r@0=ހ٠�ˉS}r�و��FLƥ\L�8�O3� ��̎4f:<�Z�4�v����5>�P=�
�$Z^ʥr�"O���"�/zO&�I���4����ъ^.6��I��t<3m�;;g���ҟ���26��˳6�Bq�үS%=��+��r��{��'��!*�m�>x�@�B��5��	g+*���Gh(Y�)�a��q�R���h�{�N�r��4��>��5}���]^���Ǌ����ؘ�ڿ����'�J�2�P� &0���IP�N=��@���>j֐�q�N@�]�܁�&n*z�6�l�s7�'��ijp�;G$n���)c6�M;�'�6�[$V%��z��X5��aΧG&d� �ب`0�E+��Y'{���d%Lt��`b�،P��\��ݟL'��#&x�Z�Ѣ��!��{��K�5r}���ަy�W�|��@9  �,M���E%B&|-�W�H��Ɓtf8uq%m�r�����c��}���a�|8�fͶ_���8 �ؽK\"�*�� �T�����$%C.}���̵Y��h��Y�I^*��ת�<ѱ���EX%�׌47t�! E�'r|���$}L1��C�[l���7P?�y�6��0@V�0���F�-#�ߖh��ɮ��
�-�0�џ�{-�R�������Y����5OP �k2]d�0��^-x^�7�ڋ�n�Cfk�W�4圻b�J�`֯�F��S��PC��z��0�Z��kvXP�
x�VB�}�xYZ0捲`;�m8�n�%i,B�gI֦n��]bP�spɚ�Tr�M��Ok�o������&�4KM	J@�}"+M�HF�5�Fi�!yF�t)��T���k��7�(��d�7�V����X�Cs���QS����j�F��	��V��1�k^�]7�y�F��2]���w#"�p
�gc��|U�}�$L�4��ɰ�GA��t�ڗ�W�N��/\����ʱ�W���$��rL��'O�l��KA>D�P�4�ʐ~<��2O�c��4Ii�$�G�/�`��K�<N�H��?u�b�)f)��@���:H�� ޴V�^�r�
O���/�3?fȤX�EEc���;�!���~-���	rQJ�HvͼV�S�躼���:?�4E��1�H��$Ǝ8޸��1��A���s'�Ll\*�(�%i4}i�g��v�x�!$%Ǧ�q�F@R${r���֟@Pax� �	T���`d�9W�,d�9��O�Ȁ�
:J^��ӥ�gJ���2���hRJ=}��3�n$%S堚��x�c�Mb����:ƺ�3qk���D���|�av]�^/>��p��5�2;�N�]�'M-p! �^+�b`�R$M(s��t�ȓ0N����O(*:|(��A�R��[#�\�Dm����BC���5�	}����'�b��#ϐ�?�$XU	�&qD����'�f��s�m�r���Y%l�����l:	�&iƞ*���`raVxk\$���+�,����O�G�h�2n�`�p��D�?�ъQ+ԺW�q�����	@��pq���@�&I�ӣG�+L��!�?$����- ޒ�6�=M@(�� 1�IK��)(t�ߵX{r;�ӱT���34/O~<0�é��VC䉠mY�9I��?*t{� �=���6ř�G�\ٛ�@��~�\��ϑ^�$b�΀-�ƈY��-D��[Ƨ�|l5���)	��O�<�G�בj���pៈ��<��C���M�f�E=HMH�a�ϐ{��Г�DD�E���@_�
X2���N�>��CkW
~B ��Oܝ�# NК$DB�>+V��Qቪ3@����-�%Y�����V��c�h �1G\��y�k�'�`V_H�ɖ`L�~P�-Z�K&�j�ˀeTn��S��?A'Ȉu3��!c�%V�Q��x�<y��|�~���׮o�N���w~2a._�&���'�P�� T��y!�$�N���d�~QRE�;��S�j�Qy,m�Ї�5z�VC�ɱW'�}�Z�z��$f��B�ɌT1x+��[:�f	R̛�Z�B�	����Y�E�Bd���[�JVB�I�en !��?%/���j���B�II�����' ~��S�O�<��C�)� ��)w�Q�>��mV��("Oڀ� �ӨW��&�6@�"O�Y�e��@����ao�*V���"O>h;c�	I�}*�%�(bQ����"Ox���^=yb��Ό�[��@��B�,b
H(Ó_�N���FE�-���)!'�+�����_�F�z��Q�6�:����Y��R���E��`� �����Y������#5�6hE2��y�h����gⓠh��FR� L��!��77&B�.@Y�q�!��h�a�K �+2�ʓW T�1��,|�ҧ(��-h$!��Gwlܨ �B�+�H:@"O�hqU�����Wh[��xЁV�䐹=���� �-���X����C�h�;iE��1C��l������IA%�0�n�p���_\,}#D���S虇�It�(�`fѦ6�����K�E�̢?�`cB��T�C�#�i�u��W+�͞����35^!򤗌 �6�1pg�7�B(���<e9�I�[��=Z�ڕi��S�Oz��󆤏G�jҢ!73G�y��'�`+�@��%x4��ٿ\G��:�*&}"i��|����%���{2ኜ;�~	�M<Bl�����=�x"��94��,R9^ZDhJ���#KRū��0���k(.`�K!b�>��Bo׽�p<�!o�@>�b�h�W'^�!QD�r��	;g�����9D��1cmE�*&\xfC	��U���4D��0�C�_��,A�Ǩng�S�3D�@U.�ʰ�h���;uX��.;��xw�'���Vf��,ގ����	;E�I�'�����]54X��@�%34�[��C�+N�U@��'��e+�ϥ
Vnq E�E�M�>�j���\�>�$D��!���ħ�}v�9%���� gc8���\34Yj�K�2J���f���S�f,�'� �+P�xF�OQ>�cϔ19�x!�ֆ�L^v	r�H$D�hm'J7�P��ى!U�Em�����3Vʢ�K�3�ɘv�B��1(�9.�CQe۸$u@��D�u�Z��KUlV$��)G6���D�;�Zq���sT\Ѓb�.R�����ޥ�.4GR�ϋH�PK䣋z�S# �a���:k_HP{q
Ѷ/�C䉀i��P�UcՉ0`la����FH�˓T#Π�%mG#jӧ(��Y��	r@�� �膐)w"O �8�gL�/��hK�O�(qߎ]h0H�H�$�S����0��� (ښc��6U��l�r�٨px!��� *�^!���J�,;~�B/�q.���FU*���d��P���Um놴�G��<R�x�k�eV���<A�O:t�F����)g�0�Qu�GU�<�T)I�M0���RJ!;ڤH�⧆R�<i�	�YP!�#ef0�7�LS�<1G�<\B���RKP~84	�NPN�<��Q6�x�qd�r��� !F�<�1��R�dQ�1�H�=h4ᘱ�B�<�VO�w�V�@�B@=SÐ���a�<IE+��m�	���F�9��s��P�<�2h��	/���#;w(�3)Sp�<���]<!
�B�0U���+��s�<��O_�7'J}���.[�B]�K`�<A∅q�t���nҢA�Ċ��e�<����7iz�r4��4(�
��i�<�i��uI�p�e�m���j�<a��&b�� Kg.HVF\RA��N�<��#�q!���D�2f^�y�/E�<c`	);SNLxg&E�Mb:}�1i�|�<iU�S9"ijL�eǇE�Ĉh�O�<�Qd��(A! #B-`F���˜`�<��#����k��Q�a���v�<���-���͙bN^���IHn�<� �9�FøE�$��E�S�(<�""Oڭ�N��Pe��b��pR����"O�=a���X`)R���h�p�"O*Y�P�,�n���gI�i���;a"OZ��d@�7�H�{�%U�`��P"O�����٥NQ)�%S�9Z���"O<T�Ю3Z�t�Zq�ηA8K&�y�f �'�2'D�	��Rq䑋�yRj<v��Ud (
�����y&��I��y��8/�!��G��y���D9nx�`�(f�Uau���ygS����+4����q���y�	�}>��{�cK� ,�0���X��y�$�)�1��k���A����yBj<	Ș�8 �N�zo#�yr䇇Zބ��I��~��X��Տ�y�M�E���x��-]D����ė��y��y�F��#����H�	��Y��yb-ʘ�\��֙kA��	�3�y��`G� cĈ�8cF�C6)_�y�H���)��_�g��U9CD*�yBC�
`�2}��Qi�8KgE �y�D��"�����O�D�~��D��y�C�J.iP4�O9���0U��)�y���!����hͧI6����A���yBk�cSj|q�jK�7�} b��y��l��9%F7a��D��y���pT���E�t�c���y��'\�s��2ւA0��Ң�y�kƬn,�<ĪUf�tU�D��y�ĄFƮ�%�@�m�� �F�yc�	K���ׯN�V��l�&!ԡ�yR�LY��l��6W�z���mF��y� ZU��IU��M"� �e��ybOD�#z�<8�H�=?�V�xċ��yҏ���<
��ȗ\��(PC���yRK��\��Ћ�ƳW�ܰâ�U��y�`��*�X�!wf�X�3b����yZ�z�Z��$P<���+�e��\g��I�*M R�l�Ң.�[<���.W���F<\��a: 
g�8�ȓr�t�Av��y��+:�ه�~'hY�VIDu��AA��;/\��ȓL�.�;%J ?�q��|��]�ȓR�vtK���^��b� MW2��ȓ�AEDY�Ft)!U*͝#/�Մȓ,ƒ�r�H�Z�p��R 
�̆�3��;%��$ƀ���ĥ+iD���$n��;BB.�v��BJ�=�1���:+��uh�0��Ʈ>����ȓ&T	sF-���g�J(2�u��
{4<h�C����fQ�!��фȓo��PH7a��KHV�@��/)��!�ȓD��x!�Ďo~�x+W���4wZ����W=M~�5"OD�v�ۊ*o����W����G"O<�[� � ��ulϊ<���7"O�����5?/�+�99�1C!"O�t1�ů�=����$��q��"OX!W/ݙ;~��"��pZ"O�,X���v������-�TA�a"O�1�잪8�����
渹B"ODP�	O�*L�8��L�=�ұ�"Oժ�٬dӒ��j��.����c"O� Z!�R��n>5���UE�(�c�"O
<��ōP����􇙿0U��qf"O,�#��ԫ
B���I�6E%�w"OE��J%�vI���Аp<p�t"O�)�7Ć2�Qa2��/,��X;�"O6��q%�]���C�^�+����t"OPbr�J
t��8âT���� �"OH\�']-�0�!\7M�9!��'?x��͓uO�I�Y"({V�
)L�W�F:A�B�ɪ,�8a�Q�r< ���3hYlb���aE�j\f����S�j'^]�eeM����j̛n�rB�I&I+�� ��j����*���u�:�(H�.O�Ӗ
"�3}�M��K�H�����0^���sڠ��xRIĴ�R���ڸK�`P�䇂�>]LT�h��KF���d�'�,�㖎�5i�,�AL�?i�L�	�4l����M�9c�X��'�%iT)I="��BL�x��3	�'���*�A�a�S�#ܒu�B�(H>A��\�s�Z�HpoʭÈ�L�	H6	�T(*5�O82i.`X�"O0�b'J0,���5!�M�Z,hP��-pδ�r,��[���t�)��j� �nE����M޾ 	�Y��I�����O^�`���+?�A�o��J�����U�ȹ�R�7�Ҁ�di��B2J��$�Ϯ4�ą�.O�
q�L���O��#����z�p�I_�0�`$	:3r�g�2mD|q�$�Q ؕ"F۲g��Q[��D���?�1*�*,@:��dĐ_��H�a���|��R��ND��ȅr1�j�+/H.������t�W�[�N��55Ҹu,��z�s'�n�<ᦋ�>,0
�`��?�T�T��$o�D����шq`���a�@%H�.@�?(:� ��]?�@�,OZ��"�C�(�4�.+f�Iq�'`
��FK�m�L�Z��^�#�taV�z{ɐ���Ԙ�"��WF}�$ �؜�d�UP�'�F8;�]�c�vPs"�6�Vq��{Bb��W��LREbY8S��4C�S��Eө��sm�<6���w"цlV�5��4М�����7!���
��*֬D?"�ܐ���/�>X1��P�a�J�3b)mݍ0�&J)	VDPz�س�����VF�F}l����
�
vT��O�8&_�]����F� +l��2��NO������٩n\�R��+F�h�_�p��@U�5jT%��W��`���%xG�렣
�d
lҰ� �f��IdN(Jt���+8@Pf��5��8��! ��spCm�"	A+O���o�f����E�F:�H�
��W+���Eo�7��	*.@N���#��?aԤZ���
/F��dUJ��b�"B*�Z��$"D�n�0s|d�J�o(<�6��4�8��(߈<㦌k��eq�KA�6����mI0h�\�%?9����p~��{�rXhE�܋��%.���?�B��}�<P:ȁ�FЬ�c�7U�T9�cI�'0�0�č:;�D35�բ�0<i�޷\�J �blW @ZX�*U�'�x�{A䋲Xa�	+S΄:4-Z 6/\U���$]�� ���c_�J�O��y3u�ZxRw��.T �3R�0K�I\?5�L	�΋/t�a�����|
���<��|�tc�:��uVœN�<ӈڭ4���G�.@6A�![�4���sJz�~�䓵c��$?�R��u~�@���-*��̛CU�hc���x��@	I�(`��.>8�& M�Z����Č��aA���l�`���_y8�10�y@�G�f����6�H�y��xB��1K��zj�3$��M/l�Ԉ�ǼP�H��V��.7� ��v$�)_!�0^~�S��Ԟm��=�3��w±O�Ă����1F�P�O��Qy��d`{K"_;B��E�
�ތ3�"OARO ��㷩�<Z��SG�L!��qQ2��9{�0���h��W�q8lq7 ��G���yGd�a�!�$�^�� @W9k�9��C�#���
`��f���:>8��ɤ4[�b��W
>��c爠O	����:p��4@ѧ2Q�d[r�ɛ����$I��7�B$�fn���x�K��&�4�z��ׯY��Z�G��O ���g'GRA:��	o�g�H"'��wq�`u�� C�.l���Jq��A��Єˁ��x�C��PhH�q��)�)�矘�#ŇU:8]X�#]�����l;D�<��+q�n��ADH��423O6?����	0��a�@;�5P� 6 *d�F�Vx����_���� �GC�lh�ł8T��H�KBV�!�?_�j�@�	�?B62��;!�� >h����
y�(⮀�#�8�P�"O�Y�d��ҵ���L�l����1"O���p�.Sw�c�Jō Bj\+e"O��J�O����`7�H>l�\���"O8�`ՠ�l�ΙAI98�y"O�T��#Ǔ=��4#AIC������"O�%�Dd�3B*j���@(&�:���"O⡨�Dąo�}: �ϛݾ�{5"O��C0�E�HW����A�P�B���ƨa����	Ó^�<PELƽl���Hr`�.S����^�4 '�ӱY��9�a�V	Lu�@,ܸr�4����x�����@�F8he"Ѐe�J�D���d�U+���I�S�L	z�P��Q�:�@�fĭq�\B�,��a�cD�={�< (���.*!��ॣ ���e��ҧ(��YV
2x>�y
�2�U0�"O(�˶�ڧkT�#����8�d���-}�d�t{8��U�;��$\� �*� �@��7��C���⋜�%����B�e�D	9qiؤz�+T�Y�-s:8��ɾG�Z1�  4A%a�S�̢?y�@>4��$D5��ʹa � 3�U�f-����+X!�E;�T��.Z4bʌ����+,]剻jטyx���t��S�Oxh�1H�q�̩
�C�	;����'K����	e�:�2�N6:䀖d)}rj �bh�Q���{�d�c�~P)ǉ�p�ґ�P����x�$'a��9e��B��<S��&=̬1q��N�RG��G.l$�t&d�o�^�E��=�p<)��p��c�D�B�0jQ��X�֠IqRi���$D�0S	�n~L3ţ[$M_2Ms�,D�D ��$ j�B���
=�TH�A-D��J'K�3J�}��Ҩ;ܤtI�*=�oP��B��'���^�ʽܴ#����O�1 ���#��J��S��0��)������?�thO�&NZex�F I,��1+�i�'�,Y��� �$>U��V/z�MX�cA��� �Q
2D�|A��"��%��M�?
3j��TB�<��̊4 �<옵�2}��I˸d���sA^_�*�C��&Z�!�	,E�Y����Uݠ1e���p�b��O�U�JI���qOf����L[XIK"�I�_T� �f�'dl��hюlA�=ئ!��*���ełZTݘf$ZC؟\ c ^:j�D)�v �>8��Yx�&�y�Yreh[���]�4�^�\�,���R��Ic�"O�M�w*ѯ`T����t�N�;7_�X�"�8
����>E�DC�gۢ���I#k�)��Q��y'��av�8�O����`j�`ֿnr��' ���&�|��ϸ'�~�S�X�(�(���I�nj��	�'�z�3���PR���OW�ڪY#1��%o*x5�'��d�7	��g�����C�T$y	Ǔt�R���:��9�00����#�Y�Q�؅s�2B�I$W��E�u�)��Xe�)L�ZB��L|�%�3h�h���U�7�&B��͸ i�@.p3�@�۔P��Շ�n@�E���U�\N�0�KK�m��h�ȓ��d�b�V�
AHڗ��,)\�ԅȓBxdP���G�������z��ȓ� ���O�"���#0�[�J'<d�ȓII��r�À��q��/Rw�̄�dڌa���^t�2%�2;b���ȓ*`8�¢I̧um����<��(�ȓy�D�b �s��䒡iB�Z2q��+�zѩ&�!of� �V?air���[��L�$EC.p�� �!�>h
�$��Qhr5��E�(�d�c�#�\\�,�ȓ��V�E�������Ea���[]�e��J4/+�$�tj�U|:\��S�? �%�ӂ3(1�ىSGP�M��A"O,����]$2>=;�>\��+""O�1�뇴3(�P Sf��6<����"O���b��0:=����ft�{0"OH8��7ؚ�Y��g��@i�"O�d�m0���5��<��XC"O��mU	6Bq�Cd߲�"O�J����y�f�2�IW?`�\��&"O\�h#��$$�T�$J�*��D�"OD���nà���j�
PX�1�"Op=q��S��DU+�)��H#���"Ols��[�Q��l�Ub�V/�4�W�'u��R���(I��SU�Z Sߔ�s��Y�.~\d����53�`���'V��B���&̍�`��0No�Xd"Ox2�G�;7b���g�0H�Ti��"OD����	#��yxƄ]��,ɫ�"O�$�1��9�+Q��o��	�"Ò��&��eNX�T/�!`��J"O�0�QaD&~����^�#�0"O�mK%m�zd.R�4�����	=�HO��$�jJ�)]@��J��3��	�P�L�
m*1r�S�'���#7(��	�>RR&�Y�@�v�5z��`^��+5E]y��II�uMVI���ǴNc�`1R�٬Nn� S�Dդ^~H�'�8��� ��� QiX�6���+DD�1o�D	�윏��	�"�v�q��?�i�&i�-0qȒ@��|8�FL�1T4Tb�O� ��ƃ	6cx��
�'LM�"�U� ���3�Q�y�5�'�@ �P1��ȻN>������g��\ 
�1p�=�&o�I}�B�Pь��=E�$�ٔI��[᧓W�����%V;�y��Qz�����k +En5��'��:��S��6D�@Q�MB��p��l�9���'D���b`?M�$[E��7���3�$D��z�Η�Ń�ć����5F.D��C���$K:��6Ʉ*Q�,㑃-D�,��B
u��C� D�E<Ը!�+D��{�Wz.���m��9�s)D� ��]Y�N@{��[<��ܢЌ:D��8t��;����v�X�hk|�@	4D���V��)��1$�X�
G.�c��3D���2 &4N��4�,�$�&&D�4�ܮPHv�;i��v2���, D�@ㅚ�!����b�/� 5��<D��)�O/ ���G�}+J>D�@���'ܰ(�t$� g��3!/D� �"�Cy��:����j1iG�8D����+�d����)F�_�n(�B8D����{"�sD*C�Wn���B6D��	� S5S�*QZuk�x�zMh�4D�@q����S,�{�A�DR��0�H7D���f1�`1yӦ��wnt�9�*D��p'�4dҢ�IF��C#V��4�"D�ل��=L�֤��D;OW$1�1B;D�xzCb�6?�[�CiP�H��]�v�+D��h&�1��,a6�A$��2�*D��J֬�.q*���B�(7�`;�k<D�����{D%CvmT�,	�pc�'D��+�oCC1�mb��M0@���r�/D��A�ϖiEyӧ��	�hi���"D�dZ�`��zs(�j����N�;ь?D�\�C�4;E�1{n�IlިIRa>D��c�/E8�T����@�1�$R�� D��x�%O��y�Q J8�j@�d�<D��˥&�P�Y{@G�%��q"	?D�x���$<�L��7j�
���"D�ԲSDʡKR8�C�' =]1�@9�D?D�� �,�cIR'@ܸ'�_�;h0]�"O pD�87L)b&��)h�`��"O(@�f��Q�.9��� �cHfA��"O��t��h��xsm]�F��"OP�ڴ��+����,B��P#"O��hR���J)�İ#)!CR"On}�A��	\B`|(CH��T �$B�"Ol�cCa�c�6�.�R�"O�m+5`Ҙr2v�S��)t��2B"O<�+�L�"ר�*S-�� 邭��"O(��@@�.Ka0a!�,��E�nx�`"O�Id�A�!���d��,ժE�D"OV�ť�)4AN`���]��@t�""O�QukA�+�.��0���{�$]A2"O��%&�\��y� $�lI�"O� @�D �
0�շF�n��"O̚�Ojb�pѠ�9&t�h�v"Op����84��ҷ�*B[�9�"O�͠#�%~��)z�OK�Kq�{�"O���dW�^t��0�G�ϊ��b"O�h�@%-i�n����BQ���S"O��1�ܔF1�a�&�Ƣ43��!E"O�\�gC
NRh�
 �7#^�"O�t�G�7g�$b��<�"O-��]|	v Qf9<
\z7"Oze�aE-Z�DD�.R���%QK�<��f�1N^��8alѷl�2�PN�O�<AEO�+ʠTˠ`�FLn2Ӂd�<��j�,��iQ�ķO��Hy���\�<�4 U�JMQ���כ�]Z!�D�<#;T��I�H�l��J�T !�Ɋ=s�`P¢�#:$�yb���~!�d��G:H� Q	��G|�%XCaM$i�!���m�DbpU N$]���P�����A6o.J$�ǉ$�"�⬈�y����4�Х��	Q�E{e�)�yr(ĉx_�d�T��-O���o�y�a�4�!3 ��!�HZ�m�$�yB!�O��hA�.u�����X:�yB��7D���I�S�y�,��6��+�y���c��Y$�wt�!
�Py�ˋ>]hѸv�Y��X\`��Rp�<��ᅀ.��X���'|X�HVi�<�B��1H?�Qi$D�X���[tIJq�<�b��-~l՚���9z�Y��̑b�<Bn�J�C-�?�T��!�G�<a�j��رW�U�f����a�E�<�N�-X����b�Ab0��1-C�<Q�낂r�
A�a�^�(�J���c�<��V�%��q`%ǞsD�P0I�c�<��L�[]HsQ�"A�4���Le�<q�^�k���ɵ[7Z\ѫT��k�<a�P,/���2ȚwZ�-2��p�<�̢2 ��С�\ z�|9ƨ�h�<��@ߞi��km��=|�BG��d�<�d"��S�<[#b
��2��%d�a�<��'Q����Pj��ug����e[�<�E�<E���@�OO�>�m�T�<Y�-�'���z���u�R�[��YZ�<��T�����!n��\�X�R�V�<Q�I�7%�>@����'�|9�QR�<�ʒ�9�H�C��B$bh;Cv�<�&,��z���#��yZ���*�o�<���]1x��A!�Z�m�@c�[i�<� H��î�?f*.b���C�I�"O�q�T��5@ZVa v-D�+;�=R@"O`���W"?>�Q���݇L*��R"O����$x� !�ϖI"(�g"O�@sp)C !x�1!�7:v�|P�"O��#��DF�|Y�J�9AA>��'"O@x�G�W,�X��U(	�M+&T�R"O�:�/�K�6�Y�)�,���y�"O��dʹz0��H��o�� 0%"Ox��Q[x�|z1���h�z���"Ol�XO']��#�j�2���"O���Vg7t`����ڎN�
HA�"Ol݃�f<H���ZD�ɖ3����"O�|K�!,���61?�԰Y�"O��ã��y�h��&ުb�����"Op�r�Č12Eh��_�4�X{�"O~�B�k�w��p"�
��U��"O��͕1e���G��|�n��"O^�R�)�2a�0���1[D��"O!��kÞU��l	ƥ�|��v"O¤�SD؄/�:��7d�d�cG"O��Q�@O�q��!%y`�B�"OD�qr�٢]���H FXj	½��"O,�u���V@�S�M� ����"O��[�@A ]r�@�'�T�E"O �#�$0������,�PA��"O^�˒⃅"ul����]GF|yC"O��S�/ٙ]S���D�hV4!S�"OtD�6���jF�+zh"O�!䦙�yil���*��<���[Q"O�W�� =�(�F���`��5O�\�<q�J�Ȝ��
��7`H�"U�<�RoQ�^?�E��?x-�C�F�<iș�*햅�� ѕX�:�	%OP^�<Q����wy�k_�HCL���\p�<х�?aΕ�َ8���a�![n�<�ؕf��ya�E�|���$i�j�<�G� Exp����$3���_�<�"T1"_
	i�ȅ-2��n�Z�<�p/�v�#���9� ��J_n�<iV�^>=\H��K${ܚ0VO@l�<aը GvbY�V�ψ[b����R�<��D�F��`�_/��r��N�<�⌗l�R�����;��)�!B�<6a��4�< 'E��.�uk B�<!� �2Ԝ����6I�Q��"]@�<���:a�\HV��V�~�0���p�<g�Jhd�C�F�s��l��#Ul�<ɅH�)�R@���nխg�Yr�"O�V���0���MS�P�8(�"O��hc	�	fBB`'k�#p��j�"OB��'@�
{'����7����"Oi��D� _fda"`��#�\5ڤ"Ov�zf��H��	/�tt2�"OFT"�n�>?�8�2σ%w�p��v"OeA/�4����P��/�.�8%"OH��.U
�4htC��W�rmX"O�M�b^!Y�4�QC�	��a"Oh,@�f*y��M�S�ʩH��h"OX�������H�!��9��١"OH�3�ڧ�(�!k>3TDD��"O�!aG�X2,U<�0�I;IT�\
4"O�e�.A�!G"|;6�Т=~a�"O�t���:@c4��ף�m#N���"O� ڰ��Ȫ�,��֠8"�e��"OF�6�4W Z��d
C���"O���되=��Iʱb#x<��"OT��mEsI����k^!й@�"OJ�� h���� ��#=f	:�"Oly���O����1��7��p"O4�Ra�̩	�@��G��`�Y`�"O��R5d��>z�$�֮�6��d�G"O��AI�0`���s䋡S�B	��"ǑK%�@�A�ܜ����@�P�i "O��S�-H�n܀UO��6�����"O������LI�9���E}xx| 7"O���6D��DEd�΁�^���"O��%̉z�� ���^�\ &"O�-P@f�9.5ryȵ1QT$���"OT�P���,ܪ�`��a�rU"O�D�&�#�J�(����q�8�"O�� M��]��͢��G��~d:D"O�Q��TY(�Uӵ��_�"�Bc"O6,K+ې$��<���̭:���xw"Oj�h�

�Q׌X
��
;�����"O`=��S!��D�3���r&"O�9��*֭~��o� @c�`�q"O�a�UL�0�o�\q< :�"O�hsq(D�9;Xh�U��uYH��"O"���O\<-����D�Ԧ7=�]�r"O������#;�貁`�'hD�1K�"O���H\Lߎ����\"];!�"O��x��B�^���Q5���J.؍��"O����/D�IC��&$^�V"OL�	%	S	H�r	7���T�f-{�"OSWJ�~p9K׍	�d�֬JQ"O�  G���{�8�9�+A��` �"O5��LĞ�
0a�Kʝ^�p��3"O��͖�8��agJ��N��0"Of�!WG�Z�>}�hײ����"Od ).!W#�S!B��k�LmP0"Oj��ǊJ�K����@��O��Q�"O�����T5YN�`� #��y3�"O��dO�'䙐7��eH2]آ"Ov#��2{z��R�ͷ 88i��"O�L�`   ��   �  O  �  �  `*  �5  >A  �L  �X  �c  $o  �w  p~  &�  Ǝ  �  W�  ��  ܧ  /�  ��  �  k�  ��  y�  ��  &�  h�  ��  ��  }�  ]�  � � � � �!  * �1 "9 d? �E QI  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(��I|�O���#�H�R!��њ]��p��'_��uʆ�vӲ�R�c�*m�'�*L��܉�` ��ڭ\�����$֮w4I�1O�,��g�W�b-h4��Ӽ9�HMB�tX���;%�2���IЦ�Fx��2R^zmC`� �p��#�ȵ�yRO����!�L�q�tR� K��$"% �"|���6U3��B0)зez��%�~�<)0��.)�#U��4��뵥�T�<��۞@J9������
�ĥ�F�<���R�}��%�	2a ��`j�<�d��W��aP��ۆ&Z<�j�g���'o(�TA0g�]j�ȺS�����'���G U*=�~@�g��J��p`�'X���	B�z��X3'�R�m�4u�	�':��D�K���@ W/�S<������ �\q�C1������h=�A�#"O8��N� Gv����^�g �<#��>���tl@aM�/Dc��2X���ȓp_�B�"'���BQ �萄��N5[�œ�J�lU���V ��-D}�����Q��*�	��ȴ�� �C�I�qv�d��+̅Z�����슃'�B䉌�����"� TU��gɭ 6#>��C?�'w�6��![�.v���a(3�i��j�X��`	O̙K�aX���YΓ�hO?!F��*e�@y�FP�@�XɫA0D��:4��(N���q�S�/�����,D��z�K��U�TǄ�'TI�9�+$��g0��9�� �:�����o ����9P�M���4t\�\����ayR�O֒O�0���xb�Ӷ���V�{�"OQ4�B�|;z��&T���S�pG{��	�d�\@A �K���)��/�!��>P� L"��"GBi��&K/}�ttFz��9O�I��rL,y`��hX�xp��'��+K�Q�����T��������1��]m��<)�]~��ʆ�&O`�3�X'>��1��	k}�K>!B�;q@ηn��l����yRaA�90�����Zcz����Y���OL�~:��N�8aޜ�A($}�q��a�c�<��R;/xВ��E-�:ѡf�c�<Y�Y0�����j��u�C��i�<��#=uL-R��	�+($Q�E�]�<񳋟�%D��O�g��,P�I[�<��g�&�:�r&l��G�.a��&A@�<6��_N^�R��:���� �y�<�w�ґH�yz �3�`��� �j�<i7�}�2٣QO�p����2��q�<�5�̏�xq��T,�s�F�<�#��![����UN�t˞�b!W�<��k���≨��Q &Р��|�<�ƤS��ڑ�UF�JIj3�Mq�<���ߣ��� �M�1vN�Y©v�<�q#����g�)��!��v�<ag��R�F�� �>���Вd�V�<�����Ttހ	�[\��,3aL�i�<�a�C�2��-�I��T��x���F�<q3 �jT�㶦ւa�j0I�~�<a��WB�<�S�	?sC����j�o�<�"��P�:���=bJ��&��n�<�/�"��ړş6K2zD��c m�<�6�P�*���^�B�ވ��ŋ}�<I���1�0��#�3c�R͒��LS�<�$o�^ľQ�ԀR;1�:�Ns�<�d�)0��f�g�����/DG�<i���B���UB_�&���SFG�<i���b��C�Hܭc�����<�k��FWL�#�M�%j(X�FE�<�ä���8�d��&J ��DoV�<s�T�\���9�2M���Q�<��/	�P�RfD�<��l�F��e�<���G�#�H�1�K(v�d�4By�<qB�"J14Y��͏%�B���t�<�PHZ�:0v�a�U�E��!Y��p�<A&	�W�� ���~tb|��o�j�<Y@��.k�:��m�9pt
Q�5%f�<Q�4F�(�3�����k�'�F�<����r��t��v�J�{F�{�<!ݚa��	���.����d.�z�<� v�B_�0�q�� �f�2���"O�}p�4�V%Y7b��i�!("O(h�`�lB���5�B�	��""OJ5�f炖l��1��Åw ��Ҵ"O�IȒ��&$.i�Vo>)#�ı�'M2�'�B�']b�'V��'P��':L�Ye	�#?�T�*�j����ͻF�'���'���'N��'���'���'��q��(�.mZ���x��1r��'�R�'���'SR�'.��'���'�:�`I޽f��PmK;�8h�t�'�b�'�"�'?��'b�'���'���# ��4a�R�QB�Ɣ�f�'}��'���'q��'�r�'���'s.�[ukF<7aq����`%6���'���'2�'��'w��'/B�'��p�D܊o6~Z3�E$#d����'���'b�'-B�'��'�"�'�8}�#ެN:�J�MI�?	����'Q�'��'��'b��'7��'B���
I�s�t���ع5sx����'�B�'"�';��'/R�'�b�' ��J]�<�K��ӧc%tQq��'��'0�'�"�'*��'/�'�b,!a� YH�,ܲ4��>�?����?���?)��?����?���?���� #�d���B ;�
1�A��?���?i���?1��?y��?A���?�r+�
�\��,O=4���+� W�?Q��?���?����?9��k��V�'���Y�i�"qR�)�	�~��5ET�3����?�)O1��I��M#�O�(���h⦇Vvb�S�"��'��6�.�i>�	ݟ�P��f�~�d��Vp~�S�M�ڟ�	�a�zym�[~�<�:��S\�IDL��i��.�� Ƴ"��<�����/ڧ��sU�8!�0�밯��J][S�i���y������]
)����t��r5���Z22��������i�4Ҳ6-y����]�[�Rsd�(��v��̓5Fr�Rp�����'�N���W>hӚ����� SΤ�R�'��	g�,�M�K�N̓n��.-k�̺ �QI~��{�Mw��t�������	�<ѮO�x���[�"�Y�#�V,1,dhǒ���I=F� ���/�S�GҎOݟ��	¸� �J�/V8�SmxyT�<�)��<)�C�*����c��O���3�+�<��i-��1�O�Yl�G��|2�ꙷhHQ���N^���Q&��<���?Y��Sܞ ��4���`>���'煏�\�}�"�L�m[l0Bt���b]"�Of��|"��?y��?a�t
�2T/�D]�)�Ĝ;]���p-O�5lZ/u�����4��b�����$d�*PR�*"i�͹�*X9����ڦ�*����S�'U*��P�h%��N�B������x[���<)��*1���6���򤆱Z��rF5�����	FL�$�O����O^�4�0�Sg��*�7�
#�Fɑ���v~��-W<-Ab�v�����O��l��M+B�i�F���� ��h�An͸7��!�#�H?����L�F#,l�����$9!��ɭ+ ��$��YoN`8t5O����O��D�OP�d�Ot�?a����h�3�K&3���v/���@��d�ٴFk��.O2�m�t�Ie���H#��Ք����Ncs��YN<ᴽi=�7=�TP�u�4�3ʒ���	=2��x���N4E0pe���DR?��d�'����4�:���On���{�ƥ(�	QZ̈���兦y�@���O^��2�4R�7�'���'&��5d)̱d���WF�qY1C�)\d�$����M���i(O�3@(\X�-��&�����,&8!Ԋ��pn����l(?�':���dې��a�l��ӡ�.�r�P�&#�j����?���?��S�'��Q����ANW��p0�kb��ӣB9y�v���˟T��4��'J�2�b�Zܼ}Q���<;P��+�O�~��7���EqpN����'ܾ�Su���?駟��k�(QKnD�&&�}��Q��>O��?���?����?�����	A�Q�F8c2�P?Vu�b���$ �oھj��������B�������Ӳ	I�@���$�d4{�:m����a�4�&�b>%�t��Ʀ�Γ^)��	g���㉌./�(�l�Q a��O���J>1)O���O`����,	�ʜ�׉H�W���X���O�D�O���<&�i������'t��'���@Ř	
��)S�`�#R���'��_Y}�'M��|�j�jz�/hP�YRGQC.��#�OJ�.�ƌ	*�8��O�Ę�	:z��+\#Y�1p읊/��(���_��'�"�'}���	�V�%0�U*�ʅS-$d�U�؟��ش��]���?�c�i3�O��8"b�%�3S�%�F��W�+1��d�¦�ٴS�V�DQ`�&���Jפ��Vj�E�
9��1�F5	E��D.G4BP.�$������'�2�'���'��;QG)S�����+p0�R'^����4M6�Y����?I����<1chٯ>Y��p�CE�M�6h��<�����X�I7��S�']Ԃ��o	�<�(*A%��w=j@q���h����'�z���G�П,���|�W��ا)�2f\�H�G�5b@�*� _����I͟��I��zy��r�r䊓O�OB�⩌�H!�U�����a�O�TnZy��4���ß��	
�M�S-��W��)+��K0���Y4y�%3�4����J��\3����Op� ��QHV�(�8ĉ�'8R����9O`���O���O���O��?ɘ��ي�@���@��}d�5Ӣ#U̟���ٟ@Zݴj掠�)O�og�=�����ߊ��@(�"rm��eO/���5���|�d
���MC�O��!Fm��{4Ht�IR��#��52������v� ���<y.O�	�Oz���O~���gW@c��q
���t��O`�d�<q��i�"4�'G"�'�������1��.���yd�^���8K�I� �	���S����n�ja�rF ��:���E.V�P ��C\�L�:�O�	8�?�u��O��Ӓf��HЌ�����,}i�{�ͅ���������b>=�'��6݁xFr���,5Zɢ�s�`B�#��btD�O��D���]�?�^�����~蘉ȇ��>u�^%��`�
o����
�M�B�߲�M[�OR�V�:�*H?�0dFԽ^i2i�qӈBt��{�ؗ'"��'2�'br�'��S{�j���
��$:��bo��[���0�4
@�+���?	����Ou@7=��E��=WE�<:�G�&�4�� m�O���Nc�)��&'���l�<QÅ-x�|�AG�H!|���d��<��nʷ~�dG/����4�^���%����˼>���YG�����O��D�O��ac�6	\�L���'^��
K��j�,�qQ&�JQ� C��O���'E��'Y"OHIǎ��`e�X�@L��P�咟�����h!~p���/�i$��Oɟ�Y4��9�HTbA�ֻ���ȟ0����T�	џpE�D�'n�0@ʂ�b���E�%uL �P�'M6��C�����O�hn�R�Ӽk o��z�r3ρ2V'
�##�h?���M#U�i��{$�iC�ɩU�A�A�O~&h0b'� �$��e��g���A�G�F�	Wy�O,��'r��'4k׭s�l�9cc�9j�ve�F��%��	��M����?Q��?�I~�Fe�p@$õj�$����1X��$W�T�Iޟ��H<�|��V� o(E�&�8=֪-:���4�̜H�fS@~B�1-|���	� ��'}�?;Jh����/C.A
B�~���ԟp�I�d�i>Օ'�"6-�	u����3	���P�y05!�W�j���Ŧ	�?IP���	֟�j�4 <��g�n�B���k��/ �������M;�O��Ф�����$�w��=���C�j�����nǴ�rQy�'	��'��'��'��ء�.~|
ђ�b�.;�X+c��O��$�O�0nZ�E2N8�'�F7-.��H�?�d��F��(7V�o��N��&��#ڴa5��OL�}��i^�I�X��C�e�b�Yy#�K�x��Y�T�?fTb��U�Iy�O�2�'��gU[lr�H�կ|9I7 9ri�'�I�MKdOǭ�?)���?(�z���G�M�f`�3�Öj��Ý��x�OmZ��M#�xʟ��¤�\��uBB+�~���+5�Z/�>L��.W'.��i>���'H�a%��R`Q�]^X8Cb"Z9h�4��Z�p�I����Iԟb>�'�t6Mȿa��`j�"�\#�	�,Q�+���?���
����D�u}�t�J�[v�P�`�0�j�ı0��!Ū���1�ڴ7����4��$ѕ:��:����S�[8��Do��{J]H"kN�h/D��zyb�'I�'���'
T>UHWk�m��2a�ΦV����C�̗�M�vHT�?����?�H~��Xj��w�b8� ̌U�
����`Sj=�#af�։mZ���Ş��|2�t�;���m@qQM������P���hC�j��,TF��Ly�O��c��m_�qG���h���4�F�[ ��'��'�剉�M�4���?I��?�S�0"3\��q�ŤA{����	I!��'���?���Ez�'�I@��ەM�������>o�� �O"�1�!�F�KA�Ʉ�?1A��OLD:�ǌ�>f(��c!-$�^����O����O`���O~�}*��uV���Ūՙ��H�Ɉ%^)�t8�����M�	��	��M���wr��R��1���8A!_�f��R�'��'�7MC"j�6M7?���K9at����,�"a�C k-j��n�
PЩ�J>�.O�	�O����Ov���OB���+P��pˑ܀WFy�Dj�<A��i�pI� Z���IX�Ο �pHR5,Bp�C����e�h���B�����O��\�)�S�	=�e����<j�� �߄�T��V��j���$��O�ՒO>�,O�����ٮ\:�x��
2���K�
�O���O����O�)�<���i,n `��'dؗ�*Sx���GL�ܸ�YvF��?1B�i��O�L�'M��'a�@.|�B$�����0�H�&w�:8T�i���"q��u���O�q���+2�4����VV�X�����d�O��D�O����O��d5�ӵ0A�LI�c��K>�d���ےF�nQ��՟��	��M�-����$�M%��1�@�JsP�Cw ɡ75�)�Z�ēm�F�h����hϛ����1�KE�n��s�ڎm��D(�f'i�2��@�'٠�$�З��4�'�b�'�|�e��g��R�	��5>@1�'�"^�y�4,Q��:��?��������$"��H�L�v��FѹqD�����O�6��b�|���&.	�I8�#�6d(!�A�EL�8m��n�<�)��dD]؟S��|�璾C"p�2�
6*@ 1e �(M��'�R�'>���Q��8޴	��$���'��$A��W�9������?y�.ϛ��dvy�i�\��J.By��U�S��S��e�J�m�z8l�}~b
:Bm�z�� 0���"S��"�.��K�X�:�>OP��?����?����?�����	Ї,���� ��p���b��$̔=m��=x�,�	��x�	b�s�({������-v�5�a�A1�!h����?a��5���Ok�����i���G�/���4c�B2�X$@�D>�,i3ؒ�G6�O��|2�X���"��O�[,I�Ei�<a�� P���?i��?�/O� mZ&1�	���I�G���PC�=�B�!�%Z�Z��U�?q Z�hH�4j!b�x���5A���HWf].�pB�AB���$̺�=��%��@���)�������M�̚T�C��_�F�c�Z(5����O��D�O���*�'�?�IӀ91�m���#��0�*3�?��i�VUsD�'���p�r��]�b�\��IH�(�R�gڢ-X���	�M� �'����S�[b�柟�BTo�$/W���&%��t'���
"�֕m��$��'4�'���'l��'�`�:$��a��MC�N˅NMvy�0]��ݴ5HqJ��?����O<�6�'a���&��JƲ�BE �<y���?�N>%?��P��:sAL9��OO2���r��'yu��2�ĞQybOȻv����I{�'��	 }.��ʦ�N
/Ҽ���+.E�T�'�'��O����M��*�?y�gN�7y@Ձ��2`�|�� �?��iY�O���'`�7�������4D���:�	��W\��A/�K�Ę�#X8�M�O$qX�������w���3�\*i,`�yVi��&@���'b�'���'�RQ�b>Z��B w��SCM�0���:dE� �	��`�ٴE<V��O��6M:��*&�*!����\�.m �t}����xr�'e�O���i��	%UH�!ae�0�Xq����߆���Q���P�IXy�O���'z"�*N2��0�H��a��Ȳ��U�T���'��I�M۵�Z'���Oʧ[��E1�/
�kMdX"MgQ^��'ȴ��?�4G�ɧ�)�z 8-x㨝,q��J� Tcfdq H��\�jǕ��ӕ"��v�	�D^�q1�Z{��!�?Np��Iџ�������)�Sgy""{��X����&:,��_�{V)@�����vқ��d^q}�'�� ��"�M-��'��J9�'$�6��1T��7m.?9Fئax��-���V-'����S&yP9PǭӅ�y�X�4�	����I�\�Iȟ��O{6<jW@�N�;R�Dq�@Xci�zի�#�O����O�������ͦ�ݺC��(�&Ѩy�AT�7,��ៜ&�b>9j�.�զy͓bL@�ToT�Nb��.\�H��̓@��ux$��O�u�L>I,O�	�O��#����1�2Щ|xV����OP�D�OZ�$�<ǳi6y���'�B�'���葭
�}�d��aU1'!��;t��GQ}��'i��|r�ޖWT԰��W�"�ʕ��4��D���XqA�ïlj1�8\Y��ij��Dٞo3,H����pXT��;����Ob���OP�$>ڧ�?q#d�($�|c�g�'	�¡&B0�?�@�iTt���'9�j�4���h�� ���m( ���J��9�M��ii�7�@*Ү6!?i�9��I�D̂��E#�6�*`1��T+d�Y���<ͧ�?����?���?�F�)&�]��߶ol��
���ʦ{��L���	П�$?��I�M�"�@��/������3D2�`�O��$�O\�%�b>u���(K�A�b뇻.������:[&�B�5?���}�>�d	�����E*	qDt`ta�;>��4�Eʗ7]v�$�O,���O&�4�l�]�6��./��Y�D�$R���(mBb���i)=l�p�6����OD�lھ�MC�i�\)0�P5�Z�㧌*G��=�3.��Z�敟��7#�W������x��tE�
�t 2�� l��
�4OV���On�$�O����O��?�#��<���9�i��>r`���������ڟ<j�4^Ũy@/O��la�	#`�b=R!�)F�|0teԸH�N<����?�'_�,�rߴ���0}����'J*A�a+w��x�jAx�.��?��8��<ͧ�?i���?�D�K�_lF�oڣ!~|�CuQ6�?����D�������dy��'��ӥL6�P��5T$�}˃��!()��d�����\�	@�)�W�� WZPXQ�Y.R�(�	���z�r�C0�����ġGǟ4KW�|2C]N����5� #Y�I`s#����'�"�'���\����4`�ҥZ�#��Fw^Pb�]��5����?a������z}��'!��F�F*Ϧ=XK��%<V�q�'@���Ŀi���Y�l���Od�_�|��C�5Ґ%DM�#;�<̓��d�O����O��d�Of�ĩ|:��ev�TWiNV$�Ҥ{��-T5
�����%?u�I?�M�;F�舚�L*?.���#[�tБ`���?�J>�|z���&�M��'����+�=u�, ��Jױ_n���'��R��Bß4�U�|�[��S��|#�O�ZZE��,8�n�j l���8�Iܟ��	ayB�|�"4pd�O�d�OH�*���n ɺ5�Y�r�v���%�	)����O�d9��ͅY+����	H`���©X��2C����@�S�b>����'���	�'pzlj0&A-:���v���;�D�������ߟ��	T�OM=x_z���4[��ɹ�H�4}*�m���u��O��GܦU�?ͻF,�Z��
]
p�q���)-����?�ڴ��vc�p枟Ш��đG�4�7� �p�5FڷJ�n}1ǅ��H@��Z�)�$�<�'�?���?i���?y �L&C�D����F��t$U+��$����``O���I��'?���*9UrMy�L�x�NK1@�%�`�*+O��d�O��O�O�VB�Y�G�@����ØzJ\cs��6�y��_��)��(��[m�gy��3�t�B���; d��"�Z�*�r�'���'�O��I�?A����,�Vl�;D�6Ha·c7�8+-����ܴ��'�˓�?1�4AЛ�ŧh��{�l�*��`��fޭ"q:U ��i�I�y��cQ�O�q���.�>��ш��_]=��c��,��O��D�O*���O��;�S�vNtx��ʔ�tp���D ʡ�i�'2��yӾ5���?���4��5;t�ɦLޓu�f�Bsd�x{�1��|R�'y��O7�(Y�i��ɛ��\�b%�$�H��EgT1O�x���/\�D~�Sy�O�R�'W����c��!��?F�J�A	;R�'2�7�M�%臱�?����?�,�$3p��{�BJA1"05�4��@b�O��D�OT�O�142��Tֿ7�p�H��A:H�C#&ȿ~-8�z�-?ͧw�P�����Y�*91�-�mĮX�v��8>|�����?����?1�S�'���Q:�&f�ƌ�P��M(ر�e��!Vnh��؟<aܴ��'P6�A����V�[Aˋ2bN�Ԋf����6-����ƝƦ�'TY���?���F1�!����5�ƌ ,�����0O@ʓ�?q���?����?����	�Ȱ���!V�aU��:v�Po�?�����˟���Q�s������{FFך%�����ƅ?5���S ޡwg����O�O1�ZY1'�eӮ�	�
V(\���Ʒ!¡0ĉ�
����ul C��'��'��'���'nD��rK0{'�M��B��@ZS�'��'�2Y��@�4($�����?I�����#����i1 ���R�$J��k�>����?H>1�
�E��B��#Q����jK~B�F�5ٶ��7�U��Oδ���
>����[��H��(�Z���C��E�B�'���'�S��ST�ќC? X����>F6q� ���̸�4# h1�+O�unZN�ӼÅǟ"$�)��q����A��<!���?Q��i6����in�I�t�5�P�O�|lDoէ+�8$ �E��|�4̊f�Fy�O���'["�'�2'ʆYBTP�!D��h����)��^�	�MC������$�O��?)R��J��ʎ
(�|��@����Ц�a���Şg�H���� E���(���!���  ��t�rM.O��K��A��?�5e1�D�<Q�b�'NX�Kդ!Ф	h])J�d�O��D�O�4���$��v ��%N�.��t���ʌv�2ŋpGñol�l�6� ��O�ln�=�?��4x�}�G-�Ƥ����<�@���J�M+�OL�B#���Q�)����Dq�E�M�t�T8�Q߀�Z��3O��D�O����O���O
�?�B*��b��,	u��+��!�$IE���	П���4P���'�?�b�i��'�Ơ�A�.��<punݐb:�)�5(,��X���޴�z4Bˌ�M�'rh��p[Ƀ,/gj!�4��蜵�%	������|BY������,�	��P��lQi䞈۶^nV�I�!������py��m��J�h�O��$�O �'8h}��Z�S� ���N-`.���'����?����S���	I��]d��%��%o'y���A�x�|�8�O�)���?�q�$��c�3���*���BӺ_�n�D�O��d�Ot��<F�i΢�Ղȁv+��� 	�����Ð1_/��'�6-?�������O|űC`�ަUc�@���E@ ��O���E"�6??��@��c���)$�/J%t}tq�
��)�:�{3G��y�W�H�	۟��	ٟ��I㟼�O.T�� L��;� ���ղ�!�:2����;��'"����'6=�52���J����a�#~7�B6��O��D0���	vA�7mv����n�z�0�� ���5���f�t���W�#��Ic��Oy�OgRʁ�W�Db5bI3}|Q��E�@���'8"�'B�	=�M�É�>�?	��?�!��A���J����b��b"����'S���?I����+p.X��Β4��q��k�Ф�'jH�#ΰ!�0�ɏ�T%���g�'��h�l�6"��{ ����;R�'���'���'��>��	��-��(����āS��|�����M�iL��?���;��4�&�3GT�H=�%����]��b�3O����O�Uo�n�*0oZH~B�Z�{�F��S�8I���7���;�z9!&B�u�Za��|V�������֟���ܟ웅"ϪT�`9��H��6���rqH�pyB�h�DkD.�O����O����B�/��8�bH߂,�� ���?8h�':R�'��O1���M�?�B�&�Ӯ���rK� n�D@�#��D9��: ��GH�{yB�
�WC��9�Bĝ6�A$\(uR�'2�'��Oe�I�M�q�:�?!qF��Z���� )u|�����?aдi��O&h�'J�'!�㞧
��#�%�I_�d�	@���x�i��I' m����O�q�x��H�Q�=sBK�d��a�GfĘ���OZ���O8���O��$*�3c�|h	W�	�L��Y*���&Ae�=�	֟0����?�&#z>e���M�N>��$�{�pI�7���0/��AX3jL�'AZ6��Ʀ�S~�qn�z~��I� �(�"m
-~�lbUK,ά�BV��#�?q��(��<�'�?����?�F)ɒ-+ #r0VtvMٲ�*�?)����$���C�A�Yy�'Y�ӣ	C�`U��5�N���DN� |�	/�M{�i\O��F���dF��K�]�!ŏ1o�Jei�f���$�4a6?ͧ����,��K�*�Y��[:MA�'�8�
�����?���?��Ş����eI*�+X~�e�_hh���=Π��g	ky��y���XҮO�oډ�zqI�	.o�H!A�"ez��4*K��cK%6�֒�DYB�],e��~�pk !-���UJK�Y
�0�Œ�<*Od���O����O����OR˧_-pX��M�,���U�6���׷i����'��'��O�2�a��W,I���Ǿ���B�M�mOx�m��M���x��I�R	��1O�	 �Þr�p���o�S�`�1�3O6�2
�.�?��)6�$�<�'�?�$�E,u����t��x�`�a����?)��?�������ћ��]��|�I�IU#�j�t�dhP
R�(:�`VR��r�O���OB�&�ĺ�G�.m���r�'���9S�>?���E&!|Hq�i̧#v���)�?�FE�YnL��N P�� ��Ï��?	���?����?�����O��z��#�f�Eƙ�*�|��C�O.�mڛ��4��ϟݴ���yG*J�/��xr���+�l�f@��yB�'��fӨMˀex��|4�a��h���}A�L9qH �%�
X��zc������4�����O6���OD���9�\9HCiVsY❻��5,&
˓|)�V�ޞT�B�'�R���'�r	#q@Z�.�>�ҬӌUIpٙ�˵>)���?	��x��d����XȺv錢���̎P�]�́#�����3 J�Od�L>(O������>�n%�tDO�o��L����OZ�d�O����O�i�<y�i��rp�'@�-��1(���{��yw8�1�'8�7m3��	�����������M�4o�}����B`�HȈ93���
VR��4��D��r*�c��c�.��$�����$i��'ƫ8���"�&F��d�O����O*�$�O���$�S�$���Ss��:-kP@sc��:;�L��	����	'�M�"k��|���zM���|"/�)BXՈg��tæ%�1IW�S��O�Hoڌ�M�'D�L�cٴ���^0�ZT
b!�!� ����]\�R���?��( �d�<ͧ�?���?�ÌR�vT���/� �0����?����ঝC ��$��ԟ<�OG��jS!6�Ȍ�­�(3l�O��'��6�⦩�L<�O?���e��"�
(C�F�T�鰵�\u`�sb��7��4��Ģ�e�ԒObA�S�%3�T���"X������K�O��$�O���O1� ˓} �V$A*Z��qq%� ���;�@Ni�=�%�'sb.}����O�,o�,Yb0IV�#mNjM���� #�d���4$ț��\�f?�V��0A�
Q�mF���~r�IP9���!R,åz���A���<�+O����O*���O��$�Of˧��R0���]Ere�ǔq9J"�i����'���'�O��Ob��׃;��P�C���TC�Mw�� ���D�O�'�b>U�
ϦE�|y�1@s�ؙuR����74 ��͓5w8����O"pKK>�/O�)�O���tϘI��3�AˮX��lB�)�O����O��Ġ<ie�i�Zʐ�'��'D .�>c�8闤�2C�"x����A}�'�Ҕ|�㉵�\����|e�U:�.ۿ��d^3}� -�GP�z1�)���p��,F`
h����s�(4S���G�Ot���OV���O �}R����a)S�!#?�T��֑z�٩����fC�j���'&.7�%�i��맏��ti	�L��Q|z ������4#��-t�f��F�r�h�o������ܑ�p�ߐ��ԠA�0u]2�p�HѰ����4�4���O����Oz����B��rf�o��I��  3�ʓ<c���Q�B�'-r��T�'���r���5%�p�`}i��<���Mc'�|J~*����Goj�Q�̐�/��eJ�
B&�j�&O~�;�*d�I-+�'��	$�!B(T�%P�y���%?A8Y�	柼��џ��i>��'��d��Ns�덥m�ِ�F��F�����N���yr-r��⟖ay2�'��&�m���qb��#j1�8�'�OqXUhdl��
y�6-,?IU!��<{��	8�S�ߝH�����2`S�C�TY�es�,��ޟ���џ��I֟���Fރr)�D�U�z�~�2FLP��?���?�ջiC!S��pܴ��j*�� ��O�zG,�.���醒x��'^�ON��־i���5����	)��
�ύ;?>��'$P� ��i��|y�O�2�'�"�O#a�����M��2�`@Q�	�)b�'��I4�M;���0�?���?�,��0�
�<$B�*Q�1���O0�d�O��O��'�rm��͈�<�LA���_�l���q�)W�f-~$���>?ͧw�P������,��գD$FI���;;i�hq��?���?Q�Ş���JЦU�5K��b���`��vϠ!i��I�02v���ߟ���4��'<���?��˩�x�y"��(Hc���v�HH��ȟd������'!�a�e\�?��:�"�c/q8�PZ�)>5���G1O:��?���?���?)���򉀼l�`5�.��X�6Q�T,F&vf��n>m��-�	����A�S柸p����%�%1�H�`�;:F���E�?Q���S�'	i$
�4�y
� JT����\V}ԭ_>lW�4"�3O��AgE���?�vE(��<�'�?���QԒ �F�+[����iS�?I���?�����d��ғ�U�x����g�M%ǖMRE��/oX,$8���s�p�I��M���'܉'E��P�).3��QI$��<Њ���OP��T�(L酠!��8�?����OL=��I�*y�h�a�N�0WLdY�N�O*��O��D�O£}
��!��IP�ڱ_�̵doR=��LC��"�6�Wv���'l6m(�iށ��SQ�舋��<��#��w���4���i0t�i���=�ʩt�O&0�"�I�Q��`��I��Ѹ��Ty��KyB�'��'��'��ӳ
��PSH[�;��M�S�HI���2�M;P��?����?1L~��N�ڭ�S�ۺ�9'���L ��TY�\�޴�"�x���*�lm �J��Q1�A���>1�̘P��J��	3ds���'(�&��'sz%�.ݗ.�2X�pǛ[;����'�R�'Ib���]�p�4W$؁��SQu�C�^�٢�v�Ǭl�͓5Û���uyR�'��jj��F2�0r��Ȃ|���#�B�f5�6+?&B�M >��'���0AO���8��I�4�{t�c�$�	̟ �I����ݟ��R5(O *�\#hJ�\��hZa���?���?�7�i��;�Z�l�ܴ��b��A�Jրr�Tx��]�'ЈbF�|��'%��O_4��i�I0K~ � �NL
pVI�D+L�($�_ �"��D��Oy�Od��'"�� 'V2H#q���$u����3g��'N�ɀ�M����?i���?)*���a�<��H�Bf�,1JFY[���D)�OFPoڿ�M3'�xʟ�X�5�*6x���T;R@�ip����Qb�X�GN�i>�Y�'���&��� Iêqad��r��1;��4�'AV蟨�Iɟ�	�b>�'��6�X�����.]6 =,�0E\&(����`)�O����䦭�?�TX�|�4Q}�8J�ȝ_J����Z�_�Č��im7-_�^ 7�'?I�H�PZ�	8�$!B<tC�!a��2���	A��yrT�H���L�	ޟL�I�p�O+�l�u!I-,)ꍡ5D�6�l�g�n)��e�O��$�OD����D�Ԧ�]?C�	�BC�Q�r�`Af*$s�u9�4QW�I4��q��7Ms����U�f���W���� w�@P�f�#"ɏM�	my�O,�GI8�x��D�(?<a�Ff?��'���'��	8�M+6n���d�OBm91�V/j4ܩx�&.�|�� B5�I����惡Y�4l��'9v��ק�'|�a�W�x����O�#���c�j�����?�O�uؠ�Ö`h8���!u=�"T��OB���O����O��}���E����_A��!&��acl�������.-pR �s��OP��R���?�;w;����QN�@\Y�Y|ʌΓ*o��/u��m�k@En�O~���  ����'7�ZAv � �8�0���5S��|rZ��џ,��������0�T�C�W��VO_0sP���Q"�\y2rӢ���-�O��$�OJ����S�0'�M��c��-�:e�c-�.���'{7�֦5I<�|��eΐ2��=a�f߯g�D�N]�_��9)��G~"-��\��m�	���'���$U��� �b �5�\	ز��|��L�IП��Пp�i>�'6�TY\"���' ��ȩ���:7���«��R����L٦��?�#W���	����ܴ}z��[&�_0n���I�%O`T�%�?�M+�O�<aT���B����@*B������"w�y��o�,`u�5/L8r��qҗÝ|�n�a��W�BǪT�v�,k-��agm�8HVՋ�*G.^��h��˖<c�4%�5�ɲKd!�5K�8#� �G�D����%Yx�	ɣHR��u�6�֧llJ]�@	��2�Ř1�S��6�j�%Ҋ�hL�"JW��d�Y��ѭxD���Ŀά��"�K ![ٸ��Z]n�ڃ���&��T��d��m�m �f�#$2ˣ�N.=c~9xf�Nu>a���*
��$��a68�(K�1d��@b����)�	֟��^���'\�S͟���xƴ�r��Әe;0`ߜS@�p�󄊨J.�'>m�	Ɵ��ɖXj�(6��Щ��>�l��6!�{y������<I����cy69��ȴZ���K�g&x�@��c]�`դ��@����?a��?���?gJ�'w2<D $���x��3�fS�vy����?(O���=���O��d��m�³��5�8�C�B�@��� R�C������������џ`�m�H����_`��.�	+��H�q�'|��'̓0N��(�4_V��`����-h�c�-RW6��'}��'|�Q�TȲ&����O��u'(�Lg\�uh��:�b�ꦁ��]����D��=���[�2`����F��,
C�˦%�	D�'b���Wå~���?���~-D�A��;]y���U �:~�EB7�x"�'t�J���O���5F�x� )u��3dEe9�7�<�)ԡPa���'C��'���F�>��(���摆F,^�sg/;hV m��8�ɧ8�&��	�[���ָOwT}�(
�b�U���ͽN�PL�ٴ��A9A�i�2�'���O�.����M�_"�!��R�! ��EQU]J@nZ9wZ"<��T�'7��g��:he���S;2�.� �K{���d�O��dH=7E�d�'��X�DҸV�m��*�[8%��5�*z�D��F����wh�t�Op��'�Zc�V��*۳6X!��<��A޴�?���J+ =�Ieyb�'#ɧ5�h�>�`hXa�TBR�Jv������'w�l�O����OP���<��� �Y�d��?
�69��bϘm��	B���*���Ty��'w�'���'��iV���f�*m�᭞2=$�a�0x��F9�y��'\��'k�	x�z8��O�f�zE%�9`)B]چ�1F���ش����OʓO����OҨZg뵟�k��ۣE�@�cόIc��h%��>���?����򤃈 {��O��ۨ6�\-�Ƣ��0V �P�G.�6��O�O^���OA����O5��]�L��X�d�֘�B��;v�`S��gӨ�D�O
ʓ3]�uI`\?�I���S�bDɘ�bl��J�O�R�&� J<����?���U;��'2����:��2L�p��X ��%j+�VR�$"��Z��MC���?����j P��X7f�d%9�`�8.:!�7a�i 7�O��3�"�<�}��$��d�4̲5jG�H�ڸ����ߦE���0�Ms���?����B0[���'H�Ђˑ�2��)w�o�����<(���O0�������W��|J2�[!y���b�F�W��iub�'_2��
q]:���D�O��ɼkܰ�{��A	od��N1_c�|R�KV��ן��Iޟt��"%��� /�3H����j���MK��7zFa:0Y�|�'�BR�x�i�-��%Z&Y&����E�м�F-�>�dK��䓭?����?�-O�$1�m]oT�,�AN�0���W�����%���	ӟ $����u'A��oB�|ʷϝ#5�d](�L���M����O���Of˓���b1�԰a�S������~� c�Z�h�����$�l���$�'A Y.m~�(Q�M����j4E����	ɟ���@�'=Z�`��?�I?��qSvg�3�t3����K��m��@$�D�����'��%��%��S`5�a��iY�oZݟp�	`y"��c�����D�k�]�8�u�V�I��2 ���mƉ'�I��t�I~�s�֝�)�@ݒ�mQ6:pk��ĭsJ��?B
�?��?����(O�.ӥp�Ib�� 3n\�p�?!��'M�I4w? "<%>Q�����r�0K ���`�~b��O�D�O������S���^���$�@lU�P;�ۍ_� �^���Dx��	��H6�eXF�<�DYG��eIڽo����럜Iw		{yʟL�'-��� � `�Z���XpV*x� �1Pᱟ:�䲟@h��X6!��P���۪0i�E!��xӦ��3$ِ˓���o��$İ�&� ?,�P����E�xR�ƍҘ'��T���I�%��X��Q>3�F(��d��wXhxG��ey�'���D�O��I�l�J��4h��$���;>O7M��
m�I��	ǟ�'�Z��sJp>K�>���X�5�ܬ�'mȓqs��֟��I|��Vy�O���#!�n�7��<�H��LD}���?���?/O6QʕC�i�S�[	t�i�5���{�A�?�F��4�?������ON�'�?�J?!(�+�Y�v`j����L �\��j��d�<	�M��-���$�O���(Z�!WC��� ���m� t���x�'�B� �H���y��(��$M@�\pk�A8Sz�K�i���%$F��ڴA�ʟ<�S���Jt�1H��!���C��N��VY��b������O|�I~n�=M�P�ǏH<j,����0zH�6M�,d���$�Ol���OT�I�<�O�$P�ǜ�f0�ӁCV��L# d�5ɂa�9�1O?A1珖&+��2�A�\
�������Ms���D��h/j�S�4�>!פT�L���d��t��Uz��ɩ�1O��{)V�Sʟ������*!�i D��%��X�����H�+�Ms��d
"`� �x�O�R�|�fe���b!*�1,(�
ĥ� |9��V�a�����?�*Op���\\}.
�Ճ��\j	�e��.������e��?����@)`�c�$`/p��E&��6z�A�4-�	���'W��'+�?�i�|� ��?u��0� ʔ%htu�@l��]�'1�Z�X������	��u�|�V��.ꀀp��Q�#�R�*2����M�s�n���?Y*O���%�Q�4��5I��;t�Yc���z�CPʟ��M�����d�O>�D�O*�:';O�����@p3�6\��`!d�7 �H�"�j�l�D�O�ʓXe,���W?-���$�Ӡ?jn��tHH	M/~�+��4�ڑ�OH�d�O��%M0�<a�͈�������Oq0�i'?�|�ـ����M�.Oz8��Ʀ����t�I�?a٨O���H�*�R��o�p�`�5���'B򪞘�y��'��	wܧY��8�$C+i�R�5D�?M	P4nګ��Hs�4�?���?��'���Zyb�.x�$�0sc�-�ڥ�Э/��6�8z\�1��8�����d��o���"�ʳ`�䡂d��M���?q��h��5_�ܖ'x�O�A�!�N�`�n�����w�4��\� �'Ŕ���O���O����Ot���-!�Щ�Ɗ�+�H��Q�릑��."�޸*�O���?�-O���Ɛ��f�H�5�VU#����#f>�R T� ��x�����I˟���Py�M[/}R�y{��_16��YS/�C�J�اj�>�-O��$�<���?���q}@40qFg^��!�_"SG��Y "�<1���?�됡�?9����$�@�ƍ�'k�99���RڰM�w�U( �"$lsy��'��I��	�L�mp�8sB�)�F\�%��R`��h���0�M3��?Y��?.O���ςi���'�� N,3�KH�2"��Ȱo�6a��أ�i'bW��I����	�k���Iq�dJ�8��ըT��r׀ !���0q��F�'�B^��T�O&����O��d����z�m�_m qkf˵~��EO�i}�'Y��'��58�'��	�>G��':���굀Y� 0Z�
u̟2e�inXy� �)cB�7��O����O��I�r}ZwF�1�G�i�j�n�i d�hߴ�?)��>@͓�?y.On�>u8
�	S��!��ڢ>(�@��|�`Q������ǟ8�I�?Y��O,�L�@�v)�Dq*$jH�KUp�0��i ���O,���O?r���Q��N�|�,	��N@��l7-�O���:�FA�ej����O���f��+WF�A�Δ�b� L07�#����^o�?��	ԟ$�''IV�XƁJ854<�'�Ήn\�Ln�ʟ��N�8��$�<������Ok��).�j��J\57��CM�:���<&|������I֟���˟��'v���	5,p�0��,D*�#��	zt�O���OʒO���O��un����@��	���!U���<	���?������ Eb<�'bX^�a���@����8m��\�'��'?�'��'���%�'�x�)���Z�Jl���#32��6�>����?9���DH�l&>5A�F�Mt����(��K�����
�MK�����?A��_��͓��:Rj���Wu��؂u�P�oy�6��O`�ĺ<!�]6�OS��OBj�c3G����LA4K�Z�!��(�D�O��d)%p�$8��?�w�=,f
��cJ/�f!�׉fӬʓ6.�|��i�h꧳?���c��I�bY�㵀͕|����� &�B6�O�$�'\����8��=�Se=��K7E/Kx)"��$�.6L,Y�*�lџ�I�`�S;�ē�?��̙a���� )�O�r�!�&���lݎn|����O.�Q�O=Y�(�#! (�I�!���	�I� �I�i6d��}��'H�Ė�I`Jl�q��F��=����(�|Rb��y"Y� �� �i�5���[�xS\�@�é_`�`*�yӼ�d�43idm�>Q�����+�&�(C�D�s���qIF�n�g}��I�yZ���Iܟ��	hy�ۦ<Z`����^�.;��f	/Q��@�#j6��O��d6���O��d]2}��E閼7�|�Ӈg�BL���s
=���O��d�Ol˓]?�5y�:�zA�EN�~Y�[���"z1"��x��'T�'���'ՔQW�'m�HjĪ�5jT<5`�ЬI.��&�>���?q���к,�L&>�jE�
Fc�0C*я9�8P���S��M[�����?Q�?�ؼ�����IH��)	���q�Ұ��lާHF6-�O����<�d%K$8��O���O��顁	�6m��9�/;m�	�!I0��O���δJ��5�d�?�{�jD�J[����/�:j�>|3 "s�Z�|~U���i2맯?��'e�	8F:Y�Wϗ��L�i�$�/4 7��O��L*=�D&��0�S�u���4mA{e�h��6�ʤw�(�oZȟ@��⟐����'��i�0 \0p�a��I�J>�3UIk�Y3�1O:�O�?I�I�pj$����C��c�5YT�)rڴ�?���y��<9M�On�d����
�� `��r�	X���t�h�Z�O\�!1�Q�矼��韼&a�{P��C熣fE:�IK.�M[�'�ذ�x��'r�|Zc�xԻP�S.\\&�I�4�x�OP,qV5O���?�����Jڸ� ��ߢ-[pz��ʨ~q�10��TڱO��$!���O�����aX�2�!0}�\��R�� *T2�դ�O�˓�?)���?�.O(9{Q%��|b�/�c���02�E!,]0�jBi}"�'L��|2�'M2�&�y>\2��Po@(����!��%3L��?���?�)O���� �]� ]�5���y�TP���A�E���4�hO��dV:fv��+}�o�D�a��HN"6ġ)܊[�'`�X�x�\e|D������k��Q�8 �ά1�Z=��E�e*�O���!A���'�T?AC��b6�c�#�>d6�y�3�f��˓
WD%��i�l�'�?i�'���Kdp�d��p=�4���KO2��?�l$�?AH>�~���ޚd^1�$EB��T�Qł��y:	B����ߟL��?��	͟�O�֤B��E��p��D_�_�	��{ӂ тmJ�11O>��Iil��c&�:}4��I��-��ز�4�?����?a�?���z���']rC�+np���ݽf%��s��7y�c�0�bd=�	˟h����T�1iB�Yz��d$�,�ʜ��,\����4*b�'��Iȟ�$�Л�e��$��qj�a�:C����-58� ��\��Ο,�Iqyb+��J�ܜ�V�z�Tp�D̠P�񠤤�>/O�$�<���?�~E�83D郪S�Nxr�wG��{Ć7������I����'v���w�m>m{� 	b0������:`h�.l�ʓ�?i(O�$�O����� ,�Ĩ���Z�hW�0�7LH?e��l؟���ԟT��SyB�+���'�?	�n�6
�B�!�T$2]�l &\�V�'/�I��	ݟ��0�y��O� ��Tҵ��;B������M����?1(O�`��D���'�b�O�"  # �-(M1��OA���ŧ>!��?�\J(<�����?����^	�2���J�8n-��hiӘ˓0g^��F�i�B�'���O#n�Ӻ� hT�VGK�4	��AH(X�\0� �i�r�'�� ڞ'�]���}��E �0�3�J�(�bp���Ϧ�"a@��M���?����_�Ĕ'*(� ���cy�@	]6���baj�6HK�;O.���<�����'�`Qq♡#}�̋5�%Z�%��/g�����O��D9dv
��'}��֟X�(U� 0!��j^�t�G�rDn�ӟ��'ڈ*�����Or��?ib�$W(���)�F�� ��iuӔ��
�= ��'��I͟L�'�Zc=���K�; Pv���`ųqj�8�Oph��=O����O���O��d�<Y�B���\��U�u��d�C �-xFP���'W�]���	ϟX�I>r,��t#ؕ7�@������}�D��۟� ���Y*�NH��)�	!r�@��SJ#f���b'� oh!���#�%�#)K�C݊M���]0^IqO^d���X�'Y�H���NV�Xzf�H�����R�������To�hZWd�
�$`*!��3�r%V���Q>!���(FR(�p�Y[�����c�8���k��z�� ������ل_�9	���#t��)��7R�Œ���h�<�@E�/���G�irh��������p���#|�%�2�S�*�3��˟\�I&
��~�S��O�x��9��� ����֪4}��w���O ���,I�F~�,C�l� �q�I��I�J�O��d"�I9�	�p����S��+_��2���M�1O��(<O �	"�I����BF�&c�sR�'�"=á�-z�f_�\Z�j�%�0�����F�>�y��Dş<�I����iޅ�� y��f�çW#�A��ٓ#�{�Q��c�*��@b>�OF�k�)ޞm�2�����1J�T����� �C}r)��:0��}&��HrDJ�Mq��ٔ�ʘGgeC�Hß��'��0���|����H�b��c��h;~mz%� S0!�$� ��L{!l�7�4�����	��HO�Scyb�G�I3:0����)#6P�c�T��I+�	-zH�'���'1:�]֟ �I�|j�+Z���0�Z(S�*
�*^���@+���᱋�(r̢��	��J�x7fٳXЄy0�L�)Аa��@ց���t�Te�	ϓC֙�&G����� ��@�ֹ�e�JП��IA�'�O�����$7H`qc��1 :̜[C"OT3�0[z��jB++��(��T}2Q�h,���M���?�� ���-�D	��ːLHD�̭�?I��X*��?i�O�l�Ғ'	�5��'E��X��^� O$\�d�@��8�8�S���0s�Z�ē��h��,Qq�|ՙ0���l�XI��3Dy(���Oz��O$-`Ũ�}e�X���ɓhyj(XRƲ<����������M���9G���W\v��3Odn��C�9�ʟ�C���fBʜ(��	a�����1�Qh�l���34�%K� �"O�,{CM�:�4AB�Q�A�Й�"O|��FI_�^�X)K�J-9
�DA�"O)�'O�bX<	��K*$� P"Oz�s�F�.|�Mk��%���"O\����R+ؕR���L�|-�0"O��E�O��<�(F��$#a&�S�"O
1�VA�D����U�5"�"Ox�R�/2)�NqCS"��e5�@�C"O���,�t&2��ӊE�9�PH2t"O:)�$E�Egz���J�B�$���"Ov9T���h[��xc)�!���"Op% ��$Y� a)���m�r�"O`� �F�8� ��g,�%F�����"O��*���z�H1�)҄��%�"O�$�I�2�A���� ]~�D��"OP0���?��X
���i�-��"O�P��dŴw��9��_14���"O`M�G�X};��m� L��"OΜ�3�ċBn�(gI�G�^XJt"O�y�뎳K��SW�hx��"O�H��$T� ˂p4���`Y#"O^��0�I�'ttS��O�R6~ld"OTpҔ.�{�!
l؟%�Đ��"O^�s�,�i$���\�����"O���%H3��p'�ёj��p9�"OH�r�'d0p�&HB7i�R�X�"O�-Be��
tS&����R"O� �x�
�6
Q�}�1�\�Y�`��s"O$x*��!l��]Rd�l�`���"Oƙ+���(�|����1�P���"O�#%$�`d&�@�OJ�l�ptk�"O�m �["D4�ű���)R¾��"O�`#ҖA��ũ%�o�h��"O���!�Z�f����@���C"O�jB�H�!�HiS�h(��ˀ"OA�&�۱8��1ۺ�R�rE"O\\��/-�������^1pF"ON������&� x�`Q[���Aw"O�eB�Kx�6I�w_�T|�p"Oh��N�&�����K=�I��"O���0+N*����`k� β�Bf"OD���KVt�4H�'�ĆH�a�"OH�YH���]yԬ_	Zƹ#�"O�آŔ2;L;u\�2����Q"O��jL	�.qTmb�������"O�]��|5�1�wM��|Ɗ�)�"OP��&䖯T�@�[�n�$9��s�"O�u!E���K�F�>�� ��"O�a�!�]7�a���,�0�"O�a2�hا8WF}s��)j�X!��DL/�� G�tmM	�$:%�/W<�a��ʎ�yR�]8�|zJϘM��48���i���A�d;�g?	�ܛd��;��ϥ2�ZZEF�M�<A��/k�$��ᛜk��9`�(���vj@��0?�s�A`�U�S&�?��"��3|O�Y�c-�iy��$�:���5e>�����y2�۫lDy��4M�I�	��'� a��a3��9Q���8��Y$��	7`Y��#{����9)
}!�Ɂ&O�Hs2�ٚ��'��>�ɕNJ��`��
"��:&��f֮C�ɧ;^\�y��9�l��oD��牜S2L�����%�d�^��t����P�J�ȓ\�� H�c����Bӗa�,�ȓLx��*���1���1��������z���`y����Y�6��q�ȓP1��A�MX�h,J��r{DA`�<�Q��U$���p�*�qPt�Tg�<��c
� +�C!�L'4	��0jN�<1BK�hl��2��K�I+B�QD�<!ザzR�B�
�E1���5NA�<qD&��.��̳s�_�6X���"O�eRP�E$v��`�	ހ`b��""On�Q�+�G�F(�0 f,��"O�2���7o�%#UA׎k���X��>	ƪ����=R��@L�#g̗"ȑJb�H��� �bI�����~X�%�	�+шx!d�/D�*�n�z�,0!�P�|��#+,������I��=�[�dT�A�R3\�`�
�'�)Q#V�Wi�陑K�1v��u��'��
S��S<nz�mH%ɖ�R�,��K�B��C�IRI^�z�!A"%&��ۇ�</Vh�'B\�7�'n���2Ʌ�a�����V��yr���Ey��ʃ�7iX�,�Pb�y��԰qN,�$�]F��B�'�&�y�KTFD��)�ãPN���O?�y2L�r厌H�&�N��\S/Q2�y��� >���H��@Ƭ����y�˛�jgV�)���.�,����y���U�����D,+S�]��BT�y���7�����ܤ*b��y2hO���C���X���eV����� z���%!f��Y�2�K�Dц0�"O�ea
_�_.��R�U�"�"�Ѱ"O��{7@J�mF0��ҥR�zBM��"Of�*�lT�s�8��E@�4�6@ a"O��(	�!_�s��$@�L<+�"O�-0�+�$���j���>#(���"O<u1%�4U(�aC`>8k��s#�'xୃrV���q�\�L��v��J��H�&7D��%n�7-n`%����è�Hg6�^i��p'B,�D�^eq�G��9�Nd��a��A��i�ȓ^�����*XlH� +(zD�!gM<i0�"~Γo&�����	�([��T\��~�z��	� ��J��_�)͓hpb��>�O��*#E;�)`�i�#uG�q���'&9Ps�
����^�L�F��JZ)/���"O�	��~�]�%(��\v�� �$��]�:�0#�
��h���;��;0�,]��G�%��P"O�lr�M�9߲M9t.X����'���ߴi��A��@˧/Y�O��kt�D�L[)��R,B[�Ј��'�i㕇��7�(��͓�>e�y���Y,NT踱�͔�9\<�W.�j��Ą�,��IѤm��V�b��dG��OQ*#=����:w�I���N ��a���h|�I�x&�c�iͻv"�+d+�!�dZcꙩ�ӮUR����Z�4Ǜf�Rw}�A�1�RZ<P]i��ȔFF<�E�\cK.���e^�n�Z8@�Ԕ�����'Dl��A�P3��i�fT�B��`A��]$4��oQ�r�V�i���������'������LL(�%�5)\P�	�*ڨ�x�K&~L�:W��
N@Y36@B�@0���3��Ph���u� ����TW���WA�f��i�3Mء$��4b��C�o�����v�ћ"�@#R ��c@!x|��A)�㐃�4�y�İ<��@�r�`�h��=�M�"6��b�&�V��x����!�>�|�1C�8(�d��\�t@c�J|�t��ȓKи=�ALπL6���ࣈ�W��Y� ��]D�-���I*O���;N�e���	�ggb��ʕ�8���\�~�(���X=F�8{�>G���`�%�!"~l��Ql�;�0�oZ�Z춅:@�'��Hå#�a�^U S�F;H����z��@p�h��T����-E�!
�a�.^�0����2D�(���7�-�Xxa����=UJ"<��Z)eY �~ڷ䎩��r�S!�e���Z8��ȇ�)�I�T��	�eW�o��-[������I�A� !�qO?�ɄN��S�a�/�Ai���G6��H����>�r`тI�4k�����(fQ��	6�����p>vh�X��g�³C������ ��4�>�*<mږ�V�9L|�̟�Ė�M��I��Ɨp�ذ���C�Zv�~ң�=>6L�4l��~4k'��1vnfl���CF����W�6�za�n�֟��3�ɐ%�������K���8�e�$?qQ����"����X�'�AY�r�Q��OXY8���5{��L�h4>��CdU�ؑg��Dk�	K'�b��gc����_���,��+S�An��	=8~��Bbn��2p�e��q��O2EZd��?�P�@n�`�GO�RC���Mz���(&��|�fֳW�f�:�-�2d�>y�1b�q�f<y�d�SX�'�v8�4��Pp�ʠG�hX�	�
g�f�iG�'�ڐGMЩi�he8Ma1��bg	��F6�̓��`Q�}̓3QtA�6�ij�i�)rhd2We�;j� )́�p�^����d�'�&��P�2A�
��
n,A0�$v�d�N�#Dt&�c^V���BP��s��6J����&B��Q���'@�O��S/�-y��jw�ؐnfҍS1X���3�E�F�u1�f��Vrͫ�&?�`*�uC,�U���:�ܢ��L�BUUG�::ti�բ�*h`ː#$|O�����-r��/\��8q˸l�������Byb��1�21��jKܨ���%�*E���R��?[�m1"�P���?)�-�
\�ȡ̤u�X�K�kذ������<�@L[����T����n4�Ԥ�1dH�H�x�� V. V*p��H�W�h!�� ,��E�i��cm^Lp���{ �58���J��I#����7�ڠ���T�Fhg�i���ZTxZ�؅��8b-T�B(M����?a7��s�L�PB�=�\щ��RV����r&�����]�R���Q�L, �Eo؜/�0j� O��ԊC�@/4���vh�f�(��'�&�d�;���)�� E/�=�I>)�����e
� �� ��ƚ|?9䈯�2�oW�}&Y�%n2���)f�p(<�7+ � j���놺��܊� ߵl_8�" ���/w��W�՝x��\��]�|�q����!i��|�m=h܈���G�xsp0���p<a��ic�c��Ɇ+T:X$0b�Ă7'���%?a�̙5e�N]	4%�uYp��F�d�'��h�h�,�((�k��+�Y�O<���O_1OuST��2��=r2�DkC�ʫHS� �aH�6ufB䉢:��d �Lܾ3�G˄�o~㞌�aJ�W�S�!���"Zؖ��C/�� �C�ɼT��mZ���-%�v�J1�ܖ% B��* �L4��h�5���)H.bY�C�I%�U;�C�06�BЀ���`��C䉐BF�=5� pR q`"�B�ɭwn.�9��C�� �&��3:�C�Xrha&�P�@ָ�q�E��1�^C䉎7UF$٠��Nmܽ�TE:m"C�	�᪐�vO�G1�q���ڻ}�XC�I-,�D����P=x����F�c`.C�	"� dY���QxD%�E;�*C�	0H�,BTf�XN J ���C�	�
 ��`�,�L���N��22B�ɡt�c��� .J���-�&��B�&gtZ#cܾj�\ug._% ��B�	d��E� )�|-8v�����C䉓.�6a��ĒNS>�Ғ�]�`�C�ɥY|1��]�t��8�V�A;XNB�I&=24;��)S&�@��΀�D��B�#8 �cT�V�=���kp�@#D4\C��2@�r`�' �}Á�u��B�I&XS�41"��t̊&�"UTC�IdǒX��̖���r'�(C�- �Zt��Zx�I�(�o�0C�I�1`"̓�*1s���!0Y�Y�BC�	�e��xc��5{�б�C�0C�ɣq F�`rJ�\��A����X�B�ɬ�&t[vM�i�d�)�*r�JB�I	x|���0&X�[$�_>:B�1M�^T���;b<	�BG�DP*B�	l"z����{T�!Y����C�ɡ1�H�ÌV[��Q��K=-�C�ɐQ���1'��7�\����Rr�C�	�u��H'J5f�X�S�s��B�!������1޵	��]�w�C�Ɇd�L-���I�T��-��*.I�C䉷mFi{���Cа���G��r¤C�		�0죓G��;�����Ƅ8LzC�	'gj!���I�,�ՉֲN�VC�ɧL$U��f��;�d�BW��O��C��^�(�ٶ^q,�a���KT�C�/O�L��6�R�lD����N[�<��C�	�����dI؃p?J�)�
 ��B�>���;`�'P��Z�,��L�B�I��8�Ɂ������F�p=�B�	���B��ؐQ��-��$���2C�	'v�1	��Ej<��B�n� K�.C�	�mͨ ��<P��ũBJ ��B�ɥ^R.Y�+O�>���"�#�_^4C�I
.t�T�/U6�]j`�O�X��B�	w�v4獄�a�@�#a"-a��B�0:F�a�D�L
H�Tq84B�I��B�A�Q�Ū|q۵�6O��B�ɞ2�TX9e��J������fB�ɿn��Y���^����%왠9?�B��0'�E���86���X��Բ+�C䉐SK.���ѴY����Bo@*\zC�	#a���Y���펰#0i��F�pC�)� �㣌��|����ͩ

���"O*�V!UjG���r�?O�B�"d"OD��7��)C\��`蛃l�*살"O�X{%]�ȱ iT0R��p"O�H�"-�n&��Ӂ�'a��"�"O�� ��i9(}���N�y�Z"O:�����F�YCo͍4h�4�V"Om��n
��6���&9DiB�"OΠ��k��U�r8�@�9B/!(�"O�h�f��0�,��x9 *e"Oh�ʴ8	^T���� Q�&m�&"O�`cED�j�*�m�<���A�iH<!EG�G��0��1P>�����<ya�]E0�E33
C�I��,R��Hy�<�����C,�u�h|4H�(�jQZ�<��a��JNpk��c��Au΋V�<�V��W���7�_c� aѐ��S�<1*�{����zF]�� T�<���,]�B���K<czx!PO�Q�<�2�ؖ \2؀s��*���(NX�<�e�8}Y�~�pb��S�<�5˒�w����$��9Q�E
+H�<����� �Fɐ�d�d��`I'cC�<7cW�/�qڒ.UyZ���}�<9��PRC�"L�X+����!z�<YF�I�u�r�e�n�2 �� �s�<�1l�Z�i�k��f�T� F
�u�<A�%�,wꆀ���ތ�fՀ7fHt�<�d��9@	*$
�p�,��"H�K�<yp$A�1*�ys%���@F�<v�t�MT�W�oi&ؐ�/�\�<i%j_L�X,`���(_Gx��$��U�<ٰm\�j�F���ʈv4x���J�<c�&N���a�ɉb!��Q��H�<��΀3>�N8���RUR5T|�<qC-A7-8r�r``C̒5N�,��B��{bn�S��B�.=<�YBi�$~�B��9$j1(�%L�k�`�4y�B�	�	�D!j�e 
�4��"N�y�~B�I	k��Rу�+*!����P�2C䉗%h��pc�^	d t�̍�:QC�	\	Sd�����Nn��s�H0D�$�Q
�1~�K2 �.��ū�#-D�Љ���?@�����O,\���?D��Qt��x�L;�gT��`Ix��!D��ʓ��-�t�+A"��]���A��!D�`3,�<���ªE#G2�}I�?D���A�	��0���Aֈؕ�<D��KD���h�횈n9���5J D���Հ{U``׉��O�����L0D�,���F�Z�n�I���0>�$�*D��֧��ivep���0Y�P3�a'D� q�/��!RQ.W=O�l��&D�8���-L��1�R��x�#D�t�B��3[�HԱaE pOZ�;�%!D�PW��%�n��g,Ű.A��h4D���fR�!�de�����2D��K�G�m&؊��ͿS��%1D�P g���p��bֆV|���9D����Iìal�$��6�̥*T#7D��Gƚ�	��1V"I�Ρza�'D�p�+ǈ1 �R!�6+�b�h�h*D� 1!��W�R}:���+.b$be)D�dq	^�c֔X*���"0��Y�o%D�� ܸ�я^�̅�&,�n`,
"OB5゠�'H,��-{T�<�0"OX��6a��*���&/Ծz�f�Ȑ"O,��&9�YAH�3C��p*�"O�����d��pF�0X�{�"O�D���w��i�Kǿ[.z�!�"OR�a���V<h����.p�|���"O,R���Y��T�D�]2$�$@T"OD|��(x{(-��Z�R�L9���`�Рv���
�����3o+���B�.D��ǒoD֘r�ֿ=b^�AG�,D���#Y4RBB���!&RD�CN)D��"���hQ�PcQ��^��@e�&D�\⣊��x�@d*��\�
!,:q'#D��ؖl��D�����:��}��)!D�h0��[+q��u��$>��=��"D��!��6��i ���v��8��5D��86�׸H,H��e�
%�i�14D��i��
�7yqI#�I�zAZIt"2D�p��/o����q�F!/�pY0B(/D�Lx#᎛2�&�8u��&5f�µ� D��@�.�Lb��iwa��_�1��>D�\A�@�7Cv�Je�P(9�!�h?D����!���t9�� J�Ryö�8D�|j��R4L�tP��N�T�,j (4D��A���v�y��a@4q,II�D0D�조s$`�_0vQ�9D���g�/q��@��*qJDH�g+D�b���-Wfmr��ؾH^8p��'D��z�̓�Z�b-�dY�1$�i��"D�h��8v�D�VM܌>��5�s�"D���C[?$���ɛ,$f�0��L5D�l�)�F|��"i�-_����B1D��@	!WQ䀊���4^���[sn:D�̚�+2	&4p҇�=]}�UBa�=D�d��ø�=���E�<�9�,=D��n�\f���C69V ����(D�0��jį:�B�ې�J)��с&<D��0���iE@4ʊ$/�3am:D��jW�"c����'�|��	;�e�s�<���{!�x���6'`��S`�Z�<1��/��#�.ش*'&�����l�<�uIEO��t*�ă-
b���K�^�<)��@zZ=x����y�(`2��[�<�AQ%$H���-�QqHɶ'R�<�¦���4i�`"��|��@!j�d�<it�ӣ��q`1�������d�<)���u򔄸���f�h�
 G�b~��'0�u����q\��a!ʟ�D1ΐ�'�X�
��Cf<q���X�C0(��'2�ԹNP�M~��zq�Ŷ7���Hӓ��'��M� @?�[Y��G -S��'�} �gI��$�(�n$	6}[�'�<��&�#A�J���2�4r�'����c8\�R�0��=l����'tݫ&Ȃ�+E�\J�ϐ��,�	�'x�Eð�7{���F�΢==|8��'߈�:�m۶OTLr6�?�ht��'�:(c�O�j�P�cψ6`ġ��'��<C���9p'H��N�6(�X��'��Aӂ�&(p���X1Qܴ��'Dr� �C:\�L���"d�	J	�'��!R'!�@O��O'�D��'*����� ��q�hO�2����� 2zB�P*LX�KVu'ʽ�"O�DcMó�����P�"x��"O����[67���.֦~����"O�yq r���dg
�e	��)�'�`a�4aC'XVu)6O-}�x��'�x�ؒ�P8]4ţ�#{'�l��'v��RFϑc�R��q�I'kl|ٲ�']�pRp�[�&���!1`Pm@�'N� y1�����w(����X�<%n �"@R5 Ղ1K�yQ׏Q�<!���&HԃU�� Cir=�c�WL�<駅řN,� 5�S�^�H�EJ�<�U�Z$z��	��Yz�j2��Ї����@�9'�,�10��-ɮ$��vӖ�a�Î�@(yIg&W,L�.��;�p�@b��]��U�q/��f����g(lL�d�ӵmU�����yF���ȓV� �*BFP6@	b`���3(f�$����q7���2��zf��8ZQ<��{�>8Q���'���*@Jҵgi
5�ȓcA�JmI�	fVE"-R�	��Їȓ]�N�r�-Y��|��SM�.H¢Y�ȓN_����C�"�������2�5��X��R7l��(\K���A�Ȇ�}�(�� ҤK̠(`�D.Q=����^���g����KT�)&�	��wC@�гG��Q,*���L/z�\��w�r���1P;(Q�&dE��>�ȓ��æ��$-#4�Ә4�"e�ȓq��%�7�TZ�8�ޘ3G1��S~�B`�Uњ���E+@�p�ȓk;�YJtO?x� 0�B$GW`����o������,t%��b*�lF���ȓ"�Lr`J�f������GY*�ЇȓI(�c�<!|&����Y)}�BY�ȓF|�<sG�ڞU"�%�G�J+�n؇ȓ��)��HҜu�<u��b\15Z �ȓ&b����]3�9y�C�+,��ȓT%�j@t��$k f|t��>P����"�Xw�A�9Tцȓk X�FJH�O��a�vL��, �ȓRl�)������I��D�;
���+B&�S����/h���2�Ab~��*G�m�o6�D��N��̄ȓE�ḇ�Z�� �T��Y���v��U�ε<�F��Ɣ7⊍��;�<#�oZ�8��ħN�Zd���ȓT�*�;�O���D��	��(�4��m?2T�QbC�t���j�EA�F�i�ȓV�`� �C�`��Z��V�@��ȓi1� �KX+d2!�͆O��E�ȓ0����e��t���&SOm�M��)�PP0I��r����f,NZb݇�VW0 *�$
��F%����"9�l���O�*���)U�q�<UX�u�"O�y���1�\���+�\zP"O�Z�KV\�H��
:�t��"O.��,ؒ6 ЁW�f�f��"Or�[�#A~Z�8q�D�K���E"OZA�0�ڡy�>��c'+�2  "O�D�*�'_��Y�$'Pf�
�X�"O���C�H?7�
�S�K�p�R=ie"OH�IAHJ�'VXIE�C(f� s$"OZQ�r!ːI��������g��l$"O� �����7o��4fсZkB���"O�YS%^�e�����A�|�P {7"O��3��9�:�� +AL@I8$"O��K+	dh)�g%5MA���"O�3����J����n;��6"O0�S'�S2ND2|2%N�	2�d�"OZ�!�Qj(�PD�,t�h �"O�)���4�����aK!`[l=s "O"�	���jx��%\ FER@��"O���2��,m��X9�%�"h����"O|̃���*�vEJ��J	�"O�9����q�&f���L�!"O.�a��Z�����Tŕ-Y���#"O"I����I<I�V ����!"O���,ԂJ� @[ScN�i{Z%ȁ"O�-��B�o 4a���ԗu>�0�"O�����lM\���G�Ne�dW"O�����9'j�!�F9PXv�ʗ"O~�B�Nۜ-��Չ�=W��"O�\['�FȄ����P�kQ����"O(�0�D�q���te�(���yv"Oxm�Gϒu�T�eD�`�V9�R"O�t��U��%�^�,��r�g 	�y�M[�@��l�iă��@��y��Y7İ[R��7A� �	���y��1N�� 0��<'.�)��̳�yB��QR����c�.!V]�����y�g��h�z� �G��H��g>�y��$O��Yavb�9?0J�x2OQ��y��Ѓ0?Ȑ���*>G�qq�y��LZz�)k!ϔ52�B%����y�mW�����b�+�����		�y���c?���M6%��Ű���yBI�{��<�QǏ�?zy���y�UGz�����a'� 1�!�y­�8eq��q��Ѷ�W;�y�"[W�Y��jN�xjì*�y�Af����R�r�b���1�y�eXE�D1qN�Pb��K� ���y�#��9�Z<B�	�G�4���6�yҢF�_�eIу�R�h����y��	s�z��`�B
R�LH:��9�y���#ul4�ehK"[�!�'�E��yRBU�u��Q��X�_x���
��y�<�(��e�7\���[�EZ��yB��\ʱ�o+Wf���A�y"�ĖU��\��c�(Q��#&�^��y��2u+$��#"9�B�Ő��yr�)C�!��$���!��yBK[�'$Qr�hԖy�ε��ԧ�y�àG^)���U2y�P�xd�@��y�BS�b���*� ݛl��(�L�yb�C����$�5i�Rq��j��y�L.��Њ�f�eR�@� ��y�a�nN� "h@�?��D���yB�5�n-��E��.R ��V>�y"�S:sZ�������RU�<� �D�y�ZRbF%�IޮG��qQ �J��y���f�`�Ĉ��k�QB����y�
Ǥ7�m�t�G�:��g��:�y'�J����TJ��5h����y��ʶ2�X���jF��>�i����y��N�B��+�~,��٣OG$�y���H2Ptx'�Y5s��-���W��y
� 68b�G TBf�H1�bo�U�"O2��1�Ε\Z����Q��0�"O���l�,`�,��V�L�	V$��"Ofq;�"�&b��(鷅�8���Ѵ"OD��fIN5@�)�M!��<�"Oduz�<�����"ׅ��0	�"O@�@��G
���� �X�@�����"O���g��:�J�Jp@U6����"O�q�IV�p�:�Y�n��JN���q"OX��IA^W�`���R��I4"O4����ʃLK��S�!�r�iW"O�{�B�h��t�8�	��"O�cB�	�}�٢�c_%e��ำ"O�I��l��t�H�B]�$���"O����/P�R�0 s0B_����"O~�sH��x�8�jg�Wp`ȡ�"O�a*2΋%�����_k�ĉ�"O���a�E�jτ���Y��=��"O�}���
ixQxQ��W.���"O���a߻=ߒ�IsKB�I�|�r"OJX@��<�P����E��m"O���qI�:s'.�I[�D��"O�m��B��#U�Qȁ�. ���"O��H�%G�W[Ā�'D�c�dA�"OjE"ŞR39J$�ڡB����D"O�U@��֊0(HK5��	U
I8V"O^MH���$f�t���W�Vnh�x$"O�a��E�ȪР�@��Y3�"O�=J��A3_:ZA	`͐n��0��"O>py�M�9L�U��k����4"Ov�aB�O��R}��D1Z�+�"O��Дkި:�e@�����$m��"O,dc�NLS�|�c)Y;�@��D"OH��AGW�2�R�G��F�(�"O�A�'��&�@d'�6^���"O4���ؑo��`&[�R̈"Oȵ�U�O�@,:�c􄏆NF��i�"O��#��eM�����%�D�"!"O %�lNudB@˕�,J~���a"O�I�)̂e��8�bC,Y�0x"�"OP0�k�7-d�-)��I�l!��[���u�\E�l�Jtj
_!�D8\Jj��d�>:�&�3��W�Y@!�$Q�*:U�'��e�TD�򁀈,!�$���%D����a��Py���
A���N��	� B8�y�'ۨߒȂ��9V��Q�B�y�s�J튤eB0p�Љ�ς��y�k�A����Ǯ5,v*4Y�cF��y$@(k�t�E�G.:�=Z�O���yRh�	~�PZ2EV�0�*��I����=y�y�㋲-rT� �`V����y2��r���K� ��^)؄a�Y��y�&>�݃� 3^����$͞��y!:  I�3���AC���ToC��yr�ڦ$
6x@'B�569ڡRD���y�-�7pڨ4����+��Hk���y�ߴ"�p��_sz(Q����hO4��$A�`y�q0IC,����r%�#V�!��a����V�ɒj��ty�DA�*�'�ў�>�����mz~$����i�6���� <O��$6�I(m��*�e����RFV*�
B䉘n,�`+B8Kᰔ��-���C�	K&e�'�V��X)g�>l'�B�)� 0���z�手��� W@,����O����W�B�D�J@�]�B�x("e�3?!�dU> !�Cd���M֒%Z�B��&(!���Y�����(����¢A�`
�y�ɑsG�m�ŀV_~V�h�B$O�C�Ib�l�EKX�P�B�B����C䉷 ] ต�N�Y��$�_�yĬB�I���1D	N�FoJ����2�hB�ɺ
��A�g�h�6�2Tj\9bB�I�+h��h0�O��Ve�S��<
��B�-  �,놭�p�(	��,GC�I0?��Y�!d����L���V)L�B�	K��X҄O�v����N�1/�`C�� _0�q���(d�8��&U��`C�I�v�|\�Wk� {l� ��͹39BC�ɛ*�]� &A�-�, ��V��B�	~�����J�)`���a�h�/D��B��y�h��c�Ԭ �� bqd\�o~B��+Pǈ���"�:C�x�j�o�zB�ɟp��xa���R>	F�	�t;!�J�1|��h���&m�9��L3�!�d�K�R�K��Y�RX��0@E��!�$�/W�6i`wg[�|�P�7�U�D�!�
[䡺"n\><������	1�!�_./B�`��>�-@�(��5�!�d�/k`t�+�@Մ!c� �A��h���N��@�)F�H$�`(�K�+e:��+�g5D��ٵ�`��I +��C�X(�4D��0��\#{�>�ò,E�(���<�$�Ox���#B-�F�Q�����Ju�џ<D�䣅��DA��/wV%y�CЊ���;�Ovj�"�3j%j C!�Z�8��;%"O�X���G�>�A4�1^�N`�G"O���؅#�pY�F-��2���Ku"O�q��d�;��1�i��'d@\2T"Oج(nR"inޘ���ƟFPFP�p�|��'iў�ON��퓶n�4��¦G�i��`��ODQ�hڡV:� ��&.;��-J��Ik�OI
\�AD!�z,kB�.Ĝ�Y
�'����a FӀ��KW�^Ϭ��'M����L�3m�,[�.��D���
�'��ą�'�2�z�"U�Aq���	�'̖�)HI�!���W�3
Z�2�B�)�$k��Z���A|g�I��C���=)�y�X�PLRb�O�D�ɛ��hOt��Iׅ
dhp���B�8 Iq�̓,�!��Q5d�D11�~b��(AW �!򤏸A������>$=����\?/p!��AW�h�!���-A�rt05	�M�!��8q�l��fϘ'E��,�������	���?E�$I��c_v�P2?5Xts�C�<��O<#~r��̓B�։���L�j�x�R��~�<���]=���T�%��ȣ���v�<)A��U��1BZ0�� A�Xp�<iK����01�eN4@AX�ğh�<�$N��� a��ϔ�@{|�R���hh<I�o~xљF���u����'�ўX�'�~��Ө�3!�V
�R�L�(x���>�4����]=On���jЯp/�"OT�u�-
�"�R`��:p5r�"O���^!���;`n�?�����"O�k�ŵ{����$����hq"O&�ƥ� U��y��-, FН�7"O.�����0)�V�Зl�?)���J�"O� ��Y��5/�l�q��؍)$����"ON�����y�;�g�`n�*�"O��q!Ԡ`��@��
�0�̘�"O����g�s��q&ٻ ��0kG"O��:Щ���P���D����*D�X���^.n�x�!n��Gu��� L-<O�#<	�i�%]��(�&ɜ.,�k�N�L�<yb�	<5+!��*3�&iIDKOJ�<���
~m����
ӧ~���1#��F�<��-�/lP��O�"^QX\!�DJ�<��M�)�zt9��
s�ف��ZL�<W@|�$0������w�K�<�uF:�.�r�c\���4*�Fx�З'�>-���1���S��H���P�P���l=��X�hɭt��P�W�r�B�	2@��t
�h;��9���*��=�	çE�~p�&��% 2�h ��+3b�ȓwtX	��L�`�t�t� g��p��zk��r�F��O%he0���r���ʓE0�lj���x$� g��9���Dt��Ґa[[��`���8�((*I:D��E�a/�L��m�0_�$D��5D��X�- Q�J���:P20�*�f2D�dٕ�L&��BT2'_��IU�1D��A�̽&�)j�(�(����+.D���CN�)���!�0�Čpc`!D������ܨ��r�X�9G����� D�`�h�tE,| &`���tH�Q$<D��q&��3iﶭ���H�d���ҧ;D�����W$6�A�	#\�h�Bf;�$!�S�'x$����Hǆ0�i�FG���ȓY/x 蔣��h���`JI�.0�Ն�.Ap��l��9:�	t!FJntمȓ(- |B/V(R��!�� 3%@a��j�t�2���?{n%Rh`���Iq����l��M&<HTI�Dӱ��q�qC&D��&$ߙh��)03��4/B�}E�.�	e����3}���P�����3����B䉻J!����`W�f�`��a!OfVB��K���ҦH�.;��"ʕ	v�>B�T�fH"]v%� `�����B�I/#"} �&�����R�j�B�5H)��ǹ vaɴGQ��B�	1O/�iQ�ƃT��O[�~����0?����4�h���#HQА�%�R�<q�L�M�%�TK��RQ��/�x�<��l�~;t̙s�O�^�C�t�<y��̭fxH����u�=ʢ�E�<a�м2�6E�4{�UJb�Y�<I$eD;R��e��!>?���ύX�<�$�C�ڥ�a���W��!� .՟��IQ���QTkI�`�x����/NXT��-D�X
�PB�����R�1�D(�8D� ��L#oG� �f�U�6 ��5D��w]�̀�!��^6<{R�7D�d��Hꊱ�����75��s�0D���B��)F����B	Q6
���F-D�@�$F��^rU��<���D6D�졣.��D�Lm:Q��S\� �BH3D�8@2ŝe�tdJE�wd��!B/1D��!���1%H���(v�(-a�%5D��+5���8})r�G�Nˬ��5a5D�hpD��7n�2E녟u �D���1D�(�a=��8�OB�g�|x`,D�� ����\(+���#g���B��"O愸�.q�jy1��[S��d"O�=(aȌ$�Pl���B�[O�|q"OJD�"��2��b ���7���"OBAJt���[���IF�:��,�v"O��*U' &�R �I����d"O080AQ�c�͸I �J��5��"O( �SIɛko܉z�Dq�6=C�"O���/r?:Y����.�p���"O Q*dI�"}8g$L[�<��"OLh�'҅�,YՀ<H�Va#�"Oj�J��'|����B�n�4�"O��" Ȳm���+D�6��{�"O}��l�P:�Ap�� ���"O�I�M�%Ѯ �Qd�n��H�"O����7������~�t(�"Ol-1$L�z��#C�{�4�g"O�!¦V�B�\�[��őn�zL��"O��ɃK�������S�>e� "O�!����)b�;�g���\�"O����H͙����3gI+x���C�"O����ʕj� ����z��e��"OH��V�� �r�Qu�1�D0[�"OD���'ְ+�h|��bV n�T���"O(��)���J4raKF�դ)p"O�T��6I���3A�+u���Q�"O�`��eG:]�����d�,`"O���!Ѷ~yJ<�ꕼiH�-R�"O�����\���%+�6-b��t"O�;�@V�Y���VnV�{v�X0"OF0�ږ�&�:�Ĕ2I�d�"Op� ��(}�����g=��St"OvA���
x��ߚCL�C@"O6}е+��i=��Y�X<B1T h"O~��@	]3�b��d�)t�>�b�"Op s�j����R�З.q���"O��)#�
j����D�2�zp"O,�`�NB&:Й�CCp�|�6"O~}9ei�r���s&I�(
2��"O�p��$�¤�+��# ���T�'[�Ę�(o�5b#'G�#5Җ�x�ބ��'7���V�%j�r�ZT-�$lj`]��'��k��Ip5h��F*_|BM���D9�6��b�K%Be�a�Ns��	8Q"Od��L��d��#�����U�"OPP��=m:�����Jf�q�"O8�aQc9����w`P$BPu�&"Of�5��S8 Y�+O,!@�"O �c��3���`H �rp1S"O�\C��A�8��(�)��/ ��K��Ia>e�s����a�'F��g>��)��7D�س# 6a�J�y�g�0b�|=���?D�ę�j�m������R'_�����?D�����E.T�����d϶)2����1D��4�)0�H���B,;��y�pO+D�|�G���-�����J�0�i"�=D��j3��7��%�SG�K��Ƃ<��O�����G7tQi��hV`X��_�
^C�ɑ/���FL</ ��`��c�8C�	,D�,�`��Үj����―B=PB�	t��,+�J�2�j�2��H�*B�I/7t���ϝ>@�����[�CغB�I.?�V�)OV!
ܯ\
�C�I/[$81�Q��W�*9�p�#HB�)� ֭Z��@�q锘�V.�sL�ԙ�"O`�#��;��ajNۀH�^��"O��gi�(:��q��jF�^���P�"O��QvbE�l�D��=��Y�"O`!�e�5-d!C�?Z�D���"O�!�'��� EcR�A�@�tX��|��'[��ʣ��y��
�]�̀)�'0��d��L�F��ʘ,�¸8�'�pU#�X-@�tt�U-��m��'�R���FӪm6��:dg�*N}x�'(��rd^3��A��Bϓ{���"�'t$8�녾�N��򊏔x���3�'�F�0��|l�����_v]J>i�����&�������;|@����ڽ�!�z�̸b�	�6K"y26ŝ��!�$E�!0�j�j`��DN�x�!��H�mǂ����c�,��c�(~/!�DIl��9I@-�� ��ţ2h�2!�Բ������]ΤHyj�2���dB#`�`�Q�Y
�
��@���'�ў�>���A1�\�bJ�%B���&9D��Kd�A�t
,D���6)C>@��e5D�����r]p�0G���<�n�Y�C(D��H��!��;�B�=cX��b�9D�X#Ǩ 8f�1T(���2���4D��;�I�*aC,�&g�A�� �<D���U
в}��("0�\�)$�kp�:D�(��'�j�$)eb��Y �|�ao5D��U��+)� t�en�d�)5D�<�Q�<%Ȩ�"s!J���%D���Y,{p|�� �Q�h���a1D���c.�W��cu���F��|�Bl<D��խ�c��y"�{�b����:D�X��A.~�a n�z��%��"D��0Nˍ43�%y�NU���Pe�!D� ���F�-�2cT$����*D��k�!L�*3���ߏy�~�چC*D��aCb D�h��V'��T�A6�2D��Õ�����¡�"l	Rh�0D��ӵ�Y�f�0pG( �ܜ�e*,�On�ɂGh�h 4�(9�y�⠍"P�=�
�#������S�$�0���P<L8�Ն�\����&M��9���7d�8���_k�L��+Әau�y
��^0U6���/� ��S���;��l" �?��*�P��D�J3Q
̄����J��ȓoI"Iia�I�<Y� 1�	D���'	a~���9X�H�A��ߚ��լ��?ٌ�8�	м�A�(o��y��
n�|l�&�FE�<كD�8>�t��IU�b�4J�*�D�<�s��[7���`ᏜFt2/�|�<q�B޲X�BxrSi�Z��	�^�<y�ƙ���E1�]r������p�<a�Mǡ]&��R(�S���:UF�o�<�enH4�!	$D��ʌj���jy�W�D&�"|��غHR�	3!�AB���G���>y�O,tI�
mò�j���,\/�c�"OMPh/W���y��R�L/��A"O�H����֤@���W�>���"O���p�ʕ1��]�<Ĕ��"O�!�u�G9Bi+�oLc�>��A"O���3�B(�`T���HI��
V�|��)�B�Jѡ���Rp�	`$��B�$0|OD�Z��������0��8��}��S�?  ��6F��x�'_�~��"O�ю7(��pK�kb�
u"O��d�X�^�j �	D7X*13c"O��M"hX�	7*�r�ށ�b�Ix>J�-5���{C�!��3 E�O�=E���
�3c���t�Ԑ��2`̍�r�	i����i��"��\ x�����I�,5$.8��q �Zt �Q4��C'S��ȓ,ت��K/�h���Ȅ</:n����J���ˡ,�.|� @/S͚؄�n��m`�V�$�5�,d�fe��	d̓��ln���f5E+�!�x��	�<�?E��	�G� ���_s���Cτ�e��|"�'���4�\�cLb���#�[+����E7�y��E�d;VIz�˰q�4�t����yr�ZQӦ,S��S�s�6��㪌��yBjM9z(`	��� �v�B�Y����y�/�p*^�� �v��8�ugR�yR.Ƅ\c-D�w�����8�?����S��LyRs'�/��ܢ���ꘔ'��u�)ʧP��ӎ�,z%�0�%eG���ȓIt�����K�E]��q�E̞7����ȓ	���F� ��̇�5N�U(B"O�m��lX9{�؝HW
Pi�Ȗ"O�� ��0#4�m!%�&1=*ؚ�"O��p�Q,c�<�A��V'|86�
�"O��� �l�;�A�`y��!rW���'<�	o�3?��N�I�R4���95������۹�ybLU�1��T��.^�)���j#�y�O݋h���8#IE��D�3aF���yB [?*; `@ԨƸ(�9g���C�I�y����$��d�>(j���$>�C�I�T�%�Ԋ�+E���)�*V��C䉔v��XZ�l��P�y*ѫ��]�:�=�ÓCL�}��?`�СCh���!�ȓ]�hP �C��CBL��Ǌ��J��Q�
�+��0S�v�:w,��&��ȓ(���D*_9fB�!!�!M�4%���t~bʛ�ܔs�@�d�H��O��y�E���6QCkmxⅣ��y�Vg<���!e�����Fڏ�y�́�n�����9]��x+B�L"�y������ms�� P4�M���C��yr�Ħf(�"C��tꆴ� �X0�yb�>^=B-H4�D%Y�\���e��y�� ���V�W���u�Ķc݈4�.O �=E���"'�ju�Tb�=W�0�u�R�y�(\�VM���aH�&{~��3kͧ��'"���Ï��WK:xV�D���k-2D��)D�"�j0�䢃�x"	�`�2D��p�-��uH���5lA�_��y�
2D�d ,a��	�C
��Ie�(�G�.����`U�ʯ~_$�+V�Pg)��ӄ"Of� U��*&���bث��e(�"O�\Q�Q�b��jt+L(�6�P�|R�'��Oq��k��ұ8�5 �`j��t�r"O�4j�lE�y_\4#JH�aDt�p"O���U"´P!@�J0�V.H��	�"OJ�.��}�(�ᆀ	U��l�"O���'N i���DN�dՓd"O�]H0B�?KV%Aw`ݞ>�����"O��	�� �(�����aU.v��yc"O�Y���0QB�t���lؘKT"O[c��%�vP9e���-\T�("O� �<s�����t�U�F"?O~!��"O�a�t�U8@�z=AW�� <���"Ovu:�+˛85��x��	Ծ�13"Oݹ���jZnx�v�ӷ;�`���"OX)dƕF����D�[��)[�V�8��C�S�O���X!HM�[���X$�R�[�N8�
�'�x�JZ�5;0�!Tj�C�Z��
�'�RmRQ�[�L�r=���5����
�'#fd��Q�k���ɞ	*� ų�'SP�A�mM:kn�vꉽ.6�k�'tx��Q�-y� 5�hIP�}�<��BÌ����M�'T�A4��u�<��nE�$ne��CN��01�p�<I6�B+
N2�;�H_<T` ]�W�Xc�<�ĭ]�����"�[�_1��@Co`�<�1FR\�T��Q5\�ݡ��_�<Y�h�:lX��	hy�1s�%�`�<�6ɐ52G�%b��V���)�`[R�<IQ���J������^�^d�<9cB�{I�tc��D*4�Լ
��-T�����
��~�!�G��|d
,�p?D�\r���?�T��H���ٚE	=D�h��$H�E�h}� ��
ms.���D9D���	��F|Q���L>^D�b�6D��1�>S���Rf#�7	��E)D�\I��=P��������s+#D���e$�,4.>H����9^dص8��"D��Z��5HŠeI%��a� � D�8�7�ۓX
�r��ۓnXa��=D��8 M���}��ܐ{����u�:D�$�`L7)O�yC��\��^���-7D�c�/�w㘬c�f�Z���<ړ�0<	
��lɉŕ�fB�| 7�m�<y�c�LDD��P�-BV���!u�<1�U�R��E�ԓ8��d�CH�{�<Q$�?�u�c!�gA61��]�<9�� |��8�ŧA&�j(#�MJW�<�a�ܡB�4��ƙ��l�&_W�<�C�z�Zq��[�E ZUp�m�QyRY�8%��g�ę7GE+Ѧ�3�� �"#ըVF!�&V�@e	�e`���q�B��m'!򄅏i�~�3�	�]���֧܅f	!�ĮA����00O>t�&�ˏ	!��׼v����������:��չR�!��A�w�(��;d�p��ɒj&!��Ɓ�H8�Pn����,	@�O�Q!�\�p'��g�d �Ѳ���N��I{�IC
\��	i<�䦇6Q��Z P,�ְ�'%FZ�<�2̛2;���N_�RvȔ�t�T�<�bt@DM�P��G|�����j�<Y ���L��ȫu���d�d�2��Rj�<1s�� ��`th�=��ҧ.�[�<��Pcz����I6)~��i%�Mrh<1����YRL-dA.@(����?�	�'�~�v捒]����e�W��\4��'Uԡ8E��6~ID����Z�Di�'�$c@B�4!̔#�)Ӝx�l��'H�y���Nu^�Y�	l	�%y�'z>!���>PC@
�J	<f=�����<�*�����{(��k⨍�KR<lS��'1!��ͻc�fp��ְ�h��5#B�nJO��c�/�Zaj1��)��<��5�V"O8��Be\�)���
 �߄j ����"O�� ��K'c�����/9�x�"O� �aQ�HܥyN���FT�L�h�"OT�+7KN�"LP� M
�V���"O�����F�L�!����d���"O�b�(��)�\��[F��x�<��&͘Z=b	�g��GL����Z�<�U�(Gք�p �6
�p�IQ�<f��/(�\��i��P�!��X�<QcJ[7	��pٖωTRy�`�T�<!���%��:3aW�IGHd�V�Kv�<q��å(�:M��ЇC�L@����w�<��@�F��@pB�J�m�W�W�<	gd�-"�6e��7[J�aଞT�<� 뚭�<%	�!�6/`P٦��g�<I"T�t@��c҆N �%�p��d�<A� ܗUb �S@���J�`����U�<Ad�@(����6,�4�t\H�EP�<Dc@."�"�.T�0*�AxHUO�<���[5%���v1�#�kH�<	ѥ��^�,��e&�X@H�@�<kXT�IHO�<g��e	�\�<q�H�>b���r4�G 2W�)�dM�D�<��|Sµ1B��%`���� �LC�<�3��K�Q�#J8E�f��A�<)���4?1(�1���5Ն��'��t�<A��Z:D�y�@+2 />�1j�s�<!��M�)B��:��ޱ240��p�<Qk�=+�,�nʰ9��YpN�b�<�Sf&#��(�ߩް�����]�<�$�V�"߄�1�n�m(hq·�^�<q#��#:b-is*�8��jLc�<���W+�Z��Й�|���WG�<�N6C����b�;s�ji��@�<y�Fʅv+��zH>+�9h��@�<q��>M��*]�M�J�CGk�z�<!t���,�<p00N�SZ���҇Yt�<ّ�]��� 3���U�yKQ�Lq�<!�@�*Պ�G�8���E
�F�<��L�< ZI�9J�7!�w�<�@D/Q�P����M����ˆ|�<�w�-,��9ju��3���VK�x�<�@��"�*�9��#i>�]��N�r�<i!N�'I��i8�� �,;&���_S�<�fNK������OJ���w�ON�<e,J	&�pM�#��$a�)����P�<gDT%:�k��*Z����'�A�<��	�'�.m��#�$���`bJz�<QPcKִ��R.�d��ؒwR�<Ic@�k��x�̜�ePv��K�W�<��H�#:���&�X��Ej&�[V�<!n����3�#����N�P�<�c`ŋ3�8�@�R&6�P��#�F�<�TiL�(e�)��ʜ$Y�x���mTi�<�ӭ��YF�N��1`�Yy#b�<� ��*��Y9&���L�A�c�[�<��+�$$�n�z�MQ�;�Z�Hei�_�<AE�F�lL�dY�Jw X#L�t��y(Le@3�
>�-�7-pZ����J�6����񮁒�d�x���ȓ
g81ir��0Or��B(s1�Ԅȓ9lD�s�G�
{�	�B����0�Dx�#P��F�an��zH�ȓ }�	���+eq&�2gJ�k(���ȓ(*�h)C	·L��*��VT���F�Τ��i�:E�}b��ѬrΤ4��S�? �,����Ae�p�f�d��4"ORD�ǩܗV(Z�%$m�E "O�,1�(W,k*�XqaDI�`@a�"OpL "�32��u3�E4;�3'"O@$a�����	�1�HJ�2}C�"O6)pD��ʁ��/U�y���K&"O�Q�1W~���2��.�����"OL��@k%8dTS���e
�Uä"OĴ��� ��		A6{�"��'4@q����0�(y��H�u�#�'�s��0�Ay�Ŋ3?�&p"�'ע�i C]$bI*`)P	V�:.D�	�'�J�䫈�k\�P �A>8BnM3�'����
���y�D�#.(�H�'*4I�-[�h>0zgᙑ�����'����W`�{�=ӶH�\����'S� ���B}�|[�
�XtJ��
�'2z�GoQVY��Q� �5Q�^�b�'\�Q#�n:Cq����&H�5!8��'`�xѦlP#ڹ�@ӧ'n�%�'�>��M��If�qk1(O%w�h�'3F���F�D��k�CJ,���
�'�bm�� A�X̊EQq�В{c�P�'��5ã?I�D���
woZQB�'�{�l-� �V�Cި�	�'�`5)u゠ ����u�P�jZ���	�'��<��	�"h�1z
�f�6�K�'����.l9�p�vƖ�^،�[�'ŤQ���G�.t9�.+z�D��'���P�j��m(�[:!�N�q�'RZ�i�56@�uA3�[�/���
�'�����#G��\A��K�����
�'����B	@�Ln\�� �(�
�'b���6 e�}��IS�g��	�'>�����,���*�OL�1)�'�����G�̀��,��F]��	�'�2�3S�G�����W�'���A�'��yS4l*UNt(�i/��LX
�'q y�0oT�3�
9��R��0S�4D�`��/׏MmJMs�FL�Y;�rd&6D����BQz�0��uI^5N�%�"n8D��i�f� �6x�0)^?i�����4D�|�E��%��v�A��,�#�!�D��j�<��$�f����F%!�ď X�(u����
@�d ֩e$!��-H�[4b&n�F��.˾�!�$�[-P��Gɗ$���C�
�!�DV�U�@�$��Hi�+c�!�䝇�8�#eg�a�*Lے�r�!�D�c�Ha��R�8Ts���!�$|
U��n�\Κd��iܪJ�!�,�p"S/�]�`\��S�v3!�䗡k��ܸ�&72WM:%�ɫ�!�C(T���`K
_��!wj%�!�ě�z�8Q�䈑12�^Q�"#ՠ�!�$9���'�]mLųS���0�!�Ċ=�DH����5b9��� �L�!�$�U��bP|��DP1灠X�!��� [�|��Ʉb���s�
:~!򤈖?�̔�ql��
�X�i��#{!��1{r0���J�!�#�+7r!�!&�
	`b��{�<(!l�M7!�X~st4�$l�2B�d麡`E {!!�d/�`l��K?=����3��&`�!�� ����T%�u���h}��#"O�l�r���S&m;Q���5	�T��"O��8�c��-(:���"v ���"O6���0>H���*�\eb "O��)db���ppO�7;�"O&Q�wkHU���I�e��P"OИ��mȅT�
�q�� ��q�"O$\U�(ft88w`JI���CT"O��$c��|M:���.�&�j̀�"Od��dS�K���k&��:z<Y�"O.K�4A&ƀ����A��-6"Otm�QeȦlT\�d�}��i��"Ol|��KO�}"�* ��0*����"O�͒�
�
��+��ƙl��R�"O�Ր�G��r���B2�ːD�Iڶ"Oڝy H�����a����"O A�C�	X����ݨ;���"OƔ���m%�99S��@� e�r"OL�R�'ߖ7����C�21�*`�&"OD,3�χ)�����4+��a"O�~4HU��_!+� x�l��!��qJ|@�^�w��p�C��	�!�����Bt����ǎ��!:�"O~|���Ӵ��� �o�$K�>i��"O�E�V� =�ʭ;T�ٖM�$���"O�݈'Bʉ�٨�/ӫv L��'"O��X�└|�q�ș�����"O�i���?�V�#�f	<��� �"O�ذ�8fa֕�2嘨�|a0�"OX%���"+�4���^�l`�{�"Ov ��Ӛ�X-��Gʎ���`3"O<`���V�x-�AM���d8�R"O  4��g@� ���*��Ec "OzH�&���B<�H)"��"K��H��"O2d`C���v��1h�Q�o�Ҵj"O�a���+S�f=�2#�D@���"OR�#$:t^Tq;3"&@�Q"O>���B�G�F�ɐ�ǘce���"O��5�E�u�$\��xG�A e"O $�N&��RT��@��K�"O�9p�c�7|n�p �ȠW���"O&-:$a
�@/�:�h4�V�:"OL	�']a���8䈎-��
7"Of5
PnҴ)W�8	@gץp�� ��"O���P�-����EA�ph)��"O,Qe�a@1��R�fN1��"O���F��%
^�h���|�4��"O�3���.v��q9��Wm�pp�"OhL�d��������%�b	�"Ot ȃ�Yx@��7��4����"Ou�`�E.aKdaH��$@|5(�"O<@Q��]�!�"hB�|>��"OV���wX�q`��p:F��"O����m�8
whe���qDzт6"O9��f�~6�k3��h6N��Q"O`q�**u�H���֎]GM�!"O���b���|l��'ƍn���"O0���
�=6�����;ĞDA#"O֩p�	�>��:���-��I�0"O�I;5���y=da�K�7G��(��"Ol��7?H�<����"l��ٵ"O�h���&!C�,��T����D"OL$�%P�d4X���fr\|`p"O�`FF�+d�t�p%!V
��r"O� f�����bI��7c�88�%*"O<d � �  w*�@u,���c�"Or����!2l�P�J+P��i�"On��6.�4��}�fJؗ
�Ȍq�"O�����X�v%�D!�^�c�hp�Q"O���W�k���t���=b谅"O>�Y� m��aʃ�(��"O�$�� �+,�(DhCN)��hQC"O��K$��*2(]r%mۮn�y��"OIf*ǒ-���re����xQ"O�h"�b����a˔�*�d䨱"O�	�ue�l\D��g�MZQ"On���$mv`���ԝ ��]1�"O�}@��84�
��N�N��"O�d�ЯT���(b��%���P�"O��x$
�}�,Ӈ��>V�X���"O:����T-⴨�����;t"O�y0-A&� (�s��0R�K�"O� 3��U����wf��PSw"OX����>Q�s%�,*��PZ�"O>TAR�6�v�Z3�F�
�����"O��Q�C�kѸ�D�<r��U�D"O𹣗��������P���"O�آ�͊�,�<�kK?Iy��Qw"O=J%��b�����Rsd�8u"O�	�"ď�Ԋ]��
S�]4�*"O܀3��D���B5I*����"O��e�x�>��#BC,��p��"OZY��#��D��ٓGU�j0I�"Oȕ ��,�ȲUGS� �ju�"OrB &��#�P���I�t�B�)�"O<��ڟ$UԱ#�+Z�l�*�H�"O��6�p��I����	��i�"O�DH��ػ/�$2��n���;3"O���P�j��0c"�3�P4��"O�9 R����,@D��!^��z"O����o� x�H�K �9H@�"Ov�i��6n  r3`Z !X|�$"O�P5j�y���hVMՅB�n���"Oܨ��-�!�`9X�Ů���"!"O��@Ⴡ5 �@�V �{����"O���F��y9��[�n�"�n�(�"O��B38wN���m�G�0��"O�l�̎�Ƕ]�4�:<!ӳ"O �h���]���:v�4'��T"O�<�J��E-h=K5W�,)�"O�1Ҡl�r|�q㥫ȉ#��|ca"Oj<yђ}��!k�yՐ"OX�
��ȗWk:��&���~T,���"O�t�P�I�P�R�ݨm�va�"O�KQDЗ���y�"��v�,���"O����%?9(B4�V"�c�"OT���
��h����1"��Y��"O�胗�E�m/����	�;��i�"O^�r�J:A ���h�>!�pbB"OpU�t�N�:�d�"�I��|Ļ�"O���3�߆1h<��'� 8�2,�"O*Z��"!�D쏗|t����"O�����f>]��jȬ{�QP"O � /�zQz�"#�ĩ"�@-�"O~�zS!�.8�w�X MCr8W"O���G;Z뒘`ׇ�P0P=��"OT�J�I�+��}�b��1~ȁyP"O�s���&9�����)��t���"O� ���� �¤e�鍺i�d�*�"O���֜U��\��F�V�����"O�5�t��j���y���`� "O*9���O�|�j� �|q�C"OT�y󭍄[�R�iB��^
L9 "O�p��d��,e4Ei:/b���"O\����!��9��.{U�Ъ�"O^5����YL~�� A�QS*hy�"O�#4Ϙ1bzJ�� ���X8�q�"O�a2��#��eI��ס0+.���"O�h�g'��
i����Y�p�<,#q"O�Y��b����;�@��m�ze"O���)S��G��)$S�P�E"O��
d ),^��bOզ6��!"OܴY���$d��3$�J���"O��Cڈ�l�ע�C�Ic�"O�!�l�(Ϫ�id���Y���Z�"OHd�Ҁ�A
��;!�]@���"OJ�D�ƨg�s�Jۍo�6<;�"O�\#����s:Zl�
ϾU�`�3�"O2b�&�.��$��'�LyI�"O��;�G�:R�{��J�s�l��"O��(Ǐ	y��QsT$�� ;@��"OL��i�h�^Q��[�|!��"O"��'�0+������P$��P��"O��kcǓ4��#Ĥ�u{��[�"OX	��@�8'�\�!��S��$"O@�j�(}�(؉`��Zc�Lô"ODxˢ�6$������H".���"O�F��X��O΅�4Q��"O�x"r�A0��R	�>���h�"O�mz�	�:��Ԡ#ذ ��EA��0��a���H��U5I���ɬS�8La��9D�T"&ɛ�gڒ}iC�Bl%i��x���sӌ�qD�\�|K�5�t��3��	2�'R�O:��W�]#WHp�c�N!��ɩ"O���g����#�O�k�20��D �Şm"�����vd0���ëIǨ@��"���w��Y& �`,�p�H��'���q���S�`a(X�DJۊۨ)Q �R,�DC�ɔR��T��ϥb�`���\�QghɅȓ1��#�`�'<Y�H��@^& )�ȓ;X��IRB͹^�8�T�!RŇ�Q�H�aDg�"��]"�V%H��%�dD{����k��fh$?7���"�ٟ�y�h��`��C�$�/Ak�L�q�ۣ��	A?i�{���.	[�0�f٤Xhb��ŤN��B��|��i֜2�1xTG2c\�ɊbP�ad!�D�6@�d�ǯ��Z��u��#U�O��=%>! �
>hhT7�T0a�"�pu%D�,8�-��$�8]�2��%���8U�$���>I�y��TEN*���`���BDr��W����y�V�Q��, ��=���9S�I���'azb�F�j�e��34،ͻ�b���O����FڧJМAb���!��PЍ�<����DP�-�8@�D�]�q����	z��	A "��E���%̬)� K�Ji�C�`�:���j�Kfr�K�o�+���O�=�}� �kv��C�&x>l×�DU�<ɳ�k��]a�j��Ք��$�N�<���̐k�\diS*��#�6��Cb_G�<���	;�8<�B^��±�����<��e��@���j�B��ZA�Xb�L�<94�]H< ���#V����C�`�<� �����D�[��:D-��!����F�'9�*�5�+�6�2ݓ4�[���B�	�a]�y��ʴb�ĕ�'YwC�I�Z���!AA��ʕ`C��B�Ɍ���!�h��?PN�:%,T�WB���LU��ޜs�6�v�\� (�C��w��Jd%[�2��P�1�C�I20h�uc�ϛ�hy*�'����C�	6�����.M�$Zhp�֎��GT�C�I9m�(�9v"U�{�^@q�C�T��C�ɂO�Es�8���#EJ���C�I>qs� ��I$A�5�t`�?Mo�B�	?7��p'��p� i!��[��#=YǓm�d5�$��&t�*9��SII���ȓP����a�9���R/%f `�?�	��&�%��3�� ��W�i�,	�Ɠ^�x��	_�n���c��HS��ⵈ���'9�g�'`p���FgN���6��:?�>Q��ט'��K��M������Q=���O����N#�JUA���w����2�Џ(�!�CL�V5��4*�t����!���b���np�pϐ�c��	]��|!�eH'��Ι>K�؍YG�5���	�30<��N~a4�S�&ܵ(B#=��O`\uJs�á>_j)���P�+&���Rl`W!͙$�p9�+ fp�lZ_(<a2 ��b�j8(�G
�4왕�UQ����?����>[V��c�ʂ��%Z��FL�'��y�/ή�T�xT ; ��`Ȍ��y��':>�"F�6�<�W�Y�n������,d�D�@����(U�޿n�z�͓�0=�L<Ʉ�W>�F5�tǀlJ��3��Y��hd�x�͜4C�}S�jS(b���ʴ�ݛ�?9�'ұO?z�F�ʆ����\�y��iR�
H�'��':����H�
-���+C`X1:��@C����lZ^�tb��bMtd"s�a�̕) ���P��I�*F]%$�K�J��p��0<�L<g�±`|x\r7�Ȉx�6��$ZX~��'��ѡ�ꀔ]��P,C�Ry�x�
�~y$�Z��tPň�q�"�y@bD(rA����|<X��Vp`j5Q�&�#1��d��ɈZT�'��
q)(Nĩ����ĵ��Eè��IR����{���7A��w")��s)W��(O��=�Op�M��n^�:;���{
�'�����%M�Y�'��C��M�	�'�����nI,��/ �@Bl���'��zv�Εfʌ	p۸6�09���1�S��Þ0&,�UH�&m���,�)�yb�$oFT��δ��j�D6Ƣ=E���o�X���y'���ÆY,�^���H��$BƐC��Ӡ�N(eFP����hqaR �f(�h׌c?VQa�fX�p>�O<A��I5u��X���(�t)�C�<���(�~t�CAK���d�J�'H"=�OR�x��O
$4�-S��4f�H���V<"�P���tΌi# ?(��͆ȓl �)�Sn3lh(�I�kۺ���>	ߴ�hO�22�A�s�/|DR�Z'�^�L��C�	/0��)�]	�>)0a�J ���IC����V�K6,׃&S9#�HC5 7�]a "Oi��`�t	�W�)@�LŚ�"O�P�tUN	�e/ܚ,�TL{A�'��'}��R1�����V�l
H-�I��y�DE�֜���+a�@�x2��y
� �:��Βq��m�q��K��"O�<���ٲ:P> ����NH�S"ObY�N��)�j[���mږ"O�;�"��vLX����n�^��"O���kԱR�m�P.	�|��%�"OR����O��51��-!�9��"O&D��C�"�����b��*?ąr��Io�O�$L�/�	JWVx�K��t����'`�Q���S�ԐP���-iNd(e^��'"���3}2m�8@c\Đ&�7g�����#��y��W,(����`�
�d�����II��(O���Ą� pA�EYx������!�ArV<|�$�F
i�L�0h���^���/�2��K�'.z�ɲ`�b�4��ȓp����@�"�$h!t,[>4�݄ȓw�\�S�O����m_�ȉ�>��>�>Q�g�&б�`��8��ȓR��T�֦¿m�~l���
&���=9����D�+s���z�O���C�	��p=Y�}�	$<C��p��C*V��AU�?�	�'S��@DbS.~�6���.��l_�H2O��"�]i�S�'2�
-��(�
@�<qp牊e���ȓ7~��٣O��Z@� o��j��>A�ÁV}R�I�:����1_�ĳ'N?H�C�I�qb�h�0,Ѿ!bܥR�M]��"�'�\-�@A���y��.�� �V���'�2%䊃.pSa�� 1�'3�Y�An�>"�}KE*��tݢ
�'UL����-B�t&�"	F��K�'!��+���3L��$���-Ԩ��'H��B!���f�ش�� �<u��'�R(�$�.�Hx�ė�{N`��'[�D����v\0��lŬt�dP��'�v0�Ac�uZ�;�NT�j��0��'�`h�pbvL��*��6E.��'-(���'��un�
�lU�('
L��'�<aْL����|*A�ZL�n��
�'N6Ԙ�F�5�9
P�a��@
�'<ؔX��0?��q���4=�$T�	�'΄š�L�X!��{�M��Dt���'�ayS�ǨG�JA��DD L@�'�Ĭaq���G׬��w��#L���R
�'	h����]����ǰ�Z�	�'m�h�Ŝ�h8��c��6�`��'�Br���:���aV��$b�,� �',`�au釞
n�Zv��e����'�%W�D�H��q+��γFCD%��'^����ъ2 >�8�*p���k�'�����ş�j�L!�'P�r,��'z�#��H�MB��B�&�����'t��(�gJgL\8���-BZ��'?x,a���J|�EhGi�x����
�' ��9��B��0�V��#�y��'��h2i�-�2��gkI��`��',`����3#����(�). ��'��{sAӦM�~�j7�W6}�����',���2�!�.�1}�*��'�4$��Ռ(|��ɬ]�p y�'�d2a��	OD���U<Y���x	�'Ǯ����+ Ø��@N�S�R�p
�'��]�P-�2�>i��C���ǘ/�yRHu8<����� ��DQBi���y"'Hb�B���c�0@ "�.�y�o��$��N>d��0kG-��'��=H����q�(h��S�)�z�;�y
� P�T!�R�*y�FAN�+�H<�*O��i"#@�B����C;b��t��'-�*�#̇K+��`AK�"���'�4�@��F�d��0h@�ӑ�R�B�'P�I1��#e�䣒#��|�����'�ֽ9׫Et���²�\j�T��'li���ϗS(��c�ą�Yf
�+�'<�tB�D�-U��|�H�j� ܩ
�'����Y;!{�%�Cd��e �'D�IR�Q�$�S�ͽ6<��	�'}�mp�������#Ԥ"|���'Bb�s�,�7IA���e
�#�8 �'�8��֡Z�]�C���'�^
�'����¢�c:F�3��F;�)�'���&�7i������4< }�
�'�v��V��%�h��A�YC
�'�z�@�o�,;S  bT��*a�4<*	�'ĶY�6� !� 0P���-����'yJaX�R���Wh�)$ܰ�K�'J8daǌ^�H�X�X �U��6�c
�'��¶N�P�B�0���
���a
�'O��r��V%id:a���x�%D��I��)�\�x`�;V��U�4D��S'��L¼#��M�҉a�b4D���mU�a��h���0�dp�c�>D� s��U!�6T��� !��CR�<D�x$Ǚ%@B�s��&WÄ��r.D��e�;<�j�k�W���1l/D��Q���"�0s���o�����+D��;�M�m���8[<*xY"+D��k����ms\�!@����(g&D��c	4�ze��K�SǨ�I��%D�x2�oٵm8��c2b�#`?���P� D��h�����-�gGװ����:D�h��F>(�)(e� J��qb�n,D�0��"V/2�V�C`�"�Љ��"&D���֪'��U07�ɫ eTMM�<Iâ{N�(�E^&CKD@���H�<�R���^8 ���� �qmUQ�<y�1P�&�
E��5'5.Ȋb��N�<��g~f�pZ��U7N���R��b�<A ����n�'aW��&$�b�F��L�5l�˰\�'�r{R�[�\5��9�/��`5�	��'!D�0�E�(&غ]��@-7h��ʎy� �5m���V�L�O���(�Ǜ!\L��ܬ8YxS�"OpD� mH5	,�X'&Q��2�bFՊ@��Q���J�|�g����>�0�t�ϴEf����Bס�$.��ER j�=#!�P�ïؼ=Ub���i�& ���Rb-�O.�8��C�~|��.I��I��'�t`�Ae�-O��a�:ON�"c��U��	�1. xb"OZ��
�6��%��MPb 4�0�|��g*�j��Ę=�?Q;#@
�x��4���R�k,D��9�#��ML}�d]�(�@�53:Ё���<!� ����m�&�J�b���RB�G<8�B�I����k$�H�9{X�@e�؝3'ب����C�����N���&��(}�xb��#D�h�l)<O�pJ��E� C�@�Li��Q�i�D�~���f�L���ac@%D�ܐ��'Y���${����&�Iz ���GD�h�Q?�vΈ�K��ʓ�߄{�t9�VE#D�D��fC�0�qs���)� �z�H�{o2��H>q� �gyBW	8^n|�Ef�o�V�z D6�y"��	�T<`l��T��$CH2�yR�I�aB� �Ԏ�
c����˱�yB���|���R��t�X��y
� �a��/e�4A��)t�BX�U"O^jB����<�:�l^4=7f��"O��9t��QnЙr�<8U�2"Or�{b$.ELt��798���"OX-).	&^y���ΫU�c`"OLa �m�`[*I��':�$]�"OV��i¾p�t�Q�*r�nYb�"OB�e
�f�| t����J�"O�%t�?��T#��X�J�S&"O�t��c�A��%h��ƛP!���e"O@�AD�bTt䳧B܀�u"O^�S��W�b-dDsBQ?�\�9��>��f����S@)�82���aM��ˆBΞ)��"O*����3|��b��ưg�V�8��Nnb˓���rc\K�g�$�|E8G�QH�B2��gѴ=���#%�pY���P3�`�e���T����ǫ�m��19E�N\�a}���C����Ɗ�>nq6��dܭ��O
�fǚ)_����В����'l�zh�����,9�Хl5!�dP�~H�Lޏ.�V�C�4C�	�{8�;�N���!��S)�6aQeԟDXA#��.|C�I�.����!�!��eI��/`.��@"ͮ�~(,N^MQ����{2aؠq�=y5�O��0 Sc����?�g�X�w.غ��6Aa�`dfG*Zs��ˆ`��A+D��Gdr���{��i�>C��J���G���᧪����$ήV�c���+Ԃv�q����������1A��
?.�ܣd��&�س$�P���c>c���?R%�%�1�M+!���a��<�� ��6���Sk�l��	6<h�Aԟ��w����'n��Y'T��4p��`5lX@y�ד[n�0m{�N�)�5E�d�vJAd� #A�!-���Rv�(*����T��k��(9X�H�8��Ԡ{d�C���⌠���d�A�0�{RA�"l�ix��۸p�:]ðH�B!��ᙅr۶�4	�lp�'��R�d6§1H���SҲ]���!0@/J�����;�6���Oa��ѲČL���I"���Po�AA�MB({P~���'�` �I�F�0��ǥ�{F{�Y"�� ;��0[�H��m�>�ēf����V�[^�����]C`�����_��f��6p�ey��Y�>����fkKi
��B#�'�j}��'66}�'�ę���6�݄�XTa##3}��D�;����'L��x���X�F�o�0]���/~;F���G�YŀEpH��>�p��D��}1^H��ӨM~h�1B/҆R0�r�m��(��D�ם&�,qeCA��M�o�&S����D\� `��pbl� Q��h�c(Z�џ�QÃ�2~PR���$ə hp�����&]:u�s+�J�2��$�j=b�&?��	�$�	�{s\�)@-^|�
fύK\��P�P�1��?2*ӧ�ԊX9<:Y�c�o�:1�AaI4�����1��U��&/�xb�n!�q��A�8&ʄ95B��'�$����uk�`Y��D������!�l��$�ΞK���BKur��W�#�b�C�	8
���2�ڇz�LI�!��w�\�� 
�8��'�Z����i�Zh!g���x�&a�=CO�rÓ+\؈�@���h��8�&��gq4� M�"�ʼ�ȓX ;d�x��m�Ө�p#$��On˖�љ����O�Z�HTh٭C(6�5��/R(��'~ 5p �N�LI*�p�/đR���	�'u��� �%�p�!A���#�
1	�'�^`Se�˵a9�m�'�ۊ,7�@��S�,�d�V�B��q��=�V��ȓP�С{�aF� Ī�Տ�2H%�(�ȓ欪�.TQ�	kC�D�)O��Dy�$��	�F��H�6���sS�c�2�O��yr��O\BlƧ��D|1T�P�[�4Xє�ė`}ɧ���DY�P�M���&_n��[��(-�!�d�?lD~��6l��rTƎ"�R�W8h�ؽ� ʐk؞�!a�Ć@o\Q�"аu�ٱ��5lO�	:v��0>\,��c�i��Pj��K_�УtC�gZܫ)O,y�S�����=�GL�K�H2A͒�:R@ؒ�/Sܓ)"fQ�7?d��I�O�Њ�Oۓy�Е�䄌:(�b���V^�i�r�L�<	GB�y�`Ly�i�,l�;�*�t.��I��d�Wr���=K3���,�XUЙw ,�97�H�"�0��R&�h������� .QQ"�Ʋ���S�$�5���$�R�%pt�@OY;"JnPS�J�.YyR�Ǳ��������^�qC�(@�P��f��D��Z<�
��� `6mŎN}�{6�G:d�~9:¡̋l���Ot���p��^.DB0�a��'݀󒯙�o2�x��X/��-��{bW�[��v�ؖ}���#>�vu��o ��?�e/��" ����s/P�Kb�ͽ\�����F �	��ɯ@���F��>!��+$AS�����'�;"�:�?AAII.B����'R���/~f��p7��W����ߑp��C� -��h����x����7bV��h��p�p���H͜C#8jƕ�-��P�iz����cy�]�]Z<)�M@	W>4�BM5Ȱ=!ac�$�X��i��<�HE�Ht�[��Ĭi�*u蔴~�L��'$��S#^�Ҧ�ɭP�L�?����!I�رP(Z�0'�3���Pyr�¡i7Ƙ8'�Ȏ2A|�����6q&��̋vȔ�H��)z���V�1? �b!p���%R����f�'�O��5����q��.�-����Y���fi�9A1����N$>5t�	�`��i�(�#$��;G���4��pa�%�%ق���JӰs�<���ܦMx�x�O��z� Ţ$/ 6^�̰�c��n����ѯL�H���
:�2��/��	�(<z�'ʊ��į�.��ԉU(+����䘨N�.P `�0��d@�g�"��,�)0�굠 ���9�4���� �h�B��	Ĵ�cJB�C�FR��6;���g#ٻp�{P�1�~�W<��h�c^CyB�^�f,c� �~�h6�M�iq�A�F�b�6�q��ɛQ�wը���c��3�Ѱ3�Z���L��<�Fd�'e6�ڥ�uv���� M8}�P *&��*]�Uq7g�����n��Ԙ�O�S��I���_�p?��'��OdN0	��"��b�-��3p�غ��� A�
lk�u��!#'�-[J:TI �<@E �'����an�����p�g�'V�8R�����|����8(Pv�H�"�qC�i�V��=G��/�^�+�.�=Ѭ���ɜv�>equ,/�,Y��_�r\��ɫb�T�@���-��Sr�	.�8����O�}��=� d�.)/�0�2$�p���E+X��Px��׵w0��zwT�w&,+���h�Xpd�V
;Z��6�ǻ[����S�V��'^H�9�Ѥ�E� C �%}�<���	*_J�1�®ܮL���{�.�u_jd�$G�(�����ؾQ�v�r�U��G���;q��x���'��-�I�1oH��ȓM#��9A'̟u���P�3.����'}��k�3 Ȱ(��	�'ĬM�ְ�����Lx����*N~�mA"l�0��\�@¸����)3�K	�'��:�"�7�����N>"C���X�WB^��3��`�r�P6�Y�a.f�C��ծN>fC�ɱ( ���t�C_�nj�l� �ɦb.�d��ӸK
�$`�ķF���0�,�1$������y	`n݊e (HTƚ�!�
(%6������_�B$R�F�D2!�d���B�m��B���pe.�#!�$A6�杸t����)y��X?{!��D][�E��J�J���'�!��t+䖄`�+Ƒb��[����!��Ҭ>l��"`�3|��)x��ڠH�!��$w��i���)���A�ȝ:V!�dK9W�` #2OMڴ�@�A�EZ!����X�I@+�V���A$����!������SoGI�z��Q��u��'f�� cK�_+*�ɀ�S!�4���'���;AX)
�^�р�ۻ!΀���'&N�bq(�<1�ԅ�mS	r%����'PL��b%�9\�,4��jRs�4�9�'��
VK��|x��u�U/hz�a��'��1��$(���
n>0 q�'"9��-Ԟg%�0�B���
wi�i�<�eЮ5̆�c�&��}]N\�E"h�<��b�. G�Jlʔbй���g�<rH�]9�D���B(/Ќ����\�<��bA7�Dl�-�'IS�y'��_�<�e�<ܒ5U8�,9w��r�<ѓ+� �5P	�?�B#�o�<�@�I�P�J�*&��ɑ+�k�<y�fN>Ĭ$��a]Ȑ�f�d�<�� >y`��Dm�.�P%!"�`�<� ���pm�J���iJ�OK�U�V"O��3#n�25��	O�E:Z�0�"O~9�Ц^�:ۘ]���9���v"O(iY�.%4���钌_bl�g"O(��W�A''\� wG�7iV�!"OJ��#���1��<R�FֆHdP��"O��@�Y�|�ޥ��lB/(�^iP�"O� q�o��<b:�R��9YB���"O�H� Ri��hC1LJ�G�t��"O!��#M�dih��d��"O�X�R"O�Q�i�S���K�	X�2�.az�"O�D*p��g.4�g�2�D5�!"OB=�¡ѧ]�zLr��)q��`K�"O��j��c�H�@�%ؑ-�"O`s��b�(d;a��̴Ua�"O�0�vl՛	� $RdL�=KE�m��"O ���d�8��%?�@�"OʔjE�PD0���і7����T"OL���#�${�DH�Ph�:}���@0"OLlu�O}�4��w	�Of(��"O�Q�Ĕ�"�kƏ�;��`�"O�4�P��Xj�q�J�xۣ"O����OG��0"�L��~T�Xғ"OFhQE��Y�8��fi_�1~t;�"O������[�"@��häU'"\i"O��YAH0E��9� �8U�l�"�"O��c��V{�EJC-ԇ(&���"OTՑB �$u���3L0X�S�"O��Ud�/t�XI�kCW&&m#�"O\��܏ˈ��iX.J�AI6"O��֣�1jPH�Tm���"�2&"O�ؓ
�R�%�W�����t"ODm��m̕<�e��oT#r�P��"OЀd#�#zt��R��<����'шa�'��\��tqDh�Um��'�pQ���Q;e8�@H8FîA�' ���e�.>&6�����?�� ��';�(Y��˘G���r�H�FV�	2	�'�0HUL@f��%��W
���	�'=�= �g[dnX)�I�C�#�'A�r���^t�%@�T;�lP�'C��83�
 ��i:�G*I�h��'9��a���n�0�A��L�@��'����1N��U88���BM#:����'\�La��-��<��DY_PL�	�'yt�ҵ �<MH`��L�n��i�דZ00b�?����"WǤE+EBS�dS�m����3,�!�$��[`��*$Kҋ @�����s�1O��ȧ���q�j�����I����B$M.uO��"T Htr!�$wJ�HyR��	_��9���jLMI��ȕ&4�IY�:���OJ��f�TX�@���%K����O($ㆦ��.8pWb�@p� ���H3m`�U`��t!���� I����2x�}��E�!~9�y2)3}�M�'A�|;��@ [�t@��olmH#f�C�N���ȓ[�)��5X���9���	�\$�������B$����[�O����D¬5�>y��/�px@��'b�ph�έYt$Aok~�"�&� ��Ȋ-O��a�9�3}�k�^D�@*�m �l�rXvK��x�K��-�]��N�y����*�{���2aZ7�$E�G�'�ޭC�R=f�H)�R�2@�ϓf�P�_Q�8H��'�*�뎱�x�p��G@ɉ�'��yQ��v#�tk0�P�8R�q��y"�P:W�e�v.P�O�(��'�)5�q��i�g���'�p�z@�'����әs5.]�uN���.�O,U���Y�� ,����_'0�Ԝ�(ԧk�&�JG"O
�bF�׬'}��K�%C7ߤM�`"O1��	�W� #�D�zV�E�$"O�\�rm/����$�$Lx�"O�])��<=���`���z?��0�"O��"�nj��v�������Sf�<���.S���NJ�P�S'��I�<��Q�N$����\1m������K�<��P�ZCZ�{��vU�I�g�Ql�<��ώk��)�՛QK&��`�<A-͊
�� �Ο/V��ٴɌI�<A�	�y������
�@tH���J�<�w�Q3F\V}�1ٍF8���A�B�<9�Y"Y�x=z�kEY}�9���~�<���U#:��q�v�Xq6h|f�v�<�s�q�x����ڈA�J�8�Eo����l�(Q���0|Ғa	��BɅ3��D  �j�<9��^�4��=�1�L��$����,aI�@+OL�T�O5D�1�1OPd�bɐ)��s𬃩u�����'�Tp��^=�� �1.	��J@���/Q2��s���1斄����9Ny�T���~�^u���I�ͬ�?��R�7��F�y�%ɱS?�UH��a�r�֬ܯI��)�o2D��3D�T���*TI�vz��	�<PK�'_$��᳌ɤO�#"�dy
FF�*��YwgF�<9�C����A4�.`� !���*T2���@�Or㥈�;LH��qO�)��.�JUQ�I��L��pIf�'��5��� �,g�4 ��V�]u�Lhh�=U0��J E�b��u'N�7�qOVb?yX��[ޔ�R���
#��2T�>��o|X���3 �k���~*��Ow���"kOP-��!����P/�	�KB�g�1��,8��2d{�lI&��=�8��'ʔ����Y<�v���
q�O�� �à�Xxl . ���礝U�>��IP[}h��IZ�⩚@e�,e��e���N��n�j}���3ǔh�O�\U���EͲa�O�y�N
U
�i��֗0 <���(?�O�m ��y�驅��7��Ssi���
�s�������4� �3Ӊ����a�O��]��/:H*T�T�4���Vd�h��I,��'l��q�n��.�h�q0)E��b���'��9�"���F��inF{,^P�6�r�)��/�
��$N	��'+ �J$��9���?5�S�?!�����$B���+H?�z�yC�7A�|B*A;�?�!�=1����J�����IZ%l�&>���4L�8��g�PpL)� �s�6@�69�6�(G�*}EP�@6j��rΨ�'�'�<�x���d��+���8l> u{��_0M���r�*�ݷ��%q�xӸy& ��<1Ǡ+�\�bG�$D
��]�'"��#�k�vVd$>ٙ1	��-����f$�1)2ޭ�7��ݟ���-�>hM�1�RC�+}���E�(D> ���dj��j@0��F� 2���(	�1�dB[����?	��ڛ2�Ǐ6fT�J�A� ���YA�V-��<dVC���-r�ys�$��q��k��+Δ��J��1�J�6k_�-)��ζlk�O�c�wcT��?7�ΑS҂*���	�a^�;�\�K�L�
BB�6���2!3��Պ���"'�c�ܒT�4���&Z+T�nx`0��5�>�Q��0OX��%cC�3n�c�H�6��	c�~�B.�ԣ�"O4u6&�/��qW�����2c�>��B9]!D��?% W �"��Ȑ���P��1ӆ@=D��U��[��9 �R�v�J��G�<D� �u#ν<<�뤆�6yW|U�:D�H��@D�#i@E���6D�ܪ��ۨO���
�-�Qs�5D�nm�6��|k��ȓ|jt�p�/D���P���#�����M�,�x��-�ܨ�p� �'4y2͒̒<��jwF nr��ȓ�r���î:���It� =`��ñ���E2�K>E��'X�9�d�"j.�YSd�;{��}��'����u�ĸ�t��Ճ#@,�I�_�B�CQ�Ǎ_?����Fa���G@�<ɨ������l؞�YM�0<����kӀ�1�E��{Dx�1K��BDZDH�"O� ��"�{��y�����<���d��UR%�Wg��Z9�"}Z#�΄N��J�iVY����(A�<�R��o����'�em&�rLP>.O����ώ)Lx�I1C�Q>�BlM#C-X�	�\��� "�F��ȓ P��)�2%��=ذ�	�p .�k ����3��a{R.V�u,�<`���0�s�X"�p=�_
���sH\��Mk�I���^%�J�8n��9��u�<�Q%��.:ܵ9R�|@F�
��s�!�B-��N�)_F|ى���	b�Z(�򊅞k���J3)��$!��EUj	
�c��t�2���n�6l@����:��l�>�|�'�5
hpx�
?u�ui�'xd����"v��i���j�B`��g-HR=Zǩ��0>��F�f�$��-͢0k���N`؞�ITƍ�c�����Ua���jXt��d�5H�,Y,���3�����[�WG��*��H(�}�'�Z���X:#�\l@׉LE�O�ey���|�@�̖�I0p�	�'CV�+�l�PɁ�ǭk!Z�zI<���WY�J��Ǔz�D��@�H�uG� ��6GL0,��I�*��V)�'�;-�N��"�֞sDLA�Ot٘�f �a�P�`vMRxU���	�;mhH�
�d�1���D�:)�ly#nFE�D"O!�5/�-V���sC2*���d�O�x���5�E�H�b>��D㑂^�j=8����c�b�'�]�@�A0�"Oh��W�muP[�&����Q �k��Q�b��D��D?��$��S�MиهL�J��"H��0\<��dL�_N!Ca�jFl��#,*���0��(T�FdF/>�ܸ�Q�!}r�ӵ~�����&]����"e�tE}r��"�I�e@J�'}!"���2Wd�"aK��T�'D�Da0�
�)�~\��II�&��
��^ (Η�)<0��0V�� �R� 0q��S��gTlP��I�0�,5Pt���cI1h�##O%{�#��8L���`6�3�ēi�`�#6#��q�9+���2D�O�	V5����Aڸ�NE��U��2K�4�jؠG
�I�Ɓ��ߗ{�q1��js������U��u�O?Ź'@R�#� ��d�N%�t|�a�Pk�<15�E�¥itC��V �+�J�my�&Q%$NM��/DjX�����֘3d��JY�����h5�O����U;lLd%@��W��i�,�R�^��c܂��x���Aa�13��Ϗ]k��+��¦��O��Ce�L>d�?�ӄ@�YB
�K'��@?�q&�*D� Q�Kr:�ДK�$e��K�̫�X��i�-YqO�>��lλAd�Lx �ϑ|�l5b��2D�X�V ��K[�}�Ӂ�>X����3D� ��#!�\2l�$,�B�Zf�:D���v�^�N@P�پ1tp��@7D���KZ7-8YaCԎ-�~|A� D�Dj���K�Qc��U��A�1�3D��X`MK	F�(� �)$\�i��1D��0���Oy�Xا-U2�f�as�,D�@IIʩ>b0	A ��B=�	+D�z$�^��	Ҫw�Ƒp�<D�!���&B���T��
p�e�4D�ѷa'N��Ԑ�Q�[炠��C2D���1c�w�����&�-b�iYF�2D�\1���i��4�r#�X�S�0D�@���N�R�n�4̉)@_� @�1D��{�o��"4<(����<������:D�d��[�S�8ze���Ylڭ@"�'D� ������ݪ'�ĥD��}�'�6D�H�2��(�81����#8�Yc�3D�IQǉ&X��)�lA��dm��#0D�`Z�M�f�ư�I=�D�Zv�/D�`QfM�k���1g�ڑ�J�s�.'D��c�l�8I�v(\�P�m)D���d����1�C\�.�ڀz2":D�� "��P��aF0(7���]v�B�"O�a��J�R^��K�C�F�c�"O�Q�
�?L�Ԉ��^�/M�a"O�2�,��\:�5������x�"O���'�Á��b`L	b�L���"O40�`J�*���a��� ����"O�Rf� :cM|�#�#�-I�@9A"O�]2׃_H� Hq��B���%�d�9E���� �T�n�u���1O�
gC*N�0��J�/�  ��"O��y�O��H|ekr#�u�Hq@V"O^��		o�Q9�b��� e�R"O��TFP��rT�}�"<q�"OAH��+���'/�]9J(H�"O�u���\Љb��T5dY�E"OȝX�֨>ҼE�c�V�1��4�&"O��u�Ͳ�J�;�萑E{"iq"O�;v
��tf����c�s�"O�S!?��W��+PV�D"�"ON�ɑNÙ(����>c�"d�"O�qJ�T*zY6- ���,a�z�(��'.�*׹i�h�a�	��&n@Q `A�	?�>�Ӌ{2��z��O�OĒ���n�S���Ӏ�t�%ǁ���3q�
�}���F�,.I2Wǁ 
.����3o�����Фst�'���I3,�`��!I;Q&F���ҜD\v5ˢ*V:��$\�Kru����l5��+�$�$�Q�j�2<��Q^�̚`fI*A���
ç.>"�r�܈
^��q�� ��=��mO���'W*���K��Q9U]�����]]LeY�Y���Sť��t�r
��u�dMc�OԨ��`���7Á/*�P;�a�j~�Oƃ_U2ĩf�Oj~m���L�7S��c�#H��f��(O�H�&�� �X��!��b>W�O��:K�e.`� #A+H�� G�'�V(Y&�B�	3�ڐd�>E��C��2����Ƅh�M7Ş��M@ƞ8Ԝ�M1	��{v�� 2$����D x6�u�Vi�R�\=M���I�!�gRR�̓����Oaz�]�{z@����^�p��$�	�'8�E�2$�#ۺa���d���	�'V$m؄i�A�衡�R�D�\���'&�E	V�悝����@!�P�'s@�C�Ή�s5"E!��	 k����'���)�끁lc~L�2��(j��i!�'4d9��K�e�iu��_h�	�'s���AL<�Z!��-�7J\���'��k��A�7*�M�ÁY �J�2	�'O�p���4F\$i!�E߰^�ε��'�����9>!��D��V���'O0�����!t$���]z �A�'�.e� .%1���'q
~E��'bl�`� �=�B\k��Z�!�{�'-\8x6M��(,���I1���)�'�LL��
�;���O��N���'՞9�	տ��̑��J9=m0��
����,	�%��K��_�44
NZ�yr�V����mƫB�RP�,A��yb.�+�0��4C
�8���	R���y�(J	m���S�\#'�6%1�*ϛ�y��9$�"���]�&Y�YQ���y.S+z�xq��#r�H2j���y�R-$LLxڅ`��f���$I$�y2�&Y�
-��R�\���Q��y�0m�v�`/cI�G`�)t�xy�ȓ:�l�)V��1V���딭ؤz��t�ȓa䰓�fF�k�����J����ȓP�*ܰ�Hϖ$�5dN�/Ҩ4�ȓb�Ē&#�EÜ��2FL�]]@���l���@��3Vh�[e�Z�>��?�@8е�oѲL��.S�e��S�? �@h�BT�pz5@�aN�KpH��"O�ic�iF�{KF��Q #s��C�"O�4�"���U-��rR쀃�"O�D��,��)u���.��c"O��P��O�UɺLq�GO's��'"O|�0�Q�M��u �e�]�h�� "Oʝ��4�n8U$ǣ[�ɫ "O�`�@U��n�2�bP���P�"Oڀ�Q��/��U��2<����Q"O�|jQG�!1~*��A[��V��"O��R�J�/ ���#!�Ry��"O�P1# ֍�3�1�(�`"Oе+Qx��Ҧ�V����"O4q�bT:
(1��� /�n\i&"O �J�bY�a�<S� I�J�4�"Oh��b^�A�(ha �{�=#�"O k�o˒SD�#�dO�T��@v"O�#��=@�m�De�"0PH:&*OȰZ�BD���Q�R���	�'��	�\�w�!�n��b%�@r
�'��p��O��m��`񩀆\%n��
�'���K$��$.�*��l� \����
�'��ũ��Ըp���`�܆A%l��'�\�`���&I�p��?*����'a��2G�طiQ�l��+�,p0X�3�'S����㖡t1��̎ur����'�fAi�����,ġg%
y��'����6L�p�ҥ�M5�R�'�ȝ��j0�2A�eE��
��'��<��f��+�B]�da�'yHX"�'
P2d�Y��C�,Y{)R�A�'=�����D�>�A��Pz� �
�'�ͺ�*ܟOg֭��;D�N̲	�'׌�X M���@ZQ�@*?�J0c	�'��
Ηa�h1�󡖊0���J
�'x���� E(�@�&@�� â1a�'�D��n1 ��a��� \-J�'�"�Ò�_��>	��/l�<�
�'�ʰ����jz�yƬ7"��'����L]-�j� ��©��<h�'�q2�)ا|�E
4F�g> 1c�'C�I��c؀��i�[�q�
l��'h��7�Q;HQ�a�˜Y�Rx��'�@�q���c9�b��]�"Ƹk�'�aY#�ġ/xd�"A̭+;0 ��' 6�Чg�8K4�t���)r@ɪ�'���#��̷��݃G�@�J�'d֝�a�V�"S���f ԾY���a	�'�:�f�.�0I�ŏ�P���	�'O���࢚8Ǆu ����wq��'8ԉPV<\�r�#Z�D�L��'],`�Ɖ�d�me͝�9D^���'�", �ԷYUT5qg�Z�/:�1`�'6��gׅII����뒑Bf�
�'��uI98Np��s���!Ep��
�'�H�1�1Z�����̘�c|F�
�'S��&ed������/^��R�'�H�B��:�ԨSm�%&�����'��� #�M�5���HR�Ƕy��'�^�#���!%Z�x��.�JH�J
�'[H�(G#בh�:��W"y�H0�',y;�C�%~��uh"�hT	p�'���!��C)z��J��+]�0��'�69�f���=��I�ǝPꐘ��S�? 2铤�'ʢ�ȵ��� �<�I%"O(h@ �ՠ �Τ�A��J���0"Ō
$�X�I�!&B~Gj�"O����Ή9�t��"J�T�A��"O�8Ʌ�I�<���!ćE,�Cw"O6�	p�^�x�ִ���L71�l§"OR��Gf�
k�̬��hT7d�
�C"O�pQ��\��l{���2O��̣�"O�cU��,�S����.Xx�"O�|��jD� �r���`)k�tyi"O�@����5f�y�S/���a�"O`I��l�(NS�E�
(2T�@"O|�! ��i�eQu!X�	ܨk�"O�^r�Pѣ\6b2�H��!�D�Z>m��Oơ�2����$!�d��F�ig��#c�5��"�K�!�!��\z$��>g҈9�q�é1�!�dޖnH�@AK7W#�p���^�!�
��̩�	΋nZE2�	*w�!�Dң,�P)i�eX��-���J']�!��;>��I
u
��{��#F��E�!�;4G�PQ�C�\`
�$�72�!�S6\|\�x�#"� ad-4V�!��ߐ2mFAbgĊ �v��FMM03T!�䂿X���8p��,k\�pa͉!E!�dЗX;��q� �;L��E
�&#!�dHB��Hyw�� �i���;a!�:oKT�`�@�G�a0�ȉ�cI!���h.���D��M+����a�D2!�dG�r{2�蔩ޓ*��0�֟|*!��-$~���펇&��q��͗.!�D�1S�8y`�
��L�r�_�]f!�Dx����/�T��1Ü� !�da�P��v��2�z"L8b�!�dZ�N��U���V�%+S�T6Y�!��Ƞ���hY�g�eCP̔�(�!��̋s,��z��K�M�@��F��PyҮȊO��1�c,�+4m괂��y����PĜ��V��-n��ԡ��yb X",��a�u����a�%L��yR�*C,�{AI�)p@���;�y2D���1Ӣ�՞4�Ʊ��(�#�y�� :¸�ԭ�ΐ�C,L6�y��);�񫡢�{~�0����yrHC�5 �r3�A�`��1���y˔����uMX��٠�y"�hpl�ː��a!؂F�>�y�I] *l�AC,Ə\ V 
��P��y���"��(r��׵Y�⨙��� �y��¢)��Po�Y�0B�̝3�y�ۮBs�kA��y\n�dDL�yb.@�Z����vfV�q��]��a �y���9e�T�I�d�v����6MЦ�y2%-d~ꨂ��L1Pd���۫�yb@
�T��`+dC�xߔi��e���y�
!Ԛ��uk�&s�TM[c�*�y�Om�P�(� ۬!�V�yA���y��W�c�j���%�E�.���oM(�y"dģ+dr��aÁ�̄c�I��y�eA�/��<�Vc�'�hY�]��y2b��!��T���	�xh�������y��&c�NE8�@ �r��U{�B˳�y�O֫D8�A�íkc>�Ɂ�D��yR�Ro']�&�D�rV�31��y
� $0v�@�T���SA.]C/Й��"O-c�6i�Jջĭ[(5�H��"OR����ϘQ�r�ѫ�6�D�F"O���4�K�k`����S1S����"O�`[f�C�?�@�	�,$����"OH�p�����(��a��J&"O��(���(B���t'@�EW�I�"O$��.@r���� �B���5"O���u��x�m�3D�[�"O�$"�a� jC����o�-\$X�"OĀ�tIT�Cv������`���"O�I��>4Jb�` ��m�|���"O��G@�r[|���	���y�"O8���Y�P���2 �_�*���"OT���D�QB�9�O,Os�"O�ȗ�V)Y�](�D�Y�Mj�"O�|�����Rp�)rS��WMır�"O� AVF 8�V��l?Z���"O�P2�ǌ'�6����'%�Q�"O�ɺ$�� 9�l@���D	��y�"On�!�O��^n<��f��=M��V"O�x��΄�Gǖ�!@�d��=Q"OؠYC�4F�v�#�dN?���0F"O��`�'U�N���ㆡ�@eb�"O2�Z������a��Ce�j�J2"O���+��j�By���,`�bp{�"O�C��e3��aw�%X�V	JR�6D��*4��z���IS�0�X�F4D�̰U.�*HNt���ܖ'��$�1D�li�l�)�$L���V�E>8�UA;D������]#>Lё+�,t��`�e-D��*bO�� ]�R�P�?H� c�(D��3�N߮���Q�2	�!6�!D��"��Q}��q3�p��|`P�<D��S���u4�Qa�"Gx����#9D�\�҅S�[���,*6n��T$8D��[�Э
d�z��Æp!h6�5D��0�N   ��   �  W  �  �  �)  $5  K@  7K  �V  b  ;m  >t  P}  y�  ��  �  V�  ��  ܣ  $�  u�  Ŷ  .�  ��  ��  Z�  ��  *�  m�  ��  1�  �  `�  g 8 
 , C% �, :3 }9 �? uA  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e�!�S�)�Z%����� �Z��I`n!�ͷ�JP)���4�H���,\��Z��(�*�-�pZ��N���V��YQ!򤈧6��r�7Lޘ�զ�]�$�O(L��fÇ�0�˴E>]��(�q"OR��х�=~�6l�F���
ٚ�"Ö��hY)F^L��!I�l�H��'G�����MP��SR&K!J� �L4D��xÊU�l���ᠪ�D�2�ے�2D���J�p=����ސ!�&���#=D��I�b�".ū掛�6�b�kf�r�����d�%��$h&��n˰E+��/�!�d�K�"H�&�%���s�'\q!�DؙX�^,p*��y�V��Şo!��0��(g�̏R�j�y�JA�e?!�D�-Qv��o=u*@�#�\�m>���)��Y9�һ/�����>ސ�a�;D���rfʣv6<X0�ڏZ�z�B͹<���2Z���y��ӂ+X�2������0HX���$��}it�u�$��TAζI�!���!����?@�hLB����2f!��7/���O
�/nZ�:e,L+�!򄎺o�~}��	=\G��aB�!�d��=SdIH!/M�E2ne��@�2�!��
�Aj�dqE���p=na!�b�#Z!�D���pu�$*L@�� #Y!�D��b����#21v �6���?�!��A Q~�y���*"�<����� �!�ʒr�X�Q����0�_�:�!�Ē<_����eb�
1�L� #�ׄ{�!�dTJ�D�٢5�y�ī��!�$�@h����*ZQ�s�ǩ>p!�$Y2:�~���Mf�W*�3_!�d��7VB�7�ݾ�*4��)�K]!�� v��d	�A� X�������"O���!H_!5�*�j���2��PKv"O�D���C�C�~,H�k"H]p�"Oܥ�Fe؋�P$`ū�	*��1"O�xX����J�I$	�"O"�ғ%�tQ�����mt"O~�4FO8P�=��@��l�Z@"O ��҃_	2fD	����������"O>�%*��TD�٘AiN9Hy\Ŋt"O���S��� {��H����"O���!!E�U�E��lΤ��"O�})uaZv�����y��8"O����!?��fO���1�"O����W�8����
���0"O�`A��Ch��#gk�:k���R"OFԑ���l7����CŪa�Pې"OF�I����B/�aZa�R����s�"O���eN@��U;�Mi �;V"O�eσrf�Y��"�	��E"Oȹz�m_�c,�����v���"OL�e�R.��Xa��a��M�s"OصJa��4xa�H1U�uj""OT[�d�ڈy�'�L�е"OZ=�Ҭ�kz�׻8J��#�ŞH�Q�0 �6\0J�{��݁gC剷!���;0mH�P��9�T�v�C��.nڨ)�K�'6��	B��ހp��C�ɳRox��ᐝL4�)���[pO�B�I�JK&a�[q�8�h��U�C�B�ɘY�$��o���=�����Pi�C䉢t��Е�]Gv��G��&w�C�I�P�\�cG�<'"���Q��
%�`B䉥9M$ Cb���}��D��^�%�$B䉪s�y�1
Ǫz$�aE�δ�B�I!�lP8�(
2~�e�&!�'gNB�q�>�@�@�:��������-��C�I9;)�Lq6�&( �4����9`�B�ɳ>������"^��(sLA��C�ɍl(�MyG�AA��"� �,®C�	
�8�ka[2la0�0PA�C�	q仂��;�J��E�A(�4B�Im�v���(���9)��ս-5hC�	-`��j����P$O�w���7"OB�:m�n�
7m�E�~�V"OVcv��+��
s�U�/��� "O�[mS=$6N��Ӏy����"O4HI�_4��i���Z�5�"OB5	�D<Y�~�+1bP)'P�y��"O��;�@�g�I���2c4~�p�"O؅�%i�_ΰe&�Kw���"O���� �f ���e�4�h �"O��2�ݼvW��bqEF^�>U"q"O�� *��q������uF"���"O�ay�Ӓ%�z]���ָ<@�0�b"OdE�*�q��5�.��A����"O^�r�JT��Dؘ�F
s���"O$��̩U5�p���`ihm�&"ON���ǅ�gV�1�C�E�8�2��`"OH��e��?���Zf�� _�p0�"Ov����->Jq�&,|��{�"O~��h~>}�&f��?���J�"O�I��\�"z�%����0����"O�������|�&��d1�A"O���F�`K��S��u�ٻ"O� �`�@dO�n���sȬX�ԥ)�"O���Ejɩ�9�@̇�*�(��""O��ZLƜg3x4a$�.*�Di2"OFu��Ü0�����k�h����"OHq�q!2�� 	q��K�V�[b�'���'��'a�'�R�'���'�������$e�� r����"R�'D��'|��'"�'s�'���'J�8
I��H�Q������P&�'���'R��'���'���'���'��Y�mֽN^zE�!n[IL��Y��'���'�B�'���'HB�'F"�'�����ث�ByT�]q��P�'1"�'�R�'�B�'�2�'Z��'?�a��m�&9H���"b�*��V�'��'���'"�'���'���'ʈCV
S!� ղ��F3��e�1�'�B�'Z��'��'�R�'���'���r�K] ~oxH�������E�'�"�'pb�'�R�'y��'���'���9%�#I=��R�&U�\��T�'��'���'��'���'���'�h�`Ŏ*=[IҴ<'�F\h��'Ob�'0R�'���'M��'�R�'A.�R
�-nt�ٱJGy��Q�'���'���'���'%��'s��'��e;�`���^����]�(9��'�'���'OR�'���'"�'Xh�^�E�h�#	�9y����'��'�R�'x��'R�"uӀ���O�̂�h3��J��
'|��X��Iy��'*�)�3?��i;`�5g��Hr��� S7���e����������?��<�����wə,#��i��@�������?��K��M��O����:H?qk䈟m ��s�$Dw� �6�Iş$�'�>��`[�w��^�h0;����M+6�YC̓��OQ�7=��X�u�X;b"`���՝�ݣg�O��`��է�O#�@�iN󄃡P�4]��A��bEP���JO��r� ��U	�=ͧ�?�Q��A�P�P���J����@�<,O(�Or9oڡ,�b����+I6^��`��m��8~���By�;~�I�`���<�Oh�J�D�� �-�����>���擟��	�hD �+�- �8hE�-@�|c�m�`��xQb��o�}���wy�S�x�)��<�W��">h|p�b
�=0�`�GA�<9B�i�Ը��O�po�Q��|a�6eg�d�`$�8~=T-yW���<Q��?I�v*��sش���|>j��;�Z�"AI�*��ñ-�%Z:Y�Q�5��<�'�?Y��?����?��	ҹu��;��0C��M�G�]��Ц9X�I�����	ş&?����_K�y���T;p(\�xd��X�K�m}��'���|�����:{e���ӂ2*�QH�q�����iK�	!Y|�I��OX�O�ʓK$�)p�^�c�0Q�s�����K����������˟��Ry�`a�����e�ON���))�2y$�ݡq�dH����Oεnf�Iɟ�!�O�D�O�B7I�t��_�b�@c��p�n���Fy�>�;,v�#��l��M~��;2U4�����i+� �[1z���?���?����?�����O9��[���
�ҹ��L�]|�1�S�p��.�M3�c��|B����&�|��4%G�E�a$U.���c)
=��'Nb���ë+i�֓�p�H�.x���fY	 ?�M�G�Ӭj�����'b��$�������'��',��k�
�\!�L�.A*���'O�^�@ �4r�R�a*O��D�|�2 �L��`2���hڑ���m~���>���?�L>�Oۆp��S��hň %T�+Ӝ��m��8Vp�q�i.�i>a��O��Oެ�愞�N�ܜ����-����O����OJ��O1�2˓*G�Ɓ�^�*��V��wQ�m��$]��X���'�r}�"�h	�O(�D�Y�L�d���O�ZXxQ`Y������O0E2e�c�t�W�ZY���3�5{N�J� w&d�Cׄ@�?Z��	iyR�'s�'�r�'��Q>���C��w�J9����~q�}z��3�M��n)�?����?�O~��ƛ�wJ��@H��_`��̑�/���'$B�|��$���.7�>O"<�c��#V-Ĺqq�\�Q�@�6O�8���ޛ�?��*�ľ<ͧ�?�al�=t}�Bc�N�$Z<���ē�?����?����XԦ�	�֟��	ǟ$��i�4ڴgT=��eYG�@�b��	՟4�ID�	)	�¤W�!e��!�o�<L��C��9�FK^��M+��4�V|?)��D��T!ļpS�Ć�s$X�a i�-�?����?����?�����O�|�SoN!����#(ŵs�bAy(�O��m��?X��	�@�ܴ���y�Ć�Yy��4�2�vi��� �y��'s��'��p��i��	��e�sП|�c�6�t�Ə
R�8'�>���<����?����?q��?���S�~y~X�JC���a+���$��P6J�ßT����8'?Q�	�+�j@ )R(գ�lW� �U�O���OړO1�
h�E��=d|�z�Ô~��YZ���L�^7m+?Qg��?'R6��o�	Ry��H�6-b'(��_"�,Z ��n`�'�2�'��O��I�M�	7�?AU���5�}`$)�-\e^�3��,�?�ųi��O^��'�b�'����1��b N4SdQ8�A֬L_�h�i3�	Y�2}�`�O�q�(�� �\�WOL4.����k�s�]�=O��$�O<���O��D�O��?�x�C���̠%`ҡ�Α�Cf̟@��ϟ�Z�4v�@�ϧ�?qջi��'���P+R(����jN4�9ן|�'.�O��p�i��i��� RTȰt�%_�j�2�Q��Z$y�Ʌ?�'�IƟH�	ܟ��Iw��x*�(2f��q� ��JV.����H�'�r7��{gN˓�?9/���$X�"y~��%ĪS��Q3T���Z�O��(�)R"O�o)����S:s&�V�%����L�*BO !q/O�I��?���4�dڷ%r����.`.����G������O��$�O��ɬ<I7�i��XB�˒f N1��F�[%ҙ� J��44�'�~6m$�����O��o�M�R���H-o�R1@V��O��d��)�63?�;`�z���'j��˓,�"X��(
7E��`mI-J�������O���OP�D�O���|
U� �,�#��L, @  ��Mi���L%p�����&?��I��M�;/��
F���d`
8��2xy����?	N>�|R'I(�M�'ԱH2��;�n\�'a��*�Ƀ�'��ٻ��e?N>q-O�	�OL��ͺb�fiR(�%E(1���O��D�O��D�<yr�ij��!��'�2�'=��gԅ\H,� �O��i�A�Fw}�'���|�dW�~�H�gY�
*����T���$ϲX�z �7�1��Z��2���Ė�m ��[��]犖�c�d��'Y��'uB�'��>���+&��#Sd�/m'���2DC8����7�M�4�¹�?���E�f�4����Z�_�Q���BNa��;O,���O8���J�d6� ?�U ���Ov��gHZ� �E�c�L�Ka� DJ�	]y�O���'E��'�d�0PF4��I 0�^mZ�L�A�I0�M� ��:�?1��?�O~��p��(��,h�m�W		 ��!�CY������$�b>�ӇD@x�T�#U��R����L<\�amZ��䐖_`����'��'��|#PP���$�X�����7���	П���ڟ��i>%�'Qj6�9�b��V�q��QE�+���p��=-�h�Ē����?Yp_���	���I�N�T��0�J%9;��!�T�\��FR妡�'Pz�p叓�?%�}��;lqT���) ���j2�Z��` ϓ�?���?���?q����O��鰤ԧW�]���Ť|U �@�'��'�6���3��O �o�h�I�5�~yZ�N���a� �-Q32]&�`�	����EnZx~Bi��_�h���ć�0�Ma��S�L���#A�VH?�K>�,O����O$�d�O
��n�GC�@q��ϔC���CԠ�Op��<��i�PM ��'�'��S~m�r�Qޅ;0�$�"@�>?!T[���I�$��'w�r����3A&:]�t�	wa`8bo�/4Cf����4����N�<�O�ԫ��1*�}��cV���jQ�O���O$���O1�fʓ%ٛf��:jx5iU�I"j�L�����<�n躁�'��eӺ㟜3�O\����R�} .ԼC�z%�%a\,<����O��J���Z�q���%O�r�OCr�1�A� }���m�n�D���'8���L��ǟ��IȟT�	`�Dj�w����'fǮ`R�ic��);��6M��b���$�O4�4�ӂ�Mϻw���b�ʥ2m|���+�4y��?9K>�|���'�M��'���8G�(O����K�ZF��'q4���N^?�J>Q/O����O�4!L�f�8Da��˿P�X���O��$�O����<�iqlH�e�'c2�'��@9�I^�'Tv�)���*W��A���B@}��'�|rML�&s���aJ�&I�ԑ��ȁ���䔦Z�����y��c>���O���B,'��5��±3V
C`�h���O����Op�d%�'�?��
T;qjR�ڱbR����aB��?�f�iD-�s�'A¨tӰ��]�y��ucE�Ȃd���-5?~��Iߟ���ӟ�p�.Uܦ��'O��K���?j��3��xrI��d�p����'��i>�I����I͟���"o��1M���m����~h�)�'a6�J��O���+�)�O���Q!�7��e�u��9��]��ꓼ?����Şg������:/l��ADF/*��<@1���M��O�t��@� �~�|rR�ȓ'FT4X��տ4æ �F�H��`����Ɵ��sy��OM:r�'ȶ��P�2-i�q3�"�w=�m���'tr6m,�I:����O����O�$`�@�%\�:����bI
=�Ph��&H7�4?!�dK!;P�Su���ߕ3v�T�{Av�	�fٰ#TXP��.p���	ߟ�����h����P�:�ʃ�0ɺ���`���a��?����?���'A���'�?Q��i3�'��œ&�-0]��`a��4u"�8�|b�'5�O�>����i$�I�q��p�:Fh"8-��W@h=����1<�$)��<A���?����?�!��Qjؑ��E�7K��$��?9���d�㦱�"M�����؟ �Ow$x���M(X�ՊŎ��(��Ou�'�r�';ɧ�)۲2�F��a^%���k����-�a�*Iv��<�'i��D	(��b�����̟�Sp��0��`v1���?����?��Ş����%RJ�c�t��Ć8%�d��c@�g�x�	���4��'���?هG�D�d����[�(�Z�ٷ���?Y��+2����4����е�M��N̙-O� ͸���,q� E97�Z�C�<Y('6O�˓�?���?)���?�����i1r��88r�V/��x��mE8梠o�)`���''����'��7=�Z���jT�/��k� W6=ˬ�j���O���/���M�P�86m~�����\s���òv�b�J�v�X�5c���<��<	��?Y�U�	X���F���eY���F�ɔ�?����?!�����ݦ�R�c�������x�G
����G�x� �W��֟4��O���O��O�Y�����RƋSJ��ɢ���K�ז\DtS3�FA�Ӓ]C��ӟ\R1OĶU*�ɚ��,i����Sc:D�5�X�d7���0-Q�]�ˏJ��DK��݁t	Q��I&�M���w�&<���f�H��"�7v��i�'qb�'*螓sz�星�!v����S�X�Ze	��Y&���F�ZT�����|�T�����p��Ɵ��	���Z�
�L�e�_#+F,aS�Ŗuy��qӚep��O����O�������;P��)��
�Dqɕ'^����'�"�'�ɧ�O��y�W�ƩRN�c�%F�6a���!��: j��dP��F�G�rJ�S�Ey�R	6|Jl�gD�.��qر!�����'"�'B�OU�	"�M�1痀�?y��P��>��0�m��$pcN9�?�e�i�OH|�':2^�������HvB6�eR��[
 ���l�_~�IE+o�F0�S* ��O��Ѷ$�� �"a�N��@��j��y��'&��'�B�'����A�R'P��cጀW&j�ڶo(B���O��d妝;�gh>�����M{H>�!dT$���d�D?+,d�d�[���?���|��Θ��M�Oj)ŉ.X�v�IS犱\ui�(��S���'V�'A�i>9��֟�I�A~$��ӧ<(��B�+�	ˈ�����4�'~6�9���$�O@����)ϫH+WoWl����gѕHN�D�O�y�'��'ɧ���'T�(h3�+A8�{������&�6t���i����?-�1�O��Ov�9�(��{��0�@��&R���Oqm�.�P9�%_�O[pu�&�?z�	`-�ҟ��	�Mӊ-�>��	W�{��J��,�Cၙ �"Ț���?I��J�M��OX��� P+���P����!�" 2h��F������j�,�'���'t��'���';�S)n ���'ҧ_Ĝ�A�)
>8iX|�ߴ$�J@���?���䧵?)���y'%�(�	���"S��qe-��'�ɧ�O�\�Q�i�DO!~�J013�B�r=lU�f�H2�$380�'��'�i>����9~�̙�O�O�y(��%v@���IΟ��	՟�'�7�X���D�OB扝*�dƄ�blD~^�,��OX���O�Oİ�c�>0���$1OcT�
q��(x��/B���J�(�؟�{V��D>��H6S|aS�L]��H��ğD�I�$G���'�&$�`�*""��6bUE�VU�#�'�7M��N�D�O�hlk�Ӽ[�c�0:�
&�A�onJ��c��<	����DV�]1~6�8?��f�u8��>N��1���,6��r�҂ig(̫N>�*O����O��D�O����O�љF�%a:)*��9c� �	Cc�<9e�iop��W�'�b�'��O�r���W��`X�'_;�B�h7b�$^�(꓌?Y����Şm�����̖�4U$@"p'B�^�D�#��(�M+R���#Z�1`�-�Ĭ<1�
�E�e�R�s����W$�?����o�d�i>�'�j7-D�_��V/(R��Û��L۠�|f����u�?a\�d��iy�����H��H\
F$��i6霻^�n����il���s�zI�g�O�'?q��'t@��FP>�:��;�z�I���X������W��X�~%�6Aܻ$�bu�g��(nsl0����?!�fZ�ƨ�����Z��'�쓄o�=>e>� r� > �lt�D D~�	���i>��ƎWߦ��u'jU�?2�i�.��6����uPJ �#�'��M%�$�'RB�'AB�'Ϩ�:3D��\���K��Z\P����'^R]��!�43������?������4e��aQ� ���d����������Oj�0��?�)!eH%Z�*�)(��e,ٝ|�d��O֦���T�s?)M>)�Iڟ(
�İ��F�go�2��ά�?���?���?�|�.O~�n� �� �.�p�� ���._�}
v�_ɟ��I��MӍ�>�����R�� k�q��"\�4~B�/O�����aӬ�ө�#JҌ��t!�2x֠�{3蒛y�X���_��^�Ixyr�'���'���'_"[>1�"�J(y� ��Ҍ+?2�$�=�M�\ �?A��?qN~J�Jꛞwn �sCcR<���9,�ұ����>H�B���=|F7�u�ĐhZD9���É�EK�e�w%n��A��p:�dd�	Xy�'a��G
!h`���0�4��g�߾- r�'@��']�I�M�0�Ў�?����?�7�B-V�d�Ǎ�u@6՛�ٹ��'����?	����j�=iAdΆ?�X
��E'P���'}�����t��֙�����īF�'�����΀b˪ĳ�G�����''2�'?��'��>A�I�SJDQ��D�N��(BI��<r���B�iU�����'q��u�\�杧	�}J�%^#C�"��,U�$����O�ʓ�>@cش��$����-q�'d�� �$�#�Y�NI�����##�2�°i ���<���?���?i���?���A�>-�	��O��1�B����dӦ=c��	ן���ݟ��z�9W�x��b�ۦv�P��5�IIH�������m�)�(ߚuJe�Ry@�j�ǖ�K�*���E�'{.��� \v?IJ>I(O�B�#\�T&��ꢪɉ�@
@�'w6�3��DL�0P"4��G�T��E� P���$Q���?�@Y��������	�e�d�#���-��9��O�u�~�����ڦ��'�%�EMYf�O~*��K0��cIù|�$����P�6�~���?����?i��?����Oj�J]�x��N�7D	r&��������4	�j�Χ�?Ѥ�i+�'�:(�S�K�L�I��փv���d�|��'l�OwF�Ʌ�iv�I�
����/�9��v��z���Z&�=���)�ļ<y��?���?Q�d�U7*�� �PzȐrBo��?�������z2F	��l�	͟�OF�=�ש��x+1X�@/�m�O��'�b�'�ɧ��2�`��,V.d=j"���Xq�ѫ2d9��2����d��*�l�1�@�P�Wݞ*p:ä�;���'Br�'���Q��zڴX^��[��@6�N
�6Pi�&��?i�/ڛ6�d�t}��'�`�S���6c���D��/	W*���'�bj
\��֒��W�X#(�q������0q;NuBw�C�	 �@��1O<ʓ�?���?����?�����;9j$8��,١??$\{pʁN8o�f.�-�	ğ�	k�SğL��������Z�"�"C��y�B,5��?����S�'|�@�޴�y"��(	 �qeC�8}{g��y��h����O�=�K>-O��O�a����"%2���%E�X�x���O��$�O��<Q��iݘ���'r�'�,��r�\ؚ�;�bL�kȫU��^C}r�'�R�|$Z7ܪ��!�< ���0b���d=x2TC� h��c>Q���O��$B�0�e��5��x���0����O,���O��S�O�
`�r�H���tY2(��&� r �r�dp:�n�O��$Vۦa�?�;p�����^e�����)Ul�a��?Q��?�b$�:�M��O `ʗ�F��GDK ^�0E���05��L�,\�cȶ�O���|���?���?��/��ã��\�=+A�&F���2(O�mZ��2!�������O����b��&���b1A�
8��F* �����Op�b>I�&�͗�`}P�!�&C"���'�	���hQ��Uyb�_�D(X�	�G�'-�ɧU%,���Ը���`g�4X���	ǟ��	��i>�'2�7m��?�4�DI�)H�H�s��pң�\���������?	�P����韐��!D_fq��@��F��x��HN[�
 8�J�ަ��'l�*0)�V2M~"�;*��1�4�^,��L�?1��͓�?a���?����?�����O�)�+J��p#���p��{�Q�D��5�M��H��|���#���|rM��+��E
� **l�x��γ��'��]������ͦ��'�T��!��Y����r�E69�2d!Q�y���	?/��'x���� �IП�	����@IY�ͨ�k�&Ү9�P���p�'��6�#���O��$�|���V�4%�'��� h�E���p~�f�>����?yH>�O�f1�bHܿg��E�_U1�um�*���U�i��i>�z��Oj�On����W&P볮s�.Q�+�O`���OH��O1�˓)��C�8D> ��爬e�z���R`h؝J��'svӠ�O��DPo}��'���B�(Y��x���@?����'�ҧލr:�����ݦ�|��@w�I�{�j�����+;A;2��j��My�'yB�'s��'�W>�y�D�"]r$��^z���ޒ�M[un�?����?�K~��[v��wqpU�_�$+.�/vfl���'�|����i�4O�1:����Z�?����~��?����'y�'��	ޟ���|���v1j%�ʍ�j��Yv�'7��'�R_�4`�4�2����?���f@��f Ih�å�:�ڡB�R��>���?�K>9��IT�ܳD�K������A~B��l�D͓ƣ� ��O�F��	f��z��DRb+:h��]"�)��y"%�h!g��+`=�pI��%H-bs�LLP,�O���W�M�?�;
D8��h("q���~�Γ�?!��?YV�A��Ms�O��
��p��A���Z%��w���䑢y� �K>�)O����Or���OH�D�O��H��OA�Q�H�A}���g�<���i��t��]���	`�ßX���?.�v�Zw�'��D��̂��$�On�$;��)ͭȳ\H9���p+Ph"�-�y� n�f~��ļ0y�]���䓽�D`���h&aD*+��*FZ�Q-`�$�O����O�4���"�����<��e:|�X,�ҏ(�6�ă)w[2�d��㟸b�O����O����Gm�	8�ȋ�����RN���؇Bu�*�J}��#b���>��ݸe�<�[�B�%�e0��L%��	�����ȟ��I�����E�'s�U��ND ��3b)�%�����?�:�������T�'6�/���>�8��
p����-^��p�O��$�O�I� U��7�)?�ab�O�? ��V�M�����^��  ��~��|BX��ӟ ���\��ܥ�R if`L�8��|�f�@����YyRb�Y(c��O����O$�'6~��@�+Јr>8���e�ځ�'x,��?a���S�D��>=���%uX�Ðʔ�E�0E�c plq�Q�擉|Wb�ZV���(a�N>q�u�1]�}���Iܟ��I��)�Ty-a�t�@��1����Kv&%�SNC�i ���O�eme��2P���� j�Ϗ��QW�w���FPy�e��{<�������"�3p�D�@by��ٳ5��$�ufA[���+���yb_�H�	����	���	����O�0J�`ܞk��H�i�36$,J!kdӚ�[a��O:�D�O��8�d�Ʀ�{
�k����8�\�o��8�F �I�h'�b>�˷�ɦq�A6��R�G����q�P�/�d�d�hP�dK�O��J>�,O�i�OҌY2��'u�u
�%#b�L0A0C�O��$�O���<!�i1� �B\������(�2��X�B�H(4׭$J��?QT���IZ��>� �����=%t��r�S�ڴY�'zJ0A�
hV�}KU����N˟hK��'�v���?>���G�FL=D�u�' ��'���'��>��	=6U�p���>"����UKܨ|��		�M��얾�?	��4e�f�4�� q%��Xۋ� ��)�e��y��'�"�'"��ʠ�io�ɼxR�YQ �O�pj�HB�G��;�E�~%���FKg��Ty�O���'J��'�jՠ ���(1c�)[��a�D$(��I��M�бM��㟀��N��\b0C[5 5j(:`�Ԓ	���������D�O�$/��IED��a���&����Rc�1ː�jq�j�'��Y�E�N?aL>�*O�m� 'ٗ�����d	9�Z$����O��$�O
�$�O��<���i��HHd�'�Rq�УI�,E)"�UL �`f�'��6�"�I���D�OX���Ot�F��
��щ��&~R���8+4&6-'?A���.���Sr���a�``��n�r���C�8s.P+�$w�<�I��T��័�I������<�q�`D?���2EH��?����?aB�i�H�O~�)`ӈ�OV��Q��h�轂!P=A�@ta�d4�$�O@�4���klp�\�U~���@�u��P���	}u�p�H	�Kl�$�����4�����Ol����m�$,�:rr��*�d�O�˓fl�VF���2�'��_>	 b��Zd|��QL�A^d��D;?IeS����h�S�	Y�E�DjEjhy6����_<���+�)[�v�yS�擭%��^�I,Z�Q£��d�z�Pw�7�����`��՟��i>Q�ɮ���'�07m[�2��i�ILqM��S&��]^�M����O��d�Φ���py2�'�r꓁?Q��=BVqaD�\*&D����?���z$iٴ�y��'��H�Z���	z~R��9�~I���' l���!t��'i��'l��'���'3���L賋��Y̎KrDV�c�. ٴu�u����?	���'�?���y��ÈIp	C�9c2���K8��'4ɧ�O􂐐R�i��DV4�,q0 �-�@ī��kR}h�A�H�OX�S��AX�z� �$�p�A�)ʣ�0<���i*�pyP�'�b�'��(�$S*�4E���ĄLr�x t��]R}�'M��|��s 8c�NG1k*����'��D��B֌!(��|�"I%?YK�O6�dZ�w0:�(��2�Tӳ�hv!�DK�v��`��� q���K����.|���ͦ]r`
������1�M��wӈ�ɀdďPc�l�3ΐ>n��
�'�2�'���V�x��f���(z�����8�hRB��c����!ӵ��bu�|�Q�Gr�H���Y��7��0�σ��d��{0����I��:�U+0�j���T�bW��ӣ+W.]D�I���	^�)��(��CBK���b�*�uKt�� *OR�����~��|�\�����T���ԻeS(6���e6�O6Io�<d���5^y�H�(�4q	j�6�:�:]�I$�M��� �>��?��~CE:�-���4�GDT�@)��M�O��]����o"�)��2���o��P�����	�0M ԪQ1O��dZ�\QXE2�oE�Z�|���E�Ic����ON���̦�GK,��i<�'B�7jH�>�2�C�O��sn=��|��'3�O��l�ӽi��	�PF���f� c_"0Xq��. ���:Ld��(��<!��/;ڂ�!�k�/k�@�[��O�oڪ/�2x�I�IL�ԫ��^��#�Ȱ3Pr�E�����S}B�'=�|ʟ��B�ɂ�@`�ٰ��>���AL,i���(`��.e���|�CC�O���I>1�*T��\�"lY!��T�ס�X<�4�i���2�/�e"�����W����2ҧs�2�'-�7�5�	,��d�O��Q��J	�J̳ǫM��������O���(F��7�5?�RN����fy�&BAb601F=[Y��R�=�yrV�`��I(9�XX%��f��{"�ʞQ*>m��4�J����?����O�T7=�޴zDd�4o�����{��u�$��Ov�D;��ɔ)]��6�w�� �#'�HH^�p�ȋB7��@�=O�T��e��~�|�Y����ӟ8���F^��$IA�
��\�P�o韈��؟<�I@y�r�VљSE�<A�V��ex�Q2L��[�h�P�y��d�>y��?�K>�����6	�;E~Y���F�U~b��%%��40Եik.��*9I�'^�ҁ�����]�^-p���)	��'�2�'�R�ҟV47 �����-� �x���+C���OP@:��'m"-s�T��]�8�n��1��8xxT�P Jk����O����OڜɃ�r�d�� �D�?!���F$��|" ���sGLP�IPy�'�B�'��'�K��
Ja[P�O:�ljQ�ŵ1��ɏ�M���?���?H~���"� r�惦z�I:g&B�)�´�6\����ٟD%�b>a�p^?/�F�Rp�MR�������ަqR/O���E�E �~2�|�R�0����,�Kge�}�<�*������	��`�	��Vy"�z�0)З�O�A��ΞV'X���)���%�O��m�k�={��՟��i�UA�ɓ;w�!�pnJ��r����t%�mo~�F\0.A�y���A �OQ�O)6xq��'4$��y�r�J��y��'0b�'��'W��I�k<,*V�I�&,) �X<ڔ���O����ɦAz�c{>U��0�McM>����I�T4���3�<��������?���|�'�L��M�O���^�X|B$�H�6��e�֮ײ)FyhEi�O��"I>I-OJ���OB���O�E���O�de����.تB� 0ʔ��Ob��<��i�>�qS�'r��'��*wx�2K˿t��Ӱ�FP��ӟ��O��d�O��O���� ��D�0=���IV�·3
�Z�B��!ѓhLy�OlX�u�M�K>��_5%���'�X�U�q�G�Q"�?!��?����?�|�/O�o�X<Y��OQ9*7B�r��I'$%�@����䟼�	��M�L>!�[��	� �tz��JÇ��z�4��ȟ(�	4S���o�T~�D��}�������$_" ���@��vPV!!���� ,�k��9[�)���h��hCԴUBhSTB��bx&�����<$|=+�DN#h�UKE"ՒnF�ysA��.W�b<����:J$�!�G��p=!���WwTq���%s�tYfF�*���5���v�'ϕ�VL>��i�C_��p�+o��˅eA�>���C��(XQ2 �϶2 �!q�'�d1��"�<�C�C{������ �r��ʸ.8fD��-�4��3*���ݺ:��U�ſD't���� ^̛�'��8O�D�>�-O���K�m�Vɠ5d 0ur���S/�¦Y�����D%�����e"�Lr7��)2�A��r$X<Y�i�r�')�D�'�����O@��7 9xAJD�)-~x��ZB�1�B���n禒O����O>��;����"�`��r�Ja��l��<1F����D�<������#ե�0�쵣t'LO��b��b}�Y�
iR����ٟD�IHyR ���b��!R]$B���C�534�0�aC�>	)Oj��"���Oh�d�2vz	�0�fp��h�$R�A0��Orʓ�?9���?�)Ou�3���|�4��4�T�s�C�\���W����͗'�2�|R�'��'N�z�bjډx��1S%H�h�|Q�/W�����?���?I-O�8�M�Q���'��j"hF�A�vc�����b'$h��$>�d�O�d
4���t�˕3\�0}� dΪ5H�c�Ge� ���O��ed���Z?���<��'W��w��5�4,�RG���P
J<Q��?1�M��?	L>��Oj�m��
ۑN�@p�/�{
�H��4��d V�\�o���x���<������<u��H���8���2?O���װi���'�"\���#�S��,tZu/C8k��`���ƘE�7��g�~hl�(���<��y�\�x����	d�(��0���`1f�:�M#��A��'���$U}V�{1��&\񦱢��
����n�ş����<1�%����<����~�C�Tʝ#Q�D�G&�{�gX��' �Aw�|��'��'TR�R�J
�H::��Mіii ����g�P�ɴ__"$�'�����$�֘�K�~$p���k(�[���8]� �IptxK>a��?�����V;K~l5r��ͅ����U*[�֕��ǋc�꟬�IW��jyZw�H1��(��rqa��O$܁�4�?	.O��d�O���<��DȄO���J81�$yr�k<}�Ɛ�n,�������~�ky�Ot�d�Y#����dٲ�c���O��$�<�Ee��(+���"rb�a*T-z��$��[��Im|��?�/Oz�	�x�A/�Tqauc�=�B\����M����?�+O���2��A�՟��s�]`����)=,̐1�׳\���A�(�D�<����?�H~�Ӻ3%�>h�D`��5!��
u�@t}2�'��!�'42�'4�Os�i��S��0=�8�QE��N�(�!�w� ��<!�&p��ħI�D9�5��d��33
�X��n&.�����4�?	���?��X����ц�hdJ�,JC�3�G�x�@7�O���O��O�3?AEcU�m���� ��K�����j׃vi���'�R�'f�s�^��'��Ɏ�����(j�M�LC�-<ӎ�\X�'�?��'�X1�FI5Q�`�cB�-~��M�ߴ�?)�C_���$|�D��_��L�$��4 �K�,ݼT��H'��`�&�I���'u"	!� �(���z<�y# �W��{AL�"���OZ��-�	럼��v�F��0{�P��B�d�dun����?���?q)OT�)I��|򡈛�G�u���ɰm�佐�)�f}"�'�|2]���ݟ��A͊�'�����@�e�����*϶���?�(O��$*!�ʧ�?�D v�z��O�Y�T�0��K7!����d�OX�&(�0'�|���8���'�� �J�t���D�<�� ?.pP.���$�O����Z����'2��æb�qhdUkךx��'��I3Z��"<�;"�p����P*V�C���/N��m�zy��f�6��\�t�'���a+?��N�b�� ���s�����_צѕ'v��'Ӻ�쒟���N;l�E26�
iW�I���M�� 
:ś�'S�'����8�4��a��P[.|��!R:��%)���Ϧm�IΟ��I{�)�'��@���.բm#��e�$ӥ�c�����OR�d�@�v�S�$�>�%�̳uh6��w(�.c>�*��=&m��HH|���?��3�r���Ėr�����fJ2�u�i"�i&P��O��O��OB����,7Q0��6�U�y� (Зp������'���'��S�|�-�d����2mJ�/dy@��;�`PN<���?9H>�(O�W�Z�����F�#�8B���e���'��'�2\���	�|,�'J��9)�P�bB�E���\�v�oZ� ��a���?9,O�%X��iw24�d�=`�T�5�هj �B�O����O��d�<і�Ő^����0�D�d�(`g��O�I��$ũ�M+����d�OL���O��C�1O�ʧ޵˕`z6)�f	J�`]�H��i���'��	(M��EQ�����O��)U�{B�`5��1�\3&@�klB��'42�'��#����D�<�O�:\)�g�S��8�&������4���%(��o��x�I���������2�A�(n�����2�i5��'�<�'ErS���}ґ�T�f�����;�Dpc�C�cQ��%�M���?����r�^���'p��Vi̵}��]SǊ@갍ٰ�q�q�p<O���O&��2������K��1llIЄ瑥��[��M��Mk��?��x��Q�H�'w�^���ҎW�$�~�1p@�:M�pX��i\�'��ġ�����O��d�O��##PfOB Ŏ�/�m0�Ʀ�I�Y�8*�On��?�,Ol���B�*��R
'��A�D�_ ��S�U� ��w���'���'n�[�Th�B�4Ad�����@5��d:�#Vf��O�˓�?�)O���O�����ԅhP�H�u�,D��R�w|$��;O���?����?y*O�������|�ƣ�0t����3���D��˦�'m�Q��	ݟ��I�u��I�a�4U�'O�4s�(is�I�2|���O����O2�$�<3��Qn�S�P�W�X�X��䈗/K�cORl�BOܪ�Mc���D�OT���O�1�5O2�'���HՂ�4@ȶU��EU�~|�ݴ�?I����J3[ך��O�'��T#>l�<[3/KQt� o�IcP��?����?��N�<�/���?EAC�^�Kt�5��~� uӊ�6�d��i��'��O�~�Ӻ��aדaJظ�왡ۼ��P�����I۟8b� s�,'�0�}�C
ˠCʸ8��!̎�0 -�E�����M���?������R��'`a���R
	*��s�Ύf]>l�u&{����4O �O��?y�	K5�U7��0bs\9�→M� `x�4�?Q���?��Pp,��py2�'��d�/N�L�7.U�=��c&��-�	~yb]#��4�0�$�O ���%�|T�#C�d�<�`m�k�H�o�ϟh�P(�����<������Ok�L���I�,�&^7N�hE��U���6<������ǟ�����8�'��u���_�)8���G��-�vp25�4O�����D�O@˓�?y���?�0���3,&�s3+J�?�Լi��	�0�r��'}B�'H��'o�I�,%:�O����4lA��8�jU;]!��ܴ��d�O���?a��?9�J��<��IH����h���U����%/x���'�"�'�U�tA�·����O|�BbD�j��Y`3�U�N[ �y�ڦ	�	{y�')2�'��z���4.�"Q��׃M�tq�M�x�}m�<��nyҀEHy.��?����
DI�^Zr��a"яw=�Q�����R��ϟ��I֟p���`���y"ӟ~iÃ%�FX�+�2?6轒��iy�ɱ E���ٴ�?����?��'+6�i��FfY
~D= ��G*`|�r�e�����O���4O,���y���ճ+�r,IR���"���Ta�?Z-���%�L7m�O(���O�	Li}�Y��aԠ)6��8�t$ˋ>��(@KS��M+����<9��D�'�ؼ8�ḍXj�ij�C�S�е�"e���d�Or�ė�P���$������$��V,�HҒ,�,k`�Б�C �Al�Y�CIt�H|
���?y�1��|�*w�<�R��C*v����Y�rM�4^�OF���O�Ok�
,(��#$��*�B�@�E\j-��"lG���{yR�'�B�'��	��pIq��$By`9�����
��W+���ē�?q�����?y�5��h��T��U��,ŋ]y�ES�.� ���?����?I-O&]�M��|�T�һO,�%H��6^)Tp9&�s}��'��|��'B@ӹ�y"�݃�BE�0�)ʄ5I�ˀd����?���?,O�q3EDp�өЀ �X�i�:"�fmѰ)L> N�}�r�i�R�|R�'�b��y�>��$כj����1Gˠ=��1��
�������l�'&�K�-�)�O��)՛m}*ɱ��Թf��ˍW}�%��IןQA��埔&���4�:�pa�r�� �ta�>vogy��6s66��q���'��#?�	�B]��¢[>
 ��s#Ħ��	؟ȋ b�&�d�}�Ă�E�r��[F�!ꄅ���ና�%�M���?���bs�$��p����S�	�h�f�ͷUf8oڣ?�0�IU�[�'�?��C��m��a�U�vCX� �
58ϛf�'!��'�髆�9�Iڟd�,׮ٻr	N�;&�X �ے@��AnZu��P�H��L|����?��k�����
]= ���a�
4c���%�i2���]�0b���Ie�i�]�ԋ�6�� ��˴0@�V���D�����d�<����?���'WZ�H�rⲹR�����D���a쓁?�M>���?g�R�&&��@Ί��"��M�Y�fϓ����O����O8���O���-�O����ŞY��(!�X�l�`y�@��	֟��	G�I֟��'�v���4}Xr�q&/ܡz��,��/ɜZ�fP�'���'`"S�$;4�(��	�Op����E�U���Rum|�EO_<����'���$�OL��pAgʎw�&QVk�3��K��w�d�D�Oh�d�O�U(���O��$�O��$��LY�	�>[�$A '$��y�,[pK�Q�	쟰�'�$����Z@xq��Qb6�R�B�*e��Q�\���I�imT�	ɟ��I�$�S埔�'Oh:�	��V�G� 	xejM�k-�Hn�Ж'�������D��E+rQ%ăi�f�I��ϼ�M[�>!��'s"�'c�DH$�� E�Y�Ӯ�	�R	uiS�6[�=�	��?�2�2	]�Pt��6��x��_�?���'���'����qh!�$�O������cFD5Dt�J3f�I�hYA�%�I�4�Zc�d�	ʟ��I����VN$t�cd�. �^��ش�?I���. ���^y��'��ޟ�X�yt� �$L��t�\SA)J H���%݈ϓ�?I��?i��?�,O�I�-;_�� ���uyR���4��}K�^���'�W����ӟ$�I&KE��80�ͥ.����h�)�7f �IП��IߟX�'��s$�>�`�M��̙X�N߳��ř��}Ӷ��?y/O����O��4g?�P䐥`�1Q�ԳƁY�y��aoZʟ���՟$��uy2�V(����?�1눴��E�S`� ��)@B�nZɟ��'��'$��>�yB^�i%�K)ԑ@��� ��$W��M[��?�)OV����Te���'m2�O^,łS@�,˄��l�+�,y1dD�>Q���?���M1>�͓��9O���C{�(��3N���T Q<_#�6M�<9Fꖦe��V�'r�'�4�>�;DݬE�T�o\����	G�l�������%��	���9O�>���&?'��[�	D�Fb<@���c�Ω��OЦ}��ڟ����?I�O��+YEr��W�8�(�U�Z�%-���i�����'���ߟ4�����H×l�5[9��PT�
>al&��D�i���'���26l.���d�O��	\�����R��)���$�d7��O��d�O��ɰ4O�S���	���{6�Z"M����,
%�^�i��4�?�%�F$��Ty��'[��ԟ��}j$��/���)/v7��O��a�4OP���O(,��L����'5\ ��-��pb�����.��1 �"OX�3Ŧ�""���3RHZ���#��I�Sn<
�Ȋ�'�����ѻJ�~���'S�3�VЉ��:7LhDX&gռ�J5�2��~���ӃD�knn��q*V�ڙ�"��O����g��a��,�Vcź)7�A�%B���<�e/�d�ȉ{3��B�)���V��h�F
��n1$���C���Zӆ�$`�ak����P��|** �@�֜"7���X�3��9� �d�O����W*-� ȏ�P�<C�`ت$`�O<��*W��5��隷��U���R���U0?UzD+�$��
Y�T&y���LA��%DeC�B� 6(4�V�8�>�`#���ԟT�:��4�����0HN !xq'T�<Q��>��r#��4?ˠ���3����I��ēt)rx���56���p������Y�6!J,j�S���i�D���2�'���La�hA�J2c���Ӷ�R%Zl�em�
d�H�[L�e}*�\c>��� r�'��<,װ4�elM)4�^Lb ܺL�P£)�����O�U��O�o{���Ӭ�{���M�/д���O��S��~�hђ���ҥ-�1�4E�fC�I t)�1;�m�e��i�PCP#<���)zFA�&z��L�I��=�]�?���j�������?1���?)�I!�n�Ol��!�aR�e��"ʜ"�D����gӐ�Q!��
�0pk������۞~�A����.:�
}3�=5fq�	0}��P��L]� �U2�՟ў|I���&B�I�q�fZ��q*��,	�L�O���!���d�D�ݣt��Hc�a�k/!�䇣�^p� �Q�F��\j��Ӓ#F��Ezʟ,������i9��m��@3dh�%J$��'�B�'�R�=�'$r(K
9�T0�3��� ��qG��I�*[.��Q�
�O�ĤRf�?M�(� �tXg��Oef����$^�~��T�!�O&����'�ԩ>�
��:#r �M!V��'��'��'�OD���D�Pw� �p�0XZ9{�'�h�J����%�@dS�*�',=��И'�6��O�˓ S���?������84V��4#׊W�\�A�(>�J�G��Oh���O̣0kv�$��'i����_�_@��a���>�f�DyRj�.L�ʄ��:kp0��,������
���<�AI������̟��	A��# >Vxm@ H�E�8��ԅQ5v'���s��`c(u�ڬ�RKOY^� {��5�O�5%��‌�,��P��E�6��gs�$��cI%���O�'RH	���?���V<,�Dd�g��'l�b�.����w0�EЃ �g�T>5�|�	�?f,1*^/�i#@IA�c�Paq�Ky�DوA�2}���'���P$?i���`�
�K@�A	�!O���'�"�'?��:򺨸�G��={v壧GX�>���O���$��)�BB��er�<0�_�+2�P��D�|�����T��#� ۞�`�����x�m��,!��cHۀo�ؽ��(��yRi���N�i*EXt��!Ő�y"���"ڀ���H	z�H	��KX&�yr	��H�:�;3�֡i�|�3tώ3�yr��%[�5���4e���Ώ��ybK�.L0����e��-nD@��'g\�(7�U;=��-���v�x���'�P�*�(G�hXp�k���+|�Lmh�'����D��]��«�ڦm�'XnPم(4gIJ�b��H�Gk���'�nQ8a̕BHi�/��-"�'O���h	VlT�����=(�����'N9Sb��Q�j����6�`9[�'c�u���%��=*��^�3,���'��q4�5dV��ᘟ&��8�'u���47Mt�2���05��1�'QHAiF!��$�h-*�`B�4��� 
�'�@}3�m�(f�>�C�рC�DA�'A�@�C�
z���r��
J��m��'W*`j���	CWe߯G�N�X	�'��eH$�Di����կդB���8�'�4IQFMQ#b���B�3'xUY
�'�6DK�-�4
x-��NN�Bݰ�y�͈�y�4����Z{��y���-INH�5|�<�+P��,�y�`�0GT	R1�>x�(a���	�yBfX�S���a��[}���Wk	��y2ԥ1 �bPI�<ZҰłG�9�y��*��$#� VrAAv��#�y"�O�����]G9be���Ӱ�y"� J#\m��/ŗ<��U8�F�yr��A*(��U·�T��׈4�y2���4�,�c!/��!���?�yb(.g���Ua�ud���Z��yA�j�p�9�
��� Ү�y�31M+�N�x��vᑎ�y�����(Y!F̕�8z�n	��y�!C�!=(Q"\!w:V��i���y2 �'|b�i�� �(LԢUi��y�(1A���㈚��q3u.���y�'ↄ 4�ߔ���*4
��y�/ï3��YrWL�9x�yj � ��y�p�Ȕ��i��C�! �F%�y�HզR���4J3K��0�6���yB*���C%�	2״�����'x��A+7᲼����mpD�K�'0*�����Hz�;!��=_���Z�'��T�0�j.����yE�0�F"O� �1
Ys5V�`�@] B�=�"O:�Y�]�^��(���)I'L}`�"O��[��,�t��$ћ
}H�"O8"�`�^��9(�	]�Mr�)�2"O�0Ydk�>�*���(Afl�1V"O���$FX4iy�upua�C��`
F"Oz SQnҒ��83�`���kP"O�t�����s(�Aч`�PTܢ�"O�Mi�'�#�H8�QܛO �ak�"O�d�DH��8T��	Ge�(�"ONs��+F~BA�_�1Jh��c"O���YKp����&�"0>���"Or�тOӟRE PFa����"O�=X���u�.	�W��l�$���"OnYi�CA�ܰx�M� (oNh�g"O���b�EZ��9`MS<TJ8T"O2X�g��,2�h�J�%3�b��"O*H
w����@�Cʟ a��q�"O�ؙq�}L��ˆB�&q�Ĳ�"O(��Í�٨%`���&xD�h"OH��5\�n)�E��^8%��"O��Hת=2&���aT�d�Dw"O@�R����
}����2u�́�"O�f��B�p`�A�q�,���'�P�E�Z��i�CQ\�p���=l�JB�	=�8�3�	ޒ2���2�B^�AM�c��rpB_p}B靋J����~�����@8�x�a��B��)�`XD�<�eH�N�葡)اg�̭9���D�I�.�޴g6J�F��O��4gT;I���甔_ɨ�{a�'�~$�敉ca�S��]�C�`Es�ӎkZ1��F�!J�{�Fg :�������<1�n�*[�XD��,�4���7hK�'~`e�͎6:���@ ̼)��O$�H7�K�R H=��_�(���c�A��p���k��Ձ�p>Q���x�@)eZ�4R�N %�z�����1.�� )W(�S�2N x	c�A+aR�N ¼{t/@ <�vu#�]R]��s"�{�<�ī��^�,��M� j�jDh2d��+|JY�7l� �D-���_�B����D�����O�(��Ѡa��nD��$��C�
-{����a|R`�3]������1ے)
(Kf-r
� [�����IQ2�1�h�g���
�-̎uBH0ؔ%�O�9��M�"u��Ҧ�x���	/u"L1���%�1�@��-ɨ�S%F�'�T" ��U�$P��BŷE�@�H%OM��N�&D���د`�*��ӨZ< `ȸ@�[7ny����[E*����k�<t����� F*��נJ8(p����Z5jq�T�s�q!�i�;y�T�G�_�.c!�$��wzJY�r"��#���)͉/��Y{���<�4��T�>Q���V��Ja��	��@�'zf�j� ��(>��QAo=A����'��l"�/X5{��3� �et��R�Ǎb�"$��K��5"b�R@˓E���+R'R�-<��X�B����	G�Q����dߊ(Rց�<��lϪh�ր�%,Z88�5�@�*�v�'���抛�a���2Q)�%
�[�l(<q6l�v#�L�XJ*p��E�\b�9�h�QĦi������>�'b9�qͻ$�1##ܛg�`L��B�\Q�ȓ=����e�PѢ���	7n	�?!$��!��PE�(q �Da�Y��Y�y�y����Y&�𺷡Z({�z2`��a<�l��'�f�sWM�+^q�1O�jhH:�C87U��V�'[sੂn��s�����$^�u��0iv<���_%�qO��ç� ! �!�f�ì`���J��|䔽Q�MX���]�X BՍ[�N؅�A�LHsTs	� ;��
;G�����ۤt�@d3���C���q �?�C�w��Di�a��cb �B5�Zh5<� �'�^`Rd�ʁp��0�&&'0Q����d]z�Na�4>��X;��X�1O�,�BMѹO��*�Ȏ�WP�h5�'��5���W�)�p��,�/<��HX�HI�uo��1 �PN���gb����X�H[��͆�	�5����u���p5pǉd��#<����� a��aj�(4�M~�fB��B����:R�6E+ 	��c�&��'�VI��LM��T���V�
$�S�`�?���� �\%[�ht�TH�����9�(%�@d]/aE�HA"b'u)�t��"OZd��MZ4���1Isj��Q�Ux_qO��*�OR2��Q�X�	"��Q�_��P�>Wp +������pQ�8�O,�h��U�#�$U�� �s��O�o3�H��A�j5"��'���2+��I��@�R+�-�p<�wČ�yzMs6�Q�=�2͢�H�'�ڀ�s̜�A�zLq2�A�}2̠/O�\@&�ݔd�@�q5���9x�
<4�T��#����pG'��sӖ(c�m�v�`t*�Wn�e2wf�C�,��&e�>�}�1 q�v��:"`�GJ]�E��5��y_J�� O�b�RH�Ɵ��ऒ�d�����\���S^J�T�Njܓ����N�ΐP3�������I(#}��
��N1V�xZw�ֆv���3ψ#A�|a#��5W�~��,�X�Ih�y:�����	 ��Գ�'�8y�F�N��A����G�	&���"��� �H� F�\��!��Y�m�����jT\A#l��Z���� \u UѤ�8%�|�������z��'$�
!�M9�<)d��S�jB�	�� �Щ_�S&�0 F朾:��94(�K��	rg��+ ݁a�]D}��_�I:����.��~^yt"��p<I�Ǜ�,Rj�~�Lc&��k�pGD���ZL��q�b8�B'�O�9Q�S�(�� 0 �"+��
g�x�@E+@^�O��8Ȑ��Ou��7�W�Y,�L�0 �bhb�
�'�h�a�4p�<h�%���U�
�'ІP2�J�V pA	t��D�h�#	�'ߔl����N��h��L(?d(��'��19@�"�J��qƔ16�4]��'@��� n�)X2�	�mD�d�`�'�����I^�/�,��W#�U�XD��'U��a��{)*%@�Ē.zy#�'�0`⣤� �~Y�F��e���b
�'�6��k�	{FH�kȿ9��	�'�d�:5�2�|9x���wW@�9	�'P*�*�� /�1��Ԫ&6�I��'i�T8G��-q��Ri ��@��'��4S��\�y�тȞ��Lz�'��S�#�g���9�$+Gԍc�'�hS�]=4DɖJ\�vY��'�j$�p�A+ �hM8�gD#g���'u��!�O�f��]�u��V�$��'�R��ҊD��X!qEꐆ:,���'���!��6.�R�3U)
�섡�'xp��d^�	���jt�˵.p�q�'����7-0B�N��C:~w�`k�'B���%�D'��q�)ʛzʾ�*�'�:)Cc�ɰ�"H�i�&'�|0�'�\�s%U%[а���
�!*�a	�'�8��b͜	l�%�T9Ĵ��'������P������<w@�9�'�!�L]�BƄ�)��Lw��(��'�� CG4W�,p *D�a�	�'9�Q�N���,���ǮEah�y�'Č�xshALl��-�8P�|	��'���Hֹq��$Hǯ�H"
�3�'ܪ�"c �m~��B+�y	�'�fY��+��R��vt�8��'l2�##%\0��E�PM}EDD��'���H�ϔ`�����K�fR �H�'P:�y�E�>m����6�v8��'�Z<*lE(1el�#�S<-Ob9��'�n�9Ъ��+,q��T�n���'��a�.��s!l�@ƫ®l_�YI�'�:I�$�Z�*(�hEnF�`��hB�'̎]�`�)?b�D�1c.\z�'1PJ��܆�<́��Fqk���'T�0�O,w�1	�!��f���'b�\��� 4@�rKE+V�ƀS�'<����;
aF|I���<���'�D�X��|h��a���-�^`j	�'����FU1G ��I--`~`0��� �A��[�8@f���)8.*���a"Od�0�@2\F��He�)^	�<Ҕ"O9ЉԳUUP%X��C�KXb�0�"O����Mśk"�YХ� Q��X1�"O�ɱ��N�)݄@� �3f�]�"O �B�;@���]'GRJi{E"OFq�aX�0��
�+or�yC"O�����2�T�zl,Uv$�f"O���d�X;�5�fϏ47j�0�"OJ���)ϐ!G��;�$�$p||�"O���	�t�P��&v��qZ�"O����cP�-�0F�B��\��"O
�QDHnu¹V�W�*ڬ��Q"O4�����>�`�)��|q�"Oq"��	0d�		���,oɞ�Q@"O~����I[X1s��S�E�U��"OU	��R�@z����שmV�:#"O��A�h��d
g�M2�@�"O�A�ra��Z�*�Ŗ�K��y
t"O�|��W�g�p����27�"i�"O8��ό�;�He��u�P� "O^�8��ղ8􀣤��1a
��W"O ��[��AyQBW�V�uT"OV���旣�Ҁ[����)h�z2"Of���o	/jx��c&G_t8�"O�I��W�9��%��x)�s"O&hy��-�*Ղ��2she� "O�a�&�)���PtC �
��1��"O�z��=g���6��Ab���y�G�3�����l�,z�@:a�d���Ri@���`G�4��D1uc����ȓN�FQ�dU��⹪�n�^FdT�ȓ82(�@ʜ����U�P�&��__�i���6���%Ŗ1�Ѕ�0Z�5��:�v�d�R�pRd�ȓaW�u�eCҔp�k'C��A�`̅�; ������v�,����d"�	�ȓM�$T�g��t�����-~lلȓDݨ̰1��3I�.��B�I9�I��-���5�&��!�r�Ԅ�C������!9yH�c?9�"U��Isv�c'I�k?�ԫ��eꝄȓư�V�O-`-�a�i��}��m�ȓN���˿a�tE�rd�7�Շȓl5��� �}�.�:�+ʻ<��!�ȓb^hd�CKA��ԥR�Y�B�&`��uw��y4�],�Z�B�耞&<݄ȓQ����hʱ.z���sQ�Մ�s+�9���i6t��>h�`��ȓZz�y8D��1r)*��v�Z�-��Y�ȓ �=�DY���7k��LŇȓt?�(v�J�Z�f�����$ �ćȓC���+��O ��q��$j6�q�ȓY�5��⍆\��u�da��`oXa��\�9��Xtf��+��A�������),]��򈕶Q�ȓ'
�����b����AY~���/�Z�Q�K\�^����	T��@�����(��z#x���v����:E��9�Š~Ĵ� �ܝg��ه�L�� �N
I��`�4�E�%��l�ȓvʒ�;�M�;l���s"�le��J�n�0���+E�������B���g�0� �H3E@>%��O3':@��S�? ��	�!j�t �F�O�^�� #a"O^�T+�$S�B�0��I�e6�R"O����iU�4���h���W�R\��"O6��ri�2��A r�9?�Ͱ!"On��TÜ79�č�K�Q+�d��"O$��a��A�����&&�z�"Od����EI+D�%b[/fm-��"OtX�JP������o��EZ�q�t"O,����_�]�p���+��_:�� "O���fU��\v�U�(%$)�"O�r�A!CD�ҧ�!���8�"O`K�@���Ʃ����H��@��"O�e���̭�2%�hҎۡ"O�8yp&��:���%8�z9��"O�=�FԖU�x�k��ɨ0�)y�"O|ȹf��7�|c �O��"<{4"O8�0���H,^�2a��*0�.� �"O�Cv�U�W�\�ꢌ�N�,��"OjةS�A�'r�	�L�Tr,=0�"O�4��n׉Z/Vq@a��ThD#�"OȨ�͇}lt,{��Ԗ�*��"O�!�d�%;f�P��F�E�p�R�"O�l�o�"7Dn-Q+Wv�d�b"O$�3����?l�� 
�2��,@�"O�K ���!�]Q�e�"Oi*c�Օ.�h,+� �$�ְ�u"Oh�it̙;x�����W���:"OH�U߽(�e��̊H#�hR"O���!�ɯA��ʳj�pn�q1"O�j ���Lz ��j���	�"O~鞴����" D�cG��h�!�Ęc��M+eK]�z� LHUn�%&�!��l�� �PW�� TgPk!�D�$��%*#� 0,��v%��c�!��/ ��I���4^�����e�>j�!�[�B(�mI��-<��3�U�Z�!�Dt#F8A�Q�+����b�q�!�	<��p{�-�8q,��0�@\!�FI
M��㝤|;��he�!*�O��=%>AKuF�/:]��Q��C /WN�V�%D����P%5|6EK�#�����8�f>D��b	L ���Z�z�F�g=D�HC���6�T�2��<]�"k:D�h�1*��F���YQ�Tv�	)D��>���铉n�r�X�-��6$��9d�C�I�#	(i�P�����I��	�~��C�ɒ}�y����-Taʘ�d�D;61�C�I�_�僢�T8��pz��ÙK0C�IH��S�$ŉ%$� ��C �<B�	6*�lq�ؙ5��10d�NLB䉍z�E��i�+C����H'F۔��hOQ>�z�&�9<��51 b�	k�Dl �$D����`�7���
���7~}�\�$D��ǂߗ9і�GU�V�萂�N/D�,��۵��WY�*
���Ms�<a��	X�v��Aѹ6��- �e�<�I��h�60z�Ew��[��e�<��GH�h�nl�R��w�4��HDa�<ч��{���:��W/c����'Q_�<��m:���Ma���e�<�㣜�:ߖ�!�m�N�R4����k�<����A!�� %�B0�IHG�Ne�<yQ�	N_��³/WR�(�P��^�<!��èR�����Ѝ$M
X�	�r�<� *=�0A�VOn���� ��9��"O))��	�7l`T�']2D�0@�w"O`US�m�7g�D��J��5�g"O�H+n/�LXx�P$�j�"On���)�=>�� qаBA"O"��J�0{R}�ǚ$!���pc"O���i��!�ؘ�`+
� Dq"O�`�E�E�c�HTk"I�,Z����"O��p5��17��21�9c&��w"O�T8#�ڞfo�(�"�TN���"O����Z��rF�*n6ͲR"Oj�pփM�������.�N�� "Oެ{�(f���]����(O(y@!�V@ʞУ�lHn�za��
J!�d·�&�#e
P��$�T(a!��M8&�
�tIe��q
��%����S����(�
\
�	����: G6�ȓ_��v�K=m~������Thri��<��X �;0�EA�/=VGBa���~ *A�_�h:ɨ뎵]��ȓ\��AQ-V��A�6��.sW
��ȓ[B2��NS<I*�0�]1&� ��Y���s�AW;Ty4���)��@�ȓtH���?R����g��\�=�ȓ}����FdT
0�"�:$��py�ʓ|b�7��(-X�fI6��C�I3S�Y�p��kS!�DF�,(g�C䉸A7~ �r��H�)ҤA��C�M��q�!O�j�@�O�_9�#>ɉ�iOW
jհ���iv�Ej��ѧr�!��5J�������O����Q��!�dĠ�D)	&*ѐ`X�xR��!���A��2��t7�$S"�-�!���X� K�a �8T�:��� M�!��P�D;fT�F�L�*��?�!�d�~���%�)a$��N���B�.ғʈOf%��'�kh,@�5�����h�"O�M�0aP9|�H[WBQ o��x��"O�M3"ț��N)�a٪�T�"O���+]�_�(��/P�@�J�P"O�ł�D�@X
D獑�
�l�B "O��B�R�`��Ƞ�/W���x"O�@�e"5���I��r�����"Ob��C�U.T���(�X��|ˢ"O�գdl�g@��q�C?��a8 "OJ��)^� Vr�t&��L���"OBMAB9�1�fG�4:ɛ�"O<����k�HX��
	>�� �"O�}�qT)����3�K;H�.܋�"O^ثeJT����I��mH�I��"O8]2�
��w�(�`�g_ e�x�"Op�[���0-x�+!Y#�l�W"Od4���hTL�F"ԣs��"O=��5��Y�#!�6mT�ܙg"Oд�-�9��@�e6�\�E"O���g�^g�Θ�3��'��c�"O,��SGW�.��6f�R�8�P"O�1�"E�=�l(�WB߀%��*c"OfuV ��(�ҭ '��,-Z�yD"O����*LT�qe�y78�"O�m�%0aNt�(4E� ���V"O�t��m�$��\CW��mX:�"OdA3&� 9cz���M�\�Z�`�"ONєo\�X0��;���"O� �9���d?���Ak|�p`�d"O:�c��КJzi�I7$�@���"O���E@��n@�Rȓ�?�έç"O`����Nx��J�G�!Yn��"O�1jtNH�+汱-�O��9b�"O.D�&�C�Sӈ<�CKC�0�"O��ST��?���e(F�Lw����"O���2D^9ou��-BYR��"O�E��N�^��DB�ǌXV�Hr"O���B̒,n	����+�X9�I�"O�9vHR�`��]Kp�-G1d�z"O A �X˞eS�ˊ@Gr��`"O���C[�0���HS*jǪp�"O�s`�_op�]�կ��*�Hж"O�dpT��wj���O�;H�0ö"O�� '�G:/6vT��H�Ka�1"O�d �m�
pe��YcD�w-,Y�e"O�U�m�h0�毑�rLpc"O~(��
�E��EOfD�cV"O:�Ib/�&Lh���6�]�L@ġ{v"O���~�x��M^��vl��"O�U{tn�j�6���T�$t��{�"O�D��h�M�H�z�E�9c��"O09"�EK&$��k7��c^��"O�Ew�i��qo=%*l�"O����ʂ,�@���_�R8�c"Ol��'��4:��t�Ի�`��7"O��	���Z��U�31���"O���d��"*�T�Fe-%P�Y�"O���#�+PN���dD~A�̨�"O.K1�R���s��pE�!��"O�]3�K½T(�`R⠂�~&L�;`"O���eV�t4��R�An�xQ"O�Q�b&N)r������'?�Ij4"O� 1��Q1$�VÙ
����a"O����;��q��3?M�$�7"O-����<�i�0Ԍ&'t�8#"O��P�iM�AM>-��lO�o�=�t"O�@9��]�n� x��)���$!�"OJ�C��8,�4*�`��=r'"O��A�S<N�I�JV�]��Yj�"O��(3�@�bj_�A�����"O�� FX�3��LR�Ȅ9SP8%��"O���R��m����p�*0G�H�"O�]�)Ţe�X���.0 �*�"OZ PD}��Aq@E� Ĩ�"O��ra�ʍ�(u�P�=x�Z'"O�H�5(�;7�4!�eIq���Rp"O���BX�Fv:��ѡՁ1���ˆ"O��Vh�>�.�!c�0�.�j�"O0����.(Ș$y�$K6&���"Oj`���&L{$�^�4�#q"O�d���`�Q�*��m�a"O`�"�%��I��o�-m��˗"O�,K��N��@2`a	?J�j̸$"O8���`Ꭴ��m�7m�&�x"On|{�է�X/�~~����"O�|ز��9J���QP����J*)�!�VX�ԉ"4�B�j�,�)&,�]�!�G�:�h���\˄��`j�>v�!�߀a�P�5n��T��-��FO7<.!�D�<R�P)Р�+�V���`
�*!!�d9(:Dd�D!�!`�!��yQ�qj i��Cv����GM�!�� .!t�*7<j�kGF�:����"O�x�aG�>;�j��C�?$b"O��)A�\6�B��a�9h�58�"O���s�M�/��bG`��5Or���"O�TJR��* ,#Q�;v��(h"OD�e,�g� ذ�0L�8@��"OޅxI�N�Ԍ�UfQe���p�"O�%!�/�r"�"��X��ЕAb"O\@b�Mϭc�~�(�`ٺ|<Ll3"OFE�M�}[蠸p���?8�P�$"O�qS�U�0LZp�K���"OL�Zƥ�,,N)(g�T���e#a"O \s�M�|(x���昗S�9$"O�0D_$$ʬ0!qd�~���{�"O��zb�ғ5��Q���@�*(�"O�<"F���'B���Weޚ
w�qj "O(���^�X��XG���G7ֹ�4"Ob����a�Na��O�Z��k�"O�@�B�M�4��ba��A�"O^Uх��RĔ�;s`ۥu^��"O��2���1\�e��mͫ��*E"OpI��o�q�P!�vC�>8��<ɀ"O����'�<�vH��!��V�s#"O����b�^���s  G�t���H�"O.�Q�L�{�}����l�l!"OL��B���a�Ơz%ό�U]0ؒ�"O� B,F�2hLh�[9@郇"O*�b��o(>�b��.e�� �E"OF�+P��7����S���7M���"O4U2�I�>f�$��6�"O8ģ�e�d��(I�1�L�0"O�8"��E�c5fL�q�'ZM�L��"O�qS*Z�X����� v2���"O�@U�?��c�y� Y�"O�:�Xa��th�烀[;��1P"O�dԈ�D�С��z�yJ�"O��NQL>N�+q�'\� ��"O��P-K�r�t��< � �iV"O�Hȑ�K3[�v��3`��8�"O`JA�M/Y�� �3OަYip3"O�0�1eS�`�j�s��_R쀔"O���
EZdEk�R/�:�"O����ށj[(�#�އE��s�"O��C�I�<6�FHVoE�]�L�"O�ٳQG�y~�TdLH�;;P�Rd"O��b��+%�n��Q�F�!6���""O��;��[���H�1+�$ &����"O�R3��r���0�R
"y!"O��!'��dB%x&a��l�Tyv"OW	vU��,Ƕ
��o�*c�!��^�/�}�b���K�+��O�!�d�U�v��b��S�"�3JʼF�!�ڍ\��D����
�z�Q�i�!�~I��NW��t��ӄ4�8;�'m�A��뛜+��1F�/���;�'O҉+�^<87`�a�P�J5��'���J�%P�����@��J�$x�'�&�X�$�U�nt�p�ƼU����'V�X�T�^-(�0���V��"�'|а: Dב!��hR�`�)[�ʑ��'�z���tN�}����P�9�'�v�9��A$�����B��1��'��{b��w2	[�DB-��@�'�6=�΋�^�đ	E�U�dթ��� �`�)J`�b�K��ΓH�r�	`"O����`�/*����]������"O. �nV�Z LUJ����P%��"O�D��)31��X��"��U=L�	�"O���D�Y
Z9t�T}Av�z�"O�d���"�����Daij�"Ou%�Ϲj�̩�@g2�Sv"O���D�m�<cs���0��`"OL!��`	Z4�X�k�GyH�S�"Om #Ņ7^�(�M[*����"O�}�H��:�l0�T�MyiS"O\�)�=�2(q+L:x����"O����\�F�mѠ��Qa�m0�"O�iw�L���Z`�ݓsxt{�"O%�s��g�Е�$㔀l�`��P"Ol�b��+i�وu�I6��uI�"O�dz���(-w���pF��C���;A"O !�uH�GR��{�e��^�0W"OĨ��j%SЄ����G�VP��"O�9�����Ȁ�;i�{�"OH�#��+.����K	^P,Z�"O����gI?5�z�ʡ(M4�b#�"O�%ٱjK16�(����?�8�0�"OZ���cZ5p��S +z�SS"OR�{`)���@��G�Hq.M��"O��0��5��=���нF\~]s"O:���C�5L��2�.�'
���"O̸CS�E+RJ�%r��Y#W�DR�"O�ݐ�
܁TE�@�^(D����"O��J��I���3���j�T<Y�"O������nY��$�P�'eD"O�]p�I�@7�̊��Z�@�@��"ONtq�n�|Ɲ�чX�
���"Oz ��ڵ<�8�hD�U�<�l�"O�Y�2k��B���p�ܬ*;
 HS"O�$�Bi�z�r �ץ�@8��*�"O¨B���1R���'�ʉ|��P��"O^QQ&�ܮy�z�vI܋�z���U��Y�KҤIQ�i�ǁҤ{����h,D�4��=��т
:Yˬ���F'D���d��5v���,Ŋyvt���i&D�<��c��H=�LX�ǔv�@�#�#D�`#��ܪ?������ ~�����>D��&F�G���׭#'1ig-:D����S���9TaH���pC�#5D����.K������m�ά�* D�l�%hD�R�0����7^���sN<D�����M�<�m�P��9D��8&͛7H:�QdYXH�`¥g;D��1�D� u>��B U�&O�<#�:D�H���WfV��MѥAtا�9D�LeiU1"�l����(_��E�j8D����Qx���'R%7���7�4D���a� W�9�$�PC���O3D�l�%m�#(3l��`a�n��@���$D��P�j�a���A@?:�p9e+8D��;�X��j8�p��&T�2����!D�Q*]�\����>����F:D�����k̴�q�5<{����C3D�d�ª��9 R�Y�c��)eb��F2D�x�D�6�^�KK<g���G�+D�����F�q䤑X�o�Y���1"<D�X�$k^�nc֡�f�$��"�;D���C,�̬ܲ�Ɲ���2��&D�� >P�%�O78���qG
�0���H�"Oj�K���+O���T'��R��U��"OD�KŐ�h���#�f�F�H���"OjPB6c�I�@CT�y�D�"O��)T�U4 ���
{�i;�"OFh��R�M(������؋E"O�����I4 jD4Ȃd[A��(B"OR�sFFU.y����unP%OZ937"Oq��Lߍe�(A�gĹR
����"O�� �(W# �
(�Q�JS��w"O�}�D�Ԩ
m2����O,9l�q"O<����[�$�4Pa祏6~��,�!��Ǎ6d@�U"�,m�)k�3�!��43����0Y1�P�C��&(�!򤌙.������r�D�(Q��!�d
>!�V,��#C	��	t�&`�!�$L6�"���HvL(�4�I�}�!�dMS/�����%���a�:!�$=j2phcv.�9��rc!�dK�������~�ly�A��(!�$�r����'卄g�ziaa�tX!�Һ~g �q#ʷI��<H���sU!�D]�u��9�b��#��щA���.)!�$@
|�F�R��ŤL����D W?!��ǵ8�B\�E�`n
�вυ6#!��[4�p3��u� �0�!�J�41%��/�5Ƀ�V�l�!�ɤl�T����Qhڞ`�F�U
�!����+�����Am�j�*�ńS�!�U3/�.0Q����f�{Tş#z!�ć�"�D�;D��c�>"��y�!�D������D�w���Ӎw�!�dQx"KαMZv]pO�b��9�'����qA�p��} �	;X���
�'��P`b��OWf}rǋȒT�E�	�'Ŋ���QZ���X���	�DX���'q$(�D*ۚLT�p�J��u��p��'��Wi�t�HH��o�3|��I�'�`̛EʄM���0� ��� �'�r���႗;�z��0L�}�>�(�'����؂lފe)�Cm�0Y��'M����M+.I^E��J�k�F�+�'�ڬpPf�(H��MC���`ܲ���'�f!y�c�Rna��=�HQ����x��E�l��w�DS�R0;�X4�y'K#Y���Q��5 �"�'�$�y���!���J����p�)���y�&����cj�4�{�!ϼ�y�M� 5���e3!��y��%$�8D�"��P�Չ^��y��)?B��Qjd���`�̀�y���0��٨�U[�2��vhP��y����B�KLH�Eg(�+_�>���r���F)L�2����b��-�@�ȓP\�<y��܍[�F��"��'H�����Zq�#� 9,Y��ژ���ȓ\��y�I�TAذHP�Ja��t�?�
�
Ĭ�*��RuZ����u�x�ȓ�6���V�JU�A����V��ȓ���&ìIq�ț����>D.T�ȓiHv�󵋊� �L�C�K�5�0Єȓn�`t���X�D-~��p��AB���P� H����*�c�Bs||�ȓt8��ba��U�^<���p֔��?���0<� J�*��7)[�x �f�w����"O��3�E��"99֦�2X��"O>�#&J�m8���4H��=��"OPA���5:�<\PA��:/�l��A"O$(�Q
�!�USMޣAb����"O��3�$ʙ
��;5�.̺"O88�R�~��Y0��ˑ8� ��"Oʩ�B�iz⅃G��X�Vٓ"O�=@��>�<R���@2"O��1���@��vN�X����"ON#��D"V�R��p�Vk�"O0����i�XBٔ=��eC�"OP��@��076bP"��%"�f�D"O�Z⊘O90���)ɉ���"O*�E�^J� �H]�|<j�iG"O� Ab��������?R:�5!P"O`���S�&�t�L8���²"O��ӂbΔTT�5����/
y�"Or�`Ԏ�1r��	��K��4��f"O��fo���N���%b"OR��tI��@`F�����,W|y[�U�DE{���K>���k��,�QŊ�J�!�L \���2���,E��#��C7p�!�D�N��C¤Jm�5�SC���!�dC@,���e� ������i�!�$(u�ЌYRᆏ~�ȉ���,KX!�$MGJF���I�1a�P9B$�C�DF!�D�o���\3�6m(s���.!�䂘6����U�G4�pT�Qş�)�!���om�9x�-�����#�7>Z!�dY6 Z��7瘮-��� �� L(!���0F��d0�	�^��ɗAU�w!��Y�!2��P�0��`6@!�䏠
��H��[��(j�E�D�!�$َ~8��dI�0J5�TI��!���O">����T�|j��F(n�!�$ <Z�lo�? t��!c�I!�d9g����!N�)��u�h�T�!�$�<D�<<X��	U��q�AGR��!�d���R��` ��c�� �׈ٍl�!��Y x4&� �c�;�GH�^!���Mh���1�L�q!B=�6G��!�
�'��{���psd���2y!�dA�u���yW͖/�7D��7r!�d� f�@2��'���Q#{;!���w[ i:b���2�h�����Q+!�ā-fn-�4NW����i��T"!�0h�����[�ā�Hʺ
!�D�$)_L 4Nِ��aJW��%Grў$���0�u��̪ )-��`," �B�&>���XT.Ƈ~Ԫ��Ԁ���B�I
 "�X�E�k���A����C�	=T��d�Y�������=a�B�I�j�tl�0�0/�j�b�A8��C�	�_o<�a���.`��B#d�fB�I:����%��P ��MAf�B䉪G">1���9$��睰E��B�	�6�&�`���
a���؜!	�C�	�V�F�(�(j�����\)X�~��	�'��U��L��Gr	QbPy����'�L��Z��$U�Ț08-v��'�詹�%�9�h��_0�hZ�'��,�O�)mŌ��� Ձ������)�tI��a��b҉ǚ5��x�%���y
� 0�� ZR��;�i��� "OJ�y&���h �ڬU����q�'y�'��)�'���T�U�[�`+��ιk60�x�'��kG�6�0i�Ӎ^�e6\m�	�'��@)&*Z.��R���_��(�'M�mxP��S�����:S1a �'=�A����0]�F�%P�DµJ�'�j,"c�v�,+�C%=�P, �'�:�4�&!c���,1F@;�B�)���5��m���ܬ_(��k�@X�yҥ_*{x�����=W㞔#�C
�y��T�̸�/
�Țy;����y��\gZ�(V���P\ѳ��_9�yR�
X<�q�5�9;Kx�i��C3�y���'2��	 �2-5"�K�����ybO�4�|͈�O�'�8sd�_�y�ɑ8�y��A�u,��0gީ�yZ����H׼k��0�DۉsV�)��'��	P�D5$^�H���̈@��H�'�\�K�#�4k��Hd����O���!A�5>�"Ă�._ġ)�"O~�ƣ�?h=2r���<r�D��q"O2���E-|c4���s��"T4!�J�����CS�(ȧ�W:!��)D?P��F�����t,�+U|!򄊁o�pJ�ԪdtJ�v�> o!�D�({e��1!Öj��p��,t_!�������
�^X2h��.�!�Ğ�IpP(r�k^�\��1t擦s!�Nz|Y���T��p�A�R0	!򤚩':�;7%G=����V@� �R�'3��'O�0�@�Gn<b<I��� �m;�'� 1���A���p�Q&q�]3�'�Z<��Mĭ}�5�qfAfi��'��T/��.gx ����+Q�X��'2��*Au�+�A	0Y
�E��'PR �pއM�>� F��e�~�*
�'�,h��]�l�����F�K� ݐ���xB�2ĜM�&$�%)�q��yr�� 8��D��ɘ�&g�հ���yR� T�J��f
��ӈ�
�hO ���JW�ՔN�D��ĖJ ���"O�	(��4�b����
�#�Z�c�"O( Y2!�0��is�K 4�%
&"O2xp�OHg,�Q ��z�����'�2�'`a|���)A@�1H[�'O܀�7���y��G0|�����jM<A���,�yBb�{A2�ӣ���R�v�[�$<�y��Ȕ���pW���G���J�����y�ˋ�W���K%.B8n���È�&�y�
�! <@PBl0o�"�nל��>��OƜ�p!6I'΍�$��+���bd"O�!'L�2)X�x�%~rJ2"O�I�0b��-[��uL�J��"O2m�w@�!=�aaD�_��1��"O�J4�I
'�t5�@���b4���"O�ഥ�O�(��pL�,Q��"O9j6�V�#�B��i�kBU�"O"�R�O�' �	���iL��"OP�B��i�4�:a�	9LU:R"O��T��;R!h(�LZ.LH��E"O��s��A���AQEۖjD���"Oj��PN�1�2D�B$++<r'"O����7Fx�E�N�)Y�u3�"O� ��Y6N�'^*4��G�-2K���"O&(��=I��E`��[� a���"ON� j�Z����Ƈ+DP��"Oz�Fۧ��XK�Y]��ku"OX}	S��5_�P����ф0KP-jqO�4��-��bB}��3+s\��t� D�����1S��&	F�6�AYщ?D� )��.V����ĭ�UQ��=D�P���{�����ï*L�����7D�ܡ��[�F���qc.��*nx4���1D� �Q���t��,��I(MI�(�$+D�� e֛H9��Z�G�'���yC*D���S��(���A��EF���5D�A7J�<cBX��jV�Z6Ĺ⧠3D��"�ڊ.��4d&�{�%3��/D��A�+�k,	���S	m2���gA�O<B�Ɇ8R��ʆ�MSy6�8@LvtB��C ���T'&�p���Rm�C�I��>�P�dC_��a�K��eo�C��(f #�X��� J�
�m�nC䉘��l�'���r����$�LC䉺I���j �S�~@�����'�6C�	8 �dh(5�׊h��	3)B�O�FB��36�<c�.�,Gy(#,@.e;B�Ij0�t@�A�X�q����= ��C�Ɉ(7�����0N�Ƹr�o��C�I��P��ћN�J9ѿR7�ʓ�0?���8��e��Ɗ,��0I�W�<�p���|�1/�<�쪵��R�<�� ��'���5O�0�4���e�<!�k!|R`{!�����!��e�<iS���dP��X'%ތQ�|A���b�<�fF�*4�{C`̡VG��s)�J�<qq�߳?�*��`�ɡq�0���n�<Y��ǿwm�-	���o��f��q�<���'$h�� �6b��6e�j�<A�MX�4���R4E]#��p���e�<��O\V��Y!D*�D鸙�c�<	���
�b ���	[�lEB�Bd�<!���^6����n^��xi��\c����<�W%�/��DK�C�+�8=&+�s�<)�l�,8���dA
�!,y�<IRKZ�;sҝ��.ڡ?mF�c7(q�<1!�3z)�g��Ha�){DdXa�<��W�DUP0��[0:4�!Ǆu�<S[���Po*?C>�۶�p�<����,Q���M��5Q�\{�GEB�<3�BT��ɡW�Wq�Jẵf�v�'��x2!ӷ���g"A�@���a�w�<��HZ9=�0���*/�Z�Gn�<!s�ƧR�v,ԯ�~��Q���c���?YÓcƁ+��\-l�8X����j��<��^$�T�	�/l�;��i2F�ȓ2�tp'�>���҇�0sw$���#����!?R�$��eF�=֩E{��'��f%0�\���\6(�<�r	�'� 8`@�G�WYF���H�7w�����?9�����+NejJ$oX�Uv�� �F���(�d#���(�8,Z��H*	�<�!!D��إ, )hP�4i��{��9�0�?D���@fT-J>XiB��8o��Q��B8D���E��'zt"�y��;8;>��fn5�O�bb��VgO�U��'`ӿI,̇�VĪ�΋��x8��d�b��S�? .��K%|�,��s�)M��t���@�����p�X�
�Y��Pk#,*D�T��b_�e&�b�m˻��,@b,)D����l�45Ff!K��)���I%D�L���ѻl<n�ɵL�.^��bG$D�D�dG��N�f=���[z��aP6D��p���:}�ͺ���
E���2D��hg���J-����a��yNu�A%D�r��.��`˰,��c<YZt�-D��N�A��f���h��DF+D����L��O3������g�sFJ(D� ��M0\ю�$Ë/$t�Q�d-%D�Ļp�( ��%�w��}�Ht�M=D�x�f`���7��,J~d��F<D��zl�3{t}c�*�� ��bE0D�� �(J�o<� ���ɳ�A3D��Au&�'.��І�DW�t��/D�@�#��,h":]��۸�J:ړ�0|����,쬬���#Uh�����E��d�|'/�W��]9W��hpr�,6D�0AW�	�Y�A��# m`�G�2D�hۄ�]84@��쐳X3�8i��<D�Ԋ�A^�n��H�6}��� &'=D�|��."�p�BS�N�g���Cf8D�\SvȓE;�
Ё�2��݁��6D����y J���K� d�5��4�*�O��BD�˯>5JP�
�+ݰ���"O���#A#N����Z�r�<�T"O���r��;^L�W�R�n���S�"O��(Äd�dM��@��@xi�"O`�`A�%~��%3`�^#:y:��$"O�A��KQ���Pi��ᢀ��yB�׆�P��6�ӅA��m����y�F;�ݳT%[9A�fh� I��y�c���t�C� �9	�x�,��y2��2��]��&@�.��8�$(�$��'�azRM��v�d�&ϐ�sҕѱ�S�y��ɻ��������?mX�؇�y�b�9GXٰ�̾3�� �`X��y"�Ԇ'v���� *�("0C�yR@ ��Ѫ�BҖKcRYK�N��y��ߋ$�ZIk�bKCo�L�fW+�y�&��O4I"��VA�`R��[>�hO����^SFP�Fm�9._�M�L6N)!��KL㲀���\Q��c�B�"!��:F"n�A�!˷Iz�r�ʈ�1W!��۶nl���C�W�%9\E��)22�!򄒝g� I��F13��!���2�!�2S�(m�v�,w�@����J}!�
�(,NزF��5>�{��I�$Z!�$
h��P{qDƲ@8�V��BE!�$фF$�<�4��4�b�8�e��!�D
�6�>-��kG�|n�x��D/!���"��Kѥ��p^ؤڱ�{d!򤎯7�.���UgMbAۓ�$K!�L�S�:�x�eZ�IA^hbNȡ�!��#%��ze�Դ}.d!��{�!��=��*V�:l�����aP!�7zp���$h�UK:���@��e�!�d���:@��-:,��� ���D�Q���ȋ-Nл�D*K_�C�	8��$��h�l�Q��G�k@�C�vBL�2D��U�d���0�|C�I�j�{���,�T�B�=�LC�)� �X	�"�4(���%F��y�^,��"O��B���7������	x���g"O^袆��p�Z�yd A� ����R"O����n�	\���2��]:e����	a�Ot��+Ư�0@���GI�5���#�'�|�Y�H)c&x9�5h1�����'`���J�(C"����V-b8���'�Z�HQ�F)`��#H�s��@�'��I�p��
���#
f�]0	�'��Ȱl��>��s���e ��"
�'n�݈�F����P�s$�+j,A���D;�A����ף��hS"..H�ȓ[���xa�@�+�䕘.<B4�ȓP(0;���
��$ҋ�<���E{B�'G����VP��rRc��~ �
�'�f|
�(��Q�I�J16%D�h��E
f��5��V�r��i�g�?D��"�$�c|F4Xs�V	'�� YE	?D��KQ�Ľ6=}�F�����(aH:D��1�O��0�Hic�ϖ`|��(�j2D�����0Ytk��
��,��B$D�0��!_�Z�j1@O�Y�lÔe4D�Xc�Dt�Br"	�
%VD�ׯ>D��y��!*g\�b�f�cYX��(D��ᅃ�/�8XFh\;n͞��O��=E���O#6����Rը5�t_-M�!�dK�-�Ҥ��X&W�:����k�!�䈿c�t���DV����S�e�!�d�GMz=$�$�������!��_�;ˌ8�2g��o�6��FL�i�!�A�Z��m��0�� �.e�!�G7|�p!	2�ș*%�Mh� �%U��O�1�A�R僰.7N����"O��[���*&jȑ�N�)F~dq��"O�(�&ʐ�"2`�A�t���f"O�!�pG��V@@����[z4	�"O��J+=4!m�mX�@U�y��"O҃C�@�v���l˕Hk
q�B"O��듆zʌ�Fօ1,��cW"OzL�0�V��l��ώ�l�;v"O�!s�,��p��I��$�~�sF"OfРâG8ms���Q�4@�>�hF�|b�'���KX
�|PN9El��
�'?��+��־Bf�e!R=AV�	
�'^��[!H�z}��5��5�~u�	�']��B�	�<�b�+W�����x"�օT�q3֢�*J�����B��Py��ˏO�`RЋС3L`J�+�XyY�PG{J?}s�$�?Eȁk�� w���5D�(+b �& s�;�٫4ɞT�w�5D��(�Ǒ8U�r�F	�X�TLI��'D���h�7T��q����~�,0�Ul+D��j�a��?�f̈p�%���;�K'D�+�L�0�L���+��/�V}�t$�O��O|�=)�O�A����Q����RI��qx̻0�|�h̓@q.�y�(ëZ��$t��,g��'�Ą��l��%r�%G�RN����D�hC�	�XI.����7p�:|	�O�5G�JC�	Ol�Ix��˜:ԑ�&Ƞ[LFC�ɢ~�N�6I۞;�@D:fˀ�b�6C��&s��5�P�ΊT>*#@�2��%D�<�q�o�1����v`"�0CL1D�$�	�9&\4�cȞ[FH�P�4D������kx�E��^1|�6Eqs�=D�� :�����R��ag`гu�\%�e"Odpr	W,P�$����Ѥ�*`�r"O��3�!m�@�zE��2��s�D5LO�` � ���l�q��7I���H�"O�(R�ʻ<ݚx���Q��Ts�"O�S��/b�ma���r9�$"O��X!hkt��#.ʈ*��I��"Ob�$mǅZ�z�����'K�<h�"O�u�E�C.㮀Ȧ��1�]�$"OL��A  ��B�"X��q�"O` ѐG/n��%��Ѣ&"O.��@\ D�������1|nB`"O�D�a�	��٣��'��F"O2���B[�,v�l�-��!�.ez�"O֐8�.�k�Ԛ��Z;^���K"O�	�c�	\�гpJ]2T�lm��"O�"BW�U�	B@�Jm��˃"O^�XU�}���� [����'��sl� _f�����	>���kr�8��0|b�Me���!(�e�J���l�<12�n��W"�ܡ�E�H����~&l�k�o�=	�����Y='��хȓ\��	u���ht�;�)���ن��I~(R�\|C@#ϼB}�%���J�hO���DRmb�R+�FKܨ�d
�!�DЪfUXܪ���l1J��t����O^�����\Y6M����y���@d"O��nۣ;�2�����^ոIY�"O�Q��C�  @��#)V�:=�"O�@��̖�����""��dT��3"O
lҴ&��Q�ݑ Lu�XaP�|�)��3��=��B��`���:��D�C�		�>�iFM?"��l��B�&�P��I���d�w�ih��A{�<2"O̰��W�0|h�!g�?c\�q�6"O)Ä�/G�8Yh ��=MZP�""OԀ�A���X*��� �Òv��,�0"O�Qa眽\���d�KBa�v"O����k���Q��J�^����"O�a�o��Qc�����|����"OX�'�ɠp��}a�BY�����"OFd�a�X�lR�8i�>	�Ty�"O�t�%`�9yF��ubD�5��YB"O�k &l@l ��9��1"OjI�4��N}�<�
�xF%��"O�q�d	��^[�hɅ�E�Ѐ�@"O��m�5y� "f6R��P�u"O���g��n�5�6�ņq�V�q�"Op4#�KE���t�0e%Jt}�c"O�0��C��2lI���V�nxp""O$��G��Lw��s�L�r'"�9�"Opt��R�`�~���:)p���"Ol�y�EV7��a�D`^�
���"O|h�ė�=��ЉF�^�V(����'�1O�Z`�Z�\^�( R�Z��Jc"O~*�8~:���P�,�� ��"O��;��G�0�����cHp���a�"Ox,��F�>bB^���������"O�<���`6���<A���je"O y�E�Ҡ
0I�FI����0�s�'p�|!C�bvbYi0lP�H�~z��O��=���	� ,h��R?��3�8b5�	m��Q�H�N��U�O��v��K&D� A2�?z�tQ��̓R}��ʁ�%D��  5!%�"`2T��1��#@"౺5"O��bE�б;zy
s"ȴ]*4̛�"O� B��@�Zʡ Z��j1�'��58#��S��H0ܮl���_�ͦB�ɐs����A0]Լ��f��V3�C�ɝK�`�Z�"q5���%�2-/�C�I�Vx�@I�e�;񶈺�	�%znC�ɁV*�ct��%�d�V��#�8C�I��|d��&]��JQ��,��B� "������4��e0D���#����<1�O9#`(ͻ8-᠃M�"(!��+P"O�䉷g�8C�a�T��z�p"O\�a� c|�TZ���/�@i`v"O	`�C t(.�;�,��}}�E��"O���fDӱtN�m3��J�.Nf"On4��]O�d)�+O�zƜ@��"O�U��RsÈhhB���2�	n>a)��+p��a��/&=F����)D�TcP'[
ʘ�g��%`.<u���*D��zm
�6p�����}��B�-D��`��ݡK*A���L��$���)D��	�'E�r?d����f��RG'D����n�y=L���g�6<�V����#D� ��8T(D�Ҍ�I]>4ʴ��O��=�O��I��񊓈'%ѩ!�ɊK���#�Q�<&�>C�ܐ$�ל�
D`�Dy��'?�Ĩ��$^��H"`̊A��9�'�B���7P��b����J���'��;&nL�b6�I�!I�z���'��1���ͿQr�i2D�u�d�H	�'t� ���%2��Tؓ�\.X�>���'T����}.��)cȣ~�2x�'(C4���@Iڵ�ǰv?L�s��?y	�M���+��P����w( �
�1�ȓdF)`�ƞ�%����GC�p=��n&�� 0g���ų!e�Y��Ň��"�ۥ��*����1�QK�x=��5���Z�'�72�c\�}���'�ў�|Z����H@��P9������L�<�dm�siF\�!�S8r�n�  �\�<�R-��M����4m2����HM�<)񍅥RL�}I�/O�1�J ���a�<���3~�$[p����	�,Pt�<%�H,Y�C@�/\�P��p�<y�n��J_:�1փ�%C�6��#Cf�<1C�o�f����5',�pӂPj�<Q��L�{��Xjd�˝�©[ �e�<Yw˖)<6d���G�i����b�<i`-X�P�bs�Ēv1X�a�Ly�<�B"A �<��eL�S
,�`��v�<�A� �f~�B�l
�{Z28$.�q�<i�a�)�8�"��z[�b���v�<�B��|�X����sa�XcE�}�<&jɥ,M��!��#is�r&{�<9�mA����CE픫E����HM�<9tlP�Y�"�h.�+:"�mQ�k�J�<�U�
��(��͂�"J�,���F�<��m�G�|����Xo1b܀SWK�<Q4E�Pd"�q�n8��H�<����-k��s-�o|�⅙C�<ٲ��i ����a���$�XB�<��K�8'�h�
��j���z�<�u�G�ܨ�n�@|L�Jq�x�<i�ِ_���s�CY�4�@�
�r�<� p%bՏ�y�����!D9�#"O�ڷ�� &k���`N��6rp"O����AX%����%`b0x3�"O�#��ΐ�<L;eoO�/�FcR"O�q���@	%)��"I
8T��A"O�u�W�д34X=x�m�U"O�ͱ�,�T`@�R7A���59t"O�9�r��lrр��̭
@ଊ�"OX�j��R�s�@��E��"�*�ҁ"O,=fgB��B�= ��(S�"O�pÚ�Lej����I�0�aI@"O�mB�l$ yZDlڴޖ%�d"O( SC)ܶ&H�a��!X�%��dJB"O�0;�*�^4a��Wr�����"O(]�$�[g��ч�L���g"O ���f��x�ΤK$��[�^)8F"O�P��̟�rʜ�ᆎ$s�",��"Ov�)�+����R��`�z�$"O��K�!ԇCC&0�P-"���"O�{tC�'z/�2�WF/x�2"O��1Tg Y4���g7t'*��V"O�0:!�\� ~p�+6�k�آ�"O|�$�{��p�g�#i`��"O^���� �z���Y��-�S"O�	@<X�8(2��%)��S"O�e�E���u��_���{�"OhyB�X���9��80�)�"Od��JؖB������%�T�T"O����A' "}�ӄ�K �K�"O(��R�,�#�
\+�"OA�"х^p�#D�&���!"Ox��)U'U;�-��ZE�i�"O�y�5 Z�vǎ�q��1����"OHe�攂[�C�`�>�@T�"O���ډl�
T0`��Drbɲ"O �BA��~��$�e�T�x::s"O�k��݊ ��:D��'�65�E"OlMY���8Gf�j[	e��a[�"O�� #�V��4��h��V��x��"Od���!�r�d̃��Zf��|!e"O�"3EO AT��gݳO�I��"Oz��Gȝk�T��"G0`%�u�"OFe)Z�t���� ��� �'�Q�!�L>2(~�:���$P����w�U6v:!�>
̭z��R����W���|!��Gt N�pvKP28������n�!�d�) w�`DoE�	ۘ�!-�Q>!�D�j"D	�W�]4g�U0�5#N!�dY]�,5��b#[��R��m8!�䖫ksj\jTiK�n-��,A"!�dS�{��9�Pg��Lz�D��$K�!�d1���q$J�!�r��M Z�!�DD���6,CU�n�+V+ �!�d�{K�HS�(����L�����bt!򤄁l��9��Õ
MVG���pe!�$^Ȣ�hV�Ϯ H|�� ��\C!�dB�E1ʀi���iGԘro	'4!���
�2aDa�308���[-!�Dl��zQ��pM�$�6I� !�D��܀q��DE޵��H��M!���5����e�O0Hm�!i!��z�A֜NT�-��"ܝ!R���"O��c�+�! J`/��m��"Ov�q��8F�ݳ�$��G��ʁ"O� �i9��Y@��2�:�Ʃ��"O�%
�#�CeO��F���"O��%��7�B}ѕ���?���"O����j]$&G�XxJ�����e"O|!P����x4(�
#���U� ��"O��%.�-0���R�(>a��0�"O��u�T9t����7,U�Yt��Q"O �s1�̒;�L@6"łw�d8�A"O��2��:f���76m�Ȃ"Os�'մ>zNL1���N!�5%,@|b`�H��ؘ�ԭ�=!�B}"@�qn\���Kg�I�(�!�䕒D�H�+#���%I`ˠ�!�$�N�����Ŵm�ޱ�׃��!�'�L�*���d���¨�`�<�T8(�(YSƠ2\�W��v�<A�M�k ���!o_��Ţ�Z�<y�I���m��3`��j�fPW�<Q�� �a5����I�u����e�S�<��Ōd7&���͖�l�0psaK�<�⭌�f�-z&�_�+���`��G{�<�d�@�6`9˲*\�0l���m�<�QcA�k�dyQ5g���s��h�<Qv�ҭ3N�	��N�E���b-�j�<��)έ�(�i��P�s�l9�P��h�<��1@/��y��2�N�����]�<i�.�)���x���q�  XB�E�<	 (R�-�욒ǎG��x���u�<�֭�O��t���	�+d�A�D�Mt�<9���*[���Xg��T�q'�p�<9gdB=��� Ŧ�C>X��k�<���o�v4YE�gk��J��f�<I�k�<X.�)X`铈t̺�h�cTd�<)#�љ:r!tm	����ed�<�7�����Z�8�t��U�G�Fk!��$}�N-H�	�5(|��@꙼%j!��j|��(W�@p���J2$i!�$ѓZ�҉��e͑W�kI�4ic���vz��� pv]��Ĉ�y��ܜ{7�A�1)��f�J�uΘ��y2�،�쑻%�3ZÈ��
�y�l�$4h�*�L� ������y��K0" ���E��Dyr��tD�)�yB��'}��(P��Gf9��H;�ybIJ�vI���5n�B4 ec��Y��yB�Р�����mS2@Z`�K��@��y�N/6ǎ�@�B�2@�D�b��y�D��xjr��X�.h6�hR�E=�Py"N��>��Jd���o6m�)�|�<�0	�&HY`M%J��Tc�HR�<���S��,�DZ�!%�ȩ�#�v�<�@�I�[��( ��7^���yB�]�<9�Ѽ~��"�߯���q��]�<��X��4m���]p��Р�A�<I��B�cxDaD"�Q��d�f��c�<�r%�$8h>�h��@.)ҬZk�<��a�"o�6-���#�b���ɚj�<!D���!2@Ջ�G�\XJ�����~�<��!Ԡ5�u���4z��|
֬�e�<�qdQ,��S�'1(�f�k�,MG�<�E/��VW��qХ�MVPz2�QX�<�V�B��)�6��
}�����&�z�<��]�r�lX31)��H��e��p�<9�ӗK��<��	?g�j)	�M�c�<� �*G�G���2�-_5-n��U"Oƥ�T�\�a`N�e�Ͳ(����"O�a���M�g���#曬X�0�"O�U��a��Hu%E7MG��3�"O�|��i]+\�z������� NRe�<a�(ʰ,����$h�{�&�a�<��k˺_���1"d$j��x�<iFo��4��x"��x����At�<��$ܴX2TtB��<��E�<��!5��]�m�����ƌ[�<�b!B�Ø�у��g�x����[�<�A�_:r.���aL����a�U�<�u`��M���/��+�!����f�<�3*\�+�v��פ�D�2�h��a�<!R�5W�%�7"��񞄐�E�F�<�CN�5+���z���C�D,���|�<Yq�|C6�i���@�ě��^�<a�g)an)3�ɑe`l��-�]�<��G��v��-J�m5g�,!��EC[�<�0^�t����o��P���p�<��a�J�Υ؁�DǮ���KCE�<Qg�q��	G�O�x;p��@�<	g,�6��K�ۦ:�2c�}X�o~}�O��\���P�		J��aխġ�yR�¡2a��j1av	ZE���rf�	G{��O����S�F{b���.��=�9��'gFH��"���c�ǜ�];$�'�6��W�`bQ(���PS��c�'�hqq��"P�D�vi��I����'pd�2��8W�0��V��8�'w�l²��N�y�ea[���'�����UW��jU�Ֆ|^�qy�y"�)�S��p`�2�љ ]�G\	.�C䉑l��Ѧ�L�����>l�#<�ϓba��ID�Ņ&,�������� �D ��ϓ1k��@gݖ��\�ȓ,������
��H�`�˞e�ȓG��q��B/:l�P��m[�f��чȓ=�^X!s�Ζ{���{"dU�jr༇ȓ[�6���l^>T��W�1y�ŅȓN�vu*t�7�x�3�M# T���s<���.M�5��!�t	Cs�6���)�t��NH,����I�0����%i8��SU��ʼ+ L��k�a�ȓ,9 ��@&�{���T�l�ȓ�jP�fРB���U���[~���ȓr?BY�aE�(;t1p���� Y�ȓn�rJ�����0p ���y`�����L�����ŨI:�y����B������b�<�p� �>�k��;+�DrW�BW�<a��׋����D�=,8,�R+O�<Q�l��R�*�c���?\��<��C�<Q�"�0! �;s��=�&��oR{�<I�-�� �P@y��Bf��p���=Q3�	 �Z��Aa��;�AG�<)aH�
 Ѭy�`=��ȃR��By�'_ uC6�Ӂ>;vL��C&͖T��O���ǔ&֘d��NN	8D���n =�axbP�X�>��%\�$1	�,�� ��m�4�_j��0}��"�'��,:�k΁4ul�s���5=h���ē�4T���04\��R��݄U�LP0U)IQH<�'M@���r�aH�6^E5,��<A��4�>1�>��G��4\4C���`�Hԁ�.�?��x� q� s֪
&Hx*���:}���_�� :�T���f��d.ѽD�vT{7"O��bL�6b��Da��9�Q�A"OH��!㗸Q����-����g"O�E!�j��R�ѓg�ѭ2��� &0Oz���
�=�Y4�3 �6�S�fB�	L.$ᡡ$]�w��	&��V�C�IY������*-���Y�A��	T�@���.�m�ԍp���`"��#��bH<ф K� �BX�`ҶX5|�8rI�'=N���<��M���s��d]biڀ��"]@���	Dyr:O�7�:o JU)�@4]\�σ��c�<�dAH�f�x���Q�6�[��t�'Y�?�j�ɒ �����|ږ	�D�6D��c#�'	6a�����H��%5<O�#<I�k�.�"�1���%�n٫0)[}�<	a��qgFq��	�pH¦A}�<�b&�Uǲ�1���K��)�f_v���'g��^��F
�����``׵vwB�b�84�4Qf��;3��0��ܜ9޼�u�:�	�<��}Zw(�	Z�!�o�+*|ءA@�4[�rC�	!jk�	ݻ1�U�t�� )sr#<�A�Uy2�I�ʌ���:H�(9)ы���y��KX��S$��Bx��@�)��dB�	�9D�L��iۂ��C߳�B�ɬGЪ��`�W>9������*�6B�	�n-r�[�f<0�����L��}}*B�ɴZ�@�c�Vl�x�(d��~T�B�ox���xw4h��`,���d�<ѰA�e�b��ՠӉR�V4b1`R�<�����NϾ�bGÂq����CO�'z�E�tO�%��EY׏��F�|��.G���<���K�Zֺ�;D��v��֤�%[�TF{���'oM��*=Y�X�hB�+���N��xp�6�S�'}�TR��`od|��ĻDn����?)E�2O���c�03<�#P+	nܓ�ў�OeY!�"�VL�S�>;�0���
O�p  �L�-Z%#�G�	��y"I�9H��@�cK��4X�vF7�y��"`����L ve�8�š�%�ybJ��A7�����i�2ȡ����y2���f���e�|�c���ymT?*þ|x�n��Vζ�S5)���'nў� q� C��SL�����քC�D�2"O,��p�L).��10Zx�����O����!��\B��E5Mw���ԡ��!�G(x����e�����PCC�<�̃��)����2Z`�����L�D�"p�C'D�`s磋�Ip�Q�
��<�yBf��t���ZxνC�h�^8��*�+ݼA�pM̓�hO��+���vE���bK34p.!Ȗ�P��C�I�(�a5m�O�<���g��q��C��<c�*x'kS�o:���bZ���C�I�b��;Vf�nCũF(٣b@�����1,O$�y@n��w[�a�S�S3be҇�	K�����s�!w`@�9�"���U!���v� 4�R�o��P�s-	����,�O�Z����CF�s�F �%,�={FOh��+��w���LQ�Х��� q��ć'Ӓp1(����P˝��yBl�(�	�.M�.�
D�w�%�y�B�GFU9�(=z�q(G�^���O�~2���D��,qB��>:8V��l�<1ŋQ�;Jv�BNRG�iy�-Bj}��)ҧ�u9uI	�"	��bT�q�����S�? ����"\$2�,�"S���7L��"O�DI�	�&8�K�㋝a�ld�s"OjX��A�bR�@r�A�w��j%"OT����T\�#Ce��J�!e"O���Q��Oa�8��D�/U���&"O<e��C�M�@���J�3-:#D6O��=E�$�D ,Z��	\�v`� ���y�fJ�����Ҋh]���S��?�J�0�O���8�t�@�˄���Bp�Ș_ ��ȓP���� �ɚ�JVmX!�ȓvǈ��OU'Z���t(���ȓsƦ9��هn�ld�Y�Dk��ȓZn^��"=��u�0�P�Z�p�ȓrM����Ԍ*���)��c"4�ȓg��@�Ht�8�V�0:�.Ԅȓp��8�����mb���|�ȓ�x�IBJ��P��hB� �&b�V��$êI� 'd^��� 9���:(d84����-2�-4>��ȓq��K�$"ΠL�	�1���ȓ���2w���9����Tgt��f�����j'�آ�2ߌ,��,y8��FZX�Q�w�[19q����ox�C���mœ�O+*M�Y�ȓ
�0��N?`<s�D_�P3��ȓZ|i4c�v�@�������tUP�����Ւ=���Y&6y��SN�6	�_8�x�%i�{+j݅ȓ`��)b�˂?�J��f^�T�L4��$�@}xg/�\�`�Yv�\�:0��ȓX�m��,ro܁!���2#r���ȓF�����f�ƌCE�(Vf(Y�ȓe��A�K[��$�C�.`!�ȓ�A�c��J��rS����B��ȓ",�Db�Ɩ7E ����H�7Fa��{2DA��ϛ4K@��G�Y")�-��;9^A[��>G��à��V���ȓdVn�	�n�$ �$�V�R�8ܜ��6'�2�#�u����W��.C�d��0�����1p���GK*_,�ȓsP�g�+|�)�<�du�ȓ�؅��s紴����$�P<��=�6M�� �3 r�1�v�Q��by�ȓ"訛 R�	X��!��ߪHB�bO9�>	����A.���&晉$#`�����=
rB�ɂGX=��h�	Nv��+P���X��C䉉"�]�bƒ75$�]s�&�#I%FC�ɔO
m�Q�:�="���.C�I"?<9J2/����s�BcC�I<��0 ��"Y%�(*V�.��B�I#,����ѭA��({��NhC�I�SxfU���(.:p,9�!�ZilC�I?PniB�� �4P1Æ[�B�+,���6A�F
���ebbB��:`s����]F��q��'^�st�C��>cQ��ӕ�{~�QpL�
פB�	"����D cp�����0 ��B�	�G
N���딨��%2�A��5�B�I4]�P J=F���àL	�`��B䉝�\Q��7,�(�KڊhNC��� �`wC��c�tX0O�n�XC�	!�f�0�B~�����A���C�(ސ�!JQ�9�xp�@�Л�C䉑o�PEq���g�L��eBحvLB�)� x���E߆r"��B�d����"Ov�rU(ckv�����k�i�R"OFYzTM"(;v��3�(j���@"O(6I�/d�n��G�R Fc-D� H��R�p�ڄ+�(}�:��4D�d3�C<���G���/U��fn0D�
���i�ʌ�aM!ZH�ҁH5D�0�^�@�ӏφ�<���C>�2C䉡mD��G��0oJ��� U�.��C�	�g�qs��\h]�$9��Y�̈C��iL�p��lp�*�3����z�jC�	�t�qs�L�V8�ۑ�> C䉆?5iw�	9_�ᲂ�ɸE�C�I�=���b���(c���ڤ��/k�B��H�E�rC�Ѥ+��{j�C��"D��"5�ϓ}U�k�,�W �C�ɞ5:ʜ%�A�U�>ܙ�@Ji�~C�I*`�fD�L���%/��^<<C�əg��
����r�`ܚ�E�g��C�!7+��{�K�o¦H�f@'�C�	�,�u��h_�k��D���Z	h��C�	[Z�Mk�3f��������C�i�����pǤ�x�C�	��x��k�h��[��(>��C�	+Y�IGmδ���"�m�]�~C䉘{�hˢL��t����VjC�I/
V��Q:>�}���X")�B�ɓ`�����B�J�d�PA�6CTC�	M�d�'bC�Z�^)���b�B�V��ܨ��Ǐk��p��I�bC�	�'Y|q�� �!��8H�Fܩ	�VC�	k�Z��Ʈ�,J(�AQsH[:R"C�ɖN�N�ō�AB	��v�C䉙v���a��8l�8��A�{RB�	C�H�0�i� jZ�d!�*�,3B�Xt(��̝���<�D��)�B�ɝt�Թ#�P'6�D��n��� B�I+�t�'AS�Q�$9��Pi�B�ɹx�}R�F5HZ,a�6���3��C�I�.DͰ/k!eώ*H�K��=��ΪH�C�{���g�8(�D�( �q˷O���y�g� >=t�'�Y�"�,0�G�̟_z��K�\p���>�q��'X��
Ҡ�/R�8��/�9�)��_Y���Һ0����BA�\�SӃI�%�$�+CHN�.�1��;4?�����z4j��EA�����;;��$���Q�O+H�#B�T,�8��JA�~�VI`��H�(�`H#��Л"S2���-�D(<	p�Q+g�%�W%�V��XcƔK}�MY�(����5$��3�T�HU2pڜ�2+)�S�.q���o��+1,҄ Y�T�B�I-9 �J��4U�����"Zz���c O�7dŁ�9H6�%�>��ʂ�w�6d�'8nlY�:�YzA��He�IA�bQ����e��49-j2���8V:�"�̈́;.�3���"���%B-4�T����;O$�)#̓�~ep1���]O�(���8Fj�A�Q-	%�1	�t�Ǧ@nZ!Q#:�%;��AhD2��5�dȗgM
�L�Q��Y��j�0��k�Q���P�.[j(�|�7�L �T�iEL��Q�ҟ.@@��IaL%F�<`�Xx�"Odu��? ���c�Y�`�\	�Cȗ�8��鳡��8y�z�Ԃ<�ne�8����3'Y�e�D=��8��P�'�4KK�A���%���#�'ф��8 zD��)ET��(d�;J[x@ړ�F�z���$�GȠ��%��<,fx�wk+AS�O�s���?Wײ� �a�@��`��	�b�<��G�[�" ����.����Γ
���T����]*�KZ`���K�/E�<y:�n^e����B��U��9�N�I���a��@%��f
ޭ� D[�jV��n�T��	1& ��M�V���e�A�M��|��!$$A!�m�y�<��=3��C�O_5e9��!`\�48�cC�?D��IV�^��%{�aR��J�'�h�H��x޽:!Œ �Z�zG��Du	2&6�O���Uj���� �-hcmW�
%^���K#.M���Dڂ5�|�����-C��I&���&k̇��O�p
VAG�-��1�dL��|-D���ɯ}#�x"&F�+������z!P��72���j��]���pQ�εZ��6�i��K�@@2(bՅ�h���;v)��^���8�J&8K.���<a��x��IP�zH�Cd�k���'EE`�n�';N*����z}4i��E��R�����^].C䉽��aر�ǅa�X��V�>W�>��0��Xt@ �,mr��{5�Ӽ
��i���<�o�9̿S�^�,b��:�!�>�^]h�Z���=!�.Շsq�����.F`yD�
fz|аW�P.U90Б6$��E>ލ0&��D�.�x����ûS��sca¨�nH �(a��O`�:�l��q���&BS��HP���S�Z瓕��Dx��T�(�d�V�I�tC�I�&�=�/�*OVaQ�I@$$,Qs���/�<�rP$V�
l±�6#��?Qλy�Dxk�*��|��A�w���V��X�ȓy�"���{�Z����g9tOQ>d��M����>E'h�A@��i]&o�X"<y��/7�>XH2n��?���R��_�����,L�*?z�)dၬq�Z`�3��Y��i�Ή�DnFJ'��=��q��kOQ���u�֊=d̐�*Ǒ~��Q��1�I�9�,��+�w4��Q'� �"-��NA�|�W�/fʒA���,�]
E+�_�<����-w �!�EEE�&�p�y��țt�ZW��]^@�:�߆���'�缃4Jۉ)ԉ�s^�_�Z%�TjS�<�� Zr�Z����lˆ�� 8�!0��Ÿ^�THq����j�'�HOލq��=Y��k�	1Y�D�d�'��#CJ��@��-�-d��<�G����:ᡎJЎ�R��#C�_�T� 1eC�QZtEr,� [hd�Q�ŗjLU�O���h�-[_�0B�"
�lJ
�'w�xk5�ƨ!�����&%�A�)O��F��.��8�͆��ȟh4�`D=$���C�"<�Mp"O
�2�+M�Jz�T�����'m�2!*v��|�]&�d a�����g�)����Q'C�%^&����\K�|���)���Y��V&&,J���� ��'�088�bC��a}2F��άp���
Oㆥ�O���p<1��M�L-2�#������P�b��ӡ=.x$.Ѩp�!�DԈ�9� ��j<��Q���1O>��h��F����TJ�ޤQ+C>d���ǩ�s�<�`�ր+��=��n_�zk�����׶tl	�=i�+;�gyb�
"M ç�	`4�㲠��y�S�:FX���,�3e��c�L'�y�,d6xtnǏ NN�� B7�y2n���ST/�9sf�Q#��7�y2�Ǟn���Gn�8�bh��yd��[TiSካ[!�I�D��,�d��m�3����@�`Ь��ȓu����B��B�qA�G������]0 ��ӏ#�"|y��6}����:�,�rG��q�9�4�S6�j�Ey"�;�(�F��N�-+�V��c�r�	uoA:�y�T�EtF��!'�~ Aũ�� �J�p��8nyzϧ>E��'�qS�HxO��ۆ ��ō"D�HIS�_Q%�p��P"x��aI�Ozx�uE���d�	ۓ:�m颠޶i���
EN�&Rd�R�4Dr�`��8��6f˧jԄd8d�%�2�kD��ZC�$[HQk��Tf@PQ�L㟐�!�!5D������i�@	���F���K'L�'@�B�ɔkw%��)�1�
�P�
��k,�X����/�lE	K��E��'�f��F��4��6�U�H�@��
�'�ry��	i�\0��Y�5�4ٳ�h����VJ��{����
�gP�b�P�E�8�tbĈ;/�{2�2M-R������)ŀ��qhh0{����BV��)s" D���퉀X�ؼb��
v�Q�
<�	=KpN��#)� ��>�P�a�G<H��R=]�!r"0D� ���&z���eꇴSۂ�x�O0m��I�HN�)��<aV�	&��B���%�8����T�<Q�#֥\Ru"�c�>�P۱ DV?����2���U?8�h�(���,_�h�Puo^"^!��5]������pC&L���nn!�� ���r���enur���&c��U	��	�A}���b�S�J|�@���=;�-�5�Ȅ6�C䉆vA����-�13�	�F�Z~�mxW�˘�%�"~�6Ј�H#���8�|��$�k���ȓp�9Ӵ�P(&�ܤ÷N�a'���3L��ZR	;}�a{򨈁xV�P{��4a��ccK���=QSƏ�5<�d���hӎ�+v��D�>����1�h�t"O ��GOX�`iP�@��X=�&��W*ќp8oޱ�H���L��=*�z�E�*R�z�"O@L�-92�Z�#M�pz��S��t�ܠs��`��-�g?r(5J�6�ҥG��C���Ch�Q�<���vN���0G�d�t�`��䟈H�ۋ0�h��'V���MF'xZ���_+�%Bߓ���P�^ GR�6�V��
�%ģhEpw#� �!�26���Ɉ<5��0b��Z]�O��!K˚fj40Y�����aϺTJ�`CFV�!�ď�I�� R�M�<<Ԅ<蒀�;�� �t�O!wچ�O?�I�4�r8J_�0Jd�pj_8EUrC�	>
�D��L�C��U�p.۬V��	�g���U�'����˪_��]���*c�N��'��S
�!_�8b��\=o��@��'1h�B��_	 ��Ξ�K��
�'�X��աȹ�x阄�L�Mu,�S�'�j(tc�8n�@�nK�F��'�<P�ʕ�Y)��])-�P��'ܐa��cm�U��oc44"W"O�ᚣ�jn
E V$�%yfpYbQ"O�d�,R�WW���ΣI?��K�"O��P�A�y�P�bs�SR��q"Ox��Nԡ*D����J�̨�F"OV��'�K����ٔ	Z^|&�W"O>|�Ah�5S"�s�BB�1���"OR����I�Zq���[�r͔1E"OTeQ��L�Zl�aPvb��J���"O���Jވ90��GꙂ�VX�"O���6� �ej�d��"�"O�1�HM��޹B/ (J�*G"O�����"V0�"@�T;�ɢ"O��)d���O����c)"sr��"O�Ԙ��ͱA�h9(S��e��"O����$��2��Q3W�[�Ra�"O��3��os��u��U\��"O���q�ƼvPP��t�I? V�S"O��2�y�8��Ά$N0"O�]qF�F# �-��A� 'X8Ja"Of������2��(zp��"O�������Y2�����-�L��"Oj���b�3
��I�kG?|�V���"O�<J�j�Ac��St'�v���#"OnP�Ed�;��ঢ়��"O]���+8�^���4}�t"f"O��P�K�yx8�TfŮ$��$��"O���>0D��&ѺXl0�cf"O&�!\�h�p��.U�P��"Oq!l��K��� ��$"�5�v"O�Q;D� h��B�B-,���"O0�K�̂y��|�
�#E����"OX�Ӆ�
2"-0��&xp�
b"O�BuOE�'���T�R=e�p�"O�,�b���A<S*��"OT���"i+� (�&5:���"O�j�®g��TˇA@�Xٹ�"O��{R��n9�n�"0!���"O�e�@�ՏvFDm��$N��0"O� ����㑩 h	���?BF��q"O���#��W�������M���T"O��K��`P�Fϋ'm'K�"O�lx���i�ɫ��%y�"OQ����6�ba���Ȣ"*���B"O}�5�ͭQt4=��*�\f�$��"O^�jd�ʞ	 �0
wX��!�"O���S��S\:�wj�&_G&��"O�E��G�i�4�C��+B (�Y�"O�C̈�^��1���cq"<��"O�P*3��<q  �R�Xau&8b�"O�X!)�(o���`��}a,M�q"O�aj�.��6��N�B���Z�"OȸA��]"e����-.S~)��"O��k���!��lKEJ��2`"O��C��Z�P�4�÷1\�5�W"Ol�J�	T%\�s�Q�mI�D
�"O*���O�F�hL@������U�"O�� �'��P����aU"�*p"O��*�]-v�P�������"O�9�MX�D���;� ��vz�:q"O�lJ�Ε�!��a��P�T�1�"O���O�7Xz�j NHGܐ,��"O�X`B�U�;�`E��dхg����"O��3�c��?{��{�eP��8�CV"O 0���A�/��U3�U�n��A��"ON��ख़3F�ȱ�j�'{O���"O@Da�/IT�"�1A���"O0����"gO��q�	�`n�PF"O��uNǟgF~q���k�:D�"O"���$��Dܰ�C�$�xF"O�������)c=�&�~��eZ�"O<�jF�Ό!��P�@&"���z"O>���&��T�l��#K,`�z�"O̥�r�^2�1���^ Y  �"O 02M& )�\@�a
 *`�+"O�8I",#e&`����Vd���4"O�,��.ҧ<tM���e�P��y�J*J�\b5�ο�N��7���y"��z)6�p@�Y����qW`L�yB�ƌ
MD����ƚX|f�
��ި�y�F�.^[l�-Ƃ$X�� �y���/`c8��U�=h�	!n��y�(M�b��p,4U�8������y����1�`�+Vʅ�A[�A0M��y�iĴ{f8	;���:m��b����y�o�E�|#FÎ-��@��Ƅ)�y�A�8T��C`��-C4)4����>pY�xr(V[X�h:&L�9�f�b�+5���f�<�O`h�co|z"a�1�hu��W�Wl����NG �Px"��%W�2��wĔ�#�Aᕯ��hO���)�/O"���(��:<PUya ��DF:��D�ׅ2�B䉩mg��2E�҅G<j��8'U��$�(P:u(D ��E�l�S�OS����ڄ-���Y�oVD��<j%"O(����"7#6d��dϹ%�$iU�����א;���ԥ�T����c�U��P%�L�����A`+�O������j7.xyÃܚk�l�cva
�e�a!��49�C��&-�Ț7N�)o||�w�"R�r�=��`ɉ6����䉊^�UЄ��l:`曈6X�@`DJ�`�����&�V�<��׷W@*�Lͪ'	�1"@.�̟t;Ł�W���*Ҡ}���1��.��IU��(�O�0+H:��8v(P9i�1�'3b8Hb��rV.TeB_�J����ɋ�(�B$�S#�ɂ�	��B�����o�sW�i�l��&�^$+�/ø=x*�r��D}"��q�.L�b̛�v�f17�� $�T0S��\��t�B�J�HGdi3�'I7�,��Պ˅)L����S�? N�h���Ze�Q�M��}�x��O����-iZ����΀2#F�b�J߭3۪��V��=� �Q�OL�<`�R ��T�Uh� ��Y��'�HDR�$��s--|��p�6�K�rG.}cAB�18����
O5n�T874���Ur�Mϻdb�:�f���`ĩ���S��a���#d�~��5
N��D���ÿN	�8�VZ�,N�m3*�˴P� ���I�f}6p�q�'$�m:��N�f���Dd�,QJQ���D��%#�]Ze�d��҄$�SH�	��m�Р�Q�Ry����77ћ�A��@j6��\���RG��9G��:xjqA�J=H��B ܸE��9�'�g�j��4�ݮv��<��8cUc���`��;���s#���e��I�/�T�!��G4+���HŮD�r�H@CI �jt�i�U�D�GHĵG�<��LG5*���x�^�\�����u�G�!p��ɂ6� z�9:Ǧ?�O<�ː�P;3�6��sC��v7� 35NA�p�:�Xe!��︌k��2W� �;W�#?�n�d�ң<I���?n�:��	�dǲI���,�(���Rj��|ږi�E*S�U�­Q���Tc�*�F��``�t��[� ]��y�kS9jM�10F	�&���@gS�S�8��&���`�dE�!��7z.�I�8��O��nՃVe|�;4N�"4��B�%�!�DZ�=�0�s��
�r⭃�������� �ґy0�+!�.�@�O�:�#��ɆX��ݱ�틘i�.$�u��"7�����B�Z/l "��_�^��5�C���4'��B��A�ଢV(�1:���B˒*�����C�&�	Q��-�Y6,x�O�9����0�Pe:�"�,0�c@�2nZ��S+E~Je�r�ɵku�Qȕ!h�B�	��H�YGaųe������A�@��-�wZ��O�~g�2����Q>睰D���q�R���pf�o:C�uXU�ЊƘ@��蕻 �pDL�v
R]���F�A���5�M���F�'�f���U�H��]{s�� _�0���| �B%E�'(K��6eE87r$[`$ ve�L�D��oU^����%)(�9���ݜgx�؉�a�~�z�?��q�����b��'r���֥C�jg$i����-s����ȓ����)L�s0N�R�L.<��|�'7��xU
ܖ6��	�|�O�>�8@��&K-�I�g�C�P�����'��A�V��?��x�!�ۓO�r�h*�m��	Hْ`���Fp�3��0$��0��ǭi��$	F4C��0%���yN���i�.h��L���@�����(��>ɇ�YM�i�%��:@ʝ�$\y8�0	��ׁ=M�'��H}�b�)7�E�Ӂ�!_�(��1�yB�g�f�SKԷ'�6Ku��ݘ'�2c%���\5�?9QC��J^�SD$�;XP��q�!D���f	bP����ƕY�er�@ Hi�➼`��<�u�ځ5*RjHy\]C�E�{�<�CϭWX&{b�9/s�L8!��x�<Y�i���@�	qA$|���!�t�<��
�e��d!�
U�2�1C��]�<	�`I�J~2TRc�_ 41�T�K�X�<iƍ�	#��1 o�Y�@ ��U�<�V�@&p�Bg�=@��!�k�<Q���9�X`��3T�pt�D��i�<���x�`�1%��@F��Z���e�<1e�A�n��0��Ǻ5���J�E�'��Y E�i�O��[3�#ZM~�s��FTd��'cT4I5Cu󚌹v)�3�Z� EV6��@'�|��9Ov��q�,{�l��m��U2Z(j"O�e;T�C߀E��� 'p��P�'D<�q��(�
t��	�Ri�U�C�Ԃ�Xy!���7���ĕQ�,Uq���M�PE;`϶ q�F�{��M(c�XN�<��Ë9`1!k�!%]��׉�J���4�8�ǚ
v"}Js�P�zG��`עQ���k�N�z�<�E,��o�)��*N�.�0�C�,��_���0�X����h��d�5rA�dO4rjУA�݊N!�D<uъ�`N�kgND���2�2��<��F�d؞��v$�4H����=�B�@Q5|ODp�j�
�\���4|����'�%c�xM@`[�i�����؈$q��9;���e�
2��?Q���0�	a�$0�'a��;fm��0,L���Q�"�ل�$V,��v.��4"C�P<X�z�KBE�n��1�J>E���� �zP愱;���s��1h� �`S"O��{t�Q�UM�I)��x�ڬ#�Oإz��9�0>����X���f��@1F[�E�W�<�q��	x�Dtꀩ�4�B-K ��P�<�bg�4�\Ͱb,Ü5�f({p�T�'6I�B'[J�OOdh#�%��qZ3�A�!��
�'t8E��ݻc���b&�W�t18R�S��ԭ+֘|��9O�P!mؔ��|c��'3� ���"O���0(�y�*���(f�D���'����O�)LZ���I:��HD��Ze�2E˗V�F���U�([�T9u�D;�M���+R"����	$�
d�&�N~�<��'Q�!E��z VdQ+�}��M'dMۧ�� F�"}���S;}Y��޻%�U�B��z�<�M���	��)��R4*�f��P,��Y)�铐h����:y�ѱ�C�5@2vI�w@��5%!�D��~<��aT>�Y�7�6C2I�>^� �#U؞�°}~ݒ�b��"e:�Y�,3|OB���R�0�>��4\��t�e(̪V$��P5_;DB���s �yD�s�f�pt�N�F@�?a� W���(ҧD*D�y�	D�T��!�sh�u� ��w���!��z��4BӮL�j���{�����2�O>E��'`Te0ӏX�n�<X�IX Z���'�f�9�"(R}됾�e�7!b?	���U�8��$<nc��2�_6��-�"� �>p!�d�)�0H �����	���֑e!�J"��)���H�V=��� x@!���xI�@���/Aod�Q�л!!�D	�`����(!E^y�Z(z�!�D[�o���(wht=B��J
��!���K����f�~Ml!�d�!򤌲B��,D���^>�)��@= �!�D q�|Q���C���rA  !�DQ#�6��A�)/�tB�a@�uk!���:Of��Ģ��u�&9�!�+6�!򄃊h�2���< ������!�`n���%E�wzd�z��ӷ\9!�$`� ͘���.Q�D҅�|�!��K�t�½sB'�2g�zde�((�!�$��&셛��R4l��`e�E�!��8�*w���rD^�[��ߎ�!�V	}�hQAGM���tx��a�9o!�]L����%.�*�DJR�#v!��P��L�|"h�P�Y�t
!��,����P��%�F�@L��i
!��F�a&�i%�Ź���+%,_��
�'�e2V�U2p?�����Ɲ``j�
�'��	գ�����1�ѤâP��'�đP�/�)�z8p�eH)j��Q)�'O���Vm��&1�e� ��#k�V��'�8Ar���6�y� eJ���']fp�`۫x�<|�f���"dL��'��y�'t�����@<"�x��6�
�b%=c��FdВ���*�~)�ȓs���֨I�e��S�j�@Vȓ|,��$A�&'z��bo�G��ņ�z�~*���C��TB��K�<�ȓ$BƑ�1m� �� N��{-P@�ȓD���I���>"¦U�,�;|�F5�ȓ9�|�C�]E:�i��\ɲ���9ћv�<��q�Dʖ�����a͋��ɭ*811!�ڗ-����3�'n�T(8V*J�%�1��.
�GCb�'��@R�Qp$�`>=CTk��3��!㢀G9�x�ãóD��}1C�^�.��y���<E���Oz&y�C��.X���i֬ć��l��Gҷ>U:튵�f�H6�\���? ԩ� Y�N���!!+�q~d|�b�*n�a�ܴ7%f�I%��L>� �H@����HA�պw�	fD(H�̈́T���	-{����qf�4,��?�'p���e��A�𐚥
��)#Z�
�?On�d.O)Y����"��l�O��@�����X���]�d���ZufՀ4^̈��M�N��!@���.�?E��43��$��� :hJM���k�\�Rn� ,����h��	P�L>�'L�T!�A��O��T ��%-,��DkUB�I1%,.����~�u �
� E`� '�
�j��JG�<��@�[�"�{���&w�����đ@�<9��z������E�s���4
Cy�<�n��a����Ak"�7��y�ˀ=�"�����*�����ŉ�y"�O���F%ԝL��uSLĳ�y��ݬ]b>C���=�d�a�Z��y�D�.)Va;�P<���Fn�-�yR�R6Z��G 83-�)B�'��yR� ��ȠE�(� \:�Ώ3�y��H�w���sfh+J�����N���ybC� s��!1�_�:l>����:�y�$� TX��?:O� QC>�y�B. S��z��_��9J�d�$�y�gr��4!#�֢^7�`BX�yb�G%#,�u�J	�[��yP�����y�˖�g-�L�7-�Li��P�JL��y2��{�[S�E?	X9�D�(�yB,ȇ"�:��`ȯ>�����>�y2�ןc��]h���g���'r� 0��ӓ
G�麳�M=b3�Pq	�'��H����sjDs�E��*����'��{5��_d(��1xA\M�	�'�4E�5k��x&�QT/Z�B�Z1�'��,0r�Rش�$��IO]��'y����k�4�d�2��[*0O"A"�'~ �2)Q,�Qꑪ*�"գ�'���
�
�/k��Jw+A %D��'��@�"V0y����`����Q�'A��`��[����&��z1$��'����Ғ0�v���n��uƖQ�	�'�U��C���r���<���'%tL��� }O��)!�2�f��'�!S�nׯ���+u�_%&�vu�'Mh��3�ҿ��H���r�Z�I�'�����;��JDOl�r���'�r!�	�#���aGMk-��a�'�T� 3���vvpP���dM���'�zh;��ޱn�� p�	]]����'�\u��,���0��!�On��'q��A��մ9S@1�a�F�(�a��'.��S�1w�0��n��V��'����2��&we4��6�^3Ֆ��'
ʀK@n"g{.@`�ȝ�8R���'�֝�'	�����w�ʔ�D���'\�4��ҁU��I&�M5(ul�S�'� �4��OL2�#Sb݀$ծ%�	�'�hh���9b!s�N	'!�|�	�'1b,#�Ɲ�'q(��T�Ų���2�'�vTbe^�h�hԋL��-��'����ǕX( ���^�z~���'
�㥙�,���'�V��Xih�'p8,*���jԘy�!9����'���4���A�ҁ��\�z�T��'�ȠR/��[�V�����)�$�)�'Ml�)w�Gr�.��b�W(��'�� V�;VLƙ�h���Lђ�'�Bp�(cP���m[|�"�P�'���A�*Y�C��l� -Q_c@���� *�zR잙���j
ë�2��"O>��1���SZ |�eHZ�6��X�"Ot�����WZ�Z�a�Mα�"Oq�&E�kdJ �^� s"Opyؗ�T�S��%oJ"=�"OR��/��[AFI��N͡~��2"Oh�Ƃ�.l1L|�ƌ�!$� �p"O}���UC�R5�cK��Ұ]�"O>� d`ĩ4�X��`+MY @��%"O�tyuό+c�^����݁R�"O�i2'
/1�}�Ňȣ;@��"O�!�և���p�9)o
�r�"O�h��B���ڳg�<,(���"O6�	��W�q3R&���Q��"O p�peK� {�	�ޖ�(�~S'"O�d�'�ԎK����i�<��0Z"O��KH�?��K�H
�9
D@�"Oެ��`�=tԠ8EB�x�h��"O��
�m�"g��!�u�C3u����"O�H��g��1뤄�:��R�"O�HZk�	tdcv�X=���b�"OYb`B:��:P�v��`"ObicRaE�y�.!1�iY�b��%��"O����GÐ}���'�-ږ��a"O�i��Ƅw��@�de�5c�vը�"O���0��{����$�7�<*�"OP]p&+m:��jWCC0�$8�"O0��`�<�J�=�tEK�F΋�y��:beD��g�� W���M˳�yb)�ۄM@AM�zp�3gO[�ybh��x�a1��eP��r���y"�ț!��u�aF�23<}Q��y,/F�4�� �ʴ5��H[s���y�P�96dr�g�h�Hs�Г�y���H�X:�IP���i"�[�y��>'	�e[�H�s8 :a����yr�����I.�.E0ZJԭ�yB�ـ[B��!�͗r)D��`o�2�yb�F4[id0��K+d���Wi���ybNZ�Fd~�����VXp�3�2�y"��49�xl#.[;P�"����X�y��+{�H ��C�� KC�
��yr�V-1��[f��>�΍�u���yB
�"kX�QI˲2��Mqf��*�y��ؽ>���W���$ɪd;Ƈ�y���&WDt�@E�&g�H��#�y2b^
h6f��u&N4u rU��y�+�L��iy��D"�d��$�R.�y��4]eb,A�A�L�^}� ���y�!f�
U@Pc��/G.�9J��yR%U�l��U�-<�0Y�׀�y���^�]��Ť7B̭�a�-�yr9�� $!ް�	��y�Ҭ�&�	��a0��y�W���x��ֺJ�М��h*�y�V$��5i���<ۼ%�����yRRc�l ��kI�:�X%RTս�y"E���H����}]DA��kO��y2�-E���s%«} #3�œ�y�f]"?�°X�R�y��M�� V;�y"�͌F�^�J�
L�d��pAZ�y���}���>f�@x ��!�yBIU?���*���	cp(٧����yҥ��x����'EՌ[��i1@�і�y
� &I� '!-�� �j�� Xl��"O.Q"�&��OfpL���� <�r��4"O�����,Y$�	�Gir�"O\�ʗ�B�����!�.M��`;�"O�`qd�mk\)��K�p�j�hQ"O�x�aC�7��:2J��}8�H�"O�A��&�̲��Ӊ_-b���U"O� Ĥ� aC�� �bҏ �ؓ�"OR)�E�_��u����8"|�ay�"ONhp���8a]��r4`��7�@�!"O�P��+YE�68�w׋6��aqp"O���$�8g���0�Z g'�\f"O�-���)�-�n�X�e;t"O��x��ë?=0}!���&咅"O,\ȁn\0]l�Rf��5L\�[�"O�A�T=Yd�0��k��W"O 쩢��_`�a��'��=Jb"O�L�b	���UJKnuHD!e"O�If�<���È�m �pT"OXX�� ��y\��I�4_:��a"O$@:�!�4a���@�(Ǌk��@J�"O[A�ܝu��,�g�!g�B���"O��xbG�"�����w�u��*O�Q�����r1
�+�"-a�'؍Hc� aڄ� 񌔂 �RX	�'L؍�� �X�p�!��.�����'���Ч�� ���bOP�u~ `�';�O�A8Z�x�i������'0��*�oR�/�8���犹H(��s�';&9�.�0Z4��h��Rl:j�"�'�2�6n@	S�@(;aNeg$|��'�>(А߃EJ ѡj�0��!�' Ȉ3*��t\lh;��͓*�"�'��9�'nŝ)��l���S�����'@���b�-<`��H3O_>�(�	�'�~�: �Ֆ(ؒ��r���m��{�'���6�	3����b"�Ps�',u�mǡ ��!*���S�:8B�'I�)�f�ߢ����p$��K�����'���:�$=�j���̜�s��0�'��(ց�7Si��@���f���k�'yq��!����Θ�,=��'�p�8��B8#<΍��@ye�	�'8�p��"w3��2�ƚu"���',p�2%h�(s�i�nx1�'xV}��
��C���	��Xp��'°cԉ� dx��a鐨>�"8��'��5Kș/4,t���	F��'�^����G�.F(P�KK;J��x�'>VT{�$��x���g��� ���
�'�&��`2}�-�L.�u+�'��Z��XJ$r,*��@�?r$0�
�'��Li�O:/���1& �==%R�'���j�k[�G"ΐXuj?0e��
�'�މ"u�H3>4U�d�K=`R`i
�'t��1)�������P<�d�x
�'�n ��J��
9�YY���A(�A�'R8��g'ǭu��`�Ԡ>x��'�T��*�Ӡ4�&��7�����'�IV�"$<��lP>5����'yR����,CV��h�9&Hnqk�'�RQ�)�4)���[�̍u�"�#�'A���Q��*��xY%�#�(@r�':����	) ,����&69{��� �F�U�J�B�L�9"OX��)� �4���H�"2�0�KE"OD�1����ʂ%�W��Cx�;"O����  �#\��v�8lBp;"O�}k���2i�RA�V�Ӈ9�Ĩ��"O=�b�����`�N�f����"O��sS.'��Y�T�EE�BR"O�Z��_�`�L�ȅ� �E����"O~��E��n~�8r-A�9.��cc"O�����ڵQ�>x��KI��B"O�����QvT`H��<SϠU��"OxLbcCN�F�.�3��n�J���"O4"��&�F@K�Z�`��c`"O�Q�Y�H�ƌ����?�֨�"O
-#"'^:o����`e� �"O�ho�q��M�9�L��4"Ob�Z"�>�	�a/�X���F"O| ӆ   ���M)99d����'!���"O8l���ٔz����WÁ����"O� ��H�~��!ϻj�"��"O�c�̓�h�T-c�&H�|o ��"O��g�ܷK�� �&˦0f�5yw"O��S�Oײ0Ӡ�I6&�(�z�pB"O�jaL�^U��@�|*ƨ9�"OnȨ�;]�:�2 *X����K "O���İe8��� J��M�Vli�"O��{W
��Jz:���6)p`��3"O����O�m`�,�,s>ҥ�%"O��	�-A�x�vX��S=���*OI�D�X%V���C��*1!	�'����b�^5�d��W�iޠ���'��\�  ���   �  O  �  �  f*  �5  ?A  �L  �X  �c  ,o  �w  |~  0�  Ύ  �  `�  ��  �  7�  ��  "�  r�  ��  ��  ��  1�  t�  ��  ��  ��  f�  � � � � q! �) �1 �8 =? �E *I  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(��I|�O���#�H�R!��њ]��p��'_��uʆ�vӲ�R�c�*m�'�*L��܉�` ��ڭ\�����$֮w4I�1O�,��g�W�b-h4��Ӽ9�HMB�tX���;%�2���IЦ�Fx��2R^zmC`� �p��#�ȵ�yRO����!�L�q�tR� K��$"% �"|���6U3��B0)зez��%�~�<)0��.)�#U��4��뵥�T�<��۞@J9������
�ĥ�F�<���R�}��%�	2a ��`j�<�d��W��aP��ۆ&Z<�j�g���'o(�TA0g�]j�ȺS�����'���G U*=�~@�g��J��p`�'X���	B�z��X3'�R�m�4u�	�':��D�K���@ W/�S<������ �\q�C1������h=�A�#"O8��N� Gv����^�g �<#��>���tl@aM�/Dc��2X���ȓp_�B�"'���BQ �萄��N5[�œ�J�lU���V ��-D}�����Q��*�	��ȴ�� �C�I�qv�d��+̅Z�����슃'�B䉌�����"� TU��gɭ 6#>��C?�'w�6��![�.v���a(3�i��j�X��`	O̙K�aX���YΓ�hO?!F��*e�@y�FP�@�XɫA0D��:4��(N���q�S�/�����,D��z�K��U�TǄ�'TI�9�+$��g0��9�� �:�����o ����9P�M���4t\�\����ayR�O֒O�0���xb�Ӷ���V�{�"OQ4�B�|;z��&T���S�pG{��	�d�\@A �K���)��/�!��>P� L"��"GBi��&K/}�ttFz��9O�I��rL,y`��hX�xp��'��+K�Q�����T��������1��]m��<)�]~��ʆ�&O`�3�X'>��1��	k}�K>!B�;q@ηn��l����yRaA�90�����Zcz����Y���OL�~:��N�8aޜ�A($}�q��a�c�<��R;/xВ��E-�:ѡf�c�<Y�Y0�����j��u�C��i�<��#=uL-R��	�+($Q�E�]�<񳋟�%D��O�g��,P�I[�<��g�&�:�r&l��G�.a��&A@�<6��_N^�R��:���� �y�<�w�ґH�yz �3�`��� �j�<i7�}�2٣QO�p����2��q�<�5�̏�xq��T,�s�F�<�#��![����UN�t˞�b!W�<��k���≨��Q &Р��|�<�ƤS��ڑ�UF�JIj3�Mq�<���ߣ��� �M�1vN�Y©v�<�q#����g�)��!��v�<ag��R�F�� �>���Вd�V�<�����Ttހ	�[\��,3aL�i�<�a�C�2��-�I��T��x���F�<q3 �jT�㶦ւa�j0I�~�<a��WB�<�S�	?sC����j�o�<�"��P�:���=bJ��&��n�<�/�"��ړş6K2zD��c m�<�6�P�*���^�B�ވ��ŋ}�<I���1�0��#�3c�R͒��LS�<�$o�^ľQ�ԀR;1�:�Ns�<�d�)0��f�g�����/DG�<i���B���UB_�&���SFG�<i���b��C�Hܭc�����<�k��FWL�#�M�%j(X�FE�<�ä���8�d��&J ��DoV�<s�T�\���9�2M���Q�<��/	�P�RfD�<��l�F��e�<���G�#�H�1�K(v�d�4By�<qB�"J14Y��͏%�B���t�<�PHZ�:0v�a�U�E��!Y��p�<A&	�W�� ���~tb|��o�j�<Y@��.k�:��m�9pt
Q�5%f�<Q�4F�(�3�����k�'�F�<����r��t��v�J�{F�{�<!ݚa��	���.����d.�z�<� v�B_�0�q�� �f�2���"O�}p�4�V%Y7b��i�!("O(h�`�lB���5�B�	��""OJ5�f炖l��1��Åw ��Ҵ"O�IȒ��&$.i�Vo>)#�ı�'M2�'�B�']b�'V��'P��':L�Ye	�#?�T�*�j����ͻF�'���'���'N��'���'���'��q��(�.mZ���x��1r��'�R�'���'SR�'.��'���'�:�`I޽f��PmK;�8h�t�'�b�'�"�'?��'b�'���'���# ��4a�R�QB�Ɣ�f�'}��'���'q��'�r�'���'s.�[ukF<7aq����`%6���'���'2�'��'w��'/B�'��p�D܊o6~Z3�E$#d����'���'b�'-B�'��'�"�'�8}�#ެN:�J�MI�?	����'Q�'��'��'b��'7��'B���
I�s�t���ع5sx����'�B�'"�';��'/R�'�b�' ��J]�<�K��ӧc%tQq��'��'0�'�"�'*��'/�'�b,!a� YH�,ܲ4��>�?����?���?)��?����?���?���� #�d���B ;�
1�A��?���?i���?1��?y��?A���?�r+�
�\��,O=4���+� W�?Q��?���?����?9��k��V�'���Y�i�"qR�)�	�~��5ET�3����?�)O1��I��M#E��(���h⦇Vvb�S�"��'��6�.�i>�	ݟ*� *���	%K�*$*)�u�����~ �pn�j~�6�D��SI����#�l��"�D.B�"����1O��$�<����F$xg.����,$Ft,PnƗ}�oځY��c����S��yWl�#��XbO� ],��I=���'��>�|j�kݯ�M+�'>���1�G��T�P�2Gz(9��'����$s��i>��I�dpi3פ�+�PEZ+6]���vyb�|�v�m�r�$D�H���rωD���d�����v}��'�6O��'��P�ԖqfD�F-NC�H�'����p���i����Dş�i��'x0�&(d�s#��c��u�QQ���'���9O 4�7��*K7�8��F�.�  "�?O,�o�3���%כv�4�>�(q#{����́7���ڴ;O<�$�O����V�6#?��O�4��ĉ*h6�Hc��qJ�x2�F�@&>͢J>Q*O��OF���O��$�O���C�K�8��E�@K��v�H��	�<)�i�t���'r�'��O�	Z9R���Jf�D�S8Cה�@V�fE�O:O1�0�0q�Av����+S-#�н���{H
�W��<a���!y���]������>׀���_~�rуr%�.C����O��D�Ol�4���p���b�!d�!	1]�:4x�L4ځq����y��`Ӻ�L�O(�o���M뀴i��*�J�3�(��LR�4�n�ɶc�V�����p��,[�C�������*0�v�����1���[b�]�3O��$�O����O^�$�O��?�[��##6iB��7F�pT0����\���H�޴z��'�?�&�i��'Ύ,��9,�T�r� D��,b�(��F���c��|1�ƃ�M�O��FoJ7 6��J��f[L�Q׌��>��|;�s;R�O���|���?���k�@-h�� (��E�#�^8l�X`���?�+O$�n�)f�`�	ܟ���w��)^���!�힝$�,8��;��$R{}�B~�b�nZ���S���%;~��

���F�օj*��s��"V֠p��O��-�?A�c!�D��6�.��P.Ta��Ѩq&՞��D�Ol�D�Oh��<A��i���b���*��'�n>)�uEO�RN���'�7�(������1Ғj]�e�I��j�_�46���MK��iJP���ih�Ie1�5�OK�'u�@;�ֺL��Q�k��%Cp��'���'�b�'���'��d��u�N	P��ȫw��pg�TQڴ�d�9���?������<��yw皥hGj�"��F�&���@D(��7���I<�|JB����M��'���	7��?�6IZc%�� 1i�'g�<�sO�����|_������r�d�2�{��	>F_T��6��\������	gy�s��E*�d�O2�D�O`)Q���?��k�d�1$%�D�7�	�����O~��.���An8Y��b	.��E�I��v��I\ZX	��>g��c>I�Q�'��Q�	��i��M�i��.����Ο(��Ο�IS�Ok���Q$JA[q,�++/�Q�󬞝9���~�.�Pv��<!Ŀin�O�C�2��j�۹
�6�Rb����(ߴO���؊��&��leϚ�&$���:]ĬXć+9������L�T��u%�������'�R�'���'��e�2Zp�&��u�&�D���$
��Q�G��vy��'�OB�ܣ\����ϒ�p~Xr�f�r���?���3:���O�t��MB�N�^����;��x�i[.kU$x�O41*�"Q6�?�$j>�D�<9fϘ���Y����I�T�v�̙�?��?����?ͧ��_���v��ă��m�t,�~0Ij�H� 3,������M#�Bg�>����?��i{8��ۑm!�IZ$�ɻ^�\i�OXD�F��\Ҡ�	���	��� �t`+T`K$|���R7>�ҹ��=OF��O����O���O��?A��l_h��a#�B,\�&�(���ԟ �Iڟ�Cߴ7'\y̧�?ya�i��'~Z۔ K�/�.p;Ô/�Z�c�%�$���c��|��L	�M��O��شII 2�&H�oѨ+MR�q�4i��s����<�*O�)�O����OY�Bi�3`s�`���ѕ�:���O���<q�i�(���'*�'��mK��x�,�U5F��r��_~����	Ο@�	��S��.���d��GI�h�>��N��r�i��E��p�O�)͙�?A��O��	ƞ%�˙
7���fC�=Mb1Q���?���?��S�'���妕����=
�4gK/>��9��*E-N��u����3�4��'��ꓺ?)1�ڦ1���@�\�Ђ�ۂ�?Y��i�(|*f�i?�	U�Lp�v�O��'���[1��p� )�8|)>����$�Oz�D�O����O���|���5�ؕ�D�& =$s��������,z"�'�����Ԧ睐\�,H@��p�X�@���	����PyI<�|��Ϟ6�M��'�(��2��1�ƌZ���e�R8��'�XYR�.�韨Qf�|�^������! �§4Jx|�7ǋq�^��fKP՟h��ٟ��Qy)g�dhj��O����O6�d̅5�H���s�����3�I�����O���c�	�P�� h�D$�X� �Ww�H�<y���$���|��l�O���BvN�bL
�[�P!A���-�}���?���?���h����<}p�&���Z%�T�>|>|�˦�A���ޟ��ɟ�M���wH���a�7(�8�� i�;*C�ت�'Zҹi��6�/{h6�0?���+f���.DG�Y�Q .T$x�A�R)$�HL>a)O�I�O�D�O<���O� b] �,�RP�V\긐X��<�2�i��[�U����G�Sޟpq�!����A�ìQbx��U����Ob�Vl�)��<[��a#D����9�cf{\Ms#j�09<�-�B�2Ʀ�Olx�N>9.O|�Z��К����Oo��)ie�O���O����O�<IQ�i�ZL���'��
; 9�t��Ð�HZ�؊��'�t7m'�	)����Ot����ųT�[	0x={g�
`G
���	n�`~2�M)�(��SMܧ��+�c׼��-r*��kB2�c��<��?����?���?!���hQu�@�s� �E"Ri����'B&Ӱ��d1��D�ئ�%�r�)N(mWz���ObB0�a�N�#�ē\ƛ��i���K�	�@7-(?��E�v^6�H�I�$�D((��[�%"Ų�%�O��@J>�/O�)�O���O*� �/�b���	�/I7��9��O����<��i�h�g�'�R�'���<o�� �b�GN��0`eJ`���	+�M�ýi��O����5���=�}sg�0�z<z`�Z�w�b����:?�'���5��4�4���<TjmJv#��Kb������?���?�S�'��d�Ц�c����|���-MtxL�#g���:���'�"�d�����O,}lnb��x$��	Ar�H�p@����4��6�3g������hd�N��4�~�vݔ3GT��(�,h$m`q��<)+O���O��$�O����Opʧ/��(�P��:U�W�Z\� �iT��c�'��'W�O�bh��.�
D��y�O�AP�m(Ф�A��lZ�M��x��D��	[�V2O�UP�C�6q�����mm\30n��<���
�2`����$�����d�'V�U�Ba��@��۶1����''��'BQ��Y�4M��D	��?��<G��S"�O�p�Ѣ!��~T�T؋r˩>����?���xR�D�H\F���!=<��d��D�B�P��)�!#1��X��&#��$^�B�Y�� $#�$��-�2���n���'Z��'��>����M<!��͍�j�DU�$���;�B�	��M3p��(�?9�%�&�4��I�w�#_��:�.�IRY��0O����O��nZ5>��oz~",V2�(q�ӽkZ�噧�ǘD�윒V�F3y�����|bR�������ğ��۟��r���ԙ��@�Ya�b�{y�cp��0�P��O��d�O�������>$B0\x�OC?��� P��PѺ��'���'H�O1�f蓗��
~�b�a�b����ؓ ќ�����i�I��&FB!H~�	tyoڀ0n��VAΉUs��8Gld�2�'2�'��OI�I�M���C��?��H
}
щ�	����bO�<�r�i+�O0��'s�'v�W�"�X@�NS1}V��"lJ� I&X�i��	�)���Oq�&�NܦV zM�k�)&��� u/��OD�D�O��$�O��/�]R�g��.�H"��qN���	͟|����M##��|������|�A��8pE����h=sd�S�(O��n�9�Mϧ(X��4���n⤚�)�w?���!��j�b]0CM��?���9��<ͧ�?Y��?��L*5^�V̒7ņ��6�A��?A������Ħ�z�)�ʟ8��؟d�O���	��&j���;s���,�(K�O�}�'Mr�i'*�O��3MϾ}�֎J��c��#0hPq0E��=�:ܸ�%�>��i>���'h�%���p@����ՒܒO��x�䉈���������ɟb>�'��6�O+�h�I�K˓���9d���V`�)3r��O��$�ަ��?�V�,o��DX�9#dT=V/���QHE�x����ٴ4e��M�|O�V���)#aT8W*��~� l ��J�>Y�:�Zv�>T��1O�˓�?����?i��?������ҙE)f�k�.�=8:H%k`fF�X��l�#@�	�����Ie�������Sg�?;�,`Pf/�XZa�Q<�?��a􉧘O�bl@�i��V�9�~�i%X�<��q�CǛ�N��ןP�M���?t��O���|j��X|p���-J(��q�U���[��?q��?�(O��n����9�	Ɵ ���36��Д�ڽ|�Z8@�(�?�P��ܴk���x�)�37"���gW�幒I�0���ϮJ���4ƕ�f��������a�0�䘪V�g��`���c��	���D�O��D�OV��?�'�?��I6<N����+O�t�c���?ѱ�i-�YS"U��)�4���y�EE�B\�@J�c�&V��y�jdӨ������j٦��'�a7���?�P� 
�>�X*L�/�v�y�m�1��'��I⟔�����	������ߤ|�@��4M��yZ�/5���'r6� ��b�d�O��d)��9:�9��;L�jt��$� Opf��)O4���O8�O�OHLaQ�ٞk����5���|�������AwX��Rsɂ�~���s�pyr�F09��ոD�A]��N�\���������iy�z��	11��O+K��)k�Qt�ԥt�`={�$^�<��i��O���'I�7�	Ӧ�JشK2�݀���7��A��h��\N\�b��]�M#�Oz9�p+ь���D�wJ\%��E�	B�@-���2IJ�pq�']"�'U�'PrT�b>93��(�*w���)���%�_�x���`شX�D��O��7�;�䛎%iV�C�-�/Bt�A4�K$v���$������ӊ6j��nO~�MG�4ζ�d���R��%bX���lYX��ȯ����4�
�D�O��ē�w�Ж��=�F����D�u��$�O��6E����/
jr�'/BR>�2c�<4B(�x�N�W���:��/?ASS������KK>�O���ZՃ�v�(�R�J(+K�P;���U��t�B���4��!��YU>�OX9����Hs�%H2d����@#$��O����O ��O1�>�sޛ�H�	�Be0��]�o��a�FCL�ى��'^��r����k�O����7�0Ԑ�*��Hߞq�s���e��ͦ�%`���!�'h�QU��?�����X��OUdp���J��!�±�;O�ʓ�?i��?���?����򩅑V,,$�sj��YØ�YIY��X�ɕ�2��O��$%�9O �lz��h���%n�|�Q�Ռ_qZ�F�����v�)�>mw��nZ�<��ϟ�J�~�8`i�*H�ܔ�e��<���͊
����L�䓉�4�d�D\�
�ء+��2x�B�*�$�;U��$�O����O�ʓE�����.Kb�'�bJ��B.uQ
I�IN�}ð.�"��OB�'��'J�'��	Bg�}�*AGJG�����O���Vb_�e�Xy��i�?� �O�]sp�O�4cJ�B�6�zá�OX���O����O�}R�6��L��*.�E����K�Dl ��p��V�K&H�剉�M[��wռ��a&��c/�Q(Q�B!����'��7�����4OǼ5�ܴ�����nB��C��2x8I��	j���%hւA������O����4�����O���O����ݰ��I.�f�0�.��.z���6&��wB�'����d�'�D��c�s�a{3�ƌB���S��>����?I0�x��$��F�r2�ț��X�+��hR� ��(�����W"T�K����|bT���8�9A�O�$S=jA@0�G�\��؟�Iϟ�Ny��~�
�1ţ�O��f�D�1y���=D���1O�%l�y��O��1�Ms�i�
6M�<��Lr��<rr��#�b}a��M��O���Ӈ��҉�4�w�^�P�ML4�*dy���'>��#�'��'���'�b�'��<�7Ɛrذ��Ԙ
����ƥ�<��v3��.���t�'�D7M=�䕀2��5�&�T6y��W,��6$N$�0�I���0���o�Q~�J@M��xy��D�i
�b���%>��R��֟����|r[�����I��:��K����DJ�x�d8��R�(��ByBtӺ���O���O
�'u�z�Jୃ93�i�'��/܂��',<��?Q����S��E�6�6�����9���׾}^t�`�BG:��O���?�'�dԹF��1����!@���*֐v��d�O�d�O��ɪ<Iw�i|3���"g9I��4!�R��3I��5�M��҉�>)�1`!Rǀ/@h�!��	]	�$���?!@NF��M[�O����R��2J?�� ���81~�D�s	� &m�`�'��'���'���'p����E�=³oR����i��+�6- by����O*�D0�9O��oz�EAubZ]��W�ū/�fEK�F̟�	A�)�ӄ�]n��<AU�� \ˠ�Ȕ��N�lRam_�<ѵ��E���˦����4���D� 8BU0V��[��h3h�.F$��O����O(�UE�V��H'2�'�o�i��A��\�B�l��FO���OV��'�'��'=RM�r	�8�#���98�L��O&��DN��'z��f���(�?�f��O�J"�?I��x��.8F�Yw�O��d�O��$�O£}��'P1{��Ȥ��) qC�m &�Z� ��ʘ�'��'jz6� �i��/ٔ\�2�0Y6�X3�����	Ԧ�۴,�z|��4��$ǘ�R�1��z�� �dsU"��2.��7��*!��x�/�$�<ͧ�?���?����?���ـi�	z���yTIЂ-��\��M h�ן0�	ğ�&?9�Ir����vE0+Ȑs��� j��\�/Ol���O��O�O0`��p��� �d˥��"Ur�(g�L)$���_�D�e�\�1���Om��Cy�-��2ɐk�T��&�@����'���'W�O/�	�M�wcP��?f�ǸZ(�Hqf�ߵ�����i��?�'�i��Or��'�¹i�6mT�����A	tшU#�)tR�t�e�f�"���U����>��]D���s��_%�n��PjU�t������	ğ`�Iğ�Il��z����/d�E�����
\>�����?!��Lz��nN8��IP�m&�ܢKұ}d���EN,h�p�A��/���?���|JA����M��OdQ" ��>�Rԁ�Z������VQ��O*�OZ��|���?���fU��V�%�Fݹ4��z�P����?A+O��l��(��ڟl��A�h�&	�I�U,͋6QVp��e������\}��'�Ґ|ʟve�Bd"�:Ys��F�F�P�r'W6 D$`,�5R��i>	"��'���$��a�E�X�Dt��iWa��|��ן��Iϟ��I�b>��'6x6��+V��qЊ]�e�x�3�䀨Wz<M�q��<��i�O`��'~"6m]�*�x�6Ȑf��@8�lmLlZ��MK�+�M{�O�|`3Ë���J?!J� E��p�z��[6Bs,�ɥ�x�P�'�b�'���'�b�'t�S�Z
�<�㇆ �����%��_�\=(ߴk��0��?������?�R��y��Qe $�FH=�쵊�'�(SqN7��ğ %�b>���R̦eΓ(S,I�r���V�����H�.�t$�,�ݒ%��O���H>�-O*�$�Oƍtj؇�
պ��X�J�	j��O����O��$�<	��if��i��'�B�'3�q��"T-04,i��)�0�!#�Đ`}��'���|���n��d�T�[�\d1!㛜��D� �� ���7<`1�8��9`��d��d�(��-��(>)xcAK�CMD���O����O��D �'�?��Ȕ�?Z&��M:_���˲fX��?���iU��J��'X�r�j�杈*�B՛���_Zp!�I^1%��Iş`�	��MS���M��O��(&/�	�b��f��IC���7m�D�[�O&j��ON��|r��?1���?��]̸��.�km��Ī�.j�le�,O8�lھ[tA�	���It�'�X�u���s	��K��حqebi3^��Zشdhr�x��ă��`UHs��+LSh�dK�Wz��Yv�+�� ,!^��B�'��&���'�j�@",��'l���ßA��y+��'���'@"���dX�(p�4w��I�7�V���FD,����6��`��)v��$[}2�m��u��������V-p��J<{i�y�"&N�*n�o�A~Z���c��?�Q����wN���%� �	�l$(��Ƹ���'���'�"�'a2�'��ѓĊ�m_D����[,�c���<I��xț���9��D�'�t6M?����) 2LHDN�	ReN1�S�M20���$�r�4:˛��O��-R�iZ���O�����Vh�ur�G2�%:�`�%%D���'�ޓOH��?���?!�������!f��Ux��˼^������?a/O�n�>��������Il�c�'�}5�W(�#4�ҝ��$�E}2�'�2�|ʟ�e�pOI6a�&���L�;z�5��[&!�F��C��?��i>���'u�M&��z�Ξ-yD�i`��޷<�ڼ+���P�Iɟ�I�b>��'�~6-�zZPM`U(��Eߖ�a�9	2��E�<i��i��O���'Y�N����K�]Q�P��+'F/B�'T�jt�ii��9��H�O��++�p@ͅ� e*�&�� �������O<�d�O��d�O����|�2&�
;e0xK����8$�2�K�
3��dהokB�'jR���',�7=�T2%��T�Ԅ��_�A��2�e�O���-��IF�Iq6�l��q��� x-1�J�,l�� ��m�h�W�3�A��Wy�O]���%/�v����-�D��⎪#"��'���'7�I��M��g���?���?�!R-��lѡH<0uBB.��'���?����.A���L:yռ����1����'�9�R�Kc����$՟���'�
x�a�Ɗ,+�|���CC�(Y��'�r�'E��'��>I���h�!Z�
$@ !J'Ob.(�ɰ�MCa��?��&˛&�4��{�L�fA1 C�4M��1O��d�O" nZ�<�zToZ}~"Ќ&�`�(eՒ$��O-��ه���/E�SE�|�Q���̟�	ȟ������!�J����jP��+1�����$GSy��k�L�Yפ�O����Oj�����_�F�,�:Ʈ�f��q���B<eh��'��'�O1�jx���\=S$�a)�8Z��,����~�K����YVB�$bj�x�	ey2KR<���Td��7���R��B�s�B�'vr�'J�O$�I��M�L���?9�(]1R0�I
$�JRzr\����<��i��OP��'��'��Ά���{c�+�8�#��!{�X���iP�	/�[�1�O�q�����MΤ��K����P5b��d�O���O~���O��$>�Ӧ@s�UQAfA�B8p���p��`�	՟��	�M#�@�|����F�|��_�=D�Ь�xb��ïN��O�0lZ(�Mϧs�.��4�����6� J�a�iښv"0�DϜgN؈pf��?�'"���<�'�?y��?�򏙖7�����m�
G�|�n�(�?�����D즙�&C�ԟh������O�L��Q!U�bSJy���>*����O2��'��7�ɦuXM<�O� �c�oٌ\B8t[�]�!Yx�J��F��t��C2��4��a���nB�O8ѳ.P�!�.f�ǃfqP�$�O����Oh��	�<a�iۂ��D��%q��D��y÷N'^Ir�'�x63�	=��d�ܦ5g�Щ x2���A&U>� �_�M{5�i���ˁ�i ���!�2��F�OA�eЄ��H��>X���Aa4�ϓ����O��D�O����O��d�|2rOM�1Z�����
a�<���F�(��6g��]�R�'����t�'��6=��q�RKX5	�P�K�{��C�'������4@`���O2|����iC��+4O8�8U�ݜb��i�@��	�$ӌ	5��y�����O���|B�d~9�c2Z=� ���),�:�j���?9���?a+O��m�-����ڟ�I�E�d@���8ؤ ���F0@I�?qvY������ K<��0U��<U+F�k����i~�V�$�b�T\�͘O�f�	�MzҬ&b���3���VbY�V%Հ�"�'B�'z���4b�F�s�X=�G�ޤ�៼�ݴy�����?9f�i,�O�I�m����D��/F"��B�^
r����O��$�������˦m�'�%  nE�?y#�`>��r���!R���yw��\�'��i>Y��˟��������o��H����\e	���)Ȯܕ' �6�۹ �ʓ�?YJ~��;��ʃ��.Uz�&�+<g���Q������)K<�|2Q E-6u0�a�r�fU��ϧ��kPg�l~�ЋO$*����Y<�'!�� t��@j&f�:4�����H�������I����i>��'��6M��a��3a�a�$ڬ��G��&t�d�$��Q�?Y�]�;�4��ieb��B�\}A"�³:���c�D8�v���Cg�B���Gr�S���:����U֜{ +Z�@���S�Ns�<�����	럠�����Z&✕���ف��v���P�̞�?����?e�iD(г\��ش���Z�Iq�X�`��L�c%^����0�x2�j�)lz>�
P͈覱�'�E�s�$H'L�{�ق�x1#H�(=�i�	�G^�'9�i>��ɟ�͓DI%`��=Ev�@�<a ����֟��'�$7M>���d�O���|B�����8�#Վ*WF�V*}~r	�>�B�i\7-Gd�)����&6H:s�źS&��tI�4nn�m��+Q��tP���W����f�|�M�>�Z���E�)7V�iC�F�8��'�' ��tP�\�4��%3#�͒%4��K��6��q���2��香�?��[�xjߴn+�y�7
�_?�1xA�*u�飲i�D7 tT6�2?�'��P>���6�d.�"�,pcP�S�h$�C�ߛ�y�X�X�Iڟt����������O�� �n�:=�|�G��4Ir$$b�X$ٵ��O��d�O��������9w�`*�$S�=�V-�a�
)1��	ޟ�K<�|��ך�M#�'��y˷��	W��T�5��Y��'�
�Pd��lC��|2T��S����B�(Q؂/�:�h��e�ӟ���ן���jy�CiӞ���OR�Dh��z�d�-MN�P� tG�@�F&�	���d�O� ��I���Y�6�y�#��{�I)㈹aaΈw��b>�i1�'��4�I�NSJM�vmT{z���ǨlrT��	۟$�������w�O���N>���)lVX��$*�D���`Ӣ	���O��d�ۦ��?ͻ)j:Dɴ#D�Sv69r�n
��"M̓l9�v�nӌ�o�h30�l�[~2��9t0�m�S�(����ba��*��ey�oB	 j���w�|�_���͟�����@��韴3��	g��!-�?0.T��F]ty��l�nE����O���>����t�'��%c����UN����]�r��<!���M��|J~��K�v�Ԡ9�k�m�Xh Ā�9 t�����U~�9i����+��'k�ɶ5�<����W����L+'���������l�i>=�'�P6m�pO��D+im|�p�O�~����3��Ȧ��?��S����ܦp�4=�>�y����y��1z��E��t����Mk�OF�b���
����w|Y#jL�.����ś5�T��'���'B�'F�'o��:U�>_�2=�w��	3K�q����OT�D�O��m��=�����L�ܴ��[��}��#��LXi� ֆK��e���x��'7�O�8��Ƿii�I�F��A�$K�)n2�X�b O0#�o�O��&�I�	Qy�O1��'u��^���4ժBDԄ�0l/!�B�'��I��M�B
�?���?9.��(��ԛ<��zGS!�X��V��8�O����OH�O�S!z1r��b@UFǺ\�����`���&Wb��u`�L,?ͧ+������X��RT�S�3�Ș����9z���?���?q�Ş��D�צ��EjR5���Y�'kU|}#�&��4�$��'ؘ7�:��$��D�O9`O��Q����"Ş*g��f�O����8z673?�"h��wc���8�d*C,J�+@j�#=ʌA5k��y�R�����h����`�Iğ<�O&�Xf��|�;�U���Y�dx�l@��@�O:�$�O����צ�ݻ0y��(��]C��cE��X�J���蟤$�b>9����i�S�? ��8�h�$C��ե�@����q7O�Lr2��?Y�*�$�<ͧ�?���O�$<S+I
'��5���?���?)����_���H5EXyR�'۬܉PM�#Xؘ�9��� �2���F}Rce�p4�IM�I�s�2 �`���x:
6r��7:r�Ǐ��[�,��H~�o�O2���\(ڂ噱G���WA�y�`���?���?����h�~��V6JV�XQ"Ȃ�Ne� k׭
�x����Q�������I��M���w���0��!-�J1:�N'N�JY@�'s:6-�韠oZ.21f�m�I~�N�@e��NV�(uI�|�P�Zpϝ�GB�js�|"_��I�`�	��,�	˟��6D<df�ЁP��#G�&�H�Nzy�h�\H�$i�O��d�O꒟��&ąP�ڇ�(��T{�|��'4<6���%�b>���� 'ҬS��V�pP�YڲNE�CNɱ���hy"i�60��	+��'4�	 u*�z����ln�a��LA|NLI�	�L��ٟ��i>}�',
6�E2X�^�$)B�����%8¨�K��R�./�����	�?q�Z�����3ݴ/'��	e��&� Z�J�k �Hf�V��M+�O�1 ����:����w�N��E'�,aSJ�D�TvPM�'u��'X��'���'o��Y��2`����Ԩ~��"�O4���O��oZ O�@�����4��J�
�K���n��sd���3��D�|B�'˛�O�$�0жi��I$c1��Cm�L\�ȃ"a[�b�䩃��\�<����|��wy�O��'��/�!2�=H�������=���'X��%�MS�����D�O�˧\��	*��plf| ����x�6��'���8����w��q%��H��P0�eY#]�Dq����IL��$k�|C��r���x~�O�|���q��'�Ƽ��KI��&n4�X��'�"�'R���ON�ɴ�M��)	�'-�J&��`g�#���<G�Xtk*O�m�`��fg����M;R�D�\d���G܆{���J�O�3��+a�l9�Fp� �\	�z�G����O2�ū��w��@rP�A�JC��О'��	�����ܟ��I�����@��$ �u2���%@C�x���)4h��h�6M.E� ���O�$)�9O��nz�Ah�P�`2ȝb#���\���,�M�i��O1�x9�&|�2扒,;�P"���-�(3E�0!\0�	$e��P�'D�'�������'�06n�|�<uH"m�%όEi1�'���'��X��[�wx�@��㟼�Il�&�3�Ölf��d��N8���?�qX��	۴m<��b2��I7
(=ٗŔ*89 |Jq�<% ��(U�r$�f� y^~b>M���'J~<�	�@4�k��O�VT(F`X�5n8�I��X�	ʟ\�I\�OI"�=a�Y��N����b啢)�48�I
�Mk�����ަ��?�;:k@�A�V:>���E%LR��Û�!r�2`m��|c�1l�P~��?J�� ��>� �SA	?5��\�B_�kv�|�X��Sş8�������Xɷ��$7D4��E���T���UZyrlh�j�	���O����O����@b��
K�>&�A�vE�+�Z��'��6�F���N<�|� A��>���覣N�w+,�Ps(Q�APH�"�kB~��P�&�����5��'��	�|�F�cW��?
@:b�B�^�:a����	��T�i>��'�.6� �D���d��3t�S &X�\�&ē���e`���5�?��^����ঝ��41LHi{�,׾p�V�2⍥<�z�A���M#�O��$�O�j��$FF6S|�%0�JM1ܔ�y2ēuNj%��[��DS ό�1wT��&'Q�bTԅpQIJ?��H��Ɩaf:����P!��{Əda�I���8Q�:��]�{˔��'E�(gL����"O��̓Ģ͏(�FX�!#؇f�0�!e�S"F0�(�>ڭȇ��L@��E�ȁ4�6�#� ߍr�`a�V4jhR�y! D�@��ղ�,�+_5�m���x���h[&}�ZlR��	q�d�:�A�\��5r7/�!K�Ͱ��55D@���&� H�x�a�7��A��������I�Γ"`���	Ο��O���Op�W
�, *�dZ$��sn�t%�H�$�
�ꃚ���'B�'�J�j��ٴ@s85 ���5Ď![#�h��I�}�R���O��O��|����}쾙cq�	�N�Hl2&������J�2d��Y���t��ǟ����h���-0jt	��T�d�֍X�D�[hK�;c5�ʓ�?1���?�J>9��?Anv�������Y�	1C�A,��ɘ0��d~�'��'x"�'���'�Hk7�X�~��p�L�9-�����wӎ���OP�:���OR����mت i!�i2���qge�,�kU�X�&(f\��O����O��Ģ<���ߥ���ğă�'��E��%��J���#޼�M�����?��-����{�菧v-�� &��FB�����MS��?9+O���ǎ{�4�'t"�O�ڱ��,�k?�Y�KP
8��u�-��Or���[ݚ㟐�'6鄴�kQ�
 S�e��*�Lm�Py��Z�-�:7-�O��D�O@���g}Zc9��A�M*C�T!d�ڴ�?A��q[��A�����'�q�rQ�n	�,Y�D�#8�r�(w�i�Ah��v����O���&��'q�I�v[pX9�U=b�P��1�,zNM��4#@Z�FxR�i�O������Z�ɗ��r��ţG��M�I����	�p�
0��O ʓ�?y�'�Z�8'�T�So2aQ���~��|ݴkz`�'��aas�'(�ڟd�I֘͟�nRP�$�ڳB`*��إa>7��O��B�L}"Q�,�Ij�i���� -�.h�3ND*&�8ЁϿ>A1J����?Q��?�-O�T� (�S�/_9S+`q� B�\�P�'��81���JyR�'A�'�B�'��h`L�H���`��
S�`��FP����/�yB�'n��'H�	1���OV���q��)'�0j��ś�6A��4���O��O*���O�5�Gj���ȕ)�!�����ıT�T����>I���?����$З3~��O�)Ɍ{U�qs�,��H��׈ޟ�M������?���44x���@��,�'Dq)�BH,h,�%�Ф��L%"۴�?q���$$�h��O�R�'9�ħL
 ��iQ$C�H4l|k��dy|Oj���O&@)tG$��^�s ٲx^Rm����?t-n� dȒ��%�'���bf����OP����p�ԧ5&F�p�x���=`��0IV�@�M���?�����'�q��%��h�;PP��ؖa� Q��i�2�qljӆ�d�O���@�'��I�D�h����5p��(�m��-�J�4G&H���i�N��'+���$v0���K�?��E��Ł�Z�>	lɟ`����X��NՕ����<���~R��l`��΃K�������'�P ��|��'���'.h@�h[dx�%�ҍ+$�(��}� �L6)W*��'��I��ؔ'����m��i�P8w�U���[���}���%�d�	ğ���Uy��(.!��;�	;'��8 e
@8q���l(��Ob�D9���<��gʁ�R�R|ր�;6��X��n����'��'��[����N�����L{p�C��98	jl�4	������ON�3���<�'�?`�C�LhRp�0׉~\ ����F�J��IƟ,�IӟP�'(�3Q�+�	d�f� t��ӌ��h	B(Nyn�ܟ�'�������'`�{�4(i�f�a�1�%��i�0�m�����`y��K�k����$��k����P�MªOAڙ[���e��'��	�|�Ih�s�֝- �j8I��Οc�q�v��D��?�/�6�?����?����-O�NƴZ��6>cJP�d��>	���'5�	��f#<%>�؄�D	_s\��䯊�9r����`ӰYA���O���O��럎�S����h��W	�?w���*�iV�J���5 DDx����%�h��ֈ2�~� a�.+���oZ���˟�A�APyʟt�'�����#N� �RQ���	j"i��@$r˱���d���-6u5������9f343�$tӼ��֏�p�(��}��m�<�`�K.bX
$�qے7肍���x�	ژ'��_���	�I��M�g�̩*�,H����]����#ΚDy��'"�d�O��ɰ4�J�������<a�GU?6��6튶c ��ޟ��Iڟ�'H:�j��n>�I�b��?��	����J�bA2��>���?�L>�)O��O �Y�J�9�|�,��HQ�R}r�'���'\����HL|�F��/-I>�c�C�1Ll䝢`CK�c9���'n�Y���F�D�'?�'T���@ѹ#r��ŏ?��l����'.�H����ȟ����?�l"�X��B\Y����uc��}[JO���Oz��1��4�1O��9>[r`���#4<�G�]�/ 6M�<�ѢZ�F�f�~Z��*Ӟ�8��Dx���@�I2�b�qӖʓJgJ`���%��O��M+��޶1�I�E�R[����a�ަ�@�"P�t������	�?���޶,�H%Q2�u��s�"M
)oq���T�?�)�'EI*`���ĬF���3�H
q5H��W�i�r�'�"�H:��)I�\E�G!�2IX' Ѱ9������:��'�>�-3�	�O����O����c��D6Bx'�q��T��&����I�T���K<ͧ�?�O>��J�����MQ�ac�ܩ��R��ɖ	���	^��şԖ'��-��3��@`b'�;a���#Q;%~^�3�_���Iʟ��?A��?����g��Ae���q:~�zW(܂!*����`~R�'g��'��ɇ��J�O�q{e�K�vNr��e.ǼI�LLٴ����O���?���?��T�<����?��Yci�	L�����H��z���'�����'�B_�13�����OklA=�P`���Ѻ���w'�r~�v�'��I�����џP9�y����y?��P��T<H",¡R�Ȁ�pM�ئ��	ğ@�'��tc�F�~����?��'HYZhh6D�`�҅lW�k�s�T������2L�:��Iy򍒬����?U<�c��>T�����K�l��W�����/�M��?-�M���#_�i��v	��h��H�u��YT�$s%{�,��On�;O����<!����a�܈��j��>�m	���M��LЛt��6�'S"�'a���>�*O ��ɕv�^�
t�W	�(����:тt��&�,���6W�s�]<l��nM��l��iAR�';��d���D�O��	�\���#�/_�}z�)�dXJ득��� ��i>���۟��ɾ��b�B�^����7��7O���ߴ�?)%�Y�%��	OyB�'X�Iϟ��N�\��PǑ���;�ƌ9+���X�̓�?A���?���?a+O�tk��Ẍ́e QfC�ڸ�3e�<V�VU�'�����'��'�"n�&��g.
����ɋN�-��'q��'�dA3�'YW�|�uo�;���8�ČK�H߿ꤴ��鈭�MS/O<�ħ<Y��?���(����t��G�Z*Yfl���~:�`�i���'��' � ��⯟��U�? �H�q�I
%L�\�WO$0���(e�iU�U���	�P�ɴ\����Y��*��a ��A7T5��JB�I8���'�"X��qJ�4��I�O��D��T4*��[�es��h�h�4"�r�е��M}��'���'�����'���eE���FG����6��+�!��@��n�`y�)�8U26��O���O^���F}ZwN�-K�OߞM]:M�uU��3�4�?���N�lΓ�?A.O �>��b��!w�}�'���@�\p3ƆjӾl�L���������?aR�O��G�VeB�,1fd
 *��S�@��@�i���b�O ˓��O���[�r���T>.��ܪ�/C�e#t6-�O��d�O�X�l[N}�^���	r?a .PHxjt��.Ҍ7+��*�i�Ǧ&��A�.~���?������S�8@���8̰h	Ë��Mc�^HX]�0S���'��P���i��m�N��؊��	!���� &�>�E	E�<���?���?q���$�>"P�A/��� H�f��8�Z�I1b�E���0��z����4��VtL����A�l��⁋��AR�q��'+�'�RT����mѣ����*��`�`�ԽȜYsw�0����O,��8���O.���/���GURm@�I�%-�};�+�5g���'�B�'��_�HJ��B�ħVFL2F��ifH �����6|Ȳ1�i�"�|r�'����<�y��>��'�}]����Ҧ)! LF��Y����t�'��i9���O��)�%��=:�	�#0 Y����2=��'��I��)��q��$���'J�>��3�
O�4�@`j�-G	��n�gyrE�S{j7��n�D�'�4�6?9&k��0�Xs��	}��"����I˟ps�����&�$�}�dD9'��5D�?d�4���RȦ�ѣ��M���?����֘xB�''��a�͋#Z1�����/�|�$�`Ӣm��O��O>��"/ ��Ӄ�*����cq��ܴ�?	���?A��D�h��'��'��$��y�@��f��� �öE�2,��|� ���yʟ:�D�O��D^�gK��a����S��\ CS"e��d�96qz|�>����K�W1,(ՈX�,[����l�_}���/�y�U��������VyR��A�H���)>s ժ�Sy�t�4��O0��&�$�O2��M7!z�����4�6y�g�ԗ}C
A �'��O&���O��/l	i31��%�`B�*&�V8��ӄ;;��՟x"�'f�'M2�'��=@��'LL(�Ƿ6������I�\���K�>9���?����$�_�5%>�a���l���Hpg�!��x2��˕�M{����?q��?�~�s����	���9(����cL��'�D� �J7��O����<q!�'߉OCb�O�������1��U+F-�$'�2�4H4��O���̼K��>�D�?=�b-S�(ntJ�$ܺM>� �jpӮ�Z�Li*װi��'�?a�����D4�H�A��?����f�ߔ��6��O*��J1_��d0�$6�S0�v��Ɵ�(��@ge�6�ZtP�oZ� �	ٟ����'�v,��*/=�(�`�ϣ�8��i�P�۵5OҒO\�?��I�hs�!���ۊ3F�l pL 8"Vq�4�?Q��?���*@�O����� pDL���4����۩O���� fӎ�O�-��HAL��ڟ��֟��[
<�4�x���'�~�X'h���Mk�e�bp9��x��'�b�|Zc��CE��zC ��%�[<2� �O��*�>O�ʓ�?����'2�ƴD�Ռ'�,I�,Hen�iЦ�r�}��'i�'��'E��F(_�!����S��>+fÆ
{�b\���	ܟ���qy�
A1��擌SP���ҷ�����C�%�2��?	����?�x�j5�+(P� DO$��lI;oX5	_�0�I˟(�	`y"��?��( I�/67��qm	�?Z��E����D{�':�D�'�����R��w"݋vH��U�qӬ�D�OLʓu���[�����'�\c `�gO�l�8\{F�5X^�Lڈ}r�'������'Q>04�X�F���{RjؠU
BI��bgӤ�����'�inv�'�?��'
����&5�\X�@�	cJ�8$�E�=�>��?����?�N>�~�F*�	=��y�@e)]��XǦ�ň���������?ɗ'�S�r��8G#�99'ѣ��J���ߴ����[_�S�OEr�\&ac�0$N.c�����#$��7��O��D�O8�R�d�w}2^>q�	؟��ë�3mo HPVn�+3~� I l���'�aQ�yr�'�R�'δ�7E�f8�%k"Ӵe�t�wӢ�)�@˓��ٟ�&�Hіi,7���Q�/� UV��1� ���ޯ;��UI���$������IXy&L�A�9�sM��U��4���nRtI��>A,Of���<I���?��,�*e�0*�W�¹���>Y�.�@�,��⟜��П��'b���.q>A���;E� U��h?��i�e�nӊʓ�?�-O����O����k���(m����`����� �%5��oZ՟��iyo�����';�mط��~��*:J�HA������t�e��iHbQ���	Ɵ$��l_6�K�䙁x��$�Q�=�~ à5!����'��W� R"�@��)�O2�����#@� q�j�J�/��}�����G�m}B�'�b�'̈́�i˟�IJ2'��#�&	sP&�ܰa���妝�'�.��ak�,���O$���aէu� Bl(���_�<%�b&q%�M���i���'ڔ��'�b^���}�U���%��i�`TP���[��ۦQ��V��M���?a��ʦ]�З'���ѫ�x���۲��� �ȝc�`kӨ`i�8Op��<��T�'�
�£�A"Rr��F�
=!����Hl�$�$�O���,|�u'�>�*O����� A�f��V�:�3��'�"i�n����<�KM�<�O�R�'��	X�$Q��:B�->r6X�O�ag���'�^t�E(�>Y.O,��<Q��sv)O=s�����"a,^��bGY}�JU�y��':�'���'+�I*}b9� ���~�S&՟~ hL�1������<������O��d�O����)��u��4SK��y�L��!
.���O �$B�AdR6���$��=��O�O��,���A�L���J�(nT�EK�'�<�s�m�;��M��Z7`1l)��{���0��ՠg��k����M@���Y3�jZ
t�AP�JȂp����7m�@ff	�C��|����vǾ������kr��'LŘD�`ʴj�|���p�w�|�1�F4��� O���0��fȖ�6YD#`(J�l9K���!\���� �ʬ&�T���i, ��5wb�?閯U+X�@dr��N��8&�I�?��?�*T�㘧�Т� �  �N��ӡ*F��!F<}2L{���O���"$C �x�"�(�<R�ҝ�O��E*�O��9�)1���9O�����#j�`d�I�6X�1Oh��3<O,��D�V��,�W)P?$�^L	�'KT#=I�OZ�s j�c"nʶR:")��֖uy�Iן��I�F*� ������I��iޑb��|��L�KY6(������P#]���N��[\�c>�O"��o:֫��)Z.�cH��d��`��>Q���t�L�>�O�(0��Z���Ӷ�O7Vz�Aiq�O��m���i>AG{Re�7�p�ӗ���E��$��A[	�yR��}�7N۰E'�D�V#S� � �'t�#=�OX��3f�(��$�X�:�*��W�9[1�AaA��C߈��	���	П��Xw���'��k���QD��;/P�hE:F�Ĵ�v)�*�����H�F_���$ȁ2ξLY�	݄qHh9���.�� q
F�U�͐AɎ"N��䆏U඄� s��[aiݛ!;0��W�'
r�IP��r�2Q�b��c����c�Dr�:�ȓ=�xUIg��%g¥�	��16�e�<�2V���'1�XB�El���d�O���R�X�=9��W�T�	e2)(K�O�����V���Od擆	V�1Jq��o�I�oS�i8Ag�5����@�̞d� ��z��k�-�$Řp^=S��
�}�&$�"�.#��x�lճ�?���?A��0�d��ׄL#���A2�P�L�*+OP��*�)§Dk��Y�iUa�fs ��H-����;�����?���S��0�q����y��)�'D��(k���<:N�R�cɏ:��ȓw6D�1F��?�z&B��sjͅ�8�� �����V����!��:<�4�g��[�b$��L��o�!�ĕ@`$�
��	+y�j��e.��!��X�l h�]	����2��6�!���2*����ţd��(7'�!�A�}n�a4~-j���/:$�!�evИ*����]����.x�!��"F\�s��~�<ui�P&�!��e+�dy3�4-��0�CC�!�$Fb��`#gW S�I�1#�2y�!��fb�H#�D�&3��k�ۚZv!�dG&M
�A��
V���ic�惙4v!�
��B�p�Փ}���B����z�!�D�J	�D�A` w�v�To@��!�d�$\L��'�6+�<ˁo�9U!��1sH)@� O)���
���xQ!�$�+����C=�|i���!�!򄏋"���OV�4���&�X�!��!DD�1Iέi�b��D���p�!�D�4n�8�"�K���0����a�!�D�� /������c��liV�I�!����y`�R*�vla��	w�!�d/}�4U3E��Y��LA� @�!�#a84��@��xpp`C̗f�!��5)�2%K��M8j���boY�#�!��J����ZEL\��l�sҧe�!�� ��� �Z44=� 偞,�,8
�"OX��BIv�m�4�ɷZn��R�"O,��b��b��#��Jl�y�"O|����R�hiI;q�O9���sc"O�}�,ˀ$E����K~�Y�"Oh(�4��7#yz1��>`x�-9a"O�1���>�EZ���6f
��"OD���kW�GI�h��C���$	�"O�9/�;���6āDm�L�"O(��j��\�$�Z ��[Jl1 "O�qc��r����!ڷV��� "O6��V�D�.k�#�Q}�zhg"Ot���LP�RKN}a���	�x��"Oyq�0�����G�	ʞԈ"O�I��f��,y�	�	X+Z�D��B"O:��Fo��.�
�X�ɂ-��9Jw"ORi��oP�`�H�s�Ŋ+�T8"OZd{�������W*�>���!d"O�A
�#�j|��V�y	3"O0�� ��Zq�U����I=�T;D"O.4�`�ew6���- ?>�"O\ܱf�5Y1V��j�:H)��*E"Oj �S%)WԐ`��P�!����O&��TO�O���䃄rzP��O�.�Ƞ�	�'
�\��hY=7��#�k�({>ൢ$�ʧn��O8�}������t��4U�Աt�]7a���ȓKF]Y�dK!"�P�5e��!�
�ɗqD��Q
�t���ȕ�Y��s�1)�J݇�4_�0�*O�I��D0s�(���Q!����"Or|(�� kP1�݈qN`�@V��.���D����&M�:���8��(z��ɀ�y�Ҋyn6`ˑ���A���`��%l�:��g�:�g?�v#�j�P��M�z��u�q�Rj�<A�� �})V�#p�
�U�P��t$��<�b?/a}���,z�N�H��EpNXXe�U�y2���H\dff�?D�@2���yB�R�Ob29[��YwǠ)�Y�U�ȓE����̑>:����b�ҵ��%��r�x�a�6�Vę�
�1y�=�ȓ_�F�c��jR����ჺ:��h��YJ$�v�]�+���e�A5b����J�7*�3b�Y��"�P@�ȓm5%Q�'��AG�'.����ȓ?X�X�DA�5��ei��D�76�ȓ(��A��L�HG��dl;�����f ���/�Q�d�w%E�zf���P�BT��"�g1̸p��J�7�J��Or�1a�*lO����gÍ#���s��	�8��d�'�.9�V�i�P�!�t���G����q
�'x��W�% :��C7�X������$��x=�"}�#I�L��L(+�pA��お�k�<'Eո�nl�wM�	N��%g?��c½���h���X�hR4{�f�bQ�.f��e�B"O Q:��Q;���g��\�܌jp�>I��:�=���ƌod�a�� ߅H]ңFVK�<9�A��6�vUC�Jv��9�� \�<���@� ��0IFOR?h��PgmQW�<Qt ��>�\���[=��9�͌T�<)���?e`�C�n��(k�T���R�<��(M�?yl���)B���R�ER�<Q�+5���''�g�=X���P�<7�H$u�Xx��k��=�T�#���g�<٠k�p�"��dO�H���0S+�x�<���9EB����ȺfR47��u�<� �XYU�̞(�<�J%����(Bd"O���o�f�Y�j �s�"O���+�D$<t��N;ZT�m�"O��ac�1q�䔳A(�sAʉ��"O�@z�d�yX4�`�11࠻"ObЪ���%��4��8*��4"O���	?uf�Hp������'<
5��V��QE	"]
n�+�φ�R��q�'D�����7E�.�#�m�/Bg陵�#�}3�tRA/�']?�|	f�D*L�R���E�#4���ȓ]�j�`U�Q�+�Lb�x�D`ٱ�F.%�"~ΓU�h�`-ٕA)�ē�/��v_�i�ȓf�@(� �˦/�`H�r��1k���N �m�66�O�I���H�(@4 )��@
I$`��'J���I&Z����7@6�����%̊A��F"(�!�D�8s�8QꉳM���de݉) �O X[sj Y��ͻ��	E�z s��f2��T�ȧ@�!�$�I�R���6x��pC�V.F2��P'�>�M��B=��h�͸|Z���Ś<�~���o� ���:�a}2�H�1�z���njPB��f9��s����#BG�(����\�����۫n��a�UH�A�D�B��xRf�D��H���j$�!c&��'a^�j
pҠ�d� �%h"�����yh��A�JEYH���YhƌG�MӰ@O�l����KM���&	�0�|�����Á�ïH�k��Gm�@����Q�R�Z�L���!��,�6��U%%l��EI�Ʌ��r���`j�d%Zj��(�SRǑI1ZKA8d�ڄ����4@�K��=�&mk�j�%"ȭ��B�sbX �f6(�X ��:N{�{�%�&�H�Į��O��,8�,Ɋ�HOV���O��0�m �DÇ"��A�� ��'2/�����
�� Jң��Y�X��
v~m��.Y"*	�U��h�mڏi��i�IU;�aPƫq���ئ�s�)�g�+,��#�Y�t~p�� D�`@��O+x�
Po�c�d	/bD��:�h�H�g�!'st(�$�|���d�K<A�lp��a�6a~�G��	�Xb� F/2�(5�Q�
�$���O�	nl6�U�X%f0(�bľ��5fӵ�ʱ� ��5r����'8�^��'�O�1�2���OQR�ʒZ�}
	�2"O��
R�S8fh�D��2�qX6��NK�YS���54J!�8<� y@Hӿ����$��b�O������J
�"���=�uoN�_�x��{��9OX���T�+�(�
Ңυ*٦�1Đ�P��U��ا����3kYo�h)'N�d�8,1�5O�dr�.���p>����&Aj.p�����!Y�U�N���l���kz*�n�\3
�kO|�ȟ�DĬ�Th��+=� �{��~��NQ3v�x�l��U��u�ݣWy��(7B��N�y�U-����<x��Z�(�3�I�Qb�i�
üM�gӮq��܈OÂN�Q�Щ4�˔9�0��Gޭ(p4-�e�O�h�qkԋi��Ѻ����>2b��'SV���+\EyBN�#^MGy�J��	Ò�E���bJ֘�&b��~���Z]�Q���Q�yH!Fߤ�ēm*���O@~����/��UV�Q�v L�Й'J�����OE8��&�6~8�j�-=09�\�A�T�(�Ni�k�@�I�,��I�?�;B�е:5�v5 �t�ذI�iF�'��P"�M�Z)8����xBz�j�$ήVHΓ�`��%��y̓1;���#�ǉV���h���8���b��O�>�8&-��E�� ��A@�'��	� リ#R�[���! k��Z�N�����w2��P�;�b��'�l��' ��r�٢��;���S��I��m�j�S7/�_D���b���}�'a� �o�5k�y�D�˖7�ʨ��O*-�&�Ƈ/�e&�(U~�(��%��.�J��5�H:1���Q��	��X�ߓZ;���@��1MjN�:pƎ9�"���kڿJ$�Ѡ^�����ξI���id@��3����`qH�e[�)2��5@��@ �4�O@bu@�����[�焔�>�
��vU��s��5>�Hx雾Pa��?��wJ�#(t�	E��j�t�:�o�,2�n�Ѥl�$Y��x�N��P�џ��%O��Ud�H4��-FB�X'�ܙ&c�ɱBK��6�y!eEVL$�����hj�'2�d�c�Hڹf�jȲDG����'
��%`�>����g�n��M���G�(��k���������	�G��<y,�2��Abc40� -N�r* ��$��3�E#2NOR���D�2H�$<�'�F�I�l��BT�HR�'ɖM�JM�,��-��Fړ��%��'*zd�&�O��Y��[
U��jQ���x�'b�� ec���KR���?W&��R$@�(m�"�� i>���w]���D��4�O�b�������;��S�dC(i�N��!A���p<��L\�	��c���s-K*F5U���O�o��i�	=?��E�j_j(�2l�^��dK��A�'����K�iFh�.� ��M<IP
&!T1O�%
�
��XR���#i]�%{^��殇�{0:C�I+n��"AǱ�8]���6���pAh�g�S�-�~��L��l���"��C�Ɇ`8l�@r�H��Ȅ����!�(B�I;,�@�:��DvYB��ڗv}BC�I�@�����Q�f�z�����C�5�L���+��7O��������B�I$"V2m�v���Ʉ�Z�&C�I3	��ٰ�HU�s�|4�����VB�	GT�)b�'�!�" [�C��0��B�ɸ	v䁑�&T�i^N�[��O�`�C�ɤa����BH�|���c�M�U�B�I�;�z�JƇ
�=y�Z'�<W��B�	�<�D�u+X%p��ٔ�[4tC�I�}��{2��/6A����v >C�I�3��y���?J�J��޺o�C�I�|�d��g��i�
l�� ��,B�I�t��<T!7���y".[��6B䉯, ������+*)���JC�	�c@�8�%ܯW��l��.H�3�B䉛Kl����'�h�����&O^B��6}�M�R
jVr����0XLB�ɂpl!�$JǊ{����"dC�	�?1.-���֣Sg��Se�M�5�C�I06p�Ch�7[X<�rE^�7�VC�	B���䏼�� [5�q��B䉂��l*�"�z���X�_�B�	.Wbh�@�B��<Y!BxTB剟,d89zGQ3p4:D���E'2(!��L-�R�
q��{2� �C�-!�䘹ݸH�W��ܲ��&!�[N�xJ�)	~�v���ף�!�Ҫ�h�mͨ|�$Y�Γ�$�!�$[�NL���V�D׼|Q5��!�D�|TC`.��3HU�W�1'!�D[�V!��f1���W�!򤉴5}�!+"��9ON��äˡ�!��5^r8�q�'�7&r  B�/��چ�.����8Y2�C��z�	�g�$60�H8T��E�xC�I�eⰚ��AtΎ���Q#U�B�	�_��!&M��0J�i�ώ+�TC�ɨE
�q�3i��V8���>(j>C�	�h��)�B��N�(C�߯XCC�I9G;:(q�H@�>\�p�ܲ:9�B��CU$-�'��/m.1���N�tB�Ʌl�J�Fٿ5�,�Ѵ �3PTC�	)$w��"�!��# i^7��B��$uԄb�A��(�xb��U xC�I�{�L	 0&Rs�UX�l���VC�<'F$��ҳ!��%�Al�pHC��Xj��sଖ:9Q����٠��C��*jn�jq$�2~ikb�VvݢC�rq���m�W�X�a��c�C�	�UCd1S���b�NU��Λ9l�C� =\D��d�\u��6,T�D�C�����#��1Y�꓆^|C�ɒBC<p��2g�a[�լ`xC�I��Z�Kr'ʥEd)��bS�=�NC�ɐK�\p��@ \p��y
�B��B�)� �43�+םz(�3�̓�,?�E�e"O��W$	�v���`�D�v❻�"O0�e�Ŭd-�y��B��b���"O��Bw�U(Y�ؕh��R���:7"OQ��[�,�HW�
t��Z�"O�S#�\�x$�@�O��R��"OD:%��:���{$`U6O4@�4"O���w�B?C�����B��T"Ox��Ŵnv�-��O�}p�Q"O2��F<,Ld�9��(E�b){�"O�� �n�I
�́/l$�(�"O�������|
�$��jP#vf�a+7f`H<Q�Q�QD`�ۭA�<I�M�<a��+���$Q�fvX1)XO�<!�HѢO*��*R�	&!R �Jd�<aCl��a���sA�u��D����]�<i�#W�b)K4�V�~����E�\�<)���`��RQ$�CŸ�c���r�<I!���l�� �uy�{C�Yl�<!��$ǆ�z�b|*P˧G�r�<Y5i��S�b,������DW%�z�<�'�#����!YT )�@�M�<9t�R�R�B�c�����jPr���F�<A�ӊ\�J=��T=q-��� �w�<�`�{�BHX�ҹ~�pa+�/u�<�FlA֞�O[ �B����j�<Q�ʚ5�h	� ��=i0݁0�e�<�$A�c�p�	A޶HF��ӵe�h�<i��Q�f4�AX,2"�s��Nf�<�d���>)� �4u8�IdIBc�<a�e��M�.�2��?|:`R���`�<)�cRgk�ʣ-��3_H��� �g�<�T� G�4�0 �֎��*Ig�<�ъө+��K��If�t���Q]�<��-S>̴��n\>r|]� �]o�<�a���}�d��
�JPQrv@ G�<�mV�f($��c(�7)~ls��C�<��06�h��,�)#2ţ�#]i�<����G���c��	��1ӧN�M�<1#O��m��h�W�R���d�B�<a�E��^��!�Gƹ@�(Q�%!D��*�5�b�q���8��[WE=D�� ��:.�$��G?[��)&D�����'+��)׈��D����&D��
uj�o��.y*��#'7D��/K�R"8`ȡo�^@��.)D�t�E�ŝfTA�����].�e�wM'D�0����f��5�v#0]���j#D��spJ���lP�[z4���'D���s�ό*���GOO8�
�`d#D� 0��_�.�$�ӐL%.2��?D����6W�Z�C���phY�%=D��*����`�\-�����#����CB9D�ԙAn��$,�th���D 2��æ6D�B�B���(T���*e�9D��z��U�O�|چ�A� �
E��9D� ���	�XqP���#U�,�ڔb�7D��8���'U&|G��� ���C2�:D�X��Q�,\"c���0s�b7D�����U��ZÃF�Q���E4D�����ϖ.��A��:Ą��3D�ܑ劒~�l�LC7M�h�a�%D��C��մZ֬x�`͞�%�xt��B$D���D�G�@���'_��@�G!D�� xA��R�TVj5���"`��I�"O�Us�nm�8�dF�.t!�H�"O6��'KƥL6`�@�"�v�H�"O��;7eǍiP"E���U:�>A�g"O,�Q��TQ�E6M��A1@"O�B���4uӊ%r"��e� %*3"O^���?@��P"ӳw�z�R"O���S����r�(��`�Q�M!򄉻{j2�r�I)3�v�D�A
<ў���ɧS�@��2�T,K�)8����I�C�	+�x����H�<xBj� [�~C�Ɏ��CRbY);������ 4\C�Ʉ+��x6,���d���z�"C�5�|�.M=� @B�Ⱦb��;�"ORm�@��
GP����d'a&20�"O�9zu �1�qAF�57�	z�"O�)b�P¶�i�%K�A�ƅ�"O� (`�D�B����%C�9�:���"O�����W�D�c�ɱ;�pH�"O�H�����H)0��<*C"O�9��)�G��D�g
M��"O��a���6|��q�͗ 0@�au"O�1R��?��H#��(�Q�"O�4x�ɜw�2U	�)�&T�F])�"O���1�E�[�@ȳ�.����f"O��A3��):F�p��Wx.��3q"O��H�_bcX%"6Nи  �A"O�34�Y$�����:=�x�r"Od�r�-��<\�a��� �ڔȃ"O��7�~7xt�a��<����#"O<Ђ�ңw�d��R�Ź#i��� "Ol�H�h9\�`�¬iX���"O&�AB;l��y ֦TZ��`"O6i��H�OSܨ�G%�|5.�Cu"O�`��"[p�9VC��"�5�'"O����+�W�`�bF�+@���""O4���ɧ ^��wAA�4��"O0�"V��wZ���R@M�*֨�XS"O�9��2ZY0]j��-tD��"O�0F-�?��)2Ə��P|�7"O�$9B�N�j"�=���E�����"O ��u偦9�RÍ[��b�)�"OU�`*T�!/�h��S� ���ʁ"O��;���;D+�,���2\;�h��"Ov4��	�z�$Hb7
T�FN`�9"O�XK1j/J-Z6iۅf٨� #"O
���X��� ���T��3&"OѺB@�{lw�R������8���k�Y3�$�-y�q�u��,)z�C��'I�|��R�%"v�z��D4TU�C䉰1�~�T�]$�p���-W-,���.���)��!��H��2׊�
Q���Z_�C�(Pb�A U�FTLt��(х2�fC�ɍ����4.0���\�A*C�\�1�-�2,�VpD��-i�B䉣D��m��K855^��1� 9 �B�	�L٨��"�[a�!���bY�B�I8�l9���43k�BD�w%�B�I�C4 ���̍/�i�j͸2��C�I7��T��e*��z���]�C�	$d��Q�n���%I.TzC�ɪ<�: ��[�>�SbbE>^ZC�	�\l:�Jdf�P�FtP��A���C䉧%�LUY�b�^sz�hR)��C�)� 
�!��K�V@��`[��[g"O4�3�i�.��!��̎2�<��"O�1�2����]�s�ە[�N���"O6H��++丩�c�To0��K�"O�	�$L�(IU�1�H�;(Ű$"O9��)�(�h�ьB8	��F"O(((po�'��H����n�,rp"O<t�h_�#����k��8�`��"OTH��+N�ukr$����@ؤ�`�"O����J�9yS�y�c�W�\��"Oxp��ɗ#6�a
��w㲉���#D��"���(3���5�D!�F���"D�XJ&`�*385*$� /x��bej?D�@ZTI����:f)���(��A<D���$;����_�8�;a�9D������r{����!'dwJ���k8D������'䬘v)Q�@o& ��7D��������8�Ȑ�T�H)�Vh3D��:�W�Ar9�h�"l�ca"3D�  �`��sd�8$���{Nyt$2D�$j!o�BUܹ#1�͚T2)�1D�(�4�@�ᄐ>!��`�Tm*D���C��^{. &Y�̍0U�&D�0Ѣ�4��:'뇟��a�Vc"D�h�H�@�T(��D�.ds2�;D��-�$O��� S�Ц+�<�[�;D��iQeU�x:�
�o��V&"����9D���A�c.� c�$�Uk�6D�4x$n_12�<
cD�́*�:D��)��	(D�¹�P�Jez���a�+D�`Unev��Q��J<HШ��(D��@�D1^�tE@����T))D���.V+}����CeE���t')D�\���ڞ'4��q/Ņw���cu-;D��S@�T<��(�@�"7�J��;D��� ��88I�������P�5D��2�,�TTL	����bd.Aj�4D���nU:�`� �JM�r���!-=D�0z�N�&Qjx!{UG9'�Ƞ37�9D���� 0�Vmȳ	x�����5D�tR�o��U�lk��/^�E�q�4D�ة�L'�N�QgpWsY�@q�'�Z��A�C	#	��s��>n*@i�'��P/X![��!�" ��O/>,�'i�i������R�Ep���!�'ќ�����
A��qI�Jȼ� i
�'�2G�M%)3�pA��	�}�,9@
�'$�y�T�v��a �k�9%����	�'D�D��-L=�6dZ�$@�K	�'��M�����`��;��G��$���'����&B�.��s��#����'�¬�R���_�^�ċ�/9w�40�'�t�B$��):2��xec�"0���	�''���'�NGt�p�*���}b	�'�P��Q�l?T	2��;�,��'Ԟ!@תUD��9$+�)er�)�'���v�[��p`A&����Ѡ
�'p*�چ���Ix�������Uj�'XXpwAZM�p�ҰH�4{�'p�sC�@]�>L��D�������'��yYv���o.����( ��
�'�~Y#!(�y��-Y2�	3m���	�'z� c/�@3>qc��)]��k	�'�Vu��@*1��C��7��	��� ��ϝ6}�h��Z�'X��"O\���&�,ڢ]�C�����@F"O4X� �.
@��6�?�~��B"O�y���X�`+�-zw�A�"O��enYg{n�3p܉I`P�"E"On�1b��.���(��H�f�7"OHI�`k�3�8T�"�I8f-�j "OzJk˞d]0WC** �"Or�2�G?`���B��-S��}s�"O�-�ׄ�+0�����`Ҝc�,YA4"O�	y�Đ���m`��$!���r"OZ\�d�8k d�v�յ?r�M� "O���F�
;xR��I�SJ:\��"O����a\�J���`[�Z��}"O�H��	6�0R��������"O�@����@PUʔ�G/	�H��"O����o�(B"Kgf��K�Lj�"OR�@/D/D��FB�Fr���R"O�Hb�+�<X	,�i�d�}@�kB"O�|
�O�|&��Р㏼J��y"O���b�%+����+I�u��15"O��b�y�J�R�(�\�
T��"O�,��ʉ�H�XL�A'�E��P�"O�@c]�;WH��GoA:*�j|�c"O�<�0MxB�`�� 5��9�F"O��hB���f>	����?Ң��t�<)q�R�n�� @��q �"v!�a�<���_�[��e`�d��m֩r���Z�<9���OP���VU'�)��R�<�箃2��q�	�+�TD
Ţ�C�<��]�n/��a'���}�Ѣ��<N�9��a��*�f����~�<�kP�0�l���F�K�X�y��@A�<��l+~���f�5�ܻB~�<�s��1}�5h��@(=CRI�Qm�v�<aЈWt�TE�'U�A@@hv�<	c��>��0(C#`�p�[%�u�<Q��1fУ� �R�3n�t�<�W&R�q(<� ��M�XM���n�<�q�J�ˊ͊C�O]~����t�<�bN�0cl�e�e .-H�F�<�� �p���K�޵��g�<9`'�6��9
���7�b�@��x�<�5�_r��J�ʌ\�*���Gq�<��A�K�m���IP���Za�<�T�`52���N��c$$�@F�<Y&,�2>� ��		���Q��x�<�v�@�aH��k��·q^�����_�<����=H��b7$Dr0F^q�<1�H�&�2E�#��0"��Snp�<1�+�7F��6H_�#G��c�)���y��c�l1qE/"'l�����y���	�X��ܷj���M�y����>1+�����e䌋�y ��,8���PL9$nPIu�Ȑ�y��C"_qD���JA�ml$W(B���z�*$ b��wв	3���+b h��ȓlXM;`a?k�݂Sܑy~����Jy�40�D]&���B�-ƒɆȓ1�<��� dZ�L��ȇ_ԩ�ȓ1��]3�^�FY��UCs�n�ȓ����J�oX�)��<#
��ȓtg���"Qg\�0�n��#�Ƅ�ȓ~	��`L�R6�Hx�JZ�z��S�? 0@��#~��lh#O�F��("Ozx�Ď�C�l ���.{r��a"OVR�G�5#?��j��j"OB)B���5�)(���1J�5�P"O���'Hw���Pʓ!e���"O����T�X�aiU�4�K ��y�-ɞ%���S�_:z����L�9�yr�Z:d\A��1v��Y�gcW��y���pe�Ԧ�zL,$��&D6�y�B��m� c��hKȍ�U�B!�y�,�<G�(�weՓ]�\�S5�_?�yBdU�B����
&X�vc��y�������uc��� �5����yoCn5jG��).P#�"�>�y�#~h��w�~)P�C�0�y�_\��-�4E�>}�|h�Raы�yRJ��<m��Sx����F�_�yBa�D���� �Ԥ쒖�A��y��*&��q�C6���!�l@�y�aЎmM0͙���9,F�	V�U��y�lL#4���皨b������y2��B���9��	%@��W��y��"�Μ��@� ��BW��y"nܧ"��L�e�%�1�L��y"�M
�J)[g��z�x���f	��y�̓F�̃�"{���x��"�yl� *�84�4�E�;���p��7�y�aՊ$�ND�"ꜥ-� ��wH8�y�W�a�H��&�) �L�)f%އ�y��
u��C���vo�5�y�<^t8D��D�� �֥� C��yҡх~j��A�:f�,E �:�y��u����v�(P�@�R��y"O��ay`��A' Y�IT��y�kQ<0`�Ȝ�0�Q!p.�y�DǬa�� �3#ړ*�ԑ �h���y��F�o]�SAEP?3B�"�֐�yB&هǨ҃�� �hI/���Pyb��.Q�%{�CR��)�	�x�<7F�V <2�cE�O�͙�k�k�<��\�py9�c�V�����HS�<��.o�T�1�k��1E��x�<��GO
���b��|R�x��Pw�<��	K�S[�bb� �,1�H�o�s�<)�،=�l,�&��224��6�Cl�<q���9U���B�M3n!�kLi�<�vQi3hy*��"^�|�S @�<	���84d�:3�"T=��co�c�<�a�+�0Y`1�ƚ'c�)Q��`�<Ar�\�o9�� Q�M-%�i�fK
^�<i�`��(�X|a� (Ÿ�O�~��8�<����-������D�W���c��~�<YB�қ{�$����<�@Y3 j�v�<�RAVVO��`솠h.�@Cu	u�<�Bɔ�NDp�� �-���XG�<�'"˅Jm.�9�\&#&��R�OD�<qbɄ�Xp]��̊���'�w�<��A�*X�E  �'n��u�§R}�'�ax@�i4i�p��Kf�;WC��y�ɟ�uH��@A� �1r�� ���hOq���"���0U�Ӣ�G(eP$Q���'R�D�
�Jdӥ�¸,�+d!�J�!�D�5@�~�q� ,:�� �*�!� J�tu�$�' ۢ���I�x�!�� 8|ٶΝ�rܤ��G9C,I�����O���D�P[��B�nJ�[�|	do�'d!�$C�om����X�<M(d�dH��)b!���e6�����+8\��i��qQ�y��ɍ=!��th��9O����Pi�8C�"q��͡���P?j�s��VU@B�m��ayG�t�u�"���z$B�	7�8����1*�d-�q'ѿo�B�ɥM���@�h4"X�Wě\��C�	�|���!N�N]A�kF
z��C�I�u0�|��.��t4u	���)U�C�	>�8,/�j����	A�C�,7���N�4J�>���@�B��C�	�k��AK"o�qv	�WQ*	}�C�ɫ	�$�)�t�r*'�Ӳ)*�C�I��P\��i�({���H���N<zC䉞!uz� d^z$�:�(ɢW�B��	#s�|(GN��\��ت��*t�B�ɦn�\����O�yl����Y%>�|B�	�^��d0�o��q:ř?aQxB�ɐ	J0�,H�q���֩D*=�8B�ɘC�I�	\���8�D�+"B�	#D�`��ȢZGd��� 4B�	��d��Ҋv�6D�c�`�\C�I�=J��@�����X�(-ΔB�I 6`�2�GCq���p�F �b��0?��k�Q������L��ayN�J�<�#�*H%���T�Z� �x�g
�Q�<)�N cPv �蝆D�a��CJ��̟���	9,��La�$�#oB�z���#'b�?	��I	�O1n\a�d�Tl��x��R��I\�������4��PK�g��F���"�B3D��s��Y�"��'��t~���tN/D��[0C��m�la���'>�d�Ǉ,D��0'
q�h5Z��垠q��+D��`�`~��[��T�np�-���+�$�O��=��D�I�	�Kޔ���&Q6��S���<)��1[�N�h��� kP<��"K+џ0F�,�{i��b�l�)wh	:��*�y�B��[5K�,���%���i�d����D�Y�{!n�"�K(w�9��a�k��\�a�4��+Ρk�hL��7`&D"��ُM��A���&_g�	�?����~��%�/Ӓ�s��W��0B�Jx��D�<��ㅍhRb�:�!��|���)�P�'_a��O��&]�����[2�����	��y���nB����m2*�.qC��y��.Hܙ�D�@okr���	�0�y��F�l�F��C�-i����X�y"�_MH�$�	��6��43���D�?E����r�Xq����6$���G;��Ox#~�υ� �������`�ѵ�G�<QB���f|�mb�셒5?�İ��j�<��	�C6�����FI; ��ύj�<Y �"XD I��ͮ-/��Ic�d�<����1�;���H������eh<YE�U����4�S*P18�� ���'ў��'V����$@iG�ꘈ!���?����!MCz���e�԰2����"O�i!wJ�_k*��A��?+I�c�<�k�=U�ҀRă��&�&�I�<y5�W�n<�33Oͽ7U|3!�Im�<Q���*�%��g�5h�)k��j�<QҤ�H8�Q�`���b�
�EIe�<� ����D�+R����(j���i�"OJ�X�/��m��+c� �!�<1��"O@�3w�ٰZ;$��W�ݍ{��i "O���l�!z�h�#�e^ez"O���F�u��7`����W��y�@˖L�,�)S&�T w$���<Y��D���X"��[A<M3�M�S�!�D3R�*�)BCj`�rA�u�!��N�,v�)�H��Kl<����!�q��Q���B�d�B� �yT!���1V�� %��I�0�� _*sr!���<�ڂ����P�.t��"O<�R�M�smRڴLڢr�Zh�E�'��ɯNZ�H ��"(��B5��
͞�'�a~"�ԕ<;Fdx��U�
����"B��y��9*[�n\%?~��d-���hO�����E�Hqb�i��"�W$�!򄈈(y4���@�T�����!��P5m�Z��r䏾�L-���[�!򄁀u�0'�X-�f�Ad K
?���>O�\�7ː	[W���b뀪H�>��"O��)1#��@�yD��<��[�"OZ�26 �;5.�;��Ӱ$J(��"OB���Ԋ5��B��٧r< �v"O��2.@1i�aJ��H!�y"O`���E�;DDn�!e��Z:�x�"O숈v�F�]���ؓ*�(-3���c"Op���.O�vpRJ�L1Ȭ�1"O� ��̌D��XCS�2)��P�"O��OC q�t4"�A�H#!��|��)�!?�����^�tX�I��<�C��	<�T1&�Qy�8�TK�*N6B�ɡ|9
}!C�HVJ�a���*2�B�ɱ]EB�"�W W��b�`û-g�C�ɺY�`-i����.P� �U�j�d8�S�O����@�!|��AK�U�"O:�3�퓞:���8eɀ�����0��;�S���7��t��W�T����1 v!�$ �z��lc�IԜIqD)��،Du!�F�R�9�r���Z����ž(
!���A�&8y`��\<
��ҏ��,!�_.^�H�4��4.'�	@��"�!�S)FV�Y2��;���7n�f#!�-\��8��� e��%:�I4e��Iq���ÀgAab���`��m�y�L;D�pH�
ί_��ȳ	֘&q�a#��8D�(�3�1Oi���U5yy��c�6D��1gN�;�P�S��]FUz��'8D�| B�qΦ��D�G�y�dQCP
!D�|�W�F��d0"1#^�&�De<D�0;��<A�l�!���,p�����O�D;�O�P�͝%	ZH�� Y�VK~��U"O�щ�� Q��V��3=@%0�"O�5qS�4q��eC{ `X[�"O))�Ζ�r�Y$��s|�<J�"O2	���ľ9Xvy�΍>H���ɡ"OƱ�����x����lЭ��"O�r��'Q<��%��	xT��2"O�\31H�"GFC�G�jV��"Of�HP�� ������MĬ@�"O�L�	Xd����$�� P� �"O�a�1�ې/��0s�)�S�f�;�"OX�	4@J�y+�59vI��v�X5"O���K�/z���SW*�9)��=�T"O� �k���M�|!�R
ʽ+��5�W"O��@E�C.�tٸ��}}x�p"O�T��l�Q�vR1��Qs����"O��qv@�1x����(CV.��s"O�X��F�ž|�%'��j!ji�s"O^�3�.��+�m[���L����"O�8kĬ���p7�39��h��"O�XxT���t����g��E���d"O��Sq�\�,9�%�
HzVP��"O���rC��n��%�c㓔jy~y��"O\ݐ���%�x���ۑge�E��"O���K7	����0VbE
V"Ot4��$Ğ�$l�A��3��a	b"O�ieꟈ?���E�Ƶi.���"OجU�I2a�`	���.�� G"Oҙr�h��F��玀�����"O�����\�l�2P�ly*�"O�0�E�r�2Pc؂�ꤊ3"O:ȠW�Ko�l؂gh�����"O*AUD�i����Q�����p�"O�q�b鑃8@B-��)�+0	$"O�����P���(�N\$�1�c"O��R��<)MHЃ�H6R�x�"O��:#���g�FQ��G\�v0��
�"O�0���	�� 놦�,'��;0*O��� HE)\](�;¢[6[|��@
�'Ќ�B��[�"޹����Z�8)H�'}�T(`o�u�Q�����
�'��m@��'7P�������0
�'� 0���ٛ`���$�t�b��'�*��g-�,	�VI��a��[A���'� Њuj��*b2h"TΗY.���'Ԁ�FMȌ*�m����KcvIR�'��P�&�%wB��Q�ɫm�%��'�D4���V# �����˓Q%����'법X���&O�\ �F\5>˦p	
�'1X"a�MKh�r��^�?W"��	�'��L�S�[/Da�)�4!]��	�'����@+ɩO�}Y�oD�ȁ"�'��8rP��U�p]a�nA���X�	���yrJO"%`��W�=�ƌ��O��y��ƙG������%
vI��yR��	jƺP�$��(+��pQ/���hO@���� �j�s&�$�r��G#]-�1"�'���{f�Y�2/�ay�+h�\���'�Ң��`�&X)�Gݎ_
���'�V����/{�^��c�Y4���	�'�~��Rk�YU�UrS��T���'S�1���A��;C�T�M���A�'�r�*���D���U�u��Y���.��L9�F�'͐h/�0xr"OdD��dN�?�u9#GĞw���$"O�ж�B�j�b]y��O����P�"O�d��'�VM9���'
�@�"O^�`0�0EN����:f�0�j�"OZ%�% ��y���[��3����"O����Q?��z�ϔ�qB�4�$$�S��J�'@l+��+��!�p�!���09M�yd-��l�F����14�!�Ǵwڬ�iS��w�5�@=�!��Ob̠��tjS�7��K�JV�!����69	T�R/J
����-��!!�L-y��q��i�<�����T�:g!�d̃e�Q���)Wy�pp3L�!�� b1�cB�* �VL����[��YY�"Or�k���2�LI�1h�!��1�"O�Cc'	ָ�0���8� �*�"O.@�l�Uނ0!��=#spu�u"O����M�q� ��e�OgEĔC�*O*e+��^.t�vI�����,'�HH>�	�;�5� 6�tX�/ǐ`���ȓ\5�) ��(�XX��rjƕ�ȓmg����*�@���gLp:]��Z��;Q�V#~�hQ�c1�R��ȓ=b���铼v��@�e�H��0�ȓt�`lS�y����f6�\�ȓh7�C�R,#Xb$B�@�\�(�$�G{��d��&,��N�/߬U�Rƍ/�y��&7$U
	<+��q�Q1�y*!3^�p�%A�⦭y�I%�y""Ԣ0�L�4�X�n`��ӫ�y�
{Eb�٦N�j���-ذ�y���5��1�@�I�%��%)�E���>�O0�Y�@�>m�\݈��ă;���B�|r�)��8i�q�e��mà��"�y��B�ɀ�H5y�᝝9~f8"��"L��B�	!	�l�����ry����#��B��&$U�D4C͌Xh�"[C�I��T+B�W��|�&�H ��B䉪L��	p� ;_�yh��Y��B��|����τr�5�L�Pp~B�Ƀ4{���iV�;�9iw����B�	�7 �3����^=�sN�Kv�C�I��m#�c��B�\H�)Ә/��C�	��L��Ş-I���ЁoU5i��C�	�*�X�jǙ�,��逌6�fC�I�$t�u@��%G���v,�0&>C�	.u�p2,�"Ȃ1�f�4$��B��?�8`b
�T�~ib(E�-��C�I�TD����c?V50�� H [~XB��
_�`3]Y�,�X�B�@�*��A��-��<���ч,��C��Y��̲�k�ja��2����B�ɩ= 2���Ҁ5ِ� 7��f����f���V˧z�P4�Bd�Y%J�gF(��0<�!!��h ��`Z�bf
`�<�U�	\vh<�#ϒeXm�a��C�<�g΂DQ�آR,�W�tb�WJ�<��$�y��8��_�K��� �d�A�<Ѣ�V��f��`��Ԓ��,�T�<a�*I06MrI�lZ�`�My"�'Ƹ�4�L���R�͢r��V���F{��$i�9�T��3��&�ǯo�aa��!D���w�����sdF�-Ђ�Q 5D��X�\$\�Z��&�D�D|pU	rF?D���agP�>�p�R���,�
��o;D��(��J�1���;!m�V�6�k8D�<ᦔ*`��4BC+y&6�"D2D���&�[%���3 <���QpH�<1*O��O>��Vd�
)���d�B�܈{�L�^x���'�؉A�V?߂��P	gw�x�'8
�������扭v]�������y�J�#������̱Z��Ԁ�y��Z�'����ǘ<�6ԀƏƉ�y��'+9����܇{����L��y�ƏJ@:�0U� {�6�F�ތ���hOq����	�3AL$12�r�x@	"�'��{���0Q�⟶W�nJr�X��&(D�� �Ig��,���	4!ԟEXL���"O�Q��	�7N$��QMҔP<�E�5"OBiQW`?}��(:�,��.扚"O\P)X!m��aT�Y*�U����b>��߮X�*)[��[�CW�8i�O �=E��/J�VIBܲ��kz]cD/���F�� �exR���؁ŌM�d
�L�扄�N��]+5$�P��٥�	)�%���Tp�0eQ�)����Ƌ		x�L��D���'-L�(Z�PG�O���`��U\;����I�"0�!@�$����	H̓
KN,�q$]���@AN%]j�1�	�@�?E����"pF:���n*>���*�+cZ2�|b�'?2�4��`�èV=G��Uk�kخ�)Ǩ<D���G��֑�B&ʗ^���r /D�@���� cF@x���D��,D��Y��ו:��E&��D�v��T=D��B"���Q^p]�k�l��%?D�� 恝�C2Ғ��Q,l�sD�Ol�=E��N�2N
0�(��I�Nd!�N��_��Ity��|���K'���C��(V�0�e�!�$�
���s�Ri�L9�N֮�!�˖1�h��(����@�K�z�!��[8!x�	��$d��`���[�!���7�v���J7I��	�j	�!�Tf�$B�=�qu*�/�!�	w�,��F�؊6.��9�L���ry�X�T&?�xϮ��%�K�`7�)���]��R���'%t�Hf���
�:����r���'Y=ptoJ\R5��:w(ȡX�'�ba���<x�����=!8!0�'aP`@%JT�;�<�E��`�F�b�'{��q� �;6�p����,	*���'(�A���Z�8󆔀���$/Ox�{t�ű�� ��G�(�̔��"O� ;� ����El�6���a#"Oش�D̐J�(H��%��W�V��E"O�9jRZ�܊�C��L�p��'����ta��{G I���U�ON�tB�Ɉ~��=CQO�L���C5�M3JB�	�JG���5���
-p&V�T4B�I$�H�ˢm�tт�2?B�	{D�e)t"ְl1����"<��C�	h�<(��[�"
��vDЮA�C�Io� ���D�<C���� �ي
]�B�I+��U�@�E45��L�ub�h|��hOQ>� ��U�?O>�s$�ɹm>�� D�(KRiD���ƃȉvuQ{�6�I��G��'�>	D�_�*(�&��F\~9[�'@`_2����� 2��T�<a�+pF6���O�
��i"DEXS�<a��ѓ)�^�{�� z9��{��Q�'?�%Nļ/~���g+��� �4D��hf�\+@��E�#�9؎)ya?D�г��!-�U��Y[�d�+6�>���O���>鉦��'k�r�G��6�0�@�'D���Fl�,R=l	�@,,&� ��#D���O�$ �dSTKS�D^�A?D�0�N]�PFL�3vU?=
�S�9D� u V�te]�SK7��1��M8D�XDjݰR?�]�FJ��+]�QI��8D���gɭ!ڰP�pa�H��#�&9D����X�S�d�X̓cޘ[��6D��W*�%�, ��P�k	��`�� D�� �A�ֵ#��S��Ư=2�j�"O��DA�{ST���W9l,���"O�аFH�Hv�5p�A��a)t�x "O�X��<T���e`݀49���b"O�|!����lpK��
�y7�BGT����n�S�OlH@b%@ךY|ڀBWhH"̒�	�'��8��l0�x��Je����'8P �l�+�F,�rh@/<cʗ@�<Y7��r�&�8F	��P��V��S�<)�I�6^����ઓ�y#��Aw��M�<�3{^�[�Mݼ	��ə1��G�<!���i����d:Gu�}���C�<����7ScVqq��+��J���|�<iwB��>G.TIfJHUz�`"���\�<����|����6H�f�*J0@�c�<�7���͖��h��;M�D3�FI�<1Ʀ�1?��Ī��*dI� &OB�<��%����P�У3�B��ɐB�<����� �-ᓏ�<�%Ci~�<��B�
D�1r
Z�b��2%�J|�<yw���vЦ8IS�})�ͺ�j�^�<��4�0��ȎFr̴���AY�<�G���"Gʂ%92��[�<�l��Q'p�p"�̲a�ԵI�.�m�<--Ƭ2���P.Z��BJP�B�I��<(�`�-��} ���B�I�;H麂��	G���j��FK��C�	-t�va���B�^�#��D�EnC�ɆE��ehK<LF�i@.65^C�1|:�`�-�-JM���D1D�.C�ɠx���E�XGb�@���0B�ɶ(�,8���4.�&����[)y �=Q	�m#2X�BL�
m�����<����Vn���d�.%�6� E�A2m���ȓ����;c����O�+vZR���0�^͢�
F�Y���O�+��Ԅ�x��|[��!�\P $m�a��8��a�&���W��Hey�l�Y��B�	�%a*����;/������R<c�j˓��9��?�'܈Mɗ%V�	�jDˢGB
G~B���'����5��<tf��-Ժ
UJ@x�'Q�D*6���4���D5�qx�'�|<!�L�B(��@���d?��	�'�4��7,�;H��S��O���M��'f\ۤgP�,��(5��
���8�'�(�񗮄$����m�y���1��?�|8�/ǘe��C��4�E*�O�C�I?#Җ��5�-�R�X��hl�C�ə/f`�3 -��>��d��hC�n���BT8W����f�,�B�*o4UYPN�8[�qQ'g��B�	�� �"[z�Dy�
��\�VB䉄]AJ=�3��T������C�*.'
49��78��� t,���<�	W<�K���UQ@H�N�������a�<�e玙;�ޥ{E-	u���3�PD�<q��̸@R�dbŭ��?���l�E�<��HP"~͐�%ϊ#@���B�D�<	G�@>R鈡�q�լW<.�3�[U�'a�����D& ����E�_Fv]KƠE��?��'�8ؠfX4���e�CH��I���xm�O�.dЗ����6 ��(/�y���!�tY����ՀQ��DC�y�&S�}��i����"Ψ�`�΂�y
� �L���� Q�G!ϪF�d8��"ONдܰw�x�� N�B1w"O6@#��D�o� }����r�ޠq�"O�$��$��u�Ա��I�O�TE��"O �31(�W�&�p��6�T41 "O T�!�*K~�hR �6bb��w"ORm�'��`;ʠ ç�tG��p6"Opu�E8?���FI>t�Q�"ONQ�����0��C>�T  g"O�H�Ȱ>�P��%������1"O���Ƥ��$� $��@��"O8	�¯8��q
��P ��;�"O*C���!?wr���Y��*M��"O�(����@O������~�i"O�ؓ`��I� �����9�J���"O��d�6FW�I(��|�bA��!�$J.�~)���G��TCa��C�!��M�y^�Ĳ�Nݶ>� u:�`H=3!�dڶ$��t�Z!zl	���ݚ$!��2S,�h{i~;7�S�!�$%��EF�6Xc*jS��%�!�d�]v�����]sd��B��"s!�d+]h�1B��WE��P��j�!�DQ�#BBL+@Ġl��A+��_�!��%��;�N�0*Ī@��P!@�!�dG8_��s�N4Eт,�ũ���!�����h�e� ��x���t!�$-��AV��/��広'\uu!�$�/_�l���P�J��T��E�^~!�Dݻu4���'\�O���!n �KI!���.Mٔ�b�
B�N}R�I.շE9!���TBl��흊 `� ��ݛP�!�^�S��m��ɚ[#�M85B6@!�$���M�y�����P�!�d�P9�d�����"�ܕr���>�!�$	uR�<�fJK�&�4���(x�!�$Ƿo�>�Jת��+����M<�!���,bP���R+�D[$d�w�!�d�o��403���3� q��^-!�!�Ğ�r���AT�69�|D�4��!�;f�1ƪ�g���Pd"� $�!���?���c����a��{D���'��h�HO~�l� �AM�^�l�'Wryu�Z�{�&�P���41U@�y�'

}jW!��#�f��F>�����'���Ӗ��zUڢ�(5>i
�'�Ε�v�Qpt4��Ưyz��H
�'	L�ak���d���y�h�;
�'\��ŭ:T�<m�4�N�p��i��'��4��]Fu~�����ve���'"�u+A��zXV���Ǟ�Wy����'?��&�A8	�`����L���'J��'KT<T�T1�'G,jP�@�
�'�TDl�+7�q�1��go���
�']��� �8+�0�R`�;tQ�$�	�'���K�Eүe�h@�祋�vRy��'���x�"B�{�F�I���k5zmx�'��0���� J6P�S@R`��(��'<�4 �iӵ{ܜ#)�W;^u��'Ѳh�U
�L��@h��W� �~Y��'/>�;B�1+gr��!��(��'~\Y��C�Xz�L_�[8H��'(���+i�`d�u䇟:�B��'�0��#��:B`��DDC6+�k��� �D�7`X�PZ��@7�ӋpY^�w"O:�q��̩(%��"��� 4j"OnHA��Ę��-0C!�5�H��"O�]����{N"-@���1`'�iqq"O�9S�e��t!�Ī��D�ĸL�@"O* 2��a�j(Cq��+G�&��"O,��6�ߛJ��Q&��=��, "O.D���Fe�-��`]�Xx�"O\5+�㗟fl`h�5l� �"O$���g������`G=.R4%"O�ŀ�-ʗT
��ʁ �7��`-�yr�V�b�4I���L,ygN��6Eä�y�"�>i&�IP�G�D��j�؅�yR��e��	�<J*h���K��y��'���%��8.mb�a�IS%�y��Z���K�]K84�����yrK�TF\��6g�7R���
�M;�y�@	~�,�� �E0,	��ʁ��y�5wk���ED/H���r�ΐ��yrf��H�0�ě�<V�!�l[��yb��m��T���58�ސbSe�3�yr�����gD�1|�b ϙ�y�a��P�^�)z�а����y��bW�I	�GU:1�PT��ǣ�ybE� ��Q��	+�YRF�	�yB(��A���J@Q��6-��`���y⭎B>��C����jiT ��yE`��K�@6@|��/д�y��+�\�c܌Y���	s� �y�L�Ci�@�B��>�
`j�����y���J��]�m'��Bȥ�y� G	o	�T�BnT�`�@��+�y�%�`�ycP"@�
h+�i��y�^	��A�!_@=ʈh��R�y�&��TJ�9p�ʋApP�{�̝��y��E���`JÁ&"���R��yb��ǀ!�FF�G���3�Q�y���E4�k�d>�)��D�(�yB�(lܹ����`���	�y��Zd�})��\U�$��щ�y�'Q�]bs6lDӀL�&����y��تCR�T(�A�Wf��f��;�yr	�D�s�8{s���;�yb�3_�&a� Nۢx:5�%]��y���$-+j�4g�0r�V4�BJP�y�)��'b4�PƉ�3i��=�E� �y�9=�4	(�*
j�9 D���y�Ӥ`�����0V��x�"& �y���-�8�怌�ݪ�b�7�y��-J���+�[�'&� Q�2�y'Y=i�Z�͋�a�(��K��y��	�E=�� ֿ��y�`L�y��Z@�~�q�dW96!B��+�-�y�
�5��A-��5u���4Ɵ��y�E���T��@ڼ1����s�J(�y�O��YN�1x��aB�W��y2'��r�$�ߒiٚ���B#�yr+ɏ���2E.�3g���P���yB��	�8i���^��Ԩ�dܑ�yRȓ� �� `ҶN��U
�#T��y��}���Q�L'�a@7��y�Q�F�h����)A���0gOA?�yn[��Ppɀ(2\���R��y�aR1��	��&�(A����c$_	�y
� �}�v)H�N��3��#Fy(m��"O���v� ���i���O�p�.ၤ"O ��]>�MZ`%0Z�d��"O�6l_)��L�F)/}�)"O ����5��UA��E>x�zx��"Or��0Ċ;/f*}�&�@�[�V�b�"Oxk���2�X�׌�o�<�F"O��@����h�z�KׄK L!�"O� �Ʉ�r+�|K��߀6�Ν0B"Oj4Zd�9x��L"R�`@F"O�	�$�L�#zh���L�VD�X��"O�aY��K`<��k1�_�0*8(� "O����%OUf)���/-!\�@�"Oj��k��xC�-s�8��"O�<�r�
^�(1��b�1�84{W"O-9$�_�>�h�Q��w���A"O������T��W�[?Z�Zju"O�)����n���R`ߎh��EI�"O�1��C�:��h�`F
IIpq��"O�	
c/�? #��1⎛�i��iCS"Otˆ�Ѩ:rT�MZ	aq��V"O��#�m��-y�)��kp6lID"Ou���P��U �	�� gn ��"O�a���t�P���B�9�,e"O��$.X��XR���B'���"O �'5w�\�ȓ@ق"O�%@B��}.����I&���C"Oh�+&#J�T��	�Q�,�h�"O�4�#CPn�<V�$(��Y""O���"��f�p$�W tBP�3�"O����,aC�h�Q��
H�|2""O��s&��O�II�A��}vT�"Oꄑ2�6 -CѡN���=�"O�i���9������5�MQ�"ORI:���9|�ܵF�W}2*��E"O
!���/$��#w`�&T�LT�"O�!(�\�	"L�BΉ�*��M�&"O���O��I!����MZ�|�$h�"O$��0F��c/Ѱs�	�ab�0#�"O`e�rdБ�41�a��]z�	$"O�ds�IȂn������B+M?���"OR��IM�^(2��A�%�:\�"O���\bZ�lX���2�B�0�"O��PŎC�;�bc�ҫ��
�"O�a&�$md��;�DW�z��U"O"Q�#�ϓKV8�`@c�+<��r"Ot� c�T?=��q���B?.	P�hb"Ol�rǉ��#���!���I�hճB"O�(��x�a
G�(@���"O��s�ŵz��=q�/�6<�Z�"Oj)����% ��c#� ,��""O�Y��k�;d;j���ȣt�B�6"O~Q�V��Z�l�ab皲g�d��c"O��ϣ���	�H���E3"O�8h�g2Il�4?����J$D�t�5iF R2�(���<K\�	��7D���$.�&�D�s)_�F-��h�8D�Dsg��L͋��J���h��:D� �PL,�Y��&^jd����7D� YGɖ 1RTT�"	�g::���K4D� q�ˎ],��""�[ac��3D�,
t���\ȲQ�<GcH��N3D����=y�ri�kM3�o1D�x��C;{R��2�&���4���k/D�� `\1��ެa�blHv��^0����"On<��DL@���*46e�w"O�=�U%I�{�Z��v(�4x��X�"O~ ��A�r��ʞ;��t��"O"�mޠ>�<$Sc��?:9�p�2D���F#	�e�!���`�@���,4D�DIp  ~��H�`��E{�� 2D�A�N�h+}�D�^�0��c%D��b遲B۶ыũV4
*��f8D��BAҋ;���gh��Hh����5D�D�c.K�G3��k��:Y��up��1D�И��c��С� ! ��"d0D� �V��-�V] 1.]1%�ɛ�.D��V��*����ڐ{ް��m0D�@c�&�����W�T����`.D�,�������m�f.�A@*+D�d!q�B�qDT��֫Ɨ��Īł5D�ܐ�C7�5���H14*���%&D�d+0)m�
Ԛ���$���IЪ9D�`����I/�X!�nS�K'-$@7D�Йf�� �<1����&��K�/D��P�G2���vL�ӦL3��,D���!%��&4��,;�ܙ�i8D�l��Gɧ�����ǅ���Aҷ.7D�Ѕ�F�L�Ђ ��f�X(�S�5D��w��)�X� �����z��Q��yҫH9:1�g++�@������y2�I-C�
 �#2n �b)ȫ�yBb �c��I����.�(���@��yҨN�o$>	�`W�#t ��#��y�	�*h���1Tȩ%/�9�y�A�*�a��%'o?�L��h�8�y�mP�j�ͭ2r����`�\f�C�I��:�엠u��ʲbț+}�C�ɹHp�$���"np��ʑ8��C�ɍ:�����  S܊��#�T#P�C�ɗ�����2���燘A�C�	"p��iI����}�, 䌆�G�LC�	�@�����&�4�,�t�O=�DC�	�W�H��A�b�0��D!P�.C�	4Z^�����ծY�H�
I�!S�B��&q�j=�d��
��k�C�p��C�	0O��H��Ey[:�*¢ ;�fC�$,�ܘ��M�8�$|�EɈ>7��C�I��n�b�fN�Z���X�D�p,C�I�@"9'�լ���$��*: C䉉'�·�6��4P���(��B�	#<����M�A[�(Bg� #�B�I�nt}����Ѯ�0U��0f��B��(Rn����� I<RвR��O�.B�ɏ��IF.֣B'F 3�&�0.B�ɓrL>���?)�0:��%E!B��$ÐᲨ�u[�P�& �K��C�	�#톉���8z(#e	<2�C�)e�>	��12�iIF�R�^B�I3f���qn�Y$��@���NC䉋�Rl:Ri' -�VG7q��B�#_v�u�B�3)�Ui #��avB�	$� �
�Z �n�I6���%��B䉟�|RuE	b���#��>h$�B䉠o�1&!W�@I)u��#�B��+Dj����W<"<qh�f� 	ҐB�	�b�v�!˃qLX�H �LB�	�,<�}�U�ϳm�"�4�#iLB�)� حM�2,��@�f��9�"O�d$��c|��ő	�	T"O�8� �	W�.��)�s}:mi�"O�Tc��	��T�2*X�D@i+�"O�e҂^ H�2��)!Ό���"O�L ��L62$�#� �p�d"Of�Tl4~8a�ud�7(�b<�$"O&�pW�ko��
4� �8�"Oh�x��H9`�ikf����0S"O��F�%nn�����3��Б�"O`h+��ϙyv!��� ���0�"Obd����G;��"A�3j���b"OV�
5Ûq��qڅk��	<�3"O��y1�Y��eK_?G$��iw"O�@S��!�	��̟4W�)0""O��h�:V���*t*ƹ�	{�"O��vNE3�!�"Muή��"OD��U�^��$=�U�\��v�+$"O���bV�x��;F,�)T�40J6"Ol�q��CSѐ��!.ݒ�B"O��KA@ O���Q��P8�Ȁ1"O�D`�1��
%�0�"O������<�P��W灚:��Q�&"O�E�gAL府b7e��*�:R"OBX�F�K�y!��gƙ�[�I	"O��#���J\l|�Ҏ�YI����"O�U�f�L�%N ̛A�596�"O(�b�X#� �U�߼E5��0S"O�ը���G�*�gi��a*l��"O����'��5��[7�¹X�Ӏ"O�%P�	G,>.���@(S����6"O�]�!I��t� �8@�Z�p��i�s�0��`���
�͛:8�Bڵ-f��`F�6D�!$�ڲc�ȁ�e�Z9$�� �gӸ�=E�ܴ6����5�'��(���a����c��|tVx`O3�(9h�;2@ʸ�ȓm<���AoҤp�4Ac��J�A��U�<�����Z��� e�U
��	9F4�!�ċ�z�,�b �K�h�&l��d�� ��IP~2�)���^�th �v���B~vP��EZ���x�
גM	�A��M�D~~�3�єo�!�d�.D��cv]�Pp$�&���/�!�E=alh�c���Ā(g��4H�!�$�>F�FT��L� ��x�M���'�ў�>)#��&~�� e
�I��r %D�L
�m�Z����!L�;}�y�1o0}��Or���>�"fF�hy9�l��5T~�J��h�'��|&�$�}�Q�ֱ]�Ȥ<𜔢�ǇO�<2*ƩU\�kgKϽ��R��H쓍hO�O�b�+5/$_�L�tcņ?o0tb�'\Z�I��B��T�R�4�Lu�H>�O�b��>�Q���6Y����o�����[�?D��sƯ�F�(<�B����
�#8��Y���kč4���d��3x$��EE6�����ƔK�x�KP �n<��=O^��������)��j��B�
R�&�a|"�|B�Q7�	s��#��d�Q�Қ�yr��2�<3$�N�	�\!����
���hOq�ִ�W�E��PY@��!<p�0"O��Z��	�d���ś�0� h�"O�e��YA��;:`����!��\/*���06�ϓ=�d�%h�5uA!���F�t��� �F٨�l�6�!���0��h��א[ʦ�a"
3�!�� Jeh�I��?5��8 ��Z�A��'I�ɯ,�0A�Q#Jz8��SA4=$�C�	��ް0�׾w�E�-_X��B�	5'�RѸ�M�<��4�q"���B��uv(5��F�b?py@��dS4C�	����f���zc�9Q�B�hWC�Ig��!�R8)RP0q�Z��B�	�y X`�F΃BӀ��ɀ&�B�	�����,܁�ve��F��v�B�ɣ8t҉������U�����Y,�C�ɪ_ �D�V�D�tT��$Y6o��B䉩;�^��g��7^�^�3AC�FC�.?���Ku�
r^n��n�7.V"=��t@RY���*B$�Ӣ(F� b����e��L9��Y� �y*�  5s���?�
ӓ{��IW
�i6��D[$��Ɠ �aI�� I��q��/x�G�?�Qs�y���F}c�2>�I@t�ѯ��L���ʹ��=�y��N�%�|�b恉�tS@���oK ���8�Oh�+�),J`�Tc�>4?�UQ`"O.4�#��.'���9DLpW><�e"OapD��3��|`�%�9q�Ah�U����ɹl6���^%r�xB�͉:@C����Tz���2�D�Lư8���w�?��p<��G�f�f��$�@F��d�Zz�<	g\�� �����1K��!�ѦE��8u�h`��ʻ<���K��I����ID�J��8pf��
��s*�^��!Gx��'4
���
)Gw�` ���:�d�'�"��N8���G��9m�<%�S��0>�H>iI'2�Lm��עC��A2$�O�<�	ӓ�ēM��UJ��02���yA�8��IL�'�X;C �#��EPcǥ0������yR���'j\�� �A�8�3хOP�NDyxR�i�E4#tbЭ��E8qe��uY�I�����IO�b��B�V��Y��^(M���I\؟\S�S�8c�,�V&�`���T@%?iÓ�ē{b��я?N�����Ɔ�AHd�'��}RBJ=��Q��GϝQ����/�!��>���>����.0� ��uB'Mzt*FKPm�<	AŃ ͈����7�"��k���j'��n��J����3�.4駌L�5�f��N�ȥO�ϸ'��諴��>cWu��Ѱ'�F�1��:�S�d�@�&�dxy��;}{遑-H>�y"H�g����`)q��%Х�E�y�4͘��e��o��=+���y"+O@b�����f��im����TG{ʟ�9���q�����$ȵc�C"OЍB�HA�I���H�f_<xC�`��
�}�������8r��"juc�Pc�!�$H��f� E]�j�f�rD	XJ�$LY؟@b�i��#.<��٦Wa0�+�'2�O�O,aq�F4q��:d�^@z���"O�)�R��R�D�+��AQ]���'�	
�HO�~��I�$�uF�p��*	�E�����2�ě�$����GbC�ԛP��$,�!�[�
݉a�	�X8��EC�)��O7$�S��N$@*����߀�8�:�� ��y�i
*�(|�S���|�8��'���y��)�'x�F]!�M�,݆�G��53���U� ȓ�&�'>�2����]2��ȓ
?�b0��X[����@��	�<9H����dW<䈌@��1	��A%I0D��!���	:_�=[�)��H��;G<D�� �lac�@��j�ɇ�f>��"O`���-^%�� E���� "O���� (�, /�Z��"O�9G���Xl�=��4Jx(!`D"Omc3(U'r�Nd��i_�uʲ��"O���̎�w� ���_�k]����"O�iwJf��8� �]�g]>p����Y�O��=�Q���D�Y�L"*��	�':2h�rLԆ7�Ăs���Z�
�O����S��>Y`�؅$EvPr�#�2xtp.a@B䉖��x���OKpy2g+�!m��<)˓x�!"��Z/9�r��L�#޶�ēU�l����T8"OFiJp�c�x�b�"Ob,(UfX�a
UB���E�!��"OX�+�:�Z� r�=%t�<��"O�i��D�ުq��FN����0��,\O��b�T vz�+�.��\wxy{�"O��2f�ǇE�qHPL�4��LIs��+�S�S6oH�
�mE<<���$�XRj���$�ɡ|VP%8$�O�	�u�3ώA���=��0s�_
A�`S�-@>c�� "}�|��O�a�c�V������7qu0m:t"O�y�����|p���S�̋���<��IJ�'	Re��/�#0HQQD!�Y�#�'�����̙�� �>�B�=D�P���.p�ư��Q�M�!f8D��H��Y�-FܔБ*7)�&i�N,D�h�E�,=��)�𣎁[]Ɓ�n)D�\y��_�Y��i����i^�E���%D��B��V�tHlۧ�n��b$D��z�`��]@�
��ڥa)����/D���3�p�:���dI�U��C)D�B���V��G��:� ��
ahB�I���@�/MTt��It�RB䉣$(ՂGb˒�r|�A�|mB�.jQ8أD`LZl�2@Ř3�B�	0Fs��Y�ئA�n��7�֦<�bC�	�}��1�d`��!Q
�y ���v�B䉏'0�,�MJ<�0ۅBӝ�rB䉊 �pxccf�,S|��2���B�ɲ�����W.!�>�s G�I�B�I�,�^�`76�<��၅4,DC�	�Itt��%G��Nq��D�qy!�̄*����e�" ~j�f�I��!�A{�Ɯ[SG.oUp�D�6!�ؑ��"�N�AixI0�D۳*!�ǵ؁��@!��ɠ��s!���fV֐"�)�d�� ��pj!�ē&p�B�p��	��\sF�G]!�dے(q��b6̓(@���7&�H!����g:1�dˊ�:j¸��J��I!�7
XAk��:,m�cH�>L!�D��{���2�j�{����烘!��ފs~�)�Cm�2}�9��Կf�!�$�#j�r݇�@��fH\�b|!��Зeg�p�%H�)%:!,x!� �Px��gn�)�a3a!�R�|�ꕓÖ�H���z!��O������G݀!nŐOd!�$
^&��!��,SԂ  �)U!��4�F����,�4UB��G�ME!��K�h-鄥���<�� �4-!��</�,upb�D/]��1PiE,O!�ϲU`�x�J�x��$"c�K4`�1O�Z���g��#��N�f��X�7�� �Tj4OD	s�0z��Č,���Ӄ"O�7/�Q�R����,odIs&,"D��X၃��r��sd�1�\bf5D�D�3j�H#$��I�,�.I��3D�h��Q�������/k��Fk0D�8ՀB�~h.{�hX	U<�9hbF8D�hJ��ԝg_�px��̃7�`|���4D�P�&��%�N`��*t*��@�0D��h�
��=EБ[b��&����N:D�\P��D�d�� �Ę,��ESЄ9D�x��Qi5�56-ƙ/^<�g�9D�L�%��,2@R��F�p�&H�!i7D�|�EM�`�a8�ıe��7 /D�c��i*��� �4�0#,D������ �0��FL?��T�6D��r�e�t�����k�k<�ar"2D�p�uC��?�)���[�$N?D�X�Xn�|50`L\P�X!�3D�P� �ZOZ�zD*Q�*ʶh���3D�T�`��"]d���#K>4e)��.D��c�� =��9���Jl{̄ХD/D�� �h�3:aH]7� ڒ�,D��q��`��uX���:�$�:�N(D�h�R%E�pL��(g�ܴ8�)D��B�ǌ2�@�ɗ�u{��ڧ�$D�l�#��>^<�����M��h�E�6D���!�E���ы���V}���È.D�pXt�	9\�H�٫&�i��;D��x!�
@%���ؠ {�	��%D�:��_�8�$��L� \��!� D� �E �-D���AA�^��8p*O�����j���#���&p��\�#"Ozc�ʏ9P�)��L�� �1"O��ɱMްa�Z��FnK%4�����"O��1/ M��s�DT'"�~��"OJEyqk� &���;qe��8� t�r"O�m�DV?Zw���$�o�BeC"Ohd��îG�lEY��=rtl�R"O杩��n �����IbH<a""O\���@�Mvi��H<sl��5"O����\%��KT�A���0�"O&�Pt&�i�Ⱥ��$�����'�*M�EI&: �ɖoP��Y� �"�@��BgQ!\zB��2g�`�ӥ�]�~peE�*$>&b�`.O�&;,<c����k�,$�@H��7�H�FO�O�C䉟@����KHE�A�}��1�O�0�ʓ=��!���L�(�G S27�r�q�)� ^���Q�$4�h�dbϐ[��)�$�l���(�M �$�MP�JzȆ�	�@"ൢt�׺c�Dy�A64�B��ė;`�\IÁ���7�F�0���8 �D�UQ��mJ
B�I�Š�3�O�6b��Qs#�+��O��iӣU-�� L:�Q�fHc��@+S������CLƵ�ȓW�xȅgR��p�ߣ�D��O��Y/栕'�X�B���>I�q�v@ C�����5RǇ�Kh<����!�t�1x?�A��	Vy2J�Vv��`��d����rC���j�c���L:����ɚ �f�[�DܔO?���	0�T�A(�*�Z��i�W�8���U�����8�`&�@@��<�@�LBE��q� ���s��JL����+)^X�ȓ?�|y K�;-�A���n%h铍Ǒ��'$lE�,OT����as�t�Ɩ�8�A"O���֡�=>{�09D% 6U���"O���U�b���,e_4�7I�A�<Qs��<Uz���J�{� `7��E�<� Tu��l�����'��>d��"O,p�u�Y�=��೧��f��"O�Q�2��v���h��*=�����"Or]�P��!�D
���Xq>8"ON\�Q% ��9��Q.t�����"O�p��b���%˕g0`x�i�"O�|:W�
�8`S�C�Ev�A"OT8Q�U=Jzk4�چ�05��"O��S+��b�K���(G"O�x�F�·\~ʕ��J�1'��p�%"O�%�3"T.,Aٷh�\$���#"O�<b#�&��,�fĞs'��05�>Q2�=4�J0�AJ6�>�+u��4zC"љQ�ׇQఊ�"O��k��Y�0�*�oOs�6]Yb������=s�Y�$��L�g�dö�
Ѕ�L�@W'J'vH���	eƺ���B\ÜY�(�6I|� @�'<-(��E�4	�a}"����s+�<o���J�@H��O��
N�Q��A�����ÿ Y����O��−�m�!�DE0 ����:�5�U	6�剄xH��r$V&N�(hz1�.�ʅٶǹW��t���3npC�	)/��m�I��$��	)�O��⪙��~R�aĖHz ���{b�S�2�� ���Q�q�`�kG�'��?�6ӱ4�:��V�mܨy��?��C�.Rax}Q���v<��ˉ{��	A�Z�ȁxR��fh��2Aܨ4�џpg��'*���q�ʅ<r���*P�"��8pŞ�2#�f� �%���r�]d�$b>c��f
�*h�dQ����y#��<���پoz�ʗm؊rè�|
7�+�����O1&�`+�A��f��+�`Z�;����Ą3��r4��MpX�+`X�F<aC�>���^����Z��_@J�
�$:���'3*-�u�lb��=U�و�'� 1ڵbb�&��Ԡ?k�3���0/��Pp�B<B�s��2vOR�O"|2 �G/�Pa�����N8x�T�o�'��E%�s]0�$>m�� ٕ`�>�s��D�z%�л�钷�?�m�9]N���"ʾ� �3����wa�0d�ҕJ�(4v9�'���[��V)��ؤO�	����𕨀�~M\��D��}c��݆0�6�i�g��U�ԅ�	�3ezU��_0n�x ��_�S���(K��`��=:��5�F�-���[f${�v�=�y' &Ni�f�����.̚��?�q�� �T���2xV5� �e��J��
�%���'���r�Lq��A�D�W[��<Q7��#�P�8N��+���U�B�'����A;�@$>-��.J����A��5( �ҟ\���ς�
1� 4�-E"��[-L�����^�Ӏ�I
���C(4��C����?5S%¬##.!%�; wR�[D�.��My�jRS+\�P%���O�'��A�Ɖ��$BF�S�-�,��qO��2'J
XG���B2�Ե�y�RL�h�ؠJ�=v
ԥ�E���?� i҉O"t@���E�6,��><V�<
��B'}.Eq�)#�Ɇ&y(#|n��@YZ����Tlx�1,��J���$<=]��B�8��<\pjt� &WlP�"D�E]!�d ����d�Ӽ\�"|�Fn���y��M�B�<�)�SK	��!��C��(r ��=҆C�ɣ	��tb��ŕ]�ā��i��x>�B�	����z֍F�ԝ*vJ="8�B��&�f�藀�0{g�q{�LO �nB䉣9H-�`À4Q4i{��C�vSHB�	)�@�a��+�))�h�JB�ɬ[���eZ�S���Kbd@�Q�4�<�
C�Z�"~� �AR0�%��/^a�dH~�<�W��Fa���E�)I $��m�'x�h@D�L���S��y2 A$����1O�^��0�O��yb�M:?W��R��� !X0g�*�?�S�X�&�Nr1)0lO�,Q�B?�t(�A��X�H��`�'�8x������Iڴ$a��a6���TJ�X��ON�;~�(�'3P-�rm؞�a�Gշ����եQ�d��$#�(v\>�8R�8����O�h��DCxV�{G'�B_�(�� '��m8��#D����ŀ�=K^�S3��
8'���:LUd��?�~℀�m��Y�"@$����O@�Y�;!|@#&��_��PS�����S�? �D��e�2�H��3'�	� l�S�	\(ka���<w�q���;��L��%�1�P��C�����I��p%��>G��PSs�*����Q�3�̠I�� =Q6��������Gd�����T�D[�v"�9;�����h��P���r��'���B, .��1��V H��{���*�m��%�+b)��K�J�B�@��?��;�z��D�6"�XIb@���D���*&d���:��y˃��#PQ�����
v`��'
\,*Uň�?�0�8�q��)At�ݧ��@��.BYR�	�!�,zW�B�ɶ?]�d&L�R�Bc%.x�t�P�ЖOj�I�İT1����6=E���P�@�SnyrA��o�a��e�*X���n�3�=Q%��a���y&�B(cܮͳ���;/����S=/�t�t�<	���"��=6.��b�WBD��?Ѡ��<CI���F��.1�<(S��Sy�+��G�� ���=6M0l0o�}��]K��L5��#�Bv�KJ\9p�҅ ڊ]5��.�Ŵu؅�'R�ܲ�L4��4�M"}mR)O�: � 4�����=�0ts�� .Z��_�D���v��P�� WW����U.H/2�~���y��Z!�݃5�Rԉ0�	o��XS4O�=_�8#��x4��̍7F��kqŝC�$"[15�˓��iA/�rL@���Ӌ*U"�G}��7�fxi��Ky���d�<�s��?w���zp ׀!(�8f�:Eh\�;'���d%P��a�2�?���T�"�(a�B�LE" �ӥl?yG	�]�MBA�<��J�% hQ �IH�`�X����;C�,[ � �\�{�Ϟ6a%��Ud���Bjڦ�@!e/I�n��@�����"�U�"�C!#�Ze/~�\5��l��|��aP���2|*2�f�չ~$� �����p?a��P9��B�FH��$��7&Z?A&]�#ɔ#k�$�`H�{e��A�%>�J)z�(�<�6©`G� �ǀW�I \4b�ÃR�'A(�J�$��{
p��|�֮�Y���T��DOX��R+�Q ��˜���5���	n8�L:�g�8}�bBubq��ίf����>c4t4�cK�)Uw�S�3�K(Vst)S��Ӳ8�%s$�<.�����44<���-۲�Px�)�y۰,┉�>\J�qY1���ē}�������7�<yK��@�8����'G�8hh�(Ǉ�ڈ"P��gľ��	F�<`ƆS�\BP���c�Bʴ#kV�al<��UDĬi0�X T��E���d:$����2b�H�X1,Y.2��ȓ]�%	� �S��Aqa_�^v��'�FA8�GD�y�rQ��ɘ\�tD�bd��kp
c���>`�0���\�b�>��e�-X�v��!� ft]XSDX)�؊�'�JU�(]�"s�� �*�A*�8��Dߩd�KpD.�Ӭ�B`�g�Lp2 �yD>F��C�	�E���s�+ީ[ �֡k�@�I�Z�X�����!N$�q��"9����Ӯ�]Y0C�ɽBmJģS�P�Cæ�� �W$E�C�	$Ǥ���a��TY��˖T�C�I� ���3-������H�CWnC䉨;4�E"噬 ���Fǩi�ZC䉱C�y�4Ǉ�]��p��| C䉕q*��6ǜ�8�Je�L��`�C�<�,���g���u�O�-΄C�I/�T��v��AQ�"F�,��C�	*]>�3.X������Px�C�I�8�H�ʡ߱Ro`���� �yK@B�	 $�$H�U�ݤ$�6����2[�2B䉻#SZ�{��ދ<.(s�)j�^B�/�F����Z�Y.��D&�#�C�ɇm��Z¨�P��b��V(Z՞C�I�Kc��r�
[v���]/�C�	�WV�9{C@��()�HU�h�>C�	�/`��r����j%zɀ�.ōj�B��)�*�RlG,L5r 焪*B�ə3�BL��T�^�f%
� ?�C�B: ��d��Vp��0��q�C�	�6�Z����N^}*�M Z��B�4kΠ��E�J�&Vtʖ��� _�B�I�hR�����Cv��F�T&b�bB�	�Kb�<�� �iK�xR�U�@fB��	Ʉ� �V+��,�5��:��B�ɦ6C�$`AΫ^91�*k�rB�	+����m.7`]�5n�2V�TB�)� ��93�;U-����Ŕ!zG"O�I*���BNcR!�@�:�"O�#�^�$ �� ���@"O���l��M��їp�~yi��?D�4a�IѐH
Hz��Q�W70ɸ�.<D�$8q��.����%����M;D����  d��Į�8b�2�;D�8b�'Z�+x�{�c�1xMzӳ�;D�`xw���k��B�D=S�v88�-7D��{R���8�:�E�&m�Nw�2D�X�f�X�o���s��ܟ%�8���5D��e%O&F���[���<=X �Ԁ2D�ܱ`�Ԗ`�|�s�&[w��8���6D�T$$�?( ��rGby��u	H�o�<!Qi3���cBGq�l��!Zj�<����8�r���V �t�ҥ��S�<��bQ�q��yaH8rla��^e�<A���+A��%*�Z�nޝSŋ�{�<��a��L`8����E��Uc���w�<���QmŦ5��ܯ$��H
��	q�<y@ܓ+�C�KS�T���rf
Nn�<iŬ<��@��F�:�� A�<!2i �6����F5����Z�<�Gä��I�������U�<��	"}�f��H�3#]t��ĕX�<��f�0D�T�­�.W4�u��A�<�F )�����)J�w,T�Q��C�<����Hd��"	
9Egf���B�C�<��n,D�ȡ��9-���',�|�<�Ɓ$9-@�;Ё�Ų�U�y�<I��ۄx'��WjV� ��A�KR�<�́Q6�� Q�ߜH��rN�<q���:L:��#�5b�� �rA\m�<����&1�v)� ��L���FQ�<����=*�jw.
�7�Aȇ�I�<�C��=�����k�>2ڊ�� �\B��$h\t�A�+ ������8B��1"-����h���IE��"$�C�	4j��Z!˘hO���s��?X�B�/)�n1����L��-�b�UC��3<��ĺ5��Bt�q�d*�2��B�I�}�\���Z�o�DIh�/L�B�	!KMz��v�8]�<��p���6�B�	O螡8E�è:[����&G�G�bB�I!p3�p��Q;�&��q�b���"O��'ߵS��42�&'`h��'��Y�I�[o�I(gS�Ea���d����e�1B����n�Z؃#����D���H`�<����>�Bt���%�'P���CR�S�t���Hį��C����Fv+[�I�r�V�P�D1c���'@<��F��>�4�
n� ��0M�rg��P���wh<QQ�\�F>2�{S����b93���j��:Dc��2-yx�|<���_+v=���ۛs��x��I�],b�Gژv��pϓ#��qϓ�#����Gė�2��ȓ`��!(^��D� mސD��a%�L�P-�C��QY6n�_�O�I�DO�G���1��M�*��'����@[5\z��Q5DD��J�8�
�;X
�A�-OjL�b-�3}RjV�A�&�G��RX�H���_���x�R�m�e!�
�$�J)���ՎV �qF�E�k2�'��p���Y�3�~	Pw �iHJ��3�th��1jN@��'2��e�UZ7���u�m�D��'� x�7A�z�A���!l!��r�y��̠n$��Z�O�G�O���0G�5O��r��>��4�'�LC���.f��X��R�zpe���15;�Orm���Y�� �P�� j�{���6mA6iW"OJ���_24�,�@� ��[�e2�"O��a�+H�ȉ���t�
h��"O�|�Eeڥ[�T�S���!
��4"O�@���ͱ+�nTH&�A�&F	If"O�`��k��e����l�-7��#"OVa�ba+I�6M�3�Z�.�!�\�Y�����@ʆ���%L�>
�!�D�)Fb���F�O,���FL�/Gz!��цFTh���U:�e�W:DE!�d2~�:���"R�F�z	*Gʍ�`�!��-a;F�G��<�@�i
�T�!�C�u�~X)��0�Ji����p�!�P�hؐ�%�I�!�U����!�ą�L�lmʖ��80¨�b@٫O�!�䒯J&����C�F��h���<+]�*�����A�xT���(���c�/I("���D��5D(!�ӆ�d��� 7� 2R�ӢA�0y��A�<�H�M�=�|�<�)�X�	#�'V&/oę�/Y����S�[�O������%7�>�D���0�����	M�H.��>�dmU�'5�9��G�k̆��FPI�'���FH�=��[V@�Z��A�$t]#����@E��'`X �y
i�M��D�0��Q HI���DJ��ڬ;0� ##��ӈ�� ���ɂ�Ԙ]XzXh��ǈtl!�d��m�F]�F<T|`��Ԯ��}(i�&�Tu?�SCN�p:��#I~�>9��S7^���J�D�!*9�O��0D���@׫K�;����N�B����  wK2:����n;�I]�'	����ɡ
3�P��D,�D�E"��"�>� ���hP�Oo꽳Є��rAT��&GB�j�|�fG�@� z���y2��12|@�ag߼h��PtEY+���@�A��f��Ek��)]�d�����dJb�nѱ���J �NH��(�"�|c�h�<I��� ��E$Y��5
��@���d|&6�n�!X��vgj �O�|�r&��eyj���6S�� r��X����f��X��8��,�����=n�YA�Ad���`����Ö>��� �H�ܚ �F�@�����jDџXP+�;��&��tY�P4|L�6b�:'b��9Dn����i B�kr���E�����hO�Ր�-ǷY���ō0���_��M;� ��>�'2� �c���`20E��%�(aa
1���ʎ�R9bTK�.VV�:6�'b-����p
rĢӃ٦1�yb�a6}b'��Ii�}�d�-��ys���\pz o;l���]�Y�<����(��l l
es����!Z�$�a���K�ԁ�"ȭ@�4h���SH�!�D��}-���a���M�j��!���#(�fQ��b3�U���l�џ��p<�Ѡw��!�^.�`'ĭa�l���e�R�#~T�����i�f�@��f�<�Af\�J�H�&N˓3�Ѫ̡+�ҧ�4��"%�x`EdY,���(�*ek�pC�F�8� ���x��M�����jG6¶t�3����'n�u��'�3�������&7h�������9��t�	�J04��dS�
��`� K��Dx��ۓ%5*u��$�ܗ�X�Z�珼��'�^�B��i�r90c�M0��Ɂ��J�m��<"Ólb��%͎�� +pp"���\0:��oE�q}����Unzɸ�/_��{G�٬t�|�O��Ζ3ٸ��O�aA��mT��y .�+/��b�'>4Ո#�H�µ���� Jx6��'���goW�2|�gB�L�P3�'�b}�牕q�@)�B +��p�'�Mc��90�<�����) v�,��'�NhAmX �����#�����'C�Yp"R:so:,���Ȑ-��Ë�d�<=A
�Q��)��j�����*Ou��b'DD�!�$�C$T�@��#�\���	�jE����F��O?�ɢ��J&��;t^�5��� B�	j~����e�_�*�n͉tR���
Y�5�%ҁ��=Q�+@�).#��ĢH0^�K��o؞�HT��	t�����w��	3����-�D��eZ�T�>"p"O� �a��!^:-����Z4j������c�D�������#}����8C�B�d�Q5�X�+_�<����7{z��[�	ވS0�ZRڃ/�XM�g��?���9j	Q>˓v�{�Ye8�q vƀ(/ELՇȓ"�D���TLI2��m�)t��+��Ժ>�VU�Td�}�a{�iԕE�� �b� �pY�����p=)P��i;��F��M+��Q���vN˶{�BUZ�Kt�<�E �`��H���ǭ�~|BI�[�`:0	��A̮������CpV$�C�I;0E��"b��K!��A�b:��
%F�9�E��%J
(J�)G�q
��?O��|�'�
=S��r"�	Q�V�c��� �'�N=��F����AAA .>
H���T3;l�e@pJ���0>�2AP#9���2f��]c��ۑgT؞� ��1?���Kܼ����>�I�����p�݇ȓ4^��Rb��,oX46j�b��'��iI�l4@٬	��o�W�O��K�� rcB�7c�����'"ZY8D�,� 9�L��a4�SN<IR�ٗE�`:�
OH�����3���%I�2c����r�$ a��u.�PWMU�=ֹC7j˰:�2�H�O��4����	���	D�v����I;N%�XH1�(1�D��Ip�|0 '��:�ZqS�"O��PO�Ol���G+g��%���O�i����;4T-�L�b>!����4�r�S��I5<�J���/��,3�"O��a�炠]xZ��el ����>!�K�.��h�iK�7��H8�KK�i>��%3�@��G��5o�rp��)2�O�d����4r�v��f�v�
("%ぢ[	D��%��ao��P�K �P0�'��>	c���ׂڽ3�<�J���I^�>I�"P�2'���3�o.쑉�ؠB�:٦g�:�\�a�Y��$������d���Z��W��.�r�Tˇ�
�T=`�z%��F ��)��֎t�2�ғu2r,{��42h���m �s�(I�'��}�q�X$z��e��dIxNT��J<�D�>�������*6p$�4�]y�ԟxe���^):w�	��L�C¬����'L|m�ՠ#q�,P�ۧ�����8k:�e02g`|�MZA/�I��S�K�5�1���#��$�>��؅�8��xrF,x��ui����s��}�'���cw吐N����oO -���%d�&aP��,L:��䟬	J4�ɖ�R (?�呇Υ�Z�F���s�c@TH<i��S�{0���!ʃ�ov�Sa��K�'�0`B%���79�f�AAN �C^ֹ�
T��@9�"O.��Q'?X����^��ޔ�R�O8�Ѣd�>���h�����[S8]ju,?:�;�"O�5�AX�g=0t�r쟿R̫g"O�mӱlA�L��d߫Q�����"O�|ѳ�R�8�~ЁG��l�0z�"O��!1�D�ST��" Ë�x#R�#�"O�P��@�L,��c�x��m�"O�@��E�.��5��CR�z�>i�"O@ti���PV� J�dȐK�z�a7"O �BꁾT1rv�؎#ǆ��E"O|]{�/�+t�zTJ�P�oڼu�"O��6E�V�飲 :*����"O6]��	�llm���/3�:	۵"Ot��D�G���|ZRN����r2"O���" /Mo`iC�o�?	�HH��"O��!�J�|�<sD�/��qR�"O\����?W �i��CJ��$�b"O��A�+B*�r�hCBַBH���0"O��ygLz��t�eA�/����c"O����J��d(�ѱ ����Q�"OJtҀ �~*�*B�X40*�p��"O��5�Za�Š���\�H�y0"OD9;0��r��*�)��wvJy�"O�thÂ�B�ܥ�NK3z���"Oڰ���Ȉ9���$�˻%SLt�"O� ,��\���:rb�)%[�a��"O��ш<YD�	�t @�6�e1%"Or!HL[i�����YǶ%�G"O`豲�]�S0����ZF�Ti*q"OVb�D�;haڨ��$�|x:�["O��c5�Ax��y�i�gQ�$2�"O�$E��vi���\�l���
W:�y�P4n��K��FD���	M���'���j���y�V�=�t�8�y�f�z_�����-{�1����y�iف�~D�C¡�r�q ��y�W�tOtm ���	�x���,Ƃ�y��҂'��Y���u���b���yB� (RC��(a�š}+Z�7"�"�y�ȕ�4����B�-��i�ɇ��yb�V*w>X�	#�ɃT�~���ï�y�CK����rN �5{@���ޑ�y�L5l�d	Y7��*��؋VX8�y�,WQ��wm�8�ݪ�՘�y�#�D]˓�G9nڠ0eŨ�y⊄/e��Y��M��%: ��p?��֫�M[ރ�ؚh�R���k�q�P������t�j㟒�n��vJ]<�,wdP6�$0�>1Έ���O񟞝�W��rɪ����P�"| �D���t�x(��
����SA>��3G8a�DcÂ>�4T
��?r�ՉV�L�@	 ��0|
�S�P� ћ�M�7Gf) � �Pa<˓I��� �da��h�� "�WLNP{��S�ʸ'&�������O��	��E��LۗDW�P;����r����˶y��$�����������#J"�q�6���uZD�#ֻT^�9��O谀�g,w����	��T.��P���t�jt�_H�	�"[���) a~�Ş$��C.P�y�l	+%��I����?1�"7ʔ�ZRi�j�)�'��8�0�K`� A��n�z�lڑ'$}ap!!�Ԉ�M�ȟ�<�FD�R-��:���	w�i�Oo�B "��Y.s���`�a���g�S�@��:]x�Ĝ@ѬH����[�<�cZpc���#k�h�H�,\�<�..�q@
�Gt�eH�r�<#�Q)]��2&��>y ��xwL�q�<�D�R�d���D޻Hoȕ��c�<	&�V� f�ًW̏"dW^} Bg�D�<I�JT�9���H�!�8c��=(#@Hf�<�Ed����@�gV|@�+g�<�&�_;Gp�˔䑗7d8Laad^`�<�Q�̳�$�z�i�;+.:Xp�A�<q�ˆ�z��)7hȢ,������d�<�r�C�v�pk��Y�4�<�ӣ�g�<�Q�S�˼@��S���x�/�n�<I5�T�i�Xa���W�R��a	l�<�2�&g�l 8�O�=ޒEh��@�<��$��_��[�&�_�mB%�}�<� *�b����ɉ3]t`�F`�P�<�e��;���:|�p@"�u�<	���LB�l�`�	�3���
ŏu�<��iI*Ϻ%C�ĝ ��ga�o�<�Ȕ���e�v�PNZ���w�<	d.Y�uM�D0���d�@�Js�<��GK�E_(a����ZX"�HÜZ�<��W}�<�,�O��鱡� ]�<�ǫ	Y�Y9��37��Iq�\�< �N� d���'��=[`�rK[�<AP	L({�:��0��7|S\���FZ�<!֣F*n<��H�d��ܹ7��U�<� �QQ6vU�r�ÉS+,J��R�<�u��x�D�`E�� ������f�<���%�uK�l�����c�<�&�g�4�� �kW�1�QF�<� T��a�ŶG���u埽s+0mr�"O�i[g�E�D����S;z�aQ"O88��\D��b��8�0�"OT�:F
�>���ݫN����"O����I7�B@u��$4G���t"O:mS���<�h�A���nO:5�f*OzU1�(
@;�`ۤ�ƽjHг�':dE��l��x>��ƞ�7����'fҖ�i��h���v'�����w�<B@�|u)5;"}�%(��p�<��b�4h% !ڑ'�6$���
u�<���O=���W�Od&h�̘m�<1���?c���FIQ<WH(�CU�MR�<Y��"*F�Dˈ9D�4q��iH�<�P ��)}|��!�,����F�]�<��`d�r��V/D�k�̝z���R�<��)`=]�a���L@}2�BMu�<�塎�5+�i����Y�H8��t�<����8DR*�-k��y3�j�<!D�-��{��\@������Q�<	��=���#j��i�DdѠ�P�<ɧގDun�
�J��g0����%�R�<�b��2��u��M21�Ra[r�Q�<�6���`����C@	+�T �)�b�<I�fCS1���
�<��Y�1�H`�<���@,5W�y ���N�zL ���S�<y�	��"���*�Ǖ�
RmcQ)
S�<���H]�]�`� O�T���j�<	Pg���ѸP�Ғ60aDǟq�<i
;5�)���!<8Hj���m�<qg��K:(I��L�=��Q`�Oi�<Ic�x��FU���t�N�<y���	(�N��U���D�T���#P�<�#!Ciu�x����ơ���T�<��ٜ8�L��E����
(�0�CP�<D,]#oU���ޑ���w[f�<Y�HD�����R
N*��R$��a�<ٗ�W����bԇ+s��I���`�<���X(�]�H���`ΎA�<��S�AJӈ߼�er��@�<��M��\��"�:6�(����WX�<�`f�+P�`�ؑ�����pqo�W�<��ګ�@!��5b|���T�<� l�Ofj�s��٭jh 7�WF�<���ͧ����TMϦw�-t�ZC�<����4z� ����N�^��q!��v�<A����<�$����_�m��X�Ңp�<�Z6.r���͠H���#,�B�<ٴ�^�b��
ֈƲjŖ���"O��0Fe��rʇ▌<�Q�"O6��UI�?������>��)��"Ol�J�ZlY�����8��H �"OZ,�⣀�\�N�(�l�,r�JD"O�D���(Z�p��iU�l��I�"O��RW@�O��c
(F��3�"OD}�C6���*��%dX0D*�"O(]���WU,1�I�R~1��"O�I�����8�2<B�35��y1"Oڭ��@ʄ��Ps��*B!`"O���c�77J���)tbH�b"O�U0�lߴ�*a��a�#�PY��"O��t��6 ��fŚ(:~�Ja"O�e���HN>Y�4둲q8���"Op��b�If�t���DKa����"O� YBЊ>rWz�s!Ç�{DX�E"OD�"j͊'��dPȚ�b�*��v"O�l�����?dN����O'N��"O2e��ŋ,�9���[>'	��"O�{��ŗB>��
�'� �p��d"O�L�a$��4�p&�1%�DE�W"O\4
�mB4���FӖ-E"O��؄�:oA���Ճm��
�"O��cѬ˾4p�%ȋ?9Ȗ���"O�cOA��{(Fx��"g"O����Nݖ)G�t��-�t�F���"O��؇��C��}��P�$8��"ON��0!�"V~�dRDf�%0,�U"O�-"*�0�}3��V#C��j�"OXh�����$�/�buB�"Oz`�E\�u
��"����fX��"O�1���4x�"�Z�8�"OD�@��+o�D����K\�c"O���B'Y@fx�GB'zN���"O������5L��a&旱X����"O�=Z��*��(@$X$��	�"O&=�p�_	eNRa�D��X�R�Ac"OP����>/G�}�0Mǖ2΢�c�"O�y���Lt�h,�$d��)�P"O�x�ɒ"z��8�׭Ё)��I�"Oą"1���J@ 8`�FE��9�6"O�U���9i�ȠB(O���j�"O\�+�L')N��W*K���"Oz��&ٹ���y��۩Q�qH�"O�U��+�(=� Q�3���J�����"Op���U�,Ek��DnE��J�"O��@���h��,̪c��ѣ1"O�H�-�t���!�ԩ
��A�w"O�8����j�����ǉK�B�� "On��C(�?�����P���I�"O.�x��ىl��U#ťN6	�h�"O�,�%��Fh���c��0�U"O��[�-���EfN."g<) �"O�t������q����+��]�<Y1E?C�v�V%��E�xqy���\�<��ؓ=5���]��p�!��M�<��!��\����2� �u� đ.VI�<9I�Y�
�	0��W�Fa�a�}�<1I�+'��1����'/���N�P�<Q�GQ�E�@ҥ���(�8�FI�<A�l<B��yQ�㞳\�,�pgm�F�<� ��L�ʼ�vl_0z���7�k�<ٱ;ў%��Y*kЬ�!"�c�<�6�D�^\ش�����h@� X�<��sHZ�u&� ش�kb��P�<pET�]�(h{��H�iZ�0�M�<Q`��5�MI ˈ}�j׃���yrA�����ё!�l@*7���y���`����%�(|8�TM��y��
�O@�$�$�-v��8�#Ȁ�yR.��J��`d����H>�y"L�΄z�oЧn'XD�@.���y���m�H��F?�"l�@̊�yr!ؐS�i����l���Ó�yr�,.O�Y�B��&�����2�y��C<̬p�`�� �d��`L���y�F=O�|D �,U�nπ��`+�ybj
<
��T�kP����K5�yB�'N܌{�/ht��C�m�y
� �D��ڤg�FZ�%�&y�v�"OT%;&��"+�>�k��]�#����"O�\AE�2 ��@jJ�/�܀�"O|-��"D
M"� �G tz�5�T"O�(SӋ�0�8�8��͂^@��*�"OXPT$� ]älrdA?uA��y5"Or4��S!P`�q�����;��\h�"O� �b�с �Y�7�!czVu""O�{����B��ɂ��/vxH�"O� ���#�ly:�A.�����"Oty�D½Nζ)���0�J$"O|�	'X�x�Ѐ3���5:D`}zS"O���嘭�:ݘF)�+��Q�"OL,��-�,��QJVG����"OR�	�i߷=*fYjg�2Mm���"O
�Ӕ��o\�A�BO0T��v"O��j'��s� ����+U��uy�"O��[T*��@M�M""!��$W"O��ca꛱iKZP�� hq���'"O�uǅ�\R5�T�Ҹ���j�"O"���A$���e�	$�:�0#"O,2@I�7k3���o�4�:��"O�	����1^Qw�b�"O�� �GH
dx�M��o�d��"OvdP�,qb,�kGK'�s�"O M�瘃p=�|S�Gw�1�c"O������k��l҉\��ر""O���¤ЕB���T�b�HE"Of�C�F&)����b�L	'��b0"Ot=���D:'���	G,�<���(�"O�xPC'�� :f�
��޹�p"O��%��?S9�k#��:K��M�"OPp�\���D�eŽ'���p�"O���'Ѝ?u,��bQT[*�"O����V�DF��;��ՉK���$"O�	�Ć8F
�����B�X��"O�4'M�?_%�"�S�g0٠"O��&   ��   �  W  �  �  �)  "5  G@  (K  �V  �a  -m  2t  z}  ��  �  /�  x�  ��  ��  F�  ��  �  M�  ��  �  y�  ��  H�  ��  ��  U�  .�  ��   b 2 Q j% �, ]3 �9 �? �A  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e�!�S�)�Z%����� �Z��I`n!�ͷ�JP)���4�H���,\��Z��(�*�-�pZ��N���V��YQ!򤈧6��r�7Lޘ�զ�]�$�O(L��fÇ�0�˴E>]��(�q"OR��х�=~�6l�F���
ٚ�"Ö��hY)F^L��!I�l�H��'G�����MP��SR&K!J� �L4D��xÊU�l���ᠪ�D�2�ے�2D���J�p=����ސ!�&���#=D��I�b�".ū掛�6�b�kf�r�����d�%��$h&��n˰E+��/�!�d�K�"H�&�%���s�'\q!�DؙX�^,p*��y�V��Şo!��0��(g�̏R�j�y�JA�e?!�D�-Qv��o=u*@�#�\�m>���)��Y9�һ/�����>ސ�a�;D���rfʣv6<X0�ڏZ�z�B͹<���2Z���y��ӂ+X�2������0HX���$��}it�u�$��TAζI�!���!����?@�hLB����2f!��7/���O
�/nZ�:e,L+�!򄎺o�~}��	=\G��aB�!�d��=SdIH!/M�E2ne��@�2�!��
�Aj�dqE���p=na!�b�#Z!�D���pu�$*L@�� #Y!�D��b����#21v �6���?�!��A Q~�y���*"�<����� �!�ʒr�X�Q����0�_�:�!�Ē<_����eb�
1�L� #�ׄ{�!�dTJ�D�٢5�y�ī��!�$�@h����*ZQ�s�ǩ>p!�$Y2:�~���Mf�W*�3_!�d��7VB�7�ݾ�*4��)�K]!�� v��d	�A� X�������"O���!H_!5�*�j���2��PKv"O�D���C�C�~,H�k"H]p�"Oܥ�Fe؋�P$`ū�	*��1"O�xX����J�I$	�"O"�ғ%�tQ�����mt"O~�4FO8P�=��@��l�Z@"O ��҃_	2fD	����������"O>�%*��TD�٘AiN9Hy\Ŋt"O���S��� {��H����"O���!!E�U�E��lΤ��"O�})uaZv�����y��8"O����!?��fO���1�"O����W�8����
���0"O�`A��Ch��#gk�:k���R"OFԑ���l7����CŪa�Pې"OF�I����B/�aZa�R����s�"O���eN@��U;�Mi �;V"O�eσrf�Y��"�	��E"Oȹz�m_�c,�����v���"OL�e�R.��Xa��a��M�s"OصJa��4xa�H1U�uj""OT[�d�ڈy�'�L�е"OZ=�Ҭ�kz�׻8J��#�ŞH�Q�0 �6\0J�{��݁gC剷!���;0mH�P��9�T�v�C��.nڨ)�K�'6��	B��ހp��C�ɳRox��ᐝL4�)���[pO�B�I�JK&a�[q�8�h��U�C�B�ɘY�$��o���=�����Pi�C䉢t��Е�]Gv��G��&w�C�I�P�\�cG�<'"���Q��
%�`B䉥9M$ Cb���}��D��^�%�$B䉪s�y�1
Ǫz$�aE�δ�B�I!�lP8�(
2~�e�&!�'gNB�q�>�@�@�:��������-��C�I9;)�Lq6�&( �4����9`�B�ɳ>������"^��(sLA��C�ɍl(�MyG�AA��"� �,®C�	
�8�ka[2la0�0PA�C�	q仂��;�J��E�A(�4B�Im�v���(���9)��ս-5hC�	-`��j����P$O�w���7"OB�:m�n�
7m�E�~�V"OVcv��+��
s�U�/��� "O�[mS=$6N��Ӏy����"O4HI�_4��i���Z�5�"OB5	�D<Y�~�+1bP)'P�y��"O��;�@�g�I���2c4~�p�"O؅�%i�_ΰe&�Kw���"O���� �f ���e�4�h �"O��2�ݼvW��bqEF^�>U"q"O�� *��q������uF"���"O�ay�Ӓ%�z]���ָ<@�0�b"OdE�*�q��5�.��A����"O^�r�JT��Dؘ�F
s���"O$��̩U5�p���`ihm�&"ON���ǅ�gV�1�C�E�8�2��`"OH��e��?���Zf�� _�p0�"Ov����->Jq�&,|��{�"O~��h~>}�&f��?���J�"O�I��\�"z�%����0����"O�������|�&��d1�A"O���F�`K��S��u�ٻ"O� �`�@dO�n���sȬX�ԥ)�"O���Ejɩ�9�@̇�*�(��""O��ZLƜg3x4a$�.*�Di2"OFu��Ü0�����k�h����"OHq�q!2�� 	q��K�V�[b�'���'��'a�'�R�'���'�������$e�� r����"R�'D��'|��'"�'s�'���'J�8
I��H�Q������P&�'���'R��'���'���'���'��Y�mֽN^zE�!n[IL��Y��'���'�B�'���'HB�'F"�'�����ث�ByT�]q��P�'1"�'�R�'�B�'�2�'Z��'?�a��m�&9H���"b�*��V�'��'���'"�'���'���'ʈCV
S!� ղ��F3��e�1�'�B�'Z��'��'�R�'���'���r�K] ~oxH�������E�'�"�'pb�'�R�'y��'���'���9%�#I=��R�&U�\��T�'��'���'��'���'���'�h�`Ŏ*=[IҴ<'�F\h��'Ob�'0R�'���'M��'�R�'A.�R
�-nt�ٱJGy��Q�'���'���'���'%��'s��'��e;�`���^����]�(9��'�'���'OR�'���'"�'Xh�^�E�h�#	�9y����'��'�R�'x��'R�"uӀ���O�̂�h3��J��
'|��X��Iy��'*�)�3?�0�i�(�[��&r�J��0']�M�L��,���	��Y�?��<���UNu���l�h6�Q�*#tq���?at�I��M��OT��zL?-R��� 9��A��M�����=�IΟ��'��>���p	�0�&E�<6�0��ƚ�M����P���O,7=�ʤ2Ё6'x��qf�B��|�G��O��$e��ԧ�O
�i0�Dحf���k`l�![��L�v� P��m���k��=ͧ�?���Őv�(����~A���r���<a/O��O��lZ;H��c��z0k�r�vI�Y�����m��Fy�	��	�<٫O@���5T}�Ec�I1R���񂑟T��3�Pe��9擳��Y�88bkgY�53 �����*F��Cy�\���)��<�K�:���7�]:l��*$HB�<���io��b�O��nD��|����	���O#
��P�����<���?	��Mq2}0�4���a>us��l�X�3�Ϻ:7�"��N9|��sī5��<�'�?����?y��?᧤iV�e�
Ӵ�b��eª��D�����. ����I��$?��	�0V�C���qB��l��la4*Z}��'TB�|��TF��N�9�⮄�y~�� ��>h�@(�i��I�T���!3�OޓO�����ƅ4)��Y8T��.M����?���?���|j/O�oZӤ��I�Y>��`��L7z�Np9%�\ڨ��	��M�N>����	ϟ@�i��;����@�V�5 �s��8aw���F�m�~]*��!����O��a�nB�@ڝ{{����d���y�')B�'h2�'!r��"{�H@b �_�`��c^.kָ��?I��i[p��O%�#z��O�z0]K� ���N�W!P1�D1���O��4�|��i�<�G��L�ǌ��u����ǧqR�M0qLӌv��X�����4���D�O��I�K&�٤a�s���Bz����O<�:���%/�	ן8�Oz��;S�)�B�ăŏs�����O0��'���'yɧ�I@m��ҁkY�vZ襸B��Qx��q� ��7�1?�'cn�I}��@���)�?$��e�^1���I�t��柈�)��iy�b�2�x�)��~�~a�F�F0Jh��#�(�����O  oK����Iğt����I�l����1�Zt��C��<�ɍ-�mZ~~�D2 ���}
���!Z�L!b�3� A؆���<�-O����O,��Of�$�O˧"Լ�[%I�87����� >P��C�i� �(2�'���'I�O���b��n�f���6"شw��Z�_3u�V���O��O1��P4m|���1k�"�Jʻ J�<S�i��� R�����'@��%�엧�T�'j֝ST,�\K�3r��U�� ��'���'�\����4%�X1��?�&>�<���ZJ0%��"U*�$�h��@�>	���?�N>�Rm�-�=�cHń(�5�˃~~2��	���1�i.1����'Y�;�0�-�y��s�+��xr�'���'��џ$贩K�)%\��E��B2���l@��|۴b��4z+OhPnW�Ӽ��hJ�d+.DC�M��>9�"/Q�<I��?���[䬉�ٴ��䃽oN��k�O,��rd���s!�q D�|]���ٟ��I��8�Iٟ���]����H�xlL@fg�hy�Dd��Xzr�OJ���O���H�Ď5�i��!)z����Ã�]��<�'q��'�ɧ�O���PiE=^�4�@���<̐�;�T5U�����4CF�ĽP���7�$�<)Á	&�Ѓ��f��I�q͝'�?����?���?�'��U��������и���/�^��R���{�.�͟<
ش��'���?A��?t��=)bxA'!q�6���GW7f��Y��4���G�������O�� L�cY�e�T���D�'{аQ %<O��d�O��$�Ov�d�On�?�p�A��*���$k B��̕ݟ(�I���2�45�Χ�?馼i��'Z���e���'�D���"�*4H ���|��'(�O��r��i��i����ש F���fT	�N(Z�`\x��i�#I>�*OJ���O��D�O,�2vIV����Ү�n�	���O�d�<�%�i����X���b��$��3萴���*veZ�pW�����@f}R�'��O��1Me��	��9S���j�����4%�"�^	3`�~y�Oe���ɔo��'%���eh�5����j��U���'���'�����O��	��M;�JM�<~n�i鏐0���ф�F�!&\P���?�"�i��O�l�'���`�z�S��фH`����,l"�'��H�#�i�iݭR���?I�P���a@�_+Hݡ�J�26��Ų�g� �'���'�b�';R�'��(��(�LB,,�e��ݲ6SvLbشF� M�-O��d4�i�O�mz�uZ1���|�d�ѱZ~�ɐB�Y��x�	^�)� v�rUl�<�R
U�;|��׌�2;�a�cI[�<�C ¯���I]�I~y�OF2J�t��Ų�I;O�<��Ue���'���'��	#�M�E��'�?���?I�&�m�j 
c��!Mm4��5��/��'�Tꓽ?	��� ń()0�Q� �]r��	~���' H�T�0-�ի��������'���WNO�#B�z7#�*.��g�'�R�'b�'��>����T*�� �*Rv��v&��O�.i��'�M���#�?��5���4� �y��[�W�$�f��S���r9O<�$�O����R7-+?�lR�2����D#a`Դ���S{�.�X�G�:h��1N>q+O�)�Ov���O:�d�O�$���2��:���n�΅2�	�<Y��i����&^�l�IW��Ɵ$��G�xIt�"R�AG!�q*��-����O���3�󉅄Q��c�{���Jg��6n�Hp$hj�~\�'���p�e�b?�H>�*O��*nìI%V��Hj��Xv��O��d�O<���O�ɠ<y�iZ�3�'ƅ�sń�;��(�[6,g��#�'f^6M?����$�O���O��Ƀ-h����*�!���#g�&;�j6�-?9#(��@'��I;���߱e��I��a�����Bax��x����۟�����l�	˟�R�f�aQaU�/P.)� �H��?!��?A�ib|���O'�c�ܒO�S�Ą�تOۉ\a�MEL8�D�O@�4�l%c�nd�J�`��$�
K�a��L !A;8S̍�F���IZ�Iby��'K��'����a�T�r�f�o�Jh;D�
7ur��'6�I-�Mӵ���?����?,���`��3&� c/�%3mz�a%���	�Oz���O^�O��?�6����BM(�f)^V�Cakf 8�!t�@y�O*���IhK�'�ny㖈V1r��eڅbT8v�-���'�R�'��O8�	��M�e��b���0�A)@>H#DQ�N�:��?鐴ij�O@ �'��FU�1|�!�4C�GI�t�W�F�>���'YL8�t�i%���a:�S�O��1��%��Vpr��5�~h̓��$�O����O���O���|jRcT��j0X��X�J�Ɓ�*�>��임r�'�B�I���=)�j�C�ˀ�cΦ-�F�v�\���� $�b>����ͦ��Fa���垪>��)�c�P�~,�M_n�B�j���'���'�r�'9fq���W�ll����"�MSE�'���'��V�D��4GQ
�
���?��+F�;�.�L�2]a�ރ�hl��BB�>9���?YI>TcǺU�rpґ��7��,���TV~�#<P��au�i�1�r��'��
�3^~\hdM�T'��3�,
J��'���'�b���@�BM���)�-6W2<9Kw����411�A���?i��i6�O��C9�X)r� ��.3���R�yB�'���'V�aSe�i����?�:����O�d,p�׺eq��Wt��9��B�	Vy�O��'
��'Y"��)`h�Z�%Z\�\%�&��<��ɚ�M���?	���?�J~�-��HQ!��/u�l��������9�[����̟�$�b>UK��Ϲ3�M����RPi�FI�ToD~R��%0�����$�^LT��=���Z�"\}�d���O����Of�4�b�?�r�[>�?��+و)�|�"�OS1.�ȸ�k;�?c�i�O���'<r�'V�,��� �C�^��L"1OD�la<�Y��i���<�qàԟ������G�V�f�Yu�Ӱv�p�H����V��D�O���O��$�OJ�4��
\�������#�����@���������?���`>���!�M{J>9�� 	}��˧Ȝ5	��A��B����?	��|�����M�OLũ1`3?T�G�N���}���#8���'=�'�	ϟ@�������=!ة�GH�o�*Ѻ���v�����ß��'��7-O�2����Or��|*�Ȉ,��G!H97�2��'gn~⭣>����?�J>�O"�D���L�!�~�Z�e�o;����O:��0���i>�(�'��q%���w�%"�`4�Cm�5M�� v�Q�0��ߟ���ߟb>��'��7-B3������_�z�B͂0�<Qn�	�*�O��$��a�?a5[���	#�r qS'�:<�ؚ���П�#��F��a�u�S"���Ay
� EC�L�v�B�x�8Pպ�K�6O���?���?a��?���F�	M����R2�,��a] �
�o3L��֟���L�֟X����s�iK�H��&�11�,8�HA:�?����ŞZ���ڴ�yr�߷D��A$U5b��x�1�y"N�TPE�����$�O��d5M�̜3��-�T\����P��$�ON���O�כvO�Ua��'2*��m��L�dPI��A�k�T��'�I�>9���?N>Ivg�#���bAC�=�$�)��P~�$�H�����J��O����J���$-���bR�KZ��`���y/�o4~e�F�s:�J���1�"�q�`0���OR����?�;P.���9�F�Af�<I��̓�?���?����M��O�<C���1:��P畗a����`���B���I>�(O��O��$�O~���O� ��k��:pb�q�#�=⺬�֣�<�i�j���'z��';�OyR�Eݦ��a��0����!B�H���?�����S�'��)�AҗJS
�qD���-����a�L0-�.O��p��?���2�d�<�K�b<���g
ې���! <�?����?����?�'��D���E� ^ޟ�S%�L�_�������>~��
�\��\�ݴ��'�~듍?�*O�y#�J� ���Ə�-$��z�ů��6�)?�'+�3~�����&����+�"5�D�`��7Cˠ1`2B�<Y��?���?����?y��tOF�p0@� i&�|bq�]�l�R�'u"hӶ,��=���dæ]$����E
)*��ùVp@��X[���@�i>��6��-�'d�����D���k�"|oZ]�ץ�3%"����䓑�4�V���O��$�Pi@a�aЦi��{�Z`*����O|˓sy�&
�?4���'�2�O*�4k�s�\��4eW>qa6m�O�y��'Mr��?������|���Q
��p��$S�М�1��Ȳ0��g�~����ܴ��$��Q��':�'�$թ$a�6c�5Z�N�/����'�D7�@"��T���^Cd�!�/�1�ځtu�ɠ�M����>q����cl�3:��P�4���7�Q����?I�È4�M�O���?���V���b�20�,T�b�݊V�x�(�'R"�'#��'�R�'��S��v��C%ߘ+vޑoAռ�r��4@����?�����'�?qƲ�yG��K�@k C-T)xE�V�Y�b�':ɧ�OE\}I��ig�����90��A9�rq���6��d�4O�{�'%�' �i>��I<���:�	!�(� ௝�aن�����H��ߟ��'�.6MR+A���d�OT�D��Dw���R�	]�"xQ�lɶ^�Z�ؑ�O����O&�O<g��(`A@�-IT���0Ý�Ȃ gې|t͘��u��}b��R���8�(!�`�Z(� ���T�IƟ��I˟�F��'��ÄW	#p��;c �yi�|7�'t7�#qf�D�O
�oZ_�Ӽ� ��(T�~�QE'1���L��<A���dX��6�.?�QlJ?M�~�)�(h.JQ���7�|���j8J���L>�+O0���Oh���OL��OR��ӥ���ִ��k��4�z�,�<�ҵiè�0�Q���	Z��hh�̋�@X��ؔ��X$\=� @���O���9���%X(�����A��!"���,�f�P�}����'��`�D�k?�M>9-Oܴ��#��Y���Ճ�5+wVp��	�O����O���O��<�v�i(�M��''��r�LZG>Ҹ�q@�((I���D�'��7�'��1����O�˓Q�rg�V-JE����qs�¦���M�O�ͩr�Ĕ��U�;�i��^���n�ʜ:l�TIt\=O��d�O����O4���O��?���C�%q���:���@s0�����T�I�T�ݴ<����O��6�+���R�����;����h����Ox�d�O�I�(^�7�-?�����( l��r��u��j��6�	�?�A.���<����?a���?�ꛒ[٫s���gI�<��1�?�����æ�HhIȟ��	���Oǲi���-�d����I�����O��'Dr�'�ɧ��ԜD�@��٥FpxrE�/^AL�9E�'�mZp~�O�:M���{�� �@Ѡ[��2�h�'�܍��?��?Q�Ş������	7���$U�1 ���Vh^,��)�j��Iß$(ݴ��'4X듣?��8Q���XI�>y�AP�9�x�L��Q�޴��d��$�$�[�'5�˓,�J�
ub�!�桁�EWJ��M���$�O����O����O��d�|�&��ex7	�.T�%@0%�
u�f�[`���'����'5�6=�,��KM�y����@m@��L"!��O�b>�Q�]ӦYΓwZ~Q�	[� ���A�d"@�̓`��E��OdL>�-O���ONXTLR�����b̘�ft�(`p��O���O,�$�<��i@B|8&�'+�'�́����p$xEE �!D.�2��$�G}��'kb�|�o�q%�5�A�=y�hq�B�����D��V�z�ˤ�M?$f��T���!���O7>��0¢�:���`D�|����Oz�d�O�D'ڧ�?�^��!LU�(��D���F(�����	��CHv2�'��6M"�i�a��&�r4��S�m�)
��d3�
{�8��Ly��VU�V����0h�4"���&$� $���GY'~l�E2eݸR�*�r0o;�$�<����?a��?	���?!C�˘|��z��E�yV��9���⦹A��[�D������*�J�	`�b=Ah #�tkE�=�����Ii�)�s��+�!��=ʗ����A���q�'qR$��'�n?�I>�+ODI*E-+��$��-S�#�nшG�'�J7�k�N�$�M�Z  pe����	�R��&��C¦��?	P� �	ßl���#�&isQ$Z6<Z�BS��e0�ȁ����'��c�j�I~���{% �Z�	I+I`���#_:���?���?9��?Q����O-��U ��]�~$F��i�<	a�R���I�M�3�L�|2�K6�V�|��L�r܉`P�چ�D��ė5J[�'�����d\��V��`1ӦܞsQ�phFjʨr�t$�Ɩ*&�1W�OԓO�ʓ�?����?��8��@��a��O�R��T��&��(����?�.OZ�nZ�n,������@�	E��.��.7|����C�:e��	L��dDJ}��'k2�|ʟ�	G-�'`�b��l�\��}ʒ)� XԘ=�ǎ�:�i>esV�'2*�&����?}�����I�Q�ԎO������ßb>i�'�6MT�\^`J� 
�n��Y�G�5XU<�;�E�O��D�Ӧ�?�cT�x��%Y�0����Xs� 1D��|�r\���(������A�'�z@�"\ܧ>`��SC�=�X��F�I��|̓��$�O`�$�O����O��İ|b��� 洒C�L���U*�~���c�Vpb�'�b��t�'�X7=���XV/K�phƍ�$i� i�x#��O2��<��	��itl6�h��
Ub@TD�d�W(R	jf�+�p��@EA�{��f�~�Isy�O���	�iM���&��D3��kP#$���'FB�'����MS���?����y�J,9����L�5k�Bm�1�?��X�H�	͟x'� xA
��+�>����rs�!?)�M��8�`��4�O|L���?�1�X7 �2HH�B�B����N��?����?������ϟ|�
Z+R�lm�&��w:�Ej!���T�ܴQԤ���?��i��O�n�/e��,!3��#v�T��J[�3��D�O����OB=J�Jg�R�+�rFJ쟀��R��](j	Y��s@hQ
׷�䓙�4� ��O���O��$Y%涔+ ��


@ɀE���%^����4 �bH���?����'�?Y���/��s��	b6�����[#��۟�?�|���׺1R�"T�Z�G��$���=:ʨm�!����$/?�� ���ys
�O�ʓ+t�U�E'�&DX�x]R*��X���?Y���?���|",ODEl�1:�xH�I�n��2&�Y6'�~ex�ㄍC �X�I��M���ʸ>���?��6}*��Ɵ	����r!ÅaR	9Í5�M[�O<�I'��������4�w���D���v��e.�Qä���'���'���'���'����PG�X'�6��%㌃��D�ゼ<��)>�v���t�'&�6�*���.#�(p�V�ͬ�i��B�1O,���<Y�C߄�M��O���1�Śe�:x�f���s|ҧ�iL�q��hF��ON��?���?���>u��d�E/M�b�zg��mG��S���?Y.O��m�(	�N�����It��	։u�,��SEY�3B`őӠ�����p}��'�|ʟ��b���/5���A!��J��d�W��/A�M��qӀ��|�&��� &�|��gL�#P �r�U�{%΅��@Fԟ�������ӟb>]�'.�6�W�y�V�12'K�\�Ɓ�Q�aN�����O��Xʦ=&�l��;����O�=P��`�������`�+�Y%�?���?��`H۴����6�&⟖��/O^a '��B�b�EJ�_�ܡ>Ox˓�?q��?���?�����P�@lh	1A DO����aP�n�nUl�$�'�r��t�'�87=�`$pg��_ ysR�6X,4Y��O��D2�����7�b��$�X25 �p��H�H�2 %�v� �Q(��)���<a��?qb
��x�L5�kT&P�hcM��?Q���?����d���U�5S����Ɵ�@�,������g�0P��lNX��t3��̟��	q�	p (�y���0|-�PC��	�n�`��10�G�h�|� a�O�h���vd���u��f��e��Βc�t1�ȓs�Z��m��4\��jV�:�P�K��J��VD��'�^7-2�i��h-!Ѫ5�II��ɓ�w���I�<��(a��1mZc~Zw^�����O۲Ӆ!�:W�>u�jI*5trYA!(Ic�	jy��'���'��'��E�9�����NF	w���E�
3�I7�M���_����OΓ�����57��hv���DN���ʄ*`<�'o��'.ɧ�Oj�Q�N�0����f�ܥ(P��R_|��V��D!cM�|��6�D�<�BAQ�:(p�nL'q�ޜ���?)��?��?�'��$����C��՟	�mI�+��������j�F]џ�aش��'M
��?Y���?9f�qt��ŧ$w Q*W>{��)۴��dD�t�&�1�'��O���N��l��ʈ!sB�5*ƨ��y��'���'��'�"�i���FEz���L���S�*@(n����O8��Z�0�m>���
�M�N>��۷g�4u���\�|�v9�ri��䓼?���|څ���M��O.x��� ��E�lY�m*����+a$��ˏ�~�|�W������	۟���`�
��<XAn#D`��������	Hybn���A�	�OH�$�O�˧\ �e�Æ6]fy��+^:욙�'Q���?����S��N�R�6�RF�ՔP�.t�!��+K�4�+E��o�Ze��[��Ӏ>p2�|�Ƀ)�4�H0y�$�I�"�);T� ���8�Iߟ��)�Iy�cl��ͣ��]�'�)�QN,� �{�F��Z*��d�O(�nZe��T�����Ա�� ���h2M�=~%F���Omyb��N��v������'��bMy�ύ
?;`AÂ��8`5�Q �Ʌ��y�S���I韬�������$�O����H�%�x��_';h�B(zӀ�[���O���Ol����Jߦ�]�	�8Q����3�������a�Z��	��@$�b>=���J���ϓAߐ}J�)ӄ7rm�vH�'2s�ϓ5��M�Á�O@|*K>�+O�I�OJX(�FZ��x�4�&	v@�����O���O��$�<Ҳi�>y�U���� #���W�L�G�͛�O��T�T%�?1Z���I{�4��Y0ȑ:A�^h"C�S�&�*��'��e�D�F
v-�AR����˟TR��'�ؔ��G>Hzd��+�7���0��'���'��'��>q�I,B���EE�b`BAp�@�s˒�����M��
��?�F��F�4���O l]�|�#Ȑ�j���b;O��$�O��אo�B7�%?y�-\?d��IϾ{\���w��"{���q�"�$K���O>Y+O��O��D�Ov���ONUZ�O�:74�kG�P�%�D���&�<Y�i���t�'�"�'�O���<lvb����|�r!*EX�*u�듈?y���Ş*���zP�G����S�$���9�jU��M+&W� �E��-W��d'�d�<9p�Z�q�.lk�N�>E�r�81JP��?����?!���?ͧ����M�W����d���	�������8HÆ�{��ٴ��'xf��?)���?q�	�)V��
�	����hx��Y�p��z޴��ĕG�4}b�O)�O�%(Vg��xv�·Z�h=(��^'�yb�'���'���'4��	�N��¢䏿E���p��7E�6��O��D������r>	����MsO>���N�p��"7O��ܓ2d����?���|r�� 3�MC�Ob�[B`ҁ<����č;��4��@ȝr>���KAޒO8��|����?���-��{#!�6�D�񡂽u������?A(O�n�%��ß��I{��!�ek�|��\044E"w�'���{}r�'��O��D\~�p*F"+d���L�4��=@��G5�T����cy�O�LH�	B��'�Y	6��y�f��Db]�7��Q6�'�b�'\2���4�'%�dsCV���ݴ3^� f�F!F�\S���N{������?��'��V�'�I㟰��O~���yr)	S���b�R��������O�ёf�j����R���b+?I`��06$D�ZAK��QGx�'[�<q+OD���O����O��$�O.˧��}{uoћD��@C5*F!3��" �iW�ms��'���'1�O��Gg�󎑦r:���Oߖ��Ysf_q�X��O��O1��pJƄs�*�I,���lZ1�21�Ah^�0�x�Il��1��'���$�$���Ɇ�u!�D���`���Ss�J�/�axb$|�> 2w(�<��
�"���%�E;(��`3[\nŒ����>����?�I>Q�#��&��QQF/��C�~��n_e~��^(a[&�ճiA���H�'�R�Z��.����[���4��y�������[E���;��T
WBmvӀMI�H�O�����M�?������ W?��1��kl�	����ܟ�����⦩�uG��l���OUM��A�����1n�1#�q%�Ĕ']џ|���iS� BWk	�
k&���/?���i��0��V� ��a�'�<ySaH31;p�DК�p��[����ߟ�$�b>e��a��B�r��=y��Q�k���.�nZ=��䎺s���'o�'��I �ȩ"uA�h�,�0��.E6���Dʦ�# �Oş��l�s�Z�!2�ɂKS~43+����y�4��'Z���?i��?y�ˌsg��^9�P��U�j-�M��Of��Wo׮�:p�:�I���q���v�``
$(�9�>O�����kBͰ�e�:�>�Q��w��˓�?A�ie!�Ο��m�K�I,K�V4 aĝ�H�±h��;Z�F�&������Ӌ(عlZM~��^<1��i!ġ:c8�����KN>!������*�I�z;N)��U��R��v?�#<y½i���1��'-��'y��*G:�Li�M(~��tgκ\��N���ڟ��IT�)�� �mr�O^�`q�����ٽM H`�a�I�Q��J,O�	5�?�W8�$�+QZ\&��/�(;�Z��!��禥83�D=� ͓S��|D��K��H`�'.6�2����$�O0M�c��}�����?��)���O�����7*?y`�	z���iyIͦX���$��9k�M�s)W	�y2[�����<tS���&�567�0	� |�x	�޴.\���.O��>�S��M�;t'j}#�Y�`UД)���!2X�B��?N>�|:�8�M㛧� �s��Q=ˈ���"��dߖ���7O�ӳ�Z��~"�|]��	ßt�c� 4�|!�Gf�?E6������͟�������Fyk�T��#�O8�d�O��Pd� �hp� �Ap��s��;�ɘ����O��D �d���}bd�`�Y�CF	(s���)�2�
�Φm�M~�L����	3�]���R�Ď^�([�(�I�� ������y�O��o��E찰���t",�ӱM��'�"��O�%Hw�'�rLw�j�杫p��{��P�����ȏ0c��	џ4����c�,���)�'�((�c��YZ0��Y�p�І 5 �0�	�m�䓢�d�O��$�O�D�O
���>~q�a0	�/h�@� 5g�&=�˓d����!9�����'?Y�ɭ=t���ɓ�$ 8SA��_��(��O���O�O1����ҤE�T�����#b	%_c�7-�Ly��CX*������DB&,z���rjOdw�����9eP��$�O����O��4�f�ƛ'��(���5�a���+-�V4�#����p�r�4k�OP�D�O�Ǩ?�v<C���L��Jf�ִ%���	iӲ�ZӖ�@
�5�N~��;|M��YVܒP/�a�X	���?y��?���?!����Or� ȱDQ��$sA�զM��g�'Ib�'�<7��_��	�O�mnZi�IN�\�"�[�*�>�벎�CO�\%������擵ya�n�r~Zw�\aӦ�B'N*Dղs�ªĶ]h1f2l�B�	sy��'���'���WD�����`�p �1����s�'#��M�E��?	���?�)��){���=I��Uq�K��\x4R!?OJ��W}��'Fr�|ʟ�<!ԃ�.��"iڑ%��8t��o=�pk�J��+F6��|��M�O��N>�Cm�4H>h�BT�@s~�@ש�?1���?���?�|�.O��o�BB��W�K:�<ܸ1��j`x�RR�ڟ��I�M[L>ͧ7���:��@d��XF�q|�ɂ����� �I��8l�D~�(	9/�A�'��&��E�jl6�Il����;�̭DD�Y@��>՞] �	�)U�,��G�~DF��o� 
զp{��!
U2�y�(�6� �:e��%��R���ԁ�p�'�p=Q��Փx�hԹ��H6�Q)�Gͪ-�z�)D�%&�Q)$��$S�|z�.єl�8t�#�ԅ�.G���ґ:��	�*M�W��00 ؆8����b�G�Z��t�eh		������3btI4(H�C�����߈$�!��B�d2B�� ��H�AC	>�x`��$
(��l�ܟx�I�<�����d�<�d�&=S����A��(B�2/,�fM��VҖ|����O�L�����p#���oE10.�@��ܦQ��ҟ�̓K����O���?��'׮���ޯ6��s6���%����}2�Ak��'�R�'���;\:���N�va{��^6�k�p2sAn}P���IX�i����ʆ �p�2�V$|;��еb�>q���?A+O\��O��$�<��ҜJ;v�9��	�H��}H��8]���S�P�';�|��':�L)l�x���M�R�01bt���*,�e�'���ɟ��I�$�'�䐣�b>1�J�rh��M�d8N	GI`�J˓�?�H>��?�Q�S0�?��b��d��h'$��<B�i�hN3��I������\�'mL�)�~��d��e�R�0=@��@dڽ7�Bt�i""�|��'#�
�qO�"g��s$B��T�2�PB�i�R�'i�>]�1(�����l����1�84��!O*.+T�(BAP'�.$������ɄaXş�$�P�'D�ea0�>F:��`1,Z$y� �o�py�d�a!$7-�O���{��)]d}Zc `�C�o	G��h��hJ�u�n���4�?I�$�%Dx����I"��FϚ�&y�,�6��ߴN���p�ir�'-�T>�|y�!��M�����vMݡP/x19c�i;��Q��1��՟Xz�
4���s5�C$�̉4֋�Mk��?�'���:�\�ԗ'�B�O�A��[�`An��F�h(�4����č2�d�O��$�O:�d,%�������H��r��}+&inZ�<-��C�O,˓�?yN>��<��e��H��8p�L
:XR�U�'��y*�|r��5�4�?�*O� ��O�-P����<YNH�R�^�V�İ$���ퟄ%���u7f^�p�>��ΔlJ6��T��M�����O����O��v6F�j�5�t9��+e�T��׬cs��{U�,���'�(���4�'�qɑǛ�:] �b��D��n&��O���?i�A\�����O�x�E*�1*��<���9p:���mΦ��?����Ɔ�'�ű��q�^h�F�.	l�ٴ�?�����D�1�2�$>����?ט�C�&��qc�4!êai�* 8O�˓�?a����<��S�QأJ��;���Zsᘢ��t�'�r���� x@B�'�r�O��i�Y������BY��Vv�숚�lg�T���<ᐨs���'*�`���mҾX�<�8�J�P�im�(�����4�?Y��?��'n����$�]
0*�YE+�DxUAħ�X��6-�O4�$�O��O�3?ɐgӱP�dQ��@�.�����o����v�'Mb�'�yBR����	�Z�#O�/��T�1)	�lD����dWl��?i�']��{U���zu6Hr��B�t��ܴ�?�禇���dg����߫y�-ƕ[��� �: i�u'���w�;����@�'���+� �p�26 ,�S��֎|�$]�d�B����O���;����x�������Iʞ@���x�"O�|�%n�
.��?Y��?�*OҀ30���|��F]$cJFf�W�*T�A-H}r�'b�|bZ������o��a�z
s���@鱮9�'�P���I}/"Y�O
"n'[6���	�gDB�R�I�"\,6�.��şؕ'��<�N<Ӭ��Ur"��U�W��r�h�æ%��ky��'O*�`F_>���͟��s��9fo�0l�Ɖ����voT�O?�D�O�ʓ�x�DxZw���q��ְk�f ��Hז'�l
ߴ��D
�9�(1mڷ��)�O���S~2���BaF�17`�"!G��%���4���O��$�~�Sm�s�<,�!�΋K�䑙 �K���`�i.!z!cӮ���O���'��1�`��w��&aN c��^���4�?����?1H>����	�wI�P�"�(M���VE"���lӟL�����z���}yʟ��'Z��ւH8q�
�Y2�R��VJ2!�O�B�'U����:0�ԃDDL)��C��6M�O(�b�^V�i>Q��}�I;�����!~�W�7L76abs@;���O4��?��?�(O*y���!)�������m� r�����e+���O��+��<��=[��	��h���'�\�I7��oʟl&����\y"�'$l��ԟ����
Z}e�$�αaA@��i���'��O����<�aU�ɛG@W<&Ĉ�(�� (!��P�B�>���?���򄑑:Dl�O$R@W�,�, �a$S�0�o��5�6m�O�ʓ�?��?�ŮN�<�/��YH�N	� 3hq�p)kL�����٦i������'���X'j�~����?i�'-��a@lX2?Ǣ�gi�'5|
mz0V��������I%�$���?Ѹ���!~���G�P� ��!Q!e�˓j �5�iV"�'��O@��Ӻ��-E�
܂*E�U~r]Qi�¦��	П$�W�m���Jy����3$�pg��Eb`YSdO��f���D*6��O����O|���E}�V�|!!��,���t��v!҂����M+5F�<���?����O��C�5�\93#��vǌ�;�#� [��6��Op���O,��r�J[}S���	Q?A����A���FO�%s��Ѧ%&��pe��'�?����?idAM�;����"R��3�/ٛf�'��Ją�>�)O���<���kn�	};� �P�]&n�ց���TK}2���y�^���럈�	zy2�*ˤ���$J:�����ݦ:���K1#�>Y/Od��<Q��?��(�M���J�k0v-�̘G��Ap ��<�.O����Op��<y�iVs��� �]�PQ��� Y�l��,R���S���Iiy��'��'�h��'9���K�.C<`�CH��O@ v�>����?)���d�fy�d�O�KG:h��)���YƬ q��'�7�O���?����?16hT�<)H��P�c���v�z�
;8?:���z�D���O�˓T�,��V?a��ϟL��5����,�'O�z͟�A�&�a�O���ON��
�`��|����D�{f*�)3&�+���A�Ms)OjT���V��M��ɟ��I�?9�O������9�F�������(��'�囘�yb�|"�I�5n���J��@1.��e�hX�(Y��JåZ��6�O*��O
�	B[}�Y��Ô"�{����M�z���a�Mc��<yN>I����'@<����W�<���L�
�x��n�`���O��DD�:�"��'��П��s�/��$j��GD���'c剫.b$��|b���?i�A�"e�a�n>hI双(Z3"ٓu�i6B-Q�����O�ʓ�?��"Y8�q��$��,�&Kj���'j��'���'�"�'Y�^�Ps7�P2J|4��1P"�rd��Cٿ9�Ÿ�O���?)O���O>�$S�3��d" ���m��(�*�*�>aɲ�� �	����Iӟ��'�h0tgk>a#v)\.˺e ���� �f�����,O��<���?A�"t�ϓN���4ŕ�4�D�i@
��'Ø�QD�i��'5��'��I�)���;���DӔ=���%���J��ЮN��n��ؗ'���'�b�8���M��9NUز�2�ʩ�2���%���D�'�B(x��~���?��'0t�Xy�F� W��˷)Q�|�V�´X� �	����I�6���IQ��'��)�.`����և0��a���v��vS�#�(���M���?����R�X�֝�{��Y���� g�ڠ� ː1r�6m�Ov�dK/o��dNU��'�q����5��%Hu&,�@�؇
MBXE�i�����n�L���OT�d��r��'剠y�hI@O��Gr���q����Hݴ-;(��'N�IV���?A������D 6�A!"�8�֮:��f�'��'�$����2��Ob����0�5&\�5ޕ���!rdeҒ/k�ΒO<�r_V�ϟ��ꟈ	��Ǜyt��)��I���F��M[�ӂh.m��'n"�'�ɧ5F"�:,ބ��׮.\B�y�a�����^��D�<q��?Q����dӉi�܉c�\�R8FT���K�u'�X�U�BH�֟T��A��֟P����ʨE(;:���(a�'O�Xi����J�柼�	ܟ��'�½j%�b>ݳ��ާ;\{��C�Z�x�0��>���?�O>����?	����<ap�åy'r=�g%�W��&�;pV�	����I����'�R��w� �I�I�? ���g�<o��B`���y�&�i���|��'���Y�y�>�"I�	|�M	O���Q�R�Ц��I���'
~P���#�I�O��I�����RnA+ML ��`�F8��A$�D�I͟�@��ޟ $����R�	Yd`>$�8��
ڜL)�,l�vy"�Px�6�B���'z�h.?���9�d�Zr��:$�ƙ	��Aꦕ���X�Ff{�4$���}�cJЙh��-�E��j�j���e�����0���MS��?��������h��f ����R�G j��nZ-tN��q�	U�'�?Yê�4�=BFBïv�9�� ia�V�'���'����B,�����2���3S$n�4h�w&%1�m��??J|���?���~�td�.�5m� qs�ϓnfPx�i\�)˥nV�c����Q�i��r�EH�l����2<��h{��>y�l��?,O���O��d�<��+u���J�Q�z�(\�aeS:M%�����O�Ol���O��G`>&��Hg��-5��}@C�#Z�ĺ<����?���?���_�<��e<J�AЂ+V���e��.�5���i��'�|��'��Ik�7�S�8b�1�!�ȳ<�da ���u|������I⟬�'�z�q�~
�8bDً o�e#h%�$@m �l�i���'��O���>�ɖ!�����铢O�d��C�Z&?ٔ7��Ol���O��֗VC���O&�x��	�?\��ؐAX+8����ᕆNR�<$�0��ky�9�O���8B��m���,>�$�Y0GZB}��'�
�@��'���'���O��ߟ0e�"ҟy��m2CY�,M΄r�i~"_�����+�S�'+(!�່��EbE�?@��0B�i��``g�(���O�������>1A�J�x>�Q� E`��,1�Ƶ+�a��'�|�qJ��C3�pAg�*K9x{��v��D�O��$�9N���&���	ʟ��L4 y+�AFM'��*e	����>�p��v��?����?��-݃UE�I�O	���I�G-��t���'��EH�/�>/O`���<��[pI�
8&!�#�(t�%�u}�ሁ�y��'���'<B�'�剮+�
$�2o\�H&,���b��*�q)C�@��$�<�����O���O��oHKÀyP4!��h0��3�1O��D�O�$�<q��W�~L�IM*B:*����ZPpޭcg HD9��X���y��'|�'�8�+�'�t��� +'ؤ�T�_(����e�����OZ���O˓7�xxj�_?�i�Q�a��}��4�O+a��	���e�����<��?��t4"͓���2U�&���
�()а���)8# el�͟��Ivy"#A<M�p�'�?!���c&���a�A�]�j�e�	�#��I̟��I�h��j�Ȕ�yBԟp#qH�R^��W���h}� �i%�I�k9܈3�4�?i��?)�'��i�U��ޓ~h�A�7#ɪ��X@sGv���$�O2���7O����y�Ɂ:i|`�;Nۜh�u�A�Y��6�_�uj�7��O`�D�O�Ix}�[��㳇J0���c��U5y.2�*`J8�M�����<�.O�D8�����3q��zqM�6t��B��	�M���?��� x*8��]��' r�O������v����P�v�rL���i�B�'Qr&�,�yʟ��O��d^�
�"����O�^�J7K��f�<o�P��K���ī<������Ok�0l=T�Zs��
E�z]�aaθKț�'ܸU�'8R�'؆\[v�K���\��0X��(�@���Y��'��d���Q�;��H�0���j��X����a�3o˦8���V͌�,��0aq%
-<J���vt{�>ڄdA�rk� b�'��z�h�b�oЦCT>���';��7�bN�N:�aK���Ѝ3IN�Z�A�WJk�\�۱��3E�̴��u�\a��*0�h���L�+
ՈIZ^�m��H�����슰�d�1�i�,��A�'�b�'�V�S����D��ˆ+"��̑6��Zb#�!Kb� �VЅq	8���C�'av�)��ҩ|� �E���Fn8�Cǃ4]:�n�9HbL��!��>mU-���B�'�j,���?A��Ԯ@2K$�d��bȞb��UI��>�yr�'����.�2@�Q�ա�<:�B�a�q��'<!���P*4�+��¤&�t��'<��B�>����I����D�O����fq�f��{��o0�:5	.��͙e��k���O��u��,�v��+�j�Cs�+<t@ ��,ҢCH���� 7@4�PQ�"~��_����ΏN���& �h�}�eȝ՟4�IF~J~jI>QG�Hr�YgґB\q��	�^�<����@PH��fC4(� �14dv�'yx#=�Oc�# ��T�fe�租0)�(Af�'%��Yߌѐ��'j�'@�o�9��ޟ�� ��dH�y�3n3$v ��Y��?�tb�=	��ra	i-N�3ړ@dI�v
Fp�pQ���gɂ��s�'��I��B6�IS��QF{B�5���B�V,-�]�u�:�~b%��?���hOJ� @�����Lǂa9ă�=X��ȓp���PE��g\��13n��"�]� �)�.ObI
g�˦�"Ti���z�c�#��h��8%h�T�	����[{F��	֟�ɚIftP��!J�<��/F;�Su��[@<��U�!�Oी��Ӊ=;>�� �h��640<�%%�$~�4Q	6�O-���'�BjG)v+�0BЀ%�kb�/J,�'�'<�'�Ou�T��.�r�q���Q*ٔ��'(|leG� l�9	�)^�"Np!	�'p�6�O��]YL<Γ�?Y���雳-�`� .Q�zxN5�w(f��\E��O���O}!���A��	'�ʧ?q��n�;c�����G�1u�Fyb���L��p铀m���aF�P)4
�NK�)��<�2�ݟh�I��IA��J�Bq�uX� �$4"ī�*C����s��k$��|��!	G�q�l��b'�O�p$�����1���B,��v�"0�9�H��'I�U>�և�����ß�ke� JH!
�׺bi|ܹ�-�?�PȠ��?G��ӧ�)1��O�����`%@�j�>*]��[hޛE1$ ����S��?�'�ͻ]�����ŧ}�6U9��xؼ���?���?����'u�,Z��0D���]���!�W�y��'\�}��hUt���m�<Jm�����Y�O��Dz�P>Q�s��
8��2*� �,�����Yh<�Ifv�ȓ�EA�k�@n�<1���0۔P��"�x�aj��Hk�<��F�� KV��;�~�@Ck�<!�J́VsX(�FٍݢPxq m�<� דO=�ak�j�.������A�<��kU���8��/ۂ�6t�עA�<�o؝�F���f(>;�I6��O�<��!M��<PS���% 2<#��E�<9)�z�aa夋)!g���%�~�<!WkFa�R�R��x"\pJ��y�<�'޶ffhe�s$�#&~j�c���u�<�D���_� �H�A^}�mK2��k�<ɡ�_M*��e������g�<9�Q�_	.��g�}�^�P"��`�<��ØF2�\	�b׺o�n��&�c�<Ⴊ��\<�@ȶ#2��fDy�<�膴3O���%
1e��	[�%�@�<a�����!�&
�)r�H�1�I|�<��W����E��2L]c��u�<�Td	:C�jh���L�W��:P`Sp�<)���t���U�N9A��B�8D��4�U�c%�H�KVc��i��7D��F�ͷy�@t6�Ľc�}��6D��
���B�`Ӏ��kCH kR�0D�P��'N�1།ڲ���>��u�,D��
�m۴0�x#bk�Z-p�S�4D�����[6�l���l01�1D�Lj�`ƯAR���.�ͪ�N*D��E��&&ҭK���|��<P`)D�\������	C����`�(D� +R��<e��*��Z�_k.1{�%2D���g$��.��ٔ��W�ER`O,D����K�u�⼸4.E�Q�����%D�����$�P�e��d2�9��#D�<��/��,��XM7��d�7D�,��&]2f���I���א0zD�1D��R�L�_���^y6��(P.D�� G���WFE��}�䝣�� D��ӥ�FP"�L�&�zYQ��1D�g�øP{�S�	ŗ1h0�w�<D�  �Y��������g>D��8�H��*y���߿��=��;D�!���X�D�]@X���8D�$���G�%`����ܵ7��L��$6D�DK���=�Xd��,I�I�s !D�,�
L�y ��[j�xk����1D��0%e��#��\�qi�^��y�..D��S�	$��
a�
 kzY�Gc-D�� �L� e��f�x�z0K�(�F�y�"O,�c�.^�j=P�j��fKR�#W"OJ�sFW�7�z|Bđ�[3P�(V"O<�ZD�ڎܤ��b	Z/�}ȁ"O虂�fނ���⇺J>�D�"O��R���d�D3�A�-ބ5��"O&E�D�M�̠�r�����R"O�HQ�k��4� S��h\��A�"O�|���.Oo�H1�.��r+T]��"O@90w���C���E�V�,��HW"O�AE���Xy� t
= ��""O�2�B#]pp�W��Gj�B�"O��[DEK�<W�xA�Ą��	�`"O� ��N�"-\X�p�'�7}8��IE"OR���$�����'%P�X�s"O��J@A�u��8���,[蚲"O`���ŠK�"t��15���P�"Od��Q�PR���bĵ:~ؘbg"O�1Hʍk�����	e}I"Of��EH'[N�(�1�Ń~gbp5"O���,��d�H��B��6zKi�"O����$D +!��iA�*5�}s�"O:�a����ȝ��B�s)|m�e"O-i�g[�:�������9�*� ��'u)v���,y �h�($k��0Pg��îC㉗�l��틎J�����Y�Ejc��Bs�XZ}��7kWdt�~R�c�F1�[q*U�(�P�d��k�<i��μBX~��M!�D�*�c׆��$]�X`�(�޴&0fLF��Or�aH�3���x©A�d���w�'�YBFǭ<�����L�t��Um�;z��@�k�PZ�S%�1U֘�c�*��<�F��(��ѹ��_�Obd���.ZO�'0VD藁�0����g��z��pgM�^Y�y��%�0�C����8:F��Ҏ��$	B�90Sx���	�N�H�`�	���C	$|Kl��r�9R�Z��f�ȹZ a����WH�b�)����&xC|�/<�A+�c�F���I�Sq�C�23H,Ɂ'T�>H��阚�b�H-ȃ#]
*��H�E偨j�	���Ţ|�Ҥ���$[\��6!~�iR�N��2[k1.4�|��uB�(S���-�T�j�D�"측F(ͅwO��!a�߀f��j�ʟ9*�]z�L�<R��-h�\�B��Gx2*�9�H��E��1S��}{��� �OVu�cM c�"����
�f���l]�ArF$s$��)@$Q��B�t�n�3�E^/I�^�тD'\%�8��'�"�{��c��H���� 
�S	�P�6jR0k� �IG�@!|O"�y��O�$�I��5��w��v��pa�p!�Y��Fs�<�0��P�p�y$��4#�TU���Y�HS~l�
��g�L2�@L')Z���0)�z"��C�T�'[n�	e�\ '�����;(,��F��x؞��-tV`|��K�=Wa쥀5�[�`�ŉ��!Ɋ�8�DZ:8����@�x�������<a1�PMQ��q�T�I��H�')H̓	�I�!%8v�D�	�/W�H���8�b5�@�:2.�𖊘�V,��/9�ry��G=Y���$�#;֥X�mF�Y�<��j\�3�"2�oE�u�U����3-�v�P4c�v�I��ˬJ3�iL�S��
eVHk`e�73pn�8��L�8�!�dΊC֘��th��Y�P ��D��={b��o�����Z��H۷oު��rd��9��I��SpO�4��1q ��tT>���2\O�hE/�/c���BB�!<efΏ�yR���F��8t��C�!f�ɛ#X�)T����Sg8���D�RH[��0��
NQ��8�	�E�Yi`�ZTbA�vf�Y�V牅6@V\�G�/t������!t7G��l]�
OP0���
�����~S��q��| �@s6� ��� �3�Y}?����M�O.4�݆@oF���Įz
��@V�ڶD�C�	���Ȓ�1u����$
�d����>?��AY4����'�� !�&�S� ���Q��ލU0h�P��7}�ȡ��<��@0
k�{5���2m��ac��
!��{'���s
�(�N�9v���&��7��x��(:n}���6Gd�Lb��R-�OT�A���.��pa�-ȩ����ڑ#82}�� a��)(��ɨe��]�"B�I%FwD�;�B���9P$['0MZU`pO����A#᛿CŲt ׬%�)�;h,(�R/�-4�^�bIбOi�����	pS���b�*\h�⍙n μ��&�`�@�^瓻2�YP�RV��u��%�E;wEJ��쌬x���Sd �N8�\�G�!|��Vm� ��Ӈfݔ��4!:q
lxVm�=��L��I=�Ҡ��І�p<D/YN���%�E�,�E���t�':�M@
Θ��!�U�ljD�.O�y:c�L[�Z`�͜ZeR�3�l(4���˂�K
<��=Nh�ba�Y��Ò��<��}�h�`e�I�?�D���Oq�kL�:r��uK W<�X�J^�z5���!Mi���TK��A'T�|����<��ӂC>}�ȟj(�{"����B�4}��A�
�0?q���PI�q��8!�b�s� �8�h�O�QG�$&�Of<���xtd0�FG�z�B���>����f��d�3p;n���HW&c�t�K?�a�Y$�[�&�oj"�7D�h�M��&���*���/s�h�H��4�¯D)�>Y�'�Q��q���Ơ�a?�0m�98cF1�L_�Pޑ��@@i(<�6��8e Lt)�mN<6�m$!ְ>:R��ʥ>�ud� I1��ӕb�0��O�� X��Q�G�,�� �
�p<14F����y� �č&s�ay�ԑ/����\$ \�Ac6�-�O��[�!�;D��4��,�ԉ��x2iG1JQ�O  kì&�OL"\�c�C	y�a� %Q�n\)+	�'��h �)�h����(:p�y�'6��9��	~�2��E_�
�5�'(�Y;��Ҍ7.�h�'^h��'@$��2h"m"4��� ��
�'��a�k�L�������0	�'YBЃ�K�g����c�׌�LX��'�jth� ��G����T˼U��H��'�vܳ��+?�����	�v�:�;�'s"p����Xu���ғ{�0��'�R|��y�e[�d�	���@�'�0�hL��.P�ĠU.U��r�'�����Bgn"%ѓ#��6v����'��ٱN�4��H��(��@A�'D����(W�l�����&���'FH��0
_�S��@���ժ�6��'����nC�8�@�V�ɛ1B���'�>0�⤑� ��C5��#.���*�'��Y�"A(,TH���֨Z\���'�$�`Ӏפ�:�B���Td��'�4�����\Q8@��+�"T��'S���Β�cN�LC�拂L�hA��'SQ�@a�=J'�
s�K�71~�
�':�Ȇ�2$��!�'I"�H�'2�A w�ܐC�����U6%;b9��'�@�J�NS�jk�1y�M��4\��
�'� �C����jăP�'W�j
�'g ���+�. �H=�W��(a�	�'�葋D�O�Q g���
\8	�' ~��+\b�F��G ����	�'��T+���'�����	f �k	�'nE�c��$&�Q0g���	h	�'��-ʤOV?����s.W�5��'��Tq1ԙ�RdZc��&�����'(6a�QFH%�Hi �͉%K����'���q)�11������,J��	�'��L-UyXU��cX$E|��	�'G�U Q����MG?5S@T1w�
��y",E$�h�Z�>!X6h��^��y튔u�P�jV.I�A�6����y�BU�Z�FD��OA�@�F$��y�I�%j�4����A4N(���@��yB(՞R6<����,ɔx3'H5�y���LO"<�bY�ta<%�A�ަ�yb%H�PBC�7�N鱡
�y�ۯ$Z���bܾ�����ye�)2�+�(^&|Y�O�1�y�`��0��iWNQ'���E�y
� ��Jt?r�&,�'��v�<�9�"O�!(v���WV(5��cՈP��"O���ǦC �Uz�j��x��"ON��S!7 <(%��#yH���"O\ͪ�ǋXIP�E,}b�t27"O�a2ƪT(*��+� �c�0�"O�=��m�����f��`���"Oz�U�L z1���]�"O�5����9?QԜ�U�'|���B"O�xF�< I,̀��u��|AD"O�{Eɢ�"-%�E,(9�IQ"O��8cO�.x2a7F����"O������Ao�E!�[�5��ѣb"O�y0ց�%_������"O�܊6�
9CJ�3jG+z`ـ"O1�d�1m岁A1j�&-!j(9!"OD(�#JPA����"��>���"O8- tl�4��D�3BeV�pe"O�d*��%�a���	:,%p�"O2�KaL�<5Y��sa�@�&fm��"O0@�RMU�m!N��"m�����"O`����7KZ�c`�툅j�"O����B�j���u��2I����"O@8�1$��~�j�)4X�b"O���'ʐ���%1gI��<�nm"Or��FeO�uf2���P�@��9;`"O��B!�33�i�A\$/�8��"O�s�/�{fA�1����e"O�Q� *R&Z�hq��[��r"O`�VM�&*RXs$�s�r��"O�i�%j� rI0L���J���"O�0K7f�u�N�Ct#(咙" "OHxZ(K�� ���͒z��r�"Ob���T�"��W�c�H=�Q"O�=b�	�cp�˖ˍ�4����"O��qP
:V�~�j5�P�O�\93@"O�1�'�B�=���jBN��>�D̑�"O���W��J)P���-�: ����"OR�G��'��c-�tZ I"OHa��#
y���l
�,H�yQ"O��#�#�3�έ�UEP/W�xUB�"OF4h3��-O�t�:P�N�B��P"O�y��l�ZeD<R �G�nc�h�1"OA��τ-n�]j����뉷Z!��U��|���Ӊ����#,XI!���
�P��K,��ȱb�7/<!���!iEG/+��-�����!�DS�Y��[��
1�N�q�­{!�DL�Y�ث�Kɍ}����Gׇ8c!��K�ka�\i�l��e���	�G�!�d� �p�P�M'F����� 9�!�\�K<�ۇ�R3h����%Kp!�D<8H�(��ē�HH`��:)�!��5. j�RB�ҧ�\���ד�!򤙺Q�dQE�
$f��	�k�iy!�
M�q�7�]9W;D����n!��A&Dps��$��ݹ.ͳ|�!�$O�|b��P&�	gzt}C�'Rf�!�D֕]v�Р'a�e�b'��#)�!��>?��<{AkӥGd�qr��C�s�!�d6}�x##GV,Rg�4a�)L�|�!�D��U���y?[�-@i����.��$�(<��QS�i�J�E��~�f�aeȖ!"����Z/8��%��S�? �C���{�ac刟4| ��ږ"O��*��A�%�ɃtA�9� ��s"O:��W�x����ʤ�a"O�*�G�'�!����I��q�"O0ȃ�!�w
R���9�p@E"O��z`A̙m䬥y��٩@����r"O �����g�ʘ;q�ɯ�Ѕ��"Ov$	t�R��� ����;)��"OXUȳ��(����0�C��U�4"O�����.�=iE/�j���"O~�i���	8FLc'�f�Ur�"OlP�$��O��z`�	�d6f���"O��9��R� �P��5ΝX"Of��e#�
~�1��[N�q�"O�`��ePF����r��'^A^p�"OhM���a4,Çn�A)S�"O��'�s�ڶO�:��<h�"OV�C���|�<`�N]�'�X�3�"O Y"ԍ�a3T�*V�C�g�8�)�"O�8�c��e=����N� ��T"O>kl�Le¦�I	g(豈*O`($��6m\
��"O������+Z[��x�ϑ$tx�"O�$����[�LDh��X>	(5��"On�c���)vP��6I7�<�1"OB��h����u��;j��`Y�"O`�+	�3�4D���
�{zX8!"O*C�AYp�&L�9d��D!3"O6�R��~��`�� w^��y�"OjH���=9q�1e�w*�x��"OF�2bJ�%�A�A�S.���rR"O��3�O�>>ꔙٖbb�i��"O�| �b��u��(QA�4MС��"O"���F��3�H( �=�f ��"O�\�p"ܩ ����a��qj�!s"O�Q��퍗sq��i�a8&�C��y�,�-b��	�IӨe�P�YR�Ϯ�y���93���F@N3]JV=:B�
��{��\�S힤a7�U�x2
b��D{J|�V%
2�\��6(%���C���H�<y�&؀g$�����rb @�SG�<!@�ǲl�@�ړb��4��\z� x�<1�GG�K�%`R�Q�dZs��B��dZ����P��	�M�.��hO�>5�孕�@9�"�9cd��B� D�`��Z�A�Ԅ��KBD(K�I D�(ʥ*>\1�SB�14�T�D`?D����'5)h�+=#:�+DL!D�,iF�;@��3��Q�d��v�)D�l�Q�p�� ��n�=X0T�Y�2D��g�)J~��!�A(\:�X�"�<�����,���:�=0��9���z
B�I�6h���� =+��ǈ�	��C�ik=�H��aǆ'ˀ@�W>)`�C�I�^�!1-�I�Hqhq*Wf�C��{�ԭ $gR�
�*Y�P���C�I=όݸ�DӖkq�!Hc%O�lzC�I�+��bG^6�	��+�%�VC�	.��Q�㧅'bN\�m�X� C��'>d��ZE�W�20�Ş7SA�B�	(Z��u�[�U��d�"��9B�	�X��T7�
xH|���@Z�|�C�I�g�8�A��C�R�K�d�D��B��#>�x�s�� ~-��;��.C�B�)� �Rb�ǆ8�գ�KB��paQ�"O�%8t�:.��1d*� EK���%"On�����PR��Z5\AT�P"Of�HH�rx�0YD�CO���	S"O��d�=�٤EZ#�1�"Od�x��� #�N�j3�ڮ%8��q"OhDz�m�)��m2��?43���"O>�BaI�0W�����#��ku�Q�C"O�\ȵʓ�#���"N"	�4Q�"Ob,Ġ�#�`Ԫu��dú@�"Ob��q#�O�a�0�Z�e�����"O����S&\	R]���T�3
(h��"O�]ڃC�����@�-���"O؝"��
%(�X&��0�BL*�"O�QS++���Z���:�ܣb"O:��U��k�P��$FB&j���"OQ�0I�NN�UP�M�'�Ezv"O��Ч�$|�`A�Gϛ�ꪗ4�yr�IBd�hP0E*%�LMkYb���ȓcf�L3��!#x]��#�E��1�ȓ���W��G�=jD	�;�D���'�\�
ώ*��)[�W�	喍��'�>��	 (*X"�FI#|��%�':�81��B�Z����ӋX�Cs*���'�04ش�AJ���fީ�M��'� ���@�J���M|\���'vpD����Rچȑ���s�\T��'<�1�eD[�ބj�lŋnYt5C�'��$Z nC v���"5��;R`\ɍ�1��Oh�5�q$��)���D��D�\���jX�e;4�4N\ �
f��-5��ȓG�B��Aώ��*F���4��ȓy�^}��g�uw:�:�n�V�\�ȓ'P�T$l�la��)�S:Uz��HN�
��(JwKɎY����H�|�<��ԏ}��YaB��+܎������(���'�&�2A8�1{���k�GE%qx�=�ȓ��l�@��3����%☻%�Ն�3<B����ع`��	�E&]8�(%��)*�a� ��z$h͓a-S1]�$��=<>����Z:]#�p'LP.n����ȓ�-	A���N�hMˁ'��k����i��Y�#@<4�1���U�����ajy����E��IpW&V�8t�|�ȓ@�lp� #K������۠|y��l�t!d��:w �ؔjW1�J��ȓV�ҠH2� �h퀐х����ȇȓi�Q�#G��7T`���'O��P��#��XR7���-A,�PУ�	vR|�ȓ,4��E.V3~�h���d�m�ȓ.�)��H<Aen�A ��+��u��z�:A �� d�i!se��XJH�ȓ�$B/�1�2�k�$tt�ȓ��9u�ޔ6���Є&�m�A�ȓz����h�lp`�㛧ns�h���D�P��t��gD!ws����k�l-x�n��[�la1�͔C�ȓOϦY�g#ʏF�����h��Ї�3��J��A�w��4!���;U��C�I�oV�����UC�H��u�=��C䉯n8���SAs,�5@�:[�C�	�|������U�q� <��b�7s"�B�	�?4����P�U
����߹A�B�I7"b�),�W�&�cV��5`��C�)� *e1W�.p<5( ����b"OB��@M�B��!���	>Y�H�a"O���őD���3&�xaf"O i�Y� �����{��,��M]'�y��/��0�a�5� ����I(�yR�_�9�xI
@� ��+�d]-�y�D�N�����4-��������y�M?&�,���W�Π�D��	�y��Hc�����
KY2�#���y2/�X�
��K3 t9����y�O�?VM	e�Ƅ'���"P�Ў�y���"~���R*k²<;r�ˍ�y2 T-9Z��
�w������R��y�`�/b_欸c�L�\�x<Q�,�'�y�̕�2��QmՌUmB�8���y"cT1<�@c��Rݶ��g�Q"�y� ��w`$b�� =�隗&��y�˔=pU��p�e$�8�	 _�y2��(Ô�� �GYL)�K�y�fΠO:)�we>:�(t#���y�JS�y�����%:Dv��TkI��y�!��p������+�F�#t�Ƨ�y´�Y�`)�=zur��Y2a�����'-�ð�]J����@30��@��(�p��A
W�o�8
�-�q�2Ԇȓ
��;����x!C�,8�y��?lv=��LT�By0��*>�e��2�(�x��M `�@����&Jt���eߺ8�Єӱ^*��7(ݠ�6h�ȓtҤ��AC�^���f٤L1Z���a$![Ɗ�*�	Ǭ�O�H�ȓAnDУŭ�(\�Y�W��`l��K�x}zeE	�bV��1K΀:�H����l������LԻvp���^����v�$�R�kO��ꑇ�_J�	��1-%F���̚�!����ȓ6�`�Z�B�/�N(JaׅB$�ȓ^��9{#�Hk�����\�Cc2���I�<(T䗤R�RBn�$u�0�ȓ�hYH��3?�z�n�!`�,H��q! ���)H��(i�
���d��`>��х�]��Mz��]�Z�����4�1�S��:S��&��v�V�ȓ3]�.o&��"��r�.��ȓ`m�d�Po	�{X@a#@����v�T�*����K�"��j�-Td��ȓ8��͂W�Y=���ׇZ'
��ȓ!bD�@�-o�Yk�$F s$�ȓ���
�cJC�ݒ#e I����:�x;�	C5w�����k]�d��ȓu��}{s�>*�4�r�[���8�ȓA��!�U��w���q���BT��/u�	;⭅�=�ѠVh��@�����{���F�S�&��� [�f��3�2D��� KL�>z�XZ.E�Hp�0D���1�1^�-p� �??��Ɋ
-D�P� �G3 ��7��{�a�E'D�X� cAl���P��F$T>�q�0/'D�PR�R�C�@���AP9z��`��'D��; ���v�,`sN�3_�h��b&D�X�c��n�D`RCo���.��p�'D�������T�ڡI��m9��Kq�'D���!9#��!�lѦ*����'D��Nŏs7�m`P˔�dQ�p�w�!D�� ��Z�##�D sR�d���b"O���bD�FU��sI�h��-�$"O�hV%��e��\Q�f�4e��8Q&"O�� i��B��b�ʫ92�P�"OXI�3��'k�f�#��A<;)DI��"O�9�Ȇ�>���&���w�XC�"O����
J	S���,X�"O�iS�)�7� �C���X�d��"O��Pq
���L �,��M�ڭ�F"OP�4$`z�Y�E�g�V��v"O��8�.�x��u���Ʌ$�(y�u"O�����T���"�2���"O00Zd��
7�����Cx�|l�"O��k�� `��&Ĉ	Y��(j#"O�i�1�Ӓ~3Bd��!T/Oz8Y�e"Ox���*	+#� �	PA˂%kvY��"O�Aۑ�	p��Up��CPL�!�"O�y����f��@&$�4[ĠӤ"O��"�ׇ
o�u��0"��u"O�L�Aܤ*��Ն�.y6�I�W"O�M2`ܠa�`��%��(8)2�"O��*�ɑ��� �¤M+"ܐ�"O��P��֜ϸH����n�|pKV"Op�B���_��0�¡G����q"Oz�(�*�=q�>�	a��3W��2�"O.LIŜ?ik�����<Iؕ)W"Oy�r�=�b �0엑}5��(�"OX�	��"�P����˥G.*�I"O��"���ԡ�I�s>�Թ�"O�<5�ٞm�6��7��<1�����"O�t�ckR
�i��GD�.�ht!�"OB@� �N�)�
fC��rT3�"O�Q�D� 0E[��:��ݣ�H�"OR��EI\#��H�c��WC�5��"O:�Ӵ,�����wD�B�C "Ot!(B��5� @G&I�Z�90"O ���P-/Č ��E���%0�"O�бp�پL�r���FF?�b5��"O�A�fG�	y�U�&��q�-yu"Oz�В��Q�v�q��
�n�8�"ODI�Q	��s�h����v�lˡ"O0m1efăA[\�Tg�c�-�r"O�	�c c���F&�s�`�{`"Of��&�%
Zd��a#�#7�A"O���X�~JE�⡎4����"O�4��m�<~�@yu!���؈X�"OP��7��5EMdlk��Ca��1C"Oz@K��ď4�MK�ʈCF�h��"O����I�y=|��a#�&C�H��"O`� �\��=X��A��"�Y0"O���^�<a�&�:ch��2g"O�(UC�t��Y!��\-̵��"O2d�䝾=�Ri"��;'~�u!"O����N�T ხ��\_(={ "O&�� c	��Y2e�D5�:�"O$PSe\�i:�3w@[=*��"O�=Ȥ�@9R���}�aK�"O�mp��tx¸ -5V��0"O�T(W��,	ܕ�!�ן`� uq"O��A� �_�v|���
M��%0"O8��v��m�@\k�����=�u"O�0�0 ׆�Pa���{q"OYj�I�%�Pu�tn�^�h �"O"|�c�M�M�Nxr�����"O� Ι��mT�8Aƌ�d"G�(�� a"O8(83h�"xp�+��\�U��!;""O���*��hRH�e畉\Q�@"O*�sR �?Qy�Y�c,��Uq�Dʰ"O�,	1D2e�Qp���!fU�x*�"O*x�w ��hq �_�kVP�	e"O��P�%H)o��y3����[O�� �"O��Q卝L�0򭓖n?r�@5"O}�!�_2�$�f���$"Oh�E�< 	&��D�#ߠ��"O���	'���j3固�P��f"O2<�� �yg��pC8h�D}�Q"O\Q3�'=I"�9T�	�?����"O�]��7�����DSxn�<h�"Oة���*# �m3�֪`��"OP1��BԖx���H�gR~A8�"OH4��Ճq^r�y��=�R�	�"OX�JU7J�,���	J��yx�"O���T��5� �*�̠F�*�2"OF���ЄY9�a��&��=�$e:$"O�p�`ʍ�MD�Ă�e�H X�"O
m#�D�?AS�'vK���R"Ob	�UA��gR�X�̃�i:�k"Oz�RU�?$����6k�3���"O�@����
��� wl�&-�E �"O��C�eJ0*p�ʑ*��#�"O�e�Ef�L���<Q�h`�"O�]�p��YHn�h�'^;$��B�"O�\@�,�� ���OZ>�Y�"Ovq�w�N�^�T��;�T���"O���mE�]�XA���� �����"O�!�E��J@Sr�M9N�4 9B"O�)�&����r���7� u"ORA�C�	�Z�l��G 8��ܓV"O���.�1?fػ�ß����J�"O~M���(�`}+��������"O�| 5��er��N�A#�k�"O4��#i�)����ІȗVe�U{r�IW�p�B�2Z(�9� ���XN!�d�315�u��R�`@(9�A�n!�]̄����_�_1��;gÄnY!�dC!�&�b��7].�tQgB[�^v!�d'3�\�� f^#3+ ���HA!�J�p��T�C\z�&�Z�Q B!��G���s�.S�������W�!�Ĕo� q��+H5���� �g!�[�^r"��цL&���"� _!�D�Y�j���X�Z�0ٸԬҐq!�$g!0�e�!
�4|b���v6!�M 4�T1s�Ϟ|̌�ñe�U�!�$F �0��/��UjQ� d�"�!��;;ĸ�t��2 �us$Ĳp�!�T�+7$X"Ea�#R��0�1I�"�!�D� �8�¨Mt��(	�!�,E�8�ȒL
�9�U�Րo�!���`�#��v`
� '��u�!��ɠ
�R��6e�0��@�!�DN7q���CB��e��)�b��<w~!��&�ta��Ҧ2���Iu�
�t!�[�MpP��_�B����W�F!U!�'	~�z�*=C� �b0�F(!��`� �r��sA	h�!�$Ǒ/�I �@�6��Ÿ�I�\E!��:Bwf��,P�rvĬ��E=@.!�� `I�P�	�\\Q'F� ���"O�E�!�u���{�� \m�T)�"On���@;Q�lCUCJ>8pb�"OP��ܷ(��!�A`���x��ȓ[�H��_�#�� E'�1g��-�ȓj[ht�`]��̼C�P1Y�D��ȓ��*q �
z����(>�l�ȓ\mʸ�W�F�V�����un����*�ZD3��%h�Hy���h�hL�� ���"2�آL~�=�@��3��8��S��`@UJ� ��*��ܒ� ��`T��FA�d��<�w��}�l-��!G:�@�^�7�����Q�@$�ȓt�pC�H�BZ�P�`����b�<$M��.���c��Ofj�P$MOU�<1C@�F�@0��h�酆�M�<!�@�7q̙!!��SJ��#u�<B�FN���`��|�"�K�c�o�<��ʘy>$�� E֚1�=�S��P�<�v*κ}ߤA�#�^�D�sgXG�<�ŧջp�����a,nO��c�C�A�<���,��!B��#M�&M����D�<�T�,�,�%�X*à�q,�~�<�G%�9�VD�#l�!hspdp��[|�<�v��i���3��\�k5�0���w�<q��ӑ%n���{q�����i�<Q���&ݦ�X�dC�v�ri+�eo�<I�f��7oHI��%�m�PXS��An�<Q�ȑv�d�2��"|V�u��
�O�<A�F[D��0�nK�Fe��]�9����RJV�G�|�!`�݆�=J!�$׶(6W�6*|������~�=��}�I���9Y���6��2s.��ȓ)z���oҗ?0�P�/<?¹�ȓh�h\��
�}X@�����ȓuW(��(��l��lV��k[X��?)�Q��f
�C;�]�$�Q�cfvl��Az��� kִ���IӍx.���ȓE��!�i����P���F�l���ȓ:a$b���%��F-����upq(3���d4*s'N��@��&j*��B��K ��1��*�0��j�.�*�/�:vA�@��J�x��Մ�3m�� ��J�)�`�Y<��E�	~<�#�M"Ĵ)bF�ř>樁���a�<2�	�(?��&�C�� ��0�Ng�<ђ�ӻ=t0�!N�J��W*`�<)��" ��W��%Ռ�� �e�<A��3?�Ll����h�Кu*�I�<QslD��.EH�0�R��T�|�<9��(�
}� �o!��p��	x�<�K�K��8١�@�-2A�%�u�<q�ͅ*l�����,f�����L�<YҦ��r�:�#��6����j�P�<�T��"ml���H�0B��Tn^L�<QV� ��$�M21apԂg��]�<�Q���L�:ClZ-}�7��\���0=Y��WШ���	�Y�i�5ʔU�<���ȮI��jF�I�V�,�6��Q�<��횽%�A�BF�p�ș���i�<���ډCʸ�0�^���-D��e�<q�)�a�H�A��wp���g�G�<�rn�#��%��ɹ-5�`�c*\�<a��F�9F�%qg�U��Td�W��V���?�
�S�? ��%L��2�}��U;YyІ"O �5�,`ҤeaĆ��JH�y1�"OFM��+�,ڄ�hD埕1�0(��"O���¯�b�r��d��;w��|��"O����Y	*��@�����<�W"O̬h���9u�`tX����t���"Ol���Lá3�)�A�2yz��iP"O�87��	t�t3T��.Q@Š�"Oz," B��=+�`��ز��"O���Q�O>�He�\(pĄy`"O��4��J|���
T\�x9�"O^%Ʌ$A�3�
��"
��G �=�B"O~4x�oR�>�� �&�[,�f9�0"O�����XAP	����0��"O���4eI�w��Б�e�0�K�"O���J�]��4�v������w"OT2s
��E8*,�殈�#|�|ء"O�4����s�襰Vc'd�i�"OL	{�!FP���R��)��c�*Oƥ�c�&p�<ӕ�:t��W�<MS7xt0Q��+v�R�Яey��)ʧ%�� ��\D<RLk�8Ҧ��p���2IOZ�F%��$��md���ȓ0l��8�\��	�v�з����]������{w�G$ô����k��
������D��@^�%�d��ȓm	����[Ѥ���O b��0�ȓzLP!SPm�66�aCAS�6m`��[�u�"o��g��5�e �m���^h���TO�lq�'��H�ޡ��::x�B�C/i�T�HS��J��ȓd��D���7^}��fJ�D.t��KD.a��÷Zn���(�01�9�ȓLNX=3��[TZ�#B�(L����	�Δ�ר�?P�yZ�/G�I�%�ȓDf$��̜�)@z�`r��5cW���[fT�ga�I=ތ��*�Q}��ȓ"Ո0r�r!B�(��*m����Q�<��G^9��D8 I�&9��h����1ᐪ�
��\JcB� 5�@���6���!��q�a+`�OvbdE�ȓd�\�D+ϱX@���V v�ͅ�Od�`�hU�lp]��H�;����ȓWn���AI�
&A���N�Z`F���J�P���SU< ehqm^�>��܄�2&\Y�CB+C�T�����(�&��ȓ+]`v%�#$��#T�A2��e��x^e�nށ�h9S!�
#[B��	t�t�ϟN ��H�$HAE{��O�<�S�� �8jkC�4�q
�'@�����۷z�-�S�� �"�(
�'��p��
j��	��ӵ��@�'�� 3�D�n�|kBŝ"/�j�h�'	L`)s�gZP� b'\�Ld�
�'���Y��G�t�8`J�lI�i�(�	�'��Zf��\yP����ůn�p,��'N�{�>�,-�u�,�̵��'v�˓�3X"�L�e�Y;��M�'�^��CC/d���ѣ+� *tB�+�'�� 2��Ԣq`)
@Ύ�N����'�8D���d���۩M��T�	�'aY�E {x�����7�:���'nfI��*����X��]x48A�2�)��<q��u�Wȉ!��|��K��y
� �t*Ќ�y�Х;��9e�|�c�"O(�ԍB/"����"�)�'��'J�)�n�0y�#T�R�D�� V
KZiP
�'s,=	��υ�f$y�b�K��as	�'rН��!ڻx~��`K��r��<P	�'�}��痥=�:�cR"��}�&E
�'�Х`���<l� 2�A%}<�i	�'�>IJ��H��#v�B.=5nЁ�'I�-q���<� �p��h=�y(���)���&MK҉�`j�*x��L�y�`��3(�ȟ�p	��r��)�y2oT��DE!�(_Ic`'���y��`���ï�8>#�DSAl߶�y�e�iZ�)��oF 3Y8��0��yb��&�zر�B!)?��pM��y"@)A��C :	�N��w���yb�
�E�&��|������ym�+����f_�|��تC�8�yB�ƣY"��`�ـ{�JI���B2�yrKOj ac�ń*�b���L��<	��d� i�F�3���{=dyq�* j�!��3<�^aP5琙Q<L��h��D�!�A�ސ:��F<H���Q�S�B�!�N�_�z����X	�y�sJ�:r.!�$.e�fu�!��ॳ0	�?K!�D��h�Li�@B�N�h�'H�K�!��`��Ñ>�����9H!��֯p{�M�TbH9.�[�מ*[!�DZ�h���9Ê_�*�E���T=!�d	�����eۂ�UA��X !��]��i��^�le��@�L�"�'jB�'�$!��� (���8�ʍ$3):��'�z���>B����Ə�;��"�'���(��c�ʔ�6l�u�FT��'���A�BB���I��k��x�'8VY����"eV�r�Q�b�t0�'�Z� �L�:hze�$C�>[�'��UiB��f	�!��H��o�D!����xr+Z�M����oYD�$���!�?�y��>i�T�p��B5�:�Ý��yr��0q��R��� ����e��=�hO���I��GUѡ�K�;m�� ��
?�!�$�Lp�)5�\S�p�{�(+Z�!�dǓi�@]��G�!r�Bb�H�!����p/��Z���7*j��I��
n��'���'@ldP�*�)[Ɇ9r H��w()�
�'���a�/���A�`À}b�@�
�'��֍+<�ptc7C�5xa���	�'#ly���:Bͪx3��P�v{��!�'T�/����h�/n�n�Ɇ�S%�y��T�F���4�
���M���>��O�l� �B�j�X)� cܤ �� c�"O���B��7n����;H���F"O��Y��_�4�k���k��(�D"Oh�J�MO*l�d8���FZ<�#�"OʸYR(�p�8UA�&�ԩ.!�D�Fl��eEF�c�l��'�
��!�-pdiK�È�n�#3���!��<j:���˃?L�ʖ��)-!�G',�Q-��:80)xu�RL{!�$� 7��c�D�
�ı#�&B�h!��iN��`S;R���R�Æ�1�!��Z�\X���n�Qh�@اX4!򤋊�IW�,�\�� ��$kE!�� �葱΃�^�α����>Q��@H�"O�4��b[-1w��+E�Š
��yP"O*Ī�hS4��!�P�0qHh�"O�|� M�T��x:rm�m@�'"Or����ѶL�R��k�DN� �O�!�E#�1.��if���X�`<I�-D�:��#"�p� ł: (U/*D�؊T��=���ɳ�;6"�@��'D�(9�B1PD���M�7G����a+D��3�Q)8{�+�62ּ�R��'D�p)��F'��j��b��l���8D��!ǩ��	L�����3^��bc�,D�HS�/�x�8Ն��_�숥�)D�̢��N���m\F~�AC�"D��:�D���$k�m�-FbX���M-D�P�冢{'�}�g�pc*�)���O0B��.F�D�c6m�5o:m�a;e4B�I�4�h�����R�@ab%DM4R��B�I/	��4�!W+?ZAF��QzB�<*�r�Ҡ��n
6��f���C�I�gXf��#��'<�*��gN�5[,B�ɐ�0aГ���KQ�؇��W��C�I�dN��{�Ę����%e^B�I�u����'R��h",v-B�	�u�0��oO���$9�Ε�.#C�ɔ;;�����5&j>%��NkDC�I'�����?a	���b��B]~��0?��M�\Ni�"N	B���E�LM�<��+
(�(P�WƓ�xd� HN@�<ye_�'�-&P;A6�)�l�W�<�2/Z(a�܀-�"Y����	S�<�r�U/�}iƢ!WgP���#�L�<��� *f�����j2d�f�@]�<��?à�� �ZSN �s�[�<��jB�Y�vK���������Y�<�RdQ6>�T�I��T�v$[�<�0��?7�(��E&�� ���2�A�r�<����+gk�����u�`Z�[i�<��|r��C��3ZF�H���	K�<�vE X R��c�E�kQ���Q@�C����<��HB{�ؑ��O�=��UZ�Ĉd�<� �4n�}:CI�9fdIWn�\�<��+�v��r@5F[����^m�<�TL��8��<�2i5y���z��h�<�קR1#MH9�gF�I�-Z�B�\�<yw�ҁ3l ��˲^��e2�C@�<1f�QT���e��~w2�)ġB�<a�,p�j�Y�F��e��mA1L�C�'ax"�̽N[�q��X
�����ܱ�y�-[�,���Q(\��� %� �yB,ӭ|vԙ�sc-u�$�B����'�'td�R��?F�,m1�b�7~�4 z�'�ha@��%e���C�ւf�>�J�'\(B��'q��ꥄY�\)̅3�'[<��D�+���ɤQ�h.� َ�d1O����)jX��06h� i��:*O�Q���n�����W������?����II�v!�a-
�àa��ތbmT��5�L�H\���P�'MڧQV���6D��{c%�e���W�x�D���e2D���$�S�w¦L�GkU�rb�T�-D��Õ�3]��=���r��pyR,�O��c���ycS�2~��
}�̈́�ug0�(P�ҙ�,�����>�"���S�? V�+E�[��X��񉚞N�ܸ	���Q����Aҝ%�^T�w�.�lDV�'D�������A�g�%�08@'D��!&��
Tr�B�Y)H�l8�,$D�H  gG�C�a���}X���� D�ܳ��ƢU������&Ah�A0��2D�,��S�I�<�Aҥ՞QL&�H��2D�0�%f�#py�ȩ��V�w&�IQ�1D��:w�E7^�<�uÓYS)/D��[4G��J�R�WC�=3>X�k D�����H%�H��4�f`L[�>D�4�(�:Fu!ڂ�D*(*X�d=D�`���^>P���h�6H�F�i�<D� ���HwZk�A�6i�lu�.9D�,
V��P��P��C�W�^�s�3D�D�v�R4��舠�XKJ!q҅/D����R�s6���@![�P1�-D���tL�3~��*M6�BxR4�)��0|�`�&y��XcCa��~E��L�O�	[���@�6{'���#�H�j>A��9D��۔"����g�o��6D���p[�xa���wi��a�y��!D��y�j/�`��1%	%����"!D�h�����3�j��"B��&X���I,D�$Y�'�E|8�f%b� �s�h/D����#q&N�r�.Z5�#�+��;�Ol�$B�E��\����3e��kS"O�-C�g��Ke�=k���,���"O�0�ͥ7��,h �Z��8@"O��RbC��t���ōLR� L�"Od$�W#6{�>��&�<-�*5
G"O���G�X,UEAC�eR��d"OdH�C�d�&�� M8���"O�pT�L#~-���c#�GFJ1"Ot�����T�v�!�,+� �T"O.]1B���)Q�(��=O��љ��7LO:��vM�8�1�^O��@0�"O*<��E^��n aы�2{m�"OJd��%ѷt��
���� sE�7"Or�[��� n����J׎am�\:g"OD�Z���	mQ���QV��R "OD�pm�9x v���F��IӃ"O���A�7�
)��*M�H
��a��f�(�CH*'�u�C$τ<t�ᄃ6D��Q�����3��Fߴ4`�'D�z֢ʑ�� ��W6s4����+D�$*Шǅ7x~`@�cQ%aK�E���(D��P�H�S�y{�"<V��(D�ly��.��F���b] �$:D���Q�^��2)zO0E� �	�#D��Ձ�U�:���c:	��" �+D�+V�լȥ*�$^��[�'[l_!�[)�*��[J�[t��q�!�<=�ĸ�a�R�h�0�+!��?()P�mC����럖p�!�G<�`��iR�vHɉ�)��!�=z���h�aZ��S(ȸ
!�$�N��1p��?f	V�1�FA�D�!�$��_Ь��D��a�Ld�W�T:y�!�'vI�mkRaF�1���XP���B_��$ϻ\p�V�9C����(�B�I�/%��`BZ�3�jPca�]<d��B�I7R���0�ʱn@�3!J�M��C䉮+B�0ZQ
կf�"d��-�JC�)� �)���E�0L(p�U�4!���F"O�eK�!��X���$bH�~]�`"O�H�E B�D�г��Ji�p3"Or�22CS8�H�g\�uL���T�IV�O�̺5��.-���c��#(��	�'喕Q0�N䠲��~㞄*	�'dbt��
#-P0��aF��(���'O+E%I#/�>}�qcP��5��'�
(�f�Y/(N �ybĂ���	�'W�Q����aGP([%� X��'��,�M"�ժ��\:EN7��􈟺�y�ѼP� �%�
1��r�"O�<ᒠ��ben4@3�F�M���2�"O����V�yV�q�3K
1�&����Iz�i��H7X˰��2N� 7���A��<D�,�"B:�l{wGՁ:ut��g-D����z@��#�Ul�C0�*D�Z��%VY����"ξxZ� =D� j����C��E1��=jġ8r�7D���2N�%~�>��S-\���3D��b��Nts����I({w���0D�Шƌ���� �F�&!rD�&;D�x����6�h�Ǥ�=-jл�
5D���v�7bs���H�<��2�M3D��(W��|���0�φg���2ь�O�=E�E���B-XP P�Qɶɫ�@Z !��0 #'	1*�.�z!�ϫ�!��n&�	���_�tp")���!���!Y�D��C�r�� �c(��e�!�d��g��@[anK���y����6�!�ۯ0U�������j9+�ŒW�!��C��|ȡbP�}��ѧ�ߝJeRO�pr��!)9���� _���"Ot�i�Fĉe���d��<�:8��"O�4���S�u�6�P���"O Q�R��P�lc&�`~��Z2"O��2F܂$e�lC`GWbP�Z�"OaHo�0�hݩ¤B�-�.q��"O��s�G���$;1a�<�,ب�"Ob��$���X���Q�ZO&���"O�,��H}���2�oS�LX���"O�P��UZ ����:�����|��'�B\@&&��0��%I���k����'��䀶�Ҥ&x�0C�-;Z����'R��D�2%r��p���@?��`�'�Е0f  .�U��U�3K-a��x2(�5<:�`�
l���ْ�C��y����6آ����M�Z��R������<���~JfL�z�DX��qIA���	J��C䉰:�b�As��8�X���dG�ClB䉁7��{�	��I`!:c�O�+$�B�ɯ'�Qj���7�t�G�K�B䉖�2%s���|�+�?��B��;�>�'��e�PL�fjE�5Ȝ��7��'ړ��d�f00@�eGV -����a�'Xўh�<�����[Wp�+��L�*��A05NY�I@�0*n�;p��"%��Iw��%�6D�D���n���$�%t�	pc2D�����6 hQ�D�� 6��@�3D��S�1�U�����Ӏ&'D� 0UG�����@@%U���#!1D���c!V�"�P�j ��[[��R;D�@c�a
l�j=�g�Yw\�a&D�(��h�p&�%)�A��=H��O#D�� Tɳa"��b,Dqy��1h��:�"O�h���3�$\E��.s�9W"O24�1�	�O
���TK};l<͹w�d-LO�ð%��-ƌ��I{4���S"O#�o���� 6/�7:B����"O����%��z�Dŋ��_I2��P�"O�hզ�N��,H_�Y��"O<%�Rڬ���%�ػP)��"O�%��GC]&պ�]�4��E"O嚃͍�������X�~5�"O�{��Y�:xI�'��}["O�tb ��^�r��cz�E"O|,��g*b<����	`�]
&"O�񃀐9Hޮ�2v�H�A[fQ�!"Ob�����n#f�X1nZ�5>8eZs"Oҹ���8yI�yP���֌Y�"O�i1��66H<�Ԏ�$��py"O�% �� �H�R�e@hR3�'�,X �ŵk�.Pj�唘E��8h��6ړ�0|zS(�%3�PW��1U�H�Pr&]c�<�qȔ
dۚ@�DA{z5[�ƈ`�<�ԣ�*)YNl�A
�qfq�q`Y�<yE�;)&�;�/��q{�b"+TTx�l�'�p�H$Ƒ�d⒣�>$'*�q��)OP�4狣;0N�Br�<`׌��S"Ozl��cM%	�~(yt���a�Hu{��'w!�ę$�mxfb��bP��jGR#!�d]�Qdz���F�h��Q���d!�䝎r/�XSuר��  ë z_!��� IM�9�A�]4��1���9K�!�ǴlB�C��t��`a��;��'�ў�>�yaֳnr�"A��y:~�*��1D�`�G�=v�g�@Y��H��K1�	J��4��n����%����F*( �d�<D�dI�)/��qiߜ#�и���8D�0�� ",�I�.� q�<X�G8D��ش�yD
����0N��JA�!D���M<-���ã�+/��j�C$D�4�w�=@�9�o�4�XC��=D�hm�*?�bd�g�Z6s�r�2��;D�l�EBX���pT��P��:D��Ɂ���wf��5�Ў}��D�'&D�$Cq��`��,!g��;%�^TSB�&D�P����<:����E$(�V�
[�!�dS=� �	�o��E�N��7�ũVv!��Yjl��V���ܔ	$��0^!�d�Y��%�{|�<P��9 �!�$	6V�21q��Fs@$Sg�6^�!�ą�A@�D
я[�l����p�Z�!򄖥q " ��Dc#^DV��-5�!��I�H��Ś`9�I�F�֊u}!򤒋���X��F�D~t�s7I�'^!��ܫk0���Ĩ7NjI��甲XG!�Ea�����
J-	��B�A�^�{r�B�XB$�꒨�����E&�1�!�,Aā����de�$�e���!�ּG7���N�* R\�c�d i !�dF�<\�  
�
c������Tx�!��Va,��h�h2]��]�3�!��Q4�q��#���Q��;��yrቤ'@3Ҥ�8T��N%����1ړ߈�����/�=���GB�Md�%��Z�І�I�E��=�d�:0�ڷfI(00C�Ƀ;�	���=;q����fLgj�C�)� ��wo
߂�"��fH� S"O�y�%E���]c�cZw�xȉ�"O��Ko�J��F��J�ܕ{��'����qr lA�Dȏwm�ՑbcS�PsB�	��ȉ5	ʲX�k6���c�C��!xq��M=ei�(�wN�0+�RC�Ʌ_6L1����I�䂴�GN�B�	1���Pϕ�9P�Iy"�%s!򤋎|�.a�(ɶ`3�����Z�j!�؎W�بb��݈`��z���"��	_x���'O.�W��\H��D�[�n$��'�!8��n�) F,�Z�fUz�'����ьK�ZD:����Ov�e)�'\��
�֜�64��H�>��T
�'m:��Wi ��P��Kա7�^�y�'^J�7͐/��4ZŖ���X�'�-Z��U:^�"i+4�G�xR0Z��D*�XY�WGޯ��hx�G��z��+�"O���&�/��2'��Y�.�9�"O>�����n���5�����["O����A��9��]Cp�˓z���A"O���g,��{��p̂�h��"O���aF�	Exqx�íZ� ��"OB��3��3�x��L�8�
\��'Bў�'���O��Gk��("Pnԇ%p�X<D��p�E+m���EыQYX�Y�¬<��h5�m��=E���rK�ML8���s���h���D�d`
�V%�̈́�P[r�JGe��r"�y���\N���TZ6���ʕ\�x�A�<\� ��q�t�)AJؽ�F��B�e�=���ڭ�v�фc~Q�nXjUP��p�\L@�a�D�v
C<Ajr��Iן��	�P����,&�C�*�8=��C�ɰ}�,Y(�(���9yt�ڙ}�LB�I)�D�pԅ�2p��Ka/*Z:B�KY��z���9�Bl{e�L�n@B�ɴu�H���TT� �"��*ʓ�hOQ>9���C�}��s��X�#��mP@:D�,�G'�b��bEJ�`�!3�=D�� �K�*&��3�8��1"=D��Ǖ77:�Tz��7+*�����<D��[#��?P�x���뚸	:IH�<D��!s �fk|��AZ%98D/9D�T'+�:�Q���?���3զ!D�t����"�8t��	�|��,K�*>D��Q�F_:z%����a
yC��<D������A!ܱK5�:n��1%j D�\���,3��(�A�{�ʴ��A>D��
#�ݖ� 9P"cL�l�(;v�'D����_�o���!���>��� �%D���"E��^1P�#�>��+a�#D��;u�	,���j�
D�ߖtd�!D��`���&�����$�N��,!D����ʛ
˲��� 8x�2a1D?D�,ѢݙG�@���\3P�h��&�=D��"�C�P�@2Ě	f�hyE&D��!��@�/�&43���B~���0D�`���#(�J-���U�^<��g+D����Θ�C�(afkY�1f���v(D���L�g"�� �	~6H�I�a"D��c�!�u/t�p�ݫ/{||sd"?D�� 6�Z�@ʠ�)a�Me��#V%<D���@�d��`�V�Zn�LZA�8D�� ��%�	4�$�*�'
A�*�"OT��`N�<T��h�X1 �QW"Od��]�XE±��g7_�T��"O*��c�uP��[�fިu��Q��"O��g,�]����D��|��P�"OPa��lZ�$�@��é��<���`�"Oj����@$�^��O=x'�u"O�Ԁ��C�~�.�%F/l
��p"O�����%�J8 ƃ�t	�(v"O���d��$ g�4_�����"Od�3��-Uh52�J.�"�xg"OD@�Q.�4%z��땯р�V(9v"O4�4�)��#�V��@�j�"O$QPr�0K'NHH=��5�"O�4/�Z.H�Z$旭V�b0"O��؃b�t�2}��%��Y��D�V"O����N\ʪ4�2d@�s���(e"O�Pq�R���rc�C<WѤ� "O�s�G�|q,�hASh�4��'"OqjQ��M�p7�ʺ7�Pa˄�4D����ƞ�lA\�y1�T9lQs�-D� C�E�$M����`�1;aش�,D�\�����t4B��S�e��C7D�s#�Q�)��a�pG�(��	���8D�<���GeԔ��$�p��1�g�8D�G�ӹ܊���� q�*$D��)��QO�Ҍ+@�����f("D��w㇛FA<Y[�bA�?���f"D� (q�Bh�PКBܙZ������ D�\{�H57Heq��?>Ҁ�u#=D�P:�$R"N�Ƞ ��)��9��:D�t �b��v*�%�׸6���QS�9D��`0JQu@E��K@�M+� �FG6D�@�ā�:F� P!N�)Ԉ�zb'D����ťefT��Y#�X f#D���n�>���B�W�)�@��a"D��r��[�&哀L�r(,�à3D�4{%���X��KdfF21���(��&D�p�H#�^�X6�L�Qq�#D�l�d��c[By@�%��5$E)�)"D�(�5�BS�R�0�2��X-D��k��ٚ>~v��Aݱ3��XӨ'D��5Bڎ�^�K�M�n���r:D���C�y$���C.>ny�#D�t���@�(��X0�h��#D���LM�?#��B�k�4'ri�$�+D���N�-�^蚤�B���;Qe.D�t�3��m7��!�FP��Ԃ%�+D�X�V�	�Vi�̈́!/����EE+D���A	�.bv�̓ӎ'����K<D�T��LS2{eZ9�w��X��`��>D��2d�=��PSv�+@����A>D�p��n��\�U�V�7F����<D���2�zڬXP�U�FxܨE;D��r�	�mNey����P1rQC�9D�l���L}<t����M���y�7D�����٠���o��Uxy �4D��ғ��C���aW*��;} �Y��4D��y�k�J�Šd�Ǥ	!�r��1D�p�Ke��!A���%?a�+��+D�tӢ�.'k�5` ^�J���C��)D��i�B�LG	����Z�P�g�%D�ӑÖ	XሽC �Y�Pڴ@`/(D��`��N�+�9�a-�"n�yD�0D�� H��a\ w�,�فR +��Ye"O��ֆ�%2� ��#K�c��<
�"O�A�Ǯ���"}�Ynj�ٗ"O`%re��1rXx2ӭp+�p�"O�� u)W.T�iw/�I@��P"O�i�n�8~�lqe�I���� "Ov�)�^B�J1"07�
���"O�m������{F���̙�"O>	��e=D� ��`&�#��a	#"O`��FҷJ}��cB��T"O�	ӁN�:�|�3�q�:g"OJ��E	>1{p`�OF�Ma��Pv"Op���5� UiV�Z7���F"O��)We�H��H�]��P��"O@u�$M�!���*��>s;����"O��2VD�b�ɩ3��� *jAp�"O����>7��,�"�;|=��"O����,&ekDa3A� �ک��"O���%߿|�p�z�/į���4"O��{V�-b5�ġd�L�.�"h��"OVQ��k5o�튒B���l�8�"O� ��._�D����&g���"ONZ�A���	����զ�A"Oް�����ip0��%F�&(ܸ"O�����7wM���$\-K�"O���ǋKgf-R���=0
�[�"O�aYԈƵ=N H��
Ϟ�v"Oh�;!��
}��j�g�F�T]ا"ODՒ��9C��ȓ&N?����"Ob�i" ڗg�آ�G��H*��"O��@�A:���������7"O��@�CS>&�j1�F%;�3�"O�ٸ��
~T1��eͭNa�ٲ"O�Yb�A�?��إ���: �"O���#�Yɖ4�3J�o�����"O��Ӆ(]3�>Mrdi�R܈ar2"O������I�F�ˣ�4��"O���fU*@�2���g^<�F=�S"OZL���"��Pe�\`�~Y
�"O�u�NB�\��@!)N'c,1��"O<��QG��.�&9X!C�~�J`Z1"O $��#JH���r� �?�΀��"O���eC@: ��k-7'��(�'"O¹�������!��"=�PXg"OT����S�|��`�g눆c��͹�"O�hG�܅|=��<Z����"O6��K�
��H�,��<��C�"O�q����z��h�$�dc"OM�qH��45� c�B�Щ�u"O>8�SBH9*�BQ�5�$|�r"O$�׃؅w��}ca��F|U�"O&��N
-	��S��|�4s�"O�5x�év#�@0��(�a"O��I�$N�T �A�-%^ɲu"O~��d Y	11�hq��+/��(�"Of�"T�8���Z��/q�2]�"O,0ZQ�ԓdP��EΚ���`��"O਩b�.����է^ ��#�"O�I��$�1��Xs���C�"G"Ot�!L�4w�"��V#	)2����c"O��hr9n0F T��0g�:@�"Or�K5���r�
B�Ӳ~B`��"O�����t�1"�C�-9�tA�"Oġ��'@6A0��I �\ȹ�"O� H����G0'@B��E͔-Kv�*"OLlې�,���*0��s� H4"O*�R37(B6xqd��U��A��"O`M#��64�L��c�}�̉i�"Oli���	sش���B�1�r�j"O����Ù(�,���!�X@�"O}�5P�wZ �B�
@*XJ8�;�"O�H�6�J<6c0�V䉾T�d��"Ot �7fG�m��s��v��	�#"O�,��
:I�T�7�y�����"O y�`
��.�pY�dP�9ߨ`"O�����l�����K*���Q"O�Ӳ�F1k��:fg�ur����"O�ɸ���[���f��Z|�ܚ�"O<�� ʋ�v���2�?�"O�I�g�Ƭx�4
�$V�c�"O���()A�qZBd�<$WRP!"O�,"��͡�D��3�XUQ�R"O����D2(���)p�Ζ_�e�"O�i�tKC;!^��A��'���r"Ov��fi�%[�J�(�?Z�`)�"O�Y'�X�L�B#�9�,<��"OVŪ@M�9ѮU�Q�/M�����'���Y��SP�Lf�Z�)'�L�z�`E�2D� �˚�zTE#�e��j�� 1ړ�0|��b�'&��;���H�C@�c�<Iq�d4����6�c1jZ+w�C�I(�|��!���,��)�=ݞC�	�zL�٘���F$���s!��B�I)a�P���1����0:D�B�	`��t�"������9�FB�	�Y�3f'H��ڤX@ń� <b��F{��D���P
�P �CH=�8Y�ߋ�y"�B����Æ����z��A�Oh��D��a2^�i�B:vFd���a�!��U����V*�DA�9IkW�]�!�I����U��1�!@L�� �!��s��PY�̯|���p$j�%,!��n0��A�2s�H$#a�A1�!�� Ʀ
G�ʸ	��"�!��^�����IO�y}����d� u!�$��P����Ԗk^t�����rt!��ͯ9���ī��f��A#��#\!�$>�"i˅O[#�p0{�(W�X!�$ȧ����c\i:ĳ0&�KN!�d�\Dxj ,2-�^`��4H�!���=8����%�O�P��Q3$�/>�!򤖏#�����Y��]x�L7zv!�$^��("F���6|T)r�Ϋ]ܮ� �"OV�#�7xt4}h�ʣZ���"O�h�g�V�p�85hW�f�Z	��"O�q��ד;��a4��(VϬ�� "O�`i�e�6s���]{�(TYt"OP��犖��f�i�C$˔�:�(lOf���	�N�"b������"OtSl� :���h�^U����[����	Jsd�knR�)��U��oC���p?� ��;z����ܛx1rT�Ï�r���'�b<�OZ��� 
U�b���&(�Hs��>9K��j��iƨ?T�!h�D�,?�)r��Ç�!��
��m1���2$x����&�b�2�O�٠a�)^Z����Oؚ�U��4O΢=�'��O��)5��4qS	ֹ �*Y���>4���T'R4~j�ɒ��<��
k%?QN�Gx?� �xU?XN�S���s���"O��*�I�h� P��	q����"O�Ż�o�L�FIquÆ)��$!�"O�5#w���T1�DYD� d�xm�:O���� c��t��'�4�����Hܪz!�_��Y��:�v�+��o�!�
8P|�r�A^GH�٧���}��$:�I�T�?i�g/ �5^rP��$@>(h���R�7$��	��������k�5v<�����Dn����I-t�L]�-E����a��S}j��<Q�'ʛV�ԍY�2E���[��5'��9��C�	�$�9h����4�xƎ]�F�>1��I�6����k�,`i�̋!�D'�*���'ü:j	QǢ�]��y�I�	�����%t��Q�DW�$C�	l�A��TU��U�lӝ(��B��9��M0:���a �2��b�<�>a��$���/A�|�oB�SND4�TmY.I��D�>�6�{�KE+ZCD1!$oWGGqO6�I~�Ӻ��Op`�\�c�|�8���7e3 P0�"O��k�@�U�
er��N"�(�Q�I�HO^ʓVzV�Bƅ���\E��\�"����G���g��HV�!e Յ~�vAs�OF��t*��,(h��6��))"O�KD˒*$�$�2��U�u�	�"O�h�G��'hOԈp��� n,v"O>���Cզ2�� ?w �t�d"O��[��Nh�Y����,T�&IS3�'��ɧ
=�������zɈ�B�,x[�C�ɺ;3(ȋ��oPl!Q�@2��#=�$-1���0�P��1��0XK�E�z̆��D�'��i��̈́b�m�Ω&��P��!�S��?�Q�[�RIA�  ^��Y¢��g�$	���?E���5U�4�d- �u����N��(���c$�P�c?2:�]��#K0Hh.�4���+}��Ab�x�K��?��Q��Z��Px��-�ذ�&g���9�%	3�B$��f,�=S�E��iI���T�ȓi���c�^X��P#V��O@hx�ȓ34��vM�2^(I� 	N�]��e��mMV�u��$]��r�E׬F~���7�|�KQBB�]�d@��h����%�>������(B2sY%c%�̌t-������y� Sp��A����{o�$���'b�'߀�j�#]��d�)I�t��I�'����s������U�[���Ñ��hO?���7E�M��Nl"`p����<{6!�D����LIe�ߣ+D�B�&`�V&�K���kp�E�F1�m*p�y��d�����F{�Oc�OI��#6*�`�b0��.Sn�� "O�%ʲR�2���K����wT��F"Op�jW`P�H�p1Ε�c7�J"O|1��c�<���C�1%�������'�ay2�N�K���9a��p� �	ʨOzb�$�OuxX�v��wbH!�����HK�'� a(�"B-M�����J������'_a&��#����`� c/��ط��xR�'��#��!�f�EZJS�`R�'Y(�틥�������<�$���'���A7��I�ȉ��&�"91�̱
�'�~p��O8K�hY����8�d�Z��d,�T*^�[@$�W� ���n�&E��y�lP�UBҽ(Ӫ�c�%��vT�'�ў"}��+^�iJ"�S�
�FI8&N�r�<� z"�LҺ7V��BI��~�x�"O�h��@�_13��[9�Ē`"Ot������"5z�`J�8b�w"O�:c"/�½@ T/3����"O���Q�0�V(��ϕ�g�X�D"O� ů�#c�8�m�[�P$�G8O�=E�4��v����ƀM���C��y�o@.�-r�ҥ\��)�U��?�H���O���YZn�r��-S
��#l�6C/�M�ȓ;f�u�ƨ�2i�+��	�;B�X��^�["��W�.�R2��Lh�ȓE|���]'i	R@r����6�^؅ȓ]"H���gL��2�΂)�����?! ����	c�@
��O�7�^���p�ء��jo(� 	N!X�D���:L�A$ N�,��y��K�`�(�ȓ5:h+6�ܵz�0��ȕ�N�~��U�̝HA����+]~�� %�!D��� m�C��M�Gb�Pp$ؤ#+D�찰�3��� 莃e2pj"n#D���5eђd�496J˽�=�s@%D���&�9cX�[��ħE�h�T�$D�D���پt���c���W�e�n$D�x���T�q�4{"(�/;�
�/D�@"CE�2D�4qMA u��-D������.�p[��B/���S�a,D�z�o�K_԰���c����f(D�h��e;$ 8��Z�pw�'D�x(A$�;�TI����>��y`�8D�����
R!X�Q"�&^5�d.7D�|�U���ra"�� �0V�X!W�(D�TJ�fAg��RG!�B�z,Ba�3D��A��s�r�񧩏&;����'D��0�?ߖ� �L�]�>���$D�|�&���x)�K�4�8���'D��(�.�']rJI��#�H�S�%D��'�9[
��CUg�.2�@"O%D�8j6�N�cڪ|P��C�b��m$D�����>߄�	&��#�HGB"D�$;��Ǭ$2Phr�<qk�f%T�ԫqB��x�p�C�ռ��ԋg"Op�9!��1����FH�I��,H"O�`R��5G3�HX1f�`�l�H"Oi	�h%8�ޘ*�EO���(�MP'�Xm�S�'y�]�h�i�쁫��ޣy=��
�'z�br�;lM�Q*�K�i�ZPa�'ΊtQW�Ÿ���bq����D=�'��<���޵{��0��H�P �'�����IӧS8�p��.x#�"�'���J���$P���Չ�i�2�Y
�'%��e�	SX���ӵi�,`	�'��<�b��<�T`�ٝk2�h��'�����+i��%3��g&�4@�'_���̓�}��yjs�=\.�U��'��q�F	N>8̣�h-�K�'L
���IN�XU͕�';
1��'6ހa���/�TPQ�T��
�'Q��XGD˞<Z�\&�6 ]l8h�'���3�N}`z�C�����'MR��W39�|`b
�.s�,�
�'�D��͜2�9c�ǈ�r.Zd�
�',��V+xfTC��ʺb�L��	�'��p�ݲL��-@�E�Rh.���'`����s=$ V�"q?0�2��� yQ�́�-G`e�!O�F��LZ�"O�"d�FR�PC��+K���"O�0�7*
�g9�tӀ�bP��r"Od�k��޽.�v�ۥ�\�E��ز�*O2AK�j�g\ y�k�Lp��'a����m	�j��u��E�>H��,�
�'F����R 
,���b �J�"���'h�Q�B��f�D8�	�
88�c�'y�2�jY�S�\�K��M7l���*
�'���p����=�c�
+g�80
�'z�͛Ň�N0��b��	U5�s
�'�s��C#�p�'�Y.B���@
�'��]�W ��2�U)3����'b���%��! %�16����' @��P�w	��Q*�?"���'��Q�"ؿO:���ƨ ㈥��'�P����@<`k�5���|�h�'�`�F��aH�!@�Y0px����'���24G��<��+���3O���'���k�kݱּ�J᠊�z9渪
�'��t2���ch���BF䈐��'�6!����%��H# 
՜!6� ��'dZ����SfD��w��M�H�	�'��M¦Ȅ����` pM� ��'\����[:�y�WB���b�'/l�@��<y�����i��!�'$�pP�5�9'm
��(�'�D�aM.*R�pIv����"�'����F�L���y���Y�'4�(�<|!$��d"V�F.x8�'�D5�b�,&�g�:2�}��'#�|Z3�U�P�X��ǽz����'�,�т`��)q�dO�p�Z�2�'(y���u��m��%�1jNZ5��'*� �r��9#�Y��̑o�#�'qxD�"��k�H����b�
���'ff��3��J,���劔Zc( b�';�1aaT836-�b�[.�<ĩ�'���&�UW3�X+Rɚ?v
���'��km=b�����e1v�j���'=��!�ʊ*!B�: �<��[�'�	Y"�Ww�d��0b*)�ո�'�~D*���u2��շ
���'�ZBZ"N��a����a M���fF�=�a��	D ����[�nƤ4�3"��J�$��dƥ@�b�R��(j&�q�ܿ@��X�[)�щ
�'ov��ī[8C�ػF�K�t�6�qڴ�zqCG(��I00����N�/���k�KQ��Ol���"��=$!�$�*�<�A`��-mg5�"h˩i�BiS/�����P2*�剥Oc��G+GϠ�'KB� i�I�V=V�I��(��9�ۓ2h���AX:e����*�Q� Ph�/	�Iy@��]�8�`�}L�d�3���1��qÓ+&8� `�;�����jQ6`2Q���5)8��&eD�dM�C�?M���E6,*&��ץ��[J-Sv����\�
�ԍ˧e<���B��#aC���`s� �IL&|9��?>dxQ�'
���C�(�S�Ç���pC� μkV �FT��ꖅ^=2�B!+�m�r�<�rU�6�"��r�O9m��t#�$� -eV]bS��.������ȶO��&%4�,ɸ��N�n��d;�h>U���5"qD��ň4f\Ԣd.�F���"��0&xyb�A>Lx�}��M�.EX��EL�M�&�($��+�Ԉ��0][�XᤌR@CFl�28�Z�?�n˂����*�J�� �%��OH���!�U% �L��i���Ĕ�m�8�E�Z�Y�J�a��BY���s�"ZƮ��U�@,=0ߓ�
�@�'��|��K�JI�/(U
P��br�d�l� ���²�����P�g�}��s@�-(,YZ�;fþ��w��u����Ad��1$�܄Ɠ=v0��١�|p@gY`C���0gÀ
��9R
Fr{��I��
y,� O�����$�Fl�Á��v��Y������I�B�(~qX)���?��U��a�+y~D0׈�V�? ��[�ĕ��I����b�d�P�FH?q�F\�a
�Y��	6E��K�Q��O$��Qe
�ڐj�9+n"UHP�-�D9)k,u�ĨCZXɑ&�)�x��"�����S ���+ģ��W'.PD㓑&��6-�u�l��w*�$��=�&��t�g��'<� h�P*NiD á�~�P�#� �3��t�F�ĀSA����U��Q�3'��2�Ε4�9��&4���Ù-, H����%��(���

5��� U�x*��*
�8x��8�#Y�/Z͗'�����BD�e��yIr!;a<HB����ŢT�'"1����W�vybq/�	����qB!:�%)G��N $;aH�-�<�OY�����0^�q���	�O4:m �%��x��$Y'mk�1O�,Ag��
n�����C�qX�KH�s�⭘�8��PA48�8	�I��Y̠L��"Ot���� ?Ԭ;���*n6�K��׮z��1�sAL�ft�&�B�`�җ���"�y�s��:2�і'Š�HgFO��yBLs�̑���^j+�@��%>1���H'��n��͙b
�iW��+Cl��r�¹��d �h((H:���;�xe��KT�cKa{r��[`���If�H��r��g�䉐���u��(��	.�x!�	�
z���$�:�ڭ�	�(�d܂�I�r�O<a����r&�;�n��W�рu�1�n^����#E� l�hT'G!��\*F�i�1��j�2��D��"̭B��؇e��vlBNrTe0pbܪ�(���Mnt��֦��CS֙�����!��^~��$D�9'�
m�bV-A��ѵY8@@��cn7o,~�B�۟�#=	s�1A�d0P��"�nxU�d؟X�D�)d�z�2S�3�Xam\�����P,0JRH��kX���j�T��(S�'��f�2AXV�.��r^�c�Ĝb2���T!�~��@V.9�<QJ����ȁ�^�<9�
�+o�T()RR/,��!���DXy�$�L���G�Z fD�F�$/TY�x=)�<�����Ő�y���,�&��{��0JUU��y�1���d�sϟR�Θ&?�X����%��͠�gԡ�"r�C3�\ДIHcpYp�U�x	���O$[��@�AV�;	�B���	�`�K!��ޟ)���	�@T(�����yz���'5���v[�L�8�
��|����	�'�t��4dۧ;Wb�M͌E>��P�y�G;��@q��&����"'��A��,�dC�>R �	`�c��s���93hޟ3��3%�;�	�Q>˓V� #�V,A�̏:��Նȓ��D����qt.��d��R�Tȅȓ|� EA�"ǩj���Ʀ 5V�9��P}�]��'E�4�0��8@��Ȅȓ:d������6 I��X�j\�-ڬ���^~M�A���q ��c�V =	 ����0��c�}���S&�)��`$ �*4��9[Lr%QT��NR����2e�pG����x5�ؘͦ���M�N ��/:�hp��>B��Fy2�N!L�JD��l��Q��Hz��>kvhp�bː,�y�*2P 4�⍷a���HB���v1+U�A2 ,�|�J�>E��'�R}�"�٪R�P� �P���3�'�̠9d�G%+R�� ��3Lթ�C�pL�R�� �z��d�`�`�����Jcd����4>��{�8f���oV�v �i�J-q�� 5�4���+[.�y�H�'� [�(ѥq�*�b�oI���'��1��ǐ� I*�E��M�>dt�� �c$6��sB��y��ݠL�@@��h���S�'��%�TኆwZ��'M�>�	�1��4�G)`)��#H
\�NB�i��b�k�l�ؑb]3G\��c�!�ORt�6M�#�!c��u��jA;(����JJ�4�nх�ɻ2���������^���ui���>�Z	��������2u�%c�$ٗ7�DE�?�҆)7|�!��)�'9m���!�]"Aw�}�Qʆ7!]JT��A�� �Qomb6���A��`6'۟?����|��9O`M��[��@t٧C�Ȩ�6"O M�!�2=�X�� �H!6�O���A����0>��/Z"PI��q#Ձ mZ��ay�<�g̶G�%(�`��,L̤�FH|�<� 6](Fm�!�J��*�vB���I+�2U8V�S>B��QbaW�M��AIv�O�D�zC䉶6��C����F��UPD썠W~m�!C
��h$�"~ΓfH�Y�l̿��y���?hu���ȓ)M��B��/V����5xL����,E���ZŁэ�a{��+Pe*=�D��n���wkK���=Q����~���Y��n���X��`����`{���{�!�x�������O��[5�Ϡ /�O��!�`0�����)؏H� � P*�P�΁´�D8b!��M��h���H�,Τ�ՏܗCD�I`�5^����O��}��?Ĥ��E�i)�t���J�8���7zb,�Ӂ�gFL툃:���I"8����:�a{R��r4���;��U(�m���=��	^�7Ѣ�!�mӀ,8�oӥl$��R��ڜyb��*�"O�i3��+>�0�F�dg� �A�Č�b?�:����H�: ���9�Ց���o0pK�"O�8����Bd�աۘxX�����[��u�*���S��y���4{�Dh�6)�#Z�1kB���y�nئY�#TL"9�9�A�>�~rH��[bm��	$uD5�U��^ ���º'�B䉁f�Nm���6 a�}x5�#V�jB�Ʌ�����T= �� 8tgL��rB䉺���Sa��T���!��B�I�h��+���>|r1�
�#K8C�T�8���  k�(�i� #4:C��#)S���p�����*�M�9<Q�B�ɪN�ƅ�$e��I�Hx��$bB��w����ANI:/�D��gg��TC�I� �˰h@�$mTY�w��G�C�Ƀj�܃F4@*�:�E�5:C�I7!<H�#X���V ��v��*F�4D��s�H�4 -^5���� y [D/,D��;�8C0iCv�Z7,Q�CL+D�T��O%bRt�DK=r��ԢS�)D�гfPK�<��)�+��Щ#)D��Tgˎ^���
�E���x�ᴧ(D�Ĳ�&��Rk���Âw��;�  D���4��{�2����!zH�� ��!D���D]U	|�p�߼_�\�"D�dx�I���1`�,]5?���Fj!D��2�n)`�4`���yA҄��G0D����/D.�@�4j��^,B�K�*/D�P0�-�bx�LYEH\�0�*O<m Ӊ]�A$P��"�h�3�"O���_�/	�xR
@�Jv"O�a�G6*��h6�ϴp����f"Ox	JV���_}l�G���B���P"O���Aƃh��P�$�P�/�$��"Ob��"O5b�zh�6�W9+�.:T"O"�be��"�^l��
�k�L��c"O��z���<�0�Wc�O��L�"O���G"�:,�@�J�B�(��"O��i��ٕ1���P��� ���"O^�"h�0�̹�󅋾8�ܳ6"O>���#����B�͛̌\��"O����H��9iR�(
o��"O��%�[�:\�E!U����"O�p��	Y�9�S�M��E�0"O{^�8�6�W'~����pj�*V�!�䉓L��h�rχ� ֤��eU�!�$M�?:^�t$�P��My��֘N�!�$ύ���`6��k��=�@�!�$_::2d!V(��4��mӢ��0]�!�d2m�b��26����A��P!�� �t�̓��X�.��0�T��"Oސ�t��~*X��f-��7�����"O� c�m��<5�<H����Z���s"O�9#�KB�t�\�5N��9̈D� "O���K�6x�����#.�N��"Op��$(�kBbm+P�¡T��| "O��)fN_�ր`#���Z �,�E"On9���E�O��d�cŲ\�@��"OȘҰ�&F�(B������´"O����̃M[��z��74�"�ʵ"O�)@��/���B�A�f���W"Oxl��H���-4Qv�z"O��	#'�!c?��+Zhx��"O����o��
��5ӖH�?m�8�T"O������(h���b�JI)h�"O*B�Lݙ;^1#6�9M\p��'8�5�� j��%��������'/~�ǂѿK$.��2�nb�2�'�D���G�N�z��N������'�z�AR�ͻ� y�1�T2m��'z��%��&�\���כ���r�'����!+�8{��H��q���'n�Q����hʜ��c�&]�`��
�'���b�-(��L��'Dd;L��	�' ^	 ���o���"`]	μ�I	�'J����I?�9���6��X��'q��3�,�,%:�Q��Q�pT�
�'��ȵLà0��8"ȇ�a�
�'!.�ˤ���qc���Dԫe�fM�	�'�\���E���ޠ�����Y���'�p��֬_�a�z���ĉ�)pj��
�'�P*�h�;��M��j�� ����'�٢D
zJI�.�<�
�'֖0S�$־ d`��.���'r�)�(]2"m'�y> l��'�V��Q@n�z�ӝ����'���b�F��(�02D	����'Q�|2EmU,|�~�xRň.he����'��L	GgW,b��#8N�E�	�'�6YT��?9��`�2�2	�'@B����3F�P�J��7u,=��'�����(DI{ץG��t��'Drx�%gN�Y�����eɷ�)�'��@�g�J10��E�U&hM\���'���3�*���s��6o�H���'*��(G@I��0��&ܗ_)�\�
�'+�]�F��Ecn@1�$H�FO�5��'���dΝG�p�[�4o�Б!O���DV=h܎���.7Pq�m�a��B�x������<X�Vd���ϔ$H2��Ic��*D)�-}��DA
�'���D�M�u��P�Q ��LߒѠ���V-s<*�@���"1�tb>u�0dMq�����=P@8��6D� 16��5!@�u14�έ0WdxjC�O�L#��Fi��:3�<E�td�!r"H�$��Q{婧�2\���Z�u��qP���23�X�J5����P������M�)�P��$�z�(��I��h+�n�s�}��˔���'!C~�.�2P��r�J�b ���-i��Ot�@e��Z"�*�e+��%��ɸ0t9��@u�
�!f�����T�3j�0�(xå͐?�C�I� �޹�wƚ6G� �u�!.T����zo�A#����[a��`�T���O��*S��Bz �Y��H�%%	�|�ց�#����?��@�7�H��'��P �Z
9|��Tk�5jw�	Y¬Qw����]�H�@��O��H�F��-�����M?S����A#�n�v�ʱOH�f�#��[_>\�oG�o 4�i� ��sh�`Ԇ�8 �
T�&�ÞB�"`܄�)� `�K��ۦlB($q�\G����"�O2u#�a�m�(����c��-��-�6 �0�6J�^a9&�Ok�,P�+ �`)���
�GL�8+�'ʪ�9�Œ-��s�a����+�L�0�R$���dNIrpo��Gƾ��;���xI�λ}��x	���eG���n�
�ȑ����p#�QK#e[7\8+����`��z��8cŁ3$���a�X����-�=Y��$f�lA�e�ٙb�Q��/Ȇ!�Q�hBn��d�xq���e�a�o	#��	�.B"�&P�i���Y
$@�4C&��bC5�X���؏z�h�D��?M�dr#�>(G���',�CҎԃth��6�����x��ӦG>���_�"��P(Q�`��M�3`�,�\;�y��1�4�HE��)�|����T�{�Hp�
�V��t�b(���Nթ��1�>�p-O ���Ġ2���dxܑ�C���U�*LIu�#|O�hkU�C�Q�0�\r�"��8c�A��D>i a�j�+�F��>M��4A���BG�		'��l3�R��˱��-U����Պ�;B���Ě6�bW�Ђ^����'A�$PA�I)Cl�]�T����Dt��S0�c�U�t͛��@#�,u�X�|H�k�'P�}xq�N1V7��J�w5�E��FQ,n����P��>�8�'mr]��ņ����y�`�C�Hw�ֆ<RlD�K�$�����Ε���%��O�lCE�ʁ����F�]�	4���'&н�0 �8d��\;�� �x��aw��2,�T�`��F�\P���s-y��'�ZQB4HݙJ� �� Jם*�n��B%�� ����(��5�X���T/8R��(p1��lB��SPl�P!�0D��C"O,�B�ex�y�ÊtR2ى�A�".n�{�ٓ2(�G��
$ ��9�,I�'-P04z%E�E5-&=��"O�Ոs�V�� r�(�i�AK%���;�j�;�L!��|�P��Q��	>ғs����
�w]��yRa�'^i���+�iI��Μ9�|�"��z�
�q��=���)0ϵ.f��K/pm�\ �R�`Ԓ�JU�Fz�џ�!A�8N��a+�j���S�`.�13�E6��58t)/6�B��+k�q��kM�B]XA�F�<)�ZgS�\�!��2��#���"B�� .3W��UEEQ�<)t 9iI %A��� 3HQ0���D�����O�� jB NU���qO@���Y�a�@P�� iVd*�OB��#F�/^X�u �>V ��`�l�0@�h<�"��\X������ã�C�Z
$��V;J��$�/`1��X3��m-��;�L�)q�X���E�*K�4��ȓ%��]K�ƅw��dc�B��x�<D�ܙ@��pP����T/�D�ǆ�)�X�I"h!��
�tb�*�%P�r������UF��Y7�dS*�(��I8sR��9�V(1V邳�H1a>DB�ɍ9Pdx��ƕ�7e��;F)�N�4B�		N����H�فE0�6B�	����H�.�1A�a�_�W�B�	<U��dkvL�_CL1��Zm��C�ɩ��HS6�ؤ-���[Ac�B��C�$"f�]�r��E��z�-�N�C�ɴI�~в�ǡ���#�e�&;6xB�/K�h��a.J�t���:EE�W��C�	�_��H�¾�R��7����<�+��^��#~�В!�V��鏢&ZRhAu�r�<9Uj��b$�Ux�D��<�r���-S�~�����S��yR*3}5}cWN��@&x=@����yb�V7�����!T=�N�)E�_�?y��٪L]��4lO��t��&�R5�@c�</>�����'6�гB���oZ4����c��5# ��a��Rr:B�I7jZn����ڰ�Sˀ���8�уhؠ��S�v�B��#���ag�(y�B䉃X��Aa�C�*X�āC�C#w�-����<6P�J��G��'��}Y� �`�����5zL��'D�pnc����8BW2p��6�p0��f}�|��$�M�����dU&
��@B"�@�{BM .&xHt�Ԧ�9v.�cӢ���D�4C�M@�l!D�<"dㄟ#�x3��7>�%I�2���%L�HB4�>F�>e��T�As4���HL���y��N2D��r�A0@���	���z��0�� �+�+��\�)��<� ��!�˥/�����%h�q86"O�RjD Tv +&ӦzVT)�O �ʐCر�0>��j�i"H����� Y� ��X�<��˅6=6��q@�' �R�[ �T�<A�i�2 ��a��� iq0�`�Ek�'`^�R�)�r�O��`�6UXZ� ׎
�:����5D� �Ɛ	%r��ui;F�`BW�� #ub�b�i�)��<�b��s��=Y�+�.�M��&�_�<C��<�8�qa �` hˏ��T�#*@2� ��'q��{���'Di޵r���&)1
�����` � u�6�s �A��bHlE�O�co!�S)Oh�q�Ɖ�T�p˕T+1E�O��R�&	�T�ޘ��I�=F3��[�f�pB��)dχ6 !���+@�ڡ��	�(��5oڧ$r��w�E�]��O�}�"
q�1͖^>�#���>�
��ȓ'���(�2$�Ĝ��S�fN���I0V�#"8_3a{���6p���0!_2]՘E[v�ٝ��=�MY�`M��9��r�r�� BϾd��k�j�)��)� "O�b�[#_�0$��ՎY��P�s����{ 1h��7�H�X�Z�b� 9���2
t��"O¼�LJ$n)��@��ޤS�mѠL�(ĮP¶b+��s���EK�t.`���W���k�B)D�(\�m�4�`7 Y�nc��ẟhK���� �a|�lX�sT��6nP�&pbR/Ĺ�y�䋜8�`bT/Z�O�h|�q�y��6�~��d(�p��	�y�,��"�v;�Z�7��]&W)�yrn�8���Yk�? �z��㔶�y�Ő�3G�@��+$p�@�7	�6�yB	�b͆a�1�\ 3��B�W>�ybdȞ=t���Ȅ=j�n��"mL �y§Ҿ?�P����	�1i<JI���yB�+%��b��*�2ak�N�%�yb`ȧ������#��s3�]��y���^���ƒH� ��D�y�O�:Y�-��bN�͚����7�y�J7�xu�G ;	�\�NZ��yb�LiC������:ܩ�g��y�ִ3���u��xB�y���6�yr(Y�b�,s'����*
2�y,Z2di���e�>z��9:��D�y���6k���ؕM*��` )	�y���"��1�6/��@	����
�y��zS�`f��*�8-ʐ`ݴ�y�+��̸a8E$�5-���� I5�y�*A{���2�V
&8@���@�y���*8̺D�`''�Vъ�g��yB�2b*�ف���d:hSwj
��y��61�� B�6��.��y�
T���V��q/�E;_p�B�'�hJ��T� /I�Q[',VB䉁ZK� ���D���a�Z3�r%�E�ͱP��DT� ��\�Q�&�i�"M��"�!�d#|Z |�4*/n���"�!/!�DQ�&������+v�%q�A�=)!��0;E"c�	LjJ��3 N�Z&!�	5z�>�K�'O=L�U�����!�]�9D��#ݑ'/��fO< �!��Z%T�"��� >\S-��Z�!���ykw)�K��M ���0t��cJ$}Rn�b���Ԉ�?i��I ;��@��g��]��


f�I=�(xO�z���x��OK�A��B2[�
t���?T�~�д�_z. �5� �l���K�:O�>)��	w�Z���D[7|ժ�s%�H>S6�x��E�lO�q�G�Z��M�wʃF>!�f�+A��0ѥ��?hl�fnV�rit��J��M��!A��Ɇ�3� 6!wF�A��T���Y,z��ʷO��rf&t�	Y���ɲ�I)|���;�'xȢ�pA;%Ǧ��U�UNR�i��<O��SbLZ�X�\Q�4�F�OPB��q��0�XP��\6��D�ۉ��u�ʅem<��EAÈ�?E�ܴ{>tE奙�(���1��o)���c�Q_�M#�����	u�L>���4u,Ɋ�͋	7�$��Q
�	&� ��G���0h`������g�$l�ȓU�l�Ȧ�D��嫂�+>h������&��O  �L�=����]ud�-)���8e\�Pw��ʲ 'D�H��T�/7�ɘЅY>j������:D�pz���7K4Ւt�[�]c<Aѥ7D���������D8vĤ����?D��SA͗�Pp*0mz���'(D�� ����m�a,�Jh��!D��#�%"���9a�o�L:��>D��3AM�[K��1�	Řwx@�w�<D��P��\=:��°�z}�D�-D�12M�b�@-I�A�V4��C��&D���@�4�ܕ��_��J��W�>D�����-B˜]s���'U��y�O0D���F.�	q��P5č*:��%�H0D����pMr&+Ѩ{��Y�A�/D�$y��K�t@��2PIJ+v�`sM1D�h���]7~�"���d�eP�u�/D��`�ʆ�<��d��0ߪ��1D����k��ܨ'�Y�;p�h��':D����)�"Q�zaC1�K,
I�ѡ6D����ڢ����#�ĝlD�`Š:D�|��&d��ģH*���q�#D��!!�=���+&d�*zˤ�{$#D��⑮Xsޚ �[�n����R!6D���Ƭ��('fx��@0��r�>D�� /��t��l��g�
n�	�#�/D��x􀐹v��y��*#K��!���,D��#&K�H�� ���Ȳ�)�&D��p��[�4`�@�Ʃ�1'�����?D��ԡ�x
�Ycl\�VCĥӐ@*D��(�F���ڔ f������(D�|�%��8x`���»:q��U�!D���q-J�F��eƁ)���� D����a\�j�����V�i�̊�<D��h5 ��=�4!��OхJ��P��	/D�\��5F�x����(<s||{t�+D�8i�I	b��PB0�B�	�$!4�/D�x�Qұ[���[�ܘ:26�3�a.D��
�@O=g(T�(/����>#B�	�.�X�i�Ǧᒓo�B��<9��
g�GNr����NP�^� C�ɟ;Kxࠇ-X��������N�2C䉢;nP�0v,�|.�8��6� C�	W���L�@
�聒陫K��B��ܕ2ER�x��)�Ǔ�J{V\��'0�����X�0J��G8Z��h�'�f�Q�E�Y_� p�ϋcU[�'_�8�deәSX�����p�T@�'<|�3���|LJ6g����]�'��@HYD!�]8�E�t^���'� ܸ�c�;���
J9I	�'\�O�nƴ� ��Μ�
��':$�����F�"���48��'�J��-9沴���ؒW�����'<����@l����gJͽV��1	�'�>�鳅��n;���^�]�k�'e��1Ѓ1n�`8�j�b������ ������0`����Ϳ},9�"Obm����)M�1#�ܩY&p��"OBл���}��y�-��F�x��"O@�4�Ξ*o����V�i�&��f"OJP��)5�Y�A+��*"0s�"O���5�]�t�X�� �$P�"Or�1#��4Y	��ƅ�h���"O���!eH�\�m�����^��t"Oօ g.^ O��Bf��s���0�"O�0FI� J��"��j$Q�"OP��eEáY�^�W,�_(�"OBe*���W��̂��_0#q�;B"Oa�#�+���@�D�>hHԸ�"O*����H6�t��ӂ&^v�"O�Y:4�	�l}\̩��A�\��4�	�'�d��vɐ�%�@�U������'�К�OF���]iE ��}�X0��'�H${��E� �։�t�DD`����'��YS�� |�Qa'HєB�X�'w2T�$K�K�t�ٷ-$.{
]��'1�x4d��Z�L� dU*�͐�'��tu,�?"�`�OV�I��'
��㑋	%���#��׮	Ծ�0�'T�����Z>Mn(	R≓��ͨ�'�ZТ7���7�ЊffGxQ�=��'C�L;q�T�uP�B�Aښm��I"�'|6yiv��>np.Qc��_s�,
�'�}צ�sbd�H�ᗄ^��dq
�'C� y�A��k����q�G�&fr� 
�'\P�pQE�&v�~}��K�-�ĺ�'���a퐺Zr�=9�<��
�' l*D�96��� L�K�!k
�'5
{�K��A�N�ʠ�@�J�`� 	�'S�e�5��`�Ҳ�ЬH4N�C�'�v9�Ǹ��lR�NT>���'z����-�ڰ���جJH�q�'���g�=#��%ƜB�Y�'s���`��&�����#7*��A�
�'�D\hG*�;5&�q0�*�;VD�
�'��s&� �2��{�SX�@
�'��;b*�0m���� b?/l@!
�'<� �%lб'Ɣ�Wb�F�X�y
�')a��d��u.l�f�g��Y	�'r���fЭf���P��8`��'���2&O�4i�:4�E�O�)%���
�'<I�C��
���DØ�!s��R
�'%����ͅ6x�+������	�'��ݠD�7>�p��l��	t�1
�'��@��O̠
��*~���:	�'U��At��z:�M�"íG��Q��'�R�;aA�5P{�<�F�B���:�'�\�$N��M5j�3�]5��'���Q��P*������?70��
�'�ڌQw Q�BX	S6A	>a��d��'�P�b���&�����BH^H�c�'�vE�Uٵr<�DHBI]�Np��'���y�Lk���1'V#�x9�'/x�9�D%U��ZAX	PB@�'�F�ڦ&Ę=5Ь�᠞�p�����'4LQ�@�)��)�1��/��Eq�'�~h��&[;M9 ��g��t��	�'��<{S,z���%�̈́�\	�'���bD
N�	���JuC� |$���'*�kG�П�L�!U��&T��[��� <���E�1���	�34O�T��"OD��� ��"�a���h��i�c"O��z&�ً2���q��94��J�"O �E��5 �p`C�P��Is"OPh�UdZ�IW0����	uo>�Y�"On�+6b�270����[�5
�"O6�Є��d��H��8Xl̄3c"O0�{G
�s]tPkQH�@S���!"O�H��ɸ3��µ��	I���5"O+𬙧Y���S�d3�"�"O|	�S�L�.郆]b�{@"O9oL!c� �V�D>���"O4$(��Y�1	�b�MJaq"OT�R�����R�� =|��y�0"O�=��Y�!B|	�dS�#~�H��"O��G��b�|Y $��4Z��9�"OH����X��t#�3e"Tag"O��xQ�UWJ����#:��i��"O��� �x�D*~︹��"O\鹃��/.�ĺb�E�U��p��"O
�����o�w�^��%�+D�PqVJ21$�M�&ON�N����%D��XB��)z��� QF_0P"�#�'D��B�e�,4.��v�޷x��4Ag�$D��Rs�O� ��u�d��L�����>D� єc�8<�j% %G�HB��f.<D�@�烍gdL��fm
9E���I6D��j��ų)�J�i>v�I�� D��g�V�`��pI�dg1F�t�>D�LpE���`Z=�g��2�(]�d?D���Q]0Qx�|𷎛�1��r@�>D��;R��$C�
WN���Vʕ:�yO1S2�p@�J��TjF��=�yҮ�+!�fT�� F�D��e���y�$˥i*)i3�<HHd���y�ˋr��D
�79�:�l��y��_0f��Yx6�^'"��!e���y҆܇-��H�ɂ 6�p#7�M�y��̈hy���K
�B�xC�!�y"�ۚ-,P���NXM�Ty!�8�y�M�3,`�!F�\�M��x�s@��y� +�e�ԋ�RG���O	��y�#7�(����0L����eK4�y���0��jC4E��9xp�]��y�ʛ-R�9��ó	j�����&�yR�@'*��2*�K0t#����yңA��
�a�������I!�Q�y��ˊ4�N=�&�Æ48Q���y���C�A���щ��yR��mȨ���B�9�"������y2&�'J�h'aB�'�HS�>�y�*^QjℌN1mK� ��yB�$��#�I��=���PE��y����b�(I�l�KJ���@�I2�yBeށ`�h����΁�����ׯ�y�IH� i�Ο���$`�.�+�yr�M	db\�,����7�^��y�썲��hr��\b����y�ǖK1�(���H�<��F�ێ�y�� -�,\P�(�f�ӖȜ��yr�P�?b���TF�%(ż�Q��iH�Q��Rg��I��䗠0Z���e%�܁�.���!�O�{�4m��j3,STB h����EϜw����S�? �a���r�RP)^&�8@"O`LQ��רih��sURs�"O�p�F�S�2תA����5;��k"OF�8��ϲ2�p�iU�L'wFA��"O��p���>)t,B�k@�]+���"O�a��5�f�b�
�;���"O��o�;��L����i��-�u"O�A��9̤��� 3"rPy�"O���S�K+r�Ta
�a�4CIA"Op���B4
P6z$�Շ"��eI6"OT�S�'�9zp�j��6Oa
i� "Oz�w�OoL�A�̟6��p��"Oxqj��> �Ir��l� 8��"O� �����b#�ܛ� %"O�ሆ�"�(���o�
ai$"O`x1B��D���P��6lZ`���"O���"B��~U�)�cC��Ii��6"O�j%
   ��   �  l  �    �*  �5  _A  YM  �X  d  �m  mt  �}  F�  ��  ؒ  "�  e�  ��  �  ��  �  =�  ��  �  _�  ��  ��  )�  ��  j�  
�  [�  + � � n  �( 0 U6 �< 3B  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy��'���^8�'HZ�L@t{v��Y�!���m��h�U��{B����M��>�џ F�$�3mJBd"`����:��V�y���%vd0�U{N���c�҈O����N���1��3~�\�QWM�l�<Ia��V�8�a�KŮ8�B�gK�d���=�҈�!U����@ޔ#	�a��Qhx��'ʴ���W�Bg����(�vD�d��/D�@c��уo�0܈�`ʺh��E��"O�7M;�-,����.J��%K̰F�Ʉ�t������;kX���N/Mc�E�u��8�S�O�(���,Ui�"չ*���'��4�B�'4v����[�&u����'Px�+��Qe�I+��O�T�`I�K<��O�c�b?my@A�R�)���E� j�KQ�+D���!��pF(���$_�3��
�`.��C�&3lXG|BV�@ZF$ߕ1F�)�fA�Xt �(�,.�����{�B��c�	Fik@�)Z�l��Ɠ&D(���L�j,�p�6"$p`Dx2�|��)E:�A�'M���H�n�)�!�� �3VdL-0����Mִ6>`��f�|��)�ӾBA��S�ل��7�� >M��'a}���H����h_1V�Q1f��y�dޯ<y�Lj��C�82��+W��y��νf�z�����@x�"��O�"�c	V�f��TB���`�~��6J�x�<!re��t�0��LC#J� ��ʂ|�<� _kl~�B�L[��"����{�''xF�D��V����,�/xrL;P�]��y2��/��\�b�?#��(�$���y❟P&����7�$5�K��,itH��&PņȓW��E(bw�h�&D߽k����ȓ}�J$��
(f�Y��NR9��d��1�`� @�]����B�E�x}��c��:4��B�*��$g�,B1���0,O��	Y��,�(����n1>0;��P�=��B�I�_&�`��E����FMλ�˓�hOQ>�I`� {����H� *H�#w�0D� 1d±'qX�s�ݔGs�p��P��HO?牡a�\�s EM
S.rpB���'�����)}�I]�~e����%���z�ϔ��MS�'ya~2��d���Ɂ�Z�r�(H�#����p?Y�OpP��O̔r��ࠥD��l��"OZ��� 
�z��4Y�k�UG�����	\�O��LX�MBF�$U�E �$%xl��'2l���Z#\/$�u�Q�zqj�'" hcT�Bn�4b�*9�	�'���Y��ǡP145ڳ/԰AR���'�6�#m7sv�Y���q�T1Q�'�8�;��
4N�(���زle��P
�'� auE��HP\��4�X���)�'�*}�c-N0H����3W�}�B0��'�aA�E�%
�lI#(NL�l���'6�j������KU5C�~�X�'���	� ;K&X2��-�U2
�'���6�	�@:l���Ɣ6k�
�'K6bT�=iqx�����2�'�H�����%���k�ǌ�ѴM��'9��:

34&�؄Gւz4���'��|�PI�ؘ`$�%p����
�'԰	
W��6�1d+B/4`�Z
�'����"�đa>���SƁ�g���	�'�LC��"r�6}�BK	sy�
�'�حe�Y'y5��[�)\:��	�'�&I�Sˉ5�0�Q�ٱ���J�'�\ԩf��T3�C҆�5
P
�'�FEpơ�de��	%*�0�B0��'?��S�:,p
�ZT��2*9��'��=x�#S�(��*b�x�
�'?�h�Dh�d4��cM��7"O��Ƈ��[,P��P�Q�|$���"O�yt� 4,��s�P�Qb��8�"Ov H��B�U&8��"_�2I��1"O`��I��N=��@�*1,��2"O䱹��ʙq���p�o�.`D6I3s"O���w"�u��:Ί%dpB""O�Yh���7>⌻���w콻�"ON��D�:M%��sթ��8.9��"O�ɱ�ː$W�� �S�L���:�"O��3��a�jXn��=���"O��a�ܷ}J�0���K<b2�i"5"O"�b����b��
c@�À"O�@��˽>�=9��3��8u"O:dk�Oˍ_ņ�C��L�ƌ��"O� ⠲�уr��a#׷Ԭ��"O��;3 ��T]F�� �#f���K"O��qD^�2��(��Y����"O����W#44�%��B �X���y�"Oh��l�D��cDIҔB�"�i7�'�b�'���'R�'s��'���'���6�{��85n�S��%���'�B�'�B�'V��'���'�b�'�V�z	-74�H�ƩV�l�`�ä�'���'���'��'��'���'����L�#n�F�u�>�>����'��'w�'FR�'��'�B�'�4�z@��CG���r���H�˵�'~��',��'wR�'��'��'p�ؑ��µw@,�(�B��H�6M���'��'s��'�b�'R�'�R�'u0�+�'�`���2��.K2����'*��'b�'5��'�R�'���'_��Z�/�@�di�S�$Y/�Q ��'���'eb�'�B�'�b�'��'��� g/����ن�޷g�aXV�'���':��'#�'2r�'c��'Z��L Oņ.>B�#�Y1�?���?���?��?���?���?�6K#+/��#���}8I�Cc�?I���?	���?)��?���?���?9��ک]QE2�8rǄ��F7�?!���?���?����?���?Y��?Q�-�T�x�D�J�i��� �ѷ�?����?��?���?�Sh���'\R!K)cP�i�rHP�3�b1s��ʁ-[�ʓ�?�-O1��Ʉ�M#0��̢�`�K�!N
Jo��'\�6�0�i>�	��4�5H��n�@c�Ӡ���@@Cӟ��ɕ$x�na~b6���a��ë%(���$h~H`U�L1OJ�$�<���N8za�٣��^�h�4c�8qz�n�"~b���r���yGK?OĪ�{�n���(?q�P�	័����	��+��6w�8��B�x�bc��-��-i�tϓ6g�Ok�����'ժ�Щͦ���;f�-dPѠ�'��	X򉵞M�1 �A�*�@���'*Y� uY��S�8 ��"��>���?�'����^�l%�E6��,�5	B�!���?Q���'C���|R���O��8�`�P�C�V�``� �K%p_6�.O�˓�?E��'�f�c�EC(>���@�֠I.2��'�6-F��I��M���O�dS礉

Y��a�K�>C��y0�'��'�"��^śV����'j��M�)�`�6�"'|���Ay��&�Д��D�',��'^��'�Q�bD4J �*@�?4VZT� �ڴPv�����?����䧣?�a��_�b�ءC��e��I��0J�ɶ�M[Q�'މ��O.H%�W#�=y�A�L�c�*BU(%�R�S��!��H�V�b/^�Iwy�h�A[�0w�փ|��ATH�r�'�B�'�ON��M�0B��?��.؀٘1`�F�⡰U��!�?�B�i8�O`�'-�7���qٴm�jX�'��5\��S
�4�> �0����M��O�H�ؽ�����wz\Ţp�L�#pV�ꖤ6�`P�'��'s��'@��'J�H�x�G��`C�([P�A�O��X���O��$�O��nZ����'(�7�(�d�$����%��-.�`���� 5�v�&�@��48���Op ����iU�	,X�Au�Ň^b.��7���w����n�U���]��Uy�OeB�'@�"��B@sTZ�'�y��xr�'b�I1�M�g
��?!���?,���	r��{�6���"�2�DU�Ҕ�8[�O�\o��M���xʟTА���
�Dh��T�sE�*��7?����T�l@�i>9��'̀�&� j�jڅ<;(��3��]Tdh�����(��ٟt��џb>�'��6��>���Nаw�諥a�
"��-�s��O�$�����?a�_��Qܴ$HVk�e�B��,�tΛ�88K��ii�6��5866?i���M����,��g7D8b7�׬2�ك��yT���I�t�I՟���ɟ��O���U��lL
$��Ѿ�
�p��kӪ�����O����O
�����Rʦ睪i{��Q�C�0j�h��0$��޴}��#��	�!z�6�i�X�W$X@�����e�E��m�fl�$ d��[T"˟V�	]y�O�b'�|$8ѷ-ԔF�<a��f�*AR�'�"�']���M��#�?����?I�*L�x4�Q�~D�*�����'p���?y����A�1]�A`�JU��P��B~�
�>-��{�9�O=���I;j
B��!��Љ�E<;������� _"r�'�r�'^R��̟Xb����MSTb��~�ʤ��	��(ڴA��(���?�i��O�� �͑��- Sٲ7�J	,��I�M�"�i��7��L7M$?�u�Q�H�I}ݱxC�_Is������#IL8#��%�d�<�'�?��?���?Y拎�n��ז� �ЩKd�ʂg�˓?
�d]�Vb�'����'�� 	�& ��[L@��1	����?��aI���Ozj�p#H�u��K�ɔ<Rk^�ؐ�¦o��8��Oм��	�?	Dc3���<�f�>Fs�I�e��0+��PA���?����?���?�'���ɑ f����{C�U�RQzg�>ROhe�� ��49�4��'V듍?��zN��-�7E^�� ʒSB	 ��ŷvY&�
'�i��	���1ۖ�O�q���� :$�"���b82�(Z�K��`�#=O �$�O"���O���<�|�5��:^#:��A���A��\���$�O�a�IA ��OP�mr�Ʉ73Y�����3PN,UY\pK<�s�i0V7=����Q�r�l�o&�?���*fe��]���V=nC0��+����4���D�O����]nm���  ��;b��l�*���O�����M.���'A�U>Ź���x�x���'f5bH�<?�A_���I��p�O<�OM�tk�,Mlw��t�,y��P��K�V���2�����4� %��@�O����$�s'&���bR��VA��O����O*��O1�X˓	&�&�**x������4����&�2Y�����'[Ҧ|����H�O� n�%4�>����'/��P���ϛ��YP۴T��#��5���������!-���~��!9(����d�R�YP�_�<�+O<�D�O��$�O����Ob�'=�PUT��&�M�� K4`� �1�i0�����'�B�'x�O�҃i��/x�8U�Z6.0�
&G�  �I�y�N>%?ɺ&L��)�|�����6p������`^�m̓lji����O�N>�/O�I�O���٧G�����h8g��O���O����<���i(z�H�'"�'Q������{�)K/�w��|y ��[}��'OB�|�K�T�>dH���`���+�b�����:E��]A��ՂpZ1��Yi��uZ����15#��� �ǟu�*]��A�2����O��O��8ڧ�?9D5g�x��� &  P�N
��?i��i��1ɤ�'�"o����M�b\A�d��l"�є�S�K�������	ٟ�P�%�ɦ��'f4e�����?}��
��)g���A�D��;5��H��'��i>%��ϟ��	Ο�ɻ=9� ;�M j蜠7gҸ}��T�' 6�Q������O��$'�9O����ǁ7A����� ޡ { Y� ��F}��'1��"��).5jġ�W�5��s�ýbj�v��x���{yĀ&�'�4�&���'��8��R������y
�(��'~��'u����U���۴���F�ꁙ��0$g*�����7<b�Γv4���F}2�'�R�}�r��V�A���7rRv�#l"@�8��`Ӯ���1���j����w2$�E��q�X���b�k���ʚ'�"�'��'��'����'M���4x2�N6@d�Ǆ�O���Or$n��.���'1B6�'��9A�pkD�U:�!X":�1��<��禉���|b5%)�M��O��d֒
dl�r��Ϛh
���Gj��!0P=��Mx��OT��|z��?���]�(��m�s��#�dR)Y����?�(O�Mo��q,��ǟ���l�����t�@�p/X|��M���$p}�q�To�7��S�$�Ò^��ǌה\rJ���V�>���n<�x1�O���'�?�bf.��ЈKUjm��;j��lki�w>��O��d�OL��	�<q6�iSv=�vf��(�nXc,և�ză3���ldr�'�:7M>�	���d���5{1/�,a]���rP&xbI��M��i4*�w�i���/`�h���OD�m�4 ɥj�"_�7��;���̓��D�O`���ON�D�O���|�v�r���Q�Ɖ,/h�HdFܖO'�F�>���'������'ܔ6=�l��m�Wޔ���JEU��!�C���M��4!����OĬ{v�i��JCp\�2���m�<����� zf�d�*)�>���r[*�O8��|�����BpG^� <ʂ%�'w
�)���?��?�*O�l�0N��I՟��I!��;���O"<�dT,w��?�@W� ����	L<1��/��	C��%v�>��N\~"��K���c��טO����i�t�'�d�i���w�@t�Ι<��BP�'��'���'��>��I�SN4l��=#��+��
S|��I3�M��g���ɦ�?�;`z����6ud8f'����?i�dw�f͂8�����,�3��@e�$��C�P�G8~D��Q���%�H�����'�b�'X��'g`�SA��l�*=h�eۍJ�p%*�W� *�4{��Pj,O0�d9���OP}��^����Z��L� !"ѣ�l}��'v�)1��i��l�׫^�8�${ l�.s��)Al�~b�	�@�#�'���'�X�'8|�f"����rR�˞.`��'��'E����P�<pشj�֍��^�X��c����t�P$c�t��r�v�$VL}��'(��'�����`tÑh�; �3�ɏN��f��4�'q����)���	볮K f�Ƭ¶éT��s�<O��D�O�$�O����O��?	�T�QW$��30IW7����[���������ٴ�bu,O^�l�\�IBh"�h��� /J��z�2B~%1L<AѴiK7=��j�x�*�"��E��Z$3b��R�ŕ�
$`p ���,,�����䓭�4���d�O2�$�x`����G�!P�(�AfC�
�V���O�˓(5��	Z�0��'y�Q>�(�FZ�9b����^>d�RyC�k2?��Z����٦��K>�O�Z�
���DaA�Z�}�Zy0D���P9�hh1����4�B��,�`�Oր� D�0��+���"�TX��O4���O6���O1�J˓p�V��X����!�͝����Q�W�I]�(��'��m~�f�4�.O�6�W�@���l�Q)�)�6� �m��M#%i� �M��OV�
���K?� NjC`�z�����Ԇ7 ���5Od��?1��?!���?�����	U�@� jPe�w�R}�^*
�nZ�wS��������j�s��*������GA���`��f:(K� �?�,���O��Җ�i��M�h�^��E͇�[�"���B/Q��8u�^���h.�OT��|���yi�m���VjP����Z��"�I���?���?�(O"em��8�Z��'�N�|DZ⣝�B���ä���.��O��'$z6̓��$%��@���*�Hd+��`�D�0?���G!� Z�iE���'/�>��D�?�� ���܉�H0J���A�n��?1���?i��?Y��i�O
U���Z9�ny��H�?o�X96��O4�nڊ";Y�	ߟ@�ٴ���y��G#��E�D�ܝ��㵩�y��H��I�9����e�'���%��?�0��O�R� �U��P8���Ni��'���8����	����	
7�x�{����Qx�zcO<i>M�'��6mn���D�O���:�ӗZz�Љ3cͳ)8V��6��	�|(�,O��D�O �O�O+l�`$ӥr���P�&B���IԈӛ�u�I�|y�፼D�2���%��'��+�P|�V�W�4� �ɂD �$�'jr�'0�Of�I�MC����?���J(W�(pE�a�������?���i��OD��'b�7M¦��ٴ#�`$���ǥy���렁ۇ|��E���MC�O�a$�-�J��D�wx~P��K�4
��g�ŲB�p��' R�'|��'b�Q�b>	�"��
e1G/.S~6h��+YП(�I՟��4Ut�!�O�7M>�dL>L`��e � /��4Z��Cv���'� �����,�\|o�I~&�0J>�s��V���9�Glېr��\;ե�������|�U�������Iџl�5NX� ,P�"�`-a�N�w�����	jyBgv���5,�<����ɟ	r���P�,�H��R��O01�'r�ip�O�
\`�u�M�|>�nK̼����X�a�$X�18?�'k�������4��%ūn��9���� C��p���?9���?��S�'��$Hצ�[���\V�� �*�ۢ�V��4����'6�8�	�����OV}�BC�#v⵨7�73�d��o�O$ oZ�Df.�o{~Y;�^��SX���J�(�����#�\@ACC�}W�D�<y��?���?����?!/���C��	Pn�홤�&xaj���韈Z���O*��O���(�$��~W�Y5&�����)ٺ���a�b�'�ɧ�Op-��i���� Aʉ�^lJ�#񇋎(���	�9�������O���|��fr��a����pY�8٧kD���1����?���?))O�l��C)�P�Iȟ����Cm�1a��j�ygڪ]���?�7R�l�	蟸%��c�b�7T��e�uZ�,?!2����(�z�`Eņ�"�$D��?��e�5N�h�D���0����?9���?Q���?i����Of(j�d�
q���M܍'�������OT�m�f��������1ݴ���yG-��6v�]����:��l5J���yb�|��4oڽ�MC6Y��M��O�9����&�?�pyUH�s�E�P��,A0p�O���|����?����?��dd���I�eJd�	�ř��.�s,OilZ4��4�	����q�S�(co:~v��bI��@8��ܕ���[覵:�4
����Ox�C��А[��AˀoW�ࠪ�C�p�
]A�O"��POf1��4��'6�I �z`�Q% ��0ϛ��R]��蟔��ԟ��i>1�'�6�K�Z���I&@��`p`Z���Љ#�T����d�¦U�?1fR�İ�4cS��sӴ�ɀ�W�H�j	��A�����A#n��6�,?�� "C��i7���ߍe逑W|f��\M�%0�(y���Ɵ���ş��I֟��S'��JF�!#�Z�p��Wb1�?!���?i5�if�T*W��pߴ��0G��;�Ř�H��ĸ(CS�x��'��OV`��u�i�ɘ#0�9�F.�=k9t9I`.�2޶0�V��j��C�S�Vy�O6B�'t�L<f���9B%�A,P����M���'m�4�McuaW3���O8�'>`Z�rT��!��eK� �Q�~��'W6듑?����S���:b��x��� ���s�$(�@�"�bɺ9�H(*�O��?TL<�D_�+w����,Z�<�lIɳ+F$A��D�O���O��<�U�i�B-!�lۉb��@�A�	]@ k���R��'A�6�"�	��D�On��;O�,��J�+�*��v��O(�D�37x6M/?���Y>AB&��+�4�ӬDu\��㊧T٠�fK�y2W���	֟���П��ӟ@�O�(��b)-7��SA��9�Ν���hӜ����<�����'�?a���y�9OѾ0ã��Z�n���-��z�'Nɧ�O-�a"�i*�d�(fhJ�ń0@�������JO󤁦|Zh+�n��Od��|R�(�L#��-s��j��V�BRP����?1��?�(O�ao��5�V��	ğ��I�j�M[��A4)G|�;���_�<�?y!Y�L�Iԟ�'��+�-W3V��I�,�?M��XǦ(?���S�'H1�Όf�'&B�����?�B�-'� *tf�e��8cC@���?���?����?ш���O�U@�� 3���
�c��i�J���I�O�Loچf�t��	�0�ٴ���y�+�n�M	GdA�+� �2)���~r�'
�6Nr��=�&�|��p��B�F�i	w�? �`"���=R!t�Y5�O�K��i5E*�D�<ͧ�?i��?����?9�H��n�xU
�f^����t��9��dΦeR���D�����&?A��;P� �[�!�6���
do��f>��b,O��d�O��O�O���	�kC[�dk�Tt�b��D�"_,6HSZ�܋тӖ[�� {�IVyB��;@\�(��
�-YD�]	 0RL�'���'$�Og前�Mcq�Q��?�6���T�a�U�h5�]������?)R�i)�O d�'6�i��7��]��� R(Xђ FM�W�X���zӴ�7�6�/����>���1����l5x�ȏ7[�,�Iߟ��Iʟ�������L��Jg><Iv�vOv4R�c��o1\5�,O���Lۦ�b4�1�5�i`�'�D8F�%�"�_�y��p�.�D�O�6=�4� �fr�v�vJ�aπ�(rZ� ��]E�\�ŅД��$G��䓗�4�&�D�Ol����a���oB�$��G�J�
���O��PP��$U�w���'W�^>R���n��PSr��6g�q��0?	dV�����8&����0�Cݧ+�p�CF��D�	�,ԉ_V��B�OFI~�O���	���'u$�!�� C�|�9!	Ȅ(L��R�'���'�R���O����M{c�)qM�p��R�|&"	ё�G�G������?��i8�O��'o�7-����˧g��x�\�qß#p�DmZ�MSiJ=�Ms�O��+��Ε��I?-�򎁧ɐ�C�ۖMntP��o�l�'Z2�'�R�'�B�'哟o3��R
�9K ����_J��xܴ_���?����'�?1��y7��>^�C4� \n(3�h��Zs.7˟$�b>I�g����͓[6�THg���
��L��슺CeV�Γvv�q�)�O��sN>a(O��$�OTd�(�FZa�eǤ�qa��O�$�O��$�<i2�i�����'n��'��S����O�V%��EZ�b�"|�5��^Oyb�'��V:��ԚW��ua"@�
*x\\J	�d���9��T����;&�b>=�a�'���	�D뒯�!_�,�S�׸W|Ѕ��������h�IP�O]Rj�-�P�)0
$)���zՋ�����VH 6%�<�w�i��O�΋�H����jKL pA�)۹T��d�Ov�Cצ�YD�[ϦM�'�H�Ԭ��?yb����xWn�{�@��O�H���$�T����'B�'���'�>���O�Pd�gDZ^ɶ\����4�.$����?)����OO���%ʂ�6�m��bZ0rXb�@���>���im��d6��	ȬE̎]�gB�?$�xUA�+��y��iX�lԵ{�d˓^���.s�/�~�	sy�kSx��́�#'���'��U���'R�'^�O��ɿ�M�ш�*�?�dM��TZ��Ve�[�*rfKZ��?�g�i��ODi�'6�7�	�PoZ�wp�����.�T���X�>�BmX�e���}�'I��-S������'����	�iP��B��
305�5��<���?���?����?9���U�~��IK'�����
�	O�;yR�'	�pӘ��d7�������'����,A�`���NC�5��Ɍ�ē�v�~Ө�i 
*N6�x����Fhꆇ�/o��EA0g���7L!lw���c��`y��'���'�"���yS��CU�����#�)N�!�2�'u剴�Mː����?���?�,��99�c
�`�@�!��H�L��D����O���O��O��8X���a��D�5��;�݁2Zv��+	�tĮ8ZC�7?�'K���/��
����O-],��C/�6TZ��P���?)��?Q�Ş��������a)��PB��/v���v��$���̟��4��'����?��%��Ti���r�yA"Q<�?Y�S��q�ڴ��$�/U�i������9	z5V
	E��(���R�b��by��'?��'���'T�S>��F���D�Ppx3JL4~�~`���M�p\
�?���?IO~���r��wl2��♭L ��Q����0L���'�B�|������)��F<OJ�XC&�z��@"�C
+p��2Ofy �JI��?�!���<ͧ�?Q(T�`*Qp����d�/ɝ�?Y���?����$̦�)�ˏ̟��Iߟ(��ǌ��0L#DO�=��9*0��s��m)���L�I]�!T�d8P�Ƅ-�����нxF�Z�Q�CF�N?���|���O��9�e�,�Xĥ�u
6%	�.E=Dռ�����?����?���h����F�-xjA�M�:蒍��DK2Ext�DOŦ��A"��l�ɘ�M���w��ZB�v�<�1+H�b�A�'t��'��6�P3B%�7�2?��[���)Ԓh2)Y���iX������>w�ց�N>�,O�	�O���O��D�OB��	�g6��� IC>��)�<���i�	��'�B�'���y��$<x̸0P�@�s����P���듺?Y��Z����OZ,�z1慠Y���v��,iN�i�ˋ^4b�OԜ��B��?Ć>���<����S���P���d����/���?����?i���?ͧ���T�51��ƟTZ�J.Bx�zs��ҥ�(�$���?�EX�d��՟@��F~��bA5m����@�<�e��ԦU�'\�����?q�}B�;U�PP��#�h��S��.�����?q���?���?a����O�0q�u,G3_��HH��ڳr� x�D�'�r�'P7���)���oM�&�|�n՘^`�ag	N �Ey��ąm�R�O���d��ɞ3^�7m(?Y��Zo�? Z s��*��H��H�-�@q�K1�?A!�+���<ͧ�?����?��կz�ZQ,B(n"
����T��?�����D���VΗ��X�	��ؔO�l܁��V�Y�4�!D� =��4��O ��'��'�ɧ��9gLr����\�aŜ�*��ЬID���d�&���H����ӶH2L�s�Ij)Q���79�<2� ��ThT�Iʟ0������i>Q`+H�8	�'7-ЍI��q1P)I9H�����,� ��j�O��� �=�I`y�OW\˓�M��m�~2�P�$���S�o�ٛ�+a��E0�x�L�Iԟ�KPjX/|���-??�'��%s߄����M`����M��<!/O4���O��D�O����O�'	҂,��9?�hd8E�ŵm3\��"�i��*��'�r�'��y��c��[nJ�"*Z�-��}B2�?z\��IΦe�I>%?�7�����I�<UmF v�3�������S����!�O �I>�(O��Ot��p
Q'Ze�}��@���[7+�ON�d�OV�$�<i׼io�uC��'>"�''�Y�ө,f ��щQf�d�E�dFU}��'��1�d�,<U$�p �_�zz^e��Q9'i�I�J��ӧB��rKlc>����'Nl)�I�Lu��C�@�(5)�1�=���	�0�Iӟ\��v�O������0q�4���F�s����by��)���O`��[���?�;4�]�W���r�!@:w�y��?��c�fʅ7=�����%�:��t��:NF��Q��
8�L!�OB>]��8%�H�����'���'�R�'p�Y$"6z���J�n�r)�T����46�p����?������<�3Ā.H,�XA��*bm��Eo������<��S�'u����ʜ�|�BlR���9Ӷ=˦hW�����')�-z�����|�\�h��K7P��L�o��=]�$k��K������t�I���xyr�1^����O�sA�5a-�Q�AC�� �C�O��ot�N�����MCV�'��&�͞Z�x�W�F�R��H[�aS���M˷�i&�ɆM�nlZC�O��5$?���%�&�˗��w��Q�XM.V���@�	�������	d��JDP��i_~��#W)7������?A����c���D�'QZ6�&�?|! =P�)�(x�0I���x�'����4y���O�����i�	/~DB�[⭎�ueLQʅd�5+�Mڡ�;%��Te�zy�O�b�'�R"��X��=qo�3V��j�
L0R�'�剸�MCl ��?���?!-��4і�
�0��ayv�R��n ���� ��On%mZ0�M���xʟ�չR"MTO�͒s%��m�@4�r�_�u%�E�Ad�,3��i>��$�'r&�|��S	{:���S)$=��������	�\�I̟b>�'՜7M_�q�z��b�Q��s��;k���1t��O�������?�_���۴Y$e	!mҴ
��`9G
�e'�):��i%�7MN&B >7m0?	1�Ŵ����(���]�>�̜�e�@	(�"���_��ybX���������ꟴ�	��OE��0�aEf�$a���9u�JmC�@`Ӷ�(���O��D�O�����dQ��� V|(Q�ȄOJ���!9����I��l�L<�|�c� 8�M;�'P�[h���u�i>l�8�'��I�K��P���|R_���۟(a���{�|�+��OG��P����I�x�I_y�t�*URՇ�O����O�Q e	��E�*�9���Z�f��s+8��9���ۦը�4j�'� ��o@�4�*�`M�cf-y�O�i�Pd�������ڏ�?Y+�O"<�"�UT�P9$�Ҹ\�pCv��O"���OP���O\�}���D�8�!OԺM��չ[�R�N�+���^W����	�p��4���y��*+~�y���e���tD��y�x��umZ�M��:�MK�O��$ɋ)��e�׊~/¥#Tǂ�)1Չ��/�uA�EҦz�)�ɖY����[NO|�ʖ�	�8��qT���;4敁5&�U�� r��+E� e˴�Z��*�� ==}d 37��9R��}��O�q�f[Ҥ���'��	�K����,{�e(_�&���[�h��p��{IN��ꁪt��u�	S���[Vg"K�vx*��\9��0SC�=0|����m� ��U��	A,b �P%A4 q:v��WQ6]��F�+$`���y�p-�����y1S	E`�
4�Ŋ�s{z=S�l
줬�ui�>�
H������':�P���䍂w�А��' [	��ֈ\��M[���?vf�B.�l�<�~j���r���a"�'P�����N���J+�ȟ�������	�?Ŕ'��SP����m�i̊h�7mդ/���޴���k�b�n�S�O��W�ѐ���	�	r48��2��Vʰ6M�O4�$�O����
�O��ĳ|���~Rj_�l0�IIѯW�L�n�{P*�1.Zb�\y�i���'�?���?����!wT`P��[��zp�t����'��A��S��Ӭ�Z��%���5D,��N_�c���R�"ӸYJ�M�'ׂ�b�*H��D�O����O0�]~M�g+/G�p��q���Ҭt�_pI�Q[�̔'~�|��'���I������6->(��T@�h��|�'�'�	�P��O�킕F��|�X@�+īYV�my�4����O�O����O�ic�*����J�Z��i� ^	OOZAh�i�>Y���?�����dD8����O���'� �ң�J�1"T��43��7��OR�Ov���O25�F�Ot-i�Y��+�BªT���:��]�� �Ss�f��d�O4ʓO$n0Q?y�I���	|�B*�|-|�	'�Y?�2�8I<9��?i�j�'>�iT�lơ�������O��]�FS��Bcȳ�M���?���:�_��8� ^}�� ֚Z YV���(l�d�i�B�'��Qː�'k�A�O��'���ȳ&�<[U��6
j��V�	�M;�EH�	��&�'�r�'��m�>	-O�5����� �)r�]o"t�3
���A��
�`����O��wxHy:�FőkP�p�i���j7��O��$�OjD�m}�V��	M?1� ʎy���I��>X����J�"Ơ,?)� W>/��O���'e�p^Y)�IY�I��E
G� H6�Oi�'�Ku}BQ���_�i�MB�L� 5'�􊅭�R���)��>A�f�����?���?�-O�H�A����43���f� c ͊80�ح�'�����<'�D����,�^֤����̂wT�i�.�$�x�h�O2у�>O����O���<�*�'}6�i�� �T JcI�C�1!%�
�($�FT�d��a�	ڟ`�I;V��L�W���@0�	lJ��0��r� �'~��'�2P�X�2h������O����H6�^��GӾy��������	C�I˟�	`�=��.˙mC=��ܱ�FD�խ���ퟔ�'-V%[��~
��?���<g��ɒ)�?.1Px�$�@<K�d�IƘxB�'��Q�P2�ٵ��D�?]����@bD��/P,U�6]k�Jo�B�*�ԭꂹi�R�'��O�6����� y$�鑄	�z�)�#������ at*�N����O$X��5�ҭI��	�F��=GֱjشA�0T��i�2�'���O�&���D��||�@:fg_�?e U��n#(3�$l�Zκ��Id��P��O�� �0���e+��w�>�C���f���o�����Iǟ�Yw)�	���|����~�]��ܘh��Kk^����\��M�����!I�s����|�	�L �"�<h(���5	�gV��4�?tNN�c����$�'��'Ƚ�'�K�_^�%p�'b8���"�$�O�ʓ�?A��?q*O��eق��t��j[(<<5EKR}g@ $�|�����$�x��u'�G:p?00I�f/v��lA��K<�M+����D�O����O�ʓ5_fp�P0�4!)�+bؤKS흗2]<@i�^���Iʟ�%������'O"	��B��`D�9C�\�3�D�{��7�$�O���?��$P
��i�OR@��ҩ-1�LC�9M�q�N��Q�?����U�2�'&}�t#	�${�M�;02�!޴�?)O���ߔ4�<ʧ�?�����1��(x��w�$�h�#��?�<-&�L�	Xy"���O��.������5>�'�O&x�	�8�- ����̟����?��u��ݡD�y�Q�3&D�lm�4%m�f�'�	�kZ"<%>���!ҡnɤ)�U� I	r��k�@��O&�d�O8���2�S��!R���-٥���!54h�`*#]��3B�Fx���[�:�Pt�V�A�Tyʄ(��>�h�l�ğX�	؟|y�$_Myʟ<�' �A"拃D�^� )�'+Ì`�o%�|�O�B�'���?C��H{'�BE�"P�*J�S(�7m�O�X��D�i>��Iџ��'�̔�B�"`���Pw��s3��H��,ʓ�?�(O*���O���<!�V1G�����|M��j�!	��3s�x�'SB�'|�	��H��E�Rб#'��������gT�PoZ��h�'b�'M��P���Sz�	Ŧ��m�,F��a'�ɦ������?1���?)��@_٠�m�1H���ʰr��P�(����Z�H����l�I_y�܏V&��4����p��U"�莔cꅳEgO���I�ؕ'z��'^�8��'���vP a�nv��x1�I�i�%nZßD�'N�ă�p:�S�|�	�?��')~fQ�/M6)��y��d�O����O�i�$�]�1O�S59K�hYRE\?a $BCM��l ���?�D�X��?����?���/O�ɞj��Yb'�sMjMږ][H�F�'J"OF�W$L\��y��J]��D�W�ؐ&�Je��*�6�MۀAبL��V�'X��'k��>�4�V��E�#>���#JnpDQ����Y��I���INy����O�P賎�=u�W�Wfgx�#���1�	���	t-&Ė���$}r�Uw7ܭ����l���თ	ئb��c�'B(��'�?����?a�D0d���5f/gL4б�nܛ��'+��e#�>�.O����<����FdR�]�m����(�L��ǯ��qF�'�������?��Iߟ��'#���$�	�c���ҁ���\��AAP��:O*�����Orʓ�?i���?YF�P�j�l�Eꁜ�^�b�-Ƃs j]��?)���?���?9-O������|� ɏ�.��=�ʙ/h�.��tn���ٕ'�BX��������	 <d��i��
�.ŏ�F@R�gЂ}�;]x�<��T���?I(O�A	`��'�R�A���l ���DI	h,�R��l�R�$�<i��?A��0s�\ϓ�?A�'2֡��@�.+���1�N�r��۴�?���$��?�q�Op��'����ˎL~ ���*w���"��لX����?I���?)�a�h��O��Sj+��ˋEZ�`���)C�j6M�<�v�C����'!�'J����>�;eO>h
Gh��zt�{��&��l�ǟh��}����9�S�` d��i�Lâ|�3�Х~7-Q���`n������d����d�<�!�#/�t)i&���agR�ɃRW�&��yr�'�IW�'�?���Q'v�I��)������)
1<��'|��'mh�H��>�+O�$��� $H�$�u��9�U�V>�a"��i��'K� �U��yʟ�)�O��A�JF�=+f�A�(���A�h*�]m���t3�A�-����<�����Okl�F�d�ᥢƽ2���hW�_�m2�	�z�2���d�	���ɟ��'=��в9F$�x�P�Ӧ~;b5�Q�_�-�&����O���?����?�cf��_�NhK��K�tY�
݃@�U̓��D�O����O˓9�J9H�>��0�L�$Yh6XS�ĳ$~��(��iQ����h�'P2�'�BBƈ�y��3��1
=f<P	�D�X>��2't����?�)O�Q1��QG�t�'�a@m�p����
ݚLS�k�j�ĳ<���?����A̓�?1�'vẶBZ��(����%Dhjٴ�?����d��)��P�O�R�'����t�.�s��Z�X�*&�R�E,꓌?����?�`~"[���&-Ќ����)������B�Zb�lZZy���l6��O����O�IJM}ZwR�0�!l�E��8{�	�Q*��ش�?i�q�|Γ���Oڤa!�P=^<Tt;��Oz���شQ�^Z�i���')2�O�x���D
;X̽)2i�1+�T
&,#'�i�m��'�2[������Qo�l[��T�;e
񈠇�0E<53�i~b�'"l�5f�XO �d�O�Ʌ#��l��Ĉ�rD���">nd7�=��ߘt
�?�I����	�6�k���N��ڧI�S��7��On�3e*IV�	؟X�	V�i�E#����`dT-��m��)�Aͨ>)Bi^��?�/Ot���O���<� �îK��0��֖+K�%��A7C��z�xb�'S�|r�'RbkQ)���+&j�-X.���l��;��Q�'��	���I韄�'�\���i>�+ �Տ9b��Ap��"��%b%f�>9��?�N>1���?3!�<�ԪΔeM����a�-i8Fbqmۿ2��I̟��	Ο��'���c'�IY@U����l�e �H�hЕ!�(�n���&�T��럖�e��0}�� 'lj߀G�D<�����<��f�'��X�PAc� ���'�?��'�5%]�V��Xȴde���Q�x��'�R�X'< �|���a�q������S�?>�u� �i0�	���شB���@�S��I2)��)# �R�HaFJ����6�'�W��yғ|�����S+�Z�L��u��	�q��/�M{�f̀:ț��'C��''��h9��Sd�q�F^��jb�΂�5����4f��ϓ�䓣�Oe����:kl�i� p*��r5�S�{��6�O����OvL	g�_��ʟh��C?��
[S蜓b�H�k9`Ő���]�tK �9J>���?���l����N��&�a�
��1���?���
�<�A���OT�Okl�"S����N�yt�Q��`��I�-�����Ty�'R�'R�'m撌��^�&k���CbM(E�
���'0��|��'1�Z`��d�pAL�Z$�X�0�31k^U2��'�I��h����T�'�l 3�u>��5�T�<��tU/ܐ-��B��0��Or�O����O�,�g=O�	�^g� ��G-J~T`�R}��'B�'��Ir�Y�M|bB$�H��="�ΰj��+��ۑB���'u�'��'����'c�O����F�[Q�2p+I0N�:�nZ�d�Ity2��4Jfv���d��<�2�k�"6�������e�xE��B`�I����I�[!6�IQ��Bڳ�B�^ARԋa�Ltaڱc��Q�'�=��bs���O(�O�0�dR���@ԜPߞdr��U8���oޟ��I	Z¹��W�S�']8\X��fA�)�8*RMʹ4C��nZ�/+؈2�4�?Y���?I�'-��'j��Zf��|��F\)����"Z�[�7���,��6��0����\Z�+�,x��QJ�?ݢ@���M���?���Vq���d�O��	4vV-!��[�`�����fQ$6-*�d�u�H$>���˟���GR�y1��50��0�n�j��4Cش�?q���X�'j��'%ɧ5& نQ��Y��Z�犍RV%������$��Ĵ<i��?�����d :Y�x�vg��~��q�s�.B"�Q��WW���@E{�'ώ�x���2X Rh:A�'K��D9���qGP�������I@y2�̫c2����1�L�YI3�">���?��$�O�� �e�O�1b��-�1 L
�W�N�+�e�N}b�'L�'��ɚ����H|�E+\2<:X0j�&�V��q�,�9���	ΟL�wm柤�O�(��J�>�mR
�-^P�`�i��'���'���X�'|��'�2�O��]"q�.J�b�y��h�^miw�9�D�O.��Q�UvPA+��T?}���G��jIA6��>Nz��.e�ʓ T��i���'���O{z��{�K\�)��YmZ����Kr�[@���?y�g�	 �� �TC�H V��A��>�7M�>n�B���O:�d�O��i�Oz�$�|�$��0L0-�%��.$8���3&��*�oD�I(�y����O0�́;eN2ѩ�Z�]�@�V���e�I�\�	�[�� �O2˓�?��':x�8���}m�@�[�r��}��SG��?���?�q� �r3Vp�S�H�i�"I`�"�F�'��-`�³>a*O���<i������ �A��@+[^�ᥪ]}2�.�y��'���'b"�'��	�����3d�FcbI�r��jĂ�7���<y�����O����O��� �D��w�|1�^4)�h�FJ_�<i/O����O����<e =��I�8�6]�eVUr`��t�VR�,�	iyB�'���'Chi����pb1×1_~�3F�O'R�2��4V��I����	gy�`��u.n�'�?i1��+�)�7C_N0�+�@Y�&I���'��	ɟ0�	ڟd�cf����S?q���'"!��3�	^�?����Zئ��	�ė']$��~����?i��c�T�;�dM�Wo���e��l���"Z�������?$�Ik��'X�I^�
t��ϗ�e�"�祟�~y��S�x��X��M+���?������U��ݙxe�eZ!�j)�u�+}".T6�id2�'Luӟ'����<���4��*�>�"L���S�%<�Mka���b�F�'��'��ԃ�>	/O8U!)�."��xy��B������㦕
3�r�@��py"���O���+\�\]�i�1GO�$T$`j�fۦ���������u@ܬ{�O�˓�?��'�(�X�m�/���F ��hպ�4�?�-O���<O�S7n�����ٰ ��hɄ̒*$��Qc��Jy���Ʀ���y�dџ\�-ÆJ=H�f${Gcѿ�p=UO����d�B�Crn�(�J�c]Rx(��ɔ@Yڣ"��x�܈����(l��y���7>�ihWH�wu���-E�9� $��L�تfG��r�zz��Ń��pB����5;�F��F��S( ����
����U�ȂT'L}���\�B' PY��(s���iU��"+$=�� [ޟ���	>c�����ḑR��a�ɸE����V�d�bX�a�� s���$���O�Q+(�:]�� @�AG;wz��H��'�p�����?	+ON�Q�ה1<���/۱w��{�2Oz�D�O��"|Rdb m�D��Ɵ��If!^~<���i���Pk�x���
[�
 ��' �	4u�:*�Ob��|J��7�?Q�$ c�F}�ՄW>s��Ś�'Q5�?1��T�5z�OV�~Ra��>�O���Z<� E*�(,��c�*�h4l�'|�h�4�X�k�(�Kg'�~q�H&b�Jd�
��V�Zp���O���e�'������pъ������$A`pM;�E?D�����[�vI�"�_�'[b�0e8O%Ez���E� <��J\:�%PE�ʏ|/~��?���M�@=+&"�"�?9��?Y�Ӽۢ+ް�prS�\j<x3n��ܢ9�Ө' ��@��ʌҊ�L>���>M��т�'�3]`��:�n��?�@��w�-�1G����}&�P��aɝi_���'V�5V-����ɟ�'4l�b��|�����3[X.4!�F��N@uB���*�!�D�+�vT;��H�1܊jB�
 ��I.�HO��dy�+ީz7p}�TV��*��ǈ7��A���9H[B�'N�'5r��՟����|��k��vhBԉ�ljP���*`���c%H���>�
?��K�	[3R��8�0K��k��Մ�E�^���E�E����1�E���
�̞�:R�����'B�'�bU�l��f��A'�9�P.�@���k�ȳ^��x���"e2W3�B1��%���<��R���'*Y�$��>���s�Ru� z�`�C픭H�RD��?��Y��?�����h��m�H�� ��?y���sָig %:��XM����,%T�-��J6��-	 $8�4@G.7�o�685bh;�o<^TL=�'O�����}���'b��M�>���@�gz�!-g�c���	Ix���@|;|h	�.ћY�L�r�' ����4z&҈����G�v�y�Dȉ)�����dB?@e��nZ��l��q�4��|��L�	��!�5&"y��싫w��'��z�d�0�1O�3?ᄡҪJ��S�m�8�B�[�,�w�d��(�1�{����C'}���"[�<ɂYI�G��I�	y4�D�Of�����F����Έ�)A^�//��z2��O���D,i���R�Q)a�3c�kax�j7�ZyF	s�]*	�dIp�	Mh0	���i���'A�Y�}�U6�'X��'��w���K�U*Z�n塃��/��h���'�DR��7�|��M������I�-j�x3h�G�b�O�ma`n����,�X�@d@�)X��Ѐm�2����?���* �S�gy2�'�̅{�c��B��[ ��~�8�O�ba�Θ3� Y���ڋ/G<{S���I������<�Q�K�p�jB3dAp�S�<�"��
'����ȆT�ݸ�ΆK�<Q)^"x$��XD/S�'�T���Yo�<Yd%�>-Y,Hق�_�=<fĂ$�_T�<9�R�X��1;f���`Tl����O�<�Y������TQJ�+�͐bDB�	 +��	K�j�6/�F��ի1J&B�:"T�R�h�.<04,?\|�C�)� �燁(:i���ݙ,��lQ�"O����X�,/L)@�)-Sy�Ԓ�"Oj��B�{u2�9R*QkR~�#S"Ov�X���A@��iSM�T
v"O~5{¨o*������ .NM��"OxXy0o݋9�t���nǜt9�"Oik$��$e�"Y��#}��(�"O�{��T2a �/HB���0"O,mX!a�2,��[E���Q�n��1"Oj5�bc�2
�bE�D
~l9��"O|-1��^�I��|AK��Z`n$��"O�����v�Q�d��Ze���p"O`D�F��
y�SSB�+c��(�2"Ofaz�i��SB��⧈9�։bq"O�h�Ⓐ 7�ՂT'�I	��Y'"O"8 3C�)@<�X�=�,<P�"O Ak�	ͱT!���f��v�@�"OС�s`��bR��0Bnѽ_�n5Ȥ"OH�8�!8/��):q,�?Q�(�P�"O`pYe!ݓq�	��b�"OԔ،X��� �U�g���A"O��)J-e�����V�tU8xچ"O\x�#-�!O�,\���N�d�qf"O�L9TH�z�,����J t�"J�"O�l6D�(�`��(pZ�"O�<�a���i��ٲLjx0�"OB`Q'��<Ml(� P�E�FP�Ѡ"Oj}z��4U�&��E�S<�j�"O�|�!@\M�d�c��ܶ_ Ը!�"O�,���S�@fe���^�zܑ��"O�b��H�#|��ū8	]s�"Ot�25j�r5"$`�;8	 �җ"Ol��&z��!����0�%�&"O��Hq���g}� dK�Lc�r�"O�Q�� ��P�
�s�@BH�X�"O� #�i�����?9`���s"O��9��	�]��m<���"O��p"�:a�"=�?C5���&"O0rq��r�^Dr�G�,mn�b�"O�1�2NOS> J�̏E6���"O�����>���v�U�T�йZ�"O�Q����y�dݢD�ď��i��"Od�#�H�yrTq�V
|ða��"O��f
��m��V�Y�y�>M(f�'��9�VA8�O�\�oV=2�j�B��H���MSG�'3���@*�<��$�R�Y��}�(��q�T�<�r��[�:ՃكM�DT[�ij��n*� 5��8�@�����m��"����i�C�	70�Lа�,R)0B��ǅS�T+QCC�O��h����.������ļq����w�J�6h!�$S3rK��q�-�F颡� O32������Ϝ[8��	��6d"�XD@L�{�&��A��s��A��6^:��1����&І���-i�L5�9k�6D���Fx�V\*�#0$�a�e�u�ڌA?�%�am]e�<��A�d��M2�iT�z*`,�V��b�<��m��F��HN̏=�� !0��_�<��;���u��$h�����W�<��͙	N���$�1+��HG!�S�<��4���D;^�"�8�ϜG�<11���'�p�6�ڛ*�xE�!F@o�<���B=
�]$ac��tB%�i�<�qo��E�=�E�IfZ���Fh�<ё"؈_���+���b�zm�1Wy�<� ����Y�-� �1Z�Rk�"O.$�>E��Rv��)3����"O�;e�ƱV��쀆F�
i�����I�W�~<G�4⏯Z�Xe�pΑ*RD	���y����(����e�1�"�bQ�'�~2e�+�O�>%�5 ۝x�k�D�0H �$D��@�AI�RA��*�E��B�H��7}Ҍ� -�a{B�B4S%�4C�v"��wK��p?�R��M�B�ɰ3B�ł��ۀ7&�����i�<��
Z4p��8�I�0�[�?�Qز����ԭ<y\�[�I(jֆ B���s!��χM�"1XuG�O��Y�˙r�!�D�^��%�Z/�6ԩe��	R|!��I�B(����q��A��40c!�D#����0� RA�ظ���)"`!��b�N���!Į&�֔�'ǱT`!�$2� ���\0whdX�&� ;�!�S+x@p�"��$s��� ��1
�!�� Jר�3?�P�Q��,�!�$�Z_�p��̊Bt����Ʒ�!��[�2����I��&�WOC��O�ԑ
�T{��	1��N���與�Ix≐x��	��̊ 5���2��;���rQ�`(<����9I"�4�$�uƺ$r3EF�#���'��5� +�����҅��	�$��fL�B"B䉩c謍�3�΋O�A:#�̜HZ4�8���?��� �s�A�F�����p�Ap�ۂUk�u!g�\�X!� �Cl%����>�4X�6��ZP �	�v L�{��J�A4�l�[�l$GzZgd���\�`�@�Fϣ9�l��$�#A�V�A����� P"�E����;�d)��0aZuHDj��F���ڄJ��͏i-��P���s� $��R���3L �U�]�T�����J	Jy�O]V�k�� 0֊�À-O�UX����'�h��� ֖Ol�)����.�2���
�`l��N�\l�a�,O1�2���gxލ��	�wm:����'fȱbf.$4�<K�M
=����$뎄7O�ܱԯ�O~�A�=I�ջg�O�_I�hC�o��O��2V����|�+��ORܦ̘U�'|�)��_&\�͚QI^#��	�n�;�^��e��-kr���ŀ� Ahк��+v�����2�n�qҊ�#Zi։� Hw��'�ֈ�@(7~��)��V9g-=�I<��&�𳒨T�t���@��P��C�	�`w6���%<((�)%�.r�7�ބ:�� {Š�Af�A�m���T����=Z�G瀧E�P��"O��ق�.2�X�[%(X�MD�d��mH�� Í�
���@H�0��9.$�Od)���ܖ:�$pz  Ѥ6n8%yW�'��Qv��aT��o ͖u� �<m�f��RI�:pv�dI�O�����ɎL�b��c�!?đ��(��"\Dz�C�y�FQ���ݟ�b��ެ��nO���ӄ.�o��i�M
<4b(u	˓G��	��N�48��Q���O��׆�'���#v�M�t�q��'eXY�A�K>f����0w����_��!r�]�4}���v�\m�(�D]�R�֮#"��H<� �č�.E��I��-��ъX@��$�*዇$y�Ē$�(�b �QGR�R>xh�gBQꚠ�D"����K�^��8��c��p�Pٰ�A���ԉ�蛞{F�c �-k��O���� ��g�MJ�HQJ�~�!�Sh��Pæt����4U!�����p=��_��lY�m�g�ܽ-?�f��*�i�0�И]n�Z3e�\��qK?�@1nۖ� ��΂s���B�8?@��dS�Egn\���E0������"2+�iP5c��t�� u�^5"���&t��΀-?8R��E�?�)�a@^���p�ij�Sc�D���߾>��(�*͐O:IcU&E�a��e���������(�e��-2|�6KB�FhP�j�ߪҸ'��>�	693�%�#9� ��±	��a�7KN2[�"�х ����ĂґI>��$h|�18�#�*g������3��	����pB�'��xR�͘�=�l�b�)�)��� R$*�ɴ-}d+̓2-F|�Cc��Q峟 *%�W
y�����L+#N���7,O�B���Ɯ1`!B%����˔#��=R��QY��k���;>L�3��U������6[���3�I{��fF���ɆEOsd���0� ���3䖅�4��A�f�8$�M�,���=�Ɔ�K��T��@G2$��T���XŦ�Xf��|ܓ/�>��2�	#5��:�rp��\,| Z�c�M�W& W������(r?�S�g�? �Qv�@�O0��jQ�� ��v;O�����p>�PD��Z�3�˂�Mu� ʤ���O�ĉJ���_�IU��Q�O�tXr,�T�]�d�j؁��I)�"xAqfɳm� ����	�$�Sk<4�����%��|�lG�YcbIº�x\��ط<A���q�xД'���>K��x1rf>f:)�s���d����4o�����\�.���J΢,��D�x@��3$*�4u��I�$��I<ЋKI�I�dE�%8�@��7��.�b(�3N�'r�N0���S7z�.扲{c| ��k�>t����PKbc�T���p�Ac!lJ%pt���KT�l����� VB�ESO�X8Dt��"0Ҷ��@ׯdjM�ҥ���) 'e�[�tO��J�$r����׆$��w|�La��\@p.�y 	,A&(i�O����n#K��i���H�����D��:1�X�m+M2KP�(�p��F��j}�'t�RD"�_j�ֈ#�J�l�@�wh��[��EhEÑҴ8���>�(u��p�F�H-h9p�J�6'���{��	�p�K+�l�rp�R9p�p��+�X `ώ�cVJ�����~�Y��)�e��&� �($��rR,d�e��c���̓R�҈(#�R�f�l2r�O�fA ��'��0���	� N����p�B�n����3Y��;��X/w��`���&|O�):�_.xP�Q"bިq�)����#	�������BK�/P�H�#�f�P($>�N�u1�9�E��{e��I���
TE��Ը�|��E�5[تM �!�/v�&�����Q�d]����4P�"�����N?�`Sc���l�����fG�Y��K@�&#�]@S&�p<)��-%��O���ҟd��$J�n���b��g��H��F�T.� 3��G|	��¯Yn%�?�r��&\�p� c�qӰ��%�Dq�D��A9�y"I�.Yb�`z�G�������8�5��۫~T�Y a���WOʰ���M�}༼�C�'�J4򮖶XH��CN�)X� �yBF�EР1b��\�@/jh9��D;��4�$����]�)�2M��&�'󮈉0O0��ªT�c��X3�Nu-ֽ��Y
k$Zd�<��I*+�Z�>1T+<<y�,ʐ%I�/yp�V,Cj�<qw&�
~�4�#��]E��+g�[(w����'Dr��BB2k�n� A�Ԓ<�Fu��'�<Y�����.��J�0]�p���'��mq6�	H�d=�h��Sqb�I	�'޲�YrfE�[����ܲP�r���'ܞ<H�j]� Y����
CHRQ��'����щ��ff#Zd��'M&�"F�L�+H~<��B�n���9�'�0���/�~99��o�މ��'��t��b]+/���B��0W8Pq3
�'�(�`�D^n��k@�ش?_�<*
�'D������i�BՉ�� �.�|{�'M�d�mЂp3S͒p"���'^R�#G��%�f0m�+��'���P$G��fH� G(E������'L���J�h�sdB� /.�A�'�I	����t���Ə�.]\���'��j���h�`�`��o^h4)�'�b��aFL�H�KƋ�6mZ��+�'
�(�f�`C��S����z-�*�'��h0f��:4�1��8%kZ���'�ʌ�u��=����V�Q�$<��
�'!r����͆?R1�5`D�l@�S�'zZ�9 ��-M�ޠ�����D��'�J���-����u�3 �Ih�'p�FKQ�w�K�'�ԙ�ԣLd�<����$�+f "t���4�`�<����#R�Af�A�4�!`bR_�<у+םŜ�#��6�"E��#�W�<��%C3H�8��`IV����'�]K�<9!���:��A��q�s�C�<AB��#M��P�.p��W�	k�<9Q	~N���fh��7�RT�v�}�<ҫ�|,�D�^����z�<�3
�i_�7��������=�y���3HA����̓�©r��ydҔT�Dqs��@1 ms����y�ɓ�cf@�����8�ZQb��_-�y
� ����OX�Z��h�C�]nD�"O��8�c�?q���˵�W�lqY"O><�#��R�@����S�ؤ��"O���V![��y�j	�v�n	Ȗ"O�(��04S�L�*��_8왉3"O�}9$�K�=㞰C"):��bU"Oj�f��
�`5���U�!1�t��"O�LYe�%&$Pr�_�B)��"O|�@Ӊ��7{�T��*X
cޥj"O�3��%tքu��L_6^� q�"O���C��)�t�kq��#
4�P��"O����$O�M����3�ʠ[�u;�"OL��Ӏ�7E�Bqju ۼ�*�[�"O�-
G`PR��(��,p��A"O���#j��S|@t�ٶZTE`r"O&��ER�� qd�ŽtG�s�"O���KG)M@fAQT�M
��!+$"O,�+��Q�����D��asz��V"OX�ńW!9N�kE� �mU��p�"O�2��@���a�"B;Hi�w"On�ԥ�}��t��;H/��	�"O��թa2�͚p��;=2�"O�,���-|H=�@.ɀ|a��1�"O�0B�DM�p����,�� �6�)�"OB�I��`R>$��CC�8���"O����P1�FD��i�02y��0"O�q �R#O���F�_;nC��z�"O�aAG(��0�a �Y�مĈ�!�D Ht�mH��� ��D�b�!�d�K� �m!H�tiHr�ǯ<�!� �`���Ҿ|�K	}&

�'{4]��O�2�2��A�x�k�{"�)�) *Ľ�d���n�M2�ժ/!�$FS���@KX�a�O@�&p!�$�72�尕f�3�*�s�.?�!�W)y�,�fђ/��Iʳ�Ý
�!���<����P���=�0�H(!�$�4+:�p)��^�[�ɲ��%�!�䘳g#���G��hid1�UD�!��R�u�� �AѬnKpQ���G�!�>��HUNǄr���P�L}�!�d֬4&4��aO�s�*��1BB5r�!�
�m�Pm��ްG���r��/u�!�dM b{���HW��*��ua 
6�!�$V�i�6D�+44~�G��T!���ej��cg��s,L� RU	!��B
 t�Cfb�#O.P���)�!��E����Iۋ��A�K�Rx!�dZ�(	^`�5"�	:pJ	�R�ns!�V�sI�	�R�_���Q@�\�!�dش?o�!�uc8AJ����s�!�S�x�6Q8R�a� �!��N"c�@�4�E.�P��㎺5�!�$�z�$ ������%b��"N!�ī��j#��a# k� F!�D�s�0� c�+s�>p�*8D�!�dQ�T�
T�g.)��Q
7/ċu�!��jFJ��b=r����soˮ]!�$ʗ=����4�%h�x�Ig�]�d�!�$]#"=�j���|��H�f.�;t�!�E�93DAD��+�dp�Vo�4�!��V{��E2LG�]���r�!�$�,��)`�
+v�jVM3�!��ȼl9r�R a��+j���A͠8�!�� :���M�^\�����<��xD"O� �!��[�EcV���W��;P"O��H������ȷ!_2�,Yy�"O
 �W��R�d����]��<p"O� ���Ň'�ĵ���;1��h��"ONa�`��� %��Γ�0� �"Oh�	9����͒�
)�V"Ov؂�Xq(��Y*�*�ZDh3"Oy��ȏ%
h�y2u��y��"O�U�'BG�v���a.ܽT�x�҅"O�$�7�B.X�ZSM ?~��P�Q"OBX��#�i����
�.��á"OIr�\6'<� �!� &xҜSG"O:3*ˑ{R^yQ��
_ �c�"O���E�Q�;9T�{EF�D��b�"O��A�������,�ر;�"O��j�)���0ؙ&��G�0���"O��j�AL�KB�]��fQ�m�f}�S"O.u�5�˜u\ %`�#Z����Q"O�Mۇ��9kƪ(�VŒ9|4 0�"O�<��O�d�(�k� ӥJ��a�"Ol�j����:M���_?u^��"O֬� œ�("�c������b"O��˗��K_�`�¦Af}�"Or��i9���I�P)�"O�	�����$��	B*_��(��"O��kE�,�9���E��90v"OZ���8Z:����ܖqm�@;�"OP9�ƀ��$��pӂ�P?]�'1Oܹ�Uɚo�z��b�J�5�zLc�"O-k]	�D[���� � @�Qo�<���o5���kR�3���c�RD�<��LH2�f=R�=I�{� �|�<i�]+]��т�P��s�PA�<�N��g�f�K -	5d�����Ts�<�%���1��)���ԭj��$H�b�n�<���խQ
���j\�v��h�<�ҁBI�i���t��4� �Og�<�v��
JM$�1�6E�⴨Lj�<!t!�YJu�c��/:�@��rI�c�<�ǚ3�������+���weM��y�,C����C�0�C!��L��!�'���p���Q�D)�l��9��
�'��x�N�
&
�"aM3�ܽa
�'��p�\la"�S5�Q�<K�:	�'�"�PR�
�5{J��w�<<�)��'���z���dЀS �W�aBj]:�'��ZS��K
8�i"eҠ1�E"�'E���Uj!b�d���W�
0��'ؒ@���N@	��$D�5�'`�d�.�ds�%����H�
�'�pK���$pr�l)� 
�Ȍ��'�`	�e��v�IѠ�Y[j��P�'��0� �E�a1��B�&ݓ�'>�i�i�+a�-Q��1��c�'���� �PAAu���!)��p�'�����F�����c>��L8	�'2��%�MI䤭����@�a��ONA*g��9�)����)����I����xe��E1JXQ��ɞ�3ux)��"O���)0븴a�)Ćig�"O� ���������H�
�r��"O(P`�T�M������7�Z�hg"OF� R�@�q��m7�5!�l��"O� ���/%��"�ӧiu�0�"O4���a�#+��t� N�d$M�w"O��3GB�Y�h@��K;L�A�"OL��#���$���Z6�ϙ#/�S`�w�O�ک���Nq@$4���b�͓�'エ��DY�,X��R�eR)Yش���'D`4[�hޖ81l4F��a�IB�'4�M��<r���
��M��(��d=<O�Q[�Q��0d�C�U���tK`"OF���[���4Dx����6"O��)���V5@�اC�2�r ��"OxA�bɁ�.�q	U�w�Xq��"Ox5t.ۀoE�PS�҂3��;�"O~D�Sj�v���Qf� T�X��A"O.�q��Ωh&�t1�!J.g��;�"O�̱�B�aT�a���vi��!�"O���F�/*�&��'E?EQę�s"O�u�Cě�%�j��!�)���"O|��iЂ;��A��R�^!�%��"O6M����9��h��N�C�T�@"Oܐ�W�4%�����R�MVx3�"O(xhp�8R�ޔR%cڷH�,�"O�I;�6M�FTC��+^!��"O�<�� P'hn� 8r�T�L�,��"O���!�.u׺k����8(�"Ot�	"O�=:�I�NB3E�)��"O E��K�X�����зd�XW"O֠�q�=�H�Qp�1U00���"Oh�I*m�-b���q�"Op�y�%Tv���_�Eg�0�"O,B@@�>x��a�� [8��A"O�xHԡ�y��	!͕&i� �C""O���JYW��ݻF�:׊<�T"Ox)9�f��z��Ig$J�h2�i�"O�H���E
D��Z���5tS�<�g"O<�����bߚMЗ��`.��"O��1��¦
 ��`��A�ٰS"O8����
I� �@�J6o!�j"Ot}�c�"�� Dٵo#$pjP"OP��Q��.]`�e��Us��+e"O�8�J22����_)s���d"Od��ɗ+l�4���ɀw��a"O�y��/�*x���
C��h^̰�"O�I���̫I�@�JsHL0i�"O��!��� �s�(yJL`#"O�A�5.g$ͫb/Əc7���1"O0��5 ҵOQa0f��&FT�t"O���B�� �a��m
&s
,�"O�� 'i�Epʙ�W�d����"O�����	�Z��GG���%AB"O�('R�B�2�Θy��1"Ob���j�?kzB0�]�B��U��"O���1�H� ^�q*��I�q@�"O�h��m�1n�L��gM�:.�\��"O,�@Q'@�n{*�S�B^�4IYf"O���G�[ 01P�i���'�(y�"OԽ�B΁u�H%���W�&��"O8|c�B�;qt����bW�h�\]�"O,�넢�X|x(w��*O �!r"Ox�Ӂ�
�~�\��KF(~�d��"O�M7H��.x�|IK� g`��p"O���geN�8�0}2FI����B�"OE�Ї�5SrыPg˘?�4��"O��F�W����(�:y�"O� 00x��D�Y�p���o���"O��� 1�B��D	���8��"O�0��7m���[��K�w�L-�"O\ɑ! 7c�P �(Ȥڠ�§"Od���fՕZhm��;[�(rf"O�L*ĉ�!Ar�+���2>˦4C�"O�bd�Y�X�*�˦!EW4�5"O�!���/yj����,E�|;"OR,@�%� 򎨈ǯ�-(4��kF"OL! ����Y����$�>6%�`��"O(`C!�j��yBP�ʤK�"O���O�X�g��`e���b"O򩢠e:/X-���;e(HD�"OJԫE�և[ː��tjW�n�@dc!"OX�����&��4$��5�P��d"O���A:4��Q&U��k2"O,��� ��jt�viW DU��"ODpU@�8O�	h�'��4��V"OjM�'�}��s���^�b�"O.T�Wŗ3f|���r����&��"O<i� �Q���d��,@�J�H�"O����>����3�ݎ+�Ҕ�"OX�"A���3�V�sD��e�,���"O�y
td\�!Ҁ��s�U�2��a9�"O�K�#ΟKs+����J=ZA"OP8p�H��B�s����j��܁�"Oh�(�c˫'ʐ�;�/ǼL����"ONq�T��.+=h,�2����x� "O��p@�mSx�+��k����"O8�
D�%aa�0� �I�pU��"ORQsU��O5�H�ot���"O��wi��v>fhDއ/�"�#�"O|!c���ug�9�Vc#S���Q"O�KEǈ?�\�g�P�����"O.P��i�
Uy�)��.5�D�ʔ"O`ݡ��-CP�e�^�t��F"O* k� �1�<k��I�s|��b"O����+��`A�����R�]��r�"O2	ȃ�T<
�L�f��.\����6"O�aQ����dP�&b��P͌��B"O`��'�S�%)x���@˶�����"Ott���2�H�v��:���:G"OԐ*�a���pH}�����"O�0`�����XM'��*�&�"a"O����Ns��eJ���0�"O(,Q ���zg��M�>T�T���'��T��eg,|C�
�5��)�'�H��'M}\Ĉ�`� S�'IN��, 8U���3N��h��'�<��0��:Y�h ��{�H9��'��\s�H�^���J�Gވo���'���3�̙�`B���� ;}�&=�'�8��f��P��b#]X�г�'�v]�@Ɣ�9[�C� 
B��e��'b9�uF�^��#��ʺ3�|D��'8�t1�58Y�	T>NL�*�'=���$J"9Ne�:�m@�'8Pd�'���ޙ�o.��X�	�'�J-�G�9Uk&�P���	Tr���'yLx����d!X(�t��O�����'3p5�4# \o�*E\����)�''��S��P�Of:��X$:�t���'0�D�5!���0D�(4��#�'����B��eMFh�ƈ0������ �i9�R6s�(y�� �!XH9�B"O��x��<"�$pe%Ԏ-g�<�#"O�q2aC��l���+��L�8S|`��"O:�!�]�O��� �˃#Y�Ԁ"O.5zqԗ�j�y��ِSK��z"O�� �_��-��)�
H� u"O,����	}7��3/W�>�6�B"O��N��8)��kB��DF���"ObW?2_�` A�J�4��G�z�<	�n����'��;5�)��Xr�<��^w���B呐a\���Fd�u�<i6L�?Eh�ͰR�T�Jy��x�<d�40�H�^#cԍ˔�s�<��M�1u� ��Lo;���*p�<��
	�rq�+}$�p�3,�h�<aǂ�>�x]���Y�=���U�M�<�� ��:������>ro�P���m�<��ȓ$K�\XD�͔b����P@�^�<I����`��"̔�� F�@�<�DΛ�|��Q�ČV�H7�!h
@�<�%.�@���@�]�1Pv�*U�z�<����+�>���0n!��)�s�<����(X�*m� ZWF���,�x�<�Ъ6n8v��'eֵ1̬!!3g^�<�E�bzm�%�q���X��Y[�<����r{",�@�I*$��(c���X�<����S�T9�@c��j_J��Q�<���E��f9 �Z�]wL��S�M�<1%̀�A�� 2Ꟊu=䤚�CWF�<��F��SA��j��B�0gv@�A�<1���J}��Y��?V���I�{�<�J�98\�XE��/<jЄ+���t�<��l��
�,0sF$@.O��!;� n�<1��],pʤp�(�x�B��s.h�<Y��X�� B�ɉ�A޲�ӪN�<��� fF:tZr��2Qp�"0��c�<��+�)5��C�ȲQ��e�Bd[�<$]�W���{�eI.:e�Q���Z�<�b��8C�0�kC��(,*�٣�*_�<9`㜩��b��T?�cE��|�<!�#��2#��)�`��т� QC^R�<�' P�h؉$�K���,`Re�Q�<�h�Qffس%Bߢ�VPy�N�<�"�[�2��Vc�mx��d�K�<I�M�"6�h��s#ҁF�:HGI�<Q�Mg>s�N��1
�/�D�<�r-�\1�!��Kр[ ��Cv�FE�<q�@�9i�$B��d�C�n!�d[+b��������U��b�B$!�J�&Y�� �)1�v!���Q�b!�M�v��I��)PIn� ����
!�D��/��T��N�2AT�: !�ē�cF��gKN[�������[�!�Ă
{6��Ha
��qxp1(��B_!�dվs<Vܫ2L+(T�ȓ��Էe!�dR
*� �����rhX#��-	p!�d))W.-�3`�6r� ���(��kt!�d�`�6MÁ�]��QJ{!�DV-,�8qs#.�Kwx�����N]!�:G���Ae�@fA��BQ2y�!�Dι.S�X����G&��(�ԘF!�D���ܙ2�$��?���[�@� 3I!�dޠ_m��!�8Y��E��T�e�!��B@.`�KC=�� C�oJ �!�� ��(�E�&LH<K�苗u?���"O�A�3B�f�|q��L)_�����"O(,�V�3�5����+�N�8"O\��!��J��8�ǂ�K�&�X�"O�YB��)U�� r�h�Sg"O@�1�����ٻS&�i�<�I�"O���#K�-@���䔒f��U"Ov�y��������,_� ���	h��AE��
s��i抠Y\HPgB2D��Z��Q'"��c�G�5\� �-D�X%kF��
��D8f0���0D�@���,�Z�A.D8k��-�7�0D��i@�[�z��ZăĚy�^Q{Rb3D��1��Hj@��B(Ƞ1,>�K'�>|O�b�h�VD��+ܮ=a��E�U:�vd2D�8+��S"���2�ȫaN14�@�դ�$�!3S�*mj�i���V�<р�Ǒ�> �!Û%e��Aa���@���?a
Ó$�)YF�V�Z���$Ǥ9���ȓJ�ʈ蓬_ĖVI�jOn�>,�ȓV��cD?7��k�a�)ș��	����<��D�	N����/
�W�v�q*�R�<9�%�7��B�a���ڼ����t�<y�@��	&i"�B˚w�TBL�<Q�Ô�_��Daq��iz��{Ј�D��0=)&�B�����s��*�4�Z��u�<�+�)n�H4� �Q9֬�g��E�<9���ܾ����9vh��u�L�<��KZ�g?�Ir��E�~H��_I�<)��I�e����  ��Z%��F�<1a#� �����b-2�2��RF�<&�W�m�H�s4�X�a�z�!EJ�m�<��� Q&��'VI��%���s�<���M�hh[�d[��&U:Q+Ti�<)B�ɏd�L|
�h�
?���!��N�<Q��l�(���2��E��kDG�<�".��r`q�w��*h�(8��@�<��%�
�0��)��\�A��	@�<�A�0:b�Y�eɋ)W�Z����U�<�U�<UaL�"d�H������*�|�<9Rl�JL�����`�� 1�O�<��Dp�':6#���.G�<��G#/�dP6�N>a:a�s�E�<!���E�|�Ⅱ�7g���hG�[~�<��O5V�R���ּj�b�pB�o�<I�ᐒI�\�#�I9mb�Hxf��P�'wa���[f�N�ХAQi�JԈ�']3�yb��l�F���Ë�[� 0��.�y�Ǒ�?S>�V�W0X���۷�׮��O��d?�'>��3����/�p��,��ȓE�����r�@:���w4-&�h�'�ў�%.Xҙ�#�T8`��1�T���r�0C�Ɋ:W����Q{ohd����q��C�I�Qd���� &4ĺ0�J�{�C��,6���(CK�
W(��g̛}�B��NY��Sjҍ&"�YG"�A�v�?i����8,߂}`v�ړl�:��7G��bO� ����F8H��1g]�EKg��(LO�x����L��V-��2�:g�|R�'=fi@�@��8�<� �&�<�^8��'��IC�����y{�	C�k����'�(�YBΐ-~�Yc�NJ�d�T���'jD �^&#���� O����'?fA�0���x���?uh����x
� �x1���rc���#&R���h��	I����F�1=��bSMɓa\6�����<�
�T��4�#X�$�0Ĥ� {|ȇȓB($� B\l�>L(GBӘް���.���B��}��M�"� �:͇�|�"8�Ð�L=�ER#qM��I�����*�m��BK�Q=��G�n�<y�B�)#��1�IZ�@��a!�E�	z�ГW�S�EҜ0�b F��(�C�2D�`��,��I��i�tB�S���"q@1D����)��2�}�%��yz:!���0D�be��/����I$fN �kh0D��zPo�
i����2�@�[�,�d#�SܧZ���#�/ȁe�D��s�E,I7���e�'��� CѠo�<P:BCO�x��$���<1
�`T�T-i0�P�Y�t��e�2D��XW덓Q:��@��7~�Z�B	5D����,%k���%�	�z�Npa�3D�$��m˳"�@�!P�m�6H�2�1D�� f[�zpa����l���*.D�|��K�<&�EZ��-	�&�X�)-D�l`�Y6=b���IPK�.��C@*D��*e@�,h��8u�� J4A��)D�T�3G�<�G@|��lXb(D��1U"�8�R�;���FjaKW%D�HHP�O�J����нFONIA��6D�tXЃS�3��5�̎;���S5	3��b���2���>O���en!'?$��@/D���I��lDr����JD��p	e�?D�XZ��S���D���[4�~����<D��J#���\1��t��4w���db>D��tb�zaD,�4��24���) D�`BR�Of@�@fˊr��(D�8[��oR�yT��'*��aG��O�˓�� �'F
t�����@��Z��yՋ_�<�5̀�N?r���˳x���5 �D�<1q�/x�6Y+�h0|����-vyR�'Z�� �ϑ*u���kA�2XD���'|UJ˝�Vђ��al� 5�L p�'c�	i��V9w�Nj�B#`���'�p� #Fܡa�:�PR�ݾYP$I�(Op�=E�T�N6:������E[��1�y����t@"��@}�h��h�"�y�M�0X(��Ve T�i�����y�&C�	!4�b7̱7 ځ����0�y�!� P�zD�yʆD���C��y�� ��vՉ�I s�4��`�&�yBmR�hl���%h{H�a���yrϝ>+A��V(����!��,�ylH�ݼ,RT'�6A��A��*��x"瓺5����
��q |[���a�!򤌶%nv�a5I�9N������%z-!�$ɃR��!	�@Ď(�Y�1�"#!�I34���j\�D��b�Ԃ!�$ήjNxa��q�l��*0 ��}2������YB���F@�A�@�"02D�8��+Ia�������[��a�1D���uK�,'�i���P�%� )!c�OC�I<+2�R��J9J�� X�6�4C�	1y��$�B r�������w��C��.�����T�Vǖ��" �4��C��%v���)��$bĈR��;цC�I)�Nh0�E-l�,���E�6C�	5W��� e	b��8���&x}$�=��g�? H�0���JI�%
s��5d��[q"O(�w��KD���w��W^4�f"O��Bc�s�RTyХ6r@��9t"O��b���.e8c�!BRp+�"Oʌ�H+4U��C[d�ib�"ONTYѠK�?��*�C˿A���"O�ȁ���	PeBq����\��h����OJ��i��ͩD`�jV:D���}�s�Ʋ5h���"J3]i����|�	sV/��Q*j(q�S�Zl)�ȓ0|L�15�� �@�kڳ=6����X�hպ2�C&v1PW1\�m�ȓ1�F���<;��iVɞ,y�z�ȓ5���u*F)sfx � П~�f1��O�n���@\��i7Z�ȡ�ȓM��!j�:R�^�N�Au�B�	m\��@�� d��^B�	#T�~(h��J�p��-A�O$D�XB�	_��9Q� ��)0򌎔hF B��=Q��4$N�^k�a��ћp<B�	�p�
�KT��\}��ԚCU�C�#Xa2iۢ�#�%+�g0Z{�C�ɂ�Ȱ�d/H�аR���*~C䉜2_����a��J�dPQN��(�@C��$
��4@b�	"=�B5��..�PB�		��}jե�9PIX=2�nҀ/�vB�I51|���3�ـ^�.�Z1IP$-�@B�I+�4��CK!?��ÔM�>!"B�	2H�p��ٗZ6! �h�#1 B��&0K����O�-[�%A�+ՎZ�C�	F*R���O��F���R+N�"˼C�	�R�����ڏp`j�cTg��#��C�ɐHS�e���B�sF�l{��-'�C�	�;�Ju��ʎ�vkusF 'a�C�	�V� �	©K`�m��Zz�B�I<O��f$�J�t�g��.x�C�ɵsJF����~�����Q��C�Iz� �eh�NI�kC�C�	������my
���l[4f��C�Io�8�ɓ����V$U%7n�C��6y�yX D
�b�\�&�ؓ��C�%v��鱃H*r=�\z�(R�?�dC�2�]9��ݬq�&���$r�`C䉔*h2=I��E�� \��Z�L �C�	�|9�(ۗd��pŪR�AC*C䉴sk�U0S.ڔM�f���fQ}� C�I>W�^��3oUB�����B�3H��q��@u(0N �AB��C�pp�n��"x$iu�>_��C�t< ���OV!c�["lnC�	>[� � �܄S�bh3s�WY�HC�	�}� }�S�[�a�}C�	1c�^�r��ŀyX��ec��b�C�	�R=����]n�H�J��Q,�C�ɢW~�ɋ@
���ܡ�dH:3fC�ɭJ�&�"��M�]>�6Ǌ�P)���ȓą�y�l�paE_}�y`��i�<R�� �N·f�����B�m�<��)G[��)�I�P�؈q���b�<i6���1�mB��(R�X�AIJ�<�ʋ� �X)7c@+ K�H�T��Py��)�'=#����!��Ru蔊�A_<?N���@WP`B��C�0-S�\U�NC�I�u��i���4!h�;����ʓ�0?� ~!��(�%^6| p�I�Q��pBf"OfMy%�ȼ>�t�S��0��z"O��:Á��z�V�i��[�S�v�R"OȉZ%��%'���GMC=�p�Ȳ"Oh9Ica($Z4��C,�Lu6��G"O��T��
��1����!}�}`"Ol��U���r4�,�4̇
M|��D^�(��Ie���c�&Ƭf�ha�L�7��B�%j�C��2�F�F�1�B�I>P  �����).��<6�C�I=P������}/DHi�G��C䉣[ 8I���ٻUq0��i�KN$B��5XE�3��L@�2��s<C�ɃH�F�R�0C��Ea�Ҏ]=��3��s�*��j~V�b[;�h�c0D�xr�(OV���Ё��>�����9D�#��߱-�DŨ�-X�(	�F�+D��(��6s!��,<F:4��.*D�8�Sn��{@��'����[��(D�Lаm)`
�(�sH�<@��*6L*D��f�CL���36�R�j2�k��(D��+f��*V��VfO#�՘�$D��$�({|���fA�q��9���=D�`K���2�@@�HK�����"(<D�����sPb�܍p�l��5L4D�D8&G˸T2Q����di�W�3��������pe	6n&�! ���H�P�p�"O:jFD�5��('`������e"O�|y�NKs �Բ���p(2a"Ol�QG# ��ya�mR2y��	�B"O�X�I�Z���cW���v����d"O�r��˕�lb#)�8~��@�c"OPD�Ƀ$P$��N�O�}q�g�� c���=pU�(��4D�$��%��g �b >=j�J D���� $oH��i�'�\�
	r�!"D�<��/��� "�
?�� b3$D���횄CN$,s�JV�;��-D���1�� tt�����/&df�9D� �s#�<k��a����Y�8k1��O�=E���X)b���1nP�r��U�C�͚P�!�d;��	�#}�x�1H��!�dA=8��i�YZS��&�0"�!򤏷��L�g ��4�+���!�$ټ3���E!�5<�D0 A�!���>3�aH�	��>rB��2@�!򄌐4v��;���]���Ѡ֗o�!�dɏS�� �E9MW�	)��ć_�!�Č�-��E��L	�wT���#@�c�!�d\�f�u�#%F7P� Ȑ'_�u!�d\�Ojz��S�=oS����Gd!�Y�3��Lh�"��y>�q1a�ǼUm!��D� 
��72Lr��FN��!�L)}KRdp4�߻4,��3&�9�!�$�F-P5r�LV<{�y6��Y�!�Dһ �@��Q�}d�,[񉄼t�!�X�Ggv�	Q���z���G�X0u!�M,\34�µ:���# �COO!�dJ1
F�)�c.V/�f�A#��B9!�D��m�����M�8Ϣ	�G��3T!�$\�o��C�@ue�]"���,K��IV�����d�4eV.�����La��P�bN=%�!��)�d9�g»4h����]-:i!��D�s�RE�M��h�<��j�lg!�� ,��d�Rv�PGN?N�P��"O>uQ�N�5M~�˒˛�g�(��"O �2��&\�$�Q
W)Z�d�c�d>�"���- ,�X�s�R�
�j���=�O<�|��ݻ#F��=0���J&0u�ɖ'�R�D4�OH�u�� b")�`�$ޒ��ȓi`H��	jٛ�ۖJ�d��M�����ϩe��ICJ�G	 <��&�P	��G��q���U�fP�ȓf�l��k�^��{��U9QT(�ȓn�� ����IelţHG�D��i����<�2w&�<�IV6�Y৊����'ў�>��qb��l\X#��^Y,���*D��"(�)� �ITK�E@	�F&D��T��{�&��-'N�$�c�A&D������a�
{�`�6�#D�x�RA�����:3K*BffMJ�#D���B�p+d�@��J�8E(�� 4���#I't�F�b���;�|H���TA��hO�'M��$u�M��jY)Cm}N�,�ȓ#����U M�)<�F$3Q ��ȓo����YMA�O���؄ȓ90\j� ��Q-N���N�)4�N��ȓ\�z�!�-T?HCf�E�@�*<��@�N��Fäs��g��#C��ȗ'��y��� ʄ>�"��֋�4O���ڧ�8ړ�0|*!�J�)�j)���R�D�1�Wj�<��F��[_d\q �Ъ;���s ah�<1eLQ+7 �W�=y褩�j�y�<�"��!po1ր KB��F��a���^�YT�ˠi�XYB�N�3j�D��m�Z���nԙ��T����u�nG{����O��  �N��A
H @,������㟌'���'��	�P<LY@c)F3(���,�h�C�	[�.�H竓f�3�	ӂ֒C䉸�V)���BQ��B�N�qՈC䉬�f�� |�X!��N�U�&B�I$*�P4a��6K�� v����B�ɷ�V�	v�T�;2|<�V �1O����d-?��퉿ZFS�%C�6�@.CP��x̓V0�1N�%�̱0��O;���ȓmL\�V.Â/:�d0�ȝ[L�ȅ�W:BxAN�3g�z��'( �&�ȓLtđ�tÈ n1���f�-zJ@���R8��k_%����pe �����J�p|Z��7L��KP�N(����p�:� S� U���/��o+Έ��Iq�	�<9%��/8plh劜 \�`DjQa����<���0�XX� �\2n\޴��Z\�<q3,4�d�����&2����
[X�<�1"'ju�%�Te�o¶�{�bAS�<��o��'�a)',Wޔ��6CMO�<io[Y�xI���<2��|�'�q�<9�AHR��ك.�Ժ&2|Oc�$ �Λ%N�v���(B�:��<D�����>b��˵,I5ڬi��/D���r�H�g���k3��'��\��)D�dcr��"t�j����!c�X��
'D��B��;�B��� Oc����O6�=E���9-FM0ŉ�WP��H1!�$��-�0�dDA�R>���J�:!�DΈ^��5k�b
��i!�V!��F��8:�j��n��Ȁ@Ȓ2�!�d�:�����SV �do7�!�� J�ɖ�?s��4�f
0K��{�"O�u��f�$A�Z$�Q�G{0b�H��'��$�,�^�� �5� ��*M!�'!� h��/J��$��?e@�{2��(qKt��l:G�:�$�k��O�QG.�?}�B)  ς&鋇�y��X�4!�t!���RQ���y�C�Ρ�ψ� of�Ч(_�y�/���B��Ǹ�T9Р�6���0>�Q�X#MͰ-�MF��#Xq�<A�D�
�褓��ԿX*�8ʂF�Eh<�a�����4���-��NJ>�?��'����!��	*$��P
�ZZ�'���I�C�?�f�s4�D�ʙ��'�d���O����sу*᮰��'c�h���ݘ ��Pm�'tD袅f�
�@��@*��\���'��,{Wd�	K�Ɓ;�1]�ΌI
�'������d��){���
R�f=)
�'p����הs	(����6+&D�	�'4lP��_��Z���ʛ4�h���'��]�`��>}��Ua�
�'J*d��'�$�YS�Io�9р��$�vy�'��a�ւ_)/�r�����]Zl��' � ���DA���W.�t��'�R!*�;(�ܐ�s��E�(!�'J��1�@��IX�"��-�P*�'|)�A�ѻ&y�tA���!*^u��'1BE�3D�8G��daR4sމ �'��S� B��e"תL��l�i�'�x���1*��iF��pY!�'qv�ߖ8On�ϛ�����'� 2�Ì/b�X��,J�h	�'����lI�.BDE �Nmp�'�8��d�96^h�O�dH}�'��\i�Yv[����G��[�
aS�'��+S�B���y�b��L����'�����;)�>���FAڤ$�'1^MsI�}TB�� �
9�P]
�'J�kV얀-
�� �Gٞ<�����'�� ���~�����,,b*,��'�-�U��H������\*V����'�����_b���a����X�Q[	�'_|����,/IF�i����HT	��'��#+��~#����c�/D�<��'��uiQ,'V�"�Q`�I�D�v�'���#Ц�t-rm`�Րjtb�z�'R������$C��0BgJ�0*&���'��j$��hw��HVB�,�b�;�'���p�"t�.�A��KVz���'|�ݘp���!sU���;�b` �'�Ԥ� ڮ-�^5�Л2J���'�" P�E�H�����+H�X�
�'��D;�J�a�I[sl��!��C�'۞h�cNW�vQ�D�£F9m�,Vh�<�t���z���)� s0��w�<�*H�@-�y�p��1��DjČv�<yV݁T������%ʽ٥
�m�<Q��*@��}bبs^ͨЈu�<���� ��Q��k�Lc��v�<�#�>A8�����U)�0s���\�<AV*1A�`��!�S9wn��a�S�<�i�L:~�8ס��e�&=ǈO�<A�	�=@ �c�N�8x��KG�<� �d��<#��Ћ�KC\ft��"O"���aܛ)"�$B���3S,(�1"O2���a?��T����T&�ԩ3"O�#�G�<ٲX��	�Wop��"O@�&铞Z��4;C�{1l�K"OD�N�D�ΥHt�Ӑ0=&�	3"O�Q*�Q�I���yA�^^d��"OV�j%c]�M��<q�&�
u"O袵 �'���Q�ڞn��"O�5{1�P�m���r3�ެp���T"O�d��M/�Z�Bs���M��#A"O!y�E6E�`Q�R�M$Q�Q��"Or���lH2<�)� �{ކ2!�d��4�X5�L1IӖ����!�^�\��ŖW(:�¦�.[]!��˦u� @����0�Q6E��h6!�$�3(�#g�X:�$Y� �S�{�!�;�=8`�P���T�ŋ?�!�d�[�~d �f�� !��'!�$ܽHv�,;h�>���˔��!�%�f��c�.]��|�s	��!�$��8J�P1�m��M��H�!�D�$Y�oa����0l�(�!�,d������ܤ��kճf�!�$P)Mb`�2GjSfU� ���Z�!��I�����BaԜh"e��,r9!�d@�^���k  Y�"�Z k�.�Py���
qH��pb��.ܖ�tϟ��y2�S,;�F��-J7�H<��!@,�yȳ[;�=1A(ap$+�A���y��Ѝt,tx#JńA�nȚ$`���y"��l1ށ�!�M�D�#�F�y2 E%,����G�.yR�ҹ�y"��	̜�3PaS$G��"ULW�y"�� �n���ڶ�ȵ�$ȓ6�yr%�]׀��P�~1pY���k��'܌ ��T7:⌹'��l��'G�a�'�'��#��ie�l#	�'ʈDid�[l����-�)a��u��'R����U)4<:� GÑ�Mظ�@�'�J1�c�wr��7K׮|[�]��'OH�(�gZ%<�m�F�Иe���
�')��2#.�8OϤ-QE��G�`1�'HT��D�\�ذ��3/gH��	�'��� q7�|Т�y��@:
�'�}IWl��J �D�a�|��y�	�'���EȄ9j���^p�!G�+�y��e���8�bǚ@*�:C#'�y2��%P��%��d2����F��yƆs� ��h�)��J��y���!)���0�˨'��a�%��y"��4��蠎T� w�$�W��yA�)}��!EX�'��Z��*�y�H�	��,�u(Z�|T�+��y""ÿT,RE���D�~�:�͍�y�ʒ*d:�aq�[�p�,����y���W�L��A���f�8���4�y���:3�h5��h��kuD�{�!��y�aη=l��pMܵ[U<b"�Ύ�yҁNTP>��D��+j��e0���y2B@"M�,��K��X��B2�\�yb'܁'�8�N��N|9�cN��y(����ۤi̽��QQGو�y���2|YRA�:'�Dh��7�y
� $�����'f���ǨT�T�c�"OPP�q�^2U��g�(X�$yAa"O���/a>�sEl�1�&ѻ"Ot܋F��d���0��  :HY��"OX�y�O}s�{p�Q�7Z"ȓ�"D�8��qK����0����h D��3`��=i޸��&<�����-,D�T�'�,���d�s�$��i7D�+7�Z�7��E��gŊ"��`*�4D�Љ���*b��1�s�O}z���#1D��#�B�in4���G�.&�x���,D���!����()9� L���8��4D�"���0U�D"U����h	0�&1D���W�8�x�1F�-���!#D��z
V:��ɖ%�4Xp�!D��3@�X+Q#F�	G��?��Ш�(4D��q���T(8TI�%�5��l��1D�1A��)��K��rp8c
:D����ǰ$Z�U���\_�b����"D��B'N�u�tY��L�Wdut�3D�P�� \
:��-�m�)��$�g�/D�p@�ME��Ҍc�#��)pc�,D� bi����AU����Ń�&0D�(��E�Mè�5k�쉂�#4D�<k��Rgv���Q�f�q;�! D�|�e�ة4���A���9Rx��Y��2D��2�G�?n��A�u�A$�
p`0D���$OƧh�8�d� \ ѱD).D�P�Fl�%� G��(V�aKP�*D���w��Y���4dK�[<9���#D��{p)K	@��/	$f�-Af�"D��p������p���?D�@��_!�Z�CI��Z���7�(D�x�4!�PYH���H7�LJA�%D�ȘċP!][`4��e�*�|��!.D��¥���m�&�s4��
/0>���+D�|��Θ����<t~�Q�gl(D��8�@��"�(T���"��9C�$D�̋�(��}!�X� U�^�����"D�8*��!u��Y�w�����s�,D�ذ��Q
q���È�$uo�x���(D���g-��;t�8�0�؅k�z�dM'D�`�J�a�����!0H�&��R'(D��慘Db9O��sϺ H&'D�p�≈�E�Н��B��ZÎ<Q�@&D���'�jϖmSb$��]'�%D��Ks��T �Q��L3ADd�4�9D��hU���Q�lx�EfJ�B3`�6D�@�B�h����H�����*D�x+���1b(Ї�G�wT�Bw�;D�� �\"�@Л���'`��J`�5D����)�yjHZ��&=����H4D��A�K�Z�ቱr枈���'D�P`N�}��eS�G�w�V��QK&D�\r���e�03��V:i!@��#A#D�����ĆV��J�	4'?fHYci+D�Тר ��ꄃ��6О�Ą)D�L�Q�Q�Y�N�;��1O�&��4	&D�L��20j�!��K"3y�a��'D�\:�b�
w�t+��=�)cv(2D�H8C�^�YZ�� �
q��:�#/D��z2O*$��a���"GKL�B!��u&�P��R>kָ��ޚq�!�X�f����jH�}cĀ:�钼ja!�� �*��*U��E���U^��K�"O���B�� "p`q�dC�[I���C"O��ؕ	��t�z�@��.G�J�"O��q3k7`v��YPI��B�6PR�"O �i�.͆�45�TFV#�X8""O2��r�ɲ��S [�Mn��2"O��� ��(#�����Vc��"O�ä��&1���	����jZĩ�@"O����*�J��lQ�P&]�R��D"O���VU%!�`s�k�)�53�"O�<�ˇ�[^�����"y� w"O�T�p���AL!�׋ l�̠t"O�t���f���D�H#-gDHj"O����͊@Rt=it��KJ��#P"O��T�X�|�l8*Ё���Qj"O����HO�)��==�R���"O:I� �_oB -K�I��9"O����лL��[ψz
����"O���#j��$�C�H�������"O\�c׃6�@��({�����"O.� �ؒx8�Q�ץ����#"OD(�u �+p̬
�.\&�h��R"O
��။b���.���"O�(�ֈT*����2�=9a"O����F�`,�dae�(pY�"O� �'�c���8"��zIz"OبQ�'�;0V��cW�в�"Ox x�$��D.�S!�#@���A"O
Q���_�.͖|�Bţ2
�@ؑ"O$�#i�RE�5��%]<(��"Oڨ����s@6 �۲a?2��"Op4��섂g�>=B m�(���"Op�t	k�}�#ɅLJ&�"O�-:dF�M�:��G�l�����"O�͸���-�H��u���f��5"O��)EE�)���K�L@�}���a"O����'z1h��Ui�D��"O>��G/��P��bG�U*���"O*}3��<��\;���:P�vY�"O���bʇ�N��s���C.�#7"O0	k�)�m�X�&�D�b��1"OR͉������H���/b�Y�R"O����O:���;�d�B&�9��"OҸi�䘹qV�e��"
�`�r`{�"OjLc�!�r�αC�'w�HE�2"Od ��ٻ$��� �"*j��"O�ƨ�X����v.0
�B���"O�iCtAܡ�pنL392a�"O:y  ��B��M���?/T��T"O��E�ׯ<Ԝ!��"~�4�"O00"+O0l�d�sD�R�x��0�F"Od�K _�a��Qg��P}���"O�@�7 Ai�X�q$F��KI���"O�-�Qk%��u���9}T�E"�"O~�v/ϲo*p-���śO���"O����ũ0�t),��>�DIc"O8��d��oTMjRᅕeq����"OX�:vƏ�;s����l
�@�s"O�p�ۣ6��0p��Lb���1"Or}�d�Q8Y�h�)H��j�j"O@�K!�ܱ�H>#�`Q��"OX8����fE��T
'�PH�"OU'):mΝ�@'.LȀ#�"O�80��S8y�a���1=�� �"O� ��Y�D�}"��#OF.oo�ib�"O0l�'�d�u+2�M)~(�s�"O���0b[�����W���#"Oܽ����*R�fu	p�#�0���"O�p[�j8b(Œ���.���C"O��cvm��ڐ�S�T�_���!�"O��,�yZ��!D�Z��&Y�YE!�ċ�"	�5�7j˟q�X���D�NF!�$+E�4��b?���L�Z!�D޳5�� C�cU5@%Xq
�E	�g�!�@&V�<r Ο=-$^d��-R�!��>�2���Q������� �!�.�� y֦��!��[f
!M�!�d�T�՘��8%پ������!�Ƃp�6��P��s^�œS&""�!���hq�W�U�fE�`�P+�[B!򤖂L"a@u�$DZ�B�L�t�!�K�1{�(���"p6>�Flp!�[�f�z(b�-F��j˓6�!�W��Q�炌+&G��z�O�5g�!�֨�<xJS�!<�QX��J�Pz!�R%8��IPfN(BL���QeP+T!�$�_����G휛47���!�[ejT���L��)З&\!��ܷCL09xt�A�zQ$�����A�!�D��;�(h�vF؟G3����T�!��O�#Zب:����!��Q�;܊�B׭W�/�d�� ΜO!�d�)H���6���^�T�jD*�X�!�	:'@�Cg��m�Z�`P��s�!�d��	�fų�ݻ�ۢ�I�S?!���p�Ќ���^\2�G%'!�$R�$$��敊/�P�!��=!!�\���7s�&A�
�!��\��Q;���\�V�@�$�!򤗔7#�((R��p�
�M���!�VRSnI���(�v��#zs!򄅈&H�3$Xx���cKX�}h!�� �3?�zuL��2���32��%%S!��N�j�R�������Z�ak!�V� ۘ��G %`����X3�!�dםG�Qsɛ����:C��!��"����L�m�Mj	��'�^Q��GA,�z<c�P�w��)�'|� �sf��dh��d�6p�l\�'����g��y�L�7���o3����'�h �S�J�Nk:L$k����'m|�J歁:��4z�b	=\�VA�
�'W�40q��#��XQ�¿Z�<�	�'e����ۻBΒ����[�KZ��'��3'YՊE��)�0@B<Y�'�p�	A�˔i(��B�72��
�'�;�W�e�0#4��>�$D�
�'��H�R��}�a��@j��'
H�����b��`��_�@�'��8��իU�8@3u`%QnX@�'��9i���~�܄@�X��3	�'���R��L8�����_M��'�>9�я����BMι\Ez���'X��S6N�g��A����T�<@�'kRʍ� �|�Ǡ�a ^li�'gv� �� ܉P��^p]Q�'�����ͤ]َ�y7%��^��4r�'3����nK�Y��[�0P������ �Ƀ&��;�������U��!�"O���qEY7S�2h�wո�X q`"O�Ȓ���#+^8��Ѷ�j���"O���-�=*=���Y+g�<���"O|�bw��<4
4ٸU���"OL��� 13e��*�fOQ�$ x�"O�5*q�� *0�Љu�#���"O4���5�����A
�1�
�9�"Oz��,[.[�<!��A4Y[NѨ"O:�A,�L5(w��^>�Y�""O����5,�*|h�+Iİ=�@"O��KՇ�a*ڹ��ᇷ0X��8�"O�[����w|RѺ�Ƃ�cQ����"ON`j@-�.O7:Hs���	� YB"O��1�%��.���ʁR�J�#"O�YTc�)���!Iߝr�l ��"O.0��nH�&[8(���:xtm	t"O���a�fv|5a��̪y6=:b"Ole��3%q��s��a>�a�"O: ��i�,�}Q%��)]�*�a�"O����N��/K޵�6aV�~�Dy�"O��b��
�#ľ=;��_+�0 ��"O*Y�s��[E���2���9c��9c"O�}��^�v�Եz2�_u��"O�����T�n�� �$Y4qH"O��i�gX��A�T T5y1��u"O|5�RnG%I�� � -�� "O�@JA��$H��H����Z+�բ0"O:<cC�P%-^m#� ��_j�jV"O��P �77��|Am��u����"OJ�	'U�E~hYU��(4�d4bb"O2��1ƈ}�p̸BH��.��#"O����䁡!�.�2r�[>ƀ�R�"O�$#rD�
l�Hmh@k�7��`"OBcVCH5]��8���U�J��i�"O��г�6�z���fyN8a�"O$����D!a�.�[�茋'���p�"Oji�um��O�@�AA����y�g��H,rH �ݣM�-��͠�'7&=�f�_60���eEd�
A��'�Xl)5��O ԍ�s�èh�|�
�'$�d(��Gi�X��
�a6�Ѫ
�'�0"��Kw�D���X�-��	��'?:=��AD�^�r�K��dI��'#��~�r���ԓ]~d#�'FhB�G'CU���`��+ �
�'tLH� ��Y�6 �	͌`j
�'D��H1�I�g��2Æ�T���'����ϙ5�����Y�K�����'�jܺ��!��L�B��Z��p�'FZ���#OlFHZ�H
F�����'l$�A�i��x����Ky��:�yr�D'§>" ��Cۉ�ūg�\����ȓm�la�gJL$xU�"h\9t����Ik��X�[g���	��M�6F��!��E��$5��̾8�ֹx�HO�1�����Ɋ ��#a#�LD�\��/?�C�I,�Ĵ���t��X�0��Y*�4�Ɠ��ɳh��Nkr���j>Q^EEz"�~�2#��I�`p΃? $ҩ��C�ȟ@���LJ=:f��pݣՇC���%��F{���G��RW�X�c
��M "�֖�y⃃5E� E!p��;h�<�J�唼�yB� v���!$%cq�0��-���x"� �d+��U���WK-?��i""O6�[���2�<����F8���'�qO07M�U�������}B�Ǳp!�ė�y�q��A"H�Rt���U�D���p<�TG�}J�`��I*i$^�bGO�<�Ul������F������ͦ��\��T�C�9Lb:|�#�Z{�Ι��B$(aS��y�J6Č3$����O�����WaFX8m���.P(��I�y��I5Y�`���Ŏ|,L>���,D�hE���2�F	kwS%I��  *?I-O�=�O"�}f�!bvbL��	,,6պ	�'wz��NK*r��-�ˌ* �Ε��)��<A�.�� ��e�h�T�`�J�Rh<�S�zv���̐A�
ۀM��yb�֟r*䃔�� ?Y>a�U,�yB[�[lČjwi&nrlō�y���'�4TQ$(ԃc��9s'�ԏ�y�$7mʂ���
.n���6��y��$Za!1$�aȾ��i��y�ו��,*v��Dx�xhV��+�y��ߝ+������O���ڐ뀵�y��)�"EjY���XBY>���E|����nL]�����?��Q2�iO�L(���J�҃@�=���@�"�h��q�ȓ@#͓7Aչ$<0Р�	�8��gs�՛3�3yފ5�7��L8�\��� �#�	�|�xu !)ƀ/Z`p��Ӫ�֮ip���M[�;C�`��"O���� �����3$X�e"O�#$H����$���L��ԉ�"OT�8�A�^���)c���bź��Q"O*)r�O�@ň!c� b��bG�'ZqO�`��"�&Z\S#E19�c "O,�i���o�R��E<�(��'e�l��h]9hZ�����\�ժ%K2D��x5F�֢�q���[��)��/���O�c�$�S���'[, �Bǥ��eظ��V�9j0��ȓ���t���``8"(�2+`֨Dz�a*�g?�Fۭ=F�Ԁ�Pg r(���M�<I�	��vq�u�bJv����<i�ˌ<_��H6B�r14�����f�'	ў�'<N:��h$ɫņ��S*����#��K��ʞ!�b)[Gl@�s���'~ў֝O�v��ňۑ&6p[fUQ1�ȓ.��Y`*��Ԩzri۹IJ��>Q����d�Z$�P�GN"BѺ �׆'�B�ɳq� %�C�	o�R��4&�(~w*#<QN>Y�BE�,B�L��O�a�8��A��O��=�O{4�'fDT�N��)�T��tp
�'�Ј+��л���ƈ[99�z0���$�O?�	�t���!� r�1�U-N
!�������O�t���� @{I�S�g b"BE@�'{����ß@�Z�V�� �R�N��(j��+D��Bv��X��p:�GN�q�Еs2E���'��	�EFx�OZ5��,�4Z�=1���yNra���$%�S��d�'0yF,2тŬ4����J�3�O��j��	��ZH4A���3.ё�,D��:��S�S�#�Nu`����-]�ȓ
�ZD��Z�ԐV �ڬ��	�EQ�"~BU�y=��aB�H��2�Q?�yb)Q�3R&�R�m��9�L�"aP�!�� �O����v�(�A��00̠�#F�M�R���@�zM���#5����������ް?� H��g�"����a�+��qȵ"O��Ǭ��iq����͕.�n��!"Oޘ��_�д��@�w}<$@F"O�0��@I� ��#�)l����4O�����|��,`W�,K��#P�I�3�|2�x2�)ФS��J��$���I��y����$�1��~��ur-K#��'�2H!�)擓L�:-35IJ�ab���ҧ@<MrB�ɉ^lu���'ߨ!
Ь]�b�`����O�p+��ֆ�&9X�ɟ�� X1d"OL�X�� U�5��ɛ+ ܌ 2"�OD<��I7-���I��4���6��J��u�����O�8I�F��"��d��'�����'3Q��Y�H�/����C��^9�(����	5)0� ��� *t����
 �Tt��d�<Qam��b2�,0k�=?EN�5A G�<Y���ޒ-�@�L%N7�Ie�@B�<QE%(~H�Q@�H�6?�ڕ��Y�<�Td��5d,a�=�$�4�GҦ��>	�����D:��Iu�+�I2!y=!�D@Lhū$lN6�"�C�į!%!�dԴ�Xu�7b�;�Lئ*Zm!�/
��z�ʑ�+R�P�GA*!�R�(��-:1f�h�����ו5�!��a��� �CХmMP��".�!���p�}(rS٢T��� �!���|tA��*��1v�H;����p�!��	 ��7@��_^�phe ĹHo�'4�|�!�VmNࢰ��	W2>��B.��<�J<)�'b%��Px,
��T��(�Ac	�'����H�L�\�ST���S8`ד��'�h!��!�&e"ǤJ,a�^��'n���d]!l�@M�A�-I.��I<ъ��i��*g���0/�i`��� �O1I'!�D�U�8<����'.�бKr��)!�$��v= ��g�E��q�@�_��ay��	n_��R��>g���w
ś!APC�I5Ti�w���+
a7LB�o�B�I�S�@�a�E��@�`��$Za�X�'��*'O9`NW�Y��m,��&K�Q�l�'�ιH�K>O�� �!l��1�
�'�\�0P������ԎfȨ���6�!�َ`�x��� �$��=��ԩQ�ay�����'�V�ꤡ�/�IXV˔l0rE��y��'�&$j�$�31�-1a �#|�p�+N<!��)��-�L<��&��q������3OzLC�ɴb���MK����&	4��B��<16Z�׮� h؋��N�3E�B�ɿ���[cmP6PZ��Z��� �B�Ɏ] N�����LX(�c�3'�C��UA��(W�~hc�5�B�	�_�JQڤDr� ��n�h��B��#~}J���4{�
��&R+~+�B��(�ȃ%S&f��9c'�O�(�B�I�,�)9s�NH����m[�żB�	I8�}`d���2�z �W�/�HC�I:/e1�c�>[ũ&i��&PC䉄0��$��0(��^3�B�I��N���#�?$9LX�
C	 9hB�I�0�r�3�7|� <(''=2B�	�$���0D�_;zoJ��el��B�/_�n�9���;�����؊ ߊB�ILm�}�G�(��Hb ��X�\B�	2p�fx�]T,�[]���C"O� >����0,=(p��o�>D^�P"Op���iL��ܸW�_�gf�\*v"O��{���=3zR�jF/�!nUzLx@"O���!S�H��%��/\�aD�T�"O=��%u!P��ŧ\�^4���"O|��aO@h��LA�C(m�&��"O �3T�Y�G2��D'5��Ȓ"O6�@qK��vs
	fĒ�"Ǧd�W"OR�����Q�QrEDR"v����"O��GEZ?3'Ĩ`$�Y�b��p�"O.4"G@3Pm&A�u���P�<�Q$"O�Hre�iMn岠 \	T��"O����k�t
�I0 �,r��4��"O8y���LwN���`�N=#a"ODaqB ]�D�`aQ�[�e]4w"OLI ��H)�Z2gvL(�"OH�e�9�`y[���%W��"O����N�r-�L�F����Vu��"O�h��ֽ�+��_��(Ƣ���y��"٠�X�"�<5�2A c�,�yfF|�i�o�' �%2�J�>�yrU�Vި]�ǎ�$��D.2�y�%�QQ�����W��r�x�Bž�yB*t�ƅ�	Z� ��e�2K��y�À X�����E�8X2l��%R	�y�����=��KD-9�r�8�y�.�<IQE(�w&( B�5�y��	 9��F!�	m�prëɣ�y��D�_�֡@Wa��\cN3Ջ�2�y��gW��w�-T��L�d���y�!!*��$PP+PTQ�������yR�	�
�AV�H[̵�N�"�y�� ��T�Kw琇HH�m �H��yb�Θ|?���e��'C�b��� ^��y¦ŋ.�F0@��2�[S�ӆ�y�� �/�@h��3Y�>E���yR��+k�nA�կ�*R�n��g��yr�T�1?�ukB��,[��N �yR`�>� ���Yڀ`�B��y�֍�r�9��\[��<�#f@��y���y�d��ᮔ9 ��@�r#2�y�G�1CK> �5�L/���#힙�y��Ȣ	
0���� :�2�	%���y¨]�x�.H�@�<+�A:��[ �y��
�E[��e
x|��O�y�n� K��
p�ٌO>iH�I3�yb�N M�x|���܊rj�$[6n��y�n�9MG�p�FH�h�<HAԤ��y��x)�u�K�ZWt\ca���y�+�/q����V�X�F٨�BD蕷�y����D�T=�4BN�<9R����	��y��2:��hV"�)7�-���^�y�'-T��L�7�F	�^ŀ%V��y��=$w	�JdTU�d�J��yb��L =y�C�f��M$�y�A��Rb؍k��)2L��
ó�y� �YzEŤ��H�dy����y��p�����C&T��Uj��y2�M�<���jRD<�"1+�����yB-�v���`�Z |p�Dʃ�y��=,�xeh˃T���H
�.�y��� ���%j)BZ,=�r�9�y���w��4X7ʕ(?��a��V�6�8�k'+)�$ּ�(��	��`��o�3e��p��ǉ�
��B�)� �QY4Kv�&�I3Ì�P߾P�ʙ�G���IG���p>Q��	"��[pc��E�p�"�E�dx��K �]F�~����<	A��q���b� �0����g�<�6cZb������9zF$�@G�y�I9|V��;j5�]E�$�N:�P("����@���E�yA�8l;<\&��N�'��6A���#�������?�'䦔�3�DAE��y��Z4$����'~�옷d�f��r��0�:�z��
�|GX�Y�)W8,a|�ϖ�P<��z�L��	}���[7��<i��@�q !�&6�y�$��~
��h�.¼������y��M3	�~,�g̓�,`H��m�4��-dD�Cw-D6h�$���I�i��m�����l<�&*a!���s���Fǲg����'b��U���؀mU�Ɉt�BH��O三�	�8�N����E�,*���"Of�ې�C����K�+�Dƾ<��D��!�p>��ȗFز	�Q��
r؀��"PS������7"���'��`As��K{��#�W#%D��d�&@崽Ps�A(�-�#D�̩��L !w�	�Em��a�,phdg>D���eB��H/Fu a5�FL��>D��i!��;m�ɦaۯ�X\�0D�0q7h�=Zg*e%Rd��.D�@A�%)��`���`2l��*/D��)�햎g��(�qAO|I@-ҒJ/D�y��d�"�;��p�.Iiċ,D�ܫ��@V���!���>����B+D��A�,�nL͸��.m��p��?D��a�D��r9i���m'n=s (/D�(h��o�֬�2&�1ug qI,D�tK`"��K�I�7KS�4�	sD7D�0 c���p�aۢ��>t��XB2D�L2Rѥ2�� "CE�i�T�ђ�0�9��F6/���9�1f I0hlт�(-a~2�T�j���H�0m�8	�ث�0<	m���m@�Eɠ��d�&!LM���/�Ц�7*�!�D��_�Z���y�B�K�ΉL��	>a�3��E9 >m����F�d�QG@9������F�0C䉝w�*�T,�#��8���T���)wj��~D�YN�RT���{b�N ^�d�!奂�E�UPAT��?q4�XsZt����x�r�R��Z�|=��'�~r賗m'�O�	�e�X�tU@������	�`n8`��A��C` 0T?)uh ��(x2�@Ә�(P�bm/D���V�.Eu�%ʦnКj*h��l�<)���Gg����BZ0&/��}�v�˴��ad�ۏt��"��'OBD��1��H/��B��|s���E�F)9�'�a��:�'w5��
H�8�iԡ}m���Ug1���eڈ�T+˩���0���0����fݤ()���z�z�zk�y-*hG�J�a��'�׬�(ݪ��A�d�/��O��4�G�����;��:�|�p��D�\�.T�J� �O�U00��%m�f���!V1{X��� 8}�Iíf�������{" �('eXDa#J�)2��e����ͩ1�p�t�֔6vڢ}rs�N*!�H
v�~sz�)PdU���Q%L�Ї�I�K00��H��� �P��D���L�,iT��C�>d�QI�& pY�b�DR�C׼���5�����8�*j���_������"�H�����F�ސ�B��*3d R�.�)I�d,S���/�X��iHй U	5�s���u��7,Ҍ[b�G9\�z��1��z�Ґ�.��p���z��� I'�aX���<\.ibBi��+��E�� p��C'HD$�3����@ǭRNTi����^�V��'�@%e#K�p��O�	ڡK�l��JD�{�&]	dOI��|���b��e�d��C� ���<H��@ S|y�D"5+��'��ٓL���4*W;D���iБj�IЯ���?�3����F���
�dA���ٌqL�٨Tl�p�� �6�c��[a�*q�$�ĭQʒ�Ek=ZQ ���&OH�
�<O2�a��G��<����n��-�G'����aa�NP`�'��u:��\�b&>����T"�@{�L��D��e�"­��:��
f��1�ד':R�Sr��������7����'lL�b�ƪE����O�ӣrkxUc�g�� aa��\'{TuC3ƌ�r����"O����H�|!�X��Ɗ jܼag<��
 hٶ(A����}v.yI�i�4;��`�KX�j���@>:h�Xa䂁=��`!AM�/��� �&��x
��t��C��0	d�u V��yRÞ�/�$����8��Ye��0�y��וT�|`�O�D���(7���y"/[�o����V�8��=���Q��yrDV�&^vI�[+˒�����yBF?�� A��¯|�Be��m�"�y� :]��$;ĬH(>��kB�~rgY!gG���I_� �P�L�(Z$s�
�*]���T%�@���O.!�����E6dm�Un?,Ĩ�Q"OԅhP������按/g�dr���LNh��3� ���H�d-"%�Wf�va�S��;|�Lq�"O���� Q:S�� ʃD¤~zD 
�+�s��b~� �q^ B���`ީ	� �,�>a�6��`����<D���g�ν cHq�G�U0i}�y҇.�O��+�f�$y�V�.O���@T��9S�y�lA�`��H��,K:Ok��X7�T�p=���o2�W�=٘%l�4�^q
_'Q)Ṇd	0\ �W��1�R�ܘP��0Z� #,O�Y����� �NLp��3*T�)%��Y�)����dMK8��ɣ=F�A���٩KߦL���+nZ4��B[(��l�B�?B���Z���҂C=Lm����Eؘ����A,'(�s�0O� q䍙Y����"C<N�'m���]�g����#n�_& �aJG�
��B�I/-��d�!ުK"S�^�'/T��KϦS���0���s�"E/,��Lz5�_(H([�gy��
G�����)�J�H����p=�A�ʽ,��!��ߟ�s��2zP軔�?�ĉ�*�>62���ļN$�C�ܙ3�����ҍusp ɢ&�>d��Z3lA�9fqOp�1���0�d���'��-s ��et�i���8:,�B� k�n�ۧ-R�b1�C���!A���Yƒ��q�t�ZV�@�y��� l	 �8�	W**gsD�agX͆ R�Ic�L���y���R�2�ⳎB�r9T�kG�O>��?�ू�S� %�ݝ7U�p8g��i�Jt��AU|���e��vtl���D&)��]�6W�p(7g� j��	?�f��&mܢTa�yҰ�x@#?I�ƶk���OF��3(}�v3�'#$�!��|�xɧ�1gv$�@�bW\��ǋ�W�'�`PM���Z(��a?}X��'����^��'��% � ^
g2L�/@(ZY�)� ��*h�m�v����
K�}�tE�$�/��?ّ�Ң�*-�D�]݄�;��sy�$�OjQcV/��R�`��tȅ'NC0��a�5d�)b�<��xC�L�^���U�؅���9�'`Y""������*樂;� m!��S���XJ�Iܬg�<�3A��s�61Z1*̤���OY�9��H�<�P�$$�Ȉ	�@�*ky��Y��c�'b\bl��n��',��4�ǃ<�H�S퍤@
��k��0az0���A%9��`Z4����h��$��Pa�eV/]j�1��bS�:��-�t�2s���ӧ��&�#*:9�s.�* ǂDqZ -�����4:uM�T�(HR2)�R<q���Dn\h0 BL�a��Z`�$)C���LK�B�Y��ɏ	��	�>ļ@�Oܶ)P��3 _p����W�2�����i�֠��vXzժ�жE��#�8I�f)����$T��x1X/�����XIr�҉��O����6�`�Xv�� �e`��	�o$��G��rܧHn4�i%lª3����R'��IV� ��A#[����U�'�v�q6fX�� ��غw��� a�<�6L�
b����'w���8�nƠk�в)��z�*,�!@�u��R֡��xBGG]t��"��?����To?�hO,��Q�b�D5���,I�<�+�#|��a�$���ybg��<@�@��e��z裰V��?�#���Z�X���'}��)��n�>u	��ʍ!�Ҵ@fk^*Q�<C�ɐ4	��5��F��s�h���(q��ug�q��ɀ�����EP%%v���>d$��$�	FZ�↊�)�T
q�U/|����5f9�yB�ļ<��3!�!��]ZuÆ$�yn`��E<b��,dcB�Gz�!`�' �A�M�@QZ��O�5%h��'6�����"VP�zG�ע.�,�a�'��p�/��`tDJe�ÿ"�J�J
�'��H)�ӭ��!��⑩�dQ��'�LЁE&u^h�H˯	�I���� ��q�lP'� Ա㠀 /Q�,��"O�,�BňU�5 ���.7���8"O�ȳD#{�]P�aY�����"O:t��iL�L%tp��6d.��b"O��yc��!¤i�䟙l@���5"O4�㇁+h (#b$Y��Ar"O (��N�{<�a��лRED��"O:t��)�"YrP�s)�$9f|Cd"O�A��0d �ԫD�����"O������=�j麵	L�|�)5"O`�pĂX�C�|�g��!.�5��"O�H���z��3�h�Puږ"O �N����Ջ�fb��("O�����Ҟ=���A%�;Pz���"Oꑡ7G�(���#RO��9BLٱ�"O>]��̞!Y��}(��0sf����"O ���Q�|s�5ɥ�ϕnЄ��"O�	��G�/Or�	x3Ν�%�0�4"Oz4�G��������h���"O(�3ˀ�B%���o�4B�Yk�"OJ$Xweǩ��Q��/����@"O�<���ڢ{8��m�4@��@�"O�5� �1��4�j��!�12$"O.���ճi�6m!���%*���"Oj� ��\ARtj��ފ<�����"O�����ΚMXvǛ�K����g"O��!�GUV�x�L��y}F��"O��RW#(_���NڣnNY��"O|����':��hi�cD�m�<(8"OB�[�c��1�ec�ǚL�fIc�"O�5�ro L%�5��d�&OBt	!!"O�P'��!�t��@7F>��"O�m+2��[��eK���8m�a4"O���*�l�(A{%`�4 �Q�F"O�����ƾ?B~� EE;7��m0p"O`��L�4R��} �.��r��Yڑ"O���Z�pM�h����2e�,�A�"O
��%h��K®EKp/O�	��	�"O�1*�	�(t�0��̰4|\��"O��2э��̉s��2 b"OlaH�	:~�@��u��UKly�T"O橊���0o��Y6`P�F>��"On��T�ز0	�D
� ��6 �٠"O�E��B��F)�q�);B���"Op�"~'� +�&A,����W"O"hz�aZ8DI�yB��W�E��`�Q"Ov	Ri� )���wiޑAqV�
"O̝�u�]� ����iە}cx�w"Oδ���>y�J��"�Ό/W0�"p"O����R�7��]���nб�$"O�`�WE��B�в~�{�"O�`V�U�xԈ ꔆC�daXE�"O�-�-̩T���KކF����"O��F|����k��R��`��"Oحzu!C�4��hk�H^�v�-z"O�1�C�a��U�Q|�4�d"O`�s�Y�RL���ry��{�3�y��\�R��U�o]�D#�/ȷ�yB�A;�%�f���Z��)��͛��y�L�dז8�0M��Dy񠘁�y�j��8U�����J"A�H�������y��D�UAC��[  B�y���&V���Ѣ�"D��v-ݴ�ybhY:Ѧp� i��H�5`���y
� �U:�ų����"������"O��§\)J��̉�Ռ(�@0��"OF�Zv��D�DA�3��m�&���)��de�%����<��� �>Ɯd0B K'!d���@]�<���Aj`�����A�,��פ��i����@F�{)���D�uC�����-4f"��ĄĮXi�yҊX,7a,��D��Yh��Pd2��¥�����"�5<!�@�a�py#c�H�2 �>�'
�P��@ <y0��J���0��6��A�r���^C�I2�`P�I��l-k�a�t�*N@���ʓ<S�eʌ�L����oͨ|�A���.Ȝ`*4��q7g�^��0���w�f��I�ut�񓕌J����ɱ�R�p�ղSRԕ��:�v��D�3PX̥c )W��r�I�i
��z�*�)���1���
t<C�	$���fk@�GD"�'K� �ԓO&�����a"qL!�'R�b���a++Z<��%�s�1�ȓb_(`��d�G��8�Q 8
��e§M���'�D��>�f��)	�x��
�bJ1����S�<�`P����B :H�(�^��cpI��b<��$0O��	�*]�����o��z`�z׼:�:�s_��*t͑�:�e"T�[>��Y���1D��w���bd�=s�)�49���b-D��A7I 	:��]p���5�-ڱ�(D��#ǋ٪I�
d��H�@��s�3T�h�W�5(D��)���?�m+"O̼��o�� IJa�\+QZP�s"O ���$�=)#��R��/���"Op%I�Iʛ\�tTD�6
n��S"O���@��0�����a��]��R�"OlD��a�9�H��n �9=Ds"O��@bb�oV�@u��*^p%��"O���A�KU��-9�J��qLTLh�"On�P����3�R���"OX}�R�G	 �H����o�R�z�"O�- ������c�z=©;�"ON����
P�Vl�vጘ@6��
O���2�ZH�X&�x���Ԧ
�
�(���Ğ�0?ٱG�;U��� �<5�>`��dM^��r��ԅ
���A^yB��;�����/s4��j��y"��+pm"4,h��b6��DKe�'��a�k-y�1q��Y�OE]S���;�� $=w�:u�
�'/��v��,}����.5bl��#E	u0��C�'}�m�#�#�ϸ'6&$�������҈-Md=��x3(�"��� ����X.�~�)�B^�i�	,���L��t0Ҥ֊O����eKH<5�G�a��_' 1SwC�.$��`�O�>���C̆Jji�`�I�C���`�'V����Ҏ>n�ӧ+�p��-O���M�8��%
��h���� M��+�7���k��׃SOhTz�f�F<���i�N܊�
��,r���� $!*Y���Ot��Lܖ	��4o#dQc�� W�ɘuVb���K�Fč� Z0Z���dLwPl�[E��-��9�&a�BG�D��@;V ���)��o���ʤ��	>fڱ��!�,M)�2��R� Z�p��ɰ6�Ě�*�m� `I(�(���b�D�vab&eI�\�4�� �j�ʓQ�0A u�:�����5Z�!�N�R���T)��e��ɻK`Px�.�$~���F�*T�0V�<��JD�>�%����~����ɐ}�N܇���KPpe�S������Ë�;}�ͪL�,1���p�*!�UI�.z�%H� �1b��S �_�(�2m�BJG]�Tts��Qr��,{p�^�0iB��!A��\rD%���H&K���z����UU}q�x�Իimʬ��"�s�x1F.�S\嫵D �#�
-�0��-7�y���U���bŋ
2��q��k�;��_�v,R6��'=Z�{�-�~-��>���1��8 E�g*�0<%�tP�J�<�D%�^���-}�O���Pc̩l{� A� /�z��r��T1�ܑu�5��:��7�O^�������i�Ȑ]R�p��FUz�$Ѡ2���d�(p��,H�"�4"�	��H����W���h�f�$���c�Ȁp�����NT��� �9'o�mP��d(�w&��네�u�j=��A�+M��e`w2O�iW�WA��<�F�[?֘t���
!�>��C��N�'� @#r��$/*�'>q���	0;M��v��g���#���A��1(�V(דh6A{�(�u�&I�O]45(��'E�q�T��=v�Ф�O�:inV�#�@mӺ˖띘h���H�B�f��m�q"O�[����`@�`8ӆ�1�D�B�j,����;My�5%� ~[�L����8����=�HyC��I�&Q�I	s�^�{V���x�^$h��६��B��)a,ٛ�y�R�cDV9ٔ�W	��������y�CG(e��h0���v�@K� �yd� )Y��NH�{�@B D�y�@�w!0����՟B�2B �y�)!D�`�L� j����nY��y��/[3P-Ja�"Ow��[#�ǈ�~�*�
�}��I�O��p�q���IY2'V�q�����!:�Ș�f��OR��4�T:�SLޔ�V���"O֤��Y�p�s�kÃ�������Q>s���q��3�H��e��I�	���kc��1M�P�R@"O���й\FLй�kP�ٞH�� 	+��D�]~�!�g}"�$5ض ��#���
ݶ�y"մE�.����J���f�Ew�REs���������/lOv-RA�E(x�La���� ���:F�'CPu�aɰ;����i�VYH&ay�Be([8��J��o�<�+�eH�Y�Vd�=�:��_ܓ�V53�nZ�~9S��i";e�����MLr���	�q�!�d��R��`f`��7��� �ǹH��Pe�p����<)GI#�gy� S㥉N!}��\�@��5s �ȓ(L���#��!^��鐠nC�!�
H��D�:.,����a{��ʚ/��Ȱ��e,H!9�S�p=Q�	WB��\f�D�)'��*#��3�tp�҈ÿk�!򄆔-gT��*W"�EHD�G��qO ,
�C��Y2�d1����>�ٰo��e�<�t��	6�!��D�+v� ��kBA��ybd�<d�D��2g�0��d��>�'�.�	���]�����+��s@���I&�*����Ј`�m�g��9X�hi���?�F!]�Aya}R�C�(G�P���3�R���O�r4h 8`�8�>�Am�#?!�M#5M��]4�	T�1D��+%�����w��/Nˀ��Տ��0��\<h2peJ�>E�D��=x4�
	%%r��+�J�/�y�Ć�~1(��U!Z�w��(����ɴ?�$b�'�9�ax��ҏdwVPYci^E�X"�B���p?A��݁M3�ի
N:�\Xb��z�`���?	��䨓�%.➢}���{�� (�	OPX��Dg�'�R���+�8��d�|�ው�X�ih@&�*&�0hcǄk~��LWI2�q��'��D�#(\J�8c'Խ `s�'�]����>���O�O ��(�?1����׃�%��x�e�����AUKH<AT��t������i\!���WT�dE(ڬO��(�&�� nY��R�'S�אVt�'��.�5�GjӤIa�~")�]DTD�3���䨛�qG ��"�Q:�@����t�9W�>)��� 8�҅)���u��0� ҂Rʹ"?i� *4 H������.M��O5w�d� ���HI剬=��5�C�;4Iay��L�;D~� �H3Ҫ��,���#|N�@��{ʟls�Ō�4O�yC�\0������9C����
���x"�׌!hv��&ت3�aIcCD��hOVе#��������n�)v߀Y�i�)z,��ҏ��y"$�2���p�,\�XA�BD��?)���:�Ѻ�-}���̘+Qn�(8M;�C�I&s�}x6!ފJ�u��7I% ��$���c����<)$���vbe`�7v��ȑ��c���x���S���h���h��/�Zl�4"O�`P��k}�T�f�˼~	�
"OVr@�[��$%`��D�\���"O@�����`�N��'��|��e2�"O� ��a�	��?��l: $�.`;�E:�"O��ID�?�H�ټ  %��"O6DYd#VL��ĺ:�z�0�"OzĈ�� ���Ugj��~8�8�"O��8 )?s��Y�靍Z�0�"O�p�S
¬|�I�d��eWd)�!"O�d��e	$n����
14p��"OX�〨X5[D�Z'_�(�p"O֤�J�,S/T�U0j� �HU"Ob��7�ՠ)O��H��D����g"O�y��#�峂�}���"OzY��Hwo0Hz��6�F���"ONճ�U�C�P�i��)z�b�"O,�j��D5��yx���%�� X"O�����r��M���I�T�e��"O���߭j� PjÞ?���6"O�Xȅ П?h8��#�1�����2D�$��F4@`$�:�
]q)��˦o"D�ā��G�'�:���f_26h)�C�6D�0�fփ���yF��<I�d�{��7D��'ޯG7:4h��N2'Up���7D�P��� D���u`��`�4��4D�̨���
a��iHP�UJ��5D��������i���[�L��5D��P�F�B߾�y�h�$^𺨢0�'D�8BB�U�*�1PJ�M��9�*%D� �f��l.$�9&뇒SZuWo D��"f�K�Qql�8�(�� D�\�$� i�!��� 8��$J1D3D������(
�`Cp�+�l4PgJ2D�p��E�}��]ʰ�.��](��:D�L��B��7����A"g��� =D���j�}>�X�Cޗ\���%D��Q�!!��ܢ|�b� �%D�|B"čE����	�� l��/D��Y���T�f�P�g6�cCb-D�|*!��:'Lժ7�0$Zi�`@6D�|�Ѝ߸����4,/z8(�!D�����`l���m�z^�l��*Oj�T�X�$�� �d�BB(�J���A?�7%9�23�=`��Z�J�"ǆ�G%�$;�J��Y�u��O8"��Ov�q+Tc�!�x
p�˨]��I�tG[7B4d�	 _D��mf���JF�RS�Ǘ5x�j�%U�QTt�t4O|xQ�G�!V[P�B e%���{�� �x{<��UCN'l�Tk�R������dst�sy�dE�r��b�� �S~�����ԝ�uh��V�1O֙�eH��ֈ����M}�R�ـdU"ʶ�FG�5��"˴�
V�T>Y����}�b�3�� 8���0�fֆU���&�OŁ6F�7�4����p>���	�k�t���ݠ6mJ��PLzӚ8if� y4�Ħ)�~��Ė�8���e�<��P�Ri�cH2}���S��S�$(��0|�5ŕ>_�r�B��Ԏ+�\E�r`�,_R^���	'?��ŀ��0|
�L��0(��ލF���:`�� ȶ��.9�e��%����A�EaZ��)�	g3a;!�U3����ZQb�x&#Q6�y"� ����Oi��A'��v�%���5���'�2�C�'͸�3@��v�^R�`�Wc�]�'!>I�W��p�
�c��D�fӂ1��'xp���:p�@�;�eUc����'s4���!��3Z�P��/W6-�
�'��ꀮ�-2��;"�9QZ�C
�'y�I�u
�/��(�`��}_�@0
�'�b��f2��#�-KnHJ��	�'��1b���-���kE��btȌ9	�'Vhl��W�	��XC�O�9Z$NmX	�'0�����2gr�mB���V�i	�'�v0P�I�|����Q�BрeR	��� �<;��5Ұ�Y���	+�"O]�$�,Z��r ��=H��	v"O������WR-�uH ~��y�"O�i��@� hU��Z�ƻb��"O��� �Ao0Y!4��<���("O���ģ�<d����v @�h���bS"O�@�Х0Z���C@�
z���5"O�<��Ʉ*�Xӧ��	WRԺ"OPA�>\7�a�e�a�
"O��Iң�;-\����o��k�xCw"ORd�r���4hC�d�4K���W"O�
E���a9z�af	�
L���"O�I�VKS�^X�S���juF 8�"O�ɲ@��9�4!���<3p�8RP"O2sODո�#a@�'XP�i�"O\��cGG� ۠t���~Gr!*B"O�=��A9n�Yю
4;��"On�K�',��X�RmIXu1$"O&5��˞?I�x
�m��c��T"O�)��)H�8��?P� �"O�I�w,Hmz0�L�����@4"O�\07�ƍJҜق���%W���{�"O��Ǝ�H ��IҢ��z�"O8�{��M����(="�II�"O�	��nYW"�8��!`�a5"O�T��C���0Iɨ5�8�q6"O:��5i
�V��ã"�g�
��""O�12'��B�� �	
/x$��"O���1��l@�	F��XB>Ԋ�"O���GbF*<��P�4�',Ј�D"O�=��Iܩv���T ݯ3����"ON0���� @����%��%�Zt��"Ozԫ����Z��E�P�r���x"OXH���@o	��z�C�x���&"O��Kp����HСc8."}��"Od1S�Л[�D�0�&Y�l�0"O����g_�x�P�+��?.�&��"O��B��z_�$Z��$T ��"OR��J�`�t$� %j!�m�A"O��Xp"�2^�|���	��Jf��U"O��X$��F&plPի4e�q�"OBh#eCT?\bP�5k-�R���"ON�"�'m�>���)�/�h�"O -��D
�t\z=S�̏W���r�"O0��E*�f�nlHWF�>ht��f"O@5{p�W��L�V�Z'pTZ�h2"O�:��V*i6N�xw.�>NDP��"O���5)�ᖔY#��*(J��4"O����L	D�P�[4C�H��u�`"O�ٓ )�.J�s֠ܘQ�A2"O[�#��\z(�P�!�?`*�,#"O>��%�
-:bu����r'd�ˑ"O�S�Ɍ�tf�����ڽ }d9�3"O���cN�R�]h�d�~a�u�"O��9��� <
����W��Br"O�e�hY�N t3��.x����"O^�yf�I�
�\�㎃aM�eZ�"O�P��f2L�j�ƁP�|/�ey�"O.\zaD	�<`$�іAM4٫4"O,�C��}"y+�)ѹ56x��6"OzicgE�Y<ʔSA�A�x0��
G"O�=���*/)�w�_�m+��"O�e�ǋ��EH�	ƥ@��t�1"O����" ��H
NVR��"O� 2�R/�3~�f��w��Z<���"O��
��Xk���n(�D�d"O�Tat�B�J��a�!��L,��"Oҍ�l��^�[m�8W^4$� "O�ɣ$��[��]y�,X�[U��I3"O؁$O�3>U��m>�{"OVHТ.H�T���H�I��(b=�c"O�����75�� *�g^{�͈a"OJL;�NRm�n�����\�\�"O6�ӓ@�Ns�MqLP�f@@!�&"O�T�W�]��� 	�jX[0����"OH��1JB�v� �JB�f����$D���(�q�>y�a��/j@ެ: #!D�\5+� l�6$���f}�,Kg� D�`��5�� sG�}���q1�#D�l���Ɖ��Yfi
�`�t�@#D� �WE�S���{dJ-�<q�s$!D� �D�C�D��)K��L5/�&-���1D����ƐN�h5����s����%�<D�����M�p�"�V���)sPI(D��p�D�%�X��5�S�F&�!K6�%D�8Hp�&ZbQ$ͅ/���{é D�K��6>�N���a�Ru���*D����(e��4 T�]΄@��$D��[wI �^H��X4`�2y\l�9 �8D��Z�#� q��}���fiv\r��5D�x�r'����ΗZ�ЬS��2C�'%:����ll\X�m�&ZqC�I�u��(�SeGjL��qA�t�C�I
O1(�ۤ���F(ॊQS��B䉊7bpz%k�Lt-����(ժB�1�X��Q�\Ob���A��B�I��xUk�#&y���sF� )�LB�I�b�P���ߢdG�-k��?z"B�	�=2��#r�ʳ̲1ʅ�N�O�B䉐'6�	��̫OmV�ۤ/�(_�C��.7�����:��pN���C�I�u�v-��m�5^�L�1�2��C�	'!��@���7m���ҡO[��C�I�]�< Ť;B���`�j��B�I�Y�ؐ��a�Yp���ɟ�m��B�I�M2���&YSd0 #GQa �B�Ɉa�$,bd��4*�Ϛ iNC�Ij*p)P��];���Fo�E� C�I0zP౉�ꌺH�$Yy�CE�w��B�I4V��9$	_<\4e�掂&�B�	�{�,��Cb�=�,�a�Y�DC�I�I.����H��`�ћ�.ˎt�zB�)x���@d z�؍k�/�RB�I2�̔
�J�*b�="����B�	<.��Ah���/X%���-b�dB�	�ppc#E sLN��r#�}�4B��V�t��# d�@��	�kB�B�I>Q@�j���s>�50��bT�C�I�#DP���CF�!P�N����C�ɃPp����aĞ��@GV��C�ɐzn6���a�&L�Z���&m~��ē8�Ni��!�6�`dl�6=J!�1,/�Ty���z���rj��B!�0N�h5!CD}ad�D�j��"O�����%jrذ��̓!���X�"O��pCn��Ա*�HP�oh�Y�"O|`P��5R��ɡG�9P�e��"OL�yR͇q�L�[�#ϙ�� ��"O� 8����H�YܪPJ�M���hA!"O��u+�%%�Y�P��y�|�c0"O<�sPiZ��BX#�KJ?�\]9�"O2��6,�m���
��!٦���"O�e��<o��]���D��� ��"OdЈ!�. 솠�qA�?P@�"O�S3��:L2�5'��#��"O��l@p��� άm��]@"O�P��n�CW%Rq�Θ1�z�R "O�(���i��@�֯;�pm
""O�Hj����{@;�N׺$�"Of��)MR��� x�r42t"O�����ݏ	����ڑu��`�D"O=�qM2Q���A=���)�"O�$�L_O�X!r.�����$"O pz���",i�Mѕ��q���۷"Or@2AlV9}����kB�4�,�"O�M!���i<XRK�jl=��"Ol�0D�1;������ԳUpR څ"O0}���� ��C)	~�3�"O�M���, �Ve�����+:X��"O�A��ִr�4��c̔�c�F���"O.P˓C�-��@��r�\J�"O ]CF�)^���jG���n���� "O2�Q2O-7Ѧ@
�IU(uxLD�"O�U� 'H�8T�D �̧8L�0��"O�1�WƗ��L��W6=�JЋ�"O�Qq�ج�X�Θ!�(��"OR���j2V���!d��"O0a:��e�@alí@
��*�"O| �c��F�l�p�
!�Ayu"Op��N�j��*pJS,o���b�"Oܨ;�ßS�@)f� Q߲ �"OPuiфY�F�PR�^�=�.	�F"OJY9�"b�P�o�1p����"O���P���]xte��`B<��L�"O0��e� �(i���	R���۲"O˰F�<Ay�R���C��X"O��ql :e´�����N���3"O��*�M�k,
( e'�� ��؉�"O�ȄON�TU�5BF�R#< 0�"O=�SB�e &u;���+QK"O��aw��	Sh�����b���"OJ}���H�g�T�Z��ެ�"Oh���@ �`��Ş�5���"OTy�OȽ%&�q)�I�#��PJ�"O�E |H�uڕ" `�.��3"O� �d	!1�T����Q6D�R @'"O����+�\,��Q�_��)�#"O�5��ۄso�iPSA�ZHڝ�4"O��RA	ň �O�>P2���"O2�S7�ڈ ��oкxY{�"O�Z�j���D<+�-N��Ȋ"O� ��6<�&��76�l ��"O`���!ǯGʄa�mO�A,x��"O�q싾8w~0�e�O(�+ "O���g��\@�q�eBc���"O�m2    �