MPQ    �    h�  h                                                                                 �sC=��u����^��U)G9E�ȫ 2F����~6���~k��%ǈ���g�21!l!WJySW@�]�^���jr`�_x��������g��/��6
��D�f4��l=�&�+�ҹj��(q� �5�����oQp�WA�,�ClM��h5��/\�H0��[�����f�z��$�+�kx.,�Zj=�,>R�OC���Ƀ�����Ũk��\ � �h�o��$�~��-)�/�8B/��"�aN���Pރ�m}�XJ"�;�P�J�DM��Ưɶ��e�=������C&S�\H������)�)���`0��e�/V��K"7�L_���k�����#�L��}b�(��bc�����m���Ǵ�z�6��1����H"�>�����=�����tmm8�	8i �ٖ�d�.�Q��8�cyC����\���̬�$�MW�	���%����豄�Ԃ��ߚ���������}�I2�E�W��Kؐ�&�E��
��`��~`n@���s�e;��ڗ�J0f����}��:X~@ٱ�I��O��\�OZ���r1�m����փ�X��u�H�,h���j��i[/}��=�GF���h	����ojb>�P| t�ԴMZV	������ �4�>�2�J0����F|L.�[����h��Y@�d�B.����|6��;�������J�H��x x�/MGJ��Zg�T6�7��r.�/a���}BL
�Y"c��d�5�W��3]�I��xk@�=d�M&��i�hvui�fxSCm�[Y����P+Z��|��2�F�<J,t=z��E�)��91S�Uuܩ��s��\�����0<a�/���LDZ��vp����"�U������A�V�P�0~���f���(E�<��n��!l��'����)\�Z��DZ�ȫ�-�G/��M����0��y��a	?�
�<�U2�|��?�������}������(����]>>uD g�Ls.��� ���; 4��A�hV��f,a�V�Hq��E��+^��Z�wߟ�F��Z
�����'��4Y��~�U9[���� f��~��TH�ؐ��K��ԧ/gv2�])�����1n�m	��1.lw�jL��~��B��ܓ<0e�@����x6�zM��-��eɆ��&NwV�����|���# ��!�7N���,p���fȃ-����l�
D��KB�{TZ�J��Qa�y�`k�j����x�%P!9R	.�2ġ��A���[.�]�	�U�����t4W1��&#�)d!���ں>�qs�a������G:2<��t|��g�n�C\p����P�Ł(F��*�J	�Q�y�Y���dk;��p�`>����1/INZ�5 �<��6�~KH�4I2��e����k�����
�	LB��?s���
�j�r(�v� s�c��Q��fQ�_=`�a��^@$vߥ�8�5�vǫi��P|��lL���4!��_=:�P�HBT��6f�pg$��	��l�B�s ��]ا>R�\��߳`)�Rn8z��Z�^NVyk�OT�T�ߐ��s���@D�֘��R-�Ǹ���:�-�~�{�ۺ�T������2�G-�ߓؤk���9�4"�e�q�� c7�^Ϗ&���3[�[�ʠ��@���a��Aƻ֞C�'ў���H|d�z�ҒM_�Û��%���E�6�簮�b�)/����=�˅�Q`6�Ss�fj�_�[����f35���L�^����:���v�t��}��O��T8�R��j��-���e���{�+��m�8����`v�
b�0�pY�����L�>~Z������,}���g8��6Dt,q7�_�_N�ׁd���C�,��*+�B5�y���.woh�S{����љ`ڲ]8�gN:���Z���Ay�M����஁�6pq#�㆚z?��O�KL�|R��o�&��YSl;u��^���О\�$�O �x+GƇz�e8�A�(�$��9�MqLa#��pV��I� 3�H�B8�;�����v�$p�|��Lp1J�NM�� ���r���r�4�q '٫�JPRB�>&
�茨6��e��H+9y��Hg�?��G�^Ǟ� m#������'�����s�T�0\ֆ�[	I��%�rv�2�)�"�����K$��Ƃ����*�d�W����gt��{uKy���� ����eQ6vb���\>k��Ǉ���G�s�Ӎt,�@����Ou�h$�O�؊گy����J��b��ڶN��
����n����fMV��<������vY�W-�Ј��C��f���-n��ͬ��
l順��7�^ �RO�dtB�b�<z�)c��B�3�W���K�^Ѫ�Ө�p��rf�%i1�����ɿ�N�dq��Qب";\_��w_��F�D�W�g�잡^B(O�u9	�D�'<���:b<GRN"i����c����͟�pE�HpB�J3<����1� _b��K�&�v���������;�O�[o��?\%|ŴuZ�6�Ti��s�>p�ր2GW*�zl�E_�ݼ;��O�D�,HoJ ���"[�զY�q���3�^�<`Ɩ���Xn��� T�'W�h�om4�����~���A��]@�v�g.�	����]D&��7�����b�dk ɨa�����9n��s
I$PXt>7֘��nX%�0 |��	���M5΅���d�C�Ec�ԯ5J���WG����k���!\9��m���I�:J�	�*���.���l���!�A0��H���F7q��C�{ȯ�n럦b��OX<@���u�� �\������љﲩ-���<�j����٩�Д�������C]?���GWI�h�=8����S�(��l�~��.��U��d��ŭ��_o��u~�t�U�r��;��2���0.��Uɛ�0��oX6�����'�J�5��H��m_�f32^�K�!��e��+���g�V>e����.�&@n�����`h���kLV��J���b��{�-�h���Ts���/b���1X5��Z���4������+�6XP���>�7�1D_Nv�.�H�l��R~DFe�My�����	$�l,"��C:� �|���o�UzKE4����'X(�0�)2�k����9zː0�ܻ���4h]@�%!7�/9�8DD��T�.A2hQL�Cm���'��������T��G�#y�rd��0��I���
Rzv�z�Y�kh����g&�~	M�@�E�B���,��>̋���t�O��$�L)���E-��ԜKM��j���,G�E.����J������?���ޕ�[�1��q@Y���'�V���OT�gT��u�������wL����ۃF�o+T�����¢�����<�����y"����ླྀXQ��)(�mH6�	s"��y���Xr./����jc����=O���?����$��o�v�ـ?@��R?�����n��L�*���m�	�D�4�����Y@��5������E���@���#��n;PxN���Ȇ�;�h2��vf�O0����f�{~ `n��h�
��\+NZ0f�r��!���˧����C��o�8�Y�h�_j!��6/%�9�ȴd�F�D�t���7	:o坣>Zc�|;z�O�V1��vZ��d�4�a�2`EJK��.X��f�[�f�FN�h��@s�B����}Z��W��M_���f���x����J�G���5Tq%�@-�.�a��i}�N�]0E
��t">4Ld�gLW0h�3X�r�%ũ@ol�)9h��Cxhiڣnx�'(�VѶ��U�P漯×b|������,��h�9��$�9��qU0ʧ�������x�i<R�/�G��Z
Z�:1���h���3��ֶ�Aȴ�P�V���Sf�( �����	��J>����2\:��?��#��-��ȼ��Ⱥ�hһҽ���ڜ�7[,2�ʜ��տ�����pz}q�p�"�(H���日>`� "fjsI3�ϔ�	���&�BŇ4CǺ�c[������c���oPª�F�d��: Y��*p
�Z��s5�
G��`U`P�S F�~��[�B�KDK�֫���v�ʼ����T����&�h��ݝ�l _}j�Y!K�C�(��	�7a���F��Z�x	(z�آ-�����u)��6=V��m�g_�}��#lY�~N�n%���\�lq6f�J~���'R�D埸B'HVZ��Y��(�Q�kÖ#��w{x�"tP<�2R� r9��ϊ}���.zJ�d󾈷����W� v&�>d\ʐ��o�>��qεB��������2�Ht���g�n�CWc*��[Prc`(a+�*@C�,��y�\�["f����`�$��͈/đ��Ӱ<��T��S+CvI�G�eS\3������
�e7L}��?�*�^�jF�(d�d ��5�f��Q��`4��Y_�v:��8C����S����+�(@��l�_��!T��=�F��c.��v����΋$KY��?�!(B<] ^�������y3���w))�f8��U}N��Y���?���N��<\D .��]�"c��ꩤHG̢��޺o��� ��'�w�BCfc��_����˲���e�|�W1�d^�Y��&0���f�[�M��;'�yn�C��aTK�>�/����P߰|5ұz~�u��h����� У�[����i"�D����<�=h�cٌ�����wfe�������Pt�3P!�s9^��@�������v���ؾ��
��T*g�R�Lj}S&��nj�aT�{�/�Ȃ�{�`��bw��KfT��R����>y�G�E���z<�ڠg�\�6��tg$��
�N灿����r,'��*�xB=��Ҋ�w
�;SvҰ�*�`�?8�B\:gK^�5������u���ʮ�
ap,��`S?���*�nLQ̤Sː&��#Y�uu��,�F�R��\�{O���+B`�zNq�8�FaCw�_��(�Ca^��p����{7H�ҡ�V0�K^��t0$���|����{S1��Mh���8Rl��D��M<�4�q�'t�E�R����j���^f՝#;W9��5H"����^"$ (T;��z�Gξ�D|�X��T�ց}U	�6�%B.�M����������lc�4���_*�?'������f�zu&���v =:��6�h���.k����і"u���,��߮~Q�HV�#��j�ˊU'ˢ�kj�ٌ1��08��s5S���L�q���ݚvM	M1�w���;��vT=���C��C�K��j�<n�Y���5I�������n�M@d��.b��zf�ļ�iЯΰ�����ڹ�☎1�p�Br�	%DDj����d��N�M��FZ٨�N~z3w�źF�����s�܇?<^=�=��lέ�)�<�r�:�uR)����I��&Rc���(�6p�n�H���J��v�^�#�[��Y&���7΀��V]�OR+?c�	\`Ǵ<�6�i�i�g���T���aP*��l3��_�*�;�����}�H*�i ��"�
UՁn�q�a0�Υ!�7����X)��;a�'ҫ��.�46�/���`�V�A1u]�v�-_F���ZTDa_Y7qTZ��b� �����������?I_�'X7	֓Ĺn��,0�r<�(ן�Yߑ�`Ӳ�d:���@:�E�y5��r ��d��ڡ`E� kb<����":�le�嬜�I�l�=�z��Ȧ!�w0X=���hF�}��ۜ{W��]���#���L<�E�����{U?(!��3+�LW�����ԖM�Zz����{4��O>)��a��}Kq]�o��j_��1�c��yʪ�V�}Sy���q~~����s��J��F�ɺ'��0B�t��r<_^�o�d�Zr�[�������;���`瀛����A5]Q� �j��^�z��g/U� �t+��!�4V)������4M�n�������R��Lq�0J4j�bb
�h��dX�s���i� �;��XP�lZ�w�NI��Fj�b(�6S�&�^D=��{_,$_ɋ�.��l�p����F`O�yPD;�|�$�)�"4-:]p	|�'�ou(�K@Z���X��V0*h2m�����t�w��[׬E�]�5h�xc�@��7y&�g��D�vŜ���<��Q���m����B�{�;�w`j�TbG���#t��r�0Gk�@	
���U��Y*7�h<%��bx/~d�X@�V�]5�1L����mtw9\�])��E��_Է�A�K���j��,�IT�������Jvz�tw��i��4I'��x�1貋@����SVs�	�����i@��D��c���wLH$��Y�m��*��4���c�N�}z[�uD��<�����"5bk�rTa�s<ƺ�vm#T�	��,6z���lj.�X����c��n���?��"�"��$!���T:���Y�sܐ��s����I�����e�u�?9���i߸UV�PQ[�'?E���{���Ln6�r��ȃ&8;����IfbR�H��t7~����R�h���t\F��Z�+r��p���	�A���N���)����h5@�j��	O�QT��O�mF�|���r~��x�!�jo`��>5.|v�����V���� ���4ۤ22��J��h�i���� [��/��9hp�@"��B$q����.�/����"�+�����x��7�eG@߂T�lh��[�.�5aX�}��x4�
o�"��d���W� 3S^��1�@*x��:���ki�x�,{�Qij�5��P�?�ò<�(�d����,�튄�#K�9�{U�����	�RM��SQ�<�'�/"����Zg�"��l�K�h���ZA3�P2�8���ft��(�䀛�r�I���t�0��\՛��:~m-]���9����ҖK�+j�u�0�2�>2V9���`.��t}L���� (�	���h>��� �*lsd������Љh�}o4޸��^�����[+�~�{��z���1������\��f
MyȇNg�%y���ItU����E �H~�l�
]{��`K��J���v˚��ӟ��⎊������X�el;g	jB���4���~Φ�>�U�2��K�a�Fx:�[zC/U-� ���V��\?V���`�8��#6J���N�?�1�����f�1�rrF���D imB�4�Z�"e�4 ���/�k�H9�RiGxC?�PW��R�WJM`j�
���%7D.u�Tƿ(�r����*�W'��&�%d��P�($�>�T�q)�C�tź�|�
2�\t�	g(�CRv|�aI�P-!�(|�!*�[��܏y ������a�2�&�`�mE�'-�/?����H<�QI>�I�e0X��:C�y:4
]��L��+?�Z��҂jx9�(� ��/�ҧ��+wQ>�S`�ر�T�vv�8������C_B����{#�l��`�(�!�B�=���~:.��5��M�$��#2-o��KB�ѯ �3����RTߍ��)d�r8����P�7N�hPE��9�r߆"ɮ)|�����D��[��J�}-`Z ]�c�qL��J4��[ir���=y�������~�*y�eh����y����T��&�5�詒[�𭷶-c�T��~C��؞9XS�Th����|P`�z�E��."�9���[D�����Y�$C��_��
�=C�ǎI�p`f`-��38�A�3kk����9^��^���D�v��ө3����TE��R�*jX�.�,�����{��k�#zЈ6ji`�
�b�l&�±���t>t��֠(��u�? g.%I6��Rt��6̕EPN	�ҁ.���y,B��*!" B�^�i�w���Sq+ܢb�F`P��8>r:�3��}�K�2���v�Ѯ7�+p� �FT?vA�yAL@E���F}&}ПY	�nuQ-CG��������\OVl@+=Ez�j�8rk^3��J���*a��wp�S>��[JHa��q����f�O
)$���|OV�����1 TM#�"�S�f�h��(��4�|'��`VR�j�u~���ن��j�9���H��>���^}ɷ �*�.JT��Ծ�P����T���|.K	��%�	>�hR�K���<�6��w���*O;���PP�/Ĕ����u�ZM>� ����6,�v�l �k�6��}89��PE�Iy,)�֮�0��������&�о�������ט���P��s�������,��/8M7�;q�ֺ}vO���D����sC�5����n`6߬�O���������j$d�̖b��zAv�*�i�勼+���z�I�Yp!}�r	�8%w'� ~��J�N�Vu桂Z���$�މwUԼF�g<��S�" �^8�H�+�3���<��:X�RD�H@@�BRc�����|{p��tH�$FJ)e��9晖���0Yx&�*�h��:��q�*O�{>}�\�м��=�6ܞ2iJ�[���
(��*�z�ln��_#�;��;��|�H�ǭ 3�"Q�>�\��q2��i}��2ֵ�7��X�h��V��'M|n��#4q��<���Aq��]�w�HwF�����D�E�7��ffbyE ?����9���ҭ��I�ӓX�O�֎��n\�0��d�C���Ԑ�;�QO�d�*��;1(�a5��fč�"�߶�|�8�'��*�뻭�: n����X�dg�Ҹ���i!(�0�g���`F�P��{8��d�J����4j�<v
 ����֬��jݜ��o��4�_'��������������
�	���s�]�������D^3�^�(�w}��S5�>��2~Y�^�"��Pl���o� E��%�t/�Er���J.k�U�J��t����%?��|�瀶�@�58L	�[�)���M^�ɐ��]����+:�����V���W]�ϓBn���\��L��J�	Ib=����l���	�sm,������Xk��Z�������� ��D�6N�/ι�[��TG��_D�!.��>l�Ĉm�F[�&y�Օ7p$�X"���:8 o|���o�K;�.�k��Xxig0(�2�����H������fe�ҽ䦸Ѷh��
�[N67�<�B��DʜIuG7ʯQ~mi}8�]3-��J];�@TW�G)��#oJr�r0pP�ɘ
H�+�0%wYe�Rh�Õ�]��~��@i3{�x�������y�*d@tC��Q�)a}�E�L��������E"�,�wJ�.��Jс��gd๳+�����k1#��@P���xV���S+[�����k�@��K8�?m�L�ns��Z����b�O�޷l�X>+dy�r�z��c�"����-舸�G��bm���	��њ����~.���D4�c�Ń�3��r�L�]�t$��H��S��6�3�.����T\���p�sT�ܠ�ϣk)�:N�Vs�ω�k���v�EqRX��Y�YCwn1Z��N�>�;��y���f=������@�~��l���̀ \a9CZ&4r���.|���փ�y��%�A�y�hP�xj#�e������F�r �*(I�@��<
�o�t�>�|��ԅV����,��ڃb4��2V�"J�V���ڗ8h[�^f��Dh+��@=��B��-�n߲�j������S�Y.�xJ�=�W�G�j��ʻT�Ӿ�v��.��a�N�}<Hm�X�
��"�A-d2,OWf�	3NK8�۽&@�$�2�/-$���~iP~Qx$Qf�L!����8P\����6x�3v�Ͱ!,%v�o�J�9B��U�p�7�U��՗�.��<Ⱥ�/�0��*Z¶j�:K�.���ƺ��PA>�JP����Sf�"(v(�"@���gBƸbtke�\pl�5���u�-T���׺�]�q�Hf����-��2��%�pih�3��f�'}'9�4��(~���k�>A� �Rsiϊ����x�ܸ9s4y��Y�'�wy��˛��F��e�̪�˟���p�E��*�
����BI��@ˠ��3U�Ʉ�1& 7��~�Ge�*��/�K�0���p�v��´���F����+�=y��lV�}j�%��7ĹĘ��d��-#J⦑s�roxU�z��-uf]�7X��gV���� #QH��u�N�0c�l�R�x�f�8ԙ�X0���2DRjBA>Zj�@�o7ҏJ.�k����z�x�{�PrU�Rv��(�%�E�Ѱ���.pd
�L��-{4���W�E�&�;d�%����>��xq�de�/	�&���2���t-�hg��YCM������P���(�5d*6�d��#�y[�G��7%\�U���J`o��B��/�x��ƘP<@]��^�9�IC��e�#���
���
8�DL�SN?D���f�j�L�(ڒe �GR����t�Qy,m`j���O�yv� �8����*|ڦ�������lC��R|!
��=kPH̙f7�l���$�-������B�eN �Ϥ��#y��N�p1�)���8K��Kt�NgW����T�N�h%�q��3=/DV=Q�ؓ���6T�~����I�%Կ��4�]���8ϴ�3��M5�5b��T�eC�~�]T4 ŎO��&�u��d��[���1TΆ/�}Ĺ����|�4D�ѯ����l�|kzt�@��ϋ�tp���B�쩊�G�İߤ�z������=O��V��$�f[�N�l�^��-�3��q�i�^byl�GQ����iv����w�ŀ��T`%�R}]j3wG�Z	���=�{�E�~�̈�l�`�d0bm���`�@t�t�>o����j �0v�+EKg��6���t���0��NR��u���B-�,]�N*�U�B�by�Hgw@Y�Sl���:]`>�8Y�:](��<����m���F�q�p�O���L}?�
�q�L{Yܤ��&x�WYd�(u�:b�|<��a*�\>"oO�r(+8�-z��8-��y<U�7���a��8p'�9�0�1��HR�����A���*�$!5�|�2���;�1[ÊM�Q��n�	����f�4<҈'�"x�sRS�W[�����T�ٝٺ�9*9�H8g����X^؎� �~�I��>Ǿ}����TS)��w�<	Z��%�贃�Ͳ�!ʮ�NB��j 5��0�*�V7�׫�J"a�\�u����� Qj�:46����'2*k�E�����LfԄ��,�]&��k�`����ь���Kv��a�;�Oq(�3���Mw	F�¼�����l2�M�.�����q�vJ��>�й?#C�?`�`^_n;30�BF�=h���o�Ճ�Ld���b�(z�w�e���������o�r��Up<]Dr��I%��T�[,�К�oN�����[�S�N���w��F�e�Ʀܽ�^3�o��39�u�V<�:�H6R߼9���ݝ c�|+���pN"H���J�)��gx��l|���&ڴZ�é�����UOH*#|m\֪��F_�6���i�wO�o�5'�����*�$ l�e~_�# ;���U�xH�� N�
"�5��7�/qO"&�u��-�G��@zX��;�qې'�l����4��A��{����A��]q�v�c�.�zG�}��D�K=7�ϻ��,b�� �K��$���l��bZI��XE��։<0ni'r0Q�0�^��Ob�����AdpΛ�6H��WM5{z�Ĩ���Z���W��O	�9붏:[���[&��KX�3gۅ�V!cL�0�፮��FH��k�{S�`�ߢr����o��<�ž�|��1$��ͽ���\�B2w�:ԗ�J��a��N��0������$��s��]�S�������Y�9/E��̖2SPyZ�wƠ~4���]��u����@�p�0�)GtJgr2�Ǌ%�̐����m���b6�7^���~R��5�qіj��7�/^�8���3���"+UWS�e�V�G�Sֲ�j�Gn�����l���&9L�CJ*�-bH!���×��s
r
��=���~X���Z��^ⷩ<Q�����6I`��Ú�h�lb�_�T.r��lQ���#�FVe-y���\�$�"*1d:�$|4^4o�-�K62���WX3:�0Cڝ2c��尣��<-�����"�hB6�v!�7osh�[DW�b��]�2�}Q]�m$du�x��1�n��T��QG�5b#j�ruG�0���sp
�����Y�ńhr��X|�~a�@$0쳓=G'&�π�eFt�l*���)�y�E^Ԃ��h��A2�� ��,���C��+�J,�Ozu��_�*���n"1^�[@�����YV)��D�������S��zpsL~���#^��E�jM�Y�v�3��fr"��E����"뒘��4��r��s�m���	$�l�閈��.@����r=c�����{ӎM�'̘�$W<	��r�ّ����O���Uo�y��N��۽��>���5�d���縊�d��	;��EL���������n,�_N����;�i�~t�fƤ�[�7-w~�ֱ�{�;��\|�9Z�rqD��Y~"�wRG���(Ҁ^&�4�{hkz1j�s�������ȅL�F؈(ޅ�s��YmW��oV�>�#�|�L.� D2V�s��W���N4�2ј@J����K����[�
��Wp�h�&7@X]VB���I@瑥lƠ
y��#����x�뛰�G6����T"[�O.�a��}�����r
	�O"���dm��W�k3IXՂ6je@�\�MJb�?%��=�i��x����G����{�P���P��3�,`l�
D*q�9��OUaS:�R�i�H~,�	��<nD/R7��D�Z�b��I�U�A���g�Ay�\Ph��� �f*{�(1�՛=\���Ɠp��.(\]h�0��4�w-�Bn������L������O7�(h2v
�+���N�y��'}��o`�(w��>q� Ss��s��ߞ�����#�4���T*/��}�M[��� ��/����d�F�n�v ��Z&
����c7�[=^����U�.g�l&D ���~�B����|��K���q
v��=�I�z%����x�y�^��4.lq��j8q���������tB��(���BJ��-xpB�z9<�-P�z�ry�ؒ�V�n���ǰ�g4#lf�WZN�A���\�=,f�_ٙ(_ڵXgD6[�B�m$ZEz윪n���Lxk�y��x���P�IR�&ѡ���[*.k!<�u����b�����W&�adR�^��>�D�q�릍�{�� ��2��th7�g^-XCH�T���P���(��n*���ݽ�Xy�&a�,kW�T�ܷ-`*_^�]M�/5�����<{�g����4чI� We�7.��0��o��
?#L.�?�{s��j.�(�1� ߽�y%����GQ��:`�u�J|�vK_#8t����U+�ּ��!�l��k��\!e5�=&c̴����HⅫ�$��Hh�6� BM� ��[��HiۍK�)�'�8�+��FT�N�6�ƺ&�o��|�-�߅��n��D�����>W�3"Ћ���f�g��� ��ѿI���V�3E&t��ؐ.ܰPZ�� P�e]�$�ϭ�J&A���J][�۷��E�
�����&2�9�/P��
_��cq|�܂z�h����ԯL�Ǒ�ϣ���9��&���S7� r�=����==���9fVQ���e��:�3�����*�^=�j��CF�zIv�h��F�;$T{��R�7j9p���2��{�K����般��`��7b�f��L/�{����>j�P�V͟��#F�Lg$�6x��t�����N�>��(ם�e�,x.*�4B�%���w�>(Sg='���`��87��:���ƪ0��&=�����1��T�p]�E��r�?l�����L��r�$��&sLY��u���}��ݹ<�/\ya�O��h+3�rz_��8����)Źl�a'�p����#���H�A������]<��$\��|�/f��˥1�R4M�̵܉hT�^%k��*
4w2�'E���LR���ar������'���*(9e�$H�9����^3t Y�5�dz��꥾X5H�	��T�f$�r�*	�^%s!��X��4ʉs�}��������*�/�C~��e�U��X�u�|��6* �V�	��6�;5��cVk)���s1얳hWԿ*�,_�ͮ�Ờ:�TW���J��MH�<`����΍���j�d��}(���b��T:M��Y�(v��D�vEq����t�C�i����rnP��}�d�'?��Ν�ʩ,�>�d�־b�^#z��ɼ�St���Ӌ�E��˘���pW]�r��F%�<����0�5V5N��i�W3ݨJ�˔{wKQ�F��t�C���X�^.�����ޭ0Ʈ<�l:N�R��ߔ��I�x	\c�[Բ9�Dp	�iH܆�J����ڙ\-�f�&�^��ʀ����@O�Y7��\����S6�hAi �C�*/�Bq�*��Ll�jd_Y��;������|H[�� i"G��m�q�2���(̕��XZ�8ˌH$'C}��n.4�Ȍr�~x�A'��],�>�~����iX[�Dr]7B�����b/�� ���g��vh�=�?I(X��ք��n��0��y���S���՟�?$d���12VnW56\<�������2d�H�3h�뱑�:�й��}КOjҮ�-�p��!���0){���F�bo�b�{n�V�Zu&�|)���<������SHPb�O�����o��+i��ű@E�;ЀD�?Q���$c]�˜�3d-z�T'�2C��/#Sk)^��y~�N����U���������aM6te�r��� �(�˕��,X��a�ۥv��Հ���6NK5���������I^���xC�Q +p������V�4̔�u����n}Mϡ����EL�d�J��~b����ʗ5��s�d�z�܀l;�X��Z�r9\��wj�3ޏ6DP�o���#��}9�_:�2.Mil�Qľ�FQ �ya3ɕ���$'!�"��:�*|o)�oF`NK1��!(X�*�0^�2�٪�ہ%6�����?�n�9h���ۑl7�����D����f�-�gQ�09m�jV�����m��|tT��}G_�#e�wr�\0xsg#<�
>l���Yۼ�ha��S.=~uR@�LA���?�J5ު���H�tH�E�+v)�E|�OҼ�����*,3��@���s�J���
����:�Q	�I�1��@�*���V��Ɇr��h��a���e{���oLd�����~��[� ��b���^m��S��?�����"F[��od�Ľ,�">m�m�	_G�<*��h�.�Ң��vc &�)uߎ(#���3�$������'��9�
wʂ���)�=�s�ٸ��0���滸ES�G��u�E'0��,X���f4n'�J���ȴœ;5���N	f�6������9�~�ܱc&5���\���Z<~rL�������o��/`��(K���9h�G�j�t�n�f�� /�FӾ,�������VrZo��m>�N|'�Ի�TV�t`��D�P��4,.{2L�jJw���ݎS�?[��'���h�݈@s��B�6�$�ˑ�;��-���0��|x���),G�����T]謬�".�H�aiq�}���� R
��"���d�p"W��E3D�6�@[��h��%r�ͯ��i�؄xZ��B�-�Fs&P҇n������#,��*���4~9��U�H�m�E��F���xp<>A�/�q��һZx1�d�����B�A�m�P-�yDf��(�F�X���w�n�<�Z\�m��+�>���-�Q�������'v���F��#W�2gD���|!�is��\�s}� ��_�(�]��ҿ�>�� 9�s�c�π���a���../4�MO�O���-�����t��[��r_9���ߦ2�����
^�ȸ�ՠv�âj�U��y�F� m$u~�]�lI�7��K٧���v\������K^�{o���g�݉�(l�?j��o��̥�/ٷ@Г#e��\���	Mx��(z��-+R(ɭ�)�-FV���q�*�i��#����XQN_ra��i����f�����D�Y�DQ�<B�VZ Vh���쏀�Zk���c��xtU�P�]�Rl��ޔl��S���ӥ.f����$d��jb��ǄW��&jF�dH�	��|>��uq:����:{�2��Wt���g��CCoےr`.P^�(ͿA*,e�ݘ5yѩΈ��R10�7�p`��x�/����|ް<�YV�"�[/�RI�(�e?k���۱��w
��LifO?z<��/j��(P�� �S�~s�[f�Q�T�`��+�E5v��8/>�����]֗��,� lSPu�z�!�ގ=��a����b�O�`�~$7�����5�B�� Jo��.�;�ã+�&%u)�8���ATN6U��u��^���R⮺�쩽�D��d��	x��LN���;Ԣ�]��s�������.�s�I��K/�kr��koe��1C
fj[�Et!&�V����N[���'Ɇ�.��/����*|g�e
,�<z�|��zjʻ�^qo��H��,o���w:��|n�U�ǈ�,��{n�=�F��xD��Z�*fQ�"�L�<ga3�Wc�_r�^�X��U��g�v��&�D�����'T�cR���j����#F�ͦ�{����4 %�g�R`�x�bcDP��-��3��S��>e��ֱO����a/g�>�6S tS1��f��N���+�T����,���*��B|����YwvDgSb�F�s�
`���8R��:S���8b��o��Tx��.��HXLpQ��G?��5���L�ἤ�y�&n]|Y�u��v�322�?\���O'� +.z�z8��F�'TK�RŔ��aJ��p]�n��І�&H�Qq�p7Hy��W�$���| L���{�1�MTg�ܤZG��Z���4��='��q�R	�͆R����J�����9�/�Hn,���ea^�y� WQ�BQp�3pl�D"�T��B�m	8�%.]ȴ����.d�dY$�1)��q$��ȩ*`����DO��>r�R�3u����x �Kz�hM6=�4���FkDr����7������,�zͮ����N��4�־��AEJ�G������i����������8l�LJ�b�M����cC>����v@y�����/�C���VY2n�b���=s3����%ܖ���id�b7�z�pk��6S�:����i�%d��z�ypr}�rz�/%����������N�1�治ި��/� wƿF\�h�~�
���^)��<z$���<(��:ɛR�n5���\���c�Z�����p�U�H�gJ�v��n�Gk����&�(
�y���k�6����O>���ّ\L�V�|i6��i[�7���&]����*`ةl�^_��;�^��;�HHR ���"����Uq�b�:�]�#���H5�X�y˧�'��q�In�4"㣌�Zyn(A�F]�9k���p13F�DM��7����I�b��\ pw�ˑ���D�!�IKgPX{YB�4n80Ǎ���O<�Ee���O ��d�ui�,���!5�]M��$��Pl,�P����ζ�묳Z:2����еs��)��KdT!��0�4���x/F��X�z�{�����gf�Wk�偯<Gھ�̖��rE��+\.�8�����/����������4���0�;5ըZ6��i��]�c��n���H�O\��?6�B�wS��I�mM�~�o��,�� 9�����&I����t���r(b�ۗ��?L��(���d��6	W������7����5ɶR����m�^�v��Ө�o�+�Y��fV�x!��4��'[nx�9�m�G�>�6L���J �;b��Tkŗ��Gs �:��d{�'�qX�i�ZM��f���<��Z�6?`����x�ަ
��4_�!�.(aFl�1��Y�\FL�ny�m#�hH�$B^v" ��:�o�|�o��K,2͚|�XX�;�0y
t2Yo�f�$�`	��7>�ð���";h�'۬'7e@o�U<DͻP���(nQ�m������2�'/�mT�]G�<�#`��r+��03%�>%�
�xv���Y�dh�_��N �~�ct@��z��Š��ޅ��jqt����v)r�$E�C��#�c�7Wf�֗k,n>X5����J�W����
R�� ?�$,1���@!W[���OV���d���E�����@�}��ֿL�����ٸ��嬠≪O�O�酆����C����^5"�C��^c��(_���m�Q	��i����~�c.���uPTch�����l���E$��2���G7B�_C��%�m�oh��е�Q|��t�+!��gOp� ���A��%�E��g���*(�n"�5W+�o�;P��tIf΀z�4FT�mf~��}���ͱ��\��Z���r'���~��aP��S�6���%<h�4�j�t�}�=�Ȼ1�F��;�q���2oL�.>���|by��V�nV�ȉ=\���4G��2�ŠJR��U���a�[�²�'�h\�~@���Bw���a`��c�Tq��Gy�j��x{j�����G,@|NGT�ɺ�GVN.�ʒa�2�}m��䄙
��S"��d�BzW7��3?҃��"�@,��1���͊ai�<x�~��=	R����P���������^7�,���@�9S$U�N��2��>/���p:<y4/�����ZӞ��$����7�\���A�k�P��N��f���(��:�s1f��#�I�x! \A�^�&��_-I�f�5�����oB�	�f�f�2�2�6$Ȅd��נ}��T�~�(OdY�͙>'-= �}\s�?���\��<��iX{4J� �JT��������;���d��MY�.c�A���W
�v�s�����Ѣ_{U[X���> l�~��v���SK5����Ѥv7$��1[���vu��/-J�D��l��Jj.h-����jg'��]�6�x�Mx�}z/ɗ-�e���ȡ�V}���̯-�$U]#��ztN:��֊�s�f�����n��j?Dl�B�&�Z�Q�� =���k�P)��n8x/��PÑR�u��;���������.a��+�͈^�����W�&E��d�L��6�>��q�Z��`��9�K�7R2^��t�G�g�L}C>��R�PX�(��*����s�ayM��b�~M�瞒�`��ӓ��/+ë�W1	<����_*ITq/e������e4P
��L�.?���j�F�(ϵ 
�o�d�6�Q*�`;G�@��v|�8꧋���K���r&�g��l���u�1!�8=��D����ݳ��;�S$r\>����}��B�* ��I)i�>����)P�m8%�<t;NxU�<�胥���r�B������D'Ă���T���F�Ҥψ
�]N庶s��G�q�.hy�)��*�4�PV���Z��)eԒ3~�)$�@�2&���蕁�[:�)���X���N�jȨh/��%�����I���{|���z�;�9r��%e�����ݎ��Xsc��[��%���e=���ٳka���sfL�z�}����3�;x���v^�7�������ov��婟�nű�ET�2�Ru4�j��a��h�p{�yʏ���"5>`3?b�A���\��{���Y>`��a��|ԧg��6.s�t��'�pRN����2�s7~,�.**��BWj��!%wj�S]�b��á`<�c8mj:�c�|�#�7ٗ��x|���{�pӛ �(�?b'qnL,V��Zu`&i��Yub�u=Ժ�d������\�?�O�F�+)Bz�8^>z�c�ƈ�o�(a�5p�������B-pHM��ݳ��RB滱q$Ҕ1|�����K�1l��M"�ܿl��T���*4�R�'{���4Rd����v�.����H[�jj�9�ڽH	?^��˯^�� �'ѓ�*��	�'�� �أT$BY�h2�	k�6%����޺�e��?_���L�;Z�����*�h �+�������;um��9�{ "�֞�.46�h��X'�k_5�i�ϖi ��5�s,�9%��F�q���0���R���\���M�� �A��M��������`�̹���lMx>��0 �BM�v;��O"���C,C���n��C���J߆��9��.Aմ!^dab|/}z�x]�:��Յ"��cjڀᛘ5��p��r�%��}��$�k�N�N�d`����ˍwAN>F7턹�܎B�^$@���M
��#K<C��:Du�Rpw;�4$��@{c�yڲ�poHi�J7���"������c&�l���(�&,��ݹ�O���8\�����6Ȳ@i�,��Υx�D�c*;�lZ�l_���;��d�f��HѲ& �f7"=��ȶ/q �����Bf���hX����'9�
�$�O4]>ӌ�cut��A��]����X���Q�D��7x��*ib�s +n�3Nj�l�-��ֺI��X��z�nzI�0�$n�������Χw�;dAy$�'M-��5�"��}W������[(���i%3���:l�R���2�з�Ҥ]�&�!��0_�ޅFY�B<�{���Pz2�2�f� �<�\H����BJW��7�Fv����˚������a��û����e�����u;5��UV]a��������Jʕ@m����0S����@�~�f���u��m��#�Ɂ������t���r�W����&�Au�b��hEꑌרh�R�"q�,A.5�o��G�0�y&^�E�.W����f+�
���1V`�F���;�hnsa �Ș���L�|kJ��db�8��U��ks�@��0i��:�X��RZ|�*�V���#�i��6:�k�%�������\_0��.�Sl2V���VFG��yȽ�#�m$]�"�ұ:�&|�po|%IK'�d���Xdl�0�R;2�P�Atށ�����A:�$Ӽhs����Z�7�����Dݥ��כ#z�Qn�tmU��������~hTC��G��#[&�r��E0���Y.�
4�'��T�YQhC~Y�I�~+��@U旳�i���`U��t~�����)�.9E�+V�>� Ҳ�걩�,����	��cJJ=�{�r��%��L����e1,@��D��9eV:�F?b��	���W7)�+5�+:dLO�%��Z4���/����ʅ�Ę)]���w��GO"�K�wP������Imj�Z	��=]�y��.Q9�0��c6�h��{�����I�$(���揕٢��m��@Y�������܌4����&k�������)�׍����Eݍ6�l���	�n�pu�*%�;k�i��c�f���o����~⿻���l�\�Z�xr#д
/N�H�zeґU�e{�h�Aj%XΧ�x���VT�FɊ�ޖ=5�,�V�*�oǢ�>|5|�?_��V��,������r+4b�~2B�J-�~��_��Zw[��Y�h�xh�@�ghB����"��V�@���9}���G�x6����{�G��W��TӰa��$�.�l�as}(���(I
z��"`�0d5�W��a3:?��G/"@�����d7q�e#mi<�x�#�8A����PH���9_Q�it�9��,�D���9�cnU��1䣗V�7����T<�G_/#G�N�Z.,L�][�i�H���g�A*�JP9؀���%f;D(bw���l��~!��$ZEWJz\����!v5EC�-�ؼP�׺nX�݇�R/+|"f��!2A9�\�ȟu��R��}��� ��(ꊄ�ȓ�>�f� ���s�;�v܂�t�ܤ��4�Pj�E.��J�~ʆ�#E�Q/s�(s������A���Y
t�.t~��S���t�U6/��	 ��+~��/��hح��KPe �v2$v����w
�Г�q����P���Il�o_j�ׂ{��ĥ��E���'E�Ϡ!;x���z���-�3�#���cJ�VxB��'�а��g#��<~��N4 �Xb���f��Q�92Y���vD�6/B	��Z�mМ[�W��h'k��� exꮎP��RbM��t�1x�,�?.\�Ɔ}7�ڠ�1&�W��& 
4d��>�/�X>��q�A,���Tq�029�t �g/�C9��(e�PԵ.(�?*"���N��yG���!MH{��`[�rӮ�/��s�2��<,֏�X��%L�I��[e�2��(�y���5
�8 L���?����/j?�(�� 0�lꑂ�ةQe��`ֲ@�;��v\:28�1�3o.�x��M�G���l�ݐ�p:&!v��=W��Wm�X���$�V�95g�x�DB^�� ����d�ڹxp�ܘT)���8�ў�7�NӔ�����BP��O�p�,��FD��X�����D�Mڤ����^�������������$g��T����)������e�]��6H�4�;�@&R���PM�[U ]�.��^ĥ���� 4�����|��z`����`���b�ȣ������k���>[�q�<=�������fG�A��9��� �3�?��Ua�^Δ�3�A�Kz�v�o ��h�l�gT�!BR�j�>K�F�,���{�����.��ݷM`3?bY_�mS��,���r�>[o��g����N��g��+6	�t���̜J�N�IR��p�.�y,�ޘ*�c>B2.E�4�dw���SX�z�)ܸ`�^8�Z:Ib�W�u�rb#���tw������p�JT�C��?�p�L��Lg�m���e&d[�Y�Бu����	(;����\*�HO]�9+$�jzp)�8��Ah�Jy�a���p��������H�q����-}��+l$J{|V���;u1���M�� �ڞ%��%c�o94(�'����AR��_C2��I���@	t�E:�9�H�q��Q�^D�^ ����2-ʾ�E���7T��g�c��	��b%�4����Ĳ����:.���bt����*��t2����#�H�uH�	t�2 �k��W6�.t��skz��䖳�D|�p�,0ծ����� ��M���7����t�;��ן
T����u�A����+k��X|XMS=��=����v6�l�iDХJKCG���LԵn�fU�.��&C���!�۠+�oߖd1�Wb�G�z����Q]�p���AG��~��.p�)rp~�%fUk�G%���VNzc��h,b�?e!#w��|F�����)��^�$��@��a��<^�d:�n�RK��oU��I_c��7�J�p:	H-�SJ�{>���♽�8�7*;&�*�/���#���lO4����v\�S״�%�6Ç�i� �[�(��'���*�l�:�_*�K;�~���YJH�= �HA"��գ�:q;#��p�������8X�����O�'�np��Mc4��V�CFho��A8]][������fu��{MDäv7F �+ b@�
 �:��N�J���"�άPI�i]X����u�nnՔ~0=�ʣ�K��;�[΂��v�dܜ�"�gq�5g�����F���Ç,�+7���W:�T��G�c���E���K!OU�0�Ѯٲ{F�g,�	3{�Qi�ˬ��O��[��<}�N�ޜ��A�y���a���.h@��Ǉ�6h���wö��V��б�è�`|�_�]<���}�KC�EX��<ูMS��ٯcT~����IɆ&L���|]����xt���r�,�����|�1��)E�Ҍ���/��#ه�=W�����5H�т{t���^�4���%򸂂�+�ە�wHV;`<�?R����nn#�#�[����L9IJ�b�Cu��_��bXs��[�����tX�LZ�AYʉV�(����65��΀@אT�8Ώ-_���.�J�l=RDď�FB�yrB��޳�$x8s"�c:�| K,o��K"�ؚ2��X��0���2O���O��U	�m��Ŧ��h.���y7[���A]DC��P@���Q�m?���)��n��jT~K:G0�X#Vmhr� [0��HtW�
��$�w0�Y�b�h޼&�D�~���@c���͚���;�FQ�tSh�b�)(�MEJ3��Y�%�-�c��,��RQ���bJ���;#�@��z�����1J�l@W6�ج6V��F���$���ү!���<�f�\L��.�����s�(ݬ�Bg�EI��<R�O�y^"��Pe"Wt��Ԫ�_ܺ���mE��	���|�t��.�l����cQtF��!��]ū��$�*=��.\����ն��[���e�����ǺRϪ�!�Y��y�vq3���ے���E�lF��&�`Un#��߾��;�*z�j��f�to������~ݿ��t�"�'vr\�C�Z�l�r�W@�E�ħ��9�u0o��G:� �h�n�j~�3��������%F� b����l�B�oB�t>W��|�%�Ԍ:�V�7���<	���'4}�2�r1J$���PX$s7[����]�h��V@�UiB�������Ѡ�X�x�� �x���U�G"�2F
T�ܬ}�.�.�az}���`
�;";JdYGWm;�35�"��[a@�{�F �ɢ�@�iw��x+���3�n�W|P�x�T�k
G��1,L���vB�=�9	��UM����4`x�u��<�z/����<�Z��tN����
�-�ߥ�J�Ae�,P�ݪ��C�f��([���ǐ��ߠ�����h\w_�����F-�=�k���|w�Ҹ���� ����2xo�
vȺ�q��) }nl�[?(���í�>ݿ; ?g-sX���{�������4�,�@�%�>Ϻ9�� *l��{���2���w(|��Z�
o�������E�u�U��Xg	 >[~�n,�X�h��KkBp��ov�K�58��r�l�D���ݺ7pl�7\j$�l�VC��s ����8z�mC���\�x�N>z%ց-����^>���JVs�F���#���?N������:f�;G����D�qD���B�_�Z������ˏQk�J�t�qx��1P�Y�R�D�o�ߡl:԰ǐ@.WU���Y���AF�L��W	RK&���d��w����>ܤ�qKI�֕�oYf�2�2�[tT�Rg��C4�ג���P�3�(�j*��D�)k�y����l�C��Hmz`�A��O/!�'�7
<g�ڔ�m ��I
bep��C�i�[�&
v?L�?K>{�*�j��(�� K�WeK̵��*Q�z`q>��6�v�b8`��NP�A}��(.�ݞ�l$Ԣ�kw!њ,=�� #��2�����$�pԖg�s�QB�+i {N�w\�4e����)��c8R�ȶ2fN.�b�%;���t�h��K�Z��D]�ƿ*C���}�"&��ϢS�I�lӵ�����d���]��	�|�`��z��~be�H��|g;$<�6WJ&����9<[pc������v����J{� ��x�v�e�m~|�T�z۞�����ԛ�!���6�������mψx���#`=e�9�)f�+hfBe�3�B�m�3dڏ�^�+ĜnL���3wv\שU���'ÍT�0+Rk�jz����;����Z{�k��E暈�Z�`N�bԜAH@J�gl��$�>V�������~#gx�6䂾t��7EdN�f�<����,��*7oBq��o>wG�SSᎢ�P`�P�8���:Ā2�2�W��C�%��rzD�Y"pIL�^K�?X�$'.�L��Ԥ�̢&_
vY+_u�g��fa���=P\e��O�s�+ z��8�� <��g��%hHa��Lp.���I����H�@��b���x�q�v$H�|�a7��K�1"�M�������J���J~
4c��'�h'�R�d����d=��X� *K9Q��H?�~����^�I: E)���Zw���Y���y���?TZ�n�^��	!�%_���
�ֲ�1=���i�P�q�@��I*q�Q�/Y��ظ�ÞMu#����� X�7���6N���j�k�͒�_��=ԫ�i,�ݮ���'"�@�=�'�ӊ��آ��0�v���:tҳ��� �ic��F*1���M.��k��xֲv1Q�ѻ�`��CbRx���yn���iDf_�~�Ź63V�*�dLkpbr�zc�1�����ы�? �6<혫npÝ&r�t%AH���s�С��Nu,$����X�7��w7��F�:��/D���#^HؑMT��x<y-]::��R&�W���·��zc�Ѳ��p��HH�aJ��[ꅙ�X:�Ҁj&�FD��x��5p��KO�W�`V�\�ͅ�M�y6�|0il�����
�s*�U!lп�_��R;�>���HG�; �J�"3Q��~�uqv��+��8'�Y�HXF����<C'/������4�T.��H3jA�&�]I��Q��P��TD�Jg7��%�L�b��! ����i�3�b�#���vI�BXL�j�p�Dn0 0��ˣ����Y��]�}�p�dw�B���5"#�/�"��A�ڞ� 4��b��:"l��x���ҚL����!�'�0�!���[FT��Z{���F�n���3䖹;<F�ٴ��X�4�=�|
֚�!��|�qPx�gWñ};�<��l~!������z]��q����@u�'P�s��S�)~�އ:~{�p���������7�N�MtѮ�r�4��l!e̷����Z���Й�G��a�X]��"��5ZA�ѽ�l�>��^�C����=<�+��Z�~��V�z2��qیni���~���o>bL.�J�f�b_����n���s�j����X�X��X_�Zr���f�c.����60P2�ۯ��W�A�_&�e.���lx�f�*;sF=LTy�ܲ���$�՝"�3�:Z�b|[�<o�j�K�(��p*X�-0�B�2�GD��I����7��M�ړ@h���� 97�cTd��D~�����)Q$�0m��C������3\] T��6G˷�#Q�0r<g00d�����
*^n�R,Y���hyL�?6Y~�W�@��~�4�h������7t�d��^a)�GbE[��t��Ҩ���g-�,���R����J�M�����[:�����1�<�@��?��?�V���ҋ?}��MH��Z���`�L����J���G���"���,��z���=�����yw"��K���L�0*'��m �	Kl�s��oxF.�O��cl*L��Ȏ��̿�k$^v���^�X��� ?�v;��U���k���E�E�˫_=�xKθ1f!����y�E�kF���,Pnx�&�Ƞ�;�����]f_����>��~�����\���\��Z$r��ഀ�o�~�B�p��G�_�ۆ�h�j��������Ȍ��F����L젢���z�o���>2:|,o�'�Vܸ�N���<��4���28��J�yE�bn��[�F��)jh��8@�c�B��X��?�̹�%��s,��{|x�Ox�"NWG�58�#TI�+�"�.��a�6w}�4U5��
p��"kSd�y:W�^30y,����@GS?�d|`�Ei��x��c�.g����P�Ro�o�.�D����i,�G/��R�9d��U�+����⯨	�Py<*�/Y���J/Z��	/<��i��O��MBA�&�Po����f�(�^1��B2�t�q�ڕ����\������i-z̩��dȺ��^ғm�������ST2ӽ���#������H��}Ip���( 8㦾��>89� �ls!���l;�ͱx��4�e�;��s��	��;Q�G$��.�m�h�eO��*3
ʄ}Ȥɷ��W����U���= ��~�	�����#�K�?��lS�v��V�p��,�)�gG��@=|�u�l�Aj���1x�*˷{v�i��ȓ��~�9x�!�z��-��ə�kؙ��Vnz�����U�i#��st��N�u�����D�Mf�y��^n��_1D�hBB�+Z�y��b���Tk���ς^x`��P�RX\�J�;����b��.R�z�<V�����g�W��u&�Md4�ļe��>���q�pЍ�����og��2�Fht���ge�C/{N���PJ��(9T^*���s�y��͈3�q>i6���=`��t��M�/�-����<�ҙ���>XIe
5e+z��^�a��$
Z��LUC?�~y�~�j�`�(<+� f�j�$B���[Q�%�`�5�1�|vR8��iQ�������θl���f�#!,�v=�lF�;��N����Es$#�Uo��nI�B� 6.�ؚN"گ�卒�t)B�8튊�-�eN�sRm����A��m�&��>�D�j-ƺuT��5�w�� 0^��߭�G3���G���O�sC;ߖ�7r���Ų��eeS�/���Q<�18P&����D>[��۷�O�QF0���9�T�la���c�(�|�zV�Ò�4x��y�ǘ�ܣΓk�iðA����ۊg��=@���d�����_f=[�����(Zg3(�'�K�^��r���X��vzi
���,����T`�R��jU�-���c�9��{�C*ʠ�W�S�`i!7bO��#M	��*���Q>Q���~��h�̓g� �6�:>t?>���_�N�W�����a�,��.*~*�B��K���?w�SN���lg`m��8���:?�\��ɉ�����z�m~���9p��y�?�cw�HL�r�+(&ZٖY�Gun�ĭ���\�}.O�:�+�1z&�L8��m�e7��� w�a6z�p��z]�S�MH~Ђ�.�#2��L�$�K|�����{a1}�eM@�c���p��%�B4��'LpRuC��]|�nB�6�	��99���H�6�Ƽ��^��u  Z��뢩�z#վ��^�0��T�zm�Y��	|9<%���%�uȝ��0���0��$��x�*̚j��G���u�>��u��S�Ӽ �Y<��CQ6����<�k�֭���_���>����,f5=��]�S����e�B��-c���"2�����ȳ���+Z��$KU�a	9�N��M	%�O����zv,�]`XS�8C}�B��n]���w���3�y-&�������dg Qb���z>P�����틙]�ڑ&�f�rp�=rf�%[����y�<"�Np��樵l#Rfw��F��ڄj���_�u^�����|�ן<��}:���RRn��=���c���� q^p�<�Hc,�J�d7�6���3��m��&�����G�W��.>�O*'�;\8h(���o6���i��	��-;������*̿�le_`�;�+�w�sH�| �lM"��t�Y��q�cꀦ���!����X!&�J�'������z4Z�yk�e�A�[�]������\L��1�D9�7IA#���b�G� \�k���$��31���,I7�X�{��k�6n��E0��p� �Z�1��8Z��L"dD��r���5ݤ:�JIt�<��y?�o��:1w�{T:}�����q�!D��t ���!�{00[î�l�Fj` m�{�O��qߦò��Ѷ�<��#����S�M�������$í�\����X*�2wJì�����',è�
c�U>]���Z�l��;ԮQ���.�S�y
�Y�P~VOQ���\�ۖ���ɒj;���t��r�'�G�\��#h�3�A��4n����Vހs�ゝ��55ZV�����K^�ri�?"Ҹ��+��g���ZV�Ǘ��q��nd�|����*��LI=J�hb:��@�9�<eIs�/m�A6����X(F�Z�Z�����pQ�:�d6+��6?������_���.���l���Ţ�F8��y(��T��$���"�,:5o�|��oM=�K
U��U�X���0��2E���d��L"0��t��Ѧ5�Bh���� 7QZ?��D� ��qN�Qm�lY�l�uv8qT�C�Gfˤ#L[5r���0,	�	i
���-HVYqh���:��~<�@��H�5V5	@���I��3�tO���{R)�wE��Nԏ�#!��B�,Z3���9���eJN5����v:^�5����Z1���@��Q���VK�pU�Z���� w��"<��#JL �����aE�o�d�#�;0�U���g���ia��"%#�Jr�Kz�|j6m���	�E��Ֆj�.bsK�a�3c� z��4��oϼ��h�$��'��̝ٳp,�K�����˂[:՚p߶�=y��p�	}��4��z�(2���"�En�6�S���n�n���R�[�);�83�`s�f:褤 ����Xy~��*#�͝��\(�Z���r�!����N� �k&{Ң�Đ�<�h)�jt�n��"�)�s�'|�F��'ާ�W�]����9o8Uk>�|NR�����V�YB���b��u�4�=A2���J�A�Z [ǲ��y�hHO�@���B�|��k%�������nc���*�xg1��=gGr��T�&O��Pn.��a0x�}Y��P��
�*m"��Ld��bW�N�3+F��X�@Kl�0�N���(�i�j�xa�w�)���(�PyՉÊ�� b��ʪ�,¯����\9�J�U�Ŏ��L�*g�+��<eAo/�v,�x�Z?����B����#��pHAۤMP
I���ZfL-�(��6������NƵc�\��l�bzV��-5{�����r�#�n����M��
�G2.,)��]���h��2e}$���;�(����Ax>�Һ �Ўs<�=��󞨀;�UA54���6(���7��Y"�V�R��N/���S�C=߭����

%t2�_�
�����kuDU�+���Ǥ t�"~������W�K�\h��kv�����y����b�S�����0��l(j�\��1�V ���
���#ՠ94�x zc�-r������4pVi6��8]{��`#�K�?�N�F�	�Y���f���J%����D�18Bz�Zg��Z/����k�Xۺ*t+x�#P/��Rӓ�%�������.M/�Ɨru�Jq���� W�6,&��do�%� I>��q�ҍL� �M!��2�ät��g iC*���9\�P�-(T�*����ߚ5y����a�9G^���a`�3���g/�T�ü�<� ͔)v��I���e�M�yb�Q..
5R.L�Dr?�ߏ��jPT�(�� �"�[䵢�<Qj�`���,%vm58֎«�r�7��޵�SqlZ!��a�,!��=���V���1���$^�
���i�Bo�� �-0صEp�*��m�)<��8���(4N�b(����^�~��=�Ю{D��+Ƶ�!�U 32.��;���IP޺"���3ò�2������w�����ʸ��Ke@~�jiq�4�,9R&c���p�[��'����,��VM��Q��8f�,C���A|(Q`z�!��������3ả�*�Č����S�7J��<�=��ٟH��ae	f8�������&�3CݏƷu^_�����_vu���n�ŝR�T��Ra>�j0d������]�{�;H���4� U`�[/b�w��y������Z��>LX9�x���M��訿g�6�tzZ�m��N�#��k�_Z�,�U*�=�B�Vw����w}@,SIs��:��`(8e8ٖF:�����ˉ#�>�[��h���Ip�(���?N�ݿ�Lg��ƣ�&U��Y��Au){t�����^%�\�|_O.!$+j�z��q8J26������ۥ(aq�4pd��3w30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�ڜ4�y^�*г�j���&|f~o,KN��xslЗH�S��ޣaQ(��OU8p��ӳ�ę^�|�ΡZ���%C�A�R�n�X���<���.���R��_@n^��g���+�¦���,t�_�_��t��T�(�gџ�l�0����G�KA�����tf,�8��'��J}����/rĞA�ɢ��`��F�qX�ߌ�����a����:��дd��-��q��!���7'c����~ZX�ox���\b� ���y�1Mfߖ�E2Gb.�S��^'��I�d�0�s�fz�={���|Y@�.����su@��_7ᢈ^.�)W�{p� �H�>��~νU��M�ز�����
�y�Q��]�����U�-j|@�'[vv&&�/&��΂|�S8G}(;�^f�&�<4�~]��X/�\�4�Iށέm�<�	�▴�����G������Xǎ0	�h��ٺ�n�AhN�k5wȤ�ë��}J�����0Q;Rԝ����f�dJ~
�+*�#��Ƃ�ဏo<c�Ǟ@���*j��J�]���s�\D"�5i٤0���'�{�9u"�oyi��^(Z�q��O2�-P�2[�I��6/|�g�9�3_\
�q��2ʷC�6w����K�'Ls���C\��1=G/���X��G�TK`��l�q�b�w\�%�Df*��X��}�������Im)Y�Q}T�j��%ֈ�� ���:���e5��K��Xʲ��9�b�yjcp!`�%-D"����0F{EQb
��+�ٟ���}�lJ�(��Q2���B}:�fţ��Ty����M���*�l(� /�p�fi�K���xN��S�A��Ta���&8�C���������άL��_Yo�Z�RRTu�㪕�-!�=O��WbR��_n� ^�P�g��D��R�S�,�C�jn4t�a�����g�Oxl��z�ud�����A-���B�t���z®��h[=���/�#�A|u��T�͒<e�
3_0�M�L�7��!�{x�]\c(Y��`6O�ya���m�Np,������6��`(���M���̍e���H�c;������tǕ7�ƴ��ψ�eP��-�Hq�[�X�4	>3-u�����jυ_��B��!�{�`��\�*��jbr�ȋށ�a�n3�zM@I6,gG���<�aS���{3�i�q�c�>��!6��� �HI\�gعK� �1�ă�Ջh�������ŭp]��\����N��#>)"�(� r�kƋ���]^��"-
�/-vF.9�7�=ø�M3�S}�OԄ���E��_�D�#�e9�b7��<i{�������e��|u D0�Z�;���<�D����ݪ��}9V��a��YbE0�,_�쬡��cN���w?�������W���9����#pF��=p��������D��<^�mNQ0ys��Ũ��K7R���3�+��k���j�4
q�-%��� rqIR����M�d�+�vɬ}\��I���������Oc%0��Gyu�:*Z���Q �>f���G S`�g���y|1x��vKB���BSf��T�����zZ:4�K7�;`�4��1vS��gؔ�\��M�df��-nfEn��`�*x���u��QK���N�<�1-鐗���������1�C���º��H�\�[�k�b���5b��t��Y#s����#��Po��aO�Ź4~�'����n!�Ͼ����&�A³q��2I[������n:��S�h�Q�>��~���ni�!G�8�V@S�)�"�^�s�s�����,��){Z���ù�"vZ����~�Z���g���ff��on,$��"r ��'4�s�Ӗ�3|������ol�t|Jj�f�y ��'I���
l�9|��!٫�YMH�����9��7WӑIW���C�������#)\�$0>��M{%�B��ީ;"�&0�$��Fa#:5���9�u�4�f��eF>�0l��U�ލ���!�7��YY�km��3�¶�c���Ϊ���?�X���sP�MW�/;��_���+KB����b��)�h�"��rF4��-4w��Vv��U�N8>�J�_*�lŕ��F� ����;��ȇ��;�>�/�#��ZP܌qo�����9+��� ��}�F��)�e΃��}Z%�K!����x*U�S�`eB�7e�-�eG�*1��7�0	6_�?���������W�C���v����L�v�m�t?��4D��̑=�)�U��K��ڐF&Lŏ�q�d��ǽ��4�����K���^8럇njP��v5����A��\�M�I�����! ��4�����Vx.�(EY�
�g��#���Ln �Sc%�#ƒ�P�V��ZpS�;^�>aԒ�X���;���+�2�u(j[=Z�?�֕�l
w��,���-����������X�8VG�XXlBK����@#Yf��F���%��O\*$o�ұ����;S��Q��c[F\�%(Q�,� '_?q�h�L	DD�[�C��D��؍l���5�mv��hZ+c�����W��Y�N�£LM��=�5�t�uoY��M�sTtǐ�[���I�'_�Vԟu�s ��J�3=pʸ����ާa��i��*�թV�uA4D����,ݮ~�H��P�vG�<����L��.���:,�����ĩQ�v��x[m��t�z�k1B��^qx�7ß�SH�|�`6������d���ЉH2�ƶsb����J=*Gü�]�	":b@�vo��n�(w���v[R*oAɏW��<�}�۲��IF�\�w
l|\Jy�G�h��Q�t�j��+#)��[࿞�H��ޢ�T?��Q"�o�#�YƢ�e+8I�, ��>���M��1f�ў8�2O��=+Ѥ&����}�A-<aGK�Y�F'��8)K�]S��ސ)�u"�ZWGs��:���zx��/�(֐H���`����j�6����/�C������; ��)3�rŐ1+�op��ع Y�z�x삔��な~���]GOSFn^����g#$�a����
����<��8+F�+>lX_��w������A1͓rϚ���&�V�i��m�Fl��~��8���O��2��$��p/�ݨ��!qm���2%8�?'c�>u�AGXQK�Cٽ��x�_��+ *p�g>�T�1)u��WGMi{L����~�ط��!��f�1NTJ�?���3���mŵ-���
�¼�!�fĬ}�k�r�����	�\2D������������(��nY������ˮ���M2�Y��^=YF����-�􅚝�
����b�W�C஛�=�?�է��O��3��9��0R��b��x��k�tUdj�[�瀧������ʴ�iB�o@�j߉+�J	���Va��!N��$-��.Ud�w�K��B>HΖcH[��ڽj�c���d#\Y�W��Ω�(

�G�Fp�<��,�c9!贶@���t��I=T�_~��cp����ł��ʘ���)�G���k�����w���\�1Q%P�Mf7�X=�G}�>3�BaI�m��~SÓ7 6%C�%����c_��H R��Ol�����4��'���>(c%�:-�م�ςl�9�Q��b���+�z�����iF�����R}Ǳ%f���!���s����⫑W*-�
>���f�4(Kf$'x��ї`����o�ai�B����8����Mıe�%�ι�S�O�姍�R iѱp]t�1���Ƥ� iR؄_�^��g�<q�C4��3� R,��Y�w\t�����g�2l�~��" �_K�A�ݹ���t~�P*�������7��/�$�A�,�'0���5�����+�yʳ�2��/�j��(��ɭ�$��꠆�6m���,���j�6��?(L�^M�/,��PxW<��u��c���-�F���B������u[OP'C�u���(�;���3:`�ܻ����$�r\���Gh!&h7`PA�����jo!��u�b�4�n _�M�z6Y0��b���`��[{�m��U�#�P�y�C6�6�u�w�9H�A1g�Lϐ��1bfy�����>���C�����] ��Ю��H��p�5"㙴�����&I˘Vv]ˠl":�/�$�.���7�K�P�ꀺ�O�gu�&��l�nD;/e�s&7l[ <�%$�oȰB��d҉�D������ծ��I��4������$�7V��.�/��b��;�D��9$x��"���Ѥ��,�ϟ ��
��k�rE�p�P;=��k���S�E����C���}���|��sH�R,}v3�N���I�����5�z�h��Q ���R������d��{�*���b��;E����|�M0��xy�m:��xQM�>S�!�����gc��y�U�p�K�>��SSZrT��Ĭ��G����7*R`��k��S���!����,|d3�w-��@n#�a`��ą�JX��'Q����/�d�	�-V����X�K��=5���|��v:Ⰱ́�}k!8��b�5����q���YP������/@�)I�����^ʦU܅��n;tLϋX���y&�a���@2[�ϻ�љ�vn�ng��SX�D������[��� �iv��%��@�2D��+22���N�ն*ȩ���zFZ��۹P��"���"�C��Z�2g@�9f�'�o[Dh�,y"C9ʇ��	4W�ӣ�t|Y4�k�o� �t	� ��d� r˜I�_
y��|���!&�KF���m\�f<7$z�I�5��PK��ۯ��'!#K$�
��zٚ��e��KG�/ 0K��ѓW�#'�/�C u?��4�>�U �>���0��UB��� !g~���q]k:���]���n�ϗm����:�,�oX�\o�i����K��
�;�2�䘫��{�ױe��x�)G�Uh�:����rSs���T��:Mv�lU<Le>��,�����J�̡��t���E��e،sv�>���#ɘ�PI�poٵ�B�9x�鋘�P��eݪޜl�e;좦����XN��*B������}5����en��*>�=7_ź6�E�?n!�����I�UW��R�"����LHh�m4�P?��DF�O�j��"����ڝ�Lrޱ�	���gm�z;���m�O0_�e^E��L3�jPq���l��Q����)�:���[��N ���̤��y�lx���E�:���͐�F�0# H��%K?D�O���RZ��h;+�ͫ���(����:�й�0��K��ά-n�I|�6F=6�&9p��@�k�j����Dk8|����sd�4tռ�&��~E�P8B7W搜�/:!�n�sź��vp�ű��P0M�`�р�3iƥ��ק�qw:�H�_�FXM7g�$�	6��!'kF1��pb� ��??T�-��F��4S!�U���'@33,H��y�'��>��Q?�S��4���َ!$��yn�䆳�����(T`9Fc�b�'5�R���ͥ��k�� ��s>�'(�yߢ���ԉl�{�T%`�3�-�ؔ�ͥ�a�5�z}���+S�z�nمf�B|]Y#�i���fz~7"��M/�@׎���?�DB<��ǯ�T�@�М�}�����I�͔~w�ᬍ� ��i�3z*~
ɜ\�A�Y�.���jG���
W�Ami��@�u^V;�S�ԘhC��QDrk���Pn�U�0m�'t��P4����TC�����T1%��^]��P"$�uo���uA\妪�Y����n��H�I��A�DG��V�x�v,�����۷�zy[;����%Y������$f|I Qψ�I/ѻ��6�Dp]�����Du�,Q^��L�I��њ�Y���Vw�"�6O��.��i�^C>op*%�ޞ7��YE>�	�,0B����"���؅<�Ư|�������J�$����3.��wQ����jJ�F�WH=�V��n_8�혫�-Jw(C�$��V�]u�lQGK�a��_��yd;d�����&W9)�"�_l�D�5����mݏn���f�'���9ࣛ~�|�@ފ�'�Ew�Wh��Ȟ�&?p�WJ>��i} � �Y"�H���OeC$҇+�Q�r.r� �t�E�k��\�Ypz�bH[h]�Z+�-	��?U6���vǐ+'H��z.��� �Ќxl�+��
�0�:�-ס�4��Wp�X�O��iSb���b�y��f+6�E���.���*衕��L?�sEO�Y�{ӽ�|%�1.���k�@�"_�؈���)�T�{�gA O�f͊l�J�U�Aؖ���P�/�d�V?�y�m�����U�6Hsr'��&�+�/r�X��;{�	&GID�������A�<��L]j��/ϷO4�?����c>	$�+�ԬY ��E4/����GC��t��}eJF�@�XO\Ā ��m���J*ŧ�{��)'���>�b(��,q��23����o[I
��6�J��t?��:_��q�A=����Ce�]�s�K'�L�B��uy�8���1�/9<�X����y*K�)����B��Fa\���%c�f��Xg�}�c�I��I�m��Q�����%V}���M�6O��{
��5���㓲�;;����Sc�t9�->-�F�b��ƿ�Q��	���������ʟͱ�y�@�~}�z�fE����]}ن�Te�ޫd��*`����t���f�{K��x�B1��j����a����AC;8{�>>��d���8M��,Q������R���c������LjR�+�_���^ �egg���6	[-�����,�J8��r�t�{�P#g|�l���80�,�A��(8�KtQ%��,�B�X����@C%/=�A�����ZJ�����R�5���b�i/��l����[(�"����z��y�/m	��,��Y�}k6��(�M�ԺLB2J`��ȏ�c��,�@��b���LU�4�t�0�P�͂�Ū������}=3�c܎D��L3��}���!yP�`4ܩ��8j�\�H��gFn���M��6��������U�!{�j����T��l��6fs6 �*�xH�POgX>���/m1���T
�豐�Dm�E��]3���֐΋ҵ�b"v�n��`��뚢�KU�]�u�"��{/���.���7rǸC���ѫOTi�9�����^D�e�7�d<�al���cG�Z"���uD��`�#o֔����Ǟ���]�7�V�3��lb�Tr���,����"�Zܢ����B#��ױ&��I���p�U=�4�]���X�iTA���������z��f�pR�X3L�y��׊g��������B��%r �5�ROkѷ<2�d/���z����͕my�h�Ҥ���7�04y��:������Q�$>��=oӴ&g�y��澎³K�:��qg�S�{rT�U�@���H��&7�/u`I�N�"S'��Yĥ�d�?-��n���`}��,���fQ���������6y-i���4�+�������]��#�:2��� ̔��k���]��5���BK��Y�G��t��BE���J��b���������ojn�u��>�e�1�A&qFj��:y2�m��E��iTn�X�S�Āє$�g-Ȗ��iR���#@�[|�����c��F�H!�|��N�Z�7��C��"��Q�藕Vs�Z,;�g�tf�}�o�`����"���]�u4j�����|,3]���o� �t��r�攊 %SI �
�m�|��	!YP6ف��`�ֹ�t7׷I�)|����� ��r#��$�����OO���1�^�,�>609��ƹc#�i���u��4GK��h�#>k��0��Uu-�{��!Z||��-�k�E0��zd�6.��j8�*]�׿(�X�� �a�_�1Q���=;	�d�k|��f	�D�a����)��vhE�ı-�+rƸ��H��m��vzO�U/h>U�@���\��9%���ă��%�L�2}��f�u>QQ#|�iP\�moL�����9�P�+����������eN�t��^�˵ӽA�B*�zb��'�,�ӭ�\e�;&*��72Em6߿�?�����W>(MeV��k�8L.mg��?n�D9����g���3S�ԏ�˒LE���ދ�[�m�O�`HX�)rS�^���xj�t��++���æDm��;�����fk }�ʡ�*3��x��<E�ܖhL�ͣ�� Q� �%~H���~���&�Z�'�;ނ�;U4��j��i�j�F=��,�(�JZH���Vz�l��9>1�:i�sá����&��P-�8֫��L%B�D״LU�Y�[NF��%�U�~�o@�:�g��Z@XSr&�_�j[���\#j��%*�7g �S?�hTa~	��R[^x��,�B�$-el ��5i�kvr��hڿЍ*���C�Y=���#!q�~��5li}���"�G���Ԩ��8 ��c��'��Q��Ps���x:=��D�6#\aT���F���U����v��z�J�Ү� �:�v��Eט�
��"�.m٥�n-':����nˮ�)��v{��[�~��􂗧��Л��q�)����HA�����H����Jn�T�?�	�j�F۾b�j`���*Ǘ+X5��*��L|��� �����`�������p�4	��H��	�o�RD:`����i��V�65����E���'���ec�H��l4�kD�l�MS[{��C�0^�O�xz��k��͌���L�|E��E0� ��x�* �W�
���i��������EC$r
�	��eV��������Y�F��7$(�S*�I��,��M=Q �$�SqG����+R�L�m���.,��3ѧ�������W����������>VoV�y��Jd��}�������kb�>�Vݷ���ඎ��u���>�oX�X%�<��kI��M�]���4���g�r��z�$sA:��E$����r��clS~9�6����L�:2F7�|iLl���[�ٔ�ߵ����Z`�d����ҵa�TF"�D�Um9�R&���
AqoO&�ha	2��8�3���5��;'��<�ui�1���rn1 )c%��GH�X�y�D;�5
��LI��9Lƴ��s�VJtH4)m��A�)�@9�>Ϣm>��i=� �ss��Jc��9��Lp����E&�ASޑN����F���"����A^����e�W=Ҋ3E"��b���[��-�mh�V��M���ɮ��(��H`?�=��@��7�VE�;���h����0�UxQ��ԣ�T�(	L���δ.9#}@�`�2�y��G����B�P���
Q|�Tc�}ElB~C�O��[NR�LW�R�ؤ
�
Y�o}�������Yld#�ͅr[�W�@d\j��B謃�1� �md��	��n����6���L�ǒ1�b�vM`XH)��'��E��[��Pˣ��-гɬ�ԻM��ғ�C�����-]�����%�&�A����=�~��l��	h�or�W:S����Bn���.�i�Զbڿ��@I�r���%��<��#3y��Ś���������5�P=�Ι"�~ZX\Z�|^�q��^�m=u}�&XR�?�}�I�h�?xk�UF�*�sð9t&x&�_�D��8!c	W�����7�!'��s$ga�������!�Ot�M{$9��f�ҠS�%�6C�q^~'�gp�EڣM�J�9���#+'�Ѓ��F�?��?>�F�a�܋��4�TU��'���,��Ky�t��=�0P���N4��P�zZ�$�o�#��Ӆ��'��?�/F">��(�R��,��ܪ��l4sM���ʿ8������ey�u��`4F�-3l�kh�@�K�9����P�hzo�.��G}B�f�#斑����z=��H�_��kϏ�	�@��B[����kIT�
=�G>T��-���: ��3�������� �bei���*=����Ar�.��B�����W��i��4��;&a��SZ�C�WD��Y����T1qL�]'3��P����ďC7���"$�׍jT02v�K^u�P��+u����A����>���~����Ο�_�_��5��|)x� T�������O[�#o��)%�Vk�!��c�-I?ҫ���њ�����héF�(�wQu�T�^,�H��y5��Ad����"R|�O�ܬ'a|^6�3C�p	H������Y�E�hu�0�M��ü�*����nJ�`��zXJ2�e��(�Rk�v2�n�JBcW��V8n_~��,����w'��$r>b��l�*���?_hdz�c�"����%�9����c�l:W���'�H3���p}��'�*@9��p~���5�>�<��	k�)����t�%\�6w�w�� �7\�؊�
]��O[�e���$�3�0�.1�� pEw�m������zչR[gQ��k�'�����#žt����H�80zM�b��O��Wv+�	������H�d��  v%�X������b\���y?�.f��E=�F.!Z�)�E�t�0�#Ds䪎����{2}�|d�c.����@�_�_�.\�I-�)]3�{� �6�ͩ.��I�[U���c[V��>M��y���by�G4��e���{U�kCD�'F�&q(/�\F��S�(F�GHh�������a�<�]��/.374���9ۚ��l	��FTp<9T��c8i�;kV����̰��A'C	���N޶<���Z�F�ː��*M��c{�4>�����|��PxU�Q��@�h<�T5%���1�F������x��.��g����T�J,Q+�Q{������(���5���"��X�/Jt0Y� �w\rB1�#eϤ�/�ŕ���g�]���lnu(p�q�D�2�7¤�4I�[�6]�j���T_�Nrq/�� ��C�L�a�UK�E�La]3�����&�_]7/�ݘXȸ���.�K�|[�ZkÝ��\�sL%�f��X>�_}iH���I[���Uғ�r%%E��B��d���i����nM�F��/(�)�!ħc���-�%��S�48Q ��5���#�k���T�����h�}([�fs�����4���D,��{*N�Q�N<Y�#�f��K��xLBΗA`���na��H��i�8�l��R����sΚ�������yRA�b��y8C������<R�<�_�^Vg���!�[���	,M�
�X�t����>V�g*��lz���#��� &NA[���t �qm5�A��VTG�n/+A��^��~(�����D8�����r˳W/2�@>�K*|(����7���e��m7=,��R�+��6���(M��M�%z��
��>���;�c�J���^��C_��"�϶�Ps������k�b��3��ܼ���:��ϳxw�0�^!��`�˩X�jPW�vOd�U��na,�M���6�QC�굩����0k{�g��v8���m��|6N����Hw��g��*��z\1�1�٥VVY�rGJ�3
	]�v ����$9��!V"$z���e���9۹]�� "H0/�q�.��c7�ܩ�������OB�?����M5D<�e��7��^<W�*���F�Q��9��j�D�3����Bȧ����k��K?��
V��V�0Q�b�K��Z�[�P��6�H�
��	$ϰ��S��N�볚�p4N7=;��KsD������P5��׊�����R�@3:jKř(�՘a���Z���+�Id `JtR})�*Cd݅l�s�+��̓�3���R��׭Gܕϴ�y�M^e�:��1��Ѥp�Z����3G���YW*�E��+UAn�`@�3�r
4�%a�T��Y4���� 4x�@����3���Ґ��;qD%�	y�N��@�Oxeۦzң��1����E�{�M�d�����1c!i�0����~ռr��n�pST�x�:*Z��E�?*�i�!��)�@ܺd�<��'��\�J��ܱ�%���/Z{2׹LV3"Ft�f����Z�o�g��f���o�4��,m"�8>����4ӈyӟw |Ց�g)�ot��t�� $ n�Ii�
u�|/�V!"="�0�iԦ��W7 �PI@|��La�:�r��>#�o�$��@��������I�+W�0�bя�#��(�
35u���4��N���>�F0�K4U>��d�?!c����k6���¿8$�wq��-ר�X���������>ӜA;�8��q\����-z|��)��Mh�����OrO�L�V��6��vc��U8,[>~ٖ�(fz�U���J?�I����:��j�o��>zW/#ţP�B-o�oK����9t��+����&f��h�Ye�p���z�t��
:�*��Ɖ��U�����eꮥ*:�S7�6�6���?��F�|+��u�W����"��PLĕ�m0��?W�[DB�đ�)���4��ڙ�ZL����"�t�5�v�_��&�����M^Aj ����jL����3��ղ�m�8�%JQ�2�@��/� &TI��5|��e.x���E�)����0$��� ��/%G#���J�� ZC�;'��'�ʒ$!�lɞ��l��B�(��KZq����3�l��S�`C�㟅�<�A�𗬬�7�yz�8��A�BT턴�NY�JF���%%zF��o��p�Ъ���a�S��X�(0�[~[�\,(Ѥ'��� An?z7�h�L		�I;[G���5�ƭM�_liC�5��lv�h�D=��1����jYFC3�L�q��x�5�o�~�H��abk�ԭ�A�ph�'(�ZԈ�{s	ns/=�z��HN?�a}�Π����Ǫ~D�mK�����L�C�bv�ގ��s�5�.��3�t:u�l�W���2*�v��A[69w�]�$�t&+�Dfq��1�p�H$ο	�ԑ���X���uв�]�Kbjӄ��*���ҝ��@bI�RoѶmnee�wN8����l*�+� �<� �ۻ���r�ԥ��yws;��RVs�t.5�M���#/��hA�v��?���s�t�KB�h��΄<+�!*�೔�����(��ɘ�`��1�3m��j,U!7�5r�6�((�GVM�����S���?csfC���ۺ�I�ͱ@������:P�����G�瓔�lM<3e�;�F���Ͻ�L�zT�!1
V`�$��b�j��� vɁ��nk�M?�b6d���Ͷ*�����WF{kx��@Z<��ȝ��8_6��q��H���g�5�Xu�1M}���3�����v]��*�]밝�9+\��	�[��".�?�X���4��&�]�]4"em�/e@�.q!�7�u����;ꋣ�Or����Y���
Dƥ>eq�7���<���$ϳ���б�ҴHIDh֝�s Q�L57�M���?C����=V����ob}i��d��������Q��}��U������G��q����p~�=��G������8B����h"C�Ǖm�#�R7�03�NţHP��Q�l$O�e���Sy� � �R���]d��:�쬵._�MbM� #%�7����0��y��5:?M�?lFQ8Q>��\�Ff�Fg�t�y����F��Kz��)̅S�wTK���H�벿�l��7U>b`7/�s�S�J�����ã�d��-�*OnN�<`5����w��#:QUr��:�X�t�}-!^�I�����ɎUE�݈ȳ���M��L�|kLM��5�p�&�>c|Y[�Θ,�"��<W�99G��Y�l%��_�����lnFW����5��&)m���8�2F"4�G���!inrr�S�����'�b��N�i
�!�p��@�V�ON^̖읕��1� �n�4/q��r�ZJ�C��08"�vU���KLZ�	�g�lUf��xo�Tj�VF�"N����4"�����3|���V�oCLt�1m���� �6�I�8~
��M|>�.!����l��q7� �I��8�{8FInӚ��#a�n$h�Lօ�
�CGZ�ViZ�	0־�~��#r=Ȩ�H�uJ��4�#�� ʘ>#k�0�F3U-x��3��!�����k�V3�k����L��"���	��wlUXUX�ڡ�Mz՜g�J;��#���Ks��2ܚ�)R	�h����-�r~G��e�ۉ%�Iv2KU�=!>!�����	��=��X)^�(���h���)>	��#4��P��o���ͦ�9c��� �Xzmݵ���6�e8S�����@���Q*��I��|���5 �eO/e9�D*iw�7�6���?�u]�É�T9�W���ϣ#�%Lӈ�m �?&{�D�<|�u�Ѝ���V�ȩ6L�Y7���C�?�%����*s�^p5��	�j;%��f��D�s����|o��5%��A 5$O��<��u�xf��E�� � �[����� �EP%6]Q�V*C�IZ���;�3z�v�S)h�!z3����j(�z+Z Fƿc�lB�9�'��Lh�+Hz������}8�̕���%B�s޴[�Y��F�R%%�E���o�H��u��Sǯ��}e[MF�\�l\`�dȽ _�<?�;Rh�o	|s[<��!�ܾ
l�n�5!p�v*�Rh�m؍�|���?tY�r��ꈣ6��5$����w�~P,C��~���b���'� ���9s8I����=��qɯ���a�ʠ����&4��D�|Q�޷���y��/(vT�PA���.%���&��:d�$�&������v3|�[�_ǈ�zy����S_�q�������H�˔�l�� ���Vz��"�������b9�;��Q(*�G>'�A~:bx��o�8�nT)�wz����*��[��9�<ݑ���������wB�G|��;�z�>3Q�@qH���c�)���{���n���?�QZ(閧�#�˞� �+p)�,X���v�w�U�f�iS	��8]��T[+	=��1;�}��
<����M�F_j48a-�]�6��R.�)�3����sǤ�ϴ�ʲ���gHI��)����`�	=���	���9�R�5C�]��9��Խ�+�䪌1cHp/)��Xu�zR}캞}��)~�\*]��F��;�Q�����~��HV�5��
M��)mU�>oF*Τ+v�6X�%�w謵�2pAAi�w���� 
M�^p���P�m���!J��p'Ň 2�Gȑ�G�7 ۷vm��)2]�Z?_Mx>���G����{8����_���8�M��yT��Du���G�yL1�����^/!&c���$&T�5��B��*�C���1���G�9H!U�zf�W���}�r���R`���j�Mc�*��4���2���8M�������>�vMj��Ֆ�9Ta|�4-����բ
����b	6ECT��9N��wr���@��ӯq{ 0�F8b�l���t���8μsk��3�N*T�'��z�@ ���c��J�S��A%a���NܺF-���j�w݉z����^[_,��.c��d[3����/�(B6�G��p�Vl��c=���E���)t;=���~�Oup��J��ޛ?��a���l2٫��=�.q��y�&Þ̘�h�4̮/ѯ��R�\{�l$߷�E����%���i�ɨ�,_�����$ac�Ɉ,���q�8$~�a�ߚ��ޟ6��Ó��BrL��� h̑|p~䅫cw����n�!��Hj�yF��.�8P�B�zg�Z�̥��7��?�>�a��j�`ɋ�2@�)�d�dM&j�V�w�\�v��Z��� ���2�E��Q�D�����|=�Bí��31pۄd�A�PfB�Y.�{����x:�1�������؄��3F<G�i�Y����`+�QA�^X�3o��485<�WS��W������f@0����3�P��J�,�`D#����N�3>@0e��+�a|q1�����{�p�"��fėߜwVޞ?��Y�hU�����O��-h`KIB����!OD`�JE��K9d�xQ�����b�M���f��� ��J�eq�N/����������c�����C�X���N�;N;�3�B�`
���S����_I_f�a�a �����$.�[�hu�Q�}h��M�+�6�:���7X����$uO��:AY�GħgF�t�OW1��#���T�g�H�C�����\���}K�OԻ.Ta����%��A��)�������\�����Ȗͥ�嶚Woԧb)p�nx�>��Y�z�jz���tb�������%~Y4����A@�[�I���ob(w���0w*.j3�����b�Q�o��nc��w�9�}Xy*V�Ϗ'�<L1�9/k��<���/�w1��|c^��.QnKFQj���)����)�m&��O�bމK�?��Q�����!#%�#�/z	+_�,'��%k���,����r]�F8:���cU�+�x�� �T}r��<(�fk�F�s�8�`<]����A�)��3�AȆsV-h>O����ז:���a����`��t�Q.0��U.��,�C\���C ����*�ycw1�)p��޹��z�#���͑*Ig~ؔ]N_FU����Թ�������d�}
\���$���F��+��X��w7y�a^qAx����������}�0t�m� t�p� ���=Ŗc�2��>��j������F��m;Y�2�ݢ?���>���G���J������___�q,��z0T��u�;�Gt,�L �e>��~�!�����T����r���żl���*���1!ā�fK��'�r��D�Aö�c��������-��!�߁*K�����c��3�1M�����a���&*.-���Q+��^b�\MC�Pը�V���*���J�a�`�<0Y2�b��Kǧ��t����s�N��_�=�z���)�W@��ŉ�6SJn¼�;a��N��-���<N�w�r4��=��X�[3�?���c�c/d*<$�8�����(��QG<��p 9��:c,�軭R���nt�ҵ=�JF~EpgD�ߥ�.��aTb����w��=�yQ��]��u�����)�㫔/`�"��W9{c$�$��E��wC�]�i\!/�O!��q��`��$�Aeɗ���	����~W�6�)�~c#6`0���bTB��V����`��~�"c�[�.9��f3��wƕyU�V��`Pڔo�V(�����`~��W�v�m	w�+�Pj@)�Z�2���!����TjK'�w7�v	�Ns� ��e2�pM����D�86�E,s�=ۮ�џ� �3�L����`��Y�E�+V،��1�D�~�����=���G"7�Y����@Q+�h?�mU�3^)�4�0�jr����+c�@_���)r�3.�h[����D���6�iN�^�@=�|e�5�P81���28�{h���Xҵ�`���@ޭ��u�h$������ �����K�+}����^��9�|�yD9��x�u�*S�e��.9Ι���de���N�	}���&��j&5'�147ʎ��G�ۜ�UN�737�%`y6��E��A�In�ǛP�� g������]�u{A����ƨ|���+D:
����	��fS㈠�u�(:��G�uF��OFG;��f�ig)L���%�Z�Z\�3�}Z�O�P�T0Ƈ���F��ْ)(:���S\&����M�����t. �I#�c�)ߌ�nǅ��e2z����tf�e=�=�����F���8~o��"�1�����$U�k��A�0S/��,��5��3����j	K�L�[k��3X���$�F[5�W�81��jqOZϡ��|7���.�k����2����V�"	��?H1�����ZR*J�č�iI5V�Q5�s�%
���5�4�����c`�����Pkj|Bl�f��(.a0�MOpfx� G�
kC��+h���3|��"EV�N�R,xK	❽�
ͭSi�;?Ҝ���͠Ei��
�1����;�.��ڠ�6C���7�$�,�)�/6�,["M��$&��$�q��q�.#�r_���I,em��w[�#��8�p^��c�'��,D><)��w�J/�ӣE� W߆4��k�ѣ�11��+��\˻�ۓ=�d�X��%����3�q��w�C�u��V:?r�L��
��:�cJ�4���<�r�6�	5�~�����$&��:��≸L���AS���C��uȇ����gP���#B�
a�G@"��Q����9B<�&��K�?�+��O�"a/�h��~3O���v�;Mp(<��>��(E�ؠ� O��� Ht9����t;��8��3L�4ҘL,�(�V�3�H�)nm&�+�O-j9��%�H��j���c�Y���t�s��+��p�޾�3'��j��g�Sć	�����-�H��ig�A{[��@�}�,����c[��$W��mN��VW�"�$���rSq*����(Q�f�����V��G;Y;8h����<5����QT�����(�VQ�/[B���}fnL���IaՂ�{B9︡ǪL
�)����}1��Bd��OH��N�uW�$�؊!y
���o�f��i�sd���؆�Wٻ\PV/��F���^1�Z���d�"�	��������+�-�1�c�v3>��*��$_��i��ؾn�IA�ِ-�y�U�۹8�Zio�����]��m|�Km�&�s�)`%=O�ɪ�2�	NYDrJ��S{/c����)�+���N{m�Mn)n T`����Go�dQ!�`��fN�@�#-m���^��/G>��}�Z�	g�>�sx�̘��k�aa�l5f�F�
��Y�������F۵��y�8ٹ8�����ԅ�g�n�~��­��5�"&��v��%2������)n�%�S�:d�ղ����]ȚE�i�U���W@W�@��"�b�����ChȀ4��!Z�{E���j"�A�!�ɕZ1Z��Lg��fj��o�he�"�"�ߢ��/�4nR�Ӛt�|0.ȝ"Q�o���t��A��qC ��'I�
p\�|�a1!��U����!�ֽ��7[yEI� �G���`����#�d$4W��Ѵ�����bT�&��0"��J�9#������u��4˔��lT�>�>F0�9U�nd�t�!��<���kq�y����º,��n�zήN����X!>��ey�����;����oeOZ�H&�f��)�4�hɜ�1\�rJ?䱟���=v~w�U�;�>Y�D�c@����	�������O1�6i1���f>Up# �hP`�?oЏ���w9/v�/�c$����E���reR
�������Xҽ��*�d���0���1Ne�<*5��76�P6c�?3����� �W�i�5���iL6zm�V�?r�D�v��t��Y�F�2�ڔ�'LI�P�uY[ޏ����T��dyܢ�vud^<���#�!j���/������H� �`q��â��q �ui�����J�x2�]E�5���}ͧ��;� #%乒����Z��Z�D;b@!���t���m�~��%ѧ���(n�SZLu���{�l��£��>B����Χ=׬�;��T�d8Z�t��B�BO��P܄Yj�FW�%�X��/o�@5�k���:S�H��3�[��r\���R��0 ��k?u�[hXp�	H�c[bX
��M�(�l���5m�Rv�|�hޒ���K�����Y����'�*���5pox�y�~0����g6'ca��#��s��ӧ=t��p+�ϑaX푠�lE�Y,ɪy����Р����v������t�.�k��rR:0�	�rĭ��v��[q�f���	�o��П@�q|�*�#X�H��/����d��$�����Hc�ʦ�b����K�*�����bD��o,2�n L[wi���z *�q�[�<)TA۶��͊�`A�w��|`���e���RQG��Ձ����)�!�d|h�L���&�?�}Q�_�s�7#Bi���e�+�I�,$�����!�𵹪��w8W�F� �+U�@��pV}��<em�H@{F+��8��]W� ʞf�)�|���s��^3[�~�׳��֔��jM�`�W`��Ö�Þg���!C�%��<�K��w:��v�c1�ۦp�%����z�<����U{~59�]K4�F�㥧�j����e����g�
,�u��
�Fvy�+B�X��=w�$n�~�A5n-���̇�媧+�mqm]ź�������S��2(�֑��%�a��ۃ��m��2)K�?�ְ>y�AGܵG�G�F�YL_�6��0S�k/T��u�i�G��L�����[ػ�O!rA��jT�������v�
Ź�ݮ-(iƊ�!�Z�f���0��r��������`s���Vw�҆Z���q��K�������@��
�|M������S� -H<Hy-����!k�����bUAC�ȔՅ\Y�CJ}���ͯ����0V$�b5&���I�t٬dnp�k�I��:���
?���?�@�4��ЋJ�C�+a��?N('-����pwޱ{��dΚZ�[P����2�c8� d'5?-QQ���s(�t�G�ڸpX����c�E��S�1��t��=؋~�cSp+S땜N���aQ�*ʸ�W���P=cG�ΐp��H���;ǘ���ʀ��/�x�ܞ��{�ڰ$+]�Er_����Z��i�m<��@�\Y����$��Q�T�|�I�ӕ�u�~�X!�f�T�[�6�@n�߂�B>��AA/�]�~0	DcC���;5��pRؔ�vy�U�z\1P�HU���&�˥=���؊��葾jd�V�Wv�2�g�������jȾ�w1�[v�XIЗJ ��2<>���boD��!���ӌZ/(��w6}�0�0MEќ��!�Yz{h�G��ĳ�1Y�C��z��
L���G_�YaUڞ�^+�V��*�3��4Ǳ��#P���z�~��@|�s���3�$.�e�x�D��(xNW�P@Z9�e��vҭ1Ά.�φ�{���n��2t��� |�jv��h!��g~�]��yڪK�{����#��&�v�9��x�������K(͎��܎�e�>N{?ݯǋ���{j�S��N���Ζ���F��'N�1N3t�`V�j�3;���wI+�y��>� dqu�C��'!�uXlr�ITȨ�T���D�:g����&�����P�u��{:Q�G��F�IO��Q�ﶎ�gf��<γע\	$V}#O ��T-�~�3i�d�)���\C���7��MT�q����&u�`")��nD���-�zS�������t���2�4z��#�<��O�����Z�I���U�)�)���/�()I�y5n����O��j��^KVG�8qT�W�گ����pn���8.�mj�R��ś|��
�Ĉ�+僴���f�S�6	'M�Hn�O�r���P�+)��S��� A�;r��<�V��<�X��%e ����FHY\��dD;H�������߼L1����yV;��H�a�m��x�t�]9v��xꪃo�y�Nڞ�"���=���k�P�pQ=G��^Z�����6S	�}�n1s��mPo�.�QAiGO����"NE�^o��H��kx#�;�Xm�V�0;�)���y�	�M:��*J�Y�������eVP�I;^�xh��^�ղ����Qٶ_�	�(������򴙍�}gM�]��.Ȃ�+�B^���ҋ
\J���m}��WB�YHO-�N=/�W"=b�O>�
d%o���RM��jdd��ǅ]c�W'F�\h���:��1P�)�8yldp'	�b������%�W��8���6f� q6��!��.���4c�31ҧ��C�����<8��J��R�B����Y���F���%�R:��Zo Ž�'ܡ���SϧS�v>[U`�\��Wh;|�l� g�B?��hWe	��[�V���*��Ql�3�5)֣v2�&h�u1��X��i/Y�p��㶶�>�5,o���e��X����������#�'�՛�߯�s@�����=�ܬ��s���a�ߠ]N�$������
߮�����2�v���X&8�hh.-�m�.��:lA�.�:��s�v;h�[��`���@��s��[�q�W���H�ޝ���ɑ�^��y���f�� bA ���w*��KO�ɝI�,b���o���n\��w%\7��=+*�k���>�<�7������MF��[wJFO|�l0ɇ&���Qo�P���k�E)߷� �0������i�?!�Qb�W��L#�#��(xm+x��,`oO�~�h�]{�q���Y8=b�\<�+?%�9~�}�k;<���Fg�V8i�`]��k�Z��)�Ғ���s�Q|�2ʺ�j�o8����&�~`�\Z��p������Zi�Ci}��� �M�3�4�g�1k�0p7涹`�izZ���k�#��~�~�]�1F����Y���ݾ��=
�
U&�1��FZ�F2�+~��X���w�ی�:��Aq�֓���}��fD
����m���),�x��ŏ��2����U���ۿS�m�B�2e�~?gm$>��'G���ȃ�����_�bq@�c��@VT�{�u�S�G�CBL9������K�!.���s�T�e���s��2����c�鴫�*!]�f/%��5�r��-�Z����b�U��'��</h�:���x7���.��e8�F{=Mr
�"-�՞��\Hm��A-��s�݌����qbC a��A���ᷧ�7z�	7�y��0���b�^� ^+t�H]�/|�'K���V$W�/4��{@(�h�khRJ�ҧ����a�6zN�<�-ԭ���Pw�j������e�[G����c��Ldc~�����\�(J�G�a�p�ƣ��$cES�����]t
�=��~�f�p�Օ�ׅG�a��[�t��=��
��7`� ��@S����<f/�t �Z6�{�$�"E������Bi��g��y��ٜ�Y@$i�vɐ�M��˕"+�~��ߢ��T64vÛ�Bze���:7̙�&~�a1c�U�ǲۯ���P
�yN���6R�P�'����b��������~�F��$<�j �2ɓ�2H��1��l[�j&bw�mv���� ��C2���GD�M:�����z
��b9�Єln��Xb�ف8Y6������1����V�৤�;�G�nY�j��9�+��Ǫf�03w�4@���__��_���ڈ�@8�0�"�U3�6����4-�D+�f��N��T@te�S��i�1
�!���*{��*A�n�ߤW�ަ X�[2h]0��#�w��tf�5.�KQ�����W�Q�Rϲ�9lnxYU���&G�\4�W�	�N��\�e�HN7l7�P-����T�
��P��`�V�V�0NCZw3��Z`��r���>Ig�%�i ������c�Pu�B����Uw����:#�3��"?�H��euW B:I�~G̷F��BO_ci�+,��(�g��lKxƳV\�>L}St�O�u�Ti�]����I��)�CD���\����%�	
�ͭ�;-��)x�n�k���zz�0���&���!�p�X��3�>�W�Z�ݽ����J<U;���w�ɵG��F�K5���L�G�:jbpK�/y���ʢ��c͞�?N�p<�8j'^jʋN�b|���F��D���M��]��u^	�M�H��ґ.�R�|��f��iB�MV�h�5�Z�~�W$E[��`�ւ��c9��ˉ(k��l�vZ���0�0k�O)��x�.�@]Ik\|���d���({|$VE��x$�#���
�,�i�]���糒��EK 
N"k8)4��_��X�E|�7b$���v���,4�RM��?'�$&l:qFN�zԆ��7�m(1,>������<l�:e�����ܘ���+!>��>���JxS�Ӽ�
�9]p��{�kAJ��ʸ>�����5�ցԠ��}22X;�p%�R�a&��������ೡ-35�r���C=:�µv��qrx��~�����[s+��.ڡ���z�������dK�ׅ�$�W/\�l�9%��Ԡ\1����5t�drE	����N4�^�3�tl��W�1���vuǇ��F��@��v_O��f�46�����+�u���T�kkG��5-]�/�R�M�~&�@Z���=耪�d	��[r��S=f�� �s� �ෑ��.s��@��@;D�r�B��M��dY#[�������6���-Ԥ��7]��Pe��JMZ�S�̤:[qA�^˚�=��'&���g�ߙqާ�k��]�R�s��Bt<�&䷵le8Ie�W����c�!O<sL=*��Cj���x�wyM��P���r��t��Mq�^�9q���ڏ��m��M>��ѓ��S�'��C�2��g�\?f�����-�4�2UC��'�z�,�0=y�l��e�LX��:��4�X��5��LXǥK6(��%�OB�g&FJ����~R/��T���⫎G�Ss<� &ܿ`���3��۝```\�d-D#��/`ߵh���av�蹹u�M%z�3���z�B���#4���,�ze'χp:z��\7� �h%B�� ��T���omF��A꽿�:������y����� �Oi�p�*e��#lA�M�.>'mj���vZW���i�<�\3s;Nş�{CC.٬D�[P�N��|nitd]'[�P��N�GU2C_u��J~���meTX��s^DDvP�Cju��@�A���fb:��	��/E����|���x&̀����&w�$*"["C���[%����IL���2gIg�������h���݃+�n����u�oY^B�]�p�ѡ_W߰;��w"8+�w�G�O$G^^%WC-.4p1���4�����Y�Ƽ���0���*f �����C$�Ɩ	済��ݢ�!JZ��	<�z��k��JjʨW>�V`�_����T�o
:�wO��$���D�l��_�_3�d��0�Ju��Z9 z��	�lb���L�py���{o�!5'���9�A~��Z]�}�df�1Y6��ډ�My��^�2��� �#� �=2�(�w�?eƫ�$���X>�.Yf� ��eE���R<��<z�!�[���3�W��`ݾD5���H��Dzu��'e��0s+�O������
ǌ���(r!��X�eG��D
b�?[�)��yg�f�<�Ee�\.I�ǏQ`ǡ����3r�s��� �Y{Z[b|�#�.5���_@�$_�%�q	w)��`{C�� ��j��ހ�q�U�a:�����Ù����
�y�:x��U���Un�/��'n�&��R/�2����PF�Gpm��A���P/<G��]8�/V�\49�a���Þ	+iM�n�<aЋ�9��c���C�s�� ��i|D	�N���+ݬZW���^_�R�S��[�{�16�	��Ǥ��xD��y0��Ķ�hd�5M�s�Y]]��.��-f�����`R�F�d�|oJTW%+��ؽ�����E��]a��J���y�J� g�(�C\��{�KDm���Ž�r������� ��(���q؆G2ɾ@��I M�6�������x_�qW�1�H[C�`�LeK��L�����hu�N���</ϴPX�t=��o�K��Ђ�b�8�{\�c%9E�f@I�Xf�}4Ru���I�w�'�X� �r%,'��iq���d��ls�%��n#��WTQp��ϠAc.��6�3-�^��8��\5�Q8��¸��=���Y� ��$�f�o}P&)f�$��F��\���c/��	�*v��vꑴ/��f?��K/��xtā�i'0��:a��z��8 ��H��z/^�E���CK�53�����Ri�B��<k������鹿RT�_D�_^6��g=(_�̌L��	�5,u.�ˀ�Lt�'��fjgR��l����K%��(��A�.��[It�L��>�8��~-Ζ%�/S5RA�VĆ�G*x���Qd`��F[c�";���9�Ѳ?�s�(/6���X��)m_q%,�qI�S�M6��(u#:M�v�"����T�c�4W�Fi��e��kK��J����\$P�U������ඔ�%Y3C����9?�b�.�۶4�X��!� `�}���jxeYܞ���}\�n�M8%6b��+����[�/F{	L������������#6v@�@��H�Z�g����1�BV�*J~Q�՚�Ԕ[o�]	�����$Yǵ�ڪ"LX́66��A#J�a�]�k�"C?�/N�.���7�b����)P)Oj�K�&��u�Ddq0e��F7��Q<����9��yF��;:Ғ�D`��ѽ��j�Z�+@$��k��sD�JV���X%bۤ��f��˞9�i�pG���[��ثB�-Mn��O@���up\9&=F���sȚ�.�����Ct}�Y$��u����R��3bg����Њ��
����;��q�� ���R����R��d�L�\�Sn�ͫ���>�g�%p_0JI�y˘:^��iKQ��>�{����)�kg,��y��0�$YAK�2ʇ��S��rT)G�m���n��Vb73�"`ըXd vS��eت��a�(d��-��On,�T`��Bn���Q3�"�عV��Q6-?,�'Ȥ����'8�ccՈ�,���8���Z�j�uk*����5�C]:1�PY�C2������٢�%IA���b�}J���nAn�gE�T���c~&!C�Ghm2�E��e o���[nA�S!�����֟�*��BihT���X@i���Z��,��у��g�����.��Zh��ٟ�"L���G�,��Z·�gi�+f�woĝ��4��"쐟�s�4@��Ӭ|;|�8�����oa��t���<U= ;�]I��
�V�|ܝ0!o�<������D���7�8qI��ÎY�5���0#0#�
$F�h�#�����+�4�m8��0t ��܋/#�~L����u�04]8��>jt>
0BfwU��\�Q#�!�a��/�Pk�q�������"���F�@��ו)�X3�Q��V�響7���;��E��E��Z�.y�xN�)�CGh[����.r\��0��e)vP<UŚ>�#�����¡��7|��@�-4g��#��=�>�t�#�fBP2_Uo�w�k|09�fH���6ӏ�S`P�5?�e$L�-�!Ws�W��*��o�v���h���ՄeWK*G�7���6�A�?צ[������) WT�;���2�Lq�!m}]?D�(DϏ>�����"��Iڦ;�L�'�x��a��`�����n�MH0^N�8�u�j���RY�"�J5���ָ�|��G� �m�������xD�_E/!~���y��cQ qM�%�X˒t���l�ZFHm;��͔��1���?q�����(�åZ����l[�l`�hԯ����hՉ?��ݧ�� ���928�BƭBa�n���yY���F�s%��A2�PoVi�=���*NSe���up�[k�	\��F�H��:D }��?��>h���	چ�[4٣��\�z�l6_b5?l�vQh0鏍@l����Y�D��y����5B�G���7g������C���¹xW'��>����sŮ �]=��9�@Ra��`�\j��+܉������`Gʮ�Yٍ�hzv��׮)[���._��.:��A�DzSĿ�vюZ[Ƥ�ʬ�����q���PH� I6=/�^���t����?�_�]�\sbW�����*@����_,qbV�o~�7n���w;���K*E4����<�}X��ބqv���Lw`�|r���%(=��Qk�&+b��)5D,6�z�^�N�x�?w�^Qx�c����#��S�~�?+�p,6���=só<���� ���8�,ٲ��+'�v�dG}a�<�l�2�F=�c8��	]�4�p�{)��o�0�Ds%����
ʐ^�j��&)�<�/`�.)�@}z�U�¤p��C�5m��O�5�I)䈯�1�p�{~�v$z0߮�X<��y$v~� ]]�FD����n���j�w�����8
�lʓG(���F��X+�>jX�?xw�
��Љ�A� G�ȰV�&%��(���m/�D�����I���}2�~���2e������m�ZC2;�?��O>�G���YQG���\_.��V�2�҃�1��-�h���w��à*�^�D
��y����eeq*�`7�F6Cی?�i��o���W�UuI0��"L��9m�
�?R۬D��@���9���R[�t�L)+��U���o����`��D���&(VuX^}_�Gj��3������Ŧ(��@�G������ a�ơc֨���x��E�}��	M͇i�d�Y �Z�%�H��:�:_�Z�lP;Bdf͢c^��4#�M�O�g9ŧ��B(N|�Z,}W��?ln����:������O�c�=�4��8:�E����B/W��0�IYJ�xF�Q%�Y���]o��K�ƾv�S�t����;[y�\�2x������ ���?U��h8�	(l�[Bh����ͭ�Ml�;x5M�Uv�xh�
S�������
Y����>&��[�5PO��Y����H�Z������T��G_�'C���t�s��n�=T����{�a8!�����9���Y��2����C�⠆����v���������.���R�:���R�%č6�v_�[Q�f����O�:�nq\�9���HC��iԬ(��dV޸Q+������Z�be���ww�*����~��m�ub$�(o�n �UwI��Z,�*�.B�;f�<	TSۖ�3���@�gwnԉ|@��ɫ��W�Q'o�����F�)�uDDL��,�8��#?��Q��4�Sp�#"�9�̙�+��,,��ޢA��ӱ�Y��`s87��� �q+5yհ��|}��<Eq�(��F"58��]7���~�o)�z�����ssm���f�^O1דa!�th��J�`���΋b��b��~��C�aP��2����Wj�V�1��,p��2��+bz�����ڑ��$~I�]+@F�kŧ�B{���E��a�
��X�U�B��̣FV�H+"i]Xó�w� ]�^9�A�B��{��S����M�rm=���͉���:��3�t2xؑtM]�A"��cǉm�*�2	�?���>Y�BG�Ek�'Z��9�_|:�d�{�K�gT��/ui]4G���L�T��֜؛��!R�4�x(�T��!�{�O�V7ř�ή���N
!��f�Gk�c�r��\�~���@���y�K��*��`���gz�����%W��Og��IM�EƔ\��S� )x��-� ��[�����b5��C�,��e<��#&[���������T06��bn:�č�t�lXN�ۼK-ݥn֯z�ϴ�f��gr@�05��p�Jc���Ba���N��-xl��!w��҉��T�z��[0��ڡ&�c!�d��9���� (n��G�6p�/���ci�v蘟A��;t��(=��~���p��|�ok/a1�ʘ-{��=�=Cg<����h�rV��J�����`3/}�]�~��{���$ՠER����i:��i��s�led�<9ǲ���$���4��)h���AT~Ԡ��F�;�6���ÿ��B���!�N�=r5~1c#����i���t�R�   �  �  �  )  p*  �5  @A  �L  6X  �c  �m  �t  �~  `�  ��  �  P�  ��  զ  N�  ��  '�  |�  ��  1�  x�  ��  �  L�  ��  e�  '�  �   K � (  �( 0 �6 /= pC �D  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr�	p>!��L�>P^�x�#\`yq�~�tD{���O(dG6â�ߘ<����F�N�B6��~�'.>I��]�(��d_�R>`��	&D��3$l��� ��'y��T"`/"�	�|az�H?X̴Y��ǘ^�B| �e �x�@�?	hlHG �*&���ɵ@�<A&��H�'�T)r��u����`��/T�i�'�S�č��F�P�+ 8x20��ĺ�y��Y8#N�P��1�P	�BL��'�)�s�Y�1~"AۇlX<�XAL<��8h�B��.z��s��N�@�}�'fvM$��E�d^� jSG�>l%��ρY7H03�,D�������b�]S�lZ�r�̹�'i��1�	��~=Xc@ѯMb����ėL��Մ��?�Ox��W���`�~�p�B��>eBV��H�Yw�^�]�*�x� �nN}��/!D�����^����b��WL����O�B���J�l�٧�QM�H�R�ϘB)&��$:��«z��u;!L��;-�Eaș!��5z�y���6G!���.Q��G{*��\�Ǭʓ��-W��S�ə�"O^���.ONA+F��6[� j���%|O0`� �B�v�ڍq�ڂ�x��i�ўʧ`.Z��y��V�k����=y����&j$�y���^9la��&^r�8Ql����)�O�yA�B��6-�Kd�+�j���yrj�8tE�Q���T�*�2����y� G�g�j)"q� �O>&ݚg��,�yb�D�#ˌa�E��^02}RgN���'|z#=%?�j�a�/>o��rw���b��}�S� D�DjF��$o�`t
�H��,�n��1�>��p<�R�� ��x�h�&RI�$��`�<)Ǡ]�S���C�g]wh(x�ԟ4*	�)�d�p篆%%Æa��*`��H��Es��:u��n+���ᑧ y���A�^89�`�<�0��%kwL1��9MV���&̟f��CƸǬ5�ȓ��q:��Ϭc����U�� ���԰�&]/+�d<sF��4�.��ȓ׀)��[�A���Ȕ!d�(U���Ҡ؄�P��3�ǶnO�B�I�'F!�6�@��$ZB*�!Q��B��7s���$�p��� !+ց?��B�IWL����C��sT� q� Եa�B�	�23���BK�8Uzuq1�S���C�)� j��Q/�9�1u�M�I��Xq4"O�����	_��K�	��7���"O��L kމ����-u��Z`�'A�p�<iڒA�Z��N@W���H�n�<�`kÌf(����B�"�j`�"��<Q왻Z���z�䛫b(h9`�@�v�<��4W�̅RQiQ2Ć�k��Ui�<yW!R#b�H%B�̟�`�.��M�<!@�s��@�B���$����L�<A�}��D���^F?�5�p�RK�<�3��-6�&�i&+��
��XGjAD�<��F�a�<:�B!|��aE��i�<��c]!ؼ,��&�06�ݱ��i�<10m���(C�I��8�	w/{�<�3n�'�$={a��;�\��3�	B�<a���zsҥ��F]5g��(i���v�<����~9zBd��W�.��!�o�<�擰a���N?W�t�e��f�<!4)��%9g��7iC���W�Z^�<Q7�'+�𛅏�6?:P��V�<Qt�t�T<Jb��Xd,�3"�k�<��a�?pY��Ht
�*T���Kt�Q�<Yv�H6�\xa P**�Hh#�n@T�<1�
ס�ΡS���)
ֆ�I�!�z�<AE���)4�1χ(U���p$_z�<iա@6��$�9V$0�q"�r�<Qt�]%L�4�2RF�]�jq�M�m�<�Se��\gX0���r�T$�6��p�<ɓ蝟Wp��2T�a��F�<ٖgE��(
@\��2G\�<ī�}ߖ�I�E�l�`�[PK�}�<�%��{�\t� ��>D��� w�<�c!H�Kھ|&�Up�!B�q%�C��CWx� �i���-���
�B�Lu�u�4�R�i��#Q.p�zB䉾^5k�)�T�p1�3L��>^B�	�U��a���=n(��3��i&B䉺k�����Īsx`y%o�'x��B䉦*I�ӁRZt��rD�<U5�B�I�Y�ș��#|�(
�� l�hB�	'���+ρ!AVy�N9}rhB�I5���۳Vm*�b�E~�B�I����U'Ѐh�^��-�B��_�Di:rcʸs�6DY�+T�O�C�ɩNQ$|2g��E��P�a�im�B�ɭQq����S�)���sE�9SzB�*�ع#́����;��â�NB�	&��
nLo��LXg�I2^B�	;����#�����e�KO�B�;i����55�R�Sd���xB�I�E+`�A��Z��h�'��C�I�q�Ґ����/~�Da#֬��0�rC�I-�H�(�ѾSJ�ҤJɂ$XrC�I	���w@�4�>0�BL�\�TC�ɚ@�B�� �� 1�I�K�)� B��T�@-�4OW?;7�ơCI�C䉄Bq�Abe"P�'&�	���	=fC�	3/&)9��]� (���Q�G�B�I;p�i�OӤ-�&��c��q�
C�I�4(��];y`�M`�/�8�B�I�o���3 �X�-"��G��C䉷s.`�B�S٦	9TΎ�8\B�Ie�θbu��:P0��'F7u�ZB䉃>Tb�"�ɏ%�P�āc6B�)� |��V'�4�H�P��-]�(U��"O^�3���h2j5�F��o�6hp"OL,�2��9<ct�AބM��A	�"O${)�+3�y��*��U�D8�"OJy���C�H�쨰1�
U��-��'���'�B�'��'���'���'���%u&q+G���'��Y0��'���'oB�'���'c"�'�"�'�z9Yq��*g�Hr�F�A�^�ʕ�'(��'WB�'�B�'h��'�2�'b��yQ�H.&�*`�`�I=�\��'���'!��'���'��'���'�>9Q�� ���g���l���'z��'��'���'���'�B�'t�H�r�P�7 ˔�G�VC
�a�',�'}�'�r�'B�'��'F��s���L
p���M�,\���'/��'�2�'���'��'���'Z��ql
�lr��D�":��I1��'���'-B�'�R�'a��'�b�'���a˖�c��X{����TJ:X���'I��'!��'���'b��'@"�'G�@u���\H93B�p?����'X��'8��'H��'�R�'5R�'V�H5�-r�,�C�$Xd0���'l��'��'x��'D��'RR�'b<$� '�<3�)�� H8mxv�'m��'��'��'���'B��'c���Č��Z�b䡈5'�iCu�'�2�'e"�'�b�'p�hӮ���O�x`E@�a��B@���EЀ��Gy��'w�)�3?�B�i�!�B#�g�̥�T���$����?��<��mA����4�B��m�����?5"���M[�O瓩�jH?�0��[��<`����B�^%�2"/�I̟ �'��>�"6��Q�
%�QI��/�T-Cr�Z<�MC�a̓��O
�6=���#J=Lkܽ@t��=�J|�@��Od�d�Pէ�O�1 w�i{��ܒبg��
`.U�p���[�h������=ͧ�?I��)X%8dyKT �Q�"i�<�-OR�O��m�N� b���W9�A��>e�x���'Q��T}�I�@�I�<��O�9#"�%%�|SG��j��Щ�����	�i�,�C�:�6i�R�Z��(BU�D(����/�l������ry"^� �)��<� ���u�"L�MZd"%ώ�<�S�i�ށ��O��n^�S�;eպ|H�bk��vR`%:� n�����|�ɾ���lm~2=��,�S�U�H9'!��jX�ђ6ƷVjڠk"�'�<TS�' �i>y�ڟ���֟��I�f8l|�Gꐝd���vL�$[|*5�'3�6��U�~���O��$�|����?)�ɐ��h�.)�T�ZG��#��IӟH��x�i>}�	��,��aó$.���4eЁ25�c�P>?4�hoZ^~�`�B�����?�����<�/O\1�R�@�c�  
R�̴yIrd�ҋ�O,�D�Oj�d�O ���<���i������'O���O%�Pȫ������ti��'Zr�|��'���ҟ���џ� ���`P��d�M���g�zF�lZ�<���_�p:`?��'����w�����E
&O�-�bM�:7����'\�'�b�'�2�'g�>���%Ƒ&��|*U�ߦ}k`�B�e�Ol�D�O~ow���͟��ܴ��)�$����d��Yk�f��f}+I>i���?�'{(�1�޴����2$Y�Fß7���h�2Tk�Sq���-o:����䓯���Oh���O���A�r�>�Y�S2� ���ӄr��9� ��"A\�mK�f%�3g���'���O:���c�t�eӎG�|��%���yB�'�:��?��O{���,Z�N�!�F��^����-e<H���ýjw���I�?�� �':(�I�[Ij扂�<�Y�K��7�&�[B&7W� t��͟�����d�i>u�I꟤�'O�6-����yHcG�^� ���}�(}*RI�<���?�,Ot��<��.:aK�l�>}kҠ{1��:�����?Y��#�M��'hNY}�Ԩ���Մ
5k�*�N��"�M	c���<Y���?���?���?�*��HRwm̆B�� [��Ú@��U��򦭉b�ڟp�I�%?�	�M�;:0��KNn�� ���	�4]#��?�I>�|r���MC�'<*���e.�(0��;AQ9�'\6 ��������|�Y��ȟ�YV�PT���IF���D}�U��؟���ߟx�	Cy�~Ӽez�M�O��O� b���C�i0Lu 9h�(�I���OZ����Gy��m�E�T*�FL"��&?ѰK�)Y7�AD�׊��\5���
�?�@��W��d�S"�$2μ�1�$���?���?���?!����O�]���Αf;�\�q��6)���r��Ov|lڭJU1��ԟ���4���y׉¡ ��"C�_�;���Q��_��y�'d��'׼i��i�iݱP���?5Z��o���À�0Il�������'M�I�(�	ӟ���ӟ��ɷ`<0�kZ�HK���%�wJ`�'�7� �8H����O���t�	�O:��>	8��0D�B4[ΚDZ�陸m�<��'���4���$�OR@��B�nl�A��hH)"�XP�h����6��<iA� )�����?�eW�<�*O�ۗ,��e9�i�EMZ4y@w��O4�D�O>�D�O�x `#�<�V�i(�28�>�Z�V�(����UFUh�U��'�d7�1�d�Ob��'���'2 ���z���@a,V!�U�-/.��i���O�5Т����s������ 5��;B@�8�㤍�o�,�'5O.��O���OV�$�O��?yS�'���&"��F�*�t)
t��������\h�4iÊ��'�?9��i�'��]c1iL4���[4�S�M>j��3�|2�'��O:J!s¼i��i�5b��
 	�P��^'?� ��k��0:����d�'8�Iٟt�IꟌ�Ɂ}:0ٹ&�Αo��h�2"O--F�D�I۟\�'�6-�6����O,��|z��}�Bh���k�kCM�z~b)�>i���?�O>�O
.|W��?�@nFe&� ���#qQ�MrĲ��4��X���`��O�A�1���Lc���$m�x�i���O8���O
���O1�:�EH�fLӸ�b,���6�j!zv!R���'M�`w�D� ��O��$׆l4�؞�|��U	�UYr�d�O�����c��Ӻ�6Z��U	�<� o�r�a1�d�)+�
	R��</O����O���O���O~˧b44IWc�G���u��'m�b��iq��h��'�2�'(��mz�a{ �K$9,�K儇K��8�m֟��I|�)擊�6]l�<� .J~?"a�i+�^D����<���&���D4����4��&�%���S3��a!��Nv�D�O���O|˓G����J9~��'7��.wTH��`�z`�
���O2Y�'���'r�'-��Z��@:7�8y@���Y"���O�9��Z:?�pD�%�:�?�%��OM��Er
�)��?~mB�OF�d�O�d�OJ�}z�ZG���S����(�&�y���=�6�޵>���'u�6-'�iށ����>"�xb�I�k�2�B��{�P��ߟ��I�c�LnZ|~B��L�R|��w���%�3�T`Q��688y��|�^�����p�	��	��\{OJ�18������Z��-��xy��t������O��D�Oj�?��KEk�,A� �V��
���%ȟ���OJ������	/HcJ`���R̔���ȟ�3�ԲףG�����'7Έs��Ο�Ӗ�|�[�l�h���`�<��e�ҟx�����	$���By�d��ԣ���O����o�<Yy�����ۘ@y��Od��O���|�)O����O���1u�:lJ�k��1Ϥ���#��@��kr�@�	ǟ, ���c�TU�4��Vy��Or��?�la�P+��[ڬ9U%Ǵ�y��'�r�'i��'����ǚz����b��tÌ\1u���P�p��?�i!<):�OO"|��OR��*�gx<(@+�L>)���$�O��+�x��ش��8T�|���P�y�Zˀd/�%CG�@��?1��(�Ġ<1��ɮ;3����K�Ha�5�ML+�O(�lZ8������	v�D�U)D�p�1]2<�Cċ���EB}B�'�b�|ʟ葑��:����W#�Ce>H��TzHP2E遯y*���|�a)�O�I>��i�`q�\+Q�P�k��I�`/���?���?���?�|j,O�oڂ$�9Ŏ�E,���cX��8dޟ�����M#�rd�>Y��M��3ꖙ�\lI򄅐L1ֈ���?q���M��O �:g悯�2I?I��Eށu��Bh?KH��#�k��'���'�2�'O��'�哢O�a�œ�]Yz��O�<��4m��)O �$��8F�O��d��]	
�lM�5�Қk����VNR}����쟤%��S��L�	��~�lZ�<����7s/�z�dH�C�*����<9�A |I���z��~y��'��"v|Xe�j��~����kN)k8r�'��'���M�q�?�?a���?�v�H
}ˎ�Іm��z	�ѣQoU���'����?�����z#$,XU�E��bx���4[�'�}���@�t�����~B�'�00�� �z�,FE�m�e Z�<���R:|! =��R(�< Cp�A�?���i���U�'
��n�z��]�D�f,��+H�62��UMב3�\����Iݟ���d�ɦ��'t~U�5��a��lݎJIjl��∞%��T�	�?QcK�<)O��������O����O��!`��9���G@�,�&pHv�<��i��՘�S���u���'�R�B�Hxt�U�_}�(���0y�I����P�i>��	 �Gh�7}��l*PA�+n��(@Т�U���o�[~� ��"iV���䓶�d$4����ʂ8d�*q��C�Ah$���O���O��4�,˓@����4���¨��ـ�@F�HoR�1r�xӞ⟘B�O��$�<��H�R�V IEG������V�3B�	Qܴ���[	P:�8:�'@���n�+��̲�L^�HN�I����2���+�OX�	���,I�2)�FȾ�(`(�Oz�D�O�Imڿ +�+\�Ɯ|"��.)p�I�A�U8����(J�'X����� }c�V��L��O�=oR�<���;9d��YPz�G�oV��4�D�<1��?����?9�-	��4!��_�>5����?�����D^֦A��Lğh��ğ��O���QA
�4�ҁ�ӌP�C��U��O���'���'�ɧ�I �%�R=c����0j����=D� ��-�7Wv8[S���ӹo��|�	�P��x7N��G�9��'սC�^��Iϟ�������)�FyR/m�������p��L���ِ|�0
��Q޼�$�O4mZ�aC�Iݟ ���Y�d��A3��֎#�;�ȟ��I�I��)lZZ~�#�#w��=�SJ�� <�*�+T;0���ZR4M�%��7O@˓�?���?i���?����)�)����f_0fn{6d7ElH@lZ#���I͟X��Z�͟h�������5?���:3-
TNd�SĎ�?�����Ş&�}�ش�yR#L	e�Ό(G�\�]��A0�Y��y�L�r��)��Z�'���֟���b�&HQ�/\v�J`8��;L���П���?�@D�'�6M/U$���O��䍤G�FqZ�OV`�����i���D�<���(����H�?q��Ҥnk���I)�}Q"! �<���HшѩF�<|3.O<���'�?	���O����|NT�ǯ�S�"�Ba�៼������	��G�t�'��`D��1O��}QE��V�ѹ�'�(7�"�n����4���ɝ�w���S��3C��(�?O\���O���;N��7M0?i�LV((��)C'�y��7RVJUrF�H$<$LT�H>i.O�)�Ov���O��$�O� ����
?�USɋ�uZ~�2a�<!ּi~���'Zr�'��O[�N͡I�F���iY�I�"��c��/)*���?���ŞM�zJ�}��ՙ��P�T�w^�M[�OB	"T ���~��|R_��Q$M*;�0Q5�@�~;0e�t�����I՟��ҟ�dyr�t��c�!�O*kP/�S!�t����R�@���O�$mZY�QG��ݟ$�'��-�j �C���`懀��`P$�+Ư��������}N��Px���eာ>� � �G�CB�2�`����ǟ��Ißd�	���2�f�9oI�`jD�g��;�Α����O}m�,�����0Qܴ��`�Ũ��-;d���f#�|�t1JN>����?�'#.i�4���3P1̈�EH	[\���ٺ)W�kU��(�~�|�V�����,��ПH*a����l	���@�Լb���d��Zy��n�6@Ԉ�<1����ɑ>��)HV����AwE
,/��I���D�O��<��?Ś�JĘZg�͓����r�����i�D���w��%ʥ<ͧC>��Y�?˘A��E�9b(Y�f��%��D�	����I˟��i>A�Iןh�'L6�"\m�pK2/��v���S"�wC0�����O`��Ȧ�$�������O�5�s���F<��@�]���Ps��O���@4/�07u� �Ie�x$9�ܟtʓ7����Ď�5I-N[F��(0#��Γ��D�Od���O��$�O0�d�|�g�H�D�T)YW�+�t�rV��;_���%�B�'���d�'�7=��� H��m�@"�	�K&���Od�D$��	��nR7�e��!èΥ8�<�᠏"""d*�g�T�s�	�!t��Ey�'M�� 7M�
w#`�K�!$Q��'���'{剏�MC2Ȃ��?���?����o"(�Q��`m<E������'U���?������̙�$��hoM�RV��'<@��D����Ȅ�~��'�5��Y$e|�1jҨ|�L���'�6�z�cC�
>��œrN�!�b�'q�6Mv�j���O�TlZ_�Ӽ��È�L�Z�ɂ*F?:A���	�<Q���?q�6��Xܴ���яn�uQ�O_�hŋ�4C̊�Yo�x� ��E�cyr��(P�X�Ba"���S�
��jy����,	������	_�'6-�w�	� tJHؤ�����	9�S���Ɵd$�b>u�ėNK��g(�5�e��n�b�lZ���S�WCa0�' �'��IupR��֜~��� �^���I�x��̟"eߦ
��L�'w�6�@;C�����3Yؔ�B��@{�:���-A��DZ����Icy��'g�듖?1*OP�iۣV�h�Z��(��ғM�`��7|���ɝPL�9���O���'v��wz|�x�f���4�L�e���6Dz���I��(��埤��П��:t�N j�91D�ǘ�(����?��?q#�i����ȟ��o�X�	�@�8��¹(w�H�e�Q3T�'����ş�S�J`oZQ~/Гl6�mZD)�-R<\
��(���"�g?�J>)O����O����O~�#��� Ls�ib�B�(��)e�O��d�<���'Uf`���?������xdTp�Hʀ�8P�Y�<i�ɤ����O���&��?���f�`)SC� |*��f��X8X!���2?���|�M�Oj���n/R�Γ]@�Ȑ,�HW|(C��_�o|��@��?��?��S�$U���?�M�G���(=��QҪ1�f�@���Q���*O>�$ �d�Orʓ�?y�-��X�P�ߡR��#�a��?���%Dm#�4�y��'S	����9O�Z�N�{f�!��fM S�$�v>O�d�O����Ob���OV���O@ʧ
ծT�f|6Be�� E�-�M�Ҹi�HJ�!�3�b�'���O�'J�wb0���P�\��s&��2,���'X���i>M�	��%���� W\U{���5R�)���B�̓f�8���O�@`N>�+O���O��+@	
.(����a \�T����`�O0���OP�$�<��i��X8�Z����1%ؘ�9��=z��]���J.<�?Q�Y�h���T&�sDQlW�x�d`+uh>,��!?���ȲlD�8@ڴ��OȊP���?!Ъ��Z!�4�ϪsK�l�%�=�?���?����?���I�O��r���GNU�� r^�HWM�ON�nڵ\�I�| ݴ���yG���H��	�м�!^2�y��'�"�'�vIPE�i*��4/G���ܟ� 2eab�D�:`�* _�`Uj�:�$�<����?	��?!��?!"��7/[ }���X�KyJ��i�0��D��M�q�F��P��ԟ�'?U�IB�R�q�*�7kHQ8f2�!R�O|���O��O1�bt1���W�(�&�ϗg�qP�K� Ak.� �!�<�J�J
�ĕ�����19 aJ`GX	,\^U���N�h��?Y���?ͧ���Yæ=A����p��K�h�p����0r�����+Y���޴��'v���?����?��n��xݞ͋�T� o�Ueh �r�L��4��D��\4�������P�s�痎Y�bD\�.]�髒7O|���O����O�$�O.�?1)��\Q�5AU��l��i����ӟ���џ��4�@yͧ�?ad�iv�'k�ઁ�QB%T��$+H6f��i:2�|"�'��O���$�i���+�j�A��U\r��(S5c�%J��$���6���<�'�?���?�����	>�$J�-G�2IZ$�[ �?����ę�əńןD��˟8�OA �@i_�v�ToZC(��y�O���'H�'�ɧ��@�C 4A�LY7bu TH4��~���&�N�x�us�����*�BLM@�h��h�'�*���Q���=�� ��͟��	��0�)�wy�%q��5� "d��]��$����IĘ��z�*؛���u}b�'6�PI�#bNT�r�(Y%Z����b�'=�.�������������<��e�� m��(A�z����i��<�(O����O��d�O����OH�'�2]�!u<!3 Ϡ5��
��'��dA��?Y��䧁?1���yǕ�v�x��@�6-��"��z���'ɧ�OV�y���i��F�vF2�I^�E���Z���X��t�̟xqB�|b^���؟hS���8-���a�GQ_Z;'D���	۟��JcyRO`�x�!�C���Ofayd�1Ht��aD�r�"��O
˓�?�+O����O��O�uA�LA��<SA��z���2O��$�1(zP$W:2$˓�Ba��O|���9�XĨ�G!�n<���ι6��dP��?���?����h���_�U@<@���d��=qbm t�������
S��d�I��M+��w������R�Dl�xQ�x$�s�'	��'C�=˛v���ݮl ��SLRQ�B�]�Xz PJ	�>�蒕|BZ�`�I��<�I��|�Ip�"�9k�(� �-�5x���sy��i� ayR/�O����O�����dV`���"]�H鰁��
m��\�'i��'Vɧ�O�b<�g�6��ġErR�iH�L��C�J��c]�@�$�64�Bf�g�wyN�xà=B@.��e`����EY7h��'�b�'�O��� �M{�n^��?	�L�_�N����81�7N��?�c�i�Od��'�r�'����$��} ���yC��z��0ۈ�(�i��ɦ#�l|�tٟ�����"��M�TW�9���ω�|�D�O���O��d�O��d3���[��Jtj݉(��i��@ϸ|�8��I៰�ɕ�M��*_�|2�s_���|"+[er����S�dQ���@!��'�V�؉�A�æ��'��=P6��:V�T��FD�Vy���K	;����	�Q�'���şl���x�ə����2�K;|%��#,Դ�����'� 6mCw���O����|�,حm�� u�2�	��ZI~R&�>���?�N>�O�@x�d��}�@����+�.���
O<�|���G��i>����'�&�x�Ŧ�.@^��$���G�B�S`�Пp�I؟@���b>ݕ'�7�M\�PA�p��`z������M}!�F��O���V��9�?��_���	�=�p�y�'=��� /�!l�����؟T��		ئ9�uw"<���/�syb�A;u�Ii����2�L��l���y_�x�����	�������O���+<���'Y"M�<LP�KjӚ5ӑ��O���O������Ħ�ݏE�:�rdȲ+b�av	F(��	�$'�b>e��Ǐ��y�:Ī��`کE�R ��J݄qߜ�Γ!
&��䫥��&�|�'���':a�%WY� ��D�_~� �`��'B�'=b^�H	�4\S�Q���?�Rf��@*��Tc�J�m޻��b���>����?YM>�f
��F&赛��"�
�Qp�e~��?�(�ّ� �E��O�,��A��I�	�N�`�q���!�$m����'l�]��ɟ���0�	E�Ӷ4��П �����H7�`��Hl�%N��J�4PV�Xp��?���?	-O�9�����@	���Y��Ԭb��jW4O��d�O��$E4�6�b�p��O��R��}2���3@��r
��"�Q�� :�$�<���?����?Y���?i����(�L�b���.��"�!���$�1�E"؟$�	ן�$?!��F��r@�=|�)�Qo�d�T��Oh�D�O��O1�qq1���wҩR��a��hiW�˪��	�&�<9��V�$�L�d�����S9_�,���)U��LM�4"�#pTv�D�O`�d�O��4�d�c˛Fd�*�h�T�D�S̷3����W���y��h�㟤[�O|���O���H
NT(f��4Iv@�)ʂ>EΑئ�iӲ�(�	 b2ʧ��;&K�'.�t��Cō1��K����<����?)��?	��?!�����X���?���K�%ſBEb�'�Os�
(�F8�$��ަ�'���K�d���c�	J�^`Vy���@�I����i>5��A��=�'�D�
� ~�($j
�k���RK,V�e�aՋ�~�|�Z�D��۟X�	�ɷAk�N��b�8REZE�T֟���LyB�|��u���<A�����yR���O�Tr� ��8t�I���O|�$,��?Y�W�c�����9*�ʬKȥ~�H�q��������t��o?1O>��h�bB�AaTAT*z��$1Ш��?)���?���?�|�.On@oڿ*�L��������l�;
J��!�Dܟ�	(�Mc���>�OF}Y�����p'�"Ob�����?!�́��M��ODe�J��O{�q��g��n�f�J��c#.�x�'R�'��5H6��'���'��O���7L�e>jֈL�Z����N`�V��l�O�D�OT�'�?Y���?ͻ9	,�+�̺ p��r�..6��<����?IJ>ͧ�?i��9ɐ���4�y2N�0�;���+w"���ɖ�y"��C�ȴ�����4����A ,;acɏ���c&�ۍ[����O���O��5���C�Xu��'�b���̩�aM�S4p����¦U�O�h�'I��'6�'32�҄��v�`Px�.3e����O^���fޜW��7-�^�S89��D�O♚���)LR����dR�i�^]T�I�����OB���Ox��?��b��<��%|�(�"�n�|d��Y	s�i�I;�MV)���d����'���i�55�Kw��ɰ�If6�)��|�����4�	�	lEn��<y�>��+6a�Rp��CO9o��,��%WO`L37oJ�����4�
�D�O����OV�d�
x�^� ��c�H�x$m��[�˓\��#�i �������mH�h�t���p��oW�?�������	}�)擷MO�����W�8]*�ݽRv�S���b��{�r욷��O�YM>�/OH��sD�/מ�
�MM�R�z�)�O ��On�D�O�)�<�S�iJ��'����{�<� C�R  ך!T�'��6�3������O.���O�� �f�x
�KEN2��H׳x`��ݴ���"�M�qџ�����nC�更�TJ�.9i�5�� ���d�O�id��O�$�O���O1�(H�jS�E���*m��T���O4��O�o�6.p�����X�	`�?dL�˵��(��Ȓu�N�{��H$���	Пd�	�W�h�lZ�<�����Jjܼ;8���#��/vF�!a�K�a���������9OۢQ���E&�h^8����MsE���?����?)�b���̄ |�,�U���7�`(枟\[�OB�$�OH�O�ӧ0P`"��2��m�ȏv	nyZ �;\P�n���4�����'�'DLɓ�n�b��kp'HA����'��'r���O)�I �M��X�2��tp�O�D��@A�^(9�����?᧴i/�Oz�'��I�9��y�T	V�5��(ʿF���'$��A�i�I&i޴
֟��9��`�ELJ%w�F=���	΢a��M�kЌ�g�פk��� !���< Z�NO/c������ҁ�QO '5��q�s D���,�dP�,�O�`-��!ǀV�rGÌ
������3��@D���ܢ=ظp�f�R�����Ak��b��]:C�cr�)��Χ�H�W�٨)��Y��U�����i�!}-�D���14"�1a�ău=�q�$�D �������`�8a
Qu���š��%r-���Íi���&�.O�4�΄3�tt �&��sZ�)	C߄/��5o�ß�������S���<�ӌ�'(5p�K
���4Bڑ֛�Vc��|2U>�?qR�^6xܶ��!�I9Y#pH�S̈T��'=2�'{6,X&�>�)O��d��XCMT%�*�x"l���Za91�1�Ɂ	{t%����ϟ��I5Q*�$I��Z��x 0�D28q �h�4�?��.
k��Ly��'�ɧ5(�5^ �Հa�.&��b�ʞ���ď)x��O����OR�d�<�"� ���Ԓ6�3]
�q��W *5��Zv]���'���|��'�"`˛+��$��Z/�dͳ���Z�2)�y�'�b�'��I�U7h�ИO
V���!��hi�y��J�8�4$��4����O��Of���O��$���ز*�)�h�A�=ʠ�)�Ⱦ>���?)���Ą:�̌�O��*�#0.��v��Z�+S*X�]��7��O(�Oh���Ot�3EI1�I�	�DL����-3$�c��6V�6M�O��D�<qG�:!��͟`���?��ˊ	S򢌪��(Gex�j%D�3�ē�?q�X ��x�����d�������[�8%R��G��	�M�)O�B��N����I̟�I�?��Ok�s�����׻v��vL4V�v�'|�o
�B�|b��[�9��ȋ���<#V��e웶�ċy5D7m�O��D�O���_h}R\�ٗ.�m4�H����'?�ER^hX�4j䤨�2���OFm��Jw�4P#�����5�E��-��ǟ ��_����O6ʓ�?1�'�xҗ�Y��rebG8i��8X�}R���'�2�'�I�n���Je���t�\)$0L=�6-�O<)9�n�B}�S�|�	P�i��{r��\��%@��N �>��U8�䓫?����?�-O�a�Ε.PX�L:���̩�D��y����'!����%��������s�]��12C,� X��E�3�H�:ł,$���	����Icy���7#-���>���;ƢY:In8���i��6��<y��䓖?q��:d�'G��ʥ�k�j�@4�ڰr��٘�O����O���<���l���̟���Ϡg����&�L�f �� ȗ�M���䓿?��M[���{
�  �{%��=d|��LB!���i���'��	�{Y��L|r���1#��11͖,Q%��@e��'���'R��'���yZw\^%�A��� ���U�[Cђ`*�4��d��nZ���i�Ov�)�a~��҇_Z|����QT�y�I���M�(O����OR�%>�%?7-�	�bTʁ,��J9 �#�=w�6� J��7M�O
�d�O��)r�i>�h�B� |!<���Ŷ4�@X�Q�-�M��?�����S��'��_�O��ˀ�B�&���$MV�7-�O��d�OF J��q�i>��Io?)�$� +
�T��,��G��u+������\�I-������Ia?��hՇ-\�{�č��@Q�ɂƦ���5:*���'4���'�>��U��j5J��"���$"�$�5b�1OP�$�<i��P*6�Z��V$8�j$�M�Z�@DϏ)���Ot�$9��Ο �7�p���`�Ud�H$��1p��o�1��c���I}y2�'4��՟2�&dٵK?�d��&B�$6F��վi�R�'P�O�$�<)"�Lަ��Gb7휘q� <Snm��<���O�ʓ�?��l�����Ox�ڐ��G��D�cW
p�V�kۦ��?����䈵�'��tq��55���P�^,+���4�?1���DEsj5%>]���?ט�U��]�c�O�j�T��0!Jf(O�˓�?�����<��>8��χ�\�f�q�<Ǆ4�'?���(�B�'�2�'��X���4?�NY��V]w��BdF�8_�6��O�˓L�:ExJ|�^uV�1д���đ�@�4k��ƌڢ��'�'4�d\��:V��tM ,26���L�,�;�]�\kFN:�S�'�?^0
��%O*d��,��mږK�>�nϟ��I֟,��,߽���|R���?��#
�I���3�"I��P�.�P����'s2Y�0ʯ��ʧ�?��'T��5��Wk��X��Z�h~�� �4�?�������A�����|����5k5j�H0��a���'��:f�=?A��?�����D�'QQ�ڄE5S?p��@��\�R8��a�	���j�IryZw��� ��ה%�ͳ�"�JdI�4�?�+O����O���<����X*�ə ~Q�QbZx��x�"DPi�������ןL�'�[>��I�(���c��ޔ�@�7#������O����O��?QWKV��i���Rt�C*aD���Uo�T���w�L� ��IyB����Q�Nဉܽi�� 	#-Ʉ��8n�����	QyB�ؤAO��'�?A���5dC�c�&tI���:n�xr��<I��	�t��ӟ��f
l�,'�D��
�rw$k�X��'�+�<�mnyb<Y�6�Of��O��)�P}Zw��f�ԋ'��uzu"�&I��4�?q��Z���ϓ��ϸO����7'ӂ-HiEa�{�R�[۴��`R��iZB�'���OR����đ?P�]�4���Ղ���!�r�m��*�I�Ж'�� �Dص?����Řd�4��G�ӪR��l�ݟ8��ƟxGi����ĸ<����~"`ұ7�lx�B*I|��c�̓��M3�����سt��?E�I�`��h��1��B�K
r��1h���o���X��BI��d�<����D�Ok�C�Ә|��Ժ7�1��+O"O �I�6$(�I��|�	ȟ��	ܟЗ'�4�rf�� a�t#sE���0$F&��gNN듯��O���?9��?�pC�e�����|dhQᛀL�͓���O��D�Oh�r\��S0����ڂ2,!��4
t��r�i\�	ȟ�']R�'!Ҫ�0�y�%(	A�u�3iX�(%<��n�-s�7m�OT���O��D�<����f���ޟ�7��}ͦ|	g�OD�t!� !�Mk���$�O*���O�X����sӤu����\)X�Mǂ|]�\ˤ�iLB�'��	���믟���O������%^�T�85�jJ0�X���Y}��'R��'�l,�'�U����0(8��ň.�:tq ��5�֩nZeyB�p�7��O:���O����u}Zw�X���'<}�!1��:\$|��۴�?��)%Q�}�s��}Jq"�%[�D�uKƞ:d"'+¦A�v���M����?A��R\�t�'q,��� �X8"b��d&���Et��0��2ON���<I��T�'>�%3���^�Hࢋ?5��Hq@dӞ���O^�dʋ1���'^�̟|��,m˄iP�3�TY��N�2 "Xl�cyr�'D��yʟ��D�O��ж�H<arm�I���CYl�LlZɟ̨!���$�<������Ok�/;i��q���[�@Tk��ɧ~����{y��'��'��5���^^u ��P�d��<1�	�Jvvu�'��Iʟ��'�2�'(�[�@4P|��`�o��I�
�dr:���'	�I���Iş �'@<�A��s>=�`,38��S�+'�HdR�sӜ��?!/O��$�OJ���2��Y4m�Y��*L/(�tͺ�A-@\Jn�`��㟴�	Iy�^�MR`�'�?����m��ĸt�vD#�bK�9Ϟ�mZ�Ԕ'Z��'�rJH��y�U>7������EY`g��[r�;i]���'O\�,��%�8��)�O��d�6ԪC,�H���Dh�f��i�� �P}��'Rb�'s2qٝ'��s����;�=@�"�#oo����a�J�2�l`y2�����6��O��O&�I�S}Zw�X����Hn��Pd�5w^�޴�?��0�����?/Oz�>� ��D��
� |�0�S�T�u b�izpR�}�@�$�O��D�����'���.:�(�!�ˆ0�VA��͞^��(b޴*b�͓�?�+O�?���ü�6�Z�kБ��W3}��H�ݴ�?����?i0+5��Imy��'y����/����Ӝ<��,S�"6z��f�'�"�'�*����	�O�d�O��� �]�vab�c�&G ݈y��k�馽�I�^���O���?�.O����N�Z�� #lDt8�LK$U?���RW�
��c����՟�������ky�.B��Y�<=*�(��f�`qp�>)O���<���?1��'�N��$�̛`O��`΋93&��Z�K�<.O���O�d�<1��ܩ1����
Â`�Q)�|r08`�@G Z���Q�d��Oy��'?��'�$�'�}�aNQ>P����W`�O���SQ�s�����OX���O��.�<�k�[?��I9E��z%aC4o�,���-q)9��4�?.Oj���O��$�R��$�|n�����xg�*~�FГ�EܷYnD7��O��d�<�������l���?=㳈U�*�ԑG"�
<Q��L	����O����Ov��A8O���<1�O}�̉�(�:"x`)p��3$�]k�4��$35�m���������S ����X!֌�!??pt{Q��g�:�ط�i���'b��'�r\���}B�ؗv�Rt@En�#�0�qA�ަia*�:�M���?�����Q�,�'����S�4��H��˯^�|� -x���
W4O����<�����'Z:M�g�,	5 ΤZ�r��'I��'�#��'v<�����O��	��yqG�[M#$�V�L]@6��O��$�O�p	�:O��ݟ���ٟ|�W%ʛ=ň���az-J2����Ms�����a\�@�'N�U�D�i���e�
"d^鰧�h�6���>Q����<����?����?	����Ċ6 �>�%K�,x�p��;Q�Z���^�Iן0��]�	ן4�I)y�@��%k��5���)A���Y�p	��$������Iڟ��'�z ˱Jt>e�$N�9�M��m�M�6KD��>a���?M>i��?� ���~f�%���'h��D-��K�������O��$�O��\z��0���4��2��])֬��KXP�ԭ��:�6m�O��Ov�D�O�]C�;O��'F�mB��̚B�-p�N�%M��#�4�?�������,%>M�	�?-B�#2ĨX�R,"��x�bK�ē�?��x �������4��!=�D]#&倥D��e�/��M;,O����Y��)A����d��n��'ĔKPb�5z�%�֏�p��!��4�?��q�Z(�����OP�����
0%F�ӥm}pqP�43���a�i�b�'b�O�*b���Qǐ�{�5s7���.�������M���W�<�J>َ�D�'�����N'�p�눣0�:��b�q�����Op��XS<=&���I��<��4���t�^ }_>
d\��-�ڦ�'�41��~��?A��?����K�0�ׁ�}!�6TP�6�'���4�#���O6�D"��ƪ b���{�tY����wLӨ���m\�<Q��?1O~��kO�on$D�Rć�e�@0xf�ɪG�\P8іx��'�b�|��'�B��T�F�X3 �<w���1c��[��Qڥ�' �I͟D����'KDm�e�~>q#&�G�}T���H�4*VT8	�c�>����?9J>���?Y����<��C�$>�V�!�훹+�f�����I3��ȟ���H�'��:�:�Ϭ	��y벦�5y����*7?��`l��'�l�����D�ß�O<��qEM�a6��gŀFq�l�B�i��'��IfG�@�J|r����1$��J�iBh8��R>��>�+Ob��6�i݁跨��v	��b���opr ��e���O�9���O(���O�蟔��á��L�N��.ϻ#DxAr�L�9��Iy2$�-�O�O����VB}�vH���jZҼ)�4�&DP��iw��'nb�O�����Z�q�Dh��i�S�$�{g��4�@�lZȟdE{��|��'���OԪ;ߞe�G���`C�!qӶ�D�O"��3C)�����O:�əw2��G懫i>,�fۚg�`Ҏ��d��ߟ��	����Ҝ������ک|6v�(Ea
��M���8~bX�-OP��OR�|"gG����BV�ϔt����k�*s\�O�`B���l�	ß��	ny��-[%`����Xt �;�jC�����m6���O����O����5K����X3�C�#�>�{p�!Yxc��������I˟@���f����0�|��pm�-ALQ��� �4��m��@���\$�D��qy� �'�M�@�'ҠLsG�0YV�
�&�X}�'���'h�	�ȕN|ڃ!ԃ����+�mS@�a��3����'��'g��'9�ˊ}�,1%^�C�%O?k�H�	�LA��M����?�/O�M����D�۟��5e �j��//`�
�+ي��݀J<���?�%N[C�'4��X�'H���0���Sd4�S���hO��T���Ŭ�0�MK�T?A�I�?�(�O2��,L�;:̨PD��q�8'�i�"�'s�����"�S'ㄵ�M�)�6� c끉/�p6m��	�V�m����	������?]Jl9�&$ Q0�+Z���ٴ5���Gx���O��1�,]�Ę2���^ː=i'������؟��	�S$P�L<9���?!�'��J�g�C\�M�7f�,z44��}�`���'�b�'1�+=� H=�H�.�p�+uMJQ T�i�r�\���c���	}�i��Kg�ħ(/�P��.6�(���>i�	�b��?���?/O�8�5��u�&�`�S�`��a�e�C
!3ް�>�����?��T.�]B�iL�M�$��a��vA�����\yܓ7�$���/v�k��	�5ڰT��i�p�4,�+Zh!��m��1c�2_�<�%$VqO����R(� L��@�P�i2d��`�I-
ǆI ģFF��C�^�+<Cp|PB������ 4{���G@	:*]��s�4m8G�&w����H-T��=8���4vF@Q[���1D�ڄ��j����'�X	v�0���-C�d���O��B,��2r-P� ����kP����zDV,��������O��C�x����%[P�����tS>�y)ǎy�X����;�����e7}r��R��q�	��7mZ�'N����A+G����s��"E�>�<�a� ��O��hem3}�BA��?���h���d̦0���Bq��2�$K��\
S~!�d�~�b�21��"$��ʀ⋸Mfax�)ғ�0�#��'c.���گ/�|y Q�D��ȟ S���(Ko����џ@�	����65�����W��!�
�U� �b�Ŗ~殍a�
�t!��v�g� s쨴L�HA��Y#LS�:�j�3%�zl�����q� �2�3�d@"/ yK�ȏ��p��M�.1�b�D6?!֩����`�'���҇T�MA��Y&!��m
����'���ز�Κ�hb��axp)��O��Gzʟ��ں}hVNءM���"2�!9(��+Kj�~Z���?���?aV��4�$�O��;E�y���Ӷ^����#Ԛn�E�W�S�>�7	�� Ta{��=���S�t���$�AY��p���N�ID�=lO�����Ŧ%*�1��t
t�c�+�+r�'�ў��?�&��,��I � �
�v�K$�^�<)q�Z�� �jÏo؜�w��C�}��	OyrČ�,� ��?��m�b�p!ԯ��B������?)�Nk����?Y�O2��G��9m�h#����q�0������O���� ?��x���*G�hqѳg�n{>�	�TҪ�e�,;���y�gI�l�j�񄀔�r�'��A����4��%c�+m��5hc���I0}>���_!���h3�S�BNC����M�6II/)�ty&��$���'fQ�<9*O��3�i���u������O���I�'D<�8�.�(E��[�Ék����'�B�ӧOV6�5���|�'P�Mx��S�2rl
�d�g��qO�Ы� D ��F8>���t�6pN���t�Z���A���.�)ŗ>�4��֟�I,�M�����O �X���:;!Fa;�$Q�6��'���֟ ����+�dE:a�R�S��ѱL<�1� �%c�x�i��7��O��mZʟ�{r- �-z�ԈV�O�4i����<�M���?��)�b�s�D �?A���?����DI�!!����B�Әc�Nh����8͘'���
ϓeJ�bff�F(��d�� F�4�=	��[x���ԅm��ݨ�O��ܩ@����L����)�3�	1VS���7��������H�!��TU�4'�Tʎ乇)̗E�����HO��(���{���pէ�+È��Ĉ�A��e�r���,}����O0�d�O�����?�����H�3d9�qȑ<��9J�g��9��EksD.��}BAߘM��hɓ���<Eɠ��`զ�JgO
��}Bo
U�|�	��u�P��V<)��Q���?y���?�*O&�$2��N�x���Ϸ�
��었�C�I4J4��Q�ޱ}��<Rf+�JFzb����O������CS��I
(�vՑ��<�T�Q�JY�8QZ��Iٟ��UCUٟ�	�|7���j[-`���0�$�A�l��X�t��� A���x2I!V&��LƗ����0F��Ç'B;	��rѮˬCrT���ߞ�2�'��I,$#2��''Ƚ�L9�@`
�I�c� ��	*Q �(٢�<r١�+�\�vC�ɕ�M�1i�0����B�^�:$ Z�M��<9*O��"�/�v}��'n��.:k���	>m���0��%7l�@`�β!�>���ɟ��`¯7*��*���&^�8$��S��\>��g�%Z�R�`�mN.J��	�<�'�r��oߐHu�]�B�|ۑ>��gH�;&b����NM0o��`�%1}e��?���h�X���=�pu�Q헓^v~���fN���C�I�eyV�ۣJC>JMp��.fSaxBM ғ2>��c/_-_���HCHv�n�!òiv�'_�E�(�:y(p�'���'�R�e�Q��ʖ����@�݉NdP����GE�m�H��	%	J��C>��2⎨~b�\`��8<O��K�F�6Y������G�M�ua=�����|�Њ	�^��7垏g)��Чe[��y
� << ��D�jK���,l��� 7��ؙ���ӮG�n�I��:V��{�dE�a����m5���	꟤��̟�A_w�R�'���:(�L��*I+!�)�0���0O&�sħD6
4HЦ�y|tа�ȧo!���6
]�1C�#B.�h@���
 n 3��'�B�|��'�����:=H^����V�V�IQ��I�Y!�d�
[%�1��.j��H+��"]1O@��'e��
��b�O�D�,��=3 �E���)I
ɄE���D�Oj�2��O��db>}JC�0T�F�H�.G�~⪍�F�h��r�&rjXด�د�p<!׬�A��P�A2U���҆8�
%R�ǹ\�3T�i �x�(��?����D��ҝ�Ć��1�JA�kݴXd1OF���R�KtN�8`Ӑ;�2Cv�T�*G!�d����I�C�0�0P�wjH%َ}�W�b��E{��)@�u8�x���\=�9�tk�")�!��0h�F̓���b�H�sDJ��zx!�d@�WĒ�qˈ�H�h�����5ht!��3z (�+�J&RuԴ��$�(_y!�ĐY�y��3V�:�E�Oj!򄈨;��0 ��g2�r�b�4*�!򤝀7�8� �d��q`K^�!��ņ	�.8��`Ӕ*t�Р4`X�3�!�Ě�-�ӗ��nj�0���T]!�dS18��m��_�s�@i����-	G!�dϩ7L���+��R�㗆A�B!��*u��t�k��zW�:!�D�*MC���� �b/��r����!��K�Y�rq7�o�,EbA��;y�!�]�}�dX˒l�0)��,8����!򄄁p�\ي�W�O��<b�$�!�dA�AV$i�I,EU��)_	_�!�[Ze�i�E�m�8{�V��!�
� ��aK�'Ez9�FiϔO�!��ٽ&�^e�b܉}T
�Q�+D�!��/���80���@�)�F�.q�!�"T��8J�IM�I)65˱@̷�!�۹]��i���Q�P|���d�U!�ܩu���f��<Q�(XP�I.x!�]�2}���̋�C�6�"��Y!�!L� �7�C(i�4�3.�Y!�dZ�lr���E?l�p�d�Z	E!�D̘z�;�޽oTp�i& T��!�䓣GN ��䊟5|�@B�R�!��1�|a)��Q-(�v�h�(:BO!�/�tų�aY�g���SH�9k!��N�8K ��[N�"p&� �!���3����NN�ut���増�=!�D�W!��J�ƣd҈+�L�-s�!���:U��5 �H�98g�X��(L
!!�� *=:��H�n��p��U|w!�$�P�̸��	+�y)T CbU!�dO$�*�[hZ-�,A��1'�!�Ăk�x�)�o�<֌�VPc�!��NPցXE�رE�z�mߐ�!�$�{����/ldp�o�F�!� �~���͖*Q\�0�!/�)�!�ʜu7���ŠM�\���.�	(�!�d
��9��G�2p �gٲ\!��,x�ʤ� nO�N������ȥ6Z!��.Vڒ`�Bgߵ#���a��A!�ӲnĦ�����$�h��5�!��P��h�ٍW��ړ�Y�F�!�M� �@B� ޓ��9An!�$*]�99��Y�q�VŅf!��=&<-B��&��̣�c��^P!�� H�! d�� w�hk��^Ej(��"O��Q-̾�$���-*�E��"O�y)��R:ʢ��#j��;"O�E�f�K�7]v(����C�� JT"O`a���أR	� ��U�<��ܨa"Ov����Н�h�*FHē�R��e"O�h��H�}5�л&�݁S����U"OZ!QU ə�d���K�/[�|��s"Oh�ab 30�x��w�ޤM�%�F"O�%HҩFt*��Й��Q"OΝ[W�W�L��(6j�'X.�C�"O��ɤ
��D�� z�	���`Ad"O�MA"+�A]��b�B�C�K�"OT�##-&#М����{���&�'��i{�収m���Y�j� ��]y��W�B��4^������]E��)��	�C�`��&C��>���^�&G�px���T�>a3�
N'V����V*������:��g"r��:s�܌@���4�Q��/Ĺ�ff��S���Y��Pp��g$�e�e
�7��B��λ_�z��ȓR���g�����ZB͝T7���O|�5��?�~dW�G�`,$��E�6TF'͡MZ����6���	t2��-��3\ԡ��C�$"��X
ci׀.88�M�z�dI f��E~���i4j��%+�1�b�:� �r�t���
]��Z3+�gi0���5+�FI�>@��8p��!XX��Y��v�աk����v8����o�Dr��(a�^�af8�)�>ѓMG/�*,sC�YL9���q0B.U�L��/��P
r��$,U6O��E��0H|���DH�,8���M���䞮&Wܐ��V<W�(  6.H���	�Q�l����B��@����$���~��;:�a���$���c��5y���D�^!1O���@�0��L�!/
_���Z�����'�ܭa��6#.����J�o����b�A�?G$�(�\�K�υ�a^�'�}��N�x��Kd���x����ϗMn����B��fX؋�����O�pC�_\���ϫ �6���D<s<d�PCc�?	�a�9̄�1�K-u�Fa2���K�'����ƈ�{rH�aŊM�/`�c��n쌙�����K�j�a��]�f����(�$MY`�R� n��">i�$@�@d��!̼��~�<ݘD� �%���C`�|��Z%gL*Z�� �@璮#��(�f� LLĻ3�d� �Ź7k�K�.�86a��2�1O( ��ML��Pa��>ga u��-�)bք�*3��8	��0:�B�
�-ڄP��+��b-� ��f*xt��ئE5?�(Ҋ�0=�0n�6m��v��_���e�n?c ��3|4��ROU�mKvh�D�V�'Tآ�7*�����:y����'�@ʖ�;�P�.p��e�(��D�{@�DxܓO�Z 8m�Fx�;F�@��T̼a���H�#W� �B%��I��A�,z��J�' �=�"#h$�c�<�&+,(��$`��W�.T}  !�I9w-��*�dM?R 4I���Ģ>1S�J�F���!AP�tll�DI\7��h���1�Jq{�.�i�������(o��D��i�Y���8LOfY��EK�-���2�N�:���@�OLo7�ꅩ7�?J�fX��M[�m}��0�J��h``���=H�S�J�S!�DR�",����ʙ���㠊�+�$d(�J��਽	�Z;
�1O���JJ"xͲf2�<�TK�:5��� �Wx�b��';�\��KA1����$�B,�6 *� ��\��<�<)�(��v�=7A�(�,5�6g@�1�k"&TZbh�bǒ�F�x�F}2���b�RĢQ(��k�,�i��q!�A�K>���Aŋq��93@�;B�t���S��T��gA}��� ��Cȕ���T��a�a���ZƦ?R.B)
Sm�L��TҁӪadJ�ce�dI9X�B�Bpns�R��gE>q!�{󄜈%=th�A�?:�Z�s�̘�L�ȈZ�K��Yt^��C�T>#�1O^��G�DcG�� 1�H�`�ß� �����:�����'qbb�h�;f�1b.�1G�n�;p)իMZ��<9t!ŋ�Z�c"E Fa2q��\̓A���(6�ܰ28i�lb�(|G}�'�&��X�8h�d+"H(}@'�qH�Se�4`�j +DK�t�Ji���u��Lb��4T���	{���� �=9�F�K����z牍Z����7dU�d����3;#����yKFc���dX�O:��tg_,�.P�\ �dH�P�:�"~F���P��AOM>Ĵ`�S��8`�t�ORH���Y�H�RI���9O��;?�X{����L��"�^��L�'�1�2�'�&m���&s����%��:ƜS� ���'�ƝQ�(�F�Hl0�g�a��S�:Id���D�TK�[����J��8��L{����L���Y����
p��3� e*2�7���Q`,&���2#�A�b�Z�s�;P���`B
.s"��T?��$�E�D���Qi�">��%q�s�������*�R�O�D�x��Q?��?!���$�.��������k�In���ڠ)d����	O$�Z�UI�5V����м]�E0%�� ���ɬG��CD��k]v(Q�F�L�">��@�3<��u�ۮC�j�ju����r@X�8(�����!�hxE�B�<A���c���RV* K�r�YP� �<9Bf]%%� ��"W�E�
qA����h��HJ�L�\��08 ��!'d�i#W"O ��C<S�l��5�S �(��#
i0�11�F;C:2u�B<��g���6,�G�_�
��|��,�L�\͆ȓj�QŏfA�B�� �3q�EѦ-����$���{�,�_�"!"b��rU�l�E�3�hO`!Ip��Hƈ��b�L5j�v`´�JB�X�YҸ�*�ѷiF��j��B�<���+��1�M��oX���6��Ħ�g��fB�H���ZYFp�$��OQ>ט!E�z��Ǎ�e�mˤ�#�$B�	�)�,aP���0c�䩁��3.5ܐ�v�&�?1�C�:8��<�V˽~J�E(�I�R[H�P�[9��0��=�����7E� 	Vb�W�L��`��3v�B�҇�E��zA�DL��<a%T��=�S�ѭ/��. �I������ܓ�`�
g��n|sf��0�0M�*#��͖���؂2�2����~�<!�"H�&���,�QaFm�Nr�� �d�OI"�n�f����)��y'n�4-`��ːoV�/��aW����y�Lȴ��t�h��;�(1˂&ʓ���5�hP`�]�g���ҩ�C⟠���<�1�a�<cLx%KV�/LO�2f�f<$)��]8n9�D�?�u���4H|����冣�4��tKI5>)H��DY�jHu�\��#�X"\I1O��'�H����D`q���A�Z~��DX�s���:2��Sg50X�Q�daKO�<��E�T��4c���]7r�1�i�.��!I3$_F�na�q+8w�Vy�bM�PˉOf2���w�h(�v�X`p��I�%����
�'�be���W�^4�ą�=W�&0�6!W
�>�9��T#�H�q�b.�bd���7^c�Xa�7&��`� =�:\:�<lO ���C���Ѡ{ր��G�	�lzV�Կ%��I�}\��Ѱ��d؞p�'��uh� S��	�H��H9�ɴ�XpK���L�O���R#�	_�$$�4K>���'�跖�1$�L��'�
qF(�[d��p	��OQI��3?��ӛCR:�Y�/��6�[���P�<��,$C�0�ԡ�(�ܑ+V$Fh�aq��!�:��1(�&����!;=��4��H�az򃈭z�X�A�ST?!6$��Ԡ2�M��ԡ3��^�<!���>C���x�&ͣL�L	c@$�A̓�( �(�3b��~%���p&քYذ�bQm�D�<9��Wy�$���<��LH�73�@s��0}�#������/_2�1�D[�~q�%i#L�&7��B�ɡw�D8{�׵Ey��P��B�y�C��B�\X��'��`ѫU�w� i�ՀU�B���ӓP��i�&V��hK~�s���,.8+��ξ��C��-a�x4�aE�n�|�ʍ3mrb�|�ƕ)S�����7Cj��adHKx�Y�3�ʜ7��C�	XXJ�F�Y�ʡ�R�[�6"����L��T?����F��O����9"��Y�S�{��ء�"O`Ȼ���4�2E����/gP�����;�<`J�&KDX�P� �Jg$���	0e��X�d,D�<Z��x�D3 �Q,%�J�F�)D�X�ˑ*)0:Т�Хd�z�qU�$D���Cl�T�Vĩ�s_��(U>D�x��@Z�q~HJ��O6G8|+�:D�h �
�(Wƽcb���d����3D�8�6͎1W<�{`K1�xxE3D�X����	&�8�r0�
0r���Pa$D��؅PWƶ���ʏ7����#D��B&N��y�}�pM�r�~(� =D��9gKO�z%��/G7\��c�O D�H�s(9x���beGk�J��5#D�hS�G�2q��A�=N�J�cL!D�� ��sB�^���yDU� '��s�"O(�,A��h�4��@�d@2"O�3+)u`�Pᣃ��Ҵ:""Onq��L�;RY����Y�"հs"O �6-�6u�Pp���_��:4��"OIcэ�6_�B�"�mɑClB-@"O����u&���vW7Ee�E�"O�(�V��h�@a0�x}ztp$"Od��$Ř�G�f('�\�YX�a9r"O~��Q+K�&�z�Yģ�)/G��e"OZ�Q���U!����@�3V�kA"O<(˶�Xx!��ă��*�t�"O<�.�4k=�`	P�Q0g`2*Of=Jf)�Y�vug)3T�U��'��*@��$?�T�Wj�R���q�'_�H�eD�<��ř4J��I{U��'񐕛u)�?���{d���O��Y��'�M�*��F¬��sa��^*�*�'+ u&����y�DV4��5�
�'��1��)иKj�"���>����	�'{T(Ar�:><�F�K9�Y��'Jia��B�z���:�/��$��'�<�X��S�NA�0�(U����'��d���G�[��E�2#OH�m��'�z5����?5��j�ŰA�r�Q�'M�P�N̪v���f$:��p�',�T�6`��3��!�v�:�͸�'U���,G��Y#�� 6�����'QZ!���D�4<�(����-K����'@��v��"z� fR-9�~�Y�'�jqj�G;L0�����"O���
�'&=��M�wzb��P����R
�'R$�6_Eb63��Fˢl�	�'��Hb"O(nlhzU�Q+�lI	�'�pe�v�IU� <D��ya���'��쩐r^��b�^����c�'�*%5JT���N&r����� &�yb��w�-Xq��h�D�1���yN��W�1�O��bZ%���ybJߨ����& �r4HIK&L[��y���^������bły�%�˱�yŗ�C$�,i�/��% �ÈA/�yr@�c;��I��&�"${#���y���sN�۷�J0tD�r @��y2邇�,k��+|m*�
���y⯍+|
�Bi��"�i�ѢG��y�'Ȩ�t`�@�r{İ�m���yRn2ŀ�a��Z2j�z%��(�y" �b96E �닼c3P��tǌ��y���&8���6�73�Z`($E*�yr�6U&�y�n��(��=+FŇ���>��OL �xC2Q�3ժ7N��蓨.D��PoFP�Jf��/!�pY�(D� �wM�3ˈ�0mʘy�d]`*$D�l('_�\���F���R�骁�#D��H��U������Zw��ӵb?D��ȰgO'���&�L�+���Q`<D�x�U���ITDX���n͢1�u�9D�8A�)� g�p�@
Ji����6D���D-}�|�)�k�F��De�2D�#F�Ϩ
l�5S�AR�2 (�5D�<���**
Z)c[�W�ؽ�`�>D�(Z`I�j�v�Ȧ*�?���2�:D��(A�v݂PZ7꟪!������6D�� � ��<|��%.�2C��\�"O��)Q
�l5��p�ź����F"O������JB]hS���ԬѴ"O�I�#BJ�d���9vYX$"OH	H���%� �����$&z��"O�J�J�[|DL���Y���"O4e:�+���Qz���(l�ly�"OxY	tn�A�a�1�T;di9b�"OXi�e����A�F	f���V"O�mqf��,�p6��
0RLyq�"O�-cE�?rf9pk��c?�@�"O>�At�	�4 �Y	£�28�nm)#"O�J�.��L�q�O��dX�H5"O� ��ƭo�0m�C�C"Rt�L�"Od؂�5{�a�d¦9n$��v"O2Y�!##�\)@�B�kU���p"O�$�Ζ8t.�i��ӁtCN�qA"O�a(�)�!=f�]�5�Op��k�"OJ�b�ˈ���7�4c$l;!"O�at�B�F��	��/\�OHZ�J�N���������E����/'#&�i���yR&H�+"�BeCL� x�B"ˁ�y�b�!T��욤�����Q[�Py"kĎG$���s��%5�{�Nz�<Y"���-�r%8��Z�u�h�ꤤnx� Dxb�00R���DG��e�"5�yr&ĿK:3`ݢRT�iC�c��y��G'[�j�j���L�ym�&�y��'�NL� +��A�<��'�0�y��O�+�Vl�k�Ks�9ar�M!�y�@��|��o�x�N��P�ִ�y��A�KN��� \��W��y�ؙ2(<S�"	fZ^<*'�֏�M��'�3`o��oQ�����+��m1�'�i{3���%d�
E�
����'~N�0qL�0A�!��@�'ln��	�'q�eY��W�*��dPq��W�`	�'��8���S�LR\0�D-V�.8�'Ѧe��3GP"�f�S�6ʺ�[�'��`�qɄ�R�F] �ě)q�|��'7,4	�HҫA��q��⇿ P(p�'e�����'>��L�a��8$>�\x�'T�3&Ǜ%�hhI��!��d��'���Q��N��'.��m��'����gJk\�a�/�z�P	�'�idh\�x�ĭȆ��@հ�'z�Q"@�H� X���e�B ��'�z]�!]H�	2��!V�̀��'�@ 0��E�F���釠b ����x��I�(�����YZ,�u����y"E��y+ܔê�5K��|h�����y�,~�����Z]�x������'�ў�O�����Lf��a
��P�b�4�P�'��(�ZM�����Bhc�'H�ظrJ˴|�	"��˸c�,qj��:O
��գ�:���$g3,�4j�"O|e��nKiʚ=�;I��� U"O�Q�@�V;&dxxY������'l��`��H�6&��1�/W	i	�DzB�'_�ܨ5�A�b�;4B��T�{���2��e��i� ��"���L��`"O���c�& ��P m�Kv�
�"O�8���." �8�E�>]k^Lt"ODa�ȃDy8�q1�X,Q:-i"O� �����M&~�NLR�)�,O2}	#*O�x�W��j�αP�!Up\I)�'٢`j��4�+T�O!Q���		�'u`1�Ck�8F�.�8Fl�D*�Z��6�S����j�\���߫T�t�Rӌ�
�yb	D�j��!F��S��r��ɬ�y���#�l���M�x}�ħߠ�y�F�{&�d�Gi[KAB���D��y�3h���'oA�J�<�bް�yR��"^��xǖ�G�ly��˽�y�NQ�:�p�ch�%=��ݻA�̤�y�/&-��`�`N�@��xpm���yB��0���!O�1����*��y�+��r�P�!����%��h����y2� d��T[R���$��DC ��yR	�#+��h �-�� *�i%┷�yo�x鸠�ri^�L4�G�.�y�f\t��F�9|N����AZ��y���MCt��Ȍ{�Ne!��R��y҄�|D����J�i���5�U8�y�O�\X%�b�17@�a��yB���L�)�f��2���	�y�H�o������6�)��P��y⡂ryXi&���4�d$��Y��y��JC�D�IfգyF�($IL-�yB���r��3�[>�$ЖN��y������ۢh��F��Qp�Ț/�y�DD�JITp�������y%�Ǘ�y2%<L�J)���I2b�'�y��ԣg���R��-)7� �����0?�*O���g��@R�H /=Qot�"OZ�Y�ҹ�����ɱY�`(!w"O�a�e�Qݕ��P�{��83&�G�<Y�dξ���� �X� ���[�͐E�<���	0)v����A,S�ċP-�j�<��?��PW��lܬ���GL�<�1	ߴ$.P�DO0hb|��*X_�<�����ZvD�Q3���.� �U�<��+K�iߎ�x�e �w��!�ɖE�<Y��ڒk��m{�oޟU��d��u�<!
��V���!�J�z�h�#��Y�<Qa �9&b���λ_�d���V�<鑋E�n�x�q�K�%���0��	R�<����o*��5�ȅKn8ѱMR�<�'nƉJ␩��|�b�)��r�<9��D�Z�KcBżFތ)���t�<��M�v	4�b�B�D�rQieMMv�<��M�=����nB�vu���Ee�r�<AdC�~�h\H�"�4��8��En�< )�$:�E�ĨWZPxK��B^�<!�3�Z���%{Y��2G*A�<QtD[��DT�N�h>�S�X|�<���X��6�ܘ4� �3#��{�<�jF�1��p��P9#�
_�<!���T�9A"�7Bz$� V��A�<���Flᮨk2N�f]�P0f��h�<)��5\�j {�S�fm2Q��fCf�<��ݸ<2�9��.D(.(��X�L�c�<���P�pxE�٫g�B�В�`�<�⫝��@ź�Kר-t"�!%�^g�<9큮!��Ja�էB�\)�`�<�J%1�0)rM��U?z�Іs�<15�s�q��'�X�
c�<��:~���j�UIj��uU[�<� ��@�����2�(�W����"Odѱ�l�4u��A"'E�E�¸G"Ox��DF�3d�0�£]<	 �xC"Of�y�c�:,Y����$�	i�T�be"O��X��4���â�(�(�
"Oڬ��ˋy�nl1�/�S�F�p"Oje�a,��U����JB���#"O>�bF��G��+�B�+aƼ1�"O�Q1�&AnZM��V�]�A"O�$JքؽP���a�@��s�&h��"O�E��KS�L���eo�-�D0C�"Oj	࢟�T��ʦD�/x�2"OB��T��7U�]�$�<x}�"O�� �X�W�D���t��'"On��O�pO�t�UI��%�[�V"Of0 �XO�"�G�K�0�F*O��q�逑z��X ���4Y���'<�4�!�%h�Z4;�L�<WَL�'e�QA�녋b͘�`�Y+S��ē�'R`LP��è%�V���f�=q
�'(����hL�zuv��V����`��	�'8�8�oM8n��tk��T69��
�'���z�H�4H&4h���K+)����'���B�f� ���i� \ĸs�'�����˄!Ξ���Z�$��
�'E�Qdq!Dh�G"
fdQ
�'k&IJ��ܢ+��<�d;��]s�' :�P�E��v�����@oM�5r�'��sD�#/pds#�/c+�	+�'��Q�m� cH���bE�$-���'R�*F��GR�����0d��'v6��0莥-���@"��w����'m*��O�=-�xA�A�h����'!`p�v�U((��%Hg Q178����'*�X8�Ƅ?a�`��F�/6�`(�	�'F2�c�͛7�*1Z�	����	�'HL-0�Nٙ]�Le�o�i4m�	�'�L��֪�4~�nu"r♐��r	�'8,��c��4{<�����A[	�'^@,�B�F�"����@����x*�'�����ĢPb^�٠f��h��1�'O�#R�2@{��k𡏳�*�P�'��U�fN� ����j=u:����'vz����p�P]��M�?x��c�'�I�&A�=�8�I��5��(�'wX�dl��n̜ Ǧ�}´��'�d1��`
�̌�F*݄p~�i�
�'u�r���)jdc�o�|F�	�'`��陾Db6��5��ml����'iV�R��ܚljpň�âW��I�'�$�;Alݴw4�G� b�9P�'Uzq�M_4)j��vG4i+����' ��TO�0B&Y�����e����'m�u�u.��_,��h�pَM��'���r�+�G-:�O��9�p���'ppQ�k�[b�	�MZ�r�'UȔRh��d�$M��b��v$��'%��g[�j�rIP K
����'f�[�_�G6��"7Ϧ(&���'�Xq��T�`���v-�--.p�'U��DN����3/�O_�i;�'�~�ض�yZ��I�c�22@�t�'�4���;u�h��+�!0nf�'�x��LܝL� �H��$�"�K��� �qY!��!.6��]%J��""O��)rF��8@h����Ϣ��� �"OX �����Yd���	�/��ѓ"On	C�su��U�7}m�"OҤ,וl�F�!���W�L��e"O�A�iX��[��R�Xk�}�<�1���EG(\���̓<�TE���U{�<	�(��e�ƴk�G�8j�p�F�t�<�#隿q�h���u���Ze@Np�<n�%^y���C�N*���AF�
B�<�Q/^&	� �Y��$�\U�Zv�<i�T�g ��:���#IoZ}�"K�p�<��iQ�=Y0���>��Q��Gp�<�A��j>�����Q42�Fa
 B�T�<�"�J<��{/B�U8��ׇS�<Q��0X=�S0+�*�+��N�<��l2[$�n�-"�B�Ka��M�<�cGУE۔$�TL�d�tHs��
H�<�v	��<��Ţ���O�6�� �G}�<���57,D��G�`V�mj"��|�<դצsm���AO�og�,*�D�q�<���&Zm��X�Á�>���+�A�R�<�d�72��u(��_e�e�P��P�<a���~�hڇ�@� 0�]#�I�<9�mZ1j6Q`��_�H��ʅ��@�<��bͪh�⭸� :càQ�Q��S�<QK#,/�� �B�55��D��	O�<YQ�C�VT��!dgX�XS���K�<IFˆ�@ۚY�p-8[�� I�<�ǏڂZ���i��Y�U��P�c^P�<�C/�&4���
�Vy2Uz�s�<���VZl8��_0���S�<Y5e�
&)B�.�5{9��\N�<�B���T]*�S���u�TB���s�<�c�۱a�p��&EV�[H�����u�<�U�_����
n�(S��E���Wu�<)Ef�?��5������ ��q�<��LX�\�V	d��
Plxs��x�<�qj�.I�D�,�2W��u �Gu�<!�m	2�X�1sk۰�2�+�WG�<�N#�F913��Yw ��w��y�<�r��oު�ґk\ P,mzծu�<Y��h>����Y�r}"�bKo�<�O_tA8�K1�߿a&�tҕO�A�<�f�9k��JǊ�"Y��Y���U�<�Ќ�;b�[&�.��T���l�<�E�	��|H���U�&�a�#�T�<��K8M$�h1mȗn� ��u�<�6���'�L$�1
)v��u*�o�<)3n�W��:ňM�A��k��s�<YV�BК�j &A����R$�n�<a��2&�%k� ٧���P�L�g�<iCl�,-sb���^%YjY�ï�}�<a�)�Onu"Vk]�UP��2hu�<a��K�|T�� Sֈ-�7%�m�<�e��!�h��Tۗ*Ɍi{#o�`�<�JQ�*=��@R�ks��jS�B�<��BŲBT�:���A�X��J�}�<3�C�.1�� iD'��E�w�<E,�G�@�wLJ$SĘx*#GJ�<iԩ[�t0ѹ�׹o��mr��[�<q�,�p���g�2.\�n]�<!͞	;I�|@T7%}��a��<�GK��)��y+��C�����R�<� :��榆�;�jHÀB�&��lI�"O���m�uz��"�"(��H�"O�h)1��G@ ���A©A�6�B"O]bb�,{l�	[���¹	�"O^��7��qB*9)�/�%(+�I�"O�M��ʊ�d\9��Pp�d��"O��$-Εi������H^��C"O�Ԑ%NQ��@�CeRL�j�"OB�8�/�Cpz�K����2�{�"O�@���&�X�r`f[�|�x�P�"Oz�1bi�Oo��ðĊ���e:�"O����]�|�҂�?�2�2#"Oft�P���Z�Q��Z<�(�b�"O�,
�j�|*@y��J�qg8q"O ��$�?�\��hMOt	7"O.�hHm��:�i�{C��"Oji��%ӞF��t�ӛ13���"O@!���?[2p��@��Jx�"O4P�c X+��;�٘d�̐�"O���B-^b��̓V&1\L�"O��c�ł�2��� `jmZ�̂�"O�q(���hS��s�	�n2Ir&"O�0Z�%
�z�jϐ�6O���W"O�� f�5�P��ş�(<P%X�"OP�SS&�4b]bѫcW�5<�dI�"O��p� �d ]�B!��p+Vmj'"O���錵|�8rb`&��c�"O���3��73���`M�33S�)YS�'�ў"~�e-=OUn5���9g��=�!#���D'�S�O�<����f��%!ƍΙ!��r���'����łA�fP����>9��)
�'e&�F�:Q��Q�$���h�	�'i��ˁ&Q!Ox�%�F*��kR�,A
�'��<��OU�f!��k�@�1��I��'�H� �&x�V�֗��L>I����> Z���K0�4LC���,�!��S(��95�x���k#N݅K!��\��h�������mÑ��O"i �*NC���YƎY�x�̭�G"O2H�Q�:���[g#ü[���0 "O>���7
�樘4�ώ�0���"O�Aё@N�l�Z��v-�J(-J�"Op��NU� Zn��"�_�<�`��"O�͡à�mˌ-xc�S�L��ɠ�'0!�ĝ�H�*�ŕ�L4j�-� q�'�ў�>�scS)��q´��%�i���,D���סI(,��{7�֙K j	˔,D�L�S"�6uL@��@ur@��-D��%�>x�q��Њ�<���`7��c��@hs��
M#�����	M�R+2#6��]���¢U�<@�0��/8.�A�/D�@�2���V{��?53�	�C�Od�=E��4Ojq��� ����ـ�*#��lX�"O��(�d?ތh�JxizW"O�c�H����Uj
وv���R"O����%	���p4�Ս3�ZH��Y��F{��IF l�<L�g"��:K�ܻW���da!��8�N��j�
6�8�F�](>!�ݺK�JՋD���*<$������]�z���$��B�`���>{��a�ڝ�y⭍ 
)�Qɓ�\��t���yr(� 0�v����B�7�y���l�P�c���Vi��
bF���yr��� �eFU�\AqKH��x� |ɉ5�I�ba�zI�6>���"O����'@�!,���'�l( &"O�A:wn�2I�*��0��$������!LO���Nڍ2M��7�(Nh�y�"O����蝆iP"��8dŢ�"O4��)X8�ZV�X)I
��Q�'�I�w3�1rԠ�P���FǄ�p�B�	\,�}X���<$�}���҈U�y�ɇebb��J�l��@��߅=eh�O��=�y�L݊6�J��1�*�>��G��yB���"̎� Bϊ>"FL�����yr £@%���v�oi< ��y.@P�Ȑc[5e�X5�f���yRLW#\���AP �Y����k��x�'An�H���Ϫ�`��0�؅h!�דc@ +3jB�y���pr(,,�!�GEQ�l*�"�F���42�!�$ƳpC��I󡔃n qd�M0F�!��N�d�:xe+����+�h�G�!�Na�����X�P�ʃ ĀY�!�DL t���#��4X��z� ��$���;O�zU��EL��g�2���Y&"O��c̔�e�ڬ�&L=,B�4�$�<YO>�˟v�b-< ��+4h�J_��C6"O�$���
+1��D�7��Vb��"O�)rŊ��-�8���G�h ��"O`u���g�*-0�HU�xfI�"O� G��$ꤔH�GZ$eP�1"O����n+V��zT�:X&]���	J�0、�zVE��%�"n�⼘5�8D��0g�3L��%�G�d��e��!��������F#(xa"h���'�P-0�f��q�kЧ8Qo���'�X���a�#6Tp�fTB�t	��x��'7&��qB�ѓp2|��Z �yLK�%6�|[�
L<kXZ�@�h��yb�рa8�����0�h�S�yR�>z�.i"i��u�|��C���y�I��AJ:pRr��Q���y掅7�NU��gQj�8<�^.�yRş�^ώ��@AE�f�<��(��y�,n9�����,Q����!���xBI�(���S5�@9i��� �N�'&�!��"N���D;���� NG�!�$_�l|����LZ�+c�=`��@��u�`��7E9B��Bֹ͚��ȓU�\�W�sC���c�m����'nd�[�'�rQ��쒎g�����'�!a�O0�|�c�G/[�9��"�'.�e�r ��t%��,��D�s���'@��&�Asq!�f��
2�	���?��*��.uX���O���"O8:g�܀� ���+��1�h�"O�U�7O��JܮLZW�B���"O�᧧I��qv��8�r� "O��ʁ���T��WiȍQ͎� ��0LO��:��k��!s��>M�j$c'"O��qK�����C�D�<{x���"O�����ػ8�H��އ%pX$r"O<��A�1�
1�l��XQ���"O6�J3/Iej�8��Қ#?��u"O����mΛ�)���� ��"O���R�O�@�6<����
>	�a�"O,xyAk�2��v��)!��}� "O� xɳ׮�͖ш0o	�F8�"O����
O��f��V.��lX�҃"O��BQa��HHb�,{��x;�"O��{Ӆ��wz�[��f[�D�"O(k��"òHC`�=����"O �r��(K���Q4Ꚓ!�N�Ӵ"ORM{�eҌ ��8'�D�X $��"O��:A�^�X�\9�߄aj�80e"O�j���D��a�ӦH�H�ޱR�"O�\!c蛂Aj��y�F�"�	�t"O���C!"����F �)�\"O��/3f�r@��΄��č��"O���hV�k�H�RX�v��� �|b�|r�7o�,�J%�ђL�-��Ȟ�BC�	�<��)�F�V�A��Pj�C�yY���4 \\|p !�@�!�B�1bsR��A�KMD�����n�B䉲���qR��h�L�=1(P���d�������=b6���V��ъ!,0|Otʓ�y�OӦ/F�:q�E�I-�Ȣ��&�y���}P��2R�
�A�4�04����y���(��H�AU�<�>�TE0�yBa6]��}PL�7Uu�O���y�MÖioT�5/;Q��yiJ8�yҀ��]C�i����7���*,O��y�J ����ߜn�q0�jд��3�S�O,�lނ��� ��v���'�b�AT3+È�aգ�����'�)�A��'`��B~�BA�
�'�(�C����)��p`�	�
�'�%!���.G�1`�K�b"��`�'���C�O1w$$�����8Y�*y`�'DB�aV��	�l�gϖ�>��99�'�B�{�ʟ{�D�&��5BCX� O>����iý,��æ[*9���#��.e!򄂯ń#sA�#�%b��!`�'+ў�>�! iD,k7���eM��cQA�@%4D����K�\�f�I�@�s;�C�$D����`�'^2��j@��s���"D��H�C�t�`�
�E��|�0XB��O��=E���E�Z��l��j�V'�u���:�!���.N�(�3��>���"0`��W�!�D�&r�� �J	)����sM��P�!�S3Jgz鐀&x�(�/U�1x!�d��Fؼ�Q�ߡI�*�����/{t!�dN�Cl��BD�$9~t�!�i-m!��*(�,�#f��Ja��C�_3:Y!�Ӄ+
H�A�BԿ!�D� ���WS!�\�+Zp2�l,v�z+�n�2$�!��$(�B�RSLΝs�Q7䁀��'�ў�>�8&/�2+�Liਖ਼3^�$u3��4D��[p&ٞn#ny��-�5T$u�f(D��#� E2�J��t���)�Y�(<D��V�[�ie�l�,R�AE2QJ�=D�TWiEff��zE�]�C�0��<�	d��k�ƟO�6S�ɝ�xK�![��9D�0���ɯh�#M����Ҫd�!��20�pgc��*C��$	�!�!�¤=��8 '
8l�13W��J!��?D�%#�oX	!$�82�Ζ<�!��,����$��Ya썡'S!���/C�,�'��'`I�'�иM#!�D/p�3 ��"3�j��tm��
!�o2��r�j${�6�D��u!�� =������!��@[��B���"LO���՚n2�lD�ҶXs�4� "O@{�@yrܥQ,ɺWkt)�"O�!#���8(BA�U
n��#��'_�d��Zy&�Y�(�P��dB��FS�!�dK�=�BP�'�@;_����*9S�!�D�+lT�"df��$xbń�!�W�	�T	J%J<"4x��,�k&!�$@�3�6H֏�� 2��`,#Vk!�ʃp;H�Pr�`S Z&�ջ5!�dH�H`�2��?4AP k&��3!�D�>���hׂv-.e�l�3!��'x���p���#z�jVAҎg`!�$�;1�R�����X��!p��M�9]ў��S3�2$)���Y�r]{1�$m~�B䉬~T(P��5L��`�FwhB��6?�~���ǾQЈ4#p�"�R�=9�'�d��C��,w�8S`�]�v�`M�ȓR����F�]NX�bVoߋ=y@u��y���B	Ӯ)�lt�F/PS�tX�ȓ�e %'�<tb��2�֊��Ą�,4ƭ��E��N�'iT
?BNԇ�>�����`R���h!m�Nz���?�zĭ�w��L�MU�^H���j Ys"�c0bѡf(ӕ"�؆�IH���́f��@9 G� ȓM�
��T�J��
A�ʛ�T0���s����R+�mD�
o��ȓ|��զ�!�h�G��z�5��3�&,�DJ�B@��� ���iO�	2L�S�,���cX�S�̇ȓrb"�T'a��\b��0#�~t��6<�(Qc�)G�j�I�k�� ��1���Kм	�q)�#;|��|%}�4�$̲a��ND�@���wp�y(�֊s���H
0���ȓ02�x�I��y�g�J_l�ȓK�`��ƀu�0���%$݇ȓGT��*JДI3iP3�`@��t_J�7�
�d�:�ǎ�{�bA�ȓ2��s4M��i�8eK�/���ȓ$�,��nW9 �����#�0���G{"�']JH���(��A��/"�&�)
�'�Ą8Bm#*p$-C��ճq2nb
�'��{狏W!��zD,jQ:r�'�vb,� b��4�V�c	���'lX�ȓ���P��3X䈰�'��p��b��(�q�ٛS�R���'h> "�>$��|��j�EP���'���`TfD�O	�A);	��'$D@���'�� ���7E�,r�'�f�Zh��7�����N�+*Nȝ��'����@��:�Dѓ�HYWδ1��'پh�(B�L���S�FwV���'T���'1Cc�0Y�IԞ)��F{��O ̹H�H�%fK�J�K:�P��'3����2`�d�lR�[�@Ap�'����7!���d*۹W��(�	�'5t���G%E{�a�@Ã:����'XB�;�C��`P���N�2�T���'=X{�BL�::�R3h2uz��
�'"���%"C̀ �����V�P�P
�'6�q0�d�JU��kD�� �v@a	�'��9�I�#}�>Dz�O�F{p8���� ^�1@�Q/w
@��7:9�6\4"O���AH�%;v�R�Y lێ�a6"O~�0i�	J�����f�2T�$�{q"OB�
�*�- �vP�(1�� I�"OT� �JҵZ!P(�B!ۻa��ٰ�"O�5��D�)*������!*�y
T�|��),6"�p��� .�q .�K�B��%Gc(���L� J��u�A+�6oÊC䉍d��������J⣖�vw�C�'�H�a)	�.���Z���h���=��PF]�"!+{H��۷GD��j��ȓiŲ�����K��H;*f䕅ȓ*�~�f��7;�@[e�j�ֱ��:h;�I�M�`[q-�h�}F{��'9V�q�dE7%"�"�)�?.T�H�'DP���̗n��(�5�C$�p9�':�ia̚�g��H�ݠ|+�Ku"O�����N0��B��<E3���'"O�T(e��3�f��*[�&D��"Ot����Hk���K�A��u�'�ў"~j��#jkʼg�S�T��ȡ�(��?9-O����g��j#�9�|,S�I�`����^��͢e�ĸ�F� ��ϕX��ȓeN�� %��, 8���܌��A��Q>��wK	w��U��dB��B��ȓ4�|۰+Zu��ݺP�åY��h�ʓ7�!�Ǫ�\�lQ �a];�@B�ɺU�L �ˑ7�2�a��5;'B���Y����&��`���᦯˚I��� D�2D�@.e���;R �?��)�6��	!�$�:ab�pW�6�]`Ձ�=m�!�]++��
C�Įn�<{&@ěo�!�d9=� D�&CM4)m���άg�!���@=Z���EU�A�F�t�!�$�	�Х(�!K�DOj�#�L�9�!�D�iPx͒�nթ1�	C��v�!��E�i���a�����YG�!�$KtN��V�O9#cfI��%��6�!�Č�o�:��%��78FJ\�é�!l�!���/3�	��_�T⭨�'��I !�B&k��	���2Y:�9gǞ!�D�q��Zw��'%�Z��e)V�!�D�7Q��À��'����EA�V�!�_�" ��)!JQ>S� %��F��/�!�F����U���R�kRN�!�ԛF��a勅�x?�U
��<�!�$	�J�;%���h���(X��ȓW��P�����-�*��cb�.�6��ȓp�IC��*&W\��ON�O��܄ȓ]��1�%�P#�x7bK8/6&X���R��Fġ�ihm�>4
�D{��O�mp3N2.�z�8'c|!�A	�'�HQ�6&8,ap�VCC�CfP���'��(���C� t"�h�;S�T��'Ħ�{�㉄Y|Ja{GC�Pw���'M��A䀨^/*13Ðys�eJ�'j��5�	347��;2J�5����'@"#��؈w��gJ,O,�p�'�]�S��>~���� ��XY���'���ɇl�?t$I��RJJ���'8�Ekf	�B�إCC?4o2���'݆�X�f�1��#5iC!+���
�'����n� |JI��苶�28�
�'M�*�&Ƕ�>ɑ3��0h���	��� �����_�In�����^)ON�R"O��`�N�5u�nE���J�0IZHAd"O��S�,�N<Y��C���04"O��������iӃč,%��9�"O4�ɗ��#6��K�bEY<�6�?D�D{���7 N��s�Re�Q�&�>D��*��5�I�oߝy�r���/D���D�'_�(�v�ް,�P���$,D�H��c� {�@<!��@�^�� ��>D�Th�ϖ0BZp�t��8 ����l)D�̡`i؈d�B�ײNhD��p�'D� K����@�z��H׹z%<9(5F$D�d�'.H�r�)3�U�1�i� D�0rd�1[w������M�f=D��Ge�Pr~��'�ĩGґ"ō/D��0��O/��a��-GB���� D��9#0e��c�nA�	$��/;D����L�:?� iV"8��Ex��8D�8�`N#2&�$[��I{�����4D�`��D�L)��@�C�NS��8f�8D�L�ᔂmz�l	V M�����;D��be$�����.F
d���1��;D��9v�S�+Dy`VK�!%z@�D�7�O`�.��q���P�I�$�@��Y|\)�w!w���J�cg&(�ȓ{6�<	3��`M�8K&`�,B������G��l��y2�	1u��Ȅ�mΰ�ϸv( ���+9�$��ȓb����� �%�x�x$ӤZ�f<�ȓN�� ��ͳ(^�Ю@�r��]��06"�@�.	��x�R�@��h�ȓc�f�!�*ߙi+��%�L#zP)�ȓ}+rX*��/)���H�'�d��ȓt>}����4����o�<rv���,0X���V��q�# <f����P���0n̍O����!޺9�0$�ȓ[?�LZcbT:WE|MsVF^�
5"%��9^��׃M6R7���p�h���a��q���_	D+��C��J=]����ȓb����OҊx�*dk׎=��E�_�,�|�H�9{�z�N(��x�F�N�<a��ͬ� ���ʮ>m(��Xt�<��\�>��!	 #�y�C�[�<��G�SވHkWił�쐺6��X�<I���<�=��cؾ�n3�`�S�<q*�m�~,3B�ٽ4�b�"\g�<Yd.G�G��+w�Y4
�\)H6Ϟax��GxaH;6����щ*/��u��,��y�%.m�<,ĉ��+P$�/@/�yroB"V��Ҧ��*�Z�����#�y�g4)?��Ʌ*�.)����0J��y
YTY�����8!4��g*��y�&��
�� �%7��a�F�D>�y����Up��o��{ޱ�s����>Q�Oj����Ʉ*����_dV���"OV`�%\G銌��/��Ye�B"O6�rwb�;�f8�(�S��d34"O����d�U������3c��iH�"O<lH��Xn�Q�,��-��9y'"O4<Y���9�U��_�b:����X}�<�a�B�������)Ų]�ŇƓR��0#`��Ӽ4@�@\(Q�*��'/�Ek�*e0�Yj��ˋBK����'4�Psd��<vX�G%�)@�~l���� hhSO�$��ЮM/
���"O���듅c�����ʁ�%"Oکע�<J��\*�����1Cv"Op5�6`]���C�� D�~�"O��Q�2�hI�A�e�F	 "O�`���B�d�sK�2|��y��"O��A�ʑr�q�$��	L*��"O�Xj�܀1���V=����"O�cS��%��|���&�x˧"OP,p���
�긪g�Z��~abC"O�y���e򐈠SLZ�3�:Р�"O
a�i�u���y�Ȏ���S"O>�A�_[4��S��=���T"O��;aH�h�|��eZ<��%"O��a�Nϥi� �3Q%�%D�D�)#"OD9Yq�':RAqVK�6��!`"O�e��K_ƄՓT)�*u�H�"O�s��I)�2�!J��^�(j�"O.M�R��/Q��հh�*~O,A{"O���p�@�K@�<��T�`��"O찠����6*��2���	7��)�"O� ���/��,.��E�!"O�8��ҼqN�	�r瀫:Il�1�"O���F
۶7,l�擽s70�"Ox�9�瘝' ak@f2'�)�2"Oڑ�U�%@�&�$5*4ݡ�"O y�SlӘx�N�S���P�"O�!�c�Ø9��"�l�,�|���"O<��6�m����JĨR�j�{#"Ot���[
O3�E�RDܛ-�F(Q�"O��LV+reH<H��Qخ�J�"O.	���
�`r��,VvR��"O� ��o4T�p�!ɺO��m� "OV�aUjHD��eF��$��$��"O8�"-�04��-��L�h��y��"O�k���q,`�U�H}
���"O�Հ�
��=Vj%�q		�
d~U�G"O�HБK�4�T��K�A�X@�3"O�A���˛@��e����/^��RD"O�d�����%�ebw#��Ĭ�b"Od�j%��KTذ����!H���ۄ"O@���"�@pV���S�4��|�R"O�$s�P���j�W����s "O\�:d��rȾx�1E@blLI؁"O|Bŧ��'��c�mQt�"OZM�&h�@<-2W�W�\BhiH#"Ol\�҉ƙ-��Ur��1�U�"O������x��1�c@�9Q(�\��"O��q�G�-x䐑H��<h�"O�5x�X"w��lS4�ֽj(�X�"Oh��o�%EU�I�&A�_�.lq�"Oذs��	ra�ǣ�>1v��6"O
I1�!��Y����a�� ,�4�x>��rM�P���A{�F���&.D�<B�H@M*$�D-��o}�)��.,D����=}���E�r���j�8D�̐�`Z�S�nt`C� �=dB$�QL5D���C�՞c��	0�ę�=4�y�%5D�##4G,X�h� "�mY� 4D��ʒD�R�<"��gb���/3D��pkT9/�D�2��k��9zF1D� �!eȿe�j%I��1Tku���.D�H17L�U^0�2B��0�4�㴧(D�L2#��$2��x���U�4�vB�)� �� h0@����A&�
AT���"O��Pf	ʏk.���  
0+944ɂ"OpK7*�sT�ѱq̐�.(�$��'!�ܐ��ݷPvh����<	f��U	%D�X��<��r`Y�]du���#D�\�lINz5���9��H�j"D�� �!�%�����!.$0���;D�p�E瓬/���:��X�"b���),D���lX�^��'�&#�&�:��5D��"�kɯ0&����#�8b>�Z�9<OD�$?�	n�Ȱ���S7�iC�(L,)�hC��sY��`�ʡk���0��
��B�I'4S�-�dg� T{\Z�̆8	<�B䉨t�<��f��y�1|2�C䉎p涰K���<}�A���A�C�C� t�H�����6At�p���^�C��,5gPhC�ϩ|�p5a�
.8��![E�=� 
/%d�3�Ԍ1k}�?Q
�
�N$��'ҍ[��)��A\��u��SO�`r7�	��fR�)P�0|���!�l�i�)���	��c�bą�C��膊�b(^hI4��]�ȓ(<�x�*A%�*`�HIi��y��-�QibE 
Ʃ	�
���Q�BѢ��4lZa
�#A���܅���L�T�,m����.�r��ȓk����S�385S�-:X/N��� -"�%��1e^i��%�f�* �ȓ<*( ��׎/W��(�Ɣ�2Pи�ȓ*�&0�	�s�x���G��t�8��2d.-�SW{�j�c턚WWj���f=`�@%T�[�>���VC'���Et��KB�za�H�h�4����ȓDqju�dNa�-4��\S&�ȓN�4q��
�w~�P�0퉓�l ��4�����'B�sd����ʊЄȓQ�h��B*���i�K�+T�Նȓq����U�Y�x)WNI�0.���ȓiB�X0����U��c�|�j|�ȓU�T�yp(Ҵ��l�"ɔzv��� ��신��1<�>��r�?�Z��ȓ.�,��dn�.��,y@�[.|͆ȓ�=��n��!�c��	�ȓJ�a�WY�rɁA,�S�6Y�ȓ$w������n����I�i�l�ȓ9Z�a��Iօ)\��BbfN�4����E�@��d�N.T:�}�E��$�^��ȓsv��I1��1Y��������ȓ,��m(s��.:��>��P��n��8��^,�4�rLޤb�ZB��t��9� V��x�Ɇ�n�B�2a¾YӔ��CY��ѢG$b�B�I�t� �C��W�ș�&H8=�HC�ɹ ФM�3�C+=���@�J�6��C�	�f��0v�ҏg�E�a���C�	=n �XR�똞]G�R�*N;�C�I'U�V!��CAY�D�
��L�hz�C�	 GS�LҰ�S�@���(p��0P6zC�I6F�fPB��2B��A1\$h�bC䉗�\�(�3}���E�)[�2C�ɾ�M����\��fH�)��Մ�g�x�@�[8w��E���
>f|�M��L���Q�&�)��1�-�>9'6݅ȓ/+�`�+����Hr��?� ���S�? 6m��Ç�^�H�R 	�k�Ҁ�d"O����<]q���qǈ�>�^��"O*	AԀ�4D�,Sл�����"O�]&��4����&d	�����"O�B��)H6��#��Цv�CC"O\��f���a�	����6"O�	P ע4z�𮊝)�}I"O`L;V�9{L�!�L�A0�"O�Hs Z10�� KULɏ7�ira"O�M��Ĭz���@ߴG"�p�"O"�铈ݟ��E�E[�k�@@�F"O6%bE*5R��ip
_��v�k"O�=����mw|(�(��^\���"O2��s�/t@B��?BE�1`�"O��hq�Bxu�#����~ pR"OiK�����:�e�L�F�S2"O8E�W�o(H%['�J�4oJ<��"Oz�A hG'��<#�%c��a�"O�4ˇ���*n�
�SJ�}:6"Ox5y��K9���QC�6P�	0�"O��*4$ZN"\�$ �b�	0�"OԈ���"�0��e\-Q0D�G"OD��O��T���"c]2W䶴�%"OԃK�$�\��!�>@��i/�y� ��LSB$84�����6�y"l�1�V�1�ɰ)���w�E��y�3iB<k��Ŭ)D�!ҵ((�yrς,\��y���� ��a5K���y��Ӎ9N�A FˈK<$��$	���yR��8V9��G�=�r����N��y���#QB��D�_�4�:P�-�yr  /�(��F L�3G~Xhb���y���fO�CR�^71�ʌ�$�$�y���
��Iq0��.�@ ��޵�yr �Nwl��G�)m��L�y�Z��T�7�O�(��C���yh�ȞT�غl~��A�ퟣ�y��ӱ=��@��=N8�t(UIH$�y�LG
�Zq��z��J����y2n�	o�Ŋ�����i����%�yB�ޒ98,y�kǰOݤ)"�%Ƥ�yr��v-�n߇`4\3Rm�*�y��	y�!r��^�!�ݢQ߸�yr]2}���T�Ķn4��@Q`�;�y�	O�"�����c}A�6�y��ߨsq��#�Y? d�1�M�y�)V�Dg��*�X� ���p�i�=�y���w_:8Q����u�B`�C���y2�q;����s-Xm�c���y�͖	���Jg喞:������Y�y�`�2J�.�*ƊV�,�\lI�&�y� CTTL��D��W%X:��Ά�y�披a����3�+K����գڪ�y�G-Q�x�ө�.?�\��W�y�H�	,&!єa 40�\���'��y�M�/{�0���A"8��˱���y��$w�ܸ�lP�P�N��O	��yA[誰�E�*E�P�!<�"C��-i�ȸ3�V i,Qo�"+��B�ɸ;�dp�͜��qsTF�+��B�I�g���A���0�����G�!�B�k�8	3�.Q�p���R��b�B�ɷ4����d/�EeN���&bB�	>Y�@3���B�>�'j��(B�)� rԩ����QsP���p�""O�!Y� K�c{`�U$�
�t��p"OJ$�R���Xt B ƽ�
e*f"O$Ejg�A��@9H��L(d)�4��"Oj�s�� '�F���ǁS��=@�"O,,�兊/�jI�@TTux�0"O��!th�a  0Q@�]Y]�"O"D:b$�lŦX �oR&WRD@"O0�P���z��0I�+NjH���"O.�a@h!�ܕ B�	e0`���"O�X�솤>J��W�ܠf:����"O����IW���8!p�Ϟ!-�9��"O�i�O�&
B� �'Y"����d"O.rc��!WÞ-���<1��j"OxDS��N���	GD���Z�q"O����j޿Q�$����=N�PY
�"Ot$2.Z�4��Az��;O�`AF"O`HqEoM�U�H亠�)!8T1�"O.�iJ�?�0�)sE�9 <�;�"O�`(ժˏ�T� &<� �S�"O�h�Q��	N�-U���;$�7�yrjڝ�6��Ȍl�8��l���y��a�ŋ�+��b킅��E��y��iM��*���G�DPQP��y�&ɘZ��z�L�*���ρ�y����^}[�慮W�"�H��yb�A7�*�:$k7S`$$`���#�yr!M�*:i&E�@����	-�y��P�_"�U�7��@����#��y��	N<�����5M���ŉ��y�V+Ჴb d�;/��H�BRG�<���J�G\:�cs L�t��P��^�<�B ��2�T�@+�ţ�'_2;�C�ɩ�ځz�m�
 Dy���۞.VlC�ɜyv2aH�i_4iG<mJ"��9Y�C�I�,��|q��%��R�"�8�/D��!r ӏZ�t����e2�k+D��H�E����̼*z�X$O&D��"����4���L�3G�*'%D�� �ҕN���Q�cݳ�r���>D�� D�FP!p��B1``i�>D�dI�e��.
J����%P����)D�d�T� �RJ��ア�2�����+D�,+B�@�%���T�W9^�<<��)D�`��˫x�(��dԗ��5q�()D�8X��L�_� ��EqA�dв(D�l��6M���Q�m������$D�4bB&��G���	�8��8�,$D�8H6aE�*,S�ș=�@�S�!D��b��B�kl���m��W���"G?D���5�ʞ-��MX%L� \:P���=D��S#bE�6
�� �%�� ��C�7D�4	EK�,ip�H9��Vi�pd�)D����'@:	q#��T�-q��Sw�(D���uF�-R-x�W�&��ts�'D��K�Ɏ�.tHզ�3�TI�m2T�Pq�AT�)�$��(G;C#���e"O��[���<N��ggH���̀"Oj�:����{��ग़�p�҂"O� ����T>��rař���{�"O���c�3UXn�w[*[)dEr�"OR<�C!O�3v-(4�Y7y|�)�"O0t9��M�K�NG:Q{�i"O�]Z��S�l�*�.�>�4�b"O� .����*��@ N�=K>��7"Ov�0r������^�1��"O�u[�J�G'���R�Ȧgs� �"O��3�Oѷ�~! f
T`�Es"O���s�(5���ֺ$��xr�"Ozx�բ@�HT9KU�F�D�"O����2!����/���X1"O"BC��r:}�P�Cd�|R"O���߃b��ɉ^�4�v�rs"O\�R(�"-���`նq��Q��"Ole�%��� �K��'&J�{7"Ojh�Pl�;-��%S -¯�`��"O(�@��<=��2�+�-E
u��"OX��i��"�C�̓#��H�"O`4�1���L�ʗ�[4X4@�3"O&}bj�5a p�#B�qɌ�� #!D�ȱ�Gz���I7t�4��D2D�\�G�<v,=8s�E9�
�Z1�1D�!��]�>s��Hv�e��$D� E�߷0�djLY�kڌ��e$D�@(Bh��X8�#�*����ad#D�,�a��*J]`�Hւ,Y���7�?D��S�On���c�Α]7腡�� D�lh��F���كN�=c���`"�#D���T�;W�\Q+�@fۤT���'D��@@+�'�^Y����#Dy�u;�9D�<�UCV�s�9`ү��N+�8@Ӡ,D�$ccG�'��`�SI�vК3,D��JK�#�(i�*K�~nV��@(D�hapϝ�D��µ	�+fN`��F�%D�x�`�^&v�Жj���Zk��"D�pR�h�
=|0���Y��a��=D��(�`}_�=H�'@(2 h��;D��۠?j��2b���%D�H�6ǂ	d�6��oB�Z#0U�W�%D�I5$�=>��<I3�_	ac��18D��h���)G�}���&k �5D�A�e �J��e�o��Q�� D��5�E*\��U+T�'. �)�=D���v�W�J��C`b��a�h=D��h�/
�t����)�Z���R֭<D�$��]�k�H��׍ߤ?���AE+9D�dI]rF�4��Y<d���O��!�D��Q|<���#W�bXi)VhͯH�!���&��9Y�!�Ա0˸o�!��ƄG��<����;:�E�I�T8!�k4� z���1B5��d&�o�!�!;'0�j@��5'�`Q�E�:B�!�dϯ#S���'�$>{�ݐb%2!z!��
��1H�FF�B`�,[&#� �!�ƨM����M��b�ys�S`!���i�:����#��j���!=I!�$Z-��d �w�\�����%�!�$�>S�%�C^��Ġ�!MP�K~!���S>�(��R���+"���#!�ă9!����� I�eeDY�7�!�d�j�K�g��(;���b�,�!��T�-�����_+��A	��!�$ݍ{�t��"厫aJ�Dł�9�!���&%�����_�|]l5��Lx�!�1A������S tH���N.�!�+|�hIH_�Op�hYv�n�!��ɲc��ݰ�Nވ.I�,�r!R�q!�$�n��Q�i\%�28�p#�=!�� hի4��7�x8Ã*=x"OT��e�>hتi�$Yx*�C�"O\��s�p�(���:�H(�"O��R�
�[��S��V�"O�PR�O��Lz�dh�	594$��"Or�c���,<H�E:w�۪$`a�"ONx��f��6lP`���()�|ف"O���(�;0�m1��	'<:��)"_�����<�2B-9���s����e���V�OX��O�����2:����eo_�T��2�"O��ી�I���s�X��tڦ�,\Ob|�t�T�)(�)���R"JDQ!�'ɱO�8rA�9H�����	Ϻ@�M"O�٢���o���x�h��*�<�b"O\}ؒ��l�Q��}���A"OP\��H�9.ѳ��H�C�| ��Ii�O��ed��[L\�M�@�x�	�'�8��wC��,�dE3DX�2'�Th
�'44׀A�>�(�n�A��0
�'��4��J��n�J�O�?�6�Y	�'�Z��AfZk��Xz�GL�Y����#OMA�n��ՙ���=�2�)�Z�X��I�80E��-��j�B��R����.lO��'��5"V���X��I]�V*4�
듍�����,T�A��+�L�"���|��1}J|�OT$ap �8��Ȑ�kD.X|�0Y��Iw���ɓ�~w�� ��^�x�f�h����M�����,�����!J�]مF	� ~�  �¥W����G{�x�l���[+R����s���-�X��=D���c��.�H����C���m���6F隍"G}��5�Aլ���)��:��-zE�-�p>�ܴ��dǪ\�L4���D
νȴ+�m��D�O���$� ?�ҝ������J�iX�qa|��|b��8���kP
­l��Z�o[(�y⫚�Z�=*�M	�8�r aZ-�y2�5K���xC�D��q1�
�y2�>/��	��Ɩ����ّ�yr��n��|��C&N*ƵZ"����?�" �OdU�C� �ɀ#⍍s7�9�"O.̚��N$.�b� ߪ'8A�&Z�|D{��i��!���V���CEC^4A�!�V8o��h��4��aR�a��:��d���=���ٟ- XI����c(6D�� N9T�!�d�.�%9d��!V�T�� �!���P���NآB\��E�j�axґ�$'���_�^�ha�i�<kk����j(D����'��� @��ϛ�6�����)D�l j�. P��#�m��(�R��(D���C8u�<@��eD< ����� 4���� a}*�hLW�6m  ����~�<����h#�q���[�eGt���C�S��i�0��h{*l{��{���8 �6�6"O�WN˔w��!CH�
�D�в��G���O���8�

'߮��CAؗ?�M�	�'��H� ��P� ��Fʚ+�Z	�'t}� ݼWw���ա�N���	�'j�8��U�K���˧�0`�@�'�T2� �E� ���n)C����L�R}�_��S�'~d4��\.Hq!V��!J�h�rs� "Ar�C�^C@���R�w2F���L�-���C؟̣�
X��6�e��<^��D�=LOV��$I'w�)�2�?T� <Q2�<Q�	p�'2�P�H�<.�l��c�.. l[�'�J%���j��Ӗ�O������� Xr��.C��{�bE�	��e�b�|�~zǥ~�����߭iY��'�ě /��;D�@���GEJ��&��n$#�8�	X?	���O��P1$���y��1*Z�����'�X����$�,�%��O/NY��'{$�Dy���S�w*��p�;Y��t�\��yRb�1��H�a�N��y�Sj���y2�\ 0�q5��d{�����	�8�1O�t��'i,-@��vt$�C �<?����\�$�8.\��aK@�3c���S�; x��^��$}J|�'N�dp0ۖ!���a��<rZI���HOډKtM}0�!�@X�Z� R!X�(���)�' ��9z�ƛW�Ti�	�i���z�r,:d�ЇW�0pjS7y�
����M#𧒟*�<#���,W��+4�TC�'�Q�$j��'v0�!��ҖmS����ʳ>34����D�O�#}2񏗙0�=�ē��H�1/����D#��?#<9E�Ѱe6��kL(|����Bk���'��Q� G �
�:e`D�`(Ru�dO��xr�6)뀵3$�M�t\�կ�%�0=�شj��'�P�N1`RHXE�ٰ �.W<D�4aѩQ$Bht�U��.?X��� 2LO(�(C���~�8�8Q&}��_�<Q��	!+v}{K�Is�M("�X̓�hO1�d��!���>y�3�\�⩺�"O<�A�i�f�Ң�l�0U� "O1B�m��;e$TZ �5_��T�"Ol����	�����_'q�q�"Ohx�À_�)Sɠ U�Bn"\)C"O4�;�]��0����>?���3 "O6�� &ʹ���3Ɲ�5NĈ"Olɒ5 �
���B�%�r4��JP"O��26�3\�b�.C�B$,���"O��pDO��	��Ś4��;n��Ɂ"OD�	AfO�h
�`�
���I�"O4�xA�ʔk�͚`ϗS�\��"O���J>Q������R*F��IS"O
��E�A�ay��Q�ϣd'�|d"O�ur�B���(�
5�@�1"Oܝ��n�ex�@+�bP5c<TA��"O^���ܼf�¤��A�" &�"O�\g�'D=ZQ��O�V�dH �[����ɸG�1R���< Y���g��}|>C䉳	d���
"w�
��7��C�	�<�r1 �O�_��y1�e�B�#<я��?�I��¹G��	�+�&_֕x0%3D�p���d��іǖ�B��L�X��I5�hO�>�ï�e}�U�bJ�i��()�@;�O��y�m}�]���5"GRX�cIP�y��* o���$j�m�Si ���<!���� (�r��L���sd!���^��d�e�۵V v}ӵe�ab!�D�9w^�4 �+7|!�FK��#1!򄀝#� �.��N����J
+��Ic��x�c(�)(<Txa	G.s�	P
3D�䩡�J�R4�ّ%_'K�b��@�1D�@�l��.H�C: �P`�C�9D��05ir
��� ��[���#D�k���xP*�� �M�eR�h��"D��a>{ڌ
�C
`�D�BD`!D��X�ɝ�u��$-�=�8��3D��*�*2���a�K�e��ٱi1D�03�)\02���o�%� 4S �.D�`Q�d�,���Kp��������!D�� f9���]�x�>x�"^!"MZ�Y""O�u@¯@�U	�j�lW?$��b�"OȍD��]�v����X7p�k�"O ����e���z8���"OԴu4w�z�A$A�Dl�0"v"O�������| 3F;@2=�#"O���i��_��a+q�5C�*t!��I����N4�yq��X4��Q��2y!���{�R���2^0c����!�7m�޼3f�	�:i�I�c!�$�!HW�D hH \��́g�̅L�!�DC�?/�����'.x��h�>�!�_�^��Ib�+���b��҃zz!��ՁAv�TAƆ;v��ӵ�6>�!�	��a7m"j~e��[�fT!�޲N�|QZuPF4`� ���K�!�Z��A�S  
T<H\���	u�!�Ų%�F���K�O<�e�`��8�!���L�� e�!-7Tq(v,�g�!򤍥lj�CK���08���z�!��]".צ��KZt����JY�!�Oj-�L2��3	/(�����A!�� r!,��w߾V�J'�< !�ē7�H�!T"}�"(ZE	%�!�dq+R��LS�LƐ$��Es!�ė�2Ӧ��C�����0mF�?e!�$�)�zx2�&�PQ��A�>{]!�$ߗ�T�r��\t�=c6ʑ�P*!��T9��� ߉~~�hr��2�!�d�S���(��gb�a��	^k!򄂆#��H ��V��88�E(@h!�d�.�X�� ���{¦M�eL!�D�/]�
q����9@�� G�L�n�!��^��\A�K��W�N1C�;�!��Ƃv���Ad��B�]Hu�Ѝx!��MY��6��+T9��ܐs^!���}>J�i�'n��u1��45@!�DS�|�R<1�ʆ�z��m�Q(!��4�r�ɵ�'j�4����.A!�_�8���YTD)J���a�;E'!��%�������i[�23���?�1O�J�kZ+8�V�"��XF&��F�'K����27�H;�̆�F!�$N�P�dD�d�D
��h)�D�!�d1+� Dk0*�|B�had�)�!�Dז��ʷ�X�0=�5SQ���|!�DʡTH�-�L[�n�lYы^�N`!�$1\�,l�`K;G� 1#��j�!�D^.(o�����V�#��}�&C� N!����~���6G�8��d����!���=�lJ&J��?u�h�d�K�;�!�$T�!D.]{�K�x(�9RM��!�Ï��Q��e�;gǲ��c� �!��+ai捻��ȞT�&]�ç�	
�!��(��m��G�6B� `�݅4�!���;,�F8��+����d�Y�!� �"x�u)��D�4�#��Ĺ�!�y�JI��&N+}���D�߇�!�ųjz (�,�u�٢��c!�N�\hD�B��.b�l�5�W� k!�dP	s;b��҉D�u���m߁SG!�$ټ7���Au��>���+� '!�D�0sdhz�D�B�rIy��Y#�!��ޑ4����V�Ð1��;�o�)|M!�ĕ1%k[�2T�l��V�ݠl�!�� �se��0�B� pJ�^����"OVH��)�"�X�c��_ �8}��"O�����b�f �g�0�"O�Y�'��0�s��1A��9��"O:,pEk�>b��X�4�U�.��"O���-��C��s�a�`��9�"O<m��h6.?����W�H* �%"OP����6R�$[bݦ
nʥ�r"Oh\��$��2 �nH�%G�� "O��Q1�K,h����clO�=D���"OZ� �` fI^��ЎR1orH,2r"O�@���'x�=���J�~z��ô"O�x��8>&�Y�j�Lo��"OV�X�`
����9�}!"OJ�1f�S�z�N|��
��K@iX�"O��@��Ѷ�׉S/KIX�yV"O�%��kHg�2h�h�XPҶ"O�p�䅧-�qI��H�Y�<5cu"OF��Q+O$z��`��{��P'"O�Pp�OC1���q+�,@�"O�U��BQ�JY�-XU�Ȋy��"Oj�"¼Ee ���I8\�H1 "OH�	V*
n�P����?gDT`�A"O@	�傅
�lIhp;QH�
""O����.�;�r�c���D(��"O$��	J�y��!�'e�	y$�EQ"O�	�*E�v���z����9��U"OJ�w�\�Va,�P�#�^f�5�"OxP����m���� /n��d"O���Ւ.	�C�`�0_�I�"O&��u�SS�����@�D�1�%"OJM�aR�p�\m��uaR%I5�%D�@��NԮI8�,I�N� �%D��� N<)9��9�VpI�d�<)� ʔ2@��S	ӓS��x���u�,;��N�a��e��ɝU�)�$jR�~�y��p�b]�U,ĤK3|a�Ovŉ[�#��x.�&C4
��,/Q�,٢��+g��b(�g�FjT���	d-�$B'p�U�ȓC5���$���G���;5O��!�\8t�	,K��*$�J�Q��)���F�_&8"~dr�/ܧA�,�a=D��;`
��4�1/)� ���⤟�`e�@��`y)t��]X�(�#X
�ā��+�`3�9�O�+� +a��;
5Ӱ�2R���3�.h��Џ^�tC�	aB��ᔬ�?6��dZ`"�T�.�<Y�	�gN���4L�>��O�j����шw��{���u�ԍ�'�"!ခ��o����d>d]1i,�QX}^��S��?�"�<���nΞV�*q��.�A�<A���3׮���F���EȡN}?�V�6}ش�%��<�®�"Bl�K���>]��C"OVX�@�'.R�H4�K$.��6G�*;�DͺG
�_�B�	�u���#kU���ԗ ��=Ib�ĝ��pȌ�iҗc�B�p�kf��A�#���B'!�dû'�l��f��J�Ti��i�r�Q��k��	l�>�X�M�)���h�d�y��h*�<�V⑒p����$V t��@�d]�K���13��Fq��I�Q�d�-���t&�$#����n�^���y$�D(`颅дb�CC�I�H�6xrŭ�UΥ��M��B^���.C'W�^Q@U�[�:��q�;�>lZ�m�D�I�?qbխB���M� R�"ljP�#��+�ax/��`qC�i ���ï�l�aE$�t��eJ����X&N��4B�TB��8�j�榵�'q���v��qj��֓4�$���$�U2��M �	�f\�h'	��7�@��d�-O ��E	t���P#�ȅ[N�n��m떝�$͜�(�	�@˥O���ܧj�Š����0=�"��;��R!�H�
ߠ8���V4-��I��M�~������.�hu��ʘ�	9�i]�m]Ma5k�R�$���ȏd���IN;,�THo$�OB��B!	=h��(�"?ڼ�����#dҌ��V�� &D�!�M
�OR-Bvm�<h��8��\���D�2i��q{�� �Q��-d�E�F�C�bMd:�ɟ��=��)ڐ/�=��*{^h�)�I��\ڲi���K�`CkܼQ�(�u-;Tl=��Z���$		�nӬ��"�)�	c,��"4mD�2�	󄪋�g��˓����L�(-o��;�d��>�U3�M��i�2��bfX�pI�ם�36�b*
�)v䄈����-�牬$������	*�x���9;�����)�n�@+�e���o��B��e���,�p]Ҡ�v~��)�O�b�8��g����ӬW�Z+���P��9u���`�`�U�x��DU.W�N@�ƇI�J&��7J�rĘX�����mp�̂❱{� q0g�	�9�ם������ś�%*&�C�.�B}�%��C�9��+��D�;���6`���'(�&1�%M5Y8xI��->�>�����'P�h�u�{��i>��ڭ����N<QQ�U�ʥu$��!�T9�b�ry���������H�T?�B�`ވh���5/#����%Տ>��r�a؞���>TJ͈���/���I�pɢ�)����>���#@�&d�$�O���'���H��Q&?��g@���c��^�aV`���"G0P�5�u��F�T`��X��<�U��m.�$��5]���'4bV���
�As�'	���[w]<��/�/��O�Z��@JO�>Q��	͸F��-(A�$A�p��c?����I^V��1aӢ�,J�\9��I+,��0�i����O�qr�"8uNduQ��N����W�0��ME2S.�#��>E��J<6J�*�&�/V��g/̾��D�54Y@��N=z`ayR��#�^#��ܦ|B��*۱Tp:�'�(�T�f���~B�Z�Up4��+��x(���<
߶#p��$N����I>Q��0DUGD�Ii���I�h��O@iYd�ĉ(,������<d�>āH̥E&�Jr~Jџ`�p�"4�%�@���Ї 鲉�"]_�X�2�	�y��Pê��v�5��
��<��$[�aB�h�?��)�'

�1[ %�8<Z$j�X�Ct�!��xT�Y1r�Y�����'�[ rċO>	�^Y%z��|�<y֌��Iܲ	��Y���u�v��{(<a�U�Q��i*��T�
Sry�L�,lF%�?���e�'-hF�9���,8�P�b!D�<Q��:P4|��K��R�$��!D�H���+άdO#f�v�1��-D��s��QB��h��]�ipH�5f(D� �u/�)N� I�B'e!Ftеd'D�̳�b��$�"1Q	[�X�*����0D����͑R�T��UiR�X�RL���/D��Bg�Q�
S�\*�e���:̚'�+D��{O��s�dda���39uؔц*<D�d(砏�i�Դco��;h�zV:D��Y�"L�|��L!FAX }i6��t"D�$A$@�6�D��$�8���dI%D���� �:�����Sߌ ���$D�옔�\�%o�0[�K�|��@�@A!D��ңaP�f� ��UH5[�xs>D�P����*pjx��/�l�+7?D��ҲlĽ&�H5��}�\ɸT�.D����n�,��4��EĦL����#,D��(�,^1`�h�AMI���"9D����b!���"@I��ِ�4D�4�U�&~���S��-����&D�(k��
8s-Xe�Ic�q�5�&D�h�Å7`��`E@75�Fu*1#vӺ�I�&8��>�b��J*���낹9jj$���B���U��46�A��O�|9t�P�A|�L�3LM�o] �)s"O�e��E�(�TB��f9����x�(�#�z)%��6MZ�D�Dgjam�O&��zI�$�q��'?�s��#V� Q�௛�/��@٥��e͔=z�*�O�!���H߸��C|�"^$(U.ػ��Ć>N�VΊzy��P� <�r!���c㠤���K�7��	�DJ�Vg)�Q��, 9㶼P��4O 0S�-�f��Y7G�!��"SN�Y7 G�9���S靲k�!�D�/8���Y�#/���ό-����GZ(�k^<t)�e�5=�Q>{��*^�x�K"�T�q���k 8D����0��pP�L�?�ukW�<U5��K��H�D��̢�#��r�ʓ��b�����N�~X^@�an�o)|���=�O����.� ��
� ��Vظ�f�A���vJ̯
�z�*ď?l�h��'H�T�c� b���Ň6[H����dNz�2T�U�E%�@q��^� ��\�U�~�f����	�A�r��(D����\
O0��s� ��S������<YO]+zZ�Z�N�-��	�Bӌ���{�n��~}D��ë�(�ɉ�"O*����T����0��˛`�j�ax�Z=)�ʛ�H��!&��s��OI1O��*/K�y�X��m�;h���;A�'e��s�X'Zi�A�`�e�hT�4K�8\o�Q�%��b��,F�N�az�a�0?�j�;3K�2I�D�����O�гE/-a4\��E��>�d  �O _����I&{F<�0�P�F4�B�I�[���nV�"X�#	L� _~�iF�7&S�Y��8�U z�ģ|B���/Wh}����Kx9;@C	C�<it�i��PJg���1V:0�Bl��C;���vl
$ut*�C��-�8��|�<��&Z)�T�q&�6~<1k��E(<a#-T�/&�:�[�=��A9���ur�r��¨@�u�S����=�F�q��]
G�K,(����K|8� �GI<,8��0��-�D�mZ�'߆9�$"^*vV4�8�ϑ=��B�	�c{�T0�i�pUv����j��O���U!=���F,��h�@�Y�����ĚS�2@O�hJ�"O24*�b��R���WhK�q"�(��G�##/�"M��AF�/�g~��P-bѐ��X�F��}�Pꚭ�y�)�8A>�����">
�{3�S��M+ �'0����K:w�̴��.A�	����dV4z�!�D����m�.��"�cB��!򤒋z�m+�j��D�����NJ!�D/j�PIr�ةc������p6!�4(np�q�B20U�5�w�D!��2�8�a�͎eM��!��z�!�D�8;r����(��a`B��!���-	������3�����B?b!�d˓I�`pJ�M�'�4ȒLܹ`f!�D�>=�͡���ktp������cu!�"��p����g �Pf �]�!�d��c��E����*�"��p�i�!�$�`y^��$
�s��#t�HZ�!��ȫg��ce_ݖpU�Ʈm!��hѲB#�,R�0x�3+�!�Ğ%���fHժT� ��BA�m�!��
?+h� 㪔�R6�6!H�!�$ϼA��w璅�lE0�a_�!�$Q�ir����R
H���#၅��!���|瞤( �DX7��G�+�!�¤>� ЗEW7_5.!
V�ۗT�!�$�2z��;��E���
HH�c�!�D!n&5R�'�i�g��!���r��
��G�n��y�À�!���c::���^�'�t�@��	|�!�d�/S�f����l�"�����(�!�Dz��XJ�d�8j��U��e��a�!��"'-�A��K���0V�U�*_!��)�����ŉ
.�$�3���!��K�dSB4�ӏ�w�&���b֧9!���V\�P+�)ŋRt�V��_%!�*x��5S�g�~K*%Rנh!�D��^>���:�$�� �$�!�ʔ��r��	:�B���� �!��I�e� ԑ��G�Xu�k�+�!�D���z}Zӫ��H�XA!��ҞnJ!�DO�'�5�DF�O���`@(0u\!�"[�2`�7^���a凁5&!��A�I}@�Z��*[�`<s`Ǉt&!�D�� ��p�/��]��ijd��4<�!�US�,�1�����遵�N�Mr!�� 3���&�q$�(�nCT
!�� ��1��Ύw�b��QFD5s�B���"O>Q���o�yqW�Ŀ�>l"O((�����˗OŜB��A��"OFe˒��*v�<�8,�.���g"Ot[�6Tj��e&Q�xɊP�0"O`|B���><��V5-D`��"O�p��A�2AA2����A6a��ۢ"O�� �`� O@�
D��;:�b��"Ot��,@�3kP���jZ��B"O��`��F��L  ��)~�;4"O�EꂉJ�M��&LA�!��#�"O�L�%�_wנ%����F��<"�"O��+�X!M���K��P�d���"ON]�e��4u2�q�G�ٰd��xY�"O&��׊L*C>�mA�(w��1R�"O���(݄}0�Ͳ�%M�/�v��"O0�{��T
T�$hU�.$�V�a�"O"�j�+I�8r�8Y����J�z�1�"O���e� 15����
�r"O���+\�\�(��Q2I��yz"O�8K�D�2f� q��J�D��"O���o�<���(��سB��""O��������΋�S�=K4"O^��7�}�]�E-Պ$*\�	q"O�!�3N��"4��C�J�!b�$b"O,X��#Iy��È�$mW�%CC"Od�B��Z��麴$A%J$ �c�"O��̔�M���Q�Mח/L0�P#"ODؙq&�D��D3��HM��!"Oġ��i��QG �ӅT9 *Y:2"OK������7k�X�`'��yB��8�r����D��`� ���yB��+�����ٔ
j���g��-�yRo��26~��FH�	�� b����yb�-V*8؉2+\������/�y�*��W������֭L聑 ��	�y���Evi� ��*
B�@ ���y�jɨ&�*h�C����+PGY1���H`T�� LOZI�l�\|	�c�P�9�|�;��'rT�h'J*#��� �f�f��T�h�:=v�+�`�Mh<9 �=�T�$���*�"_]�'.��	Pc׊:�@�4�	X�j��R�<>�j�z� ̕$~!�DA��HݲŢ���t�Wa��f���A�U/^&�u��+�wy���'�����¡[�F1�EHQ"�-r�'��c�ɇY�a��ǅ|�V�'<N�:@�	(82:�+��'�V�I�gdQ̤Z%C	vxHM[�$E��A����a\��(�//D��t�Y153�Q9�`��x"�[6C�,��4v��l���aZQ�$8��j��iz�Z�9 :�F!O$`����gI^979��ȓn�|���o\<+�$XT�O�3�<�L�l���s�˃GW�)����L��i]�pCD�����:D�\#G�)�n�S�Q6o�-(a���HQ$�\e��e�5(IX��a��J�R�J��H,{�괠UD �On�I�2��0{���98�\qp�����i���<��x�"�nf��s��ۮ�!A�˒��hO4��R�g�^"|��*ۃM欤	p��*ֶ���kb�<�G�	3։)��P ��\D�'e�#�X�O�"y�AQ�%TH��2������(O�X1�KK�=�nǼ2B�Xդ&Nn�8�HT�<!��WHBi�L>%>� 1��)���'/��d�������a�^� �C�	(�E�h��1��YccFE�~ވs4`��l�r��45aZh�G��8F
Q�f��N���?M�hZ��L���
:f\�2���  axrj��]Pr�!�i&A� ۤ�~�i�jp0�" ��#R��i��d���������'`���hu:� �Dʹv���r� ;8\|S�f��zy剁A��H��՛ ����\�1J� `�N�X�!@o(��� ��)�*W�-�墧��OPv���O�xa�>��i�
ӓ\� �ˆ1�f����#���᥉�x(+-_����\�V��1۟N������~�؂D�F��8A��2pzP� �h���֒E��!���w���c�V(� ���a��w�l� �nκ=�v�����*i\�!��V�u��˫OTAې��R��=	)��e� Y�v��@&�L����$>M��z�����HSMӼfE�]b���"G� �s����F6PI�-]85�

 �tҴ=ADS��QV�"U
��)�	�=�	@)۔M�l� U� �8&˓mV8)�����X��υk
H�E0&N=I���F]���lB:�[�F����j�N�6�^��>7�t�[)t�&���(������WI(�0+��у9�؄n�>V��c	e�0瓘T \U��O*�<S�@��;�ޘb�J�e�$���J1�"2o��4d���Č3�tU0c!@/��	�C�^�(�y�GȆ7L�RL02 ��U�y������A��L���M?)�~�C�����Q@���5����!����'tM:��Y���M�@
R�0<]P�D�"UA��S0Nݕ��i>�r��t�d M<��LX*����xȜ��&FyB#�9g��p�F[�T?)0S.F�1��!4�:4q�@C�d�X�F�B�����D,)�	�j�"L��	�I��1�Ѵ^6$��#����!�L�@ЇA�4j	$�'?A�ǁ����dn�'lJ���cE���q�A5y��\[R�\��eg�!���P�ҐuR[�, E(Q*b�	40�'A�D�\w�P�������O+�]����d 	�鑍Q�Z)R��ңzL�q 䈧�ħg�f��f��>��Hc�&@�E{v/V�o����c�52��)��L�WbҢX���#�XH�0B�ʵ<��6ea8��H9}��)�*o � '�R׋��S�`�ѫOʁ��C�1��B�'��ȪP� �dSv��M����I.}�L�2�x�kg���'�ܥ����az�;1���Ӟ�"u��0�����'���з��.�QY�%�$~3r��baԻI�@M����U�	T4���L+�'i���`!�B��&�E��F҇�LF~ �X�S ZS����?5�P\q5�ժ�^C�I��x��R� ����D x�˓Kc���!�ӧ(�p%P�ɑ/e�v�T��-@H�p"O0��rJڃp4��2�&�$�f&#���&
�.�0F��dA��`D!Tk��p���
x��q��;U����Sg�oԄU@�,��x2%�	h���jS�H$[K�%�b���y���/"��eːQ+�
3%Ɍ�y2 �/t�̻�AQJ��8@4M
)�y� 3�,�l��Fa�0XNX	�'�<!k�C��!�5�I  ��]��'2��ǀK�V��{&��7$���	�'(8y��E3 ��a�`[	
�u
�'���+3V�����&0tb�y �']:Đ!��=~��I@��k�� 
�'��z�������b 
pl��':�@*LZ@is���
�n��'���[�n�,LV|\QdE�vȸ��'�:@��bԭy���s�ƤXY( �'z����*�<d�&��C�Q+dP<P
�'�~X#�׌U�:��FF� e���	�'E0�sN�h���S�L�a�'dv�Itn�v��P����2�%
�'�H�xA��\�	�q%Bq�	�'�T=�s�]�e�<�a�(1��-�'�4�e��R>��M�-�|Z�'S�F��b��h�F&_A�� �'iF]r��{�"��UM^�'��<��'u�8Xs ��cP�͹�hޞ��)��'���{�� =W�L���&E% fV[�'����ƿ?6� �M��.̉�'g��[� �)}���8�:4P���'�r��\,��V��~xj���4�y�&��;p@i�C&.G��}�Q��y��M�s�j��<�����޾�y�/��jlxZ�T�,�`o�y��?f�]��!q�
	��V��y���4N`��B�.Z�rB,��܄�y
� PtH��ӈEZ:��l t�J*O��B�ټ.����Y������'�]R�h�I��	�������'��(��E[D�n���cV��T��'C��q��59bJh93��VIn���'rep��(��A%KI����Qb\���>��:=�6�k���P��ȩT�[I�<��i�5B�Vk4g
��"���/�E�kv�c#a'���v���8.<���H�)S�	8E"O 8� �s��j'�;(M����@�gb}p �>	@?�gy�H�I�FI���)~Z��k��y��ńW�2ų�,�X����M;c�X\H�n�>ƾ���uf`ɡC�)�����ƴ�뉻g<	�DcD:3/��(��Hw捋"�tLi#"4"!򄊆5���8�d۟kˎEѵ����qO����C�	K^:���iT�
��s�XG�vY���E�w�!�$Ѽll��b� 8A����*���F��"�U�T�|�'sn��T%�h'T(2UA�b�옣�'"�  �N}�#�Vd�,��aZXJ�!Ԇ�0>iw���_1���ɑ1mT�Y�G\��xb4��sQ>�7O�rg��R��a���p0n��"O�e�u* ����a��@����C���=����%6�bF
�+��ɻ�n�K3J��@�ȓJ|x0�D�͠��ț��t�B)��ǇHEqO�}���&�9�F�$S$��5��7��ȓ4�ެTI����cf"Q��}��&�L��տ^�9�BAO�mB&�ȓo�H8J��@?v2�r@FCx�PԇȓsHȍ	��0%��A��,�v�B)��t̠�E���~���M_0Xl�����8Ӏ�/-Z>�*�bW�⨇��0-8&n��V�0,�l�R�Q�ȓ.UB�(Y�O(��A)�Y�ȓE��y ���%H�\�*T��p��ȓ;�1���@>@v�B���Z<�ȓ�� ���S�|�b���69������F�.j��0*��(T:���P�0��"6���9���u�hM��i���t)�����Ղժ3!�4���2�*��
�H�yBB@� /�|��;K�ɪ���}�\�@!`����0~����L�A�l[�m�%s|��ȓlWb�S�A\�t�kFNݕ	����s��} �f6�[%/�	���ȓ�n�x KڢE�As7��uL���!�H���-z<~p4�ZѤd�ȓF��t��lǇ����<y:p)��2�l��U$Y�yzT���{8�H��1}(��y�f�����VY�Q�<�	 �QV�mh#gS�z�n,�w�{̓l�H��Ө�t�LH�s.ҳ �D��ȓa{�:��ǟC�H��(�65&���/o��в�ӂ�A�3E5�6ń�NaTt�T�udX9"5��H�R�<�v��<Oڮ��`��(�8���C�<�,[�
P�l��"º.�v����x�<��$�cܪ\����6%}F����L�=mK�"<�'��	�T2R�2q��7kפ��^h�@T.�>����5k���I"rq����B�ɟ��$�L��<)LԬGM���W��2Ph@�d㓌B��I��)�&_�S�O+�jS�K;wn]����;�\D*�O�زD�)§r/�����56H���pc��I�dH�P��<E���\M��;�/dw�Y�1�ʛ{*M��ө_k�l����d̂1ؕLE�b&֣<!vB=�b� 6�RU^�2�j'��Ѡ�$��(O�Op�<���Q��h�d��~3�xH>�y��3� ZE!��*o�i�FT�p4p" ��>I�O�Y�S�dl�(6�6mC�aXA)��X@@M��"��`y�hTaA&
M�ĂM���6��L�����|j7) m�N<�� c&Z0��LR}b���o�;��4g됢�@B�		��) ���O�� �͔�%������1���t`��<�	�'(�QQ�..'n,�e@LW�d��@�r��b�f���de
v>M��隍�U���7ETtL��䏱WҼp�v���,��C�$~���'�H��t("c43�2�����	Z��rZ���0.�#�qOQ>řB��06J����8� ����OL�s���ڸ���"0�.��Z
�xIF)�\J�(&B�?ᰝ�=��'E�ɳ'�0E����iCt�Y4��4!���?�'�NA�`G(B~<e�V��a�&�	�'�<\�@��'|̠$H�ٗ`Q x	�'�N\i�+�4�&�����R�� ��'��D�߻�<����{�=Z�'�X�14��.4�<YR�N0+r�A��'�h���L�.I��A���D�'�R���'k8р�G�/�8)����A[�'m��G*��R@�!��J-{�'�!�b�כg�h���ƋS�H�	�'�[ H��5�9y��	4&�|z	�'�P����#�\����
&�֥K	�'r>�J��N�:���A ���h�	�';j�@!,D&���:AoG�Z����'N���pi��4���O��U���'��h���Mf4�⤭�8bT�S�'�~䉳��1n.n��$�`�.-j�'�x�c?$��@�ӈ�,U�t(c�'t���8n�Na�#�P�EO���
�'%(�;�H8�����
b���
�'����ɱ#�cw�݌X:Q8
�'�ܵÑ`�#g�4yuC��s�q�
�'�P���<X��9�D
��<�	�'�����N�"�b���@ ���(�'S�X§0R�9(�k	 k�i��'[((�2�kn������W,����'邼�7A��@c𕰥�Q�DXָR�'�Ab�M4�L�z�8g28�
�'V��� O5' h����X,4�@�2�'�xU����5#2HJ�㌈Zj��'��i�F�Vږ�JW"2�8%P�'�@��ǃ9W��ɶ��h��|�
�'z�M�dH@�}=�x�%ُY����	�'������=����e�T��D 	�'hyk�NY�hlT�!�D�IJ���'��	��J�)� 8˲	�{�$�'�>0vL� Q�H�Bu�
�zf:p �'"�0��\���h�$pJ�Y�'������T1��;���7V�i��'����+�n����͌��y��'v$���T�����~`�E
�'9>L�P�.z�E�����BDٺ�yB��|μA�嬜�� ��,F�yb�%-2���aE֣N�;�H��yD�n4~����?9:ԫ���y�-��{��4�
m��-��y�㐡16ʁ�æ0�U�����yr�-@����z����(F��yRř�B{�r#��&L\d�V�3�yB�ޝ)A���u��-�QxsI*�y�B���ҹ� I�\�<%c�!D��y�j�8@���a���\��A`dĽ�y��T�	t��{�ЄUy���Ǥ8�y�%,O�����I��L�7��'�y�N�8�B�"U���8H� ��V"�y
� xh�g�Xi����Pc���"O
�d	5E[ e�ý!O2P��"Olٰ��Y}ŋ��L�,���"O��spI�c�(��fD��
�(�8B"O�`�����N3NECp�ō1�
,��"O�i�uO��]zJC'��"]d=�"O8�8�œ���I��C b�ʝ�!"O(5��+> I�b[�
�*�p�"O����H�-s�mT�Hs���"OD���ʟ"A@ٔ��i,�z"O�A���0���'2\�Dإ"O�M�P(S���C�W�?�>��"O��� ��c��y$�<@v� [�"OqW�5^͢����QZj!��"OJ�ȳb�?�x�BB0{E�"O
�I%���.����5X�8�"O���C.H��Z��1 ޚw��1��"O$�(%���C���)��d���
3"O�,�s& +����9U�ܖ(�y҅ҏk%�D�dNI�SSJ��0�ȱ�y"l�2	mڄ�V_d �� �y��I+��b���h@�wD��y��^	@p��ғ� ���7�y(�@�R�"Ӣ!vp@��fJ��y�$ђ'�4�c �WŤXzk�y"L�G0���)�:��i�����y�NԤ7�{�i��d����0�՝�yB��:zX�xA��Zהa�P�$�yr�܆��)q��JY{�I��m
��y�D!2�̤��N=z`C֯K��yr�Z��y鐉9[��kUEM$�ybI�[�����;4*.�E��0�y�#�hy��s׀U���`� -�y2B�83���P"k�J��$z��A��y��'	�lې���@�l�����y�lх&��S�̅�2�ڤa��y��(X��[Y�����O�m��s׆(��̘(`��q'�SX���ȓ8�԰���f���n4�8p�ȓA�
H�enk[�(�eoO�[�乆��d��P �=Rݸ�g)V  en���x�U�"��	#�q�*=b� �ȓ�D�`�(ٌk��X1NB;d�ņ�Wb��E/��?�n!B�*I5�$!��H�r�%U!�:��α�Pu�ȓ1�H괉S�v&�,��	*-JY�ȓ1-X5IF�ې�pJl��k V�<q �Cu�r�:f��+O����S�<��,I#�r'��*SP\��PP�<QVLS�B�D����Nؠ����r�<q��ߜ*&��R��
�'z\y�/g�<!��۵�4 2��n4�Bq��h�<�RUX'ܽ30i�VO��ҡ{�<����*DZ��3�&�6���C'�\�<IQ�ܕn1* hfL�cَ����r�<��ܕjXTQU�ۃx&t�jŀ^Y�<���j���*Z�(�2h^�<���-�:�:��Q=jt�RR�[�<i�FՃ%�X�tn�?YD��b�AM�<�À�9wc�j"�B�.,N�:���E�<i MP�'��t�ufK+GX쐂,�A�<�tEҡ �4$��l�}l\���G�<V�߻��]�CBN�V�%ip��@�<9D#�9M'�q��'}`��7 �z�<� H C%�W3?rF���Q�l|#f"Ot��H�4z�
�ɐ��42pf���"O>4�%�ȅk��4Qt	D*��D�"O����^��!*� �3L�%+s"O\��*��)��Q*qIQ<q"O0�Ѐ�g`�Z���YKn��S"Oz���
.cв��@�C$/�=P�"O�qBuI�<&�N�)���o��\�p"O
�F � �Db׉�&�����"Oʜ�QC�#P���V.K5b�l@��"Oĵ��EC�E���΅,1p&�"O�e�v��.s
��rPǀ,"Tj�Q5"O5�C^� ��q34��2io�չ�"O��D �/��i'���M{���@*Oƭ�-�*�&a
W�!<��k�'�8e0�(ձB� ��f��	���'�yae�[�1X��T�X�4��')"%IT�Y��;SK�C�'���q�B�0I<�bsF	1}��+�'�>�Ɇ�A'/���P �кv�R��'�&��bMe:iÚhxq�	�'o�9Ҳ+L;$)6����޷b&�%�	�'���Ä�L�:+�x���ĕ`���"�'�t���c��k���UZ�n8��'�8����B�uI�|	 iU)&�\���'B�Dcg�4%z3R��qT|��'*]�Ao��8�����h�3K��h��'�̉����YC���B��DLRE �'��`h1��7��x"A�̊C&�s�'�� y�
[+C&�������U��'��I�AeɭH���J���
�T��'����������烽�p��yz���C7:R��@��ɀ����T|���t�a#B^�PM¦�}�<I"%[%G�:5jԋ��}���jM�<��$�	>^��8�D�K�b��3��K�<��+E��� t��&pJiyB��~�<9�Ꮢ=�� ���# �|���͟N�<Q$"IH�	�J�1�D�#��@�<��(\�'��Q�"О9Ĭ�r`Fs�<9�J`�����d�ht@'Fs�<aU$P �v��s/�H� �ekf�<�K��1S��s�Ǝq��Y��Mj�<����s���r��%^>𰙇��h�<���:�&�0�	 w��q	&E�d�<�Í�fq�]�� �V�Z,�3�G�<ar���&����������!��7�yRd��d��%��5`��y�G��p�`P9V�S�<�����y2��L
)�fJF�FZ�L��Q��y�{�\�T�R�@(���%�Y��y�k�,P���bI�g	2d�-��y�$Xk]$� �܅XA���U�J��y�S��mB�+L�M:屵���y"��u���a�E�	G�����Ґ�y��ۦ
;�P��N� #K��y�Ʉ*<�f�"A/\)CV�]��y�թh]%�"|�V��ugP �yr�t���'��u��PiԷ�y�n�4x���i�
~S�ukd)@>�yr�ԗe.��oޥs��٘���yBM̭����N��8t�#6	O��y2��� C��2.t$������yr�W� ��"�dA%����@��y
� ��fi�N�N��r�<d�a�B"O��r���'���E��VN "O��#�X�Y�`�!E�?YM`"�"OR�z��]�2
T{U#92,ؐ�"O|0�aJ"\�^ )���"w��"O��; �(@�Ax�A�"��tr�"O���ȅ�"R2nYJ"O�%�@Fޔ[�x�����l�,t��"OXt�"Ƃ�F��Cw��G��w"O&��PK� A^0I�A�)^x��"O�=9�-�	���v��{	F�S�"O�T�0f��D�d��O�"^&<r�"O<��/@7�P��5�;�݃"O��G]W�����.9M��M"�"Ol���   ��     K  �    �*  �5  _A  OM  �X  2d  Bo  
{  �  ��  �  �  ��  0�  F�  ��  ��  �  [�  ��  �  ��  
�  ��    x � [ �   U& q- >4 �: YC �L XS X[ �c 	k Uq �w �} d~  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR��D�J���ӳ] �K��F/]$	����kϊB��.p2:d�a�,��������=QÓh�D}*���\�<�{ĥ��1	bq�� U&�2�A˼m2��v��$&����
rdk�A�)!��T��ΣT�8��re�q���W4O ��Z���+�'�δ+Rh��Zc�,��D ��2�S��f��zA�QW1�ɢ�݈�yB�S��n�A��M)3|��
I�v6�=E��ULD�S��"�l�B�C�tgZH�ȓp�(8�6̎��.��7�(1�І�_�%�l�-�w�K����ȓ{��4���`��n+h,�ȓd�Y9`X�^�zQ0QN�GU�ȓP~�����+���
u����5)�ذ���
T
���A�N+���F���c�H�h�>�Io:[�M�ȓ���G���,�+�T�g�0��ȓvU�M	���}0�P;�/a�f��ȓi����P�C*r���� T/jt��ȓ7��0�R�#!�X\�4�c*)�ȓ#���H��&l��:�"?r�����na��جT�0��j3R��܇�Z�ڜ�B ��w7��1��X2���ȓY���K�K<�fX�&�VL	�ȓe˜,�ӨN�Tu2tX��ĭ[NrP�ȓ�x�1m�(H��dϰ:�����4x�M*O�����,�\��>�8� 'ְ%?�8�3��t�$(�ȓy_��Q`&��fut�@d@Ϊ>�-��qXXգ�
�?Q�����'����Q�հ <A\ ��j��#o�0��Z����-�;�`��q��-/ y��g�&]6HK�Q �/I�����"D����@�,c�vh��F�<��"�g3D����l�Z3���^2CG0D���Р� 'Ava���ƴ�V�1��/D��A��� &C�5��gļTzJ�7l-D���rF�+%�(:��_�Tl��7D�`)���6 e��@����B����+D���a"ϑ"���b�C[t�$��s�*D�pڳ�& �*��e�لF]y�U�&D�d1�-q���/�rߖ �&D����oH�B����w��JAn`�.(D��:�`
q~��Kq�^>2\��!T�XCe]��H�Z�@5h���2"O�M��4l�d�
׃��8�ndñ"O�1b�b4��-	c�σc�4��"OH�y���ov�y���D�s�jU�"O0<"�*��0@p��-b�
��"O>`��7`��ܱ� ˅8:3"O��S��=ǰ�Y%-��N���"O� &��'��=y�~���L����2@"OT�	���Q'�Q0JI)RXIw"O��KD�5�F��(N;( R"O��#R��39���(ٯi�4A�"Or�PVꜴ-c��e�؞
�����'B�'}B�'��'o�'���'
&p�k��8�5i��3O�AP3�'�R�'U��'�"�'.��'E��'�Ќ
a��R�`A!�D�K�^���')��'�"�'���'�r�'���''�y3���o��@3����3��'��'�b�'�"�'�b�'�b�'Bh�CQ�S��)en���K�'A��'+R�'�B�'�b�'���'ONI�GXt�"�J%Cۓ�8���'o�')��'D��'�B�'���'aV [c�]�DJ�)�����bD�'���'�R�'���'2��'���'��$��D��ߠ��4*Ol!6�'Q"�'�B�'�B�'�R�'���'_�	��e�,y5���U������'���'�"�'*"�'�2�'r�'������ė/*��;�)��c�u���'r�'���'\�'<��'�'�3P�)-X(�q�fA�����'��'�B�'���'n��'��'Ԕ9y�HG�<�����dݷ6�bLH��'��'WR�'2�'���'�2�'�F���+��: 4��e�e�~ ���'���'$"�'[B�'�NvӮ���O��	U�wY����^�!�Ȭ��xyB�'h�)�3?�i^�ik��M-gYV���#M�+g�����"����ڦ��?��<q�zXU�C��W>�B�b�7A�����?yt`E��Mk�O��S��J?�7�7eD�G���^�,ٕ�-��ş(�'��>-�C���
�o؄p�!u��M;�A���O$L7=�28�jS�	Y�lN1fXp��r#�O��D{�ק�O���ºiE�����\#�Q�I>)�PdN x&�$m����E�=�'�? 
�(��e$(���׎��<!(O��O�@mZ�?�"c��9��]�bKB陁*$��`��X���I���I�<�O�`e���̞���Q��٩2&�,��O��K�rf@Q���?Y�b�OTx��ꖂ��#���(:�|�q�a�<Q*O~��s�,�wfP�<\��o Ԁ!R�c��ڴ�b��'��7�&�i>9��ƚ�L>j$���S�����l���I�d��!\�`oi~R5�da�Sk���P#C
5i�E���&n��ꢘ|�U��ʟ��	Пh���|��� =!nJP�VkW� t�ەIAyrA�O.���'��'V��y��;���x�`H�IW��+����_I��DX�v�x�*�$���?��SgT8��	�^u�#C`�H�IS.�����542���7�2	��f'�'!��0�ڵ��$N0KWxAx`JVU6����?I��?���|j,O�n�<vHR��I,
�<��*̫4��+0ρ�C,,��	�MC�2�>�#�iN 7M�Ŧ�+@LAzGX�5N�i@�����+F�l��<!m��u��8g ������z���������"d�4�Y�E�0�%� ��<I���?���?i���?����,߬��dJ �L{k�p�4F[�5���'���f��1�6�t�d٦�$�({%��,OE�����&O�8�3
2�䓈?���|�E+���M��O��]wx�b!N)˦�����=�F� �G�O�t�*O��n�iy�OC�'���(M)�]�2(��J�&q ���"�'�剂�M��e~	�I�$��P���O;d�&�b�̡���.6����Y}
l��m�"���|b�'f�j�q۝��,�$�^R��|ɗ�.ъ`��ML~~�}�y��'h�i�'�wH�z�(�W#E�	�h�Iրt���'��'���tR��ݴ!�H���"e���C�
KI����i��?Y���F�'�'oh��?��o�g�����Aպ'x��""<�?A��i;z��D�iC�c>}��f͆�����j稄�I�|��e ��^@:P�)�M#*O��$�Op���Ol���O˧n��ӐgF�fC�
'K�'���ĵiʂ����'�"�'��O�ҡr��2�{%,J���c��0�� Cv�'P�fi;���(�D}��;OzaׇG ��ٸ7K��I�A�P2Ov 0R���?��Ĺ<��i��i>�I�iH��x�M�QyP!�r��>�*��	��D�I���'G:6-��f�$�O���ƣw��t��)=N� CӉ4h�,+�O�qm�M+��x��
�\�x�h˞]�l�M����іͫA�����I"�u�I̟����'���$Bڭ9\���G���].����'<r�'R�'	�>�]�d�p�����?ZZ\z��U�s���I������*���OL,oO�Ӽ#SG\�B�`���8qx8Y�R�<)���?��i�x���i���=�,1C�O��ףJ@5�����^�1㐅Py��oӲ��|*��?)���?��#���d�[=��P[�-A�it\��*Or o�2Z�E��֟\��_��֟�#�ڋx��R��)'�.�@E�[/���O���j�i>=�	�?"�O��>DaG��mdQ+ԧ\82�����-?�F�E�{e���^���Z�՗'�H��W�V��4�3�K�dY��S��',R�'�B���S��c�46�F����-@"mx1�+k6�����8I�D���8ћ6�d�ty��'���ehӒ	D��.-�`�ǣ�F�[F�Y*)�7�r���ɥw�(ut�O%��H����� �!��a<{�4��DL������7O����O����O��d�O��?�r#�T����憭V/��ٟ��	���ߴ7~��O�67�>��S�*��𢁓b��,9ԏU��2�O�4m��M�'�
�`ٴ�y���n��$Z�BT�r�L�R�^�A�|�7�X&H�)�u�O:��'�r�'�r�'̜u�c��2k�\�sgϝlE�U���'Q�T��ܴZr���?����i �W���z�l��̕Cv��;6�	����O��D,��?I�g Y�VQP�	!$ �q�LТ"EX�{`���4�֦���ĀSA?	O>	`k�	2���̰,�����)�?I��?	���?�|Z+O��o#��|� W#l�j�)\���a�GmN������MӎҪ�>���nm��*3M�~�x��*�m����?q����M��O�LS����zI?I�ê�(.��82� M|�5��k���'�'���'%��'�S��4��2(МE�`�f��'ވY۴M+z���
ش�?9H~ΓM��w44ѵF��]n��w��*n}|����'+Җ|���e��EY�4Or%�F��5d��wm��0,��1O�p:S#�.�~�|�[�@���kFD�QlΉ�!��EӠY/�۟��I��8�IPyB*~ӒaBG�O����O�P���.�(0��'���xrO1�������O��d%������Đ&��#Qꩩ�(_�V��I�(�``����+K~��`�������l�GM^#St�+6bϡe��9�I������IT��yg�W	t�� �	Q84Ś�Ķ[���f�zH�5#�O�������?�;�����üT�x�ʳ���p�r��Nӛ��s�b�oڄFz^�l��<I�:���������'ϫ~"����*'����t�K�����4���D�O����O��W�)�fŊg�r$�B�!&˓Yb�*�P�'�����'�riS���5>��i�dh�
F���h�>���?�H>ͧ�?�����	j��q�pi�:�֘;��A
@�X�'v"�0����R�|2]�H������L�{�RR�܅�@��������I���@y2�~�R�:��O�)c��Ĉ/YB�@�c�&l���O��l���$���O��d�O����,Pg~4;�� ��
œ�v�Y1G�?��3O����B+�*��L���?i���a�5N�6/Bif�!�H����|����x�I퟈�IO���D���8Yk�E*ƍU1b���?��G��f�X���$\ڦ&�� &�Ns����mO
D�&����I�I����i>E���Xʦ%�'.���K�CM\萗���4���O�X�������4� �d�O�$�`�4\�@2*d�2g%�O��d�O,�u������_O������O�rH@��b�Vy�Ř�'���j�Oĥ�'HR�'�ɧ���'���au
51���(��m�e��ϝVȌ}���i�rʓ�.�:�	\�	��`��=]zPY����"��I�L�	���)�S}y�moӮ+D�-z��tCݡ8^�h�2�хp@�	��M��2�>y��#�dls�l�,O
.�h7�Ԗv��(9���?9v	��MK�O� +%�ׂ��O:�ٚ�G�
�b��b�'����'~��˟�Iڟl���(�	l�4jͦ�����*ʹ^�����̑%�r6-&*U�����T��y�ǜ4�$�˧����:�s��&�b�'Qɧ�D�'b�䊥.$�f4O|�C�I��c���m��#�2O6�JJ8�~�|U����Q
�=�ʙ�s�EX���9���������4��Xy�e�&�����O��D�O!�Sd����q�c�SJD��0�����d¦���4J�'m���1 ?:p�� J\+�>�ڟ'J� G	,���������Hh�V����ҷ2 �E��lT�KNMXBИ'tF���O,�d�On�D1�'�?q�(ю��Qc3��"� ���]�?�ÿi�6|�g�'�ңq����1*%>h (��S��U��^�u��.�M�P�il�7MS.9/�7�m�8�	q��z��O1>�3��ѿ�ֱjp�D�)C��}�Ey�O�r�'#�'���̆-�*�I�gW���a��cД@�	��M+����?��?�K~
�	8 j-[Y֨[DRsO&u��P���ڴuB��)�4������X��t($�"X"@�Zv���(�a�R���c�Kt[��D�IQyR΋�\�p v�ͶIߪ���m�s���'�'��O�剨�MCBω��?�m�>l&�P!C�V�+�D� 4�Z��?D�ib�O���'7B�'~��Ob����C�x�@h=1���0%�i��ɡ-�� �ҟ䒟��/YV��1���9#�� ��6��d�O��$�O[l�ܟ<�	}���0Lbfd�>`8h6�ņo\fLB���?Y��C��6�����'�t6�1���X��X�V���1�]� A�F|ܹ%�`�ش��F�Oa��{�i}�D�OƱQ��9�CLׁ<�}�oD�X�,(;��'�t$�<����'��'r2�iW�ٜ�T0�GUc8���'{"R����4w�v�����?�����IU2v=|�Sbn\�����¸d��	���Z���Y�4����)J�����!+�˂��|T���5�JT��h �j�3��i>�0�'l��%� AF�����U�����.]ܟ���ПH���b>��'47-ц:z�b�N�(t���˅�r٪1���x�ߴ��'��듪?��ic}Dr�����^	�� ����?�e�ܗ�M��O��!֣B<��π �Y0�@_9B�&`7�&F����R1O���?���?A���?A����I=F-p[Ч��@���t-��o��n6Y5����ן��	S�Sן������e��#�6����@?)8�U����%�?������|
��?�6I�5�M+�'W�X��$ɒ;����"Ot��j�'K�����Xi?�I>�(Ox�D�O����-HrIn���(�g�O��d�O\���<d�i�x�	��'b"�'k: �`RM�9Q�A��9���'�'��듵?	���$.4��"�al�颥n
�6����?��旮f��-�ڴ$C�I�?#4�O���u��9a!�����]+׎��2@����O����O��;�'�?����jh	Q�ʪP-�YC '�?���i2�QU�')��s�.��]�W_h���+�-�}��=9��	ʟ��	ǟ@�!��٦�uwW�9�ɐ-�h�%`��mrr!a%!�|���Oz��?���?a��?��P|�!�0��P���`�ת��",O�l� �T=�I�P�IE�s�P�rN�8+�!��-�*=�*U�߁���OV��"��ɔ�7�(1t�4h>�vfI�*��]�U�n��0�'H��D��m?)N>.O԰[K��[D��R�PMrY�L�OH���O��D�O�	�<�t�iJd�@��'l,u#b�TB������,@p���'7-(�ɗ����O����O8��X9ci�-p�/�J��� ��/{�7mc�x�	>U}�!xڟ>˓���W���X�,�e�bYx���>��?!��?y��?)���O����/�\GZ�	Wl��b}�=��P�8�ɡ�MK�*N�|��
��f�|�4��\�Rm�k��i%��3]+�'�"�����38�F���4	�4�R+K�kYR��E��+!��H%��c?�H>1(O"���OT���Oܐ��`�:�0F��$k�C�����O�˓<��o�0<r�'d�S>���L7O��YY'�Բ4�H:2�:?)�^�H����|'���CD���$�r*�!�V�bo�=D���Y����Mr.O����"�~r�|�/�$*�`eH���
޸�@/2&�2�'�B�'����T����4qsz�a�#M8����M�Nb�(�`���D��Q�?�\���I ����4��*gr���	֟�q������Γ����4�	�<q�g*6�hD�	8! kW��<A+Oz���Of�D�OD���O�˧%_�M���ʀf�x�M�/K�d@аi挤��'1��'M��yR|���#
L޸�ъˢM�b�_� h.���O��O1��(�+x�4扁o��")��m�a�F V-OA��*�"�҆�O��OJ˓�?i��sH�+ѡ�B��ʅ��<��� ��?1��?Y+O�<m��(�h�Iڟ��'lHI!E�'42��h�c��n0�?Y�P�H�	ǟ�$�����T\�ą���+��M�Մ&?3C��3r�s�4��Od���?�D�5����+H�H�pM�,,��d�OP�$�O��2ڧ�?��P�|�@���G�}��`���׊�?�]8��������4���ygo�:XRQc�v�kWL� �yR�'���'�S��i���O9���,�����	-�}"u��r��C��(	��'��i>�������џ�I���`�&IT�]���J�|�ĕ'ـ7��"bU���O��3��1Z>�b�K�O�N�ѷiӊ��P��O�xn��M1�x�Of���ON���̘V�(�Fi��6Lv���\;,Τ��O���o�9�?�0�İ<�A��bA�G�2ʚ-��F�?9��?����?ͧ��d�]�w��͟ p$0q�e!�By*fM������4�?�J>�V�d�ߴ	��&�yӸ|��� �e�B�H�#���:u.�MӚ'V���E���8��dퟲ�.�5G��|x�oR���(���'X��'1��'�2�'�����Ӭ,*(\ahN�r�0��c�O<���OjLm�<�b�#՛�|�L�4҈;j�8=��Cw�ѩa��O�Yo�-�M�'�vLߴ��$��i��5
�<6�Ph0v� "o�uP���?1�/%��<ͧ�?���?Q�7?T�K�&�;��0%ꗧ�?I��������b��Jy��'���?#=�U���6v��v��&,t2�9n��֟��IT�)� K�3z��a�����"<�m:c��
��<S��*\�l����-�ȟ��A�|���M�T��ERĽ���24L�'#��'���T�d(޴h5�	r�T�%&bh�U��7V	��K0n�`~2�p�T��*�OR�䝖
� M�b*T�ʤ����8��O��Gi�P��ӟ`�D��T���<��G�YE2@��oXi��(�1��<�-O��$�O��D�O,���O4ʧi��cmC7Y�r���OV�|��i⵳i� ��'��'���y�Jr��Q�F|z��lS.<
Y�K�m�����O �O���O��DZc��7�{����%�+*_�,��`�$x�����%g������[��,��<ͧ�?Q�gW7F�~�R�C���LR� ��?���?�����$���	Bg�e���۟���e�A��E`���q��a��s?��ܟ���E�x�D�bM
�RGFxVa�4�ŗ��)b����\nZq�'[6���ş�2T��[�tиC��6'���[�@U埴��H�����G���'K~<k�M�J�VU���O5p?*�t�'��7��]^���O0�l�g�Ӽ۳�m�tP�I_�@���*��E�<���iT:7W��! cn^Ϧ���?a�-�*~H��B�? �H�"b�7q�敊�+ �1��*���<ͧ�?���?9���?�U(�zr*�Å���۶��K��d�Ʀ�@�wy��'��O����58��@�r��i�E+�33L�
]�v��x�$���?�Ӿ���B.l��-�ǣػ8=�O� =��u3Bq�tG�OR��M>�,O�ȉ�ڻ���Q�k,:��i"�"�OZ���OJ�d�O�I�<1'�iӤ,K�7� V`�s��X���@��KC�'Z�6�;�I���D��A��4n��6���2TO��x�̙�&�ԑa��i��I3gj��¥�O�q�N�N	%��tp7M��i�� �F+��}��$�Od���O���O���+��	~J(�����F�ǧO�r �	��l����M��f��$�ͦ�&��rb+X ���������u��#Zm�֟��i>���fB�Y�u�-X>0�@ňC�./� ��ÁGf���O�O���?����?I��2Z�L�[6�m�&Am���?,O2-oڬN������h��w��\w�R��D�Ng�$X@��"���R]}B�'�|ʟ��"EŬ?�NY�Ѭ�^h��xg*.RȠ� �}�~5����&MD?!L>ID�"�����⇯+b��A���(�?9��?	���?�|(OTMlZ�U&��I�#�\Mp���8$ㆁ[Xy��y�8�hp�O���<5k&AST��i����E��{���D�O�B�Ma����K"WM]����P����KC&�Ze#B+.HԵ�7�y�`�'���'���'���'N�ӟl�<�#v�\�=XH��G"[�,#v�X�48������?!���O~�6=���c,C�W�ذ)rG��	�P4QU�O2��-��I8O��6�~���� t�T��>6�z�{�p������A��d6�Ĵ<���?Ѧ"H�r$��h@H�}F �ɰ�?���?����ݦ)��K�ԟ��	��@�N�?(�H�P$I� 6����`�T��q���� ��l�	P��uS-D07ߠ���2Q���	���s�-s��n������z���'12O��nH�s��(�Ց 땩\�r�'"�'������R�eՓxJ	��"Skd�qh��$�438XH��?���i�O�!L����F�+����f!�C������ش+����$u��F��H����}��$�ު<�Z�bB��R٩��>a��&�̕����']B�'3��'Ė�� E�i���%jH�N��P�_�\��4=�h�h��?����?��C�2=�`0��NJ��ݡ�g�C���	�M���i\�O1�Z`QA��K�&�Ԁ�	_^`��J5[jI�䜟����Y)mrəD�	Sy�/g���h�"DU�Tը��Q�0��'2�' �O��	 �M�W��?Q�>�|�����$~���L��?!q�i��O��'��6M�Φ�8ڴT�Nh�׈�u{��A@&eZ��f����Ms�O��;X�@��6�S�ߙi��I?Qn�y!����crL%�'�|����ҟd�I���	����B蜑-�Ȕ�U���X�T���G8�?���?�G�iN
�O\b�|��O���nͮO��`�j��9�E�v�9�d�O����OD�QpӾ�Id� .�+��<+� {a�h��
��)pj��~�|�_�D�I��	��<#�T�th����/X��m:'�۟���_y��v�hmh���O����O$�'?�D�� n�x:|�1M����'�>�]���%~�(�'��=\� Ţ+��XӔjDv~)�У��N�D]*�i~�O�����R��'7@���J�?�ΘV��> �� ��'���'�"���O��	�M#A@�����,K�B� �7��*��5���?�Ƹi��O9�'�<7-96�݂��
�y�ȍ�W�Y�)�ҕoڷ�M�v�Ĥ�M;�O��Z���
��O?	��Z�\} �}���s�z�H�'yB�'���'3R�'��S�J�&���S�x���o�3�~�:޴_S�p�-O��$=�	�OJ�mz����-(�Q�Ņ�i�Hlx��6�M��irPO���i�%4�6�x��`�k�;lE�!J©���в'"v����ۤ&�B�Am�Idy�ObKJ�xh�5ɂ�N�EB�L��ÃK�B�'��'(�Ʌ�M;�L�"�?a���?a�,ɼ@�D��W�"M>�� �J���'\듀?����'�Йtn��ѥ��$z9`�' H�c��M�r踋���������'��"0�P(e:����m�j49"�'�b�'�2�'��>����a?dA�����k�FA0�z8�I��MCvkW��?��h��6�4�B��u���2Hr���@��
�4O���O��Ĉ 8O�6�b�8��
'���E�O���w��"I?�8��yɸ��ӗ56�O���|���?����?���,�� Q+7�8���o��\�~� )OZ�n�&�&��IȟT��X��J���)��<��y�C�C6/X�0�[�������$�b>�qqN$���0a�%S�ju�@%�h��SQ)5?���@,,���S*����!X<Q��R�����#IG�}BV��O\���O�4���rs��j̧�y�&��f��&E�E_6MK� _��y�)v� �8��O����O��d
�C �p1i<ul�ĪG@�o�^I�i����ş��;��*0��'��T�w��p�wOܾ�R�rǜ�}����'��'O2�'���'���Q�KЄ=�IUd\�BE"�S"��,����Mˡ��\~�h�@�O�$)�HD1rƸ=��A	���#H+���O��d�O��pӐ���HI2�1� ���g�	��䁡#��~�c���~"�|W��ğ�	Ο,��'�2b"�5���|��Pu�����	}yRӴ��������H��N�0B$5
$i	�1d�h�����$XR}��'O��|ʟ,D�E9�r��r��!�f�s��B�md*�"7jlӪ��|��J���'���&�K5
D�Q�G�q#>	�֬П �Iџ����b>q�',7���X�1qVG]U7��3��x5K���\�ߴ��'����?��H�5H�m��	C}�`U�M��?��Sip ��4��d�K[ry����őY�
����wH�w-!�y2X�������� ��ٟ��O�N%���'�J��d��'���+W�~�|����O����O|��|j�{K��w��Hj��K�(�F����V�p��ȳ��n��ymZ����|Z�'��eH[��M#�'�8�HA�W�!ʺ���hՍ=&��ɝ'�~�b�K����s�|2]���)���`%[��I�O��0�@�ߟ��	��L�I]ybnӠD)��O����O��"J�6H쐖$� T�q�.�I���D����ٴA�'*��f�Q( A�PN]�,C�'��҂�̅���R3����3��czV�$�*=�'G6^�:Al��qՀ�D�OP���O�$-ڧ�?�t�69h��A��8p���zA����?���i;��7�'.�zӦ�杹h$��i,��I S�gh��9�M�°i*�6���u�p7l�@��1^*�a��Ob$�1�@�ePj҃/�h{�mC�nL}�IRy�OLR�'l��'�b�~�@�fF�\�T�5NZ�)R�	��M���,�?���?QK~��N�<�A�mL�^l�! �B�>�x^�<�ڴ;���5��i_� T(���)�F����
�����o	�[��I2�0eie�'�ڡ'�l�'�li0j��.��p�ǋ̕R�N-xG�'���'�����Y�8�ٴ7��;�'Kb9�솂GCpI�*ܥauA{�\Λ��ds}��'c��'�nl��[� )f")Ee
9)��H�4�F<O�$J!e����'?����?]�ݮKAN��1�Q�E�j�'�3TZ��	���	ҟ �	⟬��Q�'M�� �� 8� T���,��}����?�����F�M)����'#X7�#��]�V��C�)��1��� ��M&�`�4^M�f�O/\���i���O�E���`��	d��1K� ���8��E�r�O���|���?��88�SMns��C��
�����?I/O��o�A��������ID�4��:F{�H
��ae�!��C���D�r}�|��mڜ���|��'<�^d�4\0Sq� �;���	��V�m��qRS��o~B�OǺ���_+�'N�}!�ƵG�6d!�*� )@P���'a"�'���O��I�M[���RdD�He�W��D�[��1t�2���?���ii�O ��'Kf6͏�o�6H�f�B��T �@�U���d�J@n���J�l��<����سt�����'<z|���O�DZ�Lz���(/zn���'������	۟��	S�4E+e��1�4Q'S��;B�K�0��6�ӝ/�����O��6���O�ymz�}���&yVٲgN�1&�n��G�ߟP��l�i>��I��{��AǦa�|�x�qf��7"k�T����[O0@�f6�|��&�O��M>�*O���OPLde�$v袭��f� _Gu����O����O�D�<� �i���r��'�2�'Q<�Pc-�9q5δBs�	����D�Z}b�'U2�|���X��W,Bv�ɀcL��y��'v~�#���s���O����?	��O�aCf�T!z\6|*�I�;K�X�i���O�����I��P�Ix��yG���$81V�4n� b�(�?bX�	h��ݨ���O���i�?ͻOC���たTx�����6��Γ�?9���?��#޾�M��'�ReYy6\�S$�	X�S�8w�ID,$@�l� U�|r\�����	�����şh3J�2!��;`'�[���p��gyB�j�l�!G'�O6���O���4�$>kp0�2��.A�P�@�P0����'�7����5�I<ͧ���'>O� ��N�5���8����W����a��A����'��eBRR���Z�	ȟ�}�T��7���(X���� �1�:Y	T�Oh��%���6�N*?���Or�I	�{ƌ�<��
�0:��!dO�)=�PI21k�6�?��?���?9A�A��e���h���`�ӗ1PEK��2�����5�����Γ�?!���<>b�2(�������
�Z097B� ?{~��-��0����O����O���O��d�O�Ygb[)O0L[��Ԋw`�����Y�saM�3���P��	�O��dX��%��e|�|
��n>1'�0�����`jb�T���=�C_v� �џT����0�	�|�t�l��<y��r�R0Ì�W���
�^*���&�Ȩ2�X����䓔?�O��'n�%�A�p�HV*�h�ڱʤ��3�|=��0��E�3�4�Dd[A����'WR	i� �Θ�C6����?�:���'��|����b�$�����r�y>��O�R���\8��gGs�0C��),d�`���ΑɛF�����:A�$:�dԁ'�bI���\��q�A#WT�.���O����O��	�<W�i���k�K��(���fM�����s��G46�r�'�7M?��6��d�Ϧiچ��\�	�&]�fl8勆�M���i%��z�iA��]E�m2��O��'p�ao��{*u JY��Γ���O��Oh���Oj�D�|B�DN9~Ar�ш�>N]C�K�E�F �%^#��'�����'�z7=�1#�@�:/������-�\������@ߴGo���O?�5�&�i��� ��c��8q� m���E�D��!7O�B�ї�?��h$�$�<ͧ�?)7�C���q(٥)��]����?���?����$Ѧ%���r�����hP"BF���(�W>s|�`�AOF�3n�I��(��|�=Xe�FmϫB��pQD�B�P�	�\*��#m�fDm�V~B�O�����?i0��m8�\�p�Z�L��?���?���?�����Ov�R
�-6�H�3� ��໅J�O�lZ7$�tv�6�4�L�	�N�

���#'^�O�����9O��$�O��D�%7�6m3?ɗ$� "~���z��C�c#�xs$�+ M'�`�����'[�'��<��\�퉌�`���jE�+���2�[�h۴U�ZX͓�?�����<6�c�n���V8���@ᕿIa����@�	E�i>U�i#����m�~�[ �-Hv���$>w�H�G�iY�I�����C�O�Ob�&565z�F�\I�V�_�( <����?��?a��|�(O
]o;et�2mQ$̚elƯ��0GK_�=1�I��M���k�>	���?	�o*t �l	%�*,��r0@����M3�O��p3��
�(���Μ�b����?H��X�W+V���O���O&���O��� ��=#`�9%üזA��G$~�~��ܟ��I�MK���O~*g�&�O�}� �Z
"U�x��N/"6P���?���O ���O�Ia�g�f������Y`*��8z\5W�=�h����On�Ov��|���?��!D`��٢_���W� {Ȭ�
���?�,OjinZ3I��	�����?���C��I' ��s�T1Q�\2�R�H��Iן��IF�i>��+Nv(����1���� ��EMzm���rߠ�m�g~��OI�e����n��`1-��9�&(R��k�H�����?����?��S�'���֦!����D�8 ���'EO�i��f�P���b�����b}��'g�A�b�9m��ku�ц%�ʼt�'hb풇Z���3O���ļ@�^��O?�	�J��@*v�S1&.-ʆI�/��	ey��'o��'���'��S>q0���wf�`�č�� ��|p����M�s	�?)��?�H~2�&���w���cu���N�)#�E� $��8	Q�'�|�Ozr�'�}øiS��]�K�0!�t�٩i�@4���3O6!�w����~2�|\�H�I���!��B��ẵ�m�~LW��П������IOyfh�n���%�Ot�$�O�	��Ǚ�dO�[A�E	r� X<����$�O�7��I�	$��;��L���;PH��4��������E̘DpmI�!?���?���d���?������0j�t��T��<�?A��?���?���9�>���ʌ'*܈ʒJ� c������OH0o�3Pe��ߟ0sݴ���y7�ԩ.(fxx�GGt^��'坯�~�i:r6�E��	�%PѦ���?�ЪD�%�r��U[���סR%�Z̨���h�fl�M>�(O�I�O�$�O����O��P�y"α �����(C��<!�i��Q!w�'���'��O�2�ώ#Ġ��$�ܧ���a
���	�6z�0D%��S�?��S0U�P��*� }�zaƆ�+h,42F/�8K�6�bW�Y�Tl�O^mL>�,O	b ☴K{�uo��3����Ak�O|�D�O��$�O�)�<��i�ց��'��b��E<x&�q�LB�BA �'�\6�/��<��$٦��4M �fOнF[�h1�ED�p�.��y����6�i_�	�X���O'q����xa��ônH����Ӌ~y�{�<O>�D�O���O����O��?�a"׏B��C#�J�Լz�J\۟�����|�ڴot��ϧ�?��i�'BL+.�� d0i�n\�Xea$���{ݴ�"d�W�M��'��!�r:�@���R�<�]�aBP�]���QeB�ş��c�|2R��ٟ �I؟,���Y�3����&c��-/lQZ�Ɵ���|yr-g�H����O����O$�'�T�*5��;½z�@�)j��P�'Xr�
���Nu�Z$��b��wfS�}�!�բP7�A �;j��Q3@Yk~�O�V��	�V:�'8���L�{j���Ș�S�81���'���'����O��ɞ�M3��D�4x�l<U{赢%(O7�� (���?���i��OB�'��f� �/���"�׶y��T��L�S&6�RЦ9�+���'��d����?}��6@����s�b=�7Ι{��|��9O�ʓ�?!��?!��?������׀;�P��	�@��|�q����EmZ�Mw�=��۟���m��79��w��Y�#?\r$:�)_�#
#��{�"�m���S�'9	:y��4�y2`C�_��Y���U`\��&�y�J]�I�Z��I'��'��i>��I�s��G"��*4�cX ���	П���ɟȔ'@7m_%`J���O����
PT��$> ��`�����c��4!�O\nZ�M���x��!�Vy8��K�Z��8����9��$�1��Īԫv61�$�9��s6���G(G����c�Cw�8d�'�*���O����Ox�D!ڧ�?�� �1��h{0,��W�:���ɛ7�?)�i�����'~"jb�@������p�53PHQV�]���I��M���iZ�7Y�[�7m>?��̝;�i^ �6y9d/;�h%P 1��l8I>q.O��O���OZ���OD��`C�q���jc�7�2|+%��<!�i��@���'"�'��O	r���_}����C�1
��$�[�-TJ��?Q����Ş	 � �vh�"E�H}���3S����~��͖']�$���WT?�O>�+OFysR�ѾZ �|҄����}k �Od���O
���O�)�<1��i��	�'ζ�e*P)b�x�ćW�b!�'�7�,�ɫ���O���O�쩂��1E7d� '��̨�k�._�W��6�(?��nź(z��|��;"��S �#fLJ�(Sg�%|IB�̓�?���?���?�����Ox0IّCL�J����A��R&*\˝'<B�'Q�6M��Y���+�M�J>��	�~���
�/t�M�@������?���|z�ʇ�M3�O��qA�/M��))�m�oq�t��G(�����'b�'s�i>��Iʟ�����za�A
!�P�$i�<5��I��P�'KV6���{���d�O��$�|b�ǂ+6M@�ꔥw.�R⡟_~���>Q��?IH>�O�~�cG��('�\� ��SE������)v.D �Q���4�x�(����O⽋��L+h��yx �N�S�P��1��Oz�$�O��D�O�ɗ�*2����<�ջiI �C���H���*b��::uF�X�䘥�y��'hҗ|�Oo�I��[�F��!���K�R� �@��H͟�����m��<��iCε!ɖ(��9O�Hr/��"���f�Dta54O.˓�?9��?����?�����iA� ��)�3�F�x�v�蓆;��o�.��ϟX���?іO=r��yǤS0?X'�	�k�����j�*,r�'�I՟�џ ���
Ml��<yc͎��"j��د*�,$k#��<a���!V+��	[�ky�O<��ʶT��u�r�^7Cb���Em�*$2�'��'��	��M#��ѡ�?���?�U�R�+���)ԍ�5�,�ȓ��'���?)����:@A��*���#��^�J �'&lT' �8𽐉�t@ҟ��1�'��H���p���L���yٓ�'T�'���'��>���w�pw�����ȿ.�d4V��ӟ�ݴm$�'�7� �i�U:%G�v�@R���o�&� �m����ȟ����7�pMl�R~���	Bi�''��g�KC��@e�}ߌ�{J>Q-O�)�O���O|���O\��s(П^���oQ�8g���ν<	��i[�0C�'���'���X>���|��`�����.��C K�/��ѯO��D�OƒO��OT����wa��aJ�?ĺ�ړ(�8L8�9�D�s���8q�p{$�'즍%� �'����Pg[4�A����6����'r�'R����U�L�޴*](t���Z�����љSU0��N�;�:��� ����'��'P드?!��?	�	�==(I�Ao�:�04�aaG4UkƬ��4�y��'q,��V�S�?y��O��i��NՓ����@��0�
�rᘱ+�6O�$�O ���O���O��?-�a��F��1aG�E������K�h�IӟH�޴8�>}ͧ�?�@�iUW��%H�%�8s�n�}9�IQ�	����	ßT ��W⦩ϓ�?�K��8�
�X�B	�2D�`B��i�`���O ��I>)+O���O����O�y�ǌ�]��Wg��
���s��O~���<I�i��1k��'0��'H�x���Y�fH&"֒�����5u��eF��͟���^�i>����*���z��5$r��f��|�����/Y�	�r�oڒ����LI��'F�'\�xO�4�U���J<M
t�'���'n����OX�ɇ�Jd̟�7��5!/?������O	���������۴��'����?9��JnU
�'��f�G���?���J��E9�4����Ur�g�?��'����2�<QB$9���wW�Dk�'��	��t�I�0��ޟh��[��lӺQإ���H�.nz�B,'f��7m�z���O���8���O$�nz�	��O��{l�	��HJ���@Ɨ8�M�b�i��O1�6�q KvӘ�E%!`��f������<O��r���?1�-���<ͧ�?yeB���@�R�]� L;1�B��?���?i����d��h1��ß�����(KR�� e�1��
S���)AL�p��'��8�Mc�i�rO���:�VD�&�ѓh-�Q�v�����FЇVG�ܡP�6擀TM��ן��D4\TvBN&��9f'���������	��`F���'�VA�'��wP�Ac��cښ�ˤ�';6��-w>�$�O@�n�N�Ӽs��ܫG�u
��C���B���<y���?)��O6� ܴ����B�:���?����5o�Bupv�B�/w�}h��	M�IGyR�'���'Q��'y��ƿ|�ܡ�H��h�@!�����3�MCtG
�?���?AL~��	]:0u��j�HD
�b�\�	�U�T�I��'�b>����ۭ?`���W� ��Yib �sT��l����J�'ƙ��'l�'��z \�AT��e��b�4I�d�	����ğ��i>-�'Q�6��Z���� ��ɁA�C+j�w�R�[���dZަ9�?�W���	ş�ݏw�(Т�D�p��T�R�C��:7��U�'v�
 �F]�H~��;����d��}�F�qcU5�J�ϓ�?a���?����?1���O"����F�r�H�hIъ3YR@��'���'հ7�J��i�Oęn�t�I<0\0:�Ř"�p�3�)<	9��'�,�	��S�'$vml�R~Zwz\�h�ϫJ�H��B( )4�x�c�F��D-�d�<Y��)o�mё��܀��b�-�OЄoZ��M��֟t��K��@1l�r�b�����8rM�����Ox}r�'��|ʟ� h�N��K��(���p7��pLP�1�qG
c�v�����H{?9I>q�a�=@ l���
�b�8BmWx<i��i|�ʀȝ!5��`�$�-�d`�(�$����5�4��'I��?1w�M�sn����̀�l�@���4�?!�5l���ݴ����P�{���?�'c9��R=��T �?��c�'��It�� 
�I�}#��
��T	���M36���?���?��d`l��>r(U�g��K�����.SN@���Of�O1�j\��be�x�	�+EI�@�l	��E�� �0DB�'����P?YL>)/O˓LԼ��(a^�C��8����	/�MS��>�?	��?�U��?7ɖ<�D�	��9�t����'�J��?������Bc\�H%��7#�22���ABH~�o�VQ,����iR<���\b�'���c*pdk�&�Q�ntxL۬�y��Qo���;񂗦UB�h�T��Y�Rls�N-#���O��d��?�;V�p9�ǪU2�cG��PQΓ�?!���?�D��?�Ms�O�J�T�ov�)Ŋ�V ���T�Q7%RZ�%���'xџ؛�J�	�r����$�Q�6?��i�椛p�'���'���=Ѷg��uZ1��i�6�&�9
VS}��'[�|��$�B&8��xG˓#VFt컑��?kH-��i���}U Y"(���&��'{�X�4��&`jl4s�n��`�j)��UY��Gb�+>m��S��/t(�aV`D#�rCz��⟐��Oh���O��ƞ؜���(� Y@��ŝ#Dl`�j���v� ���?E'?��]''z^9`���<��iׇ:_~6��C��DQQ
�j���j���%/R�q�cB՟����Dc�4*�H�O��6�:�d�L�}�ą�7�,��E��o�p�O����O�)ˀ39Z7-6?��{��-�C�&kU�9�6H�{}|�C�����~��|]����ǟd�	����f`@�M�L�M�Y�|�¤T�d�ILy�'b�Z�"@�Ol�D�Oxʧ1�+$ωΑIw�\�*��4�'n�:��6�}��%��'$���WM���,(���E�ehr�]� ��zŌ~~�O!���|��'�\%(���+�܍�w`/,�1��'Yr�'e��OV�I+�M��`ȲE6�yJ�eW<���S��<(C���?1ұip�O*|�'G(7혙07x�ISgLz{J��Ea��i��m-�M���C�M3�ObّWG����M?�1wCkn��b�͝Y>���`�s�$�'v�'O��'^r�'B�� �V��f(֖M3�ԃp�H�[QRa���V������?������?1W��yG��9�3��j��]B������7��֦��M<�|ଞ��M��'� �I��Q�pwjp"�`����t��'lY	������|�V����H��U�c��Z&JX�3dX��J���������jy��u�>]�7��OX�D�O���k�,O.(pe � �l��)�Ɏ��d��� ش��'���[0��<}�A��P�i�����O�d[@oS�����C���?�C��O�#���*_
�ٔ-\+��"��O���O����Oآ}��"q��s/�z�6Y�1#�@���x����O��k4�'�6m&�iީk�����[g�W0$L�=�gc�p��47ꛖLiӜ��n�L�fJ����/���P[s#�g~<�6m�74 L=����4�<�D�O����Ov��8':tє ��NVy
F��3���%�6� �0���'���'��QD/�+�P�80�M�wjP}�6�>���i#�6M�j�)�O59�ʂL|��� m�ڹh�@���N�ڬ�����O��PH>�)O�M�#&�.'�bݘwO3�ڕ{f��O8���OV�$�O�<Ac�iu�H���'���FRZ���lʤO0� p�'�h6+��8���AԦa�ش��$��n{R`˗R8W�tAQO=���P��i��	<Mo`��O�q����8����-p������Y-\����O����O��d�O��� ��Hx~�d��$&�
PD	=ߚ��I��P�ɻ�M�&�|"��K�V�|2�R5	�]���9dp��዇�X�(�Ot��g��i�'>�6- ?�e)�����l�oF	+�I\������O>��N>�)O�I�O����O�����X�ti��K��<">�3�`�O��Ľ<��iB@ӂ�'���'�S6F,� �K	'T'd2�aA21�.�g��I�Mˣ�i=�O�ӂx;�9I��+o�����Vb�9��ht�&1�f!4?�'-�0�D@(��q,H��P�� $O>u�(�X0����?I���?�Ş���ߦiWNK%G\�8�풒��ܓ�քʶX��ɟT��4��'Fb�i'�f�R7C.V$�"�՞y�1ǬXf(7�Dʦu*&�ݦ1�'#R����
�?)��<�"��Zª\�o#�P��9O��?����?���?i���	�}�� ��a�	(������M�~�Tm��@_>`��ڟ��	Q�Sڟ�X����Ū��t�t賑iM&��� CU��rݴT���c3��	ݦT(7�c���#��/0�)���?�B���"m��A���R([��Dy�O�
	e�Υ�.�g���S�/���'���'��	��Mc�γ�?����?��#L�G�^�j�mĶs+��c����'.��w��֌{�ޥ$�� ��"�T#ԡ�K�$���CQ뗐9\�8V	$��;�����C��?���p�8sP"�C׈�ϟl�I���	���E�D�'�:�Ꮾ;�z���A
�(>I0�'XZ6'�8���OX}l�T�Ӽ�n�WI$���T��p��â�<y��i�6m���Uc�)�ަY�'&�1�a��?�"Y�f���p�2Uߐ�y��J>�.O�i�O$���ON�$�O����(X�/��ŚW�Bk9B�!�<a5�ir��!�'.��'��X��勯��H�@S*�T�1�k}�r��,l����Ş5���C��;J "�,ɥ+,,-���hd�p�'RX�X��K�T�T�|�^�0�능R�������72̞i��H ş`����	ß�cyR�f�Y5��O
��p�ۆ|Yp����4W�V�ۆ��OelZO��h�	��M[Ծi�7��!H����1�ɣ'a"�#�D�3��E�|�"�ͦ	�6H�@�>9���;uvɁr���F�'��lrϓ�?)���?q���?!����O���ԑY���lW��X�e�'���'��7͙�|����O�5l�b�"T���.�K���6Q^y0J>Y��Mϧ=S\���4��dp
��p�H�TA!� .�*5�6��c���?��1�D�<�'�?���?)���l.����-
0��2��.�?����\릡��o|��Iǟ��Ox"�`B�݁-���I@.FZ���x�O���'|��'ɧ��	�/ =S�Ǐ�V�в�lř�����F�J�7�>?ͧ	�:��B�	�1�$	���#3&�a���{�R��ğ��Iݟ��)�SKyr+f�n$h��ްT_�E�0-2�L���ַT*���M���>���Zщ	��UD�!ke.��6���H��?A�Κ7�M��O�@�
Q�O��]��!�%fz!YE�
��	�'�I�L����Iϟ����I]AD���ΠR�bD�w��U�p7�B=����O\�3�9O��oz޵Q�]$5�f�Qa�o��
!�T�D�IZ�)�ӛR3:1l��<Y�ϖ�L�̃�o8]~�����<�@ż:����h��\y�O�rM��NcD,h�/e���X�h�1D���'UB�'��I�M����<����?�d�;y
���/1�ؐ0�Hǚ��'���?������D����Q�l�&��J����'���ؒ�8�f����~2�'��U��]"��a�J�M�L%q	�'�bܑ��c ة�/�-��ڕ�'�|7�&JB��D�OF�l�p�ӼSlS#I�Р�[=wU�e��<���?���6� ڴ�����U�uC�?�"��;z4�	6B�w%|�I�Yy��� !�z��uc�2����{�X�D^��Nؑ�I�����s�' ��u@T�V3K���c���
	��\���	��X$�b>�CDΈ��aFU�dt�93�"la�0n�*��)_�e�'�'���;#�l��LP�tr���e,%��������{�!����ޫ9�W+�9Qb!�#'����	��M��r�>A��?ͻ�0���U��(pÉ�~Oz�"�+��Mc�O�=��JG���4��4�wU����.�#{�|�PlK2��,iu�'���'���'��'!"���Mx&ђ�'�̘��P�>�X�� ď�&���#�'	��'X6���Iw��O��� ��øvXЁ˒hʆC�$tr�lr�t�p*�Sv^�D�O��d�O�\�d#|�L��꟨�@�k�8�Ώ/�tiWi�]|h������%��)���?I�&jl�@V	U�#	be��BW�{V)67j�x���N�����S)������?��)�f�wM��
�F>'nnm�J�PjZ<x�'�66M�@�D�O��$S���i�|J���uC"Nאu�B�G�g(03LS���]��4������'��'a�S!�-x��9VǄ�9�L�$�'���'l���T�'�2S����4[i��C��ݒ'EV8�Sˎ�R�����<i���?�I>ͧ��D�O�� <.0)��͟�fL\u��K�O����H�d7�g��I.8\�Z��[@��'�(\ˀ�V7J��y��BǨ�ja��'N�	ʟh���(�I�����q�4�$! |	�`�(-�*��q�ʍ�7MMS���O<����ʧ�?!�Ӽ�v�\cH�� s@�;>EMU4�?1������O��Ol��԰fv(6mt�s#�H� �ȹCNY"�Rlg{���g�;��D+�$�<ͧ�?����ms���(Nc�x0�b���?����?I����[Ȧq�A���������*�Ä$��IZA��R�>ɉ�Wi�	՟��'R"�'_�֟p��b�G��m�5/��R�:)��4���Z�b������)�'I��,�(d�����\�c����o�0h�|I�cO �i���*�?�N�#M�;&�l@9G�D��� [�m�:|�,���J�E���(3,���)rf��/E��Hɱ^
CP��cj�)q�&,����o�u��� �.��ɲ���%Qʨ�Ї�S!8��,y��-S��3~�<���q����9���!d怨�䇳Q�*4n�8�88���<&���RB�|�YR$��_�L����)7�̊4g�SN�`Z�͛!���93 ȧ^_�����	�K#��R� mr�c���c,p�# �&]�Ā�E*b�ZQ���Ŧ��K�h[�}r�'�ɧ5����2�a�c�� ��l�e���d��771O��D�O��D�<eK�;.�h婵hՖ>RΘ��he�����x2�'JB�|"U���`(�/{�8��L!	w�K4��n��b�@��埄��Cy��
h��S�|����d�)
�i�i&Tꓥ?�������^-p�)� x���@7
4�課�ׯS�� P����ӟT��Dy�lҁ]���~=�g�K�3��]X�F����c��u��z�xy2`ә��'>tu���E]��[�l��&̫�4�?�����d��-�jT%>����?����B :]BcGS�Y���arN������0	-��L������ȯS�P�B/��{��npy"�Z�z	j6-Nh�d�'���&?)e���1[�`"��C6%��ɨ'�ئ��'2\����I'H��p��A�� �!�����fo�N��7��O
�$�O�)|�G�Lh��\54S�`�폪-���ҷi�:�ȗ�4�1O����: � %��&@ ���h��wDPm��������,���8�ē�?Y��~2�	6�,��	=b0Y��lX��'n�J�yB�'��'�p��)HD��"�X*W�`K�
b�0�D#j��'�t�����'���}��fb��j6���$0���x�@��<I��?A����L�_����J�o�=��[�>�PgL�Q��?�L>I.O> 9�͞�#�Up�K���!�����h�1O����O��D�<i����rH�i[�X��@�*_�i�0(��+�=!0��ڟL��f�Zy�����$�6���˕��HO�L��X�+����(�	��X�'qK��)�i��}@hC�r�~���_�P�6<n�\&�h�'*V���}rL�=���p%�����@B$̑�MS���?9���?��$���I�OF��q���E�v��YU�8Ã�5v�'z��''�Z����	�	�xR�l�&�.5r���Qr�&�'RCD�F���'��'=�$�'�Zc��j��50��	�%�VF�۴�?��0*a8!%w�S�'t4@�Kf��6�����Y*��-m�'?L�Iß4���\�ş0�Ir�do�7���/ �4��2Ӻ?�J�ξ�Gx����'?��Iū|-�l�rK���t�!��m����Oj�D]H$����i�O��	�Orݒ��E�(-�4)�!۝[$X-��d�T�Sǟ ���D��H�3)<P	���%���*6�ʀ�M�} �T��'�2�|Zc�\pEʶ���DH2C�C�OUe���O ���O�˓c��Ivd\�Uy�ř=~�p �& @� $��jy��'"�'���'���r�[�5�T�Ƞ*��ݺaK��4�bY���	ߟ,��ey� �*����<��Q��>?�XDPB��p|�7M�<����䓧?���5��1��'v��h��^sy�4�@�C6Q��O����O����<i%M��r�Sԟ�hQ.�)XѰ<����&�"@���Z��M;����?1�D�zd����	' O6%3�ӦE40�8��%r>6��O����<���]�S��S̟����?�-&I�0����xo*��6F�;��1$�P��� �-�Z����%�R �#E(R, n��憶�M�)O��Hc�O�=��Ο��I�?�ҭOk�3=v%���[�#�jI�6K��_S�v�'�2���O��>����q�0	�/)�|�3�i�p�Q�	����	�����?ڮO�˓mh��3��3\����
3(���x²i��<����/��ߟ|��/��G�l�u����vI��a�Ms���?9���(��Q�h�'���OѱB*@vfUp�/8�t��U�dF'Ux�O|���OB��
)Mͤ���O�.if,�Yq�>�ʴn�ԟ�s����<��������'G5X3�}��g���Yr%Ob}�b�7��'	��'�B]��'aP%v�aj��_��Ha`�Cauy�O8ʓ�?�K>���?�'��=a���!��Z�H@�W�f��bI>��?����D"aJ�'�ZY�GfN�~fJ��#�=��0�'qR�'B�	�����4�'�,D���E�yc��@���w����>���?����dϫdh��%>uqqb�8��LGG$7!4U{v-��M������4�z��?��_�~��P�b��(��p�U��+�M����?�)Ol��ӯ��S矸�s���'A�jT�k��DqcrU9uE�>�����O|�D%�9O�n~��([���h �p�7�&N$��_�,�G�C �M�ER?%���?��O�)H�iؤ ~�c�X$U� �iH��ӟ��I�ħ�����ES�����^�d�c�tӊ����I�L�I�?�ZN<ͧ.��x`&	�F4@��D-X&_��a�G�i~j�0�'��[�$?�f��q�O�q|�1��k�%!&�L鷹ib��'D���)��)�L���7��D���)LW�H����0��'|ƔP'0�ҟl��#Q��AH�Q�Qy�kדM\�m��h����ayB�~ڌb�@�{鮍�P��RE�&�G"B��(5�4g��H̓�?i.O��$�?�"9s΁69�ty���
w�]:�
�<��?a���'�����b�
}��A;n�\Dy@d�	Em	0�B��'!rP���	�E��'v�"q��n��x�"�FA�:�m���I��?��O2|'iBЦ��c�#�H�U��MP4:rJ&���Ojʓ�?9�j�,���O�T"�Xl$
���S	F4�!�ʦ�?���?A��0���'��Yv� 2`\�(y��<ID%Ђ�b�V���<A�8�B(�,�L���O���Ɩ(Óa�<n���j�
�,�n��%�x��'X�A�g�̑k�y��� r�HCݛg����i�=Nځ��i�剓!��tk�4b@��X�S���A�H�I[��P�Fu���7)�Y����k�ޟ4HI|M~n,u��� A?ͤyS����<6�Y�d�OD��O��	�<�O���T,�	�N��T��8k0$HZ�dcӸ�sd�k1O>5�ɶq@�i� ��*Z�����4f]�%�۴�?9���?A��pw�����'��d�9
�H3��;S�q�?_��F�'h�I�
�������O��d�OB(�1=b�9#���E�r�s$�ަ���*	|ց�I<ͧ�?O>�����'\v~xД�LmPD�'��e�"�'O�	��X��ǟ8�'>�(�m�}n2#U���*V��w�߲5O���On��<Y���?1`c^�	a"$�v+F�[���бK��G�����d�O����<���qF���a2��PBE�u�Y�Ug��M����?����'r 4�"��޴g��;T �T��T#���7��X'�T��Xy��'����V>��	�v�va��M�B,Y��M�ai-�MˊR�'X�ȍ�7M� I<鄬T77�a2)��_��"u+����Ο@�' ��A��+�i�O���Ƅ��e��� ק/���j��x�]��Z�c�럔$?9��]7"`��Z\杘�*�j���m@y�n߲U�6�X��'��D�/?�c�W�z+B�rTf E��Z�Hmoy��"5[�B*�	+��i(T�NӞd|b&8 ��CڴG�0hB��i�'�r�O@�O��-�����G�NQ^4��"[�sò�l�&;Z�A����`�'���y��'�Z�A��+iRLI� �
l��&e�6�D�O0�$�q5
�$��S���K1�# A��+ܮ���ʛdn�nП̗'�t�3c��~��?����?Q�$W��u"`ʅ�8����B�P�6����'\�Xs��6�4�8�D3����eY%��*�$FDҗ�v]�X� � ��x�'��'��Q���V��2�0�gh�O��XP�P�˝Y��͟��Ik�MyB�[�oe�0��eN0�a�F'�e1�T���'u�ݟ���ğЕ'lZ�[�n>-і�e"X��ᎠWw�9c��>9���?�K>1+OΡ����O�0`ǉ(y����GjPb9.�*��n}�'���'V剒3H�QK|b"jX���qT��6�r�"���w:���'��'��I�f��	^�����z]jXP�̕Q�Ù�\0��'SZ� �O_<��)�O�����[`���C��}�ǂ�=�H�HE}"�'���'����O�˓��TM&�Z {¨�v�}�%fU��M�+O��cW���Iݟ$�I�?���O�.M�CGJ!�o�i/<l9�ٟY��f�'���y�[���It�'j��P̭	��Dh"ϼ6��]nZ�By�Ȣݴ�?���?��'%��	^y��&K*8%C���-��?6�6-S���O ˓��O"�3u��y��,J��Q�働.��6M�O����O�8xօ�]}�\�h��]?���L,zJ����b��4�\ۦ���iyr�ߕ�yʟD�d�O���L�lv����bD�z�B9j�Tm��Fo�6��$�<	�����Ok�J�9�meA�R��h�0�١��If��Ɵ���ҟ��I�l�'34a�-�Iv�M��CS%�����-V&����D�Ojʓ�?y���?QU��%#,�+ �n����\�c�`�ϓ�?	���?)��?�-O�x��E�|��F� W�$�0!dR�uͦ9;�����'�\����ğ���	>�P�A'��!�E1\�"m��M[s���4�?����?����P*�fM�O�Zc�eP�U9bѐ����$��4�?�/O���Or�$D3�<}�<�LQ��E�n��S��ʋ�M���?a/O�@�f@�H�D�'�b�O�@�C\���X�"ġ]��t��a�>����?)��q������9O2�#^��ei�
��݀�@K��7M�<y2�B
=ٛ��'���'��$H�>��O�r�{F�W -KD�JVA'=~t]nΟ��I�G6����$4�ӵp�pr
��e� ��P��0�7��%fN4l������X��8����<�aY�S�EBY(/��3A`��Eʛ���/�y��''�	i�'�?��g��U@��B;I�})TՔw%�F�'@��'�(E�r��>A*O����������o%�7�
1����@�h�<���<����<�O�b�' ���R8t��%d��d��Q�F�'���a C�>Y-O2�d�<Q���$(�jTu�$�D)D�Z9"�g�v}+Ҭ�y��'z�'��'��I�"���/ƍNCXx{�֮B�d�ea���ĺ<�������Ot��O�lC��I6mF����Cf���3��+0t��O>���O����O�ʓF�~�y�:��}�gM�h9���C�����i��	ޟ�'��'y�b�(�y�	N�6:�B��lF��連`Nt6m�Oz���OR��<!B/UB ��џ�X�x� uQ�eYW�8���蔞Q�86��O�ʓ�?q���?�����<I,��nQ�P@`�ʎ19D,�Ĉ6�M3��?�)OB5°�]N�$�'��Ot ���G�w^�Q��~5�Q����>���?���lny���9O��Ӟ e~-�Q�W��Hk��]�Pt�6��<�T�G� �V�'lB�'�����>��n���ɐ.|Xt�@�Ep0��m�ԟ4��81����^��Kܧ9�v���ձ�.����K�Aa8\m��7���!޴�?����?��L���Wy2�O�����dYP�R�3�
h�6��c��d�O����O�Rh:� |�{Mݳ4�q �		���0q��i�"�'R�ߕ&֒ꓴ��O���5���t�ƍU���Ԏx��6m�<9��N\��S���'�R�'��`;Aߟ�����$�����f� ���>#�n��'��	񟐖'�Zc[Ԥ���{�-[�\�v�(��OZ��>Oh���O���O6��<I��<%�T�R�� Lq^��mt\N̓�Y�@�'�Z�D��П ��n���ɳ�d�f²E3�z�r�t� �'\R�''�P���c����TE^�>5�ȱ�J�/ ���@��"�M�)O��Ĥ<����?���`�~`̓}����9Ak������L}��'���'!�0=(V�詟R��J&n[x0��A�5����ܗ$�lZןė'�2�'\��[ �y^>7�Ғ���k��� /��#!�H�6o���'8�U�P��fI0����OJ���r�SS��=��Xc�/�"�Q[c)�[}��'`��'�Z{�'L�'Z�i9�hq�����<[����+(e��6W� P� _��M����?���J�[�֝=[2��)��l���V!?�7M�O:��ѡ'��$�O�ʓ��ONDՋ��B{�~	cBn˿j����4F�X�W�i�r�'E��O����Y<K2�`s ��e7�R�­P�`o�o$�	cy��'e��$�V�Hj�엘*0UrV�,��hoП��I某�!�V���'��O`��  �==�b�bqG�	���:�i�'�D��)�O|�D�O8�d�٪d ��/ng ���ƦA�I�K$ޑ�M<���?�M>�10�b1��)�I��I�%΂N
���'E2�k&�|B�'
��'p�I<Ay`�s�	I .�Ԙ�v%Z���!����'�2Q���	ß(���7��C�I�6��}�&.+�,�w"`���'���'��O�-�2
~>!�jR�e^�XS��ݳ&�̩�3H�>����?9O>���?�U��?I5i�;a���I%,@/鰙����d��	�@�	� �'阄��L=��ا!�f�	[8b'��21!�Y�w�ŦI��E��L�	�JUHu�I|��:*�!��D�"��*���3ܛV�'BT���r%/��'�?�'"�Ј�'���R�kB�( ��������Op���O|xR0O.�O��|��y�⍙i�x��D�X��@7��<1���$OǛF�~J��2C���q�E%:xHe��K�N
�k��rӜ�$�O�Y =OX�O|�>MX"���ڴZ���ᅔ(m77���-+�m���|��̟��S����?��oX��s�R9iuHS���S�m��t�]��h�Ix���?��)��8Y�%�̓R��a�b��Pk�f�'��'�����-��O"���xa�/��a���Z��m �L)��=A�\0'���������.��&���)��=���W>TfE��4�?�P̒�[p�'/"�'�ɧ5���K~8S��U�> 6)���D
���H1t�P���<���?����
3�&���g0F�yQ�:go��:C��m��?iO>1���?�UcQ*e�>yIS
ЂGd��$���n�B����d�O`�d�O���Zȡ;�La(�BU�hrR� d˺[v̙SZ�P�IП�&�T�	П���~��C�.ʔ��Cf@��*!�Yx�EN ����O����O �L��I�b��%�/l��$B%{Uv೔��2RT�7�?���D�O��'@r�i�֏!�E�#d�4gx��H޴�?y���䍥_9,9'>A���?�؇{0���@&��Դ�xfc��'g����a
���᠅�4�䠸"�i��I�����49��S�� ��$��k.hQa��LX�MJ$g�Cz�	Hyr�'��O�O֞X8��,hi
�$O8�l9�ݴ!�jqBR�i��'2�O�LO�I�!R�f�kT�Q�i�p���)^��'�����O$���ǜh:�L���K8r�]Ѷ�<7M�O����O���OR}�V�T�	[?qEF��L�ls���{�@1A3mЦ��Iҟ��I�&��)����?���q�f��p.X�&��2P%��X-��1��i��Z�������O���?��4R�9	aL��a4,�kb��u����'�6�ɚ'�B�'���'��s�l��j��:��4j�Z;��(qN�pQ�)��O�ʓ�?�.O����O ��>�8�C�ػ<n�c���!s 8O���?����'lA4s�<��Ȋ�܋����Ee�4"���C�iZ�I���'[��'�B��y��"�|M�W�֚8�b�{U@O�8qX��?����?�+O
��g�L���'�|mHd*�^�`�q�C�a�ȤQҠvӎ��<q��?1��7����?q��!�X��4��4r�͐�fڥgW�2�i���'��I4X���������O2����FAqC �F�N0	 �Z�:��'b�'�RF���yRP>�	b�#�ܲ9 �U�5\�a�i�ߦ��']~l�B�l�f���O
��򟘐էu'\-N��L;��S��}�C�'�M���?1����	eyB�'rq���(�YK��`h`���zr^��P�i�����Es�H���O8���Ne�'��/�`JU�ܪK`�����?t:޴td4Γ�?(O�?��	�T��i)�-
�(0��b 
P�4�$�Cݴ�?���?��狄��	fyB�'�DC6,r����^9q�blb�n	0R����'A�	*0�^�)���?i��,r6���**�P��̕0Aư���i�B��=
`�듾��O���?�1!80��b�
i�h�0gǌ�ZC�p�'� 4��'e��'b�'�B�'IBg)� ���K��	ކ����a��������Ĥ<������?��'�VX")%���vOw��t�ܴ~4���'"�'�R�?������|JQ��qv��t��n�ԓv���A��֟��I՟��?���~r�K�Qx؀a�k����'����$�OZ��Ob��O,P2�O����O���A W��kVcI �<��M�����u�I۟��'�Ƶ�N<���5u���s&iZ;�X�@զ=����H�I�$���K��T������I�?���O��'�k�l���@[��ē�?�)OF����i��j 
Z�X�b��� H4e�cj�B˓/f�ɕ�ih���?9�� ��ɞ�`4JvM�-]f�k�O'd�OQsG"$�I�?O4N����)ď��'�ƕ��i�H�p@�'���'�2�O�S�$l,e���:2�����;W�օ�6�fa�uGx����'��A��J�@C��`I�:%�����o�Z�D�O.���)�*��>a��~�� )��8��x�"����8��'��Mq�y�'�r�'� ���%J�1��G��0��sMeӠ�D�y7��>�����k��Nyʐ�)�
;E~�q�Q}b�:��'4b�'�[��iW�ȅ~�6l2wG�:�
��#�K�����O<	��?�O>���?����k!đb�HX:�4���U&��<���?����D9H���̧Q��9�
��WZP�gL�<h����?I����?A��\�'}Hm�0
�8>�ME�vi��ɫOD�$�On�D�<�G	̢��OZ"`S�eA�g��D
�,*Uf$K Kb�~��;�$�O|���O���Ձa'p�E^�G^�c��iR�'��	q|��J|2����e�#:��Z�&Mwj P�c�.��'���'������T?cg�؞(x�u`�o��UT"��� q�N˓W�h�%�i[맽?��'-���/2��"�M�������rk>7m�OR���2}�b?A8"%X"�d[��4^u��n��G$Ӧ!��ן ���?�xJ<Q��	�L=J2��L*X��	��Ai�q��iQ�!C���S�$��ЂK)�xA�O�"�MocD�M���?���yb���tV�x�'�"�O�����%s��"��S�v�ⲵi���'�����yʟt���O
���jQ�5��i�:�$��D�v d�oZ���2�LG+��D�<Q���d�OkL�v�.0&뗏<���g��':�	Ӡ���0�I����	H��'��ቇ*E.5㰘V���Ԋ��w�F�xPT꓎���O���?����?���S1��qP7hT*�JY�g�S	W�vU̓�?���?i���?/O�kE��|:F�_�T:%?��9c��0�n�}yb�'����������B`��k���>�B���d`���E��	�M���?)���?1)O
�1���r���5�b�"6�����J;<T $�M������O��d�O��X0O8�wD��{��L?B���"CK���ir�'��I�w �j��|���O���;pllm���3�4L`��X5MUD�'Q��'�R
��yB�'�ICJ���7"��$�6f�
P�bKզ��'
,�[��x����O��D��קu��"6
R]�	�({4������M[��?�%���<�M>��$�χG�H� �³l0�f�[��MkĈY)qc�V�'l�'E���>9+OH<��i60j�����0^�P���O�����f�L%� D�d������cF�)c}� 9уɒ2Д]@(:D�l��b����$�CF�>�X�� *$�OƄ�傊+ʈ�u�!���f��7Z�\ #p#��Q��i���ΡwT�C4J?�hy���l����=N��@��&��}�����N�T0��ѲZ:��� \x��5�Jif�Kd ��!5h` ��R'��p�ԸN������X
9��l˧��7f���)%kzEd�2��'���'�҅���'��i�@4��0`	�>Z:�m����Q�Q	U�mE�Q��.9j�$��h�N�'F�bH�(�4� �<����LT�
z�l���SIu�7-ժ3pACag�U>�#� �� r2�'�D��/$n��ʵE�A����I{�'@V�ӷ/�}��D05�Q+Z�x��'�����#D��G�	K�m��'�V꓾򤊆8����'#�R>]�t���:���Va��&ű&a׍H@�Iڟ��IC}�y��E�	�1�G��?�Od��i�Î�$��ɚ��۷HF�\i���v	h�� �Hy�v&7�i�����M� ����S�Er,�GyR�Һ�?�����O��!rw�P��)�hq:"(��<!	�_�zHb��jlxC�P�1�rx���-�ēJq��q��#N�d�!�ܪb��H���W���Ip�D��3&��'��-$�xS�]8F�� /7ɒl�a�,5~,A���	h}*�"b>��
4��9�@��<M�Lœ�(��[� ��HV�=��T҅�ا����O���T�� 8�0 2��.l\�Mh�dٽOU��D�OL�S�D�	),�AC��� �#YIY� B
�'���s�	Y4"�\M u.X3+��0���HO���cAX���J�s���BJ#S;�����(��D�@פ���@�����[w�r�'�h�8�oXP����A��?�Q��'� �	�	&>�d���\M8��   ��A�"x�X�$׾*�H�f �*�@�r�C�6h�92cD�9U���=W�.��L�v�
���.����	-{�ԁ��ޟ���t�'i"Z�H�vMZ��&Ee�;�4Z�":O��=��(�'%��P�]])�9`G�"��&�'^ɧ�)$�I�`�iSi��u�8� �92�tC�	�GJh�r�g��1OjRsGQ7zB�I�b�`u�#��[m4�Ȇo�+�C�	��|��	� V�N;V��^�B��6�-P����a�2�j#UqpB�	H>FU8�3��&L��HB�ɬY{��
qNZ�$��A���c�C�ɘ_����"�?U���e��9BʄC䉳^������K�ѫ��XkbtC䉝#Ę��vU�:�b\yl"!6LC�I�EOz�1����:�L�Y��a>C�I�ua�p��7G�h P!H2݅>D�`Q���J�A��K+�6@��&D��ɗ��
�&L�0��>  ر�*O�a(�M<*�v	��
���B"O���p+��2�q�D�_�m�� �"O�����O"
eniA@���xp�"O�I;�a�+y��z����$@c"O��s��ʕ$X �����d �iɡ"ON���i
7-f��:%�4J�$	�s"O�e�%.��A�b��K�`�B��"O�͋��L�,�r�	
T2%���"O��H�[�C��يQh	y�ui�"OX��8]��	6�KEp��"O��'�з?`�k7�	2[��h 
�'��U")�5�.�;s�ռ{1���'{.9CĄF�w�hA�]8�<,h�'�M����q�d� )C4L�N\K�'���l�%�j �[�n{��	�'펬�G�z��@g�d��`��'��p����=3��< ��C&Eq�y��'�(q�%(�N��X��r�����'/J�J�	<+^&!��E,R�|���'�QP�N$&Q0`0�n�45�L�h�'9@��gJ&\��d��Dۆ;��1�'��#&	��<�0D�S��:SV1��'��h����Jj��2C�,�D��'�<�[4߇���s��W$��`	�'�z��pM��+�rI��MY��>m��'����Ά�m5�S��3xԀ�'�A� ���h���"�@�'�F�2b 8W�<5�Q*����'���&F�akb0BΝ��y��'��[G!R�>�1�*�
q��I��'7,4{�G�
G��*)�#�LJ�<9
U�|hN�9��	*� ���+�|�<�U��T��������]���Sz�<�����w��P�ӥ3�-q���y�<ɣ��2�1��	��֥Rv�<Q6��4����TUNk�1x�ct�<��M'>o4Ș3%ڕb1����+@q�<	'F	�`^`	� �D��*Q�j�<��#ȏZ�F�wgA�dFDKg�<�g�I,IjY#�n >�� ǈ�W�<q���\o�� ��F,ܽ����U�<����%x�*�q��`�h�k�<iF��3k�9;B��B�`Kt �e�<����{e�x�wIL�C$����ώe�<!��ƳH8�i# 7���
��NH�<	˞�Yɰ�0���i9:�0L�G�<� �����

ufpS�ȡ	j=�!"O��{2,O*h��q����3�l|��"O:��
��Ox��!R� �v<rQ�"OҐ�B� ю�"D$��v�$�"O�h[A�ԥ*�FQ�Q�_�I
���"O��IU�@�#�f��V:-�p-
�"OH�(��{�H{0A�Ɍ���"O���"D89v�	8�j�	���R�"Op�ЅbZ6k9�+���������
Y �E��i�d8|�2�#V��%��`���y��E�
����T@L���(�5�~�憤�D�=E��oY�{��I���>Z`y����yH�$�Qiȶ>�.�Ȅ���ɒiu�}��'�4�� ��@RC��D@5x�TU���
>g{d�	bH!:*xкTI����B䉆D^������`Jv�׽&i�"?arJ��#n>��&OȊHW�`H2���5Q�+.D�����ۚ@�\�R��J� ~<��uf,D�h�C�G�T�����FhP�d7D�h��N�/�lS�c�=�J�Q�,1D�(�J��N��a1�UH��{�%<D���F�:�Bd��a?E���ps�4D�t�g��1E�:ใ,.HB�Q
��.D� J�:M�2؉5B�.v�tI8b��O؁���)�'r`}�&��*$d�yZ U�OH��a���$A�x�(�
Q��8aZ�Q�J9[�h����?I�	�/�|���*޵��O��S&e�8u�Z
���i �:EM�`�6�G�D�t)�y�M�d�kL�`q<��P@�Q��l c��77>�K��C]�V-2��N���z�M���Ѵ�6\�u��D|�=qdĆ+v�(���MWh��Ua!�_!����0�Y(K� DJ���T�7aϱT�\a�*,�2�)�Ջb6\��?,��)j��'�L�h�iҷ{5�������:�?���Q0~�P �2kF�QB�ER�jދ@%�'��d�$�Ծ��Ϙ'k��פl�"L�6��j��N��<��+�(k�3d�V����d�4'��;Ì�'aq����Z�a�$�e�[�7�H\R��'�4��a�K�wD�Ay����K:r\��b��e�P��b�7��ٸ�򄝏2b|�qb��a��I����2�NQ/,R�fK��fV�=�)�##̡QЃ�TE�ؤ�����&�;M,8�@��[6��x0���<�7l7�Tp��@ ���2�Է[�h<�E�' ��@�� n�H|����3D�?!���W�q�8��Q?5LH���l��'b�(А
 �Ϙ'�D�iV����3�K�d����F)���y���;7?T�I�@N�*�3�I*Um����	ʕ=��`Y��Dd\L|��@���|��,<O\\�a�P�M�}�cF�>�1:��C0ML,H�A�P�f�w�I�z��zA�B2ID<�j�����?TVR��ʎ�I���G{��)g�~9j���T����O?�V언�p��Ӽ��U�C!=?1�l�}0딇Cx>PT�ۦ\h�c�&D����pf��O�M�e�Ff�B�IbI+'�|����&?�����|3��� ���y"���J��u �ڼ�@(���	$bx�	}���*J�8t�N!��(OBP�+DD��B�L��h#��ˆ�'+����(� E?�Y���xA��Z&s�@BF�G�t�X��'n*�H��͚N1p< �#�
n�����$��$�er��C,\�q��ɰ'�ӉSE:L���N�\q�"O��EI�Qu]�#�-3���x%�'��]P����Z�r�0�O?QR0�K�I�X�x���Re`�*�
�V�<	���%9�XRmV�w��貣-_Qy�AI�]%޸�Þ��p<q� `�=��m
�q��E�4<a~�A��P�_��p�ƃT�`�"�HR��5�4� ����*��r�ra��R&j6��	A,�ѓ�� 24����FK)�����F!���e��a�1�X!/����U��������
\i�ᓡH�Й�NG4u3�/@sȖB��1')��`���5DΐU��,�6�tb�T��$�Ye�x����G��,1�#�+6XhB��U��x�薔�����F��}4�$(!(� H�*�e�I(<��@IAA����o�ڳ��B��'�'�qO� f�E^�
�(q�r� 1zn�%R�"O6$#Viś��e�c(��֙�<*Ð7h�qO>�3g엏S�n�q��.|��0��,/D�tiA/�V�Q��`�l�\�#.�	�,q\��'j������ +��R���Ѻ
�'ꢰ���^�J�@��S搨�(�+!��S
OV0����}(D�����{���!c
x)�ՏR��OA�9HAl�\b��J'��	�',5�t���ORV���N�
��A��i�NPE�8}r��Z�O��)���q����'�?u7�a�M�2��OD9`�a�`����A�Ih��g��hǯ�>q���X�'e���,b4p�$l��m�d�q��A�Y.>I�!�E�}済 *��k�X׌#K��%qm�#b�"��Va�=y����-sp��'
@^IhJģj�Y�4�
�p�셔��<{����m�p�'�y�)�3n�lT��#�3GӲ�1��y�1�
A��#4���R��v��x磈 4ʨ1�Bg��L�
�i�O��SB��7z�d�'%N`�1����вgL�B�lC�rE��� ��;��=뇪M@:�Ի���!�x�����hZ��Z�{�,�f��X�,J�k�&s�
��q%��Q̤X�l7�{��3J�E�ջ�U�h�R-`�cA�kĥXҍ@4?nT�W�a\8)�"O*���j�K�*��������ҽmV����[Kj�9���*\*6��<��>�.�/CȨ���� �����L)az�'���dL+er��r��I�N�z�cuj�@5� �ͱ[�9��_)v�^��]h�Z��4���`sㅏyВO.�I��Dy�����
]������ڲ֢�H~��i�1�j�Ӄ��:��J��K
?�zqZ�ψ�C�]��
(�8��E��E{�Ii5��%QY���ψB��\�aP�`�d�AT�V��hkʧN%IF�Ob�1�d]8���s�$Q:rJ��"N#V5�1m�-�f��,�11�r�� HRd{f���X�gj~�@�A��(��d� ۰
&F� 5�P�A�C^v��C� ��	SE]�p���8�m�8@[�"N0�9�D���
�n8)`u�#h���L��'+�t��6��UK�~�1A<I;P1����e� B�e�5Y�����Gc��hYD4�X�')��Q2������-��} �Iώ;�5Ä��w�"E�R�����O �k�)+�R�N4ɒIS�Fu�P���ABÏ(r~�ŊqgL'j���B�8d��� ��'`����N�49 �ղJ�zE�FA�Y����$M�1 ZL�t�W�d������).Z48��ĐWjeK��Yn��ªʧQjd .T�QЀ���'/@C��S�qT(G��'^Mn �wB`�H�K���j���8�``�R���V����݀FbF�	��C(W�a�pN�>7~,C��
U�%IhQu�ʑ)CK�,>��SQ�K�t��S��V|��ǀQ�	�hA<(Z��<i挤:(��+˭N%�(�/�~x��B+ʯJ-�Ӑ#��2��i�p���w�<��B�/x�� ��/J�9�G�1#���R����!L֘�:�C3	 � �<��b9�	���ܴV=��ZS�P%`6!�'!��.c���`��#�*��*�U`.C�	�:ˮI�T�ת��N�6t� C�I-Vi`���~�Ybť_�R�C䉗@����hۨ)��8��"ڕ7�C��'*���3�_m��)ɇ�
#�C�	�q�8��\�y��MӲ
#J*�C�	J��l� ��-M��r�!Kg�C�"���׌W긨{7��$[o�C�(0�p-�Q쏿��HfDѩ%~C�	3��|����'.����b��5�C�I�WxrM�s��=n�6�����8y�>B�	�6�h���<�R���-Z/�B䉟M�����1|(�d�h�C�ɣ1T�(�i��L L�P0�Ӷ��C�ɄQ
J!z��O@�§��?�B������+s��� ��*^*C䉢8Gh�(B�
�NB�Do"(�X��zLD-;ɇ�f�y��q%�=�ȓO���W�X/1F"�0f�\��DՇȓz-ā��U����M%I΄�ȓ�0;�͟7&ʝ�g��z���:9�H��^�=?�1���P�a<�<��9�%1�-%wrBU�ӮB<O~����N��@��鏬#la�[h���̑@�<� n��Pu֩�5���E)%
e"O��������Ԥ�)@��C0"O�,�C59|�6��e�p%��"O4B�D4Co�œ�!�E�pŃ�"O"��3Μ�V ���/�{ 4ɠB"O�Ȣ�˩Qcb�X�#	1r�0�"O����/ ]����$�ψtR �c3"O������Rڨ���K�	C(��"Ox@Y7c5rJ(Y�VN�<r$� d"O�)���$R�����X8C����"O� pɎ+e	M�eYE`IS�"Od�:wꋁ-R%z 瞣?&�Щ"O!s��*g�"d@G�¢-"�( `"OV�8�HL!�j��6K
�Q�@2�"OX�"�aP�~,f��v	U����Q�"O`���	��pF��5�2î�h�"O�� ��צIVh)E)�
{�$�S"O@��"
ؠ	SL���%D�(��ɰ"Oj�����<�u�E�X��\�s0"O�K[�9��kY=3���6!�C_����`U�q�Fia�*Xu!� � ؎h���8A�������!򤑲qȆ�Q�A��"o�.I�!��٫6~����84�`.P5Y�!��їx���0)C/��Yyƍղf�!��=4Ӳ����+5��m1�,կdS!�ď�SSi�+�J%Ae��"?!�D��+%X�mͯZ4� fY6�!�D�,p|��k�+�(vˈ�+���4�!��<.@�Fm�P����r��fm!��M�!_����/-5��]���#Xb!�� '��p�����qk1�B� `!�d�6�r�FN�;sh�]!�D�%/�`��6��C��u�&��G�!�dL�+e�T��?J�� &A�k�!������cA � |�л�ŻGT!�$�#!��B�W�Byr�&��6N!�$GJ<��֢ėI��qD���_!�$�c��%qr`�!P6�,HV#
 G!�D@�yr��� N4g|q,�;>!�D�K܆��LV�/f8�MM# !�dԵ��p��.��XL�FA\�!�D��i�ٛ�$�)W�\b�\;V�!�dϻ �� 
6�N��8ɔ̜<p�!�dj����d�>H��\8憰An!�����%�UD��2���H�#"7�!򤑕&J	�֎��.t2ܐPI�#!�� Ű���UT��)�g�^�!�d����EPQ
�HRr��s�Rb�!�ГY�ݢ�'�l= <�ׯQ/@
!�� �,7�� &kѐ+=�󮀥y�!�$ԲR϶��엇{�8�% �CB!�d1�0E����i�x����:1!�$�{M��·"�?���a��/5/!��	�fa¤X��b�X�0)!��,����cȚ5�NLJFcgIc�'����p�|��&�^��ԑ�'� ���Y�p��FT-]��s�'�D����6P\P|�oŅO�  q�'���e(4��tī��IN��
�',e���X%���*�tR6Hr�'* �I#����oЃ?�<H2�'�Ƶ*6�T�G���^q���D�6D���u�ٶwg�1���2"z�Ѹ`�3D�� r������Sg*
�o��B�"Oģp���(
�b�n�s�4�(�"Orl@C�^�K-R3�䟴jʲ��"O�5h�'���ٲ��.㎜�R"OH-1��0_�X� �w��%;�"O|h�bN�$/�IG�W�W�j0"O:�A��Φ4�n�Y��O	1¡��"O�e��W=�Z�cw��6Q���J�"O����
�+F,XP�E��A�P`0"OVX�7.�*���*�(J\��u@�"OJ� ƯG�G?��D�t�9r3�
w�<iP�K�r���K�,ph���p�<�&�Pj\�l�S��c,�l�<�Ue�7g�je���C.r�y1`�c�<�bj�e,�`���N�=���H�Ʌbh<��kY�my�$ݰX�(��G��;�y�N�p�Tm�Ï�!S�&`�����yrd�D���H���@��3U��y�#_�pԜ��A��3�XM:�)���y��U9�.�#� H�����y"�ݱn(�Ϳb�>P{����yb���0��d�F���Y掔`�G�y���'1�� tIA�U�-X+��y`�m���
ef�8G��:ŉ"�y®X$9����ǍגKy0�������y��آ���`�W�B�V@*��]��yK�d��s�!ـfRx�����yr��Cw: �P�+r� ����y�o׾k���
��P)q�ļ[�M֑�y�^5;���r�N�b�T���ʔ �y�H���Ȝ���R%e�~D����yr�����D��7^[< ���S��y2L��
�+�>cɒ���^�y���G+P\�B��6+��A����y2 \�gn�E ࣓>*i܄�3EU��y���z�!d�6 ��pK���3�y�i�$����m��d�H-9!�8�y¬�3[���E;_Ρ0R�>�yR�6x���1�^U�<������y���&J�}�U�[,a�BA� T%�y�i߷;��`�-�}�Z��ͅ�Ps�%2k_�<��X)���|N���=�bT[�h)m���k4E��=��@-���Od�а�!mE�pH�ȓ\z��س��#���Hd�F�]�n��ȓ �jp���;JҪ����n���R��驢"J#Dm\Ѫl ^���ȓ!0Ty��R&�<���� lꡇȓ� �/�Sղ��aK�!�`�<)ŌCM)�<"��Yݴ�9#k�[�<�ƢNh.MC$�^,U[�H3�Wb�<yu�]�8HpTNB+- (�Z�W[�<�M݇X���r����s�8�
�*�P�<9��H���vO�J�q�	�I�<�s�K���@�K¬|"9� �M�<���%u�s����#�U�y�J�Vք��O[�A0�`�M�-�y���!F~�)#N�*=�Qr�n�y�K9{T
�b��O/"מ�6�J��yR"��F���a`hÍ)���%ۍ�y­;��Y�AG�x,�ٛ���y���]֪p��Y1XH' )�yM�<U	�#uJ�0M~�̀7�D��y�(7+������M�P窚�y
� �)���a�N83shQ�kܖ�c"O�y	3M٨9F��2H^�����"OxȊ��.�P���ݮ_ʰq[u"O�����E;�~��6�1`Ĳ�`"O <)��πa�p��!��o���#E"O�2Ǉ�gO��v
Jm1 �c�"OHɘtJE.% j���"K�|����"Op�R f�;S
�E:bб(��<��"O�xgP�7CJYA��ӄ>���hb"Oh\A�.V0{�E��${�}�u"O~9��(d�Тv!�U\ }8�"O�p�&��bS��4JR$O�xQ)f"O���#^-5�����<A��)�"O����55�������O>� �4"O�؄��[�
�D�ӟ.�E�"OZ��a�S���Bɛ�E9F	�S"O�`�
�?��[�"�-ú9�"Oz�ɇ16��u+�!i��}��"O��@oJi���%I�+8K&"O��P�I��8�$Jt�\�H�u��"OA��a��;ndx��L�{�v���"O���S�ߴA�ɢ�B (���"O�,:��׫-0���� �bw0�h�"O����#ߤW�h���\�Sp�1�"O��X�'��,����@��(n�q9�"O��G��
,P������sg�ظ3�'Mў��L��m�u�W�f0f�h��1D���0�&2DI3(�_�\PRa.򓞨��i���GR���$x%�B"OtӁl��zp���R����"O�p�)Y0 ���9)B��`"ON�
e�In���Y��ݥ3�HT��"O\�Xq`�. lh$�(T:/$��{p"O6�9���BN,�9�撾><�}X�"O���D��([����@%N\u*"O�2�D�)*9f�Z+Ysٰ�Ґ"O�����	}(`��u��r�Z6"O���"��'f*�#��_�{�굑"O��F��f�`-�X�4rp�ط�Ii�O�����
]j��ꢇ�5�$h��Ğ$S�ƞ%/猙���	?�]��!�"�i��
$#�H h�'9n����e��| [" j���1��
v�ن�D���e"�8rI��c/�L���Z'��z��ڈ>P:�j�j 9\l؇��8e�ТO4n|�������pϘ��ȓY�˥�L��z�	9pt�T�ȓl*����
�U7p}
%�� �4ч�H�@�`��2��9
��ExHԅ�l�f Wc�cd�E׊X�����]�>�X��
:�͒��M�D0�ȓPC�ԛ�cnX��D�99��ȓ%00�VO!w8E���+�+<D��;�+�*^��SC�}R Y��	3D��PD0�����(�+x� ���+$D��6
r�1��
N�Y4�6D�ؚQ�0Ȱ����3\rQЅ@4D��̚V�|5ْc�]\���'�1D�a�
�n���k"��+����0D��z0Z�6t�U{�bب 񆕱�3D���gH6�
��Ժ �'@0D�<��썄~~�X��CV~|��WD+D�$�R�
Aɮ�R�k�J�%D�Li4�	�X�R\�'�v��h�%D�� �,�����p��걧��}]f�K�"O�嬘`E	0�GY�H?���"Oh��Q�,5�����kO/��ҧ"O�l�a�I�2�d*1kԨ-���"OL|1T�ss�X��D-f����"O�3"eİ;����d��R�Ƶ�"O���5.؈��Z䌈ie$�A�"ORi�$Oے'İ�a�D�L�ʐ8�"O(L�Ś�%o�p���K.>��cG"O�)˕��kQ^�*�L�"��r@"O�̑fe����bs�@��L3�"OTI���<[N��a�CV& �F,�"O:y�Woݔ%��c����q)V"O8��nT�}�t{��_��"O�Jч'}�ƁK��#/��x��"O�����Z;d���Ϋg�1�!"ON�$	�C=�,���ϖ�a
"O��7e��61ްA��k�B�KC"Ov��� �̥K�H΂���!4"O�<��"��4ކ5.)c��=k "O�@�H�E�L���M� 9�fD"Oz-�� ]ar9�D̀)s�Ib�"O�����L.���!�����
F"Oʁ�#�L�
��)�	֍<�xm�!"O��B��̛Y�<D���D�H� �"O2)ЗIBZ������Ŕf�$��"O\aa�Gk���-�4Xޤbt"O�<(֫�	q(�%8�-� U�-J�"On<P�f�,H�jË.##�1i"O��',޴k�Dm�C��1�$�"O�MZ !��|<�PIE#e��*5"O��(`�?z4�d12jX%Q���"O>uY0�$�%p4ϝ�-�f�Q�"O-[��_;Y�dC%[- ���c�"O p9Q�Ft�]:7��Wmbt��"O�"��pt�x�����P8�H�"O�y�@ �0rTcֈ=Ldٔ"O̴�f�	,>��6�^���@��"O.�X�^u��P���*�(ti"O�X����)5Vd�q��t��X"O�9��ar�iGaV�f�z5�a"O(y��K}@��"cR{� ��"O6�ر��?+��k���;�B�X�"O����Z�/��)"��|�2H�C"OR��͇Nv��@J�|(d�"O.pq�����\-����Xf�i	S"O����)�(�T�`%
�]�U9u"O}Q0@�Hn9��@�<�N�YS"O��B���yE�+��(F�X0"O.�+�jD)x)oC>�X`+�"O,	�B�֧z�d K�Η�f��W"Ol@�����B��0��K�	�Pq"Oఠ��\$ � �k�r��"Oe�� �<K��y�b�E�-슸�2"O�QI��B�;�h��OP�K�,"�"Oحj4!L�O�����('�ْe"O����*Ю%K�gF<�ơZ�"O�	����i.H������z�ٖ"O�ʃJ��y �h��ڇ5-���#"Oz��ժ�y�8���2$�x��"Ox�H��A�?���y��Z0Z �P�"O�t�B&+T����Z���[�"OҨ+"��p���t)��J�"O���`h��W>��8AM��r$��"O� rP����\�Z�̃Y����%"O�m{4�Q�T|����^��i�e"OV���(�B�"i"W�ħ �~��"O�MJ�g�[ZQ���^Gb��"O"�acDۭY4�Q�+��vc��JF"O��ǆω^��B5@��GI��"Oh��E�LS�-��^$ �����"Odِ�M��+�8��6#ǽ]*����"Oک��N��Z�(�"3%�8"O|�شO[r��ٹW�Еd��[�"O�R֧B'D���d��ȸ"O~lb�G8X��!b@�0�.)`�"O�`ؕN۫Z���X� �~�n,xa"O���C'L��ɣe��\���"O�Œ,
"��Q�� ,�B�
�"OrpK�AC�&*ze1��W�~�PtR�"O���R㏡���C0$�+]@��""O���,	�*�PQש0d@PB�"Oh�S*�U�,�R�K�ifzx��"Or8���O1%�(�Y��	F_|��P"O
M��M��X�X�CG��#NF��"O����U�I�(���%N\��"O̪f�Z�su*�8ÃϡonL� "O�Y�A�	9Z8T�#��S��-{1"O� �nM2jW`�"�
q�#v"O$�5�[2w�%�k����Z�"O
٠�[9�JT9�oW�J�J��"O(��W��8�d����)O�~SQ"O���"Σ>�=����#��09r"O`Ȩ�eE0\�PE�����F"O�-��+ �.¸��c��E���:"O���	C�2����l��aq��b"OT�ʓ�
�Q:M��L�	"�"O:��������C�MԾ/�2��s"O�LJ�NW-#� �r�G&���97"O 鲨��m��ܸ��?:v�$��"Oa���Ѱ[�f`8�Na�K�"Of�3g.�?�����N�L��E"O�!�,��������9h1P"O4�Q�ǯyζ�s�iԕn�j��"O�u!1nN;����ȕ�L�u�G"Ot�Pd\�^�8���':~2�ݑq"O:E�B�uӂ�c	&��إ"O*�X��\^�D �͖.e���"O�d�����_�L�@����w+n,�"Ob��5�Җ����7޸0'�=:!"O8jC$I��8�ɛ�N�~��U"O��"W�Z<X��H7%�^)��"O�|�B&�Iֽ@d'�5��`#�"O6<���ڀ�^�a�TtB`��"O�Hh��6��Q ��tiF 9�"O@�B�Ȁ+8�A��Ҽ{Z��ye"O�T�Sg�?)�6�#�#����[�"OjD:c��W���%$O͖�ڥ"OJ+���e�4,)&D�(C(4��"O�Yh"f�R�f��䘟(��"O��{�L��*V��b�ħ�R�23"O̡3!�ُB�2]0s�]Fn��u"O�PgHA6F����',F�E�u"O�e�7�q���b� C%Uj�!g"O�Pb`�I?I�t�0��7QlHI��"O�����ڷ1x�!E�BR<̻�"O��d�_�k�<m�'��/?*��c"O����P\ެX�"_�Y6B}(�"O� 6�g�qRD����+��@"Onř���Xˡ/�K�8��"O���b��e�~�A"�
�K ��7"O���?/�9b�N�P1�p��'d%����r���Z�k0}�JH��'v��Qږ&�T ;󊛭g��'>"926oR�M�z�s�ꈵ_錥��'N�q�~ �|cC�PM,����'�`x8��7G�h��HN%He��r���hO?��O2u�T�R��W��9EOQw�<�r+� 0W�����\�:�<Z�e�G�<� +�(@��A��ȊE�D� w/�A�<��c���܋C��8N��Bb�z�<�@[�J��I%��D���"�x�<QR�P=	Ԑ�^+�z��B!�uy2�'����S�L1O���if�)G��}��"O`-�� ւC�h	����|��	ZT"O��C����r�)Ң� w���a"Ot��rd��)O$8���X��Tȡ"Op�c�ܠI&����T ��Xp�'�1O�̋��P:Uz�Yo1R�d�S$"O�d�'I�2|m��M�,N�D:%�'�!��r��
��$P��,�b�0&�!�1ajxc��Ǐf�jp1�K�w<!�DM*�r����t�<��@��M�!�DM�S�u�3�J�0` ����p�!�d �2y�d�-2L�������!�$Ԗ��8jB�Ⱦ?�ၥ�@�-��d��Vvd+b��7�M�����B��>v} ��Μi�~=;v�V�B�I:I88�M�g�|ي�eE�l��C�I�p�Z����<�*���cC�S�C�	 &��u���� Q�`�SI M@�B�I8 �p!a4���)��B����)�hC�x��(�z਱�E/˒ՄȓhJ4��J&�2t�F�(RBj���U��bM�*?����#c��Є�w_ �1b��:Yߊ �&��~V*0��A�����L��\����Kך'��(�ȓ	�0��N�-<wn�*��@���ȓ-��0� �05E��ʕ�^�=��p�ȓnC��L��Y`�?s)V0�ȓ7, �VA�*p�<ȕ�4_����	Z�'�lpkDU|l��f�*^��x�'[�ق�%��;�-3$V���Z�'��v�_'ikm!/��K��Ah�'�xd٣��*R�R�r�엪B� ��
�'�&<��m�C0���%��<�
�'J�-���!��`c�R�4�������*�'3�0�� '.B�@����ρE삭�ȓ1"�}�#�G�tDXqgB6g�Y�ȓE�"剧lE�Xt����Gb,ф�*�Vx(7C011��`���SYR��ȓB%D��BkU����4��`��eDLʔ.���j9��հ,��(��
@T�� ��ac̏4&��G�'>M��
 C]ȱyP�CU�� �:D���S/�z{HXrD�7mh�X�D&D�x6��`�N� �e��[K�%��e!D�t�H��#)I)ΑZ(���*D��Pd#�7Aa0����R� r�i3T���T͂�s�4]x�EO�sN�T9�"O�Ѣf��g���c�D:j����'�1O���܈d|�!�`�ua ��"O� �<��i��@ zQ-G;[����"OֵS�Ŗa��c��Z�8�2� "O��j�@�n���8�"WO�U�"OP�����6��ձ"���� g"O�����ȴ4s�;��D�C���"OA�ᝧ/�4�P`)��3""OTPٰȈ�4"NY�g�w{D1�"O��0�Z-[U�����"�0�"O*��R�9�rݫ��̊[�ċ�"O��{�r��r��[Mt���"O$�	R��J*b�� LV�#Ր��7"O����=FFp��=1N�B`"Oԉ0 �K*`����Q�CH���1��0LOԄȳ�^,�R胶�ğczT��`"O��X�@�~��9:��3�ؔ��"On0�
˜�:�Q�I�0'��% �"OL9�#(��l�ڝ��g�fY2�"O��ī��t% `�V�5�Ա��"O���W���)�!{��ĉjaT�a�"OT��t������U)�E��$?LOxY��S|�he��gFޑ+Q�'7!����#Z��Α>��y5"[�!�d�=B
8�qҏպ|���S���<�!�d���<��&ô0>Yk ��O�!��Ŀ��]� �΍ZZ֬�1��!�D�~�4���$B���w-u�!�\�XV��P�ʹ9)R%��.BS��'2�'[�	O�'��$���J���x��P�x(����h��ə"�xy	�ͭK���т�TC�I#����ɀ,u���%G�\JrB�I�>1���t�
�&h����
@�B�	%x����L-�&`j��^'�B�ɥj	��Y�PF�Ɇ�xLC�I�]�4��c	�I�`� �X�e4t�=�-Ox�?9�$ˋ�vD����[&|:��j���U�<I�L���HX�/���%�>m�nB�ɢV|����c�m(IL��C�I)o��jl�-���D
{��C䉋A�f��2�F9��p����C���1{é��=z��q2'��W��C�I"f�i�Cg�g��ٓG�60Z�O�d�OJ���O�#|��eL6"�0�l�_� ���_f�<��ٔ8�Q�4m�Z��KP�Ni�<��&O$a�ƹhdZ�?�����bK�<�WJ�{c������}&p�b�}�<Y�g�2ev%�rAS�0����|�<�c��YH����ק1g���	�|�<)c��V�UGS�{|���@T�x���O�bH����/��(��.
3����	�'>>�&J��z�脪Sg: K�k	�'�fU��+|CjXP 	eߦ1|B�	�v����Ԯwm���q �#l�C䉒|��k�ȍl�ذ󃟒��C�+[Έ���R<v����%K_�(��/�S�Og����a�m1z`�3�#B��Xqg"O̭҂W��L��c�B{j�2q"O��y$(���=�d�^(@^2�Z�V�F{��)C�r�����-�`E���ً@�!��òb���R��Hp%F J�O���!�D�ZY>hY�hא<��B<��'$a|"�DP�
)(F.�	\BP����'�ў`�'���R B�zZj #wO	Y��l��'K�h�҉�(�����bD"N�؝#�'�h(&��b:%�Ə��E������� �s�?>�����̄����e"O,uIE#������ۉA����"Oġ�Gm�! QQ�?GId��c"O�U��>?�TY���*�"hkq�d1�	ߟ��'�PaC���O,��a�h�Dl�
�'�x|�L�$�&)��ā�zm�u��'�|aSG��S����a�1<���[*O8���O���VA�uRL���yI�?�!�DE�{�4�t�Y�;|w(Ɋ�!�䎲i}�T ���2D)r	�+/>!�� o���Ȋ�����~�!�X����CpZ�5�$��X"D�!��ob�=Q�	|���6J�!�$��qr$�A`*5�ej/A�!�Ε*	��hç��,�̡�4��V!�$ۤ|�J}�3(�:y�=B�ه^!�ĎѨ�,Vm�.�"�11�O��d-���r��fz8� g 5�H���'�ўb>�'׸�R�)
:���L��h'(
�'�\u�1+Ģ;@��OY�Z����\�,%�T�'�9C�䎛i�b��q��
P��4"Ofx�HJ���A���ഴh&"OP�1��-cd��p�],��Ђ�"O��;�%I�)>h)6jE4d��@*s"O6p�3��+�b}T/�gs��3GOz�a��N�XA���^�S���9�	=D���Wk�Kv�L�h[/ ���9��hO��I;R�k��ūn�b:1� d�C�_rn����"F�z9�EfK0^�C�I���]��m��6��M��'��R ~C�?>��eB�ѰjS��	3�'C�ɒ&dR܊3o@1Q�����C�n���O������;$����q@)3�윰k�!��cy��A�-�5�)��*]��!�d�Pt����$Uz!rA��¸R�!�dۮ[p2%dB���x�� �!�ɧ<�$u���	6X4&+@0{!��V'!E�)�A��7c4�	��J J!��5/�;�c�� %xA��O��Y6!���!QVp���<����K'!�$؞jE~�q�ʷs3 ���C�n!�Ͻ-+�\�Bc�{��`��y�!��]%@��%@>h�ڜ[���"�!�d\2:v��&�H.C+X�Va���!�$��8*�Z���9�{���h�!�ׁ�0�H2&�F���1W�!�dK!`��A�DK�uѪ�a�nO-0*!�I-Fp�W���d��q�bcǓCm!��y�.� !i׹6�,\��!P�MY!��9�YJ3��-��fG�M!��Q/_��u���
0�x���:j7!��_�[��*��1r���rml�'�b�'2������;'+ �i:�L�
I��v�|͊T	T8gu�IU*D���ȓm����X�bQl�3��ղ%�(D�P�7劏�1vؘ���w�1D��Xp��"��p*�R$~kp��/D��YS"H-xh�����E�4%c�'D��[�G�0O��M���܍%��l�R�'��G����]�ܨ���H�\Q��͙\'nB�I�%�4�C�*ܿ,ؘm�P�M f�(��0?��l�5k
�z�!�o��19� _�<�S	ֻC��tY�oB�VB�sR��Dy��'w���'ܫ(7T@#Y=f&��x��� �U8�AŹ.�����A����"O:,H�(ԅ9��!��D�	���D�'��'�r�'�ў(����/z|JI��킛G��R&f�y�<� �� v�!�.�1��(2	~�<����U��4z��M�`�֌p᠐z�<0A�)"��2`��%; �ЅLv�<��'Q Y�p�˚%I@0=�G�s�<���ۯws ѐׄ_�!�a{��l�<1�,ĳG�D�C�A�q��E� B�]�'FaxR
Z�+e���@NԲD��y���,�yR���D����f�-{~��dA���'laz�a����ڷ��1!��l�S�
��y"�S0q�;���3l�1�#W:�yRHO���B1�î/���`R��y��9�J]����~���KC)��yR��6{Ӕ�)0/�I�h�R���y��X�in��U*�9����[5�y�M�/{�K������yRR26n�'��4�B屧�Y��y�ß7N�0yP�S=p�4Ӈ��y�ÊV�H�B��D���
g����y���0��9�M��C0�ҡ���yR�V�KmP�����:4Dj�Pb#���yRB>co�u˂�R�&(�0񢡃��yf
��.I��
�FY��C�(��<��D��t�\��r'[�N�����A�!�F�
�j,�GD�E��s%��9!��/:Pxm���K�f � V�Y�!���4.��j#H�q��5���GLg!���=Ǒ���/L�ճƍN>�Pyr�L3p�V���m��Jw�$� �y���E;2����J�F��T� ��<A��d]�<႔*B�P�h�����!�W.6��q��/$�
��@G� �!�䗾t�hz��W��J1`<2�!�dF�FX�g�"h��%��Ӑw!�D�	jeQ��I��"Y�sEY�n!� ��i����X9â�}P!�Es�T���Y\�� �"+s!���Wg�鈔��S������1c!��&B~!{Q�óQ8�����<!��	w�D�c�͆�*rP�s!��`�~��`ҜC)�����x�!��)=n!ҴnG�wo�]����<<�!��q�b����Mbnʸ�``ҼJ�'5a|��ǆ{>�$�V F�B ���,�y�D���������>o��jO�-��?i��:JŉŠޡ�Z��EなDL^���'�5�4'^4��p��LI�'(��'�J|Ka�0�����Q6u$��
�'-\���E|Xx𛖀�{05z�'��XA���bI��!.r��+�'��ڵ��?�
��Ua;jh��+�'+ܘ�@LۏJ�,��ANf���	���'p�>�I�t���s���2������X;9X�C䉺
4 �Х@�!��Y5��1_LC��v~��pt2F":��¼:LB�I�\�>�u�ӸGT��Kf�V&ʓ�hOQ>A3���ҕ  
�c"ΑKA6��+�S�'l�V�z�n��L����A�,�މF{��O-p	{��C�t�]�ѥË>���#���2OH��� nnZ����;�"OB%X5��T_��(����I�r%"O�P����h������xyr"O� �(tNB�VJ<Ӂ�F$j3�=1�"O0%����LӔY�N}��q�����O���*�'~%: (�ܵ1�H�ڧ��7T��UD{��OÎ���	�%T�1aɄ���0�'_����E&zJ�i�A��]��h�'t.8j�I�\ry���5Q�^� �'� �
 ��8;�^mkЬM�Ih��Q�'�y��K,�XA�n_�4�@� �'3�M��lL L�"��p�>.'����'�J9��'�x�k�fUxlN�*-O8�=�O��	�{�씨���*X&������B�	�
D^��X�M���`��� ӸB�	4$�Q���6Y�$��3R�*�~B�I.A^�s��@�J[��B�O�X�jB�I��ʹ��OK�|���QHdB�ɩ�6Az�d�(8B9��HU7Z�C�I�~_L�G(����*w֋�n���O��6��?E�<y"L(,~Ёakׄ�e�g�<	�ˋy�j@��C]�F�|ʄ��b�<ٗ�O
wi2XZpM�����΍a�<�wоZ���z�W�l;-LEh<��k�#E�$p�� WhHA�mP-�y�h�q�@�#l�S���U,^�yR�� ẽ��'6M8� �wh׊��'�az�f�c�B��Fg;I0��1a$����<�J>E��-�;vpQ����FQ��ٖ�y�̰B%H��W$�P��������y���;�L%�ƥ�K��(!M����x҃)g5�g;}���`� �vX�O�q���u�΅�v��B<b�'�ў�G|R��DD��!B	{aĎ��xX �c	�'�N��h_�Aj���cͅn���I����D>��ӧ8����Ӟ@�Pi2Q��3"�@�ȓj�,���U[��Ń,A� �ȓ��f�#'�2$��BH1µ��IR��+ԃG5L���hAf��ȓz���#g��a锱�W��,G��%�H�	D���'��P���6.p)B.����i�
�'4T��D�!�6A�h�L�"�'�<񡣢��M<b%As�0*Xe �' �ԛ6�T1d���A�M(T.>�#�'J�L��P!"�e�d焳yk����'_naaAbډX�P]#$��7D�-A�'���q�M1||ڳ�Ք'V޵X�'��5�
S���$���iIP�'�l�S5�		B����𦑍5F0���?1a�Y(Sr��D��W�iN��y�j��TB<��A���'
7jbj�ȓx<P����(���dԽi�L��ȓ!wj�b �X�!�j\����]0Z�GbZ���|z�F�"(������̏|�X����p�<�hO
)��L`���p���/�B�<��X)B��u��jܻr�ԙa�AB����
}�Ji�fM<^�$�b�<'fч�6X��c�<_�݋v뙒o0�ȓI>��#�A!"w
8r.�la�ȓjkԠp��T"��������]����P�k��^?i"(��� %l�"��+D�`��J�+P��4L���p�&7D�d���܄;`\l��K���) 6�'D�\k��R�t <h�$'Pb�mvA&D�����ԙ(O`X5��$��!c7D�d��� ��p"�/һ3�*e*!D���Ƈ��K�q��32��Y���<I���3� �I�� 	&J%��s�ݟP.�ѫC"Op��	8�`]K�&��5}��J�"O~��� ��:�dX�%�+Lֹ�"O�Ih�+̪3��D[ě:8r���"O�kK-_ 	���u-���!"OD"
���\q����7^Q�b"O��(J��I�<�b≲A��hr"O���I*#N8@"��1�[��"O��*��� e��u��,K�Te*1"OD�c)]<	���K�\v�س"Of�C�� l�#0/^�9jr8�"O �����(�FH���Y�����"O⥐�(��z�$��Y�G�0a5"Oҍ���2HZEpvL�~�hya"O��0��d�T��d��|���!�Z�����<Ȑ���זK��4a��݅5�>��0?yv�ox"80w�N���ㅂ��<�7k�?R8`eM�g�8HHs�g�<���ޕ&�N!�Aؖp�fP�g�<�ĬJ9>�<�הG��p����k�<��h�&������րy`��j�<1�,�!H��ȋ��e��^�<)�çj�f�I���!��XZb��o�<���AO��8��FThV\��h�<9p*ԤXgj��g��2.ҡ�,e�<�Ta�,<(1� �n����Ϗj�<aǃ_5phLrD)QtӌP�Ԥe�<Ѵ��?���
3�s$\j7�]`�<��-��.���_�|��IЁw�<�6M J�E��.J7tD�Q`q�<���/i����e����)adX�<i�o�>X�DPF�
&����TU�<բ�>0,)�f�	(�F!&bWw�<�P�յMք��p�z~P�0SMAw�<�J_65�
ic�*T1x�� �w��o�<�Į	N���h�N��)�ڑ���i�	hy�X�lD�d,FP��] ���$\�=X�З�y�!S��: �C�RN�L8���4�y2�B=��
�#�>ʅi �R��y���3��$4q($��oC$�y�-�Pf1�B�-�p����y��^j̖�q�������A�y�#O�V��Xr6W�%@CQJ����?����e�4 )JgA-n���g��y��s�N4�E�l� @9��Ƃ�yb�Ѓp����@g
j�n��CD��yB� 6����s`��y�t��C!K��y"� 06��W)�q�؍����yRN�3�BkCѰ��eO<�y"B٪ H�#3Ɋ�e���P$�]�y���>ltM�-V���s�ߢ�y�O̢O���P�S��ϡ�yK�i��q�F�\56}���S��.�y��d �(�R$)St�R�R�y��T"�x������\��y�޻0��1�6�Q�Npa j'�yR`	i��ȁ,%b8i��_��y��0�v�H`lV� ��sCG���=y�y��Z%�X��'k[�qQBtS�d_��y©$E�J�sa���A�&��y2ć�;�h�.�|(zY0�Cѧ�yb	S�*eʭsw��y�T�a��
�yb�пb��YO��oTrd�a���y��܎N�b�h���=f%���a�Ӳ��'!az
� �(Qq��5���WE��R���'`1OQ�q�֏z|�`��IQ�����"O<��U,�G���q#/�F��l�"OP�g6w1ܴЎ��|� j�"O�	;��I8x��xe�G9f���"O0I��$E�i�����G��ʟTF���ܫj����@f.9FL@��ˈ�y"���U�Bꞣ����uc��y�"�zk
�R�-�v�� ��y��= %p0Q�CA�iX��S�6�y�
6 xb�]	Z�A�R���y�dJ�"���q��V�f�I3�Ρ�y U�|��1�D��#��-[��K,��O�#~*�c���P�3� ������W�<�dO ]�\�ׁ� w(�A�FQx�|�'��Yk᠂3/ǖ(y̆2/.�B�',p�eD�U��c�&Dv{�@��'��0�2Ù"E(<=A�Àp�*��
�'C"P;�ҥa�ک9�
��B�	�'�8d�PC�Gv�z�f��G��A��'��u3���M-:(r�a
:+88�'�^e3ǭ�/)52�pgIZ2g%�
�'|��b���$	|�	��7m�B��
�'�p������Q)iֆrH���	�'6H��p*C	7�(p[�A�:d�d]�	�'J���F�P�,���!�I�T%�i�'�T��/�� �b�ү9z b��O�<��3�Z�3(�b ���"O�
�c܊X1�Q$G �aP"O(Qb`�/s�&8�E��[5�U["Ox����^%�0�cg��Ib�"O����bġvmvx�lD �b{"O� �SF��$����P	�v0ZH&"OTA���(/��m��C�B{F�1�"O���f)B6��dj�,�8n(�@�"O| H�E�p
�c�+^�H ��1�"O� s�f��a,b�B�,.A�<��"O�%I�)��%j��@�%�2$@�"O",�`�O��x�̉>&ՊQ��"O�xч��H�>�k]�#�n�3�"O � �%¯ex!��ĚX��9R�[��D{��ID#���Ȁ��l2T+�X�!�DW4��C&�./��w*?.�!��L$Z4j��Z�İ
I�G�!�D'y��q�d,GzD1�VH���!���t%��T]���R!�#b�!�D�v���a��J\qqO��v�!򤓋;�Sb"�\�䐨`��!��۫%Q�-�s��r�>��M-�!�DA�8�V�I�vnQ��Ã!��
c�p�@F�qY�%Ⱜѻ`�!�D��'Q�����c3����BVQh�C�ɺgE�`��
)X���F� 	tB�	�GZ*�� *��<n^E!צ��'�B�!A	�4���~�k��
5K�C�I.24-J�A��Z��x(��'D�8S�XctҡI���جc� D��4)���NM�5�VF��4��2D�P��i��Pq��΀�OJ�W w!�ãFB�@�2�"8�:�i�@V&J!�B,!U��
�"F�\��a����S�!�L6����Y��RI�`��!�d��B�*��2h�w�\فO��7�!�Dd�0ؑ�������o�3�!�� ��!.��(�8�G�}4��E"O��1���G"�P��D��Kq"O�a��C	!�.����&a9���v"ON���/e�t\��[�N��"O�u�䌓+�h��a�I=��c�"O2�i �
�d~�#Da��
�Lm	W"O��)�+��0�y��I�j
г��'�ў"~ҥ��A2����F�*	�A�����yR�M1-���2b���N;Q����y��� >leSWB��K��d�alP�y���-i�$����,K��!B��yR'�Yb�{�>0�I�)A�y�K��Z�:`�2B�8W;�IY�%�yB,�?_`"Ԡ���|;d�A���y�����6�2
Q�|h�)�)�y�	�
��U�E�6����W8�y�R45<�j�_(Xf|#a���yG�T���b��L y��M�ej
�yR@
3Nҝ�רW� Фux��	2�hOn���O�܄� w%���t�X�-�,�[%��2LO|=#�n�� S��Q�.A�k�\��"O�Mٴ���S?��)#^9x\�S"O`�Z��
bb|0�D֩~��P"O��	�;xf�Tz��Rf���h�"OV	{�#I TB&5�U	�.�7"O� �pፙ?�J��� � d�4"OĈ�RJ°�;���<�����"OFu��R?���fhva\ 2�"O�R��ˑm2��8���9`L�r"O,y"���X�q+T��<o58z�"O� L�ǌe��g�!B��)3"O���UBێ�^��"�Ȟ)@�
�"O�wݨ^
6؛�)�A���8��'���C�i>y���@�a�TXCᑿ>yR�'N��y� �b��p��GnS 5�v���y��U���]��.��l�&�Av(Z�yҥ#1?x�`2	&p��:FhJ��y���	�N}���G Y��bR��y��|���1�ou$r(�y�d��?�F�9R��z�d��ܣ��$:�S�On�K��;��-�g���K�M��'�<A�E<\���"�W�\���'UNe0)�'y�!�2B�'^x�b	�'bB9���B�v/>E��H��X�\H#�'Rz���hH0pn|a�!���Ȩ�'t��S�\'�q:D-�#"���
�'Θ4S4	#}r�y���;F�����hO?)R�$�B�CB"U&A�K��B�<�t)�[�b���^'k����X|y2�)�'�nu�cmH'8ߞ�a4�F�T�V4��C���k��58P`�I�S�,�P�ȓPB�DM&y���7�B�Ĕ��Bah-R5�Y�ArJɊsM�����ȓx�5����#p쬠�D�)�j���^)]�D��
$� ��4,̤Q֎=�ȓYK��I)�N~��/
;2�8��ȓ0%v��e�R�?���ㄟ+�P]��bF�qW傭vݴ!�7č?$&%��A{4\q��ڻO�Rp)�g�i�����&>|��G C��(�,�W|�a�ȓ%䵱Q=	
�(DoAC����,�\S�OtL�i��Ė����E���Â@�=~�Ad&Ȇk"X}&� F{��t鉑65�)KVi�S�aAEH�4Bh`����?)�Ʃ�?9��?a��z��y� ���c"�[����aΖ4A����"O0(�ee��BE�$ K.D?P�2"O�Y���όD8��(C��m͚8�w"O�8��$�s�Z���ٻ��`Rb"O~-2�(�9�yDC� @w� "O�;�o̗���jC@�nfV�b��'fў�|B�'Em���獜�$�ԮE7�d��۟L����->�m�I^~*���0�~��tH��!N<1�#���̙�ȓd:p�d���x��l�sx(���̚��T�QD!�� �wԎ}��:�¡:�FI�.�q$�� o=�<�ȓIٮ��	������ȓ�|���X�B?�d؆�HhĦ���_y"�|�����`E2�΅V�h�)�IEojC�I5��Jb/<;�CC�NP��C�ɫR�p�!%��!M�<��o`�~C�=���1�a�d��8�q�ZA$C�ɷ&�d�Hq��c��qCG�4<� C�I�I�Wj~$�`�զ�),�C�I�+�ƌ;a�
Ib<H��;Tm�C��o沠 ��!��[tc��2rXC�6󰐳v�Փs���颊�&�|C�I�'�@x�B��5��9���Z�d�B�I�v��D���h.ɣ%�6VoxB�I�*"D1��K�6�$I�P&�)AjhB�	�L�(����ò`����2�3~=tC�I��T�囅P����a��0~~B��j3���^yƤZ���$���	�'QR��&d�"�X�q,��2YD=y�'-�F�W%0���D(�}��:�'��J�
�1��QtKތ]>�R�'}�ะ�\�m�^a�3�K:�(	�'`<,y��I5xC(��"OH-r:X���'Y�M벥и�j�$�ҨV�NI0�'p6�(��PKd PC& H�z	�'�� I(Q����kw)? l@+�'>�Tac��*|P|��3)�5DX0���'�T�2�hުb|�&��H�>1��'f$��ӎU�%B"T�F���BF��'x}��ʷS��|k]�;I\��'g"1�G-�:\���O H
�'����E��?Va��S=,�L��	�'v6DIS���
�� ����(zc	�'||d�2�նh��k�L͏!����	�'�>�pk�K����Hgc��
�'����6�J�j�r�A�!�3�T	
�'�ıa3F�9�:9ZS:3~4[�'��r���|�bZ��	�|��'��2!��J��B�Ë�{s� ��'^d�H��ě0�hܪ���y��!��'���aD���,U���j�.} �'SX\ad&P4&�3��F�eن`�
�'�B(Ѵ��� ����7iA[N m�
�'���1a���E�>a�g��" dLe�
�'$ą�/��S�B�"7�pL��yr�ґe1dCC�.r�Х$A��y�L\�e!
�	\88���E�ϛ�y�aY��(U�Wa�:Aq0��@Ŕ�y�,�X�P�����8�x5	ѪK	�y���Q( ��Uj
���I����y��S[�2b�&`�T�4	
��y�%*y��s"Z�E�N�D%@��y҉ �����Q?=��Q"5����y�CN:n|	�eĭ!�P$Y��2�y
� &����Wj
����D�VQ	�"O��*�ˆhU^����	uO�<��"O�Y��(� `�U�h��04����"O��j$愗q�`9��V�(2�1�"O����/�0{Q�<��!`�����"O�S�/�%�Q	���l��"Ox�`�I�����JPs{�ݓ&"O6}c�oE�rDxr�߾}�&��"O�4��*�{��e�S(;�jP5"O�d� .�@�Bi选�.y�|��"O%��Ts��=���6Yv���"OrAEA�P�m�V�@�9rr�T"OjQxfLލ� �%�N�sbD� �"O>��	�8��H�������d"O���w�B�Č�D`��.ы"OR} �ڽV� ��O8-V�K�"O��T�<;Բ���dG�"O؈�cI^CZByJP$��b�@*#"O��a�ŋ<Vjz��Py|$pG"OR��u X�8}�Y�Ո�b����"O i��)�����IAF�R�j�"O>-�$��?6����Ɂ�g�BУ�"O��4� ?W�a�.w}lY
"O()�'ՎW��۶L�Rcp�е"OFmr�@F.ST���e�%U�|��"O���(W锨Ie��R�N��"O䌚�o^#��(*�㚜z�L9!"OD��D�P�V��%J�MR/�ޙ3"Ov��f�Ƽ4,��3��I���"O���SK�,F�!����g�
�YU"O���؋8��\A����5WrM#�"Oj���P;i HPJ7 .̥�6"O�y;��<e^���"��QT� �"OZ�8���W��\)ЎN,xP"O��rbo6wL�x���ҩ�0�Q�"O�tbV��^�f�Pc���f�J�XS"O
}3sNG�j������\���c�"O�ڱ�N	&i�4��U�{ҁʢ"O�����7N�v1�\�US�x�"Ox]P��H!7����:<�#�"O`Y�R�S�isz��υ���2�"OrdK`P2k�(8���q���r�"O@�+�hͳT�ik�.N����"O�A�pjԁc��k1̘�|x0���"O8-��
�p�0�j)0`�4r"O2mxRc�:#��QهG�+?a+�"O���K&\�8ڷՁ_#6�0B"O��6
�pP�E�L��Ho"O������MtVM����}��	�"O`���D�$��EF	�.p�@�"O&�h=ˈ�b%`G�
jH4%"O�� ��9\��If�Q1��P"O,4K�j�$�x|ӆ�,qE2hi�"Oj�0�����h}�"FS9���e"O.����ħO�B�����/}zr�"Ot�ȧ�F,^G���FA�-�e"O,ܑVI��F���zL�	�  AA"O�i��bT-8�J�ӡ�'�d�t"OV�+Ю�wZJ%P�i��M&�Hp"O���F����TbU.h��%"OFTb$</���a�F8R�
���"Of��Q1�Ȫ��3K��ҧ"O�	a��ф6Q�i�5)�8���"O^�BuC2'5llfW1H��s"O� Ԡ���ښE����N�0-&�"OTШ��#ZP�UB�ͪ 1�w"O(�{���t���'K�"�5;r"O̡��bG�d2�A
�9J��,:"O��z��0
����aJ�6&讌R�"O:��ӇE,ۣ"��p��\��"O��[�$l5FTPtc�g�¸;�"O(� ��h�Upb�[cz�j�"O,�¦�G�v�fx��YFDX "O�9b��\* X�F���T�H�"O�Diu�B�s �!�"�f��r"O�eH2l�*oY0]���QkP�j�"Of���PV�� �-vSX{t"O�%j�JI�Y.D��b_m6p9�d"O��BB�2[q�}�!��sDP!"O
�#NO���@Ѱ��9"���"O���m��3i0���E�� ,��"O���
�d��M��%W
�h�aD"ON(�RNV	H�ޙ�v�7�8�"Op0!��39�]P�D�*;�	XQ"Oll��ДvAf��A�G��Y�"O��e- /K�蚀���u�d�%"O�-�W!�z#�d�p�g!��\�z��m�2���l��&�!�D�p�j�C3K�-8�ޕ"!C�4�!���HN����`�;N�ީ��o2u!��̓7:ъ4	���
����A�*�!�$�f�ص@C� �phj�(�n�!��L6�J4��:&�]��]o�!�D��-1���2`�y���9E˿xt!�ą�QB��S�����`Q� *�!��Y#r��i��A
2�����ϔl!�$��D	Z��s.џ|�&�S�d��Bf!�ǭ\bb ����'t$���X$i�!��#sXm��)M�$"��d�� &!�V�]=�ēV�M�?"����
!�X-B��{E"͞���4	T�!��U�`�J�fű]8l�i�)�!��[Ha�@�T:b�Z����l�!���,\�p �U=1zX��B�;!��%��9į�Y@�c�C�;,!�M97Z�(8��4  �6��=%!��ώsed�*e�́{�@�QA`��J�!�$Y	q�� �9����G�ӥj!�ĝ�&�Z9�� ?Z�$�s�mO�!�d�� T�PiҧI�|��U��d�!�	�#lz$"5$�W||{g��6�!��Ds�D�3յ{X�h𗂄0$�!���.#>��"��BPG8��0�U3�!�$	�U�����(,4� ��\�m�!�Ւ}��Q�I�7l&̈�7�
6/!���)LBUǭX�/-�x�GG�c0!�DH��p�a��˛���V��f~!��׃�>ԣ�nD>@��vN!��G,C6�(�'K9O��D�P	!��D&RE����&�p�Y��T�i!�d�|A��5fI�1��ɐf��d�!���k}���b�/W��}�Ԏ�'=��Dy��'�������+5�mȱȕ[�ޱX	�'(��2O}��3V�_�S�4<3	�'��X�RS)B*E(1(Ԡ d�Y{�'aXp �Mܬ�a��A/0N9�
�'J�MD�X>_C�T�H4߶ Q�'00��f��0/�d���R���#���>ʓ��� `��B��)^�̴`���e4(�P�"Oڡ��ҁ[��l��²��X�pGyBj&�')K� q'Z�S��ŌLcH���(���jR)�sT��9"�A�4��4�ȓ�0qi�#�`S��[��*T�ȓ_�����DRTFX��{��pD{��'Tt�8Wl�6�X[p`F/�4��'�݁Ҍ�}��������?��*�QS�B��S͚�끠շ)st��'�ў"|*R��$���I�2@� �'��t�<�hʧb�H���?H�4[��px�Ex��� ���eϕ'e�E(e�x�#A
E^�A+�N�G�J�b�;�C䉎׊|���S�:S�k$ɖAS�#=Y��T?]Q�д=�vq��+^�/��Z@;D�x`��G�U�nآ���4.Q���E-c�b���S�L<q��!��h��,�>�li�,ȓ\L���	B}�IRrd��e�K���<�!
�3�yH��L�:���.�v}���\���O��~�Պ��A�d!�&�ܺL4�5��J�\�<1�
W�� �J��uB�D�2�U}��|B�*�g}"��,���z���j���i�>�yc�%xpI�F�6.X�D�'�M�	�'(���v��+�<oܭ|����"O&�2ǂѰg��bP�21{�I)�"O���v䓰i/\0dV2�,�h��I~�Ie��x�-�4���J�H��V���>XRC�	>;�� �d�A�'�0�	s��h��� 3m˄[ �� �'��0S�'Q��:A
��HҎ��RQ`}P�`�p�����>���9����#Lq����g�q�{�^�L�Po��9tH��P� B�΀�sY
=��I}�'�"����޷j�:53g��G�����>�#}�!�K&xpj�:��$4��0�JY��B8����eH8+A Ɇ�8�ژ�E��,��4����O=���U���0�M��a��@K���6�!�Q�r22͒ �ޅ4�Z�b��E��p�Ն�ɛNf����e����ِ�+7�C�	2poH���9q��uS҈3Z�yE{��9O�9����7:&`�n"c!����l7D��ڶE�b�:�
Q��XLn�lt�@���2Y5��9gG� |��y�ȅ6�
���<�� I����RŔ-I��H���ě��B�I,_뒰X��Y\��4�fg�&p~�B��g�i�/��l���q@e$2B�I�F�qC�/1�|��%Ԑ]�b�d��P�'��:�F�9���D�v�2@"�4Z��	W�'�iD�4�	IS��AeQ8E0��,���y��'Aܖ=��@��2eg������Bܓ���m��:}��q ��2s�igѩl\��0?����r�E�#A[�2c B��)��O|�[ v��&c]��@�υ�Y����I'��d�>Y��@�@����%Y��u��o[S�'���=�'C����H�*mL9i��!,:x�=������F��w�,	 � &
��Uoݞo\�0��-�q3,��L�c��0� Ȑ�y�?��9��V�<w>I��*t@�Xu ğ]�C��4R�� -��f����wǆ7��n��hO���D3��p!�;_�x���, �V���He����CCc��^!94�%:p1�>�����W��\�+r� G[�4!�K�1��'��3�)��U;�E�`ɃV-t�I��	j�!�$�.9�v9kC�H8	%f�bUo٨m��O�D2�`�IX5��J߂?�q�M�?)��B�)� Υ�&��+��94I�@��Q��"O@�Fa]�s�X���R.��$��"OF����KȾ�+�&�"u��tӂ�'����;#�.%�|Iۦˆ�ՀǦ!D�P�c�N�j�aaP�fF����G�>a���S3|.��*�/�$Q�0I�[6�"?)���PcR�mЀb�\� ��k\H�O���D�k���h%�9zl}���C!�D�;�V�[cFm䎑y��)!�D�i��@�˅>�x���N,xQ�`���/~B���v�ĉOIjA"C��f_��P���ȟ&�0���U��9�W ���v�Y��'�!��T�l�+�(�Y��r��+��D2��z��~��S;W�n)���O!m�	�E�A�ybM�V���2�E�gG��0%���yR�6g�YF'�-,�"iS��ީ�yBI�\�P�e@5&2\��0�y�h��ٓ�K�!�XTB�ᆫ�y2(��'\���"!���dH�$���w���O���CpD�ds�8�R�5<� ��'Y��z�A�\	��cl�N� 9�{2�>\Oxc%�B�#u�9��X�7J��G
O�7�I�(<���E_-xN�D�5���a�az�D��X�B<���tE0`˃���!�U�ØmAF��oB��"�!���2y���ʊA<�y�"�J�\�!���H�h�QV6o�n�	s���8�!�$U�9��xZS'�i�8���[�(�� ��ɔ���Fk2-(s�ŏe�t#�"O�i�� �+6��Ħ�%��Q0"O
�"��+^�*$�3l���"O� ��ː< ���#e� c��S�O��j���zJ�]r�g�?6���&-d�܆�ɲA��ā�τ8�tS�G#����$l��b�8с �7�
t��!^;+�jkfm?D�lH4�3k�i��iZ�#V�Sv�>D�T��+���U��&Z7Bf=[�<D���$B�~�<�$���p�H}K� :���<9�R�x\�,�!�� S^	:�G]x�'�Q?=� �Ӑ�P:��Β+�8�{��8D�ؠA��+'
d)pҁ�Y�>@X��<���'1����&N!g�r,A׍�8'`A���:lOFm��%W�r �)�u턣UQ����
OF6��7+�"�ؒ͛�=s��e�A`�!��M��� ����7o&�"!�Y5=��x��	�)*Ƞjv�	���Ό$O�>c�����)�ӇVz<ਖoE}��a$���2��B䉺2�@�"Jj��A��M-��+cDB�S����(q��H�g@�Җ�¡nB䉢'��d+l ��"H�s�K3=4z"
O���I$l<����[-lf8��'�:Da�S��y6���}��dX�'���R�2D�p�䢖1:��1#� R��!+1򓿨�>��V�Kň}���9Ex��Z�>O>��U��8 ��*��W�*j��z��Ëp���aAÐ8�P�*���p0��O����Ԟ!�0���"�<-��m8���fh���C䴟����'	�Sj�aʄƐ*6)�tJ�Y��B�I<'V����r( �(Eo].F���$?�S�O���:�I� (� ��(��
����4"O 8�ƩU7�L�����d��8s�"Op=pvMؑ*T�-�"f%w>���"O���V���_vVy�CE�9 �M!�"O�5����V:�;����$�4�qV"O� p���l͹l��y �M9���9�"O<U�� <&t����T�j�"O������}�e§�/x��0B�"Ov ��"�.<��V�G!>qqw"O�-"��|�P�0 �2X��"ObX�2�OȒ�;����#��,�"O:�"��8D|4����3����"O}����]���"ЧM�+�bғ"OZ	���ο~�J)pW���.��"O�0�d��W���rC��rx^��v"Oƨ�g�/,C����薓-Z��I�"O�\y�YmT B�	fQ��÷"O���j��8c( Bvd��q+R4rP"O(J�`����碚�U����"O��pSƊ7L���V;N��5�@"O8u�g��KΝ#",�:��3"O��-9O|L�qIC�R��]���yi�	���cQ>=�HXs")N��y҉��2̌�ό2�� �'���y�HܶK�̸#"O�-���kG��y�䎐o����6독 �R4� c?�y���-w`�J�[�Dը�E� �y"�#-�vE���*u������y���1�z���Je�2 �qʄ;�yR^�d2��p�T�VѪ�Dd�0�y�M�����+�%�A���y�h�%�����Y� �¡���R��y2H���SRbj��Ɵ��y�i	������J:�P��EV��yRj��h4<������p3 �5�y����F�`u�4�	���F���yR� �,N�4o
��H�/���0?��$�e�X��E	y�����a�	��,N�<N���8\��>:KP5�g��p�<���4� ���*�@�RӉm�<c��1E�h š�&Dʀ͢��Jj�<�t.�%0P~=��#(��E"ǆ�k�<�A.�f@�cBã>��k#�MH�<�0�٬���.ܳ>���I�b�<9��1BN��$�J�T��	���U�<i�� +���6��`�cT)e�<���I�d$I�h�I���02�Uf�<Q�X�,����'�(C�� �(P~�<A�	��J�Tn��+�)�m�t�<Yh�	[����%!�~�h�Bw�<9��\�;������X'��͒R�Pr�<��"k�H��ЭV�w��i��Zi�<�����@��%���=cX����VM�<9��Y4�I	c��X�\@�q�<I"���Fqaa��8� ���Vj�<ѡ3`5�T��__7���u&`�<qg�*Z	��"i�_7��S-�^�<!Ǎ��9טqh M��4S�g�Z�<a�jJ�:�V�§H�Xj|hH�kZW�<٧c�L���*�r6�-BL�<I�j� a&)�o{�4�D�a�<�C	��h�c�� o��`ƨu�<i�� U
h�[Q�L�h#D��1C
l�<�wƗ,�P���L���j�Ai�<yg�MH���	ط=����f�<Q�eڢ7���h�D��%ǖ��%(\a�<q��{�y1�$Z�@Z�zrC�k�<q%K�2|ؤp��&}��!�c�<iЮ3E$Q�q�*E�
yh��RE�<� J�uHb"�Q�ti�:+���"O��Q6��uN{&�%�M[�"On��!T.L���#5΃vz�т�"O����9c@	����'r�pz�"OL��B�G$<���#E�vǶ�ku"O��`�a��3�$yb�J���Y"O<)�)"uHvEbG(Z�v���"O�z�˙2��c��?,�Nm3c"O�4�RO�.Z���D�Xξ��"O�%h��ϴ[5��	��ɷ�B��"O�$�Aи?J,p�m̞m�F"O`X��D��'���5+�,~�J@�c"O�h1�DҚu���%�14�H���"Op�C"�ϗT�
���f�D���� "O8�ZN5��� ��Ir�"O~�;ꙻZ/���K6��Q'"O��07⎞U$=k�ˑ�k/F�c"O�� �B�:d�p���@(��'�\�a���8�Go�?w_�uzd�ӹ~d���-(D�����QP�<�0ҕ:���7L5�I�h��{����:�	@ /)n
���M2C�I�V=���*�7<`���D�@�1u�QܓU'�>�!�&t:�#Ǿ��K¡=`����ȓ�L9�-��Fiԙs�n�U�o��D��I��'H���ĎJN��W`�]#��(�<�����<�#��4f�*���»-#jXң �`�<1`��NZL�[����blF�
F�P����ׁ ��y9�A��6ml ����!KТ���xc	������%S+�~�N��w�@��h��D�;�z���K�7��i���:C!��B�&Y#e
R."����,N�_�!�ƳHu���N�	Ǥ�*"J� (!�ÁV*�Ȳ������jjqI	�'��Qc2(Ǖ��EVe�:]��A!�';��3l�	J:.�B�QWx��B�'s��XtdJ��#���v)��'�c�AK�O���8�Ǣ's����'���`$�L�\�N�0�lƦ68",*E)�G ���I�{��H�T�6\��`��,H{,���1n�>d��3}bBM�U�T��T��9������y2i'L�*$K�B.��� �~@�!X��$!��E	P�~�e/�JG����tiIȭq
bT`V���q6��ȓL�E(�gM w�T �a�>,�$]��'��<y�E:�䫒����9O�Tx�
�R�wG����ę�02��q�E �\��� �V��D�}0t͢c)G+:���hY�bX�#V�>�x��+O~ �%��[��p��4mbH�)��3>�
�� 	u��"=9E�75.μf��[	Ri���~2�k�Nx ���V)�@I80��Q�$K����i+�H̇�Iæ��&a�]j"萦O�G�h���,�8h�����h*���%�yh/6pL��#���Id˟)_�!"�K���BB��$MR�+vɔ;)\�܃g<d��%P�b�@��1T��D�A����(oV�0ż���ϣ}���  "U�Kz)��-@8�@��L�62�3(��ez���tG�A=�L�B��0��ּi2 թ��O����Ro���q	�E�N�1R4F��1��pS�X�+��Fy"MP/B��FA�4�����*)��ɑ���AQ��e^<PdF��\�Ⱥ��� "dl �e�A��xzǧ�4��(x�.��Q	 x����CA���'��.D�(҇�|���O:�n�G�oZ=�
�CD�ڧ7�(�`�����DQ�i��H�L<��~���"�F�T��LЗ#�>橙(+plt��H�}9VЙ����?��Q��T�ǃ��4��w(D�`�bBUkr��%oX� #�3�Ȁ�+>���Q*|V�\��i2B��a�:a%F
%�~U��X�=�JiC���]t�X�4�?�'ۨn��\-6\0���dTa�\H�ф�}�F��DM��w�'���z�	[�+✂q��
(:�4�O�����J�bΨ����7�Xk�
�A�"@�F�9G��yi���6k�d<%��I<7Ɛ��֊�;qQ���	��LL���)j���7e�̟$��̅hچ6�v�,��D������r-�П�CЉ�$��@��j�)f�)Z�7O�
rAƪ�ēO���0F��+�PH��M��\��,�v�I�`1��	�k��鳕��l����=�g�? "��"�A97FҨ��O�lh�@�x���%�1O��q��;��=�|�xdk��q�vM��G��7㦘�s���F��I<=��y���|�;n�ִ���W�R'�1�3"ڻ�Px��6��h*A�\	I&������D>>I�qn��Ɲ��	dR}@
Z�aC�|X%�2;���$��j��ٓ�$����;t�5�& ��/&8Y���R
�'_��D'˥u�8��'�[-d��Y�L<ѣϔ6X�>)�N>�~*� Q.�
L���b���ʧ%�i�<��CT�P �s�
�Kj݋b+Թy=qO�M�5�<�3}roF� Fꍣ!dO�x*�Q��R�ybK��P�F7y�L�3�"�/�y���^�p�����kt����AW8�y����8ۖ�!ŌX;aMZX�G�&�y��2}�����3����ƌ��y�� n����0�5��$�a)�yRF4Rr��B��˾-H����y���t'ް93�K�=�L�p���y
S���0��"%�4���F-�y��@, C
��Y"lR� d �-�yR��.YSL�����,P�hRAmM �yB�,=�0��#�M� ��%pāٔ�y2�M24%n��k�I��]4�M)�yH�g�}a��X8�� �$���I�r�����(pF�E� �(c��8�I�9O!�D0��HJ���[Z`$c�H� `2��Ob,C��!b01�1Of��g@$8MP���gA�ȫ��')b�t��A��;v��i<�����xU�t�aR@�(�Р��bުn����e����Ox�r�^�|���;J|�"�ٴ%1y�G�n�x�#l�A�<��H�+��=�V��qn�ReMQEy�`�����G�W��S�O����a+U!M�D���ĳ#��e�ǓU�<} 2e>͎��O�gt�P�lݞjF����I�<͘(�GH
�� ~�)��NQ�3�	6~�h��@�S�~\rdHI�hv�;�ဴhPM����oѭr��K|2�m� \�����2N'��@�'�.Kx����S����"9NV}�a���/u �H�f�M���r�i�b'	1c20p�OL^e����+s.��O�Ll��0�v����b�r��c5�OT] ��&n�7�>��y��Έ=��;BF��t�$�Ӡi*�<��<���'v[��� �>᥎΃z|��ƻ%.��#�u�'��!��ʶ���Ђ�9�v�����"?�1z'�¨;tzDZ��_I���8ⓟ���C>���GB�o�h��U�	�6.��S�g�����$��/\&���Ś6^�hQ���K�d�
�&r<�:1��I����.��N�6z��h�'�
9��g[j�'��Y��J�a~~�y�K��^�]3��� �|IF�V5�0��U�P���6�:��uZ��y7o�#��D�"�N�DBZ�E!?���,�4�
�J+}J~B�]�[����#�J�>Ԍ� �f
M&�	�_�Dع5ER�n�R�!�)��܎�;��	�:S\��g�.�L�E����I��<II��@�d�z�'V;����ņ'�h�AT*Ǩq��d9u��!C��l3�ݗ-1̉`4��m�b��,�O�m���!.�b�Ѯ�F���$�	4�0��n��(1��/\H؈x�@�!-�j�!��� N��M|�Y	h���"���`i��`�''�i"�I���B��I^FF�}���_J~�]���A�t�y!���}$���D�4?<���Z�=8��'�����DZ� $،�"Lސ
@s.O�X�.K3L285�9�'u���I��O�}�,�:��I%��}�&UJ�`᧍�5g��1N�jx�Y����+)@X��F\�N3�]�5�� �Τz�R���i֟x@��8y����.;�6�]�R @�")�d˟%eAx��)�)p�챰��R��p>��ެO2�Up��^��cb%5�Fa��R�\�`�'`��)V���(��G��,��=����jR�]�P��k�>��:��Otj!�B/�h���4��#[�z�H�������:`h@�C9����ՙ?�0MY0)����E��O�(c(ʫ
��q�5���	�t�����Ʀ1��>E���"4$�K͸a��]���8]q�(RS�B B�Ĭ[F�4B�$��������.և ��,��뚭7�z��I>��6�~��� ����5�p��Q�4� �+�.m��7O+Lo�t���i�!���sp�ā>=��Å�u^�O����NK���<�H�|xb>%�,^�f4	sg�.Ahhz�'D�0����V	���l��t�*qED[��I���)�p�R��O?�I*U�vP��7Q����%~�i���� h���;ɢD���/)��P)wY��X6E�a'zAɖ�'��0�RQd����P�*��4��QTi���~:.Ł�εd��Z�h��&��d�ȓB�Y��`"+�J��D�
�50Pd�ȓd���,�?}vD��p����2��x���/u�����M�}��-D�����F�\T$�Z:sa���/9�T�a.Ĵ9ӌXwE������/fI���(;��@�D1d{���a1R�K�ñS�} t�h� �ȓ ��� "�E��M �@''H��ȓr����4Cܻj$V�j��$L�p�ȓ8��ѥ�יn��Jr���x��]��J[��5��{�2X��i�.�a�ȓ*���0n҄KM^�$��~-�Іȓ&��Cä`p�QӨ��QP����䃗��l#���G��� �� ����("E�K�vm�����k�轅�ܮK�ΎJ� � D�V�[`������
�Ké[58���H0>e�̇ȓ��!�
�%`�i���&w�ܩ��*�`���*K�@�8��# I�6�z(��V]��¥�׵z�@��GְM�N���>ނ��o��I�G�)_-$��4D��r�� ���؄�ߊ�<`�'?D�غ�	S�j�!M��8�d�9D�|	rnU�Z�x0��n���1��7D�`(��'O�}�J%,qp�4D�,��!S�w2����'�,�BQ�7D���b��B�
Ѯ�#��B�2D���Ɛ�v���CH
s�́�f,$D�0�����l떼���r�X �.D�$Z��]�'~�4Yrᏽ�z�8S�8D�,��T:��Eq��Lz�:� '#2D�`He�B8tL`]`d�
;p�xp-0D����\��� ���Nx��@��*D�X���ߙQ/& ���2}d��'�$D���d�1	�cFM��d~�}SC#D�d"�G��\h��iQ�W�\<�f�#D�l�1Nɛ�8Dh0�O3"�
$�'!D����푕m��@��C&���;�!D��)��I ��B%@�;w�5�A?D������U4�Ņ�Z2�I��<D�$c0�X /Ц��.ņ5ԞY�Q,8D�|��J_���*׫��Z�`7D�"�×''�4u&ث"t��"��2D�lcB�D���������s�3D�T�@���i�	P�N�&	�3�1D���G�H�c��Gj�PI4�A�-D��ҳ��I�,Y�g$
���[%'D��a�d	�^+��R�&y�C��6D��IL0H$~ �t����a�$4D�|��FC6Br�i�c��6X(���ti8D�����ψ�D�"m�,9S�9�3�:D���0I�ny�Ú�K4��c�9D�p�4LN�(�:����_�o��pR!C6D��;s@\�=��QEʖٶă�+D�ܙ�
Q l����O�^�cf4D�P�t�Z@;��E^�#��)6D�Dȅ�K�qW����0��x��4D�ı2�v��9�b!S��p�&3D�$*d/�$D �%-$�� �1D�L�匈hT���K��P�h,D��z��.!FL�F��5f�x�!D�� &���ǆjS �˶��<�n�  "Ob��u�Z �L���?�6	�R"OX���aZ2vn��Sn�@Ű`q�"O
�!Q[�l_�t�Ƌ�ȔP��"O�XP�_�i�%#�EW��ya�"Ol�ѫd�@-p��ϙY�0���"OB\[�O䬐խ1k�ҩ��"O�R <{ذxYt�A���U"O����/�"(Cd��a�G<I"�1CU"Od�C�I�F�H��B(Y�ƍ��'D�×m�<>� ��LS�F��Db%D�(�֫���X�82"L+k9�3E$D�4��*�*Ar(;#�K ���k�O?D�0����[To��3�b�J�#/D��_{ 8��D��<��-D�,r�KY34��ʣ#
��͙��<D�h�0�B�BO𤫖��2V�~� G;D��p^�`P�"�퍼8tQg9D�0{��;X�v�Iq�I�xѳ�7D�xB�AуP�L��U�D&} ���#6D���Ԩ۱�����c��Dh�Ӈ6D��Ӥ��eF�PX�}�&�ʗ!��)y��h
�"��!(�!nB�!��{�pR�L�M�X� .J*s�!�F�w���=4��i�C팈"!�V#:4HQ�[��T�U��4[!�D\�)����M_���e��h!�	�sX��2��ǻ#H�]�ЌN!��]��.��+
 4JQ��F�g�!���3ld8Ec֯]2V=d�ZTk�0�!�0z�8 W�ǀ(%z�E��<H�!�DO�4Z���e'����Y%IS};!��ƪ>��R�K�2k(H��Ñ#I!�@aL@ �D� �z���P!�\#����\�d��ٛw�!�J�B�8�"�O�HOޭ �k�!�$T�$�9�!�J3s60R�MU�_�!�D��:�n�a��44<AA�N�+V�!򄚟4�Ј�V�M7�ˁ�,c�!���;^P9v�<XH���4:
!�$";<��}�Eb$0$Oz�(\�	f�BD��3����/��͒�*ѬуV:BP��,V:=Ȫ��I�u��8q�l��>^��
� \
B,� �dn+�!��1�Ɖ��F>9�l��ǔ� �d��6���K�6?���H?�#��+ox�*���ݰyc@9+�!�?/�B�	2%�t��σ��C ���qBc�	g��HQʁ����`�'Ur��'���"#���y'�_5�������&$�����>��K�M��MAĄ/��!�ªR(p�E�%U�|IZ���n#��D�V��9Q!��p�Q� �S��+���yp%��,ި���<���iw�LQ������mV��?�n�e�@9_S�ICvC_:".�)��-֒_���e���0>8uC2� ��W)z�T�8��E. �|�cGd6Eh��ԍv�P��ޟd�q�'���hŮ��k��4j��MCd% �	��-Ar��q�<�Ԉ�x�}�Q�2 �Fh���M+N��I9��Z���S�[��%�^?!�DW
+���9�w�e��m(?��90�'����P��!𝃃�׺@,uyRƝ��� �F��~��	Qw��6-@&<���I#&�ъ2�85<�i�BF-v��a��U�H�*@��(O�"䎇.p��1E S�`�@j�?�k��D>�-��h"wϾ��gթt���D���4bߓ[p�Eq�*�<%�%�f(��.и%����皳m�v�P��Yr�I�?aԻi� Ĩ��Z}q����Kaj8�%:n����at��xQș�(��4%%�6;[�@������RnO�WQPi�s%g~��hq8O�[E�շ9]�,̻g���<WUru�,9�|���v���˥"لFq�De;^;�k!g�$�z�+&a��UZ ���4�?���z�*�v�
�u�|�?A���E0d�1�L��q��@~�'[�1J�%�#3�qC� �<u�'7Z�� ����ͦ(�ű2�]�@u��0p�84�L�"�Q(w���DT�K
������D�3F���y��X?Z�H���8bV�Q��ן��:�⅁g(��2�=����8_ b�"RD+X4���`���yҏ�?�>�i��)i	�9��J���Q��!�fZ���1��>t�	��k�n	@@�H�[4�C�ɭ<G0�9𩂺 �"@q�@D�����#D���	�%v����|bOh�h9!���q�l��Sm �Px����uѮ퉀M	�O`� ��#�X���[�ޜ؇��)\��h1�Sa���!xD��E�M'�����ܰ���S6t&`+L����5����X�!�d�$2��� E�E2�6�p�)�6FƉ'�}���S?l�ɧ�O�h��`
UF�����:&�
�'�5;����>��t����9���0B�0`�z��OV��@gQ#ڑ�Q@Q�~^�{6"O�{���qb �Q�σud��ʳ"O���f%�L�����<[t�R0"O�$Zb�Ԏ����0g�+W(�3�"O�M��؃]:V ���� �d ,�y���7J�"��D%�U,ҽ0�͛�y��Ȯ\k2��!B�._s��h���y���e[��J�Y��飇D�y��M
'9ؤkAi@D��(��ʫ�yR���F�d̜L�4�����yR�]>	�����8ARȊ���<�y�[�5��,{0�^<k4ʙ���I�yr'�+M9��y�Oזcj�c#ȵ�y�ON;-��ԡ���]�~ Qb�
��I3���P���	(|�� G�5c�t��Ƥ�4R�!�+HSȀ��Ww�re�X)=�r�O�R5"(?�1�1O H�p'�S
1Hw�5,�}�s�'\� g�<C,Jv	
�L�PDȮT���Sa��`؟l��#	�Xe��S��>I��)ؗ�/��%<n�!��OE� ��U�3�'(���`��U�"{����"O�d��l�Zm�!	%Ʋ�V\��C��C�(��֓>E�dD��v����eN0ލ�g�nX���ի3h�O�x����	2��� �� Q��!���&��;=���Vl�3�3X($�Ck�l)��`7�I�N`,�"�\�Ñ�JM��PF�Di�-���M܇U]�*��Ύ	O������o��u���(k�줋��Q�]���!�� 1@�↨.?q3׋e����vWD��451�;'��HT��-Z-�0�VJ��Y��i#��0D�Y![M,����Y�V���r�Xoߌ=�%���Su��!(U��'>>}���)(�ǐ<jȲ4���6���H$n��D��=�ʟZ��tM�m?�yJsh� ji��%�DI"o}����d��j�̄�SOwC-"��*Y�F˓{�p<3tY�-�j�
���ɵE�Ȕ���@$�{�F_/ܶi��̩��O
�P� ]�Fi�O@a(���`��[���Nh9�2�T���$��E��4� ��
4n���Pw�E�y�^8���$k�I�!�� �K�H��S��*׬!c�Qu�)�g,נr�N�Ѣ�ʿ6�^L8u�'�<:Rm���-@#âێ*�*)RM@#��l=�T�Ԩ�D+��O�n�ƨ�N���$�yo�8rWΒ�&\`	iB�Y�����$�"8~+��@k�C9H��!C�2uG�A���Qg�&��'>I pe�:�>����¸�v4�a�*��\�n����� �ɟ8�A�l�*3�nԑ� ��!��#�$
�#�+1���JMж�3W�^�㒌Pʕ|^��-y��3�;-P�qE�D�4M!ФmCud)UF�:,�$��4�@<�JنE�~P
c��xUj)K �1+��e�'V�I�e� ���ϸ'�~���+Q��2��˱bX��X��t�r�H�E�t,��i�ҦaإpW N�vQ �G�L��0?a�F˿9��[A'�seIk��NO�'���2��	4�?	rD��VH����V�Ze��E>D�@QÉq<�����͚h��5�6�??��a�7��K�M&}��i�*DX��D�	��T����Ub�!�D�6y}��"���1�샧M< h'�蓇�>q��'�l�eΞ�ư���
.^R*�X	��� �<`�*LO�n�xU+�?r����"O�	"�h�T�h�0IT4��k�"O4<9�n�'�ФE�:��e"O"�`�3�Ȉ�s�Խ-^r=��y��w�H])G��&�N�A���3�yr��9W`��<�����Fِ�y�U�>NP��Cڑ	`f�1���y���&L��� 
Z�{�p-X�$2�y�)�q�-@d	'q�<�!k��y��8іL��ʬj�j�� ���Py�l��`��eívFe����[�<���hYp��Q��.jpt����_�<QRC��e�"ɒ&%ϨaRD�j�#RX�<��jڲ(}Z�)�_/D0�*4��@�<�ï�+%�\|рO����-k�Vp�ȓ!^\��wa�o�`�0+¯i��y��{D�*���3r�9p5JR!	*��ȓ@��-���F0�Ha�c�:�v���b �� g��I��\�f�K=rM e�ȓ&@$�VN�;F��p"A�]�U�ȓ#|�Hr� ����P�+�\y�)�ȓ��X�#W?!���ĆC%c܅�ȓVLx��'d?���%W�4�\���%֜��%�F�}�X ��Z��: �ȓq6X豄���;��r�.�U�zQ�ȓn(@�)�|�CW��!�� ��o@��8E��/tyX��|�����\���`U��IՀ!��B�t^ZL�ȓc��Q:e���$�������C�I�p�d(���vÂ8 �ɐZ�lB�I�D����Qb��L�H��$���9 C�ɵcʴC5
2?~< ��X�M]�B�	,F3��Q͍!#L�� ^C�G��	3Ռ˶j�M���5��B�	;���0p����0�
C�i�HB�I_������[����*ߑr�C�I($!H0��"7ӄxtΜ3�C䉹w���"�O��J(X�-�~C�� p/�1
���p��5�
�qHC�ɛ����f-w~�Ń&�ǰb�&����2@��� ��OFz�ceHݍvq>��!B�t-!�d[�:tЅ�T �oz�p;��Ɣt!�����dQg�bvH!��j_�^!��/! p@
�HQ-`jx��(�q�!�K�Xo�Y�ؚmhr�[Շ�=�!�$��DŴ a�&�GV���GGÙQ�!�D��x�a�!��#S�0��7�H�/!�(\��-�-�� ۣ(J:?%!�$�x�&p30-Sz^E�ΗK~!�$������U�e��VH�G�a{��!�;y��1��# �qJ�>+"��ɉ�P��Sl# ��-�"t�����K��5R���&"��ذ㞢2��.P�uPFjد�Q�b�ߟ����=9��/��U8��%dnh<1�A	"��������b>eq�J7j7�<05���QJ*}rJ��,���=�g�I�7�!��%IZ��8�.�z��I��,M�?E��dWbF�南�^�T��f��jIt�80F$�)��M	��K䩋<6��a�I�u���҄��6��O���'o9� @�,�v���TH�]e�=o���'B{B�"��h�p֝�(丄A���\�P�!�S8/��݂R���U��)՛�?�B	8�l��!ɬ/(�;W	B:.��A1�ƫ8�����<�bh���a������Դ���� D$l��c��6x�=p��O%*qǞ������'G� �Ò'�)����d&U��x�<�N�d�L�':2����O�"��i!N�Ь �����̬�ڴC�<i*�)]�4ҧȟ� ���a��O��a���}D�`w�ٝLD��'�J���s�p�B����w���r�'� �b��0h*H�P�`Y�`f��`�'+�lI�*Z�k��p�lZ$�qC�'�!�	:8�a�J��,��'>&刕*�3:X!s�ώ�%`(i�'�N�R�'E�D���8�ե�h�!�'��!K��W\*J�x�c��| ��'�0���W�����A|J�`[�'J<ꃏ�4��!�&,ɍt{(x��'�����gL�j�t�Pa�>MZ���'
���E�0K���gHח;�@��	�'9>[$�!�z,��hߏ0d�@	�'�28���'aK.�k ��Tu�9
�'!�h��Rk�0`0ϝ=E���	�'�\�:P�*�<�����l)�\��'D���ց�Mk��0�R�1˰x��'�|hb�o5��� � v�Ј��'�~�{'�q �@�cK1D���	�'��S�hA�-�"E���3>Ǽ���'�j�r�"���\�4�ې4m$y;�'��(�� I3z~����h̜{bN	��'�^1��@���>� ��ȏoM�,��'͢�� 	]������C��m���'��ĚQ�ӷD�LШ��'���'_<Y����A�p��A+C/@��'��l�7Dޞ�\�Sѣ^7/ҭ��']t�O�$M�|ʑ̄!�b���'�V�Z'�4u��q`%��rTr	�'�4��?LN�uY���^8�
�'k:�	&����uc׮�r��(	�'d��t�]
S8@3wF��5�n8h�'���tK�=f���Ӿ&�`���'6J��&��C�Б{����*��[�'~Ő�i�<���Ҕ�ܼӸ�Z�'+�٫`�ih�ys��:V�ȓ}��;W��L��E�#�E>�T���m�|8a���
�>�(����챇ȓ.����u)�E�Z<�rLZ2V)���Jm$�˧�	?�|y �Էz���ȓ<n6�Q�&�q��x r��6���ȓ
��X��DeS�]���T0!�����&� O_������+�ܥ��]�4@���6N.t�P��%zl��@�Hp��	 Lb�sd�E�w� ��(`�hBW��X�p%�b�إPx�U�ȓd���[ЁՄO��MSŅ�f ���8�\�����J�[pC�: �х�3�j5Q@�0jj�z1/]�k_&t�ȓfK��h�)I�|�
���.[�xЄȓ(ZF�2��KrмR"��6���~����h�{i�z�L��Ψ�ȓV{<���(,ty�q �ȓT`b��\���#`n�=Z��U��e�B\q�� �Z�ⱦ�5h+���ȓ{�Ʊ���f;�@�� 
��ȓc0$m�[Z<^�[�M�h�@��8��k���10�v)�w�� m�X�ȓ_���O�4��4GԒC��ȓ�z��PI<Q�t���p�ȓ*�m�鏲o���B���K�Pu�ȓIݼ��cl��Oe&aQ�Pr���ȓ0\�� @�Јdf�0�VΒ\xԆȓq)>)� �V<j�L)��(�5?h8��S�? �9�T�j�L�6�\t�:"O�	hޖ#��$95�9�Qq"O��(ek��3��@qmGf���"OL,B`C��l��$j�-��l��|1!"O"�!�(F�(/��xЁ�aۄ}��"O����DJ�THF�G1��]`"OԐjf�Y7:6j��g�g�и�"O`}���#��kUǈ,�\�#�"O�h�KܹD-������9~��T�"O��1R$�!_K ��"1��"O&=+L����d{bVb�,	�"O���완!'�y�#��%-(Juj�"OV�8�� O�x�H�@1W�|s%"O�x�%�&���I4��-E(R�d"Oj�8f.�(�VM�Y���3"O��X�L�1V�ք2�	ul.�"O�� 0�X�\�}RP'�����N�!�dA�~�1�I�c�|��u�E�X�!��4'P�9�ʜ�J�{�E_*Y!�D�������-��hjB.!���/�t�Brk�R �9'���FN!�$����áF���l�,۬a�!�Q9��U[d!C#�V�Q�=�!�DO�zC���FX�"2����D &B�!�DX�:�rl1�� ".(Z'iU�*�!��ӷ^/��K��3"
� �7r�!��{�� ���$ �����p�!�D��o�=��Ef')�f��O!�N
J�jTҷ��(ƀ1���&d3!�d]�
�%�w��((�sfeݼ]�!�DШ(�2�v�4	�!8F���"�!�đ9e�@���/bɺ�h@��!�$���P$P�g�f�*a�F�?5b!�ҡ.8pԺ�l�R����p��gF!�D�+�zٸ���:&��d `A-+!���EI�u7DN#��i�O",!�$� Rl� K�|w���
Y�K!���3����ǼcH�w��2�!��J��s楉,~oD�G)��f�!��*ArnXSpc�5~^��e\d!���="�����ޖ
�h� &I-oG!��ƚQ�}�$@��d�$� �P��ȓH�NM�rH= �
�F�ĂQ'�A��{8����m:=\���b� �tć�D9��4�G����=Ay�d��P����OE�51� RN'H �ȓ>�^��p+�'Y�!� ��"j�9�ȓ㺭�`,��b4���P�I�ح��=��I�NDa�yä��	HX=���42$_6#��@�� ��(�ȓQ��ċϖD�
4H!O۸Q�2��\!0�ɅO|��3A�ϝ!w��ȓ�Ɛ2��#鞜;g�E�2��0�ȓe>�UcuHA]���sҗ'�DЅȓ7ꔜ��	�dI�1���͐�lD�ȓwc2�����-){��D�<�X<�ȓ9��S1��V	���6L�VZ�	��,�����!XH��"/�:�6ȅȓ~]T����B�0cj� ����Nk�8��KP�2�V!k�ʚ3^���ȓS��9��M1$6b@�b��H}�H��o.^�8�I,]��s�&�����ȓ_��ӈ_�`��rV��P�t��+`P�ۦi�%d$��r��W�A'�Q��S�? ���N��6`��C��9]O��[�"O��: %��,�?Zq	V"O*uB)�#cy`P�ci���ӗ"OJ�ҷ��+���c��8���"O�v//R6��'Ƚ�� �"Ob���D]	Ն�!'L�^vLI#"OJ��%E�2+@1.�+����y*7����ŏ%���y�͘��y�#[2i)7K��R4r�*�(ɚ�y�v�(Q!V�^	?h�3�gƛ�yZ��	�BA13��rC���)
�'���d�8X�
��g�B�4�H�j	�'H`ěT�A�N�,@�7���,��'��|2p�C���H`��( �)��'�`�{��~f�A�ϸ O�y�'yT�k(����0P�f������'���q�U�6T0�@�{=�,A�'PL ���>hX��v�������'��T�Є�Z���;��C2QxHq
�'�-��i���}"��ǈ~!P0	�'F������Bl��#�?rԵ��'.����#r�E'2s�a(
�'�^���n�?"����$%$0S�'��%��E^����B	��'���C�Z���UO^���c	�'B~�)j�V:`{��P;�x��'l���W�!RPkO6G���'����(�<q��� ��QHL��'�&�b�%\�x�*�it�x	�'2R X�J@'�h0AB�:{�h��'����ga��s���x���#yM±��'��02���qc�	X���?T�'(<ЁgØ$�x�@��n��#�'i�����-�!��J�5D�X�Qbϗc��Q��2W�pa�4D���׃̓���g"��P��e�0D�)W/V�H��1��O6j�[@d/D��A'M���lb(O%a��i���/D��'T�q��yH����i�-D������t�쀑 �'i���6�7D�T����y��+1aZ\ИSr 5D���a�So4q��WD����*4D�H�d�X�Z�<��%,T(��	�dG$D����#	��X�0��.,�`#$D��B%h�P��L�$ʷ�!D���9_�Z�Pd��<Tu�m2�� D��k��.D~A�Bn�8�c9D�Q��� ���s�Ю`5�ZA�*D�x1F�>"�Y[Q`�	-8d��";D� �$�ͺYC*�蔧��ỳ.D��z�ȁ$fhD�A�c|�F�7D�\�������勝Y���3��5D�A0�D�9�"(+@�E(hf��`C�3D�@Z��Z"?�d����?afYY��-D�$��d�.I����4:�Har��,D��8��V첀�`��u��p�w�?D�Ȉ�Q�T����nJ� �wI3D����O���z�� ;���Ң�$D��9���[s�ÕOT"<�l��#c6D�T���Z�U��
�E��N.���7D�,¤��
"sl@�`�S�S��*:D�(B���7�Zhh¥,/���@/9D��� f4aJ�ӕa�z�ڑiB�6D�`륦ռ�6��m^�3U�9є3D�� ZX�A$Z�TA�!Ş"�^��"Obu��`�+3n���	�=/�|�*�"O�)����&��4��fR�\Pm�"OL�aF�[_�(5�@ ��V�\�"O���3�߷-���R"�E�b����"O�D�    ��   �  c  
  a  U+  �6  �B  �M  �Y  Je  �p  �{  ��  ��  5�  6�  ۧ  %�  ��  ��  8�  ��  �  ��  #�  w�  ��  �  R�  ��  �    � � $ 4" , [3 F:  C �I QQ �W �] �b  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z��Yb�с�5|O�"EG�;֊�R"�O�~Q:�F�'VP���Œ�'蠢DO�	J厈���4D��@Q�Ђ:�|@��Tfs���(D��`D�J�=Np�A��׭7����Q,%D��z�oV5H�r��.Q�����$D��p�L���Uk��B�����F"D����`���2����{�& �E�<D��PL��j���H�G��:f;$��S���T����t��n�����^�D��� �F��9^	�F�=[`�͆�Im�)H''��*-���t�S:E��ن�	�H���
�e�pڶ�3<K�̆�;�؄�c��v�`����֭wXވ���t~� �6XvD�e �8�HP��E��y�D�9;�px����|	J�fƈ�HO����"��aA'ݥtǽ�!:w*7�!�p��`�:�4E�*ɠ����Gu��E{���\�B��8�d
5s�.,�(�8zE!�$ǈ`VaR�킍wz�q2T�
�-!��QI�V}z�f=n�����,a~�V���J^X+ָ{�儏v(p�R��5D��)��?1� Zg#��o�2���(D�p���%HА�(��� ��Ȁ�"lO4➼�eO\;xz\���%$��1
!D�p
`f	 CHA�0���-ƵH%�<D�pZ��CX��wf �B4F<D�<��"J!���#����.�aDO-D�qU"Ո0<�i3K��$��X��0D�� @��#aǵu0�IՊ[�zl�s�Of�'�6�NQ���I�k0L�F�_3��݃�!X8Xaa}��i�d	x�Ա$o��\�j�� ��Vhm&H�(#<E��4'u��D��* a�<x��S�RU���Ms�B��D��<3�Z�V��#YRy��,�OҜh�k��Z�:i��m�N[S�'����O�4�V� �ń���/( H�"O:mKw����b�GF	ڷ"O$��$L�GE��;A��t�V"O�p�##�&6yK83�� ��ݬ�~��'�̀�=E��' �R�yB&Ӽ!s�$�DH�:�y�DކE����B�
}x�^��'J�{�A�^]~|ӄԅ<(��B'	I�yb�����1q�E�-����ȗ.|�B≎;삔t�+I'�h[���8E��B� :��)2��a�,���	�3HԮB�	�s@�@���d�j����P�B�	Z�
�"�7d|�b�KD]�B�ɝIhZ�q����*�y�JO�jC�I�ynD4�7@ɫ	�8��B->0�>��}b�f�qiA�'-P�i&�G�C�z���DI^�<�sh�E$4���(�D7�)Z`?1�]��m�|yr�S�\Ӥ�#��J>�+"
E�V��C�I7B�F�v/��q̚���2j��tE{J?�����3>k-���I���A(6D��u@I(S"���n�#^�u#S�y���>9��'��	�E�l���4�\#�4����'|��R��-Mu��;�!a*�e��'��D��EY�3�F�4���Q'��+��D �S��퇺V�N�ر�	�<y�0��+Z�yAP2ez�=Hb��##�А
��~�ў"~�Tӂ���`�[�$��iD�Rԭ��a�$��΅�U)�%a��.P�l��\�.��hǾ �8:�a_� �����B̓'@�1�F�z�BQ�M����ȓVN^��ؽ���Qp§ ���n� �EE�0��Qtn
&V��_�<�ەi�#G�L�f�I� 	�ȓ=�r!f�,`� �2�1�t��=fPH�bd�3!��,�
!H����l����JƑ@��\��OC�f�4 �� ��Q���
� ����[�����-��l@�m�!_~����$��2M�ȓ^`�ђ �8z�Qb�1n�Z���.�C���J�~4aC.$@�ȓp�D�z��

�V1�S)־�ȓM��%L��	B�� �
S"���|/���%�3-Yt��N׋]�����.�ѕ�Q�F&~���̈,M�]��t�����^�U�FӅ.��S2���i�{�J���?N䉇�����fE�,Mq�(�,D��Ѕȓ	� �� ɠ�:��Ơ��j��-�ȓjJ&]!g�B�x���blV�k��U�ȓ{R"q�N�!r$0QR�&z�}��T��a��W(x�]���"^���(�ڢFC=�8@��j�g�pQ��G�"�BG"f��lљr�4�ȓ�M�P/W>o���x5�ŕ"��
�''�#r?B��K���a���
�'\�P��mɀ)%�;���
�'�����X�v\�[4	=oH`	�'�����U(���i˺	0����'4Z��[1����p �YL����� E�����Y0�)�J�iw�!q"O�q�ʇ�gs܁�˓�*I!�"O�Y�6���I	@�R�`M�"O���# R	
R��0K�B���t"O:�!ck�a��L`Æ�'��xi��'��'&B�'�R�'r2�'��'u��W)��C�5@��J�L��'��'*��'���'�r�'���'���L�1d���XC��qՊH���'���'���':��'�"�'p��']�e���nA(\�ƪ�u��Y��'�"�'���'|R�'���'��'�����M�	`���r��k��y:E�'��'j��'���''��'��'h���@0
����V�V)qJ ��']R�'���'m��'rr�'z��'MD� �^9D��8R/�)'M���g�'4B�'�B�'|b�'"�'���'Q�����Eg�j��4@�(��4�'���'���'u��'$��'���'�ژ��-���J�_���ze�'��'���'M��'J��'��'�\];���u�eナ�'-����c�'u"�'�B�'/B�'�r�'�2�'��+I��``I ��7Ȱ5�#�'}��'��'��':b�'R�'�ʱSA��,ol`�2oH�=�����'�'�r�'Y��'zr�'�B�'�J�-9	⬱B�W&S���A��'�B�'�'K�'���w�
���O��[�G���"�|�2�:��ay��'~�)�3?A��i�BU�e���Z0d8!`%֘ Bh��������?��<A�M�	S^`aCN�#s�RI ��/�?��:u�\��4��dz>���'���5!]ZA�0��~���mS�`bc���	ly�
ff�ZF��Jo����&44,�ߴ>�*e�<I���'i����!T�(�+6��q�'�4s�n���Ox�g}���M��3W�V<O
P��dٳ2w6�a ��>
t�-�5O�牛�?�@':��|"�Ql�,°a��A���Bq� 5t0͓��$%��F˦M���7�I�(��9��������ߦP����?�X�������������glJ�
0�H\�Ũ'ʗ"h���l���^"#Exb>m���'Dx��	�Lxf��+P�N��dr�h\�$�Jt�'L�	��"~Γ��Gf��F.�9��f?i:�ϓjR��偫��$�ϦQ�?ͧL�|hh��v��$��hb�FAϓ�?i���?ib+���Ms�OB��+���L�f��:�=R�Uj�dKFUO���|z���?���?����t�'��)O�X���g ��(Ob�o�t�,�	������?}$?岁	G#��`d��]iH���KĖ���C���ݴ:������O;�$/C�Ty�����Ս@�`Ԡ�ݗ|\�h �ih�˓2�u 󊦟�&���'�]���ȈW���c��:��8�'���'�"���\���41
<��_P��n��m��Qt�!+=��������x}��p����IԦ�"Ջ�9؜sW�Lu�Ը��L&�oN~r㊍3�N���6��O�fT�E:<�$�N3�N]�����y�'�b�'��'V"�i\�j�0���I;t�:��b����O��d�즵`�gl>��I+�M�����6�3Q�\0j�.�n�:WN�$�� ڴz뛦�O�Θ��i��d�OB�w���V�`��$�[8��$��lP�`h>LH�'��'�	����t�	�]�D��P�f
!���<I��	ȟ��'�6-t#H�D�O����|���}*dt:u��'eP$`t.~~RĮ>ac�i��6-�J�)Rт	����kb�]�g��,#To�-<a/�?�MqX��xm��9�D�&6"q���39��°		9.���O
���O���ɷ<���ij���lѧ�r�˱��?��Hq!
.,�b�'�7M1�����$v�~��'-�Q����Ty�T�@����ܴ<,D8޴���H'D�U��O/�	�R�>���LD6I�бʗ�M��	Oy��'B�'}��'|bW>���h�=0�j��-j�~��o���M�kM��?����?1K~���w$�Ҥ	Ͽ5�`R�H?��<YFfoӴ�mڳ��S�''���ش�yR��7�!be+6Np��p���ybA�V�@q�����d�O��әBIL����i�������)K����O�$ca �O��m؛��?|��'��*
>?�J��>dд���ٯ��S�������ē��9k�4�?�)O���F�GuhB�f��,v~ũ�:O��D�&?h�0���LF����?�y��'��9���v���kD�)��Q��6Z�8�	����	ݟ\��J�O���<Ab�41f���i�w�����$l�I�c�<���iM�O��3BS,�����a:��3�N�&5�dxӔ m���MK�`ͅ�M;�'%�wk4��'-oj��BՏir��H�ќt�NԛH>i/O$�d�O �$�OT���O��$_�NB��!L@��t;dϲ<q �iA�M1K����'*��֟���'���e��N�Z��'c�@D�i��>Q��i��6��Oܝ&>��Sߟ�PcŅ�l,���B�zv�IR.Z�<Ϝ4�V ?y�d�z��������dV3oU�HH�`�	x�ܩ:LT��$�$�OPa{��G>�4������q�;k�Ԍ���4�d���D	�0pG)�!'`�Q�9A���X}��'���}��2�iϜw�v���.� �81G�Z,8�P7�u�h�	3�a 5֟���*�{�? ���gcD6I�HHI�I�*!�F7OD�$�O��d�O����OZ���$'�n��D�%-�(�x�M |m,�u��Oj��Ʀ�@B�MBy�'��'k�TF�U���Ր2���B�a���7��6�q��	M{(,6�}�$x�fK�0���ô"�x�&��&B!���)M�M�0T��N��h�Kj��?9��?���t�}��ÍEO�����A��q���?)-OX�n�%�<5��蟸�I�?���-$p�1���a{5��62�����D�'aҴi�D6*�S7Z^�@��Ɋg��4�CDN�;��`���Մd��y�&?�f��h(#0�m��`��?ͻ��ו�-Z@OC$|��x�&��Ɵ����8�I͟L{� p>-�	iy�p�]x�o2>�,�qT�I]����h��t�ܟ�����\�������[��a�f� ���-�b�EIXw2li�`m�Ϧmsܴ6I2D;�4��ě�&�&� ����SR�h8B�cY���Fȁ-iLz=)�4����O���O|�D�O����|ڠ�ܲ��圳M>I�sh��9�X��ݴW��e`!O��?Q��2U��?�'�?�;.	4������sw��	F��(�:aⰰi�26]ݦ����O�`�v�i���}��2Um@�EP�$�v�����,X�H�h�d�Z�c��R���۟��wC:x���,��.�qA����|��럄�I]y�x���d�O����O�p���:����-@�K^��f�O�˓�?��O��$h�lody��Ee�(Q��5��y"�����j���� G�F_����u�FM��P���'^�\��I�,�\],B��D�tg˝�?���?����?�����'\2�ޱc~���"H�#����@�+CREz�� �g��O���O���<��Cs�Jw j�y2BU	To���aT?ٴ �v�mӪ}�d����ӟ�j����Ĥ�nzd8�Յ�Npt���bJ�r�\$�'9<7�<ͧ�?���?���?yW"Q(�u�Ҋ�|��\i�m�����榡��ʃ���̟|�OB�'���CDX�A����!��)�1@X�X�4	w���~�
����	�B����T����Kw��j'�tSAaA��u�@��\�ƣ-2R��Py��{�P�1q�Q�K�;r���`,Ǖ9=�H���?i���?�$�VA�6�)(O4�o�:f���S�J"�"q�߻#�6�a$@M�:|�ɽ�M[����O`��'���i#.7m�	���fY�=��[G��#5E� q��r�t���$xćH����-?���n'֍Z�LNbi~%t��l@�D�O����O���O��+��H7�LI+bOF&<��geahj|	E�H����Or�l�j�'���'=�	�8[��*	U���h&�@ `� <�۴��$|�!Dx��R�6m"?)���:�����ag�`Dj�?��m���O�q.OT�n�Uyʟ���A�3�g2�!�B��"<Y2�i��Q���'v��'m�2Q����D!��At��<���G��̟(�I���S�D@��u��,ФE=
gIG�Z�lG)����<ͧk8��	O�	(��%�V��=hv�iѕ��q*N�������ß��)�SGy��c���1�πF+���WKR�b}��"������O� nZt��L���Ŧ1�!d�!u������C���"��?YߴI��t��4���к�����$v�˓l�,hs J�mi,�y��g�P�͓����O��d�Oj��O����|�q����`)Z�(Ҟ_U�h!!��a��䐧E���'/ғ��'�7=�8<B��M1K�P)�� E�m�ń��=!�����|�����5�Ɍ�MØ'2�LS�1��`�㚘z�Y�'���J�˟��1�|�Z����ß<qKS�t��	!F��L�:���NX�� �	ԟ���^y��{���Rf�O����O����P�?BP��%�/�X�>�I ���O���1�d�hb؝��-��M��a㎛ a���O.�Z��+(�&	@Vj�<���O���DX)�?�4�67��2�"�4/���C�/ɟ�?���?i��?Q��I�O���#X�$F��b��d˗��Ot4lڥ\�����ܟ� �4���y���x����ABJ�,
V<{5���~��i?�6m�ʦ��p �榑��?A��ޫLD��)	<
쀡�t��'
����R#$p���J>�.O����O|�d�O��$�O���BO�r���:��]�tw:�Iϼ<��i�ɲ��'�2�'t��yR$w���GF�¤������(��Fl�F�&���?����6}d��.��v	��D�	;��b��H��59(O�HH�W+�~�|�[���q��3`,��'��cC∫�ƚ�4�	����I��Siy,~�zةq��O��%l@�$d:�+N1�Q2T��O�Ql�F�5����M�Q�i�7��=�] �%ڪ$Gة �G�a�B��q��"$J5�?e&?��]91@Z�jr��
�]g((X�9O"���O��$�O����OL�?�fG߆|��+7�� YVџT���@��4<$Χ�?��iS�'��pf�0�`4�dC�1*d��.��Ʀݚٴ���NB��M{�'�b�N47�Y�����pȬ[3,ڣ��5M�T?�I>�.Op���O\���O)�GV��L�@lD�\�eJ�O*���<�i��*�'	��'�Sy��j!E��|��`�7� ���	)�M�5�i�XO���$2˔?_qR��W&�f�x��H�H��eF�o�b�'C�d�q?AN>9��t}���e�m\`	���`<A��i�l���k7%k �1�a�>IV���J=���'��7(�I���d�O��� ̝4h<!c&���BA��O��m����m�w~�N4��%����� �Z�H�SsRl�@��h �(9O�ʓ�?Y���?Q���?��򉃳t�JH+%�7"@%�q�L(�f�oZ��f�'j���ܦ�ݛX�N�SQh�1����E	ן+L=�	Ɵ�K<ͧ�?��'�>aK�4�ykT�$T(�X��%��	�����yb��ue�l������O��D�^�ʹ�RE
��r<���%hn2�$�O����Oj�C؛�hq�Iş8�ֆ�0/.t�RR�//\حhDO�'�$c�O���O|}%��Z�LL9s	BY0�Q�N
a�e�������jBwQR��<��'_nJ�I��b�
0Pj�K3�ϛN'n��A� ß<�����I��PE�T�'�0a�&��W�H��I�0f�|��'�7ٺt6�����4� ����A��I��	��U�77O����O��l��A�~ o�g~Ҥ��u���'`�	!cJ<)��	)�KN4��TIL>!-O���O����O,�d�O�!�ǋ.c<A�T�Aú�Rb��<�e�i@�X��'��'��:��C��):�q���p�4�82��B}��'6��&�󩘖b�qs�B�f_Z�:��č_�����v�z`�'%n�S��_l?�H>�*O����%[z@Q���	N�.�:`m�O`�$�O����O�ɱ<'�i��p���'�!�L3C�5�%�
C[|�W�'��6�(�	���DP����4�6�	g
U
�d� E����S���o?&�ZѳiU�D�OX���MS���tP���S��	��L�O����C��N��y���I��	����p��W��,`2�AB�ǙGO�`�E���$�OJ�m��I)\��֟�*�4��l��y�C@��aj�m!e@�R�&��V�xB�`�ʽnz>H! �=�'݈���]8� �YƍE3?�I3b�S0�ҥ�������OZ�D�O��DT"��Tif�ށ@��4�U�Rl���O�˓A��fL�d{�'��Z>�X�N�Y�9�Ck	j�!5�"?)eX��+�4Tꛖ�$�4�l�I�-�<A��2�VɁ��>}1<�A䎞�z(r7��xy��O�����[I�	Z��ހ.��[S+C�n9+��?!(OB��<���i��t��ʊ!Q��A���T�;w)���r�'k�6�;�I����즍�b�P*D��`�pX��DG��M���i�豓Ѽix�d�O^%bA�۬��dR���G�8�* [�$�=3@T��kx�T�'�B�'�B�'�r�' ��`���	I��bR�K�>� ش��A��?9����'�?aw��yעܦ(B<X�F�P4"�$�� J-���c�.&���ZM���Ӥ�	�F�3��N �G�)+��?�P(�$�OܓO�ʓ�?q���\-�q횁0P�vH�Wv�m@��?����?�-O��o�
pM*%�	��.U����j�#��)Dǆ�a� ��?�&^������!L<�Ѐ˶p��@���ϙ�V ��~~b�	�3�e�i�����	��'�W�+�|��M�b�N4��%�S���'��'�����3
�� ��H��)g|�#7��ȟ,�ٴyt��?A��i�"�|�w�.l�C����q�̍�b�YC�'26��ܦz�4�\:�4�y��'��p)f��tv��t�d�e�C>v��R�H߅�����OV��OX�d�O��\�x]�m���
����d!���P����)$w���,&?�I&c��ч!Fu�؁9"��~hn�I(O���h�"�'����lJD�>h'.� �D=r�FA�u�ԸO�6m�wyb
Қ��m�����D�>D��$-l��ى��?B�|���O��$�O*�4���C@�V�ǷS��/�p�r���<U�N�bd�Ü�y�&s���0�-OJ��c�:�lڥw0�x�fO~�\܁��P5k�BC������'0����M�J~��� ���V�R�&&+2
]R����?9��?���?!���OW��Iq��*a�NŃe���.�A�'#R�'�6�B"�)�OxnZ~�I�:oJ�(M��)K:P`�����]�I��@�i>�r�Ϧ-�'>��(e�_���J�哶M�-�#��������D\�'��i>1��ݟ��I�7�칷'	$Z5�*���40��Ο�'�R6ǇI~���O����|j��'�i��L|�9�V(K~���<!��?H>�O���J ^����ѓ72hx���>
�`	H0.Z	F��i>ћ��'/E'��0��6IK �J��L����!�ٟx�I������擖6���Iy��f�R�aU#���p�0#�&dQ�
I	@4f�$�O��l�Ɵ$�����>Is�i���F�7f�d�q���l�p8��yӦ�$�� *�6�q����]ȚA�Q�O���`ƹ�U�\:Rq���d�.�]͓����O����O����OJ�$�|:3��%P��LbD#'�2��$��DIN�ݘ��'��O����'C�$p���_2L��1��	B�a�kS
�5o�> o��M����4��	�OV4k�y���ɹ���P��#7�F9)0"Φ*��<bR��O�lI>i*O�	�O��/�P�)N6"]��zV�W<2����O����O0�LV�&�G.Q��'^��>=�8�3�M=y� }A�'޺��O4A�'�2�'�Ot� ���m�9Y"잩��cԝ��s�@-eK�lZ���'Vɜ�	���q�h�_�*��V�4P��r���ҟ��	�����4E���'ߔq����8ެ�U������1�'9�7��"?�����Oz�oZM�Ӽ�Ҡg\�}3�D
�VA"}8q���<q��?y�is��¸iH�I+ �>�  ӟ� f�U���
[�ѴK�D�gA?��<����?���?���?��hʨW1d�QD����Â�H��d�ܦ�h�ן�	��$?�	�{�Y'�+/y��T&���PX��O�}m���?I<�|:�!�1�`dD l�ޡ	&IͦFv���	���d�$(���E�8�O
ʓe�J=�U��W�<h9�O�&G���{���?q���?y��|�,O�=o�	��=�I*~���çV�P �l�wT6V���	�M��b�>����?Yտi�t�z��N�T� �ň�;�؄�E!� tϛ����cSf�����:����p�wIßWR⽐��ҍ1l4Ɋ�'��'�"�'2�'���ec��������m��@Q*�Ѐ	�<������^���d�'��6� ��_+xb��
�C�<8�<}�2n4:���&���ڴћ�O����b�i��I�V"���"斃2��]�7C�VeX͘�#�;-f��+���<����?!���?Dm£S�6��ro��F�����R��?�����$�צ̀����<����O����&j�
�(���6���Oj��'K46-��IkN<�O� ��c���*�n�{cC�9�Y���<v=� �i;���| k���$����cܤ��W�P��L�3�ޟ,��˟�����b>��' �7��
t7*�HA�g~��Qu�N:�\��e#�Ob��Ԧ��?m�>q��i���{w��/ ��Pˉ�$bEz�l~�HTm�z2�x���U� ����?��'�T�ץ�>b�ظ�0$�*��8Q�'Y�Пl�����I��p��d�$@ڶ����|a�� ��8-�7�K�A��d�O�D!�9O�nz�� [=9B��	ufް	2�RAɁ�?��4�?�O�O���Q�i�dO0_*S#�R+Ov��� �<^���1>�f���D��Ol��|��%�:x�w'�3*�j���y
����?���?�.O�m5H����I����ɇOk�
?���r�ݑ}U�����j}B�'���=�d7+�J�*r��9"����f��X��OF��j�vRQ��`�<	�':'��$�?���X7F���a�5�\��,@)�?���?�����l"!L�j�fa�a$�%�l[�ԟ��46N�����?�%�i��O��<k"����I�>h|� (Ѭ|��$��1����M�r����M��Ox�jh���&�W�05v-sC��s�e[��ȾN,�O�˓�?����?i���?��
�j\0�T�*��\��;s����DO��y���xy��'P��|ꂈ]�o)td UC�K�t���oy��'|J~�5 �"G��r�*�b\40`�4+�T��q�;���ş'в$�e�^�O��Z�f$ӃbJ `���W�js�a����?I��?���|�*O��n����'	ش#�/�]cࡑ���:�0��'�7-,�ɼ��$C������M��#]B�&T
�΁Z���5K ���4��$�.�.����UD���0�.�:��1�`H ~5�A����-e��O����O����O���-�ӰxV2�R�h]90_N���җD�f��韸��4�M[����|*��A��|��Ǯn;�8:���1a��XHtKB�	xO�im��MK�'+���4�yr�'z�`�B�ʌ�↏+R ��sG��I�('�'�ɟ���۟h���
���ŋ�=R9�׎N3B����̟��'�d7틵[n���O��d�|�ˇw��т�'s����~~�+�>���i^27�y�)���˃X�D���M43�̚�k��)?=��NV��M#�R��t���,�d���RX�U��$�Q1
�"sK����OV���O��i�<a�i3�Q���v�~Y�PJ��T�qH>{�"�'L�6�9��+����OD '�ߜg��M2�a�)-��S�b�O��mZ���oZQ~b/Χ}�"���W�	S--�tI���?O�2T0t@4 �$�<���?���?i��?�+�캥
���|I�����mE�a��Z�	ß<$?��I9�Mϻ��,�5m$l�����z{J�� �'қ�-��O����O��$�6�i:���`8�(�B-)f2�8�������&):غ�1騒O<��|���}?:�a���V)��AUc�q_�����?����?�/O` m�&#�P�������iʸ�wF�n���Ɗ&͆��?��Q�������L<a�j���m��,Y��S����-)p�U�[���|�P�O�h��krݙ'�҄)D	�qhZs��+��?��?9����zxx�¸U��;nr���`�������юH�y���M���3�?���?����4��N��Q�&<��V	p�n �1H8w��d^Ӧ8�4�?�B �<�M��'U�X	A�ơ���r���t��}�P�T�M�;��%ƙ|]��S��P����,���@��� ��� �.�.NCǃnyR�n�䨠�Ǽ<����3_�?���.��ZV�9:~�,ڲȕ63o�$�)O��m�>�MK���h�R���*
�5��EI<yP�!��fP��3����#�� ��f@�	Cy��)�^ų/�:��ƭ^M�R�'��'w�*�O�剿�M;ū�&�?9�\r��0a�EVb!�ٓ���?���?).OL��>?���MK�uPځ;'���-&�5�ė7p|@� \��M3�'���hȦ��S���������u�Cm�0Ud�ɧ������O��D�O����O��D3���T�,��@�t3@�'V:���j���I<�M#g@'��dR���Iyy�	DFN��e� �D
G���rT��A�4:��O�\	%�iU���0� �E���].%�LP�B�<Dݞ�)����?���$���<ͧ�?Q���?�2�Z���(���Ew衸!L�'�?Q���?I�h��tZ�tHB�?���?ֳ��4��-������fS���r#)��${}r�'�BJ?�4���d�� 4����o>Z	i���0&_��+@��/_�6MMyy�O�z����Z���hh�
KV�:p둿A��#��?)���?��S�'��D��y����H@bրX�m�8ڇ���]������ߴ��'��#���m0a�� �h���b�.P�6ML��dMRܦ��'g��#��T:+OXu#�l�AE�K�)�a��D��9O���?����?A��?I����i)pG��]F8�SB\3��mrFzӐaX���O@���O�����I���3lJ�xz�nB7:�ި+�� kU���4?n��.��Ɏ�o�6�k���G���.����W@&GnH4�d�d���'	~1�� �Ĭ<)��?�q�%SkX�%��L�&F�B��?���?	����$Zצ��$�\qy��';��څb�$��PC��H�L�X����a}�@q�p5m����a7�1���9�B�&V�_�|�'v���G�<Nw��D1����~2�'��"Td�"�a+�ߞ?���a�'R��'"�'��>U�ɎnK�8��EqOF���b�$��	��M+eh�(�?���l����4��i�E�8t��c�I\� 1�Z0=O^��O��n�[�T�m�<���t�"�HR��t��A��7;5ąR�#
M��R%�D.�䓈�4�~�d�O��d�O��d�vC������/!=��
��{T�q��vW��'�B���'Sޔ1B�ҏOv@9E�7 ��A�˩>���y�x��tb�<����M�`��@��i�b���*F)�]����'��%���'��I{3L06�ꉹ$��[߆�{
�f����/'��FS�b�p��Fe^�Ie.�9l�b�<�p��OJ���O�lnZ%._D-R�a�3miu���!>4*숡�\Ҧ�'������V:L~��;q,V%��E���id%�l ̓��?�� �P݌�9s��(�	2"�!�?��?�#�i6��������%���W#�"	���Rk��^e�<3s��?������l��i9�6�#?���\&􌀹�Ɏ?9���b� ES�չRO���$�T�'7�O����J7�1X1�\��RY���!�MóF��?����?-�v�ZQH�D�]�6`���P,h`�����O�)l��M�ґxʟLl׃�n�,�X +� ݖX�eĆ=���z��%����I�f?L>	4n��	�~x�f�4'�5��U<qU�iw\� �WT���R��.�^�q����b�'��7�6�	���}�j��q��%֦��F��E?�8����ڴjL�%�ش���ДL֔���O%�ɖK��Dd�w ���P�@�o���qy��',hHCW�őA{��Z�/N�ƨH6@`ӊ�� ��O����OJ�?=����!hC�����Ř"<��E.^���Kt�4�%�b>��D�Φ��>��Ö���"b�Q��K�73d�Γn��Xp1����$���''��'��DO�"A�T=��,)�Fu�5�'�r�'��X��cڴ3�FL,O�$"�e��)M(><��n��54⟤9�O@`nZ*�M����d��&V)1���8-�(�n:?\��O΍c�I8�j�;�����S�q>��ܟ�i�E�@�6��G�P�r�(D
џT���X��ş�E�D�'�.)��D� l	�184��/����f�'fh7-�!�"�2��&�4�iSte�e���q�F���$Q�<O�|mZ��Mk��)\�Ѫ۴�����(a��IW��#π'[�0mj�\�X�
(���<ͧ�?	���?���?�t葓�(I��m�(*�>9Cb�&��dO��135�<��ȟx%?�	�R舩Bl��9-
�p�L���p�O��m�3�M+���O}�T�'�4ER�
RL�0�#�/p�3��::p= �O0�F�ȝ�?� d*��<	��V%U[ذ�c':x6,�z�� �?���?	��?�'������
�,�П KtHI,N�����r(,Ui��K��y2�w��⟄�OPnZ�M;�Q�����ΌXg��H2�K�l��+2���M;�O��л�b��d�wm�@Rq�ÛGd�yP��s�x̋�'���'�r�'q��'�p郷*"r����C�
�"��0��O����Oj�nZ:i;d��'�87M&�dB�&���F�*{�Y�n�&Zv&0'�X�I�p���C��oZ�<�����H
BWܨ=KČ�~�R����'Gt���3�䓥�$�O����O����J��pK�d8�26M�5TT��O�ʓVY�&ň.`TR�'�BX>9$�$�KEj��VXXJwC8jO�I����O���~�i>q�	�}-h��/ޏ2�`�j��I��I�w��B��*3�Lyy�O���I62��'NJE ����G��y#�%�l�4pv�'�b�'k���Ot�I��M�i���@%�iQ�hk+[�Z�J{��?�6�ih�Ob��'��7�� x�tC�OR5���z0k؈q��	��m��!�ߦ��'z�IÇ��?��X���Iq�|\�UgM�e@!�wDj���'�"�']��'"�'W�+{�ra86�R��-���kR����4��Q����?����'�?���y�nJ))2a���Ue��Y�(X32
��'ETO1�8d�o`�`�)� ��zW�@=w�P��1
� &/t��v5O
��%�W>�?I�b7���<�'�?�rE��:�$���ab�HpC�ϖ�?���?���������g/Mϟ ��ݟ B�
D�8�2U�����&��e�D
a��]��I���	<��(�вg�&pzi�h-z��!͓�?� '_@�"��4��?mzF�O��d�#^#�T	��P�i1��Ir�@)	��$�O��D�O��4�'�?i�II)h@�ͪ���j�P[ ď=�?�g�i�X�R �'��w����]!�
�`2�˔ �>�{�B�+'�牖�M��i��6M��Z6-*?�熟�rVF�H�Z�qfa��كL��J�X%$�̕'��'��'[�'�h�RY�](�!`A����)6�前�M�3�'T�LB��?��'U3�ub���?a1e�7l$�e	�m4	��0�f��ZW�I �M�s�'������O�����$\m�K�鄉9���I��� ����>��	'qLl���'��x&�h�'��:����`���l�5�BL��]���I����i>e�'��6�\1C^����GŲ�KPƃ� O��aBoRJJ����e�?��^�<��ԟ��ش`Cv�3���B������N5*8h$)�I��M��O������Ĝ�4�wR�}�6��<�)�f�t��p �'2��'xR�'KR�'�,)���J�eI`�g�U6)�P��B�O��$�O �o�{�R�'ic��|�hW�J��Yp�(M1v�ۃ�tO��l��MϧCq�](�4��$ѮW�BDõ�")$��6Łm�T�j� 4�~��|�S�h��ϟ,�I`�D����<��%��	�NZ�	[y҂f���	d��O��d�O�	��T�X�GF.n�F<���XŐ��&��s�O��D�O`�&�������dʛ�[�m"�F��6�P!���U&M�=X%�æY�-O6����~�|"��R�H��/��a'
��T�_�x��b�6(��E�3a��Q����H���aM�P^����O�lm�b�_z��2�M;�o�L�ED�<s�����)ڌs���M~Ӥ,�¬d���l�MUİ?Q�'�����R-\D�a��+J�:"͇�O� �bćO�(q A�5��Z��W'thP�b��:D��ς�[�h,�PɊ*(J��g$�8;
�l�w�	9���"bE�/vR:�cȍk��(�
�%6qhiB�5!9��X��v��S��qo�=d�\$�GA49�"e� k�Y펍�FN@�l8,�3r�U��N�1�m�3x�,�j�B>-�r����4?&� ���"L)��$�n������6ዲA��a��A�>v]@1��>7<�P'�z<�=7�N�H%��B�O<��pdj�,N
$���y���ON�d��`4�'=� ;��Dk��AzF( ��^��)شNRXy������OCB�UF��l!��Zs*�eΘ�f�"7��O����O��R�l�d}�]���	B?1W�J���������ئe'�,3�l�ħ�?���?�R�Y�ک�`�R�lxzq
�B�,]��6�'jD�a�>�-O�D&���h ���ԋojfZ6�(m�4�FT��i4/��\�'��'�bU��p�H ]���D�#��ɀc�l�&��O2��?�L>!���?y2�E��8u��!`A��h��ɷC�X�<����?!�������ΧYX�I+�F��}��(aa�A��n�{yr�'��'#b�'Ĝ �%�O�TD�H)R�2�h�B�%|�z��X�P������TyBcX�EZꧫ?Dm�<$��]�a���9���	4i���'�'7��'�������
�W�X���'��X����r�Q�x���'z[��Z !�����O��$���3��S>j;D�U��m��D%�r�	۟\�	���q�?)�O֘�i�+M���q�+K��Hڴ���Ȕya�Qmɟ��I�\�ӂ���ƪ������>�$hx%�S�V�6��v�i���'�h�ß'��'��>���@3J00qMc8��I����TL���M���?Y����P�t�'��a��a
�+������7�"@YQm|��-�QE2��F���?)0
0n��}���R�ȡaG� fٛ�'tR�'�L@@�>�+O��䤟���JO�bE� �-g2�,��%:��7�Th%��������I�*���cH�5��¦
��dj޴�?i�'�5��	gy��'Hɧ5��_,�$��ɑd8L9%M��dS���O
���OJ�D�<)��A�dR$�I��
�V��Q�ֆ�"5�U���'�"�|b�'���$c�T����&`d���J{�d�u�|��'��'��2]�q��O�.ə@�_?�h��Y����O����O|�O��x��h��,Ԭ�G.�	{`Ґb�E<,�1P���	ޟ��IHy���2�J��+)S*>�>�3��צQڶ�j����e�	G�cyB ���b�~�ֻ���)� \`�:$h������ԟ �'��p��=�I�O����Br���7a�Ј�b���z���x_�p�	���'?�i��ːJU�lA�(��!ļJ8y@�v�P˓ZTQ��i`맡?�����I�ru��;�"��XXP1C�Х'�27��<���?і������4-!6�:Պ\Lx)ʤ���%n�,w�Xy1۴�?����?��'[e����&=���u��TD�S��6��L����O�����<y��$�NP:6��<��-K����X״i���'"m���O�I�O �	%�h�c-^�bt%ҧ��	�@7�O�˓<�iq���䓔?��9�������A"�byX�!�vӔ�D �I��L���P��`M���FS�f�T4¤FD�K�MC�Y��z�ܙJ��c���IRy��'��� 6�Zg�u���G��&U"��@H�(��D�O���+�I֟p�I#%����c���hTxn�%}<��FR3@).b�p�IyB�' Ƒ�Pڟ�$����	)��9���N�|�J�i���'�Ov���O���a��G6�6��	`�@�����U��Hbcj����?-OL��Ư`���'�?	��Vf�p*�Ƕ\H.]��G�WK�����O��DHH֌�B��x�e�@��񐲧��"Oʱ�$���M[����O4m @�|���?��[��;8lN=�"�W�Y�M�K�I��,�I�J2����h2�~2��Ec_�� 7�wD(���n�Ŧ��'���*��}�"Y�O���OA��C�l}Y���4v\$x�f�Ϝ_d%l�m~���?�������4F|<���ϫ1� �@ōDy�b�oڥ�VPcݴ�?)��?��'����\cNpu[BĲg²��3gՏ#H����4O�1���?����?��'�� Zb.�29�PE���Y� ��К��ǁ�MC��?��.-�x'�x�O��O��q&�P(������V���8`�i�rR��H�GHʟ<'���IX?A�M��;�f4�?W	X0��ͦ��ɪ2T��'l�'��'3�{A��kȼ�F)�J��e�$�d��L��	ğ���ϟ,�'��Z��|�҅+4��U1���7O���O�Ĳ<!����Į�.]*� bԨzL�-ڇ�P	�M������O���O\ʓ�Bj�0��)��O\�[��c���J��!P���Iß\��Hy��'��ßt�n��*
ι�r�����KD$������O��d�O��~�x�cR?��ɒ*����ׅHmH}p�#N&Ei�$��4�?!(O0��O��d�����3}�Ï&┓�(NLGV�@ ɝ�M���?�)O��r�G�S��':��Oj����M��t�r��Uw��q��>1��?��R		�����Tg��	��lڀM��j��RŬ�?�M[(O���Dꦉ����h���?aS�O�.�4CW���ФZ�`�f�/�v�'��G��y��|b��uQt���M����䬝�盶oFY�T7M�O(�D�Of��Aj}�Y�H���I�T 0ĊU�� ����M�g��<�����.��ȟ��jQ�s*����
#U���J�R���O����O��E�_f}�V�<��{?Q�꜄}��]�$ĕ�aGȁa�mQ䦑��}y2���yʟ.���O��Ĝ<�|Q; +�<p
v]��ɐ:Q���o���4k���$�<�����Ok�D6&����F�J|��1�AU�&�'�2��'6��'u��'�rS������o��F�1ke)4a���O˓�?�.O���O`������%��(P�1�&�&K����8O�ʓ�?���?+OR�(6@��|J�$�%\}��BO1�F�� ��I�'S�L�	ڟ`�ɥgrr��%K�\ѠE�3�bYn�JuP����i@r�'���'s��`�����$�����U�"��SB+Z-Zf�oZ���'�"�'����yb�'0�$��x� �@	8���4(�ܛ��'W���%�?��)�O*�$�7@�3���r�սwD�����l}��'���'�V���'��s���'S�b|���u&�'M�<o�mnLy��ΩiQ�7�Ov���O��)�|}Zw���E��#{Zͨ�OԨ7���4�?	��y��9ϓw��s���}*���b�����D�'��A������hfi�*�M���?����rX���'��DX��@�����tp��@�@��v���y�|��	�O���dʝ�~�f��$(�H@���U�E������ ��I�X��Of��?)�O�L�����A�c��?�8���4�?A+O�X��6O���� ��ݟH�r)�-5 ek����8�K��M��H��4��P��'�R\���i���#�)3������%jN.8���c�h��&Y��<���?Y���d�s�\���� ��$Sc���B��e��Jh}�V���IQy��'\"�'��p	���;_T�u�Ԁs3/�:W�D��?����?���?�*O�DR�Έ�|R�Cڼ$�NԀu�_'�P��sk@��i�'��S�l��ɟt�	M���	�y8 �zO��@D��	G�T�n���B޴�?9��?������Ҹ��O�Zc�b�{5����m*f,i5Px�ش�?a+Oj���O�D�<(�1��F3�U�߀g:x	*�o�<�M#��?(Ođ9�[G���'���O$<�a��3n�,9Z3L�<pbY��l�>���?���(�͓��$�O���'+�Y�I�>�j��rK82�7m�<Q"�M1�v�'���'���N�>�;n���ò�>S!J� R�n���x�ɕ_���	����O8�>}:��P�hʪ�Y���|�u��~Ӷ�3M���-�	ݟp���?)��O��9��({g$�5J�0Y`��"<�H��D�i?&L����=�S�h3��ӟ36\��D"�"߽�M����?���1#��{�R�\�'��O`�s'ƞ�(1���EDE�l��)�Ծi�2U��+��a��'�?���?y'f�:{�B=I7(=��d̾-����'�F����>�*O�$�<���[b���8����h�F-Y#��Q}r-��yRZ�T�I��L�	iyB �$s�$	elr����F�ŘB.I�h�>a,OF��<i���?��.���T�����+�/ `�����<!��?���?!����E�1-�xϧ7f��@@�'�T�2� 2,�o�Ny��'�Ο��ҟ�z��a��8�9	| 9���/Q�h<��b���$�O���O��0�ּ�Z?e��9�� � jՄC.0*���dA6o�"d�t�i�2W�|�I�4�ɀ_����v��K�[�pi����cL���$͎��'�BP���� �����O~��Nŋ#bݑi��"o�����u}��'���'Dhųʟ0����+��;���Ղ��H�*���M�.O44Y�EWȦ��������?	�O뎚�T��Q�ĭ�/B��j�ៀ����'��τ�yB�'���'q��=��%��-3z,����'$��F�i�ph�3f�����O������'%��;-�����=��K���6����4|��`��?�.O��?�Ipƌ ���/k��e�P�[��� 2۴�?���?	U�\8e��oy�'c��C�3x�f�A�$� ��Qd�"CR���|�(�yʟ���O����Uڨy��8Uj�{1� Q@(m۟ B �J3���<I���$�Ok,=�i�Ѧ��A��h �#�-�	~���	؟���ߟx�	Ꞔ�':�t��(�2 �@��VS�E?*s�O&���OĒO$���O�42��T�v�y�SY4�m)�g�J�L�O��d�O�Ĩ<�U��+�	�	�z8�/�t��\�KW:z���� ��a���$��y�p��Zh*B�ο\��:���U'���'r��'��]�܈�����ħ�\D�F�{�B%sPf�	"t$��i\r�|��']���yR�>1�ґ^^<��Y�J2�hXb�����I؟$�'�R �Շ(�	�O2���IR�%3�D����|��BT�*�Ĩ$�p��蟸Q�D���$���'H�J-1V��6	����2Ryliy��� j�7M�G���'��$I;?!�G@"d�� ��&J����,ɦ�I؟�u�ߟ�'���}rW����CsI�#��(�����R'��M��?�����xr�'��,����%,����#Y(��Ox��(�%6��F�'�?yPO�uKl��c�8B� i�rb��)ћ��'R�'�b�Q�J:�	����]�z �`��P��&���%�0��>���Qa��?���?� X	?\�{��'f�@��Њ	�ݛ��'O�8�D�4��˟��'8Zc��h�	X;�x���? �-��OQ�#��Ob�$�Oʓa{n�"�Y29��`�7e��Ey���Ƌ�]!�'�2�'��'�"�'+�-�W��Sq���1�~u��+ˊ�y�P���I���ICy'�XS��R�Yz@�оp"�c%n�"SӒO"�d>���O ��*!����8<����㊪/��!�r#�}����'P2�'��]���'C߉��'n���pd�α �|ס?ހ�Ҹi��|"�'����u��>�1͛b`y�.�*�����m��ş��'Q�U�f�(�)�O�ə�'��EؠQ��)�:
�=	�i;��O��������;���?sAb�1���1��MG�P�ՠm�Jʓ>7ȼ`��i8���?i�':i�I�kE��g�+Do�m��">z�6��O.�dҾ0P�/��-�S���"�_�l�"��S�P;N7
6G�kS��oZ��I͟@�S����|��	b�=2��n�R���[���N]<a��'��)�'�?�"�ׇ� D!��°�B�I�7AN���'���'���ꦦ)�4���'O8h c�d�zdA�@ѝ�ҥi�4�?�)O�e�ЈFS��۟0�	ßl �+����	S��R����Ѩ.�M�%�\���x�OkQ�P�3%�1Tt9��D�g���0��>��
<�?q��?1��?�����d�?;�8�i	/us�U8b$D�8i9�cSs�	ޟtG{��' ^l��I��:���cG <�b�8�G<���'��'�"�'���	_A��O�|��AɅ*p"�u&Ǒ+�A��O���(ړ�?Y�-б�?釣ÃYX�TC��wu��"R�I�����ꟴ���`hU$S����	ʟ��B,Q���1��3&�pK����M������?���)��m�1��q�4mMR�p�O*">�XT�3y�J6M�O��Ģ<��ڶR*�S����	�?�Ig�<Z����C_�Q�*х���M���lR�5��On���^	��7��Q��ZF�f]���i���'��`�'���'k2�O��i�q�T��hU���L�(趭S�j�H���O�<��	
51O���y෫�(^�,u��ǟ�Z`���iM| E�'u��'4��O�B�',��]��P���������
���P��4d�N�:��O�S�O��߄մuQW�2.$�������6��O���OTM`��BB�i>)�	����F"�1d�#���v���GM����'J��y2�'��'�V|2GC�<7|��W��#T���lp����ԮH�N�f�����&���P�T�}�(Q��A�>K4���,����Dr�Yv����	�����qy��_l��(Bâ	����D�ڕ�� ��g)���O���-���O���I�I3p��f4N,5#fO5j������O��D�OT�4�
a�5:�������t�hD���&�%����ē�?�N>A��?�2�L}�,����S(.x�Uf���$�O�$�O�˓H�yJ��TF&%&��4���)�:Y�	��u�\7��O �O����O樨��đ�}��@���24�e�ݔ)����' �P�X�m���'�?���u�Q�� �0$���b��nR����x��'����O�$���Ϻ@-2��ӣK.	��7��<���M�g^�6;~����ѕ�� �� 3�T~��kQ�(>�%�F�ia��'c\�ʌ��)�2h�.x�5�F3P��#�^.��h��G�7��O����O����|�H�(���e+, �8�d��q$�q�i��-���d.�S؟���AM:/w$�4G�8!����u�&�Mk��?��a���S�D�O����^6�=צ��4/\����% $c�dCU�#��۟��	���pgi1oZ��Q�_0��m�j���M+� -���Q�$�OT�Ok�$[� ���,G5!4�8���&���S1�c���I֟���ayb��/~*��$ �u�؂ G�49ָ�7�"�D�O��d<�d�O��$�- )X�ýB)�&�8��ԫ����'���'""[�h#�OP����$,��p���kS���o2��d�O�d*�D�O�җc��I+.���
z�x�D\?O28��?9���?�)O�ԘQ��\���'.���G�(��k1��>,s���E/vӾ��<����?���;p��?��'`8&H	�+A��r&L,si�Cڴ�?������ſ�\ �O>�'��dm���7��"=V�$f;kB��?����?�efD@~RU���86:p�s$Ftb4�Ii͵�J�oGy����HԨ7��O(��O����u}Zw%�,0''¬�ҥ��#@�][hEp�4�?��[�:1̓
.�s���}*�-�=K\\�C'K�:����G*����T�K��Mc���?A��j'^�L�'��iNڝQ�ˇJ�!Ȃy���hӴ@g8OR�$�<��D�'���$��1z ��+�+���Ƅe���D�Ox�d�R�h��'1�ğ��ZZ����]PN��"h��% \�>���ZS��?1���?�g�ȦJ� �b�/����Eʵf��F�'d>i��>�)O
���<�������Qh��A^,2���E�CO}������O����O���<a�%�oն���C[���H�^�H�1a]���'�RS���	�����kL���)J�:dG�Ύ�Ь�g�$�	Ɵ�IߟX�	By���4è�.?^l�s�ٿR�}��B�4I(�6��<�����O��D�O�٠�:O`�h�F�,+JH�5K��Y��&Sj}��'UB�'��I8�d�í� �d>?���Ђ�N�$�"�`���">��n�ʟ��'�'*r'Ʃ�yrP>7-Mg��xR� z�0���`+(D��fU���)T��I�@,X�#�Tu����%z��ɬf5btH�� ��TC�I g���c J.�R���_$�˗�QV�X]���u�X�E�GȂ�_J�A���N��!��V�d�T�[䇗#8pX����.�|���A�Hܠ�#@ ˲�B�I�f�<n��d*���9�|�`��B^#'I�\��Ic�b��H'�����#����8 �7E�Q�pP�Q� 0�,YB�c��
Sd��O����Oɬ;/�<��FS���\����*y(���GI�����Θ-��x�ba����O�f�'��q� -�NRQX��Z��Hұ�/+� ���4�����9�.��3J�|�0 X��4�ݴr��B ��1W����B:����a~b,��?�'�hOR�㧣�-Q�|�q��.o@�8A"O����������,X]r��<���?і'�,�Z����,Y6�ې́�{-��6Lٙas&mʒ�'�B�'���`�a������'Mn�2ӊ��W�|er���p��+����X�Hvl>`9@9ϓ,��$�e��d0q��"Q��x�V�X?V xC�	`�+�[<VP��m~�cA��-Jq��)��̟���r�'��O�%`�,ι(Tܰ�B׸X�0hA"O���sM3%B6�{3B'N�F��e}�_�tB�	����$�O����4��Ei₄0'�mz���O����1X.j�D�O�擠 ����`)7�V�s�'82�Q�j��H|�� ��ݕs|���	Ǔa��U0���DwTu���O��I�Aj��0�#Rȴ]���'%�!���?A/O��6�� 8D��r���&�4����'|OTmˤ쑖�XJ��<5�L��eO��lڗ@@�l2�F�V'����F`R �`y¯Z B���?�(��Xy��O��� ł
Mx|��",ߝ3
i���O����;� aH cX#hX��O�a��i�#_�Ԓt��*��� C����	�V!L]�BdY H�ra�Gn��?Y8���Qp\T��I;z;����>}�K��?���h� ��&BJdf�N�GK���Ь�:)�!���(<�H�+�:f����e���axR�5ғO?��ې�~�dq R�V��.���[�����<A��ˡT<�-�I����I͟�ݓn�b����(T � �3Wy����O%�I�2DL�@�)�3�$���`:��(%$�RS�|��Hq�=3}@�!q� 1E������]��剶H\���#��E�Ä8�̡��q~R���?�'�hON%�MX�G"�x��3 1��"O>LrwD�Ce0@�F���h�F<ّ���{���?�'����u��3�2苰�D�����/��~�� 2c�'���'��y���	��d�'�"J����n$Jt�@�$_��N׹4�����Ј
�H�Dy^}�Q,�w�
)�$�� �`����`X@7iÞJ�[t+T%jx�Q�ɘğd��)� ��)��E�vo�!�$�'[��$e"O}��M0I8�r��;B^�b�dD�]�,+�i�B�'�R��`�~'V���O�t�z�B�'�m��A �'��H��|r$Q�?RB�*T�T�	Ɗ�����p<1G-]D�YR��(���9���Z,xv���S�x1��[�	���bG�T�K����D��JC�I*�@k�Iy{�����$3�2C����M�"Q+� �$m͐l����,���VW���i��'�哐88��	 /���1DG�z��M��`ӟ|R�)�	ǟ<��ԍfvE�$�����|�+�A[����L�����1��>���NA�ab`�v����'I3$�Hf��s��$��ؠT���'�P1i�ɘ��O=�QT�(���#�B��U����'��@%����C��y���Ó�X��Wm���v(�x��릋��M��?��S!T�q怯�?���?��Ӽ�-�[rlV�r������+0z�
P�;O���Ӻ	������|�O�H��:d�ñDЪ%
��*�x����z���̶lƠ骋�L>�2b
�c8̝���ŠN���c�$��'���S�g�I�#4�� T4)/$Tp�A��8B�	/p*�s7��;9�X]�6B���@����"|2 O:NF�;B�Y?y�Bx��`�9�Ys'�;�?q���?��M���OH��v>1��R�O+ - N߶j�.�PĬ���C��'xGXD�q��MN��6dH�L#l*�)�X�q�]�}Рq"�ˠ9,��&݋<���(�O��8���:.���@ړP�Z-s�"O��P1�EL��b4H�Z��0�q�Ni�(}�C�ivB�'�ֈB풴	�>P���R5K�x�@�'���ոlw��'��	Z�?b�|�e�.mB���%�NQhG��p<1��O��FB!;c�?cY�9�&�ӓB�@�㉍����9�Dİ?�<����J��M!�>]�!�D:{\Pc1�ϸA�F,*���6!�!���q��M�<D�x}��O!9P��N&�I&l���4�?����)�2����"A0���Ơ�2�P�s�P2�d�O�%���O�b��g~"�UJ��qR2�ʮ���$呐��m{�"<����kLLc�{��yY��T�DF6a�'��O��O�ư@��^�p/�\A�%Ä9gTH2�y��'k�y��I�z�JQ�X
��Ց!���0<�!��c��@q��A�F�)�$"�z�8޴�?Y���?9R/��cv�I���?����?�;un)!�o�7<,�[��֓!TB�Z�y�ۈ��<	�l�r\䀐F�[!^R�b�fܓ)��9�牔1@"`:�m>�x3��[�(�0��<	��[��>�O��t'�'*�05�� ë)����"O��9����U8�i�¨_76d������(���Ӕn9��Z�)³g��MgƒM����޹8m"�	ʟ��I՟�R_w�R�' �i�L���Ѷ���C����D'@FHGL����$M�{ r�
$�V'Y�jCk��]��"�ɦa���䉦aEn��� `�:��B�T-~��Ȉ2�'���'�B[��	y�s����&C�?ynv\�'g�4�<���e���@%L"h�{k�3k���<��T� �'Uf�#V�iӺ���O���*3i�Ջ�#P6���h#E�O���Fc9�$�O$�ӻ�A���
&�pa�'
1q3i�y��h�`D `8��z
�z>5;����"�e�%�O��K4`��$R@���;�-@T�'�z�h����	Fd]��a>��L0�>����(?
� ���|�ԡ��ϒ)oYn����W���,U�@�j h��)�'ǘ'��\p�	zӎ�$�O�ʧ1a�82�"��7��Q��y�R�J>HI�����?�UL���?��y*��	0\��5���,���#Q�ܫW���'\�b���	\���B2d�c�����>1��A�S��_�<� D���4-��_�2ͬ ��X�{�!.N^�B�I��l+>Y��	<�HOf�Z��\���RC�1HR��a��Q�	ܟ��ɅA,(,���O՟ ��Ɵ�i�{Em^DJ4�R@�L�P��D����a.M�q1�$���;��L>���>;Jxp��N�U���Ş�g���PE��A�4XYEEöc] ��}&����Bҙ&$�G�C�[������g�X����)�3���	S�ap�a�F/:�q�n�!�� �m�ʮ����7d�	�ɲ��02��4�4�O*�ǧ�W�����D��� �+&A8v�ˢ��O����O2��ݺ3��?1�O��h8BEܕ^6�tpa��`=�T"��x2�ю�����R@`Kօ��`yT9�'��Z�OY.|%j�e��5�;�I���?��SDV���Cr�je���P/����ȓ3�N��`ۼ!�XMbD#07�b��<���DU��(oZٟT�I+q��(�AȤ5�aI#�$zd��Ɵ���%�ԟd�I�|ʳ�e57M*����BL�rD]qyq��*R�&�xB�
��'��ms�lX�<��R��%�����b��h�Iz�ɮ(� "S�[�d_��P�-�-?
B�	�I��fI7�fX3�舲u��C�� �M�qb�-h�x���@H�@5#�v̓;ݞl +O����|�5$�6�?�q���5P�1�P�ũ@i�%�W����?Y�g� S��ԋj]V���kEN?�O��s�E2��H�Yi8�ѧ��<?"�'��C @�,M1����`�O@�<���Z!����U�<��2�.}'�?9V�i��"}��'2�$49��� �pțE*U�1�'M����ő�}�呫;ռ�s	ÓPq��H�� $X�P�:Ec� iX΀�)��M����?��,lSa�&�?����?A�i��T��и���	��ᓠ��Jc���P&*<O0�2LC ���E�n0¨9B���,.�yR�_��Y���O�5��JO�/$1O�%�������6pȒ@�9`�*����(RrT�� V�X����'�P�i�؍{�8��'�<"=E���W{�l.��S*�5^a���p@V1u~���'�"�'�a�i�I��̧z��y��U�\�n�W�N�'m��g�@F<A3�?>����gO�M�i@����m���=���3$CR�t9P�R4�I)x�X}�A ��P��	/��8��L]:��Y�ćК��C��f���BGU)"�x#7K �bc��؈}�
L$O?46M�O������F�X�����A�(|�n���Ox4���O���j>���O�OH5��a�d��Ñ�׵o{n0���'[L[�B�?e�<c1FQ��*	�c@�
�p<�`��ٟ�&�$��X��0� 4A���r�3D�|��"\9J�P�{UNۥ!3D #e�0��ܴ%4�Q�L�'A\={�M� ��<7�@L����'*�\>�sc�џ`�4��1��@�(��f��]c�!Kş8�	�x��	
Ŋ����S�d]>�����"Y����҉�4l&}"�/Hf��P�|��4��t�j�N�d/���iԶ��ɾ���Oj���O��?�����bd��XDa�?l�1�C$�I�����I�aͰ���F	^���
���[�p���@a�'Ͼ�Ru锋@��I�%焬B>��(��{�$���OH��)�.4�J�O�D�O��4�L	����,�1s�� k6��#��4�	�QU(I
��'���&�?@I��1�L�"8� �{�ߑ))J͆�	�O�(�Z��NmaV��"U���IG~��3�?�}�I�����+�\Â�
�<qqd�/�>y��/�4;�HM�i����5e��H7�,�����D�O��<�r))�U��
�!��|蚈�4�'5���ת��as!��DkҵA���6���9���+�!�$+��DB��+�L�b��	~�!�D�?\|J��2�Th�B�ʢr�!�dJ�Iܱ�!
�����C�۳!��R	GN�$�R��6��@%��7r!��'ef�X�hj�j��K�ei!�d�q�T��oҠeV�{�˵sM!�D�K 2�B�����R%��,;!�d� A�Bd*C���W�,�+��Q�/!��J�xe��j��ǋ�\�Ze�BY!�(X��%aѓT���	�j�-�!�ܦb��t����&2`�z4$�{�!���tB�A�(�h���3����P�!��>6P��:��'9���Y� �<�!��̭;���+��[���a `�9u�!��  �+��/|	b�#��:����"O�h�Ă%LJ䫅��q�z��""O�IcT>S�hYu$����U+ "O�iS�#�����8S�T:v���"O ����:?��e� �O��8��"OLxq�K�+s�b�x#_���� c"O>��FC���ءe�W�P�\� �"OD<yū̾��83c�S I��3"Of�QdK<u��jS0l��7�3D��S�i�q�n̓w-X�t��X�n1D�� `$ݘRG�����5Ya��`Gi+D����Z}R%�4�ȕ^�ț�>D��e�ћI��0b��&Y�^��b�>D�@ E�=����V%�J�dd�ѧ'D��I��9ØL���_�-Lr�1�!;D�,ڳ��7`!ND�c+߂-�>0� �$D���,a�.�{���*�P���4D��k��C�D�씻��D��b��1D�����*u&�q!����n9�Ђ0B1D�8�c�,~�Ti�4KQ�`J�9˳l0D�h�·z�>t`��0�v�(�2D�ԣ�lıx���M�
��P�'<��.�&iR����.=e��T��kK �I����}�|�'̔kJ�� �i�@�'�w�T\�A
�(9�]��';����"C^�۱#_Z i����:3���w""�'/1�0�6E�A^r��^:0��ȓ5!0��u��>SRȹ�/�9.{\�X�X/�sU�|���'FL\�	��Wl6ɩ���/t��p�
�'t�)��˅Z�"�x�
L=��R�'W>�ڔ�ƩRha{bM͞Rr����K+$ȗ�7�p> ^�C�Ty۴S%V	����a( �A�ѷP�v�ȓm�\}�O
�P�
E���k�b�Fz�c״a�.}Ï��J�����/g��M��( �!�d�5a��`�R�ܤ#�T�����!�Z�A��ip2H�Edl����l�!�D�/.J�iTӸ_O�|ѧ�N"c}!�����aZ3u���s�IT�o!�d��$�A�(�����Ƣ�)>u!�ĿN/ұj+�%|����&:k!��	B���(_������-9P!�A"P� ٪ h�R����#jG9!�$"�YX&�=�~Ah�`�7?2l�O�ștC C���H?��P���U��uk��� q��Y:d!#�Oy� kC?�:M�b�I�����	�3��K@��: ����~�����$	�����ڇf�ҭG}bg�;�Zm� �P�]�O���íP�b%�dr�˗�}T���'/\�VH�cL�)�ҡ@�8��'R��X�NC�%JF�Gr>�3@�^�n��IX^2 �3	3D��Q��7(�y6��'z�:,���"��ɱ},��Ua@j��g���y��)� ^|B���+8bU��	�\�ZxRܘ@����b�-4�*�͒ 5h<(J䯚*)�~��ǒp��`��Dy�n4;�� ��y�&3� d�� @�L`Sc%'�y�`5kq�M��?-�r\��f���y�(F�EQ��e�P��=!���?�y"HТbi��HC�+F J�ˤ��/�y"Bʋ	�8����X�o���2U!���y�+	`@ݰkɞl��r�ߕ�yR�[_F%�č`�(���M�y2�����@RhɌD,B1��V�yr��5M@�� ��=5~pɐ�`��p<yp��t���!KR�	���jqE�
����f�6�\���)B�zBڠ��'��C�oB��w� Q�Qz���>)��C��q�f�L� �%ėB�ȓ�� J��
)���Nϼo+�|���^j�<� ��� � 1s�"�+ ������y2π
r��Ђ� )���r��	��Ɂ7,A�p���p��XҐ��/^���Ă�L����+vL6�;���&=�5�"��n�R �lۏ~Lmїi�>��"x�I3���J�4�2�s�����S��@��6�|�`4�	(e�����K�q9�A�k��`��
��^�4�*�A�'"�[S�&m,�ȩ�M�韰�u*R�u��x�i�r̒ ���J	LTb�l�0�"�$y�>�{G%��*L��'d��(�R�(pс q�D��v�١$ɒV�V��,gJ�At�4��0��/Mڼ��$H%w�,�1aJW>�,�#РŻ?Ts5Ί7���2��~���1�t�3���VX��H�� ؚq�ל!��|X"�B����1o�O�����C�����!H7j�8��>&��哇ƚ:��v��>Y &�x���Cc��{u^�g�j�����'�!s���:%�%I��W�~�*я{�R1U�p��;$���j�!Q2m��Q����2cbW�G,�}�4�C$2�u�c�G8w�fd{�
�%�8eC&�H7}Fz�3gjG�����q��7>����M�j}N��1��9��q���=0����>�8�r��~=���E�*�N��'�M��l�v4z\���(�قuȈ�N�] ǣ�'n�a}���	����!�
F�D:#bX���q��d�j]r�a��H�jeH�=��	�Ϣ�7 S2.�̚R��92��AjeT
���qo�m����J��\�XggR�7/�| @�#z�v	
��J #��0R��A9��m�p?it-��^���
&�	�,{�Xw-��F�B���z�v!��cF�+2�$Q�T�~i����O�Z��ۃ�B�y�>�HY�2Ez4{��¯H���/��$:���H�=�ņ�/x���T�C��@���4ر�I
��OȤ��T�O��0�
I�;(�娤�\�|P���r�	=#h����C�jJH���D�W�2�Y�{�����e�⌨}Ҭ�� �"J��s�J�!���G����>	��Uąy���yr��`���o��Vi��&O N=c(�?��H?9���hh۷�Awϔy�"F��Yt<|1e(|OD9�A��7q�iر�Y	z�Șk�*����*����Y(��-]$L�@����R&Z�Ia+�x���B!�R��B�tLɡ]�jȰik��
��O�\�s��7\(���E!�`���'�|�Îu���y�F��$1À")���u����2(�9FLH��iך k�#=Q�l�0H��U�I�l�$U��<O�� �ix�<����j��q���O��Q�Y�,^$T
Z���Q/��4�h��C;��	d�^u��I��6��|�D�E�>���`��J�LJ�����4�Z��c����iɴ4*��*�L;�I���;���rUO]�]m92u�,�,7�O`����;��k5̄(%�Ƹ*3L]4\�:����v������9ʤ�sQn��d�h��q@K/m�+W�ɞ[�>�����P�T����h����ė�����µ}�F���l�J`qǢ2`ȭ��$�j|����Oj!r��**�"A�¯�1A�`s��	�OQR8�K�&xԔi5m�T,��
��+�b�$F)X�c�!Z�@��}��Z̓h�QB@��;@*�  ��1(�	�n	D���"�O�!���P�� CMU[��*	�>��)mI�I��eQ�;��|�2����Υj��![6�J?C�d)�"O�T��.]/5�|��)�dm�I�R�L�'���O%m��P7�W-2�H�O�2iߒ&6d�r�5ȮpY�ܵS�,kfK6�̕����%+��\�ι~j��O? @����ǀ�05��IԎNw��A���;�io�Fq0��Q1��Gz��<�)��m�<	��q�w�]1�PM!��)X�ȑp�=���,�1O����콲�a�;K�T9�(N�����	_��Gz2�+*�D/�m?�"��;gh��jCHG&z�p@�C��iR(�q�'�1O������',����w��-��̇�tA�r�3E�2b�yr�_2`��r����b�fNEa"
%k����� ��h��	W(ڰԈ���3���|R��i����v!ƖB�|pBG�P_�̴(7��,/�bm+��4���)O��A}��AJ�	8>��aש
L�0�i�:I�3	�G8���pO���	��V� ��Qɨ<��4�n�c;6�є-ô31*h2�C��_zȷ�ծ�0=ѥM�J=���bG�,����c%[�FK��I�^��QT-Wn�Iʟ��'�l$�g�y;NA�9�Y�l�1%i� E	��}!kޱ:!1O�| %cΑz�Q�)�N�d ��R��̓A�T˄�H0袤��M�H�'��������M"�o F2�1��d۶��M��CYzx��d�5v�l�4g��0%�����	��|�'s�(9�`5j��$j� V0��N��sVQ�B�^��p>)c��� paϏ3{v}"#�Uy��i>��'��٢�����Pa�ўqҎ����-3az�`�)�h����Y�0��ᄒL8&�(���(��a��U9�<9U�=oШ���݋2L�Qp��{���E��,��e�H<c�1O�a�X#0���'j�d�H>���9CT�ӷ�-0�@%bFg���p@$`Bo�B�ܓ7LU=���=1@�������W�A���8C8Q�����t*��-(`c���a8�`@�fԌ`�lQxRA�X� -���&t�F�
b�'5
WaH�(
�d�%AS*
�֝aO>�!IC
��<	#˜�%��̀`�AS��1��&S��p=q��D�/��˨On�p��]t)���C�D(It(a��'����G�T	�)c��F/�� hUsa癘y���F�]�r���'�y��T�8�� K@��+{���Q��ۯ9̅0����17d��O>1����q�d���D�<U������LhܓN�2)��"buGj98��<	Cb	C���0!�� ����$*Fg�~]�t"R/V1nz٘���mbhH���Xbub�B���IaX���
N\2��C��
��"�I�I�����c�<��t���oB�y��8w�
P)V 5� ��G�Ɂ !��J-p߶h���6wHf4��HI5y{�y��7�f5��@Y9��� ���i����b/�%��eh��b�az���2c2�ks��)��L���1&�bY9��ۼ} ⫁���=�"棑�|�a&��y���=��
P���'��>�Q/Pp� N�� H�������xy �&�����ɾf�^� �c��U-�oy��i�E+r_:�3
�S.�����7%��D�����'�J%*D��&^�@�c������S�'b��@��ނ��Dpae�S�ć�0 MCUBÍ�D=�����1�J�'��4�z�@��h��y̧h��'re�ւ��z< ykCK-&>L��'�rd�f�6�h���@�Z�N@�#�%�mQU�(O�tآq�}rz1��I!\�^��@��4o~z�8D�^�n�t����%2ܤx�׃�w�t�� �/� ��Չ0G }�t�Оaޜ���A�Px�ϙ !����9o�x��A��dW3�ޕ1􄋣l,�8�dI ����Z�6���� M�TE�<+��Y�y"F�;H?L�s'Ó7O̺�J�Н+ⴼ����7�<x����$0ܻ��ԝxB����ܵbv��2�xa�ȇ�yRɍ�X�ȱ�V�[�I[vl���y�%��r�f�8!ȗDJ�5:���4�ybfW(L�-���7@������\��yRG��aN�`k �Qan�k��P��y�c)iL>X�gǎ>,��"�IH0�y�N�<�uZ��͚"<�W��	�yҪ��WX��3`�`Ț���y���Br�T+ËL�6ʣD���y��ݶkd��9�m^.c�$P#jG��y���L�,%y����pbc���y��-�T�&�)r	9�Dʻ�y�H:��@A� Rܰ�Ԧ���yR`"KtJ|�N�,!��D ���Py"�P4v�z\˴MԌCM����t�<qg(;M�����-�}���)��Sp�<���I	/oJ����	P����J�j�<فC��	�|�
��ẔjJ^�<�E�U|��9Z'�W�!g���"�GX�<y��G�n|c�I0A��<#unFZ�<�E4�ƀI���25}�X�f$�L�<��֔<�+��G$[pă0�	A�<����i��ԩJ�Y$Yۂ�r�<1U$�@�8�����
�.�y�<A��^g���E�Ջ?��}��'�N�<����L5�P��2_��0�jFH�<����R��
��
R�ޕ���]y�<��N�/y��Ȉ˄e��p �Xr�<i�!�3Z�d<c�a��(8%Ęj�<1�.�����f�C)��y+F�g�<�����p�3�Lu��ۤc�d�<���:M��}@�
�fC��b��d�<���F�@�&��Pxl� �X�<��d�ЭPu��c�ڌ���<��$���S�Hc�Ԩ%Ør�<�w�BR��tp¢GUTv�X5h�t�<�&��:�H��ED$R�U�3�j�<�S�/o���"$n� `]���b��f�<1S��6#��]�b��������N`�<��ܺ�6ݡDؾv�����\�<���1� JPO��e[|Ų�BIr�<I)<D|�M�r�Hv��ы,l�<�T
{L�edlԾy{�J�g�<� �#�,Po�|A�Ȟ&XިE�a"Ox���)G�%PGIׂlI�"OF�xf��'|��`0� �8;��Yk�"OԠ��	�ao��� %A�pM �"ONQ�V��Rb^��� S�ް-�"O�H�f
AwH0��$���*݉W"O��ٷ)�血���48����g"OLh�A˴z^�P���R� ~@<��"O�܀�&�.�D����R8STu��"OB�ȠJ, '*S�؜�I"O�����RY'XA�#�����"O8X�5j؋R������Wj��CU"O�m�R������ԤANn1s6"O�Ͳ2J� ��	G�õ��Bf"Oh��p�2l�T<yU`ƀd���e"O��{����z��/ȥ �-��"O"��u�N#�>���\�H �,�@"Ov��2c�=�ĥ��$LI�"OL�2"���~g�	� �V�٘�"O�8ʃ��`Bf��2/��2��%"O 0�Cy���A"N�,���"O��S�u�r��Pi�OU�˴"O:��U��wk�m ��7MB�)c�"O �R�eψp|b��g�s����"O��� Ũ~n �����V�4e2"O�qq�P�>/��A L�*i�U"Oh[��F-Nx���嘸A��ec�"O6I�a�6J�< rE�6�|�G"Od�����x羼`��K,v����"O8���l�7��0��L4�ࢄ"O�h@󋌓-�,���
���aY�"O�4�FiV$�骇c�G �hp"O6�i�+T�zU�Y¦Ȇ��ι�"O.��%��(N�*�*2H��y3"O���T)�%y*��v�8+��=p�"O��x!cC0h��3�ŋ�W��!��"O�0�q�H"$6x0��I������"O\��ċ�.�`bI�^�h"O`-�
F�5� 5�V��8��"O$�K��<I����cŒ�t0�"O�	i�̀�z��ݣr�E�@�(�"O6U�GZ�r<P�E-F���()�"O�y V��y3Ȅ1�L��q�@}�%"O�,y�mO_Wƕ�f+|��!"O���m�<�HYБ�� ��)Z�"O(تe��$PWt\B���8�0X0��'��'���h��Ö
��p��N�	^@@�'��8�A�F0�aT!�0 �����dԷk�����g��-[�?W�!�Ą1)���qEȖ%sDePeJ� �!��ӽh2��:��	7Y*|��	2�!��P	)8���X�J�
��%�9N!�O 8�>ڲɛ+m�\��AL��!�D�<2��`���_��h���D�!�D��O7j���D�,�P��2EX=�!�_�T�����C�`xR�ɸ�!��&lB̈w��4�J�ƭ�!��	�y�F䂕D�5$���0�ͻo!�E�n(�����K�����-]�6O!��.�BD�[1Et�TA���r>!��8kɒ�*���0n��Tؠ�!��%)4.T
��S#nW�t`&l��F`!򤝔:4 P���An���Л>9!�K� "���	k
�!S�-!�� 
�I%CI�
�yQB�=|*��"O�-�Ql̨*6D	�n�\^�R"O(1�3ǊC�ʁk+--���R"Ot](���+��ᑯ
6�8a�x"�'��	H���D�R@���q�
�'���FN19��P��9m�%��'���@���(8�҂�@-�İ	�'�
�@!��qM%b�  l�A�'��B���<P��*⮌�'}�b�'��BaD�j*$�@�IJ0m��=�
�'��LJ�O��{�/
_���j�',�@A@AJ΅���ۋJ[��;
�'�P�(�O�S|:��m_�FΊ���'�p&cЎ>��%�g͐I��'dzu�A�8|��Dg� a����'�v��#&�yK�_�K�.��ȓ3Q��pR�r�q+b*�-Նȓb5\h8E�!>���#��Ϥ	~����EȬ���2Z��Eb�o�LM�1�ȓt���Yg�9Fj������@��ȓӆPX�똏_qYIc�Cr'�ݤO�=�J���;q�,;�8�7�T�<qw��0zP�y��+J���y z�<q�c�W�b���'�?OB��Zv�\�<i�'�;f��	�#�T'Z[�x)5eTV�<Y��*r0̄�F���"l�r$Q�<���4<0��5lޅ#=(��aZO�<���_%f�x�e$��N�ػ �Nb�<ys�̼D��x���ۓ �y�C�S^�<�C��:zl��r���1�0˄�[�<�h^.�"��""�:ڎM(�F|�<y�MY���ۀ��K	��A�'�a�<�ҠY8�����.G	U��!����d�<�pG�R��8&�ZR��j1(�U�<1f&�?@�D�E�H���VF�R�<�w�J4��,�d��<	}(�`"$K�<�V��'%����[.SP0j�o��<I�G(z���ʥ�Ȕtt|�q��u�<!���.,�l"�!�%�_>-{�B�I�}�h=B�GѨa�R�Z�읓*U�B䉅LT����#1���්[[�B�	 q��p�Ƈ�5G�c�V��F{J?+��
4D^(*�<�D"&�!D�x���8m�m3�+U P�fT;�o�R"<���O����EU�e��IjęA1�|Q"O��Cʂ!K	z�x���&1�)��'ݛ..�O4�R�+�<���C���@��3"O0T�C&J-!x�)å�ۚq�E ��,�S��ɔ;��H�D��=%�T5����Zg!���c����ݠ$d��+eX3wd!��"a�ݣ�`��d�!4ʏ�C&!�D�=�z��D�=x�j$�4j�Oԣ=%>٘Ө�J��@�%ΑV��J�a?D�Phgɏ+1N]�Q�wF4}��!1D��0�@c�v剷�S�3�H#g0D�����6;����	>�Ȉ��*�>Q��'A�S� dպX�s��`�f��'4��{3�W�`8L P�кZ$ʰs�'���G!Ⱦ`AmCR&!P������D!�f��ĉ3�;^O�� GR����ȓ�j1���(�6ܐ -�$N~�H�<ы��	S���۔�!����X�!�!M>� e���
o���q'��fd1O~��C^<����A��jd���lJ!�� n�� ˔_O�miB�-�P�t"O4=�#k��hx<�c��8`���"O$E�%o(:¨ɡ� *�@i�"O^]I�J��O�/�&j)�"Oؙ�"k�qmj=��u�����'��	J�
풠�R�|t@ɢ��<��B�I�L��r�$�4ӆ BZ+Y"����7�Ʉm�.��I[#{�L��I�B�I�4�~%�bk�z��ۣ%��"?ٌ�)��$�4C3�D('�����!�Ą,�����"��~3���'��Kx�'_�i����'��41M�&3�F��	�24��
�'�6lC!�ǂ�6X"�D>/��
�'���a*��(�L@�c��+E�2ۓ޸'M�X���]|�H2C�F'$p~ i�'B"��ġ�pT�i��/��*��'����6|�Za�֩
�H���'��a#�\}���LM!	�n���'�ў"~
ceب �ֈ��D��KQ���a!�q�<ٗlwt��"�Hx83Wϔj�<b�W�!2��`7�ir�tK�a�g�<Q�'�"-Vmp��O�XƖ���eZ}�<���y������*Q��XF%Gx�<��� 0�( S���$7�:��5��s�<a�mB�+��a�kJ 
I��@�I�<�D��"K�=��͕CJ�xǧE�<A�h..�ŉrߛ�B�K���V�<9P���a.ap��TH\���dT�<y�H�r��Č`P�b� I�<1�-2-\}�ˋ�8Lؘ!�
G�<�
#y��dc�G���O^�<�ҍ�xvP]��e�M�,���%�W�<	�&�<b��U ���
c��@Rrk�z�<��+[�~j̃�K�-#U�����q�<�3�նj�5��N�P�v$��ny�<)��L�J,���ْ=������u�<r#Թ}�$(�7�B2�E�"Y�<Q0B4\��I�V�@�VF����.�o�<	�ڿ~��,�p�S_?~u�e��<q�7W�40�LZdFF�a!n�T�<i�F���7����RTq�u�<1���-�� ��Z#'�!�&q�<qү�9	U|$�g�J	gr!!MUi�<�Gj²�b�����T�8tNO�<!�FčG'`�2�I���]��$R�<�G,9N�h1��f�z�]��o�i�<�ΟZ�aҕ��g�n��R�h�<Q�`��Z��{j�M8�cWa�<	��	 �!�% �<�z�z�e�U�<Q@ϊF���p�c��͐ۀ$y�<ɡ�&jp.�A�!F @���7aK�<C��=�h�RA¤D��`�O�J�<���&$���	�7��mP,�F�<a�,�(Zh� �s�~�-�u��K�<�$A"kAF�0f� �,�:�S�IA�<	�O�W��U���k[�u��b	y�<r(��#`d��W,��f>�I��w�<)�� <^���K/2&7��/�yr� �̸�I��Z�����h�	�y�OT�xԫ#lZ�r��&�Ӷ�y2�M2>�V4#�T,8�(��J:�yҩ
�
�ii���2G��[A�D��yr#3.f&�#���r���I�y���j��mb�߀"��CW!�5�y
� �%�чI�W��e���K!���q"O��B��!��cQ�G�,q�"Of��b�?$���m܆��d�"OqR��S+g�Y�v�N��<�7"O6�x���"�xi�!�ī|
ɉ�"Oj݀C��7p��ʕ�*g� ��"O��
@Jβ50V5�e��TY��	 "O�< �<I����O�T�L�"O
r�V10�0}�E&I����"O$\�q��M��5cV�D+0���"O:X�d���������H�rh8%"OB	���0P;ȍAW���D��JW"OT�aM���xh�O�%�Y�a"O�riT5@ ��
w��w�nA�1"O}ǀ8!>R��#��,�4UBe"O�4:�O[v�p�J��H#dYl`�"O�e�7ɝ\�>�Sb	#���"O��ڴ,��fp��@�aP
gxQ��"O��`���	$<�E0�lJ6ɚ�"O��Ҥ��J�%Y��R�S)��2�"O1���4� ��d烟C�RE�"O�a�O�: R��(ӚQ�4�"O���L ��5?��h�c"O��[��V�Tc��s���	��i��"O.� 'oǒK�LPaȈl8�, �"O�}��:y�:�� :�0�"O�\���n�p��u�^>aa6"O���e��Y��,�M�5�܁ "O2�y�����.�[���i�"O����z�<��G�	� m�ى�"Ol����	J��C�O� i�ɚ3"OzU����1��r�+�C?`��"O��S��Gu(�35l��m1F<h""O��	�a��t�\��5d�8��r"OD �-\���B�Z
��ٱ"O�d�w���f����M��5�"OZ�$��&4l0EU'���"O�`iԁV5J/2=Cc\?x�
�"Ox�z�����.W��6��"Op]����8)4�3�O���>�s�"O��C��
��@��o.Iq`,ل"O:l:+Ng�5B�B�2�β�!��F#z� ���h�R�ȩ��	�Q�!�D��J�d�H%_�1s 1<.!�dq��y9qd��t�5�^�
)!���P��	� ���T���bm-!�:3����b�)\Q�Pm	!��Q��a��`V>H28��ˆQ�!�DM�Mt�đ4l@
�L  ��P7�!��i
 ���ܯD���� �#$7!�9o��Z¤ϸ~�~�:2���$.!�$ � �v�@��@�@��4��*!�� �N��e��Z
��3)�6	!��[�x���sk�]T�A�j��J!�D�8$�|Sv���I �$s C�
F!���C��e�*�!�z�Z"�
n9!��&<��x�`�S�S����i !�D�\I����� ޖ�Z�I:!��9/�
pIe	��T_���i�O!�d�9M���Z�cF(9�|m`�Z*!�D�7	`��� T��JP�]6!����e�7 ײS�"�<Y��C��n�f���^�>�`
ŤQ�C�I4��h��7�n0�Eŝ<��C�)� ���v��2��� �	G�P]�`"O�)Wg�&0�����%Ǆ>��,a�"O��r ���V!�Tb���ê�y�"O�e�u�́NU�	cmK�~��]��"Op�I
R=d4���-a�xAt"Ox�C��-vD�hE+%�"O� ��P���\�&��an`�"O�\Ó���8@�$K�XL�"O>!��<�b� �J7�(ux�"O
�SwB:7��M*U�Y�a�`�y"O4Y��Ag�k�AL'|u� �"O<aY��.T��d@��J75h�i�%"O,���./t��0@V:Y����"OL��g^�>>|��ӅVu7��K"O�JC���5���Yc �쑂"O�S���I�$���F�D ���"O4ͪ��R�r�%�V��]wT�#'"O�	�匄� (jթT�Μ.�`1�"OȔ8%}�1��Z�l�ڶ@�!��RA4�B0�)G4r�q"OB��`�܀e�<��%��R�"O�+@ �k�dys#���:�s�"O���񌘙 ,	����y��Ԁ�"OB�z�#�j�@ӧ�d�fx��"O���"K���<�j5(��T�`��"O�y�f��BUu
2*հdM���"O��â��(��D���)]����U"O�0�P�ոWN�]�`�[��~8"O�Z��FOx�ófHZI�%"Od�ӓ��&[�!�� Z/LIj"O:�k���:�ѐ���	<9{�"OL�+%I�<.[x����ǋ%�M�b"O�MZ��ԏbhf��e�#~��c"OнbP��ij���-2�0ZS"OpT�3���`��\:|PJ���"Oz<�Ve �><�mϡgEr�"O��j'�̑Df̠3@+�&Q*�� "O�J��Y�<�	%�w�"|Sa"O��q ��M�p��Q�
�u��#%"O8q�Խv�Τ1uhN�1��A�"O��i�*rA�@:ҦN)ar�h:�"O>=�����X�XRA�K��(�"O.S�FiR��U�j���"Oԩ�dO��[`#��:y���"Of�8v�3Id8��t<*�xA"O8��'�en �`�B73:}�"O���M��}&�A�$ߠ�h	t"OzѢ��W�V��Qj�����"O.t�q,X�����S�B�,�"O�vY|� �H$j�����4"OxE:�ϛ�Z���F���ad"Ox`k5 F�#��b5��r�p9
�"O.��1#D�X��=sf>Q�r�K�"O��k��A�2�<2��:�0�"ORUj��9:>�P�@�9S��d"OH�+$��y��y&�=>\��"O���U��bvtpQ�AY����'�B:OX\�e�Z(P�yPU��nk\���'"�T��(AKؐ��eI�~g܅���3D��b�N�?pˈ�;�낗EX����0D�P:@�'Q[6�Y�*!%h%;��,D��2An�(?8��!დ�My;7+��i��P�P�>䞝a�m�0�0�ҕ�+D��C�ϔ2D�����(>] I���(�O��)� ��K��;g���i���?d|J�3GT�F{R�'�1O��R3�wl��0]�K%"OBQ�`��$F24���6xUB(b"O��㵀��"��ԁQ���"�b�C'"Op�0ᇏTx���)ݟ5��0ئ�|B�'y~8yc�z62�1��D+,�C�'�b)�B�֧ ��qX�-#D�<es
�'���b��\|hxȇA�'I[��	ϓ�Ol�
��H�E��NK23�i"Ob,3F���i���E��t^�Ц"Oh� T��*���flZ6Z��"O����H�]¬�����2$A��:�Y�����)X()R������f`|!�B�Ib�K��0A`��� ��IG�C�	*9��݁(�J
���)��d�O�����BT~i����i���׬ΏP�!�Z1��0r宐�,�� ����\�!�߼Qۢ�1%:�Č�p�TX�!�dT�0і%�6[�`��
��r<O֔hse�[��lJãG$�z�"O(�۵�/�lQS����?���"O ��"	1!R���W�R�33>���"O� �1	��P��D2�F�I �p"O\q�Qj�q�N���d�F��P�""O�(�'�?�H��`톹S���7"O4�{�j�>f��a�R ;��b3"Ob��qL0(�8 �)3=�l�g"O*a2׉q��E�)��
�"D"O(Lx�N�6i+T��ǉ;aRL�T��3LO�����$��٢�DC�<����[�|�Iٟ��IIy�T��O?N*s�������J�T��'2�h��\�	p예4�Gxt�'WPEj$oU�NK����雙>ր��'"��G.W̤��&@7 5�'x.!�a�?c�b����W0 ļ;�'�������+x�h� LM�j��`���.OQ˵�	6LD�i�� �f!d���'��'��)�-
�k7��7/�� %�5xH��'�����L9_X�퀶A���
�'"R�R��'*� 1�2�L�db�0�
�'��\��ڲ]lmт3_��Q@�'1F@��Ez:P�Q�[_0�-O����O����_	c�8�* �T5M�IK�,Ȏ2�ўP��:0f�h9q%��Cĉ	� S:r�O�ʓ�0|b OUt�tl�sY+!{�`X�K�<Y���6+蝡E�V]m�\ؖfAI�<9&�M�IKh�w��/=�]�P$AG�<e�h�{�L��)���&F��<1�d	�r��]�ǢE>\�$���Ŗ~��b�ȠG��V-~Ȉ%�S;vᱬ*D��J0�"k�nu�̊-?�B0ð'*D����K�x� �r>��[p�&D��D��	�n�`�O�O�
��#d"D�0J T�q��y	�f��-+���l=D�tّ�YW`UӰMM�c�8�g7D��R�%�7���Qn��|?�x�6�O��DHsun�ѷ!O>m(�m���4o0�B�ɥW�(�#���D��A�,�j[�B�I�8u�dhSgԝ!(R��S'Z�>ئC�I�-f �P�ZiނZ�C�>V�C�I�&9ؠ��#��q_�q�V'!,�lC��B�%�V�L��v��e�0a��㟀F{J?��ж*>�Z�i
��5DG=�O0��$��i��l��r7��t�� ��S�? n�˴��&Cq �)Ȟƈ-i�"Ox�1�A0H�P�AI�s��iY�"O�i�ф�'UJ z�*3H���"O<͢v�:���i#y��!��"O��:��P~ڈ���A�o�ʥ�0�|2W�h��S�@��t
s��AhP{cϚ�z��B�	 O�9�3G��;Ц1Q��\7!�B䉻E X\IFG�R�.y���ع;)j�d*��r���]�(x���Q�CS*uj�,!D��R�ÔN���2caM8X�p%%D���O�=i��)&b��0ъdR �6D�p�$��;VM�S�̜']��J@7D��)d��2y����@��x��6�5D�T���$9���E*���+a3D��8��~�R�Y��
�&?�`bC�/D�lQ�H�����:h���) D� ���h@�ص,��%�"�!%=D�T�u�\<L�=�R�>"�
��9D���G�@"w��۔@;o�2��sB"D�D0%Mݑt�m���
�iE�w�?D�xZBN�$a4 ��U���g*OfM���e���3n�7N�D\`���z�O�����R /r��f�ȳb"|A�'ZLs4��e�2x�a* ��'�"H�+(y4�2�Q�RL�@��'t 3��Z����3�O�,��
�'�ܹ��f��E��2��-���'rtu����u�pK������,O:��dR�*��g��$,��hW�Qq`!���t\� b�l���fb� P!�$�v�� ��o�
3���bȬ,6!�ĝL�ɒd�j(s��;!�D��)Mօ(&#"���gH�eў��ቶ3��-�Zr�ݡAF��3����@_����I���{��J�zl�q�uI'U����O��$*�OPuBPEF@�D�s�i�~� 	��"OB�����z���7(�}��@Sb"Od��Y{n ���-L����"OH�`U�$1B�8�kڝu��O4T%�'8�Qaƈ�1*��&M<D���bΖZؑ�a,GTD�g�<D���cH��mAv���"Cz��@%�9��3�Ohܲ#�-�|=�UF�2gi
��B"O
���|S�Yb���UST��"O��В-;_� Q�c֮A�ГU"O�X"�����`!���9>2�� "Ol1���s�qA�N���ˀ,̊�?�O>!,O1��?V�B�Z*�����L�������<	U��yH0�1�)ѡ$`Z���C�<a�S�ɔ��e	N ~�v���$��<���%I�������|���q�<a7kU�S��\`�2�lt�w.�j�<e��,�T�p;W�L$�*MR�<Q���5b��s�V+�
T�ΑPy2�'�����BL�����ھ�k	�'{H��׸y'���� l҅b�'y�pAɈ83�L�*$ES!D<�
�'��Ax���6��<���ѡA���
�'9��E��h\ʭկĠ&�P�Q
�'/F�Jpc��Aj�����e�c��y��Y�~��W&��<�R%1VB���?����sS� ��jԾs|ءef�->�d�ȓnr!���<���G��D�ȓ%@�zU.��^�v����2d��̇�S�? B ړm�'�0y��:l�v���"Od@������eȉ+��Bp"O��!b*�a�8���V��}�D"O�e�g
$1G� S�Hڣ0$4��"O2]Q�Nٌ!�ޭHp
��$�K�"OT%���P�I���QU�,s�T(d"O�H�Tg�.�6!JJD&|lZ$��"OX�0b��#oӰiJ�揄KX�|�p"O�d�f�8<�D(�A-$W�9�"O*�ެ&�d��["9��w"O�RWDE6\$ܭà&ۡXW�) `"O�����Ӏ��0��d�'p|��1�'LO YcdH;O��t*�N/��2e"O���%.�S�D찆n[+k*�bQ"Ō������N�Sė�J?��re"O��a��3h����!�IK!N��2"O�Z�B M*MFiЕ-����"O�dKe���D]�ȋ� PLd@@��W>���
{�������D#�$7D��Cg��a�rZ6�A6kJ�y�U6D���4	٘B��[F͊�z���'M'�Ic�����m�줻��?����:D�����J�T�8�bd��C�Y�0a:D�$�C��Pl0�3��\_�	JbF>D�l�#Ù�s�p�G�:�<=A��<��0|��*]7J�us"�R�l���"PN~�'��Y���n���({��UY�x0�
ƣ�y"�� 2�C�g/�Sn���yR�B�v�����Ic\.���ކ�yb(�5Q��(0ħ˴r��bWH�8�y.�M�H<�g"��T�~�2�E��y�h�MA�Ib����c�f��v��?1�R��&C~rr"I�!�"���,ٲ���	� �'�Ш���B#�\
o]H@s�;Ҧ�B�%/D���&�լ��!�[��<Ɋg�-D�@S��ɄM�	#rJM3$����*D�lI1�\��`��U��I�(D�� �N��=.���L^�2��"D%D�L��A��6�@�4I��j�.�8t$!�Iʟ\D��'�lX�4��&0������������?����	A�g�dM/!�F�dc('��H�+ރP�!�����S�����xB�N�\�!���YB �)�,*�&�[Gޮ�!򤛙H����׍��J��!F313!��]����2/V�F]r�Oʅ!��]�J��̺���Y�ٳ�Nܢk�r�|]�"~�$$0w�4��/��{�b����y��>W�x���H8au�����yb+|<��AT���
R��b̓��yR��'����G$U� �l8��y���6�HB��U k1"���=�y���?V�X���wҀ��Ee_��yB��L$�-"�*>uʚ��w
��?�����t�t����Q�+���q��-_9�@�ȓ6+�M���9��R����vxȇȓ��A�m@mp�-����'Ŋ�ȓF�p�A�F\5΄��9#�@l�� ��|�����Y=4���6p�b��ȓAZ�K`�70��`��*EB�@���P��0��H� 9��i�!z�0���)]����J��|;��o:�,��fD����G�E��2�c�>O�̈́��x!R'X��@�r�O�i�(8����0u`I�z�: ;�E�4t�M��S�? �YpQ�kך!��H k(D�P�"O�i�L��-�ntBJO�P�7"OjU�&M8&� 03���*n?4�T"O����FIo����I��1( ��"O4�2'jC,.T �Rh3M/���"O:\�RaΨp?H!�Y�n��Y��'bў"~���Y+Ji �.S%(<�����[��y�n1��E��C])����"��y2DX$f��Q+��X�ZY������yr+^� ة�7l8\8\��ꄣ�yb�<U��l@rJ�X�v��,X�yrH��h?��HH�]�: �v���y�*6��л�Y�=I��6h�=�?���������8�C�_:6�R]c�lN&�85a��,D�P�"�:F� �q��{\l��A@+D� 6`�"<<*�
�j(��7D���4�F�*j�2�c�=i��A1�4D��k��x �$��8<m���-2D�����K����� �Юz�x��+D��ʴ�W�7�����n͊b˴�i��(ړ�0<�H�.6D�Jр����Jp�Kr�<s�.W�k���,�&����H�<�a��
�rѪ�/��yz5�SF�<�Nט��:�$�&,$�0�F�<�a�@+1��ј%JB	m+܅*�MC�<���Ųf����3��r���q��~�<�ȕ��q�G�=Ų=���x�<m�\NlR� 7X�r9���w�<9Fō<F���3�އ_�$A0��w�<)t�[�;�p��U�܀bX��2/�X�<�e�|.�B��^�4���Qz�<��؊���p�ŵ�Y�0�u�<)���F��)«�.A��`�U��e�<�Ӥ��oiV���˒T�zE�7nBy�<�䄋,�>tq�OF���}iӦ�z�<��ܡ}�f`���1�ZyId��`�<���$4,����v�r�a"�Z�<��(�\��ِA��  ����V�<Ia/�p+(\h���=��Q���T�<�� ��$b�����J�,�#���h�<�!�

F�xDs����80r��~�<!�	M,k��2��������Gv�<1@�Mm�.U
�&���m���Ug�<Y2L�Hw�L�&뛧�a�Ǟa�<�BlL�5x4��a�ڠͬI����h�<i!���5u��To�3ٜ����g�<�0&�Rߖ3g!�u�ѓ�I�<��)+��M0o����.;�C�I��)��l�%Nb<ْ$�(Wf�B�ɖN�L��5jJ:p�h�R�U��B�I�c�+%�Yd<�s��� �lC�ɜHܱ�a헤��i��j��B�I'g��P`0���4-�E�D
�� C�	�Z�A�U��5w��Ź0$�6C�	�aZT�֪I+[�mhp 65B�6�����P� ˠ�y��qd�C�ɻ=�4$�J9�Lqq�Հc��C䉬#@�W��4l��1Z`�-k�C��&
#xiI����7���w�F$K�B䉤2jv�I�MT��zո���$�<B�ɗK��+�>&
d%�Ձ��a
�C�:,�̌��!��FI��c��
��C�IU\���t�'8��U�P�Ň�6C�	 �d4�6$��h,� ��.]�C�)� �K�O�9a���`��Y�"O�l��Ϭ<df��0#�9�&�2"OV}{sŋ�4�B]�`H�%V��%"O�`�fԹY,��[�hϝ�� F"O����0��ehM�@i��{�"O�p���R0��ѩ'�u *!Z1"Oĥf	S�Sfk�L�9KJ�U"O��yP�B�+�R`��	52�ȃ"O��3
�#}�PӪ��5�E �"OPq�)�M��U��o˘mטy@s"O��'�UNZ�q����`�S�"O*`�TرU��(Y��2�6##"O�u�S�(!�SF��<���a�"O"�&Ǐ?�`���@ƽ8D"O �+����G�Z1�%lS�[��ؐ�"O.!rĈ��<�P�qa�C�1d�('"O�i�3�?=��adN�G�}�"O����憕SdN�zbN�[��t:e"Oj6�9$$3vF��6ps��<LO�H�秒�K�@��B�Ga���"O�Q��$
� �����gU4�+�"OL���pd5r M��1K��%R����	��p9��\���E:8B�B�2M�&�)І�g3.�h��&�B�8d�Ĺ��&[����ԂO�4)nB�I�:��eY�H�G�U"��w<B�� �r��P�Zj��ZE��w�B�	�zL�$��`
�>��D��޾�B䉼b=��G���%���ؐ`�=!:$C䉽V�<��6�	~�]��P�HC䉴I�%��П)�VT31��%GD�B�gh�]����0<�a�
�\�B�	)E����&"����f���|B�I3eB�Tb$��+�
���Q-83\B�I�"|�TGĹp0p���)@B�	:N��`����.>֕�4�O"_�C��	�r��6�ֈ!POM��B�	�X� ���0��,#" �8��B�Ƀs�аy'�Ƀ�@�̯8t�B䉩t��bf	R���X�"I{��C��)xv���Ū�?�@�ȇ�eB�C�	% �|� V���J�bd �)&��C�	��44�R�S��(H��F�]�fC�I�h^�|I�^�(
n��n�:g�*C��6j�V���@� b�ݽi
j��ȓa�Xؓ�.�(=i�͚���,��ąȓ�و&������ݶ9����)���"�M#;|�`����O���g�5[���i�A��#11�5�ȓV�p`�
�4�nUS�#[6b��X�ȓ9��3 A�aH4�u�D�=� ���B�z|��L�V��K�'?�Ąȓ�H�q��
,I4Z�r�P+{���ȓT�\0vnǙ)3�t�̇;ڤ��x�x�{`�BdT��k����+�p��ȓ	�l�Jfɋ�q L�S�z�����[��YK�
�XJB�X���9�����$�$�+V/_.v�`��"�:fHK2D�$I�fو9�thz��	������<D�\��ܻ9N�A�d���z�TW�8D�غ�ĩ$"ԌĄ»a���I1D����ǟ8jBfT:��@�%����3D����,B�BE�"!��}��P���5D���pf[�p6*�x��B�h�Ҋ/D�� .��&�B	n���"!(�6��"OZ �1O	�Wv���eo��G�Ȣ"O�%�4D��rP<(8e	ѣOҖ�h�"OLyp�[5P���N#t�ڤ�s"O����6+�~=ʡa,K�&��"O"�S%�,��h�`U�s����T"Oڭ�D&@�*�إ��7ҵr�"OR�(a�e�R0YĚ����$"O�`���C��h�#�Ɂ2�*	�"O�8:�'H���Ug٤	H*-�"O�q��)G�	�hy� �1%:� �"O����*�'?���V�L#6j��R�"Op}�$A�/W�h�Z�F[snL�"Oĸ����<}c��P��A8dC`T��"O��)��N/|�ݑ��n�ZH�'"O��3ALR&=�ȕ�pĘ�Q�hm4"O���r�Ф(i��9�c��i�`�*�"O��Ra�� ��u�P��� 0��4���O ���Ћp��2�KP�����'�0-�!�[�R���RЉ�"̲� b�È/!��Z*c^d�7��b)Ʌ.ͅH�!��,ޝ��	K	u��9@�#�36�!�dW-'�||{�E!_��UZdcD�W�!�J���������1�~�!�d��vl]�uj�������Ð���O2���0�Z�����O����T� �!��?R�8����I��@BB�uT!���#T6��3+Q�R0 컧���q�!�$�&ry~���
!.�`��H��5�!�D��<0��(A�&�ZéL��!��Ӫ*{N����wLx(Ƃ�{�!�$��j�-�Da	�e�\ =	��O����`$��pFN>G�6�7瘤u�!�$���Z+���9[����U��!�ěo�:M�a�V-$��#!H��!�$��W��1�'�@�S�d�$�!�ж[�ZMa�7L��@��#�!��ܗd��nM6R��8`v����!��N�(|��e,�(�EƜZt!�dͤe��H�mK���TD
`!�˴b�H4N� ͈ir�Ғd!򄑢3�<q����'#�"Q���.;(!�d�)��"Bj�(?4u�X�:s!�$?!�By�
Ϟ[0���럮x{!򄚖	�&���*�e�j� �
��n!�DB�n�@�E�W���H���u`!��[.~p����� I��� �T�S3!�Ė4��=k�AU���E*mR�{�!����JQi?!�q�MP�!�ݟe�F� �Y�<2����l ��!�Q;.d�!m��2��(ԫ;)�!���B��p[v��E���P�I�a�!�$�{�� D�B�tvfP�D�!�d�bL�pI�L�H&��!��S�n�1@F�+X˾q8pD
�F�!��ߥ~��9�B�{��S��͜l�!��\l
�K%��(u��h�Ə̩�!�K�B���P�e-�����H�!p!�$O�u��X&�V-[�(9#Ǯ�Y!��R�mEb2�f��|+8鴍�:=�!��G�V���r�k&�IeB��E�!�$$r)��Q��?Dd�e�7�!��J�v�N9�b��']$�5�U��I�!�0�� rThD�	(պWcP�B!�� �<��惥XS ��GŇ*(��"OR�P����bD3��8~x� �"O��X'�ܹJ^�
d��y�����"O>\�#�Y.g
�$۳�żH'v���"O�9#HJ�z�lYIA��q�"O�lUK�i�`9,	��9� C�yb��1x�ҕV��6sb�H�t
щ�y�� Ԩs�#W!iR�Ak��@�yR$a��{4�>]������
��y�d�d�)�f�Z'@�ҩ�T�� �yrj�Y�u��@�97FB�Dm_��y��Z5qL� `�֠���a6���y�㛊_`���B� FHH��ք)�yҢ�3m+�<a�@D��H��h�
�y�("t��)
�CP�4^���Ua��y��"fɼ����0��������y2�3h�E����)2H̑R�ڽ�yRk\�-`|�#gT+N�Ċ��/�yr*�Vn�:�ƙ���y�le�\�G�^|�*Ǡ�y�������[!z]�������yRBR�G(~��*��h68A����y�
tq��P*[�cS:�����y����.�����D*�rM�"�y�o�'D4ӠM�==H5
�$�y2��:���ۆK��
�Z�٪�y�	ьI:x!�G�U)q��A*v`���y�"Ь���g[�8�$L��y"N�E�:�s��6c=��4AS+�y�j�;j4x�c�`�ne�Fo��y��A/T����UJ�[9&y;�i��y��Q9$=��8U���W�JÕ]3�y2H߸�zl0�톭P�6�+����y��8-C��H	54�����jC䉅d#h ���
KB
]�񩂉?LC�I�C8����C�x��0Rm�]�FC�+=/n4ӔkC|��((��3��B�	�P[4L�G>�t����&n*�B�6]"���قl� <����Z�|C䉻d�%���ct�}�G��+HlC�	 }$8�b"�X��q9�G� LhC�I"/�� ��^���Ui�
ݍ�4C�ɯ+��1�В���i�Jۖj�C�I�*��(�!�?���C�3��B�	�A܄�I��X���. ��B�	V����L�GqN���㛂�B�ɪ����)�6uZ{0JZ�h;�C�ɵ�Rxb�� �qJl�R׀Y5ZVHC䉯�L0�0
Fj�`��@/�?t]C䉥=ʼ�N˔;�<)k��#I��B��3"�I�%,9�6{�'UB�	.M��5ۥ���'WNxT*3Z�6B�E>>�y��}�2������M,B�)S����U)	������KAO�C�I�U��J�J45N��G�,)8�B�	�<��Г3���8�@��x�BB�ɤ�P
mX�b����*-�nB�I���q�7H���FK�&�|C��.X��
>I�Ჴ��'
�\C�I� t�ic)ݣl��MQ�Ǡ��B䉎~dv��
�0>���7�ʽ|��B��%e�pI���n�&�H��	�N!xB�I�l%���@dB&X����a�2K�jB䉈N��B7@�ƶh�0�Y-zc�B�)� ���@AX�����cY�gz��A"O��q����|`�D� ���"Oڐ���:]X�#!�� pa��"Or-R"L��r����Օ��"OjP���"	��p�e�3G��J�"O4����ŢZ�X�� V�]!pekp"OT-Q6΃k��P� .S�v%ɳ"O��C ���3�:h""�V�Fk ���"O (�KN������hjA�3"O�t9���M��% �K�DU��E"O�uZ!$�$����*J�W>|q�"O�L���$h�N$�D/�"08*�Z�"O^1��H�4m.*���Ώ(v%8��"O�t��_z`;�mW� n5Ca"O��@Ӄ��+�j<��~:J��$�&��0|���A(p��ͱ��]�@e�}�<9!)T�5�M)S. ��&��f��A�<����:x�X�㰠�6e���cP�YS�<i�@D;t��lÝ߄�˅+�Y�<����oų$_�mz�D;�oAS�<	"R&f�z�㍰
ưk1 �M�<����M�*,آH+8�� �
K�<9�˟<h� � �+
�@M. �G�<��)Χ��4�%<k�!�%��E�<!rjP�Tf~�r��G��`aNZi�<іoηV����h��[��9���c�<)u��/+ �Cj������^�<�����*V����[.C�`�� �`�<�d`à1�ay����ы� Hq�<��ѽR��D�-�v�v���^Q�<с��OS��A�a�.=�q��W�<�r��1N��:C��nX��b�ƆS�<��!�0?�MyA��H���g��R�<�R)L5t�{b�W�an ��U	 N�<�g�����@��[�H���JV��_�<I�ρ3�(ٶIH+Fz����GC�<I�g[4IT,�u�٩W��8թY~�<�7+¼y�:��dBQ"J�:��B�<�s�i`|���Q�SV4�A �I|�<� ��:5�*�!R�7����A��x�<A��\D<T�4ǂ9?~:LyG%]q�<��*�9o�@�C��G0�h��g�<y6E��<�2����9��#�~�<��"�7Q�bܓ�Y�6|Q�+�N�<4B�_R�U�H�� _��"�I�<��ϟ;1=��i���H�����]�<�\�8h�2n�0�CUB�<�&�����Ɖ�yڑ�c�@~�<i�LǼUф��$';#FI�G%�b�<�Q'��z�x� ��F�rrX�:�
Z]�<�� ۗeq0���'T���^�<���K/%�b11�!Yh6�"��\�<�AV�]K J��"����1��_�<��G1��Qd��"}b��r�U�<�s�$��UR.��%�vm{�o�R�<�Fǿvf�t�J�!#H����XN�<1!�k����T��1/�]�g�Of�<y�hƟ%�lA��i@�"�vи�(VL�<�i�#�$@3c��,�F(�tD�N�<����Z<L�XǞ�O(|��c�<��ʛu]�
�䄽O�Μ�b��W�<`�OL��R��W5d���G�l�<��My�n�sEV�"<�x2�AC�<��=p0��#�0
L0T�<� �2��fW�Q��Ė|U�0I�"O$�
�J�a����uJ*Ѻ�"O�)�f"�E>��%��K9D���"O��#�V�_� ��!ێ�\ݻ�"Oj�-[�O��F�ב �p���"O�P�V(�M�Eڳ=E�J�94"Or���mC�)���7��=Hή�Ha"O`Y��E�3A�TNܲa�z�A0"OB�1�F��؋���U��:�"O���� �DtC��ƙ�B�"O��yS�}m��0�F����0;U"O�\`�[���[�M�P�B�"O����]Kߔ�@�D�ں�i!"O��3ϓU^����ү3ª�"O��"�GԔ�ce�%�a�"O޴)U���>�s�A���m�6"O�i�5+!TTq��Y`�d��!"O�����΅3#�=��C2�B�`"O^����3ʖ��6�J*�>H�t"O����Q�lH�1��܍W��I;"O�LR"C�v�z1[a	B�f�p"O,J�,V�#!�d��+���X���"O>듦 ?6M ���kU�C�����"OP��ą�2F��E�l��dՆ�P"OX��]�	��p����i�t5;Q"O��Iu�I�6�"Q(�KS���Ȋ�"ORe�4���x�H1k��Ez"O���H�7&�����#ޛZ���"O��׭Y�T�D���I�qmT�"O��6jF�"����.f氢�"Ol�e�P.�d!k�CϽ{]���"O��Ӕ�Ԑw/&X)�c�>)$�0b"OlH:q)הoR��D�S�4�rݸ%"O�5�!�I�+#�hi�֨R��H!�"O��a���-�= 6�28M��"O1��oS�P�.�"w�	�:�4�T"O
|2T`��I|�!�5J��6�+�"O$�;q�Ɩ(�����;����"O��R�N��n�؃q'��^�&tH�"O����Q��A(��Y/1��Y2"O�	i &+���߫>��ố"O\���l��M�XU8*��! �"O��)�*X�T��:]���`"ORq��l��=,0��Ŏb�z���"O@����"{�N��� W rH���"Ob9�r��^=6()�Bֹ&$	Ȓ"O4D��є$����+�
��H �"O�e��n	�K��:��3TLF� �"O�eq���=�K��̢heB�a�"O|a�3DQ�d�,9��#�� q���"O>(J��*IVĒ"Ɉ"p&8x�"O�=�EL��*�ʀ �k׼hܺD"O�5Yf�G$`N�p� A�v��l B"O����c��j/��X�/�1u�څ*&"O��qЭ/C��d�oĤv�A�p"O��y����v��5��YsJ�sb"O^@�/s���y1���<lĀ�"O�Ѹ0��&9�i���0�0\�e"O� �r�[�e�zY8s�̇����"Oa2�肨b�b���o�F(@�"Ofa���ߺ�����U>H/��a�"O��@/�y���@���66jq�S"O������V������5<�ᩃ"O��d�\9V��M��,Z)�h"O� n���Z
o�T؊ċ�/���"O(p!����)r�X.c��̐�"O�(��H�gDL1�I�%,��5�1"OL̊2� �DgԘDH�;`ą�"O�U@'��g�Y��T}�����"O`t�� =W��sqeP�[�$�h�"O^q�"��'U�0�*a�5��@P"O���5��)%cS![3,�d|B�"OfĂ�E��Ah�c���c%l)�"O}@�'M<��H�!oHO���P�"OTٲ�ϝ�I�0ٰC�Q�6D��"O�$���	�{eH$_��@!�"O�%	)�;?�p�ZR�S?lH��"O�	��	7������-I�-�f"O��H��UF��@�-M7X]�"O:y�b�@)~����C*7Ԕ �"O�q� `_"��ir��T��zɁ�"O�R�Z��t*�đ�@T&�"O&�Q!�D(0�N}C�c�u��U��"O0Q�O�6!_b@ʶ�̣	���$"O����Z �0}�G�Җv��P�"Oʌ���fU���Dgu�9X�"O8����U�MM�I��W�X���"O�|��쒶"evl�f� ��TQ#"O��CG��hs8H��%��<�0$P"O:a��gM���/�y���q"O�����G״����K4�P@�"O�}B�Z�RI!8E��R���5"O�ԲgO�	~]���(Xn����T"O��ZE�L	<
�`b�Y޵F"OH �FCߪ4�2e
dlP�C�"O��'�m��BLE�]16lV"O���cn�����5�}Ҁhu"O�e9�k�I`�
3@%P��y�"O|9�ꃏCb E�W`�4:򼵓"O`t`�IU�i$n[�tb�"Oġ�$n��=���J��Rp"O\����*��Y����p�@R�"O��
��~�2����P'���'8n���o6��@��?����'X,�!Ũ^�H��-�f�ɵ8VR�@�';t�`�y�^1c6N�.�l���'����qF��4��aV�̽0�pX�'�,�8cΞ�}c2)�V�%�f���'��h��h�Y:�������Hq�'Q�ɪ�d��{gJ��,��]���!
�'��Q���m��	j"��`�61�'�TEIR���E4X��'�W�F��'�ڠ�sB��3zIصč1K~Ց�'_��0
�/Z�vثŁ�4F��'��r!EQ&s��m�0��y��(	�'�h�hV+E�AD�]C e�*t���{�'�q�&F �D�GeB�eW���'(r��ŋ�|���S����`�j	��'�R���.H�4�b���I�U��j�'F�Ԋ��Ə)�Թp'I�LC�U��'?�tp���d[<����LÖ�8
�'���K�,L�y
q�L;r�l��	�'��l�l��FxHd��
)V]z��
�'��qH�̪Kxv�R��6b��"
�'�r1��f
pF�!kS��gf��
�'�~�Wn��w\��㮓*a�L���'$�8�����n�r��!,���'..�3KM+;���J�,�2f6���� �x�$I�@-���1CA�m�ID"O\���3���%� �:
օ`�"O ��ݿI"�i%��3	�(��"OBx)գN������NL'w�t�6"O$Z�99���J<V���"O~��B��Y�x�;Ak�T�4-�""On�/zY�f�V�r�R��G��$C!���]N��&�ǽ}w��q2��:�!�$�=,r$,�eǑ3V��H2nοx�!���m�4���Q��Qb�Z0"!��ŏ:����n���b�I!�	�!�\T���Ά�N<#k�)[ !��!i+�@����7��X0��K�% !��k��<+��A�W�������k�!��A&�uQ8�`�� hM�nG!�$d���4�
|�6�x"�I�!�ğ>-�u�S)��{�T�8*Ў9�!�$�A���ׄ˞<?<9��jW�!�D�j"$M�!(��e�,�*����!��ڝT�x�(��Bk��ǭ՞*!�d��8��%�ri^����E4!���Qǚ�{b���������;J�!�DѤE���wdٟ$�9y��Ff!�d_./��Aȁ,��M��� !�dN.zh2,(7���
A0K�:-�!��Հ|��M�gC����J���#|�!��P��x ��?�E1��0e!�ۭ�6dh�"��p�,Y�'�?N!���*wH����U�9����j3!�D�o4 ���>2���菀`�!�B�R��u�ܻ	C�Z�k�!��*f��4ab ź�
����Іd�!�d#!����Ɇ�`��̠'-�iX!��ȍ�"e;��u-�UZ@b8'!����"'M�0T�&$H��lv!���v�4�u˓|�`��B��l��Ox�=�������z�~��$
	0C���	D"O ٺ�O�t\��Z3q �!"Oؠ��ə�wEA����"\ܥ��"O���غM�J��b�X#t��"O�<cdA<4lM�gƇ&i�m
�'�����N0y�,S܄r���	�'�ĩy��Mb�9i�m�nҼZ�'��9&�ޜqH6�b*2�a��'����F�430�򂐋*@�i����6�o�	�e�H�0Ձ��j�N܉�"�(��>����,-D�L�t�~�Q�dН{�Op8�͈GNV1
7%�
M��u��O��X��R5'�ʖ�J�Q��y�n�,��'�ў�b�,'N_eY׌�m�h��C�'o2Q�&�/o
��X��9~x3�'��10H�،�u�,h9*�'�lL#&�%m" t�) Q��'��-q5��f�ry�Bi�6I}����'(֙����}�8B3O�C�e��'rҬC/;�Q˛	B>�9��[8�y�o_��`���aϬi��;)��O*�;��#}j �V�V�lZtl0/�N5��J�A�>�S�'FF�01$��2�Ԃ�A*	����/O�O?7�,�΁��[��,��W�U�����ޠ�F�ܫS7��sw'�"Ɣ�'�ўtGxrJ�O�^ܠ'��l���2�l[��y�Ի����h��\҅�ٸ'*ў������@1t�eS�7	|9p���.�S�� ъ�!<�p�kWJ�a��P"O� a��̵,�4��%�^I�� #�x�C�����Ҧ�Z;��
�g�����:$�Ȱ4ĕ/W�.DI����$.X��$�Q,\Ur��'�'o�)�s�x��NL��`�@��Z�7ݒIsA0�`bz�}bugK�a:d����G���jQ��f̓�hO1���h�hO�Z��u�3�H^�z�� �x�eB��Xe�=�~� �6��:F�M-�F�Z�'��y�K"C,�طI)+�:�2�ҙ�p<Y���
%�N�{�jQ�.�حIcE�L�p���'�J�d��iצ�
��<X
�'-nD����6��Ȋ!4����	�'��yXA'L�Őh !&�r��1	�'���p�$�~��0l�>�%%~̓�hO1�T� �o�����F9V���I"O�-�!�Cp]s���33˖�(S�Iox�p����6[�&H3��]ohѹ�o&<\���Q$�$L��O�YG|�q�"k1���Ӡ`+ ��'MZi��߫v�` ��	�<!���˛(���ɧ*Ϻ-�x�E�&)!�dM�z=��AU옃7�p!�#��g�'�ў�>���n	�N0D��ڠI��� L"D�t�$V78ܦ�`r!XN�(��!D�$k��ԏ|���>[P�0�:D�,��[+/h�M�E��7FΥR�	<LOz��J��%C�n\��˦5��Ҥ�V?�!��Q�� �̒)�Ji��*ξM�!�dؙ.�`m�F&L� ���ڡ�A1P�a~2�Ol�c��������3qx`�:2�
f�<C\�b<�(�%�2�$ �cm�m�<)��<Ȝ��2��;*�@��i�<��՟*'�Ii�b�B�I^�'��&��h��\��:���>{���b-D����E��w� !-8��y4
�i�O ��)�x��&%5�n)�Ə�|�bYq�'ғ������3���8v�|G�����-�#=i���O�,��L�G)2��d�D��4�'��OԢ}�A<%q�	��@�A�9\���ɕY��݅��a�f0H�� 48'���fڋo�C�Ʉ,c��(��8��3C�юC�I�Z>}Hf�s+�j!�R�D�.C䉴U�b1u�P�l�9׌C��C�	lL�`�
}tlzҀ@0q>�"�S�O&�!�"\�h��ke��Pq��'�qOn���i�HJ1ʵ�
�m����"O� i�)@6M�Ib0iL]�nԣA"O�!�	͘;�&�!'���S�2(bD�D �S�)B!G���g�i�����X�X��D{��v�!���:(fN0����*̪��{����>deh"�&9e5\yp��v��=E�ܴ�x���,̱L�����(c�rԆȓU��,hE��.�4x��/��DІ�(�$�1��e�(됎X*���)���;G(H�@2� �^R�8Ub#$��
���&x�"�D�Lc���C�#�~�'��)�Cۃ,�HX�R� "/�����(On���B 2��T���N,s<mH�"O���]�w��]�s�]/W#����'3!��_�7=t8AoB�>���`��H�!�D�$_��xmʠ3��y��l˿)q�}�������
�9���@�U�<�؜!�-D��a�%�|����+�n������7D������^L�(3䎁�z�Xa7D���
�R�$��kY�>GZ�;2 4D�� �BΜ7
ոu�FNJ�\�yP�"O6t
s&G�X��	Q4-X%S���P"O��[p���B��� Q���V�OH��D]2z���H�<Vre�e/	�!��ʦBo4qҷ��'����FB7{qO�����
n�:�#]�-�v(�SQ�!򤆪xIriYց��(�DXH�a����^x�������w���G�[@B�e8OPJ��dI�i�d��H�]p���\J�!��\�'����� �	��m��m�1O,�=�|⡁A�U����1��i<���'�I8��$���.ƅ;�,�ЦE�f&���#D��K��7
�y�s�a�0�F�!D��8�l�/
ր�W�K�b�&)A�	?D�Xr�
������$T�B�E����<��'�qO�2
��Q��ν:�>���Ġf���$1���  Q��q��r��i�@�R�9֬����<��OdU�'/@<��t�hPR��<��"O2�0@ I�+1�xcDHQ�:�P*a"O��!��ABtH��,**���!�'��'w�K�j�@��"���JA
�'P2ԑʙ' ����b���m 
�'a�A��E��S��s�hTBH8�
�'�0ɘed���h�'n�3��B�IX	�m�� z�:98RF��Ƥ�����	�Z����Ǖ�{����?q�E�IY�!���7g&�����D��&�����ʁl2��y��ڢ ��u�e;D��Xv�Q
_�|Z��F�QJ�y9ņ�>�I���O���$խ0�ġ�	u� �XPB@�r�!��[�n؎����O��t��#	+9v��:�O�ܨ�$H4}�4x�)ڃL0��� "O 9Q,��r*����&!S��c8��hR�9�vE��Ѻ/��K��!4�����& ,�c�"�e=~�r����x� �R�nQ�q��D��k�h���<a���$"L��1@�4+d�ȳ�ӹO�!��	4јP��B9oI�4����'�:�IR̓i���5�.Y����8d�0�ȓDIB�[�BV"+'n�H�	'V�j�IDO9k1F�,^<2i��KY�B7�4p�"Oր�6��0�R �b�S�����"Ob �M
�5��\HQL3R��U $"OH�0e��btF(��(Y: ��|�c"O��h�+�0/�Ѐ��%8Y�`]�"O�M��jƠ7�Z�S@��.��%A0"ObES�$ۖ O��БL��/�U� "O(�Kd�:R�#$L���,��s"Oʬ���C[���,]���@�"OR,P0)y5nU K�!=Խ�C"Op!S�(�Q��UA���~�#A"OdMh&fZ�$�8Ep��9��Ѻ�"O�}iѧ߽f�0� ��1N��ZD"O�a�7�Z�x���{�lM9�Y�"O<�Bu���"��|�P+X�4��1��"O�-˶���,(��#K�8"s.u�P"O��YG�D-T`J�j?*r����"OzI���ߦBwR���Hęo.���"Oxt�A��%HX�!0����Ya&��"O�r��΍0֒���@�s1�<0b"O�L�/ݶD�tY���^�@B"O�mqP`ŕ�~�	� �Lv�yP"O"Y��iʜ@�FJ�X�0�T"O  �&xY��߶�X}:�"O� ��U	�&1X`˗ǒ#M�v �"O88IS+��v>"�0�fI��,U0�"O�9"V��N��u)$Gº8�F$�V"OF 9�d�<v���@[:7�FY�"O 4*�+�1�2���ԕc_�4�"O�5 ��#?�:	��B�S*�Xq"O�%P�	�?`��(��A.�`۷"OZy)� �g�<�p��)`����!"O��J�D�.	��`A��5n[�="u"O���GU'xPV �B�W��"O�U"p��Rz8�H oRD��2�"Ol8��K
�A.��IQ�:r��A��"O��(����5S��D�t��|�"O�9)$A��0�b'I�p���{�"O0ђ�̐�M�<�l]�p�0"O��P��U�M�����+�����"O^�Ԩ�3<�hY�$(���Z�"OX�82%V��T�q�C�(���(D"O��G�5�%I�ȊY�v# "O�t�$�O�4�l��NI}��#"OFa�TO�@��DIc�+ `���"O�Z�  ��iU�b޶� f&�	\!�S�)r�� ���%�����>}!�d�2cA�T�%.�
C�B$�a�?!��Hm٦Lxp�<`�F�{���!�ד'"�PsH�Wݜ��b監Z�!�D��Ag� *  ������ �j !�$�y�tz�N8��Yo@š�1l�A��Ӹo8��(�n��y⡉9Y�y7YW�mѣ�yB�]B�L
�C��e�� �=�y"c12"h���0,,���e��y2a:7��ȹD��'9������y���m�8���-������yb&˽�jM5M�<1:��f���yb뉽^4��H]
,S.������y��7]��4��D�1^�Bh�P%�y�ET>-l,PȖÅQFI�g�G5�yro֪Z>����'I�z��ŉ�3�yr�ޣ.���l�%�� BE�E�y��.5lP�Ƈ��$�,��7�,QJ:�B�F����h��ߨ|��92�k� &�,�C�O�!�$K	F
�:lD�8����zH�ݴF���-�E�r��	$��ze`�!�`�	�f+JE�z�8r��J%�ƭ�~��Ԣ��F�(KalH��y�#����jg.�B�2��B2˸'��3�a�l�f铯6�`���oZ
]��$��bA�7��B�I�[��B �I�GD�h�!"6��څ��#ʒ k,O���Y�@��mµjI>��bd��%�&C)D�8�e��E�@q�ʧwFT�� �Y�D5 �D���hj�^�H�A��>�����¯*춱��*9�l��0+�h�r�oڻ������M'	�����z.�s�<��j�v���N���+���Kܓ{L���t��$Q���`���`�`r��1et��˦�T��!�d%+�4����&< :ʓi�]�L��� 9K�i�'er1G�,O����ƌ"�R�JЯS�����"O����H��fQ�14���P`���Q�i�9���J!��Q��I��(��Si�B��a�g@W�i���d��zp���&|�c������#"/�>i�)��O&D�,C�~��K%�Q�@�N��dj$D�� D�Ρ]Y���N�<���O�ʵeZ* �&�O?ա� �9E�����* �t�>Ա�O�h�<Q0d�#E�2l��>#><=H��l}�![�r��١�Bx���"��9���%�"����@.:�O���V+�8k>��� ���r�.W�j���O��R�8䀑�LlH<� !4���3�EIےiD�Xn�'ւ���@�#1�������(��L� � LQbhiWI�>�!��ȲHx�R1[�7<t�󓆗�;q�$��"��*���yy���'(MX�@E�+�,[@/kKX�<�j�`���DWN'(	��N?�ՠ�5!��LZ�H̰<A��44�峳�N�,5��� �HE8�܀b��$ȱ�S��%v��2��v��@�4�Y�ē�nDb��ݗ):��
!���m��EyB!���zl2�\�+8��M�,AU�آ�Y<|Xl1�"O�\1�R�[p��Cs���]R,��I,?�+��<E���)� $���4���5*��v�Ʌ�T���@c�[�Z�d���"���'�6Ųv˗�:`D���	?v]�H�e�5I3.�Bs�C���������s��m�`�ե֬U�N� ���Cf�C�	s�� �$�تښ9�� 8�C�I~��(P��}���вq�x�)܌�	�n���R�x��צ�F�ء��I�{j�B$\�غ�IV478�.U/aDN�Z�%D��Kg#G�rtP��(���9Ԧ �ɾ>��<���:z2�M3̟�v�)��.ɪ�t�^42���P*^X�H���$t~4�R�Y�bt~��6b@<��Qb�{r0�$���I��H�R��kM6�~bÒ[�Hl���[�"ʒ��l��y�e��Q����/��&tLx�ǠS<�?e�
+�n�Xg�6|6�[����?��O&vHp�瀳~z���
?��d��I�Au�͉�E�\��9�& M>���-�,��ÅT�"�x�R�|����N���� �o��4k$���>x����U��3�.'���K��P�l���E7$�`��h{��U(/8�5�t�Wyu�9�h 7}哌_I���̜����H1��^����X��؅�ahڎT�h���]�*��!��3D3b���C�m�<������Ǽn�2����.���A�B;jĻ�ꂘl�>東<^���%N�{��1°k^0F���Dކ1E�/Z�jQ"!�N�P���x#�U�l���S�@�$��8[EJ[�7�P��fOʺApQ:Q�'���(S�T�j�{�0��ʁ�H!`92M)���;庄����>�z�2ٌIY�(ДG:)��� S6�	�����H
��v��8��
i 1��O�-PW@[��6!���|�=�@]�	�����L�8U<������䦭{�z[��rg
F�7��T�� 8���ge�)��Iү�T���C��11���jZ1D��
g#�>N;�q!c��B����D�03,��J@(
���#/��a�sc�H��*M�P��6�Hza6���z ���`�O $�~�F�l}���t�S�Y2���u���p>YV+�$P㾈A���#j�
�)��x�\=i$�	;Jh�f���A��L��(�D�@������Ğ�UI�K"e���te��DM@1���J�J�4i��(O@Q&�� @GV�"�!N�F�*d��fS�<`�`î.Ghj'�w�����֖g2�o��,�u�F$4>�8A`I������#Xpxl#�����4��,n��(�U��$5?�Ͽ+�C�/����ҕD2flKAB�m�<Q�(Ʋs%��)��<0I�MK�N&�h<#W�Zp��[S�#�"H�'�HO��(7+[�z᳠(�38�2z�'��4� ��&x5��r�jȴ{�2�Hqj�4|ր�Gg\�!��d�����a}�6r
Kŗ%��d�C,hаEy�fr ���Д#��@�v��i�S I�����
a�ݪ"V�h��B䉊F�0�Y��Z�B�te�&�A�Z�֨`�h��ay4,�ik��
�h����5dA�s����P,jݸ�k�)�y��)y����'g6�؀Wꐃ4+j����ɑ1��aJ�}�p����@�q#�& t���,Ta���*B,+�OPA�$ؗk4~�8VH�#^�����C~��q��P��M�#DK�5�}�ș*gQD�1�Y +֐�T�+�hON,R�j��r�Xvh�4&5 �'W�����ݑJ����&ɜϒe��y|!��'�� �(5�$�_�B	�I"{� P*Mw�U�Qm�@�O�b�:0�!&���2I	�;�<�"w"O���/�)eڄ�;"h	=�H2�l
��~2�]�@p�X�!�R����� e�t쑁��?��J�ы.wl����@ɬ���������&)$	W蹹c(��/������6T�ܣM�
�hH���ax≚�m�T�=IP��;���Cޢ��}k���B�<�&h���t�Y��ܚ�r��J}�<ِ��e����T��:��8��+Tl�<A�k�Iy���b��!Mt����L�i�<� >DЂ�̤?=�@8����~�U"O�A��O���+��p<t1�AE�l�����Ox<rc��R�R� �҃yu�y3T"O"E���I�Ro�(+�*A��H�2�>O��	�&ϳp����B	z�z��� �U��d�E&)�{�,X�}"��ɦ�#A��Ayz�r %U�z�J�
,#D�``P�O!0q$���
 ,�$�!���G�4�`�Ϟ@b�>	Y@�I�I� �҆���Gf#���` ��i��@'ȭya��(�hA֍�x��Y�ݙB��O8�}�exz�i�F\")�d�E�Wc` x�G�TnqO�}��_ՠ����Z:Hq*ĩȯk�Ե���{<���e��&@�a{R��(TT�X`H�,��D��,�	�?Ye Č �>��8�����|Ӥ	���+ra���"F�W0�h��'fj����g}2�X
0�,��D���"��@������'2� �/G�fQD�$M�pZ���ń�/'�����!K���'Q8Lq��Zj�OVhYݥ!���Ao��W��+A%�V��E�1b=}B��PS/?�Zu`l��F�	�Ξ�6���È{B���MK3ym�EW�� t�fE��k�0����s�.	��I�e�H�P�R#62������Vn�	�.=�቗E��2`3O��u 
Q9��ƍA!�*1"O�IH�Bܙo-���"M�r�
��"O��h��4r)zU��E6��"O������P�9���P%ڭ�"Oh�adM�n�,k�KI�q3"Ot�k��2QT���U=.		P�"O�����Q�N��G�([�m8�"O:��虸Fш��ǂ�'����P"O�t�7EԾn����\"�� j�'@�����ff�Ɇe�j$��H�'*�t�1A]�l�^�)��?S����'0J���L�2��HF�e�����o�~�I<)���;g�	9 �iȘ:D�]�<�U �G<��$UlXb��XF�m] Zä8�)��\� P��aP?z0A��[	A�B�I�)�T�c�֪�0�sK�2���䍘Y>�S8,AD�Ǧ�:�����97��d1TvGζH�m`0$�;��ycf#�dp����Ťg��L�`��{�(����a�az�L?
f�O�e��g�^��"���jS�4ڠ"O�l�^�G���E
?G����DT�<@���{���'�k�f�Y2&E�$�i��յ�ycP#g�a����%&%��˞�}2�Ћ��<aUa�#S��3��5�{Pw�<y�i�)v\i��M�:K�V�p Z�<��c�VX�)�5T4���T�<vNf�A�ɰn8:qtcP�<�'nTL�Q؂	��v�Z��e$�Q�<�hΒ8F�D���	~B�XJu��W�<a��8|�0�8��w�:�BV M�<�FI�B��aB��tC�Uja�a�<���K�>��u�q*�)l��Ka��Z�<��n��a�P���)|]؜�e��M�<i���E>D<�2l�?��m�/]f�<�f��m���PT'W=9��*��k�<�" ����㦊F"28k�z�<��Ή"l(Z]Z���t��b�w�<���ɬj�J3�9ݐ=�4GH�<��j1>�=("�K�lp�KG�<9�n��H̰�O���kf$�A�<����/z�����1+e����}�<�	Y*�6�����6�5I�V�<�3	��Cp�(�Qۿ/���(�Sk�<���X�U��@�YW<��rN�~�<!�AM]wx��	ĨT
2`�R�<� ��Rqe¶��CN���@"O�0���1x &J��ڱ��"O�=X�`_�$H�+P��8�"O@iKw	D+;�4x�@
</�(YIp"O�A�C�9-�� 8!���
�+"Ob�aT@;ϐ9�s���P����"O��ʧBI+<DCU�MO$��b"O�q2�o��jH6 ۝`j�*�"O�z���7$��LcD��\	�V"O�!�!C t���⑳b$��"O&�y��#P�9���4���T"Oʄ��Q� Hs�Q&#�Ll"O�ؒb�]/P��h&1�B��"O��ɀ�j$l����A�Z�t"O"�9���/�M���F�c�$ٗ"O���0�!;I��3uJ�?]����"O���,��iX~���)8�Б"O��вj�R�(!⇇9H�3 "Oڌ�D��_�
��Vƅ��V<�7"Op�j�(I�!}�*%�B$l&�T��"O�����������l yط"O�xv- �m�ff�"'ŲW"O�$P����{F� ��Ä!�X�`"OdBv������^, r8f"O.L	��T��~�."Vv�XPS"O�X���2I�z�C7	b�|*�"OJ�X�dZ,b�:	ԍ� F�ѩ�"Ozi����^��iSmG�	���"O�ԙuj��V�t a��_&��3�"O�-��%:~�bq�T1<6f�"O�!��wY�Ͱ%'K�Zq�hK"O���A ��_���FT ��<��"O�Pj���.|R9�ৌӲ��`"O�AKv揯
����V#�VQ8a[r"Of����
�3�蹐���qW�<(�"Oڄ�F�msX����N���"O8E��O�\4R��,N����"Oj9�E�V��$�����<a�"OJ�J��}�	�0-�=˰�
f"O89�!��"3�]��T1cĜ�"O@�!��2G��H�6�\�$�:|��"O��1��ʑ<J�b�G�mf��@"O>L���DJP�5O̹\t� "O44��j՛X��1��eS�+L���"O����У2�)�r��3i����C
5:C�|����#Eȶ�b��ķH�l(0�$D�����*2�$����>~��9�RDl��trf�x:��ߓFu�u����:����۔Z�\��I,~0p��FEֵR�m�м3���rx����0��B�ɉPF�Т�努W��}��I�$��XI��y�Z�r��U�O�Z�O��Zae�S�^�C�'�P�C�1a�.is�i
~~i�S�D#?��8+���<���/�gy2$M$sn4E�D�0J�����#�5�yꄃ_�|�\�}�����Դn�J,��!40���J/lO� �"2!-��B�t�|����'�4�Ӑ�(� e"�i�E@�D�<���R�Ϗ�xthQ��'P����Uqm�4�]8dR�h�{®�6#v���`�=u��>Us�T�y�@i�$�'���	sm/D��y�.;|�� G�8����Am��̬��I� ��5�(���n`���AbĄp���0�W��dC�ɺR�p%�B�Km$�@�/P�*�6��*�D� )��=9��ȹ{�`|r����en��a�c�u��LH�f�W;�]�E��;�̐;T� 4�����4��Q�҄��"m�3&��й��S�? 1xu/4SNA�S.�
J8T2�'F��R���;�ɧ�����5(]��Hh2��21x:`�a9D�� �
�*Or]P҃ϓf<�%�G�>��k�y� �!1<O]i!��8x�ޠ�`�=�!���'c�3���DPVܠ�OW'b>43�N_�h���x�FU{�!�D�2klj� �/� a�=�Q��qM0	aD*���z�' ���&�[�yԚI�eN��c�v���*%�\��!�1,�%��[�:�P�rb�=�(� ��3N��)�������|O ��oE -��f%D���/�y�|�xD�G�z��奟����Š-0�Up�˟~X�����M���1#΅�anH3��5�ON���M�Q<���' L�HEUP3�����dM-&A��'��E�M�./���ꓨ��u1��X`��m�#�,,��b?��e�K�.Z$l2��Ϡ?���ӌ(D� �# �'�Y�L�޸Ã��< X�I⁎���2(O?�d�$^�ZH���=/h؅¯+A�!�d�ML�����3[DR�F������r��3i6�y2A�+"��L���<(M����W#��>����#u��*"�ώ&;����!��3%���y�݁<PA�JO�:�`D��y�D�}��A����To(Q5�ז�yrO�z����� e�P�e��y�I�o }�����d�+u�;�y"nI;K���*e"	��,�ٔl��Px��� ,n���;)D�Z����F�Fi⢆�Z����R�'A�"D[�e��}KD_N8�DXÓ ��9�o�"`��d����%
EU*�X��j�nc1s��*D�C�D	kT$8���-t*��5+,-B��ΟJ{pp�#IX'K��#������V���Ի1<�#׫�	=Aڕ��0>�Q��/F�(�i3J��i��]0� pp� �T*Y�Ne��_�������X����շk���g�~�hHtmG�U����F��$X�A�OtM�͌'I(����o�����p�����IJ�z,�b�a�T��RеG�<��F�ʓL*�p���)�����ʾtȅ)T#
#>YkAn��0� �ʅX�R���t���Oȴh�E�U $(a3ю����N�c=Z�⥈\H��:��8���34U���@L(����-�:�|;Nߑ�8u�2k^�K��3ǳ#��%�@,�ǟܐdm;�d kb�_�|2fNI�.��pqGˈ~�4[GUV�'_�\�cmE)%���Q^��+e��?ݪ}��"T9/�tʦ�I<Rm�S�[.ҢΦhP�qѤ#T=��3�	.Hzh�iH����@VF5˓ �DL(P��Zx� ���$Pz2H���)��,NthB�� 8��|@��C�7�dq�q�S�w�ȹ�HK�V<��D�i�����VS�� �jݠfqn�ѶHσk�~�`*Kf��=:f7��ؖHQ��(iV
\#�~R����*a-^�M>������?	m��^գ�K�$���	��O��je;GmԿY�>9s��s���j0LV6r�D˓sfȥ�c�A0X���(y�����K2N#����i��s���?��"-t�,�G�'{����f�^�}ڰ�2(�o��E�PE�4 s��R�M�A(<� ѭI�Z
�KM(hJ\Q1c�Ojy"hD/6��5A�́?�|	Xd+��W�F��~���:.7�����B�����.�Y�<�����P1K�N:b2n�䈂���b0f��U�g�v�
��JG�	�X��ԡ�� ��D��F���W���r����tm��u)*�XBh�,x�jC�	2R���c�m�#�-{'&S6�C�ɭ7�P���G:]��A����8n�C�2fĥ)v��;;jN���K!r԰B�	0,d 8 F%ܫc����6��1bZTB�	(W*�ѐ�B�P݌�7k�*d��C�I.yJ�A� �JPE���ğIcC䉐-�*X(�g@�%�6U��4��B��?��Ѣ�����R�^	��B�	%m4p�)���>c�ؑq�݁�LC��(K����!9?,�ZH��SdC�	1J��1+�1jw�\R�o���hC�	 �x���"�I��
�L�!��B�	�Z��2Gm�aF<4���=J�$B�I�c~X܃�Lz�B�b�
�W'6B�I�o=9᥎��t�K�
G���C�)� 6<iP��w|C鈷T5��i�"O���r�\7�6p8!)[=s86�Q%"O�áN�*,�T�ƏYC��"O�|+��R�RwH�QZ�C��c�"O\I	bR�&�6%���04�11"O"�b0��P��X�kǂB�]��)�)*�����O�]��j@v��Тi�!?��e��"O���Z�,�j	@�b��w��p�0O����V($���Z*�HػP%��PLjR&D�1��{bA��%bL�(3���8�i�<2�(�W��0u�Ҹ��g%D�����0f䮡`�����p� �ɗ@>90�,s��Ɂ?1^-��K"8�$�Q�N�j�!�ě�EBm��˾(S��Fb�:?��D�Յ(Z��Oz�}����X�`��r~�0u�I	O��ȓ,�f�{ЦاK�9x���d��I;j�M�tAXE�a{�lS�z�P-c�ρ���d�` ����=�`o�	
��P�,sӔ��U��U��ÕB?M�q�V"O��`�f#~}�3=�2��`�dY�0�A	�H��s0$	�bĥ�e���N�І"O>�
�HG?PN]�&b�y����C��z�P��U�$6�g?�5k�����Z����A�2x��Ke�<YINX�hbƭ��-�����<���ϧd����
�i�P��r( Z��X����*shh���>�ı�1O�!"�F��������R"Oz|� �V2Gw��1fɎ~�4� "O:\�C�O�d���5�[���`��"O>m���\�̚�(�Ă�1�9 S"Ofqha?[p4��"�{7dRR"OFMSEiӌ+��Țt��1A=��;�"O�����^3-��p�p@�+�0��F"O^���f��"q����Mѧ�y*�"O~�*Z
Ep� eW&H��"OF$ꃆ��06`�� �:_�& h�"Oʹ�ѡܳ]��8�.,[L��#"Ov��?�D�1e�<&1�q�"O C��B.�s���%_ͬ��"O�A�"n�.��i��54�V�I�"O�T��>�nܰSLGL �"O:ѓ�)P�i^Q��ɍ�9�v*�"O�`{S[�16��bF?����"O��8�J�6LH���	 �Ȁ:2"O��@�E6���g�݃/�jl��"O`Ĩ!��114������}��,h�"O���RP�*��)�!u�L�t"O�m�F̎0n<�uf�{kZ �"OvŻc�V6�\{f�����2W"O���M�>q�Y�b�ђ!�<��a"O(Xf�J9h��5�:�,3"O�5�u�	j�V)���)&:P%"O��`pfıE4dx���kϖ��&"O���dA�7���2�]0(�\�1w"O��v�h��Ѓ'#U��ҕ� "O�E��I�<{�)"U/-�TLs`"OP {���j��  `��Fp�9�"O,=�ׂϘ9�8xiW�@Bur���"O�d'��	ؖ�rP?Hij�b6"O�i�ᡃkW���2Ͷ��G"O�P	�N��N�t�q�W�I��h`"Of R��	�&z�	3��F�{�
��"O�aV�ɢ��PH� ���K�"O�E2CJW�>�xm���.Gw��"O����Fބ/���UIֲ1s\i��"O \ʔ	
^�n�CRj�j1"O�L��C"|��L��C�3Rnu�1"O� ,��i�=u�Z��B�=xZ*}H�"Ov���L��58ș�ƇoO>=�2"O��3T�Ќ5>J�#�)/%<���"O��aj��	�Ti�ǈȖN��<�"Od	b7�L,p"��ѧ�ܕtz �W"O�yђM�����c���+j�X�"O�����^&�`c��x0N�q@"O�5��B��Q< �Z&�ӅM"d�Z"O����+��\ǨtzV��/'*ijs"O��J�T�2'����^�!�xz1"O���̊�	�h�q���/P6Y�"O6aS1�Nm�&qw
ߑA\ђc"O2���:FܱahD�L0��"OMR��=k�܊6�J�j�v@�"O8M��,�p�5��E��"ɸ�"O�H���D�Ei�JG�.�be+Q"O���A�oi��e�N��`�
6"O�D��Ò��8I�C� eT	��"O�e����4��PbDl�sEnYbv"O�u�	O0Cz�|�%��'J�	(V"OH���[�m;��h�%L�Y8lЪ�"O�,!e��\����Ć/GZɹ"O�܈2��F�t�R�#;.��a�"O���!I��u�8���ßg/����"O��9� �\�L��O�)+,a "O� �p�p)H7I�m �:�"Ol2�GG�^2�Є�G���HC"O�lJ��I�8¬43���i����&�&$~���
�s~�$��(���Ӗ-&��8�]�䬐��ϱ:��i�r��c;���-O�<�O|"47O���Ov��D拪+�&|+td
>�&��AOe���')� �D�?��Ģ��Xv�k�c��)r�����ZA�u���s>	S'�D<5@����=d�nuѶK3}2iC#{ɠ��Mצ��H����Q3@�4�����B��@�O����G��T�>%?�'B$�F0f�1q�%D>?�$�b�4D��� �⌵&o���/O�?��R�A;��u��ػ^��<���/+d��`
����L&�)"ҧ`��M2Ԍ��+$ ��P-�;T�ulZ9I��$�O�����O��sӘ�6��(�VA��d���B��i�Y���(�TO�?�R��<�H�if��4j�B��J�+��I�s�$�ĕU>��QlY�G�- �G�����I��Ĕc�ā�i*�Zȹ��Nܪòh;H�x��V���5�p$��A�Z>FL��Ș���� <`���]�a��䜶n�#�H�a�+�kq�Qf"�"�4�HDK���y_�e'�(�Ak�D���çU�4�7.Ջ~�@U�擄jF�Xe 	3~�P���* m�)�' �~���Z��n�{���;
{L���ǘo��a�Y��9��OlZ��ԃ�u�x8�S��r�Y��'����d #y�{�&�
k��m �'�
q���[�Oʨ=a�� �f!j��
�'�F�j%�-�h���IQ�Q���y�'�" Z&�[?x@C�g�'z)�s�'�,���U�7�|\�L]/R�y�'y�4�"kCo6z�;�NM����'/���W����dAfE�0,��'jvP�,�0s�0qq��N�e8^H8�'�R��0}�~��g�ۼJ�p��'�: �%f�58<�a�O�T���r�'�����Ί�U�=Y�D�����'>��.�`�h�ɽ>��4Z	�'��ٙ��9��13��	8;���'�^0 �@�#����࡜8-��U*�'E�bH.)WΠ1�	�8M>��'gx�	Gn̶$V�i������Y�'�&t���͞E���dIΠ��A��'�,���ZFU:X��!̄����
�'On j$*!%4չ�N�LPҼ��� �� ��� _��*P�9{����"OP��3��Y�Z��f�U	z�� 0"OzM�4D��?8<�\T��*�"O��k6��`�MBc�ͅPJ�D�"OJq)��;=���/;p,�X�"O�!��7~hi3�n �yH�"Or�C� I����S.D�i�l��"O��Cfj�9_,ez��j�>���"O�jE��o�V�C�
K>�zS"O�ሃdȆ?��8�䘍Q��-i!"OBD���ߤP1��aj�-,~�HÓ"O޹�t�D>g����:zk�(0"O �2�Һ�&�P�oMV4|��"O�PD'ؒo�`@	�n��80�Z"O��B��Zm|x�!��#Н�"ORE�U�ћ1�ތ��J̲�6���"O"���h��k���:�L 5R���"O�A���w�A*�o=�0��"Odl�4`I}
��
��y(Z0��"O�1ˆ��`�����B	h22�z "OD�cu�ځ-��4 0aґJ<`�"OnY�D�/�V��בr
:D�`"O��X��\�	�ҁ���(p   �"O�-[`�݅a��2�J氨s"O���6��*c_��p5J�)���P"O����9�l q0jv]P�"O�5A��$JO�Iqc�!dZ���0"O�1¶Ҷbg�,��A�$\I�\ˤ"OD0�A�S��� ���]5��z�"O"ic�I�1 �Y�,�,�m�B"O���X�M��i��i�3av�4xf"O
����;@ob���G /l\ր��"O� *�d�Y��F���<��mQS"O��V$Z*��B���v@J�"O��!�Oӗr��������l3va� "O����Kb� @�ŉ�%yJ�� "O�,�PI����HՉ�EbXQ��"Oĭ�f/�6{��5s�Yd)N;�"O�|s�RI�R�P0A"��"OJ�9�&��P��4"Q�+ x3G"O�}k`�R�RU*�!�;���#Q"O�=�dC	_PT	S%;4����"O�$���١l
�%2�̿A&U��"O*d¶�Q3Ҕ�"`�>&�=IP"O�I{G�3�q��;! ��r�"Or��GHV:��B�Ǻ'��A�"O��5I8e�Z�3��~�,\�"Ol�� ���
\z���9���	�"O��!�ǹs�>�9w�H^J�Ū'"O��@ĳo#ؼ@�
^C�$��"O��b0�W;��p��w}.(�D"O@��"�ɒr��!��3_Z�M�C"O�`Y0�%[{����$o���Q@.D�p1��СM�|�a�C��b3����/D����A� Űg�B�I��{%c9D����ə!H/`��pg
$�DYa��8D�\ڳLE^
�|�tF�"E��
�*"D�d�2���7��$� )U����("D��Q�]?j!�WD"j�%x�.D���cc��h���Ui����d+��,D���gC�+y�4SA�v�[$,D� 0%ɟYApD���٭Bt2}�s/=D���5*�qy�Ī��53���*Ӂ(D�x�5��lp�MyЇ0M �ZW�8D�� ʥj���Eo.�s�%J�8<�"O<x���1"�aA�
��9��qpq"Oa�C˝�o�FD+�AR�"ܣ�"O��3�.N�Qp��� 6.$Ч"O>��lO�@���6 H��)�"O}6�Ia
��!��/�JA��"O�\�kɡkG��2ӦɴCKb�{s"O2]V���L���$UK��I "O�Ƅ�F������;e��}D"O��1�M5�*�Ǥ[m*]��"O>�h�ص?�X�9���!-x��h�"Of,I��@h����#-\L\��"O$��`�%E�@;��уpH�D�!"On,�UhZ�kC��H�ƕ�n6��"O�Hq ��;s,���E��k$�j�"O��[dC�ݠ,!�@\��r�"O�2$��eI���p�T�$��QCC"O��ҳ��*�͚wɔ�d4�<j�"O,�ZN*ea^a�����=��Q�"O�t�S�vyf��牖�{�V�C"OPPЇ��H���R/�v��"O�z���^�)�w�ǀf'��
"O�
�H*���c�b	z2��@"O�u!$��!g<���G��t��e"O��(T ^�t����o͉1��h�"O ̣��,�8$N׭&�H��t"O~��$E�-+��K��_�?�	��"O"�8�)�)8a�b7�΃p:�Q""O*�C�A�=�48�D�;B� �"Ox�J�B�2
�N����t��YC"OƐ�W?(@>\Z�ޤ�l��y�F�h�!�ԋYC:84
@�y���4?������W�MCS悫�yr	C�$��˴c����]��윸�y��'�d(���^��uz�ꇝ!�D�P��i�W��]Z~�(�	�!�$߂ �����D�##Q@��)_!�G�,U�]"t�D��l��EJ��T!�Q!���`ĩ��L�Ԥ�b.9�!�dڈ&)Hsҏ-I���;�&{�!�ː֘0r f�n&�%#�OD�!�$S$+��P��V�F|�5P�Ͽ8�!�$ƬJu��k���Q[��pD��9m�!�$�-�p] �HDZ��!��bH~P۳f�P1��8P  pg!��= 8ᓆ!�2� �R�"k!�$Z�f�%�N�g����Q��@	!�$���Ȅ�FªP�\�s&��76#!�$F�4�\[�ז����ԇS�!�$A�gL	�Iܩ/������G�{�!�ė
o&��s,h{��)b��!�d��S�F�b��`���d!�K����#jO���\�� �>y�!�Ě�O4�m�$u��hT
Ǭ$�!�H;Z�(�:�eA�-k���ܞ-�!���o���@T�oL�k� 
xq!��"Y��	�#��7����,f!�D5��q��D�H6�%�GW�N[!���5Wx�
�J1?lH�e�V!�V�'fڕ�,�=sPt��n�,�!�ǼD9,�AnR�7���g�>�!�Dڅ8-A
�Y�B��%��x�!�$�?j��I+���L�$�� �ݘfp!��ҺH>���C/z��ɕ�_k!�� ����ՆOJH�A���<OL �"OXZ�؍+�5�&T�#(���"O��z�`
�~#D�#�$�`¬�z "O�L�a��Ǣ<�g��d�ޙ
%"Oĵ�G����P�9�00��q��"O�hc6/�?1����J�Y�҅2�"Op]��/�0���#c)˶ELt�s"O8����ԉ|{b `��V�9S��Z�'�R���F��T�:Q1'L��$e(�
�'Y��z�/V!p�NT��hZ�!���'�DEbwV�4�H0��♺D�RD��'�����\�s�L���H� Dz�'��bQ,ע��1Q���x���x�'�h��(B���F�C��h0�'�6��REf���g/�k>��'��Ŋ϶D�� ���ҁw��@	�'���Ԃ	גYQ��Y/��T��'���Q�+=a��X�.W�+n��
�'Z�|sDf��s��hß.r*�	
�'�~��#ڸ57Fp��#� dR�X��'�%�&#�:27��S��_S�-��'O���n]��@j�!Ef)�"O>͋G�Dm�i��dM!p����'"OFL@�b�=B�`��f�� ~^�&"OLuHP�0���$Y�\�k�'r
����փ
�����(�	�'H�ܨ��E�#g8(Q�Mc�����'���-ـ_�Ѻc$mӪ��"O���ӥT6����D�{��("O�X��-Y�I����E�W� �H"O���a��C�4,ӃN�a��(u"O�(�@*�C'��z�L�HW�H��"O:�p�(U;nJzQ�֯�14Z�=�T"O�P����43�p:��/X����"OH�OH?CF�@9��O�VT. PS"O��s`�>U�ԣf�\�B�� �"O,�Su��=+̪�@�S��3!"OX���4p�T�Au 8Z͈�"O��aLQ�V�tYqM�=��R"OJ��K)�6Y!q��|�
1@�"O �I�P0H ,8;�Ӑ:S:M�"Oν0EN������^T�8��"O���A�'&!����i�9m`U"O�,�Ge�vH�����^�PȆ"O��Rg㗭����x�$�u"Oɱ֢�'H�4A�c�����"O"�A� �5 �*AH�ݖO���A�"O�I��͛hNx���K?���6"On]c�	   ��     K  �    +  �6  �B  N  ^Z  -f  �q  4}  e�  O�  ��  �  ׵  x�  ��  ��  !�  q�  ��  ��  ;�  ��  <�  �  : � ; � "! s' �- 4 ; �A H sR <\ b �k �t | B� �� S�  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O��jg�=Pz�Aa`�#�h��!\��̇��#=B8#���fB8%pS��H�����fȉ'�$!q!c�	^+F b�ǂ!3�v|��'��EK%�ݵXF|ԲBER�/�f�ٌ��#�
ّ���5�`��'c�6vH��C$"Ox}e��N&}A�A�3Z`X�"OJi1�Hճ,U��I�	� 4Ft��"O�D�tkI:��͠�(A�Iddi��eOuH<YS@҂+2��p�T�w޵����h��\�>y���BdlcL
�g?x<����d�<7�5�)�늁yD	�`��J�<�"]2����ܿf:����G�q�<I&��d�ɓq�:Ρ����X�<񥮀�8TΩ���y\^P3�N_�<	BdJcV�����P2.�"�J�,�v�<i��1i��#P��,+=hR ]q�<���	4M\���#���:�����o�<i���3ZJ���5Y�%ԞU��g	h�<i�-
�Z����&��U@�ɱF�DM�<����+�|�h�O��i�ʤY�h�K�<����u�
� R?
Kv ça�<���.-���4��*��ZVŀY�<��ꈍ[����Se��e:��Q�<�%��$f��F�S�r��TeXX�<��(g��K�GįDlz�iU��P�<�w(]�>c�r!�*8`9K�"O���T�W���!G�Q�R-�"OHXB�X( �i#B��)^i"O"5K!h�5��В��+B
p�Ia"O��Y�Xr�-���,�ِQ"O���j�"�U��-�~��"O&���Ǚ7�l��t,�V (�"O�a 2]`��:G���ya]�&"O2K��ƹEέ�F�� F��QS"O�%�⋖�s�J�y"nԵ'��ۣ"O�Yk��z��i�`�@�p��"ODY�̙<RE��NK�l/2!��"OJ�jv�۽;�P;"�̼#j�P"O\I�/���Y�	I����q"O�D�$j�4F  �H1e��N@b�"O� ��
�/q:��W� �!��Ժ"O깚��
=%dU�f��3���7"Oba�6� "j0]H"�sΑJ�"O촁LTf�䍐ANL�r�4 T"O�LU�]�FP���2�xX�!"Ou���]�9��]ao��)��"O
�H3 ��Y��Qo�)I����"O�u�wƓ-r��@�7c��_���"Oz9T�ȧ&u�h�IK��< D"O��!�5�6���\�f�"�"O��k�eK-fCu����:���ar"O� >��sc���5S��	�C"O���I�8-��4�nO�G���"O��X �].8pw�R�u|�#"Ob�[h>S`�b��C"4]��!"O"-���[T�]!u�v%���Ĉ�?����?!��?����?1���?����?�C��J$d�bbT*v B��?���?���?��?���?y���?ٱ@�&i��(^@i���ز�?���?9��?���?��?����?i�f�	2J�x+�QEr�5����?���?���?���?���?���?���)rev\IQo�Z��=��2�?���?y���?y��?���?���?�� A�7{��9��+X,�ᑓ�?���?y��?����?���?I���?�jȍaBN��3�N����S��?����?���?Q���?����?����?��BL�`\��ߑ�v +p.���?���?Y��?���?)��?y���?��ᖚ͜�C�\�mHP�$�?���?��?����?Q���?y��?�U΋�@�Bi@rdݭn�����A��?���?1���?���?y���?����?���<��� ���m�BE�CG��?1���?���?����?����?����?AR ��d ʽ��  T�6��'f�+�?���?����?Y���?)��?���?�֋Z.1P�u�#PR��a���?����?����?���?��dQ�6�'
RgE/\\PC񋄇6\v�{�eN"�Tʓ�?�)O1�����M����]xb�� B�av@ ��ŕ�P8%�'2�6m&�i>�I��q���S� @p�f5�T���K�����	3�Pm�[~?�ڱ�S}��[�#�d�b��-�,��`�1O.�D�<���IĆz#B-��N�:%��y�D��b�&�lZU'�c������y�ǔ���1��D	7�����J ?2�'I�Ĭ>�|B�E���M#�']
��s�R�F�>e�㣕�m���'�����6�i>q�	�9k& �`��a�����+t�J�IByғ|��w�|�kv��n�����Nd18��U&���p��O���O6�|"�Z6D��ؠ�TU�#����Ot�����G�1�t���G�J�$�(w��x� $�<{�v=j���� ����O?��6fH�ً���y\�a����Z�牱�M�&��u~��yӎ��Ӱe�p,�'e�Np����42���ҟ���� Ӣ�
����'��i��?-��"M�SD�K�D�2T��h��?3*�'�i>)��ڟ<��ٟ��	G�9c��*H6��A�F�]��P�'�\7�g4����O��D4�9O�)��L�e�=�"�Hqǀ�<����?�ش2r��T�O!�t�ϸ!.�
�A�:_�:ӎ�) ��R��By�l�3��� AC�8/�Ɵx�!dʓ2�r��M�v�"$�O(
�����?���?���|�)OFqm�)z�r��	!��s�=|�j
�NC D�J��?�M����>9��i�7��O�uʒ V��q��o��5@�iM4x7�v�l�CԦ\8E��$A.�i�	�?Mj �S���nϨ{���h�A]�n���H��d����ȟ���˟ �I���Jg�̊&\�c��NF��5JE)��?A��?��i1���^���۴��S��2��	�0"cnL�c��b�yB�i�,6-�O���eӐ������ך���b�	B�+��@b��)r".ͱ��'� Ȕ'��7��<���?q���?��M��A�}p��Q�:�.L�֪���?	������ l�ȟ��IޟH�OpA������,ѢJ�j��ON<�'In7����%���?�8�h&�,5�N$yn�`C��3�I��N�?hl�'}�֝����dy��wa~����Co��!J�@ ̀��'?b�'���O��	��M#`o�S�k �%a�AXa��j*�+-O|�oZJ�g��	�MK�/M�vK6��T��:}#�< �B�I����'.��Y��iK�$�O�-	 ��1���@�<!��8]jV�����;��=@pE����[���	ğ��	�d��ϟ�Oz`%
C��t�<�:�"V�l|J��q�8����O^��O����|�4��w�����:V�\E�6	]�OS&�z"�O�6m<���I�O��6Mb��jP�sG4�"�J�d��#���I?��X#�'N��'P�6M�<a���?q1�����PCP�����K��?1��?������F�J��O�|���|*�I�q���kH-��2dK�C��$��	���o�L�ɞW���Ԧz�\8Zӈ$���I�h�7�Ŋ(.��AB�ULy��~�͐��'�X��I�F7d]1`H�U����T�G�=�e��Ɵ �	���Ic�O�R �OOz$��jS*�3��I�:��Z�Wo�I=�M��wLz���
(a7z�:�E��@J��'T���g���U6�c����q�"x1�O��̉�l�AP���tL�&N9FE�&l
Ny�s�:˓�?��?!���?��?*�6�o�Ā���ܫMr�)Oܙn;�\e��̟<�	w�s��kT���W[�����K��� �������ĝ䦅iٴ���|r�'�?Y _�(��G�;�dܡ��D�+���Ӈ!Q��򤖺_u��k�Fy��X뛖T���r΂;`��t�M0�݉�E[����ܟ��	ϟ�|yb�k��5K���OBl�&i��/�6	�/�9'� 0t6O�Qn�f����I �M���i*��⠴IQ�$���0��,ɶ8�q�im��ݜ�`�����B��e���MA[N�� �s� m��0⡈S)~v�h��4Ox�D�O����O����O�?]�it,��M�	�E�WcT՟����l�ش�Ĉ�*O��l�E�I|��@ o��Y.f���XZ���%��[ٴ@���Om3E�i��)L|��Scg�L �0��7	;\Y��j�0L��i�ЛÂ�'���'@"�'J��'�@e���R�fR�y��#R��S��'�Q��j�4�d����?9������C$�r��#|6݉ jH�W����'���w��v�a�T�O�"^�������T�k��C$
9�U��1�@}h���oyb�w�}��'����y��Y�><4
TD�[D��	�'���'B�'�bc�<����<�'��Zj��Mz<��'�[�7AYʅ�;]^�ʓ;�6�'��'�r�䛶�ͣ��D9��/'N�`�,̯e+�6��O�p��`ӎ�H\L�xd��r,OHx�#�F��Y #�������K�צ	�'�'h��'�2�'	哵u}B��j�.T�P$	���3����4_\����?���:.��A٦��:pz��%o\�;M���7�ˑu$�q����M+�yJ~R�"�M�',h�ٕ�-`��9  ��$#*���'��FPޟ�H"V���4��d�O���ۓ¼�����&�A�h�8���O���O4˓Z��G�����'��$� Y��L�I9���C�]Vk��|Bͽ<����M�I>�7��p&�d��I�����u�x~bMS�B|2����H)R�剷�u�E�ݟ�"�'F�ԁ߳~��HsǗ (`�4�'^"�'4"�'Z�>�]�q�Q�w�5Y ���Ь��5�����M�U�
��$Q����	m�i�iA,�J�2D ��;�4q@�H��tnڐ�M���q��ܴ�y�'q����c��?u˔-W<lN%d�݃x�\q��Ԇ��	6�M�+O2���O6���O���O
�3r�U-��9���L�q��L��B�<��i&����'F2�'���y���;x��s'��g�9g�@�wz*˓�?��4�����'�?���$�"�s���SV(�N=�V4 ��.��Dѻj��;��H���B�vP�3cƠV�j-!��:��b׀���'�R�'k�O��	��M[1�
�?	�F�CX�(ŅVyH0����<ѣ�i�R�|��<����M+�SS܄+�`Ʃ~n�^ x���R	�9�M�'��,B�{������S���1�u'�w�r�8Aj\G��hs���0�
��'�r�'K"�'���'��e���#=<� �g�^�R/D���.�O����O�MoڤJA�-�'�7��O$�*܌�wJ��tOT��ˊU=��aH>	C�ijj6=�@1"��t���*2��D% H�q�k�o�d�{�`��]W*������$¦��'N�'��'̒�Ӑ`@4T���C�m���P"�'6�W�Hr�4K�m��?i����	݈)��黦D	f2kMPX��Ot)�'�p6�̦�'����?�	&�@��)��
� �L�;�NQ� ���R��#a�"��	=2�����q�\�����k�A�A�XiS��E?v�>q *��?a���?���?�|�.O��l��8x��������ѓc,���3?��iI�OLL�'�6m(	�q�4��Q�Lsf_(Z�n�|ʑm�ݦ�̓�?	���!�V���Y~2���rD�۲�M>R�0�d��6m�<����?����?Y���?�+� ѐ�K?/��p@1�fK����/�¦� %�s�L��� &?牍�M�;d��ͨ�IȌb��6k��@��i547�9�4�N���O��@�goӊ�	$��SP�Z�&�(2"�9a*��I������',���'�6��<�'�?�����4��%���B	V��?���?A���d�5j��2?�����:A�x\�8�e�%��Mj��k�>9%�iq6�)�d��6�2�H�U�6��(ՙ=;��O6�r�ƈ@�����,B_wD$�ɞ?rb޹h�t�ȴ@�ԆhcՅǨ2��'B�'`r�ȟ؀��D5x¡��\������ϟ��ݴ&e�5�'Ƥ7�7�i�u�P��^m	��M�eki��㶟�n�M[�GV\�s�4�y��'���t/��?i⠥��2��	��� /T����JRS[�I��M�*O�i�O����O:���O.b��V�G7]R'f�!i��C��<���i��A�'���'���y�K����M߮{6@}ځj��FJ0�M��fgt�F�O�I�����= ����e��#`p�A����8@*E�s��k�I�M%��$�'�0��'z47�<��2&L�\#�K7.xޜ�ũ��?��?��?�'��D�Ѧ���i���`)�&2��d����32�>f��1�4��'���'`�6�|����$	��P⑬�.6@��1`N'NuN�0/f��:�˔�I�4�~"ù���NYIe�	��S%.��yj���OF���Ob�d�O���5���vx(�E�^�~��,�bϛ�#�������I?�MӦ��}~�����Ob�YP�X(MT����B�S����UO'���ŦѪ۴�?Y�n��M[�'�b�"h�d	ԈX%M�4R�nWZX�!��Nԟh��^�<1޴��4�����O��䚂6��h��' l���kQj��kG��$�Ox�YT��J��y��'��X>u ��V2*��}���_�V�E@%?�q}��tӺ�l�p�i>���y�*�ce�� [ K0hW�:�0���o�^Q�E�*?�"���|���T�˓��[�"�9ʂ�I �qeb�*⧟?�?i��?���?�|r.Ot\l�
�;�MO~��A�s��bD�Aqy� lӨ���OdhnZ�5o`�cWl�,FD�O�"�~Y��4P���f6O|�	#\�J�(�"�վw"��$��� �-�cg�^ۜy�gA��hĴit栗'+��'�b�'�R�'h�'@�N�eT�ٵꋄp.x4q�48Yٹ���?������<7��y�
�����D@'v�Za����6�ԦXK<�'�"�' 8zy"ܴ�y�˞(*h$�Ө�r��t�6(ъ�yҢF(:�`e�� k��I�Ms-O����O��2�
�A�ЍA�(�+�K�OR���Od�d�<�d�i��0��'
b�'@BM��`5���.V���2��'!�'y�˓�?�޴r�'�Sǀ�p�^yhw"_+pY<屚'2镍wRܨ5��	W��.�u'gM���p�'��ez��:jn 9*�g�N8��z5�'[�'\r�'��>��2[���,��'�ܭQcȖ�I��	&�M�ܻ��d�ɦM�?ͻ<T�%�,E�4XN����Vg�&`�̛��k��oZ6:�\�lZs~�ݧ'�.q�S�D��G�8W�X�cꍸi�R`DU�jٴ���O���O���O���:�
��	�qNV8���
"�VʓLe�6��L>��'	���'ʄ0��Z)�!B�������<9���Mc��|J~Q��!��A��fR�H���` �
#�(��i��$�ph����~Th˓�vS�����@�8k����_K��Z�kZџ�����������Dy)p��IZ'�O�!	�ϭA�����J�t�U�F;O�n_��8��I�M+ŵi˒6�C�<�����b�ZX�4@V"IPry�akh���ΟJ�Kʸ:����Gby�
q���Q�`�R�V�5Þ�P���!0��I柤�Iȟ(�	۟��I^��XF��IX���`�ƒQ�m����?y�؛���7-���4�MI>�w�>W���S ��!y&�L�zV�'�R6M����� $čl�g~��
#�T� �8����!�Z"�t䪴��֟0�C_����4���Of���O����'0���b��.3h(A�EI�&����O<ʓ=כV
 ����'8�T>��Æ�&�)��Fؼ7֞L!V�:?��]�8�	ݦ�hJ>���?�gQ��xW�]((~�H�"�p��X��^�wKV��'f��]'2ReKyb�w����D�E��@+"��E4n��4�'���'�b�O����Mk�B�)CP6��ߊ$H>��'ϩr�Ҝ",Oj)m�_��"H�I�Ic#�\+*�T�Q� W�����8�M�T�iJkG�i��D�OBUq�"ɫ����<Q��$-	�
�5�<��RE���R����ݟ���ٟT�Iٟ<�O
F��&��N� yȀ��C!6I���cӜ|��9O���O���$Z��]�$�mޓu������UX�41A�FD=��J�"6�w��#$���r�l8����-x����$�|��+g�)K1��	K��hy�O�� H�6�-Q�9�"(��A��?���?Q)O��n���	ʟ(��#?QL���O& <I�F�q�)�?1^� �ݴ\��i;�D� �`���E1�X�:�Fį+�I1$6�q�6��_
�b>���'����<!X��A���f��!b�G�]�����П���H�Ip��y�E,B�Vb�#�H�v���D٧QW��rӐ�p���B�4�?IN>�;|�0H��E	�i��$JS�ۇP���kX�6�r�b�mڜ<ln��<���2ty`��.Hಌ�'M�0m1t�מ��	�BJ��䓙�4����O����O6��, �M�'�yuJ�sE�s��L����2���'�����'1rD�2n�7���z����`	�S����4f�f�7�4�6���:��A�.D�xqA�ƴ�X1t
 b`�����<a`��)3��� �����G��%K����N�A$�
Ae���O`�D�O��4�d˓UM�fŞ,2=2 �Z���ڭ5�&h)��	��yr�q�|�`�O�HlZ2�M��i��|�q� ..�H���χ�4��a,�/R��1O���^" a���^\$����;S]�L(`C抍SU@к3����?���?��?����O1���<*�����L�^�ej7�'��'��6픔T�b�8�֚|ҍ��"��X��Ӑ]Qܸ��OB�q��O"�m��MK�'OZAQ۴�y��'��*b��;q�8�&�c�\�!�6p~>��ɒ&�'x��ɟ���˟���3<�0����( _�؂� 6�����T�'26�(C`���Op��|��H���zh���ukr�kCm�l~�J�<���M��|�'��S���/��i�`Rtڵ:#�ɢ�.ycq'��S	<0q/OB���?���4�D�w�Zr̓1Id=@i��8z����O��D�O���	�<���i V��$A�a�x,��i�1��|�^&^K�ə�Mۏri�>��iB�3 ��+v
�!Ǐ�2/�d�� t�r	mZ#N��Qn��<��rBH]Ac�y�-O��x&��G��i� �U�>y��as4O���?��?���?������O�48���L:�MZ�&���m�h�@1�Iȟx��u�s�������JS�6� v�
�͂Q�������`ӄU$��S�?i���#yv�o�<�I�o�0����4��
�<�VNн2��dL�������OT���ET�xՁ^�<n�@'kގE-&���O��d�O�˓+8�6���B�'��l���'^��=K5�;�Of��'�6-Y¦͛O<�ਘ1gR���񎉄*�4JϤI̓�?��p��2􌙕��u3�iV>�� �1N����A4��`@2���Or���OJ��'ڧ�?I��I�	.��� �R�@���H��?!�iJr�2@Q��H�4���y'狇[3��Ek��t�)�nJ��y2j�� lګ�M�TИ�M��'T�.�(ά���ۀ �ၧm��]� ��ٳ�ᐵ�1�d�<a��?9��?����?Ѳ.�:�xi�BȴR�.��� ���Ħ��@ܟ���̟�$?��4'4P:��:[��A��	�+0�r�P�OT�n��MS5�x�O��D�O�>�J�i�
g�0�r����b�����9���P[�x��"�1i��BQ|��py®]bV0�DlұUN�)��ĝ ���'��'m�OM�I��M���J�?��L�1��Q"TeĢ;k��!҇A�<�i��O���'W�6�Lަ�Q޴<_fAS��f��5��[�5a�	�1HO��M��'2B%̧Z���S���?����4!9�leYU��9������Пt��֟��Y���6�x�mE�8����2F�1K۾�k��?��4]����q�I �MsK>�p�#L�%PrM9Z��"g!Ѱŉ'46M�Ŧu��(2pt�l�<!����1�@���H��b�����\���H$GT�$9����d�OV��Oh��GwB����11�B$�DǞ��L���O�ʓc@�栕;���'-2_>E@g%v����Fό4��(���O�p�'�*6-N��ipO<ͧ�
�А"���&�Gh�k�I���:1`Ơon��*O��C��?	p�"�D��|2�a�@lOd�<J�$4����O��D�O`��<�i����N�ʔ�qW� 
̼�q�'�<!M�I�M{��Π>с�i����Έ�V�B *��"$쬰�ha�Zm0p���l��<���tD(��&��	p+O�ӓ��t�v$�5��+���3O���?Q��?����?����iX�4�DjQ���IJ ��ei��?��Ml�,%h<�I��\�	r�s������37�͝C$���
�B�5���33��v�`Ӌ#��ɞ4u�7q�7nJ�-,p��"F�%��3�
w��b��'Nb�	my��'���
��8:]����7�]�Z������?���?I-O��m�/x%�������bTN�Y��r�N��)L7{���?iA_�$@�42�6#�=BR�@�h�*qRmB`�!n��OI`�~1آ��<i��jXp�D���?�Gd���������4����?���?���?э�	�O&0���^���Q�gS����Kg��O��o�v��d�'�6�8�iޙ�VD[w1���r?�J�n��Rߴ ����|Ӧ��եj�<��.<x�$���hc���"@��1&M� �Byq�O�䓡��O����O�$�O���T�,��ъ�c(�2��0d��uh�	*��G�!�'���$�'_�� �R�7]�Y���H�����<)���M{%�|J~����N��j^�BL�9�l!���p�ʗ:��гU� H��S���O,ʓ#�����j-i%�Ò:h��?����?9��|R,Od�nډa-64��5Nl���� ��@R�D�"��I��MC���>���i�B6���q��8��T:G6h� ��CpmZO~2D�#���ӿ<%�Og��>��� g�Ӷmo*�0���y��'("�'=��'���)�-����p���I� C�3��D�O��$Ԧ��BFvy�v�ΓO�<(�×1���B�*	�MR��:caJC�I��M��i���~���>O��ʃ:tE["��P��L0SQ�yQ䴩B�4�?!�i#���<����?����?�kSS�]��GԊr�\uZ@MT��?Y���D����(�#O�t�I��8�O��@g��$�!�B��]�v���Ov4�'�t7���*K<ͧ���J�4�n��&K>�x�����a�3Ǜ�Tk�ԁ+O>�I��?�Rg'���O0�r&E�&�[� ��5(��$�ON�d�O����<�c�i&�̈�M�2��]�%ON]=�<��"h���MÉ�O�>qҽiV�ܠ�E>N�e��I�&� �9g�m�t�lZ�^BL�oB~"�E4O�Y�S&��ɣa�J`8���~d��1�ȧqTX��Fy"�'�r�'6��'�r\>���eųzD�� I�70�|8�f��M�ń��?���?�I~�?=��w���&��Z�{ .�*��i`�zӚ�nZ-���|B���j�͊��MK�'��97ɖ!Gj�(piڪ=La�'���	rϟ��3�|BV�����ĉ��)aFЉb0�\.&
��*�ɟ �I��\��Zy����d��O��D�O����?ݺ��̈�m�v����;��2��X�����4!��'�����mx�X&��gmP���O� Z��R�.�*��:��^��?����O `!��'���ʓ]���1���Ol�d�O��d�O��}λ��p	�͍)�12�"�S�B)K��k�6
��F��I=�M����Ӽ��/K���afK�kwB����<�q�i��6mݦ���M�����?�F'� O�����e�u����;���p� �|~�-�K>�(O���O����O����O�YZq��y���5EEaX8���<�g�iR�E���'���'���R>�,A���9S%^(w3rP�P)�E�R�O�o=�Mc��x��4��/mdZE�QCZ�2���$+�'U��*��Փ?t剮l�PmK��'Q��$�|�'�t��e'G+\;�eLR-x�|X!��'b��'�����R��bݴSV���A����E/[N( j�\.k�\�"���'��'���ӛf�|��o��{Ϟ�y��^�T��lr ֟SD���HC�����?�qjƾH���������l��?pa�Ɲ?M 9��	BS��$�Ot�d�O����O���5�S�h� 3`��iz{�ƙ=��}�����ɿ�M�6!����ʦ�'�r�׈9X��"��	�is*�z#C� ��0כ�imӚ�)�t�7a��I '�z� 8��TC&��D(���^���aRcG>�?���&��<����?��?q���{��	�&�/2�%zȝ�?!����ėǦC����	ڟ8�O�m"��%'|���A��<���r�O���'װ7m����M<�'��7G\-OgJ����Z�'_0�)�șYs*����/C��u{(Oh�	߇�?���)�䓯K����,<N��D���(k����OF�D�O���i�<q�i+V�z��;��K
: j̘ӳ��>w	�I�M��K�>��i�p���Ö:m܄���D���-X�cg���nZ`�>�lZ�<��:%pҦ��ص�.OJ؆�O��i$S<#<T��0O�ʓ�?����?I���?A����<*��sF�ֻd�D��$p�j4o�=F�K�OB���O���$�Ȧ�]?1�����7C��[�FU�u���	۴����0�4�*���܈Io�,���hL�WA�#$�r�C@��(j=��I�xb�Zr�'��'���'��'���U
��H1�4� G������'�2�'�2Y���ٴYY�PΓ�?!��E�L!��ϳ<���y�Onx y���>���i� 7��o≉;{�٢D��$|�@�D7���蟬@�N�Cn�sè#?a�'Q�$�dP��?�@�&Q����\n9��0s��8�?Y���?���?���9�����R�0T20�qC��R!�\33M�OX�mZ�Ssl��'~�6�4�i��bC~��E1O�;�.Y�r�p��4,&���nӜԺ��~�l�Iğ<���m��B޹N�4m!�fE�o2
l)`�K $��&�x�'�2�'#b�'���'�V s�ҝ>W|��g�ڒ'��Q�]���4w��8͓�?q�����<iDgE�_Cn�	��E o>L �g�H�>v�I �M��i��O1�t�I��
�b^�����4�sDO
<_�1S���8h�pRL�r��Uy�ДR+��C�&�wmɁ�$u���'q��'��O�ɟ�Mk ���<1��")���q���'(��	A�I�<Yſi��O���'�ҳi� 7m�>"�=��T X��Sa��&*�&� ��o�\�I��@��xu��L-?a�'���ݱ_���#�ė�47~�07�S�<���?���?���?����؄v�-�3��>�`@�^��yR�'���v�@�J���L��4��Y'� �oZ�,�*���C��$��e�xb!g�B�n��?��������?�u�F����`�4;&h8*'e�2���p/�OM�K>1(O��O����OV��ۿ-���PC��$�f��G�O>�d�<d�iJB5��O��D�|�h،B�)Ď0�r)j�E@~RI�<���Ms4�|�'�.Ll}:w�
H��r1�_!Șm�FC�'l8,y��i�p~��O�rx�	�a/�'S��(�*�Z��U2�I�A����P�'���'�B���O���M��V7
܈��)TQ��qyC�����a+O�n�Z�W��I �M˳䚡G_8�bCt�a��7J�F�k� ݱ4 l�8�I֟$�b�����my�!�/>z���$����q+C!��y�Q����֟��	ԟ��	韼�O16�;���V.h0�q�
'M�i�t�|`Њ�O��$�Od��������W�����$_.��&��)iv�@X��M�ě|�'����j�Z�xٴ�y�b�(V�Uk c��^������y���(���I�'�IƟ�I�fN��i�薏.�N��a/Q�P��	֟��	˟��'i�7���R&^ʓ�?ѣD��f�j``���E��h0Ц��'��V���x��'�\صfV6�H�jT�B�V���Y�y2�'���0�ܱweddtU����q�@�ş��!�7Tk�!)´q� �#ҏR�?���?Y��?��)�O`�)F��2�U4!ݏ+��9���O�o�=d�$��'@�6�;�i޽���߷dþJ�C�z����"l�|B޴t���~����r�d�t��🬻��M6o*���M�b�9/ٶ�a2ؽ'x�l$�x�'�'�R�'��'*��"���.j�M��
*Z�.�#Q�ly�4Z�0����?q�����<i��ߚ�$���Ǽ�ܠ
����nN���MK�iC4O�i��(�	K0q,eb5M����`9f��V{f��Ґ)�%��$�{V���V���OZ˓)�%��՘-4֭#��P�bx�J���?!��?���|*/O^�o�`�\E���_`�Qf��ԁ`��,)y�I��M�n�<i���M#ӻika�k�t�",P��1\�P[����=��:OH���'��4���N�˓�j��_�����E�}o<1:d���bo�D��?��?���?Y����O�<�@a�P-Qʱc4m	r�4� ��'���'��6I���˓P�&�|��G�?i`�(B�S�}�ëܯa�zO�n�+�M�'0_bQy�4�y��'�~<�3���yAp,�F�D���p�'Xi�����A"�'���ȟ0�IΟ ��,��)��EĂ)�E gN��jy��ǟ$�'�J6�-^�8���O:�d�|B��Á��u�P��1N��0c"Tn~r�<)��MKa�|�'�j @K�	֩�v/ǵk�9��H$-��c�^
/�@L�,O���-�?�1�:��O�=���*���yANH!����O�$�O���<q2�i�[��I:������B4?-ȱ34�4Eo�I��M[��<��4�B��5"��L��&�A�x�A��i�B6͒�[m�6�$?�b��O�������^u�`�4&p�Q0�E�_`�d�<����?���?���?�)��9(���+H�L��6v-捋�̦}BvL�������L'?�ɀ�M�;'�Եт�HO��9���%{��r��i�6Me�)擝Aڜho��<� ��*5`�7M��c���t�4�8O�xk�HJ:�?���$�Ī<9��?Qª� 7p�ke�/��vO�?���?����d�˦�sr�ܟ�	֟ s���x;G�F#+Qqi��Kr���O��l���MKD�x�c�A V�X��Nu|L@RI��y�'_A`��7�	Q�W�d��4��Eϟ�6m�KJ]�ס�UQ���W���	����I۟�G���'Dq��ʬ��jǌ
�a�2�I��'��6͏t�˓y����4��Ha��؜MH)��gQe�&���O�6�R¦Y۴d�r���4�yB�'������?U`¢ޣ;�~aţP�0�t��dAP�vm�'��	۟��ȟ\�I ���LP���t�G�Axʨ�a��ה��'�z7M�$#j ���O^��5�9Op	{b�W�|��̹v%�=�l5$	pyr�''�&�9��O��t�O�l�qSf]=ta��"���$�	��r�ֱcR���V#��U.R�X�y�hF�_�daS4�'���т�H>9���'=r�'F�O�剩�M����?Q��ۘ�:,���S��h�U�<9ָi��On<�'7��ܦ9kߴO��]2�eI%E����R�X|�0I�M]��M��'f�&�J����J���?u�]J�P���j��`;�-C�)��}���	ʟ��	����՟��I_��ܚ�{�n�{�d�1��	TU�}p)O��d�զ��U�#: �i��'�Фs��
���s���!̰���i-����1���|�r���M��O"���D�*C��a�K�Rd��֩_y|�R��Ox��?a��?���DR�}�-L,4�t���*�xlř���?�)ORm�_�����̟��	D���Xb,д1FIDT�Խ"AL�����H}B"v�>o���S����3����g
VZu�`�BOFJ�2��зMZ`���T���A���C�oD�`	$��F��	��N2Q;"!�	ğ0�	۟�)�SHy2.|Ӵ�U⋉���P�M��)��G΂s$��d�O�	m�|�@����M��eǅ�l���'r\���@[�fu�6-���o���ퟠ@A�%#�ĮXxy���H�����}�
Bt����y�\���I��X�	埸�����OÒA�k�:E�V���Cj��9"�~�T�b���O���O��?i������,��E`�u���mт�)0Mϛ�fl�T�$��S�?����E(pn�<Ir�ׅq tCF.]-�f	���<!7 7j���D�0�����O ��u��1�J�;S:��	�+F�V���OX���O��[B�ƫ ���Iß� '� ��y���ƹvŎ ��Z��x��	��M�c�i��OH����$��0�QBZ%ei6���8O@���$����!��������O~$+�o Q�BaD�jH]ef�*!�Xr��?���?a���h�*�d�%���{�K Zn�@ #�~���i'�My2�oӊ��]8X/8�Dc&R"�d��	����8�M{r�i�7m�u��6{����=A������O68��I�*f60��cг� AH�&@Q�IsyB�'���'�B�'�N�-A*��6Cɝ3��s�L�j�� �MC�.ֳ�?q���?�I~Γt���� T<hNP�/$%�4���\����4>�&�=�4���i����S�eP�B"�	i�<���V�]^�>��d��<Qv#�y`�������Ł\�f���FR�}��`��ZS��$�O@�$�OL�4���|�f�9).���*���p�*ަX�
�j�Q/�y"m�^�R�O\l��M�Ŷim�̚B:QyTY��
N 5�1e�|��f>Ob�d�27�x��'{�pʓ�r��Sxx�@`ƾrV����E9%���̓�?i��?��?����OL�9&	H�-&]�U��f(,�S�T� ����M��B��/r�h��<��JN(+��IU�E7}�`�GV=)��'��6��ަ��?���lZ�<a�/�����e�!N���xND&Ѣ�!_8�$ލ�䓚���O����O���@�y2�EX�MM3H>��H����:wd���O����&%	����'y�S>�ka�ٱ1�=3��L��O'?�!V����4i)�6,�4�f��=xW���X�M�/C�^$ʳ"=lU`<ʡ-ѴN��ʓ�����O��H>���W��E ��\+q�,�[�͊��?����?���?�|J-O��mZl*Ip�@Q:o�u���֫kP c�Dy�b�R�� �$�E}Rnl���1��d|��ԇ3d�֡jV���MK�4	����ڴ�yb�'�R�0��?Y��Z�䛒�K'35����,A<���p
p�x�'��'�r�'���'��z��:1�'i��Rq����hQ޴U� 8����?������<a���yG�̲E@�B�>'tfa��%�9~D�6���i�L<�'�J�'tq���4�y".�n���h��^%��|��)�y�.^��i�I�<~�'��ߟ�	J����R�k�(�zQ��#{u�Iǟ�����8�',�6�J���O��䎽" �S�_��Z����5_i��"��u}�xӸ�mZ���(�E��/ϡ$XL��P�N'b�ܕ̓�?��Ł�`�J42�^�����R�waB����$1R�̖($V�z��O�^���D�OR�d�O���'ڧ�?���3(r��@(�A؎0�녶�?�b�i9x�X X�޴���y�(4y��p�aj�~ڒI��d ��y��o� n"�M;��5�M��'&bM��No���3yU<�#/�Vʴ<C$)�8K^8�W�|Y�P�	��,���L�������J@�Q���P+"h���pyRBiӒ����O��D�O:���$��n� I��VT�h�PhI��!�'��6�Ǧ=�J<�'���'12z\� ��G����I&��Y����bʘ���6:41��.�O�
L>�/O�=@aL�4E�VDD�ְBdV8���OJ�D�OB�D�O�<�Կi�F<���'"T�
��ȋB<a��*]=4��ۙ'1�6�&�I���$E���Y�4�?����5�����P #��i�2	ʍTU�T�ܴ���$N6m��'��O�>�،#@�I�g��;v�=�!�
� �H��ԟ��I���Iڟ�	M��
\�����{P��$ڒE�t	����?���Ư6�a��M;M>�����4��&�a��@6���y�Z��(�4tW��Oe�A��i�ɵ�j�b_�*����"�^�(g�,#"`�\�Ily�O-"�'�b����qh�m�@�r<�#��CO��'�剂�M�2���?1��?�)���#&�A�k��K'N�fi~�ps��0�O��lZ��M;`�xʟ�hfhܭH� 81������e%O�j����3N��]|��|j7��O�u�K>��d 5\��D�����Y:����?��?	���?�|�+O��m���:P�.��4��k�4K��+�iycr�����O�l�k�0�:�G�8�d �5/�/$�|���4q囦��.�V3Ol�$U9M<~���'{q��{��u�@�+z�IwJ��.En-����O��d�O����O���|r$b�R��
�뀱iVT��tЁ_�V��9U���rS��y�S �<	�� S�����J{�27��Ǧ��K<�'����-$����4�yb�Hn�����܁T����2��y2��Jx���.)��'~�I�4�I�yva�׎��*�I���rK�M���d�Iޟ�'�7-X"�����O��D	)IL���m[*6|�y���-R]�⟴��O�m�>�M{r�x2�L�nO*�#Q%�e^$!�+�9��$J2Mˤ5 ѠBqlҒ��98��slD�D@�n�;�O9?[�!ʕ��. �0�$�O����OX��*�'�?A!O|*$0�0��R���?A�iV� h!V�`�ߴ���y�"��oLd=�gQ7�F8Q4���~2�'���*d��i�ҍp�6�V!�)�@ �}��K�;[�����
%g�P� '���'���'���'/�'ŘM!Ž1|l��Ǝ1�P�BY�� �4�L�	��?���j+��<]䚙`�f V��ф� O��'�7m�˦�SM<�'�J�'y��K1nԳS\P����y�I��O�B�L-j/O��"���?��4���<0G��/�@T�Ձ��1�����?����?��?ͧ��d��q�(��t���5ڽ�*�#cE�m�C�h��K�4�?yL>9�R�<޴m��%~��!�V�ۖ�D��ЁÏz&��t�i��6�w�H��t�h[@�O:���']���wS��9E�'L낌�@�
J�t�'���'"��'ER�'���:FB�1���d�F��$�3e��O����On�O��'��6��Oʓd�z=���P�n�����5\��xh�x��q�n�o�?��6��㦝��?y�K��@�so�E�>Pz�a����0�g�OԙYN>-O����On�D�OЬ;��ƿMt�6Қ!
"�� ��O�d�<E�i?��e�'o��'��S�(�y�t��c�����D_rd�p��I��M�#�i�,O���R	�?;�܉����f�YP�jȠ�d�*�-��2z˓���+�O�T�O>14�ֹ1^�����3�L���K֤�?���?����?�|j*On5nڶ2X�P���.
=�=D��٨�j�@^@y2Cp�|�d4�d`}2�a�̤� `Qc!2C��!b��{�l������4a:H�*�4�yb�'�,Tj��?usTZ����F�'b�a��U�41@���
t� �'<r�'2�'D��'��S�(z��q�5*��C��!����4)U�x`���?Y����<���yl�_�8GA�:;�8�W���7��A�I<�|Z��@.�M�'����@�/ >�y�A�m��2�'�P!��C؟4�֘|�U�0��쟸#���7,?t5��@V�X�x���@ퟸ��՟���Wy��l�,��2��O��$�O�42����B�CĀ[�F�0�.������զ��4�'����s��
R�Ju{v홮<m��1�'����*gl:m*�mXq��	�?-�t�'h�E�	;Aҥdm�0X%��H��:� ������ܟ`��J�OwaR�'6��Ԡ��l�	p��#;2�d�ʕJ���<	�i:�O�Nդkl��I�J&�p��e� vq�ݦ�ܴ@2��CB$��2O��D��d�x��B�БuUIs�č�(^�Zϟ���OV˓�?����?����?��l��0�mJ�)W��{ŋ�� ��/OĤmڧ	�U�I��<�	V�s��q�Hͮ3�|!�3%	10�P�S"��'��Mܦ�۴uH���T�O����C�5�1���M�����B�lEY�^%J��2,
���'�(u'��'�l=s�lH>�����O����'�"�'����^�8	�4/P����x�����'Z*lCf��w�!���}�����_}��z�F!lZ��M�Md�f��pF�IQn@S������۴�y2�'SJ��4���?���U�T��ߥ��T�&��a��E�;鲐��r���I؟���4��⟘�Zk�3R�Ҽ�'�� �E̚��?���?!�iHXڳ\� ݴ��s,D��
�O
�8��Y���L�|��'���O͂�J��iJ�I8Ubi# "�'E䌱�`,x
� ]�,��X{�I~y��'*�'�ҡ�SՎ��v���wS �£N	�?9r�'g��6�M�ӧΩ�?���?y/�6�h@�{��y6mvK�������*�O��n��M#E�xʟ� Ne:��˱)��]Ȳ� P��JV,T&8/��@U�� ���|Z���O�|�H>�k��3��w(Ld��#�,)�,���O���OL��<��i�fQ��9A����q��0cS�K���*��ɲ�Mˊ��>a�iQ�t��b�8`��-!�*F�+�"���n�Pm��3h�El�D~�"`��1��+��%k�0�1$�Ҏ�t��,H+ ��Zy�'��'Y"�'��R>�{�'�&p��s��,
蒰���?�&�hyb�'��O}�b����F�@�E�dx@�0�Z���Qm�M��x����Ǉ@i��<O����2@F�8�]�2�ꈳP5O>-��ǋ�?�s�&���<����?!@���Z]Z N_%xb�:�Y��?a��?�������p���ޟ��Iğ����Q�|#���J7
"	�#�Q[�yu�I�Mc�i�BO�H���˼B�T���}B������8�4

�w5�Iӂ�C��u9B��ӟ�#Wc[Yx� K ͅ�k��a��F��L������ݟ�G��wk�����[-?�� Ӑ ��6G\�p�'�7�#G���O6io�F�ӼkS��#�������@M,dY4JF�<��i��7-�Ӧe:����-�'��8�R��?�x�m�VZ�֬� ��ԁc�U-T��'��I矜�	�����㟰�ɹ0ˮ1������љ��<&\���'�N6�ɇkG����O��0�9O��� �A+[Y�$��Á/DxՊ��Uk}�Na�\�n-���|j���R"��$/q�-����.d�X�a
wehP�����Y)����wO��O���H`�СEDQ�x� jUo7XlP���?����?1��|Z)O(pn��mj4���.N
�����P-���_2*��7�M���>!ƹiIB6m��5Z7�/L��K!0%�͑6Q�кi��D�O�92�fһ��a*�<9��ǿs����f�L�T���/8t���?����?���?y���O�F=�<$��TC?B?��3t�'!��'L6�^&X�h�j��F�|���fN�!0�1j5�9�b�K�2�O��oZ��M��d6eh�4�yb�'=��bȂ���Qs�j�7_-���2G�,�$H�I3��'����p��˟��	^c�c��8����m�)]4vd�Iܟ��'�7-\�'���O���|�4�����Er%e
�J�}0��WG~��>1��iu�6u�)"�)M/`���3�Ɛ2Nn^u�엩1�z��Ƃ�j9����ǟrԙ|�dX!q�h��N�9V>��ǭ��r�'3b�'����Q����4E*Z)�'+�&AD&�c�+�;n��al�"����y�?�[��*޴1��!YS �s�'��!Ό��is$6���&6�/?�#!\�	����DȊm�8*�\
&�,k����d�<i���?���?���?�.����Rf���-S�4��N��:�E��L��ş(�RG��y7�����x��S/Wh�ي� �*�Dj�Hu&���t:E�z���	c|���(z�F�s��E�&�.�;l� A�'�'�\`'�H�'���'��D1u/�*@��������I��'�B�'�_�:�4R��TZ��?)��q(�(��"b�H�"U�PwXi!���<i���MSВx�Ǹ_��t�CF6�ʅLT����^̓φ(|��f��������'	�qv*��`8:���A����OF�D�O���/ڧ�?����e<hi)��T�u�q8�ˁ�?�'�iMD���^�,��4���yJ��%5Z%z�� c #;�yRG|���n �M��E�M{�O��րE5������P�5��!>᪜ �o��G�|rU���	ȟP��ğ��I��L�QG����0#�ćIq�E��Cy� k�n���N�O�D�Oz���$���څ��L�z�t0 �� +�B��'F�7M¦�L<�|��	� d�=@�o�>��7kG/ T�G�����ެx�0��wKҒO��5�l��Q 2}*AX%l�-������?����?	��|.O�oZ�@,^)�I�Y��xH��/g�4�!7�Q(5�X牸�Mˍ"!�>��i��6m�O��"g�p�N��R.\qJ�胉�g66�>?i�#V&4#��)9�Ӗ�5@Z9 ���`�	Cx��N��y"�'���'���'���	�!�b�����?V�$L`q�t���O�$D˦��b�ryB��F�O��
Ѩ\�pn�Y ���0�`D��{��'T�6����Z��Dl^~MU;F_�Y��o�8�I!��mMt���������|�V��S៤��ʟ�0F��&ٰ�����1&z�	ş`�	Eyc|ӈ��I�O,�d�O�'%If-*���:K���%�-"�i�'f&�2���i��$��'bu��¤� ��q���O-FxJ}Vg.XW� 9�����4�.Q��vt�OD@�d"�n�~��O�o�r�KG��O��$�OR���O1�˓	���i��lt
�h��غy+\h��&�E� �fW�\cٴ��''\�Qg�vML`��KSL�!<���1�O/?w�6�֦��$�����'b� Bc.��?��1Z�d@5'�0��q@j�0|$��zQ�o���'���'?R�'�r�'��;]�p͚$�*��xц��-��t#ܴ�
�H���?������<9���yW�B�<���7�#QQ ���mu$6-M����H<�|2��Ҏ�M��'h�)���'9�J��ǥGP}��'�j�����ٟ$qt�|�]�X��˟	���.1�B�(���R��nٟ�������tyaӜ ��O�O���O��%�\�k�>��� I�@�*�P�h.�I������k�4&���� 6�2�ٵlԸ�p @3	[�����h�	���P�q��V�ӏ�⏌Ɵ��V(Y�q8T���� -�t�	"������	ҟl��ԟ�D���'혅�$�,~���)f%A(�%�OBxo�2)�Q�'�7m$�iޕcEۊ=<b�Y���96���ȧ������Y��4s�ʡq�4������ �'-��X7��\�>�C�M9xu��Q%C(��<��?���?)��?񥡚�	��uAkҽ�%� �P
��$�㦭���Dy��'�x�ӂ
^���)GN߹&.Ѕ*��W}bAm�t�o���Şv�
I��"��Ү9���J�9����+�_/0�Z*O^���_��?	 J!��<�,��ZH$fu�j �7���?)���?����?�'����=ۓ-ȟD��ˋK��Y��݊c`�Bob���4��'6,�5Û��hӪamZ�NF(�c�n?� ��qP
���m�Ϧ!�'ĝ `ɓ�?b@���w� ���.h���'�Y�w��eȟ'�r�'�b�'���'��fmX�g��9�xA��Y'q�8�I�.�O���O�n� ��͖'L$7�?�$�&����TKK�&	���3��j�%����4^x��Ox���E�iM�ɭ;;1�'HғE��%���,~�)�	ъz�"�B��Ky��'���'7b�ȫy���c��*s�B	�͌D�'Y�	8�M�4�<�?���?�.���C���'�8$��́�}�X�[đ��[�OؼoZ��M�%�xʟ���nE�51��(͇��@g@ϬJ��l���3U�R��|z�%�Of-CK>a�lΖS6\����z$�0���?����?����?�|
/Oz�o�33I�13�+FP#VN�S�rs��sy��xӘ�`#�O5l�-ot����œ�1�l�+��@����޴3s��AJ>4�F������S50����{y�Q�ɀ�r�j���yA�,Ұ�y�\�\�I៌����`�	���OZ���CnB�|�3^��U��͂�5��pM�I�|�IW�s������cvl��o��I�A� �l��:věրm�x$�b>�i�C���Γ~���#�?v�>�	 ��`�ϓZ:*�#���OI>	.O��O �PA�֔�v�h�!E3.&���tL�O��$�O���<Qֶi}؄ј'\��'J&I��A�q5P�#g�В����r}�w�*lZ��}�D��7mK;z�Q���(P \�'�`��l�qr@���dNܟ4���'��NO�i��#�
r�`�'�B�'�B�'��>��?���Qq�ͳ�nZ�:�(�	�M��G�b~2�oӖ��ݨr�и�'���&�AW�&��牳�M�V�i�6-�>9��6�%?���@.$Lr��A`� �6��$R�!����-
PL>�.O���O ���O@�d�O����	b ��%�̲8���2��<	�i�,u��'A��'���y�IN�[9��R�f�wy��+�dl��di���|�
�'�b>�z�	X`et4 �]�D �aD�F\����/?�"R<=������䓿�D�� R*�H悆Bj��Д�[R�t��O���O��4��˓V�v���y�EC�r��yђK�;'�b��n�8�y@x�z���O��lZ��M���i�v`�ͷY�� �/N�^�ꍺ"'�9�v���w�J1P������h�I�0 �\���8%��)�&3O����Od���O����O��dI�ZV�9�<��A���.UfDE���#:ҥ�K�Of���O�mZ��tA�'R&6�-�D!%o�a���$.�NxZb钄@��&���4z���O��◺i����O���&[:0�a�	�&E��l��
'~ ��+��d�V�O���?!���?��8<�,��(ɟNN�Q,�$Qs���?�`:L0B�,�
w�(�,O�����瓰j�2A[�CP
�b�T�S$*Y~�t�I��MB�i�RO����@��.�<2YP���Rd9p�kge&�@9�d5Y��˓��դ�Onq�L>!S`�C���B+�#[?��x���S<���i����@ο:��u�vF�%	���+�$����&�Mˍ�F�>i �i�^А	�>?k
�ض��	e�0��eӒ�l�.�x�n��<I��O:���c��D�x)ODi��M������T!ztv5ʠ>O\ʓ��=�,���$�k#LK14:ZI9��K�$���ɀ�qo��ʟ������y�⌓jt�H��*gV�9���ZL�6�ѦM�N<�'�b��E�d��4�yb�Y�8��$rVLR����kRFǸ�y�/�g�"y�	�&.�'���Ky�̌q�,D`ê�#� 4WǕ5�0<���i,l�� [��	�a�:���d�(+b��&��?QFQ����4yQ�fl(�$_�NV�EIu��4^����	;m�$�O�)��e�'D�.���d�<���9��D��?�a@R�6�f=4�\^��d:��Wg�<)� �1)�>ɪ� P\�n�{�-���?1ÿi���b�[��{ش���y���{0��P`O�%P��y�D��yR"c���m��M�4�[�P#;OJ�Ċ6~�^����7���8�%��s/aK5���*�|��!�D�<I����*�,�:�*��(I )6%��	=�M[)G���D�O��?)k!�:���+���'�N�#������O�6m�I�韴����x"� z�%@۰d�@5I$��y8���c�<!�d��6q����䓵��>�H�92�z�AB��a|r�w� �H���O(u�� �Q�`}�Gl�0Zk����;O�IlZm����4�MCտi�>6� B���h2̊b�Xa����
N� ��7�k���		X�Z�"��O�2L�' �t�wrl:��l���cgɏ�&��(�'A�2��/�-+01t*P��Vɇ@�����x�ش2�^ �O�6m#�d� �]�S�*i�Mi.��Ro¹'�Hm���M���q&l��4�y�'��m����"m�����%J�gH �b��:p�5�I/�'v�IE�.�1��NW�]�$S7*C�$}Exr�rӸ�X׬�<1�����T ��M �HY�"��!X"
��ra�������O 6M\D����i�<�V��%�
A<q@�)�6Jx�c5��	7�Q��<���o$���D���U�N����ܸ~�DdsA�r�x���M�˱�p�3�L�g/��Zp:
�C Q�L��4��'#����Vl�/~H��(?v2��J0�:�6M	���
5N���5�'N���I��?�J�Q����F-�~ݐ��Z��srk�̖'=�{��_��ѥ�O��'Ţy��7�G;�p��?���$Be��>@Tc7n�.*DD�b$^	V�@�m(�MK��x���f֑ �6;O�ܒ��K,[��@0��h�4O���K��?)Ӡ7��<����?aB�A�}�z�{�.G-O���C���?����?�����礪���ty��'�(њ��

���� �Q�p����f�Mw}�/j�fo��ē6?Ԍ)_��pq��N�����;?���M�1Dl�(B�X&��"A�mZ�Ll���H�D��7BM�)��DZ,SJ���'0��'���S�$��֕��@	C!^v���П���4<p`�'��6�,�i�)�����RxBu�}�����l�Hj�4/��v�d���a'}�t� 'R���|ם ?M��3�@�5L�����&]j C|�R���͟���Ο��I֟r�ɄS�ܔ��E�u9Ī�hyBai��]��8OJ�D�ON�����Cԍa@�Z.]�����
M9Aθ�'�v7MP���!O<�|*�,;�r�"�Y�"gVA�&y6`���i~B�L�n��IRB�'��	�*�� ����x" ���ϟ#�`t�I���I��\�i>y�'��6m�~1󄌌&�2�B�l
��`8� 'W�H=��U�?�`[�4��尿��4ev"Ń��G4i��2���<�U���M��OxR��ܝ������wt�x�$Nٔo'zd�#�3��1��'�B�'�']�'�(�Lڄb
Ak���m/|�y�1O����OTm���>�:қV�|2d�a�@�ځe�Z6"�� BI�Ht�O$�$i�󩎪7|7>?!��0:c��{�� ,3`$Bk_>d�l��"��O�	�J>�*O���O����O����\h�� ��L�;7��x�n�O��D�<ц�i0@�'W2�'��S�?�RoB!u�:=����$
l�:�����M׷iȄO�SG�h���1�H����1r�Y`0!�j߮�<?�'xԮ�����J�0J@���NF�:"�G"����?����?��S�'��ݦ��$�~�t!�D������Ǐ)fc��A�&�D�A}b�y�Dp�wbFj��)��I*e�ftʢGT�� �4��2�4���@��i�����SԐ�f�9,x���c�6��Yy��'��'A��'
�P>�Cc�CǮL���Z"��ܘ�@�1�M��&��?����?�O~���c��w��:'��/}ء V�T�v�����z�D�nZ���Ş.o���ڴ�y��ƴN�pAH�+U�R���6B���y�	T�Z���mb�'���؟��	�rUĜR���"-�V���}\v�����,��럐�'�(6m¶^�Z�$�O���R>M؜���(T|~��P�ԥ�:�X��OܼmZ��M�A�x"�="d#j��i��d �hU?����:u�P�d��*rΤ��h	���~�&�-5����R"&5"F�J"*"���O��$�O��D3ڧ�?qc�>-`H|z�o	�[���;0m�
�?	�i7 4�A[�x�ܴ���y�n	4}�Ҽ#�+��X�\2�d@��yҥm�xtl�M�����M��O� yt�ʁ�J��֣0c��X��B�tX|�� :n��O\ʓ�?q��?a��?��I4i!3,E�^R���C��[@�-O�lڦh4&x�	�	n�s��s��>3֐j���?j6��v	����X���47Љ��OCF�"g�8,���;e��!g�DPs N�w�&���_����`:12�Co�IFybh�ZA\�ۥ	D=%p*h������'�B�''�O�I��M{�<�A`Ժʌ�Z�N�C�82�i��<a��iI�Ox(�'��6͈��(�4-���81M �	�%��ܤm�DZ�, �M��Ol����/�j����w�-���3��C+���a��<	��?Y���?i��?���� T	\:b�M�KW�	��X��y��'�"Fz�Bl�!�����4��1HZ4�$&3\3��s�#_�� I��x� g�<�oz>%���զ��'e��a���'�l�,� df�%���eRX�	�`��'T�)�s�H��J�(�xq򰢁2?���� �!�j%�&�X+W�񟀗OP�������T�br Y o����L}Kx� po���S���^�"$2`H �[��d
DgS�&=�=8am߄i���[��3|�b^|�䈸�������P��8B�ɕ�M��f��3� �*Cj�|�0Y���U7_�f)+O`o�v�z���'�M� ����	F���]�pb��U�Ϧu�ݴu����4��$�DF(�+�'rbDʓOb�0�I�0�0T�v,ڑ�z�Γ���OV���O���O���|�Q�=f�^h�ɍ����7�B�:��D�O���&�9O>�nz��3��?B��RqטrH4������?	�4�yb^����PXŁ���	�_y6ċ�k��^4p}����d���I�hq����'1*,$�������'Q�ES�%�`�R��$�:60����'L�'U�V��9�4������?)��8�Q�G�>&�P��1Hi=�%/�I����O`7�s�8�'�����k���r@G�*�q�O�ӵ��3��TТ�Ɏ2�?���On8����|���E%�M��� �O����O����Oޢ}��j��I��f��T	f�M�z~l���GP�6E *��		�MK��w)�ht,����8R
������'�J6��Ԧ����t� hoZr~�
�� ��ӃF��1 ��3{����8z��+��|T���P�I՟P�	����g.	�EID��7����U��ny�{� �'�Ot��O�����F
h���"G�E� ��ȉ�<Ҏ��'�7���!��H����P�?��U�5�6���Ǉ�%u��仢��
ǣ�-v��-d@ԣ�N����[�GQ"t×(څO|A+�V-趥�����[�"�$Q�a!�Ӆ`Gr�Y�JۥCG*!�Q/>���5���C�l�4%�9(�r-�2��h�cj���T�T&f�B�ѓ+K 2�.��m��I�@qRf/8��0P��h�Ը;$� k�z���Iң֢��e��Ԑ[�U�|�m*!��7$AnA� �c<��jtL߹,�r��Qc��'h$p���X�H�ܑ1F̔�2&΁�ƈ�,�R���`u�d9�#c�c�@�ҡ��/^��D�خD赎�6"����q�6�G�\"E�(v����5��^}��'v�|��'w�J^�$��!Q�Z1��S�h@L��%ài�6M�O��d�O6��O��`kC�O�������c� ./�̩�3� �0L5�'	k����>�d�O��H�RV���x ��]�Ȼɉ����%��MK���?9���?y��	$�?���?�����ͷDrr�!vl�#0�R疭6�'G��'���8f����������c��)G��8W��Сp�Z�X��f�'�c��:*��'��I�?������0��y����eR��4�67��O��D�[i���f��I͖+8@�f�<|�����8z����N�cr�'�	�?���џh�'p�Y�b6�u����e�,Tk�{�ˆ�B�n��y����O�=��T	�Ԙ���A�r2��J!�˦e��[y�_�)���Zy��'��D�U����SHD�}:�5ae�ͼb�*��<y��?��'�?���?QE,�Oꂝ���@+�ԋ�2;���'?$a�R��q����'�ē�?�I��+k�@�f-E:t1�'��.�^�H�O����O2��<ɦ"�\�H��B��FpR�*c��$ ؉�cX� �'�2�|B�'���ݪ,Y@ Vh��֠0ǁ�&�|��':��'��	~���K�O .U·�4jT��Hrb��b�x��4���O��O����Oz�9#����p��+$U4�ЄR�2�j�B�>)���?����^J]�O$�	�-BY1`K�>���� c�ws�6��O�O����O���>�I�@��ȡ՟$�
1-�@� 7��Oz�d�<)��ZT�����H�I�?��v�l���J�/�ưH׋߱�ē�?i���N���Bܟ�8�G��0���U� �2��i���
t
�L�޴�?���?��m��i���w�C(Ɉ�+G2h���J�z�,�D�ORd�,5�	nܧ X�@�$�9#`�hƠC0Tۮ oZfd\Zٴ�?���?���/(�	Gy6GJZ`��?VQtu�Ҧ+�T7M�e��$>�$)���h���e��lTB£cR8A��ʝ�M����?q�<��]��[�h�'���O�R�ς�m$��qC��saf�`��i��'K(b@L/���O����OV���Rg���b��B76�4u�$�TצE�ɸ�|q�OF��?�O>��+�R�cm(=���l�&Z���':`����'��IƟ0�	� �'�H���9 ����0��,x��Jq�ī�x�����Ob�O����O�p)UFͮR^e[F�"C�%��΃=_ВO��d�O��$�<�'�N�I�bڭ`�(ÖYtA�E�x��\���Ig�Iӟ��I1����4LX{����� �C���r��O����O0��<Aɏv��\{sdX�m��ܸ��Ǣ8m�Y��-ǂ�MC����?I�}A�Xq�{r [��"|�ũ����"�� �M���?y+O��R���K����s���M�xjq��a޲E��qÊ=��<���L��?1I~z�O�z��bE��*��D�p�L��޴���6;*�oڐ��i�O��x~��5��}pS��.%�v�����M�)O��`Ť�Oܠ&>�&?7�[1. ��8Ō�%y@�x[i�<nZ76zx޴�?q���?���v̉���@�}\� A!OZM��q)G�t 7�ҷd`��$�O,˓���<	��$S�1H���N��J$ȒD@2����i`��'���q�PO�	�O~�ɕ���Di���H��։cF���4�?I*O��p�J�}��'5�'!`�����#ϩX��x��^�v��7��OJ\P�L\�i>��IY�i݉ rG�h�r���Eʎ5���9�#�>3@��?M>i���$�O�i����2�i�e5�t�dj�-1�ʓ�?����'^��'e:5��N6Hdx0���Y;V�i4�GHf�x�y��'H�IʟLHƃ�X� �8�&Υ*5������hйi=r�'�O����O���CF�;ϛ�
�5	�N���������?.O.�D�^�r�'�?	X�ډjɂ$�����)R���nk��?i�d�:T���q�I�w��ժW�	�Vy�h��ұ��6�O*��?�E���i�OZ�D��klC�=K&8�%��wcN��aJ:7�'�R[���.6�Ӻ3'`�p1���� wx)�L}��'�I���'��'���O��i��Aw/���uy�7�0d~���D�<� Jz���'L ��a�Yj�|� c�	HL$�mڹ���	�	�<�S}yʟ��iqD[ 0�Ƭ�CΗ�H����\}J��O1�h�dP (�:	zr��=�T��b	��l�꟔��ӟLQ�dٛ���|���~�F��2��A�`M�>=�6�j���.�M[����$�S6(���y��'Y��'�ʄ��+0 IX#/�:+�4pf�vӰ���?j4h$��ڟd$��݈Z`|��	�x�lq��F�x�F����$�O����O��e�()wJ�X��	�O��&� �ےk����'L��'�'M�	)*��5s�@�	b-��P�B�XJ��d�Z��0�'"�'��P�0�������d�ƕCa.�#��,;� ���
�byr�'���|b_��2����9�%���lyF	<7ص*T�����$�OV�d�O>ʓ�,�Ж�A�5�Ι�$H�Ex���P�L�u�$6m�O�O ˓RV�в���(h�d*P���#@n��sǉ`$6��O��$�<���L@I�Ou"��5F-����0{g�۹d�&�QHR����O�˓}`��B����'���욿g���mݕ/:b�AGU�����O��HC�O.���O���⟶�Ӻ3u$�Y��&�=J�P\�)G���'Y��-u��y��Gӊ	�u�4�W?v^��;PL��Mg[!�?���?����
/O���	O�D�"�%bk�E(p�S3ga,|�ݴZyܝA���N�S�OW_��xJ���$uԅ��I�:|T7��Ob���O�����<�O��p�&!B4��+܈����f#(`���Hg'֝&>�	؟���$DLڸ�ЍC�N���#�#:���ܴ�?y���	dщ����'��QZA�O i����p�0Y��$�eL�j}b�]#QRT�������	Qyb��!z2$PE�V��B�ÀS�nY"I#�$�O��$2��<���9� 03�FΗHF`��B]�B��?Y)O����O�D�<i��+��	A�AF��C�H0 ��@�J֩*��I� ��J�	by"�hy��H`�Z�I#���)�����N8듅?����?q(O�ѹ#e��d�'�Z( �Ŗ�g�"�����cV�hV�e�p�Ĺ<���?���~�d\ϓ�?1�'���c�l��Lg�*:�XU�ߴ�?����֔i�^U�OZ��'�t�R�a� ��I4���Ef�����?y���yҊ�m��^��'"N�T�C��q�ܸ4
Ncu��l�_y��3Q�d6��O����O���DL}Zw�[!�� ���H�&(i�ش�?i�dK~H͓�?.OB�>ʂ���)����HB�M�Ԩ` a��08$e��������I�?�ʯO|�P�^���GĎ\�|0d �B�y9P�i�
�a�'��'��z����dQ���S�Ūbi���֊#���o����I�ԫ6D�����<����~BL�~<`����T:n���g_1�M���?���x�~5�S��'�r�'}�E�3�?�>��!�� �H��j��dS70���'����$�'�Zc�,1�O	�_�2]�b�[PK<t��O�`�e;O����O����OH�$�<��·RY2���g�,B�a�o�IF�x�U�D�'��T�@�I�����-4Ad8H�b��t�9�<�I�4�Iܟ��'|J��u�x>qh@a#p)�NT.���.v�8ʓ�?�)O:��O���U���
jx���(͘}�r����;rՔ��'���'f�\�PX&J^���i�Oz��6�H�p�<4#�Dj;����䦑�ICy"�'1R�'�^���'��7��4��N֏N�t}����F9D�m؟t��ny2D�D���?y���2�H,%�޴u'�-XUNGJ�"lu��������8§�q����ly�ݟ8!"�
�9���#��� q��2��i��	F�y�۴�?q��?!�'3q�i��#k߬� @掍	���ȓg�b���O���t3O��d�<9��$�W"���#�ɑ7�L	��k�MCCj5���'���'�����>.Ob1x��/
HUaQ���h�������R)h����џ,��B�'�?B� �Fn�֮X�i�&a���}I���'�"�'y��(5@�>�.O0����[E�Y3C�e ��
4��]�!�fӘ�D�OL�D��OM�?���ΟT�I1g�&��#�*��ϒ0P2��ش�?��.�A��Ly��'���̟�(3G(�a�ǚ����@�]�uD�`cb���?1��?I��?	*O>�b�OѵBע�bkROx�PrX��!��>�,OB�$�<���?����|Xg��%��`Ȱ �P�a�# V�<i*O0��O����<�C!ZL�i�| 섹��W�f���wJ�W�_����|y�'v��';��!�O���V%BXTE _�(�b����M���?��?�*O�����\����5��
�H`,����/�ހ�sBO��M����$�O���Of����?�q`d��j�w���`!]z�m�ş���Ay��Z8�4�'�?A���� ��k�(�-����4��28^8V�h�	䟐�	[��T���'���
�G�-KSe�&	�,܀w$Ρ`���X� �#�F�M����?A��JvT��ݪn�B�# '�}�\)�AH�d7��O���M�\��,�$7�Ӑ[t���d�*��DlF�7T7����.�nП0�	ğ��ӛ����<a��>C�� Y�%�4����h�t@�6$0�y��'@�Ia���?ae˄N�>�"�H�C��������P5�&�'Lb�'m�y1�Ŧ>!*O�D����GL�+=��Y�D
�n� �Bp�>�/O&�2����ݟ��	���]20�e1�N�#��L� l��MC��p�l�YUT���'��[���i�u��AU�RPBa����#k&�x�&�>���M�<q���?���?Y����d� zS"�q(�<U��Uȓ�ԫ>��dj%%�[}B^����^yR�'�"�'�q�� uZ0�X�gA�b7|]�E���y"U���	��TybĂ�Y��,P��5��(G��Έ�l� CE7M�<!���d�O���O<�(�:OL����:�����R�
1���Uܦ��Iܟ�������'���Q�G�~2��C�*�/XtUUC�'oI\ɱ�զ��Ijy��'���'Q�:�'�s�#��R|�T��)��O�&�i�B�'��M�α鮟6���O6���70��a�
eq�lҁ�Y,j̕�'Z��'�B�� ���<)�OҠ��� �i�m�3��&{
�*ش���BK���o������O|���}~`M�~˘�9se��4sJ�S���/�Mc���?�����<�M>َ��ۿQ��!���,7e�!� -��M����.��6�'���'��T�>�ɾQ�4�#@%�ts2���HRC��ٴ��͓����O�⌀�_k��wA�i�'�?L�l6��O,��O�R��BM��?1�'���$�)fB��LӄD�F�Aٴ��M��M�S���'���'�>!R��EN��店$:PI�ԙ��d�����<v�b)�>a�������7X�����>'��i9b�C}2͇�A�_��I���y¨��
��U�S��\p���Z��EQ�0�D�O���*�d�O���Q�/�ҁ:�EO
)��@�B�M�WpSU�O�ʓ�?����?�+OH�����|:OP!�&r�"��	� ����l�	��$�H�I���y��f�*cŚ���9�%�� ��b#b���$�O<���O�ʓ[�l x&�������y��E��~H�%,�
)��7��O��O>���O�uJ�c�O��'v$�$�5=v�1Q�&E��=�4�?9����$��4&>q�I�?��MܵZ ��(]tڸ������?!��&Ix�����䓂����
9N�X�E�G-s(�`��!ǻ�MS)O��	���Ŧ9���.�d���Q�'�� W GhBGÑ�1�}�ڴ�?��*h�����OH��"� Q�/���
�?)����42n�$��i�r�'0B�O�b��"��I%L�<4��G�&�EQa�-�M�%��?�L>����'�0�R���
u� ��h� Q<V�r�Is�����O��S�}/�d&� �I�����]՜�Q!�>tv�Ab��2aB&@ns�	;/����sy��'���5�Ԉs)3�Ё/*�l+�ğ��M;�r/�Ǖx"�'��|Zc,����.t^�1ՠ�7R�h=�O�E�3��O���?���?�.OR��ǂIx� ��H�$�`����6Z-H��>)���䓘?!�� �ڨ��d��S3�-b¢�eҵ�.�<-O|��OP�$�<��L$��3,��J��/'ԍ�uF��r1�	��xD{��'��@{�''X�"d@�W� ×�O��1�cӆ���O���O`ʓ5�6勵��d�)J��0 �ص�<$���1M�6M7ړ�?᧡L��?Q���~ªJ(vH1���(<��lʠ�M����?	+OLh�G%IB�ß��s���# 1N�
#���$�1׌=�I��l���Rǟd��ly��np�u�2<&X�S�L(�|pz��i���'����'��'z��O2��5&I߇[�Υ�@(�:d��H[��
��M���?A&�F�Ԏ��<�~Rg"O�8����Q��UD:���W�����X��M���?����J@�x�OG2096GJ�t�b�{�c�v�Dx�t&x�Jh��	>�	�?c����)�J����� '�Y#�ʰ8%z��ݴ�?	���?Y�#�?!����I�O��ɦJ��`�fʆp���G��*?ԐQ�yB'<;�*�`��O��D�`t�IA���RAP�ǅ�La�en��T�V���'t2�|Zc
��K�'�f\�Q�G�g,.�A�O.l���d�O����O"�S`�q�!M	y��m@�JTVn�� ��ē�?����?�dpaKe8_�,D�D���>�`��q��?q��?���?�o����œ �p�pg�*'ZL$�L��M[*O��d(�$�O���	U,��i����W�ˊ�����+�$�8�ЯO(���O���<�2��4�Op��E�5JH�1�@�����c!�}�H�d�O⟘�g�2�ӄ�liH���A�JT�F��(>	�7��O����O*���/˧���&��#��!0�0�BwNKZ�bQ��U��柰��t����i �~BAD�k3P�A��:����@Ц�'`*DZ�i�꧔?��i<���#ў ���ą���n�:7�O\�Ĕ�"9� �}bq��"��]	"d9'�R�Z�����c�զ)�	ʟ�	�?�J<1��r�� >���c[-0)C0 + �A��iv����ğL��D�='��r�}@�p�F���M����?q�~�,S����Or�	(O��gi�n	�!���H�b��5�9�Iҟl���d#���UzL$`��0jת8{��7�M���B�Q�q�x��'H��|Zc�z��q� ���Cq��>�A��O
����O2���OJʓ<�Љ��d��4MfͲC�įNc�`$�FN��_y��'���ߟp�	��;�I��� )��焗 -�QPEBo�@���|�I��	���'�hU�P�{>)Q�3t0�e� H&�t��+z��˓�?�)O��D�O|�DH@���I)K45y��A#��[f/U{}r�'�2�'��I?@lfȪ�F�K�%ij���Y�w|�ٳi�	^٨�m��l�'�R�'��K��yr�>y���80�vi+rj�y���T��ܦ������'�7�x��'L��Of��Sp(	�Nࠤ?e�:,����>1���?A��`��	̓�?I*O6�/���i�䍪sF�1��ÖaѾ7;<���%�V�'���'�4�>�;-�ʼ�e�ȁIӾY�#�V>Zt�1oٟ��,/�#<��d���}��Ayr*�7fJ*��U.�M�5�]�RL�V�'���'���>1,O��K�G%��uQ��A�>Y
o����St�4�'3��)�OLP2!�Z�� ��i���[ڦq���X��0���P�O˓�?��'e��Z��A��Mq!A�!?@<�2ڴ�?�*O<p�4O�ǟ,�	y���$�>�����1N��s�R�e�ɻoKPq�'�"�'�?yH>���I?H��nA(w��+3����I�fUbc�h�����	ٟ���9Q&���#
~�V` @���A�Ly2�'S��'#�'R��'G6p���w�ҼBBC�/"`�P!gJ�N�\��O<���O����<c��
MP���6 Yĭ��-�:ot|�!��&L=�f�'���'��D].<��ɭ,c�
�a�'���@�Q���?y��?���?�fFH��?a���?�
0�8� �02���i���C���'�'�P�lr"A1�$W.#�Xȣ����$ш��!��k��~"�ֽ)����%�4
�ƫ�y2�%@\&��m�{���! �X5tp�M2�e��M���w�KQV�G�#MG�{�l�j��Q�R?`X��r���DMle�k׭wdD�{�(�LvB|��CY9D̞���Q�z�i$�� p%���mܻ[<��t- �X^ܠF�[�5x�%��W�`7@�s~�`�aA#>�ʑC��Cư,�aӪ]6�$�OJ��Ov��;;6�0�؛67 �1S�̘	�Ę��fW�10R @�
�\������Oe�'Ő�ҶL�x76�+2�I;��Ҧ�U I��\ɔ�:`֠S�]�I�x=��+�|�E�%K���݉W���2⦋�W���G/!�U�Ie~b�^>�?�'�hOYPv��:)���s�㗶U��p�"Ob��V?M�(I+�!����|�����i���?�'�\5'��xה�W�C/-؜�f$��S�
��w�'�r�'Vr'p�Y�	㟜ͧi����N�~�#���~����`D���\8�V�R����ϓ&�l����ڇ'�`٪��$utt�# m���I��4
B��;
ϓn��(�����8���?�(țt(������o�'��Ol髧K� n�6YYg�
^QQ@"Oq�����Ii& Q�1˂��M}BY���������O��cegK�?D�fN�l	�7��O��D !��D�O��S֬Sb�|K�j��5�
T�OgF�8&'N�����b,6O�!���(V��u,�*l#����#>.i��C߳.��i7��>�p<���Ɵ�Ity�Yr�j�!��*�4ੵ*B#Ϙ'��{���O� �	mj�\9j	�xb	r��Px�Bǻl���嬂��xtC$8OD�B>��ڴ�?y����݌?�����gW���V��L�+�)��P&��Or��P/B�l�v@�7�~�[>��OG�l*׋^�+�:���;2�O�P����S[����L�~ŞU��ڼS�ҹa��?�ɱ'�.(�tj�퐈aN�A	(}��ۡ�?y��i�\6��O(�?90%�
&}Yd,a�T82h���p�H�'B�^��g�S���Th�OvP�鐄Z�;""��<Ɉy2�iv�6M�OV�lZ�4R��@ ѩ��ª3yD1AaT��M����?���cF6�FC��?����?���ҿ!�B!]L����V�x����N
'Dh ۶縟��׍� v�$?c�Z'׆z4����K@/�y�GչD�m�T\�s���s�̒Q[��>5 a�<ɖ��x��#ՌX�_dT��$�^��?��i�r��*���,O����5V�\iBA$	8W��i�.Z�����>y@�D9��ɒ5G\m`��c��B��q�X�m�]��h�DP� ȲB�0G��G�� )���� D��Ћ��u����f(�ZMD�>D��2tdѦd/�=k���%8V�"�7D�,�v�A1��t
&��2M|���:D�(q� K	i(���JJE�AKk9D��;EJ��N�$ܩ&����Y�c�6D�� $�WB����#��<�D���"O�i�M�
�!�`ԌE�~��"O$˃��L�ddO�mrx$"O��.CҶ��Ʈ* �����"O�1s  �&����N˨<˄��E"O�XQЌ�^)ld��k
;Pj2-;1"O䍨C��BI9��U�-N�T�D"O& "��_�9r�"�'"I�}*�"O��щϺCd
1��=v+�ѡ�"O �J�m�#Z�|���	]�vA��"O$��H�<P�P���nH>�X��"O�J���T�f�
Q�e����"OH�!b��kj�lZ�
���@r"O�-�q`�3�L�
��a�h�i�"O����]c�>�; �T�X~z%+�"O
I�G@���@��@�s�%��"OF]�0��=�(���A�"`[d1�"O�Z�GL�?�(��`�:n^2P�"OP�p�̓.hNt)���
��ґ�"O�ْ�5�u�MP���"�"O<(J&)�6N��Y�V��yS�"O|m(�"�'o�*�Ɔ���"O|EC���+�f5�Re&k�}CA"O<�i�>/Vt!�qi҈N�^�y"OR�Qd.��Hb��kt�<�dղ�"O.C�I�\���:���,�<9kS"O�4Y!G�.y%�Ī���-sBdؤ"O\�p�ۂ/�Q@�n�3Wp|�A"O�)��#r��! �ѫ"�f4� "O�=�R"�w����KƝl�\��"OP��Nٛdv`��Ȣ��#�"O��7��פ���F&$�J(kA"O�����#&��A�"�����c"O�A@��r��B���̌�R�"O�Y�%�5R2��넏C�<��"O�0a�_9G����G�#|<��\��s�j2�S�OU��+���H0̴��Ȑ�zR,���'�D ���F�/:�W*(-]>�I>Q�**�0=�գ%���kC�V8;�A�!��M����U��Un���ŉ�
TȽ�����n8��&u�u���Ca� ��v���u�ER��i>s�'�>׶<�p���y�6��� 9D���v�C�g���O�A�>!����<�Go>���(�xIT(�<W�
Y�R���y�$"O j�jӷ?B�R��E)r�n��2�|B�D+v�az���/W4j�S'�V�lh7�{����9�n�bc*�0���\�j�L�A�<Q�"5X���#��.Q�	Y7���'�pub6�S,u$.=���޴%�hI�N3�C�ɱ��@*�Fɠ"4<	�A̘
v<�!�����i=Q�p��F�K�%n�0�7f��x�!���pf�Q+I�,�f ��PXq�'�v � �'S�Y��(�x��&į�~I��'[�0����`y��,�.i�b@�ˎ�y2�"L�ű�l�rvl\�F�G�y����2^������,� f ��y�,[�x��q䝰ZL������y��t�~����C!? �A@Ȓ�y�H�(�B�k���\r�g�H��y�e�$N��	4��� ��H���y"Y�D�y�%Q
hݢ��Ѕ[!�y�+E�<l*=c�e|��A��R�y&/wU�t�AÝV}��'�R!��'�txjL<��T0�.�fY�W�O+.7��{WJ 	����S"O� ��qG�*$:E��i��\�tԁ1@���!�0���(���)^�6�yr�Z H�����h�DB䉱T�<,��F2V�0�O�}85�'d�'+����!���R7C�&X��Ub�4=<��C�;|Ofh�C�>եJ��M����UZ| u-PU�$�1��a}R�J'<'b!��i��\�j$a#���')|��L<e&������� �|ՠ)�J(Y	`"O�̱����u^|��.��R��Eo���' ��P3��H���]5��u@ӂ��c���hQ-\�"��C�I]6�iE�<F;��h���$�打R<������6ZX����Z�'񾠻冈�i}!�$O#R)� �@�7��-B��$~X!��[=��t;�V�yL�(�A*�!�$�(K}:="�%N@f	�e�N[�!��$s\�}������|℅�/�!�$ܽP�\s�JE��U����T�!�D���t�6��%�s���X�!򄊫U� ��V��c0J!�D -i�to��V��a�O�<<!�dO�e�5k�i��,��l'��6!�ϗD�:ibpE.2�<5!�e�72#!�P�;�`���20�B1�J����y��P 1O�a����RJF;E��)��"O ����k�x`�IO���z��>� ���X��x��$��y����ӳDLd����yr���qB��Q#��G�NP���0gxQY�<�r�����'?� c�Ο#�Z "��|�J]Q�� �O�!`���Z��A�Մ;�l�%"�:��3̓- �Lڵ�'и"A�=�aې�/9�"�{��� i�n�s�öd��bE��|:P�B�B����59�Փ��x�<�{/�Q+��7�����uyB�X&\��Q��3��B̮~���`��3"��(�.!W�&��UmN��!�D�k�3���(	���u�(K ���V#L<�n��~z^�Z�e;��ON�c�O֨)���1D�z�x�oז^D$�QOV�*�̇%-(�:�h��`rJ�e��V �Ԏ��J6�	 �D�y���8ŨO�)xH�7kIzQh��Pb1h�;��'�<XT�[�XE"�G��M���P�X<BH�'R�<�x�Sᗴ�?�E#�B��l�V_8�2KY�_a��b�o)?�Ei��twRɢ��ǢM
��F��}�f	Kq+-�d�J>i�dI �LG�HxZ`*H�y¤@(ּ̉���?��1Ҥ�̚z����g�Ӭ����7�-�N���4�iR���'<�!��,��X��T2[LD����u<� �[\p�A*�P+���`�X2	VRL��	ߎxd����W�K�$�d�i~(�����G�	����
`NI�S��X�ax�C�035 qCuF��n>���+��,��K��ِJ�yA�fޤt{��;u�/$�Ař?4RjdA�@J�����-4?Ʉ@��j��p �)B� �(9�NZ���O��9��b�m.���c 6e܄8�'Wf<�� m��prF�"G��(ui�YH��	��)Yb�P#req��'R��Xr�M�[8t�P��9��- M�'C��i�a*��~�d��r^:EI��s#L ��,�G^�J`�P�,ыz��zҮ��T�!tK�����΢���/9`2p8�{�.TѨ=(�ȭ�����ݶOR�tK���-�@�b⃏,�!�$�wo&�+�
u�jЩu��%��'�z����ERs�n��~҃O�_50�z���Qn9��p�4�F���5��I�~� ��3��,���ELi7��	���Z�A��J�/.���I�9~@"|
����?�Al�9n*�!�W&Q�7��C��Q�c1�4��"'NV�_�J�b�F��)ݸ1 �cG;"d��A��f���	:�ʐD{kH�>>A�w9����*�0=������A��Ò��m��[����R��cL�sì�<X_�����i��8��ɴ+/�M���R�2b Y�*\=8�O X�"Lx�M��jj��r�E9q����o��ih-�@m;�8y�  ��{�!�D��τkEx-�6���d��\Q�K߂Δ<+�x,�2���$�|K4?�OҮ�˙w���(��&F0��E��D��	�'���Tݒ(�@��&�ݤ8WTH�0�dB�k��x�D��h�E��Tm�'�T\�,]0F����a$9o�p��ۓ<��� �% �|��2� ��a�l�'u̦�bT _'<��!P)�;&IFxP�d�
��t�ī�{X���'�N�vr̈s%��'D�So/��)rT�ٗ�4z���3'ƅ�s�FO\��C��� Mc�eg�V�؇�`H<QSF�??�@�`$��-R�`1U��=u�����+��P�&�6UޓO駻y���.�Vز�oA�7�&��怽�y�o��
N��`��[�	Z��F[|&)%���NK6���L�*v���ɕ�5��d=��p�)n��D��F�|-���,�1 �cA#|IzY�4��+[D����Ȍy��3E����
��AO XH�͚HM_x��s��dY8���8�l���H8Y��#�'k#K��1�
��<���}�T\�/�,K�u��"@>g%F�a�'c�hǈ�jxB��`��c0�*1��6h��/�J�> ;kـR��)���E�#нp�8W�>�l�r1"O4=Jd��=�҅�wa�RuBUFÃt�&�KK�tj������i�4a��t�תX�L����ҏҧ-N�tf0�O�u� ܀NpZ�i]N��[��?<��{� M�t�@cˑE����	(\O��ʲ�J"Z��������1@�� L@d�T-X�L@Z.r��M<h|B�BF�#"��a #A��N]�ȓ4���b�J�W�����؜h|J���lF��{�b�!k��̋¯ľtv����94�-�"��$2햰#A�e��?�"��#8`�?mB��YP��2��0'������͔%^хE�
S)�q�9���'!#�O�� �
7�4�j����
�^��1�A���b��E��̬}��|��H�����0��	������9�x��X�0: )lOD
�KT�ì�w�T�J� �sp�'�TU���+�DD�1TT���[>Xe�D�9?T%��)+�Q�A)�Zg�;P�[1jU�@��I��5�.OD�8���h�P��խL�_UܽCcP�@��͎.�J��b�*V<;��'ҧs��#�H�	!�5�U���*4�?�pV�b�?�.%��0Z��X�4:y{"�ڟ	�~VG��,S:]
�<�U�ߤ��g�*�2x�d��:*���I^�d����+����'��>���#�7��H�ܮu�ޠ��C]u1�l�t���G��'�(7a{�*��}�19g�ؗW�쌳��D��y�i�w��#<!��O�/��Y�!�t�L�m�{���ST�
s�8�jSM�PټB�	�?���,��C64�:s�jM����׭<w��qf�S�|4L{�c]�b"��:��\T,C�	�i��@ ����6͘�bZ���6^f0��CFY�)��<c	]�Br�	�B�����U Y�<�v��-�!1r�L�<Szeʀ	]V�<I4�p��@�A�U3Ut�D��J�<!���  ���!Z.��|�T��A�<9�kA9g�J�s��(2@=ʣ��z�<)��?a�pX9 ��*U��!B[�<�v�A�<8��ZSG�.�ʘ����V�<�bE�#T�j���O�806L0���^R�<����`C�ţ�
�5�̠ä�B�<)�"��k�P�9�E��-�mpF@�<���X�N��� &ׄ�@(��Xb�<	�*&c���e&xP� �G�<� O[]+L�Bf V 8��3U��Z�<9���!������O��t�aZ~�<!�*�7h�4�g��dǲ��NA�<	Pi�j	LCe�YQ�%�H�@�<ArER�0t�ܡ�!@�.�m��z�<������nx�i�>�jTq��\t�<�R�2eC*�{�/�R=��X��n�<�'��WLy��=+
�1r "T��	BKɫe{�)���f�P{`�;D���F�fR��Ef9#��@�S�&D�����ۼ^��tqD��4V1A�2D��q�D]�Pyd˵$�+�B�:D�+D���!�@:��0��HT�0�H(D�P�c��P�N�*�Η�C��Qw�2D��J�#��rtQ�b�+OD�<a�:D�@2�D�C��#��G���B�,:D�@y#`��t>mh�gN�|���*ǎ9D�Ԩ6��!�4��JM���`�f9D�� �5�����QZ/݄DZ���"Opt�#�35��	w.ɔT-H r"O(�"$��	lL�$�[#H50$"O�	��W
7u@�3�kD�@�T"O2���"FS� ���@�dXQE"O !oU�D�'�Ⱦs��X* "OT�:Ff���ȉd����"O8T9@�� �ġa�"���"O����&��}���@�S�s�Z�s�"O1����.�q��E�F)J�"O&e��	�Z
�Q[£Ǐ?��1"Or����=$H�#����F�`%�t"OBeS��ӫ��8V�	�C�n�"O(Qh�1�~aS�+�$d�x���"Of	ɕ�̺h�dH��%f��"O�@ȁ����֨��CW+�L�"O�aG(T7n �K��àl��B "O��a -��8��q//r�V"O�l�c垞!zR�3�M�aՐ�"O�!� C��k�(�A�Q�&D�D"O��^ �j���^Yڰ�"O�!'B����Ȅ-S�K��A"O"�aaXU:���m��>��e"OD�bC��
���I��;_��"O�kg�
5&DP�I�8i�"O��J�f� "E:S������Y0"O��A�	�RW,�맩�1-�`�"O�`�FX2o�����gS�)��!�G"O�x�t�J1q��"��X�d���'��%��+�R�`QI���0�'x�"�ڥ4O�1,Ҿ>
ZE��'�.eZ�j&WnJ�9��/>�J���'yHl�#�L9b����Ŕ;<z��+�'�N��.VS�^��G�#9�V�I
�'�~���h7m��|q́�>�,�1�'��w�Qei�I���%1v����'-T���n;FKX<P�Z�R�Z�'# 10S(_*j�kWeW4NL���'.H�F�!h�pegn�?l`��'G
���I�m�F[Fl�*'��#�'Wb�%�߇S�T�dH
�i�"E:	�'kZ@rw�%��@D�C�s#����'���УO\�.�lx�Β9p��$��'d���.��	(x�`�G�=�
Ւ�'�\LQA��l��4"D�/:4�8��'^�@i'�N�/��%"��܇5�
@�'������Xb
})#N�3,��q�'R�bI�1XHi��]�.>�Ɉ�'��h�FH��?0���\�����'s~tQF�
&wiB	��m�$P�������*��)*m�o]*��p�P&.�!�D[�c����o�+G|�2#�5.�!���dHl��j��\��a�k̑IK!��&ytֵE�S�_�a�TDT$�!�DA��9��އ9k޹�q"�?&!��#�J�$��:HUX��b��V!�DL<�.������/�����i!��f��{7��@�de#'��5K�!��2D7�}�EC�&<�Z���E��~�!��<H��en�7��m�U�m!�ď&e�Qq�B�<T#�X��
�e!��HJ���F;zr�x�cP��!�$U5'�1� Jjo��ҩĭ)@!�$?[E�8��g��y�����N͝F!!�� 4�ʖ�
>m1
�x�J�,� �I�"O���j��J� �3�G�>�D�§"O�iҗ�X����G
1�`����Iu���	��&
�����W��ECb�V'!�d���Zx��dC�R����g(�!�d�
�4\s��M�4���fN/L�!�$بs�`�,�6�@Ec4�P�]�!�d��O��h& X�G��E���8/�!���ʪ0(0,��r���J��Ҥ�!�����'�
�V�z1`i�!5�!��s.����O%Y�F@���U�	�!�߻��x��ށz͜Yxa�R1k�!���B��h��ޯ,X���9k!�	4r��3G.�5j��	��!2{!���a��8c*��:YR q�
"Fl!��o>XT�T :��!+��W ^!� ,r쵚@�N�@��1dˏ_!��@&�`��n��1(ZA��h�=6X!�V aw(qc�,ԅ3q'��!�Ps��S���T���oZ	�!�d�Z�f'��!��aSU@�[�!�$�2>�P0�0�/N��A1ae!��O�E��B4̘,i� ^7(:����"O6������O�ب!�Yi,�$��"OL�!hG�k�n�yŨ̬w�D�:�"O���a�W�*HE��҄%"O Q{ӌى\�,$C�M9~�>ŘV"OrQ;W��*H~|��q�.-�-H"O"�1�&7O�PjU��%�6L�"O�Hy�%՟z��4	Rˊpڦ��"O�I�v�ڬA�&9��J^���"Ox�6��o�~e�b������F"O�9� b��F$0�U�2��\��"O4X"%E�lԮ�3.Ǝ�2�i�"O8ŋ��NG���GB4���"Ov�J'f�qnD�F����I�"O�z��´��`R=6����"O��0�;�|P9�[)",X��0"Om����tm��Ԭ�;��U+v"O�% "�˅��m�	��l�"OHM�懌(��j��FG�bF!��y!���w�l��7�=�a|��|�#yUD9�B�?q��-�`H�y"�бad�  k�,3�|]9ceˮ�y�ś%�p� ���(U��(�A%�y2��M�V� Aj��k��Uң���y�Ʈ��!%' i~��뒋6�y2�]nAi����c�N��b�U��yR��Y ��T̀?/��Xy��
+�y��M)&8�X��O4s�̈�y� �*;[|�0�U�n`bwo��yB�O�AȾ����T�
3Hy��+3�y2e_&i��8z`m\�{��)c���yb.�8]��Me��f�2�
SG���yR�\<}6�@��?6�y ��%�y��3����)��t  B��yBA�b�j�Cu*�4�S��N��y���[p�9�&��fP[�N���y�ǘ����(�a�H��:!��yr�Ɨv��� �;=8�}���V;�y��3��� �i�#,���˥+݁�ybA'=X��5@�=�8���G��yrj�	l&��&L+}s�y���yrui��w8��*V(���p?q�O� ���Z"kY��Y��дY��9�"OV�ڦ�͛?|Պ�C�
* ��"O.I���J�V�%C�#�>\��A�"O���k�,"�x� �$
X�+W"O�\�Ǣ\�3��tC���*ɜ}3a"OJ�;f��XJ���2D�ih��Q"OXq��f���p�A!r��Y�"O
T����"�N��$E�5a���"OT��P���z:(�I��QU�h��1"O8�`$��=i��\4u���"OL���艥L������^ ,�a;�"O>��p�L�\g�i����@�)�"O�	�g��Q�X�36�h�!p�"O� #^�ZG��3 y�b��"O����(Q!�`M`q�E�ش�`"O�$�'!�A���"�!~�y�"O��Xv˝Tb�`�p!�P��9#2"O�I�� �:>�,�!�	h��x��"O|H�*?B�p��b V�2�"O�Qs��!���V��!��Y "OQ�2��'�쭁 ��,_�� g"O��`�ǅ�0����A��&дx3Q"OĤ$�ׂ?�Lz�LQ�*����a"Ob� ��x��Tp���X;���"O<AY'�T3hX�dx$���f1�P3�"O�M�OM#��� �'��+ hi�&"O��!�FYF��;�E�.5ٖ"OT� �C�-����&W\��"O�CEj��T��j!/��@�D�3"O<qb��#LŦ�"�nC�v`��"O�h��^�N��B�]��� s"O�z�$�&GS&�Y�KށE��2�"OR 2󋈾`��d럊,}3�"Ov}�0K� En�x���{�xyYA"O��IwE�=D�,="�����E�!"O��iS�s%�� ��^,z�(�"O�3 h 0i�Д7cO���e�"O�ع@C)#0TŪUG��p��!"OP�٠�ы�HJ`F7n���;�"O��� ܛ$��$�T�Hx��!�"O�ݻ�C
,{��I��.�"i��m+�"O.)�t�s��(1G�?X�2��"O$��ɒhI��r�K �8� �p"O*lhe�͊Z��eH�o�
@�9��"O<��N9L���j6ُ@+&$�&"Oz�pl��n�Њ%�¹}6��"OX�2���Y ֌
siѰf����S"O�$
�Aڒ{��|0`"���"Oā�P\8j�	��ሏ�h0�d"O\�������n��$�s3"O�����D��\Y��NI��s"O¥��E���:��_�%���"OXDY�%�(:��-soO 9�T*4"O�5cK�H�Ҍ ����(�m3"O�嘕��?�^�tOګCfH5��"Oh���IC
W�1��@"d��"O�p5�T�/	l�:Ө�� �"O�Xf I}�<4	�g�O�2Yrd"O���DaB���z����C���!U"O�B�!'&�c��$z|1(B"O�l ���	ca�)r̊���T"O�I#W��9W�R�ӄ텃����"OF�1�l�T�n�%�����"Oj`IE���̼�X�BԨYz��"O� ������3z`�H�qcC	���"O.�aw�ʡ(�+���_� ��"O��FBL_��QP+ɰG��a��"O
 	�B?�ĐuiD�c�XI�"O4l�6�@�.Mx]X@/�=VI�@"O8�x2�P�F��!QM��Y� 5�"O�(���A���땟%̌Ej"O�0��<�9��,��ȯ�yD˄�`���MD�Y�h��I�#�y��I�E�~X�#�T��prД�y2��|q���T�4u9�t !�D��y�-L)Y&���e�7��m��W �y���Hk�uB^{���$	 �y�X:c`Бh�A-		6=q�F%�y�h�m՘<�R���-��l
d��y�"I��BU��9}\��*C��7�y�J���tEJ�(t�D#�I!�y�Nn��@ '�'rO:4�r
���y�3`
�L��Ϊf$s2
��yb��*;,��J �`"(B�i[��y�KA�J���V�b�����I�;�yrlҖ(�x|��ȋ9X봴����y2*6K|:���BM�?����,��yr��"{~(ەl=m�\�r*��y"+�,2 6� ���%c��QAG�y��A�:d�9��_�f!Ӂ����y«A ,(���*ǺP�ȴ:�a��y�CH;/��ق�Ԭ(`q��j��y�ǝ���Xw��#�XH[�����y��ϛar�����{ؼ���F��Py��Kԉ�W)դk�H��[�<i3�ч3�� e�J���E��S�<�eo�) �n	���L�T�@a?T�4�G�O"��8��)A��A��#!D�<�u�Z�疝pʅAФ�#!D��H&)FK�P��P V��"*D�*2���\U�$9PiΑiX�Cj)D����րd��� �o#7��Bֆ(D��(�6q����
�_��IQ�8D��B�� �f5 c>v�����i3D�h(�Rl�TP�ڪ	�8L�R$D�Hsg+&��$�e��1 ah�
G"D�`�����;�%�R 
Su�%k��?D��c#��6�����L�y��>D��swI ITZ�Mިa���i��&D��rŃ��Lp�Ы/A�5�`ш��$D�zD��K�Ⱥ�(�=:ƈ�;e -D�,��o�3, �H5��C~Z1��9D�(��h�%3�޵���<�4Qx��2D���rm�6����'kY;>i�/D���#�.&�HjS�-	Z���(D���SE_�X��dI�f V$�m�+4D�h`!�ߍ%�����2T+�ءF�3D�D�($�%�+ɺ?X�̸p5D��	���
�����Z-|��rU*3D�$��#��'�<%��D�.�D���n0D�$ke�ȽR�Fp�0��G����k.D���E�PTX �G���b����6�-D��A 	�?K0\ �(J�ts����c,D��	݊r���8��U?S)�m+b)D���B�^�:>��Ժ��	2�'D�����/5���k�0?cz�kF%D��T
T�<DM�VMʒjA8�3��8D��Ça�o~��1��A:�L�q�:D�� Z�� �_�i=ԁ�"!|T�Y�"O\	��?"�z25"]�fE
m�3"O�0p�&E�A}�1P��Ύ+�01"O�*R�M}0�j�!\�}� ��"OTdf�5AP@mR�ÈW�D=:�"O ����4�d�K%�<� b"O�`��Kґ!�$e���T$��x��"O��3*��H�h�A�	�H��Q�3"O��"��^-n���YOF-+�"O�,�bBW�N`񠮆�wK܈��"O6HksB��D���G�nCH�6"O���,�:<���l�*1U"O��v�K��J1�&�H��\��"O�ГaB3����I�%f6I�t"O�)0K�V(@�!���m�x01�"O�5;��R?�q�07��1�"OH��5N�'`V���;fj�,X
�'�� x��Bm��,9E؉+���
�'\h`�G�9Q^Y��c�3 � ��'�`��$D|U��(�C�J�'�<9�E�':F��+g�,��`�'�pؒF��-U�+�%�"#t0<��'#$QS��[&[�.)F�k�t�k�'8�E�U�U�tƊK�y���'&|��m�aI���X't�B���'v"$b�搭}~�Xv��v��	�']�ĻBn�	�¡�U���bVؑ��'::��AS�, jI%T&D�r�',ƭ�V��l-�Xu�N
PO����'Ր��#Ͼ�3b³O��<z	�'��m!�j9�
d��˳?�8�	�'^��[g�F�oF4l(wgҜv�~݆ȓp�P5C�%xB��#1���A��l��zh
]pl��lJF-���X��Ň�C�&�@AZ+�����.ɖk��B剤�n�F��4NSr=��m�.p�C�ɕy.��� gK�C,p����gP�C��!gjt�`A�&|heE��lC�I<<9���n�;�>�7�_�d�B䉓iP9xw�!��P0SG]d�B�	�+P�}�%�U�R�,�b��B�	�pԥ7,�96�\��V�e�B�+k��a�2���ep ������NB�I�U�.���P<Ҵ�H�f��+�$B�	����]�S��Uzd	�c6B�� 7��xc��^B�~�"Ƀ�cG�C���@��ym0�!G"_܂C䉇!~��oTv�Uf�ZH�C�I$C�J�;���@J���D�١5O�B�	�Ilp�g�2���e-�#;/
C�	�#��h���"*)���.�8�B䉭L��9���"_3`�ċR��B�	)��#�'ڬ%q2��Sa�)��B䉷�Ԉᷫ�*{��tHJQ+��B�	b�m�W��8��4�	ۯb�C�I.F9h�h���9��q�D��N��C��>x��$� -��*A�q�	�#s��C�I��(}[ī�]���T$�![(rC�	�(f,��|����/��wdB�I�t��ڡ(s��2Ӗ{��C�I,V�����8��Xp�O�J��C�	�^d�)U�#��"�� ]���0?фo�-פ���M���a�s��t�<���҈G�|�҅ܓ�0`�"�p�<� ��I$�ߚyw�4�D�&"22:�"O�%��ՠؐh�b
]�0"O��)���w�^�)f�\� Ӥ�8T"O��T�	�^T�9��"��{f�	�O���e�	#�였��ޠSf ���'�
��gS=X�(��`ьJ7�{�'7Ĝ�ӧ�(���i*+B)��'�4���9�x��)�$"�9	�'���3�۔H��!N_/	��p�	�'<&,ۓ�� �b�f%R��5��'^�U�aã.EbP�G3BXTq{�'E�T�JA1@�9 ���6��q�'�ΔȁHԭS Q�#�n[�'7dI���^hxs���P	�'�.�r� ɁXHT�+H��(L�h�'$�qYƬۢp�"�z��%���@�<�QG�	��<����j��Ԡ"�c�<��!$|��0�
�z�f�p7�]�<y��R�S�� 4��N�<���d\�<ËU�V`�#D@4Md nY�<Y��D���!��l{�] ��HX�<F�בt�����51�X�dQ�<���6x�M�uH)l�d��7��x�<�%J��>����ċ�;3�C
l�<���Y4z��Dn
�K���bD�Q��y"���%�z=��J��ɘM3t���y2%�:8��B o�s�UXI̐�yr�aBE��ā��4X�.��y�d�p��Y>�Y��W"F�=�ȓ&{� G�/dC�0S�lK)&�f���e�2��_��n��7m�
�p��,b�,٧N��f:�� NW�bX\��	ϟ�����C�}R�n��i���rrB_{��O��=�}��cw�p��Kp����!^|�<Y��0d�D�!��6H����I w�<��͕$�ڝږEK�G�By0p�[�<��N(f�>R�N#O��S��]~�<ٕ�ՐO�A+pKC�b�\�cWR�<!0�I�M�:��1���|�R͡a%��T��\����+?��I!)��Y�¥B�i��$�Ŭ�N�'a���94�˴&��w��8ǌ/�yBѽ'o<����A,ı*�,�9�y"%�O��(#��:ݺȁ�*�y2KN*\�~���%�*���p��yb���\���&���ġ*@'��x1x3>�9�늕	T,�҄�R[�0��*n��e�c"M�%��C������d5�S�O���05O��c����4M�7"O�����;}�4�0��6s���sF"O�� �#�?.H诏B0d
���U�<� �4$4Ѩ��7�Xr�,Gj�<)��Bl�*�!����D��`\p���hO�'ca\E�f�:n),1�ƩɸS��ؖ'o��'/��$+��a�.%���v(�:��zR��A�<�'�:A�@�9e�[#@�y���A�<1�b�<&lj�
#7���i�<��B��1�Nh���R
��%�d�<��O�� �B�Ύ�|0ش�%a�<�� �P��©��"�\�ro�^�'�?)YC�ŪTJ�<Qw�H,c�
hz��,�d�O���<�����k����J?i�1Qj9"��1;�D%D�0롂U�v��(��Y�e&�`�"D�t�aG�<4��h1j�w$Q�
<D�`Yh[�RDIQ��
!H���m%D�� @�����g�V�3t�Q>.� �"O4�:�oN�[D�I*!�XC���b��|��'�t���l@&1:�kIe���1�'����%��3K�2H�nFX��J
�'��9���S�n웅g�K�"�{�'T�H9�ƠK�d��%F��6��}A�'�Fј��>zƬh;U�9.���"�'D�<�rB��?SDT��G���Ti!
�'M��s�͏?������6ظpH�'5�k4��h��(��.ۋpA�P		�'O萲����ڪ�2�@�<i$��'t���E����2Cۚ1ܭ
�'"�����0 9TXA�+"����'R���sfЬrܱK'U���`i�'	2@�Pϝ=�B"a_!D�ȡ��'5�-����N+�̬f
�}�	�'��37�*x&��#�^4	��в	�'
|��f5X�"�xCX�z��'.�	���:Z���b��Cjt���'M4!I&cäu�DyҌ�=5���	�'cq(�*�0��P��у/�T���'jD�� �p���j:*G���'e4����:H�\��t��7%��`�/O�=q���z����H�}�ȺN�w�h0{�/D�8�B��izr5���KK\\��N-|O�c���D���+!vXٔ��=c%d��*D�h��k��j��B��3s&����)D��X�`�'!:0("�����Q)&D�SħS�S[��[4�N��!Yҏ6D���D�;<a� ��E�|#�=���OT�=����,7��'f�*P�:��th�Ȗ�L��l�*!���p���F�_.�0Q�!��!��5n�mbfK	��Hyr
��o�!�d F� �£�@$l�0�kb*V8Jk!��S�F�J������\�1p���ZZ!�Ƕ[���"�M�7s�b�@�ʊ8Z!���2�6�;kJ�V�ڴ��O��i���'�
uY��ɝhϠ��W��9����'z!�Ğ�W,�B�ˏ$/x����8!��0va"�J�ԇ]p8��+B�H!���.��U���>2��a���|5!�$ێ� ���_mҦ����O�!�� %�:�k��>�D�sr!�ב?���Jr�7�(��K!mM��P:!����7X�����^�WP��0?���׿d+@���A|
��6�Ay"�)�'E���R4+�	q%L��ES�:C��`��:�C&?�V��遌xc`T�ȓRsT� H!x͘���l�Z��D��IIZ�:G��jC�����F�DrN���e��=�5A�C�u��.K/�����.	Yש�3��0�%��:��(�'�ў�Fx�&c��ҡ�
�����K��yR�1���A@�<3B��v&���y���g����-
��Zf�
��y�-N�[l�;'/֛nG�)��'��y�`�F:N; A�<�p(+��-�yR��,70�j�W�;g��(�.ɿ�y���;U�ȍ���(. ɤ���y�>A��Ƀ��4�&���g��y"%�)I��37nH�1%��+��#�yR�¾�R@�5�W9S����'���y2S�0�ؕ��X$E����"���y��[�h<\U�$aX9>�x1K��y
� ��	�mW�Ex�Az X�
rZ��B�|�'az����`D㊛O܍���@��y�_�0�b6�$|��I҆���hOq�
(	Ƭ�%/T��O����=�"O@ݛ�'6�H�p��Lp~��"O�E{t�]�_��tҕ��-B](�r�"O2ap!Â-V�K3�VN$�+""O��X7A�lӀ��YB�-���|b�'���#5J���O�9����6͐��!�CoI fFw�`@�Q�߼ y��I��(�L�Q�/�(D���p"�y�"Op����_ ���JˑEW8̐�"O\Dk�iU�qz0<a&I8r���*�"O5�Ί�P@����ҁb���'�:����{�&�ZG�2]�B)C�'�2���N�Ԝ�f��7V����/O��=E�䀪�f\��MU.1F�P����?���?��<�š�&EvL\�p�F&'j�{i�Z�<A���iX<��FOА)��I��K�<�Ӛ34�J��V�fPb���E�<�D��$-\��D��xU��"�Ln���?��o\XGJm\�pV��1N��5��ئ�C�mצW��X��,+�PA�ȓW��	�茳3�% VD�Gt���ȓOT�!��*B�JaL���VNm^؄ȓ)'�P�sB�r�H����KѺ��K}T�Z(���Eg��~�21��Ӓ'*�<�x�J�+[%O�2t���O�=E���/U8L#��7D���'�өQ5�'ў�>}8p
�=l�!Э[b:H4�L7D�x���KB�Z8T-E,hFLs66D��DJQE<b�ȠJ�C�Zh��2D�`��e[&�p�d�U�^�)�,3D��!B�.tY���F��$A,D�p
�呠n���i��Yʨ��$��O|�O����O��=yd�P$O�B��4L^"��}h#���?i���'p��`��ǲ�̜�`�L"]�ȓe�n��#�,hkn4diE;1��ȅȓs�D�qp���L�.�{��S6���ȓ�|\�ĤٝZ�x\suK�1{ؑ��9�.�A�g;�<u�G�ǖW1>��P<��'��"֖}k2쐎n_>�ȓ�������B�Q�"�(�H��'*�':�\"��O�1�&����hR�'��Y�t^�0�4�#���"�
�'�P�0N��_(�٣�N��y��Az�i��t���F!!�y�Gb��å��
w���K���y��H:\Y�)R��'p_��TbL1�ynH�t;e�Y�dlL��!f���y"
P��YeÖ,XZ`�Å��y��!
�h�x1��Wդ�3B*ׯ�y�	W1�s� '^�^0�1E��y�@
tH�DلbU�XO<`Q�+�yb`���lp�G�D�U�`�����y"�ʭ%H��[�K�29G�9��F�7�y�l�f�N=�E�]?,�	q���y��'c\�8j��B�bF�S!=�y҈
fi�x���tI.(á�R�yr�˨@C�9u�<j��Z�"V�y�A].����2FJ�`�@1���yb셍c��P:�(��-6��HK��yr+�1�R�`����$*~�"L��y��D!2�]a!+�$0LHM"QJ�y
� ��I֏
��3G\� ~h�0��'��3)J�9���P��8�e��g��B��%k<(�14���壌7"�C�I���ۀ"A�a�
��d��7g�B�I�wj�J�<MµJ1,�7@�B�;�*�y��(@�U	D�)c�C䉵D�@��h`�!�ʈk���H��	�j�2����Bw�B�T�J� ��B�I�'�����bv�9x7K�,���ȓaF$��B��<r�S&��t��8���pQ�F�D�����'�ń�	;��+b�8g!�ӫ7/*U�ʓ*�‡G�F�8�ird�<D�jB�ɑ*R� � W�&+8�0��1�VB�	)o�U�!)]3K���	1GđQ�����O�a0��ׯ$ʆ)W'��X6 D��%/�*B���aL�;'Ф�;D�,I��Ʃy��"�F\o���b�i$D�a�N� s�����3W\ Z�K'D�(Zq��+R�` �B�6"#X��� D��%�3/"<�p7-��S��	)D��"�a��W�@1/I	����%�O��D�O���F�1/d���T�G6`n~���&!D�����$=Ob�hA��99�n���,?D�\˓B�M�� Q)��m$X4�w9D�,Q���T��]���V^F0�D�!D���o�`�v\�ec3r��*6� D� 	a#`���� Q)Y5p�`�D4D��P���"N����iХ9X���?�O��d�Z��	Y��^l�|+@(����C�	g��\�!_�0l.i���?P�C�ɤ��H�4��\���%��v��C�	�~�h��5,Y�A�ؘ�bB�+_�^B�ɑ�y�
��M~���j�*G	*B��$>�FMa2a��M�t�B6�*$*B�7L���O�U�&����
W����z�`;�!�(�h5k���+J��	�$=��K���T�'b�QV:qM���Ê�{5ja�u"OT=��݄>�Z4y�@�$t�:�"O����4gp"��n�E�H�"O<�*@�֨�ȑ	5M/.�6(��"OL� H�h�8��%�˃�ע$H!�$�T���7m��R�*H!�I��d�!�s���	�E,q��˦EL�N��Oz�=�+O4�jU�(�| +���80K�hs�@�OrC�		���P� ٣6kbБ�FǛb�.C�7@^6Lr!/�_�Z|�����C���̘���S�S�p�1G�Ήv�B�	�O�Lzi@:2*�8Y��L6HC�so>E����?�p�Ŋw�*C�ɥ�̔Q�G��l��T3A��=�H>����J9""��ۅ`�Z���8������$�Op��'gǚWB]q�u��C"O8�k ��g(M�sI�!j�|@�"O�I���Z�zU��)�Iy�@"Oƹ�BO�����лd
>��'Բ�s���:��L����v�1R
�'�0��Ņ�\FeP��\�h ����*��p�΄�N'2�a �@�z��'w!�d�DZ.�( I�q�9��]6W�!���9�����ƘV<��	C}!� �ᤅ[����S�^�Y���]m!�DS�L�zd��܎H���aţ o!�ʳ`�b=���'`4޸XPb�t^!�� F�J�l�]6���VO^2��9��IH>y��6L����D�Z���bv-:D�����r�ԭ��>c�ĩ�Q#;D�@3fðzD�h��K�Ab1*:D��� N�}��"�疓b좥�e�+|O��<?�4�/!(�'� ����'i�i�<a�J5�h�f"_�Nn�|�<I�ϋ"dڅ*R͟1�D��a'v�<Id�(S`��)E.��v�.}@R*�J���hO�-��̘��Ņ��YD(� ��ȓvH\m
���w�r;��QRч�Ej��y�i��֝:Ao�;Lr�1���v~b���n���G�NH@�1W��1�y��Z7f��Tb�?w>�`&.��yrO>s+j��昤8a4݋e�;�yR ��	�nX�F�ڠ[�����?���0|"�$֣z�tQh�" �@��5`�I�<Y�l���x�Z`JA�(:�M���Q�<ђ�29*F�[`eڜP��x#Du�<q�J \�\�yA OH��IS�z�<�#���D0.�HU��3A���f�u�<E�Ń>�	��%4��rA�^����?9���O��2S�8"��Y�H��y�J!�DL�@! D�|}̘�rmU}8!�$RSG�Yd�r
x<��L��x�!򤀉f!01� Eי#M�r��<(�!�D/�dH2MD&=��lS���Rv!�Q�2����J�*
,"�FО1S!�-}>�`K���u&
�Ge!��Iy�ԉ�� �M�BdΟ6!�d��zU��wD�ٔ��:�!�_I����ŕ���h� ٶX[!�$�+�p�	��Att0��
�8^!򄜚R�(=�Q��xT8��f���!�d�F��)�cO/-�� ��Zk�!��úq�>@a�	�	[�`:��*m����#?(��G��="��D��\f�B�ɉj�v�Z��[�sVD�T�,�B�ɟ\&}��.ٔT��Ce[V��$Åa�M!��)�¨�!fĀ:(�'vў�>y+�&Q&eF`k�ɚ�`�R8y�a#D��5D�Xb��T+��u���qN.D���C
Ō6�Z):F��&~�����L+D��+�]��D"�RYpƁ1�.D�����N�8o���ǐ�G>Hr��+D��H���5Zz,Z�jN�~wE��3D������s$e��J�@��q %��9�S�'A�荛aa\2R!8l�5H�2�̵��~8��(�(T��X]:R	�6B�ȓ�h�uʉ��n�(���*$fŇ�S��p׭�N�������7�ɇȓ.�⁹7�G�!�D�
��(��`��c��İg�F�.�t��˷Mg���ȓ;*i$����԰�C5'#'���IS�Sܧ=|��J�g�.����l��ȓU���0���+k�D�4��TqBh�ȓ	F��+/�<p���4"4~5�ȓ%�ؐ�g,�;^�$H҄%M%�����;1"���Z������T$\��h�ȓ;�Ȩ��KX��X�▥״st������Cɸz�@��!E��q29&��$�@��m�O�,;%��2�TAy��ջX_,��'0�1ѕ�C���3-9ϐm��'S`�i��S������!<ޖ�B
��� ����A�|����bT�
�3"O��A�ӤI>~���V�O�%�"O*X���3M���Q�^�Y4q�"O���6.��"rؔ�Cb]i�l��u��m�'���9g	߯@ޤ��C�����0��"OYx옲v��(X������q "O��Z�AA�h% -��쎜G�V ��"O��k�?,(��C�ۜl|�z�"OHa򧤃�t숍+���zV��"O���"�$�p(��+
/EH�Y�d"O�	9�i565�8�aɳvA:�@���S�'u�D�I�܉g��3 \���LoRO�`�ec�urqɔ���:S"O���4�����I��]�p�	q"O�A:P�ل�F%��I_�k���2�'�ў�I�<&�T��J�y��l��M�ul�-{`�Og�<	����(�� ����"^X�<Qo˿w��� 5a�!g�Q�<��i��}��Bh�c�\*6AhB�	�K�x}0Ī�)����P�%XBB�I�/��7GB�X���Uh_�3 |B�I��m�2-ۈz`H��Aʎg�0��d�<�O��e�D���Ub��"Ӫ�q"OB�˶*?� �['����i�"O�r#Q蜄�1�_�9���"O�"C�L8��`�8���y"OZ5*t��
�h3��?ﲔ�C"O x��K/΄I䀀>Z:��9"O2Up ���x|r�+K'rf� �E�|R�'.b�'��O���<J��湊6�*����B�4P�	�'�:x���1wO�p��ʊ!ON��C	�'*�"3��n���[�OF�K��p	�'�pD�)>�<E�CP�(L��'ָTx���$���*M��d�r�'("`M&qb���g��nL�'le�A�ʅ0e�؇�ܞx��S��?Y����OJ�S�'��x��!�4A�^xa�!��E)��	�'ڲ���쓊5t]�S�C�EI�'Vf��Ej	#}Lh�n��?V�@B�'�̝��ؼ��a�*=�2H@�'@��i��χ#���%���5�$���'�T��ԍ�w��M�+K�3��"Ov�Q%*  �xP�7B>Vn�H��D&�S�I�=�֌����5o��h�ԩ3�!���!Op(�Mx%.�&ɋ�B�!�dHR |�G 
6$����Y?3�!�$�7f݆a���U���"H�^!򤝖o�h�2'��[����i.cA!�u�mi��JN��\��
cC!�$�O���QW�wh�pZ�@Ɲt5ўX���e��<	t˒�D�h��'K_>�|B�I�,#hH�7�Ù,��U"��DB�I�Rw8�#�|r�_)O:4B�	J�0�;BbJ)�P�v ���2B�I*��u��C#�)�\>(�4C�I�{V���	W�r����L#9,C�I9H���V$�K��(I��O�d|6�?щ�IS+: z��O?D��H&f�j�!�D��5k���(��eƕ"�!�E�H8p`A���aŠJ�H9�C�;y��׭��_ ��
�BC�%aG�#�-G�f���#��-�fC�ɦ"�H<���[�� TC�I6o�p�UG�
�D��w�I�T�?��� ��W%B:A h�3��ݱyL�YAD"O�1�č,�V������3D��"OЅ`��ЕM�F-��@M=!����"Opl�C��ڲw>�!���7D�k�B9g���+��b��7D����gGK�[��l��P��7D�L�Df�(�J�٥�H�@E�x�v3D�tKפ��:�SB�k�t�"	6D�<db��A��݉Uk����(��g!D��b�K���|aJ�q�r���"D��Yj��GL�%A��B�!D����=jv��a'���l�`�S�2D����]<}�⸂�dƤFJ�g�-D��cPGC =� �0���.cd \��9D���C��9�����Y9���c �8D�`���+W���&B_���ɲi5D���P���ZyI�
ԇ{��1!�@>�Ȉ�n����VWz<܂s����u�0"Ox�?Cv-��Q�L��Q���y)˘��	0�
�	����gN�#�y�HV-;�r庥��Ut�e[��O�y"j��N��W���i�y�W!-�yB��`��Ly@FU!S�q�'��y�	�\"��EL>~�ά�6b�9��'���O
��D#Ҙb��8'���BP����yRjjcuyq��&fld�qЊ��yBh�>T�<����]f�!�d����y"���v8�9ӎA�Z)���g΢�y�.�UH9cS6{8�LK�F7�yb�Sd( ���y����Dm��yr[��pe���m~�Dh�&����?)���dL܄M��J�h߼[��K���?Y�'����U�)`�ɹ���.��-*�'0B�@�fAg�C��
���'nf ��V���1AdÇ �t��'ֲ�s�4g��	�3�C%O��Q��'2D	0DŖW 40A#����Y��'ͨ���Y	M!ތ��ˏS���+H>����?açQg�	��A���fȨ���E�L���I~"d�)9�\)c�%ʁ_J:m�C�D��y���'L�:���=Y�`i��$���yҧҸk �� s
��`d�!H&C���y�C��v�R�H�`���`���y��. !,���I��/�8qеJ���yboϣh�zA+�-�D4�u� ��d ��|b�y��L*�1���\�}1�yb�;)^M��`^]l(�x�����yB�I�X�S���bM��+=�y��� ��X7�f��TQ&���y���a�$P%g۫g��x2v#P��y��r�i#$Ğp�[FJqI�ȓɔT2��C�y�f��O�D����}�$d��)Ȧn�5
 �>�
��9�ecK�%oYp���J�8aC,|�ȓv��bs � I��]�d��"4��ȓqe�%����8wT8Q!�"B=FeP�ȓ���"��Y2R	!��t�]�ȓ@
��F�RKF���%R�m�h�ȓwD��{�^'8�� [V%��6r-��Y �y�ʴ��#rE {f��ȓ���e���A�4��Տ��̄�I�֩ڵ 5��9Bd�\�0��	�ȓNӂك��:V?�hZ�ϕ�DT��[�|��#Q*�i�MǘQ�*���S�? ��"�'D�@���BL�X�a"O�����6zW�Ȫ��޼D�N���"O6���ε%�u��kQ��N�!�"O�Qi ƕ5@�� �EQ$+��ٙ�"O���ÍH&qA(�U'�B�`pq�"O&9�$��w6c��F+��'"Old�%e "�9Q�qS"Op���g����$� �5�"O a��H���3�T�P$bq"OB���M�R��M
GZ�|�b `�"O��	�����,As�D�I5�"O���N+��#T�_�e��<��"Ov�{F�2"l6�;B)C�k�*m�T"O޴Ƞ�J�>ȕ@B*��D��#s"O��CP]:� 	��(�I�HI�"ON`!�ߊS��*���=�H��R"O��ŏ�;z��I$@��XӺ�
"O������/ +���0�$����"O�%���T7y�����fRfn~4��"O>�ʠEO��
�BƳC! a"O�8#'QbN9�jܡ!Ŵ��"O&�t����V��ɳ�"O:3�b=9��(��.B(vy�Ԫ��	ϟt�'�1��tF�q���c��BQjPHCt"Oĸ�'�/l��EDH���"O�QsS�
 ��eÃY�D���"O�P��2z��usT��B�j�"O��� ��E7@���3� 5��"O\���
$Gc�xb�Ԧ�
�P"OT�q��$��0� ]�
��ȵ�'���+�Տe2����	��1d�%9��$�O���B���IP�$S���$4W B�I�tW�1�'6�j�'F�
B�"B9'�
���7�[�O7�C�I�R��ĉg�/T~�%A�AFxXC�I�9��dZUf�'��1�����>��C�ɹ*����t�\�=10����Q�zB�	WR��ضM�N%"�i���#H�B��Dl�l������YWϠe[~�K3�'D�pQ���p9���L=}NL	f%:<O�"<q ����'�=g��MR�� [�<�B&��{��q!b�_���r�j�U�<��nY
��0CAM���@���y��V	,������4��T�"3�?����h����%��B�R/_�b�j&$�?4�}����a,��#�\��d�N"���C/D�$j�*�?�} �o
.�m8��2D�k�`�^�̨+YD��)Ƅ#D�h���֜ua4�Z��pI��;D��F�0x.^m����YY�U�d�8D���/_mj8&�	%��q��<YH>Q���O$��D�b (�'�An|����'R�I :���I"O�aG�m2EA�2EC�ɺ@x��������v� 2�?a����#;�H}Qg&$�i����I�!�䞨w��*'�<y�,L�Ҋ�q!�D�t��$�fc�9��ثA@�y4!��0��n�u��<���Μf�"�'/�'+�>���l�����W2r�\��@O�t�0B��Eh��5��I�)���:�*B�	�K��b� � 9�"${r.
�btz��8�I��G{2@ѓ.D��G�h�(�ZW�B:!�D�VG�,�G��$���� �-!�d��Q�����,xpnH3Chȅ�!�� �e��L�FҤ	�+�� Ja"O`�@��C�$���r���}�$i0#"O�qya��MR24k삠�(���'z��'N�ɱp�b����H߇T�#��',axb-��W�}�D�]�V�x���Z��y�����e;���P,d��g�ǭ�y���z^d��� ٿOZ����	D��y�lQ�!��b�K��5�j�a4��!�y2��[9�3�W��PTsc�+�y�Ѿ�s'�Q
�Ε�!����2�O���bQ�t�f�0��<(��Sc"O�C�i�!�h `Uм`�>�4"O��X�f�=�
$�0���	r�!HE"O���J�v�4rd�kLԺ%"O2�9��?�"͓"��Se�T�"Oxe'ǋ^�n���S/XyA�"OJi��&��T�f�t
��K"l@�X�D��	�8��B����x���qs�A�4�C�h|��� g���x�Ã�$C䉼qI�P����喍��CƶG|�B���YcGIP
�fq�5A��B�	"h���Em_�3�(�Z/�)�C�Y-���f��:8 c��-�vC�	2�(݂f*X5/�Ӆ��n�2B�ɎZ�h!c�:Mb�$+b�2"B�I ���+��ݾ��ISu�d�B�I�{IZ$1�&o]��{����C�%9���V�F��e�`"� \�zC�|�X Ggj�N5��۫+�PC�ɒP��C&��5�2M��Y��B�I���Y*�Ʌ�欣�?A�<B䉆c[x�e-���s6�¤	<B��6����G����C�E��tJC�	�#Gi'jbx�KEᐐ!e.C��	)V�XFX�Q��i�Ȑ�`,C��^�h@q�I!;�¬#W!ٴ}�C�I�>Nl	�`�4����LH��yb��#�.=A�$%{r�,��Cގ�y2���v��*m�>���ز�yr��WZ�A�b��3��(�0O�9�y�ŏ1-8j܊QȀ�Ɛ�5�א�yr%�T���K�h�՘d�Ϝ�y"�G�H� ���`+2�z�M�'�y�#��P[���F������"D����,PK4��q�qU�y��	�0(��h�-�&lxQ�N;�yRd�	#�9!�F.1RDp��5�y�II����j�n�'�e�p�˙�y�\�i�q�Ug֯z��X`�A��y�
�3{�iq�H�<	v�QcN���y��O��z)#>Tx]�rL�6�yB�Ha��݁5
�N����
��ybl~�8|�䌝�?C��	ՀE1�y�T�X\FՋc�PE�4�d����y���\G�@yu�?DL]����y�Jt��� ��.1�������ybnZ ]C�l;�Ӫ�΅:�.9�y��ΠQ��yw)�}�&���yraܙ%����c5���F��0�y"�ʌv�B�Kq����^i��ۍ�y�LQ����+Z�W�j=#�n+�y�B'OP"���m� WP�p5H-�y�B�q���E�pTX0��y"΋:Yj�D�Pl�(<����*��y
� �lz���/䀢�ŉ�T*"O�12�C&o�`��`c� w��YBT"O�4R�T�Z��uxw�ތth��&"O�x��]=Ib����֐����e�<����	5�a�e���Y(����y�<9��)+6�xa0%��k
J���c�l�<�F"(h��5� ���x5v���$i�<�@d��H��ܑF'�"�#։�M�<�[+0�4PBခƀpsEƖH�<�P`Ls�����ʢ�l�{ �D�<A��G)�%�AB��F��"�A�<Ѡ-C8U@y�q�ɾO�r !hM{�<���1��pa&Ȁ�1Й굋m�<�v�O*GV�;q��0r�
 ��M�<��?t0-����K��m�+W�<q��.- d��hȩ9��@��B�<!�A�>3���KA��jn��zpk��<�`�a5���W�ݧ"~�ҦD�|�<�Z$~:.���s&YBծ|�<Q��4�xe-N�
�|͢eLC�<�a@2�u�$ꍀg�,TzwB}�<��oB�:��Qi%-k�pb�Ey�<��U5!�d���S�{��i�C|�<��B� b9��Ν�At��F�^�<�4�@2V\��"Ӝa!Lh� g�E�<Ih2����G=�!6��D�<�5�R�A8��{���<N���PP��B�<��EB�A�7aҴY�^U�<�%�(%@��Hs.A63�>�H5�CP�<��>8'�� ��&t{ �H�L�<��a�NkH��h�"u�>�s��OE�<�Q��'vb���l�"	2ܓ��e�<)�� �?q���(A�րYa�[�<�`l��(ؾ5\4\Bth�Y�<1��K���RB�T�>�+���A�<�E��v��Qa.S5h�@H���]@�<I���1岬k�n5!
�|b4��~�<A5k�>nE�e��R1f��(:�~�<��-m�����F��-l�c�%u�<d@���r�C��TB�r��l�<q	�-oR:�A�酿c����@�e�<q�)�xFJ4R�� ��������`�<9Ԉ���	`P��F&��ֈ�E�<!#��$Q＄�c)��<� �h	@�<�rD��&#����;Ș���a�<q�A�L60PS⍞8��1��M�T�<�.�	�9 B/�;�ݫ�)�i�<��B�1�� � ��%"�+d�J�<�'c����2 �P,E��Y� ��]�<�V��(�e9 �ϼY��r�<���݃U攠#�KK�\��b���w�<qv��3^�\a�T��>�v� c��<)2O[�{�
abFďtr2��`Lt�<I��T/D�|��F�D�
�@�&�Y�<���"���H!k��U"�遅W�<�T�L ���ll��EלYlA�ȓ%ff�0�ߡ#��uq&�ʢh{�����(it��y�ެ:�ܵQ���ȓho慡"�"��� ��/?�����N�d�X���"����!�\���I����ւK��mK"�#VX�ȓPR����.��{��k��٠R�5�ȓ%���J��$%R��
�L�`�ȓW^(p�ѿel�ч���xP��S�? �@�iWrE���Ҝ1���`"O���O�4�xqC��L�HX"OV�����\x̹#Q�ܧ3�E��"O���f�#Z,�Р%�'�>�0q"OFB"/�5^�d�h�F�!z��E�""O����A8Jt�X��%�)|���x�"Oz����vZ,jQ�������"O����$J�2< ���V��"O�C"j�@�vQ���J0\a`"Oz�q��5}��!q��BA4Dc"O�0�(����i�ЍN�2F�s�"O�X�El���5fJ�'<�0"O
�8��H�^r�y�B�s)��'"O.�P�惙_���z�а��W"O���L(>p �B�%�|Ը�"O҄��/˘u2El1�䤀�"O �:�D+jԬ���d�� @�"O6I	�Ș]t\��$�łe�����"O��؄�Ѐb⦠K�CF;����"Oz�3D�D�)������"�x��t"O|��g���j�.�CU!T�`�"O�L)aAԸq��)�B_��(h"Oh`s��	*ot�09�O���Q��"OȀ8����1�fDa[�E�l�n"D�0��矄&��L:2A�`n�ͨ��8D�x��
Q�)��e��E䪕�D�5D�	Q�� �p�;p��	���x5O D�B�a;(�(�c�I$}JX�u�#D���E�(|D�c���C;2l�!D��ʗ��;9=d�@lA-P8P��>D� S�H۴_:�:�+��Uv���B-;D�Ȑ�N��L,�&��><��dm-T�����:$h�r�,O#2�dp4"OR�X�UF+ @���[�*B�Q؀"Oʴ����%gj��,A>���*O*aࢃ�ot�<[CG1n�%i
�'NJ��EOw�颓��\j�d
�'qb�{�������G��
�'�N�H�ʞ���X�BI:���Q�'�����i[�9��膋ƫV�Ex�'����!���s���2��#I h9	�'�:`HsbHɀ(	 nԕ?:����'*"�b���:s�h��º;vQJ�'`��X�,��2q�I�%ۈ��'�}�F+��C@\�k�@Z5#<�x�'�����mA��-�g�K�J�<x�'�2����������g˙L�Z�'��A �=\+D�Pf&�&	�Zx@�'������Gt\9v�	�|����'n1K eh~ĸ%1r	:�"�'�n�h� ϛn��H���k�4��''���tC_ 6���p� ܾgI�DS�'��as�C=:زlP�@	L\��
�'}椋Q-]��v@!�e��L�}�'(d@�.��t�ҡ!�d��K��}�'�BU��O�QmX����A�1	(ِ�'���Y���]�$��]��'�V�Ӯ�v�h� ��^4��e\���<����*H��� ���L���i�&G��}���������@��A��I+^ك�7D�HCD�\9kT�T&иul"I�i3}R�)��9v�LIq� �qWH��f��c�؄�I\�����q�ӥE�F�����a?)��P1��1�D
iC�W]�<� ��E�?W��R'��\0�!t�'>ў4�n3Wтl��N$5 ���!D�<��E�=z�t���b��I��"D��j�&B��ܨA�%%fN�x�G>�OP˓���1��_i���!��Q."(�'>R�'�x�(���*R����P���;���y�>�`�3$ -�D��?�y"퉲Dr��ᗉ	�(y�@��.���OD#~s��	#*�ؑ��,"�����D�<��eV#F�Q4g��f�+ph�}�<af�U fB�<۵�C"]�n�EX� �O>��Q�
o�Q�whۗ��݈[���� S�2e�����HP��I2���5���<�;�(�2u�$�I�e�`��&�-q85���:D�$"a��[\�E�a	�6@�8�9"�"D���@[�5��1��Y�\�ڡ��H D���gNY^����?�~T���3D�ԨQƁ#`����ޱ@�L|���0D���*W)H��)��
ۗ# ` �7
,D���ƙ.
�zE ��\��'+)D�\s�n�1g���t�V�
��*�"'D�����C� �l3C*�2 �:ykP�$��hO�S]�:�k1e�\-�8�ƊP�kb������`��J��\v�6� A-C|C"�n�ş(�?E��4q����7/�)a�����?�LFz��~�b�;mQ�Di�D�<H�
ف6�[?!P�O:��dOC��n�Ix��[E(5P��r��1O\��?���JA��P�%br��⤗pH<I$LV2?,(	�mB>� !J>.��	h��,��+����x��.&�S�A6LO�⟬z&�D�K���pL�Ȝ�S�N�>)�>ъ��wn�q� ���2[Q~���[j��&%^Ni�!�@���s��p�>�ۓ�����+��s��9K���,[�B�I'R�6�!4���{�\Q ���6Y�C�	?/����bED���$��eɘ�DUz���I$�I�n��E���4(�$��"^3�bB�I,$��I��ȞZ�K'��ŰS���4�L	Qr,@.��c�Ƚ8;f8��N?I���ϙU���� E�a��-�&�)���<)�d��NْC�L�I�.L� �d�''@8Fy�Q���F4�D$�7"�6����bO>��xB�. ]��ᇌ�S%��VA�$D��o�P��h��q����T
�+4D
=b� ��'�qO�"�O>�"�'��fȅ�t"O�Pc�	ͬ|׌ԁd�)~d���&�>ъ��)�	<����s#�'.��{���fF!�D�A5��5�Ȁuwe�592���)���`vn�*T`JD�L�~�p0/9D��`��_H��;��ؙ|�@���!x� �?1�ט'Z�S4K�:���@&�Z��ML2#���m�H&��ib�́53Xg��h#��!�v�8	1H�S�O����SnS%,��rO0uf.��'k<C�Ϲ��P� U,q�ZTA�'����Ȅ�V�Jm#�B�<��1�'�s��6�P)��A�
#|uy�'�����	 0uL
q�-o�{�����&eT-Oc4x�f	r ��#��y2荿~_nT�#%[oD���&����<�OR�Ђ�*I�����m�3.8D�(��	D���	K�1[��'�+�6ذvCN\$!�����+�C���� �0bA�1�k��ħ��I�"xRa`ff�;_�썀3'��Ɠ5*r�j� fPfru��Vٖ��	�<�5�)�~�H?��S�? h�ℏǣ\ŠMC7�C���S�'��̧>iCH�h��$�T�R� ћ�l�[y�'�Jy���'��5*膤XJ`�CU@�)b|����D#��?��ɷ1�rϒ`�$��S@�; )�U��!8���s�Ж*a\X���y��C� I�#N�E��ܐRLL���M�g�Z5���?NIt�Y�!Ewar�O�q�g���̦��Q��j���'ԛ���{���U`ި Y�yA�g�,sK�B�I"1��tS�&�)a�z8 ����G���<E��B2	 @L��ѱ`EN�T��y2�>x��sLŖ_��I`�lÌ��'�$܅�I<#�n}�fi�'	L%��e�5|ߐC�-)�H|ˇ���`�`���^%A�NC��uV�}'��9iE�� �Z�RC䉃B�ja��۝'��*v#�
yvC��3k�^tz�T+D��x2�LK���⟬E{J?����o�B�+k��^�(���:D�� d�!"�jLAS�R�J�X�{Q#7D�������J*`t ���t�v�	�A6D���U���x�TykR*�oF�tm(D�04E~�U����9XM�%D��@�e��Fpd3�eݣ{��l���"D�T��E#p��� �'r����,�$��1z�%�$��}0�Y�A�=H���p?!��܄mD��[�F%Rݓ�
y�<AA ��`� ��2k_R`��I�<9I��h�݃��	�@��(*���o�<�g 'i��xjgk�
{\z��Jk�<����(>��SSÔ��ZÔ@�<	Ď̂qp�أLN��X��c����?����:%T�a;��E�}}��3�O�X�<a�B�'6�L��gG<l����`̓ט'�0�|�JH�f�PdIp懸F��]9�/IY<��85�a�Q�p܀3cPD���'�ў"|*��-,AD��KF�΍0E��v��D{��� o������:�KebK���'���$�&
I\x��BMD�9�&O�GR!�4���2�*G*>�	i�M��!o!��ڶI7l��%�+g�RD��ƛ5���gy��'� �ca!���\��BL�4�
�'��d�`�ͪ�t|Yʈ)t�p�b��$<�S��b���&��Htb8 �jɛ�y"��]�@����%,�q���mZ�Q�Q�"~n�$2. I��ژ!�4���H�P��B�I*�v�jA�Z�rrE/��.�B�!�T��N��&��YS��h���	v؟�k�%�;9B�]��-��kM��#5D���1w��үO�=9�'�J�<��.�
"�9��K^j	.��#ꓢ蟂�3�@�$v����$9�(;�"O�l؅���.%.(z�OD�+�aЇ"ORT��oÞS;�uZP��fQ�"O� �[�v�`��P�Åh�au"Ox�Z�)ǈ{��K�%*�@}J"O���P��	4�H*����^`A�"O��GLΟAJa�s	; �h�"O�ț'30PTH%ŏy�nppE"O �qf �z,Ȅ��m_�N� �;�"O`\#�#X\4(P�ވ(b���"OR���������wϞ-T��"O�P�T�*8��i���8�<���"O�1Ɂ�7k�vd�qDH#h6bUc�"O�T�q,V���-�Y�
� �"O� �Q����4X�HJt��"3r0���"O0�pqBD�D2E�sѱII\�
�"O�L GlL�Y��M����RJ7"O��`�śH��Г�+�:^$��"O����Z�0�٠�, �2�"O��s���d� 0���(�n��"OmS�Z�&z:Uб��\~�\R�"OL���ώ�k�6	�ݳjl8��"O`�x5Ș'd��"dH�N��s�"O� K�G��d�"�� �k�V\@�"Oh��AN^��y8)^-1�<i��"O�A�a
�$��
"G��\�\H�"O�Y�W���]L	���U��P�"O�Q�EW|�P���!8,Y±"Ol:s��2_��d��I�%}���"O�Hb%*�>����e,z�x��"O�օ�Aײ�� ["l��p�"O�<���7Lr�m�`�,	�"�`�"O�	A	������Ώ�ʆ��`"Ot����DZf��\1���"O���uk�m�F���<d�p��4"O�E{�%F�Y�e��.C�f�(Ɂ"O H�#R�_u�d���ƉC�V`3�"O
���A'+���Y3$^H0��"O���gJ. ����~��Y�"O�L�"e�X��Q��F�-5bΔH�"Ozm��)VT�bd�3�W�Z	�p�"O ��Aǋ��4X�m��E�  *!"O�ya�/5$�p��6%��i����"O�=�`H�6ލ��ж�`�"O�I!`��5yC0$���Z�2���"O��b�S�)F=��I����9�"Ozi����S�ڕ*0j��A��Ը7"O� R¯ײU0��ɧI�E��tV"O��	001@�0���"2�X�"O>���Y�+�2� ��=g�T�"O�]���T6~l䱁�ѕ*{~(��"O� DȢ3fA Ӎ��`��!�"O4���D<Hf�a̙{�rܙ�"O8I�!͈�c�f���i��t�$)I�"O���c��_�����G�2p��"O&�s�B$_��=A��:X�ƕ0�"O�l�1"A�RXÀKL�[��|qu"O�4��I 4E2z��'I�����"Ot9Xc�T�s�,�y��6$�*���"O����/I�z�Icg��$���0""O���Ǚ�3 ���Gm!3*5D��;��l#��3W��v2��t�Nm�<�"M�A�"�QQ"PM����c�w�<��J"f��e�Ň�"4��x2�	Y�<�`C�8�J��U�E8�| "�c�V�<I��R�qf��IG?Pxyn_P�<�ևp�Lڦ�;?�B@[��N�<Yw.&bǘ��G��81'�L� j�R�<1�eD�GcX��%I0M)x�����A�<1((�~�S蛲�Z���&C�<9�$DOǠ*5aγ+�~a�''{�<鐏ߗa5nА��)�H��g��J�<Y�H�|,Lp$`�{�2�Q��\n�<u̖�3yl��т��T�1�G�<!��DNl�i�R��\|�<Ac�2|C�E%�	�ڨIIwL�}�<a�i �E��r�]�	i�U��";T�����Ԟ�&�q0k%c�ˤ�u��I1,B�qO?� t�9�aH:�d('��
޶��P"O�q�H�;l֌@��lJ�Q��X �Q�\#B%3+BY��Ʉg<p9@�գh�Q���P��N��$!@ȁ��,��!A��"7�s�Ԋ0���u
�'�mq�)_�y���k�͇8<�J�+���_�u�����Խ��OvĔ�K	"����s��3�����'O������9���F�� "U,���4:��B����lӧ�����UDX�z�	u�D����p<qQj]'��'#Mi$iJ�7�f�h5��\=X�OީI�ㄨ/����
ϓg�Dj�˂D�i�ᇏ�z�'�����CO�S��c��r��h�������n���x�"�=n��7H@h<��	L�q�����Y.�( !�B�W̓�<,q�b��ؘx�k�*��IN���۴H!�Qr�dH�hݤd����D<���x����ϨEMv�"w���Y�����iO�:$�:t��/��I^��M�p+ҭ���rƯ'�xy:ed������}�qO���/VU\�!���C.���c_�����4 R��'"e:�ΈO���AM��~ (�Ofe)PfÛ鸧�	ڎ|9[p�S�RO��`�*�2Mӄ�9��ʄBoRT �'&j��� O�������'j��0D�P㡎 N����5
Qt*P��p�g}�O�fI@�ƅQ-r�8cC�Lp�˓	�R��!fB�D+"�\"��$�۸D�� �R��RJ�ϓN���kĨ-�)�'$��YS �
Z�4l�J�qM���Oa�b�U��D{��;�c����#�����p�O$�3R��,�0=����T�upR�Դ!�����O&g�yiP�x�B$�;�q��N�L3������#_Z���-a����$�Ԋ�Px�@\��` �H� �X���n��<��i� �(!Ҝ|��@��8�=�S$FFykD�$���KEI�7����-+��7���2��_�ZT�Q!��5�L�#�N�.��)�θ�!�����S�O�Z�"rQ�`p�8Q���-In"�
I��YҬ
]��t�eB�k�OZ�]�W�C�p��܂�m˝Bd{L���u%9��8Ǔ2B��H5��E�
��SM�K=�lx�dڋV���5GT<٨2��l(�g}BaLn.�J�	��80�$ՁH^���됯%^���ɯ$	N1���s�0��4g��X�G`���t�䓻�ē�Mki֑K�6��D��z}���5{�B�+_2\��a����L2�p��	�e�h�Do�(��DO"S�@��%l�|����!e��O�1Mo�\¦��(5!v�	A"Ц�~RF�7`9\�Y���	���c�4q �W���S�ȁ�g~�O��C��	e|�	f�}YK�;&����&!a�:yh��	+D�a�D�I:I�e�IOw�����I�y��h�Hp2�S��ɪ��};�옮�P 2�)L?s�c�\�{q(�'23��Qt*�7{ڀc�����N�P!��C�+�8L�h]����(�)�F�"a�:��t,Vu���1Ï#y[L�S��M�N��,��쎳9��%Թ&Uƈ���H�<���q�!|QX�3�N�����|0��38�@fF�)RK��H��'	�``r�Z1 �(1���`͚���B�,�%S��S�v�Tc�L�/>(��%�� x���eʐȂC���TmD���x�A� �J(u��'���O�BEƎ�X �$��r�E3!�X���0�%�M
xs��ڑE��m��o�>!p@ۂNў�tl���$�n�,�����$�.Y�h��<���ޑ~�|I2�"PH�2��Kƥ(���O�q�!ݝ@N���/_ *�>���Oil��1� ;�a~���!��!��;����U��;_s��A��0�F�5�>=8�[?%��Ϟ8����O.�X��"MT�A�hD�[N�p�C�'�*�hr旇A�:��raĹl��X�pe(Tk.H��v��2�E�=�P�5���+]�E��k�Q�2�[�|yaxboZ�kZ<@Ҧ�v ޟ]�6�Q>?�B����@>Z�YV+Z��yRJޡRm&i$ğ;��e0p��1��$Ȉ>tZ=�P@�
f�R�k$
Md�O2\4���]s���9����r�� �'(�Q�%���]�������a��lyע�']� �㵨���1�Jȗ��g�O�<�aᏠ����'ʨ2����I g�:��Ab�V� �Щe0mXQ	̖�p�ɕU=�� �SF؞hR�M�Z."�Q��׿kNɻG�;�ش����F�t�f�~��yBYw6��t��9bJ�`����7���+�'�h�؀��B!8e �.�*�Y��'ٸm
DB��b`��Z�f���;ҧ'*Q(���Q�H��e�e��N���bÂH�� �?-\���O� )3$�رd�(3͠s�j���D��f)QԊܓL���'�N�:��}2�?8�Z�!V  2sh+2oG���kp��+B�<y��4!�,`��TH����7���� �x�}0AK�}ў�)AB�15H�� ��u�\��˃�'�� 4ږ#�"�"��'׽�<+QL�cH<9��� _>}B�x�2}�l���E�%.�����d�v��E�U(U#�;��Q�R��c���=�!M<+L���'�b�[քD؞$����AH�iZ�iC�E�� ".yX�h�����_�V*��'Dh��.[~�P� � �
H�������w|�����"�Rap�"�ZuH#J/D�܊F N4.϶I�Ն��i���Õċ�n�dۢ�[Xf���/��^O��҆��6��	>����S>Y�x ��� M՞�y��I��hO�%�ďV��R�$�7#l��BbX�L�z�h��.]HQ�&M0YI"�#҃Zd�<ɂ%D�k�0�'ʰ#}���rb昪� �r&>��CG&]��D){\%a��T2`@�5 �-qh�`�q%1��$�'탕{���m=Q���������@ݽn��j�'˴@�$��O�y�
�7 ��2���K��AȔa_71��T���΃��Ƀ?meZU��� Y�u���bMV�����-\U�T0� NIa~B��&�	+R�ɼ4�6�1�&��Y�����C������A"lY��05�pɽ6�4�I�h�OE0u�4gX-~����8v����$�Mw����MQ0o7���Pg�~�s�Y&K�ɠA�Y+co"�S�+�?e�� $Ҕ��O?���|Ν�����,�R��1��-<��Č/��q9�"�Xd�Q�#%��� C�!�, �%ʀ�A�v%h����}9��чnp��$�E�i�e�fm���R��-*�epA��4cCg���fA�L|Γ)n٪©�EBy��G��Yeq�3b�a*�m"�O@q��g-d�`�r�|r�`���+?F���R�Ȇ�M����n�?9�lN�3�^�{�	_\������_�r":}�
�֙��G�OF|�v`�*u�d���ʲ��4���{�(j `�8�8�1���p>��D�*޽�$iT�%��񃦚�'�@=	�GC�t�2M
��I"b��?�� ���Hs��!�n'N��4�b"Oj�YD�� �`2�
�R �!�'vD�H���$7��P.� Hz�yd�����Â�V'Ҝ��[?��\�ȓ$�p�F)�2W�tm���ָ�v�4j��)[�ֵ�~�S!̗a���I0h@\7���y�@��ƚ64�8�F��q�S�'j��D�䌛�Tͮ@+���h���"bJ����Q��J5q�T����,�0>��3Ŏ��F���f��L ,e�`#�kV�p�Np��ƙ�?a�p�W�.�� �O�t}[�dY�@�A��5=t��Rߓ(Dq�3��>����� :���0H�I��f����j�ቢv����*�,f20���j�O��X!`��.���c�@G�օ���;8�%���ɀx*��@a�Լ5���g�M	#� t��b��N�� ~�ؐ �^>�Gx%U������o��Xs GWF	j��.�Ic�O�a@T�U�n �3�ϳ?�@9SGH�R�\X�@8B��(ӓH�s8�P����3A"yҢ�V�Dn��d��OL�	c��&��8�H�C��On�XT��9���&8���t�M��|CH3]!a|��C��l���jJ:f�{5��,&�؉��E� �G�`�!g�����#-�^H��yB��$�>;V�ٟ?����S@0X��MC�b$�0�>�wt�n��`	�Q�7��S}�y��#��LhuO���%��7U
�0Ђ��oe,��׭���ft[�-� (@��Ų'������k<���I/%��IF���.���o�$$��g�=@�]�Df�6&C�	�s����Ce��XX�MJF�E�0|�,���Q8�ЬKv�^�O���5�ѕ�jQ�Ю�0V:l0
�'� u�W�߈r���GL���|�a����� qG�<��'�gy2��[x�{����ju!jq��y��J�b��y0M3:��P�\�h���	��O�\#�#lO��A!�ԱX�z��Ƭ�<���'$�)��gξ!����i-ҽ:P���
�L��b�.*�����'���P�b�{���җ��,/�ő�{B(֖��T�GDċ��>]IGh�/Ip:��%Dq|��w�-D���$A� D�1r�K�8�pH���N�Q@ Z��l���DɩIG�M�r�H�i@:03�P��!������j]:�Q:ǧ�6b��
)!�����'3�X���޳f���뀈Þc���b�'�P�aG%G%3�Se�!	]М��'��A�A�j�5�Tm�rؖI#�'w� ��s`�Sd��#cj�'l�@�0�����A��0E#
�'�(FY%G��=+2�
�|���Q
�'�`�I���}M`�J�M�z�1)&D�� b`��ȉ(p�V����ߎ�h42�"O �����n�qo�H��y`@"O�DB�fǧ�T�)�.WA�Xis"O ���U��Jݓ��
~DI�"O^��:��лC�08���"ONb���10�r��5n���ab"O��y��!g�nd����z�
q"O<�)��X��L�W�G"r����"OT��g>#1&�{W�Fd�1�"O�I��nE�i�������=�A`�"O���@�W����3\���Qs"O��Bc�1n��0��
x�2�"Op�d�Y'/�p��N�*>�����"Od+��c#ߡCϨ�q�j]!�](4�`��pF��2� =���W]!��'Q�ȣkC-{��H�"D�!��M�,
|| ��O>�e���7�!�d��-�d�$HԛB!b�צX��!���^CJ��u+U4
�-�t�.Q�!�P7JD������a�ٌ^�!�d�r�I1�ح&���r�� 0)�!�$S�6ư��P�
(`��ip!�ޡ!�ټE~�!���	~ö��EG�`]!�䙺HwB�;%�M��ơ҈&k'!�dтV�b<h'$6y���� k!��ޯ��Yb��%s�M�K\�	�!��
.C�B�k�(��01B2�D9!��X�&-��!�������,�=?.!�D�>>��xᤈ$~����+P�t
!��>�k��X�S$ԂT̗�!�$	�"��\y`��s0J-���8$!���A�pH+1·$)�d	Q�X �!�M�0,���EnA�5a��MV�!�$��F$�I@Jj��CVfLz�!�Ā7�^E8F�|i�1��Le!�$R�#t��C�"����ac���q�!��JqZ����:�%�M#�!�DN��J��s��+s�f�s�,$~p!�䃂8���0r�q��5iJ�`f!��}���s3k9D0��8ǊT�!���F����vK)>�rt��&�!�D��<��<a� O��0	�LBT�!��2I�yg�<5��yh d�.|�!�E�JO�Uh��� i�V�[�!�D�n�"pCp�6qdV��q�b�!�
8� ��.�C���'(d�!�DR>Mcp��dk@�[:2$��g*�!򤅘Q�dMHC�z��0�+Q=:{��������$͙�Fr�Y��	���A0-2���8u�1H�V�&�P��u�!S֭ـ8M���ʀ`�@���QP����v$�􂇸{�����\��D�R6�A��,�(��ȓ>�@R8 |%�T��Q�$q��cg�M�4��� ;�)� CR���Ɇ�锡`�H�"�4W�[|X��"J�Z`A�0+%�R�i[+����ȓYi� �	@��ԎL�<�,��ȓ^Ԑ횇�͠�5��@G7Ype���ԝ�VjR��qk�!E�"nЅ�U����,R:x�2�ô�Ɔ"Q�M��4��-�U!�$.EV��O(����pI�F�Ͼ�(A�(I-���ȓ��Pa&)�$Y�!䄊*e�FH��S�? �E�*���i��էP���{�"O�r�b^�I���s���=T�4�;�"O���CS�����e��}�n�q�"O@�7؆���j�P�jhAz4O�e�1�L-Ƹ�������A��zy���V>P::!"Od;�V�+�6%�&-S*A����^������5N�T ��ɓ85B����� �f���E
���2 0@rƨk�zM*4�1L-��H�$���'��9�"���=��m� 7H�0��D��h�EA���O�4�Z�n7b���#"ƓyֈD��'( ��MM�8�X��,]Pn�xشbж�I�ǖ�?g�ӧ����dۆV�����2��YQ���y"$��Y�,�Z��A5a��s����d�#U�5[���
��<1VnG9�����A,�
�r�vX�xE�U<j���Ṅ29����E^jtEԇ�!Z�񄔚b�<��.o��c�*L�,���l!5
L2kv���	3t��Q����A���rS�L�V�!�$�)��xP/S5D��R�O�wɛF�W �U����@��s� ��P$�?�>��HɀG�,8D"O⍚7�T��͊�g^�V�t��W���l�&;�����'�f��᫁8cS@(��L��!7�H�	�Adp���V�u8�1Q��]�A�>-H� %:L`PQ3�>$���a!�$������ɝ,+�,����f�Yb�x�ɏl�q"�S�)��:��ɘ��A�tT,__^��DE�3�ɫPi�(����^���[����R Iy7�d�+����{�����(�蔊��Ȉu�~ŠQ�"M$����1C �G�B8���I<jZ���$E�X��R Q�!�$�dr<��@R�B��Ö́"⦩;!�GsyB�?1���}&�,�$h�!1mL4�T*�vz��V"9�`:D� �R�3��X4��� ���ZȄ�h��9V\�M��ɠ�H��� �
	8��A�Mƒ��$T�\�@@J�`�`2�
_J�
3$�	G�i�̈́H�q�' I��	T�S�O<�Rv�	Ad̬�PP�=�
��I��q���.w�%�u�G�O��{�C����&�
7Rj�qN<4�k����p��1j��F�()\�z@(��-�LQ�꟢d�剡*T���E��I?�.�N�[���왁BW�r4�9�#��� y��>�O�Qp@�Q�f�hA�ߏl5�[���� �D �.�W�O6m95Dxɧ�[@��I�
��t��)��q�p�c��ҷx4�r7�'�p�@�ě$m�ld�.0�-�"и�aFؘQRF��QK° ��9��(l��)U���&�	oR� s,�hⓅy������V�V3c�FZ �OT#C��X"��A�IU)�10nx��!ł��M�� �#z��H�<�4���
�5��y���A�  b2���'f� C~���q�B�6%�(O�	CR'����i�4d��<�kH~���<Ĉxp�\ g*�l5��Bm����ʂ��-H��/�O<H�b�P,C,����H%iN��K�&+��"AdB�9M�L�FĞ� �<@���.I8��	�oF��wZ�Ċv	XL�L�����wxQ�0_�����֗����W%��R_,Mx	�*cvUA��Z�z_tm)Ӈa����'�N��ҋ�(-��O�~]�W�_	2�aфG�R݆����|/Ќ$��+pP]K�fK��u��q� �@�E�C�. �d��9� �O�%��'��$>c��Xrc�6ˠ4(�A�\�9���<�F�P�
8�K�g՘#��0�-��Ij��g�I�`�u���y��`��P |���AQMV_��T�5�.J�@���j��r�h��GP]y\���O�3���4���O�D�Ҡ���p��~
��#�� %Ǻ9Y���ob���	{���Գ,�)IP�Q�dQ��F<"�B)۱Xr�X�)kqO.�N|rD���Ua0��+!�*���:O<�S%�=@����D��.n��lZ�%�,�y���8A2�OB�6��C�8R9���s�8<9/�w�0�'��yhRD޼"�Q2���E�>����1H����&s�ԉs�O4D����˜�N�t$�m�s�P���>��u���#��L��~R	O (���C�D�t&��q�g��y�)U1\&�'\�m��u�7��?ё���*}�]�&�<lO"��B��0.;&����but ��'�x9j��*W*�lZ�z�1#��;h�6��P �m|�B䉈}X6	1� )��ƯڔpBV�P�B����x"�S�Z�l35b����qb��C�)� N	q�V'.�~�QqJ�7{�.5VȔ�"ba�"�'��s��c&a��<��E(ϒ�G�\ ���$D�x��.��$�ӏ�7j"�ٶ��p��dI���q#.<O��z�EM�$+4hg������'j8���~�8��Hҵ`���L�G[��O���R�1&�&�2W�F�V�ЈO����d�#�(�"��Dc^0n���80�ذ
���� ����@c�.��
ۓn�p�v���*"���q	|�i�6O�A��eȔ�x	<}J|�@�$m��z���3��݈�Qg4�R��nB!�� �@p�`���?`����[5��*|����-a�` �e�N�~�'�f� ���GE�	?k����2ֈ���ٌnKV��:���	�Jv��)S�+Լ��1�ȜU��IA�>y���O��:�m�Ê�
��� ��AE��:Y��
��3Q"q�(p��aǬ(�|�I�J�O��r��ObQFkN1Pxh�ӓ�xA�e��K���@DHŠ�`a̓[C䌂ꋏG�Pҧ����~��E���\RV����a1�� �L `�L�0"Oj��+�l��)N�\�M�%�>yӏ��3 �t�p�ί_Nf���B#}Q?Ys�MT�W=dl(�E	8������"D� �f�/�����%A:�,B���zd�؂���J�Zҧ���ǺY��$9���P�uP�.
<�y�B� >��`��n��_>�p����~bFt���aǓf��K��=~Ozh3� ��	��t�R�;�O�����c��������Q���YE��'��EQ!m�<�3o�R�P8�m��X��I1P�/<�ri;�'�21����T�'��P�x����3)�
�J! W[>'�a~�m��H�@�+w��O��\X����H���0�"J�C��E���n\<��I�|�$��q��.45.!�"���w��=9����
�rB�+�I��H��F���to�W� ��F^D8�(3����y��
+��h8r�^2E�
��ף��?�Bʊ�&=�c�y5>Pq!K
�h�����Z7��!��p��M ��%D���vB��}�,ъ� �6d@��DF�:n+�P�G�R,K�X#�D�@a:�'�O����ݳ6m��X�;x~l�U�'|fѕ� (?�v\R!$ěh,�D����U�
�q>*�(�b�7&�S�aKH��Wȇ�R:(��J�hG{����%�QL������ӆ/��	�_&lP����b+^��h���!����^(��<sD\����6h��l*��s��D5z��AӶ͑���>-�#a���RR��n>�S"�Z�<q�g�V�X���W;]�XHkСtz�[U�U,a�v��5Hŵ�O����dMjzH���G!V" a O-�O� ��'i���8�XL "a���x���12 i�	E��p>����-hj���0�2U.�:Q�W�'ZВ�f�ϟ48s�ҮT�ӅJ�F9Ж��A7�I�gΎ�HvB�	���04
�uj�� ^5��{��A
�}E�d��<f��m�F�p�j� 7��
�y2 ?�0�����?e��!� �I��a�Sk
���>�p�d�`�W�NBt@��i�b�∇�q��l�����UaA�U��	g̎��>5ـk�a{r$R�>8$��'Ĥ}r�r��W��p=q��Y�HD�զא�M�VCD��	��s'F0��
f�<I -B��f��
f�Yx��N�2�"��2�F�Fr}����<"����J1sa���_r�!�$D=EY$�"���(�ҳ���V�+T��-G��'ft@F�,O$,��
.rb Iu�3'���#"O`���mZ�A���VlW�v��	�3�)޲U{�/�n�|��ɗG�|c�KY�,L8�XӅ[/l���dM5�\�v�$[7��U8-ƬXͦ�z�j��5wjB�	�[� ���ZNZ=�R��w�*�@9�@�@�Z E�W�O"T�si��{�������@��% �'�\�.4:��)�b��hP�5��j��^�xP�s�>a��>qB�}�H��CbO�x���E�m�<q�Ԁv�lD���7;�2�)C��x���.��}���)L�d�� �\�,�BL)���W�NC�IE7)�vk�i�*��㇨O~>C�ID��������T���i��G.(kC�)� ��JS�W)�PQK�Y�"O\yEC 2�<����@�[B"OZě�f��OT(NO�;��l(�"O�R����v�8�㵣��D�B��"O�x�@� M�B*����bD@��"O�� .�A	�!��{���!�*OlТ"�\<w��}Z���h�����'0�%�D�	G�D�04cBd! T2�'�DYp��
/F�d�+PȢ�)�'}p�;�o�6`#�|Cm�]���P�'������L�=i2�""�6�F9	�'�ɪ�"�YɄ�p,s�z��'|-X�
://�ѱ��Ĝ>cpez�'����I�5�����I��*S�4��'��1"A�,T
���1�G%]j�8�'X�)e�1����𭅇^_֝q�'hR�����<�`!��W�DM��'e����Cp�\�{�R�LU4��';t�j䫅�!�`�t�����'���9 e�K����ƛU8�'?�����شW�~p�UI!w�d;�'z8e��c��|��e��/;^t���'����e[�.H�e�SF�:ި	��'kJ��Q B�z��񭒄 ��,�'̒�4b�D�t����z��	�'K`m��Ϟ�V%��hG6"�<�'��q��� \�n���l�S����'�
��M&>��%���]�Ț
�'f#�ԧ&i8��"V�p����	�')<|+�#��b�@AL<$r"���7BB�*B��zO���F�9q[�X�ȓ,{��+��_�is��F�-m� ��bYJ���"Y7@Pj@ lG���ȓh��)	ʃo�ݓ��ttx}���̱�q�ͅE�IK�����ȓ]� �r��-~�d�w�Θ1V:���m�D�+Ui��.L���f�C�R��ȓk����eT�/ޖ�k� �4�:��ȓ!(ȂD��O�N�A�_#A�*���_���$�O�֬	�HR�(M��+:���'�0*���;eń����aN��B�7+7"���(L�?"n%�@J���ا�O��2�]7�v̛���c����'逼A�C�,-&ɧ��L���(u�)��
��r9�<)��>;����%�Pe9G'���X�((Ů���z\�S��-l�5 �R툜�O,܄ᓴxޢX#�"H#�0tzO�+\�DL���u��W�^��}rN|�K�)Hm&\�A)Y	t�j]T�A�	�t�hY	D�R��M0���M�K(�9[@��H�,;�f�.
�`�� ��@b F��6�tX���R
��W�G�R8ap��0�����p$xШ�œ6H�	 	{>�9�FM�^�����M�){��\���H#h� ���ݖ���M��<E�D�J��:U��
�$̞�)��
5�pq�좄B��OFT��Ӊ)3�HP��L6jR0�A�1j�Ƙ�"#τU��ʓ.Ū}�'G�ά�D���țg���7'ytΌZy2O�!~{ܘ S��4_?�1��@��%��y<0��#ƘO���OzdPG#&�)�SU(�i��m�r vă��Igw��o"����G'L'����T�:j�X)�^�!�d�<�PL�"A-�hKf�P��!���N�>����Z��0U'ݿ4l!�dޓu	VyfD+�4 pƟ�%h!��޺!����n C���P:R!���@���IaO�M0�����+8R!�D�653�M`�%�$~-p�`��~;!�$řu����o�� - p{�N+!�B�=C���n�|�������#"+!�� �`
)NM��M��H�%�Na�"Op9���U��}��[$`x��6"O.�3eAؗ>K�%Ju���zG�� "O��	؞����e�4n;�q"O$���Y
U��r�� ,��Yh�"O
�{��H���Q�M��V�"OH�r�/ '$��ɴi�6Y@�v"O�<锠� sPb=���o����"ON�c��$Sx�-�A"Q9���qa"O����Ċ�4��(Q O�y?���"Oz� %e�";��Ѳ�78 Q�"O�L�oa�̀i=�L#6b$\�!���0�6���H�(�y �]M�!�d��u��;$/A!F PD�<+�!�d��~�+��� 	����Dw@!�X�;Z墳��IPu��Ǚ�%!�D��Bܠ� �*�n��sl�A!�D Ft��kݐkB�A�&˂��!�d\�4\X2l�.`��3C�<s�!��+f��u��#�~�(��D�!�d^=Ƽ3f���B���#�^�/�!�dα��+���sâuq�I+�!�$��`z,����[�^��=Y!��)�!�����2+0�Ь��^�7S!�ďL͢iR����܁NI!�$�I��m,b���Ҩ�=	=!�Đ�k`P� �o�X�Ah�#M!�D�9(�����\�Xy��@X�M!��[�M "����\$4l�U�􅖒*1!�$G ��	��OȯBk��P�;$!�$ʷF\��*�K��#fqx��=!�d�Q�4c��.{Z�%afn�=$!��g�z�cq�E��|���͆�2!�D�4U�0yIUH=�H)�uc=r�!�d�0e�P���n�">�ҍ�hP;F�!��P�h�%F�G����eh\�Gq��$ʷW�茒����M�`O�6�y� N�?��$Ӈ�3D��!�ehO��yR��k<V4IRDǣ":�3u���y��B�,y+@�Ps
�P���!�g��VB�T���c�}!�d�1>�,���D�Y�� �Eˮ@!��Čt�I��	!�d���%�;!�䈐V���3IF�$|$��#Ε!�P�s�l��gY�*f9K ��7!�$�:���q�N�~��r�-�K�!�
K�MB�FR3q�N)�e,xd!��	cܸ�S`�2Z��(ru�οc!�DY.��x*c@�5!� �Y�,C0)K!��B<F%���"�ʙ�U���JE!�\�,��p��"9��4C���:y5!��ư�U��M_��D��a���Py 48"0hQ�LZ�~m`�T�yҨ�/u��I���OFx����yboD�?�F���H�&=�v�;PI��y"�E�I�l���"G:�LQ�����y2�H����Z5�?9���؅ �3�yb9
�8�)&DӬHL�a�C���y��ήW��M3� A�<��mM>�y�ўD�P�Ь45f<a1�]��y+0"���$�	�3mt9���8�y�'�n�!�9_+l耵�8�y$ڎ�xp:*
M� �ڤN��yb�PV?��kD� C�ڠ��	��y
� �q�&�8,T-qpl� R{����"O8q2�I�Z{�l��n��ɫ�"O`�hI��@�,�2艛w�"��"O��Rq��^
�t��D�Kk (`�"O�0�fd|(�)�I̢F���"On�Cщ�.���r�=fy�h�"O~H��h��b5$߄[e��i�"On�e ��I\�-��(	�,�F"O��r�%-RT�!��~D�q҄"O~�2�f_�?A����G҈Z�7"O.d�Ή'�\I�p�ϦN�A �"O�i����-��"�H��)LH��e"Ol-aw�P6_	�Yh�F *~Sr]��"O" �V�Z�p��T2 &9`�"On��삛t�����D�MuLMBq"O�`)𪅬]Q���/��L_�A "OT�X���Ze8�W�@�w�XX�"Oa!�gG�L�@9�� Y�(!�"O���*ʈr��C��L*�F��p"O�q������Ү����d"O�Y���n9jí�`Y�"O��J�C�*(��!�":ڎ��E"O`����R� ��p/ɐH�&��"O
��2��F¢�U��;�Ҕ�f"O�L*�
��g0��M�M���"O�����#c����c��b�5"O�� R	���&0����!����"O��:r�;p���1Q왉z�d�Q�"O���0�Ɠ.v��I�#��;U"O��3g�?�VA:"��.3����4"O\�UC��5-��cV�Z�ƨ�"O�S�✎U��P�مo�0��"OX)��'�86j0�"���9�d��"O���/])S���P�@��r$��"O�Hr�(�@����m�?KL�!"Ozq[6n���@Aw*��)и�!"OZV�Y�Z�� �B����"O:� ǋȡQR�Y ��X��"O��q��J�O0�@y�d���Y<�yR�v� �Td��{�Vy�5���y�F�3<��`ȎF������yB�u9���s��8�ir�g�0�y����?�M�͖4�ʩ 4G���y2"��YĒ�:�(O&)����T�ט�y�˥p��CB����~u�f`�9�y2��[��D��+ O��y��;�ybH��Ux&�S��n�x4���y�L���j�����0����(��yR'��Q�]ѣ�đ~yp1��gא�yb�Q"7��"鎤	�
Qx3����y���g��9�!"H .���Ac�y�"%>��q���1ɒpɡ�� �y2G�4;�%�dK݌(��k�:�y"@O=$<*ŋ%L�4�e,���yr�6	<��	���+0�8�#��;�yrMՈ,�u]/#��X-B9�y"%L�yv���Ch_�d٤͟�y��L7o8R`�!Cбe�z�4k���y,�N�|� ��>e�x�yC.�yr���c������g�I�C/\��yb�ǡN�rM�4'�R���5��(�y��N�����FFE��i�d���y�M@�
$	��d��Cv�E�T6�yR��(Xp��]*?h����+�y
� �˃*�&�e��(Q	Y��h "O�}�B��<{Ҫ�*�'	7�p�Z5"O"��o�1~���� HkʬC"O�]��ݝ\�"M{S�R�t]�� "Ot����j?xM�ʕ.3A|Q��"O��&j�"K��©[�K9�x��"O&EH��P?S��4H�B�&�^]�W"O,��m�5Pr"�
3AQ�\�F`!6"O�$�ƩsӠ��Ǡħ]f��	'"O|��T/3FƁ�C@�1&c���"O�a��ͧA	�ȶ&E����"Oj���H�(}�b��BRR�؂�"O����j6>z����Q.�v886"OĥE�9[����Z������"OB�!P�C�\�t̓����"�[g"O��
7�U�@⮨bP�L;l� +�"O9���ݳO����1�߄im,�u"O�����qڸr��
0l`�@�"O���`�ۚo^��J-ɛ �H���"O�|{��/����Vk��J���[V"O����僮�pA+�lh ��"O� ��菈GԸ��dʁ��F3�"O96�7RN�Z�	�E��|��"OFD�s�ιXݘ����H6�dP�"O�A�(��Jg|�JB��'늬{d"O5��	`����%���p`S�"O6ͺ�O73����l�}�B�X�"O$t��#�* �Q���!w���C"O&) �al@b G)u�P$z�"Ob��$,��N��Z�nS�\�D-t"Od�ć$!b��R�K4���"OL�����,M�"-
�h����"Op���Jߘ\7�k��ɴYZ@��"O@5Y�)�b�B [��*�j��"O��ʂ�ޞ[��pU�y�`:B"O�s�'�'��� �����@�"O<��t�\�0��\˕+L�
� �@�"Oj\*Wo��r��#@�?H�"O�5���`v>������`M���&"Oؘ��mǱS�$i�OD	Fn�v"O��ҮJ�2(5�.�)-"�Xe"O�ԑ��RA�JPx$��.��&"Ojar���q"C"��`0��b�"Ou�sF%���n�"5C��p"O��K���PzQ[Ƿ�N<x�
h�<y��.b�Z�y�,۶���S#�c�<R�O$R@DЀaM�ܰK���K�<��Ɔ�R��9:r�K�^�C�.�l�<��`��B>Y���M�6iTh�I�i�<䉖<@X�k�oPL�H�8��e�<�΅;_>&){筛�_x�`�K�d�<����E�ҐH�̈́89jUh6�
Y�<��S�&?�T@R.U����Cn�S�<	I��H��0! P�4�����e�<�-�0٣����ܳ���J�<�-�5>'0<���5xV���,m�<�B�]C���b-E�l�|ԓbC�<�D���ؚ�^V���HW�<1! �u$f����I&XB�#r��U�<���V$ @  �P   b
  I  �  c   '  �.  .5  q;  �A  H  MN  �T  �Z  4a  xg  �m  �s  ?z  @�   `� u�	����Zv)C�'ll\�0"Ez+⟈m�	�|��:F���DA$������%\�U�b(\�f��d	E/P8cꔐ�gH3]��%Ib~xݮ;�p|��'q��Yh��A�Ժ@����R��a��3|-�M	S2�@�S�X8?SjtS��ղ"�0��� �-����$H�z۴�Gc��Up@�KBT�R�B�K��Ԓ[�H}��[K�t���+T�в�4T}���?���?Y��'@&��k
�"��
�jvy������I�MS�I�����O��0�*韆���O�]#��Im��iB$����Z$�S�O\���Oz���O,���OT����'��Da�hq�Vc\]�i���(x��>�O��� !R���XV9�℀2,�듨O��.�|�Xї?Q"@�2*cv��'��1� a��O�$�Ob���O��$�O*�İ|b�wG��hǩӧ��d��C���R�E���Ks�d�l��M�����v���@6G(:�����"�^}c.¯;v,qy��W?�\�Fz���w���}��E��H�"�KG�+(�ǅR5#T�9J�B4hܮ}xS�B2�MkD�i�V7����)��U�m%�B�T��9�%��&� �h����o�"�l�UG���!� y�1��U	]��d
	Q��8�4J<��eb�pUÎ�v� ��w�ߗvO`����9�hT��
�v�`m�MC��i|���:s��{e%^���iG�
���^:��jAAU�bY`a+G [|b�᥅���X7-��q��4v����FX���Q`Y9@j,���K��x���d�F6tH�P��#��&��x�B�`�$T�	m�D�1E����$�GP^P��#��4J}h�GLn���5���<�Ia� ��ش��)l���\����j��g����'���ߟ���?��@�_�H�<`�@%�lZ/:��K���G�y��N8 x�ቒ|�`�s�4���R���hH7*Q!8�zi��o�5)���[d/2O�Iv�'�l�<1�%�h���!f^
��'��ߟ������?�|��'��|�a!��&� ��7��6�y�N��6�-WdJP��j
d�����h_���7�*�	I���?Y��3S�����c!���	�.D��-[�'v^���W(k�}�`߫mJ� ��'o���a �f�h�eˁs`���
�'p��[�[�}���B�MffX�
�'b~�����0'��9;�fC[]��b�'�ƈ��aH�g� -��N�FiZ@���3�x�Dx��	S�|⅂���(��/ m�C�	�/��=zgU!2�5	���	+@C�	*8uBZB�`����7kGtZB�I�Nz`iiq̓�ކ�S�̆6gLJB��2l�zP��/;An��Ɂ�&GlB��'l
fQ��+!9�K�O��(���{���	1f|�����"�c7n�cNB�I�T+�)2�卜��������C�I�w�hB���+��PӁ��-�C�"C4B��7�)��tk�-ʏ>߲C�	�Hq�a�����x�/[�����Cg�Xm������w��XaCjZ>d���eʟpC���џ��4)P˟�����\����\��mm��	�D���w�0�Ӈg+F��pah��.7�}�	�����ׂO8p��Ȃ��Nv�C!gS>h %�ƒ$�>�#&�M��I��O��������  MR�	����4b�{�AӼ�Vp�'6���ӼqO�aC��/j�E��-\7l-6b�@�'�>�s޴*T����JA�	����'iЃR)@���i��'�R�!��^�O:��k!c┡A~���눶c]:��� !D���#�w%�<�bF���d�f $D�X����A��Ȗ�C62��S�E4D�L��ė6:�Ԩ�d@/??4B3�0D�ȺR�S�:\���&w���#�2D�X2�A�9v�1《�>��a����'��{g��?�������}y"��|<�H{� 
�x0���$D�����4�e���lZ*6�H�j�� *�	�OҒ��$��2��Lp���7U�QZ���z�td"�o�[��`�6�n�0���Otl�uL�,����`Ԛb�ɠ�kg�h��'����Ș�?q��?!WA��%�Lɑ�[�o\z�)p����<�U��׾���87�	;Ѥ��T�#��	��M�A�i�ɧ��O����D಴a]� �.=kaN�9(����O��������uy��d�$����R*w��D�s-R1 �
9�򁁇9�.Q1��B�����K����	�b\&Y����*6�V��V�M�	E
��g�LuGv���l�Zb4P��Å0ej}�4�˻^x��b�,��X
��'��R�'��)gJٰe�`��\��0	�'̚!�%��}y��٬ifh�M>Q�i
�Z��aJވ��' UQ3A��l;@��B
�5]����Iqy��'���'��l�S�V `6k�%Z�N�� 8h�K��^������!�z<YU�'�R$3$�.p3>(��e��u{��A�G�Te"r�C:����5MC��0<ї*ٟ�	b~����e���b�%�(\Z�*�ƒ��䓩0>)!�C�{�&��E�� H��S������x�6yPUm��P���hdjC�&'���Ay�!���6�%���|�����쨖�*�n=k���&>Ċ���?!R�.R0����G>*�4H������K�aI,|����(�]�#���KFO�Uq�,�G�L W@�D�d�H(5��`b�⏺$�d�A&�z9�'/��K��?Y��Ik��@�կ{>|�ɕ��A*��r�*D�H�DΜ�xǤ��` Mgu��q�,����>�A��̱]����'LA�b1���ڦ���Ɵ\��>2� ���c۟��I����IѼ�#�9$M��� �PwZ����XN̓T{�!��I�-gD����J��lɑ'^C&b�p�RD?LO ��3*B<���Y �Ź?�ɶ�2�$Ÿ?����V#[Jh 2��,6py2�mN�DR!�ğlb��D�,��X �&AY�ɯ�HO�:�Źu�R���mHl�t�a��.ĤL����������Py���4ЪP��5����PH�z�B� *�pqAR�^�
�(&�� Jaz,7E��$*�H9oV�$�B/_�u�` ��N��a�t����	�0=y�ǜ�L�|u��ݐN�@5b��ܴ/����I��M�*O���O|�d�O��:�Gؤ[������"��b�CH�C�	V�����	�
u-�(U+M&V���O1oڟX�'OZh�Ӥ{���$�O ���,ᤈ��џAF� �B��O��D�e*���O
���<���P�f�C≹b���iG�֠c1�x���`]bŇ��+t�̝�3�U���z�R,m<"<��ͨ)U01��&?�Q�)O�!hL��c	�qO�E��'�R �<ѡo��pH�d�V����H֟D��ן�?E�t�� 8 �z�G�\�X�;��T�?��!���,I�t!�D��Ē
~�bEZ0y�6M�O��d��$7�L�'R�'|�䂝y��M�4D�@�
]ƈ��A2�B�' p��À�
���O�|����x&r"�&�r�2�����^�|T��fC�:��Hzw�u/����\�f5d���Og�����
�S�$)�P%�/ȦU��O�MR��'F�7��٦i��k�O>֝�3�8�5!��!B��J>����0=�L7S��Q���:J�MQ�L�W�'#�"=)V(ήD�,�哞5FY�P<P���B�����(�B��O��d�O��D�LI��4�V��(��r��5���񧉁�P�1�܊7 c>c�hP���Z�3�^t�r1�/U��zm��9��
t�Lc>c����\�T_�<�O�f�� ��O��I� ��䟘G{R�Z6Op>�p���r|v���C)�!�J9Yr���T�rp�z䊑$c��ɉ�HO��my2����T�u�]�#R��*6���Ւ��E���ԟ�	iy��DKȭ,�`��O?��ka'!����Ǉ�ZP����%G����M�`9��c4�X �$P+F��
3�P��d�$V,D����O�b����c�����`d��J\�@QM3 <��'uў�Exª½k��0"0}�=8G�_��y��7kd^Dqw�
�q�h��!	�����X�A�l��')b��k�!Q#0�<�f��~�����I%��3��DW(�5ƌK_$��RQ%	� p٫�ē�BI�ȓ{;���G%��_��{��҆R�8��ȓ[E�-�A#_�U6|��a�L����ȓH�"c��-��2���2c�I2q��~�ŏ��&:Fp�AI�+5J �S`�r�<�Vn/`��B!�;T�1q�U�<yf"^�@�>���ՠ�H��v��y�<!&aη"��Y+��N�k(~� �hLA�<������6����� <EԄ� -v�<y��
w)6M�BL\y{�y�*���\�`�,�S�O(���r���3�O��L�@�"O~$�5,�;;d5��ÛN.��Ҧ"O(]���9�~���ˏ�S#��1"OR5J�c�2{.EKf� b�4�b"O����J��LX��u�U<A�ޅ�T"O�L#�,J5Y�0&��"�f�Y�X����/'�O�����Z�!WI�|��Ru"O� R�"��͘Y�DTq��H�!�`��"O�$��J��:�^eh���\k<���"Opd�V�0h��)R��VI��"O�y{�h�)^�PD�Se�
���D�'An�R�'e�1� E4TV��2�K?U��5{�'�ҝC�dZ(�`T��/�S�rd�':����F�*�6�hE�ƊJ;n��
�'n����L-?�丢�C2J5Z	
�'|�t"6�*�>q+��-ELri
�'S�@@C�9Pt9P7%��c��d+]�Q?�#%��B����3�$9 �� *�!�d�$���!�o���r�I*�=�!�D�$,q�'�B�e�\ɠ6h�	J�!�dKb�=�Rˉ�>���ؒ&���!�d�5]��� *�U����̉)(�!�d��;ؠ�BE'@ZxqR����m��nҥ�O?Q �F,*���Cm@,h'*`��&�i�<y��Yf�4��UȄ+l�PxFf�<�D
�0T)�7�Ƒ���f�_�<��+��:l"�p��4�	��-�s�<хKT�Hq�l����'�m�e�n�<4G�6 �N���ʅ0�n�*r�Ty�		��p>9���)	r���R�x���ɱ��{�<閃�=����e�ρYW4����o�<�O�j��K֧� �
2��`�<ѧN�r5$�I� V�.CR\��QV�<i�F�k����ރc��h�uNx��#�뷟���
.��HA.��-:JDB�,#D�,�dJ�	�F%a�Q�pj@Kю D�@�.,�TP� ��#�0��1D����%V�9�M(��ēG���H',D��c�ŋ/�)PIC�H�Ѱ#)D����BQ�e�FA)���!�R�QF�%�h^�XG����()��H�B�:t率�y��6o38�����I��m�(U��y"�WP��=�Qf
CgF0c�DƤ�yO	#X~��#���p`X@cS/�y�*�* �r��2iq�b���y�&M]�av/űT�&Q@b���?)#�o����4i�A�F�-�I#��� 9��9��4D�xC����������s�z�3�,6D�T(���7(�t�i�جQ�g3D��B�ց��p��K
u6�Qq&i1D� 8c@K�x���eF>@ lI)�;D��;/�H�Xqr�Ŭ.Q���<��*b8�\�jM5m#�,a䫖� 1����3D�ȣ�Yd�\�f�?�:@k<D�`q���w�V=8�� &!��=�-D��XlR�J� ��!IZ
^ �22�)D�;E�&+�5�..b�0��!)�O(�	�Oĵ�ކVaΈ�7��2du�	d"O�ѐ�N��(:���Uc��k�"Ozl#r���h��f2b��b"O�����+�"C�B�:y\���"OBa��瘉"i�mؗ 5>|�p"OfZ��9|�8`zUA�v(��
��f}h�~:��[O����х'�$�X׎Dt�<ɒ�
p�p1�!O+U���KMX�<1�F�P��� ����Q�*�R�<� �bcX�0]%(��a2�Y�<�"�V�-��4�T�� K���vK Y�<�I�bCte��́�e�xyDA	؟����(�S�OH:�[4�]�	NU�pF0�
i�#"OZxY��S΀ R�ʤ9�J�["O� (գDIOQ*�$Y��\�`�<P!�"O$���虅)[�D@�g��2��"O�Hq6�Nحх發m��X�G"O:�j�D��t=�����0� %R����=�OXؠ�њ:�
�A��^Q�U
V"O(��ӅǯZ�z��
�Q��� "OV
Rn�d�ހ㑞Z�D�[�"O��cňș.���Ɂ R���M �"ODm:�iޓi��9'!�4!�J�˖�'t�0�'U4TZ5�CI�����ߧAX�-B�'���J�EJs$��MR�"F���'�F,郺J2	�G���J�)�'�hh�Ϟ6mb�����X��ҥ��'��&����R�˂
{�d��'��|�$H��q�F5ˆ����ߜR�Q?a�#FU	C����CbY<��5�=D�P���@�^z��E/& D"�X��(D�psC�G�V^��� �e�ţ�$D�81�KW~�<HKqe^1e����'7D�S��+6�z�� ����94H)D�0�� +<���SD����R���O�L9�)�Xta��n��K�"�q`�k�!9�'��⁬��h3�]Ao�iʙQ�'�T�vH�]�u�/
�)�=S�'�~B�8���#fP8yK�'���ke��l��|(��T�u	�A��'b&`�3Ǩ|��x��j��,O���'А�ꄌ��J䚔�p-�v� �'z�k��e�)JWh�)(
P���'�(���(k�D������5y��)�'��!j��8-?<U�5��F��'��ʓ��$tb�)! kO�R���mh�A��<�M�!R<6�ɣ0.��n��ȓy��!d�1�����D�<k�A��<�D��D�J�造%�"�*�ȓ"�j �r�A<d�d��"NxV⁅ȓ/?�0J�ś+� e�U�d!��KeNdpSBP:	X�=�A
VPp� E{r+�&쨟�t�L�*� \��� ]D<���"Or=(���g��|�A��3�0 "O��aa�F>��p���0&�=ɱ"OH呰lW�a��m@���-"�@��"O�h���%q�"]�s/RaV!�dA'v�=�4�L2���FǑI-2��O?1P�J�	`�Ձ%�?��C&l�<��g*Q`�yԤ7�x[R�]�<�P!_)`��!,�6@�n���k�U�<��Øe�򐻴��43�BY�4�j�<��H�S�H�C�14J�%�b
Mg�<��/֥)�a"�̰g��L�Q_y�kV��p>1@&J%��xÐl�O�z�ek�r�<YG%ë��H� ��*t�B̠�Gn�<�6�
;3�����  9DDYr�^�<)c�����үC�I�δP�*U�<����67�ȥ�CK�0dz��P��{x�$8�H����1�)Z�(�b��׭x��5�3�;D��16㔿\��Q���
�`�%��"8D� ��蛅F^̤���?����6D�hp!�9Y� 0֬��s��(gm6D���ŀ{E �R� ���'a3D�|#��XI<��y w�|���	>ړ �F�Tn�_���P�΀�f%p���y�e]<y�O��f�����y��\�Z�Z\0 �S+da*�1�K�-�y
� � A�Τ|t��Q�3��!"O�$q7�K�?����-Y�h`��"O�:�I�/Z.\���|����'a�Y���Bl>!` O���l �-�j]��'i �31cA�1���BSH�8;�XM��'gf=��$Q�3Jl�	G�-B����'.�����^������J=7p�hx�' ���6���H�y���.���c�'�0Ep�ჶs|���/��P���.O0�W�'�&�Jʕ5�M�1!�%?����
�'^�Hk�Ds�&�����7�J�i
�'�b��7K�X3��Z�!�'�E�	�'�0����  ��`�i?6�V�	�'�>���.����II�x'�x��I�f0�;V�ժR����E��v�܌��R�t��#L�5����G�dX�ō4D���Qo�)������IȢ!��-D�Ti��];5Dք
��G��8��t�,D���j߰�PQ.�\l�1�)D���Sdp݌�+r�í�@�&�e��F�ģ��bn��	�ND�
�4�80��"�y��O��T����~	�,��y��̃ :�2'���h|	�sB_<�yb*�$O�&2�dS�]�����C���y2O�e�!��P8�|cscڞ�y2�Bf��,P�)�{�b���֍�?�f}�����m+tT�U4��W��DnUX�L5D�(��r|�{��և ��`�3D�ȡ ���aW,������3D��)��U����0m�o�TZ�1D�41"�[�.�@�/ӵM4U:�)34��؃犡"!��z��J{���`hֈ=~Z�)��O(�	c������v?Y�O����JOK �� A�a��`�`+��(��ȓX���r�� hl���0�@؇�ZX2]�V�:Z��{�A
Y1��ȓ#^`�B̕�a����D蚌.� ц�Y�l5s��T�@������O�d��YZD̊�	C��)�Ȑ�Y� X�?iĤ�{����C�� ���"<r���bY-[��B�*h/j�	ݜ�zYS�he@�B�	�ߚ��e�F�(>�]� �8�rB��+3k� ��B:<fD�P�f;UXRB�	���VM�6v�����es0B�	�=��9�!M�\��x���'`�]"��IA��~2C�(1�Y @Q2H��g���y�k��,�� ��m�7�
����ך�y��B�p(*82F�7/p0a�ǁ��yR	�@����' .�@���dӛ�y��G�B���/�5O�h�٠�y2bW�?j���e�Βs�������?T�d�� ��%�)L zӠ�.]Re��=D�(�Do�F= Y�Ѧ�4b�L1;Ղ:D�8yc�[X�� �ľ�rY{W	3D���� ��S�,���H
G����i<D��hq���I<T�t�L>M�����8|O4(Ӓ>!���J�����>���J�m�<�r�: *P) �N=b��<C�i�i�<I�"_xV� kv�I�I�T{���h�<�]�� J0-�&��DjKa�<94�2/�1�U�KKR|�y`�VC�<����&k��`KU�<<j$5f�C�[\81ExJ?	zcB:Z���+ܢgݖ�y��!D�\��HK�G���U#[p��Q�"D� Y0*ٱ&��trTO�#Z�����5D�� �9A���	־ ;�j&�9��"O^�wFڢiL�� i�6_,�R"O��$�Dpp�L R��d��Qg��OR�}�^DN4��NO+6XUYo�nL��`� |{�E��4	0YrG�L8�r���zC�<P���Р����D
h)��|�k��H$�``��Ȅ�t��! ��1шp(F��N�8��ȓ'���
�{!X��0�H���Ɏ~U���ո:S�(�E� +z�k�/m�!�V93���S�� -DVu�AN��w�!�DM)N��j�G��W.�(�ClʍIz!��6I��P��-�q�P��
:h!�D���,�Ҵ�g��(�)Z&Xџh�jT��M[���?��O�tE��i�p�+VȔa�pe���/������?��u���Y�������;Z��I�>5���]���O2�0 �ӗq�&}ؖ���Ia������<�,�z]�����Orl�y�n!�� U`���j�'��5�d*�;��ԉa�:~ 5���I�&ˬ����
���D�P��%���?������|�����܏�fК,Ќ,dN�Y�L�qlџ�����E����Մ�..�<m��J i�OvAВx��I�\�
0*� ��µ�ڷ5U�	�~��7���|Γ(�2�vR�d��%�3\�eX��� ��$\�	H��-��OlS爖�M�z��� =7r���O��NL?���9O�ْ��Q�ќ�{d_H�8SS!ҬyG���F�l��O�U�O��Gӕ[d�q֫[�Z��J��~4��O<���S�z�D��wJ�>]��9�bťo���ɪz���'��'�f52L��۴Z$xq �
p����h΋%�z��'!�����ȟ	�O�9,��9:��G�n���G{?��v�T>�ɇ}��xl�i��j3V�U
��\�t���F����d@�sJt���O&�"��ɖ k���Y�A�7��P�ju���d?���L@~ʟ�DÅ#��H�YW6ip,�$ϼ�SB�W:(�"�RC؟t�4$�|���ړo����o1D�H� �. ?J@� ���(�h�X��q��D�O��?i����|��|:r��"��K�52vƜ�6�Xm���%������O����4���1��\�����aJ�E��Or�4�)���Z���B�(�Q�\�K&�&B����u�؟V�J����C�I�d�咱��0��h��B�PZ�B�&'�ܱ�X�@)�-�q��B�"0�J����V�� 6��<_u
C�ɻo<!Y1���*΄h(�)hrB�	�i�Y�gش �UK@���H�C��:�����_��H�``�m;�B䉆08-G�̔M\�bG�э�6C�	-t���w$)��1�G��'l(C䉅O��$y��X/'���"
�4C�I�>� r��* p�{ �L��⟜9 ���%*l�c�dR�ܹƁ؜	$6��bCD9(k�M�1��5���n%�D�sڡ��Y��ҝu�x܁�d@	3X�˲��d�m8�
�R]>��׻Gj��.��r9(�]�[����"�0�:��WBR�q��&I��hX�� �̤A^ܡyJ>�ê��Ӥ���H�5�T�Al�V�<��	�$La(L����I-�)��MP�<�V#�:	څ�vGN�B؂<����N�<� ��l�,���͆Z���%�L�<	� �d����u� �#&حj'�]�<q�e 3exe' [|�P� ��\�<Y��
�X�ڰvgEuŌ@j ��N�<A�E��L���! <:q�U��RQ�<�"�� Vd}�@�8U�<���@�J�<�N�B���!)�1uF��fH�o�<	�+�35M�Kq��-3*�����m�<�P�Sd:f%��L$(�XhpD�g�<�n>b�l]���D�Igb�m�<� �p�7�� ��d�ᦝu\�}��"O���A,LC~ !0刘pA �k@"OM1��R'�)Xc�HAP@�"OH�K���+X���"�H��ӈ-A"Ox�р�Q�Hh���Q���@&"OB��WS�眨�$$WV��-B�"O���S�*����艮I�>���"O��`�E�&�RmJ���k���ʆ"O���֣�9R��͂��ú-+����"O��i���
 j��w���P�d��"OШ�T��0i�<}i�!��&��0�"OX�tS&#�)��݊E�Vp�"O�ѻ�"F�|���8�@ê�Z�"OZ-T����K���N6�!�$�H�TX#�OS�?�h`'�ΩO�!�Ѳ]�i@�YN�����+�!��I�����W�V�pd�82!���
!���&OJm�P|��NO!�$[q���[��C�H�٧$޼U!���U�(���V�x�P)ႛ)o�!�$�~&�,(��)jo�lxg�Ҭy!��>xb`qAŉ��#v �J�' 'g�!�dE(3�� ��H.5c����Q:6�!�����Z���Q�ti#7�>!��^<7�d���������!* !�S�N0ɂH!{Rrhp�)^�A!�,1��K�aS�86D�����nX!�^�x���;a3Z�ꐊRQ!���R�ƈb�܊J��A3&��� !�d�7?����Apa���N��"Or(����#t�(A��7��ܹ�"O��5d�>�
��ekՃR%�("O�{�#N�+��ܳ�	ճ��Q"O��U��7w=�T�b~�>�1	�'�i��H��ZAT�Ȝ��8��'P�et.P����#NT��>���'UH�Z\C�v][������'�j�r ��RI�њ�͙���^�y2L6�cV4^"�8� T�y�,I�H�(�8�a)&o�|A�l	��y�͈�)��H*���o9 �+pmX!�yRFx�`<�`�	�j��T�W�?�yb�X� �Bt���f6lhqw�C��yBN��9�H�ň�T�� �J�<�yb [.8K�hg��RL$�Kњ�y2�گt���U�J�Z ���+M��y��eY7kK`�h��5�	�y�F��$Qa$��<�rQ��u>!�D��	|h� �ӯ3o��JǨ�$+!�$"9�
]�o�,�R �Ǘ�!!�$ȜqC���j�0���p �[�!�$�l��YQ�dDz��aDEQ?!�!�Y*N�;�k� Vj�F��M�!򄖧��ɇ�%i�i:W���\�!��g��� ��V�+����Vv5!򄅰2�楠��*#���f�52!�D\�O�&5�4�
V%Tq�+ӿ !�_��r��DL�^���HN�6�!�$��N���0ڣ:�$ha�fӀB!��P�f]
��J,V�����N�!��y�~�(�+ޫJ��0�#�9�!��C5=5�$����	���1!�(!�d�1	Ae�U��`E[S���}�!���{a�P��̻vnBP��M�5{v!�� >}�$�Ϟ�&�KPfC�QYL,�R"O4�!����a�4J0�M�hU�;"O4Z.�:M)�T�ë
�Y8�%�"OX��L�PX��x@�ȼ<�,��6"O,
rHA[�`�� ֨P��� "O|M�2jV/�@j�K>����"O|E���aeVq8r�hvb�r�"On1�ޘ��`�b�J�:����v(/D��b N]/V|dKc�
�4�Τz֧.D�l�&�L�l�.x�+9
1���g.D��@�M�;V-���>r�EBG�+D��s��-W_P )@�jŚ�9T*D���fK��б�si]�i�\Ej��&D��3RNE�KRL��nZ;J6*1� )D���Ԝ�Ҡ�b�L�q7��@�%D�`�޵ �d�G)ߡT��c�#D���d��>4a�MG�&d�1@A!D��t�_�l����O�FG8t	`�2D���#a/lY�p9Si�9qw�څ/D�ೂcȄy:�p����򒉡��?D�h��T pi�+��%�vu���=D��㕄Z�G����̇�r�d���9D���s��)~@ZQIV�Ǻ���<D�l4)�	<�dă�d��#!�s��$D�*6b�{y:�e��>���X�$D��##ᙬZ0tPFeP�^J|��/D��	WnƦ!ζLZ��y�� ��.D��Q6�$"��@Fh�o���!!D� ن�L�����鑊f�H0>D�0#�M�@@�!L��ԙ��6D���D,~�54$u{v��1D�DzE�	T���9"��:I�A��i"D��	��_������0S�,�8w�:D���aD��D��c�Ci�$��'�-D�y!�p�`���@Ϭ]�,�g�,D�B�a�@qL,{'(5Z5�\Ȧ.,D�����̡w��˷�ϊ ��$�)D��{�-Ŏ
{T���
mB�8��+$D��a5���Zg��Y�+�9����c"'D�D�V��/g�d�&OI D�� @W&D���� aN�Z#F�+����#D�L�� 
�B��B�<>7tB�3	 �qw�Q<D "�N!@�`B�	0>�I���ߦe�F�⦠�w
C�	!<Α��ee\�ᛲl1��B�	�+�b�3�ی^�ѻҪ#
��C�ɕd�F�8%d1F�b4���:�C�3�z��-�� ���+0��q��B䉄xr aIS��f[��6	�Z��B�I�E�FLѴjȪ���	*��;Rm&D�K%陆y����'׉t|DjR�)D� "���$VJU�H=LZX��)D��b�.AS�d��ԇz�ؗ�&D�tyT�	�"A�4Ԕu�`�J�`#D��	%/�5�L������	q:�{��,D�<��"ݺTOVUK���&b�R�s�d.D��1�+�,!�H<���G93��J�L)D����)V�?����U��-(
r$:��:D�zf�pD�S򠁅/�`Y�f3D�h��7!��ِ��I�Bp�Ԯ2D��5!�i�Nу�%G&���"$D��[2���Y����ņ�+k�i���=D��ƠJodz��v�_�i��):��;D�� ��h��M���[�cb HI��&D�� �غ�̉%yξ���Q�5�|	�"O"�(d�ւn�|䡧���"T�%*O4 ����j呠J�,S�Pa�'���� �_̐��S�t9�l��'��Hd�Z�����+W5k�89�'x�#���m�&9H��(b�	��'��� ��P�#�8cU���is���'��R�� ���-E�h���'�1�A.tB�rS`�=aټEc�'��I�*�DIӢ�<(�}��'�	ƣ)Ypm�G'V�� D;�'��!��_�,���c�BT�-�5��'b�����;��-���?[���'���τYe��!ffe�	�'�@�X
	�\_��PҸn84��'6 d"2���"tuyB��Hp���'�8���ɀS'D�oB5T�{�'g�a�t�̽`O4MX�2��}��'r�B�)����8eS$�X"O����Mg�~H��HM�cA��p�"O��Ҫ�q�b��'KF2AC�"O�r3k�-���U&��s4<L��"OL��j�T�B��@�p]A"O�E��j 3�T�C�;C32�xP"O8p�çc�ցD��()�Љ�"OPub!
�y�,1��4 	�ʑ"O�I;u�3q�ĝ�3�
I	�"OTѦaЭLS(�b)A�&��Ƞ"O\�S���n��Jw���{��b"Or�B�Ǚ4QI"���ڪ{��8�"Ob娕��7;ʾl��m8o0ԑA"Ox�[���J��i2F	]ʙ�C"O�,�7gň��\�C�FCr��"O�Ͳ ��|�^�!75�.hxc"O�QH�O�)M��I�����p"O�墐d6�~��ģ2��X�"OLaʖF)X�hdb�O�����"OP����L*�u+���kv\i��"O�`S����k�6��rVhR@"O���'|(��)F��c<���"OD��W�L
\�t�E�M@� �"O2�0�������s�"O���e�=z(�J�bO�r��P"O ��BY�aP� ���pq��f"O\��e��y�ܵ�⫗;r���"1"O* �.�!{ƪp��T
�0<�!"O�32�ڶ�͐�l�;j�h"1"O����B�	��m��ʡ��IӦ"O��3A&]�E �U��s���c"O�)�%�=�%�%{~e@ "O��Y�ΙlB69 5O�&(�"O��@�`ȶ<��1��M5➜!�"O� d��K}���j�2����"O$������P��Bj���HA�"O|]�Bg^�dHf�	�=A���0"O��e�I1p�X�� )_k��И�"O��ӑ�+D�L��^*s�z���$��p��e��I��\��!ZV"��M>Y�)��u,,�ҏGNϘa/A!�C�I%U�b���DV;�^`*2iY�~Z^B�E*d{�D��=Gp8�
�C?JB䉩Vèl S��jQ�u�eMF�4�0B�x"�7aQ�� 4`V�d����ȓX�ưK��C3G�~}����UׂC�I�,蜝��Y�
<Ȧ)�'�DB�)� ��� <_^ݛ����Ĩ�"O"��f�tX0�q��O��tʐ"O\10&��f��<`쐲S76�g"Om�hb}�D"T�Cք�Q"O����(Q)B���b怚�L��8�"O�Br,	'0;� S�O6h��d u"O�Q3���af$���%�B���"O"�z����A�
tq�(}��4��"O�1� ��=$���s'AW�oӤ��c"OH:�V6%���rf��.��8�"O\�h��5���P���E��Y��"OL�0P�j0��u��~Mj�1�"O��E��uB�E��Jj��9He"O���QB��b���k ٢0�V%��"O���/��2x���m/&��x��"OV� ��m��D�&P=���BD"O:�"u�"H�#��!b�pa1�"O���E�ҨQxXpd��~��x��"O�h� LN 0	�.:�0Q�"OP��Rr$[4fY3|�.I�t"O�}x�O	zptˡ��w�xL��"O�A����6�J�k��T��"O�i�wj	y��bFĒ/!�
!R�"OT�nV��`̩�˃ ���"O�"��2L��T��!� ���"O��JD�w��)��HJ�\hd�"�"OFp�p��y26Lۡ�� L�\LY�"O�I`F�Qw�|zr�.K��a "O��h�4<�sE��2}�8��"O �W��z��%���0JZ�Q�"O6`ba��"<���֮��n����"O�Q�׮^849�e��̃�O��[w"O��!S�B�l��mhC��@��Y��"O^���(��_�Z��Р�A��p�"O��GN��B�H�#'�/1�Ts�"OYC7b �TZ<<��gUh�x��"O4e�� �*b0�YJF�ݻ23 Q�"OF��Q���;���P@[�0 Q�7"O�dz�H�
	�dVf��Q�]"0"O<Qy�W7X�HX pˀ��J���"Oa`��L[2�	��˃m鶌3"O�p�T�D*/Մ)�(S�S��=��"O\���E;G�b�J�e�=K\@��"O�0B% ǩ=������ȍm+��c�"O�9�ˍ���]�l���v"O�H����Q���`cc�x`�-�"O\��%��SG:\��B� {S����"O����@ֶx9�<
B�.I(��"O�q��
[�q�(#���}fN�"6"O�e����(hJt�" E�!J��"O\݋G��
[R`��'Y@�4�R"O:ݡaNL����6&ȨY����1"O����Q;S�8ݣ�5�B`"O�qr�J�A�
-�����8�(i"O�Y��'7����f�{��8�"O~��veJ$Y�R}Ӂ���r�vL�"O,��K�7֊`ڒ��b����"O�iB���:�V��ƴB��@�"O�8���CD���E��"r�� "OL��T��"�-���Mu��`"O$� �1���k¥�)?mr��&"OX���u
D��4%�6��I"Oؼc��
 ~�XZҤ��Tz��x�"O�Y�V��*�Lа�K��}aF��"O� ��s��ݷ4@�E �!�9��"O�baV_`r��%!�3��hd"O<�⣣&К�q� M��Y8"O0|a�*�q/h���iC� �t�`"O(��mH�&��:9�����C��y��[>�8#�/��7m��qC'��y�ǉ�1!�U#P��(2��h�!(�y�
��ZJ
M�PN�0�
!��C�y��S�q�US񩋀0��ċ���y�$�;trd��ڣxʵ����yRJ��`��7j�.x�%KK��y����EF�PBpXFn���y�@ r~���$��8j�-º�y�%�pH+�-$��`�_�yJЅn��J� �O8z]ۃ��y�)1Gp<�Rc\"H���C���y�o�V��B"M;T?�옇�C�yB�԰9�
!ʂ�ۛS� ��V �y�!�0`��d:b��b���6#��y$��8��q�Ę�s�>\S�NE��yrh0'������[�_��Tɤ����y��]E��<�e�Nv�E ���y���D}+!��CX1Q����y��U;-!|S�h�5xx�P#�FY��y�gX�LDXE� K�{��ct���yr�N�K��UH��Y�\7�u9� �&�y�I�*!s��`��b�ޭ�7n���y�"D�lF�s�V�E8�6C[�y��5�:�@N�7�
ث�y@��iq���Q3[J�uW�P �y�^4��Hs4�
$j��aV���y"#�y?hUPqM�r�J��.�y�C��|N)`��h�d&d��y��Ԩ
f =Jħf�%QmS��y�R"T�!�C3b��
4���yRĔy��u��b��E N
L�!�D�<w�8}z2%ܲ"��9"�'�!�d�=X�U�%`E�!�=C%�-0>!�$_���t|QQ���
%!��"���f�	i���@�H�!�Y[x����.3[6쳂&�o�!���*�-Pt��ODaZ��S�!�@��d� �#-@A��l<^�!��];OE�xz�F�@�*ȋ���8�!���q�REC.���@{U��R'!���9����.�+e�le�� �c%!�V�@]�UC�O]=_%�p��K�P!�DU�]$��a��:r� A �[���'׬)��Ñ�
���)���$�B�`�'����5�ܩ�E׉ڭW�0���'#�ձdF��@Y���
�U��c�'B@�)a�;5n�UA�!��`�ꐀ�'�܍2��\�Y����!� !�X�[�'TQ9�-|n�9�j���.��
�'!�U"B�G��6�+ৌ�I2�)�ȓp��Т���yy����߲�8���%�xHۣ�P�P�T*B���s`i�N�<1!AP9H�����F6������A�<��Ǐ�N���6b�bTP����R@�<q��͓)�X���F�Y�i�qj�X�<�u)�(h�^��3Q;kE`|·�V�<��K��&�XJ$`�ko��Ё�T�<���X�Ht��e�e�J`
CP�<ٕb?h;������P���`�Mk�<� ���ߏ������0���"O(�9f���-@Rh��n��I��@9"O�xX6o�u�����K"\��5�"O�������	�C�?j+J�ۣ"ON�C)5P��0r���%��HE"O��[�ݺd��[�@J�n'�<��"O��9.LV����G^قp"Or8i�	�-.$M�)b4IhB"O�I����j� Y�WB�[�"O�]�Q�T�tpM�g���H�t+�"O��5�&K���&��a��Pa�"O��򋃴 ���J�G��B�X�`�"O�������Z�@DG?��$��"O��'B^� t0��E��l�� sB"O���Z--ޘ��B�ċp]��a�"O֕�c��<ځ�R<�B̀�"OJ�`��?dH���߉%�ڥ��"O����ӸP��Ћ��Ҙ_�V<��"O�$Ó����S#A=9��i""O���4*=yH�)���$��K�"O���#�X�I��%ڣTHG"O��#���\�[Ӎ�:2c<@�"O61c��	�b��T�"0:�2�"O���`�V;-0i�LmGR��C"O4�����W�xd��"�e�H`I�"O��f��Cg�uI��A/ �˗"OnI�v��,!�5q�Om��,P#"O�u��s�&EB���'1z�Sw"OH�	&EO�k�������:C��C "O�@ )�I�R�Ab�fx�Y"O��HeE�3V�.��5�B�5k�X�"Ox��$G�&�8s��� ��H�"O����K��k�\�0���/�=x6"ORXB�ǁ���5G
�A'�p��"OR��@��gН�tŇo�zPK�"O��q�ԱyxIC���x��,��"OD�p���YyX}��� ��hB�"O� 2�!�BX �)X?3�0tK�"O虓�)�:qp��894�k"O��`�醅�\�q3��b
h��"OJl���5Q<8�!΂N� =��"Oθ�#��J살�ƠG�U���c"O(
`��y�XD�Շ�$��4��"O�$�g��UoƑ��'�2����"O�y���2T"���љ@�6xh�"O=!�/��!�ƌ�PoZ-�$0��"O�P����Px���V̀X�"O �ѥ��,�Ғ-�(�ĩyE"O���%!3Iz!C�cõb�V)"'"OBu�!g�Ck�P��K�b1�)�c"Oܰ*æ"c���&/�&|�xl��"O u󀣆U�9Z҈�3""^��"O��+�S�T�2Q�h��of�	��"OVX㉙�rV() W�K�V`�E2q"O2�xY���fG�5/�y�i��yB/���Hq�]68��)���Y�y��ԁ+@���脂6�<���eӫ�y��c��ݠ��� 5)2�8R���y���
\���:��	�5���y���";�����h�,1��EQĂȜ�ybNX>)���f�)�v4*�
��'{��J�
S�riI�L�c�H@L>��W/R��TsD�ck����"Y}�<1A��/Oo����6��A@�<1�E�P�F����9v$��p�G�<� &eA	]´�!�K�`�H-��"O��3��G�K�Ĉ�I,S�Dp�"On�2"B�7A����:/��\��"Oִ�V×1C�"��7�@�x1"Orhch��F��TR��N+1��`e"O�l�BI�WͲTz��=��Թb"O��*���G>��
+��'3�2"O�weUh�,a�*ɅΈD"O�u`˃ er>�8�KT�FT�s"O�p���]�+(juP���[>����"O6M#�e�a�u�#J)3�	�&"O���#�6(?���͜�3Bn�H�"O�eH5��7@�e���B�AQ����"O�I�W��\�j��3�9=�@aV"O0��5��P��A�ԢU�}(�0"O�ty�(N(u�L�2Ca�2xj��!"O"D����v&����B�5{�*�ٵ"O��	�0��Ex�aT�x�z� �"O��	����?�vB��6M�:�	�"O� #R��\ȼeq�$s �`�"O�0{�k�b�����2g��q"O���%*̚�d��bh�<��Ԫ3"O`�s�k�s� ���C�*�A�"Oܜ
� YTm"�P6�"�ԨKp"O�<�@L#U��A᥁V�f Ae"Ox��򌕡ڎMڱFM�'��$X�"O\\�%e�	�40�C�Y�$�t"O��P�NI"	�ݱ�aX(1s �)&"O�\R#���a��l�/��QT,�!#"O���6`Q�h�y�e��w���Ys"O�+6��o�@�e'P;/Ŋ8c�"O�q8�Cc�Z�YQFŹB�&���"O���E�؈X
}k�j�,|�v"O��c��׮~^T�� �(�s�"OU�B΀63�Rp��S�2ٜ�h�"O�-U�5H�[�� 1�H��y&�@�h�т۟����>�y�L�,	� ���*�j;�*��y�M�
��U£��r8�����#�y��>W�.(�@"���`$����y�DC���a ��5/_����%�y������a	�+a�*��"�yҫ�T[h4�� ·0��3�W��yr��B�qc��U:���Vݢ�y��&m��E�$ϖ4�&� ��-�y�F�Zba�"�O!!*�U��j��y�
C�/��9��ӳ
ȕ�S�1�y��@?�� Pp땰w>Խ	 ア�y2�Ν&�Ā��Α~�0)G�M�y��@";��T�3
�%���% �?�y2��&lp�Y�#����Ԍ�y�Y� jN�X��KsdM���	�y¡1f@PE!�k��D�$���y"�'ⵚQ��1f]lY$l��y)���Z`�#\'v������3�y�a��hL*�Ǯ@�h�z�i�	�y�Ɔ-v$t�a����4B4�y��j1��(5I��T���èW��y�䔷O�E�'�Μ_�`YP
�6�yr ��35���dB�Y���TE��yR� �
%��9f\�]E�����N��y�Q�*rԙ� ��G��@�
�1�yR�B�[`�`���е.�m�WF�'�yi�L�4�3��݇$a�8
p,���y
� ��8w	J&<�{�dC #��!��"O�c�e�j=�X��C���P�"Of�3A�R0a�D�$醙�><��"O�	���w�����	�Gz�U�!"O��z�F�� �ʂ���n��"Ot4��-&k�9��㉇S�4a�"OV�B0�2%P�}�AA�,�b��"O��p��)��z�o�28���à"O�+f%2�zJC/X�V�x��"O��1�T�iZ�L0��y96��"O��襀��7�<d�`"��t�3�"O �T"�>�`Yб��+�,L�"O���B��-ގ�YwE(r3H� �"O�dqP�R�kn-���ڌFE��Ӆ"O�9�� �3�	0��OK���"O���eS_�&�����Bz�)%"OX��sVu�NM�$CL��e"OPl��-!cjƼ�A��I?��  "O٣�셷[P�H��̲<>�}R�"O�dk1��#����J�>O� ��g"O��0��L�X��:��@�l��g"O�0a�;#.j1�7��f
��t"OH�d�X&?�~TR��BIJ$R"O0��&��R��ɐw�\�L�l"�"OV��m�jڕ�
�_��K�"O���aC�r�t`8T�Q�M�He�2"O	{�BկT*հ�]�N�~���"O�1�֦��s��b�@�E��DQ"O\�Yt%�8F�"��/a��"O(�µƏaڤ����0D�$*�"OTܛ"k�B�}�"@/W��cq"O����iͭ[Ad��p!'!�E�q"O�ִᷮ�9�K�6Е�"O ����Q9L� �%m\�Q��0��"O�̱���*^�> ��Ɔ)�� "O�}�"ɒ�'���j�L�P����"O&�����t��D��[�j�"O���g̷0��cJ�H`�u�s"O�9j䋎 j�v��W#I�+�^�C�"OƝؕ�ՙ��(���E%�ꭙ"O���˲Z�: 9��5f*HI"�"O<�
�j�	6����
�mkH���"OB�����0��	��튜}O���"O��w�Ar6�8���S0
M4x�4"O�I��Wm�\ѲJ�ve�բ�"O�����
Dh�a��ݨH���:"O�!	��]7m� 8$�� �hH�"O�X�0)��.�,XԄϛ��%C�"O�e{b��x�%���-Z��X��"OD��&��gʖ��g�5F�����"O�(�ʻg~$[Obh�@�"O�,v�V�^{Ա{1A�T��� �"Od!�!�G# &HЂ�ݢa��Pr�"O���f�2z5��� mJ�?�V��'"O�,�s���"�`����W��O;��$&�S�O��)�5�G5`6>��6�ܕ"'2���'.fp��X:p´�Ue
D��'H����B�0�\
��O�3݌a��'�VU[C`JIt*�	95a��q�'�$q���<�4�E�X��a��'�@Ѻ��<8���nP�	��u��'@�ɳ"傩++
�Ȅ�Lw��t�'Z!C�,S�&������4mh�Q��'�YRv�E-�L��bNؔi���"��� &I�b�,Y��I��C��}����"O�`�q$��;�8իV텼Y�ttB�"O
Tra �*��Ĭ�4o�@s"O��a�IS#Kf��5kK����BE"O���[x:��E�&�X�"O����#R'0��s��@�D~\e"�"O$��$˚��@I˰HǕRn��E"O��[�ܬjr�V���us��B�"O"�Qާ2*��ugɸfg�@�"Oؕa�? 4���0&ǆ5 �$"O0=�c�%���!p/���y�"O�m�#F8X��<����;B|�%�f"O����H�|8pCǂ;;۠�8`"O
��D��}+�����N�N���"O��Q�C?L���5�ٔ^�F�!@"O�}�LW�,|%��l��b���Z�"O�a�(��o����p����"OlC�\��I�	��
�����"O�:��P(��lk���- ��H�"O~-�eE5y���7i��`c�<��"O���pE�9b���s҈�@Į6"OL�b�^>$��,�bH�	b�R���"O.-���:]�Pؕ�<-��E�0"O�}#k�O�\p���
 bJ���"O��9�ˍw�x�����[,)A�"Oʁhҏ
�9Z��A��C�y��"O�TSp	�90�Fɹ�a�]�ĉ3A"O~4!!Ĕ;'�V�B#�M�p$�p�u"O|����I�p8���w,SQ"O����ݫN��e�%��_:hr$"O�8���ۈxS (�%Z���"O�`��b���(1Z@XL�� "O$h��'sI;��F!ax0�ʱ�ŭ�y���;~�aJnɅc�9A���y2&�� �.󷄇_�N����>�y��F�'/b����ɱ�\X ��y�垮F��\�%� �'>y[�V'�y�O.��{�J@�d�Y�y� �4X��ҠH�M��9��0�y"���*n��S�>��HjEa\�yRJ�5I
\J ��= ��($
9�y2jРH������ڃ*O64���	�yR�ˀG?��ش�͢�t}�Eꈃ�y�. �:u&X��(�
u�� ��y��˂H�� K@DN	D�&)ѓŗ;�ybM�6~�F<�f��P��Q0��M��y���!(� �1�
F�b)�*�y2��?�J��j�P<ޝ�Ζ��y2�Ӯ[�>��V�_%xq"PG��y��4nRx�!��|��}�Q��y��E�<��w@�!�|]��AK�yª�;h�˵��c�b%)v�O��yr�FJ���s�̃]���#F��?�y2�?O��mP���.U�(����yR"��+P"�GG���!Eǎ�y� �e�|�5�Ufp��N��y�,�]�Fx��$�OӚ$����y"K�C�����#D;j3����y�G7P�խ:	����꒬�y"Ɇ�]".u�F͟v�P%pD���y���.����Q�&�d�����y�b�=*��r�i�u{2�5h[&�y��HLXr�Z5Q*8��'I��y"E�M���I���+2o�Y'C�y
� 
�� �Y$99*�G]*k��e"O��9�c�&��c�Z4`EU3�"O����k^���s��OA0�R�"O�f)�"`&}���'3.I��"O��pb�Lj�ld ���t��6"O��j�ED=<݊�e��y�i"O*}J2��7?v����
�!h$i "O�Y���5��ݛP��j|"؂�"O�x����kV��yBƘ6<� yr�"O`H�'([�us� ��̓/_���"Of$��ۻ=���`�[
{VvK1"O�%�5�K5����/Z�T0�"O���#��N6�<�aИ��d"�"O>`�E`J�k�H�@@ޫl���"O	G��{�.��m�aM�E"O�0YS�ΧY¾{1��)��1�"O���Ҫ%v6u�+Ƭ7�Ji�"O�h1r�߁s��A[�J�/T�JU@""Oک�Se�qx�5JX*�~��"O�}��j�?T� l��)^��L �"O��aсŏFW��ǩN)%���a�"OX���FP1MMάJuH��9^���"O61�tb\�h̑K �;�X�"Oy��!+t�ƹr���)j&l��0"O�31��$D̶Իw�$.&���"OF�9��P	wb��� �v�$�Y�"O�Y8�I�u�Ԋ怨[�X,��"OR�[bx��Ud�i3��U�<yd&A�a��!�ԩ�N l+�/�U�<)wA��h��țj�	c7(�	s�y�<��e_,',�����Syb�1lK}�<1u
Ҍu���*p�o���EN�<��d�,��m��+Q��XL�e�QU�<QP��-4$.�S�͉Td�}Y̅N�<IA��%`e��	�kԂS�,�a3!o�<Ɂ��17 =���B56O�9�/R�<AVD�ef���'3t�X����M�<a�+�>����)��x�<�
���E�<�0�B�=U��&��%���g��C�<��Ð�6P!
B�<C����.�}�<�cƜ0z��=K�Dk1���l�z�<��
S?�Z�nY�h�����]�<�5�t����K9l̨�B
]�<�Pm�
P������GNn,���Os�<�F�ױF�T�K��� <%�Bg�<�Sa��#���;AܑK�A�&ky�<a���.H�A�Шғp$�)��Sr�<����7�����J�XHᅄ�p�<��OZ"��1�ף�q>1U.B�<YR�	:@>�T1r-��*��1₪�{�<���AcY�PG��Ԙ��i�]�<��E8co����ȓ:4n��c\�<ysM)h�q�P��R�zxq��o�<�Tꑹq��u����|��G�h�<��D�*n6C�e�%B&�)���j�<Yg*��1?bXp�ߞ6�8��Pf�<�e���N�Ό��Ulr��j�$FN�<Yr*[�;��ℭ�a��=��DD�<�t�ͩB.��fFS��0���PB�<�Rn�=Rt�ՂaI�3Ex��)dmA|�<A�G�%����MU	*v�E��Tt�<AćP8yÔq�"(�q�d�{��V�<e�߼HX�ɠ��?�8ñ�S�<9�I��M�8@Be�Q']����W�<� ����@������^|�!��"OX��R-�\�e���.w�P��"OL�1�+���Bb��s�0�$u�<���j���&�Z�REs�<��![d;�����#M��Pjeǂq�<�QH��W�	� �Y�*��$�S�\B�<�щ9n�͓�ϋ=�D��%�R�<a��S%;�2M���Z�r@XQ�<��gR8�v���Ɠ����g�e�<iq���X�T) �e��Q�͑^�<�s�� ~����#C�d]qv
�v�<p$T*x�>�aC��"< �F�j�<qC��+MWf��$��[�r�����d�<!�B��	(@8b`%��XB	�b�<y!+@AXHs��)Gg�p�fPb�<�]�T�z�g�:x������C*�B��u�.�#gBЋ<����W��B�ɷq͘`0��7ǚ�3҆ʼF�B�	�Nx����%eD����Ԑ]m�B�	'K
�5R�b��-,��y�n��M��B�I�m�ڤ���Ι�,��M)QIVC�I�d�(=���[!t�)IS���C�	��D��i�G[lBR�52]�C�	,Li�����X�h���="6�C�IZp��sL<'���j7�Ө"�C�ɵؒ�k�R5ifȑ@S@�P�~C䉣r�����}��y�g��!H�bC䉊0Ga� c��jfK�OkC�	;0�J�ZW�Mb����ttC�	w�8���EV�e����0I)��B�	h#�1fD�'M�x��$�k�B�I�#el1S���kq��k�W>3 �C䉐_�v�;��ˇd@K�?P�B䉆@��4���YTΕ��Kl�C�	�.�Кn�~J�D����<˰C�	�9C����΁|� Arف��B�_C�Q��.��\l�H��/�.��B�I��=Q J6j�Sê�lZ�B��!FyhЉV/���PD�#��4m�bB�!A��)�ի��*���A�`����'�,hH���\��`��� �`��
�'ojx�"�և�d�ʰ �qG�@i�'�Ҡ���׬!�^-P'Uk���	�'-Bd@�o��T0��率MR^(��'nH,�U	-gZ�X)ˢ���'�@X�ds��Y��CŒ�c�'β�A�TY�8���+��6�y�i�a"�]ہ,�+�Er��J��yRB���pR&
Ĭ �t� �a��y2C2������ל�D����>�y��V"�z5c�d���c��T��y�A�
"L ��M9H�Ś%+��yR�(nD���n��Ĭ>�y��[P�3�!�?X��2�̚�y�N�F������h�b���aJ��y&��=��T�eдr�*!P(�(�y�ѻt�$z�cЅdL���$*���y����\j�3���^M:��.L��y�Ó<)�Q"�ƎZy�D�¤F?�y���;[�Bb��W* ��Z(�y�,�`�t���ĺJ��ܹ%ɫ�yR��s���u�LHe&�5�y�J�=4|����B�:m.4�=�y��*ŉ_�^��iq#�2�y
� N���#W�&�Z�l��OA��RR"O�]#po�Ex�I'�T�I7��;"O�-��'r8kr�W5����"O�M!��Ҹ~�jr։�v�^��"O
h	����4Dpq:��=yv���"OX(3���,�J]r/Z%L]z�Q "O&81V<Q'r�Fo�>[8b�:�"OZ�9E��n=�={f���8��"O.�
0h�I:�������X�"OH�Q��$@H�|!rg]�i��!9�"OD�J%Z ��q���Xm��W"Of�s1�޲DrM�-�?<�-�"O`� �G�;90�AON 8@�8�3"O<���^9j�۲ ޽@<:y""O�h�C��U2ܜ��٨q�Ȭ��"O�`��74.x���]8�`�"OzMdC
GZ���d�ۥZ��
@"Of�q!	��0�<[�ޖ1�dز"Ol����բip��8�ʴ�%"O�����9v�2qa1�8w$���"O�!ٕ���~�NPs';i:�"O������w��L(Sl�Og
�B"O(c��"�f 1p��:_�hʵ"O*�0#"X6-N$��U�C]�hB�"O$R���qPQQ�eD`���!�"O�����|�t�	VƋ�w��A
�"O��QD��A�rYP�ϙ?v��"OZR��E1@����Z��v��"Oؤ"Q�D��� ��I3c���"O��q�,�!
b�� ��$���"Ofl�S`��p��C�я;��I3�"O摺M�<e�@"C�8T�pJB*O����䖲����ƅق <���'���΄����P����ui�'8X��G�J^�m�Wf�D����'���apC�&Ode�t�D6"O���O� Y��`3Ah, 3i �"O�� �ӝDn0𩓾B^XБ"O6m��� d��U/N	-f���%"O�@rn�=+`��P$<6T�z�"O���ED+3PP�҅�`"���"O`�d��6_&� Ӳ�/@��"O�����^�w���#hQ5t��}��"Od8�թD1eJ�9��8m�Xe
�"O��� ��5��!�T�ӀT�U"O0H�s�L��rB*.F�vr�"O�-���ܽAmDU�Ԩ�0z�I��"Oadj��)gS*&x��"O��s��:kv�s���zT��v"O���b�[�@ h�Ď�UB�pV"OB!�����&%��yr��)pj�	�"O����
E>e�"m�AE%s^���"O��bFL�?����.�
]-�ı�"O0E[vbӉ|�P����ѹ,7~�C"OZ9U�+=�d���T��p�ȓ?�]1R�Ю|�`��'�/)`�Ԅȓj�"�9��"	�Hx"��F�n�l0��3_��i�/N_�bYR Pyޑ�����2&��@5t��$��sD����;��x�Ee��Ab�TbIHH��K�ڱE]�9�9�-ԨJ�q��w���B��܏M�| �L�D�� �HK!Ƅc�D�#�����*K���`'V������ĎІ�S�? � �t�bLx��S:��a"O�m�`aVA�}86�M1�ܪ2"O����!`���@���"m0����"OX��Pg/KY�eA�)U{&��"Od-�%ܰ|��i��,r�ȴ�I�J�KV)e���	�9���@�G�# E3��RU1qO����9/!~M17�k�(c�=Z(4��P�k>��
<k�8��CE옔@"�-e��y�,S�"��燏�")���#A�i0pM�0��|�:h�b@��J�5'Z�6=4�PL>'Z�Y�4^y��'��	�� �Ss�-
��D	~d��0��iL�O,F���A�Xبӭ�9`��aR��Cp�󉶩M�R�i��GXx�>�{���\ ��kG#�<�~���$��� �'��i>�C�4�ē< �d�6@Q�E40+����C*���@�]j̕�O���Ɋ��ݓIX��}Z����{��EUcp�q��VS�`YA!�b��-���A�#hfY���Ѵ(Dё��4�r�dU6�����ЛNI��-d�&�ɦr�A�O9l���M��و��㒪]$�ujVI�&]��;1�^�~��'���'~n�1g�8��(SU%�!ĞM؈���[۴����]w�����2$�D8��\�l*����<a��Q(va�v�'4���ďyDdP�b,��"����_�N;,�W��:��\Y fŐ~6��O��O\P2e�X�Q^�����׏��܈Eh	%C�J��
>_,��q/
���i���|�wH&���K������)7`yceN����M��LB�����?Y�ʹ~�'"2�'����	�L�,R�⋇L���S�E6�yB�����˵�>�0�t�Y�>nڿ�MSO>�'��,OL��t�z�q�K�30���4*��xh���G�OF�D�Ob��� z��$�O���H6x��.$���7�V�b��A�(����"�E�I��ʂ��)9�����I�/�X%�A�A�}����G���kP0aKX�S�(�1�(Op���K:'�lCƍ�%&��E'�K���O6�=���튘)2@=���@!8��a+�4�?Q+OJAm~��BP��%�����\�}|�<p�՚2!�=F�{���6o���*]�N�D��]�۴���֜X�"@o՟�'>-q�D'R���	��P�/��ğ��S��;�
���6����ǮȠ(�X,x'��Fg�G���1� � �� )*ҧ ����0�ʻ�M3�n�-:oJI/XI�b�^1tbX�jB�ڥB"��B���&��J��O��n��M�����)�+!R�ݪq��Ghʙ�C�ڞ)�b=۴��'��"}�ISO:`p�GO���d��@O: ������Φ19ܴ�M�G®b�a"�픒j&Qb�b�g?y��гc����'`rT>��6kC؟d��ǦͲӈҎ~�$4��SF?�5��nҬ3��Uє��x]�7%W�b����N��D���������'�5�a�T�Ia�Z�rj�%���L��Ms� 	(�W���4�\<8�!��I�����{0J�|�1/����E�#G e���(I�n�m�61t|���OvynZ럤�����6HA�N��<�cs�18��
��~��'�ў0�>Ѳ>d�1BI5z��@0��s�'IN6-Ҧ�	��M+�-�i�Zw�*C�^5y�X��%iB5[q-3��5lO$LZ& �  ��     {  �  3  W+  d7  WC  KO  [  �g  �r  6~  ��  Q�  ��  b�  �  h�  ¸  �  I�  ��  ��  7�  ��  ��  g�  �  ��   �  C � � � s m' �6 �D L �Z fi �p  w d} 2�  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|`I!'G#\���%�T��'ItcbꀀK<�k��̥:O��'������Ǝ8�ݓ���"J�S�'y`=c �d���	%�BPiV��o�<)E�I�M��c�Q'��I���k�<Yb�`��s4��/~�����M�e�<Կ��رD�E�?�t�Жgd�<��j�aZ����Aّ'�F�r�b�<��"���e�ďfe��ѣ
�[�<Y �{�<Ԑ�[�0�Rѳ6aE|�<�ǆȕP�,x��H�o���ۀj|�<��\��!G	��lhP�qI}�<�cێ�,����ޣ��@�#��x��G�<��Fъ��u��Z�JQK�%v.1���� ׋� ^r�Bэ]lr"����Υc���!� �u�e|���ȓ_�}�㧟���\a�R�i��p��>�
H�?Дk ��t�Tلȓ*��5�&5y�d q%G�=QG>ĄȓGq�E@ÀVV�p`!��[�H�h���s�`HqH�Y�T}���ńi��=	�G$D��@1ib���eG�6�,�r�o�0��I�&��p�W� =O�AH�� ,P����D֪���8"s���G
�oºap� *}�C�IYW@	Pd]b��10#_� ��C�)� R"0)R�o"\�"e���v�X��"O��� ��)" u�g��w01��D|���On"�q�Z"f����m�,v�M��'�n9Z�HVYڢШw��)�8���'EИ�Ei�
G��Q�L��Z���'}�ݹ��f�i�6�F(]枅�ݴ�PxBjTWNX�Q꒘L�L�yV���=9���P}r�'[:��ƌ&)�D��h�X�� �'#I&�;#*��iYd�&ъ��Mh�OaV�������W���hc�!
�'�0��L�Hz1G��o2&R,Od�=E���N�T|v�8��?q����bI,�y� �+v�.m֦dVA���8�y�k\�0)��Jf�^�4��2���y��M��dX����Ua�uz��y��]�h=&O^ӎ	�n�/��O:�	�M1�8i"��OE,��*= ���F�B�@R��qfz؃���l�<}��A���}V�̵C��E1R��>Pe8�˱�f�<$�ץ:�f�f,R<�-�5�c�<GnX�w0&�CP��|�%C7-�\�<�lH�E�>��ߴ5nݺRi�_�<���<t����6(bf�2Ԭ�u�<b@A�'cp�*ŉ5IY	S�JRp�<af*V�o0�|�����m� �2G#\m�<�W�%�je����+\�ޑ��+��<Q ��g5�$�����|��G�Nx�<�3�Z����w'��/�(qˠ��}�<�6�F3n䬴����z��+�n�c�<���V�{^��uIPn�6I���^�<!��T�bh���Тs���"[�<q��>w�I�e�l{mH@@V�<����B�f��qT`��GP�<q"��:C,bT�! GI��b�MI�<)��U*5� �PB���'���A� MG�<��DF> U���K ^E�$j�DF�<��G��8@�M����r�~�e��m�<9 +��e� ��1 d�8F]d�<�@�ȸT`�8y�FB1�8D����[�<A�\�[��(���qD=�6/�_�<y���g,h�ʘ�峲��q�<���S}��h�BZ�\�ಁEy�<�e)ϢW����"�L�k ��eMr�<i��G����� &_����l�Y�<Aa�ڱQhI����$$t����I]�<"*̈�PBp�4]VTaUY�<� a@�~-D@�c@� �}"R�_z�<Y��נ9�Ւ�#W�|^� 6NKz�<A���$4�R!�Ҍ��a�\�<�#d >m�V��(�#�Hl�<�H\33��A;��؆���i�<i�i�1=���sJ��9����e�z�<y��|vH�i�d��P�P7	N�<��a
�`��fkB
2F�ԐW��L�<�ѦR��D�}�Nl(���B�<�E�̒zr�ዀ��(p� �M{�<��IJ��� ��o�o1�Y���p�<�#�!� ����6�9x5�m�<��l��f��/@&T|�lm�<�!�nŨ]:�)����ɤ�o�<��͹A|������>�(C`�`�<���=5~V<��)	|�)����W�<����='����C�]�������m�<q��@���v�Z<� gU�<� eI�j�x�\���X�~c����"O���a���I�ŲSK�W)L�`�"O�Q��P*.�	qT�F=��"O\	a�M�=BT����F��ؽ�"Ol��c.����2���M�N��"O� �d��Rr�LQ�ٮz�#�"O2��f ����ʣ	�1��"O��+F�(%��q��,P�(��y�"OL-J��Z�	��B�	X#�����"O<��uAf|�jG�T{
�k"O�i�!ќt���$2e��"O&�)U�+��x�A��:RΜ
�"O.��P�N�^L8��f��={w"O~D"�lإj>
̃$ȡ��Z"O�\#�� ,8&j`ò�*�L�!"O�Q@��x���qNש.͊x��"O�����t�~���M��z�Ȕ�"O޼�K��)��ae셺ib�qV"O��	D"Rd��ݛPk�2B����"O�����.`��9YqD�"E�0p�"Oa�bK;l��C�3^�^�[q"O��Z�E�:C��4��16��k�"O0Y��g�����f��7�l�4"Or�*T��O&�p`R�R��!��"O����UCeD��ѾK��Ȅ"OJy���Ԇ�4�8@ ��Z�<�g,�J��CsB?����Ϝp�<�7�FG)8�z���T����d�<��/ӿnjf	b$�/A�P�q�Bc�<aR�6:�V-��O*|�ѫä�v�<��a��H�tR#�Ǣ��!� �o�<��i	'0=�A
6c�����Bm�<YVC>T2��I3y���A6��T�<s�(!�ܛv�«xC�HL�Q�<9�B��69j��Βx2EAU��b�<��Ζ�C�dd�s�	��Ԁ��
e�<iT��Q��s�
!��!�(�b�<A%�E� ��<��G�p�$)E�`�<�aZ���c���'x�q6D�v�<!��:O�� ���MC��]a�gNl�<�Ï�,����[�17ɕB�<�e��-d���X$iB��X���|�<Yg��PW�����?}��(0!B�z�<	p�M�Y�v�C&#
�&����@�X[�<�4�6�<�����%eZ �6`T�<A1�o`MCa憖=h�-��IDM�<A���-AD��֬
xv�9�g�^�<�Q��v�h'�)Ԕ�v��V�<Q�e�H�~�耇B0\vQS�Z�<Q�^#
d�}Rff	�S�X���R�<Y�Nɟ+��$�6�A=} �yCP�y�<Q1倫,{��R��84�t��S`�r�<qUf�Y;�9���.d	�ˉn�<!�K�2.jZ	S��,=�ƽ��!�N�<�#.*G�`�'�֣mފ!�b�G�<钦M�#����F�#�&ؒ%LHF�<��,Pf:��(���E�nEL�<A�N�"w;%E��6��eh�^S�<���/C?�u��חJ�X���L�<�%
'H`lK�O�&����g�)T��c��)}�2E2�[5����C�5D�h3�1ĥPD����e�5D��:���=x(@���dB	z+�����2D�\kr�:Ǥ��a!��^�L�z��%D�� �e#P������+��[�]92�z�"OVaG�Q6m�q�?����"OBd�w��;2Tt�#k�6���"O<I[��˂c���[��ݍ�����"O� ����	��KF�
�͈����'��'9��'��'�B�'��'�0�
4��	(�T�'+��h�>��u�'[��' �'���'���'���'FY���P�?�pe"a �"M� ����'s��'��'X�'��'�"�'�<�Jvm��v|���"�m�<�s��'���'}��'m��'`��'��'�\-��7�81C LF/~L���'���'���'{2�'���'%b�'����$�BE���.zǐ�$۟��I�����ϟ�����T�������ٟ�`q�T+.Tc�7$��r'W��(��ޟd�I����ß��	ş�������(�5l�X��Eˀ6�>�x́�� ���`��ȟt�I� �Iş��	���R�MB"U)��K�`��&\Y�A�ٟ��	�H�I�<����l�I��������wKJ>�8�E$��[4,c��A��4�	� ���X�	ȟ�����@�����@&��4m;aÝ/E��CW�������0�	����I����IПl���������bz�܋EK�8��d�	ǟ���⟼�	��\�IΟ���\c7�+&tt]S��j����� �L��������<��������M����?��b0sԅ(0 ��x 6h@lO�{.�������������:Ձɒcj�P�]�dS��U'EN��N�6�4���O<
�-\RU���"��T����O����Ŵi_���|���O�c�vQj����c�Ęro���<i���1�' P�$p ԅ=����WFOT���i̳֚�y�)ʦ�+BFt��7�Up�q�a�X?\��	ȟ�͓���,}�X6�u����Ə"~w�m`��f�B�+�g�Γ7)}�����'��)�ѪQ�[��S���	��'��	E�	#�M���\̓(�p�$�ǒ<����M؅��쁊�m�>����?��'��I�F�`x��kE2�R	B�Ì����?i��� Nr	�|j���Op	#��W��)�N�(���ᄏ n��s-O2ʓ�?E��'�ФI�ND�1U:ђb��)�䥁�'�v6��sS��2�M[��O:�K4�4���)"���u�d�`�'S"�'���Z�a	�����ΧX$�D/Q2���s$�;C��°� �
!'������'�2�'S��'^fy�E��* �9��M1��B�Q� ��4P0�)�ȝ�?����)�O8�$�!=Ҷ �d�qK����&yԶ`�'26��e��4-��O6��O�JD�CT�f�%�̝�qv����R-,p�!��'��-��gWM���B��H��O�l",O��C���+���*$��c�����O����O����O�)�<Ӷi�:Qӑ�'���ɢ	�,�P��	�$\И'��6�9��8���尿�شZ����`����$C-h��c5	� ��ⅹi��䈼x��!�S@ן��e#`���0��))�ΰ� CB `1�}�UgJ����Ox�$�O��D�O���*�z^�1���Q`����!����I��8�I��M���|��q����|Ro)rI##!L~HL'V�{�O��l��M�����!۴�y�'��1Bp�%�`Ȗ��t��Gd	l@`l���l��'D�	����	ޟh�	�d����.�'T<x���k�q������'V6�X�
����O���|�c�M�nmā�f�z��y:5e�o~rϺ>9c�i��7�۟\'>���-�Ⰰ�D�&<ln��~�H�ۂkθF���#��ry�O��	��'� �+tl<,I� ��F�t.8DHS�'���'����O^�I��M;��A�Y��ň�a�6`�B�QM]�'�0���?i׾i'�O�5�'�F6��6�`xb
�3S���T$F=jn:�mZ��MÆ�۳�M3�''�e�RK����"p�	�r�qI�Nʸ%by[2�E�(��IWy��'t��'xR�'�rQ>{筂.��p�w���В I�(F9�Ms��?9��?!����0���w��TI��A^���Q5|�䉡��O6M�]��\����h�Q�h�d�ɬ-�$��B#*|�Q3�}N\�ɺZ	 ��2�'n�$���'9R�'�&�h�
�4 ���ub�]S�@�@�'�b�'Q��K�4o�x���?A�3Y�%"v*��PXqd�+v=`�rê>!@�i�7MQa�	�m��sDk���0@��c]��I��x�+N�t#*I96$^fyb�O�ر�I�x�Ҫ]2 4H���B�D���k� �3v�2�'
��'-���HZ���� �V�:�ئm���A�4|b������?���ix�O�N�/���z`
��8�=���(?m�dt��o�6�M+@���M3�'�R��$^L����B���$���G�$��%d�>J� ���|2T�����,��ٟ����dyA"I�'
Qc��2r�d9b�GyB�~�ne�Qf�O<�$�O��?q��hں��@�H�-c���"M=��%�f%{ӞX%��S�?u�S�rJ]��î9���`Iϋ@z�M ���@�<�''I!#�͟d�|S�,�!O� 0}����GpE��A۟l�IƟ���˟�iy"df�Θ� �O�Ha� 0�����>�^i4��O�0m�S�>l�	7�M{7�iJ�6��'v��2�J��#��{�(BO#�%�scl�V��ן�Hc+�� @���Zy��O<� �0�F�{��d�VM/Bs �s;O��D�OH�d�O���O��?��͒~������Y�iѺ4p"j�����ٟR޴F��i�'�?Yb�i��'��@�2�ˉ�4��5)Z�K�n,��Ѧ�sٴ��w����M�'�>-
��J5@Z�)��)��&��Hȁ��\� �|�R�L�	�H����l��%}�X,YG�ӜV*)�U�����Cy��t�`�x��O���O��'j��q0��$2�5 �ӊ+1r!�'i$�5�F�tӄ<&����?i����qڐ�C8�R:s�*KD�p��<�6��'���ʟ���'��	�l� x	�I~f��p��0`f}��ß��IΟ�i>y�iV�����'0�7-U�*���u�
%�p�4kք+p<��ɰ<�ֽi��S�d����$��8��9�E�b�J�`���M3�i�� �ƴi���9��ḱ�OT�H_Ll�p�3I�����NF�Mk��̓���O~��Or�d�O��D�|*ӀĂm�h]$,H�8׀��3β"����2��	ߟ���v��'Q�6=�N��t���K��Q��+G�\ Pg��m��<y-O�O�:���iE�B$lT��ph�&�HuF�#T��D�j��;��@gF�O��|��x=��+�J�E����%Ѿz�Lq��?݊�������%b��gy��'���{Ѭ�Q��!�Gpp>!i��$�o}�}��Uo��<�O� �()-�R9�f�ՓӺ=j$���r��*7n�exT*0�&5d�(�����)E�1֌8ae��M�����O���Iٟ�I՟,&?�*�ၧ1���imB�]/|��yy�FJ�v|J$Z��'��7�E�/.�ʓ�?	O>��Ӽ���K'����	Myk(D�<�F�inF7�Z���ʢ`
��9��?�T�7�b�	H�6�\�U+ԎJ�@3�D�O���0I>Y+O��O���O ��O��#��?(�����/V;[HPu��l�<Qs�i�,!K��'�B�'I�O����:v�H��ID�m�@P��][J�-!�V�m�.�i��?E�	�W;~*S��"yGb�{���b
.�
 �S�2~�gŌY�T �Oj�ZL>�,Of��pD� $"ޗdk����O���O��D�O�	�<�g�i�r]��'�T�z�CE�;D���-� ����'6��O��Oj��'R�i�R7�|�pa#�NƐ���>����a�����ɟtzBeX���$GNyR�O'�� �y߬Yi� 7`!J
��y��'$�'���'����;6�"��Ō6���#��L����?9�iFk�}>9�I��M3�����A� ����ѱ�@pV�"d�$� �ܴ���O|䓣�if�Ɂ54�〭��".4�2 ��s�@�sPn_��CCz�	qy��'�R�'�LW0=�@x��G��U#��A�R�'��I�M�E�ў�?q��?�)�,�4�[.�n5��"�"c�<�䙟Xj-O��DtӶy%��)��N=��h�;��Xȕ��b�X�J����t@!pK��S
���.ri�=��C��?ɥ�$}Zc��Z���	J �"ɺ�l��+�r�'�"�'���4\��+�45ߎX����Ϡ�K&
n�\&��?��B@�f��X}"�l��4�G�xЊ��m%+C��5�D¦�ش�E��4�y"�'$d�f.��?!rZ��ac�=jC�
���)_;j�0e�ܗ'���'Q��'���'A�0f#��J���>����"=^���4�������?!����'�?I���y'l�Y�Ɓ9���|�x�g�^��6������L<�'���'4�V�zش�y����V�,� 7��'z4�'Ϥ�y�ςq1T,�ɴx�'0�������Ɣ놡��iv@I��ɞ�b�����L��ޟܔ'ψ7mE���d�Ov�_�����ȨM�>�#��I���㟼ɫO��l�1�M� �x���2 �z�c1�F$;��1ul���y"�'?l䢳@�@�Q��_����Cl�LV�L�"k�c̉�šM"�&�1���`�Iܟ$��ԟ\D��w]
y3���1 
Q ]�V���r�'G:6��<��	��<)ݴ���?ͻzLV]���;nE.eq����,Y>L����hӼ,n	��5m�<�������%�j]�k�ؾ���+2���@��������O����O���O��dR�2�R�Q�Pʨ�1�C�(mp�ʓV��CFR�'�����'D�iVʂ5[v���u�P�D��b��>�$�iw7���'>I��?	9BA��W��:�"ED�B��8#��y��@xyrU'φ��ɡ��'��'JJ^	�ʞ0cB�"��=4T)��ԟ�������i>Y�'ʺ7�̹_�:�dH�'	af ?q�d�!B��Z��dRئ	$��I���D�ئ�[�4!
�� mC4�X�gE
Q��c$�ΐ\ְ�і�ih���O�ى�+���z�Φ<��'���gȁ~���P6�ڠ[߾Rs��<���?���?����?L~��'^2�����I
�2�
��u���$�����?���M���$����'oҙ|���{aX�O�=��U�+L�l6Lk}R�x�ڕm��?��[����?)u�G=a2���R��hy��gM�Q��AB��O���N>Q/O�I�O��D�OR�;6 $q쎓a �t���O��$�<AB�i��S'�'�r�'j���OS��'Mz`fG� 5�L��'R┟P���u�޴'��O~��c�;&��X1b*� Gx�@��"ar*��uj�O�iQ=
��]��?�/O8}0�A�-�0n�_!Mqꠃ�O����O���O؀��͑R����O�������U���T�Bb�<��,� �0 ���	ܟ��'y��'��6ƌJ�6��릕���}�>A"��p�Y�@���M�i5b�%�i��؟�<��)�:���O��� �a蒍M�7�!���,@"b���iU���'�r�'���'���'v�S�@lh5�eg� N��'dA'%����ܴ
�����?i���j�'�?1���?�;�\�+ă?/����Oҿ8b���c�ie�6-J��m�O���<���e�@6��l���,}�<�� ͑"����C�k�Dʲ`��H��Yy�O�R�P%��ȩs�T�%)��B�d��\���'t��'�I��Mc�a����D�O����_�I�b9c�h�2D
fx)դ*�����C��EQ޴ȉ'��Hz���i�>-��H�e:Թ�'��Өo����������?����'uh��	�S*��&Ȇn���B�c�8���ş���ҟ���m�O�Bj.л�
,���{a变���c��3���O������9�?�;�u���D�<L�5�I�9<������b�N�lZ/� Tn�W~�
��P*D�Ӷn[�)i6�3�^,i�S����@��|V�h����H�	П���Ο|2�Om[���s�=v���D�Rvy��m�|áe�O��$�Oؓ�����e���9���%��P�eU�|^!�'�,6�Ħ��K<�|�愊�MRv�FD�J� ���6/���I!� ����_���B�����O��6��a�tDM�y��]�� �U���y��?����?Y��|�-O�!o�����	�hn���!Bl����Rn�R��I��Mۊ#�>� �i��7������Ӡ[{�"갩V��V���X���%o�D~2L-b�����H��O�'���x��V!Ū���Aʁ�y��'(��'<2�'=���Cd:聁	�?g�v��U��8�$�O������6dw>�I��M�L>�R�ҽX��-���[�,$
�ұ(��'� 7- ��'w%�l�~ҥ�z�āc�G!1H� P"ҕZ����L�ߟl�|�\�<��ܟ��I����ŭ^�`c�&�� ��[���ԟ���{y�Mnӌ�"�b�O��D�O��'?1 BэC��<ɀ#ܾ!l�'� �1��f�Vx'���?��B� |oNu����l��yǩ�,�(@g�	�|�'��L�A���ݟ�'aԽ�f��.y9I�K,MJ��'Q��'R�'�*@ �O��ĲaR��_w�\X��-�s�V���/�)"�����z?C��	v���K>ͧw��7O7mى_0���eX�ú�r4�G�/�l��M��ƿ�M��'�F .��������S)b@��@D\^�Xs��ѐ��D�<i���?Y��?����?�-���b�Ł J1l(SB%�I��9���	�y�����V�	����~k�Y�	��h�i�E���O�e}���"�><�ll�aS�M�ii�6m_^}���N ��1O*�:b��
7�����`�,�b�9O.���-K"�?�F�2�d�<�'�?I��
�<s�)q�|�Ĭy�ă#�?q�i�-{��%��čڦ	��F�?�������1B�Xͫ��C�)��4"���o�	��P�'�L6mB����ڴJ��%��+���(x�xKr#�?a$�ZQta�ա6~�D�|*���O�D��B*9�����k�D�z�N���?��?I���h�~��oE�a�L�+T����GF�\lh�dڦ-�`N\۟��I&�M���ӼsM�S%�ӓ�3�@}1�'��<1�i�Z6-��!A�e�Φ���?�
Q�2|���̋G�t$SAO�@�ީp�MS;W��yN>i(O����O��$�O��D�O��aH�=#�Դ� �,[ضd��I�<QB�i�!˖�'b�'h�Ob�I<5/��a�b�%|:�e"�ΤH���4כ�Gx�p�	[�S�?��	�az搨D��&s0��g	\��/�?j�Ĩ$?	w�*g���T	����D��+�(�s�nU4���@3*�1�\�d�O��D�O$�4���	#�&cOExb�5��\�r@��^�R�!Q�҃7��n�����OR�nZ1�M��E�vA����R�����
{<��6�Ư�Mۘ'��d�������/������1}��d�D2P� hg"r�xA̓�?���?����?Q����O[�hpiT4H�(��'��"���:��'���'~�6mϥc��i�O��l�\�ڶZ�oG�>3�U��l
�\1�����Ħ%R�4�?�3g���M�'�"ă-�&�$��� b��iH�$P�.D��mo�'��i>����	�T7L�H���g�\���G�Q6��	ğ(�'At7��$�$���OT��|
�,�8[E�Iy'�&'@���d~�L�>���i�7v�D$>���+?ix����"
x��ڵT,��S�W�>0 B�0?��',8����!��r�d�1��1xܹb��y�a���?q���?Y�Ş����ڦ�PCQ�5V�)RHάG���dI�2K=���xz�4��'��Xa��k�n��=�'C�[�&e �W1P
�7-�OP\�A�y��IΟ`37����K ?)Î�+Fp���ìif	�,��<	(O��$�Ol���OJ���O��'J����j��вC��H��e�e�ie�8�`�'r��'��Osk~���@�o���)ł�j��Q�O$+��plZ�Mӟ'@�i>��韄G�ǦE̓�Ƚp���x�⥓���'2�Nu�
��	�l�O>}*K>.O�	�O��'cд&���lUl7�Y��L�O\���O��<q��ix�RF�'���'���0R*@�uw��@����Z�%��c��~��I�M��i���>1!��V�@�� y��҃�X�<��[�UP�"%(�9�'������sr�'C�*��<�Ь`�P�=�S��'��'��'�>���X�q� FW9d�aÑ���L�����MkCE�3�?I��)���4�nU��<�,��$i��Uh�l��9O@�o�3�M{���Ν�޴�yb�'���I���?QP� L��af��d9dā�,;���$�$�<ͧ�?i���?9��?��B�>J�`lZ�.�9�Q)���d���͂4��̟��	�$?����&��M�2�R q*��.�ef�Li�O�8l��M{��x��� �W�!be��*G���*�b�����@����ɩ0������'�^'���'ƀ�3��Y�Y��H$�J�Y&Nh�s�'-��'3r����V�L`ڴc���!�%c�����jh���N�}v�T[��:y����JV}"�g���m��M�E��w.�@���g
�y:�gѹ2T��Sܴ�y��'���*g)��?]� V�x��ߕYK̶�F�ӳ�J/:�
�"�{�h�I쟔�I����	柬���lC^,���WI�8u�Q3�?a��?�e�iɔ`v[�@��4��J�r��t�Ӫ!��q�BN�L߆��ĜxB#|Ӝio�?�ʡ�Qɦ}��?��l�"��x�d�[�X�m9�	I�z����O���O>9+O����O����Oδ9�c^-L �Q�d��̰�	�O��d�<��i�4���'J��'J哇l��R5�!D }G�ֶ]��R�ɞ�M�սi�R�d"�	�,1頭-	u�9�u�� qю� ؎���C�3P���bw��O|*J>���r5H)±��K��#D[0�?��?����?�|�.Oxnh[l�ie�b�0���[$V��RU�۟�I8�M����>a�in�:Ӂ�%Y�10#S�`3zeC&ofӶ�d�$tt7Mh���vܔ�1f�Oa��Ҏ@�'F�[2�q�3�C�������O���O$���O��$�|���OB�lE���P�~a���q�Ѯz�F�2H��	̟L'?��I��Mϻq�|���D�*u��=ೣ)Q����'O��>Op��?�����`Ǧ�̓>J�\�C�ƲiD����"�͓>�)c��O�,�I>y(O���O��['�F���r(r�L-z��O��d�O��ľ<װik�0�_��	�Jp�����U
����%8+�JX�?	fW��ٴv��6O��W. �"ůZ�dg��R�h�X��'��@�@X�&���ʋ����ǟ���'%�|�����}p�+O�kcH8�S�'mB�'�2�'w�>��	�DZ4P�vm6�0�`�>l�ސ�I��MCai���?���$����4�XY� ��'W���~ �u"�0O<mnZ��M���/��Yx۴����ir�' ����ș�:
�{U�]���(�u�:�d�<�'�?)���?����?�JѴ	Š�y �=u��b��5���MŦI@PWy��'K�O@b'*�,�˙�!F�)RĊiWR�̛*dӌT%�b>��D/˕��d Դ4X�e��*��sЀ��ocye�e��e���1��'��Iu:UY׊�O���CuF�ap9��ɟ��I���i>�'�b7�U-u�4�dS�H�|lA���/!�<��C�Z�G�2���ަ��?��U������i�ٴh3� CC�rO(0p���)2�E!��1�M��O^�h4E^����%5�i��(�6I%ha� �ڟA�"��b2Or��O0���O����O�������L0<>n�§���:B�{��XG	�8L�O���Q��Y���ay2�'�rU��Qa-~y���"D�q��Ph�L��M��_�l8ߴh���ONa�4�i��O�(8$�K�4��g�H�](8hڄF�9e^VX1�rV��OR��|
��?���G|h
�e֒7J\���>����/X�?�)Onړ?6���ϟ��	�?y�]/-���8Sb��L>��w��xټ��̟d�'��i<�6K���?e��K�U9|��Q��*�>4ڳc�9ʀ4���@!+>�:�#��u�i�O�U����"�
-�Q"�˅ �^Ȩ���?���?��-c��|
��?QT��.�4-
0�&�2ՅB�\���'<�'���'i�a��Ш?O�mZ�O_���pA�_������q�؅�ܴ�6��R��F����Q[��t�~b&E�	.����E�spXЖ  �<�*O��D�O:���O����O�'^�Us g�5WIw��?����D�i^T��V�X�	l��������#%�3W�2���3	Hx��be_JV���c�@��R}��ċ�*S���:O&�K�aA'C�Ĺb�lՊ7�|��F1OtR���*�?9r�7��<ͧ�?Q���?�4�C��*��X�À?�?a��?q��������� e�ڟ��I؟�9u�X�.* Pr%�>>�t)�f)�X����`��Ozam��M���'��I��Jub���7~�����j"�+oD a4�J2b�8H�M~eb�OH���n��H�ۥ�� �*ѯbn��s���?���?����h��n����M�u.dI��L5l�<��T��	����L�I �MCM>��Ӽ�E���.�~11�GuDr����<��i��6�Ѧ��� æ%��?w������i��GH�!*���$'^�A�	�( N>Y)O����O���O2��O�K�mՅ9�:�G�_�TIi�@�<�!�ip���'�r�'��Q>���wԞm�V��7�nHѯ��h�Yq�On�m��MØ'͑>�	�W�ƠA���xPL�G��dS����n:?�%�uͲ���4������ZX"�� /_�\�0Hk��2,�L�$�On���O��4���7˛��ʴb�B�߼���	eeO�=�z,��Dƻ�yyӾ��1��{}��g�T�lڝ�MC�O�<d����cN0n�豗�R�iƐ*ڴ�yR�'������?U�1[���S��q�J�Us�5�D�U�:���i��v�\�	֟���ϟH��П��`��z�]R��G�T�bQ�W)�?����?a�ih� �O���g�^�O<�QdG <���Y�JG�o��|���q��M�iT�dm��E1��2O����16G� &��@�Z2���H1I�ap,����=�?I�m6��<���?���?��Ȗ�*[V�s��@�<�QA��?	���DAӦţ�c����������O@i��6�@����{$~�I�Ot��'�z6��%zM<�'����]�a���K��L�6�4+��t��!ָ*&d$�.O��i��?��2��\�M� {�뙤K�H	�đ��n���O8���O���<!��iW`��� �Ȝ��a��k� ��KS����'5�6-2�	���d柌 ����M.-Z1�_�b[��(�LȦ�)ߴ$ T!:�4�y��''�%c�*��?)ۂP��A��_�М1��ǥd@J0�t�t�\�'���'$R�'5B�'^�L~(C��>�ē�@!
�	�4M2,8R(O�$+�	�OJ�l���I⡞������E��-=z`NݦUrٴ�yRP�b>�0ק�Ӧ��a�� �jT0gꌀ�N�>*���f��`�2��Ot�K>�*O�i�O>���C?	"*���Bf���4��O���S0V�&�˓i���'T]�D�'ERF��g�nIHd)�)&��P��۠vmY���	M~2�']���o�jt�'��iA�8#j�B����6qp�'�B"�1eXi0h�����埞�R��H����h�r4�g�q��e�P�i���D�O��$�OB��1�I��t��/Q��Nؔ~����d�-/v�p�S(^���sӸE飥�O���N���Iwy��y�D�V���'9t����)�y�lӐel���M+�D��M{�'��cǠP:��SV$��Z�b��w�l}����@�j�W�|�Z������`�I��(L�Va&U�	öJ Mt%�fyRs���(�<!����'�?��E�16�����'��i2����Jͻx���M�r�i}�d/ҧY$��#D_%&%JF咫n8�-�Q:eB���'�p�P���U�|"_� JR��)��TY%),\1h-��P�I���	ן�Sayb*�n�$�')�I(��L>aF&��T�Z�O^橊��'t�6(�I���d�O�7��O�|yE���G�X�0�ǐ.�������1�7�+?AG�
+XJ��4��5��-��I2B�3WP���"W�y"�'`�'x��'�"��
�o���St�ԥJc��d
:>��d�OT�$����c>	�I��M�N>i�ĉ�p��;s��h>��;�I�WJ�X�D�ٴQx���O���i����OJ%� ���G��Pm�18���W��8n�p�)��լ�Ozʓ�?!���?����>h�3**:�N�`KC9AX�����?)O�`mZ#�6���ȟ ��^�4�I�Eyd�g��ˢ�B�q��tyr�'N��'&��O��4�5�H�yg��M�69�1ŀq0R �"[�>��`X���ӌ#���r�	.B0�A:�"! <ԺU�F�|������I��i>A�	�^��9�'�:7m�&4G�X(��U%0:TK�ėvA.H���?�M>q����dG妥��!R,Wx�}Q���L<�1X�k���M���i ���iN�$�On�r��Ψ�ќ�4x&dڌ �����Yx�$肀l�ܔ'W��'Lb�'�b�'H��?��&���*&�Q���wlz�1�4<���p��?1���'�?Q��y׍A7��}@ ɖ�J5�L��睛&}6����I����4�R�)��حHGLӜ�IJ9ʐ)������e���6���	�R�LX0�'8�'�\�'�2�'o�A�sN���狴Mp��2���?����?)�����ڦ�8�mZ��D��ȟ�Rc��4���1IW��#"bl�ed�	��M;0�iON���>���B�j���đ�X#��@����<���NK��D �5���+O*�IW��?����O�-�@�ۈ<�*�a!�;>8�̻f��O����O����O£}�;eu|�����&EjP\�6��6\��8��0�&�C+K���'�6�&�i�Efl�&Htɨ I����ӂ�o� C�4<�֏a�l�� Ab���ԟ�b�mZ:/V��m1k�tԋc-��u�f]/��$&�x�'���'!�' r�'�\$Z� ����ju�\���Z����4OĬ���?a�����?�c,ҶY���H��� Yo� ��?*��I��M�¶i��<�	�j�����Ȁ�hHjNe@5�4{[J����L��5h:�P�W�'�%�\�'�n����i	�U8V��%Q�����'�2�'�����Y�ċ޴��t���]�d��FH�f��2@�s*e���6N�����[}b�`Ӿ�m)�A,h"2�Zp��5@��U��� +�*�l��<���$;d��"D�d�'A���h��[Pǉ�f����!��Eq�$�{����Ɵ�������I����%@&P��Ђ�Y�:%�[BB�5�?��?�³iü�O�xӪ�O�"��\<bs8�@�%.ff@0p�a���'��6-Ŧ��Z�Vhl��<�� ��1h��� `�r.�/~� �iN,*����䓏�4�p�d�Oz���n�|-�1�о#�ْchQ�qx����O�˓ƯvD�$j�r�'��X>�s���>2P�)�`�,W�`��.?�RP���ٴ*j���,�4�l���uoƍq��נe��,��D*�zH�<-��6��<��'E���d���eD>��N�-P��u�C>G�nq{���?!���?a�Ş��d]צB���<!U*�B�{��àׯT~B�'y�7M0�	���I*�i��;����ʯ�j��	��M�F�i,����i���5:���s�O輦�'E6���K�r�i�M�v.Კ'�����I���I�� ��L�4�X#*~H0HL�Q"m�1��)��7�ҔDHH���O���7���O�4oz�]� �Y�jR�.#b����5�Ms@�i���>�|�aǋ��Mۜ�� `Y��Uܸ˶&Cv�p�5Oh��s�Ⱥ�?�2�.�Ĩ<����?ABn 7Z�`Kٲ6�5��D�?i���?������Ц%{eH�ޟ�	ǟ�i�C�D��Dq�ˁ%l7F����	X�%��	�M�׼i��O��qFe�2u@-��A7D���Q�;O��$��hOn����[���S*7�F�������<�0���ִl��Pz1e�����I�(����`D��w�� ����
?d���cXIt�0��'(6��#�~��O]mZJ�Ӽ�a#ߙ;`6�G�0�Le,*���=�M��i=(7���r�|7�|���	J�6d�U�O��ۗ��X|�D�F��C��Ź�'�`�	Sy2���j������D-r�b��� !������dK�v�2�'g���̯V,4����\1��w�|�'^6�	Ҧ	����'������h���j\D��G��3DR�,б`��-�,O��s���?1��:�D�<A�J��'�d#7�M�W�@ ���q�<r�4Z�,[��+�T=0C�]�C(F�ڑl�8d~���'4���E}�iy���m��Mc�Ƅ�z�	r%�1%7h�� $o�~]�ݴ�y2�'�X�����?$^� ���u!��M3w<�*m�eN���mq�p��� ':����l&8��w��L��I������M����C�(��O��Z�ǘ9G����� iy�x��oX�,�'T7M֦I��i�>@o��<9��d���YS�׉\����` 	�B��Ϗ�# b����䓡��+���}Z�K�䟱T�\���P�^Q#<�C�i���c��'�r�'^哲D��X�R��25���8��[�n�@�uJ�I��MSѸiT��d)��T����Z$t��"��w��p�C@�T�vU��� �����!�O<�BI>i'�K���\�4�#y��q!RR<i��i�e�W�Z]���`��;��������z���'^
7M;�ɟ���Ŧ��b�";l\"�@�$i�X&�L�M��i�Z��Ҿi����O �HC���2�F�<AWGN����e��=|^\�OV�<�,O����O��$�OH���OF˧m�X��,_s7z�(�(P%�Q�W�i�hb@^����w�S��*����3��&D���I�/T�� �J�xF��kdӠ�	`}�O�T�'�f�ƺi�󄒍(���:FD�I�zP�F�]0��M�EF���
k��O@��|��
6ٹ�B�7˶Ej�!� Z	q��?���?	)O`�lZ�X� !�'��	=t�ĕ�$�AU��Z�"!	�O��'��7M��M����)G���RF�U'w~X�Rn�+0��O�u��['_ے��0������L�BcV�)�i@�4�TDA𬏩4�6���Hԟ,�Iޟ����E���'x6�Z��^�(���^�
<.ts@�'Ӓ7M�;Ov����O��n�w�Ӽ�+T�X7��`�i@���=8���<� �i�+P�?y�J���M��'������u�S�Z��Jǋ)�d<��'ܲ,���|�^���՟��I��I���o�U���I�t�Jw��GyROlӚ��k�<����'�?�a
�$ at�ᒅɎf��\H$�[�	��	�Mku�i��0�I�����a��ժt0KvĻӁ%��y��M�^4�	=�
h�S�'�h�%�d�'�(�
����w~�LQ�.��C�,���'�R�'����^���4.5ju0��]�d¥�L�2���5E*�����JʛF���z}�'yӔ�l� ��Z@�I��٬��z��øn�r�o��<��Z��t�������'���&c�Ei�j��*Z��'K��Lj����a�|��ǟh�	�4�IΟ���W�O�i ���NM�57� �cA�;����O��l�6d����z޴�?q)O�ͱ#�P�'�bU�7d�8	��x���'��7����]�� =l�<1�dst͙�i	�-�v0Y@�$���i�8!���d�䓠�4�����O���X�'�89Bm�c�yᇯW5]��D�O\ʓN̛��C@����ЖO��X9��δ.����9%�jp��O��'6b6-�ڦ�Γ��'�"�_��hq��+y�(1"�D��]1`����԰[qʵ�'�����4k1�|B���8]ڹ�C�!��i�fe0O��',��'J��$]���41O��;p�~���f�:_$͛Q���?��v���'2�'߬�I0���L'gD���ȓL�V0�1�8Z��6��O*��s*f�~�	㟤q*
!E�D�'?����.�!�@ˋ@�� g	��<�(O ���O����O�$�O�˧!�f�3J7p�����T�>��i+Rm�&�Ѣ���'B�$�O���'H`7=��!p$_4�`�'$=
N�ɐ�ܦe��4ٛ�'�>�'����$�M��4�y�R�x�r���$5�l��oӭ�yb,4qh�Iy��_�̕����'� T��A���p  �|[Hժ��'���'�\ :�W���ش`�Z<��'�?���c�e{���9���⯋=��|)���$�O�w��&vӜ�o����D7a\��Ajg�p�(��Y46����O�1�u�[�v��D������4��&��� �I
3y*�Jf��)Wf% E֟�	��4�	֟�$?���)O���-�	! �:s�	.L1x��&��5n��I'�M�'	F/�?Y��?����4��(���X �A�"���Q�II�6���ɦ	��4Zx��逓Q��0OZ�d^��P��'��p�)�!���*5m���а+�d�<�'�?A��?���?yQ
N8z$![�lY%`�L
Eo����d����������	؟�ӺO�������1T	H�d�|Y+��.�Z����X~�'���j��&>����?2�.� 8cd�B%p*� � &7h�IC6P1I��	 n�*ӆ�'�j]$��'�^ח�	4D@9�M��d��ܘ��[���	ݟ,��4V@�	Dy�zӶd����O(���.��X
4ሂs�m����O�m�ڟ�'��b�>1��ia<7MS����B�^Z(�pcE�<9-�F�')Vn��<Q���$(�r���8��'�$�k��������};dj^9C����0/t������ڟ�	�����Q3(t,��E�5IR�M�,@%p@�Ȑ���?��i��$^�x��4�?�(O�7��)rr�5��6����ڦ���O��n���M�'��9�4�y��'z�X
�h�I���R��(ԥx�ϟ&E����	-E��'��i>!�	����ɹmo�h ��O(HZ|�;�b�!q�28 	ڟ,�'��7�P47N��$�O��d����8CVr�jT�Xj,\Պ��	�d�O������|�h�n7�ħ���H�.B�V���储b���Ad;T���ds	� $?	�'DI��B��MI��RկD�Bv�p�t��+E�K���?���?Y��|R��2�2�C.OvAm��ޅ�>����ܚI�"]�c��[��(�'p�|��'{剿�MV�Q!�r�
P��2���h�*YQ��~�,��js���	������
f���./?1��6}�r�����*V(��Y!@��<�/OZ�D�O��$�O����Oʧf^�{��=&��i�O� �hw�i�Q��'R�'����Ȑl��'��w�lUBQ��$ 2m� ��%&��Iv�J�l��M�A_���?=��kE|n��<�����-k3��*v�M2�N�<i�-S�#����ߤ�䓢�4��l�� �H�?g�N�Aq焴B�����OT��B�k�ʓ[�&��3x����'����%^�a�5E�u,9x#'·SS�Q�`��Jy��~Ӧ9nڅ�M[Q��i���=|�	!f�(`���#?YB�6@5����f�'U=��ߦ�?Y7?s]Сz�
�M�B���I�"�?y��?����?N~�`Ƌ�|B�&7�$����+c�~�e� "@���,��蕯^���'�'��i>�]�Tv�-����q2Zmڦ6�.���M�f�i��7M_6#�T6M,?餍S�5d\�	M8�`8�AI�q��1@JE;2���yI>Q-O��O��d�O����Ot90W���`��7��?`�N%aG�<�4�i��PR�'���'��D��%���'K�dU4u�(Rv,�g�B��Rh�>�3�i��7�Ȧ�J|B���"�IJ WV^�8��ɤ	���C�ͳ���R`%Vi~b���f"ȱ�ɫR�'#��!90�1����$Qz�YE낶s�\���՟��ӟ��i>��'nd7�M�
�� �\�B0�\6& s!��
�馑�	x�I���Ȧ��4 O�f$�<���%,��X��(@B��&t2�(��i0��O�H�����3k�<Q����Å�R/.s5&�4����<)���?���?��?����oЂsƅS6�� <*p�c�R�'R�a��M@q<���D
����yy�����;%F�6@vX�É	k�O��l�7�M��,��#޴�y�'g�a�!!&[ϔ��g�d�4����9P0h\�	�?9�'1�	Ο����\��	D�
���"�?:���PA��#q�	П�'�d6��Z����Ot�Ĳ|b�I9H��̰%!��}��ɆD~r�>у�i�6��p�i>5��p�6I	dK�-Gb�&��g?�	g.�m�ZDp4AVay��O=���IY��'0�HbҊ� J� �핆Dp@p�'���'�����O��	�MSw��._��$]�/.JB� ЁQ�������?��i�"�|2ť<��4|fpyK��5`�m���\� "d��&�iV6�8|6M}���I�o��(#�O�� �'	9Z�灧 �Q��� �~��'|�۟�	͟`�Iϟ(�	f�4m��Cyܬ��HU'D�f�	�e���7-�����O��D:���O�,mz���F�?�H$����qN|(���8�M뷷itO1�<$��v�,��8�a���c/؄b�Љ��	�
�ZU�'��%�P�'f��'}� ����ҥ�8]���2�'���'|"V� *ش�l�+O���8-�y�dcPri+'ї:B��@�BE�>��i6M�v� Y��E�A� q��9!a"%�:�IП���E��r<��P2��py��O����I#��ԃZ�>������5@�ەK��'Y��'br�S۟x��')'�,]�b��^g��ÑD���ڴk%�H����?��i��O�Ζ03���5$F�e�D��dU<8��˦�Jܴ.����E��6O���LO���'<꘥�T��%�Q�ʴ|<��FI߷t�69argй,	zk���b��-�W�0[nMk�#��h����Kعh��|:��Ʌ}�b�p���J~L<x3�ø-�p�yd�a $�	�FǄ9��{�Q����GÕTB:԰�HE57�<�����P:�<y��?7�Vԣ��
�Dy��N~o֨�#�F:d� ��Q�A��A6�5#�t���zqR��7SHh�9� ��+'
u��)Ѡ��F��u��#S 4���@я�!���F"��?Z��B*�@���e��rI>�*0���Ț`�
V%D��TC�6]pT�w�i*��'�"�O��Uo�Y�d�	+
f8C�	�#' �o����	��#<�~ī#�%����
	8���v��}�D�M����?�����x�O^�!�P#�΁E�NC�e"w`u�,���'���y��'��Y��^�j�&��A��n�Bu�0���O���H2b�&������Sf��n]+t�*M:TX!2`j��'���1$�b���IʟL���S�Y�3�T~�4�O�!����ݴ�?ae%Ϟ������'&ɧu׌C�.�m9�AF &B��1��ѱ1O���OR�D�<�3j�]���iTΐ�f.R��$��)&�h�ҞxB�'�'��I�0�I�׀ 0�����B�Ru��?I"�}@ciQ��?���?!,O�p��P�|�p�x�>�Z��F�A&\`��[}��'vB�|�Q����>D됍b�TYу�p�,q��*S}��'@��'p�	�U,x��I|*d�H1{����so�=�����
�kH�f�'z�'��	*K:c?)مM�;[Y�Z����x���S�ad�����O4�rݚ肑����'t�\c����i� %d�<(4h�4`�K<q(ONt�c�^ҁFE39��a��	;���·Ӧ��'U���e��8�O|b�O�X�W%��
��׸P9�]p�`� mZ|y2뗄���?'?7�\�WQ
M�E�ެ.�I1�(�*;��F� )a.6m�ON���O��)E�i>�"o�aur�)�ՙbw6T�$dʳ�Mq�Ku~BY��$?�	���FK�<3nH��  ;Z�P,
� 4�M����?q�����x�O[��O��*�D�B5F��B7hlt,��V��'78i0�y��'yB�'$����Q��<��f��#�v�`��jӒ�d�<�<5$���ڟt&��ݯj}<%���W��6���EA�e���\��<����?a����!��\3�?l<=�P�IaҢ�i��O����O0�O��('z�Ad�A�,��b�TZ�Ty�C̓�?Y��?�*O��H@���|±�M�f<9��$L�� #�o}�'WB�|S�h�ã>)�d	���yc_8.uV�b��O}b�'��S�(�I&b�OF҄@�}=��	`A+,R�:e�]�j�r6��O"�t�	��v���+��"[d<�C�=s� 	��Ԅo,��'v�	��� �k�m���'�O��0�4�7\��I��/P�^I�����8�	ҟ�3%��#�b��'�R��+�,P�p�R(�=-/p1�'��%_B�"�' 2�'v�T[��]56�H��LB5�n9��ʗ�@ *��?Q�ޗ(Ab��<�~�bj�%sF� �]5R�|���]ަ5S������֟��I�?5�����'�,-X��P>2�Rd��U0&"=��o��E�@�531O>��ɐC����"h�(o8#��K��L�۴�?I��?)����4�����O���Ggl,��$Q&G¤J����*sn���yBG1���H��OX�I�X����E���h�$" �b� D��,O�D�OB��1��=A��\�ԻR��� �ʌ�d�"�?��I[���_~��'8�T�h�I��n%Y��:��0�L�]Z��)��Vy2�'Fb�'H�O.�dБ� �� i�j)��){3&���#.!�	ɟP��VyB�'`�\�!џ`�z�G)k�z�M��#jd���if�'nr���O`d�P㐿'J��B�66H>�����afx@Z�(����O4���<������*�R��Yz�OA!;���#��t���n��h�?���z?��1�Q[�I�RtA���^�o��H�ύ)^J7��OTʓ�?��i����	�O��⟄�
tK�:�Rtր�3� iі.�d��?�p+R�*ұ�<�O�~d��g��	&�"�Y!��mɨO>��b�X���O��$�O����<�;9�.����X7���DP17�p��'�bK@	}tD"�y��$%P�%YH)�L=F%J :��M�0bF	�?����?i���(O���O�-	&aX��A�4�L�z��P�J������7b�b�"|���J��I��A�ԉa�e.{PU�i�b�'h�m�+j��i>������x�p�� ��]��:f�M�*���z�	��ħ�?��~���:l�L=Hq�Z'~�ELO��MC���Pc,O0�d�O���3�	�F��eZ�G��+�`�@Հo�O Ż6�����ɟ��'B�A$v��jة+<
�[�NO�-��IrV���������]���~2�%�ҹ��#s�Z��s����M[U��E~�' �Y�4�ɋ��}��U�@�q#���L�HIVnQ"�lZʟ����?1�;F@mq��
ަ�pD�0zD��A��J.T���B�>Y���?+O����
i��'�?	"	
0uo>��fdS.��Q��=F���'�O���4p[n�Bטx"hO&.���[�v������M������O��B���|���?���L�\��ԋ)��x�(~E�9�����O�p�Ae��-�1O��=��u�R�H�_H��q��,MrV��?9����?1���?9����.O��ZI���"7��<]��!�$�&q��I���8�˙N��b�b?�B��H=P0��*��M�ZI��iuӶ�� I�O2�$�O0�d����|��M����a<yk�Љ�lI&<�(�"�i`�sրR�Ř����$�Z����^�N�V�R%��0O((nZ���Iʟ����IAy�O*�'�$�P�ly�UV�?�R4R��>o��<��ڦ�OSB�'�dU7`*0��A��X�Bx2��=��I�~΁�'r��'�DW�6���[�/cb���\5���B�"���??��?	/Or���x;��q�M��'��d:!�B�#�aR���<����?A����'��懖���#��#.T�,�q"I�[Z�Q�@�V���$�O,��<���7un���O�X{Q F8_�>�`Ҁ��H�A"ش�?)��?��2�'��-��f_��M3�h�8<M�HZgHM$)�h�
t}��'2BQ�H��
W���OY��[�s�օ�Eh�Y�<uK �|��f�'��O���~9���x
� p݃7�B�>j�b'S�n�p����i��S�p�	&	��ŗO[�	�?�#L֗[��1�L�:"y�$煀��'l4o�����y���l�A�M��c�����%wU���Ɉ|7�a�I���Iʟ�SByZw>�����/.8�TY��*[�(J�O|��cz�\#����_�>�q A�>�l}��.N,6�&IN�2��'���'2�P��S۟L�@�˿[�X�:�F3����B���M{�cE�r�7�)�'�?�u�	�x�`��'�h{����^����'�r�'��k�Z��S��D�	o?y��_�bAH��!�#jY" YG�Dh1O$�QB�d�ß ��e?�����:���ЋX�;�D���%��)�IAyxU�'���'R�M�T�!Okn4��_1T�cX��0MS�xt��?������O�l�똲`��!s�\4^zȹ·�L����?���?1�b�'�b�/˭t� -���?i�$m�&M�{L!��O6���O�ʓ�?�����4�
Y�.D9D$�8b�� �����M��?����'��B[�UUq�ܴ:�DK����p|�#FT ��'��'���ȟ�c��WN���'$�](�(�p�R�b6�)Q��$;v�y���d1�	��4s�i@[�O�9`iڬYEP����^b�\y"־iE^��ɊB��	�OZ�'��4��6�
4��(�8�.%��S�d�b� �ɪ ���'4�~:P�X�	^�Rq.��8�p:d��G}��'�$݁P�'��')��Od�i����Ё\>2e3cAS2.��C�>��R�4h��`�S�'Ov�"��Z��Jɟ�6�6�o;L"b]��Ο������qy�O�R��(�БB�!׹)CJ�b���-a��7�"��#gk�S�O�]�=n�	"s�M,kGR���$�ͪ7�O����O�����<�'�?1��~�J�8����Wl�7J��h�ŌH:TJc�<�AD���ħ�?9���~��X�8((I�@�F�re+P&�(�M��uy`.OT���O��;�ɯ_�dŋ�*8�T1�sᛑaN��L�QYPe�c~��'��'��|�rY���$q�PN׊x�Z���;��Ħ<������OT�d�O���-[Fp 3����e�h�*�;D�1O��d�O��$�<i��\����'H5\mP�]�v0\@гlد|ڛ�Y�0�IZy��'+��'��Xq�'�j��%/4l���N�/�0\�k~�����O����O`�^|��#T?��i���Po�"[��)�I�1��cЮ{�(��<���?���$�hqΓ��i�|H ��2&��
�l��6|��޴�?a����%Z?��O���'h�$�Љ!������H*X
�0�Y����������z�x"<)�OĔ���oM�'��p��e�+o��ݴ��*�to�ğ��	���S&�����]J&�� Pp|H4�Iv��+c�i�R�'�����'b�\�(�}R�%�&*���� ',Y��6i�즁�6���M���?�����[��'i6QA�[�&��YhF�_�Jn��rio��񗒟��''�\��7[���J1��7��]�E��9��mٟ8����4hu期��ĸ<a���~��W�S��L��+x� ���ϵ��D�<)T��R~�O���'��ԓ\@}j�(k��Ax��ФL�7��O�l�b�v}BT���RyR��5&�/_L��V��`U]	��G��M�Q�P ͓����O��O�ʓ�n=b)�L��j��"-_2y���3\��Iyy��'��	��l������D�<s�����2��i!��}���	Py2�'2b�'A�4H��˟Ok�5�C˞�RH��&�q@ڴ��d�Ob��?���?�!�	�<1D�dw�����,T\tu���ѵJ3��4�	͟P�	��Z&F��M���?v	?�L�)�k�8��Xh����&���'���'��ޟ�T+z>E�	B?abaO��I��	��Ͱ+��=���0�'�m�0I�~"���?���5�]�a4z�V���K� ��xtX����� ͓���Iy��'��	χ<�@�#�k�� H& m��W��� ���M��?	���R'_��]�n>�}�جJ
�HI��^ @���n�ϟ��I#e``�ɺ��9O��>���X>�e��$���@�C4�rӔ̫����=�I�����?u��Od˓M��=���Ү���s0!�,|�h#�iB�%!�'	�'���:9[�����(@#�O�e2�%n�ҟ4�I�T:�iF����<���~�C$E$y�į��r���`�Y��M�L>IP&@�<�O{�'-IQ50�؉j6g�!D�]�t�>ǌ7�O6%� ��t}�\����ky���5��P�@p!O�h��B������ ��<���?������g|���G vT�ㄨG���0�b��_}"R�@�Iuy2�'<�'``�S��2vL>���,Q�x�r��Ǐ��y��'���'^�X>牖9,�@�OEp�9TD-$�� ��?]Y�K�4��$�O�˓�?���?��L��<�s�ɉB�*��$���o��0����Tc�F�'���'q�Z�d@��ȍ��	�Ok�ΎH$ b��&�4%�1LF��'?�I�d�I��(�T�c����f?!��	H.�*�4.�YQ$�Ѧm�I̟�'l��d�~r���?��'Dp+w:mH�2���TlPST��	ן�I18�����$�?�ñ�КH/��ɔjq*hf�T˓��f�i�"�'.��O+j�Ӻ��_Nh�L����(��A�g����	՟��@{������*�3� $P!��7]��g�NWbABf�i�,\��'bӤ���O����
I�'��	.rn���Ar��a��^�%%�8�ش d%͓�䓞�O7�����Q��/	�L���1�76"6��O��D�O�yZT��D}�_�d�Iw?�^�Nً�!�;s�����'�8���k��?���?��#��5r3�)�2.G.(�	]ś��'.�SF��>a(O���<i����F�p��:Kұ
�8jE�Pn}"��y��'���'Y��'�	���ADDY�`�mb�NG>c�b�;�����<	����$�O���O�b ��+>d= 1T cO4����D�X/�d�<���?�L~�@��g��i�O��6��_R�5���Q�x��Ty��'���'�͒�'�T ��s�X#���V<���&s� �d�O����O��H��WS?��i����m��G2AJ>0L��t�o�z���<���?���9�D�̓��i�#�N��O��%eF;f���c���$�O�WT"�z�Z?)��Ο�ӭWT����ϙN}n8k��g�z�I�O����O
�$�\����O����O���'{��x�`�^9[���@c�W��
7�<Q2lNm��檰~���ћ����ƕv���k�NĈ�xT�i����O�Вp:O�O~�>�����&6:bꂨqd��F�g��);�D�¦i�	ß��I�?�I�}B�5SO���FJfV��G�Ȕ~�(7��{��8�2��8zb� ���'k���i���'�����b۸O��D�O����H��.E�:�R��wl�6M=��ߔW���%>-���L�I�d� �h�%ޚ/.Ra[����#�>�x�4�?n*��O�$&��ƴ�����*hD�閇[0J�Q4V��1v'd�̔'��'�"S���F�IT%�N�2e�,��7 6��L<q���?�/Ox���Ox���-LQ������2A8f�;�hI�W�� ZR1O��?q��?Q,OF�����|
6#;�8���6ΦyЄ]��ɟ'����ɟ�k�ì>�d!@
�P�g�Q3z&mQ��~}��'��'|�?)���qN|*�G�:\jL�ȫ��S�-�F�'r�'9R�'�L�C��+t@����.ƾx��	 �$^0D�v�'c_��f���ħ�?�'|@Z�a�&S��r��6FV���x��''��!�yr�|՟B��閒4К4 �'96����i��I5�:���4"\�ڟ��S����}wf��ר
:jL�u��T�`����'���O��'�~��&�41X0�	i�����

�M��L�&j���'���'��b!��&�i��5^�D����߰@5L 8۴j�H������O���-�6�	`�B9���A�)s�6��OD��O$z!eQS��?��'���+���#P���X�L�:-H�}�c�H
�'%2�'5��)���:��sZ^	�Ӭ�a\�6��O�tNk��`��l�i�Y��G�^�P ����4B<ҡ�<6Mi�Ĕ'(2�'_S�j�/M|P����M6b(>���n��p�XP�L<����hOT����6dLI�ͅ�]�Ȃ$��Ӟ���O��D�OR��O����|2�Ŏ��?I3EށJ~�̂��ˇ��ѫ镎sn���'�"�'��'�2�'����O:}�t"n�%�^�s�I�
� _��� �	���	�HA1�D�D�'�Nb��D�}��B`R6Er�qb�jӚ��2���O��D$D��1Q�xr�	 f��	8��G�s�>���ꐩ�M����?a/O�����s���'���O���pR��=H��u���VB��;֡w���E��B���1U�Y����_��zS,Æ".P|nZݟ<��GH�!�	��Iß\��֟$�i�y�dX�����R�Ͻ�Nȹ�fn����O��P��FH1O��&�s�FR7-���j�&@�o������iϪ���'���'�r�OhB�'�品7܎%A�+�D��&ߌt���40�&�k�S�Ox��+
J�PQOC2w|�j��C�G�f7m�O��d�Od#� l}B_>!��ɟ�(�Ǯy���3�� F��Q�֣��'NV�(p�|��'j��'�晈��N�`\�C�� $z�P
vӴ���baLʓP������$�`��+O���<�f�X~@,���`�(��D�8������(��ܟ̖'�E�cΦm"����	l8����L
388U8��']r�'V��'��'W��' x�X�jF�j�\ Z�fձ*R۔�Q�cP�iS�OL�d�O*��<�Eo�� ��	�?o�1�qD�L�|��f↻k�'��|"�'�r�ȉ���ʣ-[j����.f�����6�I�|��ܟ��'x���E�1��˖Ybj���A��M��.=�x�o��'���I�����?���?�vQ'O�@[F&��&�6��O`�ĩ<���:��O`��O�E��,\�6��V�,/"���*>��OF�d(����'H�P���=KJ�2�2Y'TnZ�\��
P`������	�(��UyZc�x�:�.�+��$!%+�`w$=��4�?���`ՊYGx��	Z� �>I����c�0���фH�BL��Eg���Ն!|OԊ�	HK�����D�<����U"ON�� "H#�Q4�\+����փxQb�OO���pNT�@] ͨ�(\�����[%�l���Ӊ.�%*�M0O�T�I�#��q�!�R�X�̱�3%M +���Z#���D�jDO$g���#J	�9������W�L�� H�2w��Uz<�v�A�B��a��ƈ�i0kV��Oh�D�O�������?џO��8�p/��ה0�2��\iT���:�b��C+B45��@ՠ*5"?�m�6c�D��5d[�[Y$�svA�)�nD�V,�RF|�)Uc�T���2Aˊ�R��(��b��Q��#5�ؽp#���Fhܼhr��Q`�[bh<�u�Q�q=��u3!	B��P��M�<��䌦
�<�04E�/Zt���eB̓%��IFy�,�)vN���?I���*4@ּq�(9R`�3[?�?�����?a�Ol��iŠ4 Ⱥ�+W?q��R�]`T�D���&�1W O��p<�K\0�:���d��I�ߴS,.]#�j�>:/"Q�`䂑?���	+�����O:ʓj~A���� ��EI��Q��]�<yߓG�,�`���L}�� S�]�u��l��|��&b���48�GK�Y���`a��yB[��BĄ��D�OR�'[�~\��O�-Q�Lրo&�� >r?� ��?yV�6o.aS�E�`vV� ����|�į��D"*u�p�ӝO�=;'��u��޼~@�z��\O�:��r�(ҧ�rp�S��2B(8�ɞ�m\���O�\p�'���ǟ��D��>+��t��֤V|��J�!#D�Њ�#ν5���!E��?��t��f OPFz�fB.X��!�D�l��W�ܛil&듎?Y��;\hKv�	,�?I��?y�Ӽ��X�k��	�'gU�({�q���ǻ|��U�5��
J���xF�<���L>���Ϧw9�GW {�|iH@j��~<�L�b�ܙJt��N�0�l,�}r��eU\�I;^�2�)*1xA F���|��R~� ��?�'�hOb5	����O�p��F ��F ""O&�Q��<hhꓥ��ٜtbǐ��+���?Y�'�л����PTa���]Q5���ڪ[j�$9�'��'���m�E��ͧCĆ1 ҈�J�,%��j8y�pXW�I��ȡ���k�$8�ϓ=� j�f��M\���M�lqU�H QV �Ǉ�����`�b�G|R����Ed�:N�(m
���"���� ���`��j�'��O@��v�H0��p`��9p��	0C"O.����F�1��m����/�n����$r}�X�,�N?��d�O�[P�̦��x�
ܡ$�� ���O��$(Y����O���2'�`<���S�4�B���'N8b��ڶOjά��'�T�0��B��@P��K��%K��O�({��!0�T�p�C������'��lP��?/O��H7o�Έ8�W5>L\V�d7|OUb�#Պ^����%D�!;I8I�aO�m�&E0��*�V�À� Nc�	fy�
:7��OR���|�&�R��?aĉ!�t���@+a�@�����?�Q��0kӰi>1O�3?9���	�2M��k P
Es��Vq�߃pex��?�!4��l�����FL�A'���)1}��?I��i�
7��O��?�Eaڽ�t��3V��m��!=�	�����I=[��xӦ&Xx[�}q�=8N���$DI�'_",��X�,��pgBN�#6��*�b�"�$�O�̛M�r����Ot���O��$��dD[���k� 3KR>�����*�	����i&��@.�-K�@�}YB��k8vB�#�y��Z�1�X�}&���g� ���V�����M��i7��$E{��,O��$Z�z�&/z�B�%9l�C�IOt������|f�  _�DW��>�HON�'����:4$��v��=y��9A�.F$/=��3ugD3��d�O��$�O6��;�?����JN\�b2dD Z��!��: �Lp�R�'f�h��CG�ƴ
`@TT*�3ƋH�iT�rG�_�Z��E�Ν`��aqGPI��b��?IO>Q��?ُR�'YDmR`c^1Q���.�0��\$���HC1G�����0-t��<y"[���'r
�`d�>1��+B��ɰ�A+=l�Uie���d�. ����?Q lE��?!������ͷ2���y��U�ʤh�� ��LS���jH�H)�H�Y2��8�����t�� G�:EF�Q�`%=�p��#U�%3�t�TcW��t-���
T�'������q��&.�>ae��$B.�0�c	� M�B� A̓�?	�|�9�gԞY X�I� ��R�B݇������ a􋐥5�z�ˤ����y��d�>�}�'�p]+�-��yV���ũY<P����'�2%�ac�>bY��Ia�1�
�'����q���y�
�>�de��'H��!�.��8Z��<'t��	�'� �ӳn\?�zY��C��"��m��'��e�&(i��:c$�*��C��� �Y�'ܡ�V��:��hD"O���e��W�l��@�JM^6��"O ����!+aBe�0�Q�	��di�"O��*w$G�4�i1�b�)�"O��zq ��K+�����TJ|���"O�p��T�e�^�6�I�yX]�"OJP�b/D���Gc�\	r���"O�MP��V��E҃Z�x����.D�<�SDI�[��I�lZ[e���h(D��Sr�4e�� %W�b�y�v/(D�\jc�у-2�Y:��զuoҐ؁f%D���w&G.o�:�zqi0[:��#*6D��Q�@ҫJ�q3�a�^lٗ�1D�H��ԆS�Ex2W(y���p �$D�Hkv*���%�Ժ01��p5D�HR�`�"?�P	���T�P~� c��&D��� ��n�����<\r0`a�&D��:�(����- ���;<�h`b��#D��g�I�O^�\ɠ��I?4�c� "D��b	��n�HY"r,�	@2���?D�HAf#�Z Ld���$!-�xDE1D���L
�I݀�v,]N� e��"0D������k�`�2⧇�S�q�O)D��0 ��=;�X�Ch9"����3&D�Hb���/�%�B��Q� %D�p8.C�9
x����!<� l�d7D�`0�
V�����5I�����'D��Ε�BM�`��fʍ�Z��o)D���r��G@rhn�)(\.��P�%�O�q�PSw�*�Q 7%ZA㒇�&l����&��S��sU�n��@h�n�-L�r;	� $~8e�ւ�z'��)F8Dx�)�(g���v"҆}��z�B^�ҍr��@�<��5�,���r��-C x�������BMI jLDI��D\p���΀�pT���H��;�D�Rp-��	A�iT���tc���M��y7 [�]�4m�v�>$
M� �ɱ�y�@�PO��B��X����`Z����
�'8��WJ�-- 6t[�O���@���!<%4��X�(�eÛ(�ZDBϽ6��q�7;�O�;a�ʞ��g�$p,�`��7�<��Se��<�a����f�9w�R={��)���/��f�<ڕoP9xr������Fx�+�E�0;2'ǒ�`�q�N�_7"q�U��C1�!Z����F�
��U /r�:+����	O�JF��gÕwӺ�
ϗL���l��5��}:��R� 8l��$	N�NV�Y�oӵ7S�sޭ�
ԚxQ�ܪ�|͋u�2D�4�3�����+�@g'���4$\9Ha���я2�T�q�&�(�B��]b�h3L=�r�'�����)�\s�aP.���OS���^q#���8��bS�\?:��8� K�g�ZQ��IRm���ˏ1��y"����Ox}IW`��zq!���Z�r��ɶ.\����شC�J�� N 1C9�Lyd��+�T)��^O�i9&����x���K�Bx����?�\��m��K���2��w�P�q�ą!Hf���?L���9��=�L9�Bm��p����y��4=�$��d�;^Kt`R�IP4�yB׆C�(pZ�M��<�Da�T�F��dMx$��d؊UNj��K�OZ(qX�A��\e�`�RW����C�O�����U
6�H���m'�OR��A*�=�@��'�=+,��*ˆ
D ��(��@�+Ȯu�Z�mS%b�PB��M �I�I��H<���).�
``��D�D�A�#<�2��8�h@��ڶ# ��1���i}B�()z" ��l(fr(�W�
<���/Ry"L1X�:b�b>�Po?U���v�
;L��Dk)Auv�Q!��?w�-���L�4&�_^n@Z��~Zc�}���D�����0�/Fb"�ˤ�;���L�"#|�'�,!�U-�w|����T�h������ē�B�sqW�Ժ�˞G}6�	�Ӽ�k,~�f����n����.�F��'\�x�%,+�l��Q�zuf!Ad�E,B,���%ơ�M�GW�`�l�Q�����i�f C��T��O6$
DM#M���j��E)�����I3�PlJ�
�,�I'R�W0�a�$�V�hR5���r�	�Q�LA�cE��0����E$���&<��er�I��"��h��$m�.��dp�A��bd�i�	-�|��Y���R$��f��|jԩS?$��{�	�,M�ONE�!�3?��	P#[2E�C�
�/���2�� 4�=�@�<���5t��8�a��y'��NE�EQ�OP9� �[���/6�(�Ԥ:<O �Y���vj(�� ����ɻ ��р�Pk����4��?��	ͬxQ�C��|b�&�-�$�aP�x2M�"az2|�JI9*'���󦏤�0>9���w�$욢E��qN<(�.��;�J�0ǡBZ�3�ԣh"����D�Ik`=z��d���ӵ`[����/W��@������z� "<P�+A�I9Q�O��N�Ha�{~��M��cD�K9F��0���Ť/X�0�`�9�䚉MW�E~b�B�z]�@�u�7����&���*ūӍ���r�ɪk��ٍ��ywC@6]@)���/[�	˄��3?D�P5�O�@�EG� �,��M׽tPu��4����;`S,��Eǝ4�Pt�2O�-jѠGc+���+�zʅ�BOZ5z5	����@`��
u�0�2��]?a4g"�T�Y�aΰ)N�D�f�'q�T��j�Iu�E�#��if�(˓a�)�BO·YR�!�U&޹J>����I�%<�� ��_\��Lɋ9>��XF�#�OL9�w�A�1`��E��5o`F�T�x�'+^�� ��	Gv�9�6���T>��u(�d�P" V! �t�d =D��iCmΚx�t8;�iׄ&TY��չvT歋CB��#vLdZ�b?����˼�c�A�� �WY�x,B�XU��H�<9��@�F���є疦.��1�g�ʿ3z�m��}���Ѝ�qLX��O&"=)�@F�5��dx���~�T�#���Z8�P5���
$��m b8�&Ə#+V�Ѩ�͓ \ P$�iR��s`�:�O��;r�K?7:�be���Eښ�� �'Z���<Oz!ň�t'@��U�$l���`"O
hbBA��Qi�'-ހW�(��I!�(#~��F�#dl�AR/,0ek"o�m�<1���R�d��E��k<�Q&	��<i�@�������	�tk�>x�0Q*��!]jqB�"O��zЌ�@�Y�kN�KBҀ
2����b+�^���J�GA��d��@CT��fh	�2�O�$��I�O�p���ؽ>��H�o_�f�&L��"OxsŢ�2g���*���:��3S$*	3���#%���?��S� $\Y8U���E�|��4D��������U6�|Z�"�	K��d�`9l���RǬ����V�I���W�dE>�"~BÊ'%�&٘�B�Kl�Qe(�|̓ C|��(�>0��QF��Ō �`,����U�qX�o��yR+>4|���'J�D��SN�(��A�aC¥�����3X>�:��
�`LG֊��%��qr�؄�TuR#���k���htH�
�* �'4�
�f��N��Y#G�B!s�iѕI�
@�B�8LO���4�˦S�Ta�<OL�`�b�)w�>=�&鐶��4�B"O�%�f�ٵk��Mɂ�G�n@���F�jP�S�Y�o?Q g��,��qGI>/�9�)#D�Pa�J������Ó!ɜLx�  b��Ѫ,?�pb B����d��pD)�78 �����F�!�$X�|�J� ���,���7Ւ���Et�^����'	v�kԏ�?;��d��JΰS:�*ӓty�e�gَ-�@5ϓP��!�NG�9h���r�
fj�d�ȓ}����p�thSl��Ҝ��<)�l�� ڌ�g�YI�OR���K���Ռ֬{��6IK�X\1O��)��3?��'�^�2H ©W&U ��Aa��w\��,�F~���6�����dq�%Z�`U-]������g�
��\�<��0�'>x�M@	9��qQBk�;"��ӓH��5͜K~B+R�p\�a#E���R��g��;�yBo��9��
%JF�Z��E�'�1�D�p|J0#OɁì�+>[�W��y��=r(Hْ1��(
\�E����{���c�yr�����I?4-j�K��Os+j�R���'i�iy�`�� 820I"oV0y�~EK��s��J
�M�*ը�M"Tz��`9P�j��hO�ĄK�b�O&-��A͑y�����U\��Q��"O$$�db�qX�|���K�p�V �R��J�t�F ���O�\�	�)͌#A����)a��x
�'Ƣhzծ�:5��@G��W�����,��Ә'�����𙟘�%�$$q0�8p!�d,�H:D�@J���y�z��Ċ�}VB�:qF�0&0��g�&�OԀ�g�A4x�H�HL3s����"O� �p�"����P�V�E
�@DR�"O��#� ����r��\��@�"O���KM�.��ܢ�(Q�*m����x��P�T]�82�c��ȟ�P`�܆5�p����
=4�1qq"O��RR��&��M
R��7T�=)�
(!��P�'g�;��$�3�$�7Rr��GIMv9�Qr�#r!��?T���5w�����k�z)���*ٰy3׹i�ўb>ݡ����GȰqjҏZ N��p�v�&,O�A�T���
9��]�\j����s���h��#D� s���#\�¹X"�(y���j!�D�U�����!� d��?����@�a����|��U�V�!�d�P:&l���T53d��E�� ;QJ%c�T~B���E6fb?OҼ1d�"�,yY�9N֡kO����N��2���Dt��"O���t�[#�a}�iҴ'������ܼ.�R�Yb��"�<i��Ի}Uh��3�Ga}���\��ҡ���A���yrZ��lr��4��I@'
��y�Ty��C��p7�!0�& �n��ȓ8-�|��b]hl��[ӭD�w�
i�ȓV����T�CAV�0a��Q���X�ȓ.�X\i#�B���U�A��(��I#Dxc�ֺ����@�ESa��~}�h�b<�ܔr@��)H%���ȓg����7���)�&!
@�L</؞Յ�]i� ���gxL�)������k_ h�1퉄/�Z�!%-�99`��J�V$��'�
4_8�ɇ̋?�LU�ȓJ�m���ԓ���9���u��ч�c��9&�U5a���C$�V̇�$�,��Uʚ�}��-��������ȓI��`aS!�,��pR�݋p����'�N�Ό�)s(ɽ).̈́�Q�8�8�*I)|�����I������B�`t����P��ıP%<���a༵�w�CDS��k�����@��ȓְ�$Nf���6��ZU�8�ȓt��,�V��:hU���Hά2�C剠;�Jx�ï�yE��gΓ[mB�I4�x4�$\�>��P(B�P:`����lL(qQ�V-(���`&B�!�B�B$<�k�ʕ�[�j����$!�$]%E@v�I�Mݽf`�Z�O��nZ!�d�k�*P�O�V��2�	o�!�$D�R��Ν�|Ru���޺8,!�w�u�S�]?�{E)w!��!�J�y�hE�R���c�J�>X!�d֠;(d����2/|��'�3�!�\*�\E8G	��N
@���i<!�Ć�"b<k�#����)�A+&A"!�dQ�t�-�!يxЁ`P	F�!�є4�%3��
)�,a[�j�#zo!�dӼh����-@0�����i�3X!��5>~��I��xzh�yq��9K!�$�&�N(�� -��칱�45.!�d��8���E  �U�J�fG�'"!�DD#n���T#¦v�� �rL˃�!�r���H �Ƣ}�����?o�!򄆺G�����X"L�H×獉|�!��O֝0veJ�9��ɲ���!�ĉ&AT�Q�Ve�ezRd�Q��!�U��V��&�
pW~�;��=	�!�d-�*Y��4X:\�c�l�U�!�dی~"E�&�&"��M�`!򤓓�<�,�Eĸ�gk��tg!�� ��P�jK%I��A�C(n�^i�!"Ozt�"l��:D��IVr�b��P"O�ig�I8Nά�òJ�#�*�y�"O|Ă".$��!�0�ؒ@r*�Ѵ"O�8b2&��`qaD��\��"O����{6�r+T�Hp"O@�hD �]�Pk���2C�h�2"Ot�0��K��Q�*`�iZ"O��D�Tq�tд)�+Y�r|:�"O��PL�B|���߃(��"O�}
e���~�B%k@�N\�Uѳ"O�C!7#�f��lC�+�t�	�"O��e��moP�"�.B�6�4"O.�qc�b���1�. |�8�"O�y���5����C )`@qA"O,�鵅��,�ź��&T�R�"O u"r蛲`q��bg��7����c"Oz�2��V��B��G�.z�"Ofeq4��Fε�eoY�#�j jc"Oz��&�$��3n��((8�`$"O�xf.
�!��Tb��
���J�"O�B� S�h9.Th�AD b�$P "O�Q��ᅿBWb�;��Y�5�"O��P�+�kИ��dB�'�� "O�!3�M�W��i�%䍵K���R"O���cG�"[��KS�{�ޱx�"O�	c�ʡ80y;��^�r�f���"O�����4+bu����{��)��"O �p�R�5�"q+Q�.�� Ҥ"O�8��n�5X]|�p�ʏ�&�ܑ3&"O��P����q<�k�o!p��;"O굑Έ1gj�3'��@��S"O��iq��e�8�d�ھ\��ٕ"O��iq.�5c�<a���X	�mx�"O�=�RH_�9!l�^AF��n���y�<=w��֦�a��L����y�E�&M^�c��(�K`-��y�ېA��i�o_#��@�����y�����r�
*�W!ґ�yR��_*aR��D=9�F՛�$Y��yB�8|�Iá!�?5q6eEoɻ�y���"!�X��IF@��`R.�y��	�@05҆GM�oV�+��ѷ�yBoȾ��<J��8>궥X��3�y�`��=A�o֐��9���y��e��H�FM
~����5����yB�ׅ?�`d��ܦ @��^��yć�x����-B7,�&���y�)C".��%)Rj� 䩉��y��P9��-���6m�a!�� �y�/D!�xR֏���vl,���;�'���"�3���
iUֵ9�'��9�Ē�}l���͟�P���!
�'���K��L����e�Gj(�	�'��P�Y_�Z���X83�^-��'�l0�C熑M��h3�	�':�~��'�Z�3+�e]� �dP�h��P
�'�t3�,��5{��AF�	�Uj�}���,�S�T+E�l_�Z$���U� "FJ!�yBBǱmMb���Ҹ=$ƇR��y�J\�+T������0�j���y2�S2p%����t)��AE	�+��$)�O��!= 5�U%k�G�P<��"O┰�FbC��X��~́�T"O� d��eǔl��e�C*K7 ��"O��2ÂU���3Ԩ��4���"O,p�ʁ_	z ��L-b,���"O�	��;�xh��EF�B� 	r"Obe�)� 4�ڥ27��R�v]�@"O
m�&dDoXƱ����x��%"O�ċ�e�,��$�Ta:X�a�2"O����@�M6�ٓ�o!Bδ�a"O���B:&�S�n=h9���"O�;7�	�2��2L��y�9i"Ot�RԣHIA���k� L����"O��`U�ӭ����Qi��:hr�pg�:�Ş��`���*A]��BAL�f�ȓGF����ϙbD�r��6)�
�&���ɭոqK���9�Ht;���[�B�	�V�H�d�lӥb%f���bK>D�|�
�:�q�aC�U>�9 �>D�D	�/K$bD��4R�Q:�yǩ=D��� �0ZڦJ1��'+@��d=��U��ħ9��@��/:�^���ǌ�IO�|�ȓ`(�0�1Ɏ�Z�.�#��Gp��ȓS�(��$< �|c�f�I7����N	�c#�#,z�Y� 3VH��%D�PqMCQ3��$ �:@��87��"GD�(�����	`���ȓk/^q %��*�J��?<����Xؠk".��v��
 OХ2��$�ȓs�݊�g'4�q"��#	
X���:�b�a7�\�",	k�
.�h=��ql�eQ7�ͤ�~���SG��х�}�f+��2�YI�Uu� ���	M�ɛ"l29` [�������ɺ��B�ə`�*2�4[:��˄#lB�I�p�R���aX6�2|�2�B�u�>B�	�#1��JUHM��
��ѣ�g�6&�DpD��I� �2'�5s�?D�t E"�6P/�AS�W����3D��yW�
/O,XQ#����A��&1D�X���
`bE3`��a
,�G�0D�؉!ȞN4�m�vl�K�+Ђ:D�(�CX+u�0��D�_߾M���6D���fh\$@�&ћ ��7ͨ�*�*D�x�W�Ֆ<��Sg��jAy�g&D���@��?]����D5PPK%
$D�p��UO���I�
;o4�RD�!D��B յVq�d���#@s ��+!D���FO��$��쓽o\���h9D��B�)�Tr�$!d��0��	�$!*D��Q�F�I7�<���C;((��3"�#D�dJ_&x�8��p�Dλ�PyRo�n0L�J�o�z�Rhd�Y�<�GS=P�Yz���[F���KV�<��,X'q|$��F�b���gm�<��
+I��e�R�Z�D�UHq�i�<٣k�:�j��r(�C��`�d����?ф@T�x��a�#��+D¬c���z�<Q孅+���S���$h��v�<���Ė��qP��A	~�,:��u�<��+^�`�2U�۹%��4��	�x�<ena8�3�1<��BKJ�<��� %6�)R"�_2G�4q�7�HE�<i	߳v>�B�d�x�����HJW�<��Y'��� �$r����
S�<i�͝�I�,�B搥"���7��K�<� v�
�ME8+*`�(ĉߕ(Ez�RT"Op0G`��#̀��F��k.�5C "Ovu��jL(/���j�F�Y�"O$�P���	���8�d�2ulE""O �P�n�?9�U���ܙ5�E�"O���e" k�,��P��7�X�A"O�)�&$�,`J�R�m�r�j"O�pPAH�n�����RhL@�"O��b���=id�#�e�:3��� "Oz`$)�&{QF��P�@���E"OJpka%ͳ%��y pÏ�h����T"O��X� ^�ìh�'c��<wL`��"Or���.�bS܋%�Q�S��4"OF�z�
T!A�LŲ���
E�B�Qc"O��FA}L�cԬp��H�P"O01�AaC6Y�Z�L�yn~��s"O̡��͟T)��	��*i��"O੊U���\	v���XO�!�"O���CXK	@Kօ�Z�Ђt"O�=p� )2�&t�k�*>,�"O�غ��&�N�J)�D$�)�v"O�Q�$��(���tG?v8���"OtL��F\�F���g5躑"O��Cc�+_ 4	� G�M&F��W]������g�.���ܭ�������2<�C�Ik�T=��+�K�ic`��L�C䉘XV.P҂Jˢs�ڄ�W�B?4nC�S�9�iدJi�HyP�B6{o�B�ɚR�$-لhW8s�J���d۵��B�ɶtR����Щ�&�r��ّ.D�B�I�]��JO�>�xQ&8e�B�� ׂ��'�W8��8��L�B�	IT<�C��#�V��EG-MhB�ɯo��8�l&�F��kE(~ C�ɗ:�%nԒc�~���hőZ�B�I�{�\�@6�T4bR&`����B䉈B�ز����@x��ݬ8��B�	�*���S���^�^L��m~B�ɨ<贅3�eāe��8�L1�:B�I*S�Mj���Y��\�5/�2$B��7>����LCZ����h�xB�	��P���Bv���!9��C�	�/��%��gJ�*��H���hP�C䉍$X��! %������U�tGDC�I�!`����"����O�CvdB�I;;�(D(d�ȎAz�;slA�{T�B�Ir\<K�$1M1p��VA�!$C�B�Ƀ�T���D;X���[1(��q�C�	�;T�!C�Q��Ƀ�LD�
�fC�I�1�Dxx�G48i�����o�C�ɹD��ؠ�>uD)���]�XC䉚`x��$��?NY$�z�
, ��B�I�V�[��0 ���� �TB�%&`����L�� YR,QU��C�I�l��k�/W)o`ʌ9�+ҭJ�B剠Nl�L:�hݼ7��I1���.!�$�&($2LA)ݤ+������ֲ+!�d1�j�����k.��T��"�!��Mr���BꀇHZH3�kߝ%�!����.r`���pT� �A�)Y!��Z�ok.�Gm_�A7X��M��$ !��>k��A�o�^m���@!!�d;"<5СƊ$�Bk�� �!���|�ɓd��1�l���D8vC!�� ��(E��DjL�{��fJ�b"O����%J�|:�	��0>*�!W"ON`�*�)@w���mQ����ѡ"O���g<$�~Mx��[';�|��"O(���(��6�MH1�S�E�	RP"O&m��
	]��# V�쬘`�"O@g�3��0�EU7x��!s�"OD�a��_:����E�M(3�4��G"O�`���ŶUPpD��  .{����"O�R�I �X�h!�>/[X�ʱ"O���ŋ�e��<��GB�����V"OD�
�J�/#.e[RfӘ)� �r"O\Y�@�;OP�kÅ�LаD��"O�ʴ�]�I��a��.#E�Dt"Of����7B2,�.	�A�Y�"O��;�م@z���
�r�B1d"Ou��i��ްAW��7v`XX�"OѱTD_	-U0�Y.ƕ,ֆ��d"O�e�����h]c���D��ݚ!"O��w�#.j�	sQ.]��P��'H
��������VD�WJ ���'�|�pf�v|ⱋv�ދJ�!�'׮�c$�h@�Õ�Ğ5�=p�'�<��S'�6mN��J����-�V�1�'�����k����S�nD.d1�'����c�#1V��(G>���"O��A��Ɔ2���q�	w٢9�"O�Y�� ��6�N܈uL\�q�R9��"Op���+��\��t���Yr�j�zR"Oj���-.m�F���7�� �"O����^�SA�t���\�.�X�"Opj��G�N*���@��P#"O4���cH1,e�yh�HF'%q6"ONq�WG�� �4��%g^!1O�=!�"O^�zW�!�ʠQ3�[�;���X�"O�l�� ��G!�K�۞y����u"O�����
O��ce+Q:�6Y��"O���0�݀1FR5RA�m� �f"O�M���W�ygv��I�,�"O�Y9��T`�9������e:�"O,�@P�A�Y�a�2�6"O�=�$�Q>a��M
��F7�4�v"O�2aP0%L\�a�Q'q���"OX�I��֜À�(e��2$e���"O~A#7'R�U�Y�pIKÈݴ�yBDȗ��Jǯ�79�ӏ�	�y"��_R���T��>2����i��yfP�BL�2C�S��})�fɟ�y-߂�b����"L{ĝ�r���y���&p����j	vT��uG�=�yb%[�|w�fME3rdXx��b���y�l��Z� ��h܏dizQ 境�y"��2Z�.A���`�=�a��>�y�C�-C+�̛GA&dlQAH��y"��+$�
l� z��OS%e8ЅȓK2f����R� �p1��p\p���;�bW� �w눉�"l((�2���bYs�돮~R��Ёju�LE��@|�݈�%?9 Z���nY0"�B��ȓ':b�����E�4#ڳ9��D��`|B�aa!���;�뇯8`h��ȓ��lY��*�d;�H��tWnl��d���Λ!n�R��͇W�d��A�8� Y g�{�o�� H݄�S�? ���hʌ7�JD;�3	�����"O���q��x�q╊�Ltx���"OnH��(ҔuU�	S����iqFA"O��:�/�A�t���H�`�T�"OT��a�+v܊ {�Eן(���A�"O~����@�IP2�c�i�:1�`�C�"O���$
�-%(U���!d`u��"OB̚�B2I2����'�
A2��"O�mѤ��|��ǠK�P�0y{T"OdAB5-����:2`̵T�&u�0"O�cC_6��,��mcH�7�yB.�&!)���ġ4p�4�Ҥ����y�  �{���K�U�i|�1��X%�y�bŊ�H����-�I�2���y�Ú�km��J� �UO�h���T/�yb��?(|b<6G	#O� ���k��y�퀉l���� C�Z_D�z��ْ�y��H~t(m��*�#H����3�V1�y��ޡq�)� ��</�h�jY��y"
�?m6\��w��&`���B+��yRQ2)�䔁gЦ�@Q���-�y�Ϝ7AB�i��e
�@�*Y:�yҊQ4/�<�"����-ۀCŔ�yB��b񲖪�3}5� i��y��|�����w�Q�H��y�@\<C�0�`�K�n�f�!c޷�yB��#a��R��2���;����yR�T�~��dЦ-�r�H�@��yBΗ�MO �Ȇ���1�~�������ybX!&����3��9�v}��!O0�y�KB�9�����?ʨ-c O��y��ٌ
4a:'㜣Iif��f �y��J2E�������*J^���H�!�y�-WFҠ���ϊ$8H�TKL��y�ɞ�xݑ!���M88��a���y�K%xn&�Q�.˛������y�b�#k��9��כ�褚�JQ�y�[m3�����@uA�ǹ�y���Xvع�Uj8�^y�W��&�y��Ǉ!�D �	E�3F���R��y�J�6?
ڐ���)�"���!�1�y�oV�
MX���#�H�F֦�y� ��K�qg��� �b� 3
é�y2�C�B��p*Գmr��!�X��y��jX:�q��-5B�����X�y�bàm�J���$#h40�J���yrR�7�z������,.CEHߩ�y�-�=��b�C�A��&��y�gR�Y�aFG	�b����\��y¯��$��ŉ�8<,P��Ƃ�y�o%��F�</���(g��1�yb�ȶ ��A��ޑz&8lk�G�y��+Ir����7vj��#B�yr	�0Wr�<���(o>������y¨S%K�$�;U���	��U��y�&֙w�z��C.�E��JO��y¥��v�����HEt �D���yb��L8p�I�ރ	i| :�Q5�y2�W�0R��qĀ�Q�BSMC��y�@&Z!r-�h�4�xՑ3���ybMX�Kz�8R�/F�;�rI��	;�yB@�)&�2����,k�+t���y�
��U������*���3�3�y�I� e������;0��I�����y
� 
�Ɂ�Í^�P�K�o�<%L2��"O���b��N{@�����F� ��"O��1���7?z00��|~�-*�"OD���ϗ:4��D�R�g�8�S"O�t��\2 ������eg�Q"�"O��Ǌ�+��=�����%bP���"O(�`wQ=���!��0�8��1"Op�!�č}�dH#�k��n�����"O;��/H}�ǯ�L�J�Ie"OR���)��-�M�<�P���"O�X���5�F��*��Y^�Z�"OJE��Ο�|��Mb��ʍpV��"O�a�ė+b�s�%�8���c"OH,�K�8�@�DS1Fz��A"O
m#F���PH��AJüu�
`��"O�@�l� �ؼ'	�Q�h!�v"O�� � ͝;�L	IF	��8;���u"O�1q���U�6��w\�/�<�"O��Xv��3w
TS0�Ŗ 6L��"On��%��=�FȨ#bQ����Yp"Oڈ �G�K�fu�ԂN�i�ƑP�"Ol����Z�q/xա��8�����"O�X�m�%���&*�ʌy�"O:p{5![*�:�B�\*_70h��"Oƅ;C�� ׈M����f*v��D"O��K�@'8Z5Ò�ӑ��l��"O:�s���9�zt��j��"Op k�%N!{�)pe�� ~���5"O��������~@z�	��r¡ "O&;��ӘR�������zDXh�"O����X,�Y"e�P�=*���"O2�A5L��fi8���.r�N�b�"O�lI#�%(ߦ��%�T����"On�`��ظ&�:x#`FV�)���G"O�] Ud� j|"M8Ee���"O���Re
.��C�%�l葈�"Or�%I a���G �E�U"O����E ^5SCFt]���3"Of��0,,c�x��
r.�a��"Or�0v�J�ظ��X����W"OIk҅�.gv�8%��p?��;`"OZ�C�	�&wY|Q9��#/4��)%"OJ�����. ���CJ�~#^|@�"Ot J�C	�h�숫P�^�%& `hT"Oz����b���H�S�	X��r"O���r�j�q�j�<#`�A6"Oܝ�Agɂ#?Z�S���ab�"O���Ņ�a���� �'mmD �"O��+�-��E����3 ��@fr��"OJl����2��\	��ѝ(��4*%"O�H��%�~pȓ���h j6"O*�*��0�Vв�+��v�𬹲"Ov��Ǩļ��Bshӊa��D�"O^�3ca�y�¹j�&ה{�䩰�"O"i�\*֠B�@��%�:q!��A��y�,�9��#��\$��1��f��y�,��<�~E�3#���~H ����y��ڹE�1j����~Y�5�B+��?��0eL�Dئ��dX��ͪkj�� ���x� Z�/8���G_�xJ�(�E�C��y��=C��ѣ�j�F���ħ��y���9I�2]�t�[�DG��C#D��y�)��Ҷeב
�( ��"�yr��=|�pFK��n!p)�a"#�y
� ���V:b���k%����	F�'��ߖ5�ȣ�k�Y��Pg��'WoBO���1
70~V�W`�)ՌV�<	���L�BgϼS��@��P�<���+\�RQ��Cޮ+����c^b�<9� Χt��pqua��C��(���_�<�6� /"����lI�$l�ȓ�p�<16E��(����:r�bl��n��p��]aVѸ��3���[!揲q�T`�IW<iu�)tV�yPK�7���b�Zb�<��m������El�R3%k�Ƙf�<12Ɨ�?r���a�L��1�G�m�<�Co��'��q7-��Q�`陷�k�<�1�]�昨��˂W�
(�㡃O�<�0��:� ��5�MRƬ�9p�G�<Q�!�i�<�8r��pH����@�y�<�f�_C�M��I��4l��y4)�J�<��A�)��]��ۄ���!�m�O�<)�$@�Y���Q$�m��0s�E�<a�o�'�")��Qj�}�@�l�<���i�쭹�j�0�B���f�<1e-ޞ	NH��� r\f����^�<���V<��d�i�p)�5� b�<���<A�f�q��-v("#��x�<�%�P�촠�V�Tvz�A�%}�<1�g�%D���RE�&�})��r�<IƖ� ������Y��\�Hr�<�d,�
8�$B�1@N��R��D�<с͑[q�e:�lL�7�ҥ!��BC�<	��!!ݸi8�n�JG<�I@�{�<�G�I�xH��ɅS�DP!b�b�<Q�U�N02i��I�?�tQ��D\��z���O�t�!ޡ��M����?,�Y�
�'&��Y�� n��ئK�#)ӤŃ
�'b�eA�IS0X����%`� V�L�	�'$��cK�6�� ���\��D[	�'����'��.W�L1P	���D��'Yf(��֢E~bg��(�0�
�'&z<�ĞEJ���.��ey
�'R"E&���M!��S�&fF��	�'X� g��|��p��ETS��X	�'��#�aM����B��v���'HZ�rW��2�����ޘzt��'>�8��mP���m��������'_,a��OT���th��)̶}S�'�2P����G�l�l*������0�~Y�-�WÖ�|{�acg��6� T�ȓH{���d���TȰq�֌v4t��IN��@q��22����_D9���ȓ7�d%��3	��q@�čI��܄�8��䢥�q���k�ʁ7�<0�ȓ��N�f�xk�e�?m)�h�ȓ��1qB��
'����My���E{r�O��h�ҤשH0�!y�d��	�'��iȵMx*�sW���pPֽ"	�'Bf���(�,2�2ұ�B�a$"��'�N�# C٣b�Y�nG�Z�ڈ��'@�!�c9|M
 cї)?HX3�'
 ��B�Ғ0������P�U1"�X
��O>�!hEê�c����@*"��i>�#��Z�u�ba�%�;��$O9D�dp��^�}��ݒ�U���pk�j"D��{R"�>*���A���iæ?D�x��	}p&8�?�~U��;D�� ���&?:֩��#C�p�b"O	��K̔��Y2(Qo58�"O(eR�Ȅ|d�a�^:������T�O�V�s`��x����"̠1���Hw"O����+�1{4��N�;I�ִb!"O�ř�9xː��a��	��Ih�"O"����*H�!J�O°{�8 "O\���̨:�F-�!��Wݘ�Q�"O��1q�ˁQQ~}�珖�Y����"Or%�j�=T�����Lʷy�(����A>Ap�mFg��	���U�u��)D��2g�"^~hPԁ�*M�jE��f-D���+�Sg�E��c�(}0���.D��֩��p&��ӄB�#$
����-D��z��Ь1�Y��F�c��D�4*O"M�t��DX,�y'͕"�=0��'�1O�� ���[�jM�����)�d�IS>�Xp-٩�N��B@ЋjR���B.D��aSe�U6 x ��?�4��!.D�X(5JLG��Y8&��q�^R��,D���� :x�y���ڗ4�"�+D��ᶪ߀K�N�GO��<�:"d(D�C��ˢJhj�y��Ct�� +D���PA�
e���1q�h��	$()ړ�0|����FQ両�2
�r!��N�<񄥛#��Ԡ��+G����P�]t�<!��m�&����ɨ �h�*t�<���N*]X��k���!dNQ0��s�<���"Z@�A-�(L ��PhWl�<)g��2G����ל@���Qu'�h�<�iI=Ɋ�ځo�2m_DmiRa_a�'�a�$���g��wbt�b�K_�b	.8�ȓ�� ��-�3Dl����	B|�p��C��H��-B)����!�<�J��� �d���1��G�D�.�"݅�)�H냪E�x��[���8<����ȓp��iI�n�/��ys��FbpA�ȓK�j�c&L�
B�����¬arn�D{��'�?٫%%֙��$���E�S�:}q��'D�X�oі\�
�D�6� �C'D� *�i�<}��m6EN`k����O$D�`��ő�t�E�Ŋ c���!0D��b��`��ʵmC�"��<��M��y2O�����+G+'��5����y��G"B>�أ�Z� �p��š���hON�b��ʿq��8`N>�^ �4Cן�y"��;��M��,�0�|������ya��X��oU&o.1R�G��yF��PeS��W�~di���&�y�C�*�I�q�HC��
VHZ�yҧ��4����H?��e|��S��%𧂅77�`"MD2k�f0D{�OѤɲe��k� ��	4��'1R`�� �4#�TS$c�!�z�<�Ď�z�C Gc�x��6͟r�<!3T]�Tz�ZKK�a�r$�H�<��9kTU;�(9ڊ`&��H�<qU��;;�`�"�Dr_����m�<�W)H�;��:�Xx�Shl�<9�O �SMj�����Na��]�<�f"W 
�*<Ȳ�ԗR+�k���X�<��jR�"#�|��/A-2�T%�C��<Ѧ!N%M\�z�Щ �t@0R�M�<t%ܴ
s�mj`a�9�IA���w�<� Z� ��B�H�тټ`�8 R�"O���Q�K�7n��@'o���P"O��(��B�c��6�ߪ!�(��&"OP�h���T�(۴�ΐ1Fd5��"O����ѫ(8$��d���6d�F"O��3v�^��]bg���E�3"O�dB�@�
�
�	QY��@�2"O",�V� !@|�2���^�&��"O����/.%��&�ʢ`p�i�"O��h6B �t`bux�-��W����d"Oz9)T�� ��0�d͉!��C�"Oܬ��Or�ꜣ�΂<f��m�"Oz�s��?�1��N�;E4�Aw"O|l�D%C���U��$�"�7"O
l9��J�ETxX"��~v��w"OA�耥e�]@�
�/��\�E"O8q�`	��l�GGʡ?�0 ��"O���]�
�*�Ɂ�J�򤜋"OB�*�$�Q�X�
3�0e�P���"O��#���d���w"�%ݾp�"Odق,�u��1��
Y4Z�q�"Or`�T��@|Ơ('/G#�q��"O��+Q��~M�uA��	��"OR�F*A�dר@�$S'x��)�"O"�;�O�&9@0��lTc��D�"O�ŹaeT�D���ŉ�Y�NP+�"O�h�5��rk�NU�McC"O���cG��	y��0��M+HU�U2�"O��RlF�\>�m͎*OD�9�"OP=a&%J-.��`��^�GARl"u"O؜"�LE�e��p��)ސn%r�E"O�%�dRpb��
�C,���"OJ	[p��k?,��R�J��Q��"O�q��Ӫ"�|�gF�	f���T"OZs��.&�zx�Ŏ����I�"O�	�M��(�y�B!t�H�G"Od}�1JB�H.q�ƥ�>a|h�"O�\sĞ�j��r�"P��Sr"Oa���T������?]�����9D��;���(h��9��+s�jA@-D�l%��hk�*��G'N�v#',D��SU⅊!�p����9U�4m��a(D��IU�F�A'��[V���=2"}��K'D���fBԘ[��Ś��K$��A
'D��  % �ng������5��qJ6�%D���d� �
���Cj$�1��&%D�`�!�(~L���fBƽ������"D�d��(�׈Y�6��4'�ri"�*3D����aA
z8.�xq��e�Z(� 2D�lbC�:N���qW�+U����p�+D���q,>t\&Y��$M��ɷ�%D�@����Oy�쀕��g��ڗ�$D��D�S�L� h{q�̓�hmi�d"D����w�a�O�;`�)���2D�`�E�h"�$Y6�3 "���=D��!���nˌ0� C	hTmZtf�<���?�M>����|�zt+�L�_�0 �a�=7��C�ə!��,�4��,_|��` �ϸMTC�	�Z �7ċ2,��y[��EeDC�I�="p ��ędV�QҗKΦ^�C�	�-zpچ`6$��0�˕j�C䉨V���ȷ��|�Z1;��L4u�FC�ɷ.����F��p�i�O�(P%Rʓ�?َ��)A�V��	B�J�:jP�csH"u!�� �p�g&J=D�� ��<[ܔ�A"Ol ��,K�y����g%ЍD�L�p "O�� E�Wb�е�ʰH�<Ÿ�"O���T2��c��8��+B"O�3FCo�,��%�����"O-�¯��gg�쁦"L�;����'�1ODjq�'��>]+���1�L�S噫?"N���i�<1cY�(�lI[V�(x������I^�<	�)��b��I���\P"$j�	U�<i6���V��Ӧ-����NN�<ل�Q
?��Ƈ�%~�U)�)�n�<�p��8�q�DӖT��O�l�<�$�>e��S�K�V�P%i��Jk�'�?�³,,P5�t@Q���twr�B4D�l��'P50,��st��:Y.q��=D��p�`D�B}$(3a͝lO��"(9D���Ņ�rB�y�� �0@t�,J$o8D���M��&`�)�����z��1D�l�U��7��H�ge����2D�|�t��5(ʪ��2HK�wex|��-5D���GJW�Z?��K�,3����1D���E�T�V���j[��$4D�l9A+@;��ҮZ�l
�\Zd=D��;Q(G:|(*�#Pʗ$m�<Z$-;D��:���4`�h\�#Gի K�2�.D���*ݜrID����ѩ� H:�+1ړ��<�Hu��C�|�MC�[�J`�w5D�P�6m ^��"n�,;$T���?D��Y�#г��@ţM��@PU�>D�Ⱥ���!ܦ���nħ�r��r�=D��ѥh���xXFnA�-f��u	<D��i��3j� e�GC ��0!�;D��p�J
o�����\��:�%�O����u�6�qNF��<�k19B䉰F�&����Y����P�A:V7�C䉺t���`�ʚ���A
��˓�0?��J^'< x�(@�2�Ak�<��,�*/��Da��26�B��e�<��eT���ٺL��h������~�<��!R�qS�e�sn��XD��Q�G�}y�)�''�4P���0�6`
�J �Ba�����#bɟ/eĨp���%ĺX�ȓ
�TaũsIVQ`��ة~.��ȓz >����of�}�#�_Ά��ȓ?��A�K	�L#QzA*�[j`��#��U��kN�a�z����w�R��ȓ7����Q���V�I�B�9�|��	@̓��
�\�p<�1࣊�0D����tށj��1]��#�Z�=��Ņ�W�Z(�E!����Ǆ�L`ԇ�,�=�C��	L�`T�W68���~r��� $?��T&��<��Ȅ�.��)I�&=\��(fjD�=�TQ��B~�y�PE��!���6�Ȗ'�'����y>=�͉s�萐#�R�zIQ��3��p����B����}���E"n�"\BP�&D��
E	�-��H�!A�6B��Z�m#D�����1�j<jE(L2ie�&D����AZ�4G�\8:�H�6�$D�䫲GUrA���p"�<HҰHHA�'D��a�b̽s5:`�V��b,r�ɑ�#|OP��!�ٮ!ܕa��B#�4e�|�Q�E{�O/�����}�Ja��f�~HX)��'	���pLJ�稜ʧc�4,FP���� �yC���"nF� �W:>�(1��"O�t��ڍAV]Ac�8%���	u"Ophȃ ř?@T��5 �h�c�"O���ԯS {PƜ���.���&�'��<i��N���Gnو	�va��<A�r�S�(%�;�B�	E	B��a(�iDXC�� ]��8��
�P"�pV��'�BC�	�~,�eȥ`Q�b����M� C�	N��p��b��Z� ˴��e��B�	�C>4��; �P=(s�	b�B�I+2�R�0���!�Fe�#Ǽ%����d7?�&Ć&,�aӠ!�Gc�!Xf��R�'a��힄I�*d���X7 fL0*(�y��ŷ/Yb���G���hOP��	��s*V,�f�4�ȌQ�(�t!���#:T��
��7��B��I�!��G4[_$���	��y��	���>LP!��1ؼ,!%�M��FT[��]`ў�'���|�eC*6���j��H#?e԰` I�U�<@)R�J���@K�Yv�Q�<Q�)Ln�]��c�]�`�6�MJ�<	HH?i�1��Z�=`�1��H@�<�&�'�͘��1>�I��!T���F�<N����`Cl��貑�7D����6���Q2d�8eX�$�� :���3��h��Vm6.2�|�R��)t�ڒO����K6Q��x� ��[��ڀ�(r!���2
��)H�R2�p7�{����H��6	q �I�`b�0{!�$�J��g9x���
�=O]!�DN��e�"�K�B�¡@�n�!��%��� Q.�o�F���@�S�!򤆿[�E�Ū���ʹs
j�!���i�tЛ�g۪?��l9�I?�!���w��'s��U@t(��^�џD��۟ �|2ECE����@6� �y��Q4oCc�<�v�9t�U��(���y�$�_�<�Vo��uZU3"��f����t��[�<��$�*,�ţ�G·y��i.�m��X�<�B�%Qч�/�ֱ�@��ry�)ʧ=9����\�J�D'
WƎ��b������3�n�@�������m�E��x`�i�I�����U�vC�Ɇ���%A�D��&"���FnJ�����ȓv��0�V�%!���F�Č'��]��u��sr�B?Jހ�S�֢Dq���I����<!�M$��1�Ĥv���,�Y�<�������'R�Rt�xw�	X�<1�G��U��M%�p�#wFR�'���'�1�F��gJ���)ꠌυZr6ySq"O�-�A�E�4�l !���eZ�][@"O%ZVB��4|���KJ7p�<��"OИcT��o�
�&�Īq/�ᨒ�'#�I�.��tYס���܍�0d�pm~��hO1�:�	9R�Re	ƀ�r9���`/��l�$�)�����ջR���h�ԥ"#��$(!򄒲
k��;��N�6��!�uM��[!�ο�J�k��S`�;�N�,]�!�dɛ�^ ��.�.O���V���!��Tw4��c؛u,2| ��P�!�d
�&�I��b��P�x�!�D.*p	�P�A
Aᲈ`�BT%8.:Y�Z����I�R[ę9� �4b��Yb2��z�B��3#��2��G�0���"˟�G$C�)� j���� 0<v�ӉR�aƞ���"O��q�aƭ|���0�D�~�d�Rq"O����U�/Q"��E�\�l���|�P��%�8�<� ̔n\bL�1ő�D��u�������&��L�&48Bm衤Z,$N<��ȓ}Ҍ p󥜐gt^���-�*A<���o��=�N�70ڀa$�E)HΊ@�ȓNz��z�݅~bB���̌�v΀$��)��T��8:���:��h�zx��.{�XQB)n8�Ш�dA	z��X̓)�8��]'3W���(ΦJ8L�ȓqʴ)���-��e;��A#=R���Iv $"��	�}S`��G��\�'_a~�F�' �ē���d��$�W���yr@�&	��<	��:�p�iW���y�LB�Jn\;wǭ��8��9�y�ş<|��P���˳m��]!r���yr.��2�墒LJ<i`(�ٔ�-�y�>e�Ŋ�]�ٰ����U��y��Ի)�}�B��(	���SU�:�yb+�?�I�R���,��}���P��yRd	׀��v��-�E
c���y�j�6]�� ���B<W�}�sՑ�y�@�|��8�":���)���y�;��H�%T+Gn��խܪ�y����� �$��bk���g�G��yb�P�%�,�	��<p"�U�&�yEݻPb��#�K�[K�Y�UM��y���zQ&pKJZ M���� ���yr����쐊1v�u���C�d��'H<	�*�.\��p�t�Q�m����'��*���"o�L�	�X�=�����'�p��(I��}Zү�h���s�'}ԩ[GcU0U�v0��ē�sYZ��ϓ�O�Iv�(�^��j�%u2 Q"OvhH��]�kYJ��uK��1�N���"OJ���$��`c�9�&,����`�q"O~D��F�j��\�v+]�"b 8k�"O�\��ɟ��ԑ ck��)��"OHBw�ěQ.dpC�J&N���[�"O���@C��Z���(�1��'�b�'���똼�5�>�@��S��Rm!�D�!�(53`���K|��rJ��[[!�d�R@��9SeS�&4���E�J�bQ!��245�Q��n�	,x�L�ŋ>:A�O���D�a���œ�9�NIs�ي�yo�kpd���KG6|�Я�f�6�$�<I5�����f���HV��J�l�Feɽ��m�ȓ���(��)G�5��iV J��ȓ,:��cM�BaC�ԇHe4}��H�&��e��[�U�$���|c���#�^8��
�h���M�� d�?���?����ƣ~�4���4:9n�2�\�4k!���,Unu��K(8|3��S�}Z�2Oެ@s�|���M�Ҏ��pFƍWhAcB�l�\C�	�kD����E�U��Se뇑g�:C�I$9�����@�Y���
2�h{fC�I+*S����*ip�Ѡ���FH4C�I�+c�q1���6�l-��웣L�,�4�'E?	9���/�X|(�ԲXkji{�(<D������!z@b�N��t���;D�� BLI�S���R�a�th�gA:��/�S�'R�(<`0��v)�U��ՆgB�T��M��aK�S/i�P)vd� ��D��S�? r`�MJ?06
H��!׃v�>��"Or�;7 �L�� �-�´�r���O���2�'m��q�]������/ήP;�4��L!J�А��E=8�"�' �TȄ�W�jܲ&�ærV�l
gHnA�Є�m̓U�v����gdP�! �L	Zn̰��
x&`"&��y|h���O�kM|��*�ఁ�NF!f�ʵ��f����q!q���2_L���JT�X���ȓ�<���N�+�6衑L%G
���?)���0<�s,�5+�$��ϙ��
��ě{�<���U1#�Nc%瞝�Up'/�R��`��N~BoL�:����H�;n�<j �];�yB��A� �s�5��t�B3�y�/K�zI>��F�.:Y�M���؀�y"�NSX(����pH�B ǚ�y2��&�U���q�E�e��?���p���ѕO��m�å�5�f��3B+��0|jri�V�h���G�jA�T�<�@�G<	K�s��u$ޜ�6��L�<y��_�C���"JԼv^N��c�O�<��a�O54Ѣ�a5�p|��)Nr�<�ƃO�Qa1G�+�H8���H�<1 G
	��q�*
0k� ��#N̟�E{��)J�j���"ڥ`D2����M��C䉚*�� �	������B�I.1�Yr�L�B�
���@�<�B� W��qQȴP�� Xe�ހA��B�	�%[�RRGK71������^/ ��B�ɗ!J��Qd\�M���J��dwJC䉃08D͋��Z"zAta���>8�vC����U1)J�Fo����L p
bC䉕B_���B��șp��X�kNC䉴Yn�e[lt����a��5vB�	8��#҇�� ��l:�,E<B�	���ibMG�SܮLx#�ڷ
�C�I�H~ɇM�\�)���)�NB�=\�����Y\R�����C�B�� (9ణ�*��8|&@ەg�
8�B�	,Oh���JV�*�<�r�ܡ~��C�	�)(u��gSB BD��%��C�	Z�6�;`-�5	�0��]���C�ɀ����ؽW~�P��L��7��C�	/��&n�"�X�K�g8��B�	01O�fVx`�y�7ĳ�B�I5Y�ȣ&	�C0��cO�-tb�?�����Q��J%!p,l��E��'x���"OA �Z�a�����DjD�w"O�ȡ�C�*��E��$�%Nɦ`$"O"��w�*kna��b��&�l��7"OB� v�]�9���a�|��8*r"O�a�$P�s칻��3�8}�"O������C�&s����M������a�OP��Z/��%��2seK�v��E �'l(�y6��ir���B�5\y�4x�'%���h�#PĖ���K�>*j c�'��X���@;P�3I�%��9�'� � ��çQ$���B��5[Hhb�'1:u(&�S�b��%S�e�%�\���'�z$K���q-Dy"t��$l�Y�'����(l ��P�_�B���'�N�$n' �&8m`�p�'q�mb�P%<e:����&g#\�'��t�����R� �3�eƩ/�.�p��� ��6��]� {5)N	 �.�G"O>��D�NlS��v�6I�r�Ұ"O��g��0G��0�O
�܍"Ox�t���� ZSk��
��"O��Bu�B6dց
Dd�1��d�t�<���H3:-La�)�T���%Ft�<9Ǩ5jC� c��j�.��Tk�<чc]�[؜2�,�7[Lx(�(�R�<���B�~ٚ���<��Q�M�<��E+F��  �ؐ-g�D�$�D�<���x@Sb��{��ԂtBID�<�#L��t���1gѓ::-C!}�<��Ak"y�D%Qr���{�<��0κLp���rrbq�1́y�<QF�żBV���!�>Jl�gd�\�<٤�GB@#�C�P 4#T�U�<Ie�1$����qdN�.���ҁT�<Y�H^i���^�z��UR�O�<)��}��ȧ���,�8i�N�<��E
kn)	$�܇`�0�Y7L�J�<-�i�H@��#��5�ʡ�
D�<	sJ36$	��I�j�A�<��'֐���#�o�B^�b,�g�<�sg�8OE�)֏^�L$*%�C�o�<	�A9#kj8��!aY��c�o�g�<�BMP�b��*pf�!>".d���M�<��(��U�Y�3����3��D�<Y�"P7����qdJ?��HR��i�<��(O�y�3M��q�W�K�<y��F�ɒ�/�tI@���BI�<��`�n�bK�D��!�p:`�]C�<��GI�j�挀�J
�.��42`�{�<���5�^E�"\�V���i�ɃN�<)��6O�}�VH�;4)�$I1)�a�<�-�kj����ӎ�HJs�<��DLF1�.Éh~̻!�Mp�<�g+G�Q��4:R,�]}Z<�lVh�<��BA�)�TQ�MQ����#ro�z�<A�E��T)�-"��T<1�.�r�<�&E3Md�5y����^lD�(�l�r�<�f��_�,K�AF�:X��G�l�<9f��4zM3S�׼E��% ̓b�<��Ù;��2�o߂LyT����v�<)6"K�-��r �<e��IpC"�u�<��
m�p�H�gR��!�}�<�᭞�`�p4)��_#C�E�0�v�<�C�M!C�L:�ˀ����H�r�<Y�������e@�J��扂i�<�t�AG�%�	Ҷ'��وV)�a�<��ܛ_)��pddE�e@l��&�I�<��Z��f�����+	��H��M[�<Q1W�o���
� �����W�<i��B6OM������w�Yyt�R�<1��S�L	��� ܮ)��H�GK�L�<����,6�q�`N,R�9���I�<� �	v�����ۤv���'�I�<�P�ם:���%��ecT89R�B�<iE)�  Мeʄ��$mBF*@{�<��F��" �����Vd2#��O�<!@�G����'�[�ԭ�|,!�D%j�H��D�x���؃��:n{!��C�DDx��0'��� 傱I�Dw!�$M�)�6�҃m�-@����G���g�!�D%=��% Y�r�dRw"�`�!�� ��p-=`�j����P1y��@$"O&�{!cȯ_t���e)6��h�W"O2�	C�	 ��=��S�\��	�R"O���r/��Da������wמp�"O�pJ���Z�H��Ҁ ��8�"O�A�g��eI�I�BW9e� �0"Oh:�A�)y"���dAC%QE2���"O���`MI~��Bc�/4A�RG"ON`Y��޼7ʄ�S0K/+�9�"OFmc�K�R?��V�\8.6���"O�y��L=�����̮<3�Q9�"O ����V�$66 �r�F���"Ol�(ƀ�N!T�z���;T���"Oذ!�
^5Td�*$.��%[�"O2ԫ�*ʐ"	�% g�9+iJ1��"OЍ���8-MH�4�ˤ`�B�"O�ˁ'�,�`�K5^(�0"O� 2�D[�/��p�6-,N��I�"OJ<zpF��̴B`Jʔo7�rp"O�M����-F|Ha�Gꝩc}m��"OlP
���67pL��c[��Uz�"O�8j�LA�6,�Y�r��?�R�i�"O�+��]-"���I@$ɢP�@�B�"O��ۻ&��`���;h����w"O�1�'�z����|`){�"Oz�{1���x*��W�wQ��Q"O��ʤ
�*O���(!���3$�5�"OV�b%�L� �r
W�w$��"OP�����3ҼQ ��)j$����"O����̰58E��.]�)r"O�+�m��,���Hc�Թ  �R"O	M��pٶ��G'�k\�@�w"O�8�(N�h�,8c%DG���"O�`# ?:#t};A�I3*��iT"O0�8�#L)L��AXA�>_0!z�"O$�Y5�ߘO�������u<�XA"O�2 
��Cj�D�4��1w��"O�|��o�C+���q�ܒ�B��"O8e��!��8��`�?N�l�C�"Oΰ�0��j�N�{��6:���"O���C��|�L�)�H�<&�C3"Ozu���S	5��S'� %*�"OM��ƛ�tE�  �Ɩq�<�c"O2�(� H�`�ޜ�ec �P�9j "O4cv�\�<�t��B��!��e�"O�@�1�%��A�5"S37R09R�"O����*E<��XHt��92��� "O��k��Ν7�eГ��(`�Lg"O4H�ec�,'�F�U��'mZT�e"O\	���}=�8��H�z�P��"O"$��Ȕ�t���S��, Ү�s�"O
��G��A fy��X�5�,(PD"Of�0W.ա�(�Hѐ;�� P"Ob��"��@�f��&��@�:��"O.���bHs��o
�l���"O��I ;;����=Z␛�"O\�P���j�"$0d,�i�M(�"O��!a�rV���Q"xi��"O�yrA�ǚ��� �	ܝif��Q"Oi���*.j�Xڧjי_(��ɡ"O@���<&x���f^?N h="O ��u@1���2� �qlx5��"O(��/Px5f�P�akP�|
�"O��9����[ԪPAQ�}�B���"O� �<��c�$Ȉ���W5<��]�"OzC��h�@� ��Z�3w���7"O�t�dJ�K�`�0�[!=[����"O�kc	O�NKZ-�fM�~DrEw"O�)Q,I	>�
u9��B�a�<{B"O�m�+:fڮL
�ӸfԂ��"O$�;���"�j�c�0���T"O:=q��֣Kc����I��§"O�phh�R�8�7a=[�HQ��"O�Ё�
E�D�r�O@<�A�#"O�I13JӼ��]�W�.���c"OT!�*9Ұ��"�.] C6"O��C�O��\�x-� aL�+Z�a�"O��)R��S���c��
MH=`D"O@i:@) Q�m�D@ZL��qA"O
8)�#D�|�Dl3���5oaz�"Ov�ɀ`�Bd!��.OiV���"Ot���˂Ja��Ο:QT�:�"O~��sa����sM��8T��"O�$j5�A
Ǝ\�1掵�P��2"O(� 3��!	����#�_/PWhd�"Ot�@�n�X����W=|FZE@�"O�������q��^.�AK�"Oa� �' К���.F���q"O:	�$E��|������HT*��"O|�i ��]^��j�^����V"O�H���^{�n�2ՠ�'�b|�"Ohz��5�*�R3O���Ќ�v"O�`;#@�T]��b����"O�L��x��p�P$����`A"O����
�* ���+�� ��x��"O8��㗾$t��rbD$hf�ó"OF���S��q��ӓjs�}Zf"O�s�I �E̎L�4NC4N���(d"O�p��!E"$��I�k�� 0&"O��5���i�"H8���ASv��t"O�%�Ga�@�X ��5t皡��"O��0�c	� #�ʠe�r�찛�"O���7e�KĔ��%&V�?����"O�)ؠ�Ո/H�����H�.$�"O|���,S�{`��G	M�@"O��TY�9T��C�Ґ�R!"O��
���e��\k�lRD�h3Q"O��`S�ϼ���3a�ìE�~3"O�ę���'>M´�U
c�^�#�"O��g$���rt�ƩX@�h@Ȥ"O��A�B�1�\��%2kL\Q�"O��JՄ�_��!Ӫ�="�ބ�"O�pS��1:��H�j����a5"On��!jڻj��R�h�&G�����"O��<&� �1	��o��3�%ɤ�y�),p��K��92du����y�S ���M5]��2B���y��3�t+v-D�M�������y�NGm������Ƚad�$K��bN>����#D�c�٨zI�p�E'��KG��"D��1�R>g�Z����Ϳ"���$D����c�" |F�q �J�\_�:c!"D�$3�ܻ&8���#�����!q�;D�Hە<7��xk�.
p��q�PJ:D�@� ��*����Ulw�sN6D�c�ۺp$<�THշZ�wB4D�4"鎽V�,�*�H�	B�Y�c�-D��Y�M֝B���QcN�&z�u�g 
F������ �MQ��������"�r��4"O:�2�ʁ<� �4E�I�(��V�'�ў"~bE��x�\d W"�
��)�ud���0>�O>!�˓|z)@%O-M�!kňu���'�����ա4���Y���R	8D����R&Z�l�2�L�l`¨ �`7D��ѯ�t��P�
�2'7���3�$<�S�'&RliRc"s@\h�A��v�$�����s�T;rEU3D���阦u��R��:D�Që�08� p�5�.,�ޙY�<D�T"T�}`l�9"�߭'���#;񤥟l�e前��	Ղl3���d��o�d�Qvk
9�!��sք@�K�*�z�9
�y��c�1 �)�i$g�dc��y�TB�#�w��y��	.}E`��o�"�ɃC���2C�I�A��:�N�nQPd�r��3QyZ�O �=�}����`��ؘ�KՑh�)��f�<�WA�0��$1]� qЍ�|?���'>�I�<Y����~�ņң��с��#=
ny*֤�{8�$���<���li�c��]��@����v�<1$�K� Ԁ��f���H.ɹ�%�m�'fb���)3�6)����9�5BdŞ�0;�7�0}R�>%>c�d:A-����×s �D���Z���<E���x@�A��!�"R`�8���N�EՐ���HJ z�j]|c��
�a�{��l۟@S�"�"��){T���|ZI�� �N���V~�rG/�U��Xbu��<iL]��|$Е����2�� ��c�v�YG��S�=��탒kX aʍ'��(h���)�� !4�TK� ��zz�y��\�t�����1�PI�q$V*f���t�ܾB�I9�d�÷!��X&r1�׮�/P"=��'�1Ot�M��DB�*լ�Dp2�.���t�ȓ�2`��N�x��Q͉xP��ȓ/���bO�,vL��QF�$��+�	"cե�\��7&;�2Y�ȓp��ل�$/�6�C���!#\܄ȓXbt)�&Ƒ5�ԭ@�*+���a�VղP�E�$xĥ�,�~y��	1��1&�6TB\}`d��-r����ȓR)^��`b%e��8�b�r���ȓB��0r��-(|0 ��>0�J��ȓT���� ʕ&���T>h� �$����I6\H	h��� uh���#)�C�	zkN���A�/E���G����C�	�S�b�{e����8����8$���*���'�a{bE�01���b�Q#H4|<�u��X�<	E�� �����N���l[T�<�b�S�Ҥ`�]���Y�Ԥ�M؟,�B�8@"�]�I��YPƆ
��PI�?�ӓK2�0Xe'�O�:�3RF�=1�j��ȓ�, ��
Ã���(�É�	��Ѕȓ�taH$2I�P���Ңo.��ȓ6�tP����=ڎ�  ��9�"���	�'b0��,;r����Ssq���ڴ�Px� �}��I�-^�0��)�G��yRO���:p¡�½)�����I[���'��{RŞ rCB|qg.@Y"��y�VI�  �牡,r�9`���y���#V�����m?h;$�{G�I�Of��hO mC�m��4��EP�f�J��U�b"O��;��&,��U[�C G��\"3"O>Ȓ$l'u2"\2$" ��ph��'R��C�C<���0$=$x���� P*T��'��'�d#}֧� �$:�^%P�΄��ˡIF��4�'�������$Y	�*�#����L
4�6D��T���<��t��mf�p%C2ړ�0<��A�F���'�(zZ �!*�}�<�7�B"T*�8��E��(4�)4�ߦ�H�^�4��IP��ĸ� ?����$Q�=�C䉬,Ѵ�J�-\�/3Xy΄5��b�����3�N�5Y��q ��0
��B�ə�X+��֡P��)P�*�p�.���d���A��Q�_�T/��`g8OB�O�ʓ��Y�p���+{P����=ZJ�I�ȓg���LCs^خ;�P��%�	�HO�O�����/߹vTҘ���M/{�Bei�qo��S� <�ĭE����H@(� =�ȋ "Ov�t酱;��iQM�=cy��"Ol�	1�1K*��3�T�ʠ� �'j!�dݾA�h��Q�E�y� (91�@!��Ĳ'�S�vkp����L<*xt #�C�	�j�x�Aa���s6��~���I���I�)�L<��8om�4��mΞ�Z����k�<�`�C:yV�A	\{,���p}r�)ҧZ]R`)�ݎ#@���%&Ϊ��ȓ;. 0��X|��@ץ;��ȓBl����c٪{�Y0�'�
$��iܓ��쑅�1��0��HNM����ȓN��ѵ`���ǌ�]q:��ȓH�Ȗ�ߞ%��̑�-r��	�ē�q�qC�K�|xk�脠(�hr��ii���J�����l�|* I�o�!��D�<�JXkB��"_�1�n]0s!�B5	��H��焒%B��AC��/c�	]�'Q�d�=�FL�y~$���P
T����R��P�>�ь�2���.�\2�p灉V�<��b��I���[@���҄�&�JV�<a��OsO�p�Gڕ2$�A�*�Y}S�����V)����� _޾=�$�ɬoh�B䉒+�9+���y褥ӶJ	�~�������|�w�W6"$�R(Y�+lP	�2⓵�p�2���H{��P눐Z�Bԙ�"O
X��,�)�N��Y�Y��"Oz���FM�>oa�ר�YL��"�IU�����{k&�17�^�AUH豱C�����'扛�H���!H�z�R &$����`� ^�dB�	1bz0���b��?GX�V#U�Y��B��.������L�#a2)A��M�)ZΒO>�=��y�ŋ�!.�!с�L��l�b��0?�(OX�9p�T;u4�룮��N�x"O��C��"IB�����bH�`�"O����ʏ	���%��,:��"O��b�)�+">,�2���$�|-K"O`E��T�p���6��lҐ1�"O� ����kx�����"8�2s"O.�˵'��m���'�*��"O�a���q�]� �N(>�ZY$"O�JJ�1д�n��D�e"O�Y���֙*kP�����"d"Oh=��(E�i��}�`���_���ɶ"O���6�R�h2z���B��V�6|k�"O(ʰ���eHLS�֕nO��C"O���bOƸ�T� &!\?�P'"Of=����B��d��8��p�"OR(�&*�C�0��ah֙l��"O��aE�S�z���"���.:�"O�``���:����&*
����"O� ��֥ѶE$@(��D~Ԙ��"O
9�Aj�Ef>��c��6R��4"O&|G(S~>��RDö9l���"O�HqS��}^��[�-�FP�"O*Y�1��,*��U薏��X��"O������]�ڠ�M��"i�U"O�$�#�I�V�X]�5�O{'�m�2"O�Łp��)5(�S��~��
�"O�
 o�6M�2��M�1QI��R"Ov��!]Cxe(W�J'��(�"O*�P��M�8r4�aGF#0�<�+a"O����#�*� b'	#a��k6"Or��G�!�j��唎s0�,�@"O���4Af,[!"S(O	6@��"O��j�g� !���)v�?	�Ub2"O>er��ޘL�0�CW��# d�"Oz���v6,�JLG���X�"O��B��+�譲��N)b|�R�"O� ���I�rӂy��X�H����"OrM��
�
զ��.Y�t{*��@"O)�*J)^z��pCJ8D�r"O��ٳ�OH0����.U���F�0iz�H:�>�t`Š91O|Be,�4M�b�{��(z��eۅ"O���%Z!rc<|�rm���*Z�"O�ʦ��L���#!�7?8	�B"O��q�<H[�Ɉ�#�n�Qt"OzX�D�[�o=`�{�ݔP�\�`"O�8Q��6!]��R���J���"O �jԡپ8��ܣu`��0���J�"O�ݚw��=)Z��V.�|~���"O��d�S)���@l�?(%��6"Of�J����7�̱8,ԏJl�j�"OL8@+�
[@�@�I1t�e��"O�1�ƈ/d)���.0r��5"O0<��e����@mZ�}#"O���e��#cD���I^��c�"OpT�Aȼ5?�}���x.� `R"O+��J5x�B�-I.�T �Q��K�<�%J%9j��5T�y��	���h�<�U߸ry���Uqjeia�g�<���	�e؞<�@�
4��<ᒮFE�<A�����z�nT<K�t}ؖ|�<��!**�*�;2�Y��AQP�<�e(�)s��K�lD�.d|<�E/�_�p�G�9d�a}B�L'M� ]�@��3[�n@SW�J��<�`��Z�hLKg�ʖ�y�e�22��/�I��H+Sf�<1cJ�*9f騔�V'"����Z�	�OG�q�ǉ�6cD�J5�S(��@�-�	y�搸��?7bC��cK�Y�G�2��4zp6D�L�	�$�"}�y!�Vqk$,4�3���j[2չ���Y���CC[��B�k_F� ������"̺u'n(;Ʃ�
V!>HЁOZ�o(Ĥ���cA 1`"b�
]Th0�'&ꮣ>9D҃'&���� F�.T"�N�b@ �����Z�����M̏^�uq��/D��R��I<��	J���"
����F*D�P�s��!9��i��eƀ$N	�=��O>Ҡͻi����7)!(Wh ̎bRXɆƓI޸ G��m���0V�O�>�zy:`Ex�m�
a��<�C�V%Kڴ84'Q�l���=�W@�r�$��dvאNS�a���'ry*b#��|ۀ�Y=�y��nK���(R.ӒJ�LU���y�iX�'�<9�4��%i���[�<OZ<( � {9V��Ň�"�:A3�>1���)B>i:��T� �Q�oF�v��ے��%%`H�`p �&^���*%j܋&�d#[`�#�b �I�zfP ��˒<X��>M �f��2�t@S�c]�`xl1`#�$g(�ê�7�	0�fF2�eHr��3��S�18��?�}ra��5%|�m3�-���uQ1�ڦ�H{��^���dEx��M��IŨd�P��,ģ�����;u�9!&i� �^b�@�9#��c��g�B%� �!	�➘xJY</I��'-v�gC�	7�����D���h��@�<?��E	���@!�oy(C�2��� ��"5��-A����v�;$!R%!1�X.T��Rψ�kX�K2b���'��]P�H�PAXP �k�u�\sU;A��%�E�J�|��'�s��J�
��Ո!�\�e�����3	�t�0I���ם내��@�O�\��-ӹ�<��N�;|��� k�:��g�⒨�� Yz���\�W����L)h�3+ 0<���g�
/��(�4��9�,���K�|��BnπM+jʧ)�r�YBJ�˴⁑4+fʛ��d�(���d&5S�jzu�ϓ{/�@	���M��~3剃 )*�S�ˁ2j~�Р/(��)�:4��v�ƌ��Ң�����k�1llܠ�@��.�1��	A��M�f�I9=�|�5,��n�:Esg�=l%��sc��Y�d�F�4��/Uv�QO[2J���� � M�mx��à8��9�dM��6�E�re.��#K�BN��	�o²jP�]��!?���d̜�(8�&�i��8{f��s�h6 [N]9�Z��n2(]4d�o'�!hͻf>jD��c�FJ:`�O�F�3�CL��}I*R$���,;F5�H����,Q��H��\�cD�4��jrQ���	¼;@�;��� �>$!�b⮇�oT�Ӂ��NP����*!�f8(P���D�VD��h`�L�t�=���2�kD&�E8萪O��6,"0��<��G
͊��ǆX=d��-
+O*<��X�?�R|����nx�t��LZ�J��JD��9��ɶȪi�tnX0;�BX�Q �iq�X�Q��M����Jݎ}�`ahEϑ���� �	N���ň�HR�1� /� ���	��	Z�A_26�	D�9�5����!%��'���|=�s���v/�L0��0�n,�W#@�A��	7B�')�)����z1�3$�ϐu)�@ "�S"����\�t���30���ɹ�D���$%�,Q3@*q�z�����~� a㺍K&K�1"��Q2��ܶ@�H4x��a��5sb*�&��}�mDe䰝Sk~>Y*�,ܴE�R����UP�g�L���:�$^1O:tA��}T1�tOY+M�q9�#���y^�6-	R�$1�4�%;	|�
wK_1�d0�G���KTX�3 V(u��930� y4ۄ �'=j�Z�y��U�Rش�@�L�F�L�2 �'�^3�-ۏu������xuZa�'ڶ�x��Q<B�X�R�-�%�D��h�˅
E�Dq���S�����Z 8�T�U�{�<�5?���O�@E�w����Fn�G���+AI�2�`H��>�%e_0
O~�1��A90�ICg�Ǡ]Z�	� ��P����C]7s�Z88��ʹgO�,0�de���:�"O�)��E	_m M��	��^�H@Y�o\�ZT����ѧI���5��P�������u'	'&v%q����+��<U�^�3M�Z��q��|��ytoD�'���z6�V?�R��')ٹ}���Ȩe�n����-z�����(]	��:��׽	�Dܲ��@9ES0�A�.�J�y�h�i\�8��ʇ2ጩ�5P:�
�*�-Jt���H�!�; :�ۗ��O�8F�w��S ��y�z���sx��q����Z"�$"P@� DR��6"c��ubM�B9�%L3l+"�9w��=_(��`�A^�<��47�RP1B�G l�rj�<i6@a1�$�:��x�L�pL��/vu�lA��	�n$��$�&Z�������X�vB��H�~Xҥ쏮u}�@)qNȖ�yW�
4�tx���J���cT	�F��dBX��q�#͹��3��:Xn���&dўjhԜ� �=D⚨�L�jK��&ƌ������8]e��%�lX�*�$S��sÀ2Y^��g`-��X��0�1|cXVk�����`N�,;$���c�ȍBڞ-�$��2}�Z��3�Z�:���@tM�Kڐ8˷�I�?!���pC�O������v���
�Έ
u4,�t�	+t�`	OY.4h���ǂ�H�������s��j&ϋ}:8s&+F�<$ r���{�h4 �JШf�ўĚ1B���p�F������,"��#��9���r��;H�I�3�<��#�� �S��A	!���p��:�ļR�*�B�@����1���b��0ud�4xEi�����;OKU��U����?���"/ѱwa�$`eIyݡ��C�)���s&�m����:�$D��Bæ!p���W����lyP0X �M0���+
�My�OH%Z ���
�����A�@`��@�#W̈p	^.�\D�ڑLN)B0��	��蒉AAb�9�T�� X� �Va�'A!�EDPXU��dM!o�d��@HHhD�U�'VZA��dL#kjm�'�G;��c
A�N>����WJ|�HdcM�g�
�$�H�vQ�'h�9U���C���'I;H�I����O�b�8`d�P���<��	�K�a�돔J�p�h�D!S�����*�OE�@�$\�z��U2��t��4d��O������!Б�q�GOF�\�T�y��A��#������L�8egʫuV P�rmnӂ]
��� ��`N�/_��uY'&�@��OU�\����ZٌAb��+>���%�N�x��@��,Y�?�ʃ�ߡ[%�ر�8���y�#���'h��9w1Ol=��
$��QG��}������'tրR���wcP��`ʙ_~@2'��&
�ƀ�{��Y ŗ���R�G�"H���q�H&Q%�1�C剫!p:<�d�_*ĊlE�	}��p)"�����i#�D�$��a!OX)b�T���4dF(y����m��aףM�As��!dH�|ʲxِ�Ѧx�Ā����*~��O�Y˨�,6��"=��'Bg�0�QN�Kp�"C@�os>X6A�9l���"/ۥx��JSC'Ekµ��X ,�En�1@kt@д(�Ox#��4M��)[FƅO��W�Ё����+/q�i(K��_t�6�ԺRq�1+U��5�z�`C��X�SŇ��RW�l� *
5��	A��;M)�T�V�O*���M�Ukb|���ş@��b3Nt�1ufǥO*�TD|�H��4IXX���<QDҁR��9S�p��4=D6�Ed]�B���35��2BL|��DR=UMƩT�:R�r6C�e�YB�b��>��H�f��*�kѦؤ+�y"��:�+Q�% �5�`��N��h� ��="y�Q�����9�t	M$Z��� �R'�-� �YI��\°�'(a�� ֐+�0`aC�^�H)��G;�ў��d�8(�]��D�,^����(�n�D�֫���AΔP�P+� O�`�:�+�٦͑�Bh��,U"xpc�M�-�$�a!1��MB�I�3\��袎	9?zY�E�`�<�ʎ
,�3#�&Y�Xb��Ĳ^��Ȓ.ɚ:8ty�ū��w�L�pC��>r� F��088�qG��7����1 ���y@���a�x����$E��]�@��t�4ݺ@�I�q�F�;�Q�?�a@�N�-�P��<�I�S \u�2њ �Hu�X�o��Z�!��;_�������>~�%�E��+�a|bI,k����kf\��`# Lݕ3[�A�@5\1B�9��7 ��]!�Z�wxt�#T�b�p30,�3X�qG�Ƿ߀ j,Q4��KH��!`��1���'����g_�@�h)�'��0�wa
�>��W�	V��`h޴G�>h	����[��yr����ȱa�C1z�5���]'�~����O���fk̾Un���D�Y�vt;t�|�ĆX�r|+d�>Y7�Z�z��C�z�|�#0S�zB\��ڲ�2�ed�b>u�w�ĥNԠ9C��QG"�pF�zFP�T�$y!�m%6eJ= �A�0aۓ�|�̩@�6q�� X#e�N}2æU�`�ȐD�S�>�2�MV<��@R�������݆~�li�	H%v^իQ�)+�azrkʘPZu�r��QX�� �.a���1%��5*��]Kua�	s2��ʚTRU�J߷SV���gB-`���5�Y�tL��b�e��!>ph��J��Px�l�:4�(#$�#�v5��Β<{W�5rS�
�1M�T)����>�ˇ�!3�DO'�n�7N>P�9bsaJ-,�:jM)H(4�VӺl:����(4�,��@�[3H��X�J���X�ڈM�Z��IW6}�<�/��S����8v�nI����#��hU�O�J�Kg�6��\(v�P�(7iD'S�Lx��'X����O�<���iβ�Ce�)�2��ʓ�N��$���:V��0e�"�@�[��Uc�Ȥj��W\�JA��=c�NW��3��y���d����"�5D��\⃊	.rz�v�(��lD+�&>���ra�)b�����H�6B��x��
��vb�R�N��O�ĴsV����\Y` ťq���.�L�>���C�P��=9A�ؠc6�0�>�>l�j���	*�a��0�ہHB�W��i�i�#e"�9`�B����H�M�!*ذ�/��I�,�Ódk�a�{��y�ŁY?A}P�3�ϣn�}�D�&&�P �Ճ���D��;h��4���@�n 'D�.��/	"H@�'��u�X�3��҄!T4E�p=��Obx��	�*m����-����%�%�^�:���h�,B�.�딏i6@�1HV#c�|�@�'ި	�^٬��d$�u�٤\!���n��"`�< pR�Hו*>���@(�^<�c��� �n]�q�:j� �Z�i8P��V�+:��F�*���W�W��]� B�@��������q��L']��PDʧ	�J��@�'b�@B��̾@�t�'N���D�ʛ{�T��aګqXD�䌛K`p��v����b�\i�l�1�%�Z��v)�m��& X�1C �J��bH1���]LjEZ�f���z mF�6z�e��&pc��K �nhyS�d�|���ZWk������ʍ$F�9 \!%�U�$O����ڹP�zIB#��T�\�1�I"}�UxQ�:�'��$lȞ|8dJˏkDੲ�פxw<@Ҧ�)�C�����ad�Z(��Ȇ�cMZ9�0��%S:\J�ţ?�`t{V�����9���&�V4�sȇ�gGB��LN�!V6@r�>�d���O��d�1��H�@ ��	 a�b���/����Q�C�+����F�9J H��Ua5<�����fi|�C G�H�Y�#����R 0^, do�d=2do�G$9#$n�)h��X�ǪN#l�N�P"Ѳ@����.O�q�JI�5��RU���O+b��aMB?x@���S�����B)�6лg�A�(�,��p��I$x���MC}�n  ��C�#�<0Ja Q/f;8��I[?4
�(â�b�#�	d6�%��!%�("���c26���� B��!iKD&PZ׫),)H�z��2���hTbE�t��#<�n��QPB��u��f#v���	�7;�,�cwς�06	"%BG;��I��jC:s�:8Sc��W*`����5>�6����23<
EB�8�����Ɓ�v=p7�[2u���}�L�ohMzF�F� @`��iޛv����$ @�	�b��C�1o�B�9��:	�����(7���.T`ܸ�S���
�l�2\�i�X�i�����y���D��yzf��W�n�V�30`�	�-�$blk�8Z��z�L�iY[����BG��ch� �q�|X!2�(��胉+e�uGN����%�`#�|�*����u�d9j���#5ƒO���0N��ȃaa1o�1@���	�t �WJ?�9��Yw��Ɓ��aܰe��n��D�[��ÊO�_�~�r���&�V�C�D�>� ���5U���<��OF�1_�����4�U��E^�x�V��V�'4�T� %;]��w�ĸk�ze��c�7Y�}��e���L���+��
?�d���9\�ݩ�л5�j�H�J*���E�]�)��q%���#U�8!bZ�ɱ�n�..�l���D�:m�Dx���\^Ų���-J档���Dr͠�ő�(�x��^;n�Jd �@V_V�̒V�ʇiUv�ub��р=R�4)e�ȣz�B� �'$�-���MR��I�?5I���*`�������L,�I',�4{���
��̑��݅r��I��<m����O@O$�iH��6~�OTq��D��f<�8�F&P�z\�hZDT[Gd� փ��mmE���H&gFPy����d6�ӶƑ�z^�pRF��ZF��)J12uLd���9׶�����
7��<s�g�Y�:�#_ܓz~ȩ��>SX���	\�%n �V��@dr�e��?���bbf�h�tYS�!��4\L�҃�ܭ'c�&o�6@T:#�U�:���Jҩͩ+Ӻ<j��>:��x��%d���8[�R3Lk@A��e��!��鑱E�0cb0	��F��H���1�\�B��Q�L}�t� HI�}:.��-�Pf�D��5��l��0���"�(�n�H�`93���2���eJ�Y��a���ֲq�	�j�;_��%�ܕM�p%�!�9�L��JINL\��f.6p�c�5��L�d$ �,��[�b%?���j�ONX���.�$яb.jx"�CU��(�Gj^�E��xV"%V,�a�����rdڟ>��AN*A|�ɩE<��h.$@��� r�P;�(�0���5�]2D�^�#@^p)����HOa�⃞�M�b��o�� UBə&�"�11�1H#|�q�U/��Q"�R���F>>^�0�扽HdDX��^@Y3��ٌ{��ⓢɺ�����'���X�n�zp��2%���;B�X���P{� �b/nr�ݥO� 1 �_���C'��j��XD���Θ8Y��r&�<G�z\�΀̸'<*��S��'r����@U�ORV��)-�`�G�-6a�6E��qr���RP�h��Iv�g�dO3gF� �� V%��]a�LjZ�$[6�J3,
d�X*O�aE��O2�Ð�F(��a�IC�����"O.���ɕ�&��iC"E�#:ƽY��'�X�p��	7&V ��I3>n�!��.S�r����g���n=��D�	Gx��0��� ���)C*eNވ An��jun�RC"O훳��-\��Dˑ8�"O2I�S�F�\� ��m�.	h�14"OXA��]�n��,ÂkĕF
J%S�"Oz��G)�0G��U��ʓ!��P'"OX1A#���rr����càZ�&�3�"O�D��&/�(����7��1"Oj� Ư�,2Z={҂�L�Ќ@A"O<�p�N�W��q�ҽY� 0��"O̕	Ѡ����BjY�4��3b"O<����P��4�R�sv���"O������ȡ;E��ej��aB"O��X���rb��(@.K.6�\�:q"OR��cS'\�#���Y���3�"O�����*8�W�A ~�J���"O�Y�`4i�U��c�+�R<��"OtA�@{������u~��	�"O�E�5�_�g_�Bv��	GP̍��"O�	�@ȝZ�ܑ�䙀W��LXe"O�9#�l؈	��tс:�݀�"O�[kG��R9���Ē�h�1G"Oر�!.�0-������z&VH�"O�m3���<<�T�I6j�:,0mٗ"O^ܘcԫOt\�j���
��"O8�rJ0u�Ld[�%�&}��y""O���0/��9�Z6a�K(�T8D���$ΖN��\�թ�0w�*�R1�7D����7|��(��W�o �Ғ))D��Qc��|���D���mi��8d#$D�@$⌆|v%�Cƶ�bT�%D�4����y�FT���%cqd��$=D��:�m� �ܵ��J/&�&-��?D�L-R9�V�Ҡ[�AЂ:D�{���6_�xԛ��P,����>D�(��	o���k��>�ƼJF=D�1�&�7c��� �R*�֔CEc,D� c1 ѩJp���P9m�R���m-D����*��Oq����L�@�����*D�Z��V�K��9@ D�-�P �/+D��C��Ь��3���0l�,:�-D�h���.f�!ȣ�ְz,�B��(D�<K0D�>$v�!H�<1�A�u'D��qA
ߵf`	�)['2�:��c�%D� Q	���� I2`B: S�e(#D�4��hd@ى����zy�hQ D������/p�P�Ӱo�"u:"��t�>D� ���i���B�"�J�:�p�A!D�����w��;�)��2�V��a7�=ð>i��D0}d��7N�9J�4���.�ux���.V�K�2���n��<y�ڒR8���%^?X��JAw�<����x�^Y�#Nx�I�(�p��0!������c�x����*zP�tQk��/J��aL�W`�C�I���a�&B��<��X	LN)�P�"k$���a�Ÿ�4�3�ȿ��¡ #�������N���
e�
 �`��@XB��m�?V�`��H�F&�Kń�M�r��-M.�U-� V��}�5Y�axba-h���$��
E���*��ֆ&B^��쉄
X<9!�M�C��)�':���܋��""B�1�>�s���
�yBk(!*f�I���(��V��K�'},�.�0(�fM��]!Ce�� SDX�R����I�ʸ����{ݼH���Ę����4l�)5`�ժ��49D����
H�̴��,{�qO��eNۖO=�5�6Iˀ[`�����'�~�K�����!G�6C��5ᒣ@!H^��#�a̭Y��x���G+5(��>G�Ȃ��I,}P8eq�3O����G� `D��!���v^d���>c�"���WHK�6\��Tl��4ςRnJ�x��oZBV��kV&����%Ü-8	�?�!�ŧ �� ���,�g�? @����O(p��%;����=�(�0E9N���2Qɨ���!�!0T���a����		}qؙw5�t�a�J2�P�ABD�(f�C�0 c �Hy��8���p���/B�艋�$ӆ��9�u
�O��2ĉ^�	@(7c���Fu�q	A5\�,�C��H$:���r�*&�(��� ��m�O� (妼J��& �M??q���4�a ��ڼ){�$�ܕ�����`���CvcR�A�ҸY0��*��Aϋ�e4$��i剼.���n��0i\8��O,56����k�lHR�h��ц V�I�Aܞ��a� J�Ա���>�x�)����%�P���u�ݛ�z���Θ�Kwd=�螄uܱq���yb�s��a�᜙�p���^?�[T/��S�HS�v�:�QiD�*�@1�ϊB�,)'
C��D죂a����x�(����
;�T��c��6-Y�fQ%dp�h6)_2G2(���� g���`��!�Vp@���'az�@vI߲��DI�Ek,<�v�ڊF��1�MF��ѻ��m��� !��1�`6-�9{�D�e;AHB�?e���P��y� p �4Y�n��NŎ]4��k͎*��t�EM���Bذ��X�"��b)Oz�#�׌e�h�3�Ĩ:d�䕿'�n�ٰ	�	cM��PG��=�^�sR�Ɵ�b�(�q���c��>$�l���iV�aJ��0�(�>�����Qd�H"��N�*�� [�#����'>E�@Nj�� rf�ԇX>�>!���Z�P�Pd�`�M�07ڍ�ǖ�>�J�E'��D0c�{sb�s�[!S�Vl��13Бᇇw�8��_=z4��M�i�A�@H����p�����2c>� <�cRJ�F�&9����
�;��`}R�A�i��H�GagH�A�
Ī(�HyR�#�S��H=~�T��Seԍr)��8�@�<PŜ�'�E�9T�'ǚ䛧��	?Y\�@'�X	P�CE�_?v�(�yg
/_Z��F/]K��3w�C�r\�����m���3�4K�
(���@9O��堁�d�x�b��&�4� P���Е��3(@4UP� �s�0��Z��,�B䓄)K'��"C�H�jמ	g��AI��&�'� ACR�tJ$(:s$�`�OȠ���a�!z��@#��B���S�[Hb9�')M6g�0��A	�3�����W�������ۼ�.�
ΊP�����5O]��Џ<������<1T%��@:���I�u������łX*\YZ�0p��,��HP�^4��&1�v0[�(�O���@��]&Du
#�*�ę/ZXj-p�a�.����q!�8����{��{����(@��Y�7��s^yYVc��P�y���b��ꔣ�`?�ae��z��}RMC�}8��'Vypb��]�F�Y�d�'�P$��Ob�ru�&D�yG���$ɀ�W�R��0�䛐t"̑���0&���@��	ǜ���B��ȓ�䄲�쏹_��4K@��G�&����M�謓5���$M�-�������o�y��A4MI��6����S
@�a�A���V�f��3��'�J8���O�0��hC�,ݯf�"������C�O�u���F�ӛw4�9���ۏ4��HGL�,c�:��<�*�'>��*2��z���w�A�'=D���F�ZO2�`�Oc���ĝ��QB"�Nz���x����|nα�3��> ����w��	#&�৆����<Y �έ6�n�X���04�$	�mF�<aCHV��|$#Ӳ�vT���0�z���21�<%뇽i�ġE��::΀�	P��6^<r��'�0���d�9T��es�/5U�64)�l@q'�{5�_�3�u3U�C�
d Q;Q��y[�/��W�&q4��t-�n��B�G�
u��L{�&
a~"mA���,ঃP()f�`�I?L��ݒ5��9)�� �f��thZ�]۲��W#Q-!h�P i��I��O�t`i�O<`Y2Ə	���aIt��,�QA)F�M���'#�8)��pn�m�̹`���n3�-QǤ��0����]�0�4���C[qK@���D^;o�ܑZ�I��r��r����R�vVL%����B
~:'LK�Z�<�@�ՀI`�cd��r���Ui�pZX���DC��G�+.������B�d2F�D{CQ� ���"��ˬi=����kP3� ��V�����a�,S@Ry���R�)u�	��J��'�v\�� ��S�����ᜭPH@Q�`,' X�Q��D�Qo�A��/T�~�h�
�(�<Ն�*�H��G(�)2���y��D!Sj�U��O�)�u7
L#1x�$r���v�|`FI��M���_�U��`ϝ�����	T�,�(��C�-@��ِ�*�J��J<iC��OD���C	�1����7���5���dO<?��SΟ>y �sslQ�MA���I�0����`��3��
�i��0r~x�CW*��	Cf]:��\;S��];`���k�1EaQ�KT��;��|3v.Ï}U��Z��P�M���f�$̰��.#��`aܷ��C�ޟp@l+	���6t��U�K۰ �jI��A��ʝ��MF�i�Q���v���~a�bH���޵�QM��m��%[`�	g�H��Ҍ�"��`J�MF1	�܄@�MĿ*���K&�j���f�F胢l�?!��pR�-�1�ތXfG�
<Q2`̀.��ء�i�7�Mc��%C�y`e�=(�V�W�42Tx$��[���3�� k�|�8��2|TAv�U"M?#e�٥n9f(;��U�cPR9��aipS쓶7��[wª�j�)'�	���a������уK���M�0(�4O��YP�ˁ�8�4(Q�_���E�
[�������A�شT lH�,�+3�
����>7}����G��6�*#��Z��=��o��&�^����A$�D���R/d~��͎�d��"ȵI� �B&�V#9���)E!�X��)R�dj-�3��a��b�bL���q�lA��a�0Kƒl~��l�c�فh���`f��o�*E�#H4:h�	��j�%C% �´�e9�!K��P�Ӡ�jiң�iD0l�֢� �?	�,IpBx��dBo*�̧@�(p���F��d�9l~f�;ڴ�c�C�{��P7��xL p��24:d��W�	w�����$�	��##!CB�}�2MHC��)���;0d�6.ې�XT
�(G��#�I��)� ,ݘO|̀�e�6:b0}�P.� �ƹ�!��)W�Q���
�������Jl��e��=o4}��4qCn]˲�߉��ل�Ԧ���x���7/�����I&���8��5,�[(�n	�\T����c_#H�\�r+Q�q뚌٥�K\4������(�1�N	]Y���%�L�+�i�6�SsÅ)�s� :S�uD{�!�O���HJD0A�B sA�d�!��n�VN�P�%U�-�T,5���P!G	*!z���Jp�RP�о9ReD�vV@-��k�q� ���OU�\ '`�EwȊc�D!t��+&0OD�I4��-:�Z$"����g�Lg�ԝGrؒC�D w� �k��s� ���AnM�#�ȥx�$\���٣�~bN�
�0��V�~|v�D}�6_x��������5B�� �
�Y��W9ٸ�����?X)�Qq�Q5Yr����ۊ~�����Bٔ�7턪Gu�H-�5B�Dd
�aZ#V@�RG
�0>��":O�T�W�XT����O��0�$K�'���Ł/*�4a��nӒh��τ1�0���E'/:�9p$�	���!%�-�L�هK�! �tb�'[��*�[G�'8<�0%�R)ar�uk�HW�{�Xу��S@�V��;kf�:!o�*z�vtrA
%S�谫V搬�r���wC�\�uF�V�1UL
 O����M>u� N����M��k�i�6����V�)�~%�Q@ĕC�$�R���^J�����U�JL���+V]���X^9� ��C� �����	�9��΂�~g%�Vh���'f-�f�9	���! [�o�<��GF2o�.���Kϫ����%�%/p�5I������u*�=_�M�rǜ�7^��iq�'�&��fGN�.Т�`�#�'<�z	��n~�h�ҍK#0<m�Sl�N�(���GO6-֪�@�Ó%9�b=�$쒝l��D�R��t2���*�>y�'E�P:���G�Rup���!i�|�3�U� n�p��fr	�놓8�F�IbF
G�Ta8��n�d,�CJ��!l� `��ϣ]�������V8!AY8�Hã��=
rDa�نi�Sh�k `Y��tk���ׁ��oGV����n��87���x��dĹh&lqp��
q`��O�@H])��mPe�-h�y-8�ɶN���\2*A.�!l�9W4,M�Є�Z��-�R���qC�<�
=K�+G���V)�3�^�S��0Bdl�J$!X}x���W`6�b�����Wp��0��ȭ{	@�)�k��^�n�(ՇY	&��̲��Ğ0�v��EVSy��«Ȭ} P�0Qa��m�HH��JΗ4�ȸ2ǅO���(���|�y�'��i��sd�D?gX��я�$|R�B�f��D�H�sF�T�r�)"�Įa���n�=bV���o�59��p3�V�Lg����*B�z���[�B��MZ��O"L9�vK�S`�XQ�dZ��th�$�?V�"Q[U�i�h�b��*��H�gJ]&o�r�"`�5*�ɘ�)�D�	��JE�jR�T?j�CV�� �Y�t�P'�_�}tXq��+�Xy�5ꆌs��]�w�A�0��d��v�=�ׂ�	2�<5+ ��DB��:��Y�z'*�#J�3��<	�c�l�VՓ"䀂zzX�
��V6N5�6n?,I�'�-���Ku�Ԃk�N�Ӣ� ~~B�
����j|�pu˗*yJ�)���T/L��j~�@ M܇T�*H3��|<�˕�����IXu�B5Q{���'���p�]�l���e��}��,��@ۺ
ˢ��w�W�N���� ,s��-�Ǔ^� �҃������$߰lw�yt�U,Q����éj%��`�@�D�2!%��%b��GD;��B�G�r��R���'VA���>s� �˷C��!a]�J�0���'D��d�++5����N�w�dH*`��"O[&�ʂcЊ1�6U�Ӭ��x���p5#6XL�p�7;��e��oM�'2ph��$�ɦ	�r��6bT=���=,�@4�M¡.���S�F�!%�x��.�7�"���2j@zB�>)�J,(��b�q:4b�:_t
��aժ,P"�b/ʓ.�|"H:^v�?	�$m�S������)kF��Cq�ޘI� \����ܐ�dZ?���4M�R����QɌ+nL���+�L�@��ŕ\�P��!i��!%�,��|_Zy�E���@`*O�I"01Q���"J�ԳB
�8"�䘑��f� �����=Y��b-ϛ%�S6��r(�˵�ɻ$����q{��W����&$�/0������(���ɯoA��2c�m�V�M��S��ɒ��X�6��5�&*���� R�/Z�Q���hC�p�R��H��;��4BU�3��\"GJ�9��#<��P� q)JRV ���L��^���R�q���sG@E�i�ؔ�H�3�>%A�i۾r@ ��(L��D4�0�Sr���['@��j�v9�b�m}B�
 D��t��ӎ}�k���E�EH�+RC���i#�&
���\+$��2�ڽgiP��c��Hd�"�"��G,����Ů>@�y��W.w#��
tb��bbJ���DۓBp�qZ�@y��B�(|<�����*v '�B�:��B�9:�,e��bW�pY�Hq����yiB�����D����*��5��32��.BD�\1a-j�mS`�='�\�B�D����R!�]7��O6��ŉ�N���s׍>ut����]X���T��8q�>�7G^�K81�u%�N���[��¿w~�%۴�S�\UJx��m\�m�\ ��/͗`w4y[�}�ԕ�v��"/��`!6�w�.��|a���42�@x�M		�!���ESSb�C�H:	��d��@�2o�Bh@e�>1f��󐩊�-�vhDV]~�S�I���L���B.hr q�F/c�:R�Ū�(��<A���>���g�%j��)�jC E@�
�I�ip������޴퀂iT�9N��:��	�-�Dc�m[/�^��c^*%ؒ��"��O��򉔯:K��2=�.1Y�CX�O�L���(�b2��pM��a4��T�E�|�u vc�:V��M�N�S1wx@�&)��q�`E� E�<h#��#(m���A�S��$ r��6�4��)(r�X��$M�$Hs3��D*?Ϭus�N߰DH%�c�?#^��c�۴1��=3DQ Z4^-�C��*>΢mS.��CG�5#�?&D��s�X�0�1�`�^�ZF�sa/r,��`�m��	����Մѿ#
��=y�h��h�#al�m�E���O�"..Ej���"$��c�5i�lS�&cB0z"II�2�]�v �� )"Yb�@eI�4䉚Ĥ]ہˊ�?*x�Jt�۩rt���� �qO|pQƐ_QZ�y���"B�@��sDF2i��5%իf��=�V)�$h$iz�(@3 �r�k�l��]��AӤb�ˡBѩc����^���)��A�g |ت8�f,U3J�n�g�vG����i�Z9�Ԏ�xn�l���"yФ,�F���w��Q��I��o�ܙ�B�CL��uڤ,�@�i���I(����ą���	�n�܉��|��DE�t|Ґg9|#�p���$�^\ƥr܉�b��(��yq�O;:aЃ��>���ɻ9c���"�Ra�)mQHtJ�K�0��$y��� .
��&�g�'':-��Hئ=��ETl��jшX�89`J��0�V� UF��U���k�Sy�C�c�\�2-J���LläL9{��(�@��1�N{ ��p=9���#P�� �#��0���#�L�;��iR�HH?i��ǃ3}�j5}�̣1��':`���W�8ʧr�n�SlC(����-�Ky�i�=���$>躈���c�"|���#� |8��Bs��A��
=�:�!BK���$ڮ�T�?ӧ� �U�m(b�~|[U@DnZ�ʦaY�#�ܔ
&�G7��F����ŋad��4�� B�8�e�=|!�D�d@;�IʷAu�Bd�QmR@�0��p31�g؞��	5v����H�
'Fdӷ-�O(�����y2�@�z�N�R&P�N�((�����y��A�j�<if�;
(��`��yrBč@�,�x@(�+.��Ћ�y2)�p�����X!�4�PNU7�y"oT�J�"�s�͉=:L�B�	�y�#W<y�@���	�gb:�y򥎆a4�����䈁�JN��y�ǃ$���y�U4\�@���y���2�ju[�hB.}��PՋ���y2��O��C�~��Db6o'�yb&�
��qK�v��A��^��y�'��|\��a�߂SEl���-^'�y"�L+~�:$x@nI�Xb:����P��yRl��r�R"��M����3���y�L�1��4r֡��FH�r����y�"�8~��0�Uc̟�X<� �؈�yb�5W�$���Oɧy�V���J�yBn��y��H.�c7��wL���y�A[#-�L�`��(Pr8��i۴�yrn�4G6�LT�R�Z9˷��yR*�0N9^(�t �J8��+��	�ybDH=�tF!F�x�rg���yBj���܀{�̃@V�%��#͗�y��ۂ`h�|B �
�k�8:a�P��y"��+��kt�G���dP$T��yb�N�.3n�����49��@�N��'6��8E��7v��x��G*9��9�yb��*���8A��)��k�EJ�=g(���̦� E�w��L��O���s�c��M�bIɐ(,h��!v�_���y�I�)a�%M?1�a��A�<|Ɱ�� ����К`v��0ყ��c0/��*��	N~�S����1F������R&z���>�k�YN?�"	p�N���'g�á@֕"~���Ç�'"ќ�{6����ӽi}�x*��?�˱`��?ŋ�t��ܜ+
�b�Axh���3F��ɱ� ��Fa2��� �<9k��OȾ�,X��p0AA�AxJ̹�̛��k@� P����0|R�B�S�x;��<��4PA����� �z�^Գ�`E�Ք��c��-��?=�PbW���Ah@O݂r���!���$t�Q�X��) w�Q���	��:�8��W
"�V<:gb�w���IL�P��Zļkç��� �.�O.4�
�W��]��u8�|z���0P��/O�>�`O^�p��u.�L�iha�4�I
�HOP�Ov��I��O�D��b��ږ���"OzLR�m�I!,P�π�tX���"Ot�I�`C�w�2��!�M�yF��+�"Ob�Rŕ�@�0M���	��h	S"ObqHx�N�A��5���H�"Op��a�%g����� S��"O�5p�ѐ��:�&��JP�"O:L�$\��P�^��`C[��!򤚞=�&�9)YOe�i��K�!��ֿ
���p����u�p�qG���=�!�J�c��9���C�, �3ˋ�l�!��@�"Lib�\(�%̈�O��Pj	�'l���V=e��A�匃g|��'b���͙�8~T!Gf���Z(��'�4�J��A�fB��hcN��
�'��H9 
��2��m3^aF�
�'�=J�
��̼�2CB%@�8Ȇȓ?�$�i�ٖ-���H\k��P����i��WB2�/�V�<��ȓo��\����G#�d�[=Q�<�ȓ%�l��a��D�ȼ{PF�6H����Be���I9�f`��I�2Y��h��S�? (��@�ыF?�XI�k�1L��X@"OYcvdD�B�>3�埏@���"O�%��hN2n��!B%�ئBfhz�"O��E%eA~@zuM��zM�}KV"OP��BU.e�8��m]�3HH��s"O�H�.F/�"
_�vA�iQ"Ol��]�����Q��3G�<�c�"O���G,�F}��fʔ!�N�H!"O�z�I�8O���Wϛ�&����C"O,A{��0@�X��[�I���C�"O�ٙ 9K�|�:�LM(��U�"O��q� �
��8��(`h�\0a"O�$*eaH�l´c�-Y?No�x�"O5#v�O)Z��	3fZ����R"O��X�+]I�T:��P�sC��Q�"O�9ɰ�ȃ. �d1� �c+^x��"O�-�G�S5��[��\�X��"O�5��+�.��@��� ;8{Fq�A"O����A��22 �1��0�"O��D�ΣV>�LѺ�R�'�R�<I�g��g�R@pVl�j�F��bTM�<Y��݇ctts���uv:j���I�<	��5s����Ҕ)a䑱`UC�<aR�Ɛ;�P)GI�~Hhq1�Y�<ђI��KX�4R-D���D,IY�<�v����q�W*��)b���R�<y��3g��	�fՆL�M��C�u�<yg��-��и�">b���hf.�x�<��-T/s�������+s�] cKr�<6�����4J4�F�9t웡�g�<	�k��e�zh{qm��y��Y;��{�<y���?PXd)�.�IS�#_m�<�^�(M�]0����VPyj�+Dk�<�@'�P��V���q&�d�<	��ɯT�`(2�Ǌ1e��m��Tw�<A���kA������T�n��׭_[�<)��M�J�;@`,c��Y��P�<���@6e��j�M(*Ȝj1�\Q�<ٲ-�4�H���U���̚I�<逥K!�a�g	�0r�kĂA~�<6φ�$W^ݒ'�D�؜�W��v�<�g`ڕ?c�	J�L�Q�<� bL�<٥@ֶ�t����[Sӂ��F@K�<A櫒����s/D$z��p��PF�<�&h�����q	�>vź,H$C�<�,�� �ۡ��71+��	�|�<Q1,�?�P�"��+AΦ�Z� �{�<ѐ�"<	j�,]@񣔥�;|��C�I�Z����E�?��Ǝ٤[�FB�I�2�`-cקI>�6���/Y�%��C�I�3:�3��1��yib, i�C�I HHYQ��AT��J�)�
jFjC�I�p�� t�g�Z��^�txVC�	uqj�	��'^
�Q)a0~txB�8p�����$^À�
&d!^�B�I0@��Y�a�2�V�q�Ɓ�j#�B�I�etx��f�[j��%%�B� y�hy� ��%.N��F�Y:�hB�I_x.A��k�8�I���&T��B�	�n����"<.�,X:�/Z�H��B�YJ�P�\;o
� ��#�dB�IU>N�r��"��1�-��C�ɾ�"xQfB�+8����F>�C�	.PW��1���~8��U�E)�nC�)� �b�CHS�����˓�3��<RB"OVպ�:�μ!`M R�L�"Oi��a�%��٤���&��5�p"OrQ�`ǆ"Obв&\',�J4�w"O���k���,���	D"O�����Ş;���� �(G�"���"On�{�]��M#a��Me����"O �jN��hVx��Ed��f@$1�"O��
�G!��L�|2�aE"O$	��C��h����(�h3"ON��u�0qx\0+�#B��<J"Oj�Ck�J�ġ�#�b����D"O����g��,��M�k���s"OVtCԂY4�	�4�N<h�@ "O�L��"�-Gȭ8��R��]j�"O�x���̉8	��`���k�h%�"O�չ2�V�hT�|� ��9C�<�B�"O6 W�ȏ?��"��:F�,��"O cG&��rs�ak�`\�i'�}��"O@���a��>�KrAȚ^7L���"O��8�(�$+��q��]�K0@m�"OR���P>��BP��j/h��"O�u0����"	��f/КX/B�
�"O�Ĳ�J]�8�ʱ��$�!z���"OX��c�+r�*2�Y��a��"OZ���/�p?��bJ�N��mS"O���Sn�nͻv��'SlJa"O���䘐P:�E��m��|��4"ÒP䃚6����ԘfI��"O���$E�9ª���c�uX��Q"Ov�����pD�`1$!�U�xb�"OP�"$F�]݊�Ò�NXp�-�b"O�x9b�@�P�-*�*Ғ%pp��"OP1jO��&�0H�Q�U
^`)d"OJ!��IH�^ ��i�I�&���8�"O<Ԋ�ȀEBq9��zبp�"Oj9�taײVC�T C�8o����"O& �爇��YT�W�Ak�4��"O������I�J a� m�ePA"O��U�͒o��)2� G�����"O�Y �-�"=�m#.S���y�"O��O��):�!B�Ǡ
�R�J�"O���L�8H�� "��6l��ҵ"O����ҤK7n�*�"uL6��a"OV��E�T��Es2AHxd��"OH�B���3321�$̴A<��"O؍	!	R_-b�fŋ#lΞ1H�"O�Q��		7#Rȹ��P>d��G"O2��t��uPd1j!��_��B"O\��K<p\Lu�p��-m�^��"O��(7	�W"$L� PF�D�X�"O.1��%�r>h!q���P�����"Ot�a��� #`*��R�ċr��QB&"O�D��d�&^94��4��x|��E"O�="�E޾qD>E�2
�c��	��"OA�&I>�<��	�6���Y`"O�4Sq	.L�:���� 6P�z�"OT9����9�b��rm48��T��"O&�륁��948�;1�-Rp�� �"O�U�v��eȡ����M<ДS�"O��e�+ �-��46c"O\���W�a��LQ��߰�6=k�"O��������Q���1��`�"O��r��_e���bд:u��xc"O� 1�B��@@���H�)[�\�1"O��3�����Af(8��(q"O����N0=�Xǀٮ3z�)"O\e���ƅ!+��k�A)#j\�	�'L�b!��.!����#��0�(aA	�'t�����L�:?���r�\4-3�4��'����*I��⌘�9\_�r�'sR4��	ߚ+'$�SA��b���'��Pz�C�%&���h˦, @��'�j���g��K�4T���,�:`�'h��Ły0��S��E?���J�'H�rm� Hvh���#�3�$�
�'d i��E6�,T�d�.pƙb�'���ϯ+j<�9t P��B�H�'�rd��n�9A�Uz4dG����3�'G@1I"��zFu�` E��0�*�'���&���@_ =�GF^�v@��'=D��%���T�IbLs�J��
�'p"�"��,z�Йf��ewz�`
�'V$DJ7m�"!�2�����kT�PR�'�<�� \�@ie��:^�\��'d:H�4�âs����(��3j���'��y����7\�f�UjÄm��D[�'E���Ӊ�1�V�0�S�g��'l��x$��/�U���� lm6��
�'����v�[9j��ǅ3P�:
�'F�°	�e��X�O�>tƉ�	�'|N]k%,x�!/��t4�"�K�<a��8��]C�m�����YD�<�Q	�b��P��;M�D#�@�Y�<�j�����5 �^���r��]R�<	$BJ1;J	 !�	.����WP�<�7kC�Zt��ʒ!ц|8)��q�<Y�ƙ�T݂�m\�TWd��*	o�<�G�Ի��2�Q37V9S�,�s�<�tكB��m�%�~E�ԢB�F�<�@�P��h�b��I�Ҭb'mD�<qG��\��-��k��� �d�<�p�8Y���h�M �)��ENw�<!v�QP|@HCPϸ}Ćؙ�bPq�<��JT�a�����H,H(���D�E�<9w���B���p��(	�����DB�<�&�W�N�^��呢R�N���u�<���F]�&��#� !dX�S��x�<YS���(��1*j�܁Q!C�c�!��{G>	2c$0Seq�a`T��!�$	*\� �.�)>Pi���۴�!�T�_����g8Ezp:Q��2�!���8��X9\ֽ`@�CAo!��(C����/Y`�8�2�!�,8!�$��\����D�m�*D��� N�!򤞢[P���
�&o�����/C-_�!���<,*�J⩔:���GгD~!�D�h���׳C��$�Є@2
!���dE:4
�L�=\��L�d�ټP!��T/l�"��UA��~������!����d���)���;cq�"�*_�I�!��тh���I�{Q&x�0*���!��[�l@2CZ�+����'O��7�!�d�J� �  �P   g
  F  �  ]   �&  X/  �5  �;  5B  vH  �O  pV  �\  c  Qi  �o  �u  |  ��   `� u�	����Zv)C�'ll\�0"Ez+�'N�Dl�6x{3;O�1"�'"dE�>2��EN�%�D�j4Ý_�ց�Ф@�n���#!��a�w����CG�?�JS��?e3�f�x��x���4~�ABA#��j��5��Ėj��]�s�??����ƞ��u��|@�t�'oT�ɡA�T���,w�Ɲ{� �y^VxBt��O�4��a�|Lc���I�P��П`�	ݟ@�I֟0i&ˈ�	�$UyYD����㐼m����O,L��E���	�'bkۊQ1��'�r�]d��ÃN�
V��!BP����'���' ����r�R��?љ'���n�u
����j�8�^�s�@Fu�r7O.%��U5���z��GO���	�S�Dx�O`�����>����,j��8�p�F���,k�P=O%r�'��'���'���'���ɼ��h�Hy���!�$������\��4���'jӒnZ某��4J�UD�i����T�'*��i�Ę�.Af,�q�ކkT(d��+ғ?Y�0{r�7g���	c�34R�pʃ&� �С8���#4�0�3�X8i�hl�McҸi\���O�.9X�2eĈĊvF\2!������3�0��w�h�xz6$B�]t2�s�-}�����D3aBRh�U'^���ݴKl����N�vXY�	^2
p� �T9vв��4d�l�`�v�̨n��M[�%�
X��U�fov������#��#�k	s�>���,�):��:R��<"=�0�ҟ���`���n�n�Jxq��ϑ	lLq��M԰b�v�^�F�����;�|�;0����?QQ!�	c��c"�ոS��HF���?1���.�x��!�^�p��S
ݖA�����O�DS����m�h�d�U�[���s��T���D���?1-Or�d�O����$,�� �5���أbUئ��1,�v7�1�C��,_�V	bbm����]Y$�m��M~ݎ%�I���hh���Yj� �K(�X���ûo��'�VʓpS��xb����FX�U%��<H��ȟ4��`�S�'�y�H22�0Q#-��=���91d����?�s�i$��Q��}0Zh�q�G8?�iX��z�f�R�`�����@`D�c��$F��J�G6�y��TR\q�Q�IzQf���yҤ�,[4%���C $QdM�a'�?�y��CtЅ��E�%Ja!y����yRBI�0,j��#=p������yBՏ:�8��gJ�/NR=ˠ���?Q�g�f�����h��所&Bδ�%��D2��{s	6D���i�dL�*�H�MS����2D����!b*QX� �+W����	;D�Ĉ��*S�ؘ�R��hG��з�:D�� �ȓ}� -kW�)���T�=D�����.�\�!�*@KVa`�<��i�U8���6
��/7 z�EߗR�6�{a�<D�x����Vq�1�⋐�2��Ѕ.<D��y�	H0COT�Z�!)���,9D�`�c_�n�\���ُC|�=���$D��3T�� {y��B�jB#]�v��F#"<O�t��LC���I՟h�s���C?B|���4�lx���ڟX�ɣPx0���ş(�ɁeP����Ԧ�.ϻ2W�Q?|q��%� ��H��7�0<�Qn�5OFա���%߸�4N��ȴA���2����N�Otʘ��*0����OF\n������ ��&V�ř$K�_�h�{t�:?������(����QBE��qR�!��ec(`����>Ɋ������U��>|�dʧ�F�>��)� ��M�K>	SJB^E�!��2�O�8Ͱd�@XH��:��f,���U"O�#�<@�f�����8N*"��f"O�LHӃL�["pʂ �
���"O�A�`�ў��}���A(���"O���$N"��x�㈪[�`�2�"ODɸ��/�F�k2d�7 F)�bKu�ГO��C%����d�OF��<q�	σ~���-��!�a�]�J���$�i7�6- Ei��K���|ʂ���P~�� ���/�p#��,��J�]� �`�7���"�	��$X��'zNA+ O����4r�) E�qʵ�iv��N+ l�Ie��\�	ퟘ ���.���sE���`Ѻu�fNgx��P����-:QJ�≁�l.r4�#�O���W��@�4���|��'��������1	I��ir1�Qzĉ0���O����O��d�<�|''E�d��Ȇ%]�xb��y��J�2�衰��G[>���4�B�`��y�J�o���WBA�=����λ���یKCT��`F*(��t�7�G9]txEy2�W�[](�To08s
Z���E�$U����?	��D(����ڜ/4�Eѐ/�V���ȓH%5�&��(����GB�mx��$�ش�?!)O��@��@�S�)�jAZ!	F�HSCh�/4�����<���?��Z����D���0;⍀�=
� �I��@��Cm�9��ߦ_��I;��'Z��#�	�0�v�;�ɗX�FMj�\�{e��+!�ZD���Ƈ�0<)�"����Ik~��@��Qx�iQ
� !���Ӂ�䓟0>4��a~*�[��m��|J!g�[��@���&���^�����*��0�	oy��S	��6�)�I�|���Rl�@�S:B�T�S횴Q��h���?��ؽ
�r��s�L�裭]��?E��#�2C�f=�W�_�9��59�L�����x$Mj���Z����n0ڧ-��qB�0>�6��p�a���'{m ��?���)u��H�����F��	`tp�rW�7D�s�%ѱU�lI��A�B�D8!��4�;8�>}��G�p��xE�&!)�T"�b�צ���Dy"<��d�'��'0��
� %f�!o��hD�U"���!�@�g���o�R�`&��`�g̓@�>�� ؠ&J�p��7v,%M�!?{\��"�H0�J[�g�y��J�ÉY��8jP�5�V���4�?a�EhP�����,OZ���O�ē7]_,���D��/��h3�K�w�B�It������Z�Լ��>t��˓	�����ڴ�?�/O0��ۆ
�؅�uǈ"Z������QX�w��O��d�ON���ƺ3��?Y�Op��%'ȁT��T��bU3�V�$-��xR�Śf����I�.m6@@�R ����
�'����W!��y�6���0����?�q�'��}H�g����1�`�=C��
	�'',�Z���}��4�УZ�9���K>q'�ir�'���qn�~
�"���	��ޥi�@Q���֫]�~Q����?�#��?�����ԣR9fSj����9l���)E	DE葧�@�O�2�Kv��6{Ge�J�'���w�7S��7�S�ZB�L��@ؙNּ��	Q	a2zM�tG��SaџD�6��O4�l����*�lՓ�W�dX���s'��;��'M��'��H��瞑p�r�p���,;0��Ff�'Q&���`�K�<�@�^D������S|�p!l�؟���f�T�F5zo�\!C���qT���3���)+C2�'����S�ռB�.�O�n���Ɔy�I�JÆ;�`���鐽��d�=R�0F*:H7��SI�H�����d��3�O*�!� ���%>��r@�J5Qf�h��O~��e�'��6-�ʦ]��P�O��IB{Î��0@q��l@L>���0=�G_�Aڸ0�O�_��)S�ɀw�'r�"=�T��N��\�� ֹ-�I;��>��A�����d�%�����O�d�O��NuA t��k�f��� ��w��1��rf����'Z��1I\��Ϙ'�D���^W㐉JT���
tL��)EN�6A F�'��I�Y(��Ϙ'S6�`�-�Kb�[��_�!q��i������jc��'ў0��h�/YHDDV��d�J\�<���&t��A�^�D��ex�Oy�o9�S�P�����4V�����Rz捓�Bˎ	�5��ڟ���������O:��1Eʅ3"�B�◦�_X�pA-�!9-��"3�ȦXf���g9<O"<���L�r}k��IlN�!o-Z$.u���?@�D q  8<O y�e�КN�ހZ�5.������+�'�ўFx̂�r�;��4X���=�y҈W'~�	�h� ���3e��&��A�IB��,y4��'HfRA�ŏ5nW�U�2	_�3t*Ň�y�*���2ΐ�Z͞���I�ȓ}�d���*����� ��d�BنȓdjN���A^'^�L����*?����'��<���k[4��_Byƀ�ȓt�=*�KD�=ޭYZ��\{��	Y�~���	��!��J�^A��b�N�<Y��O;�~�զ�@+~�@�RL�<�Wi^�Dʂ�C��]���� '[`�<��FʦS0��E)�d�z���]�<q�L�z��,�u��44��b�c�<���&@��dʤ%^�BL� �័���5�S�O�T%	��(�& �CeY�Lt�+�"O����%|T��$dR�R<l\	�"O���-N�$��LYe��2K6�t"OF�Ӳ�[�(�e��A���R$"O>-�����LO4�I lK�,��c�"O��J*%A.�L��i����U_�D[�,�O�8���,!$(��\9a�:]�&"O� h����0A��{��L�d$�"O0,�TnuN�m#����$/#�"O��[1�C�F��t&���).y�A"OfV�yL��:¡�v���е*�]x�l+BŨ���+lX�):��26�s�+D�0��,i� ���M�>[��5�%D��S���$:�V�H�CĹj׸�K�#D�����&(e����Ő?p��A� 5D� BVgş���Y�)=2�����(D���kB�w�"�T�̱&n���'�%ړh� 8E�4D��X��@��,�!(j��RU��yr,/y�����`Տ6��p�Ui��y��^�p)�MFA��e;8��h_��y��Y�8_��{�j�c��Q@B �yR�ԃ\ܽI��0^7����iG��y�;wn@�i��HZ�r�����?��Kd�����i�4 P�ꎉ�q��ng�	�bo0D��ɤ$� �8x�̯d��`�0D�L0W�w�Ƭ�0�H�4��S,-D�(�'�98݈��t�Z�U	��3`)D�L{Cώ4Lp-q#D�2!��3<D��+ѣ� 1�<�q Z!U��8�E�<	s(�8�0�+^;bo����#mT�ܑ��4D�$ǆͫ�,����t�~��@�2D���$�P䩛��ʮaI���C>D�q�:H��R��9��4�'F7D��V�I+�p���D>w�<�#�?�O����O�Ԃ4�#��!������H�"O2}jU����)
#A��6`��F"Op� %΄�D$��s�<	�p "O���EV��؈RC0c�$1�"O<2�!�-:����gC��h�z5"Oਙ��V�"V.�
�Q1�H�퉇G���~���ʬGU��`��vw��8�i�{�<���&2�n���K:	����Fy�<�WjA�X�8� c�RjpL�pc�y�<9"��!�������z�D���`�u�<���I�O���h$m��Vg@Ջ1��I�<��d�nT	!E��(
��[V��Пl��*�S�Od��ZSo�������X�f�LYbD"O,����x<�MH��P�
3�"OhZ��HM�t��-���B0��"O��A�O�+QpQ��+O�C�1qf"O�0��*	hI�������A"O&�0�\���P�Ч!�rq�\��0D�<�O
(a���]�p8�-��ra�4�"O@����՛.�z�0�KSX
)�"O-sP�67�,���D�7:D]�"Ob� �.�:B2 �C -_�j �̫"OH��B"c岑�e����0�'�8!�'2D�1��,F��Rg�U a����'鸘"s�Z	�v��f�\4�]:
�'�B�����')
�� r�SC��	�'2h�2 E0�!A���(4�޴��'�FYZ�͎!� ��sٕ0�j��'�DY��E4��|RÙ�/`�������.�Q?�
ġ8� ��qΓ�@@�J��9D���@;b���s�&V"+����7D�<
��܋'\�`za�KC�|��J7D�@)5���DTT�*N�F��g&4D���(L8_,ѫb�N�_6"�hI5D��ʦ���M9��u�N�+�@��O�� c�)�jBQa��$� pS⟆y05B�'E�l'!K֖�Q���
c��D���� ��p`�F�%�N��%�����B0"O���FH��vUD,�`�£R�Z���"O����)t{���U�R�{���3�"OP�Cl�$[�X�X�͌}�C[���*�O���[ �����G$}�y�"OnMJ��Hx���A��V3Iwr�#"On���#)@0�aX�pmd��"O<-Ӵ?�<��ٸ+V.�Pv"O*����%
�ҝ�"Z��}��'�2���'c�=Idg�x��ٙ��$}��j	�'�.|r*� ���@��@�~9��3
�'vd(�FO6�����(!�����']=2V`�&_wx jd�6��z�'_^D�2�1ܖL�f!�eD�
�'L�!"�%6�\��g�QNY����l�Q?ىC��T�ۂ���6�l��� D�,�/�*|Q�k�Kl���� D����.�<��`.� I��()D��"��X?|'z]�(�,��xWi'D����ß�'��,���6~�ƭH#� D�T�!�C6M٘ ����Ё��6m��I��"~� ��k.� Q"M�=��ah��>�y�iM�V���X�KK&P��=�yBi�)�J]�ƃ�DNp z����y�(��/Dų�G�$Ce~}�R��!D���d.E�(�t����&,��DH;D�D{I�=J��h��g�=9�PeCĩ�<�U��`8�з*͜b��z��+O�^,;v=D���0L5W2~�a�A�<�Ȁp�/D�$ ��N�Ri�t�޺����4.D���G��}�$������"%���"�-D�� ӣز�ؖΈ�u��07�*�OZ����O
�2�hݤ6�0q0�֯CFܨs"O��v![�;
`���-�v%��;�"O�ujp�G8��U�2�7X�m"O�y�"������/]�T�"���"O�5@��nגx���_����"O�L�(�)F��YB'k̯A�N0X5�	7A�Σ~J5G̎I~��AB*Z����@UA�<�r�2f��(��B�l(�A���@�<y�Y (��!�,0s��]�#|�<�A�'QI�t�`l��!1Z�g�_�<1�Qb��L�7m�%=��P�p_�<ـ�����0m �N�P�A�������0�S�O�Y�@Hn~R1{F�>VOB�	"Od��.}gX�م$dK(T�	�'<pqU�%3&\ŸԈF���
�'U܋4'�P�����g������'�:]`�O�;-̮��D�I۬)�'*4�Q�j��L���@�Ď
)�t,O�e�'�ЭaFlƟR����'���<�A�'�$Q�AC�f ��v��3[N8���'$���	J.tRD��F��&�`��'�/v��E°�V�L^,�@�[6�ybϕN"İ�)��9�|��p����>a�aFh?�*�XIV��RMQMC��!�Kk�<y2b��[7�����s��t9���h�<a���&:μCc��:��41�AJ�<�#��$��x&�3MH��Ip�<a����1a���O�.zO��@VFAm�<��`�:y&x��a�)J�⬸��i�'X�̣��i^=m�*�8�?������4�!�DϗCZ1�w�^85Kcc]f�!򄄸teN���ߵ&0��VIT$/!�� ����ʝY\d�
GC�#PMA�*O�y7"ژ5��(b��!^�&8#�'E��B6���W�<���!24R��,�aFx��	�Iw4���U��޸)1��\>�B�	�+�b �a5t���A&0=C��<(���A�*U03Mظ{թ�d� C��1@��(į����`$��B�	o¥��b��R��� roG+߄C��!c��K�j�;C���(�j�F�
��	W�$աcd�~3�d��8DC�I?!U`�Uƍ
2��XB&O;#?PB�ɺ[��HSm�M��]��6~�B�I%9l��yr�*��\��b��e�>C�I�W�͐2�+MGE1k�:Ya����C�&����-eK�,�%i�� ��V�Qr!�d;g������6N����@�f!�$6,֜�`���a����@���!����3@%H� ���g�Q��!�$E>ܼ��@�0
��ȣ��<0!�$�"��QjuI�>A ��p-Z"ўtsSo7�'yrм�AM��@:�;E��v�ẍ́ȓz�м����\�h�+�y����T����w�"u�0�R.O !�"��ȓjZ,���+0 #4�D3~�=��+� ���Z9��x��Oi��ą�k\Lpc����i�2Ixta����ɈIT"<E��m�Ԥ#�!=4������6jB!��> 
B��k��z�Yr��>�!�ĔO
� ��g!Θ���D��j}!�D�6P�օx���G�fɐb�8+�!��31d{�+�����j��
���v�h�)�C ��t�D&υi����)}"f�^}�	`}H���	ɒ���q�8;}���L$��B�	Ou���G�v�� hdʆd�C䉾o]@���b-* ��@ư+��C�ɰ �8�����;t�$�1�lC�^��C�	�Yy���"�&�p�W
qP�C�ɺ:<�{ֈǹ=,�)F�n
0⟴8 �>�S�I
	�r CT�]�y2��p�l�*�!�^�i�h�Y����1Q�X��[� �!��I<Z�ƌC���L�r�bN��y�!�D�>���'�L�,���	�!�I�a2�a���/XڤajA�B�!Z!�$1������i�V���Ԉt�L�x��*�g?�ǚ;�m)��O0q	P<�c�i�<��u�<ٳ���)XAP���LWd�<)Į:��BŠʌ>Q�DxD��`�<�F�"_ʮ���F+�ȳ�Z�<yS/U1V.)p����%b0���m�<YVl[s4�kק�3cp�+����p�,�O����u���a���v8��r"O�a ��[��]K6#J�_Z��P�"OV��7A��D��b�*D6B���"O�]@"�\�B	���1P'"O�`Aׯb�`Y���S�e�
51��'��x�I�4I���dh���^Hq� ö�=D��"1ME�7iF<��\]����f>D��{��Y�I?2���ܵ��]�@�/D�<k�@�=T2
b�&2hA`��0D�2Ck�.��!��#V�(aX"k3D��t��B�(�&X�$� A��/�ɟ~�"<����*,�5E��|Y�ˑsulDaU"ODa��-�'E~E�iʋIR  5"O�В�j�
Y�֭cBA�K�@�7"O� �H��ȍ[�QC���2@^���"Ot��V |D� v �4��"O���P�ނ�lA:�I���`�E��O�}�Pi���7k�]�l5*Po����ȓH?vhCѦݶ"B����b�;\sv���T�����.FDtƃD:e��Ȅ��@����4��I��J��ȓs�6�� ��%+�VQ���
���ȓm�ȰcH�*uFxH�W`˴>T�I�Dy���D�=]0���I�ysF�#k	�C�,b�h9XV��g`\�g؉,�C䉀&�	ȗ�F 7�5J�׏(�nC�	�E�D��,�6!؎��E�w�JC�ɧF�P�F��w�mztGS�e�F�?	�KO�[y�f�'�B;�n����F�}񊑂����S`�'�
iۧ�'r��'��0�U�'�1O�I?3 ��!�.I�pi��4iѝ�ԛ��(�$8���g�Ȑ�ר4ú�E|��?7��J� ^px��6L�1g��g�!�$ȯ@N0l�Մ��D%�aۤ @}�}R�<!V�	Hz��w�B}����NCy��'Ҟ|�Oҟ��� �}:61C%��6��w�?��y�>�b���,J �P J\2K�H��+��I2>O��������K��� �ᅿN�)	2k�����~�K�����|ΓPon�)�˅�BA؀���S-{U�5�W����C��S.��<�OLdă��3Nݲ�HȀ�i]�\�D�C���U?���9O�5+���5Fbjm��nZIl���2t����u�Ot��O�P�*5�H�)�8Hҥȼ�Fq���PT��O(��&�S)-C$��7L���e�L�J���I�MA~�'���'�"AL�Lyݴ6�}J�)�&Q����sAQ�x��@�'�P=�M�\p��	�=�Vpy�����DJ���%U&	�AOʘ�O�s��S	!?I&(ʄ[jL��E�ߡ`>^���hې��L�-O��p��O��$֙�H�4�x�ʟ'�˅$�B��#�
^?qr��g~ʟ�d� F���3^���.T6��l�~e�*�k؟���էj����$�+4�$�9��%D�(��$�]�2��@<`��]N~Ӛ���O�ʓ�?1����|���@�`���I�(���2bԽo����'X��~����i�OJ��"�( �@���@ZqFT��lM{������?�'��	�v���+FmG+��E����h��C�*Ja��X`/F�$��-�ĈR�p�C�I?X����#M[���p� -��B�I=g�N�
6-�~�p���lҜe
C��ʤ�r�.��|�h��A���C�	$��,�s��>OH���m	�F`�C�ɩO��� �a��3,l����oqxC��/���ǁ
:w�p �A��1c�C�	�2��+��'I���׺7��C�ɣ����J�$�����@��w-�#<�&�)� �;���ٷ#2-GX�:��	D�<$�r�a�e	/?#�er�G�B�F�����P1KqL<��Gԕ-��� �5b&h�&��ڄE��CC�R�ɰg"W�0�h@���Z�P$4��	qJ��i`	�"�T��EN�f��)q�%X�����b���������i�����ʐ���`�	4�pp{�
��THa���2�H��+��G�| �l��xJ۴~<5�@-S1O���E ܸ{����'�R!ǐk`
���� �T>e�O�PE�' @�戚�g3B�M<��#ΤDɂ�"Y�"|�7O�f`�⬋�ޖ�I�F}|=k�튀��	Dk[�)��'4�9��(R�F�qӘ�D!�Ӹ=����a�/CXP��	W�B����CX�h�G�ޑDkV S�*W2�`�pT
3O�PFyr�	������iK
��8����@Ǯp���OZ���+�.A��B��O� 9�&� Y!�յV�~X
'e8��Ô���S!�=�9k�l3�ʷ��!�d�<[t���LB;���2a]$:�!�dN%�ZE���մZ�BȒ���!�8P�(Z��Џ ��tۣ��x�!�$�3%2�DH�
 '�X�jD�ȱH{!�� ��80�tL�!Q�\�V��u��"O��M�IΩ�_� nV�k"O�r�
����A�Y�U�(��"Of�jk�?d��A��R�T��"Or�zWŕ�Y��X�#_Tr�{!"O�����dVB�B�ߓ*&��4"Oti�%/��$Wb�(��L�6���"O���4ER�)����<STdɦ"O�-z�"�6m��X��FZ�dC"O�Tȅ�͇~�4�k"hK��( �"O�� aLB�u4S!n�*�<��"OR�C!�/{{�SO>�U��"O��a��U�������ҁ�"O���4̕�I.��S�Bԋ_����"O�����!�6�C��$%Y�@�1"O>�C��D����0�;"倈�"O��!p�̻X� �cV�1S�� ��"O&��C�\�4��լ�7U���0�"O�l{�jݚgE�J���6T4"O>�`"e��v֖R�l̺ٖ0��"ONmrǈ	)a��d��[�0y��"O(����31�i:�k>tC� �#"O*��6b�6x�l���jV�t�`u"O��r�I��p-8�󲉘P��Yc"O�e�0�,fP�R��i� i��"Oޝ�/l���d�t�p�@�"O|0�B��q�NL�qB�@���"OpL�v���\�\�*���"/zMaC"OxQڐ�%i��00�!�3>�*l��"O"K&bX�~�uc�Ќ/��c�"OX��0�0[�����J`�r �f"O�8h��߱(�`�d	��83]��"O��ڲ7�Fr �G2�H#f"O��zЕbY���Nۋ�w'*D�+3��p��Q ��H�wH�1�)D��3@�C�I_�h�l�J.����'D��pC��qfT1+G���87��sbm&D�D�䍄mv�#ѯD�rL��pf�"D��z��*N�y�pj��6�x[��!D����AP-F�V$ha�?m��0h >D�dY[�p�jV��&c�j\!��.D���Љ�4#�,�K1��W0|��-D�(�A�J�`	�p��%L��*D� d��)
�t�I�UBH@H�"�4D� �T��l���S��0C�$�N&D���pL��o����#������0D���s��j��c�/ѓ�e3�L*D��v@�9[�p���!�[f�)��&D�,'D�9�,5q�.O�23|��&D��JB��8y�P�p���\�N	��9D���#��	$z Ђ�G�
����Ro6D�����_�Ři��#��CT�4�l!D��Kэ\�a.���E�w���h�)D��4�8Uq�L9��Êm!�M��#<D����CT������B���%&D�8�A��Z�xR��*f,81�g.D�D����#Vb("Շ�
t,��bC/D����	�QMQ�ወ,� �c��?D������X�Zĳ� �:(Ԭ��(D��)$���\���aK��q���j'D�0��A��n}F�@��0���&D�|�C�d: �(���4-�&�Y��"D�|ڡ&^�x�&�؂���0��05	 D�������Ra� 4�]z��?D�� ��R`�nl=�#�7V�N���"O����]�s����d@�Eþ4�`"O�y)$�^��1��N�� U8�"O^	I�`�55,�c���4{���f"O4P�Ō�f�~�3�$�.
u�S�"OXe�bJ���Z����@�;�����"O�	��.+Y����G��eQ�"O� �M�M�P���
�6�j]��"O���7�E�I�5	�%3�N��0"O<�)���	8������K)�xɁ"Ob��⏒0<��B�����E"O<UH�섉lVDm��e�9h�"ࢧ"O�XZ��.8ؽ ���&@:��"Oj�3��K��c�I�TQ;"O�ij�G�9r'�{ C�1Cm&-�t"O�]C�*%S:<1ɰ�V�$S�ɂ�"O��@f��nF��bA�eJD� "OV��ρ?}ڎ��D�߽!A��f"O�Չr"��!ӦH�D.�A��"O�E"�ɘ|y@H�`M7�(���"O.��3G�?C�J��g�ߔ(�L=c�"O,m{�Q;<lty�#K��u"Ox(k֊2u�� ���V��[4"O��"�]*?�n�X�k}�TB�"O:xBd!��8U���TQ���"%"O@�6�ԹH��Kj��U!4W"OL�k"O�g� 퉵*߻`s|��t"O��X��	BD	S�@�5)��eQ5"O�݊'�q&e�qϝ�sT%A�'0��W@��V:P�`֊�%��k�'�p��c!�;` �����
.`P�'a8<*3g�4������?f��ec�'�|�˖�R�U#v�y�%]�b�̐
�'�"P�G߇4.0����=`�n-�
�'f�hB3��v��EScΜ D�!��'��9��Sy�@���#kz��'�(�A��2�@H`��- @���'�(z�"�<B �%�B-ܝ-���p�'����0�\2Y8n%ౄ۸YxD��
�'"F���0Q8ݓ�� ���'��d��d��J�� Æ��ְ��'h&@i�
�/�@i�@�^�����'>)��ױBF�A�ާ%�ظq�'��P4d�ZZ�M RN?#��ty�'	�;ǡ�&}@��f�1 ^~�c�'�;��9N� cf�+�l\��'��uy���Kh<����|$���'H�9��C	J5.��ݬn���:�"Op�;$��[���)C�R����"O@�QNO)1��iA%Ɉ����C�"O8� GYn>D�5��zO��"O��x�� jؐy����2B2�bC"O��d��:;u8�3 �n-�pf"Od�+b�W%X����Bc1W���"O��#	�;������Y��A��"O��0����DYBH �̝3w�X�"O ��G��\42Px�ˮdZ�\Hr"O�S��42BT9��$�e;�@��"O��ꔌ+��U�b0� ��1"ON@xF
��X�p�;G��ja"O����'U�7Lb�&T�<����"O@�8��
�[ ��`k�,V��!�"Ob�5ɟ�{"9 �#�
0���E"OĈ����$f�P�ɀA�� a��"O� ���G�"
~v��!H��"��d"O���F9���G-;��(A"O.<���=>�8M(!ëk$�	�1"O0�W�D�T�"�	�.m����"O|�G쌽,%蠫��]�(s���"O�L���Q{!���@C�e@��"O����W��Qp)��@Q́R"OD��T$��r��E��(]Xq�"O@u
�h�6s�]{�B�2G8�"O��I���+v��}���jU���"O���b��KH�9ڐN�S%�x�T"O���
�S 4���,�&�1r�"O�X�A�ޖsT��2D቞���R"O�p����F� � τ`�p��"O9�&�V܈��	]�g8�2�"OdJ�Үw��8�Ɗ'��"O��#D�~O�}*dݷ\�8�B"Ox����+��52u�ě��]#"OvLfƅi��a@� a�BP"O�$0��<5T�|ðE��3���Q"O�B�(�%;��;��]���2"O`1�`��q+�	�f,����"OF���晉�dhX��66�bH�v"O��٤�0�Z4��$ڿP�XQ�"O�M��*$���V��0M	0yRQ"O��e�!�zM����	���"O>�u(ȹU���၇̾fE�0"O\\�bƙ�t0AAG�c�r��"O ]�1	ѕ@���b�X�p3Rh��"O�}3`����a��REC�"O�bT�6u�\�����B���"Ot�"��VGM���`��$���u"O��`dBY@$�P���9�9��"O����K�~W
�QR,(ע�0"O$�k�MF�I�P��%�ӿb��)�"O,��/@�!YA�f�y��AQB"O��k���^Ͱ(j��![�H�C"O4�1$��Y<-1��3L�܍#�"O>���ƙ�^�أ��Dp���R"O.�H+I�D�m�$\�J�1"O.�i���#K�z���Xm����"O�a(Q̍6���.ZW��C"Ol !���=�BS�T�N:�s�"O^@���?jf�X�%ݪ(�u�7"O�UB!��E��R�e(D��"O�	�@�v@}�#eQ�T�Ă�"O�%����z�ة�7�]9c&$%�P"Ot�VZ1~y�Si݋��zQ"O,�`�I�>�=Hg'�GHE9 "O�4�C�L-D��bئ.���@"OJa�%N��E��� �E�U��d��"O,�Ʉ� �V�,�A�J�3� u�"O 09��CE_�]����!O��c�"Olx˅?	#��o,!�"O��
�
g#�X��bi����"OH��f�5����W�[OY��e"Oި[���3�4��֏UV9�	��"O\��6�M�G�jƎ]�8��a�"O��P���c(:E�l %O ��!�"O��&L���y�e����$��R"OలC�?n���c�*G5? *��"O(���aS	#�6�30H���ebv"O����$���.����0#�\���U����m1�2p�=<OUs� (V�"(���\#�Ѩ�"O� �5�#�<W^��E�Y�0�Z�Z�"Oڅ	f�;.��Ic�����(��"O��FNX�#�6{#,���M�B"O��#P&ߝT�p���c�*}��"O>��i=w�I��L�EHB�!�"O�P�3ǏP��ȟzSDش"OB�U�L�e\~�Y�oȡK<R"Op��J!%Ţ- �՚܎��"O�����nIRE-J����F"OTD I�#	] ���M�2%ĄH�"O���dͶSȆ�;F�H�K�l���"O�p+W�)+�yz��9O��x��"O�8�Z���b�@�iy
�'C���2�2Y¬mJR, �?��2�'��pԫ�;��a���Ǎ �ʝ�'�fd�􄂓s
�%���Y�\��̠
�'9L�C	\Q���I�6Na$-��'��UB���1,a"q�P�.��'5P1C��1InJ�0@�9y�j���'��)�OG*[���%�b�'��s�Q7\�jF�ЖL�:d��'�$��J'�M��~\�y�Ks|����B�a+��gș7�y�C�3P����:0~n,p%:�y�,B1z}Ҕ���J/"��kӠ4�y�0�ێ8�,�Ҥ&VX�\���'KZ�GK\9!��(��i]��,��'F,Y��U�&j�l�w���Y��%p�'VXHy���B�+�$S����'g�0��¶ʮ0BNA��N}��'s�t0�(�ر�tD���Q��'l�Q�p�W;{���g�5{H~`H�'�D�i4	^������w�օ��'�6���5Y��`�f#V#;�0}C�'�Jk��Sg�MY&�;_�`�
�'�d��䌌16&	�`
�8����'i�@Qc�u�QB�'��*�"�i�'�,� Q!j�d��Ktp�H��'"d���S�h��A,ܧh��E��'f �d�XY�H�۰.�("����'�nV �2Wu$Ըe%T�,4z�'��]sV�+��}P�K;:� �',��W�BBF��4gK�U���'�.%�-�#�uH�	���K�'��	ն� �z��	6Nej���'�f���%�
�P���G�^��'I^X&1F�����gпH�r�'��x�p�ʥR��l����-,�0��')(���f�eI���p��".��'�F�Z�WE�2I"�(��n:XŸ�'tY;@��@T������n�8%R�'��x�D�1�.IK,x�"�.�d�<Y�h�3rr�1�d��|�"��H�<�7+��-p��YGcކ+e�zb�M]�<I��jK��u��<4{���0F�\�<i�C�!ZM:Ģ�ޝ7%Fx�!��`�<� ���}��}SX(��ox�<���:ʼ��Q"�l���-�N�<pA�4�\�ze�G�F\"�iLq�<��"^(A��;f�������S�<�%�%� �WO 2��miU��m�<Yu�e�`����A�N)��Ol�<�W�`k�aiĄ�W��©�e�<As��!��U薦�O��B��<� f� c$\0y���Gw�"��"O�b$�Z�&&p�3�?6��\!�"O����׏"�� �U*��4��r�"O�����/wqfQ`�&�4R����"OX��,WT[n��� �"�䭘�"O�!�1��6&�*%*����r���+$"O�V��!iI�I*B�Ӊh �4"Of��a�zX �ۣr�V5�"Ol�#��6�e��M <�$�r�"O�܃�f��}�88,���ah�"O���� �[���[B�N;dE���"O.�R�ơ/(԰�`O�~�z9�"O��b	��&���C������"O^Eh�+S�MX����4�z}��"OE�6�T;_B�6˲��p�"O�hA�mB4GY����c�)���w"Oll8�7{>�SţE�r���"Ol�rǍ�{蒽�$��uш�y�"Oj]���%�N���/M�R�̒�"O��
���Rj��T9_&�bw"O��P.W�Ѡ�ҞFޅjW"O�@���
f�2�˒�B���h3�"O����)��Nb(Y��O��:��'"O�Ռ�>|[����C�5�ݚf"O��Y%��15�����j��%B-k�"O�B�����<:ǪY'g2��r"Opt��ɏ�$t�7��A!���"O������N�9�㰴�"O�����O�~1�b��;�0�u"O�9��أ0,�%�ł�U�Ċ�"O.�"�,ޠ~*
�J��Y;|Q�x(�"O�UkD��>e�+D"�9A��&`G!�#9��%��J`�dD0���!�d�7{� I�+T�`7��I�T� �!�D�_ִ�Y����<̮�I��	}�!�D�@�]�7YO,���u"�!�&R8f�{�@̧- ��;��^��!�[�.��� �4\%��)2z!�dI�f�Jh �,�
8|౒�ٶW��4�R���|� ���|x�R��m��o�[�<�q�_���i햝_2�!H�<����vQn��I>E��oN�;��Sv���0�����y��
`�@��2~�> �A����R td���	 .B6���X�j�,ۅf��ӧ�Y�a}�_2Jɕ)��3��� rB�j EP	:�
O*��!�Y�+�1� )K�,�~�S3��/<��T�K�4�$`�IBv�Si��kP! �/4��Iqcܴ&�C�ɳ�v� &��$ �������F<i�`."��L �B���Z�)��<Q���<  �Q�d�3f�B�J�A�<��.�j�@S��9t�����ɠ�:�@%��.tUZ�A�Z)>9��3�@~�z�c(�V�"�%�$j�|��I
ْLP�n�7 ��\u���SjR�t�*�s�i*���Q|%a��1�lA�CeJJ9�e���'Bh�§�Y.��ѱ��i�(�:$�~"rlP�(�N!>��"t�m�<���9%���礕�j<ܰ���
p�j��U�˟?�ZH���[q��F�T�Ozİ�`�n bB�ٻgЄP@b"O�$��eъl3@)֎Q))"����[�i���2��!m��&�{X�n*�Et�ٚFG�3G�|e���EY��i�퉏l���%Em
�U�ѯ�.bE�5�L#<jn�q�I$%}� �V(Fd��P��.ű2Xx���бz�LX�7�IS���AM��TG�a��K 7G�D��Fd�NZ�b�A����
��v"O$������W���l��f��!��I�K��zA���H�8j��K�>���=ݤ�2�T/W��0����P�>B�I�K������L��}{�'Y�`{t%�pͮ>Y��˛}I�٧�ϨO� �(�h��	h'˒6uZ�Y��'kt�U�A�mX|Yjp��i��
D���u4��ق͇E���Q��Az�*i��)ȑ+4x-:1�8�uE�3���y�'?y �%I E|J5b�<�H��)D��A�@���i�S�]�T�e�Tè���PF��jmB�I<E���O�d��2�M��oK��S��;�y"�Ō!�l,1��[�%ZH�C3�����ɗ˴���nN�p<����g:� ��	(=�d�o]��Љ����|�1���Cr�1� N1�2DG(\ah<�G�Ѩ��uB��D�`��}��r�'F��C��n�t�5D��
0ܳsj!f�C�I3j�䕒��է9(���$��C�Ʌ$�\�ґ�Λ/������_`(B�	�?*�`�%�?�. �F =
B�	
Hj\����/��Z�2ep�B�5$By*�����N|�a
�Z�C��?B`��ͼf{F �5V�dB�I�[Pj���g�B\��� ՜$P�C�I:S�B��́�`@~�!�.�%��C�	�F�X��A_2V��q�*�B�	�2�m���ď|�x�"�=7�B�bz.�۶�9b�!�5!E�CT�B�	)4Ƥu�֦Z?ji8���-nC�	*~Q�9#p�@�/0@Y�iJ�.C�ɼT�������ੀ�b��$C�I��^�b�eB���L��#S�B�$s������&�R�Aˈ�'ˌB�IS��c�zs� V!ˢ4�PC�	2J��k����9nU����O2C�	
fx��"f���2u�r�]-$C�I�_IY��T�9��H��պI��C�I3waX���@A#w�(��P)R�tV�C��@�Ɛ�`+��&�h�t�E.bB�	hJ���BK�"r<�|��j���rB�	�r�Zx�Wc�#�,�R�O�QDB�	MU�zĦ��~2ZyC"�OAvB䉚O��	�%��(]
��4�@�C�	,�P��,'{����o�w��C�	}/>��v�Z�-��\�E�!}+B�IE$�A�)���C�l[�n��B��w��9G�R�]?z}{W�bw&B䉀v:��F�M7vD�'/;;�B�ɏ#��|	�*�=�����B{vC�		e��I��U�J"���� )L� C�I�f���� a�8g8�y��@��T�B䉠q�`kI�C%���D�$�B���TÆ���=�xTT�F!;�B��;|t��Q���=�p��;"��C䉃:����d������?C��C䉿 ���0��O"�3��s%�S	�'�0�s3���O6.��fbE�znٸ	�'����E.9��;wl=l����'�rA����R���C�h�4d��M!�'h±�e��h�1���Oߨ��'���a���g�^���A0H�'�-)���(ۼ�RV�@3)J�Q��'Aj�%mTZ|���p���՘E��'/�U��N�1K�DI!^8�����'��h�0X	Sz�%�톕{����ȓo;���`h�0%Ҿ�9v���Z}�ȓ ��5�TA�jCx�RE���*��ȓ$"�c�:3����g83�2��ȓl�  WD�
(��K�m��1�ȓL2%CR�:K�:�Z�b��o�R��S�? �	j@� 3%�8�����xR�d�W"O$\R�"[���j����-�@"O��! S�O٪x�A$̈́xӐ%3$	�=B�������>RL�5	1<O`XuȐWP^ �G�@��8�qD"O��A�i���m�d� C"O\�p��)���g�R�3���2�"O�A)�<�5�խ���˥"O��J��R�]z������&���;�"O4��wDҩ9�J�в��%(fr	�"O��0)K�
�x��� �{��)xW"Oj@q��C����U�0�L��Q"O���G�
��7%��IP�"O�,�0�)����Ey�X�Zc"O����$�x��,����<{�=��"O���-�X�Ti_,�W"O����*s���U����"OH8����"�$�!.�e0ph�"OFd[��I��$�̃`H
89�"O�|3wI]�l��1�1,[EH���"O`������8��t�ҥL16IR@"On���H�9ON�"e�����"O�S(�}!� �Q�^F�>��v"Oh�5ɉ�E!rl�C���@��e"O��	�i�;��S̘�X�d�B�"O��f��-aP� &���3��5j�"O@�14䅖zp\��r�O�O�>%�S"O4�+3MJ�}K!(R(P���`�"Oй0ҤM �D���Ѓ`�J��"O�YY��I�N ��ˆL���L�9R"OȜ�q��{">�K⪌�����F"O�+5l��y�"�1!��0b"O��ҡB�4�QC�Ƀp���`F"Odk(W�9����F;c���)�"O�IY#C�!s���æ[�V�����"OT�EB�����'w���"O�,3�k��a�D|ɑg��_�$ب�"O:06�M����iAb���""O栉e"^�f��L�L=OFqZ"O"5��lE.�U� L\�a��	�'"O~Q������ 
 �6�P��@"OЈ*��E+%(v�{�o'~�R�R"Otxy�C�%X|H�Fo�M����"O~<Qg�I-i��������|(�"OzeSv���y�h{B�:Xh��p�"O�URB���b|��m�\�ĢA"O���.K"A��t����V���"OzͰ�d�x'�0�GV�GG�I��"O~�eA�Y �x1�+e��"O�%c�N�H��� ���.0�X9B"O,��1MΜ{�QI�@X��E"O��P�旆�X,RW�L�h.�� �"O��Pw�1!ܔ!
��4_�Ĳ�"O@)葢_3�(	(���}|���"O��bs���OC��{BP�h��}HE"O�ӷ�AM:� v��8Y��xXS"O^��Ù�#xzS#�3V����"Oԡjg%J�;�Ɣ�Cn��hNb��#"O�<1� ��[)z�[�#�[=����"O|�j��x�S󢊾9�J�+�"O�(����%�^�� 6>�}0s"O�	b*���n�藢G.��h��"Of�g�rBp�!c��s#"Ovl�u��H�|��r�V�PZ�"Ob�����G*��Rr��1���0`"O� ��	��*8�8:��A��̺�"Oܘar(H��,)��I $��)Bf"OT )`!Q.�50��QOi��a"O4�)'�7>Rֱ{A�܉zxp�"O��  �&@�"LU\���7"O���D)
������nA��Ѣ"O�����Չ9��m�M�)9,|(�u"O���oIk�\%sː�.m�A�"O(���	�|��l���
P��:"OF�"��5��pG�V��t��"On5��9O"�J�!�>@d�"O&��� �H0���14��A�"O���ʜ�`�pE"pM+(+n,�"O��a"mޙ#n<,����(!�"Oly��(��D�$Ҡ���.����S"O.t�pi����A���Ix�8��"O��;�F^ m� ��ӣ{��l�t"O]�q�]�?����A�t����"O[��YT��0���%��>�!�d	�S^ZTb�dA�e)�AcA��3D�!��
�^I[�Kر ��H�L�#Q!� !DY�Y0��?!�>��e�],d!�êJ�d�eOܛ~�8<zAf�N!�^#8�"53��1=i��h�=!򤐁BH�0B��a�\�-�	_:!��26|�%��3R�x �U�
�5"!���BcșҴ�ԵKnQ��)X�M!���|7F��A�t1d��h���!�$sƠ8���L�d��P�ح�!��]����������t&��C�!�^Q[$1P�ϕ�9�`a�E�%�!���
A�]�O�FԂ�1�ùn�!�� IJ8���kY�}�D;0 1n�!�d��Smt�@� \�����.,�!�D����Xɵ�."S�Ar"�,*�!�$ߨXTb=��AJGn�a@C�s�!�D�����T�
���z`n��!�$ʥ3���'�Z�|��8��ѿo�!�dH[�b	p��
Hpr�a��gx!�M�N<� h��o6�\�a
J�p`!�$�8_
<Ț�씺C6
B���ca!�ē�A}�{�Q!ФZ�M���!�D��*p�93�[�b6KҰL�!��)�����U�^�8�t{\!��:P_&�b�8M�ܰaOX�U<!�ޠq|����>O���e0"!�$��ip�P�M������{!��1q~�"��YN,��
v!�$Y�[g(���*f���h��N7U!�L0|>�X!�l-hf� "0�Ȉh�!��50��y *t�� �&HQ!x!��rr$|B#c���	��(Or!�Z��8��#oۨv���ㅁB	m!���+;NuQ��K�Yb��f���M�!��:)�`�s�Ú�\K��s`G%�!�䑃PM$u1��.!�e�o�	t!�DP7\d����f���AD�'qc!�$j?z�㰍�1ٖ�f�<eT!����$�W��1(����
F��]����̒�.��v+���#�?(����"OH�aï�"��r�
�h���"O@89dk.K��\ �8i��	�"O�QW"�O8:D���yI�p��"OؼSE�ME��]��&�V�:M��"O� �8C ����T(rl�%�ؽQ�"ODr 	�r��` LٟA�2qp�"Ob��U�G���2�k�t�n`�"O<YA��?Z�a#$ŋ�t
9�"O5"��X}2]x���[WF0��"O���	w��\!���4��x�"O�D�B��:�FūW+F:Z#\<��"O^d�se��!��$i��/�d"O�TI��Ԏ6o^=��'����W"O&���/IKQ�q#E&�V�>�)�"O��Ac��*!|�L2�"+nDH�S�"O>���Z�Y���d�M]���"O��a��_ :ʴ�%�8W�I(w"O L3��!3����M^��M��"OL�V��m���'D�P�Č��"Ol	*�0R�(�L�'xٌQC�"O��ɚ�;��5�� ��,��[e"ON�zWɆ��rS��7Ny#"O41+�Ј� ���a�0O���""O��� �U�*R̐�@�Ӕ���'�R0��F�tД�⇭
y�,<S�'�@����׺E�������h`k�'N��	�"3��$X�X&z �p	�'�r4I2❆!	�)�WI` QK�'C��2�n?j��M�v�������'Q��r�	��0�B�!L%�`a��'��ti���	~�J$� [�9[�': !i"�ю\ɣ�֒]Ǫ9�'�H�;�P	�&\!C-�`�<1�'d6 #3h�K��-��\?SL� ��'�̨S���|��i�. �Gf���	�'���	��G�I��`S��S�&�	�'^�I��l�9�DL�a�V�4`�'��)�F�a��i�D�;Hi� Z�'���H�"\>K��������'�H����=�ڐq���
A*y��'zd��$��;0����F��@ĲlQ�'�Z�	�g7~�p9AL�2:b$�
�'GҀ����N���� K�7�ҭ9
�'[����&	ʡ�F,B7���
�'6� u��(q�(�ɑK�)�F�	�'��$K�5A�E��f;,��"�'�.]�QÍ[�|��. x�'�<ӡ�E�Q*��aJ�
?r	��'o�h��B�<v"`�F)	S:B ��';DpI�iV�v���R����'��}����:/��	���21d�J
�'�䅉�FJ,�  A�+��AV6E�
�'�	����n)�,Y����Q�q�	�'�НЮ̙9�ʀCRjL��!�	�'�&a��Q�Iښ�B�?̮(��'Sj�J�Խu��4��oٙ4@!�'
�ݳ#ֈN[��z���3���'".%`$�$@�|8RgM�?~2vI��'���3D]�W$�F�ּH�'L6`��$4`�A��,ݡG��8�'f�8��A�V�0�?9�fy�'d�=��ǎ;�Ԍ�VhA).ƈ�0�'�u�!��\q��A6��&2�2\�
�'W��'�ֵl�``��-0���	�' FD�Si��x1
��Z"%��=��'�t��*|�@���9`�X��'�D��P
 ]G�X��,�z��'�=ae�Sqz�hao�<|�N4C���  �hRaچ_Hڴ�4a�S��-�$"O�P(�H��*�4h�Z�D�ك"O� Ɯ�tT�l P�~]J�Q�"O�L�ӌ�9�HP`���9\L��1"O��x��ۆ�z9�&,�f��-��"Od��3�*��U�#l�T���d"Of]��$$6�T����q�S�"O��y��ωT� ���F�@�"O^�`��7�%k��9M��mqb"Od]���3 ��
 �Q��r"O�!����'>���K��S<�����"O�p�ǅ_�8���R�ބ^sR(8C*O"��0`f��R%���H�T��'Z�
�I
�}/�h1ր�,s�]*�'�(QJag�FV�$�D�??�Ȋ�'��I��T�t���4k'���i�'v:���.�ҭCR��Q�T�K�'.�M��ѭ	�5Z�#1xs�T�'9���l��w������B&-�(��'H��#�iÆ�r!A�U�����'$X��B����Z�S�iHK.4-��'C�)�I�@wBU��I��~h��'�|qXW�0�=�V@�3�@�
�'�>��5�	_M.)Z�f�'xĮ H�'�̜K�N��pBf���ޒh�T��'�ڡ��J3�ڦd�,{&A��'��Tb�W[ѼTi� T�p����'�rMpT��!c��qbU���e�.�R�'g(�y�d
�h"h����J$� 3�'P�yG���t�08T�S�@d �k�'��`�K��X눜c���;�h��'�@};��Od(J�`�ߢǔ��'=�l��n�2����Ń�4���(�'qn4 �N�enXlKL�0N�œ
�':8���(5D����X.(�Ub
�'����1��(YZn����(hA�
�'�x$xwo�;X9�)����&�4 [�'/�t��M�/2+P�����/cT�Q�'N*��7 ٯ�`a!aٴu��EZ�'�~ਕ�ڵM�>M
A	�g�P�9�'G��ڃ$�-L����w!�eB�1�'��p�	B� A���H
H�A��'D�DVS�8\�S�
�98"L�	�'���b�^�/:D�O];7��	�'1N��L��Pb��Î>.�.�
�'h��V���1�f�)�љ�'���åM̈ft��E1!1����'�x#2��+UO�9a�HND|�X�'��I��"͒�R�i��?;w�4�
�'�0|23�m��SDf�7�$y
�'4�X�$�R>TDʱX�)��e�'�=J�(�$c:�YZ�"�%j�\r�'R8H#6HU0<�x�vً-i`���'7����)d�>�@�[��J���'�&�{wg�l���*� �>I��'���ґC��C ��ʥ ߷$�U��'O�Jt�W�#��e����E�T���'��M��$�$F�1�㔱<cJP�	�'�n�k�`Z>I3�ʕ-Y��
�'�|)Aw�ژ}�H%�e\�,�e��'	��������~�R�N<;ڸC�'�t�!H�R7�ɁC��7#��8�'��kc&ʇ�\zs %9��)�'��Q��%Z�� I`H�\.��	��� )�Un��o<��)7g����("OzM�E�Y�jF��!�|��J!"O�����H�&��Y0���?�~M9'"O����;+�@��QW����X�'��qA��JY�����O$v��	�'��!%ѥZ ��[G`	P�k	�'����(Ɩ���1M[�7���'l��kw�F�uv�ԭ�*��A��'��֋�	G{j�z�*۷9?�-�'���3Ѐ�� s�ޜ{vZؠ�'2��¢!G���狒n��}H�':�`�ЇQ���Sg'�/kcl]B
�'Ty
'�A+�r@צA�:���
�'�䠢 ��rɋ6��I}�	�	�'��I��L?B�Ԁ��ŗI��<	�'�xHV�Y0� ���ڐr�'��5���A*�;0�=0枼r�'�b�3шA2�^)�A�*��8B�'�
��toH�h4 �w�'H��'¬�v�ƴLx$৏M�$:ؐ�'Vft��fɳI&�+"�(P�N�+
�']<𠃂[����ËI����'�P�ӧ){��a��l��F�v���'�.Tɐ \}˚⭉-߆���'� �[b�CZ�q�$��'1h�@�'ۢ-)�i����{x�y�b;D�<�A��hل)U̬��|�s*&D���#Ȕ�GѮ�d�N��h��L%D��Q���*,&�c�Č Ai&��D�!D��q�E�`^L��<e[1Ç�!D�����CVXH��8a������ D��K�\����H
U�����>D���Qiګl�2Z��D X��E0D��a�1�d9�_��
�3� D��Qj�<O^�آm�8�6-� �=D����m�5,��E ��.0�.���
!D��a��L�&vzub%S+h�"��D!D��r!��;c��iۥ���Z��@8t"3D�,��,_�xa�xR�V�=<�,�&H/D�X����;~`ؕhn�Rj�H,D�$@���4���@gm_�!(����-D�(�],N�"ɦ��:�B�bcn-D�`����?��@�rKI&���� D���\$L�1���Y <��2�E9D�T��N� `i�$�r�RZ��i�8D�$�'
[?FH��"`���f����:D�ܹ�؀l���R��W�yx�qg6�㈟R���B
Z<0�ڢ�;#[*��"O\�xЈ�1g8>D�Pd�0!zՉ`"OT�"C���V���Q#R�;r4�G"O$`�R���H���G���5�"O.q� �p�f����?y8 Q�"O6�(B+C�6��]��g��kr~�h�"O` �@R�d&piŽ�ÚYQ"O�1J�䍎"F�rlK�\��8�"O��V�̏B�p���	��=ʡ"O��ª�<{�%Yu���⚨��"O~�
���,�𬈂Ղ1܊!��"Of4�B�zr<Y$�{��y� "O4t!�g\E8����7P����"O�dH��	�Y	�<Ц�ϼ7�$��7"O��I��
y"�|�f�Y�P���"O���R���>HR H�`�<=��8Cs"O���C˾�(�P�������"O� ���_�!��Z�.�Y��"O���uj�c0��� �)p�XS"O8HCp�
V��W@�1~â<	"O��觢����������"O�H��o�.��űvM�*� 	*"O��9D�?�Ѩ�쐐3�H���"O�{�� �� ٲ�N�J,�)5"OH42R�P���8uȟ�FH�3�"O<�)�0E�8�ZR�פ'||�	�'����D�ԑjNF9*2�X	-��TH�'\r��"*J���b*�p�Y�'��i�t�X.fg�HJ"!O<w�.�{�'��ReB�W�BT �=Q<��'4�L���ql�x���x�N� 
�'���N�
GqtM8���qzr2�'Ϯ���,Y���4��h6��J�'��8p��i�v���&\0\4,��'��p��(|�: ���'$��'<,�����K,��%�(M�:͙�'�ށ�Vb��s�(�!T?�p�9�'��y�[�A�t8��=U���'m��`l��9Ǌ$B��D��-s�'��q�k"�P�a��B5����'�����ȓ��ء0a��7���2�'d���:h���#Bh��'e�A��'b>]����> [x�� �U�!�x1��'7��A��E:MȮ��A�1F���'["�ʴD݊?�9Pfb""��j�'a��@R/��(�"W'�XXq�'���I�)	�8
��@
G���"�'JP�s�$��	�i�@� �*c
�'@$��f�]�}8��Y���4�hY�	�'夕����"Ѐj3%Q�L��'�`�r��>k��S�c�1k���'52�(��ǿ����i�����'�n�7�O$::XK�ҨI�~h�'��-[������	4*!�'������M�ܐI���#Y�	��'6^Y �A�98��ű�R�Bˏ�y�O`�̍�����^���.�F�<�$�I2<%L "�鈏x	��Q�.��<�����4,�K�
E�k<��+gÕy�<I���'�B9h�Xp��5_���ȓE�,�rP��}m��Q���9�h)��^Xm�rGNX}��e��5���$D��#$���Ǐ+o=@��C��a%!���`�5�×���Kdq!�$I�'p�Lq1E	�t��u��/GV!�d8_a�ѭ�6�2,c�� x0!�RЕ���#H�ظ�mX�V!�ć�$�J���-��-�^�	M]	f�!��)��5�h��1�:|ٴ@804!���/2���r`
�;𪉃'��6M!��4Y�慰�'��H�qr(ǥ\!������z���7�X� i�0'!�d̞�^��G��:w�^��HY�5!�DԔpx�����+N�@C��Y=w�!��W&m�lYR��C:Bw )��FS�y�!�dE*�tQ���.��9#g虴u!���;��Q�V�U� ̑���:/�!򄈻%H�r���z˪�	��<F!��W7#)�e�`�D:dR��Eis!� b�a�	�uI��Kg�˭ �!�d��!_F�kv��+�؉
t儮�!�� n��g&,v�k5�Q1"O$�3���:"5��z҃O�T l�J�"O�C�տ[%@��dE]2F�P"O@\�R>%�8e:wA0T(1�"O��C���W\����ȕHpc"O�c � 	�g�Y1�P3�"O�V�}`a��G>� �)!򄄛1��8����y�ʄٷ�׋d!�(]�s5��w���j��S&S!�ֹ7���+"�͡��I��[)!���i/�л��ˍX}��r�=/o��䋭�2���4���s�􈤷%me��!�f��i
  'KKH6i�U�����U��@�v$�WA1�S�?�NM���ђ�.\f�E��[�#�����>R���I�(zw���r� B)1"�o��GR>ט'nq��
Aj��p���e
Q'75W�KqӲnϟX�O���M�Ц�%\?��p2d�������
y?�����>�4ɐ�\RA	S�gWдw��r�'8�7���E%�dkG��Ԫɔa��Ȋ&��4nta�$@��	�0�h��4ݰ<��J�to�	�����_��q�(�:�v��t� ;������,���On6�Ex�c�5�d����]�7�����BfAP(��r���Pm(N��誟^]r�(�^����i��$��Ä�|�d��!�>V��dC��T�?�glF!�?���i������OP�drӾ��1"؃<�$�Qi�(KƬys"O�k�͍,�~ �A�Y z&pj�X0�M��iL�'��d�O��g��%+�9:�̨ ��Y���ՅVLfΑ���ȟ�
�ZzFLq��M2T�V�##�j� � �#�gy��֪[�Szٵ�	2-(��ʒ웮VDf�1��$p �\x%��Jт�������
4Ɓ�nc|Ƞ��&+(&�$������O
7�Je�h��%Zv����"��iK�D`�4�?�)O�$�OޒO�Ӯ,��Ѹ�D���`����CզB䉚��"�AF8]�c�ar�ɟ�M+U�i������4�?9����iH�_�|��?x�>}���b~��	dJ��������<B��@��� B� N�~��>PD@�C�B���!�*/�r�(�� U��<9���R�����"��0�U�g�.�b7.��<���D7~`���#�n���n�"��#�nm��П`��4�?9���9��E�"�b�AǍF/:x�lc�I��Mk��@*��<E�N�{�|-��a[�z��H�2�O�o��M�40���7i�Pd<�Qf��>q��h�ޠ���if�W���?�%�����ŀ<2�,�'���N�BS�������E�(Gg��1���0��!�J(�S�?���AU��=�B,�kбe̛��R�"�&� 2!\�Tܚ7m]�Qɸp�a Z�:V�#�˹|�1�.�h�DγN�6��˝+C��oZ%M���Ʀ�`�4�?�Οv����oԳ3?���v���ԙ&lĕ���O���dF�i��n�/a�R�paݟMjQ� bݴ8?���|��O<��hY��	b)q�hzC敡r6�h�	Пĩ����^=��ȟd�I؟X:[w���i�d�ItLF=5N�#�N��b]�	a�/L�q��p[�V���(*�!��f�iF�`�!3s�|"��B4�S���o��Myp�U�o�: ���1�i��� �p�a��j���f��\�H�@�����c,_-����� .%r�P���?�"�?�?1U��3[L�gyR�OD��9��\�`�֮fn�1�J8Bp��G{J~j���la��	�!-A�'��6'6\⦍�I��M3�>�e����䧏56�
�] |  �&M���9�fGObvt����9!�Ę�+�3a[:B_�Q�H
sE!���	omp�*F�VD�P.��!򤎈�6���D�T&
E�W-�.�!�����䚱��p��E\��ITy��|��	K=%!����*��>��hY��^9!�ʵSJ�����L�.�p�A�]�!�*\�>H��X3]P� �/�-~!�dRK��%b�<9��s�.�'q!���1J��1�%��l�rtzQ�Q�pl!�\2�Hz�*^�;�ѯ�!o�ў���ӫ1�Z$��ȋJ+��dN[1'ȓO���5fl�X�蝴0箑3�,=�!��G&�2�a���*M��x�$.[�t!�D�r�:�@A�VS�t)�'£�!�d��DM� $���'f�`�!�F��y	��OL��1E�:�!��,U ؒpkVEd'es!�i2ya%͌ke*\��(�*Vj!��)���lִN;���s�R�qY!�Xf%(���dAR?����@V&G�!��в_���[Q3t�脡6B�l-�ȓ6=�\�)-Y��#F��`9$��ȓ.�:|�v��. �[�/	�E�B$�ȓQ���gßee ��$�φ_0��ȓQ�E�mV5L�8�R	�n|Da�?A�Q�.�X��)�H���ʽt؄ȓl9�$f �5�:=�5��6y�Єȓ?���ϒ1�2P��/`e�E��z]��IR�;`S<�d-{�t@��EJ04���;z��������6�ل��z��5�ģDh�M�q#ĉ1֜Y��0����Iإ-�e���O�ą�'�YGN�&���ˠ�L��ȓi����j5+vDK��7e&��ȓw�D�bpnD�*{����e�Je�!��<.U摂���\���j�/g�!�߻e$ p��D>=��t���D�!��,x�qp��'C�\$Շ�?g9!�-:��,�!�<al�єgX%6!!�dO�G���-)r`�!9c���2&!���T�
���&ю,�H����_!�Y�L�s�C�02��1�U�[�!�T	�u�5%�'V�4lUӝ`!�� ��J�-��ad��Ғgԙv�8��4"O8 s�I�R�ZM��/"����d"O��A��G�r~|���ג;���k�"O�y�펳Bd���E�
)�4ٲ�"OҰ��j�%Ed���mPAp"qH�"O�2��D~taa�l�#g����"O2�Q�iWb�j��À�-dȭ��"O(H�e�C�v������ǽk[te��"O>Y�5j�J��� �Π1U^<	`"O^�x��+���S�ߚ��IS"O^X)6$^�t0z�H��,�"U�7"O<-0g�4�����:�`�5"O�QP�a�9 �1R��&�TM�g"O$)��KʞC�J��V��=s�(Aq"O�E��L�%��<8Ci��MU�b�"O`�Y$��	H،��%^�IE�U"OQX �7���˴�եr?�	8�"O*=��ɵ7�VĘ�͌�t�=Z�"O��"���8�`q` /��[|��"O���IW�.#V���Y�LvJ��S"O0��l�T�.�JSA�&V�����"O�P��n���ڕOF�g����"ObP�u*[��0�]
bBp�j�"Oh� 4D�<\�>9�Rd����0"O`�i�bJ�iS�}Pv%ߜK��M�!"O��;EQ�����pj_%!Ö()4"O��P�C�y�@!��h�-�E`�"O�	L�tXەf�?7� Q�"OV�/4XT����l<�8���#�!�	-R��	�&�'<el�3�P~�!�Y
����ʈSZ��Ik�5!!�D��@�B
U=p:�% U�_!�d��2�򌃀� ]Д��N�w!��ԫ)�N��e�#&�"\�ğ*!�D�-�<��'��A���a`���!�6�J�P$�qÂ �\!,!�d_Ql������7%O@��F�z�!�U�|5@�קǎj�@P�K�!��3*+�� ')�	��q`�@��*�!��=��b$�U�L�&�`vn(q�!��
��ʞ�rzR�[�a�!��+	��\�����JHF��l��n'!��m�L8��~م� �\�!��#���M��tK�`\=2!��$@^A�ڊ0�d��N�!�D�0Wp`���j۝6�H�q���#[$!�G8'v�`�@��A�b��g�Q7�!�ĝ!O1N�R&2wֱؗ��`!��{}�pX���߀Kn>�� =D��h���/3�ر�S�L�3V�E?D�蚗�S8/rF�aPJo߬1S�m8D���l9w�I"ċf�vk"�4D��iF��	�٣F�?$��%�u�.D�Ԙ����۞�*�ͷ��y��)D��JRȄ�f4ӥ�
� 
�:�5D��Y��^�+����Q��y�ޝbӮ1D�0
s�}4�L�&S;��usT0D����B#P)�QcT��$&�M('�/D�d��)҄B�ZLp叔-�n	rƋ.D�X6�]Ɣ,c���MzNq� 'D�,0 ��(�@���h�i,Ꙣ�"D�\��0B�&d�#�2���RS�3D�DzB"��!bƊ�U�h3�&2D�H���zabkȦ5t��N$D�� j��5�_�G 5��F�:ʄ��7"Op���MG�M(v=	D��
e�3�"Ol!�� \�A�`2���*I]�9�"O���ȃ7?ܰIS�ϦzCl`� "O �Q�bB�@�Q��+����"O<}������]h���~�C5"O�	qP�8�� ��n�M>U�4"O!seP0zƘEC���kH���"Ov���P�p��0ȥ��%"a;3"O�	C��+s42�{�$�{R�*"O�G�E�.�X⭇�)��R�"O� �M	vG>�8�D�g^z0)1"O2�q�A��c~PHa$� JT"�"O���'��DsF��E���db��ѷ"Ol�!�'�1b�ܕQ����Z�`���"OX�!�e�,��� q���P�a��"OP����H��L���[�D��T"O����+X��@��"(E���"OlXR��(�^D���VB%��"Ojp�(n�bh!a��-Old�x�"O6`�ET�ܠB�
�`�"l�F"O��0u��L��Ys�,�=b�%ڶ"O��DH)K'"��D�H�Qr�"O�h{"b��xe�m�&?հE��"O��W��3_{2�d�9VR���"Oz8꧌R�gp`�4-��=���k�"O=j�V�1u昺3bD6z�	�"OF����Q�\��(Da!uo�`Rt"OV�â��^����E�:QV���"Oް!.�40��=r���S�Y��"Oh}Kdȋ	z5��� �%R:�#A"O�숐�3Ua����J�V,�ػ"O��`��gL {4!'` "�"O�@x�!�!J^B\�7IĤ2v��S"O����ai�KA�Rx�1�2"OX����"s�|H`gGC�zl�� �"O�9z��΁Y
���.+��XR"O*�S����;�� �)�F�F"OH4p��ܪ!��<��b�*��E"Ovh��C\� πi�5��6��`��"O�P�`�|ݾ𺀅R"g��q�"O��1���
���K�$UG�hXX�"O�=v,�85�t ���D�����"O�,k���<Q��� u`���"O�9VbY�09�	��V�`dڵ�ȓJ4а�ݤ/fr����C�>&ԅ�t+8e��C�2�H����n�(�ȓx �P⥢',TRa�NX2Dt��ȓ:!�����{�x�7�0-_��� 7ƕ�#��[�0��E0Aᜠ���б�b��2�l��#�
T�ȓS �PH�#$�@Xr䘎J��e��~T�M��Fa�0���B�@��ȓ:�8��O�-"2a��ff���%]�����,:�Bd��� 6>����YQ<;�܍jZp�W�Ѿxw�)��\yr��/H"� )JDJƳh�̆ȓ$��a�娖#p+����Ͱ8���ȓ,�H�[��T*~���`֯`01�ȓpp	��D�n>�)a��J, }���ȓ9���X�'Xfb���[' ��:A��盀l4^���M�j��5�ȓ/�R��A��(�
�j��k0X��7�(1b�JԧwdT��S���\�2���S�? ����E%7V�����;,�U�"O��x�"�#{9mD+��r}4\ f"O�IR<CZ5���X>g`j�z�"Oح1�(A�Lqc%PX'�[q"OD�s�Z�%n��I��D5��͑�"OrĠV�^�y���I���Q� "O���-�&�,,)C��^�p""O���1��i����wH�+	�`"Oh�z���3�
+��A���]H�"OF%�Q&S�(��I��,D� d��"O����Ηr�m:A�F�+Ә���"O�y`/��v�Ȱ	@BX0��<�"O�-:1C�2���D�L��`�!"Ox��V�ٺ7��P�H���{�"OT�a�n�;E$p�JŨ3���"O
���>:���ȧ�6.?�(c�"O�Y�7'�/�t( ���1�1�"O4t�����!��������u�"O���ωR�~I8Vj
�fy>D��"O����M5'Z��bC	!X[����"O�T�!E�,�����+2E�)�"O��;��B����6�T�U0���"O&D��Eʞt��(tJ �"O�y���֬Ys�-����Y9�X�T"O�����.=y�hK�J9,l�'"O���&��	4{���K�  "�%s$"O�*�ܔ��``W�+���B�"OFp`D��y��()�� �_�!�D��yb��A�*eߐi92���"O��A3!���В�C3���v"O"Uq�n��=E���bKS�.�bt"Oh��a�L#^��j�d�vy�s"Ox�a�@�F}Y���&��L�4"O$P*��R���@��2���"OX�j0.]�p٢�k��)`6.2D��ϓ-p��di��{���"D�l��=>�<��!��8*@T� A+D�P�ŉ�!hZ$�b��M>j��",D�8�0�+2��0��b�E�x��w�+D�0X��	/�z-�� ǱY<��&�+D��9�ӎR�)����6���%D�X���S�7AR�2�G|��(�ǋ5D�(8�n��Tk��17O�j%����B)D��4
_�o9�]YGMg��u#cG!D���E딊/��z���L�Z��5n D���͆�>,&1���=~�v4�J!D���o(?N\��I��vO6�a�2D�ܑS"�@�D�"	�g�F���1D�������R��"K�n�$�!dI0D� �C"�\X�9j�	�y��T++D��cC��$S'��3�I96t�w�=D�@"��[Zi�G�',	��{�A;D�@ɤF�*G��M��L֘XR-PW�:D����hR�Y>r 8`h�k�j���&D���F�,n��bP��(bF��#k7D�X%F�5��8[Ѩ˗*��Փ�m5D�����.}81"�+*ru0�'9D��c�ݘb�6�#���!u8�a�8D��@G��#g��z�)�2]��-*D�`r��E�Z1�MK��
&_NC�	!U�T���b��%v��C1m\�� C�I�a1�Ԩ,G_0��� �چ-�VB�	�K-��Յg}hJ��P�B��@r��S"H�"����C�)� 6�Q�!L"1���)U�ú|��	��"O�`{�NE�ȵv��W���a "O:��¥�m��0�.�jE�g"O��ٕ�]�W�H��-�� �B�J�"O�� �-�}|ıC��O*T)�0��"O`x�I3K��X��"O ��t��C�0� ˑI�m.�y	�h��}�1IC�M�n��OI��y���v8RDt@K�j����
�yr���J�킅,�)A'�x����y�Ha{r8���2xD	J2ߩ�p<i��D]�Q]$E�r��&NԜ���/�!�Dּ%�ɀ)�7l�Y !O�}!�d�?�@���8{�
���N\!|q!��u��<�s%�._�V �퀧4p!�� �(�(�Z0@P�e���j�I����xr�ɴj����)�1L_t	 V.�x/�B�ɡmu� b�HV!r��Z����op���$ ʓH�T� Cī#��-��
^�-�ȓOVv`�!&	IZ��TY*sL��$�hG{����{YR��@�Z�����!I�y�,�	V(�0�u��}E�a��L��y��D* ��$ZЄ�%Q�*��O�yA�\|
�е��9q�8I�M��yRB?z8ň� Y�
9���y�ᆴ��橆3#��R	���yR�i4����|��*2��6�y�`C�p��I�jK�?���y�E�;�Hz��՞FPT���O�y��)�'v���#6�����E�k��Ѕ�}��8�HݱD�	ů�r5�ȅ�E���P�!=HxP����޵m�A�ȓ.s�P E��1$�TY��	�&��ȓ N�q�@���_�(���_�pmZd��%}���i��Ę���C��ic1(̮w��c	�'NnhA1e��r
Afͧ�h�'� 7��>��yR�dA���<���˦6~,�A@D��|b�x��X5���H�F�P1s��c�h�IGy��O�#?�wI�l�$ة'Ɣ�}�J4�b�v?��\�y0�d'!V�%����
����񉯍ē	�$"RdE�H���*U�:�ȓ[��	QC-���2uD[�*�B\Gy��|*%E�3��\�X* (�сB��t�<A��� .�h�� ��l���c���hO?��?g��l� ����t�E�G�c���4��I/WG�A���C�*A� �ڐM	�C�I�aH� �vm��0��Rh����<Yڴ+�	
I4fT-�B� ���0���|��r�S$Yl���6�%@����g�'���b��7n]̠{��M�>�b�	
�'��@��hX{Y<P 4�=+�B	�'آY"փڎK��s嚍2�<�	�'�bŸ3&^)[d̹��B(U�y���2U8��5L6)z%�N>��?��'�Ą�eA��=A&Ɲ=o��'�V��֛+���u�q ���$Ϊ�~��	YT�t�2�8H�R��"��@!򤌲0�J���M�r�'I��d�<L>�O���O��xuAJ��h��c[Z���1�h}�^��8C�'�$���J�PAp8j��%B\nؑL<���D=}�W�\ט�Xt�_.3]��HT*���y2�L�fcx���G�0Lei�g-�O&��d_�}��#&m�--X�h�f��a�!���|$� �-��%r.��l!!�� ���2Ί'��YY$&A��`�"O.1G�\�hB�d�ܜ̺0"OL@C4j�T�j��܉�$ �t"O	Y����J�ȀCV �- ��'��D�"���2l�#e�c��ؼ@q�{��I!C�*a�Z���t��eK�SK!�d�x�q����1���aqOѳV/��b?��B,�ŞSoЩ�A���&4-*���=�	�� �"0�G%S$[^2�k��0jt��{1��C�/�����p�Q���μZ��|���3BH�B0ެ��f��1�gN<N}��z�D�X(i��
DN(���A'[��AB �3n�xE�����L
��*Z���.}��ȅ�B�q���0�!E��9���	}yB�X�� d��9�-y�.�1�yB
ʄz�b:�d�<4�;sϗ+��'F��;��|�v뙍O��wL`��p�WtH<�eCͰltJYؖ�.F*=��W&��'�ўb?s��<eƂ��D�Ű\&�I�!�&��e�>q���e�/7g$���(>�I�T@���'d�zR!� ���O�y�襚�
ۛ�yB��?'���P��^;oi8 ;�E[�y�� &H{ �p�H��1X��:Ua
��?��'�l���mBL��b�I��a1��y"�Y�lx`����i�?��=Y�y�,��Y=,a�J�@DBP.��O�i���޿ �Ό�ef�a�X�ƀ��8j!�ߤD)�#�+��9�T�Ei��( xQ�"|�e�M>b���ƇD�$�ZL1��� �hO?�ɼ�
ѳ�B�72��`̾{;C�ɜ,T]��4.� K��5N��Ij����ԍ��d���2�MO$����(LO�㟈�l�7L�I�� h�^e��!D�\{R�N(%�~���ݲi�8m
R#D�0���
�M�X�c��q�\!aV<D���N[U&���G�f��`>D�A�&�;�\��tJ�j�n��"%=D�$ ��N�A�����Tj	{�L6D���Gn�e���q(Ϛ��q�c6D���E�٦�id�Km���4D��J�7�`QS��U/Np�<��'2D�X*G� H�ʔ(���h�:%crd-D�@���A� 5�-� d�'T2��1!*D���"�R�&���@M
�a�Xc�'D���#��-4��
��m9�ıQ�!D�3�+�3����%���"8�h*D�<+cg\F�F+���y�T�Fb(D�$z���T�ֽ�� �?N��3��#D�H���֫E�Ly��"E+S���1��6D�|��A8qޒ�b�%C�s����5D��g��F�� j���� P���3�O���p��P����R�o��Y)t�ȓo�2� �� :EZ��AX�~"���^�IAg	��ZTk�":M|T����-ipJ�T��)�A�)nn�لȓIYX�pO�<���*N�}���7b(
砙����{�n�u���b��)��pz���pЀU���,&8C$1D��iG�Kwb�+&��=���`�$D�4���n��0�qD�8���8D��� a��a����` ؤ��aN#D��ȳ����P��ƭ�#z�V��F D�(�w�I��>�Qb
�,0����Ǌ?D�� �Q���7���H!JTd@��"O�i��,�,���rD��=�p��U"O�4 w�ͳM���Xd^�z(�"O�BV��i��Xi!�^�`̀��w"O\���#ܹB1C ̐)�r�9V"O�`b�m[8���r�.B)��Ö"O����������Ǹ���"O�8���'j���ĦH��(��"O�ub#^�U���wlU=�<x"O�帖��J�}��HW;5�yr�"Oly"�#�6�T�;R- A�&���"O���@��xj.�`k�V�> ("O����(C�E�!�/�h�y�$"O~��w��jW<�f�@;}Œp��"On9;B`[�\�HY��Oթ
�H}�""O�<��0@�2	�G�Ȩ?���0$"O�\��P��Y���E[#"O�p�c�΢K��j�n��_ȌK�"O�H��չQD���#MR��v"OF�a�A�`Jx��\1z?���1"O��a�b�J�Å�d��Ё"Od�`E�S��0�D�]�Ѩ�"O� ��%Ԯ,v���M�"�`"O׋]�}��¡��_���"O�81��̜p����BU� 3L=
�"O��JwD�+�(;tK�	0P*$"O����,F$J|iI+��Z��s"OP[����<&��G�=��B"O�PA3�^1Yp�h�E.|�D�q�"O�L�����9x���<V���{"O<I�A_8a�
�yA$G�`�T�"O�P0ЋM^�PEB܅"��}� "O��0p��7
jFQK4�W���0�"O�yi�LF�!��y� B0f�Dk�"O^=�C��8Ȩ 2 �F[^h�G"O$ R��gS�-b��>X�p� "O� 9�� �ͱ�F�P]���"O"����)>�,�b Br��yR�	>< ��1��+-�P=@a�A��y�c��j覕Y#�ڮ,i¤�Sb��y��
i����d�Y/Y@J��R��yb`N�X��K��_�΅����y���n���k���4-k�a��yb M;8O`򥣂�[F�#�ր�yr�X�)۷�C�Y(B��rD8�yb��� h ѫV�J�i�Nҹ�y�H37*�;�*@�Jt�t)���&�y��VAD��T烃C���Ǆ�y��+;�B�	�a�",c�t8���y���{-0�A�	�	1�Nd�7` �y2i]�!l�릈
���S�냱�yr:���7�
g&D(1�D#�y����]�U�CD�6"����I��y��Z9��PV�F��Y"b���y���D����V��p�D����y��p�x���ۙC�$�����ybjL�U]��B�N0>���+�y�j��c��1�0p��(��Φ�y2ʂ!ZH��
R�`_�T�'h#�yrώU�&xA�
=^��P�&��/�yr�M<O�,����8P��2�)���yZ���؀$F�C�|��KG��f�ȓ��19�/b󲅹c�G�����ȓN�fz&��S2�I��<v��<��S�?  �0&Wa��H��E`��p"O.`0�IU�^R̔᧊��NƢ��G"O�@�6��m��\	�i0P�|Y�"OȩX�AI�xI3T�Ձ2;FU2�"O�*4Z 7\���`��"��D"O��صF��&:�|��a��mÕ"O�)����?c��-H�aBS����6"O@R��"�x�reU��vA �"OT�0�(q����E��.��I��"O�Q�E3"V�Q;AK�<�:v"O~��ӈ�#}t�yX��P�K�24�"O�X�c6l`����^4R"O"A�f�A< �:]/����h9!�W��	"D�� �ݚa�Z�4!�䁄D��'� ��=bшGF�!�)\T�z$�8)���1���F�!�d �`Xꖮ\�[sj)���r�!�Dٸ	W�(�b��;yz�2��1!��O��<�s�J!B��m��8!��Ƌ3ȸD:�I�m���VBЊ@�!��X�ĉ��I�d�b0���B7�!�C��,q �!F�g�<X�" �WW!��Kr00@#ީ��DK#�֞�!���'��)�g�t�Ȣ�	�H!�䛠j�8	"2�ܨ��ȧ-O�-E!�3�ҙAg�1)��"TL�K�!򤅈{  EV�c�r�ӆ�z�!�^�^ .����\:���W�W�!�dB"%7l�ˡ3lDj����M�k�!�$F�F�UŬ�(�v�cBD�T�!�d�1[ Fek0�*(��pA˻v�!���J8>�'��E�V��O�w�!�Z�t|~�I��D�?Y�Q�RĆ1%#!���Y$�q��('@
����?P<!��.��i����?�����.?!���%;r�1��&�]���0�CE	f !��2s��M�q%K�d��Z�(IE+!�ĕ60_z���H�d8�����Z!����M��E�0��Ѣ$Q�:!�'4���#�JO�j��5ʥ��!�M�a[<0X���5�d��'f!�$Nh��X�"L�p߆ a�e�4b
!�ċ:]6��prB��I�z�Dv.!�D�f>��Ġ�dBȉ��<L!��
B���C#M��b�Ӊ(9!��==g���%ǋ�))�����ԓ%�!�$`R�&mU�f|�T��ܡ�!��� ����)V,/�P��&�-v�!�$E���AP
����@0b&�!?�!���Y��،����U�?�!�Ϧn�l���`M�b�]��ń�Q�!��g��#�D��ʄ�,*�!��]==]Ԥ�U�Tz	�]Z�ݑE�!�Dո1>��d2`��QC�ѼJ�T�C��+BbIN4fɧO�DS&��ē7�|��5�͠e�ŉ��E>D4�鉲K������_#��y���QsLh���Zi���ǅ�<�ʐ	%W��3�^�@�Ld��]���X��O
D��Ђ�BՓ ���'�`ͱU�E+$�����>,��y�\���^��H��!i(��9�ts��f��B���~�����'eC��#�'@1Z���׮���Y���>@z �5̞��ɨa��%fG��3䇠���S�&@���#5�z"o>[����!���ѥ����4��
�@�>Q(��#��V���h��Od��� "Z�<`��Ov���"Γ`Qdxڗ�Vh��|����:I�m�A)^�\=��2�N�����F,0��<�4��Y�0��B�l����(Xh�5`/�����t�٢r��3>����5Ҏd�I���TZ6&�;N7
��C�=n��찀,�fʡ`L���� �x���"{pգ��īf�t!�fI6I�!�$�(I�a:��Q�y�����ۼk���2䛤g]�ǚ���{&*O�Ijv�Іy��� �O�A?bl� 5�8)�~��AL��?���=dV�DJ��Q4i"D�Ao̶z�����&*U�& ���d����~��Z5�ؐG���Mv�I5"L�Zr�J$Rц��e,�--��?!���3.�\e+�j�0Z�*�-��z���ab�"7l�+ע��Qk�t	�G��~��ݹP��b�D�?_��D|�`� ."�ito��P��̲k	���Q='@L�3SkҬ$",H��<A�S�O��v B�6�h�W(0Ј��S�#)�B�|�6��AC-�O���B�IHF�� ��Z|ֈ���)��KXyܘ���.���Ф��$������͹
��K�d`5*D�D���A���x�����2��сr��\Ux�{"��%s���
��\)3���e�!D`R����a��ى��9O��Ґ� "��P@(w�P�I�"O���Á >L&k���(���:�)̯;
�s��B�%6 ��N�E���ɮ����@Օd��+��\�&��D8#�r���mì� ՚A��<t���EvF�:�$��̱��=�O��
��C�<�7hX=d���;5�D�s��0م�^�
@��P1x�"�'���_='lp Ja&�$9RЅȓq�X)pፁ!�y�`j��$����H��4@�aܥ��Mj�!\^�O���Y�h�a�)�����i,�!�$K���dPaē�8�D�xl���Wxc80à��B4���F�u��%#p� �O������7�Ў����ڜP�9�aC�&G^��"`��5�[��Ԝ���6�B+
��aC=,Ox�v-�'T6m�8�mx��U�>e��q�%�"��O�miE�4��L3Ta�SI�ن�9�DlR,;K28�s��*/�R�s����O6�R&�%Zs�lx��ɝ,���3�y!��p��O%qPԭ��ꋌ=>�bʎ48�X7��x?$���}��q�,D).�=8q�D@�$��&c�F��'L�>��+W p<jdk"c� �K�LK�gc� v,Bk[ f��+
�ce��]H�'����+��=0��#ǙE�Ź��-�~��#@I7~��}� et4Q��6l��{��2z�:��'b��TqB>D��-��'=4�U'��&�=zG��Xu覭'x-܉ҌM l�O��iSD͏,.
��@M�0M�R�O|j��Y<����<[�4̲��N��Xs�5�!��!>�l���/`h0]�SA���`(R8a%>�"��>����O���&�F�P��%�?{z��j4�����tY� E?W:��g'�)E���h��DߚD��Xc"�9�fȐUa��m�oh8p��V�$�$I2�l>#>)�e��f�*)���G�I"r�Ze�N؟�HV�0�j|�D��m�'�L���j�2@��Ñ�I=%�\P@��d6�)Reɚ&U��k2�(O���9B�0a�d
�~L������(6�j�!�,��WJ����=����G)3�t�q֌G� �h�z���`q�A�1����#<)2!޶7H���$'�'\�|��Ū��=ֹ�3�^�:�q���\��E�#��>���3��O?�� l�3)v�бF)�=n�^��v!Ğ�25�B��j�ɧ���Ǐm�I��eq���WnГ35|�	�A�#�޻DG����'-�ɸ"i��YI�1{�{�ʱ�
�+/�р��
�+�.�o�R�ҍ��ʰ&:���r�2�Of��M8OR�9�2ӬwV|@�'�i��m��x��'���R�Ƈ|By�7)ߘqD`�'�ZA��Z�!h}s��K-֜`�J������;[qO��(�լW��i���ջl��ň"O�}��`�(.��y�e��.'n��"O,����,h���ڴ< f%3"O� a�nT�)m��Ą�<���9�"Oα! Ֆ)z����c�8�<�1�"O>�K0�_ i(p/^�Zxx�#"OF�!5��%%F��"mߏ ��$"O����{�@�ǎ�GU\a[�"ON�1o��Q�@ C��$1���1"O�M��!�l�lt �F�k7�<�q"Ofd!�%H�-�B\He��*
���"O&�*�#��"e�d�J8���"O��mS�*�xs����>۰0[e"O�9���[��x����1s�|�3�"O�cs�ӷ(��a�J�F�tL�w"O怊q��/�����$�uع��"O��X��T�6�	��BŘUi�܊�"O��I �=d�n���>}�i�"O�  �X��F�c�H�� ��L	�1j�"O���2B��Z#�2�M�W�����"Oh��5��HH�h�E����8�"O��b���7kz�L��j���"O"q
T��X���aR��G�8�3f"OҠ���@�d���XÙ�U���"O�st#����iN�j�jt@�"O��Vh�.d������0A�A"O°���	PI��I�ʠ|
�"O�B�	�]v�Sh�z���[�"OfA�D�Rn�^|��G��BL�4JF"O����e�sxl��"���s:<���"OR,3��%V�8"֥R3�	�0"O4} �(����QD�g��}��"O��R�ƿ[K*1�tD��
G��� "Ob��у��`S� *��ͽ�T�0D"O�5�%S�12�H�#�0,h�"G"O�Zw�?:������0Ѐr�"O�=ɆI#aI��%�;�p��Q"O�1-J��d�r}]�goA:�y�l�"��Mɡ��1���@�H��yb�_!�Pi��ʡ2M��@���y�.�W��
�5/H؈�HY�y�AB="�q�[�7��PI�F���y�g ��h���ӼT�z���.�y��A���G�Rez$�%���yR��B���Zt�^������E\��y���DCe����
�(��r 9�y`�4!д2���+v��Lpb�B�y2�N:(Ӛe���n:L��#�*�yb	&7�<P��K�n?P(�rl]��y��H6
;��#T�*��=Rk�1�y�j��-�H�*��P�-����T���y�圴H1�r��#j@��j��yb	��-�9p��7&��,�ҁO�y�CK� "H�ʠ�eC�둄�'�ybdI�lO2h���G($�z�;ѤF;�y�#��2�$��c��N�������?�y��U�$x۔$$Bp���F��y��Y!T�ex&ȂC�X����y�>Rpe��EX�{�Z�y2�4��@�ɢOV�ȰV̞��y�J����8%�OL�=�����y�R�h��z��CP�j C�yR�3G�z%���]18�&@��ݓ�y�B��yC������h��! �yb��9$�$����U:��![�cJ��y�����eXM������Lsg����' �@�)�b���#`
s����'�y��y��B6IE�ocDx�6A֨�yB�D�DGSj�ӆBR��y�ȅl`rEC2����!11��3�yr/I�B�V�c,�f�c�bN�y��ݱoHV�qǈ���mK򦀖�yr� �leBCND�}D-����%�yf@��,9�Wz�<\ĭ��y"��g�؇��6s>�qk�MC4�y�&�5|:!p%(W�ib8����y��f�P��#�kp8�1�E��y�N�-j8��D�dW��bm��y��=J���&U��`Ep"�J��yE�6#���hD&ÊՌ�p����yR�@/`鰸��MƘ�R�#����y�T�Z)��ѣ�٨Ќ�O�y
� ")C�A�r(��͝H�l��E"O�m�E�J}�(@��X�M����"O�i �: � �2k�@�\uY"O������l*\k�	�]-��"O��P��4{K�͂�hPV�qs"O 	��D�=�~\� �� 3�x"O���%.�	��`$�M��"O �I�C ����eY"���k�"OZ�j j	�A��iZ�d��d휡� "O0�䐛l��0`�C64"Px��"O�1q��n&Bq�ϝx�lj�"O�!'�T�B2nT�S ݱnj�`"O�m����B��1�ÀByN��"O������`B$��0�*
nD�	2"O$�5`G�+BD��lU9Yn��"O����/L��0��߄iKlAx#"O�i!U��E�����dY�"OĨ��"O ����Y �d!`C�3QM�"O>�ƣ�y�V9��p^���B"O�+�[�&�p�j����-$Ԩ[t"O� ��T�(��9K,��$Lm+�"O���R(��+WB`HAi��^ؤ��"O� �tg��%P֐��	��GZ���"OT�a"�S���sE[�0�:E"OL5yԮ��nN0�4S'�A�Ǝu�<����Z�Z�BGb�Q�IcOX�<�ӌ\�Yl`ũ��jƒL1�IW�<���5#�Z���*X^>hQ@�RQ�<y׃�u_
��m�EI6M��CQ�<I��Ӄ
���*I�G����Q�<�v�	ۮ	C@O5c$��X�+\I�<)�+ܳ1&0�ď�`��)��|�<�" �,"FX� 
���ad��W�<a.�w�druU;W�	����Q�<Y`c� �ƚ7>���ç��I�<�� "Lxr��'�E3,FZM��n�<�eCR�6�@�׍\*h�4E��i�<���E>:�>��4�[2+�x��~�<)Ҭ�4����sl^�
=p��r�Vz�<�v	�c� �$��w�<�aHNw�<��,[-L�@$qF*��1Ւ�,Rh�<1wC�3]Ǽx�u���v����C䉙ܤH�!��1'�ܺ#A��! �B�I(�*�	����d���l�HB�	�� ����2f�i2P(�0��B�ɱ!���Κl���@;3N�C�ɻY.�a5��P F�ڸ|C�	*�X+mئS�Y2��3g�B䉙,;,�{AH��{2|��cJT�RB��9@��t���N[�$�����,XB�	�7� b��n�8��Gߐ:B�I. �P=*AG�bEH�+����"OR\8�.ǐT^�yä�,E�8��"O�%�OZ���D�T�"�r��A"O�U��|�� @��j�:�A�"O�S0��vu��
Rj%�FUBe"O��;Gl0���`���d�8Q�"O��i��;�H��T����b�˝'ؔ�P��'-J	��( O�$�(0^�H<YM�6L$��ZG�ȅ!��1GW���3D�GΌ���j���Qc��Qwji�� �|��P!�	4��	�M�;E,PL��	t��,�1�G�4�9���=(�'�daH#�M�U|LX���f6����H�F�S ��w��is�°^R,��c��U��p�I 4U.B���e�1�ӱ���f��"0a	��Pv�2=@�bFƔXX(HIn�v�*=k��aB����;A�@<tN��b�^�gz��2�'r� 1� jm�E���F��4(UM�/{��9�F\(B�$�H�Q���/\�;c�DޡJN���h�����Fߜ�C!��'h��BG��$oUџtSF*b��KTJ�t��I��dдM���:u,׵��̊E%�2m�  ��m�n?V��.,��A�UA(O`�"@�V(@�I�4� {�z-IS�V��"���udD����J�fU0���$,l�h� W��H��οA���-4Z�it/� �B�	����Z0�2]C@�r._1��x� /ʫ F��E�+��)C�m����
��0^G@��Ү���.�c��HP̈�!ƥk� �|��
f�x�`J.`�-��
��e	����1��!&ۢ��AJ���:NH���3�Ahe�3��u�Ǆ�7�˝$\l"5�D-UG�K^+}�0�)��Df�xt���#��e+t��� L�!��C2�\��7C��I�	��ZTö:��DۖfP���U,����W��I<�W�x�B�;- �����U:�5p�~��K1�VYеk
�5I������"��H��.X���I�l�T`Ҥ�
�K�G^`�z��v�	�FZj�Rӆ�4Qrİ�8P��<�����p	�o����,����Px��ފ B�!aC��*	��q�ra0"�� Zҟ�� O)h0s�@�ly��6D)fL"@��?j�J���!�"&iz���}U� �_�X�<J�V�4@$�7yz-'?�TI�#�,p�z�����n�-K��-�O�Dyc�A��S���!F���뉥y2��AD��>V�����=k��q�p�542x[�5~�џ؊���sP����-K��])>'��Ae	Ø���E��y"k�^7"y`�ѝ&Ru��C1��䎣9 F���E���)§;N�K��hb4�!v��x�`��[�@��)�.f"�aǔ���|r���}&�Xi��֘_SnɈ�l^#
�<��c*D��l��=�$�B��!dH����2�O�)gCIA�7m��+T(pqfջ\��i������!�DؕO�
PS��J(I�P�GC�����#��1)�����S�<�m�u���3�T�kDlk�C�2f�j͈���4hɜ�7�B5+�!KFM;oRT���<a���O ���٤c��Z�a�y��r�"O�P	��
��Պ���x�~�
��'���0�ܯ}�(�g�'UF�kTb�9.l�T�[�>�$�k��υG'"%���1<�0�Q-ΆB (-�'@ `�x��m�9G�p�i�}��CfK�m���%� �\V��U�ETW|��դ9�	�\��{����E����
 �LY�c�5��-�̃/��D3h���hְ��)ʧ^'�%`O��׸E������h�Y �,�K -�Ty���͔����Ƈ�<渐������{$�Yq��J`�3��){��UR�(�#9?f����J�!�X��Z$F�6�S#G][��?q!*�+m����"bp�����=��أ����r"$O �K�D2�0$�b��p�P��`��7<��I�g.I43��?Q���D���*wi>�I��[�4����U�>�=��۞)��t�s%�+��yl�3>�ޜڇ��,#l���7`�D���w����7"_*{ӧ(����� Վt��k3�LY���m�
N
V�XG��}�)��8BDሜr�(�N~��)0�"��	2<�(	�`Op�3�ɗl~H�J�+�\�y8�!�1����$KnxF�t-�6J :���-Q	JE\�%$��B�8`��y��������!���aчiF��I�f�LK�ɲXz�[V���,,��I�ޙkA B�	-�耀`�˙ z�����j�R�' �`c�GQ�S�'s� ��0C�X���9R�W�}��!�ȓ�f��c�n�|�iwcBn�܇ȓg.���t���	�e)`��L�ȓd$��w�cߡR2���IJ�^�!�Q��29)r���� )�i�W�!�dֳm���a�\9k6U���ɷ�Py��<������g�ޝJ�ៗ�yr��'Y���҆�\p��#aJ$�y2	��b����\W��q��GA�y�Ƈ3l$6�b+�L*FQ�q'ȕ�yr�,=c���7.�*:)x�J��y¥ʹuOd����4 �B�G�2�y��[� ֲ��6@�2�����
ƒ�y��B�5�\��ӧƌY��Q"ӠC�y
� \���KS	��z�m["W�hC'"ORE�®E9v�X�il�� [�*""O�x���R�x��ͪiNTC�"Oxq����R�1����Z(���6"O���X�.jmڒC+���d"Ozj�.\�Rz8�b�B�M�"O~�hUn� � ��u���:i�"O�����T�y���!>��A�"O:%3��5t�۳���{? G"O
�z� �w>t��1)PE�"O� r�dէzXT(�ۨ^�*�cu"OR����8J�|���]�e�$"O�hC
�>_m3ԿD��1�"O�Yڱ,I wb��t�Q�J��a3"OB͂F�@�e�$��PS9v^�
D"O,��#z��tb e �H<f<��"ON�[� ɣ=Q���q�r.^`��"OZ���,��5ڲ�].a2��""Oސ�"-�3X�j���
�;r��J"Oh���� �@8js� ?����"O�Ěpj�5s���B$��A�t�B"O"|��2D(�B��\��<5�"O�e!ԧ� #4yPƯ�j��5�"O����n[*ʐr�2�X��u"Ot��dOG,a�����s��"O�9�'T�9�( 谌����Ҕ"O,hS2F�9~t��fN�J���"O"��GO�rT�5D�7Y��u"r"O����n�-j2��򢘈% �}�"Ov%�V$L7 ��"��&35��i�"O��8b�
ẉ�@)�' �Y��"O�-��\�B��y��& vd�ѓ"OZ��ϗ}
T8����!� D�"O��� �v�zW  ��T;�"O�u8��
>N����W�4v�T�C"O�Iƀ2?b�1��]�#otlR�"O h��E;�B�Ӯ�F�N�8u"Op�p�X'~�zm�7L"�%$"O��׃�25����`�%k����"O|�;�M�#����Ϛ9�r0�"O ȹ���e!�P+DP-��lI�"ORy
3.͹��(YC#_Rc��7"Oh,� ��s =3���Nmbm�%"O��`eJ�&�TC�fP�\4#�'"�Ii'�@
T���"M��R
�'R�zU�S����=���@��e�<�ÍR�h.ź&)�Q��ٹ6G�]�<	Pk}Ƚ�bܘ���T�<��)�'g�z�lF�Mt��ira�{�<�p�8���Е���o� ��u�<�E�=��);��IJ�R ��:D�T�$G�;�x�J�	h��R�B�	 g讴�#��'^�x H�-<�B�ɒj� ��sAI
�R�� �C�I_��q�c,Ȱ4��a��B.[�!�5o��A�� ��b�إɡ��_I����9�����J��X
��=��	�4FNĳrh� ���#w�Ef�`Rp��+��� ��߸�yr�i�O��O8�� �("N8��V(@��JL����>	S�&�H�çrb�Q�u1:<������	�ܔ!7�$�	�ސ��S�&� ��iך��lX5�é}�O@ѠJ�Ӹ��O�rt`��\JϮ|�T/IPV���O�Trf��'����8�7(���-1��ݬ1������V	q��\(�M�������w�>N~�8$�	fJ����(�j(���C�1Oh,D���|� �L�e�=\%
�!ciT�w��u�"��4�����De��.XF�$�U�k0Υ꣌ۨ>N�Dps���G�^��*>˺��+O���Ͼ
��\�ㅅt��Qp&\0i�裀i�����8`1��?�?գm�!�D6@��\�L����x�dܳ#���QΎSt�!�ߛ��'	�z�Wn��xV�Q� &E"��yBh�,����$�Ђ/^��a ����y�)�M���	�:$R��Y��Y.�y�*O =`y�3��)"8�A�!�9�y�%�� �8�����):�����y��F?d��"�� :+R���aD��y�+�	��t��/E��&d����3�yr-�09S���:s x�/��y�^l��Pd�ӄ	���F%��y�J�8������՘�PNѩ�yr���^�D=���I�I�<@�7oI5�yR��@�b�zt,��H��q����yR�~1�����99bekP!���y��4��HAF`@�a�m�G���y�.����1���RI�0�g�)�y�iW
T�ƅ�� 7<)�!��K�2�y"��=�,�ɔLVB�U�5oC;�y�����}
D��:c����H���y��Ц}9�H#��Yv�L:,=�yr�ͥT��Ro�1I#��8���yRc0_�`�!�RI��Qa��W�y�$�r�MϠK��� ����y�-ԝM)f��2��D"l[QE�%�yR�. 'ęY&��l	�,8�JQ��y��6�D�@��)h�mȡKJ5�y"�7�ݺr"B6Z����Ĉ��y�IV)�21Yv�U�Mw|���`h�ȓH�$H+��ݽ5W�8�`B�1��P����!�Ds��Tu<��ȓT��[�L�Kd�U�s��C\T��ȓV��Ai���*��R2J�y�����x�I�+U�h�XB�Q*{a���ȓ;w<��5�Y�~5�@{��ȓW���k���^����!�[����ȓq��Hi&FF�?���C�5y��P��U���r�(���g�/9���Uڐ�2v�ЃC����G�,]�fA��%pɓ�+6P�踋��Ʀ���ȓ]N)��%�6$\�6�D�%\0��1]T�CE�@�m�p0�b�Z2� ��� �z�V>j��1W��RM�ȓyR���,�F��a�ԺF�Մ� �� Fm_:dp�C�.W:X�ȓ^�Z��Q�b�ܬ��8\��\�ȓ�������U�!�F�&�����Y�x}"5��$r�$�P�Dɀ<q�Ї�o�e��	,Z��r����t�X��9J�C#	Ѣ	����nK0r#���ȓOE����=���*S8ņ�f-�5��� �{w6����]�ȓa���!�ߣ{�T�a�u�t���]B}�!MBl�|Hr��/ꝇȓu��;V�ϲ@|8��ļkX�ȓ#d��f�		VH��Fƴ1�����zSp)C�썟d6J�	���
�\ԅȓeR<%�VB�6f�ѓD��~�\<��P!��7O5fq��L����ȓ **Wi��N�sP�h�@�ȓ��p�d���d��n���:=��S�? �e��Kl�9�-��[NU""OjZd��x���",N�:E�|��"O�5Z����qă*;C�s4"OJQ���e����t�!.rP�"O4��T������Yc�Y<N5�)"u"O.,��m����e���O"�}�7"O���̘�N�;v�1){� 1�"OF��F+�(Qp�̀d�.T��"O�f��m����a+�K�Q��"O�]k3�^�E�����
ߐT�*��$"O��Y�F�fzZ��i�M���J�"Od��e�D�\`.4Ph1Ƨ��(�!�O 7 �T��C̄g���V�(ie!�غ۶9��F� Å�;yt�4"Ot�@J��q�-ˮ} m;�"O:���LR�_KD	ZE-��1� ��"O����f˜<��l�*���"O9qcE](�T�P�ЂIݜh0�"O�-�Ҋ�0l[2��׭_���ա�"O �7,/�80gȬwrt�S"O*a����b���Ӭe�$A�"O�	3���h'�=î�m�n��!"Ob@n�!yu����40�����"OB)�4��v�u8���=!���w"O�qR��͚4I�5ٖ%�!@���3"OrY�s
�D�ؒ�J��~��a�"O��Cb��Z�ll���8v���E"O�%P�B
G����F�@,e�}�"O���&J�6/0#6�S2�\��"O��rBU�a'n�
&��#zvP��"O��PbÎ6p��単'm�-�e"ON�A��Y���bLK4/k�-J�"Oʈ���	V���rhM0h�C"O�U�㩀�о�2*ީK�0s�"O(pŁN��m�'ę�0H��Su"O���G�R�xcx�B� �%<>p` "O�t���N�T�9Dʞ :3���0"Oryjp��W,V��0*S(,�k�"O���ʛC6*��i�1v�٠"O^��3!F���#�'�|�F��"ONx� �H�R�B����	�_'b�8�"O�e��@[70V�yq&W6]H1 "O�E�a���?�0uZ%�6����"O�rb��N���9t���20h�"O�Q{�b�3�����9v��2`"O�)wn�N6ެ�4G;_^��7"Oz�q&�l P���Ҥ}]����"O�u�+
*/��<䀔*]*��c"O�I�!X�2gj�A3�цvU���"O���Ô!{S��	��M\	�F"O<m�eŐ&32�ܩWi[��[�"Oڵ�E�V�p������
���6"O�}��'�/lH�Lz�f�0R"��"O�q�!$Ę> �E��Fܗm�@E"O4�)��k��%���UkHp�c"O� �욄~��B�=U>`"OH�آ0�4$qv�є(8LL�R"O��Jh�uY��n 5�=�"O�����Ұ J
�С����q"O&���$a�d�Ӱ�Qm*���"Ol�r-�d��Xj�E� /�91w"O�(�[���A"�?,Y�T"O൚u�4Z��Y3�ƭ8 R�"O���p�\/���gc:�����"O� &yY��Z��y۔�U�\����"O� ���,�9 0�E� �.uD"OT��卐	8(`٤3M`"O�=���\5�ބ�n	7%�"1"O&���D�4:�:���^@{�"O*5�g��3O<`1�N?;�ˡ"O\4 f�>��0 ��W-R�G"O8�!"R�f� l��sl�!"O��)���0 ���#H�&�HV"O>�p�� ) �E��W���0�"O���d�@�q�|��4��'��:�"O��"B��6|L���d�zH�(�"Od�9��S+g:@�i���]��̘�"O���D��[�J1Ţ_9{�h��"O�y�蕋 �<x�@@םt���qB"O�X`g�(�n`��[�>r���U*O�h�����9��0qe��^�p�'��L���>\P�X�`�+o�<4�'�:$��
�k�ޡ�w6��iq�'{0�(2�֞=g�a��8A�pHa	�'\��D�h������8	���j�']f�³�[�c=����Y#5���'��I��;sF�Q	��K	Z� �P�'����˘�x��*QIжU�4��'ʲ$�Հ1n���0/�� H�ݩ�'���s�X� *�����!)�h���'� ��(����@�pd��s�'�؜���ɻ5̺0@b�ƭe�HM8	�'$���	\0�p6 �2\��Y
	�'`@��%�&�@z��X�j���'@1��˅|��m�WjK�NG���']�ʚ)T�9���Fv����'�(P� Z�L�i c��(��"�'�,PLYq�$E�獉/s���{
�'�lJ�h�<A�����q�,�
�'�D`��A34���h���>~�>m�	�'�.ᘄf�܎�7��td:��	�'�40���%n�h�������y���_T�=óOX߼h�v�U��y�	�6�ᢷ�� \�*ţ��y� ��_4`���@7,ep�K��y2!R�0�)��L�/J�PL�2���yb&$�
d�T��/p����G[��yC
�*;��A��W�#���8�����y�(֥��骱͘3XJ��M�y�N߇%�n�2��B! J@�� ���y�h�v������*f�Ax��O��y�օLJ��03�����e.ό�y�BSp��d���X>�F�	b�M��y��H�>y
�̃3u�,!�)�'�y�aI$�pݱC�!V:B�k6N��y2K�>����N;S0{�l�
�y��P%��%�b�`�n�Y"�T��y��R	V�Tl:�錑+H�����y������AV�%�j�y�C�y�!�Fw`5��3� �)��!�y2�.��j�� %�p�a���yb��d����/ǀE�������y"��%f�B�	W�_��P%0�a���y���" 	J)�w'�%jA(��ӕ�y2掉x�dC�$U
�Dp��c��y��u��]����{gΤ/Y�:��ȓ5���b�&~���ட�C���ȓM8z����i�|��Q&N	D�N8��S�? nl2V���"��!"�范H��]1E"O� �P!=I&���l�17��"O~]K#��/H�@�X��X�G��9�"OܹاAʳ	6�8����P,�z�"O��@nY�9"�B�Rx!�ɋr"O�\3)߶T@E*f�� Q}����"O�U"�Fʘ��2ta�'Zv�ű"O֬he���v�ȱ��O�7���Q0"O�]I��2f�M��Έ�9��S"Ob ��� C�\�nH'k��ɑ"OT��� Ao}�u,]������"O6�Z&L�/�reꗬߒwrZ�"O�F0�@sEVc4`]�"O\�I�q�P87�ǿR��� "O�!Ȗ   �P   t
  V  �  m   �(  �1  �7  ,>  �D  �J  Q  KW  �]  �c  'j  ip  �v  �|  T�   `� u�	����Zv)C�'ll\�0"Ez+�'N�Dl�l|!9O���A�'j�e�>=<%
�ǁ �pp	�JQ0K%:����V�E���r5掐9��"���H�A��?m30O��?���B�[,L�7nI6r�diq��6j��L�I	th�� 4�"���O7�u ߆d����'4$UJ��´l��̱&GI9�b� Q��v6=I��Ofi���C�oڦ�×��Ӧec����� �IƟ������b��Ld�`@2��4]3l�#&lڟl��Z|�a�ݴ����OV�Y�a�J���O:92�*E�h�M�5�2 @Ѝ��F�O��$�O"�$�O��#��O:�Z��'A��Ə{�6!���=��!�s�6�Oh牺E�x����17z(!@ F�U�,��Oz�	=��90�?1�LL' �z��[ N�H!	�O���O����O��D�O��d�|��w�^��`@��5��)�e��,��<��?���v� �o��M���W���kӐ�o%�M���-`1�(��q@�re�� ,�͂��I���G��^-Hؘ���%r��)����'X�����Kd2H'O�",ڛ�Dk� �o��?��"#�>9)���?��R�I�8:IZ#�O�,$l���4x����W�X#	X,�ɢڍ&LX�C�g͸YB�1ґ�iA�6�DӦѣc�8SQ���"�ʳ[yp�"�+�W Th��
�SR���ݴ��/uӤ9 rټ+W^��#�5_p�+�B���IxA�ַ,X0���ԂB�$h�*'�E���٦!h�4E[���
�0��K�.�|YBe	�PA汘D�űb�TC�'�=V�"t��H~���BFL�6m)jX���!	:�!	�Od�Ё��� 3���^�k2):�I6"�D�O�����:Dn�}��h��@��1c���'o�5�f R�?�,O����O�ӶS�� ���Ǉ{d��B������Ǣ1ˮLX(<=d�B�(�v��Pubs9}��2{P���$6�t1xh߈J�M2�H�R�L��A�@��'Φ�r[rIc�	_i�D�3�^,4�����D�Ix�S�'�y�*Q�ZUd�'�@�o#�Lr@����?�&�i��˷�-�͂�M���v�0&�nӲ��S�� Z���B�K�	��$�2���zC��$%��y�kD�WFܘ�F�n��ʓ��=�y�g��ei���#l��Ysȗ��y��|� �'Ȇ�f�08�W�yB�ݛ��L�4`�s�  "�N�y��޿*�Х��'�$�ĚD�[��?Q��U�����<�t������ވ&Z��:D�(�&��KB��y��$0 ����#D�؉����Ř2�G/I�@i�ք"D�Ę7�T&m0��[ �b��5D�Hd�"$���UĞ>u.U�� D�ܳ"+V8k�� ��A]��B)�<�t�x8����C1d �ܘ�hU� �<D�ĸ&j�=5��#tN�☉�4�<D�D���M!z.~�z��3V6(��;D��,�:B���xEh�[�r��D9D��3ufG�x�����H�e�T�۷�7<O�eA��I⦥�I�XH5��q�� K�^�x�����؟��I#"G����Ο�əW�0�#S�^��y�P�CgC<�cn�[&.s���>��@�O�����Kf\ <w�|�2�]�Q��1���6�JtSn͍� !1�͇[&�B�+I72�0�?�V��ߟ��	��M���'� ݐ��	nh�G-rJh8,Ob�D$�)ʧvf!q,��z�%�5�_<��E{��I!�M�T
߼b�P�+��G��$t�Z�9����|�C��j��``�D�HC�ӯU�irSI�tAV���1D���`�f R�X�I
ILc�/D����LN� ���T!]�V-3#D�8�����3V�aK�Z�-��02��"D�`�B�Rd�y�b؟&}&�xF�-D��ӳ0+.���l�"����6����Y$�p9���?�Iٟl�ISya��Ap8p���֘u�"���@��bô�s��'_$�7�V�j����rk�|RR�d���Ny:���a���b�8Ɇ8���=�����i�>&^c��iQ�y����'o�-����/ɰ8K�Ɵr�����i$ʓ4�Լ��e�矌�I��I��.���¬��H]L��AT}x�����P�~��S ��[nE��I]������e��4���|��'���ߺc��4�	�U�@k%'�61Ξ,�Eg�O��$�O��ī<�|r�! 1n"��2!�n>�@��KX<@�(,{�u�����E�\��y�*℠�r�ـ1(��g��:2���cԈ�A�-1��A�N�y�����c�%���"#L��({�TR��?ы�$/.�ZB/N����pD�Q�l��ȓb[��`/�HHP�CE��6�%�`�޴�?�+O��(Ƀ��e��ȟ�U�:�j��3�X�|o0Y2��ԟ��	"g��)�	���'���s���OO��SS�O�0_��� �8hTE�0z,�b��P��	��'�P0���D��H�SצC�( �����pgZa����nr-K�Q��0<�
�ğLcK>����'v��C%��29��m���E�<	$m);�A�	#15V�B,HC������
oԚ��#��xP��޷9x�'��p��7�M�O>�(�����)Q�0x�!�I!@�HbV*T�c���O�T{g(L?Q��m;�.�1g�,��)�'y��;C�}�
�Ӱ�*\�'��šT��bl^�33�N �>E��/��"�h��Q�7D`�5A2?)������	h�O��D�"�X��ƭ��҆H�\�!���J�pZb� J�!N f������V�O(���F�ݦ�!�ݶ�U�ij�W��k��?���ߟ�IiyL	K�2%3�F"j��EJ�1< �����(d����m�(��`��D֫d��8� B�Z�����T4$�c�(��;E�$:��N�
ݚ9�%���:�p�8�'��L
�e���ę�7b�u����i@��'�B��p�'V�dU�l�	�D�	�1���;�+�8&��Ѓ@e��i��ȓE���@DIƵ$�N@P��S�jҽ�'(l#=���i�S������``��A�W9��4#��DU���	ҟ���񟬗��O�����֐r�IZ�.������7v�����A����x�6<O	yBG�I>���`�:Cz�tm�_G��&��hkDzG!-<O��D��_1�P�e�-�x��~'2�'aў�Ex��l^�yA�o�j"�CU�м�y��X��P�ra�$v0�ȴh� ��[����'��7���B����d��y�,+B@�l�J��3FP4�����O�T
�(�O�$s>Q2a�D�&����"܅����I�"$r&C��C6��E�.	����D[+ ���C�  �ݡ�H�OT5s�	��V2T@@�(K	}o<���'������?Y�O���Q�o�R��@)�"[u8�)!�|"�'aaz�ʾq�pI����@ޢ�Q7m@���?!��'"jIRq矟R6dl]r^�����d�<yk�1�'cRY>Q7�ޟ�`��;<<�i�S��q��	����8����Zx�;sژ�R����?�O��ӌ4�z�RT�q�|!� Z�PNN��\���ů+�$�ߴ�h��8(£�g�T�C&ӊc�8Yb���:Ч�O��D>�'�?AJ>�!��L &29ٵ-C=�y��L�.������L��������OD5E����~0as�ƝQ^���NV�L��	Ly�Ö�h�2�'1��'-�Ɍkʌ�H���#.��=���6�lĈ�΁tWX����C����ɂW�g�hkJ���/��\�B�Cb��w�వ�]0�����i�$��U�g̓FF�X;��L�z�E�c�D��f(�O��$Ŭ	��ҟTG{bM�����3q.D !���W��(-!��s#V��#�FYxެ�d�8��I��HO�)�O�ʓ\�S@�>R� ��� $��`q�����?����?�������
5�)����RN��X!�É6n�&��A�BE�@�S-�[x��/=��H���� 
�,��!��>I�t��O�oQ�����v|��Ưov9���S�<�9�P1T>�IaA�'���	�'OpU0�Ɉ�\ޝ���^�@�m��'&� W�ݳr�����M>	�V���?�AWd*�AD�3�ԙ0�(R;Z��]�W��m�<r��.0��|�%.�6~��F@i�<�f+n�Š������i�y�<ѧŊ�O�$��W��/Y. ��u�<уhHI�$�6�N�~`�{�s�<)&������b�K���8�(l�'Ott���D�J�rL����)MV8E{�bN�u�!�Ĝ�L����i� [)�����#�!�D��FlJ�z�!�o>���c�R�!��Ә<�Z����>\�ȻҢ�Z!�D׎�	���\�]KN�{&#�!FE!� ��+ei�}I
T�U�����͓ �O?� ���>,��A�f٧c\x�k_s�<�P���JX�ka�ި�k��[s�<1e
��')�لgU�|(��Ts�<�u݂YE�R,D_��@�b�d�<�B�hi�d�rT�x@�bb(B�	�Z��蓦[l9��0���9�H��N��I�5����Su���@�^�9	"���S�? �eJ�$H.(�
�K�3��tئ"O�d[�딚h���@0���f| 0:a"O�h�9Kh��RlNEt�J�"OR��ĭ�?7\d�PG�ާ�\����'�0�'8����ID>k��Ku�NA7��1
�'�����CG��氺�9����	�'}���W'�(�AY�1��c�'o):fG�[[b�[g��,8�	�'�̈i���,�^��K�5$@d��'}�P�6O��y�w��`nV0��D��WkQ?	�i�?|!ئ`��*��񲕀>D��z&O<�<�x`�	/�6l�g8D�8Z�L��?��g��\P����4D�<���d���S-]H{��$E-D��hg%��!��!�'f����+0D��J��M�v/����M��~|�� �-�O$� �)��m�`�Y�/���nML<��"O�ѹ�@�g���5/��|F���"O�J4��a�5��F�xZDD)�"O&8sGl�6Er�ԦE,7y�j�"O�`q��N ;&�I�!�I-" �Q�"O���F���p�hhg&M�w@��RT�<bTN"�OH�y���!�`*�d�1/�YAr"O&}A'&E0$�h�+E���A����"OzXYS�G)w�l%;�S0k�.!��"O���C)�����U�+3����$"O"m�� �|�pQX��/	�X}�'^����'��=�c*��Lۇ$E�Y||ez
�'�(qLԄN�ޕ�FG��M(&	p	�'�:(�e��5��%Z��Y�E����'Wr2�C��6�5��[+9����	�'�@�B��Q^P ���ϯ2u��c	�'�z���/	q�"ݰ ���%yh�1��$O aQ?YI�O@�Ɋ�k�d�R� �2�0D�p�6�[VX@���8 �Y'G0D����%=\<�1�^�B�@ "-D�pYp "#vu1'�Тc�̀��8D�\W�b���O�
��a@��$D�Au�EU)2��jL�,� ڵ#�O�ɪb�)��r��rC�	�@Y��M�"i�ȍ��'p���d�Z�����u+Œs7:�Q	�'�f��SD����K%-$g�޵��'.�������1V%�6� 4��'ID���m�)l�|HD�?)�2�"
�'eN�:0%ņ8�zYQ��^+����,O���'��Y�����EP퀕���r�'|$�iw�W�c���� �[<ā+	�'9LA䈹$
���B\���H�'v�i`g#�1f4 ��c���	�'�C)������D�P�N�6�	�1-��_R������&��\�%ʄ�<�T��B<hR�ۆ�� �d�T<���ȓ|a�l�CڍOWJ�Y҂�H�N���Ct��IA��%x+�@7D�t9��"OFq�c�=|���B��-;�|$	"Orx�g���9�����ᑭ �$�F��.c� �~�% ȄX�ЂI�}�A(�M�<��X�H� e��a����LS�+^I�<If.�Z��1�3(��=�6�(�BI�<�H[?A�{ACB@��C��^�<Y���'g*�S6�J4m�IY]�<�CF*t F���(`4ɩ��؟�[��#�S�O�݊�H���I�	#=_��k`"OPհ��ͧLfTE3�m�>d���at"O� ��:�F�M1�����_H��R�"O~�+��#|�����	l1nxÕ"O� ���Ǯn�f<��  }��"O�����GF}\���3��ܡ\����#�O�����1��5o\�H4�i�-6D��25��$�9�p��'f��u�3D���cV�;�(5�F��T����.D�Dj���/Q�ը�ɀ�/�i%�+D��AC29�|���(�/e��؛t
+�O%`��O���&`�t�ȫ�F�lo�i�"O,)�Q�ڳd�A��#_Z��:�"O0�"EI���(@ZE��cT0A[�"OB}zq��^���i�$��2tEQ�"O|=+4��_��3&e��#|��`"O��K��*pTRa��*6n��@�퉍l�~�� Ck6-Ƀ�ԫU�œ�	�p�<@F��u�xҕO-`S��hk�<y�DZ,p��I�� �S��p�	l�<�2���7�4)�Ϛ&.�5d��j�<�4`�0<����3FC\�
����k�<f��=c� (V"�c��-�D�埀*ĉ3�S�O_�h��T��<�`D2`��-��"O@!�Bʉ�U�����	����0"O���eG+n��UC���r�R�x6"O~���	a�d���c�`ݎ}��"O����� �����!];v�ޜ�"O$��Qj'WFUj��u`|���S��㢆7�Op�q`˾�a���B"��"O���Y�o�x}Q���4�Ty�r"O`�8S�áxꥠp�
-���+C"ON���c�%�-z�/x��T"Oʸ��˟#w+����L��@ڥ��>)1�Z?��gٳL:^�o�V�TӓaUO�<�E��Q�����6Q9����h�B�<ђ�	(պm��e]���!�L�Y�<9E���s$���2��#/�����a�<!�� �bi��o�*���Md�<�b W�s��8��R����t�'/T�;�����A��l3-T2��e�E��W�!�D
@���H�ɞ�;}����;Y�!���x
6���&��j�h�b�-H�!�$G(XfHè�-lyN�y%!˾D!���#�A�E�8�a�'!�dK�9��P�6�B�i��@	���d�:�O?�
��_a��1��4��}Â�z�<1G�^�|dICg�-���r��r�<��%_����4�H2�0l��� r�<)���܈\�l� 9���(VD�<�uDQ��h�+�=
�����f�<��W�z<���3�Yb�2QPt��cy��p>���M�H|l躢�߂/�pA��G�<���P#����񤚁U<�	I���E�<�叕q���
�N�<�H�H5[�</ʆmML9�ƻZ� D8�.�S�<�L[�.ܴs���^�D=�a��Qx��3�f����Ā�k�$��T��+=-Ll'@(D����@�~����g����$&D�@§���iBd�BJZ�k[u���8D��ˤ��6l�dT�%��$�`��0D�\K�I�������tY�X*A<D��K�� #"�0J���!-V�cm>���G��R!k���r-�<rDB7�y"B� |�D��0`< �c��y2��h�!�v��U�d��Wc���y
� ����J�o� �)3d"�ְ#W"O` ���ѓS;z�C�B�6Rt��a"O|�3RO6@�Z�W˃2lL����'z�����S!Q�>�H�N«z!l�Qw���1�ȓ3,t\K!�āw:p��r���g�JІ�#�Z�#�y��邖IЁ1#"���JӾ	s����l���H��ˀ
F@e�ȓCV���F�*ZU@��Q��\8��u��3u�0:a��A!g@3F;���'?y��r��1�C@�~FVXS%����@�ȓ}�}*�A��D#�����Q�ȓD�άG&Ӕ�\ ��!Νp��)�ȓ?�؁h��S�t��ꖪ!���ȓu�����(ÜD����-����I.r�`�ɹz��,{�jղi�2@���H�
�B䉥A��D���%0PZ1'f�RC䉿Wa�P����:^,r4A�B�	�|���ʥ� <�1�`B��^�|B��;T�X|�D�P
0iw�v����2D�h`f��8]�줱�#��PK0b1�:�fdF�tK���& ���IYC�|�Q�S�y��R��f��5�A�Swl�Qa�*�yb�
!.t퐤b�J�����P��y͕�YRqe�Z�k1�:�Py�T9&Dk����~�X�-UH�<As� 
)�(:��_�~�I �`ǟ\k�N0�S�O(���F(�Fa�"lԆZ-G"O�����=h�� �O"VI�P"O.p��k� N)��+ǯ���(�#�"O��@���>b)����;����"O�%Qch�C���'$ )�#QO!#��x�"]�C�ė�D��'�O��'���'`>E�r�O�����?m;�)�#d��ZC�
s���ɷ�oy�'��'�n�ke��`�P�@�9Yc<�4�8$["��,}�X��1�\�X�.�"c�	S?�͒�&s
��\�4�
y5\���i:���a
�ԈOh}@!�'��P9<��	rV*��x�h}ڷ�K�kl�i���	V-�2�0Ę��S\��a�1�'�Ox��'8��#�P�2� �1T�*`V�9�)O�Ag���H�#�JyBV>E��ʟp�Ȏ�\c�)B�f� E���"�!PߟhH� ָC��cg	Q�"r�M��S�O��0Mu� ��/�:B�m�'��ʝ�&���
��,	��?9sԇ�J�()�P��$7���u%n�Ĺd��On�$6?%?�'��0� �E#B$B� H)6�r%��'V�P�����T���� Y7�E�]p�'>R#�@�,0 4ez��ؒak�,S\ے=i)O��ʇk�O����O��$�<9���E!3%R�*hu�Ć>|mJ��4��]�i.�h����-���I@i���0N�-�A�N25���`����@�E�)�j�RR�#Fx�&Ae��<K�ߑ_��ur2*�?��d߾#���'�ў��Z��}��"�< <
��dP21��	�Y�mK�)~f����d.���.�HO��Opʓ��bfM7��p�"�υs�,�����?& ֨�?9���d�O��� �JP�/a�9ↁwT���!$@)[��U �غ^t��@�s�b�YV�K���1��m�k��'x(�܋�쐆./���ϓ{+�\�	
'F�� % �6a"�j4k՞O�@�Ib�'��D�v�X�~Rx�B���q��� ` D��:p��mbl�pr���\E �R�̼<IB�i�Y��I5Gҟ�+eD7�q�E�(5�M�
� ������O6�D�O�\K�b�1}���2Ə�7�(��i>M�ӄ�!Z���*⟢1��Bք*�r�K��Ӌh�hZ�@����IG�z��B������@/^L<��PV��O���9擭!��zA�A5o�q���-��C��0��K�6�R��w�׊L6�=��!�OD��'�v�U�_�����+Z��A�O���'Jv�1_���O���'��<8s)o-�1L�����'���QE��~��F-#5�R��7;�(,�я�}\\�pG��|��/�U�ħM�?�i�CZn�O/^�8�k����.D�E�\�`�'�БH���?��O�O��)� ~��6�a��� �޺h�s�"O���"[�?Հ���(s�Y����ȟT��R�Ĕ�48�EU5W��H
Ѧ@�Q��d�O�Aj��̅lm����O��$�O�L���?�+��������0�AՂUԊ��ӌ�_N��(���&R5�Ο���Q��!fuʰ��iHc��-T�*���E���T�@U�`���g�'�q����D����p4<��Of����?i��Dy��Ӕ���jP9$��8Wht��DJ4D�4"%L?AL
}S�,�e�	r�C�O:Dz�O���$RB��8�4a�0t��ڳ��:���P�p?�ז9HHi�'$^{��; ��]�<�4��<;t�"n��p$�u�d
R�<�q!A�<�v��1��%FP�7��Q�<�gBR�/�fy��Lν\�&�:���S�<�%FA�D�L�3#��� EW�'#�1mwӊ�O�KP�*D1���V�m����<����?a��{���I��YL�Q�M֜�y�O�$D6ܪJ�^Q���T%�Tȏ�$�X�* #6/Թ�b<�Тڒ;���U��e�v�1%Hz�E����M�6�ȍ�$�\��'���'��ڃ1klxS1.^t}ڨ�/Y�Y��'���'��W>�GxB$�`� �A����0�� c� ���>�_���4.�,5�8�T!+9���I �<I��3��&�'%�Od"�� ��2h쵢�.'Q�H�r@.O��=�b��P��D�R��.=�s�U�Ep��&�ܣD�'��S�H���ԧ�q% 4*@ʏA�|�hc��ΌAs�S��':�D
�(LS���
�IH�F�%f�q�'@B�'�p�J���H|� o�>;>��a@��/����Q�X�'[���B��yBo�&s���f˙ft��C�l�m�,lJO��O��Y �(}��~�� v���`�	�g6����� Xl0}�IV*���c D�^��-p���Y�(�2e�O�x�5�>ƛ>Y'�Iu�d��U�����WI�i�W��Z�xb��<E�^���[�O��tr�'q�}���N�l|IA�趟�s�,}*���(:��ɋ|Ⱥ�E�$�m��Ae��<�'� ly�m�<��'��eF�t��F���Yv�V�z`���ǯ�?yh���+k=?��y�B�~%����Ts�hÝDm��̙�?Q0m,�O$�r�P05\�8�&�	9k��B�"O��C�͙<)LP���&: ���%�i��Oj˓���Oh��Y�<���s�E�$�U��ѹ4,��m֟��	y"L�~I>��%����>X�$a�̷���RpN)�D�<!O>�~����?{@�h;SfQ=hx�� bN�<9���a��M�Rc�#�Ԑ��SI�<�f!�,�@���(�lM���H�<���QX���`N�(�i3��B�<!!�ķ+���*a�H���	��~�<	�iϮ6�����F	4��T1@�N}�<'�J� �����E�YlU���x�<	g�T����%)� �%�~�<�Ղ��29[� ϳa'�}8#�r�<��ȗ	e*���˹���xLAj�<	0@��os�p�@·5B��USh�<�3듇=�Լ�r��9��,����f��ll��i�K�3#.�B�l�c�Iģw�Π4@�#V�^�:&�āy�����+] 4���%k�m�pl87iM�
�
��F�5bΎ{��ɛE�4p,R> w|(���W�d�x[�JQ'm��s�aL=_$�y'��+�,r֍ӥ ��@q�\�-Nz��.Y��i���H��ml��9|Ze�T-�
nְe�^���x���?afă jcy�R
F�|���$���	�~��lGF0xT�$���5�YY�	�&q��	@�Q��pӋ�U�OFT$K����=��0�g���eZ��J<q�� �|��4:țv�'D��r�P�b¤t'�a/�14M�عv���O����،4���)�'@� I�#!y�x��3�h.��Ån��M�%�f���r`����Z3\���'s���P�eߤ��E�W}���Y�'��e�@�]gN8t$�>F��'V2�*���	Gdށ�#���;)h�'|���"��{Lr1��jɒ.���i
�'׺MzF(��y%���[�$O.�	�'&�@�*�G$� pM��T�4�*	�'�j5��CI�A��L�wY|�A���� �����$U�h\KDmыV��9��"OV$[��
)�����iՠi���"�"OJ$�w�@F�}"�.̯R~����"OP<�PG����TC�mIU[�a�"O4�i����`ܰG�]�<"�u��"OL�{C�Q�1/>4Xc�_`�
�y�"O�i���ܒ��GA6��y�4"O�����Jnb�8���7Q���aw"O��'15�K/,�4!�-�y���g��	Q�ϯoM��:��W��y��حms>�z���� � "�Q�'��)��� G�i�@!W�JX�y�'���{"�j��Ȍ�vX��'Sb��%���Ľ��ィ(��B�ɢ[~@qr�[!p_�4� �֯
�jC�	��V��*͆~j
Tɓ�#�dC�I	����Q�%����Ug	�/<�B�ɟD
��0*X!$�Z�,E5X��B�O�:�a�ܴ?YR��&l��B�"&m��+�V�O2��6n��a��B�I�s���#��8IL��Ї!ϴ �2C�ɺp�X��(B�v��({Z/cF1��G_*%8 ��
1֥�\s6|�ȓ6��YAƢq�F�pU��;���ȓ&kXMa�LP,*����!O¹\�݄ȓuPS��ӂiv�Y[�n�+����8�yw�7g����g�-�v����h��nW0I�ɢ�V#;G��ȓ l�c�ߨK�l	+�G�m��]�ȓ&�h��j߶��WMC'R)dȆȓ��q�o�2T�
`� X�p��ȓU�hh
V�%w���Zjh	�ȓJg�	2G
Q�Kc��0�2/� ��Iu�=H�e�1��1�Sj٬X>��},���ɜF��0�UR��VT�ȓx�*�R��S�!�d����om���dx��a`�� T���B�R
X�� _�5
Tk2�:P�"�d�ȓ*��t���TxX|��KN�*V�ȓY���w㍢	��H�d�&�n��ȓ8���0�C�(<`a���7ę��k�l����/M�g`Qz��Y��6�<�ga@�K|Tpqv��E'@��ȓf��s��
]�i��b�):"lM�ȓo�rh֣Z�X{�� C��&p4���ȓw��yg�ۅ:����WB9�n��ȓ>Zp9�6cK�0�� @)
D�ȓ	���G�
�ib����%n��ȓ(O�Ygąx���V\:Y2a��gv �����i�6YB��4̄�|b�I�1ס'α ��N%�����Y�Z�W*̈́�V0 &D�m�d�ȓ�A#4�3<8ܳb]9"�b�ȓY��	8B�U�.���`	4W�d���8������ד���(`���j}�ȓFH�aäB�o*����ł��昄��j���n���H!����NC�H��U%�m`3l	�ab��4蚣?�$��R,l-��1|�ܝ��Z:]�e�ȓ���S$� ��ȣ3d�(�=��8��
@�L9u�����Q#z� ����u��A�m�x�R+߇4�؅ȓ�H"lU�t�Y�ĉfd�a�ȓ\��`�6�S+8�l	n�'�y��S�? ���R�'R�)��	�0T�"O!�*,�|S�D�&=nF���"O��`h/�D�h5�']T�%K�"O�:��$&)pq)��,s����"O*�ʕ'�>-�.V2I[��8�"O����քY�Z�v��s���y"c׀]����3�X� E��1Sa���ybya6�O�RKtl�$D�.8�9k�'IB SW��/8��]����:80���'rDyi!
�C��u��OIbE�<`�'L����O�=0S
	�B�CU�9�	�'34�BÃ*
���aB@ 	�Ł�'��AL�=F�Y鰢\.v�,}�'0�H���9�,1eL�,l`�M��'R��G�f;����V�g$vX��'�����φ��]��.���'�	2� AvUY�(�w���'MlP��K�&!��D*�����'Ix}� �8(�8i��> ��K�'ςX�6	սc*��$��F^�̊�'���tC.>����TN�!i^fܑ�'AVEr�C��U�p��Df�P���'W,8k9�z����S0
�c�'lآd-�z�.F9JlȨ
�'�jXhaE��d(}���أDe.�	�'6L���F9Z:X1E�/<{n�Y�'�R�r�j�,S�^U���'4�-�'���[�
�r�c��#6O��'���@I,G���:/3�4��'��E᫔��-r�� ����'��4��JzD*�����Y
�'p��V�}����s�%��+�'-�|��(D_Wpqj #��q ��	�'�"!"2HU'=���y���M�IR	�'����e�]qD\�2×:��=��'���0ॊ|��ݸ�m,kJ�Eh�'A�IщɆ#�Ș�!N�\��50
�'�`ҁf̬9��h�R�E ��}p�'�i+@A͂��(�5c���'��� ����:��� :� 
�'ƨY# ^P.�5"�.�Ш
�'�LP`6Bֵy/)H�K�y���h�'jj)�WK�<��u v�M�^�X��
�'� `�!�S61��`r���;C�P3�'��=y�HE�L=���?e� ͨ
�'���B���XZ��g%����'���ٳ�F�����0Δ�k�l\k�' f���k��!^���qN)�'����5���Y�j�C#���jXiJ	�'~
qJw�S�}�0�rH@�
�2��'�D�g�D(K�"�x��\��"�'U���E���(V6Qy�c X���'�jܢ���W,0|;�Cځu3��3�'���(�&T")�Z�íR���'g��KO?%Z�}�tb��Cr��9�'�q�3�ɂ(�Nu�C��%q]tp�'s��a�F��	T@���P%U0���'0��"C1N
��p5Z6��V�<��F�6[�����t�RR�<QRoX�`Ӻ��"�Q�C��O�<��ɔwu�PӨʆ]�t��ae�M�<Y��my$���cq��0����G�<q�m��_{H-��O?'����G��|�<�%�,��r��J?H��qj%TP�<� B����p1(�i EK>{�@,�C"O� ����"V�)z���8w����"Ot�s�G_0�8D��^�Y�=�C"O����nJ6��1�����]���jC"O��1��)x���av��d�DI��"O$�8c� 	k��|q0IH(c`6���"O*��,�-��;��6>:Lb�"OĴ[6
Fo�E �,�craY�"O�\ 
W�6��Ì[�v�6���"Oj��t�M*pQ�9��M-
sp�#"O�����@%_^,�T ֎)S���"O�!�o����e+�l�q*`�cW"O�Ē�Ǖ /�1��k4�F"O�L!�/�=Sen�k )BT��"O�H��GK�K�4p�GW�y��T#"O
tB��N
=�b,��� ���쓠"Ol�&`�5[�Ջ �]+�K!"O���p$��-pF��n�_l���1"O~�凡k�����:]�eK�"O�,RD�C�R��0�q�;2�Ⱥ�"O�����X����[��"O�aV�jTb!;u�_�RZyq"ORuA�.�9�� C얆=�1"Oxy�4d���`E��Ri��"O�� ǋ�Q��|"�R�֤�d"O��%g\0��}� ���WS����"O.�
���+9��Yٓ���)h*M�"O��+�e��,p�j�[��F.]h�<�w�P%d�!�@��^���i$��b�<�aʕ�/@�i�H� ,��h_g�<��G5X�<�їHR�L�������N�<��-ݎԊ=2��ݑ\b���iK�<������*���-@��4� @O�<��vkN}�hH^D�z�R�<��Ī/��Ъ��8t�J��ZP�<au(uq�XR��Xc�<:�F�D�<Y�N�;P���J%]�l�WnLF�<���T4H,:�c4!��&<�yRE�<!VaV�|�Je��LM�rrq�"nN@�<�'�K#D�T�(cS*�@k�A	d�<��)"E�U�4���~6F(b���k�<�������%�Z�iV5�VHP`�<��ނ�4 � �<Ar�[Cm�]�<a1G��:Ԫ�Ǌ��j8��̘c�<�aZ�2�<��!#=�ji��b]�<Y�� �V�t�D'B5\0P���]Z�<!cf�*�r�hG��{�h�7��|�<I�ċ*.3���5��Aj�RD�_�<i��H�>�t0#� ����Ge�<A���?�����N�Cf���� �a�<��g������*i���K]a�<�fX�-��(�s�UI+jD�u,�^�<a7F[GM�L"Q��f�̀���QX�<�#��%? ���(��Kl����l�<aD��j�`�����LP����]m�<��	71s�EQ&�-�djck�o�<�.�*b�b�+\�C��k�<�H*m{����틜���p�h�<ᅋY+qP�s�!ؘ~��;���`�<Y�ո3���g�jE�q[��AC�<A���4"����Bޔb�r��a�{�<馋ʳ=ebg��4^��&�P{�<�S��u����JD%DX�b��*n�YŤ�*x��TcB�M?��<�����E���)"��"FC���g�<� �<Y�V4�H��aBKI��K%"O(��e�H
<,}����N�8��r"O���2��"��$ᕶ	��Y��1D�[u �4F�D�x�/M9P 3l?D�<)�-�	"� �`L7d)&|���=D�캁Mǰw��
7@�k�+0l=D�@!��O$s��A�b�C	k�P��:T�L
2K� ���:#�Я8'�=��"O���B�=��i!OO�nx��"Ot�z�ڿDa�P�G.tr��"O� 條�Uߊ��&�!5z8Ӑ"O�E+&�T��CE&Ĥr��I�S"O{��0`Ý�@�K�k�"O(��1�
��5;vZ4��"O0��7��o_>��Ǝ]82���d"Op�Zg�U$�����Zf��:6"O���U�_�<yR1��$}���"O�@���]�0�B��jx��"O��4��9/����]3"O��r@"O��bFւSvh!A��L(yL�Ě "OX��"ၹP���DN�$��09�"Ol��4L7�qJ�ʚ�n��K�"On$  �
k��d�'H�P��u"O:���,,KZ�Jr׻"�|ّ�"O�m�FÒ "��������P"O��0C�؍���c�E/Q]P���"O�噇����(�M���
M�'"O(�U!��|�'�͜w5�3�"OZmyv��nmH����>{,$�x�"O,8��;]H�ۖ�ސPXш�"O��r�� ,~�Q���^����"O�T�B�+������ǟ9��i�"O򀺖`Bn.)q��<����"Oj}p�)	�Vq�$�I��h��"O�Yx3G�%t�(0�A�L�H��"Ona�$�«���#�2tԱ��"O�ɫ0�И'{֙s"��4,���Q"O�m��T!%�d��d�,�8 ��"O�{C�@6a�歙u˖7:�F��"O�����/ӆ<1���kd���`"O��A�*�S��IZ���e����"O`��&F����;$`M�x5"Ol������hd��*�LR+��TH�"ONU�d�(\���a��L�	? �s"O����"b�Pѡ���R!���s"O��#S�ik��������[r&��t"O���6��"l�H��ը�R%��"Ob$�A��.�r��t��A��ԘA"O����IN�E�|\!�$�x�l,D�`[f,O�)%��'�:Vq�m���*D�ZQkM,�Ѝ@�"2y>QHT�7D���E�^�2��P��R�zU�&F4D�lJǅ�2,�B��0C���L����%D�4"���&k�P����M0ڀ(�#D�9tEX�H��@ p(H%fU�H�t(<D�,�`
\=P��#© q��@#7D��
�W�5�5:v�A�xp`��ǯ!D�p#4�I.i��Y�E�%�.D�D���=F����i��"E�.D��� L��?�иՆ�|h��#+D����x�<�Q�C�*�J|0�º�y�+�Dp2�ǐ'Ac�I��y�h�=V�z@ۡ!_7o����2B
%�y�̞�?`�� �DIe\��L��y
� dz�G�!]�42�m�%�^q��"O���O�c|
h��Aـ�D���"O63$�Į3��Lc`���n�u@v"Ov\��϶ތ<X���xv��"O�4��H�$F]�g&�6 (�x�"Op��MU.X�D�3Х��xoX���"O&LKs䃄?\-�q��-lm��"O� �0�V�Pr S�-�"\b���"OF���#Ft��@'Z��%�"O^���k
e�3���B��7"O��q��a�X`m!e��h�"O������`r� �d�
���ss"OA��E�C��`J碊),���9"O~Q:�ƒQJb�C���O�~��"O�j�KM <;�)��@Q�^��e��"OV�J`�����@g�T�����5"O
�*��9�h��u��u�ȉ�"Ol�a!n�`?L%8s�َI�pbD"O�(	�ֹar2\����/���*�"O��hU�4��E⡤U�?���a"O8��J��i�
���y�ܵ��"O&1"ծF>�p�$F-(�L��"O��8vNI�oHt[�ŝc`���"O(E�� �.d��:�*K,:���R"O�a��"�J����J�?�F0��"O�I��PrR8���I����"O�MX���9r��)�!�ƃl�xĒ"O��b�G��Pt<���Ĉ�z��aV"O�}X�I��7�|JU�����@"O1��j�<K��Mqqȗ`,hA��"O*m["�Sv5z�(��O9�n4h!"O�Q�"Κ< �j��{�%�&"O�YB�կN�ڑAg���j˞1µ"O&����
:����m��k�d�x�"O�T����P4%�!�ε\�Q�"O>�� ̀ݾpu�	xpt�h�"O�C� &O��@�dȽiu�}j"O��J2�\�_��4@S�N!<_�,�"O �c�l>� �r���t5�u[�"O��I@�1�l(�t-�	*5k�"O9���C�� ��!�I"���"O$A�KN+R�ڼ�$�
�jP<�5"O^��H/}ώQBR�u�d��4"O��#Aդ,9�ТU��դ8��"Ot�S��R,
��T#c��h$1�"O�A�//PҼ-����aex��B"O��%�-�|У����)����T"OL�i$�O'��)iՠ�v��Y#B"O�ͣ1��[��ҳ�	*p�C"O �0��\4I��h����2Jf�K�"OJyPT6Lw�$	�Ɵ�O��ل"OT,`CJE(}"�p�M�}[��X�"OrL!��ҏ/��Z�E`�a�a"O$�7��w����aA� R>�|�$"Op2�O�Dtp��P�z��)�"O�����+�F�  *),�P:�"O��צ�}Z|X�5��#?< ���"O�\˒�ę&{���)@u�"O)ڥ㚼-���t̜�CN�X�"O��9���:4�R�J9Xn�܀r"O��;��:��%	��"!��M�"Ol�
w/Ι�t! ��/ ��+v"O�(����D2x���W�L�P}��"OV���kP /u���v�<�����"O�  �8A�ڨtk^x� �
��$k"O�D�S�G� �c�ƚ.Mg�X��"O���A�[�tnb���W�
�"O!�
ەO��#$�.~�L\��"O���EJ��%�^�h3N�J5��"O.��9w9N�j�
"	4���c"ODT*C��(rl��#�R� ��r�"OD��B�/��8���L��Zu"O ��&��AŐ��@�ʏ[�Z<�4"O�Ic�AS�[P�
E�_�|��8Z�"O��p6N�)���aP�%~��xP"OxqꥭY�F�<� )F+_4�l�5"O�⠈N �BY(u����$"O(U�T*��=|ZT���=.�9�"O��W�4��$��c+!.�ԻP"Ojр�CL���s5��l�,X@E"O,%0�fڸ�D [
Z̨"O��˃��]|P�X��\�ޮ0�U"O��Å���Q�$İ��4"O���e�*=�5��+!9ر��"O½!ra�E%j4#P$��)4��3r"O�؈�AH�#H�1�ѺA&�A��"O<��! ��Z�.y�!Y�u�y��"O\yxSJ��U{
�����uH����"O�) �T
f��A�%J\J�"O�A�����%3�	!�mʓsd �"O�p!�I�4���#�,�'5c~=P"O�D�`��0(�ޱ��������E"O�!j���`�B� EI�<Y�L�#r"O�Ӗ��]�B�hO2u��"O�]�0�E�U	0OɞzoL]C�"O�0�D��U���"OX-Q&�����Xx�+��"O.�0��Z���U�hY�X�%"OL�a��K܄@閦�v�Ly��"O Ű�잒?��Rs�L�7;l`r�"O�l`@ Uv��c˞q@�X$"O��n�7#n���g"�Z�
�:d"O���ʅkl�Q��@�+u�=bd"Oܡ�����p*`J�~u�)3�"OPmXU΅(DLJ���,e�4�&"O�-&��;:��@�SM���"O������n�8j�!U�Q.}Z�"O�)4�l��D��Cv���"O(=�T䀙o�Y�'�]�� !�"O(3'D�,�|�1���'#V�ɡ7"O�j����Y�)#�t (4��"O�!����+D�l-��8q�"O�)�5lG�Ρ{Dĭ�����"O�X(���2)N���%D�$����"O����s@��$�:=ִ� C"O\p)��+gf �zbk��Jθ�"O�E(C �;@!���Q��!Qk��c�"O�M��!S�
(��NP,w���X�"OL��B�V��x� �V�p��1"O^���G�`���G���m�""O�K���gM(����1W,4S7"O,!�ń�|�8Y@�'Q_����"O�%3QC�?;G�\QC�.MK@��"O~�p3) �lwT|cv ɛT�ڥ�w"O@�TNZ�
��ī��[�D$J@"O� .Qm��Bu���h�8�KQ"O0��OW
�$� թC�F@�2"Ob˳O_	��A��7����"O� �Ի����l0�'A�07oʽ�V"O؈��&# t��9q��"OmI��Q�^���nE FT����؆d�������$b@=<O�l#�%o�l9vg]��d�6"OF���)h� r Sj�hHc"O�V�4g�64Y H��k�r-�C"O�����$���4H�$�jjS"O��@Be�"n
��F<,0��I4"O�E2DۘrtiyU(��5+d"p"O> ��?����2�V�}7TUJ"O�!�BS�%���@�z�1�'"O�Q�I�"�D�$dÀg"p�@"O
mS���94��;UBiEZ�"O��gF%XZ�zFl��Ld�"O�Ҡ�����J���+n�q��"O�x��$̰*4��:R
�ir���"OF�y��מNWոj��9� �a�"O��Z��N �>����̆t��\��"O��ɓ-V�<sV�J@�
��¤�d"O"����-�����M�q�̼0�"O8�*1ꌍ|r�q7L@�cȈ�1"O�a��9>҉����-��xv"O"$XPFZ48�0 ���E$���"O��P��:&�����<Z���BD"O6�p�E�lм�Kw$R�*��(��"OvI(ס�r_�J��В�:�f"O~��-] Z=�:!�[��BL�7"O�)�@��[Q��h@�"~'8�8�"O~s�Y�c%��q�\&*
��F"O~]sb@�#���d�v����2"O�x�t�9@Tx��˭9����"Ojja!���`���\"R"O�� ƀ׃u�t�#+�/��d"Or̀@�Â!ӐH�'	��=�q!2"O�B%�w�j��1AF�euD��B"Oa��^sZ �)r/@Fٹ�"O�Y��$��u@ �k��L'-.zD��"O��Z֍�5m�xaI0&(z(�t�6"O��D-� 5p"���W"Oh�) ˈ�2�!I�&#?ܒ�c�"Oh(��V�yL�*��҉sf��*"O��󫊹��|z�q���[��yB"�	 �p*�"Ϭual%�6�L5�yb���0
P��Y�m����&��7�yb���v����Lh��l+F����y2��K���)�H�2wɠ��
.�y�� �z!���]	Z��@&KN��yb�����p`�E��VF��5� :�y$����X�؋�E �Ѽ�y�Q20�xKt�ó�8��DC�yBi�85\����
�u���Xf	�yb�Q������R>k7P(㰂ݨ�y�C@��eB�6c�-i`�S�yC�lH��%�W׮����y�f�T',��'ăU�&�Y��
��yi�
��9B�]���$Ή�k�!�DL�
~=�&�I�|�)#_�R�!�:-�>��CMޯ_v�2�5C�!�D�%G1k,ӣ����U��'��Ep!Dg�2�KE�"zƀ�'�����Ŀ4�P|h��^����
�'<�u����q�e ���	.�|��'� l���0ឤ;64���'�8i�KFU�XD���)���h��� �L��=v�H�s�=���d"Ol9���)$=�E��f���H�"O���4GKs����c�� B�H��"OL�[q��?���ӡE �|��ɩ�"Of���,@�Z�����P�5ã"O@h�cJ	���X�J-g�8��7"Oֹ�%�t�:����`�r�"O�p,��)On����$~�0<�5"Op\��/a�u��Eçr�.iZ$"O�\0��M&4b�h�u%�~�|-��"Oȅ�5�tkbB�Ē}��"O��2�,��u���c���T�d��"Olh�
�`(�� �K�U�j��"OZ]h7K�
h=�pujҕ���c"O�����ԇ,Z,���+�f5�	�W"O�L`t ���D���E-*�Z�"Op*�;*�4����VfIr�"O��!�ӷa���X$�]2Hd���"O(��ԊB� 7 M9���3�]�y�'�,!c�=c$D��*ӡ�y�#�/Y��cE���7�p��S��y2�ù?�P��-�&:�r�3#)�3�y�mTA,��K� F|�{�L2�y"�C�8�E�D�W�|��|�lۛ�yң@9�<�r�B�9!q,-���@��y���5�R���JW*�rx�����y�/�!) ��ʒ\�P`p�0�y���*u�,s����BO2Ya�h��'O�i:q%�:Y�jU��+N2Te,�:�'7T��BP���<�퓄Wv�8�'�����B�΢|�E�Ҟpd!S�'�.����}�d��*L
r�p�
�'^Θz$�2��a��G���r��
�'�C��;((��J��b�2�'��,�ܲ0��9K$b�J�а�'Z�<�gDC9��Y*$�
D[40��'ᘩ2�A0U#��T��3D��ݨ�'��|�����ɨî�@��P�	�'�Z(�Q#:5hXaC��	#��X
�'�Z���F�'e�$ܣ��0����	�'9* e�I!���!�:���'����˒w�t���XG|0�'1.\B�E�hÎq�&	���'�^R���(���f÷~�fb�'�"@��h����[V!C�&I6z�'�x�B" -G�&�c
��'Hf�P]����&s�T�!�b�<�2�V<PZ��iW)B�T�UFEX�<���E�"�� #�|Z��i�W�<YU�1:[R�d��4 B��x�<�P�ޗ��wL�2>~�+��A|�<if%�(q��i�$�.��u0�{�<�A#D�b��.G*m��e���a�<���Վ@hl;��J=R�H�cPh�Z�<!G.R�F]��-�q�,T[K�J�<�Gh�F�����\���IG�G�<I$V8Z�#u��G[�`�M�D�<	aL�]�j��qF�8�lt�3A�v�<�&�E�K@kw�W���عрAs�<��.�<U���*5�,|��y��Zr�<y���}!�uʓ��1Q��ckHm�<Q'�Hp���� =�9�a�n<Y��v����7,�(9�H��,L��ȓI7P�c ƓX(M`���C�)� dm���*�����E�0!h�3%"O�A�EU�	>�=c���/41��"O���!Ê�*	Z��ŀ,�Tj�"OTț���1	�n3C��!y����"O�� �>oo���v��91&I5"O�M2R
6��@��ŀ ]	�"O4�C�JJt}{a�[�LZ�HP"Oj�¢�W'"�����Z�I�"OX0�Am�;~F�s����BŹ�"O�D	!f��Q��-����"O�Ix��S)�2E�♎�����"ODi3�+�k�D�c���!�"O\�Cd�ahA�⍚$2�R��"O ��E*R���9hEl�(0��p"O2�K֋N#q�Yp`ȊQ0�$J"O��K��q� ˆg�6(P̡d"O�RU�R�$�����GS�9�T"O����D��)ӧe	:jeS"Oza��әW�A1���5�J��A"O�(�0�`(V3u�U%�j�Jp"O��QK�i��\�%��pn5i�"Oh���9>n8�0���\j��kD"OB2�Q !�Z�Z��ƞW�Y0"Oj����L��6)h��ՓR,U��"O^���>:y�`vB�D8S"OzHZЇR/DY�v`D�z=�ua"Ox|`�O��p_!���I� >��r6"O��f�0�Ι���̸p�2lpa"O�I�̲6D �@��2��u�"OD��R�ʳA�N��%��A��=�2"Ov�
��.����љv�I�7"O��� ��|��0R�V�6�$�rb"O����h�ly��/����ɴ"O�Uې狠{����T�T��f"O�h���,��,*�n+S�,�h�"O$�9�O\�iT�a!�7�ؽ�"O\=q媚�>v|�X�Bμqp`��"O �ɲo�v����5�;kn$:�"O�bwQ�M���(�cX.~dܭP"O���2�דV{�$ ��K#gh�SA"O6�ɳHB�	S� �Ƅʃ9QUr�"O|��0��8��T��[�@�X�"O(��G�+2]��Dώxx�	`"OQ�a+H2=�P�˩t�@EA@"OTm#��:����C=f�(�X�"O�1���(14��c�YN�W"Of ��I�VL�J�aC�uB�	%"O(@ق��#��%sr *E�e��"OQ[3��8'Dp#!38TX�#"O~�%��!j~,Ђ�R�u(B�T"O����9l�d:գF-|��"O��� �&+*4�7�<���2T"O�1�5-��z���*$bJ�d�H!�R"O��{�I�"��Xp��9���Rf"OX�a#&Y.'D�jsς��(Ӡ"O���6'��J8Bea$�Z����"Ob��#��xEV���^*{�l]��"O$٩�Mں(غ����G��9��'P���X=W���6�M3.[����'"�"U�]����&�*��l��'���^�X���B� a��H�<�lM��x�;��	M�X3��i�<qED֩y�攙 !�O":��f�q�<A��T�L���ρ_�hA�c^p�<� �$�����~��$2���,a2�0�"OBU�Vٸ>SP0`OA$GY "O��gK�txT��d�w)dg"O�PTl� O%D���U�\x�"OԸh�<��%b�59bR���"OXk��Ì1 ]pA'P�p��ɧ"O���+Y;/�N��	? 2y��"O���́D�j�95�[�M`�"Ovx*q�G9Q���
�C tX��"OjIc�BU�wb`���\�kp�`��"ODV7+5p��(�.�!�&M}�<qѧ\27R�z� �R4��Q�Dx�<�"�y�
�I��E5���)UZv�<���\�\a�ኃ+.|P�U�\M�<Ɇ�k�HAk3��*��8���L�<�U�P�&�r|��2=Th�@�O�I�<I�o�0I[���cOE����sh]G�<Y`� ٬��� ��� mNo�<�gH��RsA>=������n�<iD��KE䐙# 	�{����O�a�<����h�� F��12���G\�<q��-DF�Ҕ�Շn����p�WA�<�'�9��b��ȟn�Jt��|�<y`�V_���ɶ���0}��Em�<Y5h�5]��7lLs�6�+�&J`�<��� |�����@�b, ��G�_�<����i|�A:`!�u�(y�eL@�<��h	qޠrr�T.)�̉��-MW�<�M
(dtY�
B�V�,r2H_i�<�E���  �Z�m����e�<��f\)2L"���	1Z���`�<�R�̶.��qӅaY�_$0h���T�<Q�MIq$ryCg�G#m��5�v�<2F���Y���V�����Rq�<y��GuˎH&�^�H*�<�R�<B䉚�Nt�E'T�7Z̸���һPC�I�_@d@�gՏ:\�Vd�4Z\B�/;�(ً 
G�oF]�Ąê*�|C䉭��!(%��
�vɠ��.]�C�I�g�rK�>wN
|;'�$7o8B�
8�dpMK��p�B��T�FB�I"0�����^(s�P�a�=�<B�ɾ<���䒳 �!Zn��"O��q�T�f'��6��.�@��T"O�9���'|M>$���Ys��˓"Ofp"3��$�tq)�ˋQ�$��"OzD���˸D6~��	�8૕"Oּ��΋u=��FgL"=�,ё�"O�	��Xa&*��`���4Y�`
�"O�e�u�^�F�<T�S%��8H0��"OfH����#Y0��s� *6lG"O��Ѥ)!�N��"]f1��`#"O2��(� {6.DqU��5,��"O ��Ď���HЗ�9�"O��R�b\F�fm���x���p"O��+��\LRK�j�C��\3�"O�,��4Y��h �#��~��X3"O���C�W�8�n��#D�"�`5�R"O���G��K*�hWa��#�<pB�"OJE�I�(*�(H"Nˣ�����"O��Ɂ��zYt�X���/�J`@E"O�2���Q��-C�b͑ �Q�@"O���P�,D�(qwa�O��g"O�\җ �
5���� Lt�F"O� ����MQR�jTɶ(��m��"OJ��#`_�e+`00bY�A�}�3"O�)��� �\��&��f���"O�t�k�H�00�C\�<4l�X�"O�Xڕ�m4��0D��WKVY�"O�]B��F*���8�a;|Gld�"Oz`xϊ<���0�a�� Iٸ�"O�1k ��u��b�5�>���"O.}�d#%�m�2a+ְA�p"Oȹ��h6���RQ�N����2�"O:13���k����NH�k���j�"On�h�� �4+�ٲ�!D�j!��"O�-��g�����̎�-nl��"O����U�|�hT�d��
X�� !�"O"	y4��P�����IZ�d�R�""O��i5�ԝ�8�h��Ȥ�R�S�"O��8B��t����'T����ړ"OB���m@�B��A�%U�;<���Q"O.U8aI�n��i��E��)��hB"O�Ӈ�+e$����8_ =�`"O�$!�n��aZ:��1�^.m. �)�"O�ຖ�G
%�24t��@&\=:�"O"�C���PX��a��F�/�|	"O�U��H��6l3aƳ7����$"O:��
64rdT�`,v���W"ON��S�d�0��T	C	L�J�"O<y#a�E�X�aj�>&�*��q"O�͠�Xs�%�I��@ߞP	"OR)�5C=�$�y#��*4��0"O��!�)Hs�D :��R7QI�!�"O��E�wH���g����p"OHy�FE+R�*@k�f�|���1"O��sB)��ELҘ�ӅQ�i"���"O<튒��&)`���G%.Y��,x!�$��<�#J<
�.!�t�
��!�J�V+����(�Űj�(~�!�D�D��x��� 3j�u2b�i!�D�?.0�I�3�g�T80'Vx!�$��k���y2A�'kl>�	�Ɨ!�D��@Ѽ��J� z7<X;�,[6!��,��zTOڱO)x��*��W!�$��u�60�����ZS	�%(X!�!h:��Ё�M<	���4hX��Py����nE�5	í_�}Wt�������y�"N�5��q('`@������yG�:~`��'�Q�:��a��7�yBM��Tx�*rmߥ\*��q*K��y�,ǦB�Xڗ�ɮ%ܮ���`E��y2 �	iU��ڶ�R�L}h�0�
E��yb�Z�nM|��=MS�u��Ӑ�yҪJ'Ebeq��Gu®�i�A��y����T7NM���ʲzW>IY��ۇ�yb	-:Th�[��a)�P���y"$ԈP�*�AJS�XE�xצ��y U-`�\�j�ٖ|��-)V�V�y��${�����`�"���e]��y2�����!�ĲY�D=���ɽ�yBL�lC ՘�CD�Kj�,����2š�$�<c�tx��AEw*�paEO�co!��'1rq�櫗8([֭h�D��_!�d<����.T^���e��	\!��:C�ZT��∨so�SFĂYP!�$E�y�ZԌtm���!$БV�!�DE�8O����ԫLVF\��	�9\!�� ��f	?���@2 �ic�"O���'�^�Zen��J��I��"O���W���jE�Խ6,`�"O4���dC;}o��Ӄ�x��4"Ol�A& �k'�1�T����5�t"O�h±�T�1��F��s�jAB�"OZ��t��;c�!�Ty|�`"OtuiT�ؽ8���J�GN�{��"O�|᥄T3P�(�@FMχ�@)��"O����	<��P�GmЫA�@�4"O� �ыћB9�A� ��LiH��"O��rŉ��8���L� Wؑ�"O �cSa�=c+�>���V'�9�yb�N���r��B5`p^���iI��yRA=�<��A��</�H\���:�yb�Ps�&m('��sO�\Y㠏��yJ%W;H� �S�\�J�	�۾�y"�~]N
򋜓P�}�#)���y���(gb��-�^fX<{V���y��Αl���7�J�e;����\�y�a��8�4+G�E#Z��)CR��y2�O�
��YC��'g�p+�mМ�yҊ��vB�40��z:0`x�N��y���]Вx�)��]a���S��y�ݲ@�x�Cv	)Q(��"��y�� CT���܉T�����)�y��_%T�8w�>x��2��� �y��I�%�T%�*ţg'@�g��=�y�D��U^Dc���m����&�T�y��L�A$��v�X>�y��6
����%�O�s|:��E���y�́X;.�飂�y�l����yRf��e��L�1ɖwn�8u�0�y��q|R����
�ەc[��yR��w�p�*g� "I(D;����y2��WڔE����_�Ԁ��9�y�GE63��D�V�	.-~�GM�,�y�`�0?6H�pa����8�*�y2b��6$��`c�V�-&n����Y��y�/|�N�j�k�`�i`���yB;l���O@>\7�u[a�-�ybB[i�*��^#}��qk�-B2�yR��� � `��z��c���!�y2���e���/IA��
C̗*�y����D�H�.�%��Y����y2�X�+�IxtH�a Q?�y��W�l�6=au`�0E!R	�V����l����27d0�Q.݊�ȓ:f.˷�� Y����f"m\��ȓs��H������elL�o�ȓw���`ƠT��4�I�3���ȓO4��dh _��`w�؝N�RɅȓ;q�L��O+��y�R�M�%�i��?�����8�%(u��U��x��P'F4r�Ø�N���`�J'E��y�ȓ{z~t�����41�a���9f���ȓy��� e��	~���KG�Ha�ȓ'� �q䂓�wI>	-�<�G$R�<���!�����|Y���L�<��X��ё�EK���Ї@	M�<	 eX�=��M> }�H��OD��y��X9+����&��.an�j��y��V5�4��b�,��ؘ�'A,�y�b�S�� ��<�،h�D<�y
� ����N6���@Ǔ�-�H��#"O҄(���#E!F)J� �+)��u[�"OF�I�,�)B�@��S�^s���"Oj�q/�:T���׋� ;��t�"O0������S�1��4���K�<٠(�dO���� 'z�N���*�K�<Y`��?/ĢijW�U"l��GʕI�<Y�g�3>�=� �S�V+j7n�D�<e]�=p�U@ѥ�[��	c�L�<	"H���[���Z�м�0��I�<��#(f@�{�ͮ;
�}qC�C��?)��"#�6�>E��'�(�鐊U#79�� � /� �he�R�2�X�㐣�6��đ1��V��]����Ͽ���
Y���6O	o?�p�c
�㦙�rm�������G��.�z`!PJ�s��5��	N��]��A�8�D�t��49��'`6�Ҧe��k��M[a&A˴��mH�Ig�9�mf?Y���:�S���]!���!�v0�`)��(O�lZ��M{J>��'�u�ޜ{��Yj��VQ�6y��M��D��mbde�d�i�ay�
��U.)XF>r�lأH�?�.�Z��_h��u�D�ǎ���*��,	��d��3���:�&�@T����E̼P<���i1wq��K&��9'1LcVU?9��HR(�(��O��@P��$a�!P�.���m�Q��̟X&.�۟(Sٴ_"J�gy"�'��	�f����^>�u��)�T3,�(.Ol�����	��-)��è.i���݃l���ikL7�Od�oßț`k��?��O�R�K�nC�}����Ca��u�q��7��l�G�'�b����
�KmL$���JF�\�|����d��� �'}��j�,ZP�'�2F�4��2�)2'\�l�[�&�{f��?|�� ��8�^h�6��"^��OD�Y��'��D�k\q�ށ�F�ɄC�9r�nO v�7M�OPʓ�?�*OLb?= �iE����{@�^�c��{�̣������T$��KѸ$��)c�)T�>�(�R��A��#{Ӹ��G說HEmZ��M������w���#�jͣ*�*�`�kV�q��@��Ⱦ)�����O��d��4�@x��n��*��=E���q�1�OV ��F;@r
1��&u�q�����͉���x  ��}�f̲W/N�0ul��Y��K>J+jA���1�ɭh;f�$Eަ�޴�?٩�X�{ѬH(A��Z6�[�*����$��d�)���d!Ύ
Oh]�7��^��c@�6�O|�o��M�ܴ9��]����'w�*�1Dd��8ŌH��y	���ֹiF�[��S�?%��ؗ%�:u�ac�RL�X�!�ʆ}<j��ѝ
�l��%�l�d�#�S�?���:I/l �c/A�*��Iz�W!�Ht �x C_)I5�4� d�e�|-@0�1`��\c||�K� 7�q㯗h����4(ތ�	�LZ�4�?����i�|eH�ޙX��D��o<J�����'��T��E{*�N}�ab�]mZ�,�*0�.���ɶ�M��i��'=8�9���,�Ձ֍k5r��t�Ucu椛$�՟h�	�X�.)R&h���\��՟���
�u��'G��.ɂ
��E�U��('�#"G�A�L���̑�\'�x�c& ":�D{���u�����qJem�Qא�h3��u����b([�C���h���:*AY�_?�se�J�X��O�$a�e�|Kd�ӏn�u��ӟ @�aIԟD��4��gy��'���k�*�fȮh\��$gL�k���<�˓K 0[���q�Z��0"����b�`�nZd��?��S{�̦�;s   �   K   Ĵ���	��Z��tI�*ʜ�cd�<��k٥���qe�H�4��_?8<�q�i��6m�i�����X�p�Ո&�J2m#0�mZ�M�@�i�~��v쓞�䜀A�]����u����흐Pd�ZF�v�	��{r�D�'�N|m����$��AA��h���:5��M���6�ÑtI�˓}��J�pd��"b �ҔJG��Ȱ����:Q0�8~�t��b�0#���/O��8�Ba��Ɔ3�G� ������M。Bk?��O�x`�'���c-xB��	�]�
a�����(�8�kF]���	����`'扴7��8�DU
�E�K: *,��B
��$ߞ�O��#����8x���Kv	�
_w ���k��F�Gxb�w�'����'nn� ��xD����L+�4y�M����ɮ8qOf���/WWN�7䆍MA�P�t�i��Ex�I�'L�#!�Ʋ�B=ە+Ӈ��tq����'��|GxBJTd~��.'�Iᢋ"~ �h����2���OZp���F�`Ɔ8����~�T|Ps ��!���Gx��RK�'mx��	����5�<�p��]3_7�L�F9�_��D��xrL�
�5ZG�\�Z��AK��~��E�'�v�%�8��'��������f����I�LD�5X�q���OC�����	�OF���Ӻ�,�Mu�)��M!�FQ���K�θ'\��Fx��j��In�B���x	�a%��,��ɭ :�����I�,v��T��x��ˢ%�B䉹Q�t �  ����f�0 ш_����'_��z���I�O#G�S.&��&��;�d�$��.�y��'|��'b�'�2�i�?4�,�J�(	�ʹ(�M�<q�\��O@������qUkp>I�	�M�N>�r[iM(6��5%����!����?���|se ��M3�O�\��A/uX�١�/,rqѳk�Cs����'��'��I���	���I�t�M:S�9)E|�Q�T�U��������'�j6�^3)θ�d�O��D�|�7j�v�PG�*+b
4�Ip~"g�>	��?H>�O�VL�#v44:u��S��M�Gb���Q�醊S���|:���O�5�H>Q#��{�|���"{*$[�._&�?����?���?�|2.O2d�Ӆf< �xW!�4p���+Z�!h�1`҃�<��i��O���'�2�WV���@$-�}td]�qگ`�P   �	  y    �  1&  �-  4  W:  �@  �F  9M  �S  �Y  `  ]f  �l  �r  &y  1�   `� u�	����Zv)C�'ll\�0"Ez+⟈m�f�`�	.[	��D��v�P�o����#e��5r)���(�>^��9���:U�$�S�fa�|�;,t�����F�&����a�d�h���& �P��ڶ$�J b$��+ym��:E�ұgl8�HޜҜ[`��운ៜ�dG�	Q$�S��
=_������R����k�`��T�	��f@��煟QC�- �45�@����?����?	�.�����bB�cL�;#�&{be����?���'{^�:F�'��'��0�Cܦg�~��T�F3�<h3��'�:��A\����,�r|��ϲ��'1�韶Ђ@��#� p����w�ͨ��)�O��ɹ/*�-�Wa�{~�b��97��꓎O��	�l�=���?�[�4nd I�h�Ĺ�A�O����O����Ov��O8�Ŀ|��wg~�1��2;�q���NC2��w�fMq�4�o�9�M+��z�V*lӄ�o���M[��eO�Aq%aʌô=�e�Ѝ^;�J�Od�F��/-",�Tio�[/9Vnc���	�lr��	�47���j��(o��?��S.#�z�2!a�RU^$K7	Y'F�0�!�M��!ݴ}�%�m�r��<�� T1p������'��s�Ȟ,"�#d��80
����'	"�'c*��ճL͊�o/�<�XbP�'�2�'\1�ZՁ0���81���2¢v�5�uQ�DE{���Z�V��cA/6 8�R��hC�D!��?����˛�?�#�؇R�0h�T�Dlq �O�˓�?������ę3:vrb��+-��3��i��Yb�B����d/YlD����'!�ݩGfK/F�԰"�&�-1�B�>Y�x���[�*GN�ԏR��0<����0�ɇ��Έ^V�I�ŵfе� G8��'M"��	f���@�/Q��U0$*I 6��#�%�O�}o�.�P�
�c��%z��O�AJ��ٴ��'ߞ�f��1�ՠ� ��j3"�0_A`e�t�<D���BKI [*�ȡJC�6���+?D��(�J�k�^�Z�HO?:Ī�i1D�+���v��HQڵE���K�#.D�dysgD)o�Y��ْ���-D�8uČZf$�H� D��-9���O�1S��)�'!��  �o�!j!I �d�qC
�'��q�� 4XU���E*J�S�8I2
�'� �`�)��9}��ꃰG�@e		�'^��B'׳�<Mp�j�
Ba����'�,a�1�Č6�0!� �'�BY��'���#�F���ʧ@��8 )O��s��'_hA�t�Уj^M��kϥgq��(�'Sr�h�Äm%0��\����'4�0���L� ��C�ՓL����'��1)�C��Ix\X�xv,]9�'��@��G��ł�������ϓ��H� �i�I<� ����Y�k�� �l�(s`��$�<���?�'|̠�P)������<6��f�BX�!ǝ�@Ԣ�J�ꄬ�ax2&W)� ��#)cI��'�*a���W$`�٘3��I>��ZÓa�"��I�d��4�?�+ɖ_%�0 ���g,�\�p�^0����O�㟢|��
*I�|��E�Ĵ; £=!��d����#7%D7�25�H�"Q�D�d$ŷ�M�J>A�	K�Xy���O�j�3�L�ҥ�eh	XM��80"O� #%���f���b�ƍ�s.�-�'"O����DQ,n~��f��S��4��"O��C��eq�݂�R�5�\\#�"O����	�̑�`-B�Xs�ȋ�"O x[�@� x�����>}~�	�c��O��R���2�$�O~��<I@J�0
�0)���b��@ڲ����:��i
�6���^��%�|"��DT.L�d!@"M�s��X�*@&2k5��Ȍ2C8�d���C�`���s���Z�'Y����+�>��cCB3Mf8��i��ʓ����{�矬�	��)L�^�����H��L���yx����cY�7'H�C� [�HT���+Q���Ŧ���4���|��'��d�w�`�HR�S��B�j��J��t��O�$�O���<�|��#ެ6�D���	�]�93
2��8`�Y�O�pa3£����ybkT?{��͛@c�H�V(���2$��s�X(>R樨���||��B�H�9�HMGyR��4.�DY�b��\�@!&f�������?A��d1v�8�S@^�
Zxۖ�R�l�ꈅ�(0�M����1�^PBaM� =8�%����4�?�+O�5[d������O$^��t�,��8RCg+衹	�0h�1Ex
� �;A�Ғ:�����M�B#��!��'�Hdx����8�֭s@�"5a>LY�o=3�ax���?�ԑ|bl y�\j!�D?�
� t��$�yB/�P_�=rrQ@�(RI����?��'ƺ�sp�9c�p�a��%ՠ4J>!�
�ԛ6�|�V>M���l�Ť�Q/ЬA���0���������#��쁃�,�^T��S�O��B��Ҡ`�*1"ScS9 �Q�O����@K�2k��X�J�n�ޢ}2F�����l��E�y��� �_m~bC��?����h�l��>`*֜�2��+KĘ@�G|��B�7/������8Oϊ���QG���?���Sp�|��׌�CTh�G����mZ͟D�'�P@��O2�'J_�����­}�j�je�օ��x"��X5�X�Ti[�<�Rk�"v�|�<�')��5�@� �=x�50�,Jl�<H�%��<A���@�|\�|�<qW�G a�XeX�/��Q[^� fɵ�M���?�Jˋ�?��'��$�O����O0��V \_Z����G�F�Z2H+D��j�D�H�Ƞ`�;?��L�'�<ن�		�M�����̃it����ɱl���� ��\�X�C��O����O ���<�|jb�FF��a�R�?��h��+S�lD��YQ�)�l�Р(ì��yRB���Yb�Ouc�Q��ʄ�R^�U�� ��y$�W�8��y�f��T���ޏ|e�r!�D�(,����?q���!��0T�O���L!â
�i�ڵ��u���{ՆP7dH���!���%�0�ڴ�?I+O0i��W�S�
���0	H�\1	��2&�$�<���?���|d��{QƉ2f*���j�����_g�nIC3F՘K�.5{���0<�FԁƆ�v�P-�<p �����bA[�rd����kĽ8�n-��I�
�`���O&�8M�<�$EQ�+�b����
���'����O��x�hQ5c.���M�O�F<��*)�Ol��I)+:r� ��� �g%A�p@���<	��)��O����'80�����R�6i�q-҆f�&�+6�'��Y%���i��N5F�	9g(�O>��G�� ��Q!iβsl���$.?A��S���q����m�,LA�����o�V�F<EBք� W8;�	y���D�O��}j��=�f9�WA�<@b��@ɞ$GyF�*	�' �Er�.�.y�.�;-�G)�i��$�E�O嘝k�'V�{|С��kY�c\R�qf_���'�
��'}��':"Y��y&�T�/b�]Ȅ`�|b���D쁰T����`W�?A���{�^��|�<��!4Ju��I���0HP�tMUZ;Ԫ��R�?�q�~���|�<Y����T�Q`a�Y
p�a��ʟ��'�2���?	��D {`�I���F�aX2E��:(@B��!;� �C�#V;�Z K�P�$�.�'���'��Dg��)�d��!l,ƃ'D� �B�Of���O���<�|:��ٖ�Q��#�C�P��AX2n+8(���|Y�i8g-Y�
{�ymH?���(+����C�]V=&��EB��+ܝd�@L
ϓ+2Y��� �Ȍ#��Z#�}
�K������u�'��$�5�	]�@ �Õ�m� �+9D�@�1��<Kq�+�;��B�7��g}r�D�~���7
H�Ѧ��8�X�	f����!���. ��ਃ�4Qr�1`�4�!�14����1�#E����D)0!�D[�.�9�c���:Y�e��,!�$�� X�mȡo�HӠ�H!�A�h�dP��܀b���˒	Tq ў����%�|T��w.�}\�M���Dz� D�並�̀!�Di��^7�(Q*�?D���`		�"�S�D�+~�c�B;D��7c�"/5ِŘ;,�h��U9D���w�432��J�<Dy�,9D��wE��4�*�yg��5C�����O��$�)�'z���2���}դ�ʗ΀^�b�R	�'Q\]�T�C;܁�g�	��2	�'1`��#A�0�d�pb%zzb�x�'�<ѣ��A�-���2%�X�w�X܃�'yH�PA�Y��(kT�Si㖕��':,� �Ξ/(}�=s��\�
5I+O^	j �'�rU���D�
ԙp�K�V�I
��� �l9RO�**䠡��o��*w\l�0"OH�`_,��:�q�\d��"O��u- 1؀`r�(E��1Y$"O@�����DW�I �.O�^f��F�'��D8�'Z��4%�"W�4�H�:Z��z�'��z�oG8A^���n �X�"�'J�H �
�0���!L#�,Xi�'�r���)��-j��)(N��0�'o0����R�Uޔ���+��.�C�'���J� ѧ w�d����v���ZQ?%rb�7!��p�c�(7�bl(�(7D���2C9d�E��� �LB��4D�|���֘yF���!I���(��@3D�,Q�GC�8+��\5,F,��n0D�����q�z�#3O7>D2�I-D���3C��~V\͚W-�6r�&|Q�J�Oڵ��)�'	��*P�	�g̼���G�m~��	�'��'�+���#e&�Y��'���x�(.@2��R�&*=�Y��'�<����!�@=!b	XxV�8�'��}���tt��#�XAR�I��'iz�f�K�JK 壠�\�4P��)O���c�'>�y@%�*&4[p�&c��'���!Q��kޢ�"3��5z�`��'LZ�J�뒭i���qB��<W��%��'���aE@��Hبec�bZ�N`H��'��A5�ݦ�N�h ΖB���c�=kXM��T�l�FK� �xē�"�De�x��vANy�Qcׇ�(��D�dy�܆�ERTqS�\�(��;P�Җe(�ȓC��y��V:;g�EKr���<Q���0g��+% <M1�Jq���|��l�ȓ���"Ȣmg��ZP$e�^F{�ǘ�����j�J޴~�j���?�q�"O���§��%t�`�Gy>| "OQ �+O�2�t�%(��g�Qx@"OT��F�ѡkJU锄�:�LY�"O��3�ŕ?<仗�AM��Y[�"O� ��<Mr�,�,B{2�C6�'.v�Z���S4%���Ao���8���� g.i�ȓy��T��8�(�"��ɰ�*(��yuTE	��ڙoN���`B7>� �ȓ3����0ʁ6'��H��5 Pl�ȓD�ҹ�cK�Kt��fЭ*#2Ԅ�%_.�Zɟ0:�t
�%�)"V&`�'�>C�(Il)��$�p�n\jV V.}�⥆���qx���}��'C�+g㴅��s��Ñ��8܊���l�'r��	��7Cv ���:�z�Ph˯L|���ȓ|g�Y�S��?HLѷ!,O����ɓ0R��	7�ʰ��۹P�x�PDGU&%'�B�I1UJ�� ��^D@�P�V�C�I%�|����>4p��[��, � C�i�� ��b�b� ��#I:V�B��W*��6C�b�$��L47�C�	�v5h�dL8}�)��	4���=Q�@�r�O~ep�OHgZ�@�������	�'+J,�d�K?=9$���#.]�~���'-\��A�W�C�&�g����'��m���ȕXڨ��č�l����'5�I�s�[��%8��9c�VD��'܀Ի�+�/p*��`1M"`�h��DD� Ex����l�L�H��۩0�2 ��0�C��*bB���Eԯ��5�v�U���C�)� XT+���&q.0��䘂B�Ɲ��"OHᨐ?�6Tr��̶�ƌA7"ODi!S �(�$!cabGpuxJ"O����]�$4,�3�vwDIqZ�,K��0�O\)#sB]!x����AC�jA �"O�Ma�f?��<�ċ�<��<y5"OB��� F��q�t-k �W"O`TL�(��� b|V���"O\ J�)�]�T���&8Tr����'��Qx�'�"iP$��%W�	0ē��z�S�'��q6��V+�]���<i��Q"�'Őy���̼T�t=�*��Pb",��'Č�1����ּj�L9��'*Jt�SF�p�q:��"G�9��'�lq0x���QW(��Ap*�����_�Q?�E&�IR���f��t�d+D�8M��W̶���e�W��L%D�(!��D[����E!
#�p Qg�!D��ׁQA�i�E�SѠĉ7� D���îA:Zz.��V�1Ȃ<Y��:D��{3�
��~@qAAl�H�	���OV����)�'*��� ��#q�z����>�
�'��<�E��L��h'`�ؼ��
�'&�l�o�5`�С��ܯ��$
�'w$XJ3�O�
�5�U�B�'\��#�'v�𱄁�>i�VtB�T1���B
�'k"�s�JV�u�S�D��ya)O���#�'�$IHaȋ&vR�a`4�B�?Xܽa�'J^u�RfN%�v���m (b7��
�'$��3`�$�
q�BB΄cT!Q
�'zVL��OCp�b�ֻV�m�	�'�-JU��0h6Xi�Q�O�G9���	�8�FD�z��͂� ��L�Lݟᜑ��~������\&3�.YX�$0�Ԙ�ȓ�6�����,`���́:k �Q��Nu��Q�N��	�D/�6	�L)�ȓt�V����u�N͋� ʆ9��I��U 8A��VOb���Η�ZM��F{�J����ݒ�"� 	����C����:+�"O��
Am�8��
F=,���J�"O�DZ1�M4!6
����_l{r4�"OȨ�qD&Gt Q��S��	��"O
�Zƅ]P/:�1��S�"�r"O��&��EYF$�#��>w��%�6�'�������[b��sʞ�/%���')ҩ7�U���~\�`!��i0 t�`��WL�������Ԏ�+9�f%�2͋=TP���ȓ7pp[���=ڶ<� OE��V��ȓN� �c"�4-�$��	W6��)���<�S��_8*��9KP�2#���'V�	�J���i0�����3�11I.��ȓ�؀y��18��9`'ߩ,꜇�Hnt�)��+�,�����$puFx�ȓFW��A��B!Z ���bMM'i���ȓR�8��$�UZ#���B,D�,����;�t�I�q�p�0�ĵt���#��yB䉻:n,��g/�DkpmS`�Q�&/�C��>s40�9���b��*4�C�	 #��BE\jk��z`��xzC�E��Ӊ�E�P����F�[�B��#]�l�"��P2$& t3�mF�"�=���K�O{pB��,�(��"�\�H�'
�	��f�u�)!e�K�^`��'b���I��-#�x)<��+��� r4Xe�RJj������*\Dp�&"O^L��iȻ|X�q��[���E"O�Թ�BC�,������%m���Z�'�ʩ2���S�U�P����%2���U5�,�����q����5���m�$���t�j"	R u �ы��Pm����V�d���O/_��y�bK�i��B�3(����Տ̍��h�'�o:�B�=7P��Ȑ�#a��!����ʓCqz���
�,l����)v�p� �C�c�B�^��%#�66���N11XB�I����T�`��TQ&_�SZ�B�Ʌ2�~��X?h)�i�p ]5H�B��8zpm␀��p��	3"�~���ތ]r�D�<Xv��Q�B�H��uB��':!��]�S�\Q��ҹGf���o�3 !��Ƭb�@���Z�,
����E!��^9gc(P��!Y�c��u�!�DQ�?U�(2Lp	F��,!��ΌP�:8�1AX-}*�z��X
"�ў�I��+�'o�����*�!y�	ǥ3P1��^a�\-��d��%�yHLRӮ�`�<�'�*o����g�y$
��C��B�<��H-��� IS��E�<���ыFO`�4�V	2��%d�D�<���TD�c ��U�\X�l�ǟ4��.�S�O�V��k��0��,�d�Úa'Ԕ�7"On��ud��l_t!���Q�˲"Of�� (���)cmM�-����T"Oj�@�=;z����S�`�f9qV"O����&؛s�N#�܊OU�d���E�饆X�uyh���O��'	�'�8�';��˟���D�Y*.="Li4�?���3l;D��sJM�Z�41RС��;ąHP�9D�ʄ��	 �]`f�V�{���S+3D��x�o(tX��t���Kw�yP��0D����,�*�0Sr�
�T�v��2m)D��	e��"&� p(
�T3V�i��"�	�Nr�"<��~,�b�Ƿft�`Rr�B�M��L��"O�Ҁ��70Bq8�H�N[�e�5"O�P��j^$	��HCҢ0Ue�'"OL����تS�1'ӆ,���"O�Z�ő�V�xd#Ւ<]�"O�̀��W�Y�L��֠�u��
����OL�}����}��?� v�؝8j���ȓ0����fސ$ �$Q%MŅȓ'�RT��n�r�8���}"�p��(�	����;	yF��j�V�����@N�jcƑs�r�j�m��L4HՄȓ�܀��˅'����؄-���ɷ7�N��d��MH ��@	=�z�4��!n !�d	 g���BL[;���*��B!��4�X�����YC��0|�!�D�
����3i�%L���BE3I�!�dC(o�	4�X�LƑRC�@2,��{2�Ö��ɣj�|� A�]3�$
3�!X�FC�	�|�� �	]=R���!�Y�]�C�	�V�&`JE���0ɀ����3��B�	�%x�J� �*)�l��G��~�vB��A���pmm��Q0sB^h�fB䉸R���83ɗ$)|m����P���Ĉ�e �S�)I�>7*�!3�����p�S���!��D�І#��-�,p��+<!�#��)�e��T�f�{V���Py
� ȱ��Jyz�h1T�Y6`j~��5"O���!��-R����q��0%�ʩ��"Op�9GÆ8Ҍ=E�@=c��W�H%�O4�}�ke���A%�e-h��Wi��ȓ5	�1�ʀ+]�D#��=|v��v�b��#`�3b�:����4�~B�	�H�`AEQm{ܼ�wES/��B��8?6��q�<YD��'C�B�o�X�I�
�T�R<�a��;��dJ$;W�~�خ-�"M 2@�9^G�-�ЯL�ybN��DX�
2�$I����_��y��5�ĹHP��-f~U�b�,�y"�R��Y� �d�!!�)��{�'��e��B�k���P'�5Y�`��'��Tzg�@�Έ
���>3R(B�'�P�C&��U y�F/:���(�'<"xS�F9�Zu��%�V�-+�',� \��fq�N�JaT�p�'Q��+����P5�ըF2CP|i�'���C��ܬC�����^2�@�+O���O�O�6��A�4��N��bU���v+�B�	���� q��9b�(@4�S7_�lnh�ɭi1�rm��UoxT���O�-R���)㖟� �'�¥�L���<Q�kÃ5����T�L)v]z�Br픇{i�@��O���O�tz��>�6���ʖ!�5zU���#c�t�f�J�ծ��OΠ���h��>8���2v��0U82%b�-�����>aT�>���Z�Y�4�T�P�jiD�ۢ>�t�1��?)��Vy�����?����#Mf@ ���d}`}�c(�� �t�;}2g-}Ҭڷ���MsG�?I�*�k��=T٨��c��my�����	9�ȟ�){Q�)b�6mz�NF9M�@�I?�iT�T>�I;�6�����TG��{2�"׈Q�>]"�̟�����Zg��$<%�>����qEE��*X�p�^őS��OڅH�'�~���O�s���3����u�Ш ��6̄�b�F��O������pYU��3;,��eo�t�B9�ȓ[������.m����?|S�o�x�����<)��?)DՇiJ�EJ@AՎ!���E#ݛf�'rT�|讟
�O�iQ��Z�o&�e�w%/*8���M<�*O��O��:�"S�ԩm����?D�dI'"Op���	R�G��5�FJш!�2"O��t�S���Zn��/�<q�"O�`B�J;,k(yc'�8�,+"ON�ꑨmVe�U�!h���˵"O&͂Ƣ�|��	T�՜4=�"O�+�.J�
�8�p��x�̈e"O��wLΥ`&)��*����0"O�:E���C�F<�g׍g�v+D"O�4SԆ�:Y/�Ty���.D�@h'"O���0n\	m&�\��ًw 0��@"O�I���@�<�����<<(<E���f���y,ġ�RA�c�5pl���ߛ9�j�3��ѣvȄq��ͣz_�|K$�1�0mʷ OIN�l
7cŬr&���3�ܹB$0'�½F'~����+1����+Μf8|���h��Am���ʜ�FB,�@���̀3�4�BW\�(+���r�I�X��}YW�8�йZ#�>+�C�I7\��*��<6�!עI0�hC�	�SEb�����	%����(qGBC�	�2�� t��l<��˂B�&Y�C�	%I��%@��8����ᎂd��B䉒 ����k˲G����,X�C�B�
|A4��t��uC�Q��B�	� ��:��G��+�fڀr)�B�6B>���c���e�&�!]�dB䉊l@A)"Ę�A�GX�#�B��{����c���dh�	��B�I5h|B@�眤5�n�+�枣0%@C�In�LA�� �j�G[�)m�C�)� XMh��R�>`��"' <�H�"O2���#�
9ȑ�2*̍4j�K�"O pz��L�
�h$���\mi�E"O��y�(@�l�8x���;�ظ�"O�pf$^'4���H�iЃZC�qC"Ou�4�B�n�����;4:��I�"O��M	'���4K'��P�"O����Փ%BXIC�J�(t�YX4"Oћ�L��/b:���eZ�X(��"O�d0s�Ԭ��cMz��\�t"O���w:Y�5��H�~0��'=����E��Z���Ev�a��'r�ȋ��S}�<�a*ݘ?��43�'�\�X�)��,3¤��s59�'�8�C@R�>���`�12� !�'��ؐ��]��IJѥ�:/��P�'C �z# ����A��,! M
�':|�cA�Ōi��3�iHq�:���'|�0Y�^*sIʱ�ũ�b��A
�'e-(�c���
�g������	�'Ӹ�Z��N�Cv�)4e�)>�X���'!.��V)� L؂鈤*���'��T��+º7�0Qq�f�U��Y
�'0��!4Η�y%F�����ܼP
�'b��Ι�L��KgS8%O� ��'����OZ����x6k$�*�:�'n�yb�O+7�R��r�x�'�ʸ㓨��]�\%Y��^_ȉ��'�"(��_
��ɺ�Z�98D��'&<@�C.�1�v͊��)���c�'x*��׏��P��Z$M۟C��p�'C�Ӷ�·8�L�V曦A/D1�'w�,B��O�0T�QGW�4�ʨ��'S|lZ�L�Y"-�p+L�/P�d��'��$n���H�iQ)~�p�'j(r�ɧG2-���w%zE��'nPa�N�ؑ;4C�kj����'��܊���|���;kb��0�'�r=����t�5��2^�,P+�'�J�aw	7WV"���+�=R|6��'B����� =�8m�R���U~�{�']6��g!^V�!�"f�M�"|��'�(d��Jőn��uF�!D'���'M��'�R�D^^��tK�=j���'5Mq�� *q|b��4��$-���'j��0�%�
���蒹*fx�
�']$L���X�Z ;�
V
1���
�'��� ��v�TbҊ9(��hK�'ǚH�C�_!r� �!a쑀0dX�'M�x[bՅ`D��( �_�l�H�
�'Ax!Y�L��>��-�T�tb���'�F���B�:�EpÌ�)i�H
�'�`���M�T>MKc�"7��a��'[��%����dpRh8!�5q�'�^0k���U�`+"P�f���'�� qao��|���u�פ^}�	��'��c�Mˬ[ ��i��\�����'H�9��'�/J��P�4aZ2SƮ��
�'tJ� bUG�����%J�R��
�'�j�iRǛ�E�ܔ;�cU�F��Qh
�'al]xU ȉ9��C"/ڡDq��
�'���#��ٚcŞ-!��O�E�����'�.)ġ�7��P��'U�z8(�'=
4�@��*y�,�O�4Me���� �I�
��tK �*� ɅpZ|��"O���B��g��M)g [��P�P"OF,;c�D�!Q"Q�v���j'"OЕ f���yπZ�B�W�F	T"O�t�Ӈ�xrU��'�){H��C"O -�4f E60H��)A.��"Op��4T�/��0�@��,�(A�d"O����N��Z` �ӳ"O!�W�J���g��P͙�"OFY�T�}�d\�%�%u`y�5"O����`\�#Ԥ.az���"O������:��X�%,7��mj�"O
��7G̸G>�� VO����"O:��V�����E�1�P���"Of�%	�Cn"<�W��pb���"O��e��OJ0��$LN��yv"Od���^?���P �b8�l�`"O��A3�#W�X�r�U�8��#"O�ef�M)(DQ��*		sE"O�i�$OCg��-(%��[��"O޸��S� ���O��J��4[�"OXE���,�
��@N
g*}*S"O��R�$[(L�T0�f�ڝ9F�c"OxD0§��n`�A:$��|�`"O�m K�g'P�e��2�|d�"OB���NQ�(��ǅ�Jg���4"O����f�%�l���G&bSp�T"O.��JE=�P��ʕ�\7�"O�!��A+N�$ ���*1b�"O@Q�ªQ/@=�!��h�.��+�"O�Po/X�@zV
H	��,�"OVq�)Eޜ�P@�ϊ"&�q��"O0\�D�	\JIش�\���q"Ot �b�%  ��GǞ0�F��"O�Ibc��g�X=釨�%i����"OƠqgc�(7�и�G�L�����"O���`D����A�/��(�.� �"O��1.V7��j���;f�≺&"OܩRL�|�D�X���/兖I�!��Ƨ}H����ϾX�F�K�k�5w�!��Z�C��]P��D*=�J�! ꊗX�!�=O�Q�AT�o ,��K��!򤈯I܊��娕�|z#U,t�!�M�%�(-�r��)lYy�mY�=�!��
3^��+���B���fĆ,�!�$J�w~�4�T�<*t�rb㜺w9!�� �1�Fi��g��,�!��y�@X�d�޻�̰���� ]�!�ğ�x���-�-0@ ����!��Q�%g`4���	�{����.ԗJ!���J�L!6�Wh.ġSKN	T9!�u�,3M��@ �ݓ��ް�!��W�X;�52v(��pD�9O�F�!�U1���3 �X��]���2h!��.i�b9X#I�b��ЫG�`!�$��w��t��b�Ttr �$4E!�Ē�9Wn	���@��e	��Pc!���`��3���� ��P�qO!���x�Fuа���-0�%�� �d'!�$VjJ�d�⚖#vb�� �[�!�$��	���%ͅRub����!�!��  �i�Ξ%]x��-Y�A!�d ?�bxÏ��gH�	;�F�%iC!� H"�r�'"i�\,�ĦЀp�!�� �)�W�ơt�Z� CB�'��	�5"O��p�}�z����{B"E�"Od隄%K�	gZ��P�+>0
�"OD��e���=ZE�ِ~�P�*�"O�z!�I,^y�%���ޥ|C:��"O�Pp橗&x_l,s#b�x<���S"O
��]9����7!�z:���"O4QcSȔΨ�;�	�"Ap�"O��SG�:�����S	p�͡6"O@��Ν�<*\9q��b��i3"O�d�w�N��ͻЩ���`�j�"O�u�2�W D��c$i�R0�! "OD����̬�4Ej1	Е`���6"OZ]�R)ֶBL@�U�\
zA$i9�"O�	ёѶ>�&E
��01y��"O�|	&AW;1rQ��蛪9���B"O\��͍�2)��:��"U�b9 �"Ox�`�!�	Y����j�6�J�A�"O9뤩�IP�\���[7J��1k�"Oz	j6<0Q�I�3l�	�0"O�)AI`��M��C�+����"O4m8���'��0����0x�j!"O�� �K�yH�a�(�.0P"O�|qHRrr�č��[�*tk"OZA+��phYz���(���"OP� OA�2�����iN"Zr a�"Op��S�Љm�$�����2�b"O�|�s�Yj�l���!�'ذxQ"Oi�2#�WP�x�B��t�\C�"Ol� b�̼[$d�a�Y�n�X�1�"O� ��f�Rl8�8_�|���"OP�	�1C&�0�l�u�^4{R"O�9)gl�"!���r�y�H�b�"Oԁ����4��i���K�Ql)�r"O�l������b�]`r�e0%"O���Wo�!r�Lٹ�P�yc���W"O��:g+U=\1�͓q��75�`�R"OX��3<听��T��0�q"O��K3�l��D��[�<,H�#�"O��ٴF�4n%�� �o%M����"O�H��+�6�䜈���"b����g"O<�+r�.9u����g�����"OL�P�`������˞x��%"Ou��H�)o���G*S6*y�,��"O���m�3T��+B�R	�0x�"OLe�ׅ�>}A��_�H��"O`sD��?"�q� ���V��\�&"OB�KQ��>�~d�t�K�eV�ezg"Ob��Uѻj��{�#�^Fʸ�"O�� ƭl Z�B�?B���"O4�a�-M�]*��T�3R!8���"O�T9S�=I&N|��@؂g���"OJ��Q&�<�q
èW\0��"O�ݠq�1�Y���_G���t"O�2�E�;ֆ�à��$[��"Od��g�e��B�h�'?l$���"O}��<e�P]��'Y�n �䛼e����7�%�`)b��-%�'kfy��N�;:8�Ҡ*Kmw�0��'�2�"R"��_U�������<Q+�'iА��*�N�15��&���'��a���N�&FY�e?X�Vx�'%Ri��fp�c�A�P�z��'}2�#fa��vx�0b3���B>l �'�����U�"
ȱ�c^���J��� P�H�*݌W��$�ْ/����e"O m�s�Y_uDЪ`ކ�4���"O�z��ەm�<�8�M�Z���"O��"�X#��W$7D	� "Of ;3o�6v4X'%�aQ��"OPTQw.I G]�2�$/nW�<�4"O�Ec�(x��}ң;Ul&H��"O2s��%)��d��Q�c4p8@"O� ��P�<���D�C�A�"O�ݰR�%���$� �lz��Q"O���rR���,֝+;��#�"Ob�@7���+K6�;6fz+@0�#"O�Dp����増1\'�� "O�� �iT�i�
����F�-s�"O��JC���`!>�'@#_��"O��hw�ʟ'B-+�6]t��"OЭS��B�z�y e"O+5�: ��"O>EQ&�U!R&��T��,����"O�1R���61I���Ơ�t���P"O`уQ��+���FM�U�|���"O`	��/61P����_WpU�V"O��{c�%&C�=#́?{Rdx�"O:��O����$S�%�*�Ѵ"Od������H�̟-n�B�p�"O�q�"�Zkh��bC�*X����"O�����sE2M��۬?�6��"O.�)��қO?�0��Ñ1�֐@�"ObQ@�6y6M��l_:�d�H"O�{�m�%Z	��؅�s/.�h�"O�)%�hm�����%#X� �"O�-�2h[�nb�ȥBR�a
��+a"O>��@.��z�n}3�!ФgR�
�"O�}(�M���ATq���t"O��9`�0 ^��QS�K�C��\
#"Oh=i�D
 �jH�4N�:6��t�S"Ol���bV'<�L���#G�*$�"Oz����(E�,���I+7�Fp��"OT�q��_2PNi�㬎�J��l��"O�YY2�/H���k0)��y�l�c"O��)�N�*<����J�<a��iS"O�������<�0�X�5*����"Ol��f������Ve�-Z5�"Of̃��@:01^��5%7R�� �"O��3�Şd,���g!ԝx}���"O����B�$CnH��I�!c���"Oj�Z� �1F�xų���7 I�!�"OV#Vo� ��ܹ��ŲHL�`y�"O2e�_�F��0sL_�O���u"OJ9��*%|̸�24�N�\����t"O��T%���i�S�S�1����"O>���M�D �*���GZZU"O�iHυ�q�Ѕ��L���"OشZÁ���RԎ�:��|qr"O�� ա7B4����_�
�ʴ"OD�j��G
j�=*V�q
t��)D�ةgOT}^��3��;o&�pQK7D�@z�)�=�Ff��n/F���"3D����P'8���("�0G-X`(��;D����� �i)�З�N��IP�+-D���C�{"��X�
N�06����&D��	w�[)<TM!@G?f�����j!D�tc�HD?;B8X��虽F��F!D�HS�L/B���C���q�.D�l�#�8d�l���R�{�LC�i,D�� N�{L�;@�°�Y�XAs"OT�j��R,������.�I٢"O�l�A�D-
5��2�NΒ"6��Y�"O��+�ƙ|�@=�t͋�
��?�yb�����x�,48� ̛����y�D�v��s���g�J�;��4�yB�Ƚ#8�a� L�`�ĕ���L!�$�"G"~D�ԩ��S4���«_�!��m�e;��S5��4�ӭܮd#!�deB�гP�ߋ	����U��6&�!��]��,=:�f��[�~]��mT�t!�dC=2݋�N�'�e"rbׇ|�!�����s�*07�d��Xu�!��_6:\��3Ҫ�7".�t	CDܐ5^!�DZaj�BVU#�4h�U�X�4m!�D�(>}.|[Ӡ��id�#�N?!��.+hQ+p	��
e#5��!K7!�䖛l��Y�b,Ź��I��ϗ�9�!�d�G٬�cބ9�
�ۀ)��!�$� F���B�k���`�5<�!��:)�`�P�:ZXa��9u*!�P#0z���xrX�Ju�X�,!�Dλq~�V�{�4��O�/!�J�EݞM �c���0!�oʱ�!�D)E�d�%dB�l�T8RANJ�h�!��I����;�8��7���n�!�d!%Z��e�����>Ct!�d�)�"�+�>,&�'�^%.!��U�7
	� ��t���7⎷a!�$J�`����T&��Z�f�iE��!�S.K�����gǾq�c�ʎRT!��>6�R��-;za!�E֧�!�dڑMP�	��<>�����4_!��ӍC12@j�^�J��u�'�<A!���9k,�!�R�4*�iD�"DN!���,X�Y��Y&< ��2��;�!�JF��d*����Y\#s�Ͼ�!�D�n> ��I)Mx����)�$f*!��[�P�!���m0	��!�dӈBӢ5��� /�Lв1/�K�!�d�+�l<ђ�����z%��!M
!�$ˌ�X�� L�<�"ܢ�$[:U!���U�ti3f[�<"��� Pa!�֮K�F�Ȁ��l��D�'d-N]!�$��!:vq�6(|�X�1�++#E!�$��j����Ĝeגܚ��Q��!��1v(壴��}�
�uN�C�!���qc��k䇅�**$����4�!�d4S
�<*"ۀ:b!��j]+U�!��_@R��,\��Z3T�q[!�=Od��2/UCg�Qg'Ũs�!�"qr] &#ѦNU�<xd�e!�䁗\�>Pj���0F��ݺ���]!�d��q~�j�.��-��}��/��v!�D?�8%)p� I�H�ˢ(T�s�!�D�9k���C�нW
D	�'퐁"�!�$�2L|2����;�B��V�$�!�ʃ^3�Mi7H��8鈱�_1~�!�$�
eZщ`F�B��%����3@!�\$;ڒ�Ѵ(א���P�ۍ"�!�D��gi��b�c	�4�p��1����!�ӝ~T�4��*W�D��"ؐ!!�6gp�q85"�/���G:MV!򄍧\/�탑B��X��P�D�!�� �����k}�P7�[��T�"O�%����8�:�1�	ק_�>�)�"O������%i"�̪pC/d���"Ov�J�e�.	�(�BIBL*�0"OȤ�Q��*N�"��§�_Hb�"O�ܢ��H"Tlfd�%��q�zQʒ"Ol��d�(`^�����;�"O� ����+�
 �"%X@2��"Oi��ڬ=��p�eM)7w$m�"O��	��=s0�T��ݘ]�}�"O(���D�F��)�L="YȠ�"O�b���Z2Ç'�1d�F���"O�� FƟ(1�����ߩ+��|�3"OP���G�?(�>l����\".k�"O0p�D�>b�(�K�<n,�!�"O�����
<Z@�Ʉ�/X9""O!��h��/d��aGh݃�J|��"O6��A��
�й��/�h|6H�G"O�aA�G3��q�r�Ģ]��[�"O, ;��E�|���B�
�VAڔ�6"OB�!2��,��Qf�-��R� D��9+�	"�.	�	�b�"(13.D��׫X1.��,S� �e%\�Ê+D����Ձ]��R���V*� ��-D�l��΁���-I�`�/V(���-D���B� 6p!;��'WUB<#3g9D�|)��@����� ���
��bG4D�t�䒺q�$���6Zu�`�� D���EZ�M}��3�/ˀA����S$0D�T`Bc\�/��d2n�3Rr�@׉<D���6#�D���d\S^Q�O<D�d����,�i�@L��5�ѩ:D��K�K>��e��E� @$<3�C3D��뙑W+P8�'%"�p���<D�h�G! k�<A�fV�X���d:D�:�D��H������ms��;D����'kv��0k��H��9� -D���w�S�B���f��!� 5�P�.D��!q,Z�H>ܻ7ϧh�\Y
TK,D�y`�  r�s]Jf�S5D](IH!�2�<,��@ßM��]Q��T!�<�J��郉I41����X!�:K�4U�6g���'"���!�$O�5;�@�3�.�:VΞ�z7!�Ĝ�9����ꁮ�F "��H� +!��;.j��@ օvҠHs@��5!�DU;��͖@�Z�rv�.M,!��@0j�(92��650�5�'L��N$!�DD���}�c��0, t���_!���qN8��D�+�����^�!��!zqkP,I
�<;��+?�!��[\��
é �c��dˀ�0\�!��[�)�֑�b��r���3Á9�!��S�,d��O�w|t��� d�!�d����BڄZ]�m�W͏*!�d�-R��r�˃=�T���L	�<"!�č$il6��g�G�	�����67
!�dݲ.�QS����A�F�I�0!�D�4h����B�W
dT&u��fٝ�!�$��n���'��T���\-!�$�P
|qg�Y_B�`#BqO0 cʆ�.�l�S�(�����|��U����f���hѩA�y�o�,�
ȉ���^�P���C��y�fH�L$N-� h�.&"�X��Ǎ�y
� (p��V�(Op`06?dI�"OZܘ���?yBP{e��5B3���"O�@�c���v�-*���F���"�"O��BBmªa3ʩ(��̸N	�đ�"O�p��h϶:b��1�]���`"O(Ihu�^�z�� �.@;6����"OЭ!V G�=��D0�BY�M�FL�4"O�,��[�q������3�nh�"Ov�p䪐�WF����n���8�"O�\�U��*���DT3��	B"OjM��BH=� �a2�G�_���ɱ"O�!_&O%�7�ؿK�B��7D��'W�au6�3��W(r�4I��;D���q0􄺃D:Ehҹ��6D��)�ش!�\4Z����<�d�z�	3D�\25Jɴv�xJ��:wf���)<D�ܡ�C¤�d�aŠ0�l�SE8D�X�A�L��eɕ��,�i��*D�y�Ζ2���B��"`<+��(D�<7�]&=&l"E �rM�D%$D���
çc��*���=g�V��
8D����ᕫq�2��ѣ��
�J?z�!�dI�v����M
B���3R�ܸ�!�M��AC�"I>Ա pgP�~!�B�H��p0�٭��եT,!y!�dԡXv�ث���E�p8����=!��J�,l:q�����
���j�!�M�#B����e�D�rAҀ���!��Ė��={7Ή?j�LQt�8:p!���<�̕x�'(~���!��&iP!�dZ�=���Be�H��J���@G!�ڭD����ǤB�7�H Jd+!��Z�:�r c������ƨ�+a!�F�)��Cʓ|���&� !򤒏 ��Lb7,e���"��#!�I�P]�� �X7C�B<xG�1!�!�Ν>���'>y1���Q�U�,�!��T���Eѧ%)NB��E� �!�S�-��� ӈ�_"\i���.����3*��`G�	0e��o�+Xv���gM��HD:�E�4��(Sz�ȓ84|u��>� ,"G���Tȑ�ȓ���	#��2V̱��T:
4�\����E�ю_(p�TX�d��;~+BU��Cj�q���{�fYa�8C.�Ʉ�=���оB��
�f^�y@�������o]Vl4�'���-+�x�ȓs�LE��%Hd  �NBK��0�ȓW��CQ偋lej@�<߼�ȓVN@�L���@u��F��P�ȓ^
F1
�B�4;.b݂��x�t���m30�`\!��sƮ�ug:�a�<D�0q��U�,����1�H³	9D���d�g��A�%(� l��5D�0I"�E"��5�OS6}��y{�B>D�pBM��z�(����F�*~q�)>D���a:|k��KI�F�h���;D�Hrq�J�-���1`�X$R���*:D��;�L�
f�f���G>H	!h,D���TC�0a�1,�9ٰ}��/D��uCI	;��q�c��~�p� �:D��P旙�l��lK1o���Xrg6D��*TbB�p�a/
�D.R�*Q�2D� ����0]��
$�H=s4y:�i0D��  �X �Ӡ��C6&���d�P"O���!N��UBV�ڎ}X���Q"O�CӪ�'=u>��M@+��LІ"O�x�WnΖ.A�u
����C.��"O��h��E�xwj�q��̒i�$[�"O�(�A��.�*�b̪"R��4"O�I[q`�$pw�)0��N�k8�X6"Om�V�?UH���M���JC"Oxa��@�E8w�&5Y
@15"O���h��1ƀ�ҁ��uH^Y/�!�DM �M��ʉ^X��B�9WL!�ą�i�, �t��<��-���T!1�!�dL=Jì��`
M?���c���!�$�N)��#���.E#ph	�R�!�S�@j���d�ܣq<G	U�!�ǜr���q���f�5���6p�!��P?���q��^�Ɲb`�M!�DQ7M%DԠ�\�L�6#A�!��1N� �q(��j�6U���Q&X8!�ؚ[6u���G�I����0��RK!�d� Ov�80AP�V��cv'ف:$!��O�G�VP�3�á`0��� Y�!��<͜�!��?,T�� � _�!�dܛ3��d�AW�(Ʋ�)E�h3!��A��ّ�F��X���A51!�d;WjL0�W� �E��]�c'�*e!�D0��Z��/S��(�wF¥%�!�,��bo�znt���F.Z�!���Z�pՃ�o�2ET����S!Dq!�D(M|U� 瓡G�|)��/Y!��p��'/��A�(�H�<cp(q
�'�*��$��3P24�Fi��h!ԕ��'0�v�Q��= �%	,(��4@�"O�
�C�ji\t���`�d��"O��y���<b�@�q���3�<�5"O�	#�ćr5J��㜠l|�8`"O�mr�A�
^�̘�qLP�|���%"ON�2��9|���C%Ѹ����"OЫD���6ohA���Y� p��"O^�ڔ̛#����O��a"O�+�n���U�Q�}�f8�"OD ����B5�5y�ם=����"O�|�QOZ@��Y{�j�7Ƹp��"OHL�V��
$��I��&��"OFUaU(5��|�U�9v��9�"O&1�W
'��q�6���"O�t�e T�-�Z`�+�~x#"O�YB���nRNѨ�D�<4�`@��"O`���K�l�V%�EH(,��Xp"O��)��R?
_��I��\$Y*"O��x�%��ƹ�I;h��"OR�jǨY�3�$�SC-�-\���d"OX��"F�.4�n��-
3(�Rh���'�ў,B`�O�h<X�����5���rN4D��jB. ��
x��.s�i��K4D�p@R���'pL�@�aİKx��Z�4D�D0�X�X�22#��aq��QO0D�P�DD�0E�5��fԾz�,���(D�	�-\r�8��Z
��*BE
�M!�dW>���K���[�.)@Q��-FA!򤟷�"��dM��Y�xT���I8�!��Ux�X`Cq����4�̔8�!��Ty\6Ar̀5I� �}�!�䎬���p��&��ئ�>�!�� ʕ�4�o�^=��nU�1wb��F"O�}{�A^(d���Í�it�b"O���E�}xN@	�ne:�
�"OD�d��w�h< 2kF�nX����"O��jB�Po"^��d��IC����"O
�)b�[�"�R��QbU.K2<	Q�"O0�J�I2 ���a �<*f�`"O"q����\���ؕ�
*��8�"O�8��-����;@��.o��!��"O�h��CX���� Z_�HD���
e�<���ѯuO�y��D��|�a ��F�<��I#���k�'��:�z����|�<���x����1��bQȬ(��y�<�'o�&X��Xc.ĚD�P��(�p�<1ѫ��8	0�r 埛�f�P��a�<��lS)`��i!V'��$`��H�<�d�/f�)�#@�.R}+���F�<�Q��ED�u���-0�:}CF�HY�<���7H�D�A2�yg)�k�<	�dJ�r�x�1!E@�T�H�2FW]�<	�
֖o�xQi �C�5����<�#�ּ7���Bn�fL�$�~�<�)����k��	D(1BR[}�<	�,=0;Z�P%����e���H}�<�b�]��H�ɓ�W?��aK�d�<9��@C 8������6���i�<A�F�hǾݨ�$Q4R9J�F�h�<�G��5n:6���h���ご�y"-(NH��ab�	`&����Ƣ�y�5��Y�M�VS4��〙��y2i��-�����B�@�1ևV�yҬ�/�J�0E�8b�Q�l���yJh%��2�W�*��L�0J�i��B�Ij�@;"I��M�<A�/��>B��(����0�2Q���c o_�B�>� 4z�HL#=0h}�r�S'#��B�ɛ|���A�@$�w�,b�B�]?�H򳋁�j�X����[�z �B�	/q��r�*Шz�0���c٣'|B��C�^ �%��)��E�,��B�	,.�ތ��d(~QS�@� \�LB��!*���bWI.x�B���/+0>B�	���|y�C1u�P�Sl��I[�C�I1Q ����MT�������z�|B�B�r�h`CJd2䣋�VnB�ɼʶI�`ɂA��	b�S�[�RB��0B������83R�J!���VB�	{��aHD5O#��ȅ��2G?*B�	s~H����ni���SF�1P�C�I3�ޭ� /��NI�5� ��tTB�I	d6J��A�)\-\� 2n�g�^C�	�\_�M�UF�}*B�B�,�>r�,C�ɢm�]P�����f�
8*C�	�4���FF�
-6Mr�N�=bC�	�9�((��Y!6dAr��PC� k����	�8q����Q�C'�C�	�S��u��`�5��Y��\�&2C�̾�P�Fn�UYr�Z1	/TC�I6K:)y�˶N<���,\	N&C�	R��a���H1]ɦ�K��'F��B�	�1�����i� :���y!.X�7��B�I�Y�pA@0��+lThxkvK��4��B�ɈE��T;�/Z�9M,�,�%h:rB�ɧf88�Ʈ�9g{��:Gn�>9&C�)� �`�VAP:��������A�W"O�{�+ITT�[�c
EHY�@"Oz�q��60l��&�z(�l�c"OZ�@�����m�����=(l�"Or4����������څ'��m�P"Oڔ�%��y���j���	N���R�"Od��2�-	��ȷn8g���"T"O���P�N!E���LA�r�T���"O���F��$�|H"iL%ޒ�R"O�EH���0_����W�x���"O8��⋆�����Œ�%��U"O<$i��x5�4%S}��p9�"O��hF����j�b�1y���i"OF0�r���`�в��T�e���U"O\�� �ŷ�2��j��A�٨�"O  �T�Q=@}zĩ�H��>DY�"O��1��G�3`$ߦ�dH[B"Oz��GiM*@�#��8���"O��n>�~��P@]�|� 43�"O0ĒQ�Ы� 3�M���r"Oȍ���Օu^��Ռ-܆� �"O�P��n��J"�9P�]�qk3"O~��5(��P�ZI;!*�.^��l*q"O`Xbc���D�9�	S�b�8��"O
l�&L��:���%*�EP "O������G��S�a�RB�� "O�$[Ch�9_��(b��)�L��"OF
wi��F���d�P�8�ʠ�"O)rT��{�����v��z@"O�̒R�.8:ȥAT&��z�r�"Oh�8������Ő��P��9y"OH �"*�t�F�#UB�!C��aC"OH���]�A��Q��a��P��0�"O�Ap��<=1I������2"O���7�ؐ$_(�S�b�N����4"O^��v�؟�<rq"�)w�X���"Op	jt�ς;��	*S�Af�"Ś�"O��X���?=x�a�H_�ώ���"Od=Z��0�|��gS5��)CD"O��3�ߡwҴ-���@�=���zS"OԹA EׄU�J1K�dƀ���Ò"O����h)���lB� ���"O�X�̚�;`��:t��C���5"O�ihE�HRƤ��"V��e�3"O���6싊&1V𣂍emf�"O4`c�k�����gk��ځ"OZ�bea;6����$#P$��"ON�u�םiO�9zՆ�,ML���"OP����'vbMإ��7���"O
��ac��]�H=k�D[u�B�"O��*sE~��#�c>�1S�Zc�<Y�a���x�83��	)�"�u�s�<р�Իd3��h�BIH(�xva�G�<D쒅%���� ̅:o�ːO�k�<I#
6o���C]�u:��d�<��L��@��D�ٿ?�@�3�`�<)��C�a|�ey2i]�q�`)��AZ�<I�ęs���m����p%_�<�P%Ɲ-��%'�bq�uGZ�<��k�?sF>鰥%� C]���ADR�<��E4G|�����8hk���T�<i��_���剌1���� @[�<�����&�@�^�L?Tس��*T�������0\V���o<U���	*D�� � A�~^�L�^1j���"OԽ+�ؠB � ���Ww�ŀq"O��"@ޭ$��3ģ@�wy�e[u"Ol��#�a�Ҡ��i�3[��Rt"O΍�r�]�6�H5x��_-@H��Q"OF�p�YP�Z�ʘ��YA"O��i��3Q(y�Х��U �X�"O�0c� ���h��J�����Rq"O����Pu�܀����ZyJtR�"O����j�.*@I�Ӂ((��Z"O�q;@�
�9C�]J�BN8,2��"OZ�!t�<�^!i$Ir��zf"O� ��'�MN��	j&��1ʇ"On@P�I�5��*.R8F�6�V"O� $�ўx">HT�� &�)"O"%���N�M����K�6u��"OI�½��ջ�k�/Y�܉�`"O�!/M��Xr2�̥#XN��"O�ݲ�e���X�	U�@�K\Y�"O��!㉝P�lʐ�T�7B �r"O��R&�9P<�d	rh��"OJ��2� �aM(�V���D�U��"O��;L5ȁ���1@Q��H"Ox���kƷX��eag��{3����"O�h�F��^o4��M7qNLr�"OLZ�E4X�Flh�E�hPq�@"OD�+�L�lNf-IF��K��"O��#�ބN5�TȲ���X�;�"O
! saM|��i�7��|W"O�$;W��(?�H����Z�V�hb&"O���&���M��<�t
�y�dl+S"O���ѥ��?Ğ1�ܝ���F"ObD����-W$Y��GO�H��TkR"O>�����:Qx4L��M�"����E"O�h��H�'B��<�I�/���P"Oʰ`1͈��M�h,�⸈D"O�4iF)�'��T��'M�}�ĵ��"O8�8ĉX4A	��V��*
m"�Qc"O8R2�\8}�\�!�	"|���"O.���-��2!'�@AP%3�"O�Kt�D�Fq�]H2h�V�,$��"O���ǣV�b�b} �)��It"Oڹ�b@G/�h|���8j|X�Hs"O���2��R-� q���;He��8"OyC�X
32~ع��<.V��	�"O�@��]�\����F,��I&���"ORt�B�Z�:w���U��)z4�"OpT���.t]���mO�0� ��'�p"�,��Of.�6L�Ri�K�'�V�a�A�K@P(�eד_�j��'������{���*���I
�Q��'����o��q:DH��A۰;E֘k
�'��J����peS��W!8�|���'��% ��ݷ�����ˉ7��
	�'����? �0Kci��-0��Z�'��(��J.0�J�`\pn�uX�'%I���Vs:��k��աbN�!�'_�I�
��E�X�0���'Z$�x;�'yR���ב~ʴ����G�}mN�k�'�jm)�_�S� {�j��M�P��	�'�"�I�ΰ0!��>(�#�'L����F%Pq\��Q�B�`-����'��i)�&���Q"D�X�4�p�'��*cB���8�"�1W�t���� |)�r�[5~2 ��tB�3�Ly�"OpciW+�����Qpת�{�"Ot�˵/
�/� t�&��71�Υ�0"O��㎐�M�p�{v�Ƽz�E8�"O�m�aF�-���@��F+}��u�r"O���p�X�nX���*G��ٵ"O|��AT r�,��өd��2�"Oj���8`�~	��iZ�X2#C"O��  1�h���h.Zwn4K�"O>(!��-1���!���>�D��"O~|x�l�6��$��ˉN���"O��GD9pqVp��e��R�RG"ObH ��(,Zy:�Pt�5P�"O
	3��z� �ɖ��*_Pa�"O��ijQ	V�AzsGF6�$�b�"O� �P���c0xYP �58�h{#"OVIh�o:[�f�qT����؃"OVj&Pu�^e��&D�b�^�Zp"O�5�ah�D�����
" X` "O�yu�I~�=(�MW�+zLĉ�"OVmap'�0�<�Q�]ecf�Pe"O�����\.c���
]294�CP"O�<�r�9
׾}�G�L�^Wr�9�"Oв���_����F�C�1��"Od=B��c�P�w�K+O��`��"O����#pn�AS�	��5�"OLl�Ԏ�����X|+�/��y���:fZ`�p'������5���y�șop����@ߕ62��H�����y"(
	[�H���M�6�#d��	�'"�����R�G}�H12EGH\ld�	�'�aP�ώ2|�Lq�B�ר:R$Y	�'J0��2o̒R�%� �Aփ�j�<��GS�<��H�H�[Hvܺ�'Rj�<!��S�:O2e@��DF�I�w%�c�<��㈥[�4���S�F��p(K^�<S�Ĭ���Y�J�(4}T%9k�\�<��\ �&�B%�\'!� �h��
~�<	�Ό jX�E3Ū�=')nuh�g�w�<QE�A�YjL��<OC
�W��o�<�Go�� J��Խ!��P:��Q�<�'d�rI��B�j#��U���UM�<�B�#��PK݉iή�X&��K�<���\P���ɤ���B��؂��H�<�R
4-h�8�'b��QiKN�<Y�NG��Ǫ��fJ���bEFG�<��L&�.t�Ql�Q��pP��E�<��#ܮZ&���g';7V����<��'E�k{�d�0/��I�4XZ��}�<��d �E�� �L�Rj� �a�<�B�E�`MVM9�lF�N��F��a�<�� ePP%@f�ϞV���xR`�W�<�4*Z��Ɣ���\�5���"��l�<�"��2]���'	��2ސ�+�H�C�<y�6Q�\��q�z6�����W�<yF�ʎq�jDʓ�> ��W�<��	�&-�2�{��t@n9Q��j�<�HC;Ģ�1��I�J�(1QQ�<9v��e�pRDC�9�b�
īP�<AuퟱH�R@�5���K�z���Q�<���7�&�#�͘4ǎ5���F�<)V�QJ�A*u>Ƽ$��]�<	c�F- ��
�g� ��u:S�W�<��II�)hL"��ε�Y���I�<� ��#��WR~����/(s�5W"O�{��Գ-`ô�V�E���"O���'��i��e�V&(d"O��%!��=}N̻�d� /FX��a"O>l���@9RY��15$�uB  w�ßXx�fP�v����'K��T?�{�%R�$L��BF3.�IS�ֿ��� ��?i�<��5�dN ���r�`ί~ʽ��+{>9p��
k���5���D� ͓�O/ғ]�E&��%0�`{�G�h��ᤥO�\(֩�6�� 
HF��>[��"��0ʓU�	>�M#���d�icą0�/%ް��CV37��7F�O`���'ATm0�+K0Tf�	��-
��ɨ�����f�R7��{,�!��iX�;G�]!:���(�l���4�?�����i�0�����Ox7���3Pd(����c�69AeH��e%Z�������Jj\����V�H�k|��A�t�O�kF�9?�I��0� �ɱFK	T�F�ʃl�5{E�\���Mf�TD�\c�4�C��F�D�8� �>���ߴuJR���՟X+O�4�s�Vu�sa�9\�pl��[���P��O��d0ړ��'�NhX-Y����$�=�	9���^轢2�4��O&�n'��Dto�"��#�g��g����	ğ��ԁ��;�fE�	ҟ��	��c_w�R�iTЋ&�ݔ<$�ZN��,�4�$&X��ӄ1��M��şLT��� �O>�����1��4I�b872.Ta���%jJ����ɖ-�rb�f(�SY'Db�Pz���*w,���R�p8c�h�>y�L�ܟ��	���?������r�8�/e��A�r �7Gt|��'�"�'�ʟ�O&� Tf^����!�;s����l±�McR�i�ɧ���O��	#E8��`TF�	vb�X#(
\	��
 lѽ<�ĵ�	ğ$�IꟜ�A\ȟt�	ڟ�J*�0aQ��` L�R�iS
�,z����b�H�z����o� i�d�Ij(��
�Bذc�n@�Rs�8�Q�קV�6<"D`3��   	*	A��k$H�xeb��{$��O�53Ц��S]���So�9|�&�����im`%�x��˟`�?�O{�h8e��R�Nx�G���pE��'4�"=E��_p&��k6��y4��&��9�~b~���lZIy��2(,�7��OL��~R�M?mv�rR�:LK6��RM U�)Ц�'���'�B��瓊L���I�'wN�8����|
�BٴYt�h�r�.2��b�UX�'� �(���1*7��8v�V������@�$�l������p���Q!|l��(N3c�4����On���j��)�TFݾ�8%���� ��<h�D�2�?9I>��S��?�"L΄���ҢP�8����,K�`�'��6-�o�)w�ڝh��ªP�T�dd�K> �*@�iA�DC���>���?A��x~�U����?)�4{�|���� _�������w�y�G�ϰX�V��V	+ڸ���/A���'�����ט0h[hxe�S�s@��1mP�tAt6�C�?ǔ��S�ND\�;����S�ll���s���磖�l�%p� �wS]KAcc�~���'646��ߦ���~��M�Æ	�O�H񪙽��у�m?����?���$�Ob��4�IRm�F���+�?]�L1�u�Vb�Q���޴؛V7OB7��O��%�g݁1$��lmdMPqL�/f �Y6D����=��$   �   J   Ĵ���	��Z�ZvIJ(ʜ�cd�<������qe�H�4��_?8<�q�i��6m�M�X\�W�]�Cqj`�Jʦ�Btm)�M���i��F쓄�ؒ+��I��+X�
)�G��چ/��3 �"�{b@f�'4mZ6��h��b]BzP�{����1���#�-��#�@�� ���(6�ٱJ�\�E����A�eLIY�ĸR�BXC���l��&�ğ�� )O�i�8_��	P@��V��я��s�H��,�M�'c?��L�Rɺq$���튚R��ɋjt(����Lve(SMJ-VX�Ih�@i"* �ɿL�D�E� �	B%��[�J�ℛv󤇠�O����kG<��ga�8 �$Ւ;�EFx��\�'���'�~]�0��H�`�QDR8Q���cI�<S�ɚ'�qOz�� M�'��,�GE��"�\;D�i�5Ex2%�K�'B�xx�o]�,K�HbLD�-].�D����'::�Fx�N�X~2@�����! �'���q���� �O�BL�7e�� 9S��#G8���Ό;ĀDxBlGg�'̈�ɇ�T�ҰP�;.�m@W�	�@b����IR��'&2�cJJ�r�̓��[�6 ��'�*iDx���Z��9�~$�! 2-��E.1��p0�̀��?�լ�>A����e��s�T�O���;^n�5B ��1Y�}s�4��@A�{
�}�'@��O��)�!�:b��G�>�.IµT�l���I�m��8�f�A6����5�؅Č9;fe2D��h�   �$ J](P�y�~�i�,/D��R#ř"}l����B$~it�"�.D��XvhN*,.��Á��f�F�r�!0D��"���;���s�Ɋ � I���3D�`r�� =���cv)H6V����d0D���q�O�H`��DoS� ���/D��ZU.�1@�|� �Ȣ]y�\sq.(D�h[�F��Yҵj�h�S%�'D��y�e�C��\�g�T=�=�v�!D�D���ߜW9b�j�#�8 �Yڔ	?D�ԣS͔T�J	��ϑ�r����c=D�p(���'TVl�����20�t-pө?D�\vF�FxMa��E!R�45K*?D�lcc���lqR�PB'���[�D;D��a��M�_��H��_*I��|#&�:D��z`O�}f�"̟6���ˢo7D��ʅ��YF|�����	`��5D�1��Ȕx(�ڟ�΄q�i4D��(Q�\�j�    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �   Y   Ĵ���	��Z#tI
)ʜ�cd�<��k٥���qe�H�4��6_?><�'��4f�V�R{�4��#��:��Zׅ�J�7M�ܦAZشIm�$=��[y�!+3��	�� ����摹&~a�灑� 2q�=	�((��6mۻ|\Պ����&��8zկK"��ɦ>���í��$g�	�Es��{��o}�<��H@�,��X��g��"���q@-3�d�#.8�|Rc��r/8H�tEL2td��Ҝ`C�����eӠ�y�����?���(S���	n>��8s�&�#�K�.�kLE����`�!$&6܋��[&F��D���%�1�+���ʎy�e3��|`B��#Q��� ���y҅x�'���Fx2,�!�`�J�d�!;c�_4M��#<q��,.��
���sՍ�*s��5���8#C�%�O0����$���'�b�8'��%&�֡�$�[_�)�4d�"<q�#��n`@�j�%�2���/9|:�E��{�q��"<$. ?ɓ%N3	�X�h�(�Y�8�k�D6?�..i�$�@+`k .dlNXAB[*8?�Ai��ċI�`{��Il�b)8c�9���,F�I&��'ݘ'��HFx�-Wb��	���� �E��qS��Ԅst8�	(f�Lu�x��Q�<�16Nv��y�ƌ�k��X�Y��� ��Oȥз+r�3'lę���E?�d��F����4^u@lI��X�Sބ�a'�	���X���>	�㐏%��p����#F:�
b�G}��a�'M^�Fxb
�!.d�|����.L�Q$�ڛ�y��A d  �'w^h�aC�qĜ��퇾<����'\�t��t�Rh"0'�"e�����'���ɲmҬ]7R����Ö��y��'LpD9���G`^� ��!����'���!�!+����O�}2���'������@�Vx�	Ѡ��sh@���'�	)ad�	��]C!�ޤr%Ƥ�'�����1[����CM��byT�0
�'���@O�l4b��ܞ%H���'q�i(Q ��ݞ��b��.� ��'�:e�%G):����ХF"�F���'��(�RL�"JB����Q���'(62�"��0�JiC���4`,
�B�)��,Y(`XfmQ�g�]� �B���<���ߟr^�[��Ѽ ��ˢ���!�Ĕ,,� �i
&]��j�� M�!�D%��P�MB��5���K�=!�,\    �    �  �  )"  m(  �*   Ĵ���	����Zv)Ú'll\�0R�P����=9pn\�Ёba�#������{�<I�d� �t�Z5$��vT�aN�!@ i®�,]Q�����E���I�A���0�2rTƌ�&���L�/xP�A�^�M� maf�E�m�];g�0'h{G��PZ��xv�Ӳ]m^X�S�a���N�y�D�{�e�>;P`���H�F���;;��ac5����$����72>���)ӹ-#����O����O�e�O1a�Ta��x)���g�%i/J��T��<��F;�"9��(�<1�)ޗ1	4iY����@���DƎ� ���ғEt���0 S���?i����l}B%�iU�`('.�(���x��[=�M[����p����.�|�',2�O��j��֝'9ʙRF]]��e"O$��nں_�p���M��Զ8�D�iL>"=Q��:�?a+O�q�JV�W�`,�5�@���#Μ�q�L|��,�O����O��������?��OYy����
4ɷΔ;o
$�06�P.�Tq5�'i,�P�'	�@ƪͷqº��f^�$ X��	�'X����fB쀀o�~a@�/j<0P	�'����`P�����cb[d���"	�'�PĂB��qr��C�[
_�\Q�O�0o�{�I<H`$4`#ϫ�>����%��6�(]�΅Q�.ų.pA(�N\�;�!�F�a?�d�t�Ŷ32��j2#�8�!�dQ�P��5&��O*Bx�'���!��P%V�-r�*E�����1�!���$-�<��)[ lzP&<p�!�d�Z���bH��O�%�UJP}�!򄍲a�ĘJ��Y-D� i�&�F�A�!�$o�9Іeh�4sƆ�2.!���KFB����7o��Az��ѬV�!���(Z��E	�Κ��;L�!�d�Q9�Y��Q2� V	F0�!�^��c�.$1��¡�$_5!�_7r���R ��9HH��wa��!�䓢.P���f�7}ĸ�1 O��!򤟕o{zH���3b��u�k�!�� +$���BP:�ԩA�g�7"OL����TV�ИSD# V��A�"OB�16K\:[E襉P�^�a����f"O���6O�W�x�A5��&�z(@�"Orqh���?�lP�B�m����"OJ|Q�Aקh�h4A�k#z<��6"O 
����$�!�*�
0kx�"O<<N�K+P`�)@(fd�$P�"O��1V����&���I�J��t�"O��3`ţq�`��3�L�g� ��"OX�2�,E���1��]$6�5(�"OΨ�6�W�x��D�@���Iv�@�"O��*�ON�fX��L�\�r��V"O���t�>�BX�%��X?��B"OnqbG�3 ���΅~-L�`v"O�����?�H�+Nʋ!t@X�"O�h#)Ux1�/adܡ"O�a��ኌE�@I"T@�08V�*"OJh┈	� ��I� -n{��K�"O�i�Ȋ.Y���'��Hq�9��"Ol� �T�>�kS�B�<i&œd"O�3a��w���`&� �D�-�P"O2(�VϜ	��!)���y��ږ"Op K�d*���cN�h|�b"O��Gi�E ���G�&wr�y"O�(x��Ї-��A�m7:Y��	T"O��4oW:Ikp��&mݥfhv��"O��2��$y�P�Gb��!e�0�g"O���b��n�ި��a��b�P�p"O�m�G�DaL�,�T T�Q�Y��"O� ��F��2q0�a\.gLh4J�"O�STB�'e�z�ɤ�^��4JQ"O��Ұh��3�x��R�L���(&"O� ��qC�k*�N�b񺡊�"O⥓��,6p[ P�몠q�"OЕ���n��bv��,�,)t"O6��#�ϫl�4	I�@�#4&4J�"Op5M��]���A��Q$����"O��#�S-?Q`S��!@���"O�L����)l��Z��p�| s�"O&�i��ϊMܑJ"	+:�@�d"OnؙJ�h|R8ѓ��ȍ�"O�*a��q�F��al��)���"O�l4Ɲ8920�qQlا1���1"O���NZ�����6��}��"O��dlL�r�n�x'��XN@ڥ"O�Xz�턚ؾi{�e� ��u"Od�!�%�Y�r��2x,��e"O
�ݝw�>5�@՜*_��ӓ"Ot�[QꌁJÔ(�v��[U�x�"O��{�L�~�ш�!'F@��"O�*�C[/P��a��e�VAh "O��9��G���Rk�5���Q`"Ox|�! B�Ed2AH$�}�\غ�"O�̘uBÉ7�H �3�X<8��qp"O���"&��i�L�f�Q���8�"O��ӂ�O���}*'�N�\�]��"O�X�`�Cq� ��%�4�D�F"Ox�Sq�>R�`i���\-�4ye"O� !��C�P�TU�E@3N�ࡁ7"O8�a�P)�0mN�lJ�Ѧ"O�����=&{��tɅ�3Th�� "O.Ѐ�I�$4n���G���P�"O6�@��;YS^E�˓G���:3"O�D����cJ�hr�<Fq�u"O:�3l[j��H�f)N~���J�"Os�6�9�"۳�L���ի�!��C!=8��#���l�ZxJ�^�\�!��7N}k�PY���`RV�!�$P4v<��O(�h�3���%N�!���'�E�����ĄA��M�sD!�D�,N^̀¤Y�1�.��r�-
@!�d�$}d��"ݣ`L���N�-�!�A�JH�zvm�i�N A��De4!���.:��S�&iތIrs�W�i#!�Ï2�e
3�^�|��a�R)�!��3O�S�a�$���Ɇ��=;�!�$J+$�X��d̆f�Ya��$m�!���b��}Cw��.X�=��$W�!�$�Z,�PAP�ۨdX����'ƅ!�!���,�@� #S8~� ���QzY!�ē�ex$�����O��7�/F!�ě���%��F��ꨈ䪁��!�D��(�@`ؓ�ϫd�\y��*�0�!�� Hb�8���O'E@�-����8�!򤋩;��xuAX�7�J��wl<O�!���q,X�ת�8E���ee�#�!�d�'P�D� V�	��*֗�S��ń�d�`8�JS�#u♘u�k�ޱ�ȓ+���P����|,�F$T�I-ez
=���E�$�F� (�|���<I
���_���*!�>9�IǉX;�,�G. &j(��2eP[�<!Ѣ�5�ʜ�o��F�@Y���^�@X���>R�z\G��%�:A0�璈F��X�B�yK_�# �u[�A��
�.SD,Ir1�8JI���D�d���?�'�b��5h�,yںm	G!ժ5��
�'1R�Ё�
o  I ��R(A,~�au@�.]h���$�*����� ȁ�Wkӯtq�b�L1�����'?A��!�)x�0�Z��2���FR�Ql$��f�Բ5��K2��2�y�2F��܉�Iь L�q%�G����Y���+�BܯXF�<S Ʊ�(�@����#y$���.X��	�"O�R��Y�rQh	�&疇E xe�g����+�� )rnxZ �G�:�1�1O|H�R�רW�<(���G�+�n����'{|I�VV�"��혰ژ� Z$G B�`$)�cͮI렌[t���az�I��|�:y:�!�� �Na�Ƣ]���O�t���L�`NQ9��
�6]�`�c,�M}���r�F�6�ؠrE�ځg�JB�ɬ8;��f����T ��k�˓i2z�V�@�#�@��3#ޮpg ����)E�!�!��F�d���G��!�ӱ^�~���Aԣ:���O4Z8���<�D<U���Z}@ᤝ�T�S�R,��Jݶ%(���H\����C��R�@��(y�@�9��׫@ެ�5)ŎH������|�P�'��A$l�^����)Hu.M��!{��B�̠�ʩq%`�
W�!�B靚>�"d�!�o��d�"�G�<!��.?�1G��.�u"�aUl~bV�t �iER�XM���>ʧ Y@��F
A����F��
�؆�W��\I���#)�Iצ�<|��p�ܵt�X=p��>����O������	S7��@F8�����"O�MI�5-� �Q�~U��)��ii ����8`�p �
�9�4�ԯ9Ft@��:YGjŇ�ɨN��C#�X��y2G>)�� �c�FS�z�b&���y�I�9x`�)� K��^���bq@	���'(XRF��Ef�"~�T��#
x� B��-h� #.�d�<�`
D <)(9�&�(eZ�����L&@�|���~���$�-in�R�B,
��U�󭏓E�!�d��|�	AF��h�-B�|��Ǘ�`�a~2�^�w�R��1�D�@Sr1���*�y"�\]�� ���0L�
T� e��y�OE
+D���&DO!P"�����y��B&)�VXav�@'Xu�� H�y2�άN��y�ՠ'�VY��͏7�y� ��H�����xI���y"�I�q$X�P	��<_f�!2���yB�+T&�(gA��7Ų��e�� �y'��q�	�-Õe��Ȕ��yr�2E3��P 睹(���aǥ�'�y2�ռ���W��q� I��ǟ�y�mS$����lM"6X6�:�+�8�y2�Ƀ+|�L2��-���k刎�y�ʈ_���ң,(y�na$�ɴ�yO�0[ 
c��e �y�`Ҡ�y���-C��#q!�/y�0`�I��yFZTEz�1D�E���Yf�B�y2�̱a���+��S#!=�ʀ:�y(�6A$�p��W� �.ɻT�&�y��̄Q��,Y��V�d@p���y���r��x�d�@�K4	��G�<�y�A�=P��j��Trh|�V��(�y2�\:3h���feїf�!F�G?�y��$`���v�`�И����y�K&N�d�
	a�@��bѨ�y���@S>a�5�S�X:�yR�ĘP���P�#S�h��	��yR�U�V9�����H�����N�yR���H9�d�XW��M���]
�y�K�1W��&�%N��jq�Y�y��Ä j�Iy�Ћ@+bQ����'�y+�3y樢c�/�`@ ����y�Ȉ%,�I���w�5�/	~pB�I+<�4��ՀG�y�� �ψ5<pB�	���E� ��?WI�a���EB�ɦ4pv����:0�j��Pe��N��C�)� X�0���'�f�(�����$�e"OЕq�/��<̈́T����5T���3S"O�5��۸�)�eᗕT��-��"O���!Ȑ:E�� O�7�uC$"OFЁbI
 �>D�F B�*x9y"O�к�E9)w�Ժǭ %T��Bp"O�Aխ�	\��U$�:�2�i�"OޱJ�o�+�L!�����ՙ�"Oh���O�����Dハp=�� �"Ozap/|��!�B�@3Y���"Oh��M"� |�d�S`"��s1"O��	gZ26�0Qk2LT:1*lr�"O 8i�	�Gm�QAPC��5���ۗ"O� �"KƧ=�(�[�'�p���"OTU�ҏ�d�PP�s�Å?��y�3"Oh9'��x�v4s�
�-��@x6"O�⇨��H
��XҦ�2�Ɖ�u"O����l� )Τ�c�sS���U"O����۴�R�Q�J:!I���W"O)a�jWUS �@J֋B$�)2�	w�Z�� mXr��$ �G��6�ǀ5�ؚ�O��etDMs�nģ@!��N��Zb�Å/i��i%L-H	!�̅]l񕂉�Wb!bL
�!�Dϳk�|�H��حy��!jY}!��>�����S'Mu^�q�)�9_!��A�{tp]#ӁQu�4x�j�!�Ė�1�\�F�^�~7�5��J�!��Я`۰@��0�xh���f�!�dQ�o��q*Ò+޸Qss��!$�!�d�9>�H�a�{Ί�B�!ʶ4�!��«@C�{��ќ����+0!�D��N�� � Z�@�B��s!�D��`q���wM�%�䎅�[�!��i�Iy��6n����-L�!��.�<�w�DՀ������Py���"}ΒD����fQ�u!��]��y�NB� THq ����;0�Z��y"�
U�+��٠ ֲ�xV(]�y��?��h���a�̉�����yRM�:)t�B*�,�dR��O��y��� � �h^�!`�[��yү�!���Rf�	d��������yb�;C���!&c8RH�@��y�`�iM�AP��mn��ke���y2o�~�̔� @I�bm�P�e���yBeOt��Y�LٸB���-Ԁ�yrϛ)O���k �0	�B��t�\�y2)\٢\�D��*B�rW�Y�yR�$o8��ІO�{*DZ�L��yB �	n�H�C2 [I���7���y��V</v��$h]�����M���y�O�U$n=�c[�R�hSV��y��&��uQq�4L�du���?�y�A��I/���G)�I��䳲�S)�yr��#�T
2�C
l ǠH��y�/Z�t�z|�v�߀:��uZ���y2��o	thl�3FƠ�#��G|!���a�"e(��I	)W@`�Gڠxq!�Dn>��(0�M[��I�̲o!��/q/v����&�b��!�ܓR@!�Dݤf�����Z�SD&D �ax"퉚4�(eХ��6�pm�bP~�jC�	VD%���U�$U��)2�C�	�
�pA�ҮU�Y4�qj7�KJ�0C�)� �@�RXw��J�lء0g��`�"O�a�nS�)�>��kX(b��t"OfѠ��K�Om���R77�$}�$"On;��%W�@Y�d�[y$<�f"O�0��/�2�1ƦP�Pn	�"O�$*���0t�[�e�}pM�g"O�h�eo�4uxD�%�I
p+w"O���)Ā~�h�0u$�8	�RS"O�,���jt��	a��]��"O��Qd��`���&j� �S"O�����M�~>T�[�B��zU�H�"OL�*�.��c"[�qR�E��'J4��[�x*�`ܙA�l(b�IW/�y2͖+[�t鑦b��lr�ډ�yR��'x*0	�o�5Ka����P��y�F�>
��!
7ni����)�y"ŉ�'��-�u��k;��Z`۽�y�"ˮ2�0�	-�j�2�ϓ�yҀ�0P��1�)�%�n(�!bF �yB�� h"���g�	4�`]���\ �yR�D,�� *A�)+^j��yB(ݤ=�DjS�o}UP���yb!�_6Ҹj2�ЭV�FQ���,�y�k�8Yh��#H&�����'�y�-ֵ!�`|�0|�r�A�8�y�jX�o�0��PȷGT����݂�yѢ>>X=�� ;�����	��yB�C!X\=�w!^�.��Pq!D��yr��t�<�S�"�|(�@��y���]"$�hhL�	�kL��yb��놌�c��5YShaX�݃�y�J�A��c���M9xt�ĩ��yB�վ d�s�/��GY��Ʌώ��yr�<�f��0J�n�n�zE��'�y�i����u�\0w��ЄdB��y�@W���D�w�� o�
�����y2�7^$Jت�
R�g�θ�-��yb�G�8Yxʍ,m:��2���y���<'R��O�7-VH�T
��y"��=�`�DL�p��1�y�)�I�	��[2��Sţ7�y�JL K�p=�C/�?(|D�����y� ]�p/�|ۡ��62�l5KB��y�	�WԌ=��#�~Ad���ŉ��y��.8�
���4g�"��ܝ�y�e[  a�@œf��@�%dJ1�y��ǀ?���Iϊ����3ujʂ�y�2)�p`N�:]^�"�FV��y�!c	T�b���B]�U��+ �yҡ.k����U!���h��"A��yRυ'��9i!�^�� i���y��[�E�|*�K��k�̽BB�#�y�Ç�m'U���4;�ɛvFԱ�yB#�8)���
�<a#\9`���yR�UR�lH��D�ѕ���8B�I0Ba	�pe��#*qA�璸]��C�I�.�(���˻	������I5 B䉴oTP)s%X�|��q��@U'
��C�	�>�jt�W��?/�,`�'�onB�	 5I����9#"d�c�NbB�	�.̄ �I�j� YT�Q�P$�IR��л�'��Cz��
����*خ�{g=D����c[)o�,����RLA
b�(D��F��XKh���/�ٹ�I&D�� ��f��=�L�T �9&����"OH��3HH�"�4�a��iʍ�1"OAb7� 7a"<9�F�&qN�UPr"O
٪���'�L�
�Y�D ��"Oz�KC��$A��)��(�'�&4"O�d"�D)e�F�sC�W"L�^bQ"O�00�NN ��"���&X>x�B6"OdT�Q'�<(���BU��}A�}R�"OzmI"�^��,� $M#b{P"OKۖO*��wD �"�̉3n]��y���}��F�6"Xx���K��y���
�`�7���Hp�z� ߇�y�!�;n���R�-;��XS��y��KZ\�s!\�$P���-�yr#��<a��۵���	#�?�y��H7r��-K�J� �B0�o
�y(P �����$��ٙBA�)�y@���u��\ b�񨞠�yB�ƨz5P�H�D�7,%��
�,�y2J_��h��U�'2�I2��C��y�j_�wvJ�Pq�N�1��Сc @6�y�N=�RH˦�>����� ���y����q���S�V�3���;V���y�R�?��X�D�1��D�d����yҨ_�d����W,O��A狽�y�
J���9 �d�	��x1 ڔ�yrj ��^#$
��mE�@��y�DY<�
7��8\\B�{T��y"&��;w�(��hG�Xjä���y�	T50溱9�,�7R�*����y���%����1P*b�IĒ�y�
�Ա�_6m�P2'�&�y�e�1pəRIH���@y����y"�ݬ:&MS�b�87�D�CI���y"J��q �4
I�M�R�-�y���_^�H�/Z�'"q�g��'�y�o�"f�´HU�Ң.�537�P�yr�;���H�G$	�Å��y2 ҋB�8�����&f�����ybX?y�v��呄�8����y�O6eL�!�"�~BP:�Kέ�y��z������ds�͈�y���Bt,��a��`���@��R��y�k̢Kh��C��3X��#�+��yBlE�_q�X�+�
K\I")� �y��N�[�^@��G�1DFMB�o�2�y2HD'`��<{�dҷ,�B��2�T�y2W�]u6�с$�#�]�0� �y�WD>HɣG�ϴ����yNE;Nv��C�
�
�RC�V��yBF�� �LzdF�W��B��yB-��[� ����|�D9jҋ�y�O+p3�42C^� q*q�R!�yr��j���a�2X��p �4�y"O+��@b!�0��(�����y���<Ѥq �F_9i�&$��e���y"k j��l)f�Fc��MC�K�-�y��&P򩺴gH%[��YA�j�y2EǚInQzᩝgB^t�6Ɣ�y�gJ�F��ьv�f`��]��yre��F�H�"ŤM'$�NYҵ�@��y�B�8I�<����Fi�5�G#�y�i׹I8,%#qC���d:%	�y��F9K� -j%$�fd�!ʺ�y
� �x�k��E^&{p@�=F(�X'"O>�#�h�JC����)
zh�|��"O�,+o[�D��Ѹ�.Q;ZSZ�[p"O�|�O�1A�� �홨L?���%"O^�!�-�y]� Aި%���+1"O8�8t���su�Հ"�Q�j�pV"O�(�p�݋�sd�X@�$%8�"O$	;E�()4̤	��@8��P�"O��*�1��Q����Tn�X*G"O"�[��ԛz��y`N!J�%��"OFt[B֊~ܸ�A!�#���"On���]4s�ASB	W�\�18c"O�iV'�
^�ܸ���O�t��"Or�ɴn����51D.��AFu��"Of	9Ń]�2l�X�Ы�!W@$��"O��z�nU�YKl��o�kT�:G"O0�u�ƛd�Va�4��?d���"Oҙ��G¤_U���nPQ��s�"O,�9�B\;~i���.ŎW5���"O&�IW��:����L�0F.��:f"O0�"�(�'|�E���P�0�g"O�!�3*Y T+*�  ��7n��Tb�"O͡p�9%�\9�>(P�3�\|�<���J�"���kW�ԅ)�te��ds�<�uc[# *  �   M   Ĵ���	��Z cwIJ(ʜ�cd�<��k٥���qe�H�4��6_?><y�ʄd�V�k�,h"�l�A���օ�0267���հش=�D8�IBy2 ��E�@F�4mBԁ@�ϻU�,u���:$c �=�G�"�o�6�"eZ�p��7O�|�	3��
;2���<&f�J$a؏U�Ɂk*���Ȏ;q�I U Bd����:~�(��(�,{� .��O|p$)
�=��'�D��*ʟ?#�PȓNUoO���$DlPN�o�Z��ΓC���͡<q�O�e�P˩('ąm��6$>ax��L���p,O��*��J�)7�jC�䙲��Y�y!_3"���Ƈ,5PVN��yb"�w�'�L8Fx"c�J����f�q����w����#<�)T���%sp�����T2����&�W��O�)ێ��J���'�L��I�=f࢙R3#���:ͩ�461�"<���9�@�&9;��Ȕft��CV<�����O�H�� "<A!?A�͝] ��pON6$��s2�Ly�B�'����?9���JU�tȃ\��~t����2ܒ"<��a$�L4���H1*
�i��G�9kp��l\= �1O��	����1�ē:,�"vɉd
�yY� �%G, ��4NJ#<ف&6�[?Q�L��v<�k��o�z��%���\��P�l��O*Րg)"��'H*ם�f��`eύ$�R��Ʈp8��=	W�(�S��'�$�ޟ�B�kB���<���O �Ȋ�� �O����
��~�z0j�	Z�iR"O0�p�  �x�"OfY��IE1{�%���L.P]Z7"O�Y�D�1 ���)e��H��"On@S���9Y���s�ıS��T�#"O�$Ѐ#�Հs�a�Y[�ъ6"O�d��J�:�I1�E�$fИ w"O�)�9R�� pХ�\�հ�"OHu{�̓Dm�1h�d
<q�z�{�"OLx��Eƾ( ��uW���qȒ"O�8�"��V�9�2k� 3�ڑ�D"O��xs�Պ ��0Ѣ��/�u!w"O�D������� E�5F6x�'"O�1��/V�F8��Q3E	 "���S"O�li6�z0n� �_�N�P}�"O�QP��s��k����	�4�y#"O���c��0=v"�'�+���X�"O��ۦi6��yXtf��l�h�(�"O0�AE�(X2�9�c�D�.����"O
�X��Z�h�xQ�)*�����"O�}rd`S�tC19F�5uk���	�'<6�c���#�XI�@]	E�| [�'��Ĩ�� >1��bc�+,lII��}�65���1)���
���x�D�1�x���K�Q��(��|iL���E�'%��a����$p!�}��{�Z�@�J�8GR`����#����ȓ^ځ@��<����R	�Z��ȓ2�J�x�d�[m 0�M��M���v�����L@�+�b�{�Hs�⑄�N]�99��K|���g�ѱc�*���AfLZ���4�*Y���Js�@�ȓV�b|9���>3��c��+�D�ȓ8{�I�D���:
��` ����nC�O]�H��jR*�>G�B8��[ݬ��JB�8!���Jӌ��L����ٕ~�lHI�g��gl�%�ȓ	�^���)"�>P��I�TI�T��*�4{���1���iE-SL�&��ȓnf��jWdǠ<��v���ڝ��y���v@�H�̩��f�yҲ���^�5��.�!����з=����Dr��bR�Y������0��ȓL~zP�g� ����Q�܅3�>e�ȓ&"���oH�w�L�R�SC6Y�ȓS-$�K�ʈ�x�P<�3 \ �"���f�`T(�� tX����"�h=����k��EAd)E�m#"퍟D8���!̪d��<Ԯ�btGA�Mآ�ȓ!���Pe&���f/¬	�"h�ȓz��iҡI[���Y�͒#e�Դ���R��ī=;VX��oWH�@l�ȓ.�|i�2o��R���a�&97�хȓq��з	7_�u9;Et���'���wnƕ����V1B@�ȓc�8Eǘ�<N�� �$ձ\�~8��L)�I��)�f4�ɐ��*|l��ȓf<�mԤH
da�p�j�t�&)��� S�LEB��'�8�L �-�
4���� %J��X�'�\��¦�v�:ɬ�'q�Hs�.�4���[e"��H�(���� ,�� y*zX �"O� \m2�-�5��\�Aˍp��Ȼ �U��,�a3*H���)��<��*�?`�����W �6��l�E�<!�͊6 �t�� ��.��)�����<yC�M�Dy�­=\O�����9�
�`vm�y��	��'�����O;3�ra�E YjN��'�K�f�^0��y�"@�lQXt���T���`�!�4�O8��f℃\Ӭ����)�3d��c
�w��Hq! ҠZ!��77L��r�8k3�I� �*X <@�C՚*�`��N�"~Γ^
T�
�W/7:��yqJ�i�Q��9������Ϙ ThY�p t��I�y|��i�'B��$��F����
�J��ez���a|��
#Ḑ�e�ӣD�d��k�d�5	�F2p�a��'׮���AQ�W��-��������䟁?��u������(�8PI�Z7 �h g�]�>m(q9"O2h*B�\�^��m0F��7o�@Г& �Ĺ�uH^���)��<�Q O/OK���8*����\p�<�B�Sx}� ��]l��t����l?�3`E�-��h�e���G�EU��� Wb����	��"1��'��r��>FP"��'��P�<��'�l���%�	N��Cw�I*���'��mV�B8'����JJ?���S	�'�d�"J�"h���8V癈Bh��'�~(�����<�P�됞w+bɲ���^;�>9(��W����S��0d�]�oK�!�$��P_x�T]�d��!�n2p�]��A'O���hQF�S�R('��O����6Kv��(.�~��7"OD�8�P��%��x H���@@��9�s��Y[JT�'�T/{��I�^�Ԉ��;M�� "pD�8l�
��d��E��9�m (���Q�F��"O��`c��)c�Ԥ�sB�`���'�ea��JSB���AMGG�ȓ�}��2 ���K�e��( D���79�O��b3�_��$�k��D�2Vz͙	�'�L�
�͂0Jz�p��@�(^��ao�+�<(�$癀�A�����7
�,�I.�\�șw��К���P+Rh�Ј5q�X	�']�L��;�7��i�����!ʗK3N�p§<D'�u��-L�T�d��'~2�k$�ݗ��	=l���Sႆ$"�KfD��4�4��d��9s2���}��!�L�$S� �i��%����T�\�1Кt ��H��B�J�K�I��q
�'�M��`\��� .� |���B�y2N��~�����7h�4��h�-��wȏ)7�e��[�I�a�$O��CBڇ#�Y��'/���P!�z�b���J*�0R��Έ�T�'O~�ҙ�AB�#-�����|�l���j�(� z�w����5F�h}� �G�ۡ�i	�'����Ռɍc��X"w�Y~��e����Q�0��H&t��e��j�_x��H�,�a��pz�
�y��M��O$��%HBaJ��׌Ϝp�D�	�v�<1��]�\;rAS�B���%C�+'H1I£�.C���b�ه^4�͂"�$>��bĬ�+S֔u��	�;�6|b�˔1n"ɚ�����RjȘل+וO
�eKpi��L�r���J�nu������� �ѱH�y[c���N��AcJ�sH��'�� c�؏wZ"�&#���s��06Z�� w�D�@mօA"�9��(+EtP:�Ɲ% �䑛wo�U�A�'X-(���V0$�~�K��5j�}���C; ��q�РxP`1R�M�^�$�c�A�@�1��E�"6����O�r�(Ѿ,��'��)��Y*6�����[�:��э��d��2s�O�iC�hj�DV+pB |{
V�t��4��2;�:æ��6v�b˓>���`,;,O��[��LUߊ=9!�E,����V�t���W��+�nK�#��1��ն`LL�>i��'�M^�0���i��(D���Ñ\��	1��t�M;�-�H7�������s'N5 �l����c7�>���I�F*B+�? ��K�*P<�3$]�|���H!� "ZM ��UJ�<T����w�^	W 4�����X���۰<�D(�2zz���g��n#s!�J8����j��x�2h�L�A)8���@-?���`5B��7�е� �"O�5�6
Ͻr��m �B��$� �Ap��S�I��h n��Py�#}�k `t ��������
B�<	D �8i��xK�i��;��ġíѡE���v+w��b�����H���G3�Y$F;Yy!��H���j ��n'���f�F�W��	���,���Vb)|Oi�DꄖVy�\��3a[�j�'n�2�ٕ �V)��i����NS�R�~dpG�(�6��	��� "�zv!���Ԉ"�O�rU41����)�Tҷ�Ա�h"}���0@|��70x�y�@Q�<A�jTXP@�`��3$g�`ƬZ7�RE��EU�dC�I�k4Q>˓��8;��8�����[�&����ȓS0R|����l�F�rQ�R� K^�l��u�rm[�T+n����O�]C�:�d��qmH�y�{r�֝۞T��g��������TO �ք�`l��+D���
W>Z�^-qg7p&��@�+�I$V�Y��蔯~��>E�	��}��KH8RP@d"�L)D�����P�����K�_&n Q4-�;}_�"����	N��~Bi�)H�M�1�[�nɚ�dņ�y�k��(JDO�Y�X�"P%ƍ�ybI�#F�=���'eĂ��-
�� Ϗq��x�?L�9��q�$��P7Qф0�W-�7=� 9��-D��p3̝���,��/[� ̼s'�&D�$����r��8�X?�)��"D��:�,�
1�����?zٔ@
C�>D��Hǝ3^μa�`�fN�ɛd�>D��h4(W�s�� �Q�Jt����+D����$f|��f!M:L�6'D�l� �$kVӃ��.��ܙ���� I��eta|Riؕx30q	AK D<�u.�0>)�`�.A�xa��L\�{��4S)����ۢR�\Ʉȓ=�B��� zg^9�4���`�|������	�g�O6�#i�|�ӌ�i�:���k���y ���G$!B]B�nSL��3+-i��5��Q�FĮ8Ѷ���=�Ъ�ZL��~�� �u�+@�؊��U�U��K$U�.�H�㉒V�R�3s,�Uܶ�sPJ�<�h̀6m3~`p�A�V�W��X�!�'��`#��`���I�$�N1�
�+���@�+���W$��W ��V.��+0^�' \i��8|�B=K�N۔Q~�H��^= �7��!��]G0-��&R�}��ɂP�ڠ(ƴt�DҁXa6��G��-@����X@:%��O�"�+���M7g�q�r�U(:� �  �J�5�az�j�A�X̓^j��h�DηE/���d�Q�0�~iI�״SC�|;��N
�`�ח�?)uϵF+����!����'���t�է,��"�h�Z���L>)��CX������@RU�2'ت�2ԐթK���	�'��<��Q���l� j��G6�?��l��$4q�FI�G��y2�9��xV��j�Yv�J�T&%Ё�ì�1U�L�1�H��b�'2b���<���iÌ  �tR�R�z�rP��	\�2K��j6$C�ɽT�.� �GD�wdA:\XK��ζi~<����dB������r��d�V!��? Pp��z?1Ǉ��=�9X$�O�(�x2�݆Y�=�`"$,O^�0��S��<kܴ
i��T\- 	� �0��K����^}��ѳx	,e��Oqy��W
A����Lr�I�0a*W������5�8Od=ڥK��`e8�4E���˷��G�b��� M 'X�]�I�(��H��1��dQ��K�:�Gr���
�FY����آ;� |�b�A�\Y��E�Ơ���K�O����N�R3d$���S�|�Hَ\N@ �vb����?�Px���o�2�90��4��"�+1hn��iқ���.�,��f�n�>�) �n�D��|�n�7\�
��Q�R0[�4XE%FjX� �c�$c�
�y�Z���
Z*:���.�-��)��Dl�^Q{�4q�ص�M�"~nڮ/,� {Ce	,���@�
x�O��!���z���	Wed #�UNJ��#KY'��I�l��lj��\X��y���K��ģ���en�(X�ě6k-���=a�u�'UN�u���?K�`c�Θ	9�<���9D\�%��'�MԋόO�����,L��C����h�~����]�tY�� E�%n��!�CA"�!��ŗd�`T!wj�( �sR�A$D�!����`�pP�
�����NS!�#�ڝ��I�O�
�����%!� w�y�$�.Oٔ"t�)P!�dӃZZBa*QkRC����c X�m	!���+z1�(I&r��d�q�@�K!�$�φ�H$h�03�� ��34�!���~�0��6.ǁj��\��n�>}�!��
Y�XXcCY�f���@�^�!��O5��e��H��S�Ʌ�e�!��Q�Pd�O� t�,�!�� �P�c�P4"i�Տ�mX	�"O�%8�mR�#���0D�٣[�T�4"O����BOS$�q@!4��"Ot���B�*�3R��K�Q��"O<�����H?��� ��Z"O���K�#b��S`�C�p�L*"O,}ᔯ�N"&���Y0X�hٵ"O6���(��:�c7cP�P�XP�"O` r�F�M��2�m��~��4"O�i�ӌY4̖�a6>�%lO��y��ا[�����Je��f�A��y҉&0���0�(�NW�����'�yBL�=�f��̩~e���b$*�yr'S�I�v�C ��8`�ĝ��y҇G-"B�D�E� v��yF����y��{��er��}b���(:�y�Cԛ3ʘ����t�i;�H�y�䞁,<���˜�\�*�:!�R"�yB	�t���Q�"��U�>i�`���y�%�u	<k�њ������D��y2�/'N�,rC Ս�&��Rh ��y��I6O��2���3}�e:3���y���7ܮ%���
5��(٢ �:�yҀ�j^��CP� ����=�y��`��aϾ�����&5D�p���70��d�68��-3@l5D�hj�藇:�%�Y�^��c7E<D�p�bF��\v���f�U3��L=D�L{b,ښ,h�
�'F}�)ju�=D�8f�66t�k� �[�4�91F;D���2��y�ұ� �U>4��#6D�Ъv]�K��Spd_�jt�27D�D�2�Ջ@(�1�?�ѐV�3D�x�1)�h�EJ�C�	��a�#:D�����6W��+"ݍi����%<D��3�IǢK1�\8�iO/� ��(9D���ᄝ�nM�A� �>�ꠘB�4D�ԋ�^W�����	Z����S�2D�3�N
h�N��`�K?v����2E3D�8��4�>���"ǖ{r-
�#1D��(��&Tg��9��ѿ7��(��.D����dE�xAK��6�zܠa*D��!!��DX�X3���8�T�r��5D�8sB�'A�$T�C�^�^sD3D�����ɣP��l�q��.���Z��1D�أ�hK�WX.3��D=D�� 	T�"D���a�v���y��^?Q��QBn5D��	�Kфej����Oe����$D���M�\�x`�R�(�j)�c#D�h����nn���e�!^��1Po2D�Tf�alHU{��+*.=��3D��I��3s(�ّ�E;7P	��.D���𤘋+	Rܱ�dB�y4F����.D�$1��Þ*��ذ��/�:��d�1D��{w@�C���� 1T�e!�5D��qnO�e��&� �Xc�'D���N�9Ʊ�P�S�<^�`���0D��١�.�R���]�~zu�WC*D�8����&OC�i�O۪|i@�o+D��x6��	"Q<�i���6�HA��c&D��&$%=T��Y����0��Q�3D���A�G�7k���*
2����!2D�`�І�F��XЂi_+���ڤ�'D��h��߅>����%�ڷ-{�)׏(D�� �I�F�"�S�]�xK�0��'��)@ �$*CI�&g�H�@��������rd"D�h[5鍽{�ޔ1f��<Fl�\���"�K� |sei=�H�(���n1(��q���$�ʅ��"O��� 6��Irp��H����oذ}g|Y����)��<�qN�xd-��/� w;��T�Mx�<��%A0��k5\6����U�<q���)���a�%3\O����#ˬE����F<�)�C�'�,���X/�L����fA�A�*W ~e 		�	� �y����:ij�l�6l4� ��OM�@����&�(��Ă$	B
d�^�13��0A��S�"OY��� ��!�f��()��Z�Qf��`�H_#��)��<� ��1��E�$�~5"(��G�<iW�^�x�<��w���e�����`��<�g,CzXr�`&J=\Op�z���i�C�?	X��q��' �U�r���!�� �C��"�����m0Bԓq-��y"BʒY�H
�k��b}�q����Oꤢ�� /����$Xk�@iU�4#2p�R �Y�!�X	�����L$T���ψ1(����Ѐ��*ږ��L�"~�|�����U P�j,$�@�ye�]�ȓ_Q��X3�ʀH��L˲(H2f�h�ITP7��Ű=�`���&����!ȝd���
ҥFX���5��	B�E&,���L1hQ��,�$�y��؟z3�]����3�����ą�y��,ݔ���'Q9#,��C��y"fɨQb�:ƂAA���p�dѥ�y�Nʊ��6�M6.P�@�K� �yԀ)��MΫ_�`�Wƌ�y�EM��J�ΑLHμ���A���'Iʴ���R�S�'9
�*�̜<?6�H�HD~�Є�"�R�ʔjR.��cA����FQ�o�m�ɱ�LE��Oq)�%ά0���Ɖp�IjdO�t�&B�ry�s�,�6d�!�#�Jg,���_���>�0@'6Z����i�NR��rA��wX����RM����R�h�Ԣ�=E 49�a�0u�i%�-D���ǤK
��[�	ξW!�PL*�S~!� "�Aؕ�M��B4�c?����t|�9Q�B�#x0X(��+D��dM>Q����F���~�᥎I���+۾Bjn諁H�[�vb?%�Odhk�a�0c��x�5
'd�HO^tЖ�&]�򙛣LA0m�SÁ�n�tQ���߸8�P q��<0l��I�� �ʀ�ߒW�(|`j�"F!��D�>&�lm�� ��D�J$1c��$/�=��"�Pn���Ԑ� |��\s<�󌅠>�f�34��k�(T	�%8�\ ��-����Y�L��:U�ܴ��D���%8t�	���%	��n_�T�t��-�S�r��B��!�D߄V��;�lK�(ؽȥ��/��!y�� �θ��`�	YTX���o��% � e^@U9�NE/,�^p��O�������y�<H�E�-�H��I[wZ�)��]�r�hR�̣i&t��Ռ�iq2��$�'3r��C��^����v��	aO�eb�'�;1)���2/����:�i��Ǻ:R��.8L��M���h��ǉ``�(��ďi߈i��.�|�h�o^��ZQ��N�-e�bL�a`֩
�ꥨ�'St: ����UA���d����V������^eo��za�W{Sv@�O=��]Y�F��|���w�N�x@Ư~a&މ|"�=���h�@�@$F�d�b}	�'�Y�]�և��QKz�+��gv��eˑE�I�fr���%�1��S�~����e
/���[q��*=�џ(��"�/��aҖ/�2|�������@cœj�>�����$�h5���|��]$�l1��I3+������<r:0�E囚g�\˓C��`L�j`��#u��j�|#}�K�P��u`�"^-vl41y�<q�H^4{H�r�)R=Fp�	��E���yy�G�)6�"�sTg_�)Xȭ'?�ԛb��)zc$���lڨ�`c�)7�Ћ")�kh�IW�#3��U��ʝ��=��!Vv� $S�e��P97#Q�F���	Y@��ݰ�O.OA���fw�3cF��y2�g>�3ǓQ�F���A	��y/�q�^u$_*1Ķ�X7-Y8��'�n��6l|�G��됇@��8�Ԧ�4,�Y)6��5�y���-b���y�m�.[�`�V+H�+B�B6l�����:PQ>�S�? 4i���2u�Y���S(~��M��"OHI넀�) <)��,P8.�>4�4L|�R	� ��ă�|��qArخ��r�z�"ܷ.q�C��c�X]�� ւA4���	��y�ꝌG�P���/?k@�ywa���'"����N�P�t$��Ӿɪ񙗨�f`�8P �I�C�I-+�.���O+Q�paF�5N��͊m�X����*O:�K��Y�TA5b¨]�s�Eܹ[� ��!/D�Ќ׀TZ]A���1�lӘ�2��@(,$��J!�'���5S!`Z@ڥ�9$���
ߓ\_T�S��^-(�
6�M�cOZl+f�4t	���� X�Be!�d�t[�����P�S��[ i�O�m; aL(�R����0�`�F�uY�2��2o!�ċ�ٰ��jVH��C뙉'�̋��J�b��OL�}��9�xd��M�હ���,�� ��$B�䓼r��K�F�MB��ϓ|B6����>��=�B�CJ��yI���N%fmb���C8����Ʌ�F�d]��Z���n�=Є�G��,2�!��=w�A��@��!Su�ǅj�!����ad�@�G�T��b���!�Ę�}`^��ŝ�D�{G�~�!��L�cU8a��O㪬�T@D��!�""�I2bo�7٪L�m��\�!�F!L|ꅩJT�i�aPSU#|�!�DN�!].@V������Y�K�>X����VP�0��\��@Ӗ]3�0�$stم�0o�*����̟��gJl��%냯K�l���Ǐ,D�P��/����$q�M���4��O q)`�ϒ�~�eϡR����G��A�O�B�QG�j�)�)��n<Q��"OHi�dI�0�$0�%gG�e0��7�O�@i@sJ�Yw~�Q�'Q��Pb��h��Sq�{�+
�TXђ�,ON�����`�*z��05	�`�E�5,�M
pj�aB�$	 �&�?I�Y��N�)v�/lO~ęU�(d�#��	/s��a[��r@��\�����ȍ=���0�����)�Ŏ^3j���[wb����s�,"�
4v(h�'۸��@k��`pC��P6z\6AX��
�.���F�U]}��eaנ��+C�|J��y[8Yp�w?ęz�^!6F)ф�v�p�(ӓ��`R�*f���A�U1~�~m�b�Q;��QwkI(�q��ו)n��î�p�����'{�nu�Bf�
>���<a�c��98������i���Aov�h���/Q��P���N;O�!�֌@
�Q3���*Bl]���J27زP�s�^+-`M���x��8K���$?��]�
�8�hy5�?ZA�b%��pf�8�S��M��ȂX�<Q N�Gx��r�����
R��h�g/>k��,<�y��E��CL^�1�
O�%��HD�RV� J��J:�L� o�m�T�J��ȠO��{A��#���ʖ�ĬQT���z?�o��A(~K��M��8:�F8��l��F.,O��IԨ��v6��48�]�ʲ�����[��0�$k�K�S!�K�I��= Q�Mcy2�E�+�8�� �a�~����V03�@���oFwVO���e	�<����4k��=�e,��R�:�q��t��}q��n��
���S5Z�j�@��S�\��e���I$�'^:h*��A� \t��#�Kuh�� �B'`i��@�z=�ԉ4�W��h�0�ӼYa�ѻjP�6��m��_��ć1�A�fAV5���u�B-v�ب�E�$b4Pc|��b@g�z[I+���V4��'���S�*�t�@SN��*]3u.�9@Z���:-I�Jܶ��V=9l �$�Kc���!!M1Λf�G�	��� Hg�ӧ������o#�#d�����R�@������z����0|J��ǺC�l����}�̭+���^}r���7����4.Qx����S�}��9"�)��;�M0��P�{�qO$�p��@	���S���\J�@�{� %��i�`�B�	't�`	T���qKʘbC����">)��N-�ȣ|T�<(��S&/��?hpP�,RP�<����7 ���)��w������E�<�e1)�2�+�$S�R�١�%�}�<�a��F��KvC�K2�a2��}�<��JC����j��MG�%��a�b�<���Y�FE6��dɚP�P�
Z�<��k�$��$C�ޛ0��@e�P�<��8y��@�<��UX�+Q�<� �10W�'%jl����ш,Z�`�"O�"�S2�|�2�S�6� �i�"Oޠ���n0��a�T/��Aiu"O�����ОMU�-�BgM �X	�C"O���nV�>�y�#HA�,��"OpP��İ*:�X��S�1�65!!"O�#AF�1vq��"�����"O��J�DL�ð��ʆ��I��"O�\Ba���B`Bn �?�luӴ*Od�Kg�[��=���27�8�	�'��]�df�/;Y �*F�%�"��	�'�EG�D�i����/,l��@�'Ǟ)Q�(���L��ō"e�f�#
�'mx /�fz.��@�>^�0�p�'�
�p/4
��p�G\!y>�8	�'��i��W�� ��g���49ڽ��'0f�	.$r)L��e>Y����'�(���fϨ��i�Dȣ;���'��ar@Z�,� ���5ː`��'�t�����]�T(�A�.[w�Mp	�'��,	��R-Zwba1�W_����'�j%0�ƈ�3R@� O�W����'à����/�8�d�E)�)��'u�x��"ε��*P
M�:"��'m$�Z�Yuj�R��F�2�6���'����cH�,���fX2%$ٺ�'�6T37Jͦi4"Թ��(:f�'�~-���$(�F��$C U�&���':a[�$��n���\ �����'�~i�e�֓M���1허)����'��k��>E|�a�`���_�4��'@ �*�͂c��tBӥ֟C]��a�'����`��7���z��;�8I�'�L�鷈:w�ā��$֪S���
�'4���V�^<�%� �I3��˲#)i:��Ë�1-����|Oȝҁ@�Up,M����<u?�]��e'
�y�헰+�����������L���fɊ�ohy��,�D5��ȓ<�p0C7HY�{@�T�Hr@�ȓP��%��^� ���F�e����M�����G3V%�-�"NQ��b|�ȓ*T�ƭP���ӧ�	����<�ÇGI���O���J�)V�@Er�Dd��
&��'�`7��؍�'���B^w� �3?�')�d�$�4J�f<���V\���kFA��E�,OrE���O=L��W%]�,(�hT�g�B1B��T�|T�	U���(1��	�fǓ0��	�M�d�8 ���@}rh�6i@!�֡@���	Ll�OE�Ub�H��%v�u��h^B�HSd�V���Rr�7��%���O�?�yPƋ4%�А�œN�	�1Ad�L[�@I�A\8�'���	ׂl}@��"l�,xԜY�)�ZQr)��'�,Ô���Mx^Ԃ
ç)�R��G��jѨw,S�R�x��Ż�~B�=c�P����+����O� J��p��cyp%%�����8=|E�X^M%�����۞r��d9�����d��K�UD��!7(�<a�kFy��IZ�a�J����w
L����تΦ����,��	�'�8<'?-8I~�6#�20eb� �q�$�6"
�h2И�0#�V�m�;a"��}n:�+	�{Q��B���=�4��/O�V������������|xX���S�{��@�b�*wU�  BF� @�h���OV��'@�2S�W�?����j�|_�<еJ�xg(%�@K}"��.U[��3S	I%���Z �\ �+ZGjX 5l�	C�D�$�����x�f�E�~�>q(7���>sPF]JY�@��`��S�p�^3�ݠ��Tb�ѩ��\:�!�$-]��J�O 7.5ry@p��
%�!��/1�X��AӑL��(c�'�;e�!� 
g"�9��L�S�Z���O�i�!�d�>.(*yJR(�8φ(K#��2!�� ��S0��?iT���J��p��E��"O�)pE�ڸ��q
���7����"O��!���o�T�ZB���8k"O>�`%o��%���($���mrX��"O�I��ŨN�@"q��M���ɐ"O�h��K��P���	��=A���"O�;��Έ@r�� ���0/2F"O�%�`����	�b�:"W�c�!�ٳBl⸒7/��>i�	�v�ͧN�!�_�S��`��-4hf��nE	2�!��4d!�Հ�m���P�L�!�FY�<=�;U6����"�!���I#���'��I�pxQ�B�[�!�P�R��A{U@V�H�P�����&&�!�dUz�>�o"Z�&H� ��!�DX%=��b��&Z܈c�.Sk�!��-_$*w[�byI��"!�=~�,���@e>NEZ$��'p!�^�@�Z�0��L����-z!��2�`�"�F�SH�!#g�<r!��3WO��j���a>��B#&�:gp!��w`�t%R=r{7JB-S!�*W�|{���-�T���F!�%)�����_�m{�@�fA�$)!���{���;rT$d ����>Yj!򤌆@�T�3b����E���]K!��[�R��!S o�w���(r��y�!��-?���J>|���T%�?F�!�d�.���g#R�tx�U	��aK!�D��_a(��ԁ̏P�ĹQ)B�#F!�כ[� �k��(��	1����m�!�D����4#P ��0Z� T�A"[�!�W�y��q����O�@�	㉈�!�L:o�.Q�q��6�D9� ND �!��0-PZ���ʅ
����Т�!�ĕ�GjLfB�Ut��qɅ�!�$=xޑ�a�: �r��6)���!�d�&@E��
Ԣ�F*h��P탄b�!�D�>|�t��$�Ux��<�!�d�F������'���ǂ���!�$)3��c��-Y4Re)G�N�/�!�]%o����ʰ*w6h`�R�y�!�$�?����ӛjZl}��`	J�!��͒Lŋ�̃{���@" ��8.!��LJV�P�b*��e��rr�̇%!�DÁZBJݲ�	�r���3��|�!�o���`$Z�t�0#� �!��4E@0�#���4#�aD�!�
'��4��([c`��+VN�a!򄛙R�&�3&�8nC�11�lS6rP!��VG;Pp��M�P*Z}��J1%�!��Ǟx	�B�3��*�jѵF�!�D[>Y��ģ���0FըQ��O�!�dNcs�HA`��� ���*�!�d %-���1&a  �0�RW��*U�!�Z�4�& ��LSX���g�<q�!�d:9<�5q��4v��y��Z?\�!�č��b{�M��	�R��фW%�!���}P� �`߇�4M(���G!򄀃=F$`%FP�d�8����ZIV!�A��� Ʈw�y �\%SS!�$������-�-a��7L����R�5�r�!mڹ�lI��y��֬P��D�!��}ɦ�9&ڗ�y
� �D�g�ʁgF` ���!j.�#�"O����Z�<M��$�UW��Y�"O�a����"'K� �C�<o6pI��"Of8{�C�>�j&�<`%pE�7"Oj��b�Ēx{�HE�]�5�Ekc"O�)���\&0�@8����2�`"Oz���ߋ�2��v��	� �r"O:����
)��|Z�#	Q�ؘU"O��q��#ҭ��E%Җh�2"O,���/�`����#�+)$ʬ�C"O���D� �TK���d`p�"O�)sW)��Z��#\K�l�"Oʴ�P�&�>�I��k�`���"OΉ+��ԇX���X�^]�~@BW"O��D�ϯU�����KW3v�� ¡"O����n7����٢#��	b&"Or`z _�
�xE�s��r��a"O���&-L���A��_1R%09"Ob<�'gq�0&j�1��I��"O5�$�B�E]�e*ѹK�}��"O&�xD
N�0i5d�xS��i�"Op�P"i_�1��0��P�'<L�5"OJ��t�V�H�� �%[��§"O�|ђi�"rHhׇ��pҐX�"Oа��C�$���ǔ$��u�0"O<���gÈP����2&�-�x�W"O����
�HO�Ar��W
)��iB"O*���ܧ|X��{��Ü)�X��"O��R%́�#��cg-��#�V�iD"O��qv��B�Ѻ�픛"�d�S"O
d�d&�6��X�M�d.�qW"O5rc�7>l5!���Ѵ(�"OH Z� ˕)��`+2%��[�t�"O��`��8��ph�a�z�Q
d"O������(���OR����"O*��uAH8^�~9��d	�\�R�"ON�"(�;��	t)�._�,5�"Oެ���3�j��'y�.�C3"O|��n�r~���`��;m`Z�@�"OB�+pD�>ڌh9�k^�r�z�""OD�[�N�7'��y��a�t�"O��*���k���U�/b	I6"OȰ!�f�,J�COQ_���V"ONI�S�ޟSs ����g��%"O8���K�{�������|�� �"O0TZ��H�sm����K����"O�%���()���F� 9�(d	P"Or(���f��]��Z�7�P�q"ON`��c�d�YC�k���*V"O]���H$"#j$��l�E�z"O8���ӎ{���I!0�d�a1"O�l�kȗcGb����kYr�qC"O֥�U"���Ait�X?�ũ�"O��{��ѯ2�@,	��̵P�0�"O�;���a�U�� ԛ=A� A@"O$XV�v�� 7�1|���	�"O�`�ǟvg�t�U �V��e1�"O������4C�,��(Ȱ	5�u��"O���#�X�{�����@�&y�D��"Oy#畑 ���'�D� \{ "O.Q�C�Q3
�� �wE�]1֕��"O�9 D_�"����]5x����"On\�g���p�L��N
��"O�FI
�phQ���
Ҥ��4"O� l!pa��	�d ����/��9�"O>�"�[:J�0�"��s��A�"Ox 4
�:|��1uDFb"O8�1�˞I���&��d�)�"O�n�*��Dh3I�����OժD�!��Ƞ@:ݙ�l�j���0��!��Je4���J55�Bu��D�!�ć�?Qr,�g��*�	`d�!�D��V�@кA��"*�j��D�!�dD���1,�!�F��UÁ�_�!�{G��6AN�/^Xj�!�H�!����@�Bd"\�f)`���4�!��V�j��M��-��`p�E/�!�$�L�Pq��C���=;�D�F�!�d��Y� ���
-'��I���P'Oޡ�d�$5�
�p��:}J�`Z�A��y��� i��S��O�]k��i Lӊ�y�Cݽ|#�K�,C�H�ɛ��V0�y(C�nhct䔤R�tH!d��)�y��]1�̀a�ڟ���
����y�%����9�ԥu����D �yb��r�ŋ�'o(D�5��-�y"'S���p�sJ|H���d7�yB�NFP��e�)<m��(�	�yRlZ�r�B6E���!�ϵ��4��'���@eD�1=�A+&Ɛ+lX���'�4��̗�xO޸be'�	r���'�^�J�V�9�rk�/�+�:Uq�'���QmѢG] �td�3
z��'�*B�@"�@�3JC%����'w���fȀP2<�B�+U��(�r�'t�����W�������Y��)q
�'^u;fE�9}�0�K"A�����'��	�n�?w����B��<C,�J�'����a�Т�F�5����'3���@�1��`"6��,&e4p��'��ԁ�Ɍh U��X3�Xx1�'ǾMA&���S�X!*����h
�'֌����+U8Ȑ�tO(u \0
�'�����.Km�D0�	^<t�X�	�'Bh%7��w�pT��9 �D��'p"����X&���#]&Q�;	�':�`E��q�<P6��C�
�
�'Ѹu`Qfխ	e�l��4�\�	�'a�})΄1l��A���W���\�	�'ox9��j�T|ma�\�_���'�x,���	
 W���b�� Pm��'J���e杹��,bả�f��i�'$�����6^����C&'���R�'{�E�biB�{�0��#���P�
�'�B\��c�%#� ujG�H4���@
�'�Ι*�@Z+L%�D!��-#�JiB	�'�xe����b�~l��-ƍ!�P��'"����L�e�h��2l�
eI�':Z��aش"*���e��j	�'l�idA�O���A�0$�i��'��4�P�	��+�F�#@*�@�'�D���Kj�^�"��Dh5��a�'JhH����L�Re[W⑴p����'Lb�"�	qF�]����#��Gy�<aw�'\��UrU'\-p���AFPt�<� ]�L��@��E���m�<�4��0�6i��[0ޘ��#�	f�<�2�����dE��)Nq��hM�<�+w�   �   �  ,  �  �  ,*  u1  	8  "?  eE  �K  �Q  /X  r^  �d  k  _q  �w  ~  W�  ��  ې  �  c�  ��  �  '�  ��  /�  ��  [�  �  J�  ��  A�  ��  ��  ��   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C�>����鞿6�!d��x�^��I��~�!��
�l����v���:�9a��:uZ!�L�,Ƞ�#g��UԀ�e��t�!��v.qc�ʁA�P{U�C-h�!�DD�x>B��cG;c�lK�,��"�ayR�	� Q2���F��u�t��� �/��C�I�Ld֘8����D��T�U�#�fO��=�~bh(e������M?��m���Tg�<� �������T�����R�g��dR"O���ѣi�A	�͖<|l��"O�ȁ�N��SO��µ'�#{u�L�"Oҕ�sGY�>u�0@�'B>]ԕ�b�'I�O 5j����)ɲV�л�"O"}��J]�P#JLa�׊R�Q�֓|��S���O��Ḡ/��l"�88�n�:!�D�	�'X���P��u�҅� D�l7�<��'{���6f-虡4��	.�<�R�'L�Q8�C d� ��욯zA��'a�l�3�F!C����4},0|ϓ�O�4 6g�'���z�h�!�P�R�"O�$Kue��Vrl��MΈӲX�S"O�!X$�ZD��z%��B����C"O:0���b�V�a@���VĪH��I8�\��׆pT����Y)i3	=D�$�&���;�#!a��9��H7D�|��BP���x� 脖~g�T�#5D�H��
�Kh��Fo�Z�s#�'D��)F�^��$H�/ǐ'��(#D�8�\�.V>���bYO�9�4m%D��3"�Pq�f�2P.p���(B��$K
~%x�b1Fb�la�CN�.��C䉮T��[#A�$I����(��AC�C��H�XtN)qH�!!��A��C�IHh,����s�6C K�R�jB�	����#塕��Z����}�B�ɥ~�� 2
?<�[�"��nZ�B�I)&�ĝ[uj	�%��a��;�hC�	�f�-� ���=��d�E۸a� B��;}�܉�e�1(��1��ġ=JB�I�!�\3�oԾ�p��C2h�C�	FxXz�g��dp�Հ	c�C䉇>�6���a9yVa�W�vdlC�	�!2,ҧ�?U�*�����5�0C� XwZp''�q�1c̀�ThfB�I(wM��+����k�I�@�ӽ	LB䉆���F^�=*Q�@GB�	�4�ܵ�!�� (Yv	`s��7�B�	?s�r��d����hj��I(8�C�	�g��d,�(M>�h�h��q��C�	�TTx�5��<�� ��&��C䉿[.� �� �a�P��/ԌV�tC�	3F�!wFY�b �'NV��C�	>=F�m�FǵxZ8U�ց�	tLC�ɦ:�p�n[�u�ҴY�!ӣd�BC�+;���U&�<b��T�@�����C�	<+A����Ǜ �R�I�.ݻs�C䉂Ԫc��T/T.nL���ܴS�B�	->�N�9�N��T]@xËZ�a��B�I�E�Ĭ1� ̮j��� A��'�B�I8[�2�r ͫ���TP�]`tB�$�0C$�!O�偷ƛpuNB��]EdP�o�4'��m
D�ُ9.2B�4$�t(*d�8X�}cRd�+DB䉷L�T���k�2n�i�CE�[SB�ISQji��6��{@��/'�C�	�sϴ�;u
�?�X�:b
��~/�C�I�F!*t��N�:�0�h�-	NzB��<�C��3}"%���CW@B��&`H�ܸ�Ζ)��p��+� .fC�	'�n�x�$t���2�I8�^C䉟2�F�@�╧Nt��q�ŪXtB�I15D�"� 0h},�H���yA�B�)� ��aF�H=�`z�aN�'b��v*O��xc���2�~�0����}��'���� 0����
Wl��*
�'��ԁH>pxcG�o�����'\za�2mF�3��H��ˀ%o�����?)��?����?���?���?Q�=�q���-xpB�ѧ�B�j��9��?i���?���?9��?a���?i�vD�U����;�Pĥ��?P����?A���?���?���?���?q��S�x�+��� &�h	���#OVlI���?���?���?���?���?��j�$X�գ���l�o�d����?a���?���?����?A���?��(b���[tu��+�B�h�J�2��?���?����?���?����?a�I$>�K�m�����Bl����?��?	��?���?i��?��,�lyGm�1��x����n��,���?��?���?���?����?��g�x˷EǂP�C���'�
�C��?����?I���?���?���?�7ⴹW)>��
A�������?	��?����?i��?����?��s��A�N &)*�n_�a ��0��?��?1���?I���?����?a����*��)[�|��� ��r�J��?Y��?���?���?y���?Q�z�(��P��
^CB�ve��A�Z)[��?	���?1��?)��?�c�iC��'�:�i�ƩQ+x��r-dԙt��<A�����0�4)�f����s�P�p��&�:�S�C{~��nӘ��s����9��S�Z�A�u�_�ƚ-��՟�R�(����'Z�	P�?�����uc2&MD+0�ѯs�du�����Of��h�d�Uk�19�A�v�R�q�2�a�����#1!#��L�'Ad��w1���G�[	7��%�ECN��xM9�'$�?O��S�')����4�yR���B�@T@��)T����pM��y�9O�����ў�ş�%�dȌ��#QV5���%`�L�'�'67��-�1O�0�vg��k��Lץ
�ؑ��/�����d�O���u���'|��Gw��Ȃu B�}{�O4�DK�1
>	���I.�?��H�O\�p�n߲iM�:Q�F�Bc�m ��<Y(O���s���$ޑ6��$ѳMyE��uOv�`�ٴX�t-�'f�7-+�i>�ꖉ Q2�8��Q�'�a���o� ��ß@�	�ED�n�q~�=�,��&c�<hJ��~KL,�&ş)���#�|V����p��џ�	џ�Rp�N
W,
��IV�LH*3��oy�u�mIB��Ot���O̓��d^��%D�8Gr��i���Hb�Ʃ<����M��'L�>���O�;5($s �� �h��MM�Kx�S� �>��@jhy`�ьO�ؖ'c(`�C� ��,��D�	H��'/��'�����S��ݴ`� 	�@F��	�/􁻂�D3`.d	�Z�����g}r�i� 	l��tK#�^�p� �G7Y~���D�Uo��m�^~�닥�ܠ��w�'ojk�3=� !e��!'2<)�+�T���O����O���O��$9��b�.Iy�$:?F ���>/�(���՟���9�M�$)Y���dNߦ�'����M��d�di6�ώBb�(CUFN:�ēM���Fu��	]YD�6�7?!g����(� 
����s���?�Jx�$��E�F�$������4���$�OX�$R)�e�5ᛧaU�l�FnUd�$�O�˓Z>��.M�\��'erZ>�05#�+$�����LDA�=�l)?�_���4 ��v
&�?]SGKE!F�:�tB��@¸��4u T0h�I3���|��`�ONd9L>9����IF��Q.2�Ψg�ކ�?a���?����?�|"*O�$o��Zm�U��h�r����L_!h��I�������I��Mc��B�<�4w���E픧��=9� S{$��sǿi��7mC0H+�7�??Ae힧����3��[�j�x���,Ү��qe\
�y�P�L��ܟ���˟(����ܕOΰ5���m��eg��$��XXmq�(x��-�O��d�O����dD٦睈B]�a���q#~-�
ӈh%ډ�	��
O<�|z��0�Ms�'�ص 7���NcHLp���A#��؟'��)�4Ǆş�$�|rW��S��k���FTn��"��6%�Rw�\�������	hy2�{�T�*�OF���O��.���P�C��Ii�r�Э8�����D�O�7��]�'e�:D�P�1R���i�d�	ǟ$#����2U#B|~��O2P��	�x���0'��(e�(ј	h4&ז�"�' �'E�����"�!�3����^�qo6`x3�C���4.G~�S.OBl�l�Ӽ#����Is�y	V�A<e�L��E�]�<���?��i0�a�ia�$�O���WJ���!*�v'z���n�4���2#�F�RUp�O���|����?����?����>4��D�5����LN2,.� )O�o��+�m��ȟ���X�Sȟ��G/�-?�н�d��Y�b�*�(C����I妹��4Sg�����O���H�3U8�UY�� Q�YggI*Ly EY��d�*\�n����*h��Of�(2��2�K�4�X�d��蚘���?	���?���|�+OzUm�
INL�ɺ/?� IRa�8:x(�cC+��H��	6�M#�2$�>��?׵i�\��R�*1ՎQ�G�N��Q3#7��:O`�d>Bf�Z��Vb�	�?��=� vmS��A%1TCV:l5t0s�4O���O6�D�O$���OZ�?ᘡ�.n�Ȉ�ɇ8�Z�#"��Ny��'_F6��+5�)�Or nW�	&P(vă����j�*@M<	���?�'hҰaش��d(<	��E�ϢiR�|
��G{J�#�C*�?�&�,�d�<ͧ�?a��?�U�O�"ߘ8{V�5i���Y�	�?!����������ٟ��I�� �Oh�I���.�J�*��6�&��Oܘ�'R�i��O�S'Y��YA`�<1B,�!!���t�Dy�eo�()ں�s�:?ͧZP��DH���bd��q!�M��1��ɮ�	���?i��?y�Ş��d�ͦ5q���$u��j���v_����+^5A�X��'��7�>�	���pӄ�b��;L��6ʍ[=���EOH��P�4*;r�4��$��X;~���'��5��]�5ɂC�5{��W"���Iuy��'�R�'���'��[>uP�Ɠ�e���QBOϫ�j���gۀ�M�Q�?a���?�H~j�v}��w�"𠱩�
,��(�EC�g�ԵSv�b�v�l��<ɪO1�0�1�}��ɡv�j����W�Jq�偄�qUd�	�js~q��'6H�&�����')n���J�X�����V.TEK��'��'m�Q��"�4h`Bs��?���'�N BT�O9z�*q��@V���i�B&�>Au�i��7�WC�ɤi��9:R�II!b��2
F���*�#ϟ�t�D�|�c��O�D��0��#�d@(5�pBvI�(]�
�c��?1��?���h���$Λ<�f��S�[�8s�Ao҉H���Ϧ�P�B��D��:�Mk��w�t�d��3[˸p�WlI��`�'F�6m�צ5�4}��`�ܴ��Y L�6 ��z�v-c���m��!�@�~���cB7�Ľ<ͧ�?a���?9��?���1]lM)eeA�S3���r�U���dW��M"q�ןX�	ڟ�&?�I2de<��4�E_@�y���إ
��IY.O~�Dr�>]$���[�Ş_4�ځ��o�(M�wӄ#��!���\����B��f�	cy�
�nH����K$t��Y@��f���'zR�'��OL�ɪ�?AE����@g�ż'�� Y��'g�@H  ϟ�a�4��'����?���fk�QθZ�K[vhrYyA-V�2�h��iH��e�X����O�q�d�N�& S�b�ײ�0�����Z>��O&�d�O����OP�d1��R�L0B��7�^	���->t2��'$�ix������?�j�4��7����N�.6�6�`F���\0�x��'��O �Ҥ�i��I	T�{��&L&�`��ǌo�� �p�ؿvn2"Lf�	y�Ob�'�Ɍ�J�4�A()8[P�ԗ���')�ɮ�M{����?A��?9-���(��Ģ|.��S�D�	���8ѐ���/Ot�$g�\$&�ʧ�"�c�X�n-�HA��:G�2�#��D�$�N���"}~�OT��I#z(�'���3V��VT�[r�ϊsjV��V�'sR�'�����O��	��M�1%KmȾ� #Z/��
�!��zF���.OT�l�`��/�Iݟ�w��	[��ٛ!ǆ�}�\E
\🸠�43�pڴ����H��Ÿ����+Z>�$��2�r�U�1�D�	my2�'���'���'��X>�WDF3Ӕ$��,%s@]A����MK����?���?�K~�F!��w�h9c�[	T�V��W!�_wZ����'�2)%��)��+��6k�� ���M�p�!�'аC��б�$r�����#|B�H]�\y�O��Dؼ�p���f��سQ�Y�4��'���'3剸�M���I��?���?�sd��l<dK�C��L�2`C�����'��ꓬ?I��H��'V�Hq*��Z�,ʳ��)+:(	(�O4�ٖ��(J P:`�IN��?`��OF)x$$�3���Ԥ�<�l�`&��O����O*�D�O6�}:��4&Te*��4k�t��0FS!{GR�(��K��f�ɸB�'�J6m3�i޵����u;����$þ���i�j��������;ش�R1޴����(oȤ�'|�8��6?��H���9$i��*v�7���<ͧ�?���?���?���=|&�u�aE�L��%9uFY����Ӧ�1
	�,�	���'?牝T�d-��!V1b(�3���>�P�S�O:�mZ1�M��x��t���k�$	׆��l?�0Y%ˀ��T�aH����Q0�����!"ؒO��.Ɋpk�@��#J�����|���H���?����?��|�/O�oq@v|�I�E
j�!�J�� �VA��ɺ�M3���>����?���i'H����?U�zh!π�(�S2aWd������lA�S!������ld�Beǡ�썣+��H�B4Ot���Op���O�d�O��?���E�`�8����U�3
d��b�Gϟl�I�d�ٴfy ��'�?��i[�'&黳��-������
�i2O�W웦�q��\|6�+?q�ȆD�ШB���3#7�#�윀r���H�O�9;J>�-O��O��d�OĽ `�����)��� ��E�g��OJ�ĩ<�'�i���<��柠�Oz��(�	�H�Ĥ� d�zX��O���'k|6MS��i�S��du�|B�I�Z��"�F6Q��	V'uSB�RS_!��4�P����ָ'?2�h��M�8�h�A�.x��	�'�^Dt�/ƺڂ� ?tI�	�S�~�-Дh"q�A��Q=�P
�e��5<��@�쟃�С��B�ncn���@NR�iX@���HvgĐd<��6错;� Q3�O�R�\� ��e��oP�yh�͹pT<"�̟E�V�Q�'��0��̛���4/���H�B ��A!"��*��Ap�,�8���f��[���,o��kf"O��g�F8�(0_XeX��S���pT&I�c��'v��f�7��ݫd�L�y �E8F�F��q�Ȳ ��k�� ��D�F�[�|��`�`�����N"r��4���Ŭ<a>�F��e�A�!��F|-�FDN&aI?:<z8H!E�bXlaH���-H(5*��.$���%"�K$�� �c�O\uP��� >�6q"D�K�9C6�9Å�O��d�O�,�@:Jy�nW���y[�IG��������X��#E�k���Jg��)�(O�<s��*�� �	�Y�"+$�r���T<E ���9P��a�'Ot�'r�D����?�O~����t�z�c^���´c�:��$K�����?E��'��	�-��`8��`��,�>`����'�'�����
Roâ:�&����O���D��P䊦o�m�R Y`+'4!��թ	<��!�1Bz<�ꡨǽ4!�C&��A��;W Q�pHߋz�!�$�2��|�Df��| ��J�AH�Z�!�d9�Z=K���bg��%��br!�$g��e��m�� L�9�4BƃXh!�$Y�f�T-�5���B�XZt�@�y�!��i���`1�Q�T��
C���,y!�T�{V��%/���P]PP��H!�D�7Ul�@���h����Lև!!�䕘6��B��Q�چс�AJ�r�!��4 Vl�$J(P�x;6�)=�!�ě�a�H�8P�%�9��$�x?!�d�/&�b�F���l��S7@�!��+ێ�(�NA�+"*Q�� �2r�!�d�Q��"U#H�a:(PoZ:9!�$D6~=�UJE�N% Q��՟;!�6NS*���	� �'�n�!�$T�r�p�ra@A���u�<&!�DQ�.o
��'�Z#'���׉�2�!��� �@��A
B9��-Q��|�!�$D<��y	d"F�b�^1"�m՘x�!򤃪q54����YXX��l��r!�ĝ�[�6��GBY��{�K b!�DZ%�X��_�8�x@�%��uK!���*N����(����cӶ28!�"z��Lyˎ��jd��O�_L!��?-h�D� [5G���V!�䃠��(z�SN
}S�f)R!�ď�{��S�'߳7J���Q�T M!�&>�$����
n*�U��O[d!��s�<�)��?t�l�ir��RL!�){z���n�;u�>��Z~�!�$M�17[Q��E��yұ�л�!��g�A��{��I�V�z 衇ȓL��air�O�E���Ƃ�4`�괆ȓJ=�!�*w�x)�JB�d��"O��bR!JZ��݁B%��g}t�KT"Ov����&��)���)���z�"Oh�wM�0�p!��u���(r"OL!	R@>R��a��f١��R�"OvL�7K�e0�����ߘXՊ�s�"O��%� =hV��U�nӪ�2�"O�}x���ј�cW�W�N�V��$"OR�ă��3`ٰ��W�N]�a"O�Ps��ϻT
�#
6`��m�V"O:ԃ0-� &���cJ���[�"Obm��a������#��BGJ�k4!�D��N;��h���)eF��b�>!�d�#"^ �B�B�B �͠���EG!�l���k��W�H̢I�'d�>?!�D��Ji`��Q\�,�QB�?.�!��C7'�8.)v`m�7IM6 ������ i!C$µu�p�n�30���"O��A�a[�F,,l�-C&�nyx"OB�0d��2HL�x3���eې�"O&M f�G0
8���.I�bl�q"O�xcGE�X$A��+�|�"O�ѣ�FG����Q�N-SC�q�"O�B"��@=�H!W#�+vEp"O~���X61���g_�"l��T"O�8I2�й_Z ���'˥����"O��Zu�h�挠��� LN-J"O:��чѧD�9�4i�#7�t��g"O>��C	}_26'Y�<%R�94"O��B��������ܪR��A�"OL���"�=p',ac�Ϗw.c�"O��!��8M�H��/#����"OR,ٗ�qIr��:E~0U��"O�+��"���bg�'5{�LJ�"O����n�S��qq�JE�MD��T"O��
'� 
�Xx)C%'�UI�"O�p���*3`�9Վ��.�Pl��"OD8���܇pI�`9�&��T��*�"O��Y�,���N��e/�g"O�yg"�/v�$�H�#]�*,d��"O|��p�Z�1!i�R��A>�y�"O(	榓�]3&�+rb82�"O��sVk� j�M��K^�K�j��u"O��!��r'��:3Ii����"O���Ǘz�A��s�^(�"O����o"*469 G�HXŪ��C"Oĭj�DI+!����'+�=�S"O���0��zڂ�Y��Y`�y"O�!���>^��)UD�_\]P�"Ob]��HV�+�\y�RC�]�։)"O
�fE$ }B�Ŧe���"�"O���5�V�?�,����Xئ�	 "O��2��������#��9��"O$)ht+�0Vs!���'=���A"OVy@oϦb$ ����A���"O�E�N�`� BfݿK�zE �"OP�A�'8Z�����	�$;PLB�"Oބ2��ԌPW�p8������"O��� �]�%�X�* (V!�@��D"OLb׹�V�ز@��*_�P��t�<A%���}{�ms����"i�4�]G�<9�/�2q���K_=b)x �fQo�<1�4a����ڒ!|�4��Q�<�LT�P,h�!bU�P�:�[��q�<	�	.XP�S��ňb�y�"��q�<a��ݒr�&)X��
�d��f�[l�<�I�7 :fa�k�8���ʑA�<���6N��Q�g��V}�`�+�{}�Rx��	���)a��FF�_�����%8�O������<�N�LѤ0�&mj+1�o�<qS�D�;	�-�DI�D@h(0�KZC�'�rHi�0�k�uc2�1*=
��� �2���O�����G��d$}�ek�.����N�i��O?�ɝDB%�� I(�:X�R�2"�JC�r�($K����
�2#/�0J�$��I�D;�@��$��#��lx��b�ߣRt�Ň�&v<�p���A	��$�\4 ���O���b�(@)*�!�92A�Ѹ'�J�D>�Hr�'IH��'��Ip�/Y!*��E��Oƃ��<ȶC �@=��D\��yr˔;1l`5��D�zH���jS�W7L��&�ņR/>�ZmE#)�M-F��é��9�����S�? ���Q��
/3j80�(�7 rg�i�JX�mV-ǰ>���(�$ً��:O���x�@K؞�Q�aǵR/p ��$��z����Dd~)b����w/v���S����c
�(�b��iH8EDx�	׃H&�����T�9�lyU �4;Sn�b��E�T!�䄑(�� ���L�H��+�l�N��b�/ �' �>���8�pv��~��(�c��*Z�zB�ɜ+~J���Ϩ]�]�Q��(BP6�_�`zZ��R�lCP`\2H�8���I@��%q�$?lO"1K ��d���~h}�1��0��q����7�^��ȓ�$�s��JzX)� -2B���?�AN�Z��H��I֜4�ԑ7'Z�M��L!�Cě�!�d�%/ND�,�$�l��C������թH��b�"~nZ��ҴB6��a�
	+�n�vC�	��`��=%^� ��j�L�@��+��'��xb��U6W�B�`��IM��u1�D\�d0OD���64����*5���r"O�-��/�;l�����!4�)��	�dm���):>@\�a�܄0��IBᏑOb!���u�<�&��?A���z��׬]�����p�=E��4�p�C�\H�I:��N:;�&��s/�x�ph	�K�E�G@]�#�U�'��[D!��=�0�ӗ:=zr�- ;���c�JX������u��6m�p�\��E.k~X��K��^�!��,&I<tXf뚾H��@�d�Iq��H�Ee�D��>���!��Rq�TKc��D�e�*D�<�U�76���ӵ�!.l�`a��tӪ���
LK�S��MKCE�4cBᲖ�l��)Q�Cg�<��Ы-�E #�^�^	�`�g�WN}r$(a6���d��U2QТM�8X@=z���)~4a}��3<��I.���e�Q� ����G;6B�<3ꜰ0&EG	:�i{�Oq�"=�!L�)�?�"�D�.@1C[�t֒��<D��I��J�5�<��Z�G�8T�C�d�4\����w�S��Ms�F	����B�_.Q�Xm���[�<I���-Sr��{ �. ��f�Uy2��p>yA�\�V<��KթH'9bA`D�PN�<iDh�c���#��L0lJ�UN�<A�nX�����*	(�}���J�<yG���'Lx�D�E|�lp@�_E�<�5bz����!b��{�����[�<����m�V)*hj(�S��S�<�Qn��6����'ԦN��Kf��L�<y�Ē�7��r�*�96�飰��l�<�`�ƨ!��I�愜��A�Ġi�<Ap���/�:���J\��xp��l�<�ҦȂ[F����	-[<�ي1̇e�<��f�l͚l8c���j¦?�B�	�nw���#�Y4U�2aCj�i��B�I3&�I$,
�-P���_�`&�C��8c2R��E��x���T!�C��0,-��ȿ4i�ZV�Y0`zC�Aih�@�G��BU���=@C�ɑ*`(�j>>Lr��?��B�I� p���+9�d�x�N�a�B�I��h�;��E<� ��&L��Y�6C�ɷ������( �I�C�	*n͸���e�	^&3C䉁?�b�r�o<!���� 7)לC�	�Yޚy�FK3e�l�h��`��B�I�i8��W�5=���;��B�I�U��Y�v�?A���HԤ��L�\B��`���JgIka4�Ǒ_!X"/$D��� �ϠVbR�gL@%Yܼ���/D��  ��nR5W$V�b��b.Љ��"O���a17U4 �0́�S%�	��"OPi��jY�W�<�d,�?~ZI�Q"O�`�-Ϟ �R��g+�5�@��"Ob4z�,I�U��4
�)Z�3@"OXM�1��X%Z��6� K�l�s�"O��ƒ3>�
���a��I�:��'"Ov$ ��2j���f(s���R�"O��Y�,ʙ�
,1�%�YkX�F"O ��'/̀���CϩR~i�#"O�Yڄ�ޘ\&�\Ygτ' ��sP"O&ܰ�
5Y]\��c"0�&@J*O�S������sV�1�`S�'��񩠄�3�1U���K��XJ�'A��0�*W<@� ���ِ@ 4�
�'ۆ�RO�1`����OH;᎘r
�'BYʴ���V������I,8�ƝS�'�^գr�[�k��Ea��ڢ&@��'�ڙ�D�2<���ϳ~2�!��'����F֟N�,�AY���K�'�R�!B��YD�k�i8~�V�C�'5�y���΂2��ᓢ�Vs1z���'[zDZ*��z49��4l��@P�'چ��g�#+VX�q�[�d����'m
�A�#�~Y�P��,1��`�'W���OA�J|h"��<�x��'͒�R�f 6'Yb��`Ç ���'%��IEOQ������V&��'Ȣ��g �4b8�	�	��}Q<���'8�����'�� J� ��@��X�'#�]s���|��Q�eEm�X=k�'�h̹!a�ڎ�C$�� TT�':���ʃ��,z�i�)i&���'�8��w	�>lܴ�C���̴��'�P\�e-JBg&�h�]:!����
�'�z%�S-S�H����s�ܸ
�'�2�Fn��'�&9�v� .�ab�'-�)S�N�Q�;A��-l�έ��'-´Ҷ�N.@�q`#�ؘ\��\3�'�q+���S�9+��T"?3\���'+n��iNb����8��(C�')�xpi_H�\�h�JP�/a ec�'
,� gV3A{&����(�$�Q�'5���˖8�vDQe�-ml��Y�'�8���"L�``Q�
�����'��2&�Y�2��{B�]�;p��'o���@�6!iQ����*���y	�'���b�# ,M�I0�����I	�'4Zy�AOP*L!z�C��N+9æ��'<�:6�TE u�&��
i�	�':�(g�B! ���R)�]!Ԣ	�'�"I����첢k�,�F���'ў��f�46A�[�&���j
�'A�8*gC�Vݦu
�ψ4#�<z
�',)��	(%)�(���t�9�	�'��XC��O�>	zU�O�X�`S�'$��23H�x��q�����v�����'�xY �#�+�"itO�$�@	��'V�]3�EE���������'���{��& �������"�A:�'�v�9r�
c`�0K����;�' p�AAǌM$��06G�=Z�'����`�pE��b�ŋ�'���	�'$e˓�S�i��%*�iZ���}���� I�F��&v�"�R�P#
�[�"Oj��nC��X�Q-D,u6Mp�"O��V�&���;����"O��R�l�b� ���#h����P"OԚTm�)=�@��bQ������"OP\��&�	]������L�$�D"OV="u��BRx��qC� �����"O ���aֵ���K!�Y�?��Ԛ�"O�@� �ʍRQ��yCAʎ�ĸ�"O�5Xp��_���Q͕�K��ՙ2"O�8��&ڋ��	P���cܤ`��"OJ���gUHD��p��Ы}��X��"O\���])X��-��c�F*a$"O����7
NLm* �_�/�(p1�"O:�!�'vH���l�(V,�4"O,���ۈ	5�pr�˅Mv,��B"O6�K�ʚ20[�l�-ɚG^�l:"O
@1�LD
J��h�U�R�ոd"O�9B��O��KӬ�&8Jص"O�=���L6D�B�"�N5����"Oܘ�@ ��P�N�"F�S"O�l�0N�"��9����I�1��"O$�s�@9jEBT�@�r!^���"OD�r%(T!Cv`u��hs����"O���H�r���P&�V1'�fi�&"O�a�Q��!zZLD��ǈ�A߾��"O|$��K8=�d���۔a���"O�	�#F�h׋�iqL��G"O���piX�R2�I�kÂ>il�0�"O$)Iq���!�/�CGt�JV"O�%#ծM�mBdXc��Qb����"OFk��N�WP� I`�/O�̊�"O��;p'�r�0(ʣ�
 ?@�p�"O��@L�"Q2�[�14��p"O�;3L��(�����:@�y�!"O(x�b��!%��l��0�y�r"O@�5圐i�<���L�;:VFA�P"O"��Sn��`((m	;<h, �"O���af�g�Эj��J�Y"l�"�"O�hT�\10Ą�ɂ��+#"O�l��0W$I�E��P2�"O��t��@�R�3���(��J"O���jLo-������74�,C�"OF(�UGaJX�!Ƣ�C�]r"O��YR�F6�
�i��B(�fd��"OB���cT4(��e9��9æ�w"O�Y.�1%��b"%D�N�Ľv"O���Ǝe�����CM'��H;P"O�i@��Ff��$BɳC�����"ON��ો�V��a2���T�Bh@�"Ot؄��W�yC������"OB�[�d�0 ;�92 �D�g�%��"O�2ri�I��i���oؔ�""O�i
�_��+��@� �|�jW"O
�{&�P1����V��
�0��"O�M	6#�*�N`0��2;�,�!"OtQ�Z/�6����
�Ŗ� �"O&�`1"��.i�gh6�fe) "ON��e�F'U�.�7�¨B��P�6"O������X͊5
C*Řw�40xP"Om9��+�Ui0�_�R�8��s"Of9SV(���-�!� |�"O��*d���P����qm�r��s"O�����4Pz,�r�oΌ��"O� �H���[�^��R�ΎF�!3W"O��Ѧ�;&�
�ٳ�(�����"O�́���P�����b�$�i4"OZd  ���&�9�����F"O��Z5t� ��۵62���"O~���'�uN�� Ê2M0�)�t�'��D��(��h�$ �O�r�=�ȓ;�$	aTd�V�4�PR�6��	��y�Z!�ܬ#R��R��?4"�}�ȓA�ָ-9 a���]�H����aJ4D��u%;\E:��CA]��-c�*O A�T���X�n���n�{���D"O��#6A�JNԥ�$`	�Iѐ��r"O��@���1��(q"�;V'��ا"Oj�:" �>e"͐�A�u
� ��"O�l�r#ʴ<�L1b�<_�	�"Oh	�I:6<f-i㠎�;��u�"O�-�T�Oo�i�f�Y����S"O|ܢ�ˌ5�~��u�ژf�e""O
pA���T�p ���6"O�����K�AA���dR�0g"O�����.���#�N]��r0�W"OFU���&�~�K�B�~Э��"O`T� �B�q �C�CK�"O�T+3)��|�U"M8[��-Y�"ON����.EcDq�
B��d��"O�0儋�R�TÁe�p�ޭS�"O� ;���f�$� ���c���X�"O$H�C��A��U�BM��/N�T�"OJ91$ܤ	��X�ۿD8�x�"O4P9'k�G�������MJN�`"O�IiFg�;D��d�`G�}��"O��@��Ne�%"ǡU
M�*D�Q"O����B����a�����w"O��" = L�Kp/E20��"OVԓ�I�|P�=�)_�Q��"O����Ίd�� TB
:fni�"Oֵ����@�^̸g�@��h"O���CBT�M� �����"O�!�MX-P�fPr�^]�k�"O���D-2rc�V��T��"O��k\/���
�k �5Kd"O��a$��>ܡ���%T��"O�q��b�b�nm�w�[B�4��"ODmQ
������� Q
�I�"Oڬ��@V.`���
T�9�I�@"O��9��\[&@��R�T�D"O^�y�]�+@��A�;Y�0�B"O($�#շqæt���܇��y��"O2aԩ9� 8��BÑ �~���"O���a��Da:�h�n~���D"OxB2��!@������"nl,y�"O� ��n'A|&�BP��P_\�rS"O��>y�bG_>S"��"O*@q"I�l3���#��?I�#"O���R���`��	�m�F��"O��	��̑�nА�핳M5*$�"O����ڦR@m��˕Y n��"O8��`I/M����*��jT@$"O�1�E��d	�
4�J,W�H�+3"Op�P�ˬ�ܘh&��&>�(��"OP�Zq	�Sb;�抣e6&�U"On��g�K�j�BE�P��7��J"O&��螂(�J@/���p���"O� �s���v�F��4�i�<�cD"O�I�$�!0��Q�#G݄}�&�#"OQP#֑��y;�^��:�h"O��[���d}Ԕ��>,$��5"OB):_2L�!��_!:>�0i�]��yr�4͈U����(�l�w�Z?�y��@ld��0拷�쩓VjP�y`����Ҽo��정��$3��	�ȓ"B���R�%"�H���L���ȓ,{r`�3����t`X��_8��ȓ��@cA� �X�w��;�l��ȓdx]p%�C�uH 8�I�b�х� ߆0;AGQ�t�:t҂*R�B����5Z'AV�&d����K7Ji�ȓ˰!�IW��l�Qj7�^Ɇ�b�D�l�!((�֤\
��ȓc��U@�G�t����T�$���m�(!��$C �L��%��(�9�ȓ.�T������`)������ȓ��S�gU9��H�&��[�x�ȓ6̨�cង���Q7-�k}4���POZW�6)F ���F)xp"O���D)BtH��aID�� �q�"O����k�Z	��u)�#j稬82"OR�y�F%S����t� ���"O��p�=c1���ǈ�^����"O޼��-*�� ҡ���\���"OZ���ָU�^�� �ȟ(��͊�"O䰊$j@.K� �ׅ�$�|��"OD�Dm��U��d�#�0�w"O\�`'L��{H�Y�գ�?�Q�"On�Q��؂Y$<�h���;:mA�"Oq�3����}��- �"O~�	@����Lb G�*e~l��3"O���rd�D �{@�P�� P"O*A��OȥoX:�"Q3���C�"O�J�r�X�2�O�����"O$$c��_9>T@��:��4��"O�=��qk������ 8/L�Z"OF��Q�.~�6�!WԌ9(ܼ:a"O&%!����|M"lJD�ۦ$P�T"OjĩE$.A���ظL��|�@"OT|��9MR�b"c��E=L�+�"O�H�񮓯6��H��E;̹B"O�@1�ޚ(��9@,�S'N5��"O���e�9F�ܤS�JX"^�ٻa*O�Y1T	�Kba
���}��y)	�'w�Tѣ�D?8]ڭ�S��<�ޑ��'f"�Ig/њtb-1$E�np\m�
�'&��s ��#w(�f�S�_���	�'d���cԋA��j60T7	C	�'.�C֕B٢������FrB		�'����.�2�r�dK.>���Q�'����6Nͮw�x���S%v��2�'b �����)A��a�NIG�)��'ly�%�ͅs줼S�n�	b�8�'����*)����+�$K	z@��'���H�+�.��8 TI��B6!q�'��@�+<7\��-%A(,E{�'���q�œ?BG����8����'���#��ݵ{�H=+p�X�B���x�'���@�u)���@΃DJ�q�'�j�!C�yG�a[�셞B�ȩ��'���@�ɢL�QcQ\B���S��� �E�$D�yj`�Bc��(xx��{T"OX��a��=3>�)��R!No(��"O@�x��2������MW�@��"O��[�Cѡ}@Uk�$n>T�"O�l@�O��P�����vak "OH��V�c,�c��h��y�"O�CP��c��4�;#���`�"OD���R9"nB��w떈Y|:8�&"O�b�������Z` x�e"O�a2���Y�T�CҨ�!ET��3"O����\����-h1��b�"O�d��	�.�dd�m�
�*p"O�`����tۤ-&�C
�����"O�}���8<pAx ��F�D�6"O440��]3C� GD��3�|�5"O�����DIP��`��d"O��YW��l�a�T�.�xYې"O�����T	�e�3��&\Tlp¥"O4��ꃪn��@�B�F����"O�-�r�W�4������K	1^��z�"O|(�fm��V�6AW�0%4�%"O�R3������!ǰxӈE�c"O������
�z�ՠ�&�F�#"Oj�bs� U�x��o�~��x��"O,�"���>@�$����� ~~e+"O�9�^:(�b�Va3zY��#�"Ob 3eτ�	� a�t�<K$(qQ"O���p K7Z��H�5C��2DT"O��� �E�_R���X6{���X4"OP�+�j]3X*
�`��3��4��"Oh�i]�M���WFP�q�d��"O��B*�)�\�H�l�hH�"O��fhϮ*>,p� <am�5p�"OʱӅ�V'i��J�O�_V�T �"O����2Z|�K � �[�@ �""O2�SƬ�I��`��O�O����7"OfL�UB�%Q�:@1�b@�+����s"O�	*�MVj�q��׋j�޴�@"O�=�e� b��1���_����"O�=��,�%�
�C͂�_��1c"Ot�@`�H���Dk�
�Y""O!12��{����I�y�8��"Or�b�F'uK��qۓh s4��ȓk�����7x���9dN�r
&$�ȓ@)��pm�;���%�г.;~��ȓjhm9�HU�D��Ap�/T��8��ȓr<���ä��F��Y�`e�zهȓ/0��sa�Ia�Qn;ꅇ�&4��(7&M@�	qe�M2*$ҽ��|��}�G��&�z)���O�*��ȓ����9-�)�RŖ=E�r�ȓi�J����o�й�A� �g$��ȓ<$��b��3?`ģ���2#EDՄȓN�B�[��+"��}SU�׬��ȓCe�[G�:]]6�9�_�c\|����BcO�>etT9j���!UVh��#3UA�#�63^<4�H��ȓj��<��@7/8��i��Zk�����a����1LB�m�#$��-f�`������2���`k�9����Ĥ��z"���.а*u���AB������W�L�z�MĆ\ڂ))�-P<Gt��ȓ�����Ȝ�7D�u���� ��@rL3�O	�)�,����Z�D����S�? �4�El^%��1�5�K�
���e"Ojt�7A�3W�<��!�;z�Ѳ"OJ��'B\��i11*�2K��"&"O6�k(^��lC�iY�wH��y��E�D���K�V�"�1D�·�y2N_�B�L(�í[G�,ȓ�'�yR�0�p���DU.	|d&A���yR���P�z�z&�S"}�r�b堆�y".�v��Hۧ�ֺa�]sD@G]�<�al2�ꈚ���.)�]ҥ�}�<�h̰/A��/��p׊��W��a�<���U��h�G�	�t���5��t�<�j�=~J\,�A�Ğ�j4�Wlp�<�d瞽"��#R�v`���p�<�Uf�.>0�B�6^܉�NS�<)`L���z`�Γ[(L�+�Q�<a��	��lɷ%�n0���`NO�<y3�M�i��h塌����eEO�<!�Ay��8���?M�;a!s�<!S!eȆ3���2u�EH�<q#�'LCT�PSU�|�l9��N@�<�VO��ZTȄc�~8Șb��u�<�E�j�����z��0t��t�<᳉S�W��D���]�B=���m�<PB�']Vii�eƉ)�d��c�<Q%1Z����^�t�����A	E�<�w� )�x�	���`*�H�d��e�<�&S2��8ɐkK��4hRi^�<��@��N�t�Cϖ�f4(A�$S�<yeK�Jn6e�o��a�N5��*�t�<�sg�=c�`�'��c�=a�o�<�%�3y�*-�Dτ�6����#��l�<��-C�>Q�JX�n��]�3 �s�<�ӌ�#�P� ��I�tlj�kHU�<a�Ӽp�ذ+��@�1�萫Ӂ�M�<A���O���DD^�v���e�o�<��i%~.�`�ǋ�4{bPk���g�<�v�G8ze:�b���h_^�(�_I�<I���8Z!�ѤX�`+n8xdF�<�P�Q��2����M/��1��-VI�<�nƌ&����큈G� @�Z}�<�7���`9��ˡfQ0+ʰS%B�{�<�1o�D�U�s���P9�9{�k�v�<A�I��8hZh�$��X̮���)WX�<1RK��l���Z2�K�̈���Q�<�⋕{����U��c�:9���U�<y҄�=th�!j�fW��F�`4D�O�<�W�P$b$ք^����aV�^I�<�7�G�*�<0a)�)pnY�BO�D�<��I�6j8t��3J�2�����@�<�3�Bj�zͲ����*M��Dh�~�<)6�" �V��"-ON�!�À|�<YSN�>�V��	ؐ`5>�q�kSz�<��(X�Kyl��ve�"�F�+��vx���'LD+1B���a2U��i��d%O���u�~R�"�ܞ����"O ���A[>��X`�DK�{�La��"O�A7C��}�D���D	U�� ��"Ol��� o|����B�R�|T@�"OВ���3ZJ�h���7x�x��"O&��m��c&Nb�� �"O� 8��� (j�|Ç䒽pC�d(�"O�P)�l\��J��7ߠf���8S"O�,���!���a��3 �LI�"O� ��*w`з,�Ā:�D}�
���"O����Nɼl�������E��S0"O��b OԿ4���a��܆&��9��"O��p� �w[�`��fҼS��=��"O����I��$	h%�랖D~���%"O|�X� ΰZ�� �C
jN؂7"O�9�
S=k����d*�Ch�|P�"On�y���3B�P�Hu��}(��"O~���)œx�.q[�	E�m�"OY8��	,J��PfߋX�e��"O�u��H�(��a�ܳ��("O(�!�&�6�3$�0i�؀��"O����$\���t���;�"O8�ã�+|�L�*���g�2�
�"O@a�vHc|�dC3��|�h�S "O���6![�g삡�$�&���"O���'D_� �WD0A!��z�"OD8�1�Q�!,�TB�$<�L��"O,��^�K��L8�&O�B�09"O~i0D�"�ZX�ͬ%��$�w"Oj�R�k_�
]y��X�U��0�"O��R��9x�t���mI!I���U"ONA[%iEo��t����F�0e�t"O��4��uD��	8*�Ќ+�"O8xp�G�^��uږ�\#�*�J�"O�<kQ�ǒ&����A.^����"O��@4�Z41F��p@R P ]� "O�0J�$��f*T�ϓ.Cab�S"Oz�P��� wΪ��mΝ����"O����ʰ;2�ē��I�߼�1�"O
0��D�5��������c0`��"O���g�dNԴ	0��F'D|�"O��C'��su"�B�Ȑ>E�}���D(LO�YQ#@�	R`���OL�~��pI2"O����\3$I�yXh�f"O>�86��L��xKfΔ�_Z ��"O��p��||<���9iC~�S�"O4��I��"$��l�>O*��� "O21�P(8�rt�LҰ5z�A"O��A"�Y�T��@ ��-qX@Qw"O����홻%�Α)�(�̄$#"O�	� � �BZ�g��d%
�"O�Y�
�8b`XR�o����!��"Oꉺ���BC:IN���uH��|�!�$���`u����={B�h:���!��ğ��q�.T".�=��'_vz�y��'�1O��p�� /�U�5�?pQ���"O,�**��l# �85�I�(J�k'"O�d�D�m7p�����O=D�)g"ODLi��ЗA��UJ�8_�ԡ �"O􈈆!�@�V�����y��"O�LS��J]b���f�lp��I�"O�Jq	�.i�r�`��n=�I矰�	çrwR�Z�!�i[���G"Ht�ȓ]T���\�"�T%#�E]�^h��*�~%��H1DD�q�Ӌ���ȓ?���TJ(
�.�Ag��+�ʐ�ȓI&���C+|���x�$ɉ�p��ȓC@`R��}�"�
 �̯J`��ȓIW��7�LY-��{SL�@�0��NNl�j��2G��	q!I �t��Wԍ���?ٴ4`�%��!��ȓt��k�cUv���OU0�z���}oj�"�拍��S��Lc/Ć�S�? l��5�\?�!J`HYgܽ�"O>% �b|���  IN��"O.���п7҄�SL[8 />�q&"Ox%A�#κ'e�]��N.X&�m�"O0GD�.�t}hւ,X�+�"O< �s�W)�جw��k`b��'"Ou2�o[�\�D)�gU
\U�� "O�Hx�ϋ!V�N�B2G^�{��v"O� R�c��{��P��&U4��"OƝ٠"U,I@ �PB1n+���s"O�����	/6�;�B	_"|��"O��U��,�	إ��9�T�0"O`�S �Bs8���DJA(�"O�e���B�m��|��@�y�n��w"O:�����
.����!J�ē5"O�TA���$�|�*BׄAН�"O��ub�R0�};�@C'�b��"Ov`"�,C�h���@���Je��T"O�<If���%0$X,W�`�)�"O�y{�/�Nr��A<y��t��"OTH���=�l�ʦ8���z`"O�����%�Z� >9ҒU�g"O>�Z�Ǝ�W��@���:�B�2B"O�q�5�[
~�l�o��a�i�"O�P�ii�J��-�t��I��"O2�b��]t��X���M�W"O�6�P�k���z� � h�~���"O�d(	??aDٳ�P>Y�>a��"O��X���(�lh��،s����"O&�vI`; ���"ĥy>�m�"O\����[��<��!ޮN/0��%"Ot�4�/}t�z�� W�HI�4"Ota�s@͔=R�	Ǭ˨#�$�j�"O:�q�횋P�E�ԋO�S5V���"O�t�����Q8�%`*O b���"O��kM��0���2S��0la�|��"O�9J	޷T�
���ac�i��"O
��e��G�ةq���2va\T�"O�Lx�N%t�D0#�֚"�(�"O�,�C�0����b�,I���"O<�āU�A'0�:Adçy�`��p"O2�aɂ�^��[f۷NYf�i�"OȰ��$O�<ĔAS���-��u�g"O�,�B�)�2R#�.��hiw"O�������)�7�U5-��Å\�T�IK�S�O��\@� dB��qgX@+.%`�'���`��оRi�8Х,�=�2uK�'6�=b Nؒh�E��O@��;�'C��bBN�T����\i�'����,�Z����#M��6ܢ�'5����A�.7ɰycE h�|8�'�RAGӏނ	�2�ŚtQ��Z/O@��)�)ʧ�B���ΧYT�\���]1�\��`�L�¢
*(�)��#!�\����Ar&K>C�f0Ɂ��8a��ȓ2�(9w�D3mvI�]�UxL��ȓ7��X�e�.����3O�J�d��ȓ 醨��))}�� b�#4�ȓ|d
2�ġ:L\d�t#�$t��a�����1Vz�@ �I�g;�|�� ���j����Z�.�#���)���0��I�5C�T�S���i�l���.�X@�򇉅n�N��e��%je"T��\����:�� ��"byj%��S�? �y0��]�N���Y��3jq����"O��p��p��pJTA)k@����"Oa�	[�L����t�� \949`'"O%�C21Ը�Ue�8s���"O昀� �i�`h���!H
�"O��i6!)ekL�F�Ն)��
�"O$}�512��C�X�x�"O0	g�<~n���`������'o^��Rl	�<�݈��Z�ER$�'Ђ�Z2�� %��T���U';Ҭ|�
�'�t�ä���P@^�9�
��g�2�:�'�6�P��W������oM�S���'5j\: '�6[\��q@�$��Q
�'8��*EC�#��ps�,��t�U0
�'d�esv#�R*
�1/��a����	�'� 0�	�<Q��a�0h:	{
�'Gb��U����|%i�	ۦg�e�	�'X��+X�jy)��C�k���G��`�<�q&��|�d��̄/ar��w�`�<��0��@��,EK�q��I�Y�<&B��6EtM:3��#u�X}�֭�O�<ɗ��8V��BL��}*ZQ �g�<I4˕�>�`� V�V9�eA�^�<�e-td�(�7��^R~$��+b�<!�9�J���R/k����/�u�<q�gȣg��Z��7��{�TG�<!$M� )J��7�LZ8�q�Jh�<Y��m���郞��u��m�< dY
.���՛v��"���`�<���T�k��xVd�C=h�z���[�<Q5�
6-~B�&����dB5�DP�<	�L���p���_@��r'&
u�<Y"O��'�p��ǖ@�䙥��i�<q���VQ��C!7�v�Y�UJ�<��U�j��J���b�(؋#@I�<���P]�ڔ*��ܲEQh\e�Nx��'?,�(A0�P����L�t��	�'�:(!�*1�^]���L�3 ^H*�'d��j�%�	-�d��p �~���'� ����\�ntc��_6�L�
�'�@�!�d��	�4�i'�F8.�F���'t��%�A!~�J�f*�= >��	�'{���,Y�?�P��2m����t�	���'q�}��-U�{�Z� �jQ��:	�'e<	����%>��������'���R�ѺH�r٣R���߂���'$�+���"K���pO�#un`��'��쁣��
K�2Q����!V����'p�y��B�3d�-��%�* "�xi�'�%Y'h�(@���kR����бr����F&L���qf˚M@l�b	�I�!�d�>w/.�㔦J�tD6�"�d�L�!�@e�Y���8�1��
�g�!�d�Q �%������g�&_[!�$[�9t���_8i�V	��b� 1!�qt�4:TW�U}^�
�AG,# !�<, Q%@�@l�����F�]k!�A!��	�a��wX�m$ �`!�d�SH��3�o�)BFpcc�݌Q!�d0g�QX��@�E�Y��o�?H�!�$�#"�2�ISbB�u�,8�h�%T�!�W�A/�=��مg�j��:&�!�i�jYZ�D�� ����B5�!��Օwa6��2�C�V�z䇔�5�!�� �᳗b��5ߒ0!��	�HQb�"O�-�C��;J^Y��	�6uԴ��|��'`az2݋v,�(j`L#S)p��"`��yr�Q�:���H���`�1�F���ybg�L��Q`��]��0�@�yB�."q�[��A-���k�i��y�ᗃz�%D��y��Q�:�y�ʂ8621��J�=qo�)������OT"~b2���K���"e�,v7LP8RC�K���0=�di�:Pڈ	�"פO�HX�g�G�<q���^4�� ��"���P�B�<�!I�P�8���5x����z�<����r�`�u�H�H�@Tq�<�M˕R1�9C�냒QK��v�R�<q�,:(l�h� �3��0p��IJ��?�	�'6��ɰ��B 56\�^�VA�u�ȓ��h)�EX�k���k��H:l����Q��ab&g�HR<�9@@�l{PU��z�P��J�W�8��c�<@�z���J%`������(����|���ȓA2ĉQ�>&�pR��2�:9��a̓2�B��n��^`�Y�Bl��s���G"�S

��4�֛�Nu��!0ԨC��4A��bG<k?}S��Ò;��C�Ʉ����hU�`�1�6�O��JB��<U���Zf#��)JDK E��
�FB�I�zx�} ��(5v�hn	�c�0B�ɸP�$i���@4A@�j3�\W�ȣ?q��)Zݶ5`��� xr��v&�"�ў\��	�h��@��"��e��Y��H�C�I �ιc�E�K&�� �K7 TLC�I/�␙EH 7L��U�E,N91 C�I8g�ʀ�+n8�%JᏜ�C��2A����w+��G<��iwꎲL$C�I <>�� ��ɿ]R��gE�����d*�)wHh #(��#�8}�"���4B��H !&�����4#�@'��F{���G��U�
e�DBG�������yr��L%��j�W�y�t`���ybAA�.���9C,6�x���OX7�y"�@0\$4������&FB�Q��y�&@j������JG�$B��S��yRf]�l��j��F�@# 9䎏��y�)F-(E�Wh�9d�RC˝0�y2��m`�i��s��1�@ŜpI!����Х2��P�V�����I1!�Ğ0L���A��޼>��qR��#00!��&:b�Kdș�l�8,r�&ײ*!���]U�u���� 
u2L���; q!򤟦j�F)�4k	�+c��g#I�:�!��P�pi�a!�*U^�ab�*�!�DǑP��(qb��o:������~x!�$ԭA�R�z���@1��ի�rh!�D
�\�D�!��*�Ä�
]!�d��aͨ9�����F�I�Ĥ�(p!�d�=�vթ��d' ���eD!�D��=���#���rg�}�g�!�$�'s�ࠃ-H8v�%���!�
*&�4��k��a�@�;!�$#p��0hС,w\���b�5�!�$؈��D[R)��|S��^!�D�^FҥJ�Ê*"T��.� .�!�$X�t�L���iǷR"dU��ݖ{!��DRm �h��jb�\R�� t�!�� F��eG�]��+r�P�BߺQ1�|r�)��;9C|eb����}Ė1B�N�=Pq�B䉡;L~�Kw�Ʌ$����&U�b�rC䉍>�4ɑ�b�h�A�D�h8>C�.6ta@�8W(��2.TD�JB䉳OW0a��O۩b�I��b��H}�C䉬,�%���_ݞ��Ev�C�	�
�n��%#%W��sD����B�	�>�~ɓT���,����H*B�	;��4��1QɢȰaKD�2�bC�	�@|d8b���M�dI� ��B�I���Ű��@�i�((�%!��_HC��> ��`c`�v�(|��e�?@�dC�Ɉ>2|�A���-W�8S��G,Z C�	�1W�0$퍫]]D�d�<;hC�I�_��8UK'Z9\!�w쑝Q��B䉒,M:����O�Y-D�d�B��� ɝ���E(�p�!�"O ܓ2��,Nɮ�	�f���Ca"O������6�L�#��o�ʵ�T"O�:� L�s���9Ab��v�"O`���e(Ǣ ���Y�#%���"O*�����p<x Y���!��`"O��CM�R�.mbBBW~826"O�Up�(��
1 ų�(zYj�٧"O��!��q������qQ��'"O�#��J(lb�j�)?=x@"Oj��GhO����J�wN�Y�"O�d ���+��ݪ���vM��h3"O�%hf���5�6D��M_�>���Kf"O�YKV�-4�Z|a@ύ(%���`#"O�Z�Æ5�pq �����L��y�N�&n��hs�Y�5@00���!�yR%o�U����.��h�Ȕ��yb F���P�X/Q�*�RC���yR�O�ѣߵ7m���n	�?��ȓj�l�۶�?z��}k&ÒGP��ȓ�|��$��5V�I��N�P-�܅ȓ7�*��(�i��튑˓3+¸��ȓsن8��׆G����E΃-�<5�ȓ�|�)�#�R�"!д�]�f�4��ȓ4��3�-�B�}1�ȜHVDH���t���A],�$=c�ѠS�Ņȓ#��Y���I�NRTc����fQN-�ȓ^�b�	�lQ%<�"��p��E�d�ȓE ��
��XP'V�q2� 9x5�����l_&=a�t�ӱn�0ͅȓn{����C��$C�
!���ȓ�T{�瑒2�l��.60\�ȓjt|�gP5
�����pS�p�ȓ)��P����]3�@nRY�ȓ��@���;J�0;#��/hB��ȓ4ƜeK����/�4��Ƣڭf}!�d�20:�k�F�[����E��/!�B�kq"5*����(�@yZ�KM�!򄈱�$�JP�ݯhu�al�	!�d�9mԖ;oO��eHG*	16�!���.-�m�L�$& ��)_�*�!���=,qn�����{|��G�ڟi!�$ܫ,u8�:b�Ѿ���P"�,-!�ǌ�
I�7��<|�4��Вtm!�,:�*qm٧/�|��ʞc!�ɇ;�ҕ+"� B�8Hҩ�<a!��(V�BŨS��X��C��!�� �Ũ�kɚ+b���6�Ӡ8M<MYW"O@-�Eh��GKv9�rG�2נ���"O��i�A�~H�po�����U"O�	���U�� [�+��<��#"OJ���B�x���j�
v�,a3"O�@�D@؎h��p��RchP�@�"O��w�Eb�xDk�K��;^raH�"O9�S��TՖus�HB�~'�u;s"O��kpH�(<8�ၰ�]�I!�I�&"O8-�嬅d_&I"�e��8���Q"O�,[%	� �!�V���H�x�"ON�c�	�vt�aI�0F�p�4"Or�#v�ӸVa�h��4-��P"O��ÀFO7j�qJa��C"`��6"O�\��I�5�~�� H#C�d �"OD5)�(C#a�J�Z�'��{IV1a"O(Y�Ƣ�5b"�e(� `���"OZ�SKX�Z�L�a��Wۖ"O��Վ��!.�"v��=~��Y#"O���G���X*w�3n7\��T"O��B���72h�]��)��J��k"O��ӲSt�&	��(
�cb"O �Y����L�"I�3�^�S�d�QQ"OBM�Ph���)r�ֳ%-|�P$"O���Q��r0Ec��� �|@"O��p�o�!F��Q��["d��"O��sda��%5~�`U,iV��z�"O:	�Ɗ�8�dI�#f����("O
�	���PW
�2a�2��$"OH�J��
3����hI7O����"O�m��LtP�Q�Ι�Ol,�&"O*@� *��@��y��5�"O&�#���u��Y��?�:��"OސZ�I�8=�ԐR1S�c��I�"OJ-r�䇓HV��S�(����[�"OL9�J	�<���sG�$�0x�"OV�@�d��4p�#���hն��D"OPq֬B�G
��T��I-�	Y�"OF�"� �5r�b���fܬӷ"OĴ+$F�f�*B�T�M��z�"OzyX�遛b��+u�����"O�T{�O� ����G1Wt0�"OzH(`�'xl)��_�n>��#"Od��!�3�0�� g��u*��[S"OhI"� #D�p91���h�1ZW"On���V�r�d��hȝ(�vT�"O�]�4��X�,���fٝ~�Dܘ�"O��y��ٿ#.t|ʧˊ;*T:�:"OL�C��,�LT�mְgO��"O��4d���M��,Ǻ2O\Y��"O����W ,D��
C�s���+�"O� ��,DE\d���JT����"O���dE� p ��V��3r5��'U����H�\"8�W焊G.�"�'��;զ� qu.��Z�j�6a��']�E�#�I�h�<qc�� ?\M��'�v�wr��[�a�-B��e��'�V�)�咇�L�iT8<*�Ը�'$f�A򨃤y׬EA��1-��L��'H*�k�j�2Cl8�ʐl��+����'����P N!�00�*Y�[	�'!��8��
/`��2�� :M���'匕�. ����-"R.��"O¨r�'8b@�y��Ǒ
o)�e"O�  �8���a��m�fm��&Er���"O����e�z���8>jZR"O�P��k��t��cf׉G�x��"O$ �g,E5/N���E� ax�"O�Ay"�B�gߞ�sd��RE�@A"O����J��<�h�JtC0JC�Hk "O�T�`E�S�4�b��S>H3a"O�}�� T�D��騐����M���"D��C�`2K������`���3D��ƏZ��H���G�����*3D��4AŏJ�"P�H��K
�Qx4�2D�����/�
Q������B��/D�|����P��e�Z-@g��h �/D��e.ڵh��LcF�� G�4i�f�-D�(y�OZ8<�zq�U#�$��1D���� 12�\�k�`Q(���e,D�$���8z���a�S
����(D���l�|3fK��l[�Hj��!D�����R^¶���%> �����#D���qkA�ل�C�(M1�$����7D�@�#�8q��,
7��:M�����/9D� �5���]���pǆah��9�j7D������%"�̹7�Q]xHqAIb�<�C��4KO����	ژh��嘥�IX�<�dK��d,��tǜQT�MТ�K�<��"Q�l��8fbN�{ɂ��cŖI�<Ag��������ܾ!O�aA1dC�<��fJ9����*��I� !@�A�<���3�xx���]��]� ��t�<��KM�=n	(��X4�셁D��m�<���A?p���8�������`�FA�<��)N�V�nY( ��;H�`Q	�A|�<��סFDv��@!�Y�||q�)t�<���#$WH�PԎZ7w"�9�t��m�<�1d��[z��33��3 ��1��Z_�<i"�Ȗx�bݢ�hX�'>� ��^�<	4N�n.���[�0�3��Z�<y�[58�p0��_�:��SG�Z�<釉*k��ɓH��8\AYcG�X�<1�@~,ze{�Q�Dw �j5�X�<���ԪNS�0� ��&,��i*p�RQ�<���9Ąl��`	";2���b�<���-�*ɂ��8�(��Da�<���V:v�N"���\���`�r�<Q��U�=@!�R/�G1T<��cIo�<�SfX1_�t��$�!��aE-Hl�<yA��2"�h]�Sh���ܙз�A�<A($E�JT�6���9>�Ҩ�t�<9�!�0Ĭ���}%�蔌Ae�<p$�(taPo�WR�YHԯ�c�<q�j��?]d�!@��8�#��Ut�<QuCM/xn�:����B׸ZrBنȓ4A�¯T�$E��Gɝ���ц�=�����m����F�%*��݇�i��A��HE����b�j}��S�������HT�֖�<�ȓ�X}ÄK�.��V�ۑ ����ȓa�B���i	�z��ro��\&���ȓ��\@�ΐK��岷�P����ȓ@�~-��%P��Ja�R%�"���J+ � �\�6��cI 3x ń�L����L�#�&� ֹb�&�ȓm���Q(�7y��<�Ңa!2kKG�<!���ް���ܸa�rQ
��<� L�3��\�N�6�0���
@�*���"O�\	��T!'wv=�6�S�-甬��"O���T<B���$I;ֲ��"O�qQ����.�4 �Ï�K�=C"O��S a]�`}�QJ������"O�}�qg��H��t�#m^5k�F�Q"Oh�86C+%B��*BϳYE<0��"O`hHa�F+M��G��� >rX"O��y�,rI�.�'6,�B�"OPu��G&��{�C����"O�8R��< ���C /��&�T�`""O��JtL�QJ���sC�i�B��"O���F!DV��1)�!A3i��
�"O\�`5䔉S��d�b��A�t�Z"O`D�s�  �<�#Qg*��"O�}���C�OϞ���AF
\T�aP�"O�:iƲi��˳.[�L��\Z�"O,����
U_�di D,�άZ0"O41{7��=h��\�v��+M�����"O����'ބX*:l�R@7nLMB�"O���P�#"�pCD.O�@�az�"Ok�*�T ���,�(`� �"O�0S�쀑*���l�)!��3F"O@}:�����(�j�"�X��"OZ�{n
'?�D��3�:���z"On��T�X�M��<�2�H*�ZA� "O\T(&��OA��îP�sr��8""O��	P�Ln"J\���> ~�L�!"O��j�WfT4 �/�Cw���"O��	h�d�d��\q@��"Ov�{�l��б��o´e"O���)X�G,d��&�ΟCC�i	�"O� :RO�@_,q�Ǌ)d#*�Ї"Ojh��Ę��M�G�;��ӕ"O��r��l6��@O,�� �"O
LP��e�<D@��O�I:6�"O45Ѕ,g�	�1@\! ��� "O�@yU&
=�H�6	C%-�ŉ�"O�P�M�8 (�k��L�G����yB 	�{��k&n�>i�ⳇ���yL:Q�V�X�M)`�@����8�y��\+%�\���]A�q9Gj΍�y�/���>4`#.�V�����n�'�y�aĘx�����B�K^b}���y�MG<l��ٺ����7 ���ì�yB.S�"`~m�2�A�'^h(B��y�c�Jp �V�ܣ@�)�w`Q�y�˓X�|�`*i囶D\�y2+����`kC�HfB(�	?�y�cͷSF���$B�\�������y"hZs��86G�4Qh�$(6��y���2%1ܵYV��Q��p���y�D�PY��1q�F:r0���ǋ ��yr��pv�`�G�ΘcH�j���y�n�+����_�	�V�CF�Ȱ�y��4y\!��/�t 􀸶�ِ�y��V!+,���M(�j�UHO��yR�2�ޙ����M��0(O��yr�ɥn0�2 �ģ%6 �CJ�y�I��P�yO��V�@�P��y�ؖ6�je����V�V�IQ��?�yr�S%{�x���Fz̈��C��8�y"F'F<�d��	ۛx��+�Ɛ��yBoW��ָj ��s��Њ��[��y
� �9A���lm(�"R�75�V"O���b�
\�e!���/2���"O P�2��3������y0 ��D"O�J��U>/N���2,T��c"OB0"|P�8�I�$�����"O.�#%L9y쑢�a�x�� p�"O"u�"	�W��qb�5f���""O �Y)P</�\���}`U�B"OT�p$Ӯ$T���Hp]�I�7"OB�2U(�/3	t�1g(��L�j"OĄp�GN%���7�˟i�(�"O�dQ�\�D�P$8���&DX�0"ON`���ȈR�l%���q��� "Oੁ���%'���jg-��z~�s"O�{Ť�.+bR���KN	�\�
�"O���`�ܠ���{Ɗ��z�|�;g"O��C��;a���ĩT��8�"O��ZNV�IE�u�%�{{4�@"O����!��K���7@Y�0��"Ot��gM���9cK�J����"Or�#��V$��8;q�V�}��0�"O��&�Ӫ}5��@C����"O�qɢ+��f��t��*x�Q�"O:ɚ��W*o&�!8!�Nr^� "O&��1���&�����4�>��"Ot�A���BA"�3�6A�P�"O�嫓A�[�������s�T�a!"O�$v`P�Fm�`.������"ONi��j˧y�Vŉ0(�Q��p�"OҔ�1?hd��'H�&v�>��"Oր�F��Z�z�S�蝰0���C�"O�)���eu��*��|�bT"O^��1�[>Z�X���*P���Ec`"O�`���JL�� 8n��L a"O�<�F���F���j�3�(�!"O���AG^�Wc�ˡIǊ6�h	�2"O&AP��
.mP�9 k^�t�5��"O�%�����[;~490����z-�g"O��cqA�p$�8'`�=,����P"O��`�T�=~~�#�nWC�DP�"Ox"�Ƴ&�RkI� ��U�7"O|H��	�	:�t�8SJ<~|yb�"O�p��4,Y(,@�	���is�"O^��6�I-�b��k�}��	� "ObyQ-S2�$M�$
S,���0"OD����u�Р 	� Y����"O�@Q�NݮQ�ҡ��D�B��<�"O$��ڸ|}�Y	Ą�	c�p
�"Ovc�Z�l~�	w�E�Z��"O��fa׺n\��P� 
4O�a��"Ob!K�����\4�y$y��"O>��W�(6P-0�ȊA#x�f"O��z5O��[�����Q�D+S"O��b��w�y1�/� �@���"OH� э~��Y�Go�?^@���"O�!Aō�O↼��]�r��"O"{��&�`���];(7�՘�"O�A�@��s�j� �_A�yj�"O���򥗦#��Q�DH�[2�]+�"OΨ`A��!%��1BÒ�*x��5"O�!���#J�	�C�
����"OV)FL�0��8CU���V^�:�"O8�Yp-߰� ���r��P�"O�-�T�:���m��b����5"O� �HqQ(�9k0�qZ��	:�i�"O0���MW�t>�JCM�c��MXV"O�T�b��(7>�k1�,	�h���"Oҵ��ӅFO�(
�㕋\�} "OjD�r���h7��եL�"�@u�a"O"i�'(�6ڪ��n[3qў���"OV}sv��;Nn�ڱ��:�0�{ "O�,�iب%\�x �g�?,���"OD��iG�$`kw��W�PH�E"O�9�B�^�&!A�A�n�Ka"O�� �@C�$���o�RO��"O�i����0Ce����hs�h�+2"O2��(R�~�Aᐭ�7ۜ`h�"O�A�� �Q��{b���(��"OT:�ё'���b�k�;y�0��"OP	D�Gˎ�h7J��pLu��"Oz��fI�B�L����Q �}��"O�I���c�� �bIV�:�Y�"O>\[Q��`�~1�*G�V��tڤ"O���҉DN��3�*K`aZ	��"O4ub��ǡH&�E�C�ܿ(�
y�"O.��5/ ,:��S�³T�|�zU"O�ɲ �T�]��K3Q��"O,� ���BG�:UdM��㛝M�!��Q�e�)��2<r����!����,bqgI�V"�9�UA@�)�!�@�z�����."�<�QV�\�fF!�"sr0	WE�e��A���&,!򤜎T�,$k��#LlZM�$D�h!�DTi�ɻҨ-u0t@�c	�o!�d���F%�G�!~�(p-�u�!�:��I㋚�$��ݘ
�!��A6x4,�td��tm����2U�!�DK(\1���1�����	J�!�ė*U 	��ᕗ^Ķ8���e�!�D�&�2- '�C�0f%��i��=�!�$��UL!Pc�{�|��)���PyR(�2hX�Ls���oVZt[b��y�K�-Ҥ8���� ^����� ��yҌ�/KW��Ӂ�#Y1Q�R���yBۭ�jԙ1#���^yyb����y�o�(x�F�TjW0��bsB�y	�=P���&��7b�R�U>�y�BϏ3�>Գ��.�@�����3�y��G�^�����J�z1�ᐅ�y�N0
0ir�Q�t�0�
�����y¥A-G_�e�Ǔ�@jU"����yR���Mn]�蕊����m�y�	�n�nDj��T�xϪt�&����y�D,K n0��_��iㅅ���C�ɳ;6+o]J"����=М��'����,��;Q(pk0���a<�-��'~�y���[= ( R�l�V9�
�'V�=J�a���5c�
QǬ8��'��i���0�����J�n{�'�:��@4I�5�ț1�3
�'�̜ia ʔa�j�3%A>�L83	�'�� �/3����`K?Nꈫ�'�j�b�ǚ�a"� ���=X���
�'X��j�>��P)�$��|h����'� �çh(}�|���ʿ��9�'��X�Gc�"<� �@Ջ,%@��6�\,0��
v{R�{WFMx�t���A�S.Ze������
9Tԅ�S�? ��� P03�V�Y�ʥ~ȢD"O�]Y�>Cf�="ֆ�,��9q"O�U�d�'4Z����W��aI�"O~�fiH�A�����?4V$�aG"O|qiT��~l�Y�D��)@v�&"O�(�F�2*��lY���
GL
��*O�Е��h�\�2!�����
�' t�Ϙ�Bb�R�G���{�'�F5���TG+���Wn�D��EH�'@h�ȝ2�}�PKM�oԎu��'�㍐�j���V���a�L@�'t��S���0�^/X�ੇ�=�z܉A��_�� 9�)̓\8���ȓe�ĳ��ݑl�<J7�&k}� ��H��} Ǭ�?+�.4HS��1$���JO�(ɥE�a���a! �B�)��{�kƎ��@��F(��v� �ȓ:7I�D)?Ρ�lV�3���N���9�+� +�6\ G�
ݜ���7}���O	�AA,�Ud!��@$��H��|�ׯ�*���`�ް�B�É�h-@�={��ȓz�� ��2N��ȓ4�K�7,�i�ȓ'>�X��&�.��P�7�(I�ȓ/�,�:6ףg���#w,ӈD��H��#;�8�V�ɲA�sá�WFE�ȓ$���FB��>~l�ȓ%�RE�wk��t����@&ي4 F�ȓ#\ �#/T�� ��ʚ�=�޸��M��Sv�- #���Eك&�0��ȓ2�b����]�Hf@�k�ޣ:'t-��TT��2���@�"mN�ϪلȓdN��'e�6)D��B`��n�<�ȓV�Py2�@%њ��Z�&X�ȓV���H䀅'��⡦Bv�&��ȓ@&��e�
�E��D�ԅ�i�b̈́ȓ���[��U�vפy+D��a��M��wܱ����	x�����	�lhD-�ȓ6��zRh�i&P�
)���ȓ����ȉ�>�d�'AZ�!��l�ȓq������7�PAx�aF �q�ȓo���qM�4i`�mȥU�VT�ȓs�FH�ŬC�[��҃�|�p��PU�U����%�ԉ�K�(�ȓ{EN��Bo�%����b�ԅ<�@�ȓ?��p��/�aB
09!� �:����z^e���pNl�(G�P�V��ȓq�0 #Տע4�����]�@���$����
�$�3�mQ�6�����7,.�P gC�:� � �f	�Wo���:Z�x;�� "
�@1@��ދJ��I��t��a%�{�8 `�/e���ȓK��1����>�\ccL�S����,�Ry����9j\�����[X�L��x����#��<1ؔ�#B�ftZy��g6��glD�&�����iiL��ȓL��-��I$;�2��ӧ�1H�8<�ȓ8��,�&m]9Y��{7鋖Tr�<�ȓ�|#��=R~�!��̝'��)��&x��&kϛ�n	i���7��ņ�jb(W�q��_`���ȓD�\�����	KO��	�J��XXY�ȓ|A�X�&
(	r�
DK�+TH��g���c��d���"�)NC�)� H�Cdin���ʇ@ƚa"���"OxM�E&Z���ŠL y�]�"O�|�7��.z�`�`�C���"O�4� \�s��Rn���"O�M���źdp*����>/YĒ"O(L@�o%r*TYc��.K��j"O���w)w� �	��ݕvWʬS�"O��	��6z�Ljn,(3Rp��"O��4�_0}yJ�X�M�]�"Op��ԨV�7�6 ��
���K�"Oxx���ʤ��"C�<d��d�v"O�XS� /;r��t�RHan�b�"O��0�zD@����8b�����"Oha�7ʀr��Q��c�5�Ї"O��3p)�	>��V��	v6�2A"O�y豍ƓEk"���HT�kKr<k"O
��玨~Z2&� K,�%�"O:\ZB��	={$��"&�D� "O̫�Gk1P���n�"1l��'"Ov� Í�}2���  y�^��"O
E�I\�p�|�R�"�2p��"O�0�@D���u�P�z|B�"Od�����#���`�\�
���1"O������%ML���-�f�D�0"O�����\�f`C�e
�Ph}3v"O��a�!�5[�$5�%���d�K"O���E�B�\8:�8�ҮO�!��� �zQT�V�mN�ř��%$�!��6i�5`%ɔ*Lڑ�"��M!�dC-!6h`�2�*���nĊP�!�$Y�5�x���VϜ|㴇��^$!���(<"���`�8
�E��G�T!�H*o�j� Ì^�;��<��Ǖ�b!�7O�h��bV��zi�A�p"!�D��]�p!�H����$�s!�d�#=��;EF��U�8�p��K8	!��?%J�ɷ&��tg���虄n�!򤁯7-��!c�X���>�!�D�hC��#���4 �y/Z�(�!�$�	��k���s�t�I�!򄍧.0�Ei�A�cj�� ��^�!�$�2]��C�MV2HR��s�σ1�!�� �aN"��$GW?�퓐CE��!�dI�H��!��ܣqB�I�#�g�!򤅧\��тӮ0W��%¡��+8�!�dMH&�2'�
�Z2U� L�n~!��֋	xt�b�C�ww��(p�$2w!�dC����PWIi�X� �H�,w!�$I�"�z�x�	 R�X-�al!���Ȥl��#����'[H!�䝬=��q�m72�P�0�O��x-!�$��j3���B�� B��j�<��N��k�ŉ�f�:��.���ȓu�������r1��+~�*�ȓ%[.C��(�D�"� *-�`���th8�J�˘�f:�*��@?9C���A��=+�F�9ڎ���7T�B5��@�R�����Vd$�+pV����dUf0���9�0L����N�ܥ��-�d�t�ӇWv��ۤ@X��2-�� �@@�gI�L�J�I*�LV��ȓ ~J��R7U^�9䞼����a�L1�`�-���r�ݠe�\��
��j �øG���j�"^��Ȇ�S�? �=���� w��\��:��(�"Ol� ��;gj��#Oэ�&�P�"O�"UA���r�C��|���"OPD���� 6)2���U�4�A2�"OD��@/]"<�"��6�ˏ1 �ʴ"OH�yA�L�$��f#��B2 !�"Ol96(}�2���#M�� 
�"OZqɠeF�9��[�,ܪ#�jK�"O��d����h7&^9!U�
�"O��"���ifB������K`�rS"O2�$K^'1����}B^��"O���G&@=����±)b !�"Oz�
r��x<��q��f	l`��"O�bk@�^�na����,*��9�#"O��ؑ��d)�B����t��f"Of��5�Y��`���#*yXa���?D�h�@A�$*�h�3i�.-� K*D�\���5�p'ҝ)�6��'�&D��R��EN=���c�ì�(��!D� �Ѕ�g���BGhB5����!�>D��:gA�OLT�DdV�U���
P�;D� ��	�&gP�C�O<B�\M���9D��Z�/�ѸT;� �<�~�h@�8D�:��ߣP�^�q"��*v�p��G<D� ��IC�s��$("����<���$D��+�AE� t��(ǥh��z�f8D��s���S���s�:Fx�p�#<D����L�S5AH�o��&����9D�<2'$�D��D�����b%D��i2�H^%���G� �ɤ���7D�H3R����V ��L� px]�0�4D�ء�ر�6m�#I�>f9�w�0D�P��G k 0�	F������;D�����y]�ah�1V���$.D���Ȃ�Nd:|��aA>�d[!� D���C�� k�@q�dA�ckhQ$T��r@�Ymmh�9�-Q��8�a�"O�]��m�C�*�@&�E<�0���"O�<�o�&L�B�KS%˹8c,��'�(]"�b�-V��a#�P'iL �����!����-�4>htER�H !�!�D�3/�DC��|G0A26#�1�!��V�^&Д[�͟mMLu �i�){!�G�����z$vx�&�H�!�1 ɡbә�4��!�DK0~9N��A�ث6-��A����!�D��
,+wl�,SPa����9�!���k�"urF�	�L	�d��6*!��XlN�SQ!c�h(i��W!��6庵�d!F�p�^�z��Y,d�!�dS
��[rW<���H�H�+�!�䚥N�z�'$?G|$�A�Q�!�D�?C��C�,Ɲ!�����a��!�d�-#:����-(ʮd��C�:+�!��$An�ȃ [1{�����Q/Za!��W�/B00n m����!nİv�!����=D*�"��7(�����!���z��9yu���������5�!�$FzN�M2q�I.W4%y�ϑ�
L!�ė-'�.)����AD!��	�'�����ԬM"�p�"a��R �3�'�����"v��e�"k�U5����'pԁG:=���AG�ZM$�ϓ<��ag�V��D&y���$	�e'��Q
�qs!�d�?0�����=s�ء�j_�1��'x�\���?	`��� ¤��.�b��tp�f�{�2�Yr"Oڸ�j�((4�
��t��SPbͺ)�B�,�(�9�`$�3��ۗ{2QU�?MH��A��T�E�!���y��2�PR�x�yeÉ�A|Z�:˚� �5�XX��(")�4�HX��G!F��ط�(�l�ttᥓ�A]�)��jb7Ÿ;��@�0�2. }x�!p�<9Dh4`h`����`�sy�ᙇwPh�#'���i\
���(���sM�x��9�!��8yg�`X�kA801�EC��(u� ���
���3#޵Wq
�:�Y>�<�Q���ű@��+��Lkc�UHX����F�0F�ɓ	�6�]%
֣�x�Z�I[���0[@y9E�Vc8�:F��� �n{��!��Q�$�q`P�3|4��Q`D*it�=�Q ����ƅ�m�}��K�+�aҴ�y�X��z5:Ƨ�
���!3���I�"`{T�	1	Q=Lxu r�l��ygA�h�(y��צ�~Ma�.�yb�Fo���*�e�}����BX+�|���kX*AP��W��2$��Z��o���Fy�D_P��\k K�pǾM9ҀS���=GL�'.�7$��U�:A����v2Z��Р�bt���]ݮMr ��a8�	�g��ed���tn�uK�����;�I�Rq�U{�F�����3	�j��0;5G�?�°"�m�:I��ƑP�qҮ<D�4J ��p���I�MK!>�ٳAi\����bg�C֪(��iѾ��-j ������@ߙHY䵰"�=4$Q�4�w�<!�.Ҫ�q�#j׉(���g�֮$�6����P>�h�����-{�r�"�Nҫ|��<YքR-xh y&��z�Z�*���i��L�QC�������M�P|+��c@��'�Q�]�p���4U�"\s���:�p>��	7�8�RM��-:2�ã�b�ũaϐ�H��6	U�o�"X�a��I�qQV0I���6y�W���!�$�1\���C�e�,�p�E�H��<�%�^�SU|��2�M�qU�U��0��O�*��;�Z�����8����ɞ:
8D�ȓ|���Y��Cf�\�RaB:q�,1�7)I��* �)�.0�K��ӡ|���aP�"ʓj� qK��ͥYIH�yb��9b+�!���j�|��.��c���JTMA0m~�����<C�(h��
f� �vN�-ւ!��"\X���6nA:�I����	�=�h��K�<�r�F�v�m3� N���謟FAY�R$���@g�6#���D"Opzt�})�!�0+O8�a��v�|  �'��)��D�0@�P�J'§�V��MXa�c�#d�n�(p���6L^C��-�h=�#$��$�nM��4��l�R��=E�s�5-�֘`n�ٺ���N�.:V����#'	P��ӟ��{� ��wj2�9�M�,9��D.� !=�A��@��.A��c��,A�	
�� l ���(��Aѩǒ8Kh	Ex2�-#�hɑ"����Xgh�����ah��oOЄ�B"OH��&j�>���Q��V�{OF�T��)m�2��͍���S��?tR�5�Y[G�\�VM���Kv�<�R��98�N� �EXr��f�p�<9�*ÈJ��X��A��\1AM�q�<3�ސ[�����QQ�t�E�n�<��k=\��)�i�?�`��RC�o�<IM]���yqh���e�A%�d�<��+7~��W&�*8���Dz�<y�	;m��*%a��e�E��`�v�<i����j��+V�!xvB�P��]l�<��Y$n�: a2M�"X��U�� �D�<1ǌ�'ǘ��T	�=��9�	_A�<A�L��:�F�R��W��ܼ�F�B�<S�ױt!��0r ��4�L��M�{�<�Ģ��d�!�Αei>�C7/JL�<�CG�*F1��޽r�4"� O�<q���6eFua����%˕@�l�<��\5?���WI���T[���T�<9�+��d�0�`ې'��H����<9@�ǈg�(�b�ě�88E  ��m�<ѵ$��t�)�:F��DX#��j�<	3���Nu���7�B0MZ ��De�<	�f��$���� �,.�n��i�D�<� �LsE��L����_$~E�T�"O�(Bp�ߡ}��;uF�"x>��HT"O�,)����r�`[�f;7��@��"OS�%�7임 �ޯ*����"O�ڲ�!H�<٧ٕ(�� !�"O.�f�A`�
A��#�R��Pq"Ol�b��9:�c����SV��"OB���N�3�hX�!\�.F����"O�Yє�P�_r�Y:�[�i� �"O�EZeH�3~� U²�4@G��92"O�@��·W���B��A����"Op�ۢ͑(`�,U��ѓ\���"O4|�r��$?,�1׫�3d����"Od�I2j��c�RA�F�D���U�G"OT$��
k皔 @�PZ�0Y��"OLU��ɉ1�$�YBW.(`ڒ"O2�[G�܁`�H�(�s���e"Onњ���b�CF�ߠ��D�U"O�U�����ؚE�<1����"O�$3�ț����yb�5�mk@"O�P�ԯ�'���!�G��d4�@� "O2,���8�}k�� �"��"O�Rab�,C"���1�
��F"OX��Ī$:>D��d�=gPI��"O|l�w���Lu�����ˉqH��;�"O���M�:5�Z�{� Y8O�ܰR"O������>Yu����τ�s4d��"O��yc�A�[(1*M��f?��T"OԠ��9K����퐮z� "O�<��"]3\�j�P5LK.�IY�"ORLr�Z��Y��k�#1^`���"Oh���"3hȹ�)!p>zź "O,Mkp��.%�V��F9Ctp��"OJ�R� �v�����G�ok��3"Oƅ�.7DQ���Z=�0xg"O ����?10�V�J�L"�["O�t ���[�$���&חV���"O�TYюW2*h6YJL[��"O~���Ht����#*�=	�:��F��'w٪�ڍ�	�Kd�)c	;D��1�HٲJ!�d�=j�����˵ l*p��ԁ24@ѻ��I?��gl�|�'�$!Ă�V�`˅EA]3���'@tB�eV�X_��4�I:W���b2j�E\n5��刡LA����	�`���!�9yYDT�%�խZ���d�*r񺜀D� *Y��ۖ L�.�![��P�4���0�l��*���!��ېI$
���F��f�'�$�G��	<"ђG��3t4�F��)Pu��h�+��nO<�Ò��1�yBh�X�vq�F*��t��1�&�U�x��8�厗�n�t�CG���i6P����L>��n�Mc��i�%�v5D"�(<i��n�|P��B�p�9g���Sa���&��pҘ�`T·�q%���G1�������!,�!��Φ/�axR�ߦ<� �(�mX�z~$])��a� �`�T��h���� �̵!�Orh6Ι	\͜-JT眄wU¬�Ɲ�<C�N8澨9��H��!���s���xAAaKG�]0��IH�~x`݆ȓu�HCu@Ŋ-�b�&�Qq�A:7K�7R@�ಯ֟[k��(�G�f�'��.Gf���EW$B\F5y���KV��.Dn���*݌?�n1�`�S�6���X�����C� =(5QC	��<���(D�`��ƥC�u`tp�Bs�$�F�6*��kC#��w*��ʳ'��w�u�%�]�
�ڡ��-��\�Ɠi�0�#f�\��%���R4cS���'���cDMZ�m;D!�m^]dΜ ���L�`��� ������	4�!�$�T���x��`�
t��(q�dG�Q��!��0LƠXLC1�ĒO�`��iP�l(��u�$=�0
O4]�$"��v��9�J'�%��^�8
�c�N���0=� �PB0��=`��ls ��6��@���'���
�A9��T�sF-����4�Aa!�;{V\[�H�I�<��g��&�h�Rp�7
-$��M�ɃoR\v%[�}����$^m�Ojd�d攈c���6L:f�����'�(9�Ĩ	��`��Mv�6*ҒEJ�b������ � ���ē� ��슰(�@�"^sBh�Ɠ�*y��	��.u���ՐEi�y���R�yԒ0
щ��
�Z��䒠pL��/�I%z3v�zr�z�#�	�Y����<�g+R�X��<AR� ~HiR!��Z�<� 
:>��T ���,��g@J��@�c!�v��d�!(�B\8��^�y��.�>�I�)Cy�~5`��ѻ_y���ȓw�@��"{���×0*k\ ��_��c�"�$h�"��%l��<�ȓR5B�+�)n�+-"n�`�Q�"O��rA�I&��óLs˜u:&"O�ѡ��՗r�`Q豮[�w����"O����D�?C�Z�;6�]<��m�T"O(��q�Uk8�R%�
2����"O�)�'f��lF��&*B�*�,1�d"O2p� �(�X��P���w�1�P"O��%�47�`1C�,B
M
2,��"O�tt�2T����A��q�	
v"O �Y&k�<������&h�Q"O�)3a�)Q6`	aC/�zeb=��"O4%����302�{�,�#zEΉ�q"OdS�l�s$r)c녂G���kG"O�p�����*zpu�j�8st��[ "O�}Y7Q��R��d�Ot֥�W"O�̓���o0~e�`�!P�D���"Or�C�ʁ)M��l�� ��p�Cp"O�q1�
�z᎜c�H� dy�xr"O��8hB�о����/fb��"O�a��SC�F�pǫۏXfN<��"Oΰ��a�;%���bQD���� ��"O����C�h�:T+vĞ�[�z%�V"O��r�N�0��X�	Q�a��8�F"O,��r`�#k����ȗ~���f"O�u�VC�;pF���7a^}��"O 9���t�Q��V	)g�ċ�"O2|�2%�Z�8k�)��at����"O�EPT�D�MZ�И�'6P�{�"O*�s#�V�O�u��ѯd����"O�,Z�M�:\�,p�Z8iT^Lq "Oԉ�c�����r�.��N_Z4��"OvuZq� wƴ�'��%ʐF"O��!ਛ/n6\X��ſP �q�"O�]�Q �4	N�� �M�[���4"O|�
GEU�lf�8�ϳy |T"O���I�W���J�&ů\QFy
A"Oh���zҥ�g�[=*�b�"OP)CD�B�iu�\�a/y*�$��"O�cg���>���J�oT
P��"O���P�Φ0��уM�7
�4��"O JN҉�6�Q��D��.�"O^�8�V�Z( @8t��ag���g"Of�7`�*�`�)���W���4*O6����ܱv���
�V�s��1�'e���C�	���cϝ	�f�S�'E��1A`ʐy;Z��1fye����'�Lِ�cwJ��PPѱ$���z�'�81j��p��m G�A;���'��cƊ	#JR�0:'@";�$�H�'|~�DI*%R2��fG?�h4I	��� R�Jt*R�|.DT0&�,)c!y7"O�)�k��v=5��C�?ri�t��'<=��׿��	%I�.IC1�O	6xձ��� C�I=7 ��R_"�8M42[�O@�ib��jg�t��Ef*�0�g��p�y�o��g?�B䉺�Tͩ�)�?H<|9� iU�(}��Cq.U\~�a�+W�T�}&��W(��'���"�1g�h`��+����Ø+}N�H4�>H�Z��a&y�h����GE���K��Eʂ]$t�վ��b�&�w�@Ah"�Ō��]�J�q
g��V���o�J�E���W�<Av��8sD�!�w��*��d�Jgy����dL���"�>,�����	�;|:%q�Ƃ+H4�`�C�f�!�����[d���o=�с��D�I�t=apAڸD��p����{�Z��]>�<aa-��u��Y��)V�8;�Xh�KsX�H��D�5d(�y���G@�F!�g̍.k��s#,-X�`xxU�|��`��	� F���+�e���p�.֊YJ�<١%T�&J�ۥ�c���(T�����O��	�@�&�����6VX���'���w��9\���-�8ĩ(��x�ց[���1%vd�q�I��E��w�rd[G�hW����Z[(�B�'��lĄP��* ��/��u�h�BI��A �#I��R˟4���o�'�Fi��#Z@���j\�t_TX��n��Y
W%D�n�PE�+�!l����@a��q��i��d��%j��^�I���P����&�]�Ipu�fb�f���D�l3�v�c���8^�:܂��51�l�SSY�@�C�^�(�V�%\}�PC�I$	��`��b�K�耺t�F !<U�`om�"A�F&S{^a¢���.Y���4�sޅb0�U�Z�b����u�j�#'=D��hB�+�G�4���$LV�a[^�8ⴍ�t#�/�J�z�cF&G���0��J8 �Kt�X%�@����5���d�9,Wfܢ���6 H6��t���c��y��̒�{�Թ�L7nH��Cv��5Y�$!��I"c�(��F�Q��q�%W�DB㞰����'�-���j?L�j�L�)���0�O*��R�Y�8Ć��k�?T��yC�'�8�"4��mA�XId�<P�zlƩҪDL ��$�B��kE���a�0��~��x���T��sƞ��vg��F�D�b �,D���-̸v�]����(0��A%i�t���;'�i��\Ӳ��Q�����9r�Q���'�~<�
f�XC��b�7\O�	A�%r�����D�thVH� g�iؤ�8��^)d�,�AFĦy��-�K8���q�_�jQr!���U�Sjmke�#�	(����`�f��}�����dȨ�k�t�]�E����ȋ���@a�
�yҬǙZ��BF��Fw.`['*5p�t���.��`͸5P'��v�:M;���k���-�!��
$qiJ��nD�M�!��G�E-D��3�%Ji�A#A+E�3�v�S���<�@L����5�Z����D|�EA�JZ�#%AC�Q���rPEX���=	U͟/S�����AKx�Y�͔.J�x�t���WZ���	�N��	a@v@;��Qfѣ�I�+id�#<i�;.ƈ��F�Sy�O��Q��{�>4��f�!FX�];�'��!q҄٩dH"���Y'7�F��qO]&O��Z�Rz�)�矼
��%�����_�q��\��$D��+��<,��9GK�h�
ݛQ�"D�P!���s�v��@�eF�89�� D����&Ǽ_v@��n"tMR)� ?D�\#�FݏB,�u�p�q$}�cd?D���E��:�\-�fC�S���ڷI1D�xB�ٰJ�=�[��40��L�!�$�PMz�Q�Lϔg�MjA����!�dJ�Oc�)(e�ǝ	�����x�!�dӪ}G
8�D�=*Y>ݐ���*De!򄏛[ǆ�p����x@���&�#?a!�$2�	����7DT��(�84U!򄜫YP�@! 6�������:G!�ĝ3��Q�m��<����-�I!�$<vpƱ�5J�7)R}�흽P�!�YGB�뵁9?�@�\%�!�H�Bx�A��� f���oB��!�^X�u
�@�N�>՛�?V�!�� H�8#�Ϩ.�������H��"O<�YS���@6`�2��<���"OHU�A��_`��,*	�}S!"O��#L*RL����!��n���[u"O�YA.��U���ˁ,전�"Ovyc��ppSS�I49��"O�x�/�t:�h��%/�Y��"O�AbU��eD��
Ts��,e"O�)�V��/)�(b�j�3��J'"O�aCP�2�2H1		��!S"O��0�ǻ�P(r�h3�a�R"O�3 (D�/,
9�ѧ�M��@JB"Ore���L�D0 -8�������"O0DR�����|�*�G��w����"O�����$��xYW&A�T����"O&)�e��x���%�����"O���ូ�Q�O��g�d�q"O�<�P.�DX��J!a����"O4��B��}*8y-ȈD�����"O��FYp���B�M�)
@}Y�"O�i3��$+,PP�6&�p�\}��"O�u�b�ށBl��)��J�
��!�"Oz(c�_�}P�Z�gU�_StJ�"OĘ8@��T$��D��@���*W"O>�s�cI�1R��PD�rQ�X�"O��P*8&�,��Gʞ		@�qA4"O����ZTX��2G*���"O�T8ң��/�QF���]�D"O�,)��		~Z�$SV�F��rA��"Oĉ�J��^��c��X�A�p�&"OR��R�!Z���Ыk� �I�"O��"�ŽT�^�:dM�/r�6(ʒ"O�	bu�R��J�.N_UR�h5"O���Vc#����l��s312"O\m#�L�6m|<(ؔs#f r��>D���,�w�	j�&Gu� ��"�:D�X �/���Ƭ8��?
y��ɶ�?D�8� ��#~[1�2>K���(D�䛃�[�^(��y�R�F�����) D�9d*��/,���BM/~HD��s�;D� �a�Z�H��5���)L�f�2�9D�xa`��b��[@\5B|<i��:D��ۖ�nz�8	d�� i.H؋b?D��I�eĜi� [��W!FdLB�N/D��b�ؽL�V��'l�lE*D����.F��Za!�d��F�z��&D�hI� I�6�J�k�*L�
�����$D�x�����T���3rf̂,D��3EߏN����K�B���� D�$�A��2-��zW���8��<D�xs1 鶴�5&ݝD�
����6D�4ĂT�-�-�]��0��8B�	�z��L�k:@�J e۶)FB�I���p�W�eB� x�W�$:B�s��$q&���8�p@��9SB�	�H�vE�C �Q`�����Q&C�I�� I�bذ�d�b`f��C�	1ne�zs�é�����`�=�B�I�q�D�1l�96eHAk��A�O܀C䉩��L3S͜L�N5�C��m�~C��f��LD��~���&�6QMjC�zZT
�3M%���o��bgvC䉟s��3�-^3k�U�@�	/~W�C�/?L�H�c:&�X�с�8�<C�)� ���T´C�uC�m̊��l�C"Op��3�;v�;Cl�{��љ�"O��Bu�ҏ_o� �,�p���S�"O�]��MތH/tS�!n�x"O�����,
�Y;7l�a/�ę1"O��hW��(F��Cu���[!"O\���C.v�I�'*<���"O��#�P����"�$6.�2�"OI'$D�z�x�x5!D�h����"O8k�@<DZ�$����<k�"Oz�J��;|C��r��{G�!"O~)	��F9k��|���SJՋ�"O<)��G���6a����aZJ	Y�"O��B2�;1�A�a��"���
�"O��{`@�)�\��/iwԜ��"OVؚ�+�b# %P� ���2"O :D�4K�tض���9kBi��"O��jo�������4m\2�ڇ"O,ܰ`Ʌ��89�����9ؔ�"O!���?^�ҁr�(�Z��<3"O`@�C��6}�l��B"5���@"OF���2 ���K"�A�!���j�"O��ѱ*�+g(8��oB��� �P"O�}��͈���bcy�"O�0ʷ�3�:�b,	#(_\�HA"O@-y!O	a�)4="D�[�"O4X���}�RHt��'�]ʢ"O������Lɘ��ۋ�I��"O��Y�A�|�*�8D�� #��Mb�"O�\:U��+��m��'�(�� 4"O�]����`�ҥt�ɉ�X��4"O^�Kd`�,��m!0e�F�V���"O��"񥆉|��,P��FPt�xA"O��' �:�Zm��E%29���"O��A!IQ�����4]-r90"O��V��'�\����w0�{"OVɋb�-���c*�j�$*�"Oh9�Ř>*�����
�z�����"O�ZÐS����rE~�\��"OL�y��Q
��ue ]�`�D"O��4͵EO��aD
 0��k�"O&�$R1=t.��֗S5��� "O$Y�a��6xA���1<�
�"O�E9���$(�9�nO$_>.<h�"O��8g���M����a*ļGJ���"O�E���Lrb�8��U;D� Y��"O�x6�ҜX��a㗢��� �2O2���ٵy&$��1���$�1 ��ɫ*ϒ����,@�X�$�V�f0B�I�.�BMjs�_&?�����('3ZB�o�n�x��=*}�����L�h�C�	��� o\��Z-)��Ȗ����(?q��U�~}�5��M��`�<1ԌˊX��-q��UQ�H�1U�
w�<�a�¢��@` "�k���S&)�l�<�*j.g�=�.Ԫ��_e�<ɶ疼KpxH2'UM�ܐ��J\�<�rُNHcƝ=S$pZ�bRX�<�g,֢?%v���G WE�	��nJj�<���7h�� ��DP��	d��b�<rDث��E�2�r�,^j���E{�G(�����"	�2��x����u��<q�����'v���yU�C�2LP<����&WQ��9�V�4I��ا(��$A�أx�}z��Z��76O�9�'
1��?y�>0nԐK: ���E��E�f^��D	�����?� ���Ԉ;?.�Ivcէm���Z���H�'
v��i�'`��p�A�&��Ua�.��Oڹ��i>��\�`y��S�/ت�����!pz��%�P{7��o�S�.PX�g�ݺ>��S���'�%�'���a���ӟcԘ����! �x|S`�ٿZ�>����(O?1�WDϺd�	�	��ł�"ac�<��?3mZ��kMe�2]
4*^�<Ys�  ���'eV
K��,jEq�<�%[�M̆���d��#u�� ��v�<Q�O q���A(��(�6��G�u�<��d��*��=�t�zA�^p�<U�K�N�0��q�5JӁ�v�<���%(�p�ڇ�w�p�³#�r�<A�čA�Mh/	s$��+��s�<�0�\�P�2��@�߂��!BIW�<�� Й-�0�c��,+5�CQ�<�AI b��e�,j�x��&h�<�r�S��Hf
�*�T�#ĬNb�<�p�O��t���n�"t�ƽ����C�<!4�TPj�!]:�����=T��J�M׊GP�[��(1`��,D�$��h�4���CF�0_?��;�+D����n�?U��P�a��t)�	��(D�v�i�ê���j,�+^Rܘ��'c�0�����8�ʹ匊+j��x��'�\	/Cd'���Tˉ8_(rt��'[D��@�1~t��3����2��'��Ĳ7�ù^�003��%Py�i��'z`a�� ����oV�xXҁ"O�Q��R��m2���e{�"O~���
Ւg|��f�OV�8m��"O��{�jP%H���S�|x�0`b"O��"��t[r:�o#O�\"OT��c�޼G�D����G��};"O<� "Q�Ԁb�G�K��9��"OF,KՇU>�\tq��2\{�"O�Dį��@�y�i�6)�NܢT"O�3�Z�i�D�V��D�aW"Oz��S�L� �q�����p<�"O*Ⱥg�?}�x�Zu%VT�\y�"Ox�Z �I3"\���� ,:̪w"O�$U*.�:�c�@�#m���@Ot�<���4\ܦ�S��R �e �iF�<�0�<QLxPc��X���t�C�<i���q4�rD�O�S$BY��|�<���W|�qhEF�	(�\��NJp�<��-�8vA\�����f3�4��YV�<IuaN��{&b�*�n!s��\h�<���:H
fLЙ�4���Ίm�<��@'NO�E�D
H<�!�:�	���S?�b��v�C�!�d�;�Ԑ˄HG�a�Tat(��=�!�d�)U:,hF���p����>�!���f�p}�$+̀{�d�<D�!��;�p��C�� n��i�cܓn!�1y�J�" ��J�����4x!���+�ΐˑiBS����T�'
!�B�=^�yжK��+�>i	��I�X!���(}���#T�2]*6�1a͌!�σ.2 ��ߒy���cj<'!���x5f�s�)^�+׊ZD�C�{�!�$�|O
͡P#�M�E���	>�!���
�3qO��e���1%�ՐF�!�� �,��l�0���!"�M�!�� �4�se˥H�N�s�)��aQ*��"O�ɘg�ωS��E�O�{1Δ�@"O<4BfIE!g��0���DЀ#�"ObT8��Mӄ�x��>�@��"O~��@��Jy����(��+�"O�ܱP�GC�0��0[ɪ1�"O.��"i�&E��ð�>�.�k�"O@з��&/6��j��LĲ�"OX�C�jB
8��i�>��9;@"O�ҥ�%HcV�۰g��i�DQ "O��`Q��6Yd��(��[�B�Q�"O�lySǅ\��j����\���p7"O&��`�M:����83��ɉr"O¬�0�)[�X��W �F"F1��"O̙��A�"_ܲ��ɪ��/E�yrN)
Ll�����	�~�� ��yG�L<b��d�BVI�`������y�
ڀe�$Qum+c�<ēE%Ԍ�y�X"�YG�C-^Ȇ�B%O*�y«��l���b%l�;f���8 +@�ybM�2<�LAbq�-
^�,��
�y�i�d���r�9|�´3G`�?�yr�7|���8�h�KB�K:�4�ȓ_nq�1�ѷ	N$萦�+O���ȓh0�"�����['Z�9[�̈́�~s��b��!�r,a$EB�2�:Ʉ�,,x2V
����i����%�0نȓ �%8�mX*���V�R�5����!!g	7~u�����ޒ
��-��{��T�&̂��ʔ�We�)-�l���$�.y�p�֨Czm�f)�r�L��t�RI !��+;�4�F��ni�݆�7V�m�"��Q�F��e�%���|g�� 瞹+�A�SI��j �i�ȓ?�*	A%r�lx�Ğ�_v�����s�K�����E���i�`���-��1 !��R��72)h͇ȓP�Ј��ŕpf�u�i�	hE���(yy�B��WQ�|�'���8�ȓj�"�Y��XZ�P�(�*n깄�~�*����	�y���TBD<XSd�ȓ*q^��m��h!<0�&��k���ȓ���1���{��)��ί>M(X�ȓf��" Z�h�b�[�wX���G����׋E�7���$Ҽ~�怇ȓx\t�h`-��7P$�s6"\"h��@�.��b��	=�|�U&�5��}�ȓ7b� �I��T}��	WKP�r�J�����QCːx8�6�3A��9��b�� ϞY�at���捅ȓyŎX�s�R�q�X�x��A�5����^�bd�d�@ ��bBi��<�F���elv��S,�gꌨ*��� �Ą�a7�$
���T�,l�րB�4���qr|˂̀[w��!����y�ȓ	>ژ:�I�es���.�(Y���ȓ_nD���M�8�%�P�ը�2�����cGGD�J�, �Rl�ka*M�ȓNX�z��߁	_$��jӔR�\���0���g�TE�4��c%��sC��ȓ_=4�RDwfe��KW+E���ȓVs�T[��?/����R/T��0��G�r�J�
aĐe��@�7rp��;��Y!	�01�A���S4de��S�? ���O�>+�TMc��	3LY"O~��#cP�Qy�tP�h�
N4Y2�"OJY���N� ��8�i@�dhm�"O�e#�AYN	��&ޮh슑�#"O0�a�k4m�~�c(ҳ
s�}��"O,2��D1,a3L�:;�Q� "O�u�L�� D��e�"Qƭ��"Oޭ[��/�>�D��RW
̊A"OX| f��&q�8r�M|<\�P�"Ol%�r�-%�uʢ�!4-"�z"O��pʍ1m��M�D�A � C"Oބ�IJ�,a��Cm޲|z��"O>�+�(Ē_d���'LJFRF49g"O�8�FJ�{A���*�<1�=�u*O<e�#���KO�M���f���
�'=�Q��#�o���D�r�ؕK�'*|H���M�5vјU!�>�&P��'��%� �!z$t�����G��k�'��G��%�����a��P_�eq�'�����	Ю6u�� ���I�H�0�'���Bl�=���1� ҕx^��z�'njQ�#�!=�TE�F(H�;�xd�	�'�0�ڲ R�,\�+#��?3���A�'��[�l�;ޔt钣%1�XZ�'}d=q�OT(+l.������(Bd���'H60���̅
�;�!V7%:&���'�jh�C���&<0Hpd��(��k�'&F�;�Ζ�5������$���#�'8
0��j�c�m��5p����'�,	#���d
d}8��ye�a��'�ӄA �"G>���mϚ{��IB�' �����C��V8��d	@�G[@�<�&�t����7P��A��x�<�b������(�i��8��ae/F~�<a�fG�`Ɇʧ��
7�N��ZA�<ԅ:S�6}��A�npj���g�s�<A�o1p�u�0
8�l$au�Pl�<��N1Rm켁`!�%V�p��	B�<Yq�D�06U�a)N�q�v�#*ST�<�E
�
A�]hP�L+"pP���P�<��ŋW���	��I�x���+�g�q�<7b�'Z���he H��b��Øm�<9ԅ��K�\T�F�ucd�`��!�yI.~�8�I�G_
���
��y"�,7Cz���^?B� tH�hܒ�y��7C�\����F�"ȑ�V��y�%SA.���J2Bi� � �D��y��b�)��CR�:����ǆ2�y��D+v�^���AL;�ptYrb��y���	�@ب��S�d��ac�B�y"	��j�Bd�T�^�`J�J񫑈�yRf�.j�1F�G�j2 ��֪�y"Ɏ�=�e���K%��M�u���y�fD=���S�H*O˒���I��y��$����hKS��� �0�y���[����$Ets�ّ����yR/�=��Ҥ�O.W2�4�_��yRf�D�n}��K�op �	��y�j�)5�n��FJa8��K�AR��y�Ȁ/I<�0eŔ�{�`��P�y����f1� ��M�k�hI��ˋ�y�oA'!>������dq��T�
��yR��zGJ�B��n��1����yb�?%�R �7.������y
� ���ЂE�'�X�+�.;��2"O0z'�T�[��U�K���6�"�"O�dxV��	�^A��*ɡe��I�"O�A�VgV�m��u��	�$DB$� "O�=��E�#���
--�\ �T"O���biQ4j��-�t� V�z�1�"Oaa�bU*�RP;6�� ��٦"O��X��ǆe=@
�k�=� P��"O�I��6l� A�0�
, �JQ�"O
a�� �Z����g�'g� AI�"OĀ�f:M�T-3�
�[�\�"O�����Ǫ?��^�D���4"O��x�
   ��   �  g  �    �*  q6  /B  �M  zY   e  p  �{  *�  x�  ��  w�  b�  ��  �  @�  ��  ��  �  ��  �  w�  ��  C�  ��  d�  � 
 G � � $ �+ R5 '< kB K &R Y \_ �e �g  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE��DG{�𩊺9hl(&���洠�H[HGQ� D��݃nĪQ��E;^ҡh�;���0>����t�L���:$�0z�N�A?������Fa��d���<�rf0v
���A��
B�I72���H�A8|�J�8z�'A1O^�=�;c�`гNO���7bێ
ޠ�ȓa�m�'�R�:�,6Ή�aLR|��ē���)	,b�ga\v�P�	E���C��%+�ؠ�U�.���0�ūYLC䉕q�(���#�/�m"2+׵��B�ɝ#��&M^�p<�رo�4�C�o�����-(��qW�R�Qn�C�ɱN�<A�0�ߔJ�H��"қy��B䉈~������Dub�ֶB�	�CcΡ�����	般�
�;o��B�I5�݉B�I�-/��{l�"{L>B�<NQx%��,:Hd@���(r��C�I&yp�	u�E�RI0����Z05�C�IlC$,�'��^b0z��r�~C�,���Ѱˊ�-�Nhir �&e�B��+v�qӁ��2n`�� ����C�ɐY�0Q���@�<�A�#��Q��C�I/'=�d��J�>+�"��9�C�I`|�y�O"H2ΡA5�S3��C�	]}�ѹ��b������10�C��8eJHjfE�p�^���֒h$ C䉌+����3�7J\6`3�Ԧ��C�Ɉ Ta�˜)��ۖH�!h,zC�#7�h����&���^:>C�I BDBuA"��>u%l4��>/0C�ɏs����� 
�>t:-�O��B�I
I�6!�ό�Q��-� Eη��C�I}�������9]��"��ޢG1�C䉩G~�z� ��w( ��pG��C�	OF�)��J�x^H	�H�[|B��E*ޘ��C	[S�UB6��lq�B䉶sE�H�,@$˳G�z,bB�)� 0��F�I$K1�i���?7>$j�"O4�����.:����EB<6�ڗ"O��f�?��X�����^)����"Ot��������� �J,��k�"O�lw���7�� 
��@�P�:��"O�XG�ۅ ��P5i3"�p$ش"Ov�i��ĝ�`"TE�"�isb"OPE��zhr�����rG&hJ�"O 0��-� L4���= 5��P�"O88�G�Oo���QF��v"&�C"O@MB"%b�m	�j�7}f�}��"OE�ƚ0rH�����y�pғ"ODp��܁;�P�ѩĦe�&"Of�9e��,���*	�4,J|�"O¼i"A�|���S��%*q����"O�+���GJX����W�БB�"O�iR�������x7�bD,���"O�e�4']QByS� �"�i��"O@ĐP�!ifl+PZ;!V0,��"Oj��J]1R�*�P��Q!7�y#"O�ݹSF ;�zh�oԶ B`�9t"O<�32L郳��)$ى"OT@;c���g�p���.[q�$ S"OT���&v���A̕�)jDM�f"O���a⑌�Lay4��&}� �E"ON����ȚT�PR��@$G�FŁ�"Oƅ����U�4��c�:m�$d�D"O�����b��8�TɃ�x�4tZ "O�<� �'����ɕ6���@�"O�q��O6�:$�Q6m�vP*�"O��b�-gA*����ԫb�^��E"O����yp44�R擄h�\M:�"O>�2��J�>�N-���_S;V	��"O�tp���vB�͡�
?=�)��"O]�aiW�lsN�#�*�:]lE�"O
����@�9�T�;�cC9G D�"O~1�"�(1�lS(ŗ���X�"O�ᇀ.K}<ݐ��4�ذ��"O@hp�(^�{�r�1�ײf�~��"O�D[f퍛^��C��Ո�40��*O<�7T����z�(O'�ei	�'?,�CVś�>�uHuK�3�x���'L�@��+���ű�1*tm�'-�؛�m��M���
BoŀM�
�'M~��s�Î.��L8�C(��%J�'H)�%��|<�@*Uk��]��'V��z�H��9YT��>u��m{�'����ıYa�u��Dʤf�r���'/|��bO""r"u�HQ)T��	�
�'cn{���$��ts��<t<�
�'x�dqM6��]r��ˣW: �	�'��0�qLB�Tc �y͓�w{�c
�'�(�$�Q�w��4a��k��`�	�'� �;� T�~�,�F��j�ޙp�'�`Z	�ұ��Z0#$�b�'1xR�B��C$�H	-N�/�n�!�'VHI�B�y�F�{"�P)�yҎ�,u�����E�:X��H�hנ�y�@���h�h���R��`21�7�y�ꓼGN��!� W�9�`͒3�yb�M�UZ0z����*\��"��y�a�H�v�B3����(V4�y��0a4t#1�W4��ax��Y�y���7B��x���/8��l��y
� �8���,�B�!$����"O(�h�톤&�jE��Hތ-.J]�C"O�9�se�������*\�"O��S1*��.����˘�|��x�"O8�:&U
RI �e��V�Tm)��'���'��'���'��'��'�<�k� D�s�jm�$jұ�ZE$�'�'���'e�'�B�'���'(4�7�Z��,SҦU�m�����'�'���'���'
B�'Q2�'�@�'
H� 0���P�\, X�P�g�'��'k��'��'&2�'R��'����"��'!�E�/�S�va1��'���'���'���'W��'R�'P 9:�fE� ה�kH�!| ����'���'�R�'�2�'�r�'*��'��D��
Wì�#��ư���'3��'�r�'hb�'���'R�'=t���ˉ�S�t�J<���q�'���'���' "�'�r�'6��'�x���Ӎ^���� �o�&��'2�'�2�'�B�'���'���'�x� �N8-�����P�G2F���'���'Zr�'O��'�r�'���'B�!#D	�1��Cwא#:����'MR�'h��'wr�'(2�'���'EQ�B�8U���b%��Ͳc�'�R�'7"�'��'��'���'�N�C!�B�]��@�1��x���g�'��'���'���'I�'`ӫ�iG�˒:���D8	��Bt�P&W6�ʓ�?Y*O1�����M����Ox�e�X�|�� 0�˞{�
H�'S�7�0�i>��ퟐ��GE4$U��7\�ZqF����	�C�an�P~�2�@���@��ʈ-��%Q!� Luc�L�!�1ON���<�����)Wܠ��&�v���f�g>)n�J�b�P��^g��<�z�ϛ	r�6�[�N�Ŏ���O��y}���ʛ�U8��0O�aD�d�6Tr�cT/o�\�Y�:O��	��?���%��|���]H��؏�*� �/��{d����(�D���CA&�I��
I�p�E&V�T���+	B�6��?�X�H�I���ϓ���q���+tB��sF��rUd�'���lj�j��1�c>mb��'0ޕ�	�Wn����.]� 0���.?����'-��"~�Vd6���3!n� ��L$�P-����j�����@ڦ��?ͧw^4ı��Ԩhz��[�M��?����?A�Ɨ�M��O6�S����W10C���Uz+�|���L~�O���|2��?Y���?�ifm�2 :U��h��|%$�<w�iUR�#P�x��k����SE��L�f1kP��5@V�$J!B�����Q��YB�4A+�����O��Ĉ�8e uR�
S���!A�Ui�І�$��hH� q$�"k�N~�A���$4"�@��e�+��@� 4��O��O��4�:���!����dR�
֎� ��RZrx�G�ϥ�yGyӸ�h;�O4�l��M�i�rY�7b�<9�b੤J��|[D�S1 D�ao��;O&m�R*`�����4�OpF�C!�w�@}�&�Z�Y9�u�t�N:}��ъ�'cR�'d��'���'j�RM��"��!76s�Z5f��x�B�O���O:�oZG�P����b�4��4��1!&�M�p�*���ܷd�"!�x2$}�oz>AI��립�'k8�b���')����3�Ġ�o�8$ˊa�	�A��?�Mk.O�i�OX���O��HcƆ,o��8�&@���F��%e�O�$�<I�i��;��'3��'&�	}�`��-ģG�Q�Fg�#9��������M5�iӰO��韈|RG�J��򁪕��c���K�D�'X�8lcq�(]��I�u� �ʟԊg[��� N"�Pq�CD뮑 ���:�f��Iܟ���ӟ��)�SFy�Ld�|A��+��mI��pdlH8A� ���B�&�dʓr웶��Ix}b}��!�T튬G\ JR,<>�H��cE�q��40����4����jt(:������Z :"��.�����N�8HR�4��D�O��D�O~���Ov���|�p�Z��<�Ǯõ3���A��(���@J>G��	��x�´�yw�I�Q�C��*RNN���R�6�W��)�J<�|���H��Mk�'P6��Pg޽k�$L��fЌ%f3�'r䵺f���X�Q�ؙ�4��4�����3?�,���Ֆ90v�x7c�;���D�O��D�O����Hܸ���'��K��/(�\b"!ן��%PPlϝX��O���'�6M�-�O<Y���M��x!aK��Z(Y⋟Y~�BB�z�z�p���<��d�ĺ����O��R�e^�͐�!/n�j�{��Y�b�l���?)���?���h���$]�� ��B��e��P���I"��d�Ҧi��ݟ����Mӊ�w��@�M	{�8:��5l70ݣ�'H��iad6�Ĩm��7�2?#�����铗v�^L���+lNLp@����"�c/O�=m�cy�O���'���'��H\:�v��ɜ9 l���4$��(��I4�M���%�?���?�L~���E�!�N�[�}'��\�p�شE��$��)����WR�\�ƌ#�֯7y�8Z�ʺ��-_5�a��'�:D�'�~7��<qT��t�@���.!=��*�/��?����?I���?ͧ��d��{Q�����Jܫb^Fyb2F>H,Q��q�8@޴��'��������Ox7�ΧN���PP@ƔWa����!J��m�odӚ�	z�2��Ce�K���yq��ߟ���:(��=� u0GG�V�QY�D֝d�~��:Ov�D�O����O���O��?��������ƫ
�@�%,����������ٴqt��/O�4lZy�)A �e҂	]98� ��K�#�v�
L<b�i$���O����i��	)A:���oǽ�z5iA+�'P��D�P�
���Ay�$sӚ˓�?a��?��5S�l���g���pC��%��)��?,O o�2@E4 �I�L��P����q�-@�ìF�Z��%	����XD}"Mk��5��z�)���V���
Â�/V�bD^A+>P[$Έ�,Lر+O���B�������4�p�a��5l'�9P�ݞL�*�(#�O`���O��D�O1�r˓��ᓭi�$�[fɀRV�ԪN���Ȓ�_�ܳ�4��']��\N�ƭ1MZi���ʇJ�.�2V@�B���u�Ʊ��+s���@�D��Lk,O<ت&�,4Ψr	\<%d��bg���'���'[�'�"�'���"1"1%e��kK� 3gD	�b�ڈI۴/u�(X/O�D$��+�M�;�X��T��8 �� P1�iB�T���'���|J~bdD��M�'��9PECJ`I�<��/ך��ə';�LvDHџ�iAZ�ؐڴ���O��D������Ȓ)U8x4��Vl�p�D�O����O��4O�ƥ��j��'�"S	7ö�Q���\��MQ �/+�OԴ�'�7�B���'�H�PA�$i�8��U�.aN�Bc.?Љ*N�D'��.��纃��Oh����� g\;R#� ��ƛk���
���?���?9���h�"����bBP�p%��	F�(c��͚�<�]Ǧe����_y�cy�����n%��R��D�y�t("��ˬ@��>�M��'Ǜ)�I�ƚ� :V�K.A��LH3��0Ɓ/qb�R(	�E�q�'�J6ͷ<����?����?!��?�A*��}�%ɚAM�8'���9�(������ן�&?���|M�X����7�֌�AlD	<�Ѫ�Ov�m��?�I<�|�D��4bl��'
S�@��	UEN2L�ɓ!�G���$�<����PU��V� �0� �hy�����W� ��4��l���������Suybbp�D���ORu�s&��_�.�6���\�l�"6Op�m�G�	v�I�M���'^��Ԣ$�,lJsF�>� yI���*�"�2�i���$,��1�O�Ҽ�'�
�}�5f��������?t���BM8�y��'�R�'r�'���	Υ�]C"�O>^�J�#t&b#��$�O��$��	FId>��	5�M{O>�E�&Z�ur���08L}��'C>S�'�6��ަ瓿���n�B~��0MV�d[���51<�ST�&sz�7�
��tX×|RW�����X��ڟ(�!��j�#��B�6!�q� _�r�'�I;�M{�j_�?����?y-�F�"�AL>TٌE��f
%(��6����.O��Dv���'�����<�Y�/Y -t4z��D�m��:�ɘ�V0 ��L# ����?�p0�'��$���Qͅ�B4��b�X�ӐbE��	�������b>M�'�"6-4�6�I1�-����g��x�(����O��DK���?�Z��Bܴ"�~�Į�HĊIB�3HP
��i��7�ĝL��7�`����!w�F���Oo�i�'���F�����fa�4�گ�yR^����͟L�I�����L�O��I��`Ga~����H�(��{���ӣ�Ov�D�O�?Ux������$}d��k�āBI.i�mEa����l�L$����?��k�EoZ�<	�(LoLH�`J%K�btoք�y��ͫI7D!���n��'6�	�P�	�n*A��M��8S`���*j��I����柨�'�:6�0Xu>���O��$�'_�l��f X;
taz7�D���<b�O��m��Må�x�etU ���Y&�L%s$��7��O�2��a�n�m�H~�B!�O�m���snڹc�J�`�V��A�&Fu�����?����?����h�����c����C��y�4˴�F[�������9C��џ����M���w^@��L5
L(��	�}ډ:�'x�6�ɦa۴�.��ش��ēq�f�C��o5��z�M�po
i�e��/R���Be'�ĵ<���?���?���?I
"���$U�T#�D��������٦��J����Ο�&?��1h��m#V���~����#�(=Ĳ��.O��Dd�@�%����)����w�� �uTf�RG�I�^[]	W�<��jL-6n��]����D8dhP���=<A�����,CJ���OD��OZ�4�X���V�!�R�5zk�m�$AC>�`��	dd�,y�&⟜!�O�Pm��M3�i����'I5�@a�ѽV����@�ɟ;���Hw/�(z���L�����f���5(�F�œy�
� �~���	ԟ���ǟH��Ɵ���E�8!���L�0���"��/�?���?yñi����OwB�y�ԒOZl�P�Ϥ��HP���@�܁���v�	��Ms���T�7M`�֕��ئ���q�D�i\�Xp��g�I�h���`ι�?�%,�$�<���?����?�` �$a�d��#�ve��CBe>�?����D ަ���J�����	���O�8�`Ӡ�&S?�4;r�P�:� ś�O*�'"7mEǦ=pI<�O~�	g'T^��pG��6��(��Gpp�9�Cʹ��i>EI$�'�VT&�(q��T��a����7�ϟh�	����I��b>A�'H6��o`(�4���kK~D���-Z<^E��f�<�Ĺi��OfD�'o 7���)��I�`��C8c��&*�n��MK���M��O�EB� ����<� R �rN�L�D9�`��;=>��f?O���?��?9��?)����T+`�"3B˚a���-�3?��o�4Dd�I��4�	S�������ˑOM+L�fX��*$e�2�㣭��\����~Ӯ�&�b>M�#���͓ubp�@�8Қx�i���Γ> ]�b��OH	BK>�*O���O\��7���N̺�f˲B
6ɹr��O����O���<y��i,TK3�'���'P�cq.�:N��՚ba���������}}r�@��{�( %�Xw�;9+��B�G/q{����+?�n^�(S���K���'8W��J%�?�sh���J,�7�ܨ3��z���?Y���?����h���䔧$O� ��&NŒ);J fiV�$ ٦	Ō���I��M��wM^̑ԭ�>\a���Uբ�n��<���i�^7�릕����ɦi�'(Xu�����?�Ĩź+�F��Wm�;G�V�{�#��'��	��I�����ܟp��?�����J,Q�(ɢ7	&	��'�+���6âm�����	n�s�����~VTµ
��8�Y�������4*����OY�!ႏ�%���B�NG�'��1�n�W��4Z�l�G(X�Kk�l�{��sy��;�>iJ`���VL��#���Lb�'�r�'��O��I�M���L&�?)�(]�T�>���,�B琥���%�?y�i9�OJ��'e�7�
��YܴpsT�;�b�2��AsvGN�p4�u�X��MC�OT��H؝�"&%����
(��O�v�*�Q��H�p�c7O����O����Or��OR�?1#�O�2
gT�Z�h]�g�R�#�$�I���4^9v��O 6m'���A�4�Ы��,n�\�v�@ �M�N>����l��?)��Ħ���?!D-<6ib��c����K�D�99�ʍ�f�Or�	J>1+O��D�O����O�X2Wk�O��4bĪ�{sm�O0���<�Ľiۊ����'\��'��S23� ���(BD�aʔ+��{]��̟��	M�|
�F�\�M�+���ܑJ��H�am�<�TC����9*O�ɓ�?	��!�$�
J����-�7P�� �D���d�OD�$�O:��)�<�f�iTP�ƥ�(�D48A`Eo���a��jXb�'�L6m4�Ƀ���ަ����<s���3��R���Q�W��?9ߴN&� Zش��޹qz���',��ʓK<p$₉/�~��cJ+bR�8����O<���O����O��Ŀ|r4+�+�P��%m�,X�æ�%b���D�r���'t���Zئ�]70J%aѨ�&��s���*`4y۴-Ҕx���甲䛆?OzxH���m�b�,Z2�&� 0O� m��-�?q3J+�d�<���?�r/�mL�i���O5'p�SD�	=�?	���?����dئM��K͟���ڟt�ud�1)��C�N�)<�$}(�,�W��Z���ԟ$�I^�ɲ���B�ɐ��B��N�A�
�`	`�҆� �t��5L~����O�5S���h@6��u�œ��<��X؟��ןD�	Ο E�$�'�&�9�E�V� X3A.��$hPm�v�'�6m�M'��0��4�4�L�"��yd�	�F��t��6O�!n���Mk"�i��K��i ��Y�}���O9���� �:zfLx1�H7��� ��l�Py"�'���'tb�'�nO-vG�)�FD�'^�����J����
�Ms��_��?���?aK~�����C�Ѷh� 0!WG��^�%T��I��M#s�i��O�)���).c�}�uN=�� X�[9��Ǌߧ_/��c�|�F,�O`��H>.ORݲRL��S�h+��X6�8�c��OJ�$�O�d�O�<)ƽi���8��'#*I�t� �Pd��*Ɂ�*��'P6m9��>����ҦY�ܴ���*�";�ν��)��xE˟ndM��ij�$�Oh�ǍQ��'j�<��ԿSr�`Jx%P��&s��*�T�<m�iy��'v2�'�2�IN�}�๡I�R��I[v��=����?���Y��v��Qr�	��M�M>��"_�$Τh�� �=�x̹�gɤi-�'�r���$(�	؛ƞ�`c1*�![V���e�W�D�����W�,�6Y��'ixA&�L���D�'c��'�D٨�JcЉ���2HG.��'D�U�4��4I�9*O��Ĩ|��#E1>��QbSfɸZ��Lb3$�]~b�>a���?��x�O����4��pi^!�t��N͵/��ؐM���2�O��i��?)d�0�V2_��kb)��z��i�IG##D���O(�D�O���<�W�iX�%ìKn�:P�C��D[�'-Za��'��6-5�I���OH��2c��`:��Q` �2v]���O��m���lZu~��o	������Ovz���%.���,�#r�܁�'��	���ȟ��Iҟ���t����##�n�C#@ ���Z�cT�
��7m��Hi ���Oj�D?�9O&�nz�aq�G+1���#��?�p�2�������}�i>����-����L@ЫK�^�C����7����
��N�O�rK>,O�)�OƀC�C��	PiB�W�,�T��O��$�OD�$�<� �iѶA��'@��'ǂ	ԣ^�@�Q��IH�L��@�D�j}ҍ~Ӏ,nZ�ē2�tp�.m�푦'�L��'ܜ9�C�[�+a�h[���TA�T[@�'t��اh�!��X�&BP6*��PhV�'�r�'
��'\�>����P,.�c�/��c�����ò(lz	�	(�Ms�ŕ3�?Q�R��F�4�\�u@ƾ �rыaKϜ25� :Od�oZ�M��io>(ҵ�i���8m:�J �O�� PiQ���<9t�Y��| k��<��<!���?���?����?1���`��(Q��A*m�d�DM�����I�#K��4�I�%?1�	:t��Y�Q��xN.屔���p)�O�oZ�M�g�x���ɜ�G�TX�6*E�T�0K�o8�J X�@E&�剾i�
��'�,�&���'�Q &i�"-NJ� t,��~n@��'��'�R��D]�(kڴFS��#�mqȨQ��4x�a��<D��ϓI��&�$Gm}��'��'n��n�`�J�*�a��r�(�&b����� ���3 �$�����yp4�͵ ��xs"�G� ˄��0=O��D�O���O��d�O��?ŋ4��5u�nI��Gx���A�|y��'6�\-;��S;�M�H>�`�0,���{�D["Pw��v�ۖ���?��|�4H�>�M�O> �3��~U�9eDB�GS��uK]�1������TF&�O���|����?9��)sbź���~-L�0%'������?�.O��n6u�`=�������E��c���,�����EB�P����@B}҄`ӛ��*�?��&���W\�[v'I� ��B#��*lz�x��Ɨ�ex%����+�ٟ�	D�|n��	������0�d��jZ���'���'���DS��:ٴ�<��1NՄH�Ĝb���-���"�A��?��%p��\_y2�iD�5:�f��
:��qd�)��! 2�zӐo'�f�l��<!�3��Tp�蟘H�'ʸ`�	݁F��]���\�5R����'��	Ɵ�������������Q��G��p'恹#���l�(�@7�	#.�����O��D:�9O�Xoz�i���ҁV�kQ������DA�ޟ���p�)擂y�t�n��<q�N>f�� h��#完2s�\�<q�*�{f��˨�䓌�4�4���^`�3�[�`�P��W��''����O(���O��W��F C�r��'ibn�#JQ�����C� !����>��O��'���')�O^q�G��E��5"��*|�LPz���,k��=*g���&$�9+`�&��� ��36�^�sN4�Șq��G۟�	ޟh��̟�E���'T���r>�AY�7*	���'��7͞`����OP�l�v�Ӽ#��ç�.$�7K֚=9b%AN�<9��?���i�,��a�iW�	�pW�O>Fhݦ$c����:_����$��A�	{y�O���'�2�'Sr��&\l���E�)��}��f�$"��	=�M�����?���?�M~Γ�	�� �aK���aB](f�޽h%P�������L<�'�?��'~�l �F
�<mIU��a�������#m�`�'��ih��H���|"^���� ��hp^AiQ�8�x� 	������ğ��I���Ly�kӚ!��O�1���j���Pǂ�GQ�y�6O�TlZ@��}��%�MC$�i��6-�,Kad� ��q |����pN�Ԣ��v�.�hD�=v��|!K~:��8`�i�qc�(	$XY¢�3M$���?A���?����?9���?a�M�����8�!Eb�'PH���%�	5�������?�ʵrb7:�I�WۄU��`y�͸E#.L�k�,I�� ,�>�6M:_��$�O����h��T�g� �ȟ4h�kQ"�� U��s��@����)F��1B+@�J!2�'���A�'iZw��	��F�$�O0 �B�,<���E2Zx�Z"�O�D��E�<�7�'q����'�?���)O�{��c&���&pgB_�7J��ӟ��'��6-ܦɯO,ʧ�b���+1X�j��يy�"E�k�<H��ݹ%����'z��J���8'�|��֞-�d]����c���# 풔q1��'���'���Y� �ܴ4�ڹ��W5^�h�栁(qZ��á׫�?���9���$�C}��c�ڡ¥��)D�z��2�GH�����I�U#�4U����޴��d)@�<����O�v�hj�PeJL�nX���	$_,@�����O��d�O��D�O�d�|b�&ޢ>�Ьh�hQ%BFVȩsK +3E��� >r�'yr��d�'�t7=��1SAʍXvΠJ�jŗK���ab*�ߦɱٴ7�����O\��]t��6Of�qK��%Z��#Wwt�C�:O"��-���n��~y�Op2K��U�a��3A�B[SK�'K�b�'7R�'��	��M;��� �?���?�*��&Zr(��D�m�^q���̡��';���?�ٴl��'W�E�w���s����"�5���#�O6(7)�F1�xs�f#�	�?	���O�(7/4>����r&��(�8��/�O>���O����Oʢ}b��r�X}qǒ{{Xm9���K�]��$?-$��'O87� �iޅ[s����(��j[�]Op�2��}��شBu��w���i�im���,���0$$��P��Ak�5 ��CQǓ3 �zD�l��䓢�d�O.�D�O��$�O��d�6�^�y��ø�HEEɒ,>�5J��ES�*I��'$�����'�E��'E%-11*��&f�Q�v'�>���?q�x��tAˊD:ƀQ"Q�X�@��Dل�v\JkL������!/p��0�H�O|�M���3
+�ċ�C��5���?���?	��|�)O��lZ�9l�e�ɍE�@�ZT'ÖL7���m��*�D��� �M��j�>���?�i؄l0-��K��R�-�@�zs)��6_��<O\�D(ro�����i�֝���C̖�S��J3A����4�y���	�����ܟ���쟈�:��؉2�铈��p��,�?���?��i���Ocr�p���O�m1N҇!vj���'�13��jǊ�V�I������?�B����Γ�?y��Sx�? :�W�Ԗ9ؘH7;5��Y�鑿�?᳠-�$�<�'�?Y���?A�(f`���C{��zCfJ&�?!���Ҧ�1�(���������O��tQs���\�1�V.؊�i�O�4�'x��'_O�)�OT�@�@"- P쨠솝'Od���̰&D<�����I�?1(��'�$�����щB��ea�ޖUn��0h͟���ן@��ӟb>e�'9�6�C*ڸ�щ�� ��-��� L@�e��O���M�?�X��	�s�l��*�L�Jf�� �ɴ�M����M�O�u�����zK?-���'ut)(AS)�v�襪`�h�'���'�"�'A��'y�@��Hy�j��F0�f���a�K>���	����@�s�h �����:e��)�E_�s���F���0!ҿi�*�O�O����Ǵi�dN��=����<t�Q���Ri6�$߃7*��{��M~.�O���|z��qaf?&�B�C�� 2� ��?1��?a(O��l�B#X�����I�eX��%� 6X���Zb/I/|  �?�P_� �	ޟ�JJ<����o��P�-ŔcB����A�d~�+Z�)l�xpD�5��O~���4-�BAT�vU� Ȟ����acoѺS&��'���'���ş|����t��U!ѧ~)hm"R��ğ *�46
!�,Ojqo�b�Ӽ���8(2�@���]��Ě�<�3�i�86����ApD�ʦ��';�bukH�?%7%�)�F�i��ʤ��9D@G�hR�'��i>e��ן���П��	9(�hy��-�*0b�-A7	O�}�|���9g#<q���� (�(��蟨�I��MS*�D����ܑ7�O*_�\,�A��~��	�'���'��O�i�O���²f�r�"���5*�ɻ5��+�Rq�L����ɻ/���v�'�='���'�������9���	栚UH�E���'_��'3���$W����4yȪ��%�Zͺ�ǣ�8�4Aı�JIS��x�&�d@}�/bӦPn�M��ёyH0y��#�<�DA�i��ȁ�4������2��LF�����_�@&�V��L�w�M�IQ�D�O8���OD���O.�"�S�T˰��vB��5�f�kÊ�6E�μ�I۟��	��M��n����٦�&������a3 ݨVm@�#I����x�I����i>!��!��-�'� =zd@	X\�����d�щ��S�#��I�OX�'�i>����t��N!��Ņ�[d0+�/K#�J���ҟė'�d6m_�&ے���O��d�|�u_�4.ز��0�,�DH�N~�>����?iK>�OX�A��	�m L���.��}y� `����g�D���4��ͫ��7�ғO�p4NB��jue��!x����O��d�O����O1�L��6�O�4��*؍~����%	{�t���^��(ڴ��'��ꓥ?)�d��O'�KՏ�r�2�z�G���?���[zhP��4��$�	.�z�������i�ě�F-P��QF�$pRD�|y��'��'�R�'d2]>��v�w�|���'�&4Cݲ��M#�hگ�?����?�K~Γ;��w	Yy��BG:������o�����'��|��4�
�F��1O|���ቦaæ��!FǺa�f1x�6O���X��'�B�&������'����v�0,�D�gj��P<Y��'R�'�bR�0�شP�*����?��z�|a���e��*�⃥?L��R�>��i�|��%�dPyj�Ȑ��_~@\�5�UO9�ɿ���&i���-'?�ˆ�'��	�I3�\��4��Y�I L�B����	�����͟���f�O���L���!�8[��Y��4Y&��dӂ��OP�Pڦ��?�;n��XQ#�?�h8���Pע<ϓ4�fey�2�m96m��<���jo�ѫU���X��Č;ph�c�G�,t�Yۖ!N�����4���D�O����O��dF�| 2��X��hK�� �T���F���@LuR�'2r���'K�3��g6�؛wOV�dk��in�>����?ӗx�O���O��%����'#�V�����,$��)f�҃ApJDr�O2,�Q�X%�?��;�D�<é�t٫gk�kx�Jr�� �?���?����?ͧ��$Ϧ5zwG؟� ����r���5��Tq$�q�ʟ�A�4��'����?������b*��mד?����AG9�P��d�i��OJ�X"����'D����?m���}Q d΅����ɉ�0>��ן<��⟈�Iǟ��J�'C�H�Aw��|y�-Y(+�f���?���fmߟ���禕$�Q���@?�M�g%�.�&EJ�R��=_�Km��I�"�6-5?)��\���XQ�`3#���&�c��TK��O8�iI>A(OX���O����O�X��H8�a5�i����O��Ĥ<q��i8]�E�'"��'��S�TM
�+ �]�nT�f qb~���	5�M�T�i�O�ӫ!�b���OE<) ,��j[��6���(YGμ��Y@y�O�l5��dJ�'���pڦ	ތ����"|�p�'��'�2�O���>�MSЬ�B��Ћv.T%7�f䒆J,y�����?I��i��O��'2,7�:|,r���.(_����G��oڮ�M�3d��M��Oz���/����<�7�a6���:?�A8f@T�<.O��$�Oj���O��$�O�']9��i���3�\�ÀJ��\��W�iݢ7`�O>��O~��8��QԦ�]&����#>��ف��	0�v��4-`���/��ɐ�W}87mn�� Z!+��͑������b\�"�8O��AN�?Q �<�d�<!��?)c])y����A�-+ӾAQD�N��?9���?����������џ �	ʟD��JUh¬V	cސq"Nf�gC�I��M��i O|9H����`��i����2���#���Ӥ+�?X��d�%G}�7Z��G���h�QZ��k"��G��`�`jП��	�8�	ΟE�$�'�i�+�������n򘙪��'��6͊�0X���Ot�m�|�Ӽ3 ��81$�$��L�<������<q#�i�b6m���Ԯ馭�'�L]2s�W�?	�,�F�T)Pǩ.�+s"��
��'����<����	������c�^��C�v��Q�a��(�@�'	�7�5]��$�O���)�9O�<:B;��hqL˖P����`�`}�`�tem���S�'g5� ���-@�D���JF#\X�j!��	x@�Q.O|u(���?y�'0�Ľ<�1O�#������+)<���E�?���?A���?�'��D@��ݨ L͟��R��,c"dݘ��	A���K6 �ϟTX޴��'������My�x\mZ�n�h���N�Μx�M�3����R ��Γ�?�v�N٪���������h;&5ٗ�D'EJ84��	D�D�O�D�O���Od�$ �S4Z����U��Ye�l`��%&DU����D�I�M;�F��|j�;���|�TQ$������"\�p��Ŧx�JO�mZ��M�'G��ߴ����)l��ciѸ7Dh0�
x����M�;�?�q#-��<A��?q���?A�`!}����,�
�+m�g�j���O�˓0s�֊֘B���'R>)��H�0H㴐
����	zO%?q�X����ڟ(�L<�OV����ؘ Ϻ�����`dfYV%�1P����	��4�� "����O�A��)�3������C�D���*�O���O�D�O1���S<�V�Ih����Q�
�J�8�cIm:u��_���ش��'�8��?�'
�39p*8aǙ62(���sB��y�i����5�i=�	�8���C�Ov�є'�t5#� ��~�̐+�G��u�f�'�Iߟ��	������<�	e��凹}���	$GN&��H(�NְM&6-�%�����O��d+���O��nzޙx�o� 	�Y
�*��-:�9j�	�?�4J�ɧ�'z�e3�4�yr������Q�D/���Pv���y�Kڼ�H��		e<�'��Iϟ����
�\�
�<x ��0�C�mE���	���	��'�7-�8�$�Or�W��b� ��9�Zx��ˆ#a�t�p�O�o��M{��x���:y�������=a�E�5ǁ3���N�z8T�K��`�`��|DA�g���Ē��F���B(l{`�9���-�J���ON���O��$:�'�?)�!�!R>����r!����*�?��i��H��'4�b����];>s�(R$�`*�i�(5h,0bf�o�(C�4/��
m�LSC�h�P�Sh�]x�������T�������������C�����D�OR���O�$�O��$����`"LB"x����`˓x���c�5p�2�'�����'�B`sTg]�aB�i�&�	h@F󱃥>��?!J>�|����3HN�p�ƥ�Ւ�m��0��H���~~��&w0t��)}�'u�	,n�n�tC�;$��Da�H��	����	ԟ��i>��'&6-�v%f�D_?` T`wGs'x���_5d���Ʀ��?�PQ��9۴^כ����8E�J�m.	�"�Ń	
�8�U�*C4�7�|�@�	G��1Q��O�\�'J���w�$D�d!�9T�@0��Qª�9�'��'�r�'�"�'u�Ԙ�B�� |�ڜ��-�q��,�O��$�OxmZ���'�T6m'�DI/g� �x`��_d̠�5��ِ�&��S۴m�f�O��C�i����O��2f�?z�tթ"��l�D���_b_���-rƒO��?����?����
�;�f�Ni �k�e�<Z�f�����?�.O�mo�=#U�A�	�����o��l�8��cV�P7j��ږ�߾���b}���܈oZ����|��'%������ Y@���<U퀭�S��UD⅁b�7������@�ғO��M6n[҄P6� �?�΀�2A�O����O8�D�O1��ʓ��&ܖs�$:�$�68(��2��� ��,0W�'N�Hz�⟐��O.�mZ������þ0����&k�vl���ٴ^���B9ߛ6���`��2���kyy�ň�v'��y`�6 q���5�yRR����͟X��ܟ0��ݟ��O�xe�F�P�P��dITB#[�8�+ rӈy���O��d�O`�����HĦ�%��p˖ʗ&B�-��h0e��i[�4؛��0��	)��6�g�T����	h�s$P�x钕�j�� !A/<Nb.J�Iny��'C�� s$�u��7I�|��Eѷ.6��'���'q��MSr�����Op�y�b��ɠӀַ4F�h*��7�����dMæ����ē:��MR ��-gQ��k���V4�'̢���Y 8 (ғ�te�ܟ(B�'a�[i��^vJh��+��'(�Qp�'��'��'O�>���/#�zu3V!�@Ɯa��B�Z���	%�M#QE�3�?���
K�v�4�Ҩ���¼c�� ��B�Pfh�31Oj�o��?�ش4	�-��4���Prd��'҅Z@���F��|�!�R�LJ� �4�D�<	���?����?A��?�֡�$a�C���0�F���F�-��D���!qj�֟��I̟<'?��	u�����!�%*q��"O�
$R�:�O���{�$%���ٟ��V��� x�J�-ȂK�l��oGr�0����ʓ5�5��$�OP J>�+OJ4yaO��.����C��	�ֵ�BH�O����O����O�ɵ<��i��(t�'��+����u�D��XxR�AQ�'�P7-�O\�Ol��'"�'��Y'�4L��)J�6��ds�7]��i���Of�bܴdX���"?������"cĿv�$�Ц*��:��p�Ԯ��<a���?q���?!���?	���&òq���C&�RG�rec�"n��'�`o�L�p3���W��5$�<��K�-�N����Z�%[�kґ�ē�?I��|"�����M��O�H�	��.���2�i�!P6����J1v�!���T�$�O���|B���?y�<�(=���W�>n�����$�my��?i*O,oڽ����ҟ4��R����{�q�LCɐd�Q<��d�E}b�qӴ�nڇ��S�d�8P��mâǧv\� jt&��బi��6�z@*Q��S�;��DW�	!%Q�]�"g]G�\�+�+{�0|�I�����Οd�)��Cy��lӬ��V�̤BT*UE֎Xi��;����@T��
6�����NyB�iG.Y0@f�%r��
!c��3��Pp�r�� nr<n�k~��r���S�3M�	6s$�%;��Y�"�D� ��8���ry�'j��'�r�'
bT>�椕(k���;��C�6�A�qd�<�M��Dۿ�?���?����cf���/7g�8���$`��y��&�,U��nڳ�M�2�x����G4ٛ�9O<��D�]��$��퉍O�TH�2O�ɐ�H#�?�� ��<!��?I��D>.lµ 7�@64�89�׆� �?9���?�����Ц�SE\y�'�2�C�?��EfC�%� �H���Fc}B�i��o���?�d
_D�xaX�X& �o8?���G�F@^�P6����'TDL�$ނ�?��a�	J�͸M.E�P���<�?Q���?���?a����O��1DHD�YUH�
�N?L\��Վ�O�Dl5Q`ٕ'��6-�i�mk1J�,ɘXC&J֕D�8��z����͟|�ٴ ˰�
�4���%"V��'V4�Xd�ԑ��$�L�V@�]X�k3���<ͧ�?)���?����?�aᒮ?���;�a�w���h�T���Uͦ}z��˟���ܟ�'?�ɠ*. ����E�2�[��B !X��*O�Dq�%���^�I��ؔ�����Q���ERsW�M��LaP��l�㞪�2�HX�	kyB� :UW���(�>���17掖w���'���'~�Ow��<�?q������x��Ũ9�PЙ��M>b�E�ȟ�۴��'��ꓜ?����6o�7s��Ũ磐*$��!���}FP(�i=�I�W	�K��O>q���T�}F������|���
��Y�o��D�O���O����O�<�8	aP��ʘ~Ru��O�R�ލ��ٟ����?�p�}>��I2�M�H>96�֏`n<�R��i��I�V�^�gB�'�7٦�ӵW�]lW~Bl����-�RB�����+�F=����0Qa�|�X�������8���ʐ5� A;�i��q;��ӧ�����	sy�Dj��bRe�<����򩈤��H�ć�F���m.*������d�O
��d�)"T,Z.���H�j2?��E�cV�C�EP��{������͟,�|B��5R)���#��3slɪd�Y*�R�'��'Z��R���ܴJ7&=C�I��[,E+GK� &�L-I4�3��H��?qG[��o�;G���C�NG�z4-C��B`�r�{���M��@)�M��O�%��c�=�d��<��i4icА;��P�B��=<L%���$�Op�D�O*��O����|r�`��Px��h�d�y:U���,"!�V��5i��'RB����'� 6=��eCRÉ}��ZA��h���*��a1���S�'5���۴�yb��,r@�+���-ԑ�pa��y�bE����^�'A��ן��ɉty�d����*d���aE�Z�������Iɟ�'�87mˆ@HB�d�Oh��q��0�Pϛ�)C`��P��x��O4m���?�N<9W�^gYz����HR��� �����
2#&��ϋ;^��:��;���%M����v-��%"*�� \� ����Of���OF��7ڧ�?�@� S�Bhk��:%W��3�$�$�?)��i�>QS��'$2+o���杞~��R׌70�T���Aܻ,b�特�M��'P��IU�e��V����rB\9-h��K^>�Bb��L0$�D��/i]��$�0�'-��'�2�'�"0O&��Q�dr:c�ڟ�R-��T����4+o�q���?����䧥?���R:y(�� fs5N��m��l��矘�����S�'S���7O$���K�p�,M�D�%��p�'����ß�ᔔ|�^�(5I�	�
�I��E:���p��'K��'�R���DQ�h:ݴ"ﶼ��qv>̓��XPP
Pˌ�;�z!�jf�F���Z}�'�r�'�r(�dF�=	� Q�cBWzp4%A@Ñ�X���=O��D����x��~�	�?����l��v�[.-����㙂"R��I�� ��Ο��	ğ0�Iy�'w�����$)$Þ=��b����I��l�	џH+شE���s/O�9oZv�I:o--��C�+�.�+#NV1rT��'����ϟ\��>_Ԛ�m��<)��u��8r �L7�T���"%2-9�D����Ծ����4�$�D�O@��H�Tl�h8�,ʚ|��|���B�2��Oʓ2t��P�6Z��'r2R>𐫀c��4�Q;'����5?	�Y���I��%���ϟ� �Y�v���f�ZY;6�T6�,E@���B� S�j��f����?�	��'�V�&�X�ᩆ�T�q��H:K�&D���L�	ޟ4���b>Y�'� 6�!%���`r
1O�lhs��0R���3�J�<���i��Ot�'�B�L?,��e�g�I�m�D-��"t2�'�~@�i��I�r��IrB�O�!<�����7�|R�d�����d�OT�d�O��d�O����|J�jͣ'Ep����	,Y�@y#'�a���	�7B�'c����'��6=�d{���./"`�SJ d4�!c�+�O�� ��	I�946�n�\s�D�J�@<9s%��J2(a��u�|���3R��RF��Vy�O�2!�B��$g��'�)Ӎ	}4��'q��'��ɸ�M���
�?����?�D΁18�T��o��" �C�d	7��'���(��ӎX$��zN]�P!6Oͱ	���#M ?�BL�C�"�����'S��D�2�?Q+Z�ځ
"`~�a��?9��?i���?9��i�O>��1�T�)�^PX�	9m����k�O�En�%8��(�'��7�=�i�997��B�� �4k�<4�|�cLc���	�����!CC�n{~b&�4���Sܔ\ɤ�@,b,�,P)֣ ��(rѝ|bY��џ��	����p��֗5�Z9*B�A�<�%�v�eyB,m�Jp��m�O �d�O��󤍮AZ����P? �Nd@�K�P[���'�r�'�ɧ�O�x�#Ù�,5N���̈&J` ��A�%����O���t� �?��&���<!�*��p�v�06_	O	U���I��?��?����?�'��d_ɦ�i1��� ƶ:�NQ�@NC�`�X봬r���۴��'����?���?9��̘����dȎ<�7��%)j�%�޴��$ހW�f�@�'��O����n�zV�Y�Q�(*�@۔�y"�'���';B�'����P��B�(4_�E��ǋ�bc��
a��O����O>Xm:mM��'a87�"�d�CZ�d(�σi^و���w�|��'��O.f���i��I ^״HJC�.4l~E*K�=�~�0D�	 4ab�D�ay�O�r�'��cXu�m�G�",u��8����)��'S�I�MK��պ��$�O�ʧT�޵��X�?�4X�U�Hi[Tn!?�V_�h�Iڟ|�O<�O�4 r�F�v�b�#�:9���WH�4GZ�	�a�*��4���+��RD|�O����E��F�>�h�L]"l�H�OR��O��D�O1��ʓ����,Z!��
:�X�����=����W���4��'�X듄?Q��_
J��iF+ە�:M��.��?��h]2��޴��D�+TE�������=$���Z� �xd��n�L���iy��'���'���' 2[>)PӈG	։��`Q3b�� ��$�Mf)���?q��?H~z�u���w@�Y�c�
��8�#��(x��xY�'�B�,��)��,��6mp��q�d�&�1[�͌$��b�t`Bd��D�r-i�	vy�OBr
Q'�*�K���b�!0��֕�b�'Sr�'��	��M[��J1�?���?!Q�������P33O�� EFC+Z��)�h}�`wӎ=o����x�C/L�	��A�B��͓�?�`@ې?����+��$�����C�6�$י��(B��r@ǯ+i�!�ēL���S�)6:�y���Kx$���Ҧ���gyB�c�l�杇�2����G�D���{�����	��M���i�7�_�
�7-z���I;FQ2,{A�O�2x)"B��3�r�3!�!T�����D�ay"�	8`t�b�'MA�X�tG�Uަ�k��fN��B���|�R���5�>���R�	@�bb�&0�����M˳�iPJO1����f��\Q��Ն��::�0��G<}�M��ɲ<�� ��-4��W��䓬��R�z���1�敧`�Ab6�Iefa|b�w��0�t��Oڌ* Ή�5�x�б��8P.�;S6OНn�O�!��I��M[%�io@7MF�8x�!	�n'8�08sӨ�O/,1@6fe�B�Ax.����\�{I~���v��c�پ4���� �M+z����?����E�J�H��
s\H ��/�����O^�m��2!��Qכƚ|�I�|�$4C��(�1��i�>��OЄo��M�'z�ιK۴������P#����B��E����Pڑ�؏�?Q�=���<i�ZE	:���⇙Cc(�Š܆|(�"<�R�i�*e�$R�,�	F�d��=`��<��C�8d0��8��D�Dy��'����)�T>�Z���EEڔOs.�tS�#F�E�����`ۑM�D����������і|��8i���S�);6�R�ccB�:�x�
aӰ@勍l���U�W�@Q�,� 'U����O6�l�U��X-�Ʀs�MO=
� ��D1
KfĲҠ�0�M�g�i/�)!�i��I<�� 0�ODf�'���S�1ng2`S`�ϣ&�� c�'��Q��:��K.|D�򠝥yL0����_��M�S����$�O�?]�����A7�M�%�G�	h��c��%Q��"~�h�%�b>�k��զ��%k�F��,�:s!�PN�J�ɁŠً��'*��%�ܗ'p�	�=�u���<|m�""AH�nBZ�����	B��,�IퟄZ�� z���ȏ�N�vĊP�Si���	��M#a�i<>O� ^�#P1I� ��E�0>͚U���A��K�p�F�ūQY��r�2��˟�ò*�({�t������@�zB�.D������2{�Ƒ�acU�#v�IQ�����4
�̨)Odl`�Ӽ��f��3�|�j�dɜ�,�z��C�<9�iM�6������'L��	�'+�yXŦW�?�Q��S$.�ʄ&�*k����C���'h����Iҟ��ǟ��I�Lj<�c*O�x6����s��'�7�&[�4���O��4�9OjE�B�ʅ��@�t��7��Ȓq�g}��'2�|��� �)�\�K���VWЀ�&��P~�%a1����B+���c�uA8�O�ʓހH��u�1䥃�}��1@��?����?���|*(O��mZ�L���Id,(p�#;T��u3B�k��	��MS�b��>����?I�\�(Q͐�3�j,����9@��H
XRpXo�c~"�[
I��E�cܧݿ��@	63#�4:M,5�8{���<9��?I��?���?!����T|��AB�2N2��0c�4i^�'8Bgz����5��<��ix�'U�p�vL�s��0�l�_Hf��|��'(�O�(�{�in��0�*����1���$)MT�J����W%"�/ZX��ey�O��'�r��9@@=���W3*���;� U���'o剖�M���V �?A��?�(����r�N��^t�bm��h`:�����O(hnZ��M���xʟ�	SoĞ3�t%���-o>���@�4���i�L"k4���|�C��O��pH>Yы�,rR�C
^�<v��¬�?���?����?�|�+O�Dn�+�ƸY#Ϛ�q҈ز�O	�8�xHL[ya{ӆ��.O�7��1�f�yC�˿'8li�Q�`�mZ��M#k̛�M;�On�9S��>��<#bV�P�D���=H�i��C��<-O"�$�O����O����O�˧M+$�z��l����FK�Ĉv�i���p_� ��g�'F��w��X���J�:C� +v�@�x�(oZ"��ŞdGĩX�4�yb˜�*� `��)әKhંA��yR 4��MX7a��#(�0T�҇����r�ށ�H�q�I�p�H��2���Y��	�i�,!����BM5���SE�_����@c�'$xDb�j��j8��+����TY�跅H6����(1�sPU��[W� M��t@�@�RW�Q`��J�� P0�+ON�"�I��@O0��p�B��,}b��4%�
m�a��٬
H��(��t'�����L���J@��� � 	  M�W�&B�Z�Ȓ�(�R��Km��8���)�Ρi(L6^aJ����C)�1��ie��'��Iz��+L��X��E[�5h�%�!j�<�d0�d�O>��Q�ݱOf����H$VѸ�,�9j�<%���i���'V�I]��aட����OR�	ڷ_ؚp���C�ɺ�됦\9^�'����៸b"�S�����͊C�I�C��D_��� �MS)O�����ݦ��˟L���?Ѡ�Ok�ÀD-|�C��&({lL��J�?؛��'I��^��O��>�fUE�ҵ�+��v��$�6G{�`t�(����������	�?K�O�˓,�Ƀt�޻#x1��c_����S�i3�l�f�d2��֟�: bЪؾ�uդ	�Fh:�DU��M{���?��9q�*\��'�b�O&4����+��X�` H.��C���F/1��O\��O^�DD{ޠ:'��*��u%��^��4mZ�����AZ��d�<!�����2嚾f\@�`!;���(��f}hÕ��'�b�'�2_��bЦ�P��:�o1|�����@ ��O���?YN>���?v�E?B��P��R�B�@1��m��U.���?���?Y-O���K�|��Q�����t"U�`�9@Ŧ5�'2�|"�'b��).�b چ�����B<V�hl��cJ!S���?	���?�,O�P�ժ�M���'���r�ߡIF�1k5"77̬ @�c�L��,���ON�D�&q�J�|�p�J�`�l��� ���d�#����d�O�}�hxUU?%�I�H��+��5��)�3Ve�i����oz��O<����?i�O�?��'��i��GN��҉�r�H�d�<E��S���b
��M[��?���"eS������㜔+@����H�:8�7-�Ox��G�S�
��/�d(�ip
�o��B^�"�.)��6M�d�oZΟ��	���������|�S���=a��j�d�.�f��)H�GR���s��'��	^��U�4�I�0Bn��#�[(|��#O��-��4�?	���?i@	��P�����' ��@**Z���Yj�,�b@���O���'R�	:b��x�����O��d�O�dPT!�,
�8�Je���f�w`�˦m�		l���L<�'�?AI>�6k��r�Y�Z}��*4N'c�֥`�Or-����Ob��?���?�-O�(����<&�H Q'Ńai�9���J-^�'�4���$�0��u��bANP�3@=7j<������M������?a*O����4��Ӡ+ot	���ͰXl��q�藕!�6��<i���',�7R|P7-K�_3<���k*6�28�"��6'�	���	ڟ4�'�,XHE�5��wp:(q���8r�w���?6��oZןt%�x�'N.���'��'X����lƄ$֨�fV ;K��o�����Zy�eH5t$d�b��k�%n<��oߢr6�d�4.�,�'��=����	F�V
s�������
 K|��������'EZ��C�t�H��OpR�O�H�=Ѿ�H1.�utԸ+sh��|���o���@���*lq����I�O��I�|n:� ��u�n{���B�3]�F� !�iM�Y���'n�'7��O��)�u���~ߜ˧��1yU�rANJ(D���)��E����y��iطGɚ�",+�ђdcоP[�<o�ޟL�����vJ�]yʟ��'�a2g��k��E �C�W_"�jGO"�I/ׂL�H|����?!��L沄(������\u�X7z���ire�kHhO���O����<!�@ލg�Ȩ����J8,IC���=���'�� ��'��'��'���7,Z�1p.�fc��)q�� ��a��ՠ�ē�?���?*O$�D�O���(L�'0�1�c�Hg$�s�L�D����9���O��Ĺ<�e�2)�)�2S���Yn�PAj�+̌\��������S��zy����҈�<s��|:���2o8$R�o�y���?����?)-O���B��G�S�?`�y���Z���!g�?u��t�۴�?�M>�,O��
���O��O�`�6ʑ.U�h�� �q�!ڴ�?���J�Q1�q'>)�	�?��{kr�
b(��X&Ol�H�0��<aW�¿�?YM~��OI.�w�X��h���1<%\��ش��dI�=�mZ�����O6��^~¤�NI�!�̔�MW<dق�́�M�+O�K$��OX�'>E%?7-�fr6�R�aٞPe�MhT�9P���?X�>6��O�D�O��G�i>=��i�97�����,�"Y|Љ�I��M��@��?9����<���PsO�;8K�u��g	���������M���?���&�|�)O�C�dԀH*p�Y�d��D������1����<�بm\��������2u�%u���BY.D��	|���d�r@ʓB���T�{��yb#5G_���Ť9;^��\��r�ϐY6b�x�IDy�'� xp�lķY�����Œu�^D2p�
�W��	џ ��]���?��'dnL"p��S��/���k�46�P$�'z��'5bU���������\��+�Q�R�t%���d�OJ��(�D�<1�C�?Q@�ӑ#��3��.'h%y�͋=��IП��ɟ�' ڬRC��~��#��`���B� ��6��K��E��iw�P�\��ȟ��I*s2��矄��>U'z�!�ޡ[�\�r�_��u�ܴ�?i���_;9����OR�'���J��_����f�Y&H><��3��A��ꓓ?���?�c�X�<y���?����4KE1n�J��H8D�6|!�����M�(O �äa��]�	Ɵ��	�?M �O�n�/P���w`ݢ`kd#2h[dq���'�b@��y�|"���&_f�M+C�ذEq��86(^;K]���.i֮7m�O����O���u}r\�2�nB�ڽ�$=�(��d���0�>����R�):�<1'B�,% �"�d�N U�i?B�'�/�� [L����O��	�-�rD3G��N�P<;�IP�$6�O�ʓl�:��S���'��ޟ�����ܢN��!�e"�>k��izR
U�$KJꓒ��O���?�1-
й���yѢ8 P�٫r�l��<�Át�����D��ҟ<��qyB�X��0u#S&�!`��&[�����>�(OF��<����?��t�$�1&љlx��Q*}0��P��<����?����?)����D�D �Y�'X����U�ͤ42H��3��\�n�]yR�'���ݟ��	�`c�>���M�J(��ʏa�2�ڑ��馵�	͟��	ПT�'Uh�
⋧~��6�de�כGzP��o�j�����i��Y�P�	֟��=	x��It�Ă�?1�xb�������h�q���'�Q��4��%��I�O��D����X�c�-8\�=X�@=  B�qELJ}r�'�'��q��'�bP���'O8)�D�RS��S֬+gb�lZGy�+�'f��6-�O*�$�O
��
S}Zwy CRI���,����Ȧ�ٴ�?Y�<� ��4�����}���[�C��D�6IКɐ6��˦�Z"mX�M���?y��ʖZ�4�'�j��c�.��Pj����m���i��P��3O��Ļ<�����'{!�oN�J�v`��!&&��ݱ��f�j���O6�$��w��$�x�	����ȼEG�iaw��U�����d�&�O�xI7O��ȟ��I؟\�LY+Q|�p�C3$�x�bK�/�MK����y���x��'RB�|Zc�(U֛z�P�� )&&�A�Od!�?OB˓�?����?-OD�Y���-3㠔�E0��ԥʺ�&����0%���� q`!�o�e�v��-Z��,��G�=GXR�	gy��'���'��ɦ~5�yh�O���Sfk��d 
cІ� ����O~���O��O|���O�M�O�)�g�}�XQ*kۀ6�4�u��g}��'��'�	)�b� H|��a��Z2���]�i���	�"[�f�'S�'�r�'��}�!�'@�H1�����4�Bc[=�| kme� ���Ojʓ���P��D�'��$��*wV��q�`�c<X`*��GEBOz���O`�Q5��O�O���+�n�1R��2�R���m 46�<a�KI����B�~
��z������ß���(b���
_)3�{Ӕ���O
@�0O��O��>��_8?�%��
�CY0�Ġ|�T�A�'�����	֟ ���?��N<i��u�b��raǺu'P��0�Qf�,|K��i�Ҧ���|�(O��D�7+V ɶ �K^�A�	��0)�\n�ğ��	��`"� E,�ē�?���~� }�T�i ��)pq2��̸�M+L>q�+^�p��O��'�H?� �� P�Sv��9��iǢe�ҹi�f2>Vb�<��C�i�����z�
 �0)�8�v����>1DOV��?	-O����O��<�T��;W��b���$��RV��$C)Ҹ�G�x��'�ў��%PuT����"�C�>`e�� D���H�Iߟ<����ty"�T�*��S�B��Y�P��J��҅m��u����?ъ�d�O�0��k�OZ��3�_ ajDx�)H�_�$�y���S}��'k2�'V�I�7�0�2�����_e�5�
�a�"`���Q�>em���L�'���'����yB�>ɗ'��x�XT�r�t���V٦��I矄�'�l�����~R���y��h4�����=��P�`B0.��"QV�����t�I#���	^��''�	�"-�ΰz_qV`p3��,6�*�n�VyEԴHab7��O����O��)�l}Zw�b< ��"S��l���E��
�4�?I�@Fx���֟>&kd̅���(C
�=���a��cO�7��O��d�OH��q}RV�)��?:@HS���& 1b����F�MK�I��<������?��؟H�C�"�*�k���oƞ!�E��0�M��?i�'�U�1V���'���O����l�' �@�X�L�d9�!��i9�IƟ,2� |��'�?���?��LQ�<K��+)C ,�q�*�3���'��1��>!)O8�d�<)��3�^�g�,�Sg�`i�=�4K�B}bK��y��'@��'���'��	%ez�Q���`�ذ�i�4<�&*��G�����<����O��d�O\���B�p���C��o�RMiQK�,p��$�O��d�O���O ʓ�-��;�R<��kI�t�J�R�>9e;�i������'��'���y��W�5� +�O
6y�؈�)��lʶ��?����?Y.O:�2��[��'�8�U�O3�$�Kw+~���Q�z�(�Ĺ<���?��SK���>YĪ��6�XU�@�y���;����E�I�ė'�JykU��~���?I��6��,B�Ծ.V�ʱ�C
]�(��\�0�	Ο����q�8�'���?1�"M3T�栁��ȦF�eB
wӦ�8*0bQ�i���'���OԌ�Ӻ�`Hɹ�,l;�/ԁ岥� ��-��ş�xw�{���IRy"��ެq̞,sF��-J=)��ܵD����S0en7��O�q���m}RX�`c�bA7p`\(�pCF�y5F��d�,�M+&��<A-O@��;�S��'��qMy�1LG�x��ȸ�Σ�M���?��'dnĹc\�x�'SB�OMh�ғX���Q��=���Q\�̖'&��O�	�O4��O���o�.l�p�Z�2y�f�\�R,^7��O�I E�f��������\��5I<% �b#� �E�k��I7��DqX1Od�D�O��D�<	qeǕ$����sh=�p�޻]��X�w�x��'��'���Ɵl�I#L��]�	ŶES�Ěr��8zxa�1�I��p�I��h�'r���a�}>5XU�{
D����/yD�+��>y���?������O���6����Z[J�[iԚs�\�B��xD��?���?!(O���a�NK�S��b�PVe9bȒ�Þ=�ʥyߴ�?������O���ޙr��>�R�
:p@V ��o��p�LJË�����GyR�'W( e�'*��'Mr�OD�1S5�+G��-(�ؤO�0��,���O �$Y�)�X$��T?m��n�.�)Ĥ��'.�#�cl��˓D�F8	'�i	��'�?���q�	�?P �Q�JK�Y@��!.˿2��7-�OP�$MG�b?92
�4~��E	�f�%C�x	 !�O����	\�|��O ; O �@ÆM[�%O2�yr)�2+�"���$R�iԼt�&x��^'L��L���G+3�.��8?5��bU��T�#jѶ`�v�SC�N%	%��nƟF˜���(	S��2�?.�N���M<�z@���K/X-C3l��Z��`i���G���r���:9�z���=n>�x��f)&��Ȣ3$G��R�'r�'�z���T���|����+,�J�V�Q徽+��V�T���S��7�q��V q���1��		�B�2̓�k�Ɋ�,�C�H��3͔�6�.�B���<9t	ɥ��UC/�{DRM'�H[/=dri)we�5\���H_��B�d�O$�=��!؃#��5X���K܈��`fh	��m����W#H*��Ezd�
�" ��<��U��'K�q�%kӌ���OVI��ի4�Q�S�1h��!�O~�D��`%$�D�O2���:xp�w��m�	:@G D�d�	(ywD���N~P��[�:E���X�8���2���UnB�G�0T�P`ڵ--�C��'(<B���?酷i���h��SO�,��)����;$������?E����[F�T��\	 �V`A���K�ў"~P�i�vت���ZG�xar�́*>��G�'副C�
� �O8�Ģ|2aO�8�?a$+��y?��%�Rq�!��P�?���Y2��X�Oi@�����~X*�z˧��`%�T�0'��q�� �O�邆�;��)��$>��"}"u�!.*�J�O�M� (��u��^�4�r�'��>���0�(4!�,�?=4���L_�4H�C�I5��Ջ^�]�@��3�G(o�.��ĂW�'\���+� `��P���&x���>	���?q
!~��t@��?q��?�;0v��p/�cي����SJq gC�=���@��'0d�p�gə����S�? ؼ���)4����`��^���h@K�T�х��x���y�q��'ǚ��D�s�"�BPeZ{(�E�W�'�	57��4���=	����Un�/d���#�G�!�E�U�T$(4m��� :�K%UI�	��HO�Py���={�����C6窭Z�nC Lf0�b�d%-�"�'�b�'���������|B�S�c�r��0j��*���W�%~�B�/�:��͢QK���<���1aP��u���	��ڸj�T�i�0]P#����<QՃ��[V��ԧH�*�vER�ˊJ��X�	���E{��D�y�`�z'F'N��`��@�jO!�&09ba�!�����3�d�471Oj��'��I�M�D���4�?��h��x f
�z�nM�VG�
��+���?i�
Ȥ�?�����$�G�tϛf�$T�B���7�ߢ?��r� *�p<E�9L� �Y�I�4����
cO�(h��B�%p��!�%~��x���?)��i�*7��OUpֳT��g�0]3�p� A
���۟��?E�4��F������;*-feI��7�x�aj�`a饌F�uJH �%��,�h��2O��p�`\r!D��?!����J�~,z�$øP�|�SN�#P��՚��+K(���O�,��� ��!�5%̣f"�裐hE���dY>Y�A�5	�F�
4F�*L@�Q�3�!}RL@)f�d۳aH�1X��t��l��>�'j�*2 B����U�W&e��2}ra�+�?)���?Y����O���4,�l AD�2{��Ĺ�\̓�?9
ϓ 0�%`W�ug�SG�Y#�A��I��HOf��UeL�_xt��&��f(O��D�O�����u�j�`���h�~����?�!�d�0&��84	�1�d�(I�V�!�d��1��1��I]�=�;GO�|�!��߶9��,l�B����	l�!�dH5O�0їOلy2 )��bE�p�!��o���b�J�e?~i�'�"�!��
z��0 ��
(Ă]k�a��t�!��B*0�東��	�5�M��ޡ(�!��7H1���h[�7����3�)=C!�dԼoPp�"p%��=�0�C煛<�!��߸^��ۧ��}�Z�"S�5Sc!�dF%S��["!T���
Ef�kP!�D�b����dN�:������F'<!�d�Lb���,�:}�J�C5!��"|�4�t��8i�2�ʷ��+!��5��y���)�~���!��m�!���v��y{�o�@#"�y�!��� f���.N�f L�k�,o!��Jz��e���04�����/�1W�!�6����!΍�P�����N�!��"�ft�Xh�z�m�*J�Xy*�"O���o�1,jU��B;/l-�"O����	�`|�E���!g�YHg"O*؉�@�zʀe�dG 7fx��"O*uu�TKf<��ĉT:��"O�E������*5o�?8�Ait"O<d� �Р�xa�N�&T�UK�"OR�
�7�'��"��=���ȓO7�YWN�_��Y�/�_Nq��C�R �tI�5`UPn;C�V���UqWϓ�5yj�a��=Qi����Dݲ�C#2��ٷ+� ax�ȓi��h񉅱!,(5�GNP�BO������1S&Ӻn��	�lC�a#rЄ�7@��P�ђc��J� �ޤ�ȓF �z1�f�	c�D]\ค�	�(������ր��^���ȓ&U<XxE�хQ�2�lS�[O��X�|��ԫJ=wn��ي&�����?86����5���0��_�@�m�ȓjr@��D� 	_x�V�lβ��a2��R@�$b��Q"i�mT�|��S�? �t�@�x��I��f�f�ة��"O����^�!(��Z��=a�"OTL�r,�-�H�Dm�"t�Z��w"O��u��:��ĸs�
�f�x2"O2�褨���9��˜�k��ͨe"O�ݸw�ШV���!ԫ�&�|m[�"O�,#��`����,9���"O %��e�"��M*C
ՀR$Np�G"O�1��
�ih�]HƂ81�	�"OV�[%�	%3>�-�֠��L�HS"O2�b��>�`�� Aԝ���B"O^P`So˪f����'��=V���"O;P	/�f=A�y>���"O\���X�,�V�4\��"O��
�ƕ?_n�P�6&��`��"O&�#I�em�ӁC�Boڡ���8�l��)��������#?1�RuV��!��VI��"	ftZ��'\�D*D�>0�>E�$L>h[���u']+2���Y���(�yR�V���� h<"�r`JO����|Lx�h
דj��!��|���� &�= �A��	pX�УnW<��h�H��K|nE����4-!�D�eƺe�B�ܢj���a@�p�Q�L�Z���'�����;JP�x���2Y[���$�I,1��ㄅ.�O�m�4쏮g�r�1��R��to���:&,��'���$&���,k� /ah�U��S�j�Ѷ"O�c���������K�X��^�t2�O��M��]�5��H?��cʁ[z�X�!����D���4�O�XsE��-C�5zC�	�����×<���(�$:}��+q���њ��{R*	AM�H�Bϗ!{��r-�
�0<)�E�j�	�VA (
1�N�$U�yR�����SEĪ��$	��'0QAJ�P������!H�\9��D+R�
�k��M���+��f��,tnz�BƏQ�c��Є#S@�<��˽uF��jN,5�LЗ+@y��^�=��`R�A^�ِw��x�OC�h�C��*�lQ�w� 2R�k�'�4�s���
UI�`��5��r��)s�� ��M#"��fD�c�nU*�1�6��	�'��M��ώ� q�1���5����?���GȜ�%Ϯ RE��!|&h2������8���s�	��9���J��}��=s�e� ��<��Mw#�X℈_�<o��s�cK~��r������0V����fT6�?��&�-"��ɫZ��K*��p�$܃{�L�x�Ol����K$8�@1bK�5kc�m����E�gh4c6���T�����SX�v�I��?Ac5��$�`�Ʌj�*E3 �`[�u;#O�%���JjY�R!N{�6s����YX�33��%	UbT��l�G�xX��S�jX�V)^%;6�O����J�(��Y��ͭtpް2u�'J D#�-�(0�n6�ל7���9��űIՄi(B�z��Q�E��(�G�'Q�L��.\�WZ����-`̍��zm�I�BeH==�����(�McF�m޸-릯��~��O�iP']� ���Ļm��ʣI*H��!�7N�=lB�#��T"���!�޼�D�Ҽ�8�E'Z%F�x9" ��O.�i%㱟0��!�?!�yעٵ�b 9sW��X��p=��OL�@�ċE�&WF�cND! e�!�f� 8�:Q;�e$}"�>f�Q���H�)��!�@�w?Y`A�3-Fʉ��#�@ેe�M��4d���A�d=�f��� �t�H!D>zYXdIדw����F$��}�v-�<�	�(�T�CF��/g@���*ߣ7j��>AƥNhN2�� ��U�
��U ����b,�L2�a[�A� �N�A­^?(�2�<�4���[w�0�dt����g`����8�q�'e�h��M+e9uj'���he�UF��2 ʔ�Pe�@#�rb�!�٫\i�m5A�/J�>���L����$�����	(9O^̐��ϥ�$�����DW�l�'2ړ�$��w��Ic` 35��[@��[�P(�竞�*)D�k$,�!F��L�<i�$��m� ��>>�Ȩ�JD�B�`��	P)�g�� �(���C��6m���æy���t�a��
Ɔ-"1{�(�c:����h @y��8^��q"kP/:�M�
��!����g��#����0�ř�l؇6�P�Y4���_�\!�II�iH����V>�5��Vy6�td�!DhԢ�G@#�@ b��'�@�X���'E<�i����~m`��B^7#�nDAfEذ�x�0>�
�+!M��P�e��m۶���@���D�	>��l�6�O� ��;���� �L2��ُa�bT �cƤm;Fݺ��'O~!�	^�&l�5�ƥ_�&��ED�vA�Ӯ�Q��y�F%
��t���6�����#\O P��d�9Zf�h􁔡w�x3���H��	o��bL$*���9C��O�Y�,�f'��'݊�x�L]�i(�0HA�<�dʝ�/���	b��a�v0�'#&�H��H�`fH0�4F��a�O���n?ͻU������8'fd:�^ h�2X�j@PH "��p	��r�@ߧP<4���d≞!xi#����H��qOPh�a�%u8dr�d�|Ҙ#p�'�J�Kg��1T�t�+V,X8-w*0/�괄�d�Z�"E��	�9�p����&F�P5
�I��Z+0� �N��t�Do(� C<��-O-�M�͜�W2�*����'�B�ɖ1�������>OX`�ƞ�a\�ɟʈq�}��I��p]��3�Bɠ\"��*�K�:
�!��4#�P�C$H�n?�Ȁ�U�i[�']~E�ۓk�JX�tQ�"�b��" ]�?�T���\�4��%d�����SZ8�ȓ2��l�5C]4%�����-�Q�|X�ȓS����WOJ�l�Xa"����7��ȓ�R��Ƃ�i�.t2�؋C z<�ȓw�rYct�E���)��K>G�p���pr�=�@DP�sd1Y���:Xԕ�ȓs�#2�ˡS�D�xᅔ6/�@��	]�QH��s��<��(SN{��������6��N��q�#wd��ȓ~��=���|D��&]�l�=���^��7��3 ^ցӱ���kvrA��WD��K �)?������Y����ȓ,D�eK�,�0�UA�"킼�ȓ�d Fd==(��¢ ���2�E��m�
��t�IV冼��77�Qk�@��D �� �4 BD�ȓ|�|:���<c{��kLk0^ �ȓ'f�$WL�u"͠��#oy�ȓ$@��J󬝊*��7鑤]�����*��bb��'��	��^�m�y�ȓk0�8E�C�<h�%X�EV8�`���f��	����e(�I^�s������\4���]�(�k��Ŝ!�X��%Zm���8� q���t6p��ȓK�ʠ�Z9:����7/�.jj5�ȓ7�Y�dǓ�?x<��DA�ІȓM�B��1�H�|�I�� ����MC�LidBɬY����t��9aD��ȓm|h�U�
~��Y+�ݹ[� ��s�p!����lk�Ặ�ŲI��e��|8�����S-ظ"��+PZ��E6( �Ƃ��>-��� �8�J}�ȓX^Qs!�*�\�a��ρ.�|�ȓ*t��	���Iy@E��r��ȓ+䘀l��]��9��Խ3�̠�ȓJ������R74$I���0����7�y#���m�6�	�wР���R6N(�R�W�r����-Z�^X&]��lC������D��@��OP�hF4��3Y��&�'H7�H3�����ȓ!��Y��<젷��*N!���k#�\��L2NE��͟{���ȓ
�z�B釓?\�hi�����a�ȓ(T���`B�|��Y&aC*
X�ȓw��q��-ϒV;P��@b��;𚕆ȓOG]��پ����gD�'!�����𐨧�O~�!x�h׎
���ȓa�E+��  <d	�E|��Մ�xȘ�갋9C݆e9d&�4,X�y��S�? �5Q�.O�ر3��AF궽H�"O�U���e$^9���=P�p�w"O���� �8y@�"T4��4a�"O�ap��-sF�zR�_?<Ă�"O�M��-D J���H�A��^�F�ʂ"O����&R��z�h0�J���"OM�P`@z"�(I5OU�b$�G"OB��V.�\�F����
�-�@"O�Ĺ��.+����n6_f���"O ��Ĭ�8_���U�fMx�kR"O|��A��}tb�@V�B�@�u+�"O�X'���н9��<t^��t"OrX���V�/~��� �ư]el���"OR3#H����e*SH䅰"O	 �FL#.��a���l�ТD"O6ǂ �	��| ƬP�"O(A��NY`@�i;_�P�{u"O|��I�p�HdP!V�H��"O@�����+��(A�"PRA@`�<I�)׻R����raפ{ | �p��\�<�����b���-R�*e|XQ��V�<�D
�I�81ٓ��)�@�2�
�{�<��(�'~|ز,T"<@"çGt�<����k�\MPӠ��T��
FY�<�F��X��=P��-y�x!��R�<9a��x� �2
A* p��R#�b�<�"���3�\��bݩkY$�3�Pj�<	W�D,h���{�jZ�=�`��φf�<!g(±C�vɣCeU$(Zd�WDh�<ɡ ��U����� ^�8PI!�g�<����9���Cb�DE�bY�6)�K�<Q�f�+R�z��fl�m�0@x��K�<�ć3D�.Õ�̝r*�X��/�]�<�cEJ�S��[���j���t�<��E7bfP�2��
M=���&�{�<�a��,+X4 w�z��4r�%m�<�W�B�x
Y�F�}G6d���X@�<� È@x��*��C�vְ�ҍWw�<��Z�q�"��x�mr���u�<Ƀ�ޒ2r�90"jȭ
����#I�W�<$���&���M�{(*�)T��T�<G�F(C\�`I�f�~�Li;��^F�<����.X1C�Uy5@ ��B�<�%��YG�	��
�(��T�áEz�<���Zt����#iU6�ġ]`�<��(��"����-^6�� -Y�<!��U�wB�!�9{(�k��`�<���N'U�I�(��2+l4�SC�<�@��-���y�
	h�0tf�~�<�b�4u hA���;NqL\��"`�<�IȮKN8��sa�[#�ث��-D����f	��8���g	|d��++D��2�m!h%=�5�ۃoth:��)D�<��7md)*��ÑP�j�I�N)D�,Җ@�6>��7a�S}.(��(D�Ԑ�S�i����T��9a���0e%D����L>�L�j�#� �ʕA��"D�l�ë�*z�H����V;|�fX�!?D���C4�2@u� /��p*N D���0en$i�e���	��J�*D����� ��b7�O�U](I�)�O���N44QB��$ p�$�F��(~m*B�	�W`�:�3|ʰhZG
��8�RB�ɹO,�hC��" ݔ|kf�Q�x�RB�)� DP��� �R� � _/wX�x�"O\���k�PZR�HS��&��XjF"O6�1���,kq���kn���"O.`Z ����+��ӛnf +�"O�Bɚ�Y:)P*7��$(7"O���� �dM��7q�%S"O�D��S�_]n��d�4�d A"Oh,�b��J&v���_u�Q�"Oz�Ae�p�kĎ;0GNh�"O�ݻ���"�R���i=�V"O��B���xh���F��#w �k�"O��8U�
L�ʉ�`\�s��)��"O�	��m8x���eW�R��"O�)�7䔾+����e�$nq:#e"O��mɕzg�X �WHn%��"O|�9���]H�c֥Etk�"Oy��2)bB�B�A	$rCL)��"OB�Ra�����"C�A�iB8(�A"O��I�ԁ(BW��,F9l�"O���$��mN*����G�΅�d"O~�G"��pIF=��L@(yfl���"O��8J]�}c.��t�â%W�D"O����i���(ѱG]=KK�DXu"Ol�A��ې
�^d���9.u3"O��UeĂl������ lH!"O�	�J2u�I��Z�%��y�"O>/�
K�)��&ԓ �,�"O�]��K�>�� �"k_�v8��0"O�lق�F�}�ۗ
�\`]�"O�(2C�
��m��۩i[8̳V"O,83Ae�+���ѦBPߪX7"O��$��9��QKuC6��}( "O���G"�%ULA�ł��*�Y�"O
)�p%�:b�B5"ą֬��"O\�Z���:�*�북��T3�pj�"O���g��!$7�	�%�7\0�yȡ"OX�y���x�樉vF��A-Vy�"O�h��yT+N@-z�Wy�!�d_`0��Db�o�lR� ��!�dʧ�\Q93��1i����@��G�!�$�.T�U *�Xc�nV�\w!��&pD���G�r��)8ጉ�g!�d]d?��W�8�!"B蒩 ���ȓ=#l5��皪y~ʕ���G�tP����1çfR�W�Bi�1n�+8l28�ȓR�p� Tf��A?0�˶�U3R�<чȓ
��L�W��8z��o	��t�ȓ^������g8pЭ�����ȓK��411������>M��ȓ'fP��ahM
T�:0��6�F��MS@L2O�<�V"�
�v9�b�Ph�<a-�j6��bn�]��凊O�<5+8��9B��!~7�1I%��d�<9�-����LQ�e�`N45���_�<q���'���Y��O�!��pR��`�'��?M�6��GJ�,٢B
�{3�Б� D��񧫍'P�p HSM�  �d�D��p����<Np�X��)M�~fLn���8���EN(w��6�͒E�ȓX��E���E��MA��A*	mJz	�'q�����k� �I�7|ژ��'8̝�P�6вY��c�=m.��k�'��@jt�C�u�
+�-�.nY$b�'���UaN5<��S�L Ĕ����� `�'��I)j�ye`ңP�����"O���eƵON<��f��<S�"O�hp!�ԀD&���Ϟ3����"O��ELNЕ(�6DyR�p"O� �@^.�`�!��+i\<��"O���/�[����$��6���"O��J������3.��v�@�P"O`y��'�,i��-��I�Y��"O�`:A.��_�ⅹ�k����=�"O��(s�7��m��/=���)�"O�̑2MH%RxP���]�#�0{�"OP4��L�g�FMK��=a���:�"O��(�jL�zp��d<IF ��"O������o��j�:J״u��"O�U"���b��;�b�m�J �3"ONu�ӢZ�BDkƣ�=}l�Ze"O���ܓj+��DH�s2H�"O
Y�R$݄�C�-�)s��)"O~���ĉ�eU���bl�i���V"O����烺#�1�� %�`�x�"O`E�#N�`=�L&�ۛ#��Ȼd"O���G�1��%���<�"%"O��`���2D4䁅�|��"b"O�:׊Oo��P;$�Оr���iC"O�I����E:4� f�/}|I�"O�PEI�\[�
����W"O��Ǉ8��<��B��.�}Q�"O(0��BܓW�P�xrg�R���"OƵ2gJ�L
���ЀA�� �"O��FM�z�:�F�V�6"O	��� ��|� ���44����W"O.Փ��+Oc�UP@$��.�����"O�Pp�B�H�Ќrb�O�_ctf"O؁�F�z!�T�fL��s��x��"Obu���zPZ���A�8a����e"O��o��ct8�0���?�ܘi�"O�415�I$�~�n>S����t"O���Ǫ��̠ g�{�ԩ�"Of�Sᔆ(�v�4,@�~��b3"O�����Ն4�P�YfO$_j�=;Щ�D�������+Xk����i,��A�I��yC��
�*�Bg�Rwx����ȅ�lu��ք�q�r�q��i��Y�ȓCa0��d9v�Y��Ƃ�Z���!fF!:"or+�u3dO�:��чȓ�	 b&έjh���H�h��ȓ�Cw���T����G�6]���'?ў�|bn?` ���J�HG�P4�NY�<iԉVq(Y�VÑ9� ��b��U�<���Ô}��R�2��x�/�S�<�q��/B�XhA@:Zb�kS��V�<�c���)@��k��u���hR�<���Ͼ������]�b�����#�G�<����,�Z�
e�χ5s�J�m�h�<��(C�N��Ա���Fy �z��I�<���C!� 劕�Y^t�p�nKA�<1�D/M��@��d�*���b��u�<�I��ODF\1�H߆�����F�r�<��JÔ[��P��x�l�4Ho�<A�b�,7`�y׃ �{Y6i+4˖j�<��Ĳj*��0�X�}�T+ �h�<� A,T��ȷ � #k�9��E	h�<����i���Ї�;(��8 �	g�<)p:\��i�1K�`���p�m�]�<� :A�h��8<���C@�q��LP�"O�%��e�2s`d�s��V��`���"Ob���dߞctFI�wF�!|�F	�"O�A��jO3eQ-�BK�x�8�B"Op A��:
�8D�  �,�S�"O$8�U��l�H��W7��Eɇ"Op�B�H_6,ڐ��WF&ŪP"O�Z���+ �h���8�0�"O���e�ц`����םCF�"Ox-���23�DM{��M2���"O�!Ss������u�PX��A0"O<9�E�Q�{��3e����0"OnM1�*��-��4��@ tp�"O��K�"�	>
8:�d+f��b�"O�uh��*�;0��0Ud,�"Ot��u �T\� 1&b�����"Ob)B��0 kz�q�K���	j�"O����:J��Q+�PVt)�"O�YBѯ^�2�����>jG�z�"O~d�&�9l
̴x LǤk4�	�"O�`b�P�^�Fɘ��D�B�
;o#!�D�#50L�E�E��yR�X
!�dZ��5��R���;� ^�{!����	�Ѡ�c�_}�*��>=�!�܇F 9#��YτY��i	�	�!�?
 n����6\!^�q�G�J�!��B>bL8!�� ��v��1�!�-5����d��-S�&�
��O�S�!�ė��]�mB�*�J��"N$<t!��_4
Y��U�ŵB ��P� �!򤛷)B�����*\��6Q0%�!�$\�>j��WFPbD|�b�'���!��#>z�!���'4ly{�L$Z�!򤜛2P�Q��+/��gϵ7	!�Ğ�)/��q�T�N�8���f���!�$�����J�!�'b�0�uH�;m!���:or\3��2���&��02�!�$O6�L��*�=+��E��f�!�;}�V(��`�ML�$S"��0!����bXh%��5R48t�T� 8!�䍹_p��*SF'���Ҭ1R!��4V�؍�M�=m����4��5:3!�]�^��iՃ:u�(BE�.?I!�D�0�Р���Xp2��s�@!�$C �=�!d�+%J +!霂E)!�d��#��0yR�%MI*�ôE��	!�D�X�^m����"�8R��(8�!��~���PjP(B(�g�!�dߨ	�\P����?�{Ĭ��i�!�D�\�X���i�\Yc+^�Dp!�AZ#� U.qߎ%�G+��FP!�D�)l��#J4ܦ�3�(M!�Xd[ziZ�e��rɌ���X-?=!�$]% P���cI��� j��-]%!���BI^ SӇͫv�Aœ~�!���)@Q�wױ��L@s�G^!�]D�&m�Sn�p�
�!%%�5A!�$mǮ19�H�,����7aY�R.!�ē2�Tx�ʓ�e���p��DG�!�D�>(�)8 �_�<����P\�!�Đ25B̙S��(s��y��I�S|!򤒂:ڂ��S�-TF���\�Ni!�ĉ�\���h���TOr�ˁ�<U{!򤇺!q�]��!��LL�X�&�*Z�!�� �"Fg�%/���0�b���,�p�"OJ$�Q!�n���P4�k��!�"O��J���9O��c1a@�j�A�D"O91���sI^��󯖮\p-
�"O �@���:N$$ٴdGxn�Cc"Oڌp�ό'd�|rg�:g���4"O>�XO�-�:�s�j�`1~�	2"OV	�7�ڇt�N]ȥ�!W$�Y�"OvTE�\�/0L�QSe�br��D"O`|�#�޷0�
��ccY�*�� y�"OT1Sb��%P]*t���Q}W�"�"O��B�ȕ#V� �������"OZ�H�"iʬ���3Iv���"OZj��M�-����`�]5p�("O$�5F;S~ܽ��&Wm��@bs"O��1����`r��re��!��Mp�"ORI���u�\4�s�� �P1��"OFh�&!߉6�PZ�/R�ݰ0"O
I�LU�B�!A@� ɲ�8!�DN'+��(юS�x"�y�`
�S!򤁧I&.�+��Ld涸9v��? !��%Tp2�k�� ٺ�xwe ^�!�Ā��zu+t"�- r�jG$�=Q�!�D�S�>T�@OH[x�3@ꊟD�!�$�r�@�3�8Y����(ʕ>l!�DT���H�mX+c�~9C2-��Y!��?V
��hdaJ<~��˵�I7P!�$��~F���A�V�3^���q��8?>!�d�{��E�D#T��I�b�!�ލ��QYg#޻*�&�3��+!�Ѯ7�D�z�H
� �zL;pGF!!
!��9�h�ɟ1�^��l��8�!�D�`(Àk�9d�,٠���!��ʒ$hT���ͧ3����u��m�!��N�Lu�q�F눂y���0��|q!���	m���KuA�fT(Æ�OjY!��ʕ?ϴu�&Z�&-������V�!�D���lL1�K}9����Z�!�D�.0%�Y+�g�+e��q�wn��Yy!��5�8=��B�Mɦ�	҇�,k!��)W̹����x���`&э~c!�d�*��kՀ�,>8��cFZ!�$O�8lJ�� M\��M�É�+{c!�DSO�J9AF�4Ր��r��6gG!��$z%�XP��$%�x\��Θa6!�dY����[�I i����E�$k4!���
M�.8�A�/"5*t�⎝�K�!��U�fA{ϡU�L8���T�+�!����bY�eFp��djs!��_�$�,e��^=O�H��cc�+B[!�$��A��� �cȗm̤���@��!�Dh�P!�fB$�e���Z�M!��H���`�u���2Ei��=e!�$A�5{��ʅ�Ȱ_	�i*6��aP!�D�,+,���FC_-9c�� r'!����d��Ek�%�t5���Si1!�$� ��}�#C�!߾�φ0!�P�1⤼äʞ��,���� c"!�URN�|���-�аM�7!�dF�3�$K�Ǿxn��4͏D!�$M�f�B�τ{kb8�f�X�!�D$]��$jBd�s0ɐ�-��C!��#U�@���h�d�CD̔�o�!�DG�yB��$nʝ�~�h�k�	�!�� "�J�G���Jv���|��L�'"O"���Y�a`6�f
WC��"Ol�·n�+ �:H����8�2�q`"O�hi�
��[f`�c�'Q	9�ri#e"O���F%�,n��U��Į;�nȳ�"Ox�%��*����!��v��q"O��W���T$
�V]eD��0"O�L�WB��4 ��)���"O(�@D숷ͼ����I�
��ur"OJ�ᰬ��L�\®�A�0ؐ"OH4���V@2x=�!�H$>��Y�"O�9`J�$����B+խs��aؑ"O0tc� �4 ʕ9!E��x�rS"O��P�$o�a@��7D�4Y"O�%�S��*'�~y��"M�R �"OT1ye��(L(�E�T�V��"O�tq$[2F��e��Wo��9�"O����=mT�2c��	Z4tЇ"ODe���&W튅�l]2<���2U"Oڔ�dGS�}�0M�Ş�Z���"O^B�#_�.>j,�g��1+�\Y�U"O�X"�G77�LS����]�Đ�A"Ob�qd)ɿJ���JF�-6���yR-$�l���� q&a;r*T�yb�5���s4�
�dt�|��G	�yҁX&�j��2�
���5:t��?�y���CTQ�e�m@
A�6�@��yB��k�I�/�k}�)��k
�y�E]�d{fEe�~�fc�+�y���-���e�aɸ�r�IW#�y��\fl��t�X�T����j��y�.�R/���P�=�j�R�H_��y�X5P��zr��6
�
]��y�
�S�)�E��%��;V���y","{I,\ѦcQB��)S���y��^HT(g������G�y"�LDa�@ a,���9�yb�EX��� ��1e��5���y2�X�"�x�(�&$��U���5�y��@�y6�
L�D��!�yB��#j)���O w��I�!��y�l�7���a突���Y����y�JL9L��\2�	�(H�B����y�i��g&���˨q�JԊ#�>�y���6�Ih ��*!�B��"F�"�y��Z�D_LYr�nѕw� ����y�\�{�xpX���$(��-B��y�/޾/�ơ����m�b�Ig
���yR�i�J  `H�b�J��	K+�yrP�US"�i�^\���w��y-ܪaY��� �)��,P�Z��y��ˤ4:�@�#.���2�ֲ��'J��?):�o���X �Ħf�j(@cJ'D��Д,�*���C��(YĎ�s��#D�H!�釯W>�ڵ�Е$�x���a#D����E\�4�0���B�Z��#�y�,�ak�셏~v@�J�T;�yRm1=߾蓤�nz�%j����yB� h��J�DS�m��q+�<�y�ň�RNFœt͏�3Q���DgY�y�o��.|C��
��L�)�%�ym_'�:Y�qӸ�8�)�� �y�f�
V���ڥ<�h�S��y�;p�`���E�5�xH0����y
� d$QƞP�j !!&̿E�ȉ�"O��S���O�bx[��C;	���p"O�q�R��oWj��ޜwP���|2�IN̓
��|��LD�'W�iP�eԤf섅ȓ�*Ly��8S���)�ͬ{XH�ȓ]��ᨔ� W���"�٨F�8@�ȓ
&z�y"*Շm�>�q%��� T����}�DJQnh��4��($�Ňȓ�༁"��ng���0�Če�f���/�2�IC�m���WƈD��	�'ў�|�e��'m�����m��}��d�Ḡf�<�č�� X� ���pl'��\�<9��	�N��A��$"�R@�CK�\�<)1O]�%Nv����$p�\|87l�U�<Y ��>B��9iB��K$�Ɖm�<1����h���
��)��_�<項X0#� Pr�6"�|����H�	j�S�O��=��cٵ_>>m�1�vY� �"OTQR�'��;���+2��YIn���"O<����=v�Z(!�Iƅ�!��	\�Re*Q�B�/��:)�@�!�dy�R��቞Z���Œh�O������m�z�A��bK�<�a&�#@=!򤄴��qr��
$f9���&��!��0yD�*�$1���!��P�FOj� ���0J"��⫝�F�!�$~3z��T2aPT��CK�%~!򄏤P ��7Iے$N�0j�KE�j�y�ት	����U��!Ԭ�SB�U�K��B�ɲ�R����ðq����FcU*k�zB�I90n�g䑭@CjM�e�T��^B䉁"?�������#x��b&��s��C�Ir�t�����?h���bZ++��C䉄}�i'B�$��!�S��B��&�jF��F��V+Сm�C�ɊX�N$�g��|X|�N�`�O�=�}�a
MO
�����ܘ|=|�i�e���ϓ!��!k�0rCVX`Ƙ���݄U�虥c2L�2�B��@���ȓ�|����Z23잁zw&I�f�����V812�ş�>���z0��2����U�|��&�U�V�tEBq&ݫ�Lц�&�ޙ0F�,.��d"1��'cBDP%���	z�S�'GdZ��40R����u�B#AԈ��yc�QkMX.m�ސbuB�`�詄ȓ�L*r�@1��(��	~U�H��- ���i�}lF�P��X�,��ȓLTm��)�,'p����[/g5r��ȓrn���E��I1��t�	���D��I<���f��Z|:� +<�V�&���	v�Sܧ 7�Qr�/4Vr��bN�.zB8��d�'9DQ�Y1� �kw�����YTC'D�|K��˜n/Ȭ���]�o����M%D� 8��(TŢ)���N23�؁��"D�D�S�&���[��N�K��2("D����n�g�H)�d�� �J�`�O=D�<��^w9�U�@  �.!я0D���n�$>A�m��펏G����+�����p�N\� �Db�n%�śq"O>�+Q��~hR�(S(����"O����"��@؄�tHG�y	N���"O�9#�⅃8��J�I"	�\M�"OH��h�>V>Ap��Ġ(��K�"O�A�s&3+�R��E��)B��"O� �,���S�Md,9#��A`�@�'J�����C����P�Cu㰝HD�?D��3��B
(Բ�ӗ� �'�����=D���Ċ"^�i�*[��L�f�<D���G'݊Y� �x)��a�F:D� K1�W,#��L9/\��R�6D�0�&��:fr�jU�e��Q�,4�O��C?���GKNg}< +u
>z JՖ'6ў�|�VK�t�H@e���&�+�#�q�<�!�H�	s,� ��u n��lk�<I�炒8�^E��GB�X�h���h�<3��f�-�%k�:w�x�PM�I�<#d^�=(�-!�A����@P�<�PA�">��i��	Z�9v�rx�P�'J�܊3(7 �
))��Lq$��	�'x��A���q& �V�ùN���'��ة�h�).V@�,.#<l�A�'}|����ڹ&͠m�5b���*���'K�%0�w&y:��4�ȓ)ބ�G&N�}���R��U�F܆ȓh)����ߦ\ �lG���K$�<�ȓy�lM��G��C���h�5�J-�'�a~r��9@h�e�R�'>��6�֘�y��H04�(gボa�@I� \�y�m��0���/L��i��y�+U{���W"�
G2��X�L��yBcB'ܬ	����34"�� ���y"dܽ0h1����/)�"�	�G=�y���"LyLmE@ͻm��D3�K��y"JQ'~��E�R�҅dD0���A�y2I��z�'���bu"����0�y���!=�B#�	]_(�#�^�y��X'.��MBW��h�������y���	��D9�'Ϩf��xER��y"C�R�D��7,��uz��pc����'az���U� Hx�+L�?u`�@���ybχ���k���G��]�.���6�S�O���-WyG�u tcѭm1���'v�@���J�@ �d�h�U��'N����R F�s ̏�=���y�'�bPJ3���C��0y��Q2�ةH�'(��R�k�*a�4��&�T,Y�����$0O�Y�!�ʓ �q�S�%�h���"OD�Iॊ�o�j|�5�Ơ!T��|��)��E6D11��52�e�vm��mr>C�2A���"� $F&M��d�B�	M��I'`�}�M�s*
�F�C�INX�qY���+_�Bɲ$��>y��B�IC� �i��o0�u�v�����+�d�O��?�'����7}��榋/ n�
����يBQ�a��愵e]v�K������'\ў�<�4�֡Kך�3�k&Z� ��k�<	�l�H��P��^���P���d�<YcDO'oC��H @C�:�= Di�`�<�ǨW�k��3�,�!/r�U!CK_�<Y�(K.ߢh����8@Y��Q^�<	��q�)�n@.k,̚&Ɂsh<��b�.sg�P�cLL?�lYA����?���?�L>1�����bC��V��@�T�q%�r�!���I���9�	�,Pu!���!�d?!d�!�.���5"���PU!�$�L�*})D����Y��$8!�$��q��u��������)��!��D�R)��[��P��8�נO�!�� ��BuC�&hֹ��I��pPҒ�'�!�$��:�PrFN� K�BQ�����0!��J�d#h�c�
�Vu<,�K�!�?S�LV��ZH��pcC�$w|��ȓr����+)��1:�D�
A���@�(�G���p�@5ie����܇�a��1:�ϝ-I:����̂'ˤ��ȓ_�*�m�-�`���=,A���	iy�|ʟqO��z���5A3+K70H0�`�}�<�e�/Z�əƊ� 2=�4�!e�t�<3���V�@�^& �)DIV�<	�AՏ\΢̨�H˗dD�Q�H�Y�<Q��E�^+n$����I�#J�q�<q3�I%(�K��n2�89QN�ph<F%��A��Bĕ24y������'7az¯�K��{K\9t�\�A�(=D�`@���;K�PXs��)9��8i8D�tQ%��E�^��'�9AeVI�SB5D��y�ޏ��1��=0ڱ�F�.D��C�a�5WӀE)��.]J`�P�(*D�� %H9K�ȓ�@� ����=D���q�� +>�%��-�(-pE�:D��zEK@�Z��Ԋ����9gTeb6�:D�89��*%��h���6��H��*D����L]�=�X��L�G��p� $(D��2Q%��v=�� ���) u��"v�&D�d��ĳWs�h�� �:= ԕz��$D��p�B�(R��C*�: ���: �!D�M@]vٻc�]	�܀ d!D�"�I	^���ICƟ2�T���"��?���	�N�!�5F�,7.� ��2~�!�D�I���rQÞ���<Ŝ=�!�d�	� q�e�C8;���;G㇈&y!�ǪQ����.�a���Bh�	!�d�+X�x|���O�ux�I"�� �W!��{��)xS��J����\�i�ȓL��ݰ�CJ�f��y�Ǡ�^�D���l>=@�G �E-Rو���M���� D��Pp�YS]��G�� j��|�j?D��e,��N�B����&�Nd�נ(D�̓TC_!"��y����R,����9D�|���sbh��m�V� �Z$o8D��(@�D�:�x�e�%��aH6D���v(�c*�=�tm�4�ݒ#��x�"<E��'���{��
�ٚ@ɝ�q�2"�'��Dc�k۶�'#��Y��l��'��	�Ũ!l����^�J6R���'�m��Ϥ
X>m�pK.APı�'�:Edaڔ)�δ,T佹����yR�ѓy
�Hf!J+^����w`E<�y��['����_:E�X1�5�?�K>����蟜�1g"�4"���"Ӧ�^d�w�0D�@�mX�/Ӽ�
')�(�l��׈.D�\�AB4:ON�
�`� Y2 +D��H��":�btس�ů�6q�g�4D�,d!�z�z�@��G�i�X����1D�l���L3K����d�"�*�3D��kbj�x���	��T?����2�Iş4��Ӝ$��	�Am�����K�h^$G
C�	 R(��[�Ȕ�B��BS�Z�L�C�	�h�*�tH�|���D`�"i�RB�	:?EI�-�GjԤӷ��E�B�	v3�HEi؊R
�arGAPFC䉹-���q�4z)�ⴭ��qW�C�)� ����G�
e�p9��D'������8�S��djV8!%`W�.�@���͇�/�!�Ď6ӠLk�̇�y�y
���,�!�^Y��Ȉ�7B�z��UG�=&!�@--J(�!A���Db��E=p�!�āXY��0�c��u�|[bݓ(�!��]�T�P�S� x̍�!�3>f!�D �����ĉT�d�ptJ񃉹@F!��6\	J��A׎e��ĐP#P�^�!�A�Cw���Ck<?�����BOD�!�$Wt��"�	ȸX����N
	�!�D�)XPt�f\�>����F)�Vr!��6u�<�Ӓ3�\�	��� :g!�/K5���n�<a�gû�!�ە694���d��Lc"< �d�?!�0[�4��r�R�P�~� C:G�!�DӐ*9�Q�0 �┰�=o�!��Y'hpt�@f��DP !�;'���d�<w�������=���`(��z=HC�I�0 D��a����MJ/��fC�	�@��r��><��q�R�0Y��C�I�R��K�M&$�`��.b��I�"O�-�A	Ћl�v�R�-Q !b(�d"O~�i"��A�H��΅L*@qI�"O�taC��s�̑s���:'� �S�'�R@˩,�i��� �~y�t ��!�DҨ^<��Rō&	̵!A)�0�!��yB)�k�&u��<1@f1P]!�$�a�d�c�GӰx�d(��]�9�!�DP������N,�ƍ3�,�4C�!���Bo&��Ǥ��s�T@#l�� !�ď�%2�(��Ϻ9�2�]����DH��4�f���)��9#�<�C䉆@�����-԰(<U�G-� n|C�ɯ
���Q̓�ĉ��LZ�6�zC䉜1E^�RÄ4��da�L�K�TC�	�:�|��D��J�����*�	9��B�I�E4R aڇNyv�� &�&k�C�!�,��f�]�J�txj$,6�(C�ɓ`�4IG���@���g���B�ɴ�v��&M#)f¬�C�^԰B�	���LA"(�)T�1�_)XӂB�	�q��e��$��p�ٞ���=�	�����ƣR��*)P7�D�4�m�ȓe0�2�DE�~����ȝ9NtU��Sm��7��/h�%�dK�6g:|,��dP���Տ]3%���1��S��\��E@Tu�8��;�ՉV����z����2fI#���(G�$4�����Ը8��,f��e�t�G;�J�Ɠ0䩵7��L�D�?MΕq�'��Xg����24B�0A:&��'��,����]x��	G�"����'Hx��Clc�b��*�\�3	�'�~X8�L�0z��1�R+&]J|��'�����N�P��4�բ:����'���a��Ѻe[@�G��/P�I���?!&�A $���̴f&&�bF��y��&�hh']
a�	r���y���-:���EM�R���������xrE�.(^�HQ�	ښx��ĉ�%G#b��Io���9F��!nv��G��T�t on�<���0�@$I��L
L���O�<���)�l�J�Z��"��՟�G{���1� H\鲅��>� �r�Ȣk���"O�����I&�$��c���Z�"Om��fV!&7�iA��J@rN�sO�xY�D�C�������
4?�j���O
B�	�#v&�E̓i/���DH���C�ɿ%���)�/jؘ]Q��T�v��C�� dj���ŢC�P�ybO��B�$m�6=�3`�!.v�@aV�irȄȓ6����S�zth�6<�9�ȓ�p`���ުDC�EP�%�1�5��Q�w	��&����1�![n#�P��AK��+ϐ
^���Ňу[uF��ȓh��)�GC�71�p+��݀r1�e��	z�'�d��a�_�*p�JR�}� ��'�D���p� ��l�rK�5	�'<t��ٗ��L��Ӆ6��L�'��=as`Z6#z�4�I&&����O氛2fA3*�f\ #�:���)�"O؀���`�p�#o�<9�"O��a$gͨ�ց�#V$=�@U�$�'���:�D@R�|Jt��%�([�4|O|b�,��IR	Wi~M�"���>h�� 4D�@��k�9�Q���]]�8�Q0k3D�D��E6�&�q  �C�6�+�o,�����Jd��I]>)
�� �$�Ի�"O�1��4 bu�� �|��H	"O�M[u�;�r�ه8�X=b"O��c̎&��3�
]>�r���"O����P#��v
�(-�D �"O�"e�x<ssdD!���I""Od���L)1d4�Ӏ�P�YQ.Y��I��@F�� �	'7<��aئm�6�Q3���y��
#/���أ�0zچ5@�I�yҦ�iM�8`�;t���AN]�y���N����C�%m��d1��Q7��'�az��,c�4m #W>X� �%�Ķ�yb`8f���KK}��(�UA���y!ؕ:eb�����u	&���y���X8��B��D&l����	�y�'�"O�h)����6G��IcC���yr%��/��}8V��%#80�ks�@�y���@�.��c����Q����D�O,��-LO ؑ�4K�B�I�ޛ*�PP"O�3 ���1 XA��!P(i
��p�"O,Pñn���A+q�T�@%�8�"Op�JՂU���b oM�1�Ĕ�"Ov���터z,,I�s/�6-�(H{e"ORB�KE)1^U����>P���"O|��#qn䑹���7�
��'"OR�@��Mж�P1��4F�H�a"O���"�PB;��Y�Y���"OF��M�f#@ ,�F��g"Oj5r�A�;.Ad/rQZ����'%!�d6`^��A_�wۨ	P3�@$+�!��'Fn��ĸt��"Q-�.S�!���\v���4�TA8��	�;!��(G��:G�|��LA��d�!���1��Uz�ë^|��8%���5!���+v�"�y��Y�w<����!��D;~���qB`B�S3qB�N��!��FR2|�F�G'ft%�Ҍ�9�!��RS�*qF�Xb*MDZ�!�C+�.8��`�. f�����!�d\8{KxHZ���
��I���s�!�� �1v㇞�x�ʴ�M�fH���"Ov��7�^\��<�h�8GJ�1kG"O=P,�/y�z$1�e^[������'����kC7^�T�&NȜ7�`����<щ���&������IRP�!v E�I��B䉭g՛���!0�;���m}�B�	*�����)O)~T�I�5NB��B�	�]�HP�Bf_yi����@���B�	k*BY�a��"I �%8R�"O�d�mթB��DaP��+i
�7O$M3�C�lp��BEZrX��2�$)�Sܧh�:E��q�8#l�zl�ȓ&浺㏘r��5HQ�ǝtzTtG{��O�h݃W��9B�	ڲ�ބbG�4j�'�P���U��J��2)Z�R`h�'�Ze��A̒|Y@�C��#	���'����?oV��"3Qb���'��E�r��yظ��u�ԑG T�K>����i:z��hZg��u��������_|!�đS�(�C�(#�t� ۿqU�IA��(�x�@��K�G�܄��jF�@���"O��$ڣ#�09*$�V$h�T�g"O�4��j�4,ČsaǱ-�>(9b"O��a앝s���*W	�m�mb�"Oxف�IȉT�u�@�Ї"v��RG"OPx5�[3(Vd�j&�W>J.p@"ORlB'���E"� q)?b:5��'��'�ɧ����R�eQCͨ$YB*G��P�.7D�4H���2�ʌ�Aߠo��`C��7D�P�W"%.H���=)~�!�L(D�l�`�!�$�!Th�)@p�� �:D������9$F��1)�	A��Xօ=��*�S�'P[BPz	_�u<N���f��LA9��~B��i���5:�^�SԈ�"hΔ��۟ ��y�)�=�x��'cASӤ��c�C.�Q	�'�0U�p��$��}@���%�J�'$֜��T�<�j"�B�.R�		�'@6� F�� ܐ�{�f�~uzA��'ڮTjEe�j��2v��{�]�'^���C.8���ɴ&�%��x��xR���_H-�c�ЙnP��T՘��d�O����O����O�[�Pa#�DM<MβU���!��P�0k��BF��)�� V�QP!���v%.�����/)78!�GX�pp��:A$���F�T�s�!�D�j�� QĆ	Ԣ�f>��{2�^��1 2�	�e&I��{��T�j,x��'[.�Hs� ��Oآ=��
ɻE&��<��dŁ�~��:�"OHh7(�*D��1���+���k"O��)F"Y�N^m�R'X� c�"O��bᙼ)�X5��?]�H��"OBA�rIIHu 1��n��&;D��ћ|��'�az򃒝(и���D_��� ����<����'jxr1 �Z⭚d�>�	�b�'�a�t����ЬݽE��A�W!�y�휆<�6�[���;6@��K�M�=�y���g�F`��>x*�m��c��y��@�R v��R���ZLdPe�+�y⯄2E뒅�GcR�U���B���$/��$O�1q��++d�ܚC��x��p1��'"�󐤋=(8E�
��=	��>�	�|��M�O!��j���K.`+�͑h v��
�'�R�(��<�vqz0AƺM�:dr��� l!�a�<a��4re�E�t�y�"OP��Q��:ʤ2F�����ӳ"O�!�U#T�2h�8�$N��>\���"OHxQG��\.����B� ���J��'m1O�k��	$C��qɶ"�lY��"O���R(�N��%*� �{l��"Oh�)��Ūq*$����>V{)�3"OX=C�����S���yc�� ""O�M{Bǚmz�dc	�Ue*%"O���C���H�8<���I-_'�)W"O�ًW��t��3b��(�i��X�����k��hȤə�b� u4I��'�@)!���6��ݙt� ���'� eKC�V&ǖ���΋�}���
���d�2#[z����M�L��5Y#++D� hG�>jV,b���0�� K��'D�8+��[�w/t�z$AIj: �	%�	X�'j�I�m��[��I�g��(&�
�>B�I*n��[��P8 *�y�JBE��C�	3"��$g��-st�B<i�C�	$K~<���ƌ.崕pE�މd�C��<@R飠�2	@�	�cH��>�dC䉢(2�F��7k�ӳ��}�jC� 	�J��@�Q"�
@ U�2U����d�O��mS�T�f��C��ag޻"v�C䉉6��J����o�a�!��ӒB��, &�rc�� '�]����2	0@B�w�DqA*������2"$B��	�(Q�v!�@�¼���P;��C�	7�>e���_+��Z�%����C�9pB�[���/���A$��"���d�O��$�&�N�r�ǜjFB��r,��f2��D$��S�m�<�Ȍ9��\��  :D�<Pe�1,�b��N��h��C8D�
/�>U*СZ�`G6��'5D��`QK��"M:D!Ǩ^�FҰ� 3�4D�����9�$\�����?��m�'�0D�( ��P!�F�acA����j�b-4�2Dn�R���N���<#���ן<���4+68��Z.6��+�*��z�p�����)X�~U&)ɋJ�P ��<D��P�l����p�G	x�L�!/D�0�7������JY�`UM@C�?D� rQlx'���"���x��)D��*e�M>�R@qD(U+9@�;A'�<����/u�vT���y��d
��ݠ��ȓ!�\���lB�c�H�`���)���IaTU�,ۘr�6	�2�$;����d^��/Q<~�f)r5C(��ȓl��t�EG 'pxy:�BͲj����ȓWdi���,����Ĕ9Q�݆ȓh���P#_d:�aen�7DyF��'^ў�Dx"D9-�B�H�J�
�1R֧Y2�yB�.�0YqB@T�v#M�yM��*�P%C0�C�8l,�QC �,�y�������0�����-�y�Q2�����)�hx!��4�y���7FU|YHu���*$ I�7I��y2# )�ܩj��6dw��8�?	���?J>���$9��XB`ϒ�0���Y	�'�x��Ō9v� Pq�M|�l��	�'l���Ҏ�]�Ɲ�EY�pk��'�n0��g��+i��ar�Bb�pв�'��	��`�%Ad�9j���S\H�@��� ��;��[�<��Y�O]96��4pW"O"5�r�M�[X��nC&m_�` �"Od詠R�+�x\P$�=vl�ը�"On�TD@��FC�*;^`�d"O�ұ
�8���h�,^����"O���`��u�u&�N �Au"OQ���$��ô
Q�J.�y�
��:�����!Gf"���
��yBJ�HM�%���j����V����y��	q����b̓e��œ5��yRK��]�yz1*�p�r��H�7�y�Nޢ.��-c��Y5mp���D+�y� �;��q���Ӧ8m���� \��y���Nah�;@dK�|,e��i͈�y�`�/T��؄K,��y$l��y�F��S� �Cd���
B�Ac�M�yR��E��@	cX�1[�	�C̈́�yro̔�2<��n�%r�(��Q��y"l�0w���`.,n�������y2鏦H�6U[Vi=a4���KS��yb�9�T�إ�X]�A�����y�"S� `��;��G���-5Z܅ȓ=\�X
��L�m<Z��Ú+�贅��L0EN��	��c>5J^|��Bs���L4������2iLq�ȓCo��C/�e^!3Ш�F"�ȓ`�"u�Gk�)<&^M+���H��<�`�acF�.hk�;�� �Tj�P�ȓ9葐�  nK�@X��C<����IJ�`>����JĶMsV5P�,֜KɌ<�?�ӓ�b��G��7�q�eM�3���� ���i�K!��24�X�����N��q�х�� \�p�n��9�X���,(��S?f;�أ�&b�x��f��H�3NB�}�:p��fU�x�Xu�ȓM�~���W�r�r}���S!GʼX����${�QW(�Q�Kl�><��P���O�0O�ejUL��$Ėa��g̾)a<8��"O$ �Ҍ:�*�7��#uT�Q�"Oph�E(Z�W�4Lc��6+7� �"O*�@�h��� �&J>�B�"O��a2���+fb} �G�B<��"O��P/�}LrHA��m�]��"O�B�ݞ�0�Ā�*H�lm���'r��'x�dI�vD�A�iɿ}�|�����'�a| ��08$GBA�4�H�vaɡ�y����$-J8@�M@�5h� ՠ(�y�ڳr�h(��"������y��W��}H̓2V�)�iÅ�y�H �pt�**TtJa�W*�y�A�vn�A�C��P������y���:�$�C���I�$��y���h�|*�gO$&�U�dn�#�y�n�	A�pP1fK�� �l\�yB��
q;:zq�$
����FL��y�M���(+e�T({���Z6�D��y4�.�3W/U�y���[6�ߕ�yr���u�eb�Sl~�hxEN�.�y�i��QD��S��*`L(�z��y�KT���c"@ X����j݀�y�Ҏ}��M�sDHKPN�r ���yB��.��@k$"�/��b�թ�y�E16A�2�X�V�&���8�y�n �%t&4 �hY-M���E�B-�y
� ��#� �%�n��c��pŐ�y�"O���2i��C��kdH;5^d�qA"OZ�����2'�=���OEQ����"OP���獧t�PpA�&ǰH�ak�"OV�qĂ�-���x��
�p��B "O2tX��N�%@��3�M51n� 3�"O Ee�FHx����̀y�@4*�"Ov�� �Y�|�*J�#Y�k�ք��"O��CP�
1��<��L]�]��� B"O�5`��;b�&d��
����IR"OL��V�ٸj���S�2O.�A�"OB����:J.@�����2:.|j�"Ot��R�ƒ�J�SLc�a"O3p��g�I�3���(�
5"O"�X��SR���A�U�|��e�B"O���C�Jă��	3V����"O�m�6��|u�7A�&�a"O�q��:	�D����l p2"OB9��,^�Y�t(��/�i� �F"O��Bv`^�X6(���E�d�"O|�4���MlJ�[e�^� �P�"O�rI,6��u�#�`�ш�"O����L�J����`�R�|YV��"O�Lr�Ɗ�?�}��@�Y2
)�1"O�� ��p ��D	/>#v��"O<�{�@ �	��R��Ű	
<��R"Ov��ʃ#�Ι62����`"O��:Q�G� �L�f,0z�U�U"O8Hj�'�/z"�Jk�xy�T�3"O:5��R4�lzD8f1��"O��p�3r�H\��A@�eM��!"O�8��JS����	W*�'�&�2 "O���	��S�(j֩��\��]�"O��[7�	Q�1gnH'p꾔�"O�)�Њ֮�{��C�@ڶ,��"Ob@f�Ȅ@nҜ���!<�-�5"O��:����U��$aRU"O�@���6��ekփ�����jB"O����#˷	,��	����P�b���"O���&l�ߺy�eC5}4ZX�%"O�,
ã��#ⴱ�����<�Y��"Ob��/��b�0��#W��d-�s"O]2F��![��	�e��o�cE"Od�� K�=
�d���K��Vp��"O�MB�ɖje���ͺT���X@"Op��-B�y���ƤI^�u8c"O���5��to,��A�T�8Ke+�"O�]�S� Qt����#�����C"OJ`@�g%��DzA� ���i7"O�TɃ+H%��۷�f�l	��"O�h��L�q)ċگ����B"O�����ѢZ�P,�fMM�8��L(W"O��!�w��h���P�d�L�"O��C��ڴpQ"# �;�($�"O2� �B;hd�DHB����"O��ҐG	���ƣ
1	5d�PA"O@0DK}�ՉrcR;���
a"Ot�هb�o��Ac4���9"O&���Z	V����1☛	����a"O
�X@�s�8�W'�	�r}2�"O�Đ��T PQ�M�p��Tn<qs"O|R2�J�@3���oKtY���P"O���MȩU�҄��\����0"OJ�	q G`�b9�������3"O� TX�pg��I$<spl�5|�(Pxw"O(���T6a��Y�@��� ��c%"O*\�%j>,Hy�Q�K(�����"OH�s��ȐQ�i fI�$��`d"OD��ҨǳfP�H5d�5K�� �"O
�a�Q�����;x����"OF,XQ�&@J�`��_�WPb��&"OFkU,$,�}zd��,1�Ա"O~�@�&�$Q�R�!r�ڽ@!P�30"Oȹ��I�;F�aSCC�.��"O �!5T2qe�p@��l�R�`�"O�����E�j��- 0���H�9"O@��+1����a��)�(p"O�!�F
������֫P3�"O�P
�B�nUDA��`��/(�*�"O:�r��̧l��*�,߱)7��U"O��1w��2<ܘ�CԦB�t���"O.i�#E�[���8��Ȭ{��ak�"O����A��H��0�������1"O:)"�.��1ka\�|�șQ"O~drr	�6�*�a6�	xL*��"O�@"u�;>
�M��]9#V)�f"O(qwJGC�(��-���
a"O$ ��+�-� %V�O�T��"O\h�O,])�ҤӘ�%{ "O`a��46
0X�%��0�����"OF��D$���P#ĺ �JpBP"O�Qu��15M�9VG�6�4%:�"O|�3l�8`tP�#���	|��H؇"O�ia��ڥl�PY�^4���"O�\� ��e������kϐQ"O�t���*u�d�T#!f�q�"O����O�0�0z�!�z����"Ov5�vϭ0��aq��&E��4q�"O\��Q�  N�Q��P#E��P�C"O�*���TX�iïP��Ũ�"Oze2$��;#��run�~�p�7"O������*�;'��bf�h;@"O �r1C�,y���X!�֘c6e��*O�Myvj�n4�zb�ǧ#ޜ��'X�"Si�5�V�;C���M
�'6�ؑR'цh�Er�	XN���
�'~l��%L��jMT��1�P>L�V�9�'��i5�V�L/�@���@�~1��'-*XCP"(Rl��" ��@���'T�P7�
�uD��R���93��a��'��Q��B�q~��dǏ�2��@��'K�h�sϐ�%i�)j�U�,���"�'�� �,țT�H�iTKR�5 ���' ��Ĩ�6f|r �6
"a��<��'��(�Ѡ�T���za/]N��� 
�'#�k�iL*2�@��hH	BU^��'��zvk#~�z��"�ɚ,�A��fź0����vJ��+�=&�N���e�.D�

*y�ѣ:BV&�ȓM�NT�����Z�
8We��ȓb}h�C��!(�>mj���[� m��Xt�E@��/A8��,�3	V5�ȓD�r=�
��(�p�Ï�W�h��ݸM�/�1���E�L�KM֍�ȓ4i��@�7/!�q[g��)(�:���D�`�I�
�fM�(�j<~Jz5�ȓLYԩ3dʣ^��!�)B�+.хȓ#g����;���R�X3p�Zy��S�? Q��u'Ԁ@r�Q�8�\E�q"O� `F��
{}"]:�ژ�����"O m��,��d��� ��+B�k�"OT��n�' �Uڢ�7D�)C"O����]9-@��N\�C%�"OpȫCo�/?�i��_�7��"O�ma����F���q���)수�"O,U	6$F!8In�:��֟UuBȕ"O���6�Y44�\0��7(mĥ	W"OH!��_s�:a�@5lk�ݢ�"OJ����>j��+ں>{�l�$"O����'�tDPU���(�З"O��is��7
n�|"�עu�t��q"Oڰ6a�1o�QP��ϵ<���S$[��D{��IU|�*i���n���J1��$c����W�#�pa:���?<t��	�y���c��ÇC�3I���ծ�y�1.\ع��;i��H�cm�:x��C�I	.�| ���V��
������d)���-q.��f/D�9��ِ��sFB�I2ly@�nH�p�bQ��Zc�B�84.�����Y73�rd��W%~�B�	�4��G�4V ZX2�o��:C�%��7(�	:o>�@e�$��C�ɮ@��`HR79� ���U42�HB�q[��Cp�Em&�9��X��B�I.h��Q s�������B�I"\, (�h4�=01�F�h��B�I�r�i����`�t ��e�V`|6M)�0!K9v$����C��5-��$�%D�D�F��>"v�@#�F��	���>D��A9g�z抁
2׮�(�B*D�s�S7"D~���@y�����&D�8�OE�R����
lq3�$D��2���"�В&֋I�<�!�<�G��>a�(M5�0�۵Ԧ3���@��4D��(�-�LZ�uEL�O�2���o�<��g?�S�Om�Ě�� �0i�ի�HݐP���y2��K��{�('$Od��S�
��O �=�Oj$����[��5b֦�(� R���/��>�k1� #������0�Jb���c�����D�#�t�XÉ8]����Va�'9���˦�Fx��)��`�V���΅-�L(h��ș`�!�ā�H�bШE�ك'���jqň��V��'��gܓZ���K&�]84�E�a%��^8��	�<���B�:���������0��Ay�>i��hO�T`ShXh��Z� a򤨡�A��O��@p�j�OZ�8!��'#���7G8T&��'�L8��N�M�6�T�W�E �'N������qO�a���� �@�ʻL&��"O�,ʥ�X�du��y$����0��x"�iPa{r�]� F��(��~.墠aο�y���r���;�`�3JPH�����>��Op#~B�b�7[�~ȉv�!$���(���V��hO��ŦAE��hʲ�b!O���#�<Ʌ�)�'m�Jtk�&��v88����'*��ȓI��-�s*x{�>X�7���6$�&�$��(/���a�F�x��&��)2C�I��|�0A1^zQ@�ی'G�C�I�!�r�#���ڠ�a�֥}��B�G���*�چ�fQ���g��C��,)�)D�;�<=�W�[8�C�	gBu�$.  6�01X �ܪ!�h��p?�fㅫ��3�KȚ��D;fJ�eX�`�O� LՊ����ɁD��3�h�"O|HQ�O�SF�� MT�G�m+�"O�`��q��i5A������T�HFxb�5~yL�ڠ�W�� h��J=�2Q�ȓ1~�T9RbѲ`�0����g ���ȓl��z`��)�Б�k�-OG��	p�'�"<I�4��(���$�A8��_�r�i�ȓ	1�����+6�B�s���D�'ў"|Z��"qT��g� ��a�#��E�<AV�ǖ+?�Ѵ&M�F��P�dA���xB��b�*� /�,��swρ�hO���I���h���ψ%Kz)����'ݰB㉋i��[E�	��ѡ��ѣo����hOv�<q�+ Y64�Q�cS=2F��Q�a�TX���O4�{�A��d@���V�C��@VS�HmZd8����}�vZ�e����rk&D�8�WA��X�ٓ�-�>:�]n#D��	�.(�2�h⃕Q4��ƫ.�O��5�CBI�^� �Xa, ��m�f�	Z������=����/�haH�(�O��'n�S�3����2ڬ���A1��%^!��МQ�N�B4TF*�B`Í�+S!�DD?؂H9�bT�� HX+m!��]�3eHA7�I�cD`,�%$ہUN!�D Nx;"c�)?��s��E�HC!�$��
2��
s%��o��(2g����!�$��8[��P��w��xp! �C�!�Ă.>2Ŋ�2JX"�j@e!�Ę�I����+�
QJՙw��1da|r�|���`�XRe�� �{��6�y�!��'��T�3�դDn:@��&Z��O"�=�O1<����#TuZt1mM�c�����'�D��0*�f+RY���]���
�'�RTj��R�"�H2Fw����'lA���<s���� �n#���'$��I6��U����a�!^/��J�'<t������h�@G�Qp���'��d��1����#�	�$�/O���N��P\���Q��u���� 	��}�4�pg�5 ��1�/�/:��B��<D��ᣔ8B��ȥhN���9D�8�/ղ	��}ؖ-W4��y��&9�lZ�#}p4�f%��{p��%/ݳR�8C�	?=y��aM�f?<�� A�'Fv���/ғC
1ԭ��J�`q�L�?xv͆ȓ�n] Ԭ�,A�Hl���V�x�'���2�)ҧlmfa��C5N��M��*�X܆ȓb�7�
�[�!�H�0�vYiN<��v=Z�C9H4��qF�rL�=�ȓ� ���F���ܐ�f�A9H|�H����
�V"/Н2q�U�͇�	{�'ϴ�07`�^�!d���dĀ�'�L�R�_ZF:�i�����N��'��C�ER�T9�!,�u�t��',0@�����B���`!�R���y"�)�H4f��$eJW%�t�z�&�� z�'��uY��*�,��ˠeY�D��'���s#�T7b[��A4'��K	8y�	�'n����`�bC���B�<a	�'/��0L��|�{���,=�$�(�'�I���׼V����I�<��$��'t�# LS> ��(i�$@��� �'E��hO�O;���� � \�AP�5��3	㓴����B��8\� Q�r����S�? fX�C!G8^��yhVA��s�"O&���Y(؆�kaȵ"2�a;V"On�@�
�9�xЛ��1#,z#�"OXl����)mJ,zC�1�]�g"O(��桗j�� ITA#m��S�"O�i�,L�H=�' ����qT*O�`s
"%�P�B�n
�(9�'��Ik�)�<Y�\P|`�ʊ9(ҊmC�H�q�<���4L\��aS�[�ut蠴�i
�'{ܼpl��<'�S��ެ\�t�ӟ'�ў擜ٸ'�fd�'E�GLάa%'��.��L��"O�ɫ�C�4m�Q�F�#�9[54O�<)�����"�/j�,��㏏Ad����"O��맫�26Y����6U�K�"O~L����5[6�Z��
n(�� "Oz9B�"0�qI���9_��`d�-|On���шfmЈXj�eL���"O�m���ʩy�8(*1薡��q�A"O��G��l��K���0��l�"O���� �b���E�X|hD"O�@`��ɍ��9�P�K�b��"O��h���4+�A�Z�P&z$$"O��I�	� ��08B�ڠ"O�eR�K"ª���R3m��"O$a�ѭ�2l^��Bhp �"O���1a ,vǼ�5��5�4��`"O0۠�B�� w��7{Mj�"O(�1�N\,�� Jw��6	U���"O�PZ�Qxd�=�C��(��C"O���!N�<ޥ8�"�m�W"O�|;E�L�M�|�I���K��¤"O���nX�j��xpgiΌ*�V|�"O�TXF��3XNb���K=��Ӄ"OJ<� �� H�A�v�ϝy� �#6"O���mP�*)
����і8�"O�5��J��u:���:kĔ�K@"O�-�p#X�M�p]3�EE�'���K"OX�S�l�?�9�#���?`��"O|�Ɖ��A�6�?B	$]j�"O����.[�����=D&�<�P"O�t��K��xE�5�����"O�]y)��J`��x�����"O�@� �I������/�8d!C"Ol�1)D*07d!�1E���a�"O�(A돱R'�<{�����!�Q"O�ͪ��P�&���I6� ��D"OJ�peʃz1Z|��I��O��1�"O���p�<"���a	ޒD�A�`"O�9X1��=c.�}�a�	5lQ��c2"OPP�^�Hzè��d�k�ᔃB����1a#0���0�'�*`˳�C�}#p1B�G�	�!2�'�Zu��/mwDHkTjN�x͠I��'˜`ǡ7�Bmԫ�}�`݋�'���`��V�"�$u��K�8M�D��'mZ` �D�.�f ��&�><���'�����ȋL���9��!bo���'{ �x-�H�,��pH>nD0L8�'�N�W̉�j�b���gY=[���'�􉡀F`:�(�&�]z ���';b��T��F�P �pn���'eZ5ϖP�����-[�o�� �	�'/�L�7��Hhh}a�A�o�� 	�'v��em�;@`����]3f��e��'�I#A���*��q�� f�T2��� �г�+�17��A������"O��iЌ�~��f˅�j(a0�"O�]@b�Z��$�!)�>�%�f"O�����1�N�SΞ�$���B"O�|+��I�]���7"�^˼�!2"O|1��b�3c��\����\��"O���eW�
j�+'�ܕ`�8��"O���-�#���9��=��tZ"O�X�cĞ	R�w�N���9'"O$ �ꃍ^��@O�9L��Q�"O���Gj��E�N@ӲO��a"x�ӣ"O���R�B�i��O	� ��s�"O�ՠ����g�����*J6��"O�T�"
�*s�]���#��1[�"O�����R�48�Т�i\�;��j`"O�9:R.�@?�
�ݍHV�E"OЌ�L�}"@0��l�x���"O��c�.�n�4{�,��R0d"O�9�N
H��ҡI�B��h"Or-�W���*jꔂ��<PM��"OH@8�J��<�2��`��)4�� "O�䠳DիQ��-(#�6z/R���"Oh��.t��wM���0��"Oj)
�e�7e_`��E�1�ܥ��"O��S5爃ij�<ۆ�&(�n(��"O:�0�/ؚ9����,�54�ݹC"O(|r���)+�T�s��V�/y��R�B�V�������,�����C��u�Z-z��4Z(�􄔻R�)�N�T��NL�T��x!�4olB�0��"D��B�!�Oe,M�G�ǀQS
�r�>�	 RY�J5��D���Z���.!�@� ��S�!��pw�@���$Ͱe�R���JH��*�{�������ɶŰ� �̏)4�H�H�_�eTLB�I0AEL�;v���L�`dJ&Z�a��	+��=`$�~/R31)��jS���-RU�Ü�0=i�I|��'���S+T(i��107 ��p��'_f��([~�q&S6m;�p�{�I�7g]�O�Oj��9�MW=F�̢0 
�fB�TR�'g�LcM�2:-� ��Ver��'�4c0��,���',��@z�$�'D�M1��k�B�� Cdz��
�'nt){���!w<�h[�"^���'�����CFB����%��0��'���@֩�"���i`I�L��q�'��a��nQ_ۖڒ�� tp� ��'�d�㦙\%xUё)�
?V"���?W ��f�m�H��nQ��08�6�Z�h
Y;�"O�Hp�	R)l�\�3���/�(Oȩ�F'BO�Ni+���\7H����7@�\��u-�QP!�������[l��a�,��!R��!+�s���H\v?����OL�k���j��@
���`���"O(Ex�I�("Xq!�&V�l�װi.6�{Q�D�)+���
ޖ,��xR��)��0�"��8\C� ��ē_p:� �(!��*�9r`g�	$X94�iI�㍔	C���A-L�b�����Zx��pC��W�K��+S.��V#�\8"o;�	�\&�Ǎ0J��h2�q~�&>IA6��oB�B��:f&I+�!8D�L�/D�
:�S�-�H��w��5b�R�� �8A�ެ0$Q�x�ң|��O�l˵���v�&(p�ōbu���"O����Cy+Fx3 � mkX���?9m�'"E�YT-�ƦQ"���G~��Z��[�,

�F�*G,��0=Y&A�G+X�{��=/��Zq�Q,R2��
���"t+�
� ���'~�1R�8�@iP7�ϕ(�J$Ç�"�X�!~�PI�b9Ӕ,�dB�	U�:�3�ן��ݲ_d���d��1�u�)	��C�	�����Ғiɀ9�$��мy�@�8�&Y28E�P(��m�����;IO�!�'��� xI!pˀm��)�X'�0i�'�}�t��,I^͓AN��DՆx_&��V�� zj"�$�?bI@A�'�S�m<-��� ��O��@u�ԇ~'�)�/Z"?q����d��;R������y�H |����~�x�z����	[����q�p�D$�sG±P@�'HԼ�d�8X8H�Q��X�D4e�#��8@(���'��b�8B�D��[>B�A��ؠF0qțw���FF֮F��T�I��]e����M�p�:�E��hk� [4S��ij�#Q>S-��BNY�
�y+%�''0���[.$㒅A���5V��Y:���~�'��Xr��?�T��L�Pa�xY�j��-n�ѡ��"y���/�=���ْ�J�B	�T�?s���Ң�Ӽss.���eԠ���.��]R�]���$W����7m�6i��D�p�½�' V�6i붊�)L\ @m]	zr}��r���ӗ)K\0��܊|nI����o��E��F��v�r뒟SRn�ď���Px"��}`���R��Qc���r���G!$e��9U7!��$1w@�}X� �[P��yBIL��5V�_?��Ca��wކ�a`/H�	V�����<�5ɑ!�jȑ�HƝ(�>�!Pk��b$�F>�v́"��xi!k�(gܙ�*�4�p���'�00�qB�6N�^��SCؔ�. {�}E��Āؓ����n� ��`Q*���	<
 xt� >}\��X�Ƽg�.�z�+Ƶ:�����$Sh�k��2LO<̉�-L
���cFˀ�f�U"C#C��ڌ�,|��b �ءC�����B�5%~�'/��?D��rk��8��4��֤ ���j�� \+!��,��<y��Be�^��bEۿzl^ɒA�NPb*� 6�+-S����u��#��|���S�T_��  �I���>��G-گGz؆�>�YÅ Z@8���V�št��-- ���g%��Io�x�9O����ɪ|^���Ói�怠B	:,��E-�>"����?�g���r�	A��uZb�O��ب���	!O4X���]a�r0���[�bT�� ��E<1c�J���(�
;cR�k3��3�$���+�i�EIÖA!&��X,��1�B���3T슲b�A�B�Ɍ.~�0Ꚉs��c����k z�1t�;�)�'7p�L
$�Y�B�رB/��:�ȓh���bPo�<�* �����)�HC�IsPP �5yHtԐ����PC�I/ �K � x�ԗ]m.C䉕F����F%S0,��j�ү]8C�I	Z"�����߂$�,|���Q8y�B�	�'6�eX�/�c�8dQ'�-o��P(�év]���>� ��⧛T�<a�f�o�2�S����m�9ÊSm�<��n-L�� Dg��/�@�tk�d�<�x�<8��W�	� o`�<�Wh� �p$�Ɋ.���pUhb�<���#�L��a�Y���sQlW�<� ��1�]��LH�h��9�d��E�<�B%�yD���aBub��U|�<��DM(E#~��I�J�!rmI{�<���@��$��L!o���is�<�ʏ=~���
�L�0URb�i�<єd�oq8���Њ�52La�<� (O�J��q�O u�\���� b�<A����� �ۧ?T���v�������E�I-G���"�*��q33N�;:?�C�I�ʒ�z A�c�q�D��	+Bjc�x�4�)@qO1�ȼ�"�@0x���="�|� ��'T��Q'�w̓x�H`iC+��k9�9�Ǣg���I����YR��|�  I��t[1�� 4����5��D��mjŋ1 :��	��T���3J �3��K6%b��"O��.gH%��[0��#���dc�ԋ����y3��>Y��V(Zy���^}.�猌>0�~��'�*}�F
*��)��L����	��'["e��eB��<�`�%ĥ<?D\:h�O_2��qJ�
F[JD�SE�W�����OQ>;��Ď���
1�_'E_ʡ��(�><�;�E�}���i�Q`��|9J���ɐ�?��K�F��Ӡ>un�7�"��$X�VDԉ��.�<%o�:d�%>�:n���aP�����S�'��B(�j�C٢B^͈�&M�8�`�ě�?��y��)N�)`y�DeC�鴵m�4a�a#��#)��DP�'7��!2���Q��'l2���cO�yʨ��i�1Sp@��'�:ѐa��_���l	?
�ց�G5-� �%-�C������\+u�Y�O�-���S:��k��,����΀('쀷2>��E���\$\X��]1���(���0�� z��$��if��VA�:)�\=�b�G[��wTj�Bpe(��dM�T�������`� �eK<17�I`�di��J�{gj�����#04c>���J�1&H� ����51(�05��H�(K��K��L�%BD7�ʁ��#�XC�UZ'@t{��*����`"]�3F�Sr�DA����#��I��F�<H>���
1c��r"�t31�B/�Q�Z�>6�J���5$��
�r���ӓm�Ɉ`�YS4�59���Z�)��ɕfh@�Ч$�cR��(�7�d�4��y��]k�gB�p�ș�J+D�|#�a�@q�ш� [OPy3�/�$�C����"F&��)A:D�p�賎�qKd	j��++S!�d_�/"%`G*�y���K��ߺt���=��/�:����Ib|9g�R��4�1g$�;�C��$q^���B�){��[�)�=Q8�C�ɖ<�9j�K�2V�X0��G<y�>B�	�!H%p�+����q�sDH�X�B�ɱ&�D��h�h� -��G�XC䉑v^5�FbW,N���� Ӧ@�
C��6&�x�:#n����4�δ"D�B�"�>0k!�.��HP����B�I* ��yK��(A���Wčw6hB�ɽV9��v �h��oK8.B�I�	�<Ȕ�m�|H���>�:B�I�]u�]a� )s8�rEID*�2B�I E���+@�6���c���h/ZB�I\6=����.d�
2(]>I�B�	/h̸gd�!@"����"��C�	�V%����)C�>�m�DZ1C�ɷV�RƧ�=A�xMK7f��T��B䉷b�J����5LJn�xg�$��B�I4�,����N�~WhSG�hC�ɓ"W��X瀂�>�Y"�MsIC�"O��u� �	<��1��_�!����"O��qg���l�ށ�v�H��a�@"O\���@H�e5LHg�XI!"O؀��gX?@��x�@䀱\�R�1#"O� (���p&���柃<���"c"O�Q�4NV�U3p��&h�.�pp"O��p)��}_���% H�i�>-u"O.Ec�
҈0�lA�d�X7.�1�v"O�5`��4HK� ���TF��Q"O��2w���E��P� ���'
����"O�x)�o��<���(K�P���"O>�K�ATT�yXu!�������"O�(aw�H �-!���EӪX�p"O�1�B���I0���0����V"O�ĉ�E�.^�>4�r'šz�I��"O�	+Qb�8*�vA0�H�/Vlz��"O0E �@@�Ga:|��_)3T=d"O~:����X�b40�Fݾ���"OLԹ+m{E���eEؘ},L(F"O�H�gF5A'�y!�O�#��%�0"O6�+��L/6*�����ճe���ȧ"O�ШE���t�\�7#A�r�Z�7"OM�FM�,M��}�򍐙%f��:�"O�2��x ��lE q�d��""OpR�@Z�>�8
�IW
�H�"O&����
��"I���R�	����"O^ܸk/fnU�� <��xU"O��QJ8D�uSEF�>b��T2�"OAS�H�`����� N�g�ZqP�"OLM�$��Ճ�o�,g�X}�"O�qg�	Dp�������)ǔ���"Ox �ƉH�Kθ���;I�����"OΠH�MA�}^�U͇@j< "O� X�+F�;ZP��7LBoFh+V"O.ܨ��V`���c��>����u"ObU)�=Y���,ģ>�ҝr�"O�tr�nA,J�،Q��`�~`�U"O�P;v�͚̄���DEΌ�xs"O��!��	:A�h�B�J_���+"O�S�b�.����vd�zzY��"O2}p�F��CX��"��(
b�C"O�ْ �E�_���Z���$)EL*�"O�ʅ'�"��!�ī\m
q��"O.�q��a�f(�S�ѩdoV�U"O��s)޳S��SjQ�P�0�"OTu��b��%� �㈀4Q<ȩ�%"O:ȱ��>n5r塚�b$�D"O^h�S0n)h`��M5���!"O�ĩw��f>�%'B?��q�"OL(����,^d�K�珗(�"O|��ԤԆt�z�@7� ����"O���b�Q��8�蕃P�Rh�<�y�K�������	��"Q���y��Um�PM��F��H��g��8�yrLQ`�lTF�@�{�(�c�ڴ�y�l��%JUI���|��8�s����y��J�5r3fM�w'���kڷ�y�넨V�B<� "z i�	�yB��bS=�u ֟k�2�څ���y��#}*x�a��1`�L����6�y�ȨO��i�1�B�;z�[̆��y"�Hy#g�=�2�C���y��;`d����B�֑۱��y��U�><���E���Ȱ���y2��/�|L�W ƇF��<x ����y��قP�
���ʃ%������y����X˲iW3�\���ߪ�yG��5�Աq���>L6t���ŕ�y��ʯ��d�B�E�	C��Ò���yR��\��x�iH/�J�A
�y�	��pqд�,β{�Z�2��/�y�One������"�L�t
��y�N��V�V���$�2iJ�����K
�y""�^�D��1�� �SL��y2$�=*�P|q���9��p�����y���f�6D*���]��tC��yb�	 t��Af��rp����y�̓91�(�s��v��H��\��y���$����F*e{F!q���%�y����!��އ$��irȇ��y���]V�\���Մh����O��yL�u������2{d������yr��h��u��ER?����+�y"K%TG
�k� �&R�B����S�y�F�y_
�p�n�M�.-��m4�y���V�`�{��LˠXX'�y���:(xY��ԃs@ � @��yB�D�Z��M�'�y���҄�y�'˚(��"t�I ,�6�sG���y2�  7�|`��1j����DĂ��y()���sPe�:��xb5��	�y�� `�����ϲ�Ќ9��N�y� DІ|�7.�>@����G�yb�94K�Z'�h� 0�L/�y҈���D$�D��j�P0�+�4�y��~�!"E�d��9pGh��y�G0��P��^��ۣ�D��y
� �����VlXy��O�	#o���"Od�Ѵ��I������zY��`q�L��L�=����O�1pӋ�`f. 2�L��T�!0"O��8�`@�Pl �D�Eg�p3Ѹi�@���!��|��݋~�T��� �ky`��H7�p=)�Iڟ@�9��e���BxCz�B�A��f �@��>D���vk�Q��u[3���t�0�ɍŜL�Ԉ��Y!?q3�i�&	5Re��N#��)7� D��K7"0^q�HwD�c5`(!�߹r/:)�EG���!���q��'	Xh9���w�	�@O	�/���Y
�zH,u%o�.�b GEF�T�P�� 7z\���٤u^81T�A�4	��I��j0�F';J:�3���[����7��;v#��pR�NMq�h �B3|�|�[Wb��ph�B5n��3���I3�YS�O&l�!h��KI��ۂ.�l�֍(7�B������پ)��X��k\
w�6t���:IL���*���λ|�~(�r�
rP0=�d���Vi��MF�\�f��)#A?67�D�D�@`��ʑAP0d��C�ź�3�P�t�~x(��L��ɗ(d��qnRk��Q"է��H����DV�I��$�U8-Vܨ@�Q�.T�|I1o�8}G�xc��ӿxY�取񾑓��5"^0��ቀIAt� �!Y :�Ƒ���[�>�nc������,\2�abL�b�#��>n�肅�S�z���E1O�l ��Ι�or��B�M���xҪ�>�}
�K �~ݬ�� ���J�~�S&r��w��*�����ꖃ=�Ajw�@���������" �"ɚ0N7eѼ��rb
n�<a������#Ɯ�!�\,����67
�`��Y>f��Z��3l/y����R���p���B����k��w��� ��ֺ�X}a�2lO<�r���*,J�U��(�5V�����S<ja`3�ҩI�T8��E��y�#�2I<��t�c�1UjԴ8�,�i'�DJ,xc�.�	�k�!"ꔨip�Q���IrCHΑP�H��� G7��q�jű*��0�Q.pB�	�\-<��d(U�<��栈������/J�qO�']����>���:b!��&�6ܰT�M�$���j`"O.D+��Φ8��иC�_Z �P�P��c��!LqOQ>�)A��!��勊 ���)�O1D�y�F��]w<�hԻ�^щЫ1D��ѯV�9r��S5�٥n�
iuJ/D��Z�%�ҡ(1�P�),��0J1D��h�`��4�v`��ѽT$��p�,D�`� ���3��@�f��� 8@��&D��#�!���lèQ���y�Ӆ)D���g,V$ �q��<�h��J;D��4��Wf%�N�y7���J;D��R�a	a���B׉H�s$�!�f9D��&1d�gh\gMXi��ּx�!�_	E�pb�.;na��A_�Z�!����œ1KF%C��D ^� �!�F
5DÇ˞�@�������p=!���"hW���G��ԀA�`*!�DϝaܜM�*����Ta�	!��oG�u�"�C@1�(��L�M<!�d �.��-Q�)>B]t���:(!�dL&i�F`�IȄ}T��:���<!�d�
P>�s�\� ̔��H�^!�I�&̔��S��������!!�D��-j�02�ݤ>
�`�$( 4!�$��T���r7M���<�$∰7!��z�H��F��{�T���b�O�x2�<��}�<A�m�: �(Q⊧1��9b�UkܓX�9Ê5O���jTq�T�ר<=w��+O�\��Z=?uғO1��ɘCꕂn�Bn©d<̚�C2R�T=�
$�O�y�&�*< Qˠ$�(��A:�'�Q�dɾW����,rcǡi��I��IR. W�D���/�u��!aǏZ���i2.��,�1� �s������>M�`B���*�'��>��J��>E��M\��dXj�F�	�����D���Or��)H#W($�K|r&�`nf�:�!L<|h�� ���e��y��4Q��� ��g�GŊ�3�[�<�s���#V��'�P���,��G�NP�O1��-��]-n�b�X���4{P�Q�Э��p��V�ֈ��?� $)�ٴ5H��m�_�M0��#P���6C6L��E�?MSF-F^�q�>���^�Hw0�jV�׀�҃�A ��?��^�M>B��F�I�b�A	V>/D�XGcoL�����<�t�г4}��Z�� ��
�` �B=0L֣?a���l2�	���O�<w�a;3@��.&<5�@�D4c����ONpB�ak����qO|�ZU$�}2���a`p5q2��hq��B
:�>�R�$6�_�^) ��(/�4���
�l�ZaВH� ����
���������sj��Δ� R��hj��ݨ���O]�xZ�V̓O�h��F�O?H2��E���F���z0TD��iI�{��`��j��Cu�K��V������+�O���4	�!S�V̑��M���a�'�H�kA�^ 2��'��=�ڔk���֫ɼ Ę-Ғ"O01�JòvnU�5��	����r�x+�V�둕|���n@̜(���2L�H�(����y2戉}�� Y�M��F� @coϲpa��4��'�x�g�DS}�r�0��z�L�Ҹ:�p��AĄ���,��k`d��^t8t��KT�lX`�Y5V=p�JTƂ;j��ȓi���*`� �	��� �=x.��@������R:��#�+�?f�\نȓ7�j�1�c�v��̃�G�,�N!��6lV�Ʉ3&;z�e�dZ��ȓ$�����;S���X��XXΝ��%�6����Z�&J�@I�le���ȓ[,���BB�Ph*�SӏϘ&<0���D6�єD� Ne\@�ӽ��ф�"�i���[�>�;�N�9I؄�\.���p�% �b�:�/�43��ȓ09�@�{\(�
��Z-w��ʓ ���PG��<���r�'��WL`B�I���	
|����'(�C�+c&�Qq!삓D:�%�Ё@u`C�I18�Q�EΌ3e� �Vd4G�C�ɛ ��TB�H�����c�C�I�NR����J�$I%�A;�C�I3|�p�V��|R'�<	;hC�:N�ұ�c3��4��<A4�C�I3H>��@U�R�$3�H�d�tC�ɗ}�!au��3$DF|� a~C�	1?w�|(���gZl����92C�ɯu�H�z�jD> zPLP��C�ɀ$�H�G`Ҥ2�
�z��\�	�B䉔T�ً��^	=��QHf��?;'�B�I�}�pd"�	8|~��2"\�dC�	..���hQ��oC�� ��۾Q%.C�	6� �9�/2���q�ŢH�B�ɴ#�phr#]D�2A�P�®g�C�I�y#����/B+WN=�"�\�$��C�ɇT�Y�Ɉ�b�\��F!��C䉒�{u��$�p$�a�Y�k,�C�I�@�>Ii�
��/(�G��%t6C�I���{r])XN��Ҭ�2C�Im8m�.�#�V&��T�C�ɂl���P�j�E��؁�G͇O��B�	�ֺ��VOfL��ڕk�F�2C�	�5�D�1M1 �h�f뉾&�JC�I�S�!`,��c8d�B0/lNC�	����&�P�[�R\��I�uN�A���fmY�%��[�Z����2
/�	1��H='����""U��!�I&�6X���Ɯ7�&L�Cg�}$!��yFFT񐫓�&�٢N�T�!�̾VƤ� fG� �䌱'D�=~�!�ė�q6�y����r�!����@3!�<2b�ѓ%m�7<oDԑ�a���!�� � `@H6R!�J��P$U{���p"OX]�O_�"���zQ+ܴu`�[C�����SS��� �����u�.r �V57�hbf�h�TJV��ClQ�`Ø&gt���%d��E�ᓵXd�	�*!��-C���8^}z]�5` ����-��d�
��Ň7�r��#[F&��BM�,N�����=OZ7�_�M�Չ�9����		T��hHa�?E3�-8A�Q�v��D���[$����)�'(^p$s0��$U,բe�,Qi⹊�%�B�BB�m~���u>er1Ύ6?Ӥ�+� �R�����l[�4`���b�aR�^Kt���ӟB�A3 �r��пF���4;i��@£WN�h>�{o[%m���E��;zȢ�:�3����zɠ�2�Z��	9B(a[S�.t��pf\ +��C�I?K}��RUc�$lw�z��-8��|�xB_7y`�h�f�.����ě�y2��kXic�����HAԐ�y��@.eN��P���%�F�%W��y`Ě>��@G�,��;���y�Aɮ���Q��qRP�$��y2��6,�)E	�r���u'�;�y2��6VЈ�P�eɸc����I��yR�2��J��)odH(�@�y�c���� ��Ð(Q�H|Zr	��y�K��ZA��B�HԱQ�4�y"K�%�p ;�/�0/���*��y�n�=���,K�N��aЌ��yZ��y��Qz�$)+����.$�B䉽$g��#W�ϣ*U��[�(@8Hz�B�Ɂh�RL����'Ki&��s	�1&�FB��5v+���J0�*�ddI�h��B�I�EͶ}IE��/L[.��r��+Y��B��#缑(��HFFl(Z�� t�B�I�Q^򄊦�Ɠ$�.��@þ��B�I8n�<�;���t"�YG.�r��B��=ja�T3t�#h�H0���Lx�B�I�=�|�r��F"z
ZyP�Ɯ�+�C�	5ª���Ҝ�`1��h]�dG�B�	�N/��u���^$	�-Z=J��B�I(]5h���и �Y��L$P��B�	- O&l��EF�0������\tB�	�o�&=��B�l݊W��=,DB��MU�!�f�!i�
h�wh]*EBB���@�E�\+'b��#Ƨ�;{�6B�ɪ�<��ˏ�I����3[�B�4_^D��U�`>ʖ�\"I7B�	(
ol�id֖".�RE,� �C�I�a�9���؛|�q+`�
��C�ɼ~Re�b��t��re����C�In�n��Mʶ:��(gEU,B�C�	�H��X��BU �X�o�8X�C�	 [�^hRoW_��0�U�\Z��C䉀���µ`�	&א��u�({C�C�	�o�Ż��Ze�X"��9d{�C�j����$K
=j/jT�(Y5��C�I�[D
|�$�ԣ}�\�	D$ܬsz�C�I�2P{R��C��:�fڄ[HDB�I�z5�}�Ec�T�.qJ"&�(L|C�	�d�ć3z ٢E.��>3tC�#F���s��� �`�+̀LXC�9�8���W>K��؟J�6C�	KKv���(|�@AJ'a�0rV<C�5�X��C�X�9��E�b�C䉲Z6FHxG�G�%Fr	rF-� z�B�	:LIx@�ћuh� �˞�]hB�I�9��jB�0J[<-��]?�jC䉹'0؃�O^���҇�N�l_C�)� N ��bǊSv�kR��$Df|dh�"O��"Eҝo���K�u5�Jd"OVu@wfH�o�le���L�-����"O��愙�"䲔ꁄ%
��"O��W�ݪx�hS���N���V"OX|���f�R�bw��'�r���"O@�R��H�X}��� �$N��"O���U�>Ӫ�{��I�1�� `"O*�1�� $�؝�䨛�(�ԝɃ"O�	��@C8`;��,K��Ad"ONM�6�+3VLᖁ[?�r�q"O
�c� N�/��`� V�� ��"OTh�2��,��4��N�c�����"O���ᨁ�v���-�B��0�"OV�	DD�%� u+qK�8g"�"Ob�ѳ��F�LA�ъ�+`d�"O�E��:s�P���Ӕs\�LK"O:�� �ځX��!�u����0)1"Od�Q֯�<}�(*$
������F"O�Iഭ�9/��	C�#�V�&�z�"OQ��ğ�J ��@�I�x�"O|LzVO|oؘ�j�(}b �6"O���O�k-nLB����N���"O��an��:ghD��$�� �"O<u�ѠΠ>�V��Э�!Xx*"Oޑr��76��b�L�98o0�{�"OTbv�,v�t-��AD�d��@��"Ov�X��ߓ!:Ѥ�[ ��Pr"OJ���m��D�.���Mp��dJV"O�ؙ��׳+�����*b��tb�"O���L9 ��d�V����ڈ��"O>$�*X-�r	�CC��I�i+�"O,�s�	91�6�p��E�i��Ujv"O�L�TG��$���*�Mڝ�<A�"Op9PӁ������1lS�7�2���"OD��B���X{�Yt R�8�`b�"O�U�񬌱=���8V�5�h�{4"O�"N&AĞd�wo@�S�$(��"O��cL#z��)��ǐWَ �7"O����ճ1��I��)H�yo�t�"O(��Ӿq�0Ƞ�Ρ~k>,��"O�բ�n��FX�B��
A�#�"OЄ��[¸�)p��a����"O@�{�)H)0�.�sǮ����=�"O�%�ą+�X�C���|���"O�剧+�{#�4�2�LcM�9�"O���ucI w�� "K�8B���"OF���A�J� �ʐ���L�X;�"O}�t.����B�@(L��� "O"�DP>O�5s���4X܎�rp"ON��"G�OF�t�rC~����"O�8��Ѧ>~�b��I��Qz�"Of���
K�iy��J5z䠫C"O�0�A��cj2H�UO�Y$��8 "Od�Z�+w+�f�dc\�+�S�"Ol=���v�]wDI:��YӴ"O� qd B�&�X8caㇽ!��{�"O�Px�"��)o���FE�8ڠ��"O�4���PZ �LAf+2?�� ��"O��9Ǧޗ1�-���.	�25"O �J�����|`#Dɝ�M�����"O��XF�_�ϼ�+ǈ��2�8=��"O �獝S��(�- 3��`S"O��I������kr�Q >�J��5"O� �H���EVʹ%A"��RX����"OXs��
���1AO?*1D���"O�E��'R	m���I.�4�����"OfM ��]�"�D+#-���T"Op�abgȀ*�p(ҡO$Zb%
v"Or�c��QX���☉BQ���R"O��ԢR5^6BS�.�--���s�"Oh8	�Ǘ�b_�<���H�;���x�"O��"�@3 ��S�ev��P�q"O��K��\�,(蛄cG+d�X�!@"O~��(�"�����
�r��2"O�kk&<�h`��C�K�vM��"OPD!UL_s2~���b�����C"O��1�"�Q����oU	����'"O@R��)�����E+��͢E"O���C��{v�3�� C_x��&"Oҽ�cMS�t���P�E+P��"O�C$.��Ǌy���Ю�aZ�"O$��6g@
k�,�b0̀�cR�*�"OzE�Po�+�����ʉD��у"O�zr��7+Jo�47�V�H�"OV�	�+�"IѴ�S�L�#_���"O��@/���mQT�SGJU��"O(4sk�6m����(�/(� "O���oޢ,�\��ue���W"O�$q��C8qu�d@Z�#U"O�������a`�i�#=h�C"Oj�)U�����$�A��(xQz"O�`�bg:b=!&�O�ƉS"O~����')�]K����F�h�"O�l���1s6��c�	j�}�B"O���k;7��̣��0_@I3�"O��h�*�B��� E9I�My "O�D�g �:BȐR�u)��
�"OVDH�+ɈW��v7n5�"O*\8�G޼�V ����1��"O�D+��W�H�A�J0i���y�"O<`�7�Ď>&�8F�ɤ˲](�"OKW�M:���b�4A���1��y��+W&�}kv�H>��sbֵ�yR$K�$��/����y�톓Oi�4Ұ)�'=}��a�X �yR%Z:�b��I;;{N���ý�y�F�1n$(ʶ� cXvHӃB��y�Q!C���'��*��0�B��y�Ô#J���d��#Ԥ���ױ�y݁M:��F���1��nH��y�'W�{���獟 ��mڷ�_#�y�!X��� sG����Gi���y2獜&�<�K��\�NU���7�y���5���c�FߏR���fȂ�yR
_��!��!ȉEO�l
5J�8�yҢ9R��}@����?��8rCE�'�y�a�?)���΂�>�,Cc`�1�yR��(}�9��/�>r-�B��+�y� ߐK6\Ȱh�jB`1�f�ϝ�y�h��.�*�A�F�bo�y3&M��ybfB&[�
�Ǣ�-S�t;�Ř2�yB�[|4����6[,�{���yr̾)�>�R�^2�y�X-�y"��1>5�iX!nƟV!49�!g�:�y�	�ޡZ1��D���f"���yRm������	 �xY��KV��yBDځ4�� C�� �&%VŲ�y
� ����1!g��Z��"��l�"O̹gL�D���p����씩�"O�y�` #D��1�/�:�P��P"OH@Q��)o>��m�*:�VE�"O�5�V��!�h�3���[eeA0"OnP�0��O�p1��K�TTN!�"O�	X�P/�0��
۞`?�\�"O��p�Lޚ^-���Ɉ;&d1��"OX`R�o*��B��n �D#"O��ą>²�
��T�M��	�s"O�Y5e�&B��:�͕/�␲�"O���e�)Yrp�P1�R��Bw"O
�����y@"��J�hB"Oа:Fn׳G$ �+7�{H,26"O�5qQ G9$2\��C�!2
��c"O�p��I����C��1\�C�"O�H�3�]6"X�d�T�0�3"O�ڧ�P���a"��u��Ru"Oּ0T�س_�	"�N34�X��"O�5��N#{g44��B^�M3�\�"O������5R��"�@~~$�#"O1���\���'X/DH�\cD"O��a!��,ʼY���3�5"O�XbP   ��   �  W  �  �  �*  �5  SA  �L  X  pc  �n  z  ��  Ǐ  Ö  ��  ħ  
�  ]�  ��  ��  #�  ��  �  ��  ��  F�  ��  �  ��  �  % � Q  {! �* t4 �: B nK �R >Y �_ �e  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m���'�Q�XI���M�\ ��cI
lx�2�>D��c�&q��KQʇ� z�d�D�<D�����((�[E�/_���)��<D��8�ǡ��!D�'����?D�����9'�[歌!����=D�L�끐Gp�u�C��:r���ȵ`<D��1b�E�E����b�3&�����#;D�� c��R.0�@�J:=�t��(>D�����ՌJ��]d��	����V�:�d2�S�' J
ssc�+@����!��Y
I�����i�M�+L�u*Yr�]��.faR� Ĥ>���0B���H��ȅƓ�x6�S#VL]A��aרub�'���A��/$2pt���
T���'���c,�.������]* =A�'��k���1}�`�����]��!
�'pP^
DL�q�����S����	�'�`y t�I7��Yy �_�O�~�q	�'��`+p��`^�����X�;�$��'7�[F�2PJ20���\(�ݸ�'k@@����%AtY{'ҽK� ��'<ў�}3jݼEG�!�a0w+:�) �S�<)��*H�@����-w{�M�W$FS�<aE�*�*�����C[D8���N�$��k�XC���`��G]���b!D�t�@NX�Qd\x2�I���c@'*�YQ����i
2~_|�b�씻)^e�U��9H%!�$[F
�(�����8h����'nL�e��'.昉�d 	+��]��'!�1�5J �8�^��F�#)�q��'�ȍ�աQ ^��H�� �(��'l]����
�\��ՌT���P�';������@;��b$�?_�P��'&�3 C�D�^]�6��XZ�'#2����H�'���p��6VO8���'�@��RA�aX���lˊMgP�
�'�B�Qv(���fM�7`��'��Ik��4($q[��Q(=6���'�����Y0w�<P�RŎ1(�A��� �Y[vDJ[t�#��#:h�R`"O�\3g
Υ6�q�J�V'�-��"O
���h��m�`�d*ܑ~&z�v"O�|3`!��3��E*4�G.	�����yBJ��U���� �B2"�Y'�I�yB���G�� %l"�:}:�@��y�@^�**���"�7|��	�ˌ��y&�%)�""�!w���K�J2�y"���i-��i!^�s��H��y� ��_4��.ׯZǊ�SU]0�y�`�%or`ň�DV�x$d��yB$A(ڭpn�$I���Iq����yr��-]��Kc�ٖ>�b8P0[2�y���5^�س���
<%����D�y��F��P�V�=.& �� �Ң�y2g�6$��2���u����	G�y�οq��nc:�W�7�y���f��9)`i˚|�-y��L��y��R�N�B�3�!� *	b�+��y�N�} ���` �~�~�p%�;�y"F59��haVfqR�tR��y"�9*x�c��g��� u����y�FȦc0��eP�[���`�-��yba�a��B۲V�œv�J�yG[�5�|x�D��I� � F��y"�	R0��JL�J
d9Ď߫�y⫆)Cs譐G*Q�ʄ� �
�y���)AB��Q`C�D �,ź�y�"��6%*ɤ��p/�T��	�y"�J�1�����R7f�~Y[� �y��w���*$�0ff~� �� �yb�i2��*bT()s���y�醏�	�8Z����r���y���-G�4(�\�~ z�"�P�yb��Bq~�i�jQ�^�R���ؿ�yR
����'��Xu`e�bɛ&�y�M��^��@U"�/K�4���̸�y���'J���2C��B	zdA��yB���٘�W��N!�@��#��{�-�)87J�3��_lA���ȓ	[�)2�-C����H�&j���+��5 7N֓N�D�JK"`$B���^�����{ �t���BtՆ�z[>e1# �O8�ّ�HAe�$��`Ê(J�'0�=�&�>.��l�ȓ)zV��CN� %X$��.�8Z.b܅�+��)��A�Ky@�5e�2t�$i��7�H谊�A+�L8�M�g�D��I�( �fD�e��k�,T=󾥇�0Q�}��MYMV`��ڌb�Ve�ȓA�J�{���bHLi��C= |!��0̌	GG"&t�'ϛ7�Ҝ�ȓba.��#�!,J�mra���Zs�E��AQ@D�A��E��ա%� �:o޽��
�U��ʤW��-k�&�#>T��,3�۔��}�f�b�
.�T�ȓ'��T�e%I�b�pY$���vy�ȓ$������P�zj>Q����$Lt�ȓB��������s� �q�A�H�r(�ȓAW����W�X�j�*��<��|�ȓP�$�k`��i�.�ңi�|�n���- I��a��qr h��Tхȓe}z�3�MG�f��xZrE��U��S7���c/�,Q"ύ+IX`��S�? Ԅ�GM;e?��ʇ3��"O�̫f�3\������Նn;��""O�5���I�Jo�"�f-�v���"O5�4M*d����͘6��M˦"O��
��U�z,)b��z�A
V�'_��'B��'b��'t��'p��'Qx�Fe!u���1L]�%*a�'���'*��'A"�'72�'���'�l�0VH�,6' ��CS�Li�J�'���'���'��'��'c��'�*����BR6jii�&Q BazU�'"�'tR�'�' ��'
��'��#�%D�I�|�G��{�`=ig�'���'ob�'QB�'pR�'���'/��/<��(
!��Bj���'.��'Yr�'+��'�B�'H��' ��h��\q�-�'*�".t��Q��'#��'��'Kb�'GB�'~b�'-�Ut
d{b�iG�;t�ˤ�'�b�'o�'m��'m"�'~�'�����n15� "QD�2x�� �'"�'���'%b�'���'(r�'�^��GP3qf�9��ҩ�B����'�b�'�R�'J�'���'�r�'��	�A�jDf�ǈ�,����'%��'��'f�'r��'���'+#���S��<K�K��z������'B�'�r�'
�'���'�r�'ȹ�u,
� ����ڣC
a��'���''��'f��'�2�zӸ��O�Ԛ4*į����_O(N�a@ my��'4�)�3?!4�i5�u�,Żdu�L���_EئP�RI݁���L��e�?��<��[B䩩`��W�h�!�((q�.����?�Si��M��O�ӫ��N?c���\��a­J�7m:5ɵm%�	�0�'k�>!�P�Ms��p���N�T�u�aC��M��,\̓��O�p6=�Q����4m�@"�ũkD1��O��j��֧�O��Q���i���=&�e	���K��A�v��2Nq�dz�ȸ�n7z�=�'�?	S"ٜ��r���(>z�-0(��<�(O��O^(o�)�Dc����R�>���0g�תfb䉹��Z����Iޟ����<��OT:e�؎���]5l�
�QC��,�I�R3�%P�&�S9R2�����K�iD1Wä⡪�!X�x]����zy"X�X�)��<�S��s[�1c�*5܆�d�Z�<���i��H�O:Lo�u��|����`��ӷOG�� H�M�<	��?���KVh���4���r>�H��g��&=b<�t)B�C7X�����0���<�'�?a���?���?���F4;zr�{#���|f��%�Z���ċ̦�&��� �	ߟ�%?�	*�@f_�+�1����P���O�1m��M뀑x������iQc"W�H℔��a�2]�d�dH`�N+[&�E�A�L����I��/���X��T勢�*i�
0�E i���D�O���O`�4��|��)X,G�BEYz̓��D�T�ʶÆ��y��a���Q�O�nږ�M3��iբx91�>=L��,�/2�9���L��>O���E��e�bU�2��#H?-)�w.��f � ���& �;��X�'B�'+b�'b�',����"hS�;MT�6�[�D2QP��O4�D�OΥlZ�j)�'i�7�=���.����Ӗ+� !�`�vz��$�@ڴYc��Oհ�ָiv��3(�ZF(_ 6��AR��Y�M`�*p�(d��$�<AE�i��	��p�����	zPp2BEB��TM�AǏ�B����I��'�j7͆�8)r�d�O����|�w"���H�k�$c�:\��k�K~b`�<���M뀑|*��li��8 p�����Z�bϖQl�G�aӾ1�'|���
B����<�;H:�"�ʗ�I������&:�i����?����?��Ş��$�ӦE*�&G�v�4�x�����Pu�M�Sp��	͟4�ش��'b"��Mc�.��W������ ;�J��� V��Jz�I���l���W�Z6m�t�+O�"�kόP^f�)w�[LR�uS�DA���'�R�'!��'���'��ӭ�PY��(�ఈ��2v��4n	�9���?9����'�?!���y�!�X�\A�#1Rj|��.+_07��ԦM�I<�|b���"�M�''xe�W:x��k���q���ʙ'~��w
�y?�,O(�n�hy��'2�	�������BƄ4ғd޴���'�R�'g�ɲ�M3V`��?��?��iהh*4Z2C�C ��Dc���'�d�>i��@f�	$��rb�(C����.I3]�ƨ��<?��U�p�<��49��I��u�o�f?Y��]t�i�)˲y�F�`�MI�?v ����?���?����h���S�>	:�(�cO�G ��*�IT7�$��Ǧa�.ٟ��I��Mc��w�N�Cf �$�L��,K�4̡�'��7���1�ش'>,p�4����4�`e��Oذ�C�*Ey�l\�7l�A�¤Y���ٴ���O���O����Oh�$Q�q�@J��	+ܲ-��@�1Ax@˓6�NA���'i��闀*��!JpDF/�(Da��¥���'r�6�
ԦU�L<�|ʖ遬�Jx�q�E�6+z��4������4e~�I'A��`Ht�On�L���Q����j��;&,񲐤U
)���r�ȋ���I�(�I��Sgy�Cl�R=c�%�O�)+F��|���  ��XW@) Q��ON�n�p�$���ݟ,l7�M�OY�<̒$��#Z(J�X��LW��mr۴���3J�{�O�I��u���� ����wR�i'gNS��57O����O���O����O�?9�pK�RA�u3 �]�N��<����`�ڴcwr��O�j7-"�$�?<f]i'8;���p�&�8�1O��lZ&��$O4v�7mo�P�W�P���ٔ��A1R �R�t��,��A�O���PD#�s������O�$�O���CC����&�&?N0T�=3N�d�O�ʓNě���5G��',RZ>�Yp��"v
��X$���X��y���=?��X����4j���=�?e��`�2���iƗ���ª_���-����?m�N]�	� ���0y�Y����Ny�Ok�ޤj��3�l������㚂V�����O��$�O���ɯ<96�i1^�2�wOV5�iZ��N�3��V�C]�	��MÎ�i�>�g�i;d�mTp��3 iE�!�	:�ovӤ�n� x(n�u~2�p� ���!�剮!(p�"��Y��٣�3���4����O����Oz��O����|�h�0if�s�YE3���G�)���~j��'�������]�2I���� ӔHVȻP鎼-�!۴tW�E2��i5dv�7�c���G�V	�<�L�_*̴��Ko��P(�����iyBB`�
˓�?i���b9��.���2���e���!��?���?�/O�to��D�`�����<�	s`�����_�J�
�%L	#	�4�?�R���ݴ ��V4��C�n��eօ1j�b�C�#j����UԌ�t��G����'�,֝*K�B�O��H!4|��Pˑ
���)Pd�ҟ���ȟ��	ܟ�E��'�J����Q�Br�E�n�=*�����':~7̓ A��$�O��nO�Ӽ�S�@;7���\=>���W���<q�i��7OϦ5!$D�ۦ��'yz�{��?	hGD���!P����Gv�<+�ϔu�ɘ�M�+O�$�O����O����O�`-���f�l��c"@6S���A������'I�����'����Ѧ�<8ê�)�d�=�t$0`l�<���Mۖ�|J~R��MB�NU�%���Lw�Q�W�ڊqC��TOT ����q+����S�v�xE��^�ز>lWN�G��<N�8�����l�������ן��xy��uӴ�rL�O�d���!~Rj�hW)�pzp�Ck�O�	n�m��[��I�M�ձiA46m��
�^��iڸ#x`-��Ϛ�<���rVf��kN���B�|u�,O�=���>q�ԃ���{���B܀'8O��$�O:���ON���Of�?y)��9!6�1����b�:&�Vy��'��7��in��OV�l�g�%p���Ƈ*o����j��5#�PJH<1��if�6=����Dq���K
�ȡ�Gar��C��@¨�5�Z�.�t��W9��d���y�'7��'�R�'��U@B�˙(G !��K�ip���'/BW��ߴ �$Y���?�����"?��<�C%+"U�%	�M*��9��QߦUP�4-L�����(d�|<[��N�;uLp7��- "����Y�z��4�ν<�2��-���;�N�ӼS�U�
� <��n�*lh9ZfB��?��?A���?�|�)O��n��i*P�щ��0GB�ڀ�0|�jĂğ\�I��M�"j�>1��i&�J�IQ�Kw��Dg��2�n���aӶ��_�$��6-~�@H *�'E�.��So��uw�'���[��V��!d`6�!�Q��?[���IΟ�	��	ޟ��OX<m�p/�	��U���$]���`��u�.<3��O��D�O�����$����u�;��$XI1�Vq��M��|J~�`���M��'���:��.�x!`���6'��I�'u~)���ßkÖ|�Z����韠`�������R�b!�Q5�����O����O�����̓K�b�'|�-2� McGA�G�z�������Ol��'7��¦��M<��FC�S�8 ��T�T��(�l~��:B�FPJE.��O�@L�I���ԣ\�İcqlT:��TƄ�sb�'���'~��ڟ����{�X�X"�9��
�HS���1޴�����?	��iu�O�X�9]*<`m�4v� ���F2���O˓.�r4ߴ��$@*ct,K�';]��P�E��?*�@�F֗#M�Q�5I6�$�<���?1���?����?��,�$��S̍-F�5�ai����$J��I�Q͟8��П�%?5�ɰv9���E[�kQ� ����� �Z�O:�8�)��YrP%����R*Z����|O�9�"̛:��'���_x���q��'N�I�f��� ��N!�lS�ۯ)Y���	ן|������i>1�'��7�1D���LW��Q7o�*P9���I�3,e���ܦ�?�FW� ��ryr
�"O�+dΚE�T��$�1;\��i�I�t8ĴR��O�
�&?��G� ��e����WJ]�<�z������ϟ��	ß���\��6|� 3�&�+����C���Zxz���?��!�������'87�(�䇾��Rw�Xd�.[�G�?e�z�'��#�4���O�J���iB��}�6�9�d�H���k�BՉ.P0ŪBJOr]n�\y��'g"�'2��V��Rh� x��H�]�R�'q�ɾ�M[���?���?.��i ��VAJ@Pc���e����O��mڴ�M#g�xʟ���b��Eր�8&N�5�(iB��
/# X�P�.]A�v��|����OՃK>i�O�<  �JSb�;d\���?9���?����?�|r)O�5oZ��:��PFZ�1����`.�mޤ"���蟘�	'�Ms�2ϣ>I�C�,�z��Q�@$)��5���0��&@��V�&��<��.v%�i�<� z�IF+���m���Fu
�`�2O:��?���?A���?I����U�4���67D�a;�e��k��<l�s}Z������[�'fX��wV � c�\9�p��<&gjxe�'��c!��ƹ,	�6mg������N�X`�T��
R��p�,s���$�E�J@��*�$�<���?��,%a�ԥ+%���0�"�?����?q�����\��՛W$�Jy��'��%Q%g|��q��Z|����n}"�'R!-�D��X>�� !8($*t�_e��$ph<,ӇiѦ��H~�����L�	��Zh
3h
���-�����rC�I�����s�U�8�|I@g�^"_,�t�I��M� K�/�?Q�%���4:���<�@(@t��2{�0�d3Oj��O�(oZ��fxog~�D��=L�a�'�TY;�	p��b���5��A�K>I/O�?Ic�4 f�r�+�*@ll+�c~�Aqӄ̛�-�O����OR�?�{��	��&�Gm��D�¥iĠ����d�O�D-��ɏj6��I�$<@�@��>;πM�Цy�JY�''�ax�LJE?�N>y.O̙��ƽ{
�ՠ�@&c@�27�'�X6��QR��d�|X湙��_f��-�!�[�Ip��ڦ��?��V���I��i%�h����V�Ɇ%��,�n��'�t�2�a�IZH~��;V:��z���4�Zu��i^V/�i��?���?���?����O��Y��h��$J`I'(R*3A�'��'��6M�R'�)�O�m�i�6<^Ŭ�6���yw�&i��;��$���OR�4��ջ�u���l$����>|O��:�K�y���02N�]���C�	@y��'�R�'��'9������4j�x�0Ҫ�����'x�	��Ms�ߜ�?����?a-�b>;l@4�01�IK�<Y�OH���O��'��{��|#"�Ռ*����@�M� �ǈƷ1( ۴h8�i>���O�O���A8m�|�	��e&��A�,�O��D�O��D�O1���rZ����x���T+M�l-a�L�,�Jt��'��v��L��O&��Ag%Pp�&B�!&��$Sg�VdI��DE��Q2 �^Ѧ��'(�A��PR�/O<�Y�̑$'���¢'=L��2O˓�?����?����?�����)J�4f�	���\�4 *��.T+�$mڦU�V-�IƟP��U�Ɵ�����;/ىB�H����&Qǌe�ע��?)��*���O[���s�i��$F	Tδ�r��j�����.?�Lǲlq�'��']�	�$��:�jc	�;�^�ySD�8�F��	� �	П��'��6-S.����O���{�i�b�ڣs2@���nW5��P{�OX���OD�'�h�%[������D���5��g-?ysE���ݴR�O*���?a�ŘeCH��o�ftaS0e��?���?Y���?ً�i�O>� 7G�����J�$�f��f�O��lZ^��I�'pf6m9�i�aXeb�#5X�S`G�R�h�b��f�<����, ݴxd��iٴ��$)U�B�r�O�}��ꞇ=9��j�"�����r�OR��?Y��?i���?q��,^�p�t��6��x+Η1��MP*O�LnZ!_����IӟT��Z�ӟ���/�8���q�"^�84�����D���pٴ����O�ٱC�Q��m��
Gt[T�*��y�ѩ�T�|Q������VA�Ihy)R)[�0J��{k�9�wMQ����'��'��O����MAm� �?Y	S�-�~�y(K����5�#�?�q�i��O�D�'�"�ih&7���r�P�`��,���l������c���Sdv��A��ҹcL~r�;T��4j�>>�+�DL.A ��?a��?����?�����O]�}�`+�!2_�-���(?� 	��'�B�'��7-�� �	�O`�o�b�ɬ0;�p�U�3�y�7'[ V�b���IXy��ܴ
�����
�@�?,��T����)DzA��*�*-�Ӳ�'t*�&�З'�R�'��'�� ˇ� C$���I!v
�8��']�P���ڴz$�����?1���I��^Vܝ(�%W3M���@�}��2���¦�x�4v%���IZ
~:̱H�,N��U	�(�/^��0���Őt�qH�<ͧd�`�$ơ��fa��J�9f�}K�b\�8 
 ���?���?��Ş���ȦՁd�!mk�%r�k�*(��0&Fg8��	� ��4��'���ϛF�D�U|T�A(U��d�бЃA�d��lڮ��n�b~2�ǣM����W�^��dѴa� [\���/� oI0��Vyr�'���'��'��\>)��E�o�r��c�	9E��y�'�۞�M+.�?��?J~
��x���wM���H���[㦋�l�$�O�6��X�)���/?>r6�f����� )d�v�Y�@��yٔ�A�r��B�`Wt�MM��\yR�'vdװ��A��$�,W�Ń#E5B�'�'a�I��M�u@��?)���?����7y;r�+�E���^��'�,�9:�V�}��'����]2�<��%�	�'F@=�D)=?��m�����!S�>��Od���	�>���~����%(6q����50kr�'Hr�'���ޟ�F�I�e�Q��*��>֠�S��
韌��4R �����?9V�i��O�N�j2n��J�ca�IJĄ]�_�$�O�6���A3��զ��'� M`"��?E�	� 6�ʠ���X�P�'V'
���a:�d�<����?��?9��?����5'��#��

t�X�QD ���ަqKQ�Oyb�'�O�2&�/g� 䚁�Y?!�:L��*u.�4͛ƈc�t(%�b>Eh[��ثA���`)V����h�Q΋=�������Oj��I>�+OZ�)7�4>Б�j[]E4�B���O2�$�O����O�ɺ<���i�ԙj��'�@�yWM�o2e�HDj����'��6-'�I6��Ăۦ��4W"��$��;<H����>��$��9����3�i��	6~XTѓ�O�> &?!��K�ԉ��
"Z�xXnB����8��֟8�I۟��Iq�'[*Q�0(��'�Ҥ����= �����?!�:�6���	��M�K>!#����t9uoH�T�F��rd�F̓�?�,O�1:��|�2�2��1��C!v(b�D �u�x�WNg�2�ć������OX���O����A���4H�)|���v�E1#��D�O˓���#�4>��']�R>E2��N�6�ɳ��2
���C0?)�W��I\�S���ȒG�҅�F��?�ܤ�V���gH��y���,Zu�Z�]��*�Bh�d�>a�����C��ȦJF��n��	ퟌ�	ß$�)�Qy�L~���Q�A��#���t0�)����1$�˓}����^}B�'R�E�bg]�DY�T�򎚍2�$X�$]�|
"L���'wֽI4%�?�(c\�,�0�<f�X�RE��U��|#ap�ܗ'fb�'���'���'��S�o�(mhC��9%>���(ZEg��{ߴ�|��?������<����y��C�9�je[fE�:����gݬ���T%�b>Uy�ۦ��g@����)����6g΃�T�< 6�˒꿟�%�p�'mb�'*hZ!�̀)	��aM�TzdPp�'�B�'��P����4���P��?��J�V�@d�ݨ]�|hx��	]�|݋�RM�>A���?aJ>Y'K� ��sc��v�pX��@Y~��.i�a��i�F�����'�҅��rbQT�S�_��X`�B�<g��'��'�ן@��?�*Y;Fi��:�^�Zw�� q�4!t��2���?a�iA�O�U�g8@�e��]�6���L�yr�'���'H���W�i[�i�]�al�T� Γ�:1TD��W������8����d�O��$�Od���O��߅u�.䓀eʚ#�b�� �+d�d�1[�eF� [R�'R��D�'�l%J��ٌr�8���H��n	@��>!бi
66�Vm�)�����c� #xU���pHΙ!�؍�g&�-J�'c�,a�^؟4(ј|�S��K�	�2~�:��Pi��Zg�iZ �\�L�	�d�I��Say��p�qfN�O^`�SGG�tM0�@�@#2Ӯ��1��O�\n�@������\�'ۜt�W.S�"�F��f�̤bF���_(��&�i���t��Ec��Od��&?a�]��. �h
�r�dU�ҧ��hQ��Iҟ8��ПP��ӟ��U�'�t(vዃk��j���>-�%���?q��k�Fo�,��IIۦq'�p�ގa���p��R�Q��q)��"�I���'����i�I'QG�y���	2Ѣ�B%��	�3��%L{��P�	ey��'3B�'�BN�7H�:4*�`�@}�֋ĵ ���'�	#�Ms��Q$�?���?�-���w�c#��ե&��`В��(�OR�d?�)�c �&e`�d��r��zS��<�A��]!eF�b-O�铠�?�s�<�D�_��"�$I2$z�I��y���O����O"��	�<Y��i��MxUJ��`5jqH�BfI��SW�B�'�6m)��"���s���#��\d$PA�"�= �������[�44��ڴ���)$ly��"��:R
I�6�D ��B�D�3%ef@Γ��$�O����O��D�O���|�Ug���1�$�P�(̚�'��DE����'"�b�'���T�'|�6=�8� �f��0.�ݺU�>U�������OF�b>9���Ȧ�ϓ���s+6z��!z�'��͓�u��_3�?i��,�Ŀ<!��?	� _
֜yhtゝm�t�	�&�"�?���?����Ą���P�������ş��bL-Y���1bn��M[�7BC�f����m��ē*���#`�<��Ձ��FM }�'}U��(�:��TZ���ISП@ZF�'�������1@
���.��=�L1���'^R�'���'��>��I8����M�*�DY����/#k���I�MӦ �(�?��G(�F�4�!�2�O�K���kr�ɜQx�j�:Ox�n�.�Mc�i'����i'�	�89�L���OPfy� �_�#��0�,�<��в��SE�IZyB�'d��'P��'-�	��2�It$� I4��c���|�剝�?�@��Ɵ���%?��<-v�u��#U�f� �z�Gǳ�t�*O���yӚU$����8	g˟�?i���.	(a�|(1�N�[ `���O�<Y��׌4�`��O�����O'r<<jI5n~@ 1�B�zЎ�D�O>���O��4�Bʓ �&��hxn��k��UNѢТhY��ͫ�y�Kq���Hc�O��$�<y&W�lM�њb��g�n%+���0 �=��4����Ê���j�6����N��7Y�d�d�)�(�05K�����O��D�OV���O���6��Bm�!�+VZ�[$#�Dj,�I�������M;�a��|���`��Ɯ|2i�]��I���ٝF.��r�����'���'�r�D�E8��1OR�D��� h��(7�,9q��s�,K �/�?Y��;�ħ<���?���?��$(H1�-�*4���@��?Q���d�ߦ�ӆ&�۟\��ן�O/�iR��E C0���,ǒLx�b�O���'����?�V��h��\��f͚;�:I"Y�h#�Y
2N�1	h������i�������|�F7N�ip�͠ �d�pQn V�R�'�r�'����Z�,ش]��((�i���a�A�`;$aDN��?��!��&���a}2�|�6}�r&N%��z�j�����b�Ǧ͹ܴt�Ve�ݴ����%O�8�B�'�b�
�����:F��dH��J�l̓��D�O����O����O��Ĺ|���L�&!�<��.�@%̜:B��0����g��	ӟd%?�	
�MϻWȖmR�j�.<y<Mp�'c*4iy�����OO����i����,�Š�'Wm�Mr5��A�d��B�uZ��U��O�˓�?1�zE� KD��P�+���J�D�@���?����?i-O��oZ/H�e�I���<TU��i���?%��g�pr���?Yu^�a�4oK��"<�D�CJ����Ӄ$�T�h�m�>S�����}����)-y��%?���'|���ɼx�x���G�*��Y�1��4�p����|����|��w�O�����<(Y���l�@�3 I��r�e�r�ۀ��O&�Pڦ��?ͻ9 �`J�?#�m���ear���?�� ��6�ӣI&����	Œ41��i��W���rd�W"���Ti��D�O�ʓ�?���?����?q�f^�	P*�De��ʧ�"S�1/OrUmZ�}���	��4�	a�s�L�1N������dZ� ʄ�׮�2><�Iǟ,��<��S�'F.I1��=(����b*$ﺘ����M�Q�(y���T��$*�D�<�@#͏]�H%h��?�\kF��?���?A��?ͧ��$ͦ!��� Ɵ�y��.7��+7"J|ZԑѠb�d� ����r�OP���Oĸl��Z�@�f�,���k����_٦�'z �k���A�O~:��"54=J3Ҿ2��KA���!����?����?����?�����O d�����	��[�f��4	E�'�r�'��7��6� ʓ`⛖�'T�	|bT�&�&Td�GT�e��<%���Iߟ0�	G�Qn��<��O3�n��]���Y��K����C�����$�d�<!���?a��?q�܋&~��s�$ĕD��Y�ֆ��?�����]צm 4ʅ_y�'���T��	v銗G%�Pa��EW4���	؟�IP�)´���!�j��%OһU��a;w�ʘM"��*��M�3^��ӶP��D5�D	�3�b��gk��Lx\Xumݒa��d�O����Or��ɦ<ك�i@H9�c��?~���3%
�d�Ph���<���'5�6M8������OF�6�]�iIgGٟ2�ȵ�j�O����x7 7�.?�;j�mY�O��I�4L�'K
������f�4�IDyB�'���'.��'��_>���-�x���-���!�&�Mst ]��?9���?y����g���ȅEF���@߬J<0��DK��NXl��M��x�O��T�OH*D���i���3@�&�`�
�q&0̠v#�=���Rk���"��h7��O�ʓ�?�������Ċ�D��M0p+K�^0V����?���?1-O��m�z�$�'?��	�3=^ݘ���,� H����|W�O"d�'}\7ME����H<y�iQI�pX񥆞2C���1�^V~�K�e��*�g��fe�O���ɽf."���F�R|��B�:Qώ s�C�jB�'�'���̟0�	���N�
w�T0��b���8�ٴ^vl��*O��n�a�Ӽ����a3h|��Δ)q>��I�A��<���Jfc�6M(?�CX�Q����5E�%q%-�,� '!
.�֬N>/O��d�O.���O����OBAZq��>`W�Y���a�<�PG�<�f�i�M���'�b�'���y�*E4����3+�$�؛���l�^ꓙ?9��������3�e۔k�>ЃE
%�S��0i�	Q�l4�'Ťy%�`�'��$�g)O69]zH)��ߵ!���q`�'���'����X��p޴2V<p��b���a���o�:Y��
֐=0�tw����P\}��'��ɟI��P�`���{=�e �&�O��!8�D����'6<��W'��?Mk%����w�x��f�A��������ٝ'w��'nB�'��'�񟈅�6Х`h�u�ʶna�a��O�$�O�������I�OTmmZX�	Y�� ��CN�<m�x���M�]uP)�M<���e��I�.
7�<?a"+��1]�c�\�:��!���Q�l͢ ��O�%�K>�(O����Ot���O��r���=J�@"Bf0�a���O��d�<���i�^�q��'�2�'��f�ɩqo�00� TJu#čvI*�Vf���x�?�O���"�1'nh�d�P�
Ӷ�s�KAo��t�a�Ʒ~�i>U2��'��$���p�X:*��(BI�g�t�v�������ߟ@�	��b>%�'�N6�W�νa6ğ"*���3���5�n0�h�O�������?�_�\��R�@���s�M�ƣ�')�	�'�11�i��	�/
P�!g�O9�\�'��)3&�9(̡��ɜ#��]	�'f������Ɵ��Ip�Iz��$B�8��V	A�!�&$�ɜ9cyB6�@�b�"���O&��)���O�oz޹h�jŤd)���a�")�4@����L�IL�)��g���m�<� ����(Ÿ]:�=�W��ih�e �0OT������~r�|B]����ӟ�bIآy��ؕ�̚Y���������ڟt��My�hx���Qf&�O`��O�X��!I IeP���1\:X��(����$�O�D�q�	�Y@���h՝N���ӹOz$�:+������M3����jOJ?��(�ڴ�[*#L�8BJ!L`�;��?��?����h�����m�:!Z�)
�@c㜂�����H���ܟ���$�Mc��w�m��K�5k��RIH��ܡ��'��'��6M�	�(7-)?�4$�L���S�(~@P�B<�l���H�Ě�'���'�B�'���'���'���2ֶ>FтF��=%@h$-�myR|�(�X�@�On�$�Ox�?�c�[,||�c@��.�B��	�!���[ݦ)��44a���Om�5�Vز����H������G2��7��q��I_i��'���'�d�'�>uҦ`�m�*ׅɢ5i�����'_��'DR��Q���۴$��Q���`�#GL�s�`E[2�n���t�����\}��'}�	�	&\� �&�.txb�u��'F���Ц��'��jf(��?�	%����w���*���/ 6
��I4EsD���'���'���'��'{�� �^�IB&c�"abI���<	��JJ��л����I&�di���x����B*WX�(QӅ#�Iڟ(�'6�͉g�i��	�VX>�!$�h7�Q�D�Y���\�!��tӊ�O���?���?	�nj2�h6N�G��ĉ�O�^�ԃ��?	.O�o�~HXH�'Z�[>�)!�؝|Q���E�G
]L԰'�;?-����O���'7 Z}���4�x��栕N4`�ybӇ�8}/G��4�T��-��O���=Fu���"����8���O��$�OB�D�O1�����עD�E�G0]fD�ZD́�3���C��'rR�dӆ㟨�Of�$��u�����ִc��I0�ø|��������#S�u�'��i��
�p�*O������m>xi7��xz�!�3O���?1��?1��?�����	�SXEh�*�-S��e���%5��oڒi�P��	����	}�S��r���+�|D����*�[�^f ڿ�?���>����O+�h��ik��"H�Bq*��B9��.иT��D�*6�U��'��'��I�`�	��zi�r�	�9~J��s-ٛ*nu�	ߟd����ĕ'M�6-��$ʓ�?�Td�/Pذ���AH ��0��'���?��I!�'Ԝ`��`�!头aP E _�l=��O�II����!�7�g�S�\F���Oj-#�ǐ)�V��5��ҽq�j�O(���O����ON�}��	�^�bP� �pEH���Q`���U�D�	7"�'}�7�'�iޅY&L	}V���b� �0h��4-z���Ty��¬t�V��ㅘ;A��T&�
���R 4x�޹
�DS�h�^�%���'b��'���'�2�'�@B� �R�a�R:���cTP��A�4&��q/O��*�v�xm��K41���g�Q)�Q�O"�D�O�O1�Te�JJ��l]����,H.�t�
�fAx6m�y¥�T�8������d�z��[5V#8V�
�h�� ?����O(�d�O~�4�&�%��v� ��ČJ*�h#� H�Yd��'����n�⟌��Or���O�3d,���k�D P��W
��Y�`�V�]�)��L�?�&?a��
N��Af%�C�b�C�CU .����ݟ<�I��@�I��I_��!}���У.7��
p��;>t<�8��?��盆�6��T�'2b6&�۬|�昋���� u����*!���O ���O�i��;,7-$?��K�h`YpfҮc, �%��:�� �G*G��~��|�S�`�����	ȟ�O����o�)Gz�t�F�����	By�|�T���m�O�d�O�˧C5��$Թb)�D�t���%��d�'�^���v�f�&A'��')}�c��H8D�~����^.w+�в�'Y�k�~��J���4������_��Or���iU2c����B��;�T�I���O���O����O1�����&�H� �L�(J���V܄V�6���'���m�&��C�O�ilڴc��4ײ��t3Ǧ,k��:5�x��oZ�XAnyl�P~�(ܭ
��h�S-k��g� Aʀ�]E�I磘�|��HyR�'o�'?B�'XR>�)5k�/�U+���yw:�
�E���M�'@�����OΒ�t������]�"���O��De*�3�d��t[ٴ{��b1��I�=
"�6Ms�Ի&�X��Np��)ܚ�s��[�<	�#�	 �.�Y������O���^�+���Q�û0�lqbN@�X�H���O��$�O��r�F�z�'�b�[8���Z,Dz�[�ep�Oft�'
R�iF~Ox�Q��+�F��vhM�w'�lr𕟜8���;�ZHش`�}�Ӽ��`Y�D8fo��h?�(�&Щ=�*����ß��ş����E�$�'����e���㪊3Lv���'M�6�ocX���O�!o�Q�Ӽ;G�اuHl�o��[9:��`$�i?����M���i�$<�$�i�I���(��O�>��R��|��:e�����!C�J�	ny��'���'���'��"^T�t�A��)HxI��5��I�M#�'��?���?�J~�74�zeOʷH��`��
�3�S�D�	ß��H<�|�4K�`�? i�5�#(䘺VN�C^P��L~�N��'r��Ru?�K>�(Oj�kGC��4�<�Ս�%]P���D�O����O����O�I�<�c�O�����O+�!dfߑ>���Ά�y|����s`���Y}2�'�Ie��S Č�Bt�La���f�z,����FW"6<?��LB0���J���߅2'Bͅ����gω�h��K��r�X��⟬�	����	ȟ����ޗQ�&��/`�@�N�?��?闲ij�T��O���~��O|��v�� �>e����#_EZ����i�Iɟ4�i>�	������'<NQ�& ]���%£K�r8#�P�G����䓍�D�O����O��D��V��4Q���b	8��^�[y��d�O�˓b=���� F!B�'�R_>)
���z��&!��x��##?)V]����4u`��#�?�bb�h�U2�΍t$��A��/����;C���������g�|��
�n�l`�.W�Z�1#%JIj��'�b�'����T�89۴x%��6d˻p撔��힣=uPhH��H=�?��(ݛ����v}�Jo�TD�����j�4}珌�`&�<xX��7���%+�B�Ǧ��'"�=�D��?3�Q��X���2Y�}k���&�\��c	t�<�'�r�'
��'�"�'��_��dS�"�<8Q�9�Q�&?�,qܴ��@����?������<����y�B_� *hm��@
�*���i9���'FO1��XK��|�T牬V�(l��U Z���<?�I�q�Xm��Ov�O0��?q��fh^DS3�ڋq깠�H�m�L����?���?y.O�n��L�^0���L�I�S��ȹÀ�{P�`#G޳*���?5U����~��*ܬP�Ӛ�! �ǒ-X�4��'(pC�d�ǩ}���4$�ϟh�c�'���¥�¼q�Yڂ�W��Ȅ�'��'.��'��>��I��6E�1��_z�D�pD�K��(���M��bő�?����4�5�jX�0�RH�E�D�[���14O�$�<9n��M��OJT�+[��µ��5{��dyt��h�Ƙa�/19x�O�ʓ�?����?���?	�D����bQ7w���j�F\�rڈ�0.O�9nZ�� ��	�D��{�S�̡#L�95'�q���.؜Hc���$�O`6��Z�)��� +��(P�_%�P҂Fc3@u-� �n�,�̸0��O
D�O>�(O�=k�W&2��G��l��,�O��B6M�O��4�.˓5l���`��8!��R�Ό1@��ipA�,ZnҨp��㟈�O����O��$ۛ%<�0F��z|lYq�NM������&l�@�4����&�?�'?i�ݲCY�����\�@L� cEJ �X���	ȟ������I��|��I�'C����mû]�P(�'�f�����?��NL���2��	��M�L>�CjNwB89����{�ph+6��L��?)(O]b��z�4�?��T���=Ĵ����J�;g\-j
��=�䓬�d�O ���O���%Pl  G\9�Ԉ�"��-X�$�O��Tz�F�A�6=�'{�Y>!2�$�(B<�g��?y���#?e_���	R�S��^P�I��+@<a'2x䪊�s��H��� $g>г�V��9�ϊI�I�(�d��c�~{�x�#�?�����I��4�)�yy�(lӬySWh��	���d������N�]�����O� m�`�F�����0+�6���F��=��X��ay�#[�����h�Q�@���O8�̕'"PA:�#���4��ǗX�X��'=�	蟨�I���������t��N=kd�d"5�*bȅpůE]�6��[�����O��d'���O&�lz�Q��#Δe�I.]�/NJ��!��M���i��O1�l5XC�d�z�	5��] �SO��@hN�'h��ɴ
<��'�4�$��'<�'�,���'qo|���![
�KE�'?r�'"W�8Hٴi�vI���?i��3IB䱗镡}Dn�	�G�(� �2��>����?K>	�
�@ ���h	O�`��{~Z�Jp1gE�Mۓ����J?�`΀i�֪N .*tAD���
���9���?����?����h������|Y�-B@�X�V}��×1`��D��W���x���Mۏ�wX�2R���\�w��L�؟'��'��.w��&��֝ �N���9� {��A�;	^x�OI�.�#J>1/O����O~���On���O~��P�9��ʤ��V8�.�<q�igp0���'v�'y�OwRl͕�P �!��-:�$� ?W����?�����S�'~����$	<7��+�T,���+�M�S�P�Ed��&��$/��<�'D�0����OU�a��q��Β�?A��?����?ͧ��ĝ̦M�pA�ٟ  � 85k��BǷ	m���B�'��6-=�	;����O��dA�ݰ$�ؐBI��ڧ�0U�pc�O=N��o�|~�i�>.*����䧙���Iwּ)ؖN�/0��(��\�<y��?��?���?ُ��i�2�z9h1��/N�>��N�e�2�'�2�uӐ�򠬳<᷶i��'���Z6G�%Z6�#G�BK�Zu��*��O��4�<x1�Dz���XU�-c#j�+FD�{�b�� ���H� Y�8�,��a�I]yr�'��'6�F�����S�M�+z*`ؐ��=%H��'��	�M�1"������O��'�X�Gg�
 �-��c��2A��'eL��?���|u���� �]���A'dZģK% x\���$إ� 1�q�PU�����IY?�J>Q"��?42�@!)֭m���"R<�#�i�������M#��3hH� dP�pTx��O�(oZ|����� �aD�^��|����.jP 8��П�I2wH�lo~Zwު@��џ��]���Kb�\�9�*D��D�D$>�̓��$.|O�i��-H��b"�F�$
���a�֦1�3�C���I��R���y���=5ꬑ3!��7�&9�N�]R�'�O1��i��Mm�<�I2��|��튜3,����W`G�I�j���!��O��O�ʓ���W~�3P��m���N�2ax�h{�Pm`���O����ORI"!�Z?�h�6�
�f��#�5����$�O���Js�ɜm@��;5���f0@����<,�A=f͈#����M봓��&l?�����yA A"aB�CT�¡x'R��ȓ�T�[sDJ)7>��36I7�A��.w�f�Q {���'N27M+�iޑ����� *�)4oZ�dx�xp�k���	��H�I̤nX~Zw�DPݟ�����=%uNdcV�PD�� �D�<	��$	u�H��N�e�8�$��3R���
�M�4�ר�?A��?���EB� ��DXq�����j�����ONal���M�b�x���&H'2�Je���U�d̢�y�گ*��d�P�'7��I�k%��0J��o�,`�ƨׯ	��˅$G����O�F�l���V�]ᠱ���8 r� ULͣSF�8Տ�6� <�¤�j�<���[�i�pQ���&"X�A�J �N�ْ���(����������/T*f4�L[�'��� '�N.�@���[
dF�K&,�z�Ԕ�طV2��rWeɹY���g�����dI*}I��{�+��q���ѓ	ӡzZhT3�cģm�*�y��7�mJ�_�CxdP��l�f�pX�w�c��EZ���#��I4v,��Z%͊&b���0�N�TF����#G+�9�4l���%K�.Jj�1�&j@�u����xr�'��'��<H��iL�f�Ū|5��'͂�g�8�'
��' �Y��p���ħ�pa��q���'I�J%� ;Ѹi��|bR�����/�	�C󠄪���K���R'A*!/�6�O�D�<��͡S�Ow��OӠ����[�
��%b{��D�3��<9�f�`������J
	�C�̬MR�@���>\��FY�����ǥ�Ms�X?��	�?}��O,����X��`��c��PA�{Ӣ�{��QEx��t��!E\��wF��Gz͊��ֳ�M�r���r��'���'���">���O�qf%G���C���U�`D�4�
�	r�9�S�OH� J<@P�)����fu`Cf��V(d7M�O����O|�2�
\l��?�'���Q�&k���k���.x�ӌ}�(���'���'��G8r���B�G�]6�Yj��TmH6��O��˟�I����� ��5v�JuE��S���{�������^ 3*1O����O����<	��N/]�$�A�(�/�� �sZ𒳞xb�'f"�|rV�$�./N�H���Ⱦ>�NaxS�*�b���	ş��	^y��tʮ�S�wך%�5)^܌���'5L��?������W�>��������
 �x�$����	H����?)���?�,O�1�Gd�Ӭn_�ٱQ�%Uniӳķ��ՠ�4�?�M>�)O,Q���d��8]dԠv*�5j�����/ko�F�'��V��%�B&��'�?���(]�ݚ�o�"�����*.pj�x�W��x��0�S��r��)ƋrRL�X�J�n�Sy�$��>6��o���'��D�#?Y��@^'vPy�.Z3�����Ŧ�EB8(5�'}=:�wɩHСm�/B��D�Iӟ4�'�4�'L�T��q #X<�U��V$���x�$=��DM9PO�b>��I<�^�R�aV� ���j��Ӆs�((�4�?���?�զ[���|���~r���2H�k��j���x"�U��#<�G��T�'|��'�bd����\ʐ0P�m�V���Á�>#�ʒ���<����m�����d؋'�@dr��
�*�S��x:��$�O�d�O(�d�Ol���w"�$P�)@�h�" Q�m~��O
�D�O��D3�d�O����G�jM`�a��#��-i�NNm�7�v��������Ο`�'����!q>�s�^�!��e��;�b�z�$ʓ�?�H>���?�QlG�~j�����9��Ȧ_��ykC��
����O��D�OT�B����[?��ɥ�H�!w�P*�L�ĮW55�����4�?QL>����?1t�L���'2}p�o�8��򲨎�'�8޴�?���򄙝���O���'�����mR�5z����*�d�9R��=�fOL���Ob@�ӯ*�	e�!)�	����Ǐ��
�榁�'�)h��p�v���O��$֧5�ϟ�m��<��H<U8���M{��?iw$O���'�q�fȳWA�.�p �7�^�sP�i>H�	�Jw�*�D�O������'�ɱ
􌕒��,"���h�b�V��ݴP�Z�������OQ�I�0)#��"J���ڝ1�nU�$F7��OL���O(i �$h}2Z�T��~?!�"�-��Y�A��-j�+TI�0]��M>����?1�X���q�Yyk�E��!V�� �i8�H=H�든�d�OV�Ok� ��f�Ջmw�`pD��L���PY�P�C�B������̟x�'*N��$-��T�&�
�,��܀4a�aP�O����$�Or�O���O��K�'ڶmx�qh�U����W"j��O��d�O��$�<�[(J�i�7t����Z(d�|)[��0B��V�$�	b�I� ��78�܌�%��AW�:��(��
p�I�'�R�'ER]��IGҤ��)�O���%���(�9Y�J{����Mצy��t��̟|��*LZ���^�d�x&y=Vܶ`§GE�g��'�Z�� X��)�O���u��e�:��(H"�4z�`9iR/]x�I���I D��l��q�z�"��yVH����3b,�(�O�𦽗'���fӘ�d�OJ�����ԧ5� M�+��m\�e�d�)!ʒ�M��?��ê��'�q�����g؈h�b�U�ݺ�iX�)�a{Ӝ�d�O,���a'����(]Z�b5r$�� �7B�=��4I��@���?�*O(����O��3��+:��8�&G�S@�I��^ߦ�������	��x�K<�'�?��'o����:>�=C�TP }��4�?I/O�,��*�F��'���'�"�8!�|�$��W<
hGᖗ&!�6��O�,PኚA�i>���u��3_W���q�Q.5S'Ů
��5�O��h�i�O,�O����<a�G:�0d�>f�T��Mȃ2���$�����OF�D#��ȟl�ɝ|f '���[��i6�3	�b�3�Ǚ���b���	uyR�'�����ޟv�ca��3�,�jǌ�);� (�4�i6r�'��O����O� d�/b��j3,Ѥ1�q'٦Lx���L ����O��O �:\^ �������pl���l�!�`P�0���B4�7�O��Ojʓ}�"5�����<v��B��(랹�  	%A�7��O��D�<��jU�s݉O��5���斀�S��-L}���gj�+�M�)Ol���On���O��Z��ƶA��OR���J�#�^�!�i��Ib�bB�4��韄������ĵ_���Pi� :���4�Ӎ!��S�4;B�ퟸqH|�K~n��q��
Uܙisj1隽=�6�~���o�̟H��������|:w���.��e��irv��Ņ�<n�������'���L�3?y ��Q~Xuiv���)w>�q�̥W?���'�B�'V�̰�Z���I���c%i[�������!+�	��y��	��pb?)�	a?�2�
aiFy{$����b���ƦM��>U�f�'0�'��'W����A�?9lE��/V�Vn(��"�>i��"NTH�'B�'P�V���ePZ�@`b�d���$��v�1M<���?yL>�+OHAZ���T�蘒s��Q#���$�6}��$+���O˓�?IǄ���Į�0Y|�P`&O٨2�� m���M���?�r�'��?UL�4d<T�w�M¸����O�Z��-�'���'&�^��:4l��'�<�x���p�r��&���J��i/"�|�]��`3�\��`��Z��"H�Q|5�B��� f.}q�i �_� ���%��ԔOIr�'N�\c�v�A�	˪n	�p�pB�4��=�H<����?!BX,MWȜ�<�OV�y��'��&�$�	��Ǌz�x��O.�Of>4���O��D�O@�i�<��x���d冺~{�`y��H6���o����	,
���21�*�)�ӧ?��#A��1�� Y$@6M�!t|el�џ$����h����$�<م@�2��(���|s�Șb:��j�4H�(�Exb�	�O�ȈU��r�L���,�d�F���y�	�����K��خO��?��'[T�s@{����L+}�\٩�4�?!(Ox�rA;O�S����	ɟ�saS+f5�%��Ղ:���3���Mc��@>����P�`�'�^�d�i���f*�*{Y�ݸ�K&$%PKaj�>�+
�<9)O>�d�O��Ĥ<qfŉ�.�$�h�HR�&IreH�� �+Y���'�b[�����|�	�oFX����<a�F�$-=<�f �&!?����?����?�/O8�+'�|Z��^L���t
§s5��1�Ç��'q�^���џ���4f��/��Z�k
�D��Z��4oZ៤��ҟ��	Uy2�"k�R맯?!�*�Άѳ�ʛ\EtP0e�7U��6�'i�����؟t
�&h�0�Ij?!��
�v���-��	�Ŏ�Q��şp�'�r��p�~����?���t���5���Z%���q�Հ*+BU3�V����ΟP���2/��m��'���A>Zެ�B�W&��e,VbA��W��K�����MK���?���d\�֝�1����6*�l|�s#Q�b�7-�OD���'g���OF�$�O��>��^�b{3`F(S�@t� �x������̦Q�	�����?]��O��K�da9�.	0}ML�f!�&�L�Һi�4`�'��'�����:���1" rf<���'t��m�Ɵ���ؘ̟@�����$�<����~���o
�qHM�0%,��Gc[��M;���?���+:��S���'��'.�)��Ar�`�@��W�V���}Ӽ�$Y�"����'��	Ꟁ�'�Zc?: �3"������L�Y꼩�޴�?W�	�<���?����?Y�����8Q�ѨB�Kr����W�
�0a���M}�U����Iy��'���'G�X����W��q�䓿Uh��$��0��'l��'yX�����������"ѡ�k�02�x9T���Mc+OD�D�<i���?��&l�}͓5 � �8���)R���ԎY8 LB�X�i��'�R�'j�	�5�q�����/*> ���[�9Hִ�ǠG���\mZܟ<�'<R�'p�B��y��'w�$8(��k��9u��RG�D�wH���'�^�T�)���	�O������芷 -�F��E�?f�QJG)�x}"�'c��'�X�q�' �'"�i@:f(�,I*{������lo�VW���c�F��Mc���?!���*�X��]��������7�(�r�.6d6��Op��#!��Iyb��S�d�"iJ��½qU������&C��	��M��6�O.���O �)�S}�Y��;��1� ��AAE��(�*^#�M���D�<�����8��ퟬ���0p��Jta��+��Ѡ�M���?���`�4�S���'���O�������Ё�+9S��Z�R���'Q�a��O��O����O6ę���pA��(WJ��4��Ȧ��ɴZ�H)+�OL��?�.ON��ƴq��'Z�l���`w�\?�HP�Q��s�e���	ҟ��	0��Hy�^�h�p���O�aN���N��v�(���f�>1*O~�$�<9���?���^�0x���"$�(ac��2�ENF�<i��?i��?���򄋍c ���'@�h���FN{V��W��#�n�lOyb�'e�Iϟ�����k7!z��paN�ep��NQ8	�����m-��d�O����Oj�m�~-JQ?��I�e� 3�U:��`�H�Z����ش�?q*O��$�OP��Y�T�1��&�� �a'�[?P�����MK��?�/O�����WF�D�'7�OF4l�Ф]���$A	�K���XT��>i���?A��M�,͓����O,�S�h�d8rV�^���R5o�j7�<�Ü�#����'�b�'���>�;U�^(���^�;Ԧ�����
E��n�˟��I�LA��w�	tܧH5n�b�m��"B�W	��8n��򴽨�4�?��?q��kV�	Zy��1m:�U�bo�$4����!�q��6-q��<	����O��X9o�p#L��v�@ڄƐ�(�6m�O����O� �[쓈?	�'ޑy\z�D�Ժ:L�'��b��|r:�yʟ<�$�O8��̣?����"��'kT,��Q�F'BaJ`m�֟��6��;�ē�?i������1
ٖ)r�����C.�\����Q}B�D�uV�4����@�	XyK� a6����`�0�;G��1�N\�3�$�O���?��O��E�p�,Dz񂕟WWШCg�9���OP��?���?I-O�th��|�H� g���)N��>A0@SK}��'�|��'R�ܫ1��$M�_[�SL�	=#�A���Z� +��۟���̟ �' 1!	$���>(��9��Σ=ޢ̫&b�%oZ矜%��	矐�n}�P�O0|Z0b��H����N%w@���i52�'~��uM<�I|z����0b��J���iL$e��Y�J}�'�R�'��
�'��'��	�a0h��i��B�)e�Q1�&\�`�Dg͚�M�!P?��	�?M2�Oy�+�.��Ul�n��q��i��'��@ُ�$�|z�'�" �4��+( ��e�V�fc*��4C4�3�i#B�'-b�O��OP���ezNy�SYrҘ�q��2<jN�lZ*���	[�i���?I筍�"�#F{���H���y���4�?����?�Ef� #�'>"�'���vy�R7��FP ��Έx���|���yʟ�d�O~��]U���r-P� ��ɷ�\�_���oZӟ����!���?�����K� H/T��u�Љw `�W�Dz}���p��'FR�'�[� Z�bÒb��� Z&^�'"�dE4�2N<��?M>	���?afT�C�t��M4=~$�h���6��2���d�O����O�˓6YjE+�;����1�0D�0mq��VΈu�2�x��'��'���'u�(B�'>��BF��V��ylK!�4�"�>����?�����$�+�l%>��3-�3gz4-K��U��d�]�M{����?q��;C=ϓ��g�"�#��	�L� ��P��7��O����<�
ͳ<��O�B�O�"k�*�G�,U6Ƃ1|��t�2-=�D�On��%R��1�D�?yS��<���V"+���0�|���0�X���ib�맃?��V��6F>��$��\��uQ��O�q֘듩��O���(��Jd�����x0�3F�iR]�@u���D�O������'��\��epU��=�왑�oK?M�i��4D����?�/O4�?��IW~v�K�GW-d8*F�L�&5�4�?)���?�bᑤ��ICy��'&�$���h�*sÈH��b��[ϒ�mW�R]��)����?��-��}�%H��MX��*����p!y��i��+	�[]:���D�O�ʓ�?��?t�8�0��2xA�T���;���'<����'u"�'Xb�'MBW����L�c�]�5�/�r��#	��"�O�ʓ�?q-O����O��� c���d��W����Ë�3Y�4�A>O����O����On�ĸ<��m�?ym�G�Vy"���\�XgJ����VX��Ǧ�'�R�'lBʃ��y"��c�p�䄜�6����P���
ꓻ?��?9,OL���f�y���'�p�Q��  ��5�v	��V)�	���d�<����?��ag����?��'ᄽy!�K&bL\r��Ql̡�4�?!���D�<p���O���'����E<m5R�J���jB�U#`Ŕ�{����?���?!�E��<i.��d�?� ��$BA$%�Y��ޯc����ճi��ɋ�|pߴ�?����?9��~��i�)Y��S�U�|9�-� ֽ�`�s���d�O\U2C3OB�$�<��d`�7R��1)���QԼ���ȃ��M��bٲ�?���?����J���?+�<����E����b��Ŧ`rM+���c}�+ɤ�O1���dG�FxUAb��u��g�����$nZ��T�	�fP+���|*��?!W��'�	p�H���]�"�f�O��
w��O����OZp �.�j�@Is�F�*��'H�X}�L[['�{y��'7�' ��:&a_ C��u� 
�4w�yS�c*��ˏ��ԟ��ID�'u��B�̉6ղ�3u�ްPi�]����.8ɉ'�B�'`�'�R�'(h��%Ǒ�X��Mp&�ϒ���S�ѕ՘'���'$������$M�| Mډh�*�����d{�_�I�$�P�	�JEf�>�c(JY�n��7��0�dG�1�ꓻ?q��?��O�Asa,�IJm�L��B�P�,�Ƞ5�N�mʟ(&���Iʟ ��*,�	1rl�pb�	hߚ�E���T��7m�OT��;?�C���ħ�?��'>V�е$3��F�"\��	A�xB�'D�H��OD��08R"�
��9�큃�ɬ&R�6m�OR��Q�q��d�O��D�OL���<�1Hg8�@ "�3Qx��R�']�.
�lZ� �',�B���4��F�b}���ɁU�~�A�$�M�e&,yq���'f��'q��@.�4�"0����
i��� �eP.q
�І��Ǧ1c��s���<��+\�x$��e�lY'* �v�qT�i�R�'��j�81��IL���'��d�)��H�R�E��dx@���`Ex�/!�������\�Y6��5���A�c�d��i�V "D����*9��:E��;a�y��!:\O�)�Nr2\�6/�|G�d1���`\�2��Β�OȢ5x�Hc�Ǎ.��9��?k�|�C&�3m�@b'D�%�� IŸ
���,V�<�^�p�HY*Z�%���<9�
�j�n�I��� cg_���3SnS�(��0
��]C����}�B��N]L� t�ϸV����k
�?i������?�O�ii���0i���+��G�>i�f�����tC�S&�
t��#?���>,б�19[d�()S�6_Є]J�¦3�0(��ǸuH�kvjU�^^䠣�����?�����4oH�Tഊ�!�A��A�a�1O��d�' ��#�������ݞqP�O��m�o亰����t!�Y3��/9\�	}y�f�;!���?i(�iq�
�Oƨ����"�H�ƃ��h�bi�O���C�D�M�1�,,��h ӟʧ���Go�n �eI!?a\@	*��j*q��!t$i�#+V��H�"� ������!�BeP+uѾ�r>y��蟴��h�O���A���D�ͼ48�@U唤�y"H"@1d��r��	���0<��鉂�$z���k��dC^�.��!جO<���Oȩ@�I�@2���Or���O���R����O�1G�Kv*�"v_�Y+�(�4'����)S�@���5�3��ԼF���ꖍ	�*��A+uB�Uj��X�D��I�^��#$��|R�ޕD�н�晥m��aAOO,�r��,�0��O��:�1��5/[�g5|��'6		xB�	U;��i�����$@�C�u@�PƑ������H��� ���A ;IBMṡf����O��$�OL��;�?����4���u���4�i��)�(Хdڲ 4j|E0K�l؞̣�j�$�x�
V&Nr� AGn�}�(��ϖG���'��t�8���@.p�.� ��X&F+:�⅃�g�}kG�'���IF��C���{�"�(<�,I�K�J���xH�U��"|d��X��*x�N��<�E]���'�|)`�z�����O�-�򈅹��-�7B�g��]����Ox���#2��O��S(+²�3���]��`����xb���P�x�%��' *�k��;:4|J�ʰ|��e�����	�ē+T�D%��9�A�D皲1�ȓE��ULU9.\�}�b�R����:=�&��s��5PjS!BH�xo�$[��'9���6O}����O<�'lo���G�6ɣ���Z^��X'̘'S.	���?!� �A�P�B���u��I˳K����|ҡHװ�e+��D��|4RW��l�DՒ4rAiUhzO�Y��-������k��/mB	��`����F��I1�~r�'��>a��4�J�J���i�4�)%'B�	+QXB�������&h��Q������[�'#�U��� `X�|I�@<[�"�'���'v>�;�Ú�)����R0?h"�+�'�8����³
Ӹ,㐪2/���'q\}(����V�1`$[,e����'��)��ϲ��5�皻�F(���� ���9P���� IDx�U"O�!�cC�IRteN�Z b5:�"O���(�*������2BJ�Ѵ"O��A��P�%��m���R:N�#"Ov\[�f�!P~�ia�/_*1D��"OB�1�Az��r�	}!XŢ�'�jlJ��\k��9@��%���
�'o�C3o_.SH9��h6QӠy�
�'|V��t�ש��4��`J
F��PC	�'�@U6�+{�ԀIa��6���I�'�D�G	�+��j��&�y��'��E���h9jl	u$�H�� H�'T4�Woϩj���".��L3�t�
�'�["j�)�`��@��ع	�'&U�cb�i��DȐ��]�	�'h���7h¯]��Z�gN�t�\��'zd�HCi��r��:74���'���7%��X;�u(@hͧ$��a��'�X��i���TmI�(ݐQ��
�'k�A��(��h����BLQ=M&���'��X�	V�kQv��MѼ+G�m��'?	ɶ�\%��)� G�� 08��'� ���E�:O�*0���OW�ѳ�'IpXb̗<F_��Q��J�J#|�:�'��1'�)^M��J�g��G��̸�'��i�_�=-�X���݀'���'�V���>r4�� �׀\��'��ؐI�~���B��/#�'�@��6ǖ�ĸ�P�G�#¬���'d���t�ă%�8�y�/�G�R�c�'^<��E'��c���FDX(�'V2���؀�xJ�#O�A=l1��%��hɚ-x�,���0>�2�+d��p��6�Za��n���a��Q��H��Nv���t�@�Cyd)��#��
�D�3�!���0j�a��+��Q������%�1O���@��'�-���!�0'��
Da�qJ��5!�C�I�1t�3E�޸1`u��.�"��[Ç:WL��z3THG��OF}��'�"b�K�GD�$%��e"O:\B�Lh{��my��D-�hŬ�'0��\�A	ڔcha|���D�f��"�\4���&�0=qE	Oe&
e�d	��<��"K�K�����R�S�\`��YB�<���ܵ<C:k�)8����s�<���C��1��}G���qB�h�FĒF*<�]��yBF�l���Tm�?U|J�*g-։Pl$���ɘ����[��>�kE��H�I�Ic�3*�Q��=G�A�*/-���6��-[����&��ђ2��H�,[1�?O��T����,x�^�2�J0LO�q:�n>R�F9�8O�qڲˑ�&���Pf�:X�"Ol���'N�=J�E�F�'R�<�[��D�%V�,��=u?]9T�(���N_`	�`�g1D��[�J�O��hR�K�Ji>���
����d�,?1�GW���dS�l-������%
b�	�Fש>!��_8;�F1����T�,9��ζs*!��ѕM��6eC�q=�Y�vi�.B䉲"�J���F>�i�f��+��C�� (�B}S ��{f��IE�%"O�u��Kԏ^��S��%Fm�`"OZ� ��	}KN�KPK%2�&P0�"O���'Δ�-�>������`>�xr�"O�p��-�P�'䙌X����ȓ1'
�3��Q<�X�/�c}��ȓIy
����F�q�^.�*(�ȓz�rh����5��phW�}����=9�'�;�j��IM�,�*����c&ց1!�� �e˔e��M�&t³�>F���M@�٦8$�����<i��1-�aA�T��'��A�<V��)K���� 8���i�� %(��r������	
t!Dۛ;��@V`M�U�����ݺ}(�!(���
r�$8Cj-��D�>��<��� y!�D��4Tӄ)݂t��| �k]1S�1O�}�gE3$tm�#ESU�O�-�c�!����*���'�rq;H�I3�������xb�'�AY�0K�>���K���d����pg��E����u�F��� �X�F�3Q� �J�oP=_b�9��Ϳ�N0�ʚDԅ�Ɂbt�u�1mN�]�0I�V$Ѷ���	�J�EZ�\p�����PzZ��u�נ#�Z�8��V��u���,4���  \�HDH|�� �Ha�0�&?�V	�d�����mX�7؄����Oձ��	!�M�oq<=Ap\/mr80)4"O�[4����	��o�9u<��s�!�%S���&C��ox��RE�3�1���PI��RTd�ɒ�C�#�5iЭɃ�,��PRh�*qq���G�$*��s�	����Q�kC�O���rC�j�n=��'���ja�O�Ct�U�^G~���I\�m�&`��'n*�yt��("�lP3�(|� 8և
"g�9�D�!2�z�)q��)����O�ZW�3�p<i�-��!1XI�s�	}�����Zd~�v2�i��͗�(2��1,	�Nq!!��6?��$K*=I �1U�ӳ6&t ۠��(��TӓPy(<Y�
��fo��Z�G�]�]�C��m0�i��%�x��Ӂ��4H��&��I�}�\�O���K�D�p����ȑ
�(�Nv���
�K
�ʸkWK.$hQC�E�$:LPBC��R� �sBf�t�	-i.Z����a�T�k,�N���/��w+R�,�`�b�Ƥl#�yD{�I�+6rF܉$S�IX<ٻ7%�8�y"��hY}3��(m�~��"'T!����7(�����m�B`%��1��Oȸh%�ܒiC��3a�3�����'B�,�0S�P���2U"�mH�k��)ð�
7i�>wm���ą��U*FR�߶�G���e���[�2�$t��'�������ģ��2x�T��  �Y�r\�4�'�>(���B5MN���'�|��R��.�	h�~�)��P*K
8 wNN��a~"/_���A��ݐFn�a��\8���",7Ph�b6��Z�Pj�jy�̄����nBBq�l�}P�@��ސ��`�0�R�F}�F�7@��e�W�lͦ��"�
�?dI��H��� 	D�<|B�K���@�MJ��C���t?��`A2�;�H\�KJ'��@Ye�Mvzz����29�P������ν ����'�V�iי���ϓB�ԛ���m��q��a��=+�69zԻ�G>r�ԥbAf��ja��W�[�p�a�AL�M�W�Q���,OB�"��>�t��B�cwd�,m��Y�Q��ix�x���ȫ��p���B�N���S �>v���c�)h*頦K|y�� ��B���	@�>��_'�d�2�D�ƩA2Jb�'��ĨW	Y-1��Ѧ1�̓� X�>��)"��|XX@A��2FЖtc����	&%�,�0�'�v�&ƈd �k"-F:�ι�hr���P�fRb�a�+Ev�.֨X�N|��7���4e��F<C��	+1�>s�'��L�DC[{Vh��*�[P]saۤq�4e�1o�M+�f#�+.�Ӝ�4�
7�>�ĢLK�����G@I��GH<���\1*�������N�����H�XR��V���YPZ�� ���:䀈a)5O�Ţ���RjP���n�:p{l���'���P���6;ր�gk�8Ob�Y��U�$x�!gL g��3��5�X��(!�0�S <Z�d5��R3�A�O���2br%fQ���D�fu�O;��)Z���!�"�%ҳ�=o��B�	% ���:G��=�r�ˁa\/^�Q ��X�3
����Oz��v�3?�����f��E��B�*L�p�����F�<�U!�)���d?�B�(��R�2�Jː����&$\Olً�	л��p�%�?����B�'�r9�Ɨ�zHh#c�NM��U�H��l�n���ӨJ���{�'!��TH'L\u���`�1f���'��h0n�6���P@G�O�>qig�"�0t�C�9� ��'t������ {�d��f�<.)z=�A�J�o����A�~?I��An���$֯}��=I"�*���:e
�!�ʱ?v�Wd�K(�a9@��!<��y�kת0�𹀪
��p=	v!ХЖ��ĮB%wj|sQ�^S؞Tj��^�/���i�R�K�uұf݇w�0X(c�Ej�	�'���%�F����Ҁ�Ly����$�R�=�5!:�'[�؀P��N 2 ��#$#?����6ޢT3Ѯ֯j>X�wNOc;�ulZ�*����?E��t�? lt� �A8%|k��/~�}��"Ob�E�Ͼ#qV0Õ��hw$�[�"Ol�`_UX�x'����T�#"OFm)&�l��(��zu��["O.��ѦV����n�o��4��"O����L˵v�1��NP�j�b 3"O����ɸC���0�$����#�*O��)��Ѳ!�.���&Pkw��A
�'��Yk�0D�R�p$�s0n��	�':�k�
{�8���M��sL�@3	�'[�����Q֬%r��ڙp@<���'�����H�.��e���(2���' �-H�(	�Y�|����4V����'�lr�)�*@kRe��l�=:�T=��'4���X�"�@��l�Fi�,��'C6�0�	׻4] ���9���J	�'�L�3o(	s]2�ܩ/�4�	��95�F��>E��GψD�����H6�j1%�cMB��S"���D&��y2&!���Tl��|,r!D�2�Od�S���4H�"��eI	>=u�1��'������<1`n&%4A( �:
��I�E�<�'#u�����?�@�ӂ�j�'%،�#F�O:M�T�&�� ءN��*��Չ�'���#�ۗ~;X��!.ְr�M͞97�]��{���'��E��;|�dy�p��%�����eD�����'�v,r�nV&&4U��'U �ĥJ�'�"�p!��F�'�J�Ĝz}��U��;SF@���x���p>	cF�F ��ɼ j ���� `�uKW�h����ʗ�֐}	�?Ii#�,}��< A�8gt8�'ʓgU`h)�1�]X����21+��)>�.0�E��qO�}��rY������%8��zDJӚQlڳ�c�}���i��{�AϓS4b�0��-6$��'�y�#'�O�P���$J�zh@&	�K8�r�"O4�̯_-
d����#4Ȁ�$"O:�1�c�s�,3�<j@�bv"O�`I/ϭ/�H	w@,��1'"O�Es�\5�z����6�d�"O�!:�Iݡ(��]y#�P�1H�Z�"O�Y�$φ�xm"Y� J@��a8�"O��a��S��3��xLeKV"O�����(��SoGp��6"O4����־ݲ�>�"O��I�I)u��)�V��l�h��u"O��k��U)9h�r�aH&Cl��"O�m�$mJ\�T�K�/����|�"O^ՋE$E~})�@�;��2�"O� Y�j��&Rf� Mǽe�"�s�"O�|��-Xp�b)դL��P!"Ojf�N� Or91iN!q���"O�-r�Ge���f.��|g�E:6"O]�0�7b�dA!f퇣Iv�`�"O�d;ѩ�0`In�إ�h��BG"O��A�b�>��@��@�8b}��"O`(�F� rЬ�f �M1�л�"O>-2�Gǔ�<��D�ӽZ��,��"O�(b�.ݠJ� ��чN�Lx(0`"O���艶3y��kA�Rm)��K�<i$բp6VĈc��B�`c��I�<I�� l0-ӠF&"����'�O~�<���`�\�Pf�%[f� ��z�<�3c�!z �xb�-@�֙��L�<y��B1ǬE2��Oqx�{�g�B�<�AR�fH;c"T� 0!ꐧ�i�<i��Òw� ��C�5L�-"`�k�<� ��C��@��%Z��ϝtt^-��"Ov C偧�؀S��A�Y\AI�"O��Y����K���<YzY��"O���6�Ԍ����Q�X�,)�"O<���e>\�!�0�L.~=��"Ou� ]'S����@�#4��I'"O@��c$��Ts!D@�䀳"O���q�Хd��4�G��-D��"O
���-v �O��q>d�"O��*A�^����`��P���bs"O�[�l�;#����Є�"1*��0"O�� AR�v�|���Iا"O�P��e�h��AC�)�%	
T=9�"O�5�N$BQ��K�Q���1�"O�X8�k�6w���(�-X��Ĕ"v"Op��TK�!zվ�@`���fWz��"OH#�����9C��RTY�!"O�Ȩ�`A@E35OW�h?���"O�	S�% | j'��!F;���"O
�Ҥዓe9��:���7jpi�"O䲶�({F�𑠥F�t �9U"O�=��K�<aJ\[��ϸy@LCE*O�ĮQ� Y�I�τ� ]B��'9ހ���_yf�[6+�5w�F���'G�=��`N9W�0����r�%s�'�,��N
/�TPY�&�8�6�C�'m:Dc�EA!,JI� @Wc:	��'`j�Jf��-2��AC�j���'���
�o�	Diڔ��)_MQQ�
�'\��xV�������nB��	�	�'�L�a˞��H�`��8j&���'�j�eA�,����G֑EG�a�	�'p|	�#k�>1�$x��@FO?��''l3feD-�\i�6jۆ@����'9R@yvk��!�\l)�h�(<ڸ	ӓ��'z���ŉ�)G.ኂ�F�,��'Z����  wp�B݉
Z���'���D6d߲�*2�پo!����'�ʈ���'J$:ԪA&�9n�2x��'�@���B]��0���i��i��'%���΍q� �����d[P�	�'�T%1$�'K��m균��LKt�#�'�d)�싒_�hxIW��*:���3
�'�B�K/W�� ��a�\�,5�	�'̸��el�^�Ul�$r(Ԛ�'�l�g�̢V3B���A@P�bX��'>\�_o�T�և�S��u�'nXP���%{����c��E�����'���ACh;f��Da-7���8�'�z�3��C�`�%�S�ޱ��̩
�'1=sT��cA\9������i	�'}�	Ӓh_�}^�Y����`�'�p����а1��UQ�z
�x�'��J���s
Z��,�+\F����'sR�[����,m@�K�6(��b	�'>�)�afV�}��H�q_�=r�'�I�ßMp�*��4cZ��
�'�~س#(�L��Q�툛3� �'n�re<as��w$N*/���
�'����Ej��B���]%��8
�'zd3�n�p�Vy9u�]/��t�	�'#Ca�=M�p-P� L�We���'�P�cW
�\�H�#V�H�:h�
�'��@#�/�1���5��!v26�;��� d�Rc��r�|�kʟ=P�0��"OMI5��K�)�G�;��L0�"O~�h�oX<4���B����}�"O�1V`\�g�4�c�0a��y�"OZ ����nH	ԈQ���bs"OZX��b@�}����!G8X�6���"O�-90���T��'�Pp"O����&�7#/�B�,@7'Jh:�"O|t3BF�e�Ҙànуn����""O�y@ǁѼ"`�c�,W] ���"O;np^)cq� $����S�H�C�!�d�)E:����G+0�j���$��%w!�$��X�ɰ�"X�\�jT,T�!��q̖d��O�g�
1K��.L�!�D8��anF(���IF�_��!�d�:d���"����,P�)ˑ@�!��0:s��bN�b��|�b�U*p�!�DJ�ɑ�T�.�R�S���@!���HM�ak�G]�[��ؕ��s�!�dǈD�с� \	���c���<!�y�8��,X�d|L���N�%4!��az]K@C�BQ�|�E�
��!��4~��y���1V4���7j��e�!�Ę�Mh��V���ʱAr(�W�!�D�E��щ`.;3P��t�!z�!�U'�>�3�ʗFJux�'��!�̆nL��Q��]�87L�+�� 3!!�D��<��yTቝ08�U���==!���?[�� ����>+����Dх!!!����s�a�,h�!!�n&�%{2,A�v�!2g���!��<s�ibQK��?�~0s��V�!�D�&���Q�OW(=��R��T�!���1.��qA�6Q��1�mS��!�D��V�P�+ub��/�L�I�M�S��F�)��e�����Y�@�w,�?Va���<�O��O1`�%�	�0�`�Ň��.!(�"O���0E�
=B$�J�΃:\�h%
��	u�O�&�B�lL�<�e䃹�� �ȓ���a��WB#@+�1<��ȓ"��B�J8�Kt�P�z���Sd�r*סwf�Q!"�M�V���D�@"`$hdd	P#B�5�ć�xN�Di���u<�[WIZ>{.L�ȓV|����F�#>ĺ��d��I�}���h�2�Z�+�)C����A��H�TS������ 4Hd]�<����q�D�S�_�E���P�K%y��C�ɊV�f�yh����@�$D�B�I�L�&��"�΅PE�E  �C�	�!�l��G�1N��y�1$�0B�I�Qff�F�6}V�JW�E1tRLB�ɤ[�4`BC��oq�Qz�=68B�I�3$������Z1��2�Y%��C�	�-��j�/ӑO^�����$i�C�	(8���A�U�x�FaW�(j�C�	6G5�d�`��k�5j0*��^KZC�I+f��D��:�;��	'k
,M��U�p�˅ϝ�[)��q����ȆȓTt�`�^9M�D�c�˒�+Zԕ�ȓ1��t��H�Wy�rb	+&�ZІȓh�"3�g�6Ɋ�[� �mʸ��� �a@�!�=;gd�!u�Ɓ��P<ʠI m �X�l0�T	I�L��ć�S�? `10�,е�5K��R�wb�i3"O�hʓƄ�Q�Ly ��H�>s^@�0"On\��+׌k�-Y%ą9`p�p7"O ��A�Z=Jh�M�9�P'"O~�#���%}C�l�ūH�-*��U*O�E!��J+δ=�V#Υ=ӺLI	�'(�(�&�
X�Tx��J�,G��!Q�'b:�ʃ�2��	QFQ+熜��'X�0�@Ӡ1[�i再���h�'Qڐb�K��R�� ɵ�6��"
�'�pv�E's��p�hD�^(ڱc	�'��h[E*Y&[l`���+��Tzp�"	�'��j�e}��(����T�8�',�x�fX��aث �0 ��/�y�@����Ġ�����ؕG�
�y�ٌ%��beϼt�R��y�� Z>R]�"�	3��S���y�Jɀc���C3e
�x�PwΞ�y�"N����
ABhц#�*�yb� �v��$�g�$V�2�����y�h"BV�t�Є�V9Y�r��8�y��K�+�|K6jԙV���1�^��y�`תi��=Y��_-!=Z�`᫈��yE
�.=�h�����t��A\��y��ȿ��e+�Z4���+����y�)�[�F�Z��X�$PB�" �5�y�O�[i<-W�15�=jRM��y"�G!<Z^hp���1:��� ���yR��H2�9�JP�9��EbPF ��y�I�h�)�A��3.��Z�nΦ�y�mE~���v��=����^<�y2�PHU����J�;�4�����y�N��Ba�"F�� 8��	A�y�ؙ/'�0ҷ��[�`���ض�y�i�Hrv��3a�J��裕F��y�a%_�����b�.I��������yR�B���� ��j��1�B�yb�\�X1��c$��L��� ���y�ފ+�6�{��NM������y�*��3�E�E���ӂ)ȓ�yR��wljԳ�a�@a���B��#�yBf�a�b} `Q\v�a"ٜ�y���6u޴�C�,ϓw�Z��a����ybl�/G.�
��$�\`�1��yb�.`�`R�F% `!-�e�<	ġ¡h���)�}{� ö"OZD(&Q>c��@�Ąd�d\�"O�-3�F�L&�yb`պ�|{"Ov�@��d=.�E/�:%�8-�"OV5�ԩ���L"�#���b6"O�h@Edх-r�Ū"mE8��1�&"O�l�Q�хF�8��N���
e!�dR���U�����~)(R _�/!�.J{�����Y0jұ��,�Y�!�Z,Z6$홦kE?�f�0�.��~�!�C(B3f� '�ǶB�j�.�!�D�v %��dܫ5-�Ba,^!��E�k��#K�:hq�c�FM�!���BRUs3��P���u/݉�!�d/Q2"���;�]3��E�!�Da�$q��V60�깒�@$f�!�d�>hX�q����0�2=K�.אl�!�d��Kx �Z���N\T�#ݴ
�!�J� ��r�'ZOHp%	0K^�!�� �A�Ǥ�1ex|�t�J�n���W"Oz9�bO�7�J�&�*>��z�"O�M����l�83��.H�<�r"O4̱(�	S���0��\~V\�g"O�LB��e��+���`�,X%"O��IW�Z�Rq>̀�� �����y��_�f�l�BQM�2u����Pi�.�yb�3���Z��ܴs[^(j��P"�y�jD��q  ��k�LL���@"�y���тA�$Ǹy�0����yR"�rA��F>ܐ��vAG��yb�ݡ?�Hm�RQ&x�2� ��y"Hߩn�uJ�EZJ�D�SI4�y�EY�9�(�p��ڛ?O\��@���yB��!L���s�	��;���`萻�y"o
:U����&/'(�#�Ά�y�G~�y��G��.����g�4�ybk�?�e�$��>3���L!�y��ҜV��A�"�م>��X���W;�y�JV�u�6��C10������y�&H�Y|\j�H��<@�Y�d��y"$_�F ���,]�7�q��`�'1���e�`� }(P��lal���',T*C@��v �h�!��'���ӁVt*�T����:V=�C䉐�\��p*�2\~Q�P�#1�C�	�~`�X����^��&�� B�7=�X�hb搘xo*1��o:C�	i�¡���@W*M��x��B�?)H;F�Q��"�v�ޅ��B�	>� �(���< Ő�OZ(Z�rB�	�¼�Ӊ��H��ҴM�B-PB�	&�"�)'H�:���J3��TB�I(x�j̓Q)� ��mq��L�:��C�II�,)�!��%vGL�aŕ=g��C�ɾ/�֩!%���K(�B�K�/�C�I�V� )��ϣ�m�����B��.������&�8�p���JJ�B�ɫoT�y#j:l���bb.�N�B�I�L,\�s�f�Lo�m��Z�pB�7������+5�cAH,ZLB��4oG�0��'�28�,e9��R�hB��A��Q��ʔ/���ـB�L C�ɻ<�.`�WO�H�1BKl��B�	��$$��HA�}xb*�F�L��B��{H4� D��j����D��m�,B�I�i�*гS&�=Gr�p��ҁq��B�I�z���V�u�6���QT�B��1/�x���O�OB���B"C�	]���)�OR�L�q%�_7Pa�B�I�,kd+�D�y���s͘���B�Ʌn<���;�찔�	
w�C�I�>�0�`�Gђ fȰ����5��C�mM�	�s���W\)�d�	 2��C�%{�ЍAqɵ{�XqckFhI8C��?e�	��Ñ=zbr�ͅ�H��C�<0C�E��k^�1�a����C䉚��E�"(����K�F��B�	B�F,z��Q��	F�F�RĐB�	�O#�(����Vrq��O͚B�I�[~l[a TXv� ��I�C�=	��j��9r���`��]m�C�I�z�����	x�Zq�XW�6C�I�b�������8ena��#Wee,C�)� Ήؖ��;q޽2�I�G�2u��"Ov��'GG8?_v��Ҋ53T�ҡ"O���E��1W��ʂG\&~�s�"O ��eG�&���I���#��w"OX��4�٤L�`����,l�"On�)U�]2>���b�S Z%^�8a"Ope��˗00��o۽:�՛1"O�K�EB�j���[%�P!@�p"O[��ȸ%y�%"Dm�C�����"O���s=v�8�+%�vq��"O���S��Ac�P1;�d͸�"O|�i�&"��uS��F�i�b�A�"O�Y{�N�	p��� �' ���1C"O������ �pģwD�^�6�A�"OTI`���d�>% ��B�Z�~�!"O:!"��Q����ԥc�$��"O>p��-��D�@�RwH4"�8|�w"O�D�"Ր�<���Ǔ�xE  ��"O^��e��N�`�[�F��LEXE��"O�� *Y=������"$�:�"O�-kA�˦������"
%����"O�p��+��#���D��V*L�"O�4QcC #,�1P�aF s�Ա�"O�$p�B��F���:FT���t"O4 B����2�C�8���"O���o�q:T���3W�:�"O|��-o�٦�A��`"O`a;�c��C��1TM[�q�KF"OP@�Ԉ��T�~��l�}^@�Ib"O�T�EBK�,6D�kFi�.PJ11"O���6�R��U�nМ���(��k�<�A�7)���o��w���0a�\�<��Huc�q(���4��d&��Y�<���ˤ��v�W1��1��SX�<1��*N"�Za)F+4Xb})EJU�<�#��	"���-H�3V~�hVH�M�<ᡃ�����V�Z�D�H��P�<Q�M�9�:MJ�͗	�:�,�H�<�G��Tlr|8'J�k�R��	i�<��JO�A	qM��<�8رKKl�<��b�Ů���J�<�z=����e�<���J�wt�9�3mһ��l�a�<�� J&�x�(�.
�k���8�iVw�<yE�U�b�r�ƀ�?��l@�Dr�<�զ���a��i��S*�)5�n�<�؜6��HwLV=PO���b�R�<���� d��U�I�rHށ�	g�<Y�&ֱs�J�H��O��yT��a�<aq��,f]x��&�"�mÆ\�<I�!�0���0���l|F+V�Y�<i���:İ�5Á+<�`	�ϔU�<sOO�+��mi��+Z�����J�<����L��l��K��L����[�<�@�QF;%Ѿ~��p�!�X�<�uN�6\4F���M�REz���T�<1A)E$K��={�!ǈ&.�ȓ3��S�<y��fD�4�7.�lR|�&XU�<���$i M��4�j�LQ�<�� Ň}m6D��/�n�����t�<Ѡ�Q=)�0����M�dl1��n�<a#B�
2 �C�Q�&�L��V�`�<�\�Q_����#�P��A�1o�C�<)@�O 0ЉD��m�<}Q�	�B�<���H�P_�@�r���4���c��|�<� ��'E@�j4-J�b4y��"O������	Z�jձC�97!jm	&"O� 3��Si��X�J�.84`�"O&��7ƈ,IP�[�*S�}�5"OıS f�nĪ@��f*T�"O(1�v��m��l�E�
z�{�|�'��2CȐ>�P�.N*"~�	�'er����� ��Kt�خt*p���'��A2e��cP�`$䖍p'}X�'�F$K�AF��Ұz��]A���J>9������O�f�qd	X���r�P�h�� �':�SB'�>_f��ҩA*\�>1��'�2��nP�\��щ� �\j�E�
�'�b1��ʙ�X5 3��LI����'BY����9�8�I�J�=�H�q�'%�A�$@`4|��I�
$�ȓ,.0(��L� ���( 60���'�ў�|Jr)�.HN3�c[9逸kt�[D�<)� �0.�l���q��T�]>FB䉕HWΩ�!�����C2O��Y�B�	�c�ڹꕨFn�:պ���n`B�ə�= �酥U�� � �BB(B��46ҠUȗ�<h
����gP�:7*C䉂w�A�D+�!J�a��0BNVC�	�v�PB�(V�yS��$��(��8��C�N�*�c�-�Ky�,��0D�ܪࠋ�INNy��l�؉SR��O\�O��=��F�vBT������hj����C"Ord�樃M�"�"NES�%�1"Oެ�+��w��}H�L*6��ٓ"O>���D
e��p�Ս�'q\u�"O�a��P�n�4��O 'i� A "O���C����i҄(>�Z}�"ORhj�@K:r?`��ed���B��gP�,%��D{�O:��P`$]�|��+S)ܢ*#�9@�R�'f��5��?c�:�M�~_��	�'l������?���KF�\y5��1	�'y8D��lχ�ҙR�ƞp?��'��t�­�56r�;ThH}�,h�r�)��써Y��HP���*�������y�۬68�vΓw�����.�yR!�c��y�rK͍lѦ1#��Y����?��bdsE�I�zw���snM�r�i��07z��������� �D�P̠�ȓ3rIy,˚#�6�6�0B�$u�ȓc,^ X7���L���3�F��Ҁ��o��E�`�>X�(���I�/(�d�?a���~b��2<dx�#����W�4�$C�<��aظ8��8B��8v&E�1��}�<a�m��e�!��@_>M�Ȉjw�Q�<!��Nn���Y%+�8,\�↢�I�<I4��r��{���/8:���Ҭ�D�<����"I&$]A�� �� �B�<9��[>J $��F��8�1*�z�<A���JSN$zH��q��1yĆ�̔'oɧ��֜SQe��hA������(C4���,+D�H�o̜{`�	u-��2uD�h�-D�cBbɶl�e�Ǡ�+ud,(Jb/?D�0�6��)u����c,%+���*D�@���A#.��q���6� ��o<D��á��.P�|��_��IK��.D��2�II�{�H�RŊ2!�@��ū-���O�������&�<��`	�U57,y�ȓ�����`�t~�kT灱��l��S�? 6T8t��r!~"#Ӡ����%"O�c�y�rd��
�/�j�sf"O������94�лB�նIy�ҁ"O�e�#B�2B��H�"�5s���Y "O��*�l� '���C��+y��8� �'��W�Ї�	�`�,	!�eՐ/J�Z��3t�B�I,|�@��;0�Q��1`�B��,���TW=qs���w`0_�B䉛c����`DB�n�����N&=�B�ɢ3����1[��9%BL�w[�P��[>YP�n͔DY򦋆;%^L@�W#=D���&�ǋTX*\c��_�l.|ؕ�-��4�SܧY��u�e@��t���c�f�M�ȓ}�:᱀F�b� J����v ���#D�	 ��N�����Z�����0����D萊� �@��?��d��LP`�����]R��8s��?�ƍG��
�* A�(ŵd��u�7���JB��"z���s	��$���Vi���'�S�OY���5��>q2a�w�(�n@V"OT�6iN�z�4 ;�nۼ5�Z��"O��9��L�-"�rE��E�8�	�"O��h��|�x����&I�HɸF"O<�`0`?g�Y#BB�I�����"O�c�7|�D�"@	�^	r"O����kH#e������s���Q"OX���M����CA/ ��s�"O\�%��	���"�MK	[DQ��"O�h�O��ES�U	�/9�B�6"O�D(6��2?9����q�.(�b�	ɟ�G�Ԯ��no\�en�cb���ʃ��y�@[Kd&�d��H>шD��yr�b�l�TϋW��H�nСjaDC��4��Ɇh�>.�|a����>;]�B�
yA� S���7�� �C䉳y�L����)h�D���G���C�I�;��$��=R��Ɂ*�t㟸E{J?=���DT|ű0�)-!� SV�*D����H�F��2�֟A���'(D��q�	�IS�]��o���]�fn;��=�S�'Z9�Q�^&x���it�F�`h�E��(|�q��Ȫ��0��P�RF����R��H�ƨP2%J��Ā��"HDt��om��is�#G���h�N.?�����W�^((3k�/#��V!��?��ȓ���Е!�#2�5��cª���8�|�k�/A*l��ˁ�;{�Դ&��E{��t��;#�ry�� P#�\%����䓤0>ه�P�hЩ)2���b��qІGU�<Y�C��0�e��1� S� �N�<)U,�=V~��$.w�n�č�U�<���M,""��*.�i��R�<�d͠%���rL��Ku\�1�LEP�<�g˕�f�p5cӪT��0�����L�<��#�&6&��G(_�Y^.�9��J�<�\<2r��w�5FtDQC�F�G�<Ia�הZ������IO�$�@)�_�<���F�z�D�b��S= g@�p�@U�<���r@�pv� �BZ�<�D��j�`� �E�`���/A�<��C� *1��J�P!4�����C�<����?s���Ff�2��H@ȟ`F{���_ 2b�;U��3�ȍ*S�-	4B䉐|������pT��𔦕�,B�)� L<��b��%*�B�L�%0�z���"O�DJ�,U?��Y�eēu!�X�"O�l��G3Y�B'�S��*E�E"O�:�џ�n�cP%�
�0�2�"O��))=^7@�ga����
1�I]�4�p
�E{�d{$�-)Gv#�(:D�{N�5�Ԟ;X=�Sg8D�LJ��[#w�zmpf�E8>� �k6D�d�+�$%QD�����:��5�g5D�ĉ�c�.2Fe�0�5vZ����1D�`�b�7.t���o]�nӴĒU .D��`#Θ�D h���M)b���-D��v�O�<�Hb�' )'h>�k9D�� ��8c �0��o�:,�v@���#D�$x%�-i^,�fX�,D<�l<D�Pa��NE`�vb�H^{ 9D���D!d B�QFJ�;d6=3d�7D�hP4D��	��t�r�. ȡ�I7D�з��wLB�1�i��8�@5D�T@$�[�x�5u�O� ��� C2D��2"a�a��$����R3�1D�t�6�ݴq'|��u�J�}��@��34�
c-�.$� Eȣ�Q1�t}y��N矴�	џ��II��0�o�
g�Fs�� F��}
#�1D����i��/�����/@�{Ē]50D�Z�m,Z2��V��8@G�Y��.D�x�p.�&v���P�&X��5�#A-D�T8��Lu��,����"@d���,D���)q2��C��#*�P-�U=D��iÞu��H��/�10`nXg�<D��;v�O�1��L� �8*���[f�:D��ʾI�*%�B��=�n���9�	S���Ӗt<c4MI�GY�,����G�$B䉻o\T�bޟL��pf��C�B䉐F4 1 #�Kϐd���(��C��C��=cc���f:��;�ݏS�C䉢U>���@*�D�4�m�vq���<9��?Q���O6����K~�Xa@�|ư!�C"On,*��F�;O(�����L�� ��"O6͋�΍.���(2�j�^�(�"O�0!U�B,n��b��
=La@�"ON5xqaX�D��])��Q�sEp�Rc"O@\�b�\}v83�ɘU�b<�"O
$��C©/�<I�#KR
ݠw�'22�'�ɧ��tDHCl�)����eX�t��n�K�<�q�X:9'�@���Ŗ��� K�C�<F��'�$�P"F�
!8(T��A�<�r�ò8:���$��kHF9J�@�@�<� �f��͸����*�� �c}�<9RE�>SB��1I�+5�A�v�<1S"� I�Z���
�#<�q��eHy��'��OQ>���)H`m���D-#r�`��f6D� *�V�0󰭊s�X�+�F����5ړ�0|
T@Z�@�h�w'�1�����\�'�ɧ��JA���"̐���\�L�ɚ��/D�����B?d�L���+3��� U�1D�D�BF_�~~��9b�1��D��<D��Z��J�pg
�it�����9D�0�O]����X�6��,��&7D��H��J����C��G�<�&�5D��k@�D�R���l�L(�����O��6�Of�)�V1�nI�ƀ�W����"O\}��v]d����>9��Bp"OF #BC /���7��h�TP�"O� p�D��_�z$S�����2"O���WGD�Bb�)h3���(HJ�"O�e�3	B�N��SE�S��J���"O�ȣG!�jE�LX�lʡI�h�"�'Z!�� QD�0wm��fD��K@�J�!�$��p�64��ݼ9���Y�Ȗ)1�!�d�p\	
�@�r����α�!�$��Xn�#V�Y�$���K�����!�D4�P�A��H�t0�ɉ"�!򄀠���YbK�c޶���z�!��R�gb�I�흥?ԶL��D�; !�D�>�qIbg��f�n2�d�O!���24ZL*�OS ?2C@c�W�!�d�w�F] ����=�x�#uo�:r�!���>-tx�㇣M���A:��	A�!�ԓwWPY�"�8�r�Qr�	!�dU�m��� ��99��굉N�W!�DB0s�!y�o&y�ĳ�D�"!�^�8j�v� w_�Ӂ�
n�!�	�6#6� s��+?���f(�b!�d�@����R��(E�<�SUn� ���$2x�<xc�D\8|
P�y��.��C��	&ﾉj���W�8�I #K�<�vB�ɹq0��4腆�$��a�L�XY$B��(H������B	kyHc�j�'z(C䉦,dlՉńް�M�f�0Lv�C�I)f���� 9#�aa�;<��C�I�9�����=o��P�G �Q�BB�	�*�\���J]�)��艤.K�8�B䉐z�:����-!���7c݄rj�C��8AG��q1��0`��1�Ì$~J�C�ɷ��U��,�3t�YK�M��(C�&{j�`3��H�N
z�{��B�ԼC�	�V��ѳ������CG�5'��C�	I��pFa֤A�r��$��|/�C�I�~� �&��o���မ�-^�C��;;uic6a��|@��4�ҙ��C��1�ܕ@��ťKN*��#��	&zB䉦0�!��BY,IR�3T�a�B�99gb�����'~T��D��<�C�	2��d@Ч�?3�����K�#�bB�<\(|(�g\�H�Vmb��ݳ 6C䉽-�lq��A�*y� �a`P�,c�B䉹	���P��P6Y&�0�>>��B�I&��#�O�9 x ����h�B��6�1��L�*�`�[q�ʴBSlB�	"m���V�26VH1���2C�	�"��� 5�M-Tl sիD�C�I
0�N�y�]���5��͏�S��B�ɇE�j��ǧgrf����8��C�I#ڨe0d@�:Pm$�%bX�9s�C�I*w�.t�L���.*h�C�	��,Ӂ�^�=�䕒e�'|��C�I�O$]�[3�"�J'P�z�C�	�
�Cg�D��!��9��B�I�]�t��g��0("u;7%M�,Vx�=�ç\�����h�!�$�bE$���k&D�pI��ߺ.B�Y�fX�R����/D�+�g�h��	�g"U���q�q-.D��J��V��f�pG�d���SW�*D���q�0$߬�`�M6m�8�81�'D�ؓ��=$�����G�?�R�:4�)D���t�ì@� �z�EͰ����`�%D�@2��71�D��^&@���j�n.D�� lH EC��W(0,�a�R5v��Ux�"O^Ԋ�N~:ptj��Įr�$8�"O�P��@�|����PI�E���$"O�	hŊ���cu��2��u*"Ot�I�ܑXd��-�#�v���"O��C�[u�rA+Ƃ0Y"����'���S�B�q�j��i�I�pğ�!��D����$�U�p��CZ�Q�!��<G�N	(�O?Hֽ�$��6�!�X7S�0�[Dn�"?ղ	���b9!�D�;m(x�-Q�r�l���%�!�����1$�a�Ĭ
���jo!�$�4ZA�V�������aZ2qh�}��'R@�����3g$W�b��'��c!���v[�� �$�-H`�s&�wh!�Ę%���C�Eʤz/��B@�sA!��*-���a�!���@f,ԐY9!�d���� ���.x]�����^(!��9\T��UM��FC|�	%��=d$!�é��y����_��E�q��6{ў��?��y�Kl���Ύ,H�V���cܿ�?I	�'=�uC��|�L7�9kZ�3�'>�a��V��� wŀ�e/V���'�F��
Wf��apGئdRXqC5D��a����=hP���L�zP�+$�4D�̛7��"|��-(���&�6�*�h3D����W�Xف����@k��=4��� B�&���0��(B#x����v�<�wIY�.���0����[�:��'#�u�<I��n�%BdBэBԂ+�*
w�<q�,�!Gh���͕W�a�aK�o�<��j^�)L��ӖnҶG��b���`�<@� EJ$��O6+@u��L_v�<qt��m�B\ �d
0J
��s��s�<A��Ԥ��H�!��gzt����Dx�lEx�ӧvj� 5��IP̃D�I��y�)L�h��f�@ Dm�������y�G@
��0Sw�S=Q�DtqV�y2,ٓe�t��`ҚP�`���ǩ�yӒ&���C�azeZ<z�e��y"dU�r��Z"&?�ȡqFeқ�yb�¾l�ȱ���ǺY��]��䓡0>a���\��y*��$&��bw�<�pDÐb��jV Ԛb?�@S�/�v�<��@M10�T���B,~-{`kSL�<)�وK�iQ2+� o0�z�o�<�SMݨhz.��ΐ$"A��`UT�<!� ��i2a#[<j��L����v�<I�"��m[�x�d�7h�p���u�<�cC 
�(���ǴM6Z��K�<����C��A��F� d���d%D��2���+֠�Y㨚+c^d�C�#D�8sF4nH�}��I�%yd��w*4D�����/f�4�f�X�7=p�@bf0D��Тφ�ze2�a�
�m�V$D���v.��!]ȝ�,�	y�e� � D�԰��e�y��Eհ�����$?D�L�$���XH�D��oA:e
�?D�����<o��M�㥌�]u숪D#=D�T�D�D�0��I�l[�X�"=D��C�
�Eo��@�-	{���Hd:D���q�
�JR�AO	l���r�-D����F�K�|�0�aĳ��S��5D�<s�'	6F�N�@AҨ��`.D�� ���C���B��|�(H"O�d�PLŌ2�^I8��&9��"O�`��F��^�*��`� �J<2�"O��Y�N�6)pAr�_ Tn\��`"O� �N݀#�`I�R�B�;o�0c&"Oɘv�	�1���U�s�Q�"O��"�FC>R.@)�5nI�!���`"O�3 @�'p�� �MNF�1��"O�a0�4	T�)���ߒChD:t"O$����ɟ_��TI� �a�p�&"O�H�r���+VHB��=+��U�v"O" �� �#@� �J��<E@��AV"O���%Iػ;"a��]�a�"O
aA�ٚ_P�;a� �p�P��"O�E�B�H�@��ح[�P��"O:���
XE��jX�h�����"OFi(�gC!`P��egىf7ڈ��'ڤP�X<�"�&C� ��s�'Z,8���L�!�����hy��'�.�;a%V$Ј*#�L��	 �'�dr4$S k�`�:R��]Ԕ
�'���C�C�hņy�a�ߕQ����'8(��κ"�&�qP$؅M����'��@�W�Cf� +@��4Tm����'�2ICԬ3	����w��Tɨ��'�������Q��Q�a�N���'�$�Jr�-)�,�ǧE�("ցK�'�pI�a�&V���8��W&ъb�' 1�vN�.2�Q���W� ;*�)��� O�uY�ʈ�;�B�)#�AH>Z7"O�E��@D���^�4ʀbȋ�D�!�$�#�:�� 
�P��;VV!�DN8�b�;�K$ �����π-I!�$J�x��%�TC
�v�@�u�۲N9!򄌉a���v��<stЂ��#!�$�x+&t�@�H�ԩ���^�B�)�.A���X`�8�t�̎����'�V1 ��Q�G�ڀ���y�%�/%�ļ0�=Ĭ�����y��ê"������k��x8�dN1�y�ꚉ>U�x��>���R��Ɯ�y�Α�cd�`
VJĞ�@5�	��yB�#q}��8��_����D�1�y�gZ;7.�\�$d� �~�J��K�y@Os��� /������y�c<N��5J�hGXUIq!ɋ�y���K]( ���Y�a�` H�Z	�y2�C��TdYc�ϥT������3�y��8N�nM��EԾ!c�ϐ�yB�  8��&J);���0w���yHU�I4X�x�ݻb���W�Д�y��ZiF-b�&S�b�8��B,�y�L��/5��Kg+ƨT��@h���yr$�"Z�0�P�f��K0`��GG%�y�DL�R0�M�����>�~��&���<A��%^�u�V�_|l����L!�dշ,��XcM��bo2�@�E;z4!�Ę
��8�LM,f��R�B�!�$H�>�������mM.)��� !�䉕
KJ,8%@�sHZ�s��|�!�䔯jD����+��e:�H(y�!�d��K ��J`F�'����TCV�t��{�\N&� @e��K���e��r<!�dցa�Rpk����{��˃R�W�!�� ����U��rX�u��
��A�T"O�eÖB�DP!枧%��� %"O��Z��v�l�`��;�b�p���y�<�FME?{�X"���/��yA@@�<�L��Y溌�Ɵy������{�<i�S��v��dʗ9^�a�Pw�<iCBCKj�bcL�q��qS�Y�'pR�S��0(A��6��x�_�2��C ��	�Ql<O+ސ�эڽw!�d�4��I�����1h��?z !�$Ü��M�<>1CRk�#�^���"O�Ib�E/S.��f��ߺ�0"O,-xr*^�59L|��$��U���ˑ�|��'A��!�_"oap`	 ��"i�I��D*��HD�T"�J�U���6�f ��"OB�9� JPZ �2�� ko�P�#"O�%�f�<c+ -Г��S�bH�"O��)�cGl�b�
ǇV�^�jZ&"O�8j5,^{*��q �X�z�D"O�V�.:��y��-�
}�4yAP"O�,�AU ���ƍ�(^�[""O���r���P�L�,D*�(�"O����G�x�� ��K*�D��"O����O�$��a�ڎ3:��"O���ݦ���Ӿ�p����{x�`�'�xmа"'&�m��.�|����|�'ݼD�	6T��4*�SŜM��'���G��<آG�Um��ϓ�O���X:M��L�_a��q�"O�`kwn�5ː�����"O������&�p����%�e�v*O�qS㊣agR ��J,���y	��ʻ?`na/��M�� s�\"!�R8VָL8Ӭ��X���F�!���D���TVL�@-�&���	k�O��|ʕ.�0x�N0�BC30D�p	�'�(ҧ@PG &|��o�`����'/��9S���D8C��(摠�'�V=�凒>��H#C (u� ���'���4ƈ�dZba3�mߵr�����'��ԫ�m�d�␂�; 4��,O���/�i>!�<A�LE�2��$bwf�Ig�5�'�Mex��FxR��rAMCCdA; "�S ��yB�ˁK?�d+��	�5�>��FӶ�y��l���f ��%�͹fD��yR����8� ���܌ #�ڜ�y���b�PD��Z@��DE��ybΆ(/BX���cIqŇ�?����?����~�`H�>G�~��h[�O*��IS`�<�w$��z�1���.[hM�Fh�<� K�Cb�bt��*,Ԅ!�0.�d�<�VA��| 0T��>>�HY@�@�`�<��0Pz��j���
��	ze�B䉓+]�h£瑯y2 �B�`O�B��$����Ȏ�S�\���d%O��=�����}@$c�3Y���I5a�N_�t��"OL!U��:
�h��I�L6@q�"O:�`��2S���I����)"OLT����,��I !hюs��Hr"O�D���fnXi�GQ�d�ᩓ"O�1��D&3p�"4`]�Q¡"O�-�B�&{��E  �0{����4��ӟ�G�t\�Yl���i��OZ@��a�?����?��<�c{HɉSuq����f�,�"O� vhqt�A�m��Y��!,Φ���"O�8K�̛�{p���g�5�����"O�ZD�V�L��䚷�ΰ1�
l�"O��)DL��\��#��ڸE �X7�'���'H�CVB��|`�Y	V�Ԑ*�����hO2�=A���
�h�@��=�*��P��yrKz�.嘴ʍ G��e2�I�y��үT��#���t���y"��Z:�$@-Ms*ݚ�bE$�y�ɊL ����3w��U�	�y��:�Љ�pO�ڶ"����-�Of%��55���BB�9An��2X��D{��&�`���¡p?n��Lt_!�Ę$j`���3I !a'�@�,V�*A!�$ѯ|r\���
��1�4�`��!�_����c��+7 ��/a&8Q��'P�� �K��bP���˼j9(��'�`�%3/�t<����7c�MZ�'4�9	� ��d`����.6If!Y�'C~Xc�#�j:֝2�
�;/���
�'��hfIV:Z��P����*���
�'4xm�th������¬�j�	�'�Z���.r^���/M���K	�'g<�K���D����)�nHZ��d<�'nh����h+n}!4�R=.��ȓ{�^U�e�Z
/V������?��u��I�<Q����|�� <Y�4X͂k�<a��/#pH���/DIz�hy�if�<qՠ?}iP<j���~�zey��L�<y�B�n	u�c�,e�h�W��F�<YmNeE%)�4�s��D�'�a�i�P�m�A�*C������y�P-�zH�DW���3��Ż��=)����dɠ ��M` l%{X`pvf�l�BO��1l@����3`I�|Rꬱ�"O�{�	�4AU� ��D�n�"��c"O�XS@�±#[|��p������q"OT$iө��|}��)Dǔ�"�#��ID�O.���Ƭ�)���҅®DG��a
�'˼�B��ܠ_!�D�
9��U�ϓ���<q��F<�<�
% �Ȓ���yJS2#N2�Q ��4�pB���y��Rv@M�e�ē���!�d=��'�(��嚼,�AB	�e���a�'̀IąQ~y��IX;_Pʎ�� �&�'���Vm*�c�6`k4OW�<IO�^��1�QH��DX$�R��SH�<!Ơ��c�D�0eĺcoٲ��o�<A�P9��)k�"��Z|L�W�d�<y3��+�.@�C\8#�5	fKM\�<��ǉ���Ai���B��?�NI�ȓ�#�'jX44k��T̈́�F������+���bā�T�0�ȓE��!;��	+j39($A�����G{�'`��5e�<y>0�4k�NL���'�>!��ے��Y4	C"`��'��!cC�۸w�R��-4_X���'0z��c�U�$�Q6
�..����'�5��ˏ6p�L��d�޹19,9�'
Ґ+�L�D�s�!I��R�b�'{ҍ��kS�Ǌh���F�K��k��-�D:���<k��p ��ap ��@�A�<�0�E#�N��MO/{�a+QEI�<i� ���0k�(O&[�@ED�<� 8�;��1�>T g� �`1�R"O�9z�
Cxu�T!��]����%"O� ��&F�%��3�y ��"O����aM~d�
��Z~r�xID�'"�L�S�Ӧ����F�g��L��<�����������t]C��-��ES7"O���k;)�^,�vbY$RlΝ�"O�)�UًO�>}�s,ڶ/Y|U�w"OBD�vi�Hz�m�v��U�\ZD"Of́ugW�CI\�U�N<H ��"Oީ������Nu��A.͔��W�'��D*;pH"�Z/I�����kΰ.�!򤁋p�����C�7T�vH����%�!�DՙK��%��g�N�����ᐝI�!�DQ�+kO�s������ �
��P��@ld �F!�"�(����<R��ȓ�H�*a�� ��)�􂇺/"捅�t�d(�Ϗ/f|�]�-�HE8���	� �''d5x�j�-
�s� �;d�*	�'>�����w/��j�_~�� �'�@���ݗW �DI�L��TH
�'����O�� f���ONP��	�'D�x�P�[e2��!��E�C�4s�'��A���Y�ʕ"�F�w�
�']:H:�Әl�>�[R�@�Cg�k	�'��ea��h԰qS�A�G+Z�#�'��%�S0q$Q!U���F�Ƅ��'L�ar���8r��H
E� 4rP)�
�'j$)�*A {²��Ď�&�]
�'�j-걭��3��t��,��0	�'$�ux5�J	&��hê��*�����')��r�8(f�!)��&6d�P�'�PD��o�S����D��4�#�'?r8�(D+T�F����*;Ax���'g�х@]&��]�4��'Q�t��J[�nt;�˖/UGLh�	�'�zq��;Y~ʤ"��$�k�'���r�*6�X���ΐ/"���'�~��k�oڦ�z�B�}چ�R�'lX`�U��95z�YCf4���'��쓀55�4��+�p����'<<���-3�J��V8? `�':v��n���� ��47��#�'|��9�(H�0 ��T��7���A�'��p	��!,�1�J�_�6k�'�8QZ��`M���@
EzL���'\x��!��%�,bVM	.8o���'F �9"�.B~.�&���0��
�'}��+�kܡc�hQ@խY�+�-��'��dk"¼5� ��� ���(��'���m�<,W��!�J�Yv<|)�'�d��r�>Z "��Lr` �'Ll�q�	� r$nٹ��N�>'
�X�'���y #�)E�~͠�D�*-���	�'p(<��\�	�N0qͲ@���'��1ЃI^=�P��7bm�E�
�'�H�[Ԡ�Cl	��E�+^�`-��'d���UjӖ%9� XS�,Q(�J�'�����D&d��1�C��6N@:��'뎠���/e�0�p��-z�Ё@�'{t{B�8e�qY�I_o��I��'Et<����'I���
@݇l�FP�'ZN�pDA�D�|Ɋ�;o$���'�8�딅P^B���l��̂�x��� �i���=iЈ1�IB�q ��x�"O@<K�,]�JK��H�G�r�c"O$|��+�C
�+�mP,'e`��"O����@D%Ij����m��^$���"Oh=�$Oӟwؠ%�ǌ�
����"Oн�GI�5i�)T-6��P��"O�%f�4`3J�H�vtC�"OfxS��9%N}X����o\q�"O<�2�
?!�Hբ@�0!�,12"OF(aп_��%�ը�#�=�"O!�âN5-4Щbd��.��	��"O�ժ�m�PK�x�'g�e鸽;"OHE�F�4�Q Ĝ�#΄5Y�"O�,� ��'��1�L[�&M�"O8b�hύeK����{� U#�"O|X���< � 1Ă������"O�@�w,M}2q�עןaR����"O@=��l��h9�%���#��5�2"O����!�6��@�WDz52��UJ�<9@�˕(�<��7��E�H�f��G�<)w�-eW��! c79DM�RIJ�<�Gҝ	��L"�ֈD l��mYD�<���-z*ҍ���O
H��ף�h�<qp�L4R�� ����0r�q���b�<7�e��� ������	J_�<�G-�0r� �A�Rتq�J�W�<ɳ�	]��i[D�R�0�y	vl�T�<�v�Z 48��r����O�<Qq�S�+1�H3@��
a<T`　N�<	r�vd��㳨^A��	 �J�<�
�8aԅ9�]�\�\�Ab�<ـŝ�,�49�g���l�B����b�<!�^"��l�	��s��T�<�i�tfѠ4�\�\˔��K�<�˞�H�x�c ���~������K�<A�⌬A�hJ��[�X)�dϒG�<)���{���3C�N�W4�a��E�<���2Hs>��JD���I�s�A�<��D���r���8>���|�<!猌�,��ʗ.�x���x1�z�<q����E�6���s���:��Gx�<���Z)5u��¦�Ɲd��T���u�<�l\�y|�C�,��(�,��2c�t�<��.Q�j@0C���K�b,B�	��5�Q�جvT�(��DY�~�@B�	�%���R3���y��P�i��B��5_N�t�����=���گw&�B�	ow��Z�)��B�L�F�l�C�I�	� ٤D�%��A�eϺv�pC��ZYH��&B���sgc˷I�2C�ɼ\���O��G�v�P��3W��B䉳,^�4�,��(�r��t��B�	�C��w�#�8) N]x�B�I�&��t��:R���P��% nC�I�J�y�(���䚁L��$}B�I!Q!Ф`��0������̶b)HC䉉.}aPa��?�nL�n��@C�	�}ԂdaBJs�<xB݋�B����x�2�I� �h������T�`B�� h�ұ��iB�lxdC��*0~B�ɭM��X
�[,W4ڡKӷ\�xB�	 ����KA��FS!@B�I	�T*�^0}К	���D:i�B�ɒ.����ā/tpT�
�bݲ[��C�)� &q��J�- ���|����"OT�Ⴧ˞Sx�P s
K�h2}�T"O>XHD�)%Pr%�VD
�Kg����"O`8�j�	ꬄk�˜F=؈��"Of����&W'xm@��]?�M�7"O�AX"� � ��F��� �c�"Ot��LD5MƵ*"�ʇs� ��"O.�1,«GQ��#lϨT��Iв"Od]��'�1q�!3��
�IfpR"OX�P�ȟ�Y@�@i���)��0#"O�%"T����qb,{Ԅ��C"Od('F�-26���K��P`J�"O���I�r�������s����v"OJ��@e�#�� qf��kA�L�E"O�CB푪A��#AL�� )zlsF"O���
B1t���`�g���"Oh�mT�]�h<H�f-���k�"O4踤k�=G
ě�%S�e��XB2"OlPj��7_<i �e�;'���9#"O���F�@㨨a�B
�ZP	�'"O��3&��V�u�!b%6�cp"OX�[�Y�N�^tp����VPf"OH9�`�ѯ3޹
U�=��=��"O��)rLJ"k'��	pG!crސ �"O�*2�%��ą�b�| �"O�@�v/�#�ҙx�-ʙs���C�"O`uI�k"��œ�ϗ7B ��"O^�R���i$�L:�L�se"O�}ـcE�Y��q �U�r���"O���ˋ�] ��I�N�;3P��G"O��է�(X�ys�(> �3"O���^�Q2���	.���"O(i[�ː XX���h)%�5�S"O2ԡ$Ӝ]T8��F��&���"O�<҅Ǿc~�Q"�8E³"O�[�d�����AVD�&"O���d%����#������e�<)��I3(�>�óKıdT���NXi�<Ap#��1�������b��=;q^c�<��R�!�$a%���XN�FK`�<i��g�Tݺ�#F�c��!҆(LX�<q'��Bk(9Z[�+Q99�ԆȓV_fԫ��� <�$S2M7d�� ��~���˔�F<U�2P#�1;����ȓJ�mC��4p�\2�Ț	8�R�ȓ��=⣯X�*I~Ź�"�:g����	�@)e� �Ap!"�� `���ȓ2�|��UaMb�V���l[�L����ȓJh�S���9�>U§��}�I��z����j��ܒi��U��f��ȓq%�yGŜ{�uqF��V����o�b��B���F2�Ya"m��#'b���rx�4JX�y�nM	�M	O�F��L�e�e��U,�R�N��q���pbz�Yq�����x�@㒀}��L��Rb`TÎY�0�:�>��2�"O������9�ƱX0�eڪ�m�'Q��[ҮEC	��8KD�?D�����ة+�Dka��1b��8b 8ʓ x����1Vt�@�))���	 �H�o_!��*n�ٗϵZϾE`0��k��MG{���'G9��Ň63�dr��]7/ƹz�'�*�y�'�*��lr��޹����G{.��$��5
�`G��3K2�� �D}a}��/?� p��E�S)V�����fN:��"O&(�P�>�P�k�1'Y\����Du����]���qʌ:6nB� �$��M�C䉽7��(��@	g��]8cKSa��Ø'������dX?�d,>�h���F�#Lؼe�&�� �!�D
Y��Y	" �+%�p�j g5����O�b��F}�,�	��� '��im`��I��0<���DY�(�X������2"%�!��
=Y0��SQCEI<ؙzab5z�铗hO�O���|<��A��tu�F'A�!�de�N��Ɛ�t�$�7g��c�!��M�k���������f�lo��iӲ쫲"+h�()�Dҡ]���"O~���&��*a�P�'>&�8�'�1OƘɁ�]�5)u���[0V��Y�X�@���-<:�d	Gɕ��D��]������#�S�	^x:�y�ᇺGe� �$$V�D!򤍖50H��œ�"R��y�Lr���hO�I�fC�C�ԥ���3^$�2"Ov�a���Z��p�G��|�� �D4lOn�i�N��XxR��� G#7��ɥ"O�Рu�#J�̭��n@�a��"O �А�S1d|i ��:�z;��'����oQQiN�J/���A��]~��d>}��݋���hY�-NDu��'��y�ۙ+x����9%�I9w*�y�&�'�$�q��K~�x���&R��y�N��y	��)�V
}4
�[s���yr�-n?����(C	d%z��X8��']az��F;!C�h��oG0>�x�XU��Px��i�8h���;`,ZР�\�Ql\�"�'*�l�P��%I&�jS�P��8	�'6���a&Z!BUXKs� YEn��'�VR���+y"U�@k*X���~�
W�B�'��d§�K�GȞ1���	�fضD��o���ڂjp���D+�3u�R�:#�RU��	q���ʠI�< ���G�+�Z���*��(O��Ӥg�x����:^1>i��%T�Ok�B�	�j�"���j�&&@$�z0b��`1ZB�	9m\�ygR�"�愂�&�8 �vC�:HF�x�DY6~V��ǧ�k�DC��530iC�$ܐbf1Qq���`B��	yz:�P ��>%J�z&�F&I�C�ɿD�r07�^ܹ���kFhC�	�,o
�Ӡ`�;2�qA���S9�B�	7\�yY�C� ��A�d�&5h���>��B*Z��]��H޵	����FL�'��O�� �O���̓2K 6�j-Ov��A9	�'Q���3� .���:v�P?l�$����D3�'}z�C%"�P"yH���/VRT�ȓC]���u$�2�N�J(�+K��Ɠ!�X��qOL�~��t�]'w����'�ڤk5$	�p�������	<�$�َ��<O�	�Y�HM�J���Yb����"O|e4���]�a-�:��T���i��'D�z2�F7!�,I�TJ��l�����yb͙*8dstF��T��c
��M��'M$�Т'Q���x���fX�'�ў�}���.���`"K���,�f�j�<!w�M�*j��0��i�d9�%��I��HOb�$���QB�x���y��;q3�O������K����(�4m$�C�	�H ,�U��	X.ɉ5IC�d��=	��VI�O�Bɻ�F�KD$�GC�R���"O� �(*�gB�V���;wg�:=j�@��'���w�ĳw�0�w�� [>�1*2'"D���R�j���1�slI�$a;D���c��M��W��$@:��G'<O�#<�����~��xB�^�I��,�"ϖM�<�GH�}���b`� �,La�G�<)��[$F�Fh���m��@���o�<�@BX �2���<kV���o�<p��*;�� t.�w���P�Fi�<9���3$vnR�8QV�
�8x�ȓ2k��a��3��	����@I��ȓq�.�#��*H��l��h^	�D��'�a~��վ��!iE�G�y~�#'��y��ߟT��tBӠ	-<X1��/D �y�E�9O�]��*�,=�q
X��y2��^-	�%�8�� K�޴�yB�XMry��L$0D4�!r#Ͱ�y���b�ff��x��%q(��y"	�Z	��i��Ƚ>mz-�%�ܶ�y�f> iCa�	����D���y���-zX^i�sM�o�@�)�GZ2�y�oҢ;��F
ݻ!�0������d1�OT�Q�ۘ(�ԙa4�@*�e[$"Om!���[���FIV�2��P�8O"�=E�$���V��s猗I�M
�EE�yRh�WzH0��ƜCl��F�����$�O0���;K�=����[(�XV㏩+U!�ݩ��HacS�3,& ^c�!�DԢv�a2���D���9F�D�A��O�����w/��pg�>M�𠱈�3��x�E�,�TLq�ǼR�<`3F�9|���Y��`#��D�^O`���P������.���|1p��ڎ!��Ȗ/P
o�=[��<4������4:��	�⏞�{Ndh�hi���=�����<�d�d ��؀��b����W*�8�y2�'��K�昹�H��m�)?���	˓m%�7m� ��F�ܢ�h�*>�͚�]���'�~���.�X�BE�ɔN|��'`�M�� ɛ�Oq�X+ ��b�`�B.�0(>�b���'�'1��x:#n �)�L���b��9�6`��|�v~J~&����#C�V�h�Y���2��94�L��Ë�x��l)ҡ��dJJ�Q�����x"�К`�`�ρ2JX2�@�/�����(O�0эbJʑvb�	HE��'��(���ɣ�y�)W�W���2���\z�����'��#=%?q"#���fW���&nY�%������;ʓ����		0�R�a���<R�艂e�Ҙx����'�n�{g�đe�x�"��<�6D%�2�S��?Y�"QS R��!P���ݙqa�<��A6�O2�x��f��QC�[`{�@���Od���O�=�O(���`KD�!0�U��J;8G����'Ԗ�J6��6U�胐�Š{��K�'Z�����+m���Y��J,{��y0�'��8R#h04���J�\ʠ��'O���5�O<Q/T��Ǌ�J��aE"O���A	� ���-�Y�$ b�"O��r�Hfs5�����_��90�"Olv�G�m�:�C�N7��)b�"OH��B\�&i�����/6N�	t"O�M�c'F3;t��o�8z��	*�"O�7͓�G\�] 5,��
��hs"O�qdK)a�m�2l;�����"OL�`,�
]F*�k�!ɐ.�t�"O�Re�(uъq�g	��C��y
�  ����8;x�4�_.�6Y"OB��Ńh�,��cD�G�|1j�"OV��Ё�7YlR���!A>z�"��G"O�=�ե[*�Z��b�X*��P��"O���#c�*ʜ��B�[;y�Q"O���#��* {L!Λ9fɸ�"O�����8W����B1^c��ӳ"O��2��B��'%ӷ+y$���"O6<*&�̀*�p ��'���e"O@��QN��Q�*a���.PM���"O�Db#�bG��۱A�)���"O����Ƒ��d\y���
I���""OJ`�4��y�ĉ`ә$�V��"O�	��D^�ajb3�i�)]����"O�@�У��V%���i�Z���"OΌ�B�_�xT����	?,���#"O����1�n�!2�Ռv'�k�"O a�.�<rw\��A���5"O�Z�	|jxh+$MX��P�"O�}�kH�U�b��&fN�m�&��S"O´+��8�Y��G��M�����"OB�ʂE ֌<��Cqp@@�"OFx2D�X?��cDG/O�����"O䰉���Mb���B�o�f-Ơ�?� ,��F�*K�-���'����Q�q��1�ڈJ��$+�'�*`���ag�=��$д6B���'��Հ�&K�,㌹8w q�HX{�'�F|)u��=w�Z�,��i���2	�'��m���(��swa��5��|��'YV�Ul�!Ԍ��E�<i\(!�'Iv�)��[)�d���+N \����'�����̙b��	ׯbhC�'n �BF�߳.�>�!hE��JI��'Xb�HE�In��9ȅhP O����'��m��c�0[�\i�.Ç��x�'�TH��0�fP��Ȅ�6G�TQ�'��@i�&�*2��3�ı.#��P�'�h�R�&�']?�r��Ɍ$�He��'j��ぜ��
YA`�&%����'��A�L�-F+�y�RaD&�D��	�'�ި*��[9@44��Ԃ�%�u
�'��H5���*i�C�	�,M��'5:Љ׬F=3���D)�7<E�'�L�X�$��=��aB
D� H�'�dܙ�C�}�`mY � ��e"
�'<|:���nb�y����'�4����H*Z�piŊZ�"7b�p�'n��Z��ܸO�<5*��_�/cbų�'�Fl����H���p#�S�"����'|��wm��Hd8u!���!P-A�'�$�C�Ϳ0X�����
�'J�@�덜uc��E��V}��t�x1t�Ϭh�`�S��
k��$�ȓ�LQ�V"�e�.1���Rrߦ	�ȓW�NɸR� `��`ȟVC\Y�ȓu�$���?Q��8���I�P���|Xf�ʐ�ߨ]�D���.S�
ͤЅȓRߠ	aT�K�.rL)���:	/���ȓk�����'O�1Lp�#쁶^�b�ȓqF��e�M&*�T�ӡȋ�@Y��=Q��s�gX#s�TX����?� 	��	�
����O>��5�.3�U§�ίG�ɒ�"O8��ġ�K�8���oH�^=�\Q�d.m��
�'C��,+dM� ���9�
N�d�ԑ��S�? P�afK��2bX���G��P�:}j�g��e�qO8����Y����S�-��	ˇl	���T�!D��P�o�j�(�@��ĩU��� �g���V2�Oj��G�@�59T�
�m�L{��'N ��b�[D~RE;OGbU�A��/:V�Y����yIU6 �&8��cǫ%��I�VƸ'�@��,�c>͈��]ZF�1r�j�j'�-���,D������N�<d�fI�Y~J��e�Ij�O� E��O�l�WeW5-5��9��S�`�p"O�Pq��F$�ږ*��z��d��"OЬ!�
� K����2�ޝ�P�"O��tB�5g�pa��T��q�"O�4M&Ch�AI�B��'TX�K'O�2�֚8���y�o�r��Xe��9,_lC�I�vע���a���	􉊈DZF�?�6��nFxb?a�%�J�6R���m��s1&�R�l0D��)��ω	e�h��'��(x!�<���!�6➢|2�oF7Y�P�rP�ʏL2d���Z�<� ��c#0��&�̰����CV��1������'.��1&�`x؈x�ɚ���p�	��)��a��K)5Nn!(��t�4$��B�-��B�D���NW
5#޵+�n�\{ȣ?1�O�^,�b?�[@C�'��<h5��]^�	De;D�5��m�`'B�1b
J��ba2?�&�D��������c��좀!U
h��ܰ�"O}��L�JLʂ`�"@g��U"O�8�c/C�-��#�)F d?T���xRj �|��=�~��%�/w>;�d��|,�� ��a�<��J1q�:�(�JS�7P�����n�N/OH�Pq�J�M-��2��D�v��D���ط
h=3���#.�y�k6	b5ϓ.�\qG�{���J�/5s���4��C� ���٨%� ���b4�	���5*�P�j� �'YY�'�^�2u���0vc�1y�D����-W�t��5���˓)����)�KV
\��^� �朠#a{biK�z��ɛ9�.�;e�Lb�����L����R'�hP6�K��'�J�٠LR$0��В	رH�j��G1|�ͱ�O41'��b9vy�E�ދf)�艀(Tuz�
��W'_��X�B��XY�Ǯa;t}�-O2 J%�]�Bp�塞%*�X$)���5��5��+�V8��f�B�K�i�	*���"��#Z��V�Ax�&� �*�p�I1�na��'J�,�UfD�j���<�UNG]�	؁F�";?�p�@Qo�:<�|��4^���8��
90��
���H� ���|ݡ35cö��E)@�`qBՉ�=��$�#l[`P�NY��0=f��*�Z��4fW�(ZRL�ơ�|��	UIjb��b�&m~z�&^&(����A�EH���hEfG6G���p�^+m�^��"O�(���O����B��>��<�F�g�๡���,/sZ��� \j�8H6�^�M����'�z��;J�������4z�����/�&�����,��$��"\�'��ss�A$�^�d��jC~�4i(�AF��I�[衃�]o1O��n	��xH�u�]�1����I7�n��E�TIh�+�e���A����Ǿm]���s��Y�8"7��$�y��B����0=��n�p�4�I@�C&��eXgF���� M*� ����po��˅�H������|��띐!�@�i�(Rp�d�����I�'c��dE�fT���JZM���(3D 	Q�$8�P�%�ua��3D����y7���.ͪ�n�x�g'��0?���A�J	FP��ç+� �b&$^���C+�.X��̐*dA&��$�~�l�h&�v� q�ީ=��`��Ԍ�4�BN�%#��+�ןXi{�dG��TZP��|�"���"O|���N��Cei�g�(���OB�P��+H|f!�$!�=�#:�E�[�>$ `�?Uon)�b%G��P���צ]�DbΔ��:�Z��<}�v��4L'�D!�3b���o�k����'�8�9�
S���{������Z�4�LqH>���ڇ6�\�y��;:"�L��3.�tN�UH���3�,�O^A0Ј�z��z�U��(��?O΍��o�(�'��ܛ'��i�ؤO��2�-�P8LqsBK� ��u	�"O~��!���7��p��	����r�����A ] �E�=)�Ȯ���+I���uE�&�S�^h�����µ^�JU2���n�*�ST.	s�H�8U��f!�� R��U�\�-��lrF�����Ɋv�����@f�8Iֳ'�� b��CTdB�	����i�1����A��:J�x�	�I?�I�?E�$��r�6�9�܆�t���D �yB̐�CɢhQ7��`"ޙH�Fƃ�y�
Z�g�z��3�ÏX',<[Aiӈ�y"�۷+��J�$��`~P���@��yM7F�q2�U�6,Q�Ѝ��y�ɇ  �p�%K�.*�x�@�N��y��G�/��4�#��$���ku@
��y�aؒNR(-�P��/�p�)�y�'T�/Dad�މ ����*�y�I�%�Vi07�G&'�f��s���y"�Y L<�|����!\h-h�'���y"�c(���N�W�� Ȁ��y��O8WC�-H6�Ċ>��L�"g��ye�A,�%��&EѸ�K�k���yҎ@�J(�ђ B)76��L��y¨��P&L9 I�%~������0�yri�%\�Y��O�eC��3��A��y2�C�X"HU 7!j��le%S5�~Rꂹ;dT�=E��c	�6��UI����]�88j�W�y+F��Y���m���mÇ���	1r��3AK;<O��bf�� ���"�,��9��%���'��1��	
.e��P��sÚ-Z��
�F!�3Hܓ��x�)�/ac1O݇2�>�Adf��hOxi�Af@	G�T�C�����:e	��e�ԝP��Q��C�yR#Ohn�{�D�|�$���d���?��F�quX��)�(N2!��4�x"�8D-zdRƀЁs<��a��x2���F*X��,B�S���Æ?
��  ��LϛV��Wsƀ0���UX����hJ�����ΌY<�ö?�)��#�"91d�3�[z<����׍�� qo�?N��aZ�i";xC�I�'�E��O�ls<Ô��m�H�>���LR 1c��2Q-I�C����a[�N�6-���u��� �������VZ|ț�"ON�[7V�Q��l�'S�Ui~h��N�u�da)��-6m"%�F${��Ox8y
Uf��y���o���K��]�h@ �j��r�'ͥj����1�¸vOZ�2큃@H������$�o+8D�)H0c�+}�#��6�_t��
��0�0QP�h] J� ER�vt�H�4�Y��#Dל8��!�ӣU7�
�Q�7i00�PA��96DY���'/�qc��w�PY�t�,n�i!(O�Mr�!S�b����'F�����Q81j�f+��/
*�@V�%,XA�s̓T؞Ա�EK#	p�I�A����%���C�"�����|/F	H�� JR$��b+���"OX2��@"k����$FxOv(����lC�(�	�^ ���E��G�O/: ���3Kߎ�k�7D��ူ-Ϲj�)����O2m{$�}�����6�Q�v�ɰ@���Fc��&�.l��d��q��?n5�=*,��o6"�{�B]H4�� ! �L�9�t�4��*f=}ԁp��!M�j=i�I�c�|Ϛ+{�� y�a�JUSHD�����c����T�3�Nt�!�ګz��4Yv(
DI(3�Ć��th�j��i�&J��u����2�z�az� �p���BOZF?�R�!-Ϡ�����wY��qD+�����=H-ry+�H,��2i�a�	#4�pڙw���3�gC�o�����k�h�H�y�ICn�v�QH~�O���b`�LLaOغY���6�O6a	���4����5��l��L�0��FlQ��Ą�V��1���H,�$�PT���\��:�(�iX�vt����c�*��S*�����Q6f���0 (ӗ7M�\B��/:wY�� �6��D��<��43�X##�Z�J�,ë9��\�(�0u҆9br��A�,��ìL�?��{WM�#'�B�*l*;���:v��x�D��L� �� �azb��#i�� �B?�1ˉ
$�A�i͎���:���+�����@�����0�߮}���Q�KI���C�z�Vܩ6:��h���
L� �#px����"xl��g������� R�Q�P��ë��}u�5X��M�L�TA���<����'o^�P�G�+C"��5�	?'�\��0`�M
���W�
�z�K"��&.*��+V��v	��t��Hy��O\�&eЦ'`�[����J?� b­�`VyRR�_�4�|2KS�d� ������+�<���DD�=�6-iV��/�l��B�JN��#[�ty� z!�aׇ&#��)'M���n���`K\�����M�h��(OnX �Y���y��:�t�8$�  �/��%�#�i�3�	�&Ŧ��B`��B��;��L&+��C�I�'��� �X2���u�L;7̌�Yk�}Ar.�$!�b���K�p
X���JB d�E�F�õB��x���+#��<�0(��\:�5-�� 1Go�<q��ܡ�B�{��1����&DQ�<鄤�T���ڷ"�/L��h���J�<�v�D<�
����ܕq2!4,K�<��߸d�lAGʌ�{>�$Q#�A�<1��ve�h��E̠dT��@�<��AX�+F���ӣu��4�y�<����ꘘA��� ���psc�<9w`L<n���r�'A"x����Qv�<��(U,{P� rb�8�@!�h�{�<	�"Z��X�P���}�Hy�#s�<a'�ާJ�D*�E���(��bl�<!s���r����b�WW�Ʃz��o�<	��ZQJ�D��$��u�N�<�0�A�0����3�Ŗ>��8�Sw�<�^=S\q�H�9�B��m�<����xrx��f��2CtXK��P�<i�����Sa�|���"��L�<����%�p�)ڲz@�i�r��H�<١
I�@�3|aҡ-BI�<�WM�;��DHN��t��Q�M�<����� ;�S����H�)��OI�<�㌖
V*T��M�:t�A�!n�M�<��+6\#l�H1ǝ9C�����A P�<y"�^�}�`a�4%���fL
Q�<A��]�(���(E0ܔ��RC�Q�<�%G6A!a$_n�ۗmz�<��ʖ9�C>2#>$�Fm^^�<q7�ѾD����	�?McR8c׉L^�<���Sn��	�%�
H8}bi�}�<!�Gњ7���K���35	P-*dN�g�<	FU�8;"II��ҩT1���[a�<�1�
@�p:��P*M*�a��e�<�ׯN'^$\ɧ�_$e	`�ど�g�<���S�T�F�#���1+$Pc%�K�<	dH�7$ج"��B�?��pwh�@�<i2��za��[�#�^
zUX��e�<�AX�����42ăש�x�<�!B��R�T��LTn8&/Et�<1�̍����%m�-"}蜚��Av�<�'��
'�����.�k�Z�<y���sf"�2`�>P��q/PZ�<�⟫U�i+����]�k�V�<�a�ϣs"9V7$��hW��L�<9�/��6��'_�S5Yro�K�<ym�f�81ɡlǯv�~�`�\F�<�"V6v��t.�ox���h�[�<R���SyA)�d�.vlz5I�LV�<9'�߿Q�vX�P�+a0FcM�<A̟m�L a@%m�j�H5��\�<EA޵*�>1b��M�wU�)`&��]�<G�ФF/H�1�j��f/X�ת�T�<y���cŬ4�cC�i0�8Xf�AL�<!�+��E�l�!�'D�7��C���g�<Ʉ��E�8�&�F`���e�a�<�F"ǆ3N�u@ �K�z%���PI�<�ՕR�@��-�2���5BK�<)�%OL�M���I2������i�<	k�gz��sd�bg(��q@I�<�#ϑ,֠�2��"B�8R��/D�RW+�(4>��� �|1mr�l)D��ڵ!̴v��!��m�+����ZHC�)� &+�ߒk�ڣ�´��R"O�r�m��Q� l�X@A"O���f�@�It8���~C @K#"O��QA�@M�z�I�=x#xe�"O��WA�y}8�5g� O͌!��"O��dޏzv� 8�D�C��r�"O�@�3(d�(����z=ڐ�v"OE �Ԡ��	���36&� "O�}���'v|��e���T��"O� E�,J�+�o��+� Ib�"Oxh� @�j��M�B'6/� ѲP"OxY4_�>���W� <����@"O��07!K�窡C���ڢ�b0"O�5�� ~ɘ����_�$5s�"OZ-G`Σ.���2"v��"O:hC �-	��eHU��)I��"O^��xӴ4� '[Qۆ��1�y�ʑ��>ܩ�d�� �
pc���y���pHm1�T((.����P��y��\�n�L4""GM��Ɇ��y��C �TD��h�9����:�yR���g� D�@�$��4m���y�8 �*PL�.x��1��
�y�^�1�h��
R1{`�r����y�7�Hd�pj�?k�D�ȳ���y�Kر!�fȒalJ06Q���؄�y�.�6n�����Lĩ$pN�
d)٢�y�Ո.��-	� �P3���������Q�e��8wK�qy8 �ȓ@���rM)%UM�gQdT�ȓw|�9�KZ�S�Z��qǓ�f 	�'��xP�#ߜO��Я�++�	�'Y ���1_l��i�+���1	�'4���$��<f$�5E�%��#�'P2x{TۮlD��H�h+��'�varA�V�T�L�ިm0��r�z���@��y�h�t���:)�a�b� �V����o�<	�	:d��K�dUV��s�~�`�s�M�Z����K
ͮ��O^pa��.�U!�ݏC]"q8e�߬ ���W�P�<a*K�/ߤ� �*��:mD����'���Â�Z	A��	&KK���"/�6h!�ON�N�>m&\%��gA"�����@5!�$Y$ ��r����Ti���:g8�Ȱ�9*�N�{���UyZw&������1O��Y%Ѯv՞���.Ȕ``v�'�&|�B�c ��mZ�c���9R+�
|�r2� kZH�IXn,L0 cVkazb��2m���"�&�� @�����'�^-�3#9b��'q����~�����}�i�
<4�y#5�GH�<�w�u�=�E��3y��-{E-�yt�1��2^��52B�m�1��@��OE��15����N��-��k�'OM!���@��w�X����u)��)��(�A�Ž|�����A]yZw�H����١�1O�Q��e�J�DS�4�z}0'�'`JTӑKp��Unڈ&�e�6�5Il�{�E�f����@]�q㞲.Caz�L�?��Pp�;Aj�!1
��OB�2��ٍ}��'I���u��3�H(t�c�R4*�N�PW��s�2D�PI�K$��Q�c̸m
�2j4���QbI.�D���?I���;fqn�	Te���IG��'BjA��v�t@�s��RQ�IҪVSح��OS�x�#���x�2�����=�4�ȓcD&�Ґ�B�G��$��!�C�ćȓ*P2d(��G~\�YJ�ڮr2T��$ �q�b��q Dp�e��8��x���*JuX6l]�D �Ņ�3�ĭ��B	�o��8e���fF��ȓZ� ��@�-rhܒ�O@7:vK0D�(�!%D�����ƈ�^7֥��&D�� X�.\�N�J� a�ېi���h�"O-Cgћ
j��%��:�|<#a"O����ɚ�ؔ�g/�43�j�7"Oڴ�㫀�a��s�A)�޸Au"OFjp��Y�p�gΝ5!��QB"Ot���o@�/�����n[�1R��*O�|���qْ`��.u���'�: �6[��u�weH�ao���'
�P��ϖ��
}���F\��=��'� <k�oFD5�Y��{z
�Z�'��uH& <�����Y�� �'~� �,6xPXl҇��0�ؼ�	�'0���@��YתQQ`l��}\���'L�q;@�`?Ri����7be�B�	�ج	RmZ�tݺ5����7j
B�	�z�%����R����9.Y�C�	b,. �C:9�,!KV�\0L3�B�I�a�X (2�4M� k�)t�B�I�A�x	�`H!y،`��ڏnh�B�#ʸY5%C�A��0jb��(d�B�I C�zx+�
�%32bP;���Wu�B䉟�b�C����۔쑃���Z�DB�	=%Y�$8rbJ�#Lt�A��T�,B�	-]����, s�.�Ȕ̜�y�B�	�d�\�s� �,J\=��CΚ^q����
�mA��퓢G2EUL��d�B)Y�B�I;���R�ˬBX��ue�|�Y����GjJ���<��Yi[,�x!�0E����'��Dx���wF*��a��Ǧ�T���ܶ#�l�ʕ�87;!�d�(3f�樊gΌ�@0��0�ў��F�̓\L�!��i�h���T%G[�lAѤX.i�!�dۀk�MqG�]8�d4(t��/v}��r���c솃C���r���!�$��k����$h~Iiq���6�!��i��
���#�|ҡ��2\��L���]�B��7�ܮ@0L�:&K���<�&��I�h��r�	h��KU�'5r�[T�Т'�Y �
*Y��4C�J+$�H���8F.��`@�$3P��ēb��b�"��Kg�E�	�2H|�'�&�q�%8�(�k2�L���hRb�u�K?��¨�L�*|1A�BC#^YD�6D����'T.U�p��
�y|{�lљ/@�z�c�ze�gG5"���ty�7���!��I�NL�c���	b��Q��<����MT�jAI_�R
��)'��X��jM����8ݴ^*��N�\�q�S�'�V|��,:J�]�gՒ4��M�'Ԓ�L�u�7C�O:�XP�vJ�e�vi�@׹r���`)�P�	�V�0?Y�OX�z�l�c�X�~{��I�,�|yB��g��ő���<�->^=�4a&�^�>d��6)lܻ�%�M�`)���D�a���ĝ,d�:�`.OV\r��i��Hթ�cP+�(���:�f�W��1��� 5S��O���G���Q��D�L�H�T`�".a`�4K�WzqOP����*?�*"}�eaD��"L0mE���8�e�h��ɹ�2�2�	�_��	�F�_�*D8��&��H�1;jI��%�3z"�p걊����g�ND�'����&�{X�8�;+�l�r@���iS*9j`��Q�P#^^T���4�䤆�	�V�DQ��Ag'��A�i�4U�L(H��`�
�QV���\X{����'
�W	�4���O,��zt2�,={SMT	,rQɇ�+��!���'�����	��z����r�R]����r_r��s_7h�M��)M�ap7�V91�UÆ���v�ZU��l��&M@1�y�dܕq�
�	bS��B�,��'��%�/ K�UE��$�s���2vC�A
��qa��Qf���D*�-`70� �^��@��-K���b�� �O$Y�C�M+4�1��(�>���ϓ�g1�5�L�t.$��I�&�Xtê�(9ZRa�SC�h�xp���9r�8��ݩKFܛ�%��>�B�ч�s���䁾\�0��&G�6 # �sM��U �0fh�`"4-��5�j�A�_�K��I&C�.h�`�)qO�iݔ)�`h�W';���g@B 0az��K�iq��cP� ?IBI�&t�HԹ��7.<�%֤"��qj���:^�y{�B"_bU
"�[f��m���\T��9�,@��G��^!����E�](���F�uxu� ��ZL �\\)`� �e��td�E8cE;+�6��E�W�U�Y�'[�M�����f����5%ʡ�wa�0��e�e���P��DkB`\�x�y�ұ�ӹ�:Z�FY1��`�'�O�uCrË�p��`��TєPA�c7%3��Q�
���|
� �`�!AٔuR��>".A��O&�Yq��E��cABR�Ys��+� ��G�	���';Z� �`�E�@f�0#d�|���퉌d����S�0�S%K�#D�(���ޠ @ʜ;W�ʓ
fL@� ��gܓN� X�cJ�:?����&ѿHǶq��N�(L'*�30��su��2�n};V�s�Z0��h���^&e�1,��M����I�z;P�@���#H�d̑���
��cP8
q!�D�8~j�ϽOn�rB�N�-!��B*	Ȉq'�ҝR��r�"h!�!��a��B���:!��] v���@Ĉ�R2�iV�a+!���t�\�9�fF|*�ehӗ[!�$�<v��3��&Z��q���!�����g�;$\�x8�Ȣd�!��b<̉q&'��X0��A�<;c!�$Ɨ}ZNУ���#b��j�OF;-�!���\��Ad�u�nE9�D���!�$^�7ȍ��
W�<�*��w"�ku!�dцW�*pQ��D �>�ڀ"�4kZ!�D�N^�5���q�a��S"[!��e��y�GS(;Rj�Jà�C�!���?��7J~�Р�!�x�!�d �?v�C�Q j>�B��yk!򤑬9DT飢+S*Y��1�A�+A2!��E%4lp���Ɩ�Sg�II1� /!�)���[��M�~TԔʐ'��$�!�$�q�B���I�M�R@��l�18{!�D�T�l$��� �H�	���5Y!�D�W�"PF̅�`�Դ;�ö]!���l!'��]wX����(ji!��[ �H��L%��M��H�/�!��C�E�6� �/աa���#���"("��%�L!b��]�%raz��_�3+���㘋84�Q@#�y�H)�D=��EL/3�ވ��-�1�y"����$<9��й��]xb莽�y��:-K�p�Ƭ�/���"�f|��'W��ҡg�򴑡��fY
�"O���iB$ 3�q���4>���'"O�R��5{��Ăт��z,`lZ �'�^Y��.�)�[����e���@��1F�4�(ɲ�J�=_'�'�*��O����r��h@�Iæ�S����(ݜ�E��OT!��:�0|��GS�sꊄ�D,S�:$I�J��y{�I��N	�ѫc�n�s눀���KtV�����Y]d	+��Y�)���HwE{��T�"�ˬa�4� ��~�����x�w�ƅP1F��A3��ˇ{nX U�Q�`�94��<�`m��+G0�!�!-����B�\�b$��2��rj��<���j���Y��M*h��O�/=��u�ˌ�?9���(����Sk8�T�ӳe�^}[ #ƌj���rk�:z��9S�1`Ȩf��g����g)�?�	u�'B
.��2 ���l��OL=I�p�)�|0�G��c��%���?�'���ⓊM�1X�4:֋��"|y��>��0�%#�?q(O?�gCD�I+4|���Y���8p1�>z7F���b�w�S�?�;[�:���̕9;`"�� ^Պ]�ȓ��!���J�1�S&�4b9n`��Zn�e�tB��z� ��2^O�8�ȓG��\�fB  -H��o!zVх�
�$�2�BE�D#�8)�O��}�d���3^ ����B�9p�jS�
-�L�ȓ����E�C5^d�kw@
*-�ȓ_��Պ����듢Z�SF�݄ȓ]A�a���.DϺ�SGkٖ6��Єȓy�r�xB% ���+��=�u�ȓ1
��ZX���XU�όL�tن�P8�A�;�|�]�� !��6D����QN$D�C�V]_d| �.7D�H�gO��}m!&���X�X�!D�� ڄk N�?н�6$�"),��c�"O�l�T��?]��z�e�T
���"O؍�t�� ~��Mh��Т`zЫ"O<=��#T #042D_�֑[g"O�=��c�ۤq1�iuB�iQ"O�y�'c".�p���&]]8��"O�|�-�,@��Jt��;J\��x"O؀CGk���S�Ŏ9Kԍ�b"O��rd"]T��PD�!.J���"O�щ1eK�5E��I`�� �4IB"O4���
�o�ސ��^�ʘ�"OБ!f��H 0���-0�d)�"OD�#q�в1�낏T�J#�X��"O�ݲ�ߵ&+¸��`B}ڲ"OPeЫ�	;~h��#�X�ɣ"O^4e��1�L0!aÖ<<�;@"OJ�q⍒)؁�Q#�_9D�!"O��X4
Ԏ4p����E�b����"O��+���t.�5���]�R���"O�`'E��&���9�́F�]�4"O��Ї��<�)����2��C"O�Y�!I�f�Ф ���Q�����"O����̃0�����#6K�I�"O�9�T��<7Z$pB �^8�Z"O�t�w��@��� s�ʚs��}ې"OH�2�b[$`�>0ڶhښM��`��"OF����M�o� q��(Hz�$� �"O���.�`̪S�\�Z.���"O�q B��nE����̍��րb�"O������
M4݉�	�?P����"O�� �=I�� s���+(o�D0E"O�	�O*|$b��ݕA����5g^~�<y%&�
O$�KǪ����ↀ_�<Y�!�	[JE���K|::�
��[�<��.?c7h�:U�B:�~��ǚ`�<��;�����/�
Q
����O�X�<Q�GE�U��ݚ#� #R�q��TU�<a%��R+�쁰���( �ٰsh�v�<ye*�rtx��`��:�AV
�M�<��	�"[��J +�/��	A��G�<�db�+$�lH#�0��%����{�<��)#�R��R�4���R��_�<)q!��s �-�Q@�2
���UL�Q�<)�- �P�z2�B>L��b'�O�<��&vPL���܌,% I���N�<AW+;n�P�:u��\Y1aɟq�<E�)�ni`����`X����I�<�pL�@^а�u�g��9�tƎC�<)��Y�pd��`dKҼDQ�f�Tw�<)�nĪ	މ*���(`.Y���i�<��E�(}��y��c>{r.��m�n�<928@<�
B �?��x��Yf�<���ܙD���f(F��lpR���_�<�a.�37q:0+#���㧅�Z�<a�*Ӕ5?��sN��]�<�c	 `#fd�,%���h�U�<IC~�����(*����Q�<9qoW6f����%i�F)HǄ�G�<y��ݣOА� ,У2�nU@��A�<!��U�:�KV@K��GLK�U��C�IL�!�?t����-�4G�C�%t3P��v��./�v�:��޾'�C�	Z"d�b3%̤*\��C�%�4B�I[�b�c�*=D�8C���<�FC�)� 
`S� ,�"�ڧܚ)xɺF"O�$@2�1�rTS��H�b�J%��"O�r�fÃp��<��!;���"OE��#�
5��8Ƈ�n���I�"O|�$��f�^�RS\=ˆ���"O4e�3-f��$r����3"O��`��G�y@��W'�I(8��"O�M�#�ņ+E0�9f&�u�I�"O œ憐R�5#DL���ˆ"OL��&��0+?Hi�̙�e�-�"O���c��o���u�K9���J�"O��S�B�( ����	݇��墓"O�	@��t��@��R��"OT)�@�P�*cB���-��bb�2�"O�A���]+�&4�F�#>�6a`�"OT����A�[�XX�̎_�P�U"Ot]I�D��
2aZ� ��9Lm��"O��`v"]�2����)pKjA� "OrC��w�@�� �\�,!p"O4`YaN�u�ݚdiM�;4���"O4�Hr!��mA��W&0t�s�"O��S���� ��AB�N�9"Oz�J��c~2���X�}QA"O�qa�NF�WRQ(�֍��"O��e�$*��і+ ('B�tW"O:I���Խy����
�
62���"OjYyv��Kh��3�i[�Q��%"O�h��c�4���:$��$3��а�"Ox��@��V�:�cힶNh�l+Q"O�ԛR�٭c���@��
T�X(�"O�dX�L�>o�n�+0N��2�"e"O�ܙ�D���Lz�	���L
�"O��3��T����@A���x4"O��!���V~��k�*�j�~t��"O�x�3D��y��9�u@P�oy��"O��@Ts�<JV@Ǥ(a��"Oȝ�1Ϧ]�ޘhSƹn��I+B"O�ڂ$� u���u.�1�X���"O@��@`J#���9���0����"O4)BI�_�:4K��Y�H��� "OBr�&X2|	&S��  Z�P5"O�mIF��XZ�e)�����"O���G�ůG�&�kĊ��?��"Oԥs�.����9��~���"O�)���Y	)�h�$�˗�|�a"O8�p���,WK���Շ�.����"O^iHf�U�I�n�Q�IB����"O�dy�m�9Pf���i�r���{�"O�``K͗1����f���Ps�"O4 "��3��(Xo@�3��`�q"O�܁q���k�"9"e,2�Dt��"O�-+��(f�A0'C_�@�j3"O�=��)݌/o� y!��'qm�q��"Oz� UC�#�b=�"ß�:@�"O�����$H%d�����x���"Ob�
�A�}��`�Oծ6c�|��"O����)N�m*UB&�؉E7(Hh�"O�x2vh՘h�P��b�>qyr"O�� �ͭ	�TK��1#�P%�C"Oj y�N�! �u�S�H
fD�0t"O�Ԃ�$RN�P&�ع(w&�R"O��h�(/i�,4�g픝_2��"Of�,5F��� /��I�'���y�+�3s��)� �$����q���y
� �Y!�`� 4�t�REӨ3���"O$`Z��E�)��a:@�� F(�[�"Ox��g�-MH�3��H�}���"O@�vo�!]j6�3S���X�+�"ON��4�_�{������ |� ���"O��)*�`{.�r���nକҒ"O�	�J��/�-��H�A�D]a�"O��׃U b��AQ%['{��p�"O�dsGQ-zH���ƅ�+W��H"O�|�u��4i�� �^���j"O���`����;Q圲"( ��"O�a��@�l�D�dԖV9���"O�|@�L��_���X7U~1�9�"O�Ց�	O�4MS�薚^/�� �"Ox�ЅO�z) I#H�*  �"Ov�*씯X�t5�4��Y� P�"O� ����tS$,�%i�.�����"ONa��螮Xj��򠨄�?>�A"Oҹ�p邽��-��&&ո��Q"Oj�S�<)Xd�j_�;�:`u"O�� 2k�'<"� ���X��"OF���߃�$�:a��)(�L�0"Otq���`�6<i�lА"��Še"O(�S&eɯ$`�d�G�@�"O�Ԣ'@ɯV
}ٲ!^q&04r�"O�%��@�?3���i��޲fV�r�"O�1"�j�9 Mx�
�6bx�a"O�I���њ#�	�AC'&Dҹ"�"O6 3�+ҝ+��S$��7=����"O��1Qń�"�=�Ǆ_	*J�E;$"O�0a�L�/Lx�I��ރvB�)�"O�}��	��&`��đ�1X<0Q"O� �wB
%P􀐩X�M�(0�"O0S'�~b����3A6!�"O��u���&�Jd�B���H#�"O��BGGT�%�^5�kS�s��DzE"O��±�� B������&JŨ�@"O<`*ugلw�j�H�� ��"O"�@f*[/J���ĕ�:O�)k!"O�"$a�4��Q�����?v�Z�"O� �0��#4���FI:Z�t` "O�����K�4t�`	qh�T��!�"O�	v-J;.�xT'�2L����`"Oʉ�G�� >Մ �����V��"O�ۂ)1���E�=u��5��"O���+�=vzn�Rd�At�aS"O�b
��rg�4�$$�zS��[w"OX�XC�W�Πr2CW�>Jq�"O,<�V!H&��Z�l�w��"Oҳ	lO�A��߲� �1"ODًC�		Od\�ږiA?ؐ��"O*4�A&H�j�Щ�����uYT"O^�����7����,o�l���"O~h���.#���uCW�:7R\9�"O<� kƭ_��lY��7�x�"Oei��sfl<�Շ�*v8L�`g"O�D����!iev5�"�Ɣ7���"O�<�#A�/���#(	! C"O�L�u��,];CКW$uA"O��9'�B�I�6�����`ׄ2"O�-J0��,����H����"O�Ar   ��   �  T  �  �  �)  45  �@  �K  GW  c  �n  5z  �  ��  S�   �  b�  ��  ��  =�  ��  ��  L�  ��  9�  ��  �  b�  ��  �  V�  � a
 T � � w) �/ �6 �@ �G ?N �T �Z [  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8��H��I*Hă�%�it"L�B��AH<��	öZr��r��H+}J����Q�<ᕆ��8a�%HI�Vݚ�;#`�L�<�ǅG�a��P�����4S�h�O�<a���!=�Z;!)��䤒Wo�L�<I«��>Bp�Ā�L��%��T�<�􅌏i����䇺>؈�i6n�L�<1&0E@�9�7Q숨�����xR�[�wb��j\�g�T����)�yB��,�t��܀R�Lex��8YW!�dߟ}�6��-���H�HU�"OJu`�7��⦌�#7�d�c"OJ)� ��/e�:PYq�f�x0��	JX�x�(G�r�q�Cԧ?�Fp@$5D����*�:(�th
��e`)� Nh<�Bg�Np
Ղ�ݼ�;U��h���?!6�R?D��('��d�S�	�Z�<a5�K7�i U��i��U��n�k���OY�)�Ő`m��#@�YifD�b�'����i�J��8	��ʴL��ط�O�"~ΓT J!��57LTH��Q�ܜ��ȓK�p�0�A�/���qGH
ad̅�CS�`�(6`���C7��=�)���>E(�#Զ(�ͣ)�=(v�݅ȓc�����#O�`r��s@·IB ��e�����C�R5"|�d�G�Wlt��.r��Sk_�I�Q"�(��Ic� �ȓ]�~���D4&�p�q�ϧ� ���GS�-M�F���Ck�'$�r؆�)Rp���"Y�R�n����l v���;&eX�%ڪ}
}@�gd���.�ի�o�.Ŏb�Isb��/>��cu�7��DB� �#'O�x��9�{���;jh,j��å �vԅ�S�? �@�V!��\&����dN��Q�"O@Dځ�B�yn.��6�P<;�~���"O��"��Зw7j��IY�U�Xik��'��Ć�5Y&�#���,~V=*X�7e!�č �<�{���+j)�t*#\Q�P��cZT[ׇ 2f���*Sn��5�|B�I.] �X�2�V-���n�:s�fB�	�-���	/�n�����ٲD|�C�00 .�x�/��U����8l��'Zu V��/�n�zů��dH�rǓI9`��)��?1،,���,P�M�¿��B�	�@���c֍U�!9�E���C-]��pG{J?Q��OE�7���A�'�Z�X�[�*O�0���`��UM�-F�J�"O"��##
MD�yc�xT���"O��D�Z2��	84k?cc"��"OFI6l_!j<��rV�ÞN>VH;r"O-��D�%T@�
�(�:E� �Y"O�d�fh�#W.�)�V���
5��(�y�)�Y���і��*�8��K�l��ȓS��,P�(�?�����L��$Szp:%�im�\F~�cĈg��� ֋�1T�P�*炓���=y�|r��,G�yd�J#D�E�ƪ�5�yV/C�r�[ ��$=�����
�$�y�iC�d����#�14��`R�d��y�\� "�@͌0L����� �y��Bgz8�C��!m`����y�@��V؆��+l�H)��L�y�Nٖ?���S`-W �;��Z��y��"Er�rR-�InL�sQJ��y�ɽ~D>�)�JOS/&D`1I��y��= L��9�C
H�ح"�"�y2IɀgJ\RRXC���B#KW(�y����D� �aG�e��{�EW��yR@�B1UG@�V0���QN���yR��7P˺��p�I5NM��P�'�yR��%9���(�<F��xb@���y�%[b�!)A"�09R<u��m �y"�D�v/`���X *�䭩K���Py��4S�4��F�A6�b�'W�<9Ǘ y�1y�A_���sF��G�<Q�aG1`y��J�M�i��%�*_N�<�1�_�.�D9��+U	�~�gk�Q�<�w#m=Ԍ����1	:���#FW�<Q�E���Q�p������Tl�Q�<Q�j)����P�)/�~��!�K�<A��[a2�	��ȼZ��� ɗl�<�L�<q��U��W����`��<i��1 ��Sd�M,�޹xDG�{�<�� :'�`A��N�4D<�Q��}�<���ʠ5�z��ҥ�)?�0�Ey�<��$K�3��̘'4��4��N�q�<Q3�"f�x$(�-J(=�0��'�Yl�<!�]�$d �K�̖�~uCgBCe�<	�i�;���V ��.�֍j���g�<a�ʲm�JLAڿN_��9���n�<)f����s�K�q�gmQj�<��Ʉ�@��`B��E�ޕyC-�^�<I�$�yU>��֋�/#��A���d�<y�Ɇ�ER��R �ح;�6����]�<��6�<�Y��2h�}b�p�<�� I�a��W�b�|��Dm�<���$}L�%aGoU~x4�B�L�j�<�Cǯ>����@Iz�yr��f�<� ��B�!���"fe�="1��r�"O�][��ۚ_���˰�W�f$�Tc"O�Y��8N~�`�V�TD�`qD"O`t���/��=�ҫZ�z6J�1"O@�z@�!R�4�)�'�3��0���'T2�'e��'��'��'�r�'Z���Հ/�����.Ȕ~I�A��'>�'���'���'���'C��'0ԩx�IY�C���e�G?E��u�'�'�2�'�B�'���'e��'�R�'���P�FI��9�#���H�%�'vB�'#��'%2�'?��'�R�'Ä�z�-/�r5p��O�b-��d�'nR�'Q��'!��':��''��'��M)��X�	&��KĥA�9;� ���'$��'G��'{b�'0��'1b�'��a��=��3�h�)��ʵ�'�R�'x��'-"�'�"�'�'������kP����)X�+w
u0V�'��'���'O��'��' ��'¦\[�*D(?TȒ��%��G�'���'���'B�'��'�2�'�����4O�4���eɍ`Z�)� �'�B�'G��'5��'o��'P��'ƶ���֊{� �q�eA�M�ny���'��'cB�'?��'�����7M�O �+��r�/B��^�(�!�O����O�D�OL�D�O^���OJ�d�O��r�i�&���O@�jtı�&,�O��O����O��$�O���覉�	��8+���h�jlbƣ�,e.e`"����O��S�g~B'�O�Cx�\8v�Ŭv�A,Յ8�� �'i66m(�i>�I̟�k�-~j`C��	�{�,�oA�D���""f�m�G~�1�V}��r�	0Y}��JF��%�n��1���c�1Ol��<��i5M�.�!�f^�c�2��0�E�,y�anڭ%>�b���R���yGA�%Os"�æ%�`����R	�T2�'O��>�|"q,���M��'�plx���||�6�&�i�'��d���<`2�i>��y��p�� r:�G�k���ILyr�|@`�D$����>ђe�p֥Y�TEm�3Aɂ�\�O��O��	p}��"���#&X�q2��� �T5����O�	T%_)j`1����j`����14+��ٔ�
5�z	!���G:������O?�ɜU�H�k`�X�4c��̣n��扰�M�CC~r�tӆ��ӼU�H�o�/�u���A\x�۟��	�|q�KA����'��)P�?���&�S�ȼl�h�B^n�'z�)�3�I�X��$��E�N���(�¸Q�|�bћFAŅ��	���ғ ��y. U�4�D{aQ����I��M�3�i؞O1����O:���/��T��P8t��5ܵ���<1C���Iv��������$
.~9�Q��(�$]
B�q���l�a|)g��-��n�O���0
C8b2���UV�p(�z�=O*�oZP����	��M�d�i�Z7m�5FB�{⎓z��`h4���=pY�f�p�!�.ke���I~���}t")1v���-��"fđlRXP͓��?��M1*�����ެ ��PD�L&����O*0m�Cb0�'mP�F�|B���l<Z�L�� c��X��'U��������6���bغc�L3H�&�Qv.T5"*6�Pm?�M>�(Ol�ĳ�N;D��7��0%�<2�2�_ʛ���5���8�O��4�E���2#н���V1 �$1�ON��'���'ɧ�i�Jʌ���&�?������N�Qا�E&`6�Sy�O 0�����0�x���K[^��|��l��9�|���?����?��Ş��
�鲖��1aҠ���#F�:�X$��(T�8�' 7-'�� ��D�O��R�ȦpY$��M8W� s�E�O��Ä��7m??�)VC�f��4���W�`mP��u��X$LA��K��y�V���	�`�	џ�����O[RA��A1���k�k�_TV���|�"��3&�Ot���O�����ɦ�] ]�()t
ǍE��m�Df�I�����M���|J~Ѥ�$�MS�'�е��;B|(X���Qe�lI��'\�	*D�ğ@QF�|"V���	ɟ@��C�9E���p�ƒzX��QݟT��ǟ�	AyB�xӦ�Jqi�O
���O�L��@4uS&E 7h�z���'(�I�������͘ش6܉'��1�s�%� ��Eg[0}��yQ�O�AȆ�B
R���"-=�i
�?�"M�Of��b
p5&��v��~F��y��O���O2�$�OJ�}��'�$tڣ%\!Ma��ܤvz�՘�� ��b")���'��7M)�i�M�u�ܭY��+7���<Ysӂy�\�ݴE���i[d}i�i��	6=�iC��O��H��)H@�M8M���BR��xy��'B�'��'�Iʷ :���Qቕs��<� I�9V��	��M�B��?I���?�H~Z��7@��@"�&q�c�FZ+g"`Z�T����4Fl"�x��$��*�~$!tb<Se�I+7/թK��K��GNo�I�TWXQ��'I8�$�T�'^x)$+��t~b�y�I�S��-Q��'���'�����_��3ٴ@ؐ�B��[���h���I:��&O�pΓX�����b}rFf��u�IǦ��s�6kv�!#<@\B��PHۜ�m�H~	A�B8��ӟ/�O#� �|K�h��
��d�7a���B8O���<N������
����#E7��˓�?��i	,I	̟��mU�wk00�ӏؙk~�A��&�kO>	���M�'j����ߴ����;q��;Ǣ�tB�X����i*�Aq�H���?9'd%�ľ<Q��?���?ɤ��Z?������`�0��l �?Q����d�)IE��D�	򟨔Oj�A'��7m|�E����<L��m��O���'���'ɧ��[! >�r��l�n��FO	W��-7R7M��<1!�j� ���B?�M��xɉu��9,�t<;��Ӈr�B��G�O0���O.���O1�˓&3��#@(|b��B�a�4>���	 )�Ɣ�g�'2�x�"��X�O��$�'�\,$!F�G�]
�K �6%����O��"�L�Ӻ{'�����T��2���<,�)&�F<Μ����a���'X��'�b�'wR�'����]�!_�S������F�d�E�ڴUQl�K��?!����<IS��y7�^=Wr���G�ċ%%���)`�"�'�ɧ�O5��RR�i��d�{=a�
��e�ى1=Oz�`���~��|�X�,�	矠;�.ο[�"A�@6n�"$��J����Iԟ�IGym�j)X�e�<���r�	��M;\���sɎ�ͮy1��)�>	��?�K>���GP(��*:�"y�sd�N~b�TМb�i#<�� �)�'�B��O���q��,Qy��H���:?"�'["�'!���ğ��P ]�[��$��d'3X�v �ʟ��ߴ./(2+OLul]�ӼS�B=~s����D �0�$�W�\{?���MC�i&����i��Ibc���O��P5���6h굁jar��S�IBy��'m2�'0��'w	Sy!t̸�J�fU���"N�d��	��M�0��<A��?�M~�}�&U�˷ub���"����P�]�,����'�b>	A��yG�X��B\(X�1�6[��� �4��D��(�b�'��'��	5'�!Hp-'}�zLՐR^��'W��'x�O3剢�M�0���<y�&Q�xB���I<.Ǡ4W�^�<��i=�O�	�'��'D���/�p(�$n�p��(�
9z9TrQ�i��I*��%3����ߍ;@��
���\�K��4�	b�(�	����I̟|��My��4f E��Q�d+1hR�'���y��'���|�dy1b��Ȩ�4����3񩝵	�Ǡ���8�[I>���?�'	aH��4��d�4�݂'�A�<zt�ǫ��ظ9�'��-�~|�_��֟ �����B�p��r
�)u�D���Xޟ���oy��~�19g��Ov���O�ʧA(��R���E.F�0 S�����'D�5��6��O$O��=-�H���P �| ��K�Av$A�ӍȞ(��� � �Uy�Of���	 �'#^�u��)�
�`�F�"�����'��'`R�Or剄�M�	�:�����D�l.H�dfm�ƨ�(O��l`�i.����M�J�)9 �p�%�>aB�P�JO��&Ag�nK�Nj�|�	�P��T���,�TÄ�<�S�l����\�^��3�dأg
���Hy��'�R�'>��'�rY>��"*�	Sg1hCL|{���eH�M���#�?��?K~��1���w-�%���RTےD2wM��l7�AB���O"�D)��O����O�>��t�iP��9Ef�H)�N�?�b�{�1fR�Ď�*�\�A��-�,�OX˓�?q�1��H
RB�>��IA�T%�ג�?9���?q����Jڟ��4��On���O�$x�fI&dv�r�ٛ<wh�4�O��O`��'���'��'7T�����g���Hd-3�Er�'��[�D��ܹ#`�&����\ő��H�l�$W3/����O�zU.��f·;[8���O��d�Ol��0�'�?I�eE�.��i��fK�gCf@9����?y�'�,�k.O�Im[�ӼG�8l���I�80ՄT�����<���?!��kdT���4���L5	U����'���Ҥ�@8W�����g���y5`,�į<�'�?���?����?�wL�ˏ<BW|tj����P��@����O��D�Op���䅔_��)2��	?H�S⨛�1�Vy�'�r�'�ɧ�O��mKW�зg��h�G�X}���R)R�U��O2�z���%�?�vm"�D�<a�
ĭ:�%bIYY�r�F��9�?Q��?q���?�'����例97��Щ'k�)I06Y��A�i��9`�Vݟ���4��'�$듪?���?ϝ\�� ;ю�(h����'_��`�4��d�����c�Oo�O��ɚ�E0���$�<z��"��y��'WB�'6��'��)�-��ұaو*׎�[ �� mz�D�O���^���B�Mny��e��O�qZ���dF�y'C�?Vk�DY�=�D�O~�4�D�ZT�b�T�Ӻ+�(Q9�幠GY1v	��1{?���'��'�������ΟH�I9�B(pt��Qp�M"�he���şx�'57�Eq $�D�O4��|rE��)y� P�i�#{ߎ�"�+�t~�N�>!��?iH>�O�.]��"�{*4!���ÚGЀt���R>I���Ǳi����|"tN���$�d:���
2���J ���:�͂F០���I��b>��'�6MB"!~p�pUy5(J�G�$1��3a�OT�$��5�?�tX��ɖ�I�T)�p�b��f��,�l�Iğ\kV��y�u�/�<p��i�<� ��У)k@%C�O۔=�V���0O�˓�?����?����?���)ʬg�zmpiڒKJ��Ȃk��3d��oZ�ur"]�Iԟ��T�s�<q����ᜄE���YN��[�`H�f�}���w�ҍ'�b>m��J����H�1�,Ñ+'�]Hg�@��̓B� �3"�O��YN>�+O���O�q�)�	ek�[�)Y&Q_d9RŁ�OB���O��d�<���i�b��T�'��'e��`X����r�-G�P�d����$�O}�"xӀm���V�6�胤ح[�@i睯J�<M�'����ƤËI��EZ`���&CɟxZ��'���8D���<�A�
�6?�|�D�'?��'�b�'��>�ϧ/��d�����i��X�C'��[����;�M�3"W��d�Ԧ��?�;'��L�"�_+�t �7�L�j�����M� �iĂ6-�0�6ma���I� ���Ӵ�Ov&��άT���ǆB�SZ�r6��c�	gy��'���'���'��$�,N��\�d%ۯy�P1c���(e�ə�M#p^+���O�����Ă�jRz�p���J��@9��(V1$��'P�7��Ԧ� M<ͧ��' �"�d S�O�ZP���)$�1c$(?].U�.O�x��̕��?�T�3��<y�lο?^��GX7\�����?q���?Q���?�'��d�ަe��$c�d)��>f��SE��bv�5Ab���4��'���?��?��Fƣt�@��.X�5x:�U�=! DX��4�y�'��`���M�9O����j�A�\�c����CX��#=O����O^���O���O��?y�ū�Q�ڼB��U�m���� ��$���`��4^d�D�.OVlG�	
B���F���W�fu��|޲�$�t�	����"}2�n�j~��tw<QȒd��0��E&��'�(�V�Sğ`˱�|2V�b>牵ZP��,��(�����:��#<i��iv4I�vP���IW�)�)&�h³*�?F��D�$�����Egy��'j�VB*�T>!0Y j����dSlлfc���Edԛ{�0Y����n�П��ԕ|"B�1X؄麷�Y9w��HZ��U3�x2�h�v���.��5+͒lL�]����k�(��wM���DMP}��i�.���lQ�G���1#*\6H�zm���ۦ!�ٴg6�Dk�4���эq�����J��˓j�h)��D�d�*�2�@ݧ|r�Γ���<|O0�@b�ñn�HD�뚣q�I )�ئ�B�	�Iyr�'���<mz��*CNV"`0���䤓	h� ��2�M�MK�i80O1�
@�v���		~bQ���6H�u��C��c��d�=��q��bj�O�����	�v�vJO��L�` %���ax��yӴ�[C��<a��|����O:i( s��I�;D2�2/�>�Կi4�6�UF�ɐu ����/���(�D�3���\ �q��h�"]g��IH~b���O���yѨLCIU�X�ƅZ��݆*Ex�ȓ2�3rg'6N:M� �-�&���?;��$T(I'�ɭ�M���w��{s��G���[sȉ� ��'�t6Ӧb�4N��5�۴��d� z���}o@;�@��fl��wQ�i�]��f-�d�<Q���?���?����?1%Ɋ)��cF%�(���O��d�ʦY�t�џ ��̟�%?)�	�oT���&/I?:Ia��)�2zl���Oz�m��?1K<�|R�L�>��X�| J��T�29�4;#C/����"+���0����O��>�	#S'��;PY�"ʬb~��"���?����?q��|�*OP�m��8�b��ɵ$�`m�`��"w�d���~��	5�M��>ɕ�i��Di�h�+���T��@XrƘ3.����%�B�;��74?ɷ������.�䧛�C����[��Ŗ1I��y��O�<1���?I���?A��?	���j��d��=���"N�
a��=�b�'j�/i����7�N�����'�P�D���_㈅P�F#I��<o�����"�O�$%�8Dd�&��H�D�Z*v�8�5��_��kB�O�c_h�R��'�(�$�ܖ''��'.��'6����E�7ni[3!�4 �����'b�Q�D��4~HL0+O0�d�|"b�ݲu}f�ӆ�U}Fu� @Xi~ⅶ>�f�i���/�?�Qr͞�N�!3d��:�s�yy����w�IsC]��S�Dbb�Mg�DՂ���B�N��$Z4�W�2�� ������	�x�)��my��x�vT���VQ�����?x�V�Y�k��of���O�o�J��G��ɒ�M��"�8W�<��oQ�t0>hʆ�@ o-B�i�H��i���*�����O4E�'E��(V,�4!���h�Y�`]H�'����<�	x�I�H��v��ԭ^?���t%R�W�@,b ��VX�7�;?�����O��-�9O�mz�
d N=v��C0Ɣ�N��ُ9�R�'�ɧ�O3���G�ik�� Ap�H0�Պ:6���Q��`���4)�p�����(�Ot��|J�S-�XI�Ǉ�!n ����'�d�B��?i���?	(O��lZ�u�b��	����	�~�\�-#Zا!�&
A:�KVh&�I&����O��7�䆳H����Gi�f�d��$E�k���O�����\�4�F����S�Rr��͟(�CH�!8�z`��C��c�<��T$�(��������G���'W��`��X�f�T���E�<����'���Վn_��4�M��w���6C@�O�D|�3EzW�@��'�B�'i�,�rS�&<O����,8�ة��Z�� �9�$ �U��黀������8���<ͧ�?���?���?DK����5�F�F�TP�ˋ��$���u W��������&?	�	�GB��Y3���Ts�l�2��<����O��n�&�?�K<�|"Q���R�!'n�:tf����Ʈ$�ވq7O����c�����cPƓO��gM���20أ�lKUxț��?9���?9��|�)O�nڤ-?�)�	�>�aq�ǉ+H����錸c�|��5�Mc�2Ź>��i"���o�d蠐'�ԡ�e�^5ZL��1��w�7�"?զ� <�	�䧘���$���5a�4/�|�RD���<i���?���?����?������,�&KV']����GD2vJ�I��4.���O6|7M5���P��)�r���|Y�Ο�v�!%����4/��'	" Bߴ��$�(�
@#�I�16[$�XuI�dТݹ�5�?��e;�d�<���?����?Q��:<�Dd���;;Kp	����?1���B�E��i�؟H�Iߟ��OU����]�;�\�T-��w�&h��O0��'��'�ɧ�	GI�a�En�p��= '-U�>4���d�)�
ؠ'�<�'`�����YT)A�`��H@i��T-:�t����?i��?9�Ş���YŦm#�LD�e�p0����!xNv	�dݾ�F������ߴ���?Q_�lB�4o�b��r�`G�´ݬeW�)��i[j6�M��6m5?�R#ЖqC��ܬ��d��"2v5HF�T���tc�{��<a���?����?���?�/��t�i�l^��cKm�����N�m�i@˟h�	��%?A�	(�M���`$�I��xsR�-��Y�����M!�i �O1��ܠ��x��扦b��0�Bn�	c}`�+���ɒ/��P�'��&��'���'mV�J�;@
!F@�'��K��'���'AY��rش<�z�(��?����*�JS���O,�ӯ�zU:��H>��@Y�I:�M�Ĵi�O"d�	�~�:Io�
TUp`�R��l��"^�݀d�b��V�����ğ@0M�uҖ�ö��5q|�۳��̟��I���I�E��w�i
E�ܶ �(Upa��m���Q�''V7î+/��D�O!nZI�I��$a�F�ɥ�!�>�����yX��I�M#��i�x6m�N�6m7?�Ń	/ ����(rW�%�CdT1��CTɬ	�j�{M>a,O\��O����O����O:�����>k҂�j�&�#?�L��ʩ<��i���%�'O��'��OE"�ַ���ąN�4��H���� ]�v��?�����S�'���`�ϕS$Py2�ܾ ���2�H�+�MS�^��֡�G���4�$�<I��A?���@@�B!����A$�?a���?����?�'��Ц��Er��
�C�#Py�#��wN�1���|�tZ�4��'���?a���?!QgN�x�� � ��Sk�!!2!Ъ�@5(�4���Ȅs�Щ�����#�� >�tI`���0+L��V?O����O��$�OT��O<�?)�O�l��g���". (J��|��IΟtI�4I.`��'��7�+��V�V-9��D^��2A哀pz|�O����O���3&@N7=?��mYwn0�H��Fb��b��m�p`����X$�4����'�R�'֞��W*�x0�!s�^ �@� �'�"S�Pc�4�����?q����I�*��!Q��ػH�h[���b��I�����O���<��?�[5�)�h��
�@�Q�lݽUu��P��æ1��$`�K?IJ>��OU�5��tX�+ڣ7���0�K9�?A���?���?�|�(O�n�%�����T�u��ԁ0�L�MI��j��<?�Ǳii�O�@�'���L��D+)5���u��&/�2�'���0#�i��	 Zu)��I� ce$���DH�4�q	-YE�Ģ<q��?���?)��?�-������TI��Q��O��j��d�ݦ���
I���	%?��I�M�;B=D�(�F#c�鷅�0U�Y ���?)N>�|
��ɕ�Ms�'>z��욭G�\���3l���'ͮa��$Iu?)I>A*OH���O8}�" �vJ����f�MZ!���O����O��D�<Q�iX�I��'���'�0�%�C�0#��(�R����dMI}"Hcӆ����I�}i�@ 7ܓ0�X}`u`B����$a�$�� -���I~�Dj�O�����<��MS�AшU� -��"������?���?���h����T�HL8���� o �X�珂�~�R�$�ݦ}:4)�Py"d�Z�杽d|(@��4$���B� 3q���ڟ��	�d���
릙�'��| �m��?=�!)�1Zm����O;1�r��W�G��'��i>U�I�$��؟��ɍ\mJ��W��<YET��b�!LV��'��73�
�$�O��D?�9O,=�@���3��X
����m%q���?����ŞH��Ys���,��Q�/8X���m_dê�0����(��[;*��fAV��{yb��q�<�k_Xq�"/۪5:���[�X�I�4�i>�'�*���]�2�J�6\BIJ7o%Q�NYSs�Ԡ�yB�u���@	�O����ON����x��Y5G�ܜ��e�e"���ԩg��T(6� �d�>��]-8�eac⏛)�B�Y��2��	֟��	՟T�I՟��T�'as�8YC���G��׊ݓ�*8 ��?)��c�vh���I��McN>��
	9Zl�$GS &�0���	����?��?yF�� �M˜'B���� �d�&A�U8B$`է6,YUO	��?�P!�$�<�'�?)��?�Վțe��a����SҎ��ul��?����D�⦉w���	�ĖO@���D��ljb	 �Gt��4��O���'@�6�ܟ,$��>��#�H�}8N+�֫q�|��j 8Pӊ��cƷ��4�zU���߈�OByie��U�h9��͗�*�p��O����Od���O1���H���9m�΄en�=&�ȷ�0F ��V�'���yӰ⟴�O�n86�TJ�j�w�`��I�.}q���M;�����M��O&)۲����$�<)���d�l�Jv+KA,*e��+��<Q.O���O8���O ���OPʧV(<x��S79"y��n	*����D�i�p���'���'���y�{��.�X�Zh
fL߽Y9>`���R�jEr<lZ��?�O<�|j1�M�'�"$jԎ�1�8�pc����#�'�hـq�����1�|R^��I��l�#&V12 �:B�[��F�&��̟d��矤��Dy��oӮK�m�O(���O�0�7��>o A�m�*M��;�-(�	5����O���"��l� �@ß A�@� MԌ
;�	?AҞ����߰Fb>�Ƀ�'F���i|��wh�@�l��/_%��d������	�8��Z�OF2�9Ka�a1AɸC�z�BG'�6,?2�pӖ0se��<���iP�O�nAt�,K)[:aP�0�RM^.f+�D�O2���O*���!m���3T3�+��ġ�CL�%��x���\G��ɱ�k�1����4�����O ���O���**b`�!��x5ĝ��HՑB��4�"ԬD�"�'R���'�����I'*tM:D�I�Nie��>Q��?IL>�|�D����<�J�
�dm	N<~��	b"��h~2�"x�Fa���Q�'�剋j�53D@���]�-�g#:��	������i>Y�':��$�,�j�Get���Yf|�MCV��%�y��f�⟤ѩO8���OV���&I���Q��#�t2�����8�s�u�b�{���
����>��]�K#L����)AW�XW��8\J8���|�Iǟh�	͟\��d��Q��a@ט�l��.u��I��?��6}�6^�1+�I/�MK���䊿59��K���֚իԠ��La��O���O.���
6
7�y���I;r0ڒ�ܗj�:%	�� GV�����'-l��R�	fy�O�R�'�ҫ�oe8k3�X6��
t��Z���'���M�֤�7�?����?y+���eNAz�1���6�)�����Q�O\ l�M��xʟv�Ru \�7OޤJ������[���+c��@'A*f�>��|�P��O�ɢJ>�a�Ǉt�H�V�C�@aH�.�;�?���?Y���?�|2-O(m��� Ku�۬`�D@�3�G^°��#�x�D�O��m�F��l{�	ԟ�ZGbT�
��A���Kc���<��%~��8og~ZwkT��ԟT�cs&�f䀟uu+�`��7߸q����O���O��d�O��$�|��V�^yӁ/S/)�0��!�ɥXm���ݪo>b�'3r��t�'��6=��h�"I�>�ݺ� [�r��<�f�O���0�4�<�$�O�e��a�<�Iža# ��	���{�������6|8�8��O�OR��?��vc�(�+��p�L5h�	{����?����?+O��oڤ5�,�I؟���)S2����>��a�ތ.��&��������Oz6�C�z|�I7̘�ͽQ�+X3s��	P��Z�,ރf鲡$?UzS�'沍��Y��UQҧA�����҉0
fe�I؟�������R��y7`$��M��+ͨ+"ػ��<G
��pӨ=�g���ٴ���yw�H|��� ��P9N��u$%���y��'�2�'g0�:Ҷi��	�~;��ݟ�ъA�׸=���g�VX|ةQr�9�Ķ<ͧ�?���?���?!��C�s4�,k&�&qm�x��CɆ��ϦIRF�k������ '?�'R�}h��*KT��h��"'Zi@�OP�$�O�O1��y`gm�(y��ܓ�B5Z��)��R�4��6�7?Y�gL�ZH��IU�	my���k_ ���=&��q�F�3JSB�'�"�'&�Os�ɨ�Ms�R�<��کp���6fÚ �aVc��<aӾi��OЅ�'���'�2e��g��i�b�*�
hx2nT�64t��i��	�Q�������߭�3DL�q"�8��G�V��m���Iß��I՟h�	�P�����
��8�	C?Ja�1 �/��<����?	ղiD�d��O�pnZi�(�}`���3c���Z��$���&�L�I�I&z��n��<���\9���@��Un�b'�>���[�#U�����W�IOy�Oi�')"��'R��c�f��*��\%WXb�'@�ɲ�M�n�����O��'=���#k��4�ڌ��DD*C�B=�'�4��?�����S��`Oh*�-����uPxq$*��=�T���1alx��O�Ɂ��?�6/*��T'4�]�>���HD�
(bv��O��D�O��<��i�́�i�jjΩж	O�a ���䋏����M3�r	�>i��u�}h2Ț�z���n��eY���?0�&�M��O�����E1�K?9�@��J��)`+I�6��'h� �'-��'"�'#r�'~��N�V�;c���l4:S֭JiL��޴!�����?�����<����y׍��/
���p�FAd�|�eVu���'3ɧ�O��lӀ�i��� �XE�W�d�tX�Ղ��e��7O~%�$�ŕ�?y�	?�ĥ<�'�?y%���Ԙ�6��?p���	S���?���?Q����D���3�ry��'����@����M�:2�18u��Vs}��'vB�|� �WD�zv�+v�v������-~�f�0�wĎ|̧R�l���<�?�Ż+����T%P?��ۢB��?Q���?���?��9���9�+C',V��P �$l׆$80��O@Doڔ[�'d�6%�i�5�5+�-s�N�:�tE~ŢQ�`���Iޟ������oZL~"]�_�j��S������`�>yUvMy�f�X���ҙ|�V���ɟ$�	П���� �7}r	�"%��T���Dgy2cӬ� �`�O0���O����T'@f�jS���%�<`B�	ɬ\@D�'-��'Lɧ�O��de�-^$t3��̇aц�x��P� #f��O���j�!�?!1�+��<�ʛ�zcB1zDD,^����b�X>�?q��?���?ͧ������4�џ8�6���,露9��S� U�a%�̫�4��'w���?����?�e�ɓ:g�pXb-��6];cm�S�Y��4�����nPb]`�O�O��#BYf�0�g\N��<����y��'A��'�r�'fb�i�2~��
'�$\�����k�"��$�O ���Φ=@'C�|y��sӆ�O�� ,ֵT�4x1�h_��8�貀<�d�O��4�����or�.�Ӻ��$��Y�2��<b~VTJ�*M'\ �8Q�'D�'g�IџX��ԟh�I'���D	>O��LS2
H�K���	��'��7mU�
�p�D�O���|b��J9D��D�8p$���I�v~⃩>���?�L>�O�$�`Cn;L���� Ȱ�K6����b�i@2��|b%D��@'���Wl�<2��5��!�G� �P�G.�h�ݴ&�� ���F'Z��K�^�y8�����N�������?�\�T���9�T�����<��L�E.��X����h1 /��I�uW��<��	�<�rL�l�r����8�8���E�<�.O����O��D�O&�$�O�'8�j�ҳ/�; �8�P0��)��d	b�iZ�p'�'	��'y��yB�v��.ڷBP��
s�J!)��z5�˵V"���O��O1��i��
yӜ�I-��sb��$Tj�@�j�]Q~�8'�\	J��'�&%����4�'6^��̢eT�8s��_�0\�r��'m��'��T�pIٴn��i��?���K���K��Z&�н�6�J�f夼���$�>I��i�"7Zd�	�:�f١R@<!|s'� y)��9xP�p�'�M�L�M~B�g�OR���)���kRi��}`RcЭQ��:���?1���?���h���d��x8��s��"{n,�V������[즕У��Ly��mӾ���� L��c̨4�-�! 67�Ɍ�M�i��6M�!��6!?y�'�hz�i�#��d7 W�$�6U �TaH>	)O���O���O��$�ON�be� ]Hl装s��P�B��<�q�i(xi+��'��'��y2����#e�T(�0�'��.VǦ�S����a� 1&�b>���kK	�0���e�`�õ�ɿF�-���Sy���'�A�	!@�'��)\2Ŋ$%��Ts@����-p@0��I�(��矨�i>�'��7M� "���D� & �Ȓr��"E$5�V����Ĝ�1�?#[����� �	X\��@̃�Nm�m� A-'R@������'��� �#�W2I~��;l��i
`Ş�k����0�U�.�0���?!��?q���?����OR �2r�%83� ap��8�?���?�ǳi����O92�m��Oby��ģ��Q9V���x�L6���O(�4�J�{�isӚ�Ӻ��&�I���@�/ï����@J�bV�m��'P�'��Iԟ��Iӟl�	�
�v�Y@k��I�����(ռ1?�L��՟�'�^6m�e�����O^�$�|�&� ��h�hE*W)�����P~rb�>����?J>�O���2Dܮ2�H�[Q�3��HYV� 4-R5避i�r��|�꩟�%���F��"�;F�[.7��d�ß��	��P��ןb>=�'�7�������&>����"�� shL�
b��<�ֿiw�O���'B7��3Wj�!�S�0�҅r򈕨=[�Tl��M�wc9�M��Ob�2c��Z�ȼ<QR煃t%)	��!�����<Q/O:�d�O����Ob�d�O˧(��J`��k��u�u�Y1���pA�i�2�!�'��'��y�q��WL���K3��?O�00sk�E,�dmڊ�?�O<�|���J��M��'�hj�mZ/�L v��V�̠�'ئ���ğ�`��|�_����Ο�1�K_0��}�"]�~���ҟ ��˟��I]y��e�|�I�+�O���Oh=�"ͅ�YV$�8q@ϕQ�V�"�E6��+���]�I���ē�Ah�&�'b>^9�G@/hn���'�||q$�I�LQ�<��������l�!�'�uCq�� ���3��3PDN��p�'���'�"�'��>��I' س�aH�Aը�:Q�Q,4X��0�M���Z���$�Ϧ�?ͻ^u>�C��J*#Fؚ�dޚ���d:�F�O�6�E^�~6-=?��d���<�iQ�q z���$�"�y�Ҡ�,BrPM>�*OV���O���O:�D�O�	a<X��`�b�
�,8Tx$E�<�B�i�liI�Q��	Z��؟�#��\�2?<�*��l��u�SA���Ē٦m�����S�'G�@�� ����?n���T��S֎�K���,GT�˓%#�X�6��O4Q�M>�.OD���\�%�~�����1.��@�em�O����O����O�I�<���i̾Ժf�'j Uc+>�"��!��B鼰!�'�N6M2�����D���%���M[Bg�(3a�K3�1k�ޤ!	�����4��DD$l����'-�B����N >�3�Ua�d,�g$�Z��O*�$�O�$�O���6��B�8|����XN���1�B����I֟��I�M+��|��}��f�|��Z��D�W�ʬ0��ȧBeM�O��m���?�S'	mZ^~��Z����ض�#e^Q	��9u��f��̟l���|R[��������I�|��Ň"~�Tő@��-�z 2�nV�����[yKq�*]����O����O˧c��X��l��)L����']:�|�v�O�O�S�b�� �"B��&t!V�- �(MY i�8C,���@kAEy�O� ��	�\�'�<�B��^�w�Xl�g-��VOЭ*��'T��'�b���O��	?�M�!õd���@���8 �VE�7�a�6Xk���?y��i��O���'"�7MO�IA����%Ͼ4ö���HϺ@�4U�	릑81�צ]�'�X%�r���?=x$S����'7�I
����K���e*l�`�'/B�'�r�'��'�哱oT�5�&A��l�]l�tN�ܛܴx�,,���?�����'�?�T��y�L�3`B
q���<`t9@�L0(J"�'ɧ�O,�!�F�iH�Wr�(�HgH��2���@W��x����C��Ӏ���H=��)4�ٚJ��Q��R4�09i�^�H����O����ؠl���� GB>S�ƤQ���8GzP���#6�Ҧ�B/8g�׾P�fI��AO$g�vĐ3e��Թ�f�D�B�����-�
m�p9��O'��d�j�BD�V�T��8�4�$s\Μ F�F1y��Y���# �4Qz[��e�N�˲�7�[� �DgV���P�r�D6J����&��A`NŪ�H�#�b�õ
.��4�)dX��mӭVb����H�g�4�)���g�v�F�Է�~���O�ciV]o������R�����kܥ�EԿ_Ū��۴�?�J>��?	��ݵ��'&��k��������T.(1�4�?�����D�"� 8�O���'����Y�f�`Ă�b��Q$���d�RO����ODekD3�ID�!a�(��|�ԥX'g�0����ɦɔ'����y�����O����h0ק5f(NT@�;�#��G��-"Qb��Mc��?q���9��'%q�H@����/%# �!5��]��x�ib���%d�����O��D�T��'���"ol���i^o����D�	}p���4,�lPk�2���OT:�AY n1�Bǆ"3�M�wm�̦�������� ��m��Ol˓�?��'�,��O�f�l�s#J�#=���}"F�$(�'���'��ҊG�)zf�J��\����
6��O|�CI�R}P���I^�i��kք\�1BP����A��P(�L�>i��/�䓾?����?�.OJٻ��66^l`)6�]�I�\���E�::�`�'���ܟ�%����ܟ�*�_�
	��2�u]&��lv�a&��	؟,��^y�a��T����[5t��a\��,�Ĉ��RR�6�<i�����?a��R��M���"��9��	:�0����+��tk�[���	���	cyB�:k�'�?1���~EZ�x`⍂}�zɊRJ�����',�'4��'�ZLx���6�rp��	�дKZ_���'O�_��G�!��I�O6��៘dP��ڀyk��W%^�X��I g�u�	��8�ɛ:U�L�?��O�>=��k%#  u��q��h�4���-�ƅoǟ(�I�����
�����H�&+S"KfZ���ݹ2�`L��i�r�'��`�&�d(�Ӏ�>�G❮h�x  �/Â6mD1���o�ߟ���,�����$�<Q�!��*�C.�)S`��CU�G@���S?S~�|����O\�F'�%����7��(r(�Z4�R̦�	ޟ\�	U�D}��O�ʓ�?��'�XizV�*dlh�q�N�~�⼐�}�і-�'yR�'3�陛k��u��c�Ƞa�P{�7-�OA9rL�Y�i>�I@�&xF�;�ڕ����iF&(�)N<y�����O����O�ʓ;����t◀0)����w����R"�:$�'�R�'v�'��i�Y��$ݮx���UA%9P�:p�v���d�<q��?)����u��Χ~�Hr1)�:H�.�ca��-k(`�'�r�'��'��i>y�II8rIQħL�%L|��O*VG�O<�����d�O���|��.�8݊���hR�$� ��H��M2��i��ON�$�O��3�b�8C�'�0�"L<o�@��g�C�Z(j�4�?I����dG8A
�P%>����?�طE�7�XE���w��ly��-��<�f�%�?1M~��O��S���_�r���ަ{�t��O
�$��h���O��d�O����<��h$Jf�W�3J|DiRu��j���O6Ƀ6V?
E1O��҉�co H��ö�L�O�,��6�i�t���'�R�'��O��)�cϞ<�^�I�h,H;(@� BO&��!� +6�Py�y����O�(Z��W�T�yR��_K;�
Cc�Ʀ�	����Ij9j��H<ͧ�?�'��	�ڰq1x�8%ܯh)�]�ݴ�?.OpQKW/Gl��'/��'2,�H�)3�'V�J.IてBO*7m�Ou+E�a�i>=�	񟤕'�UӲ����D���L�F8�r����ȅa����<�'�?Q*O��dL�n���r��1�d���0�H��U�<A��?)���'d�6� �P3�^�,��u�EJ<Qb�!�i�J���'�2�'��U�Hp0(�-��īѪ��Չ��^�E�N諕l�,����O��$�<Q���$�"Z:���?&rl���%$h~	:B�#M���'�b�'��X���!͕�ħ��I��܆@v�ip$W^����i�2�'�Iϟ��	�5|��Id�i<{�9�ͥ^Y��!AKŢ:қ�'K�[��5%���'�?���C�Y�it�������K�ݚ�gK�I_y2G��h�2���ПH#f��/����Q�~�L�cW���I�n�	��Οx��͟���pyZwF�5���l��Po
�޴�?����!*��^�S�'H�,����% ���
�J`��n��:����	��8��ПX�lyʟ.��@	�8m��Cq	:.�SR�e����0c�"|���W$y���Z��0󔦍�p���c�iQB�'�A�y�8O�)�O�	�d��ex�iQ1g��9#��ؖ^��7��O<˓o�<x۶^?�I������ 7g?�U��k�f�����Í,�M����©��x�Oer�|Zw�̈�'�@)(z�H�f�A�4��Or��q��O�ʓ�?�n�ʟ\�'�.MJS��%8�m' 8Z$P�R��24]�O����O���<����?�!P�0+�d������|˥ƥ4|� h�����Ov�d�<����XB�O�x ��I0W����Ď�
e���h�4�?!���'��'_����M���M;A�E�z�H&�Q;zx��M}��'���'���&=�f����EL�l#giۉJ���2TE�pAP�l�͟ �'��'62+K��y�Q>�&(�+	�r�A�\%=8��㮁��M[���?�,O���HD���'9��O�$�é"aA�(ڃ�,0D�#��>���?)��m�.�����m�:|�F�Wc[�>vv��K�M[/OXU{��P劣������	�?��O���v��i��d���U�Q�Pw�6�'�҆ϗ�yR�'�r�'uJ�)��)֗E���yv�L$g��o�1�4i��4�?a���?��'q_�	Yy�Mي^���q%
�QI9�r��',�67�����}y"�)�OH�����>�4�Y0��6D�E2am�妙�I���ɓCC�͡�O4��?�'���{���~�L �q�-F�<T�ٴ��tm���S���'�R�'���0l�5��ma�O �|t3xӄ�DG��'X��֟T�'YZc�X���(�eR�Ӣk�n�*�O�X��9O�$�O���O2��<Ic!=
q&� E��)g8���l�"h���c'W��'��_��	�����#���������y!��ZW*��C�z���'ub�'��W�P���Ҳ��T"��2���Z�Η*8�X25 ʛ�M�-O����<���?Q��/W��'���yT	ƚh�v��GF1L��u�۴�?����?����dV�{����OTZcZx���N$ez�e�bB6�Jڴ�?,O0���O �dǷj���O�	&��z���B��$�υ<c3�6��O���<�.Mg��S�����?� �J�LY�l�p+I0(�t�7/�	��D�O��d�O8	�;O0��<!�O��!�`�O����q�T�g?8�۴��'�60o��I���Ӹ����N���g�wW��{G�M>���Լi���'�X�'��'���	O�AUp��$!�2 �� ��ԍϛ&�_�V&"6��O���O��ɛD}P���� w�j���ou���4@Y��M���<J>�����'
 �:��B*�8}�`��\:m8��~N��	���	�E~��O.˓�?�'���H��Ѫ,��A�� �m/�Ԙܴ���O6��r7O�ҟ(�Iݟ�Hʤ�`�j �E1U6��C����M����v��Z��'~�R��i�]�D�G)=��0,�����a�Fo���d��K��O����O��d�O�"+F�����n���Q�!��b�˕Ƙ�p�I`y��'��	���I��h󄑪T���S8�@$a�I�,Y���ky��'��'��:�f!ӚO;�HE/R���풊W!��4����Orʓ�?����?�j��<A���e+'����(���T�Tn���Iџ��	Qy�Ȟ�^��'�?�1�acvş%&�p G��\ n�埴�'fb�'�rh�y�>��Ϛ Q��;�a�m�:������H�'2�A��#�~���?�'c��}y���,qu�%* �?�6��U\���	��4�ɠ8���	x�	o:$*(�Ƙ���E"z|������'�B��c�w����O����֧u7��z8�yaD[�\�($��'�M����?���Y�<�����D-���0��1 �6KH��1,���:7-;��l�Ɵ,�	��$��	��d�<A�	� i<i�����RJ��2�
�V���yb�'A�II�'�?���@�K��ɠ���3]Ĩp4	�*��F�'<b�'6v�Y�.�>�)O��d����ć��� ���7 �Ӡi��O�B�1O�Ɵ���ӟ��6�+-L4��&��K��lNƱ�Mk��@pv�CBY�<�'��U�8�i��01 �1����bFϓo`�,Ʉ�x����aU�$�O��D�O<�D�O�ʓm(�,��ce�>��'��X%Bg�R�~�����O�˓�?���?� dN�DŶh��Ǘ`�"���� .}�����d�O�d�O2�-�4��7�`�2 _&fZ0܉7*Ֆ]E|Cg�iP�	䟠�'Q��'��@C$�yre�:!����������&��6�OV�$�Ov��<	��
,�����aA��P��۴;��M��0Z�i �W���������*MkP��k�� b� �F��+-K>U��J#�i��'$�	!OT� SH|r����@[�Vy
A)�Bٙ[~E�叇�W=�'���'��P �'a�'��I�>/P�����DC��!zf�%Rʛ�U��Y�)Q��M��\?Y���?��OZ͋$� je��Ȇ�_�g��X�i�R�'�8C��;�2����f]�w��e�(�t�b7��nAh�o�(�I�`�����?�'�Z�tq���ʿ��ᇭ׫=t�6�W5L���|����O��)�F��FD	��R�
�K�ݦ���ȟX�I^&rɡ�}��'c���VP{�R%,�x5Sw*C�CZ���|R�=�yʟ����O���A3p��}:'��C#J�#N?c��Qm���P�5ND7�ē�?�����[���$�N�C�'S5�t(�(�S}"	8��S�d�	����	NyB�V�v ��!G�N��Ifᇽ?"�``�>��П�'�\��П
4�0��5Q��+X��T!g�se�	Ry�'���'I�IN�P�O����8����j���O:���O�O8���O2@cV9O`�aΟ�(xvab��ƌmq,���c}��'��'<����u�I|�ߴ��ۀ�C3ZT8�Qh��&�(6m�O��O��D�O~aB�!�I1*J>1c�F��b]��#3
NT�7��O����<�TQ��O��OZ>���E)
j�чʙ@�h�G�;�$�O��A���D#���?!	c�T���X�t+����Da��z�n˓d(�a@�i���'�?���|W���`�;4.W�p�-�W��tw|7-�O���_,y�����}r�(ݏy$|��4)��H��6�S	�ql��H���<�����'�~�0r��uִT�VBԓ�fx�@lӐȉ���OL�O��?9���v���#K��8�b�M�5��i"�4�?Y���?y�"_=1G�'���'s���L.52ɋ�0tܕ#إ^O���|�� �yʟ����O��$��+I�]�!G�1IXT����BÁ�̦���7�P�J<1���?)N>�1#^�4[��"+K<8�Sꚼ+@�}�'�ڄ;��'��	ԟ���J�F,���g��4��`+ŋJ�vH����	����?�����?	�"&�e�GN��,!���T)�8Wy6qhb*�?�*OR���O��d�<��AU�R��iւ;��D��M�`&eY� S�Q������f������nQ^��I�~�T�������}A �[�F8�;�O��D�O�$�<�ō�[�Ol�����:s����B�A	���o�\�=y��8�@٘���?��'T"�2�%)�b�GbG;C>�)�ڴ�?I��������O���'���
�0P���&XO�-������?q��?1���<a-���?jp� ����g��>~�qh}���N���v�i���'���O*�Ӻ2��Og*,sBDӦM�ԍh�E�ަq�	şr��x��ث��$3�ӂ5[�$�#!�3�� ��֢�6-Vs~	l˟��I�ӑ��$�<s�#"�rRl� )%�[G���@�����yr�'��	Q���? "D�ij茀�¢0z�cź0/���'��'�@5Q���>�/Od�D��9J��:�$�� ��E�:��Hw�L��<����<�O�'�Jǿ/p��f-��}���SB-�2Htp7-�O�{��Ms}�W���_y���5�N�1Q��+��&Xu\ĩ��޴�M���b�ܑ����O��O�����'��q*zM�,2>�"�� %r�Ieyr�'Y�	����ş0�"�M`�*wk�]��r�J%\�?���?����$�)y�8%�'h�T��b�ʠd8Tڲ�PCڐo�Hy��'���ȟT��ҟ��BE�~굆�u��C3��$-�����"�O}��'���'@�I"&1d�������Rܩ���U�)>��$�ӆjR�dl���'���'����y��>ӃœN�Daj�o��kF��Ŧ�����D�'�|��A��~���?i�'O.���	Ǌ0�b�LL�
��8Y�Q����ܟP��e^T�IY��'����!O����U4�p�,P�6T�h��@��M�4P?q���?% �O� �VK �K��x�B�p��i\�ɩ|��?�g�/�i������5nX)#�7M��A���n��ȟ���/��d�<�(�9��J�k__{LU lVBǛ-F��y��|B���O@� %��ԁ��#P�����[�q��ӟd�ɞRG��0�O���?��'{��@!Kв ���pT�%r�Rݴ�?Q.O؜�6O��ß����@�$�4�sF���;{������ �M��'f:DW�,�'/Y�(�i���B	`̨q�K�� e�ln�*���9��<q��?����򄈃��0+7�
`@L��I�8(��E`���s}�R�L�Igy��'�"�'q����G"L��e�ɯ��Qvĕ�����O~���Ob��<��.ĲW��i^�9����e-��0�WhG�"��W���	{y��'���'g>EP�'|X�cg��Jf
$9G`� &} Y�2CzӮ���O"�d�Od�[X�c^?��i�	eJ3crk�D�=��{Ѡuӎ��<���?1��b��ϓ��	��U�t+̮K�[��,907��O��d�<��(�}��������?	��*
T�(�ޓ[�8�glݦ���O��$�O蜚6O���<��O�� #�LW�.u����bB=ڮOH�$ɢ3����O���O����O���3,P�m�&.b�j�� &
�t��7-�O��>�:c��� �u�Î�<�&�;P�Nm8�,�b�i5Đ�G�tӪ�d�O����8�&�p�	vG�}K�i̜Kzhс�
�%����۴W�$YEx����O�%X�ƞ)/��r4�Y
/���˝٦���ҟ8��Q�zY(K<i��?1�'Y���P�N��MX6!�A�J4���?���?��؏9$Z%`BG�'	��IqHɺGߛv�'���7�D�O��$?��Ɣ���dVi$k[1r���ٷ[�T�gG'�I���������'Hl�ڴl7QP�&�)1��1N�#M3`O �D�O@�O"�d�O `�a�>�ڨkfc�#|����aJ69G1Ov�d�O����O��D
p���6P�p�+�*@ ��	��ux7M�Or�$�O�Op��O����B�_�֠�'X��d+��.J$�)0�@����O��d�O0ʓ`��ԃr���	VND��CN H(� -��`|F7��O��$%�	;�~c?ћRDAG��j�F�ex�l�DKw�>���O��$�O��0�|J���?���*
>%��AW��d�gˈ�BK�� ƙx��'��Ӥ{h�1�y��:�胩EN��ɂ�J����i|�I�u)�%Jڴw������S�����"2����uI�a��sv�-��4�?��c��Fx����4����gNa*�ũ�J��K������6��O����O��I�_�zI�S��2OԈ�'�A"]�H���i�da2��d/����l�h���sS�_mV"�.�:��f�'t��'�0�R�m1���Oz����4�b� L�[�dͦYѪE%�/��V�Pc�(�IßT�I�u�~��	�8����E�C�R���4�?QV�WR�'���'ɧ5��V�Gw<�b����X��Aϰ��$H��qO�)�#"��O��8����)P^Ls�IU(B�9��'B��s��`´�cR����
���=O��1VL�;#.2eɠ�ȥYQ��Ao×"��\2�C��VY�(A,χ5�^�m%�.%\i�դ�%��,��mȁ�
<�!F��b12�S�*��	��LH���MRnPB��[�@��؄��#4Rmpef.2���D��C�i��ғN
�%���q��9�g��_��FD�P��`���5\?���4O����'���'����(�$@�,��P�Юh1P�b���_B�C#k��$�2��:�vmZ`�Fu�'���
jN�\��!nH��v�[Q	/'�栳 	�r:���7S��
�AE�2��O:��R�'��)�?��xJӂ>ŎXI�oV�`�*�Oj�����;-��{�-�aLY��'�.O^�1����p,Ƥ��L\ 
H��04Op���Lz}b�'��ӞN����џ<�I2Z:^��geY�I�p���KȾH�e#We��M8�}�'�ޱ݄T��S���'��]rA�a��L��%ܩF_ ��>-� )����J:k��O?�$��'���9e�B2�:l��Y�a���ON��%?%?m$�,kg�2T���Æa�
�݈&�(D��r�)Q��J��bN��w:���&]h���' �n8SuMUܖX�g�u�@����?CH?)��Q����?Q���?�g����$�O�I��̡*����O��}��2�NR��\�OL ߚ!�V��1���I�:X�Թ��=L���k[0�8����#N�y�G��&�:B��?�=)wk��1a<�� H�g�茳��[?1#��͟���I�'$�I���d�ʝy\vLR�(]��B��:Ƭ��ӏk:�F���$������?��'^�i�C�q��R%iU=��h.Y�$u1�c]�%��'I��'%��X��'��2��ɐ�D��5d�)�!�e*@��Z��(1��H�-q�X��	�Q"��Q��C �ZT���c��쨧 @�H֠ȷ��q���1�O"O��@��'~�*�*j|PW�_��N�҄qK�ўtFŏ�o*�JM�<g��Q�,��y�FF�<��:��\Pj�8��W9�yҢ�>I*Ofhi��E}}B�'���&MX�[��[�R�P�b�*�/"���������|p���x���j��8b���Z��������P|�l�A��d�n�����/1�Q��k�W�g\Z����4�:����AhKD 	"q���ol��"P(4���`a�j�(+X�������,[7ti��*3-K��da���<Y�	O�=�g@_^5�gc�V����Ɂ��.���q�Bl�Lh��t3�X�<	�dXo��	��H�O�B|Ӷ�'���'�nM�ƢL� D"q۠#G�k���!���RCt���.V����(��OL�b���Q5,�������ՉW�ĸW� 0zV!߰]���`c�O?�$�0=�X�Hv��.Mߘ�!2ꚯs���ӯ�O��n������O��I�[jx�k�c"�]�ŃQ 2C�ɑl1D�#F��8*@i�Vc��e�"<iF��M3�bN�]��n�2j���s�� �>�����?�‪<��Q����?����?I���x�D�O|$A�e�2(��8�i]�Z�2�"�ʃ�+����M���3%��)3�'��pkd!�� ]� �UaP�p��+ �!�ߍ;Di���HS*��䇠%!h�q�oAQ8�����̲FK�M�}
�dfӢ o�M��#��ӈ^Hތ�ai�1LtH��+ �xB�)� x!����	ZČ��'F��\쀢i�m�'���������
�16���Pğ�#��t���W�<)�a� Bz��`��]_�=2��[�<���U�:KX8iP	�3�Y�� _�<�� )	j hzF"�/h\�A��P`�<a�Q7y��� �~ hT�Ha�<ၩ�1a���i卙�]j�hyN�[�<q�FB?"����S�7��-b#[�<�R�b����U�-z���b�P�<��i�8�d �%V1�P�W�<��¶TءR���  �%��PZ�<!7�
1׌Y�N�1�,`!�G�a�<��d�*bܼ�p$��)c�k
D�<A�^���h%�<!�ld���JI�<A�f^<L�B�ϝ8�����H�<IN�8f7r�+2��R�J�J�J�<a.T�O=����*���,e���O[�<���r���&��J�z��,�]�<ɧ�՘J͆1 `�Ѳs5ԑ�'A��<!F�P��tJ%hT�9���� s�<y��G���Cіh��RׯRk�<���lf\�B�`S>J�&(I��e�<��`�8m.AT��b�� �[�<YF/M:q���gjE;��{���~�<�ەf	 I���42�8}�$�b�<iq�_h���qr��4dl,�e�w�<�7�ݛbV&��$�˕ۈ�:REu�<iPE�x��@/NآU�f�i�<1BJ D���+T�O9֐Q4�EQ�<is�]�b%��h#� m����N]L�<q����#�]�-�,��It �c�<�ȓ2ݻA��@/P�D�_�<�b����dcԌ�}Q<u;�m�f�<�Gk�~��C� ^�r�LFa�<��$����H���
�{��-��$�\�<�s��X�����3*��Tc���V�<�w�҃
�I\�0�����P�<�u��<��ذ�[�'f���`�w�<ap+�)H�NP��"�)kkֈ��I�I�<1�I/U{��6E��A�n!���E�<����~��3E+R�u��i��(Kw�<���;IH�]�%b�6B��u@��u�<���Q�`Fn�+� �P����LXM�<y�/�^>�q��'����F�D�<�p�æ4Y�A���ث"v�;q\�<Iq���U�RDH'Z��qf�X�<��mm�6�cK�����V�<q7�8���!�f�&J�58�B�G�<AV�Y�@������% ]VБ�HE�<Q���:��z���!0tXK2�h�<�C�:D.m�U�Z
Q��+�a�<�b�,V�� l0���P�dV�<q����W^�i2�P��>�(���]�<	�O��2��
u,A*��Ԫ�&c�<�1j�.� E!��
rZ$Y�cn�a�<�B�U�7)l��g�]�q�u*t�^�<�	�4e��+G���2*,���A�6:�ϓcB"�Kq꒬!�D���M�l�����I�gJ2ًSJ��-����
�&��E��<�!�=(�5DBÇ9\��R�џ��W	��la�Ŋ]�XSdm�	$h�}��"O�!0N��E*(���L�2_�*W^����
J1IqOQ>�0��Ƅ����֝(^�$�+:D������2z(aCI� |��P��*�I�t���S�? ��!�&�gö� Ö\�JA�Q"O�xT�6̶1��!ޅ���U"O�A5��H�b�Fώ$�VE(r"O��+bn˂C2!D�Ř!�NP{Q"Oİ���L(5(�Y合QO� ��"O�`6��,N��Ew&��@Q�D"O�<���A{?�aA�ņ�r�4\1@"Oh���N�	^`�s��J���T"On��1hVđ�'�rI���3"O� �5�
�-�n�b�GI6���"O�@@(\8/�Di�@�&�j���"Ob飲�@�8p6����1$܁d"O�(��j?�ћ�"���D��"O$4@��V�d����ݣI����w"O�a�(���1�Ѭ,��"O��DJc�tY�KQI2��D"Oj�áC"+e�B�钯f?�P@�"Oؠ�T�вJ���e��-A0,� "OV�2c�@��qT�^���A	w"ON9XC�j�`�IPl��Er�<Zu"O���� �A��,��wE03�"Of�3P�8z��#ۚ\4.��"O�đ��K�nU��PU�<l`���`1!�`���Rb�C8AR���c�(H��y �!�O,��H�O��#P�V�Pei��+�(�r(zs"O����O�2ݸ\���'d��u �	(;h�`��\n�l �|��Pi��ġ��B��ysG�<����: ��ڔ&�-u#P��+\˦�P�Q���f
x���s�h���a���kD�b	>��"Om*��5�VH���!l�}�2¡��1*Q0J�c�S�Q�џ�[ �,E�@�pN
#�����L3�O| KG퉆7�T�BV�z���çB��X��0��D�d����=�`�8�Cݹg⼤��U��4�Dz�i־�r����1���'?݉g J
><"P!�i�9 ���3�"D��)i
4C�-�d�L�1GY���|� lC�n؟El�K1��~���i�hܣU�!��p1��1b	�'*,�CʕGNx I�Ɗ�Q�Ux��O�9p�X�w֔��s����O:Ԣ�� �.�:5U�Yy�|Q��'rE��lQ�4��8g)]�\D����Ϋ$���&�˨3Ҵ����2�Ҭ�E8K��;�	 ݊"=�R�M��V�*�e����D�)���/������'fe�'"O�l��`\�e�0�W�ޘ[���t�i��iҨ�5}��wRs?E�ܴ7�,l�E�p�a�e� |��Ʉ��.T�Z��>��,"`������)���AܩN�$��l��1�6�H�Y�Ĝ��HO�d%Q��Hp���y��dR��I&ɑ���ȥO"�pD��?7-Ȁ
��`����%⑑!�z�"@M' AD�p?Q��
+M<�@q �G���w�  �	:(�H=�2���Tc���=h��ӊ>w̻����	�f���3���4���IMcN�K@�E��4�$_��D����ǒ\���!x��#B�C����&(���'9���O��� ��&ʶ�ZrO�m�`�	� ":,�站�m)���KfRUi��9.%�T.��.L�H��a(�g�Seb���,�o�<��ΐ�=Q�|ԇJ<P���1��2Z2@+m���@IZ#��"��� C4���	��cqy��S�~Ԃ�:���F�1�K��g��$[�+��C��܂��'^�8".R�D�z)�(��!x�m��$�ҏP9��[��Dȑ�[�����y'�'9f޴�s�Z 9���"��0?�ыi�>�{� �������%�.3ܰ��3%jy⊞�d:�q���ߴ\�^!J4푆���y�c[�5��W��X�L|�t�͜ΈO�m(�*Z�xJ5"�����>|�����53��Bc��Aſi��8[�n֑��A�e�F`F{"'�(�R��j7/��MtF��y"!�(a�q����4 �t"���'��E��4ɦ�h�� #Zyai֡R��C�dJ��p?Y@�o�!�����5Fe��A	�5� ���=�ܬj6&�-�~��H,�#�nE�<Q�9���0�g�5G:p�a�ӿsc m�'@6gj��]�n�1�c
1?�y�v�T�<�P*侟��Uσ�%��[�'��Z���i�
A����R\��1*(<ٌ�ڣ-)�@��Ή�aT�]��=q�(�g�? 9*�N�0,,�C��A�0���>ae	��M�,�!��?ٲ�ޯ(Uș�1�� ��t�f�@�M+n��T���~�
���Q7+��۶�.����c��sڰ+V�Z���,�B�E/U��:4�=�O}8�)��D}��Ze�����0i��B�KV���1>��+���1P�)��d5(��(��Y3e���v*�= �}���=jFa|��q~ppĠ�o�qd ؈wy�|w�ȋJb؉�� ���z�/ۇ1���Z���3iD�U��k�?�^8C��1>H#<!��M����φ_�Ҽs� �"���S	<����,Fx-��"F�Q?�����Hb��*��l�dA�k�?c��i���(���2�f��b�j����4��K;0�b�����2ޯl���O]P�:,O@��W�J�K��9��VϏ4yv�E��O�1�� �[�'#k������R��́Uȍ�o��\2����_���kS�.8E\��$��uy��]-;�s![W�ѱ-�k��y���P$ڶ l�'��J��"��?q+a�6d�6 9�iK�-�,�*u�
o� ���)N43Ұ���@PC�(�`�鉅%�Y#��+��'e�X�O��9d�0dĠ(��(`K>q�Ţ,_
)cUJ��U<4���L�8~P-����"v�	Z���(p��ۇ#�-S(���펷�?c���=���0���?)[�y٣��H�'��@S�ў,L���R�ۧ�&�K�-SU}�����O�*\��`ۘtX2�Rף��l����V�ʅON6O�x;��ŕ}Y@e��E6lQ���s^^]�ۓ)��!���K�[�L������Y���BR�%�������Hc呥(j�İ��D��X֤��1f��Y��W�x�&�S�	���I��	�a�`8�47B�pi2m�^	�� �u����+��nj�5$�ZV�6>?��$ŲTjXSgH5C��H&��:zFBEP�@!$,@\`P93����tk��~(c�P�ɖ;kNY�DD@�px@�qb��T�m���h���ŋ2��HkW�p����B�
�X�*'%Ԡt1v�	3��^(d�����V�ұ�t��l��x�EM_4{ Jc�#�,.���#�\�D��i,��a���tQ�#?	'��=*��-ӳJ	�]�L�	F�\��"�?|O�� �;.����lX�|i!ŋ9%LH��A�?I����?��O�5�#�.d�1#e@n�11e�h�&t���3[���f@+��>�!�'C�Y1���	��(2b��a�������<F�‰b�|b��>B��lZ7���0D�4��<��M@#���D���������iyR#+��'P1�+ 	vn]H�o�����k�m�,�q��-!�I{��E�L�f7�����1�A+�)��9��@��+]�,Y��ߔP��T����<�@l��;�RD�W�ƊRF�O��'����&+|cU�=Jh���z���J��':�K�h�6�yլU�"�rJ�/<�ra��~�`Ǵ*�W�Jk �̟���?� �x�(�hq����s�$y1�ɡ0 b��z��Ǐo$��vI��sτXg�t�|��BJ
� y9�LI�q�0��>�|"Ac܋S�ō�22��R3{y�l5��'ڊ���j	9~���O�]�$(�/��d�SL��4���"O( @�+d|p܈sjVv�r�|�b9��v�"����"2�� ,���ˑ|�t�5�F^0��ɲ$<�x���}�F�{��#l����g�ZA�Ð|��h����X�0�**��܄'lJŹb�ĥ�ax�AQ��O
5�t�����
�n
&&"O&� �퀨 �4��5%�����"OB �C��2 f����ҳ#�ν�"O��Q���/^�tA��¨~wεz�"O ��&�GU��0p��  v&0�"Oe�1hG. �� =[G�y�v"O��9Ģ��nQ��ٖhm��"O�\���2 ����!ag�<7"Oΰ`KҎf��I��dB ɷ"O�����1~��#˒`⸣�"O��80��8	Lf �!�]?T(P�jV"O0�:w#��,�����nԂ3By��"O�@E��PsX���-�~p��"OLiy��G�pR�#�1>�5"O@*'�;����h�Q���� "O�$H��Y�dwNyt�{�l}9T"Ox`�睹0ZT�teI�Dʠ���"O�@g��j��P��1�Ѝ�"O\�
##ֹ{����&� ���"O�8i7�P]�����D�>�Ґ�`"O ���f�@�%C���;����1"O��ugǁ+���+k�l�Hd"O�=y�A݋+��`��7}F\��"O�,a�(
T���:��[>|:�¤"O� �u�ł?C�H	cV�'m���"O"��� ���T�03� �{�<-�"O\I�#.Nb����Y	U�&�v"O`�8�M����QB+��L=h�"O�qY`�;<����]4i�*�"O�@(S��H�B��(DJʑb"O�D�f*�2n������*:^D��"Olے�A;X�ՠcG[�=�-�"Ot ���3\��d*�p�e"ObY�b&��<��Zu��1�8�Q�"O��[F
ݣ�Ԁ�C7L��Z�"O����yK
�wgۄJ�X�"O
�ŋ ME������,!"O:�񥅝.f���fb7Wؼ*F"O j�H�Y)��� ��.��4��'"@��$��/� �
��t|hI�	�'�Z���D0c,-yA��yR�A3g�ޱ���	�l)p��'����yR,9)��)F���q��x����y�jN�D���r�� @��]I�'_��yR(u�4�)�kW2wN�����y�'I*��t�r��5Vh�˷����y���y�����F�2n�y��+��yț-,q"�1��]B�C�͜�y®͜Dt�5��ĉ��Hhy����y�ᔚe{t%8B�M�v(��)�-�y�޺8��H!-�]����N]��y2��6i�<,"�G/u�H8�"l��y�8G� �k�"�t)���P �yR�A����J��_vP�P�Ѩ�y�KGm`�fσ(R�X�{P"N-�yRE��'��X1$��FW��(@�y��]�'�*4�����7	N)�yb��[��"� �*hI���=�y��8�`����&Ua�	g�Ψ�yr��Aa8EA�&Ux�{�ʈ��yR��Z�$�"�G��p�1�+���y��Y$&�cԧ،=�I�oV��y��S�"��i���V?Ք�	�g�4�yBߙ{&��x�LR9c6!��k�yBOű�xa3�b��α%U��y�BD���C ħĪ�U��y�N	
7I��ċA�f%���y��Q'"D�E�����9�D� �E�y��6G��@Ї���=S�Ȑ�y¨-Ub��ԭ2���7����y�CK"m�4�S�՘7��D���©�yB�-dX(�1pKI@^��e�C+�y"&�0��X�K�"=�̹�e`���y��&�vT���ǘ5?B%B��N=�y��ϟ���s�U7bl]
�߱�y�ɀb0�t�bU�<�dp`�*��ybm�/Hh���!��4�d��#�y2<���E$�"�髃���yB�/*�J���Ċ_W������y∄�*�TQU"��E��2]pi��'@���L�fG*� I׆z* ��'���h��&� ��|�V!X
�'
L�� �&B�f����H�^)y	�'�ă�샾k_\��7��C�*4
�'"Jԛ0�	>c� +bJ$4�B��'n"�iv�ѩw�8�;� ��WPp���'@��A�<RV� �.I/cFZ��'y�MqV�L0��\#�['b��d��� L�C_�t�v�� �B-IĔi+�"O ��pgҕ�xDS��J�f�x9 �"O��a��Q } �mP$���n����"On�p���g�"�ԥ'"�T��"O4�����3Un���OL��"Oh=ZBC	�[ڤ��%�.��9��"O`2cf�.3@F���s�bi��"O|9{�f�v�&��N��p��!B��'��	4xJ���h�
����C��,{j��� �Tr=����B��#S$�� �� 7n��ȩg�nB�I�?���@��؈q_b!*� OnB�	�4��	���\�d?(A�aÃ{b(C��1" l�b�۰|a���΁�K� C�I�x�R)���rP����a�97�B䉶TafL�fʄ)&в��E���C��*pP��J�0d��p�J��-�B�ɴͦ���L�2wӐ-ZTI�5�dC�I.��c"I
�5��@��;6xB�I!YY�2'�2 ^���7  PB�ɒ!mPr�_Z�~e����18B�I-g.�a�n	
H�07�B�gnC䉬���jEN��	T	�p�:C�	2����T��3��k`�̤��B�ɂ.p���%�E��
pU�b��B��q�~�c���B�����p�B�I�C�p�rp�D�m��=�V�&@�B�10^!�� G�t��
E�v
jB�I�MxU����0�!�6k\�tV�B��!s
r�y��A�Z\�Ȅ��k��C�	�P"Xad/o�Ӷ�B�[�C䉦b�!�"�'Q�@ ��_(�C�OԐX����-8�9pd���C䉀(��!aV!e��6��0:��͆�!K�4Q���-���+t^d���|�&\��lح	R���m)�8�ȓa�����ג^:��0�	D�l���ȓ[����,����Km98�ȓW@����3j����$_7����'��}��A%=j�qc��`����<�y�Đ�58rq�F�яP��E�&J����'��{�aN?t��[7Y�ED.�v��;�HO���d�%i�lS"꟧���C�@�!��@dx���h���K�iٌ{	!�$~���˖�ɝ0�:@�0"�w�!�d�F���C�m�Ä G�z!�ֵDL��N��uflT���X�6}!�Ė�V���Zcł.c�ҔHgf�5|!�L H̵���q��Ps뎆F!��'T�6d��Կ=lJ!�ÃW/x�!��R�)����W�G�2�@Xش��2#!��2Y.p$�e�Y+f��b�I4V1!���-a�4h��I7��i���-�!��Z�����a?D�����[�!�dPpH� � ��Y[z���O.a�!��U5Pj �r�J {���5Hm!���<9��L��n�[Q��"�!�_�kq�ث�&���8�	2�LM!�
a/R�����)��!���;&0��DJ�}��		6
�N��L�2��'d,B�I�&��.��pg~�����b�!�ę�jt��p#BB�*h�Tƕk�!򄍩22�J��,�F9{��K *;!�d��F����g�N/�n1�N#)!�� d���I�tD��l�{�N���"O�q����]��e�:	�@٪3"O�M�T-��"=�-jD^���1�"O���O�G��١L�G���t"O�"N4OӼ[���O���'IF���$Q����fK�B�݆�y"��:n,�#��F�$QyՊ���y�H[� uRx���B�@ɤ
]�ya�~��3cd��"�\䋤�O�y��ƻIKJ���ꕒ�5(����y� �dd�(�%�<,�~e+s�
�yB�Q=X����,��5�&0��B��y2*\)2���K����k1�Q��y"-��V�� �LH<�x�+����y��-���OG�e����D.�(O��=�OZB�EӄAE�DZSi��-��p��'S�Ar� �ZᎬ���]�}�&���'���
�n�)mx���A
�_�Z���'���sF78�T�W�[�Xw��R�'����M�Q�v��5	_�NS
�
�'��-(�`��KHXR�d��7N!�	�'���c�lU7��7�H��'Ĩ�$�&��͑W!P�c��%B�'2d��"�O����h��X��Y�'��8� �'��Q3&O��4;���yr�G�隠���U���I �yrI�W_��C��Fh|�U��yR��� 2�����3@�l�F�_��y�ŗ�S������F9:j���h�y�N�0i��=*�D�d��PR4c��y�$ٌ\j�:�U	_����@D��y�o�H�D�Z��ޮ[�6 sĪ��y��23"�Q�Ц��h-�,�Ӏ�%�yR�J� �r��Q�P�2��P����y�U�|�H���">�@-�W�M?�y�jR6~<u�F�L�:�adc��y��$x�ЈPvQ�)�+�3�yr�ߞ^��@R^2�׋�(�C�	52 |B���,~V�e2�Ĉ�q�C�:ٖ��wɪ5ʼ1���
�C�	&TZ��"Ť�'"��|IŇ��+3NB�)�j�a�ț�w�hP3�-Y�b`C��+>&D�P%8�����2Y�zC��M#�a�H��5q:��d�a|B�"~��U�����> :��+�B�ɝ4�� J�����'��[�bC�I�?�Ġp��yv��t���
.~C�	�*%jp�������y�M�-C�	2|���hB�� y���!)W_T�C�I�4��9�&�(uc�\�#(�;+�C�	�2��<c6jW8K��BBI�m�C䉫���Bw�N{㤽B�eַM��B�I
z �Bb��="φ�"���/,B�ɀw�~XhD��9����B��a B��"c<4���0¸H*cL7IFB䉥L�]�v�ɫ ?������./��گc0�jS΄�H���&�!�D������E�,-D�<�%Q65!�$�� |=H�	?Ӯ���^;- !�`Djm�D�ӸW�b� �ˊw�!򤒘!$
���b����Ң�,2!���@�����&�����6�-A#!��.Kv����ߘO���W�X(5!�D��8�j��ߖ���#cV�E!��  -�@e}�P�2��:�"OбðiY"?��x�錌(��s"OpX6)�CA�5!b��$�d�� "O`e�η/�~ɫ�(�1L�<pS�"O��#��� je���ME�H����"OreĞmz-钆Z1bX8""Of��%'&�=�bh�	j
T�*�"O%��i���%"U�"H
b��1"O����aO��Hi�,�r�3t"O��b�Z,p��x�FNS�n�R���"O,}BP�!@;<�P��Ms<���"ODppc��.��A\�7K��9�"O�m�R@n`�R��֒��#"O>i���ҥ�Ъ��v�Tk3"OD�ir)LF�P�(�3�(|Zt"O�`(�N�.�z�H�*F�D��`"O|�#k�6���`q��-F�<��"O&�J�DR�E��J1[�6TD"O�pC�H�S�lAh���d$�&"O�9cCFF<�� ����6DY�`"OJ�*��$	@@mxEᛧ �	�"Ot��"뉔pj�+�M_0"dA{R"O��q���%
���̛>Y��{�"O��aQGս0Ji��F�=�@<�2"ODй���B���ɰY�,�V"O��y�L��8�`:�f�Z`.��W"O�������)e\�ɂA�D`��b"O�0�tiFs��hXb�-bGX�C�"O|0iAEYNbv,��Q�7'��d"O,1��h�rMiqH[�n!@�CP"O80��X�obL��Թbi<$s"OTy*�'�$~�a��"�\`�7"ON��%B̦<8��I���2"����"O<0�F偵M���`%*s���E"O�	�蚪}6¥:�V�,>��"O�8Q�����8[��Cdx�"OH�f�V�Y%n�@���0P����"O��Z2�D�z��,
/8
T��"OR}��k�	l|�ܰ�*W�r�ձD"OT��-�?!9 ��٭t���"O~��7�9Aδ	�-_�ˆ8�g"Ob�hfAFEP��,��B�Y�"O�� F3�TQ n��<����A"O\L��J�cւ�qL�O,D�j`"O��P�Ŏ�J�N�,�&*�`���"OB�ק]&������`��䒣"OhY1a�y���"���mQ�)�G"O���GN�,;`��2E�f�`"O|��FC��)�*I.��Za"O:�V&7bn��vn��~����"O�aa��'t�n��TL��h�@"O|�9��??2h�'�΂ɨ�"O"L��B�
�P����qA"O���#b[66�.��m�
_�$�@q"O�9A0��h쌹p�P������"Op�2�T:|>����K��d�HI+�"O�����@*.���s͆?r@��"Ov�C%�R�)���3�*ud0��"O�`�$j��G�Fa��i�((�l� $"O�)!�I�N�������w�7"O�m�ʏ.�v�a��H/7c����"Ox�腢�"1�4(f�"X|�Q"O�-[fF�;uԄ`qD�� aG"O���G�L�=�"DQ0/Ӫa�g"O� @8��B��TP��¡Յ\���k�"O���q�K1��I��KS;f� �	�"O&����Z�l2M�6I��YB0J�"O�m��o��H��V�aQ�i��"O�̘�a� vw,(��ܫR����"OPQ�)�>`�+�&�#h�`�4"O|��"�8O������G�l�T���"O,����8*zf;	0LPi�"OQqQɆ4	���1�H�Mu�P��"O�$���5�zD�T.��lX6��e"OP}�E�*\I|t�-)4JJK�"O4]P��<m��aɶ�
�����*OƁI4=,��!��33�l�:�'~�qhF��2������t&�da�'F�� �!S+[�41-Ȧ���	�'s���͇~�@�Qch��+�'�H�$Q�)4%��E���H�'B��xAжU�Ь��E�(����'�����#�#3{����u�����'�0���HPBt{�����|a�'���h�!ÊUf��'ĞI�t��' �mZ��Wm�,r4I�*Kf���'gN�x����*�B!n��Z�z�;	�'�V��g��J�Z�1VBڑf՞��'ր�TC�x
 �cU�4ք��'��S4�ܙ�x�)��2�ݳ�'9�I�`.X�u��M�Ee�r�'�0E�5nͽf/F���H��h��X��'�H�Ҳ.�4N����/J�L\q�'l�}�ᦉ/�dL8x�ڨ�'���� j<
����Ď��@
�'��\H�d	182�GgX,S���"�',Щ�Eɘ1|�@7k�H�L��'�T� A닜I
^��̢s*n���':&�ga^=0��|kW��9�xA2�'�<! ̪-l�-{)ޯ&��� �'����Q,�.��X���D�jv�b
�' �p��fX̘��ć��T1��'3&!�F��$>�&L"v��[Ҡy�'�6�����}�h̩�5'Y����'r�G��@͜�
5��J��h �'X��I�H["AbN�I�͚6{$X��'���0cס8g�0�UL]�|����'5~�r@��,��Pui�?�� ��'NŠ���>:1 ��M�Y�|�;�'׺�����<!�psT�ќW�f,�'����"�׼~r�9XԬKTzr���'�|K�
Q���SCB�G�h��	�'&�E#5�Z> >�`�J2n���Z�'o��T+؄���Y�o��m>	��'(���H�`�0��-��8c�A�
�'���2"NY�y����O�17<U��'��17BP&'\<�y��5�h���'"�i�1ni�T��k�='�l��5D�xd`y-j�P���Қe�>D� �@4Kj�|8$�)	cr�b�=D�${�NqL�Ժ`��(r�J��wM:D�|it�,�����%��x;�k9D���w�Z������E�p���5D��6F�#Ya�0�ʬ�����4D���DF��2�-`�l�=l��P2D�H�6'�){��x	A���5�f���n,D�T�UAE�i��!àX/nPda!L'D��!lH�\|FUP�	tX��q"*D�� a��gX�xB����ʦ\��{6"O�HB��+i�����]3���"OV����A��5X�Ǉp����"O�4I�&�5�v8P�֊ܖq{�"O�,���_�3K �����O���"O�0���P�u�Jyb���L<�� "O
��b���g�d̸2A
 �lxi"OP�<.��P�"\&@��l��"O8dXA�S~!f�z�^	-Aā �"O�\!���t<�e��9���"O,L`�yD�h���=`��D"OL�r׫O�w��F��4�p���yr��-�j��RA�r�b�	���yB�͉О��"�<�F��P�=�yI�#�^1�v�$���!����y��I��}B.����4�P9��=a�y�C�<{��G�9�����	�?�
�'���Kq�˂��.ę7�1��'�&|���H_d
dBg��u`n��'%4�瓷BM$�pՀU�q�
Qq�'���O��Xd+P�	;����	�'�ƌ3u��=^zVq����5J �	�'S������r�Tkv�܎:.�@�	��')�I�6EU�0и��զ�4��i	�'=x�
��ʚ@��%�ĥŲ=+<=��'�P�H�k��I$R��+��'��� m�(-�M�s((ʒ�
�'{ ����Jd`mۦ-Vڔ[
�'{p3���?&�Ѧn��;Z��'�f��2�-�aVEĩk0����8?�6B9N.) ��-U�P3DC�x�<1�JRR������*ʔSD�Gt�<���1..�攪=*͚#fXl���0=i�FS��Ő 
C#bLѠl]�<!%m͒0؜�qG���H��&��<�U5u�V��'�W�3��,+0cC�<�񠅙A$1yt��*����2�^B�<�"�F�9��$���H�=K!y�B��+)��b��[�B�����gH \94B�ɫE�[���=��T{㏊0l���?�<�tL	e��J���F��ȓ�t����
s匝���ӒQ�>!�ȓ<(t� ùJ������7"؅�,+����'x<Aj��E�m��IR�'z@�PG`V'L��T����LpB
�'f�XB�ln���`���5<@���'�@*�aп<0R`�0�8�����'�j��[S8|S�l�2�� ��'��|�u�M++Xǡ,)��
�''j�H�抯3t⬢��W�P2}��'*�3B���kV�I4rN>�L>���)H �J`�Ć��~���+�!�ď�T�Fy�i��D��,�R�I�M�!򄈃F����V<m����:�!�
3�<��DN;T�<y�#��+�!���ڬ���@�$F���u�4`�!�D�V,Ҷ(${��9�ӽ0�!�D�[�B�)RL.A��S�l�X�!�D@0�@3w V.	44`�Yw�!�dT���UЊS�����B�2W��$�"~P*�Sh���JU/�ĕ���� �y��ŋHO�tkç��,A)��O	��y�ɷ�����`ƻ(I M{")C �y���mB�37�Z�id`���։�y
� xd�ց[�|�wk��cf"Oe!�"K�m@�9��РRQ*dqQ"O��U(ּ�go�}3� �%V���	f�S�O1��QhʩM�&�cG�E�)����	�'̝b�N�.��8w-�
L}"i�	�'�|!	��~9x��$S	�'�L�z�+Q0���2������W��y�.�9ȩ(�jF�#r�M�GMQ��yBM��}��Q�(����s�/^!�yRd� ���S刻g��`���:���hOq����q�ja����"E#4�axc"O&��D@=ɸ�K�ᔟp��A"O��A!Hٕ>�)K�K�#���X"O�y�s M�;��� ��E�F���A%"O��k�O�*S��8q���O�ƭ��'��8���)(��ԁ'��Q�4Y�zC�IM��B��+i��R�)��f�F�O���ɸ��yya�+'2���"�>j!��>���h�]�p�D!��yJ!�DXh��7Fʭ���W
�!?+!�d\���p��J�F^���	��`!�C/^B��t��? >��T�_�q!��~�Z��Ƨ`��䲦�ih��y��R�r�ޔ��C�y&��s�*K����(�OL\ �F�r���.�'(C1��"O���2U66 �"&�$���"O��qF�&R���`QA�`����Q"O�]s�"��=��[dj�c���f"O>A��BqI�Vʆ�Pr4"O�q��;L)Q���3^��C"O���@�#c���F�ԗxh��R"O��+�Ǒ+kМ�%^�N\�HҀ"O�!00H�at�[���3PY����"O�-p��T�{�܁(ԍ\�]���"OT�R�)z\�|����4���Q"O&��W�ɬ5��|�r�"���"O�qp�i�U< �#G�C�L��5"O���!�
#�jQx���<N��Hi��d3LO�H[�cYh��
��['7����p"O=����*e�ݺC��i��  "Oҽ�����g��`�D	�t�D�E"O��2%@�H�q�sH�2�*@�F"O����()���2��'&x� �"O�����nπ-t�Yc���>�yb܃����ԥT9sWߺ�y��W ���b�ʕG����'�ۙ�y��>�ZT`D��(���H0���y��k�)Rj\�S唽1f��y�A8B��� �ѧTm�4{���yf
4��BǑI%H9�b@��y��cm�@ F��H�����3�yҤ
'��9!������B����yB#�"~��@���^�'0�Jvĝ����"�O�HQ$�*-'���f��
P�nMc"O|a�'F�,WGV�z�b�=Ĕ��"OF����Q?Wt�*� �^*�;E"O�1�W�h-�Ay��g��P!A"O~�
���?g���4������"O�t�pJ3b�$-���®;�0���"O��C��2Ud!zeɇ�C�P8�"O(�ca�n�[閒#��x&"OJ娀".D�fd��Cqbe��"O|	������*����ePQ"O����[��8�A����\��G{��� ,��"Ue1�p!�]�O;�8��"O^�:Aj��r��r冝�
*Qj�"O�
�%�K����O`�Ȼ0"O�;T�T�m�D��5o�2!�zк�"O�����f�Z��bN
�4X�s#"O���F�;"�J�[`�ߞ[rj� "O�uh�Ղ]%$�Jt��4�bM���'�R��'�Hm(��)�F��p��9�b��ȓ,8�u���ƺaѮ�f�3�J��l*Yʖ�1
����lӚ}��Y�ȓf�hز�GJ>U.��&���ȓg�A{�ʛ�I�8�o�VxI�ȓ{�H�I�;T�^�ˀ��r&�,����ջS��wώ�VIF/9&��r������9�L�5�<�!i��x�v� e� D�x���՝ƭH�c�-RNfeX�%�<A���zBKM�=xR5R6�Îb\���o���j`�T�$�:tn�̊��}��;��:�������kH`����>��Qpr�	\J,��,�9-xν�ȓ;�(Ԓ�	�$t��%U2E`��ȓ�(��qa\#G�a��F
fQ�T�ȓ!���&ŚM#�xBu�ܿ^�$�ȓ��=p�S? b�`2��9AxY�ȓ-.BhCR��=㖵��X5X��ȓJt�K��Хad�1zSjЄ�Z�$[�`U�f�L����.-L옄ȓ]7�����$q.^�a3ᑤD%���37����m�	Yf5�d#�!#��ȓ
y���`ŋ�7Pv��ե�\6*���}�j�(0	P�� �G�5�t��~�)��� �k��Ԓ��;�H}�ȓv����ف1$j����k���� Z�L�5�*w��%:���3"X���Sb0���7� ��I%-�r�Dr�ӻb����l�?X����@��|VB�I (N��U&���ikG�0�C�	�Z��r�3���R�Ȥ}��C�I)5=x;e �b�f�3#�)}�bB��o�8�Ю��00���M@B䉵$s���PgB��F�o��'�B�I�d�ȡS�A�'g��%An¢=i������!ӧ��v���x��bd� �"OfH�2->#*2�a$��+�%#C��y2���e�6���HA$쐑�yR	�cD,�Kَ|���w�.�y�hӤ~p����0o󲨺fM���y��H-�-0W�ȪnM�LN��yr� �b�8���-�=M��ұ �������hO��Z�+)pP`�f�׿N` %�s0D���ǉ�2Dh �P�	v^��g�<و�哼[�@Ly#���g���[ !U�p�TC�	�_�4� ���6��<|4BC䉚7m��̟�e,j\%ҍ�vC� RZ`C	�G6���ʄ9ϢB�Ƀ'���rŅ�`m�D�Di2�$��?����ğ7Zҡ�L�o�hD��Q�!�U$�T�5�Ǖ2J��BЅ <��I����	[�)�'b�vL���&��0�G�ˏ�5��b}(UBA�<U鈙J'�
�����*�H�	�S�N�c����ԍ�ȓ?��Ā��A�E �P����0N����DTj�qr$�/a���ۅ�U���p�'����wf塣�\�_��@��(8]|C�)� P�PG�DW�1��)��1b5���'\ў"~�^�4}���%@<>E�D�
��y�/�r�<Yt@�(��)���#�y��8��bE�0���Xf���y��K�O�`�A�q�D���y�Ï�$O��s!⍎t2V�х�
�y�#Μ`D�8 ���oj�A�c*Н�y�?eC�C�C�d�L���ϐ5��D5�S�O�\�"u�\'��9�U
؆�r���'�N�+���<���(��N�#n���':�#�ɰY��L�����
�'��I�2d�,c��,>n&�q�'M�U�ǣԈ$.�De�N�9�aK�'$���!�V�
���Һ���'��pϘ=&P�����F�kZ� �'Ԭ�ie�Z<�z�X��k�f��'%�`r�1!?5P�� �Z�����'q�R(Z ��҄o��<lj�{�'���ITD63 ���Ԥ�+��i�'�Z�x>��!�����([�'�x Y�@_�[��;�A��^�h��'�6H�PЎ���Cq+D8i�`���'\��9AEʄCa�tp��P�6N� ��'m������c���cA��_�y�'0Z	p5�H�l�H�{`O<%��yH�'w\JPO��3��A����!V|��'֔�C`�Ė5��B�Û a�!;�'�����e��C�J\ID��%��UЌ�>O��X�
��_���s���&3��8�"O���"'C�Q� ���@�6Q� ��~��P�s��܊}��ΐ
�<9��^1�iM�}���
��X�e�8�ȓ(��CMG=`���zd�>Qۀp��"�2p��hr���R�M� |�ȓZ�4�مŉQ(PYr�IԸ�ꝗ'p�	b�)�Oz-�#�E!}�D�3��I�� "O-��P�ak�8���K�i��a�g"O��ٔ)�o�F���K��jA�"O��ঋ
6�����\��T�D"O�(�0d �c!�<y +�6D�
��b"O�H��� ]��L���qpX��"O8�&�ŧ�b��w6�x��|�]��G��'[~�0f#�!`� J��R�#�p��'p$�z�e�%�b�cqV=-�N���'Z �yB@�)68 t�`h3y#�-��'0�u��@G�}�H�_����'�2pXU�Ii���Na2��'|�<(b��
p�:���G�L���'�
� $���<qr��,V�Tx*O��=E�D"��d��)qf�6��l����2�y��VM���%aU�3����ӟ�yB�T��v�G81��l J��y2Μ�
A\$ۥ'ӟ=���T�ܦ�yRE�Poj����I�t� ����ڵ�y� �Xx�Q $�lk��(a�͵�y�b.W����N�dH`�(M��?я��v��<8D)��U���d<=�*���,y�R˛�Ⱥp�M�\�܅ȓHi��iٙ���ʁ�I0��y�$%��>R|��D��E��I�ȓ1-`�b0o�|��!CF\�;��Ѕ����F/�+��s�[Hw	��8�L��"R�J�e�W&��j�a��8n
�CQ��1fD��b��4��'tr��3� �A;pm��>�6`d�T�	�"O�˱O]�b���[ր�4hK>���"O��jƬ�CJzāe��GW\;�"OZxpFB�i�H!�3dE�H����"O2$�nճP�����Zv@��"ONY�P�ήTQÓ�� Q�
h�"O��w��1n�2�! ���́�C_��F{��ɚ��4��띟I��aD�G
m�!�Iz�D��+	\���+���'d�!�DP�9�k����.�4�p���N�!��}D� 0�ׯ26\�`j��!��228��+F�P'��x��hY��!��ў<:��   5d�W"�(�!�� p�T#TDO-u��e�1Z���'b�O�#>�&�
�F�.�i"�ī`\{�l�S�<�*1}.�"4� ��I3� �K�<���w0᱅�ei>�2T	�M�<�GC�)�p��G'�0�:ơ�N�<	5����� Ȁ��8sF�D���F�<� DF�,9R*玌�)uH�rƥi�<��� �E�����B� �AP#��hx���'��A��*K�X0h �${T�m��'�0�	�ÿiY��"/���b�2D��JU,O+:HT9����W��A��%0D�J0.Ƌ5v�(����fe�Q���+D�Y�ҍFM4��"E�Y]|i�l*D�h��M!&�HC��N<��Y��#D�L+6(מU��I�FF��jR$!�D(���'(��b�ݥ�H5 3��+����'��eɤ.�!���[��9(��'l8���晍`}���&	�Ԝ�'$��se[�0H�uCQ�(��ڷ�y��?M�JW$���`xG����yR��=T��L	s�#���W A&��'�az�ă16��*��9F�b�Ai���GxR��??�t��D�\�f�&�J6�P"�y��ŻGK
T�A�#X|�-딎L5�y2�Nk"�,X0Y#X���c�� �yr�M� ��][Ą�]	�d�夀��y2߾a5�ȁv���MP� �F��<��?ٚ'[�ٛ��)�lez�@��^�����=��y�ذ5&�t("` �7�hURfI�7�hO����A�'+�8����-J�Ti�-%B6!�D��
9$%�^@�Xr��Y�G!�$��b��%.�N1����(ڦ !�D©=^�E����@�xT��?f�!�$�F�B"��A� �'$��}R��81"�>�I��܅/�.���9��b�����>O�i6M�!oyY�7�Ո�R�.9��q��M-z���������y""��R�u�GҸ
(��	Y�y���`���۴Ag8�sM�(�y$�0$T�@\6O\�ˁeΫ�y�Ό5P�v���/���c��y�nM�3����P` � UF���yR�L�JҤy�ѩ.�MS�g �y��3-
 i1��#d�c��_����hOq���Sw����,�q���s�H��0"O
�!W!�1?A��,Ð}v���"O>|��Ѿf<q��KO�mv4-�P"O��#�׾Mt9�W
�yV��"O�m0$h�.�Hd�ÃA�W��`���'n1O�q���1	��B��Yr���"O6(+q&�Nt�kglF���T"O� $�Q`d�&F�S��]*��i%"O��cO�a�&��4%��d�*H��"O,������̨�3�Θ_�LX0�"O����H)T�H��a�+6���"O���$��:TM����F�ZE��"O�� PȖ�z��$ӈ^M8S"OJ��R���&�2�ȡ��v^�Ѻ�"Ol|���rl<;�.60E�I��"O�|Y�
�$&�Dq�fK�A��b�"ORa�t	@??�u�w%�0s>��"O@  ��E�nL�C�`3���1"O�p�n�?A��|��$�|H�"O��"��R�f-3s���I`�i@"O�`�%N����1vaJ�{F"O���#ūr��+P�\�`�`e�v"O�d�*�P[�m;QnB\b<��"O*1z3OB<e|[M�d{����"O6��b�/r76���,��C�0�;B�'��d��PK������/Uְʃ :?��}"����"�+@������%L \ٱ$"D��Qd���u��`M�f�=��g"D��y��D-�i���Rf��w 3D���)ٖ%T���!�H�>��K�!<D����'�Ȣ�Є��1"�?D�hx��H��0"ޣS%����>ړ�?����?1��$�κ,g"�HR��"B���:� ���y��)�,�c�L�kIr��c5�y�������H��_WF!�@�N5�yҍ\�Nm�ݚǡ��R|@���`ˎ�y��ׇ<6��
�C	`ؖ�� ���yB,ƻ={j�2šF�(Na����#�y��X�X!&�A&�86H���O\���O��`�U(�djH2c�nC�7"O�0F+M�N����N�b���;�"Orᛐ�\3�lyJ��G.���D"O��b1�W:V��B���?5��t�"O�P��E��U��&� t�"OP8j��#|ZL �A��6?h�pQ"OBu�ĪF����;Q拠0���y�A?&F� JA8.�6$���Ѝ�y���zdR�G8"���cܦ�ybCNN�!����� @�B��� �y��@1� �	��`�\�-��yn�,f��4�V�FQ>��E��yb��2��4�!��E�$xJ�y�@�4D��}0��@�T��x�Ȍ��y�̞xoм�֪O,C\yS#��y�F��s�^�[E�עQ�<��r,:�yҧ��G��QWIȄ3��e���yrҨE�I��?[�ZpYbdI��y)U�E�A�@AEvx�ΐ��y���6����E�7�&�1����y�H�5U�N�x�k�=������y��S�g%�,�� ��z����'G�y�/�'N�����Ԭ~H�4I�i���y�+u��%���ڻ��{�ŉ<�y�d�+�,m*Y�n�tq�um��y�M�ɲ��J�^Jt�УE��yb�0�J�k�]*���t"�;�y���0e�l��#D� ]h���=�y�!T���qS�$X�@`0p�(֏�y��+�< �2��9�!��4�y�mާv��U�#��wV�@�& I>�y�	+1�B�˃�ȓ#*jѩ�ʱ�y
� :��ܗ�r��Ԣ���Q��"O���	�8'0��k�K��`�Qf"O��ڶcF�ތ�H�!"Q���Q"Oะ���%�����N9�Дi"OzLA0�NA\<l��#C$/{��A"Od�ґ�&��ب`��2+�^)C�"O�H�E$�#7_��c���8m�B�"O��!�ݘx�Vj7�T,��x�"Ot�)�i^�W�`[��W��k�"Oɨ (�t��<���%���"Ob8���&Q���0-�����wY����	G���$B�	v|ZP�W�?�B�I�k�B�b�gӾ��Ļ��6l~�B�(�*�hW"8�*	
�f�:��B��0\� �Qa�K���s��x|(C��(!��"A�C�`��b����g>D���u�_:^k �n��q��Qe�1D�ɒ$�(�C �Ɔ*!��E�"D�Xa�Mg�,ɵfZ������?D��
�fM!���@&)](��9�p�!��õpL�C�-A�\�G�<tC!򄍯I��l��Ē�=��e�3�P�!���-��5�B
M
���8��7�!��6<�܋e*�#L��p/05�!�D��F�(2�bU;:�t�A1�W!S!��Ӛ+�8��Q�9�:"�Vj�!򤉁 /|����발�⁞�nr!�d��n��P�j�i���!c
\�!��L�IO�����D��"~!�T�x;�-�8�l��5�3�!�$�=7D�E����!3��i�5Jg!�-� @Nԋm�V���C5F!�
v1�r�U������aI�J7!��IX�����*��a� ��!�<_�t�c휬H�A�!�*+�!�䊧z������Mn�Hz�BQ[�!���)��M����Bk2$´�S5�!��&f=�p0%�Zx�#��'h��'��>��ᦔ�L�0Rڰ4b�K�"C�ɵG��@xs��=w��,j$�XN�&B��#!����*ҫ-�(�[�.ۏ]�HC䉖 ���0V%�<*��! �
�C��7V���e䒹By�{��j��B䉺��TЃG�gNj�����w�C�	�1mp�Z'�<-�)�蓔}<��Ot�=I�y���}�茱�N�}���ˀ0�y�M6B�h2��y���rA���y��'i4��td�0s5Fipـ!���O�4��얥 �R�y��F�x!�DԵh����#� e�:���΁,V!�ޑS~��K �ݥQ��\`�Kѕ6�!�ć;l�>���,��0��)ȟL��'wa|R
ӜJ��1���FJ��(���y�KI�[� 9�,�0?� �C��yR�]'p��Tꓴ+�~��훣�y(�"��e�<7��E�¢L,�y�%�_π�ĩ>]��B�ޙ�y2 |xZ��L�OC,Ē��F�yR@F�Q��w%�K�t1dL־�y�%?`�Ӗ"IR�<P�����y�%�rG��a,�F�
��
)�y�Jv{�,A��K12��J�%Ŋ�yRj�l̲*�˞%3Zii����y��*5�UR�L/���6��	�y
� �8��B�`Tx����Pڱ"O���%��͢%�\���@5"O4����D,��1횄lҦ��4"O �Z�n�X��q�� �x(� "O���&D3�l�Ђh��8�Ұq"O�����'4�b�_=&�����"O9��	�%B���9��\}�t��"OlhP��Īx=L���ĄEg�`x�"O�8�t�QB��CUc˲R�����"O̹���;���c�K�3Pz�% �'i��'�0:�D>r���A�؝��'�^p� �% �$�Q�;qe��'����W��1!7�yX$ЋQ��)�	�'�*)�*�(hgd�b��;RU����'2Tr!灶i�����ڏQ�y��'hX�i�D]�y؝86�Y�H/:`��'�0ḫ;�v�(F��P)�����)�Ot�y��[���N�=b�HKd"O
5a^�c-ݢ�
G�hG�[�"ON��C�[�gj1�*�MN���C�	z>	2���p.��뇂S�o^�CJ,D�P�JQ�y�beA$)Q�<�`H�TD%D��#\d]�Eh�K�0Ȏ�0PA#D���Q�ˡⰍR�Z�&�(�p-�O��d*�O�d� 
 G(h@���d��"O"};-a,���Z(U�L3�"O��F��7��rv��>g=�=��"Or�����	U���C+MOF�p��"O�1�B���$�	�\<�9��"OJ��T��V�Xh� ��	#���0"O�� A��Op6�Q�J�6a��"O��� /�!	��I���NǔYK�"O�	
a�˵5��Y�L+MLb9B�"OX��W ϲ.'v!4NXB�pѓ|��)�m)�]��hX�8��1"��_zpB�I;DA����gG!��[DE�.N4B�	=�^�YQ��'"x���D J��C�ɆP}�D[�.��;� )�@M��C�I$P�Fu�B��/{p��tjL n~�C�	>jy�Ç�+R�icgH�(�@C�	||H�q�R<8�0�#|B�2n�<�� ��q����!gLvB�I|]4������3����e �4)pB�I7N�����R��@ ��_$E�C��3��K��M�	Vʘ���[52�C�	<H$ЁN��)" ��&��N��B�I�M�M1���O����4`0`zC�I�~� �a�J��TՌ��e�dU�B�I�%:��#j�IfL%���^��C�t��49�M�*��}��S�ywjC�	�0�2�����;��yHb��p�B�	1�4�L��w��K�n
#$,�B�I�s.����d�1��a�G�8`��B�I�b隂j1�U�&@�
o��C��l��MP��V�0��%��F*�=�ç7=� xa)´&�!�ae���,�ȓC���g�]E�Ա���6;�Ň�Ht�C��8
 �mS��o�.��ȓ,ްb�	|��K�f�d�ȓ���W� ����{5b<`�̅ȓ �y�
J2Z�";�i>G�\��n��Tq!��I�V�ʣ-����v�����\xь��|2T1`'Y�o�<\�ǅ+D�t���۾A��i+'�B�&�X��t�&D�� b\�fK�E~�80��>\����"O���E��D�d�
WƷ>�.%�"O����E=r�� Eض
}]p%"O(̳Ƭ�I&D�)�.؀uIɚ�"O ���7[��`�k	b��yP�"O&Aa��S",(�2�I�
t+�Z�<�sϝ�Q6�I]|��G��X�<yvI�$Yjdp2��vT��-Y��B�	R)qKƂ�|5��yRm��0���D�ID>���R�BTC���<H6����&D��8�g��k����&ηoW���`#D����Q�0�","�/�	$�*A��?D���Vi̸8t�u�^:@��L��K>D�T���[�*��t͚���t �	7D��`3(�)B`��z���7Gh��k�)D���s��0F�m�m�|��%�'��埄��S�W���hI6ob�E�'+ח)pjB�I��¡H\�B�������b�C����i�ǭ��d3B�R�s�C�I')��EF��RE�,`�f�+i/�C��/e���fX�`m��g+ѕfw�B�I)~B�� ���yybǙb�B�	�6q���G�l���QH\a�d�=qçoܚ6E��
w�%*V����"D��R�d��``f���
-s�� ��;D��W-�"?v�h��jD�#��p���;D�<��E�	v��<�Q��.ct����-D��`�3����߆7L��2�L*D��Á���f���(ț<n�Kd,>D�����Ԟh34� ����P�X�(s�.D��X���<ˊ ��&�&:�4����!D������Cq�F�B�AL�AO!D�� �b͔'~ޕCV�B���x4!D�$b�j��I��!hVʃ5���1�M2D���vVUЄ�3���`��sQ,1D���Z�qF�=�pd��6x�hpM.D� ��-O-p��)0��Yt��L-D��2�7Eh�J��U��ku�+D�x���^9r��Ӏ׻'���@o(D�0�-�tG0*�#U&?&8��g$(D��"@l^��B��������E%D�t�#,]�K�<�*���K0�Ax��>D�He]�M�n � I�?�� q+!D���ţO'i���1qI�c�z�R6�2D�8zi�0JiB|V�̺2�v����1D�t#d�O�F)�z`_=���N=D��Y�0f�N�V����lȊ�a<D���Ԧ�$єؘ�!�a�:�!�:D�L��OަQ�[\<4�1pE9D�����']բL���]*K����  5D�*�*�b�Ͱ�ϛ;�va0��3D��نɏ�"P�e,H�C\	P0�<D�D�Aj+�J��ѭ�.c�e17O9D����k��:�lR���h1�gK6D�L mг+l��p�98nJ���H)D�H�'ڐdd���A����6 5D��Z�dC�3�u3@�gnB��v�&D�|j��Q,&uv9rQ�ÆYV��S�>D�0��DC	��<���N�a.�m{�n8D�����Ӄ+��슶G�x v�3D������p�>8���Ȑ5;`Qqm3D�4�2l�'���S�	$7$�)��#D�����q`A�l�~*�ׯ&D�� r�	/�y�6�@�p:�}��$D�� �p�ܢg7� 3;p*�J�"O����"��]"#��a�v�"O
���	L���AP�U�H�,ɓ""O�\��G�!f�jH u$�K�l ��"OhPrԠ�.i�d���G�Գ&"OA�AA�:6Z�SǨ�?��s�"Or���Ռ�&���I�>��=(A"O��
%D�;&��8���Z��"Oܥ!��<�| NŮ�$m�"O�ȁ!�J�U�^M��,O";p*���*O���l�&Dѵ*�-6��|#�'BT9��@}�ݱ 2 �J��	�'�`@�����	�w�L�g��r
�'�zq��`� ]�����3c,��	�'�1k�K�7e�����v%��'m���6��{��P \3��Cr"O����Ma�H�T��~
 K�"O�t��b����e�ve���4��"O~�yக�S�����2](�`"O8}p���� �!�9X�H-�""O2|��m7Ј��3*Q3sĄxu"OT� ��"*���	���#d��A"Of5W�Р!bj���L<Ai�x��"O��Z���g�b6�S�z���"O,��!���J,�o��yaq"OfSK�q�������/fq.P�"O��jC%�(-�EZ2�C�9����b"O(,��!	5b�<�0�䑇R�D�!U"O�upekY� 5z�`A�X+\��(��"O&造��7�V��E��b�h�#P"O�EpB*\���`)�
Z�`v"O
�2��pҔ�G�0` &"O&MrP��YG89ҏS�Mp�|�1"OV�QW&_>1�d�q�.�l����d"O��쏩,���
�/��4<Ru"O��*#%��%�"���z�"O���6(��~v@��[�����"O�Q���n���)1C��S&NAk�M,D�����A3:,h�{FO�~M�2@7D�l@�#��)���j��$6��K9D�ܸ�S��ɠb ��)����B6D��0�&^kC�}#c��A#bUc�3D��Z�ł�#�:��'*��]�0Ah�0D���t���+r�Q� �#f��-D�|���ݕ�Ta�]D�0E���8D��1-]��I%�\{L��y�D5D��:ӈէ	�.�1���?��Y�/D�Ti�*T`�F�����T.D�hKT�I�d����ˤ(���t�*D���#�U�5�VQ Bj�DP�:Ѧ(D�h)�!Z0@�(��ƓU���+BG&D��g惗|݄]v}��01d'D���D��?]�P��I�-g��h��e$D��p��W�¬Z�c���q�×7|=FB�I1-f�Ec���i�4�' .N�C�	�<��J��Ƕ&��@�3�K L�C�	=E6ik ˸Rg8Y����,f�,C䉇h�X�ҡ+�B�,EǬ�~'4C�L����M^!�4���m ��C�I�t�dMI��\�:⺼��fC9GؼC�kD>�`̛+�F�	灀<�\B�	 $8�y�D�&,6z�ä^�C�0B�Ɇjל�aw��jH�5*w��grbB�!T~�넎k�8E�?m�HB�)� �p�K�Wn��bG� ��,*�"Oz�i�Դ(��ɷ,[�X�.��"O���sd�6dG�ઑ�I�h��(�"O� 	�	KO@L�1�F�EN�xja"O���
V ��S�˛�q%^��"O�`au����@S��=$0��"O
$[���w��`��j�c|�k0"O�Lpª�#�tS��e�X�S�"O�D:D��,<l�E�+ti��"O��S!Y�Ӓİ"�@�j\���"OdĲ��֎"7f�k��X�M���"O�U����"b����S��l7���"OD!���	h�H'჉o�<""O:��g�)e�v��6�чj��U(D"O�1����Q#`�PD-(��J'"Ob��g�F�~L�"b֢$r���"O�EJС��|n|��g�P3ll"�t"O�����PhS��9nX0"O� #�JӸn�Paf_s["��"O��H�iA�Ko�D��f�PO��B"O�rIΊ�&���d"NK�m,8!�dO*]]r�I!g<�(r��[u!�D�2�*e+�<S"���qÊ�.b!�d�90�hbf�57J@�4�@�5M!�䄬&�:q�PM�e���KU�P9!�/r�V�C�eӞ(�"���	�!��:a�h6 �@Q���6�!���,�B�Cv�C%t� ��h�!�8�.$�G-Jf��c��<u!�Ğ�9FN��p�	z�)�t"�9c!�dF�N�J}H3J��h��(W, <qb!�ĝ�>�p*@,�Ύ EȘuy!�$ٱI64�P`LA�X;�0���c!�S�����l�b��9ТEAc!�+��I�ۙ/���1�%�:`:!�dP
�X7d$���bO�0p)!��^�-��̀��VRlj#n[�w!�$�2c�`է�.f���vM��~o!��2R�VIz o��+��8�4��1�!�$[ >��yjf�G.L v�`v��
q!�#$��\A7&�r�8��	ȓ}S!�d	9��`�A�S�i���̖aD!�ę-H5$!z��c�t��H�SP!�$�h��9��*�Zl�c�%�4|�!�D���d��U�D�M�?`!�dR������� �z�2r�@�E!��>k�J���b5d�����X�k�!�G1I�X�{U�%芐Bk��h�!򄍔<��+ ����r5:�i�)!�$�9Y�� �ЄY=:�J,Ҕ�[-N�!���"���T���F���֡�y�!�U�5�0����ο(��Ě�2S"!�Dg��1�J0h��-S d!�d�5?LFb��P>��Pg�kT!�D�$9��y 0R|������-cM!�GV��@��O�
�z0�|2!�	� ��B':��[���na{B���b8����E�*�r����G�1O|���˸L�hp�*	,Zi��Z�_�!���O\!s�5�v��PE[>#/�`�"O�����\g��AtI��;&�2��4G{��	D4KQ'��2�@?�0P�	�'\�ȁ0Z'���
��^}��yR�'U� p�OZU��Aʃ�
�Ȓ@��� 5a��H;6��1�A�9%6H�c�7�Ip?�~&��˶g�[e�yqA�:H��@�� .$�8�#N�66S&�ё��. ��x#��y���&�zTp%�Ģw�����^��y� �}�"M�-�$^ ��B�y�@�v,ޅ;�d�p��r�ة�~��)�'��g���>z��Q�)�XX�ȓC����P��(Y�xbg
C&6�,����aKH|\<�䛨8�q%�D{��ԧzqK�Gq.�`s�?�y���$i���ˢ�y�V���Ǖ���'��%��Ѩ�0	ӈH������3�l+D�h��^�r;��C֨W}V��3n)��?!���}�&����"�h��D�'q�!��X,�)������]z�ٛi)��hO���;��Z
n;x�Șqt���'���؂t�C� ��bd
2RLd�"�>����f�z�ˢ}٦u�*X�5�i�0Ϛ��Io��ħ<]���gi�a�$�e��1���C�)H�y���0T�� �A�T0FX�ڕ$Q��Ov�"�4�<�D�	�#0.�i��R&���&"4���%�İ��@��
�r��@֍D�<A5�n�P�I�/H.�s�$N�<��G�=mR,YF��g#��@M߹��x���m���x����L���
��F��ē��'t^��Ja�$p�(��ۡ`��j'To�<�5ꉄ���3n]�|R���&[l�<�����w���sn�m.|�U�S�<	�];4�����OwFAT&�h�<Q���g p\�4,��0P��xDI�fX��Fy��Z�s,8BA��á�L��y�ؓ��,Z�A:�U�*E����hO��ʘP ��� �0��2o�I��"O4!��+I���V[Ѿ��V��+;&!�Au���6�N�>�B閡a7!�
0kt|�k��e�B�R�,!��҈haCb�����ì8�!�d��jl�f�̴��
.R�!�DC@�q�U�,�Egֹ)�!���(�>Lx0� =B�tt,YX0��'�B����C�(ھ�!��_(,0���
�'�`�N-g����m�Oc:���'�6x�q)ϩx	�I��9;����'s��b�Չh^�iA�I1iH�0�'rR�Bԉ�8iv���#����'��� Ю��F�L�EmP��
$���d)�'m�����ն�E"��7��d���R�����*~09�i0$m���ȓ�����D�"E`h��S(�o��ȓqE�<�u��n��$+��U���ȓj��d`Y�#�)!b�޽b^��ȓ)^P��º?o>����I�&�>q�	�j�3&��j��0�a��c���ȓb��Գ��D(YlB�r�c��u�ȓ0�Re�5#�8h"~��բ�:+��чȓOR�m�UG��X^�zQ�_�&m+�'�� k�N�}�ɘw˛B~2L��'�Ή{��"�2�a���7B�l�i��ē		�!)M�EpF����>��a��hO�>9k��2F�`7�@ys��	�C^v�<��X�k�ҠS�m�1)T4x"HH�<9c�,X�[����y}�� `RH�' ��8}��>��E��⦪Փy�"�RdA6S�(��	^�IS�2aJ�I�!H��7�Ig6M�O��'j��9�~n:� !��-XG̅�����k��ਔ"ONu���R_"
q�X�PL.p"O�h[Ќ�@ ,m�!
EGl)ɔOB�REi�L�Z�r��£r��� C$}R�'Xx̀qOD�r��ڀ\�i�����'W̱Y�έt-l��LP/~��'����c!�o��x�@R]���RM>��'ț��i>�	F�i�E�х�	�=८C�#�d(TO;�$"�4,��w@���� X�VI(Q�'Oў"}�c�Ƅ3��E*��No�R�B���8_ў��G<�(O��Yw�]<��-3Q�@�v�B4�>�d��O.�� �NJ�"s���q
AjQ8�aB}�x�I�F-���E��s�=�OP�DY���A<�n!+QI�St�l��I@�'��*�OX]f6Q*ƨW�����'kZ�0!ǹ@t2�е��~���J<��4�O���3���2��I
��z���"O���r�0	J�a�5�`��p�D(O
��b�쵋P��>]��0��
a!�',�h@�"�)T+���˞n�!�$L�{�޸���!�irQ��(��z���K�+a>�
G*�6t9@ɘa�!�>��}p��4���D�`I!�d�^�I��|s��0�DG-
S!�dQ�����Æ��� 2��*ga�2>O�干o���(qA�GL=�U��"O6��*\�G�Z�kJF��`��It�O0�iӰʐ> C���l#�⸠�'�R�)`��5��"/�; �D<A�'����g��l�81�ÒH
�Y�'.�� � ����H�"J;��+�2�I{�dÏf�T�BJ<]��A�4M\9@����f���ZB.{��H`S�O7�a��	Z�O�n1�NB�
�4TS��m�2�����:d"|�%N�Q1$8�G-$
sǫ@�<���$%f�jgn���T�A�+�VC����]�,��qf�;7�B�	�N�s����gkB�k&">���iT7;b@9)E�����Y��X�y!�䔵���C�A�pXb�`ԩ��T�'{1O~">r�%yp� �c̋l�8:ul)�h��
g@���MT�)1�H�I��&z\�I3m���Dy�O1OX`�P�Ǻ'�X���$��cW��Q��D�d�>	C����3��D�؅1��Y	h�,����|r�]��(O1�`|@5�T�fFD�0��'vݺ��?Q���\:/+\`#ʛ-h'th�hO!d�!��P*�0T��<T	b$J� ��	-<6�<Οɧu�kٱ)�\l� (��Ô+�/��i�v��a������;`�Iġ�>�-OR�=�;{��0�e��>kb�'H�3`�T�Ɠ.�}��@2�3�E$l�:<��y�ͅb���O��:���GG8�0T юg�6�`
ӓ��'���q W�1ڎ�%C�*5>�x
�'���A\�\�,�I��@	C��	�'cN��%ۈ����ga�:x,��'�XE�/+��1�F�/n�@���'�D�*ハ�J�As!�_!X 69X
�'��E��Sk� `q�X? T��'��eB�jڋqb��*$h8׾mb�'��Q�� /v�|7
H+>�*=�"O0$�u`�1P�U;�-�/D
$��0"O����-D�"��A�!��E˨�:6"O4�c*��Hm���%���z��"OP`�0�^�o��	Rp�T��5��"O� �x���al>�J��Զ�1�"O�=�S�K( ��(k@��?F`�"O�e�ܯ �R�j3`�

��p�"O�@[%��n�tX���AU��"Or:7���Nђe�C!�;7��6"O��4�5aB���S5��"O6�P�B��KԈ��э_/�"ORK3l�9�=�r��!*��u��"O�ܻ�i�/�D���N�H�lm��"O��2&�C�+���`A��_�*P*�"O� ��&Z!Đ�Y��^�a�"O�(cҨ̺�h���S��`Xj�"O�H'#q2��� �*N�xĉw"O@�+��Y���*WO߀�6ݩ "O"��� �06ld���>@2"O\��0d��$���K\�6�RQ�a"OX��Aع4.<���z��6"O���� G���("��8�: ��"O���W)�=��p҃H_06e�(B�"ON��!&]�H&C��"sXa�C"Ob�����l�F�6�E��@"O~��!�Oh�2$Xba��s�N���"O^	 �ؚh}�q ��Y��L*#"O�Mr�1$"�h&�\$�8�� "O�5h��+/ @r��,K����7"O5�S�y���cr�@�6�|;�"O��6�ɟ0tPr䈉��2}X "O8���k��JH�Xj2�CV����"Ozp��"��+������	u���b�'x~H�!c<�|�{0�*H��b��?��u��'Sv�Ya���T�q'�����'�I�DnZ�,�F��j���H�'n�@ ��>)��9m��rD*��'�0�PF�>f:���GLl���@�'r���E�rl���ցo ��'�
��נ)
���sf� Q=���'���@C�r��\#��R�Ue^h8�'t����/{�ft�j݈L{��+�'ɾ�ʥ�\(T�RY�G�I���	�' ��D�L>= �1��!F���s�'E0����� T��510��kr�� �'7R@��(��v|�1�#��R��'r\�*B�Q�u�̑H�.D��'�4!i��Y-#�D-�v��	n���'F�$�-M�)��&!��hr
�'-8 +`��i0$��5�4etR�'�%�$��z��ܙ��	�T�$��'�(!���*\g�%���2C�}��'�#򣃢�d�д1N�e��'��i[@"�,q�(��蛖ZH����~ƈd3��	A��(����F�(��f�l�s@o̢m^.�	�k�+�b���+0*�+�͇�O(��ܟ�����T�DK'�F%V��p��t��y��L�S�$x=Jx��A�U!��-��\��û6�E�'MZ-`�����(*��R\�><�tA�8Ɔ݅�UG�I�����J�"�0O{(����*�1�nͷB(^�@`	q��}��|�&-���&�0���^L}X��Cr�=
�e :x\P �B�V� ��q��D�f�޽??*��%FҼ6�l��ȓO�(�!���R�r��v׾x��хȓn�~��0-ʹ�ҕ���L�q����S�? ���I��B~�}�"���d��"Oʕ7��;�5���@Ǭh��"O�q��˚|7�9��f����%"O��)7��|��R�)5O�>P�@"O.�x��\pu���ԩHS�05"O䡺���=.�l��'�!)��#�"OV� w�Lx`�����z��5k"Op��E@�<r@в�e�,5��ɇ"O��ȶgL�S�H��G��P��a@"O�Ms�F�-L��h�5]����"O�TQ��2o~L94&R2f�ļ��"O�����.FbA
�%�!hẼ��"O(ݒ�a��i^1�7��3(�x �w"O����%h�*����@ތѣ�"O|��H� 	(�DA��ӛ=�X�c"O�uA)jV�1:C,T�����"O��Ӷ'U!��|�᜛B���&"O(��Qbh�j^�d�����"Ó M7����L�!J�hH�'�vAI�N[S�����)>��Q8�'^(�x&/V9g��k hDI�X�	�'ܮt����Z.dT��#-�Hy	�'�ri�f͑�O,��ƪ����@p�'�
��e;���Jvn��KD}��'Dp+Aj��j�V��(�M����'�� ��BJ�Z�䡘��T�w\̈R�' �5����FaƘ{�+	;kU6	�'�ؑ�m���cpm�m���2	�'^����Jl̩�2�Xm� =)�'�h��8�*�i̦7h�k�'#f,���ڲi���ajQ�>�u��'{�l���B�K�n]��������'W��Z`�	76����P�"��'�x��ʉWҐ�td�=Ft5��'����� ��S�*ɋ#���'&6Dj띡��!cdǈ�����'�0d���`i
��� �9b���'�J�`�&K1*c�!�`�/L�PP��'�áBK(MR���ە;�
�!�'�9���-F��9g�������'���R��l�y�F���6$���2,���aӞQ��[P�ΰ���� A�a�F"On�kG)�JB�iCS�e>�3T�ɡk3С��Ae�O���Z2������M�/����	�'8�-c�Ǹeݬ�#�O��2�����_�4�p�c�m���)����cT5#q���uB��rlD��*D��s�ƔS�r�j®�zL�Q�3쨟�z��v+��C��'咸S��:6W^a#O�6t�	1�p��-H�D�;'���u�ݧ5�<��`jI0]���t�1D��$L��(�:	�3�5s(2�v�,=a#��.�,#|Zg"MT<��
AP&R�zGk�f�<a��}�`,ِ� ��|j��,ŉ��Ǒ� ��O?��C&)�D�	��כq'��!��C4�!�䝠bxl�U�A ner�^��$S�A�� R�듊�0=����*���L�$ "O3\]���$�k�~i��EE3UZ2���^�0~�����&w':l)�'d�Ѥgi�6���ʖ}���#����7�|�+&ʧ'MȬh���u�����K�2R��0�ȓ(d�(KAe��%�<r�F�+ Ĭ�b��V2Kb�O\	� Ŕ�(�T��K0�X�B�0.�KW	�W)8B�;�e E'�� ��	 =,��3�Q�Qp��Q��\w�u剨Xm�EAJ;<����T��^
��$��c�4ɋ���y�*{P�Q��t��@��M� JQ���g�ٔƹH�	1}����(���֦C�e��=y���0�Bm�񨳟Lz�Cۙ�X�:�� p1�!���W0���W#F1�d]�s"O� �M�7S;�#���=q谝q"Mtհa��Y0#*�;�NZ�3*������y'k6|O)�DخsPL�qo��yBA͟[J�#&n[�@0D��U���e��<h,5�	�A�d�iE�XR%؋���	>�*��E�Q�T���JJ=3l�zr�T5P�&��"o��B"� �EQ%��]�����R�@��P1O����	�f|��ꅲIe�cP-��L"��8��M�$Έܰc�Q%�ej ��o�d}2a<����CG!i�f4qa-\4g����"ON9��Y#;�Vy���w�� ��'T-}�!�s�U&9���!7j�M{B-���)H'�y� W:e���h	=}S�ђ�X�y�f���H��ð��U��J�?u��X�\�>�7��*�Q�[w9�U+�	 ��x�SщaY��k��J,�����Z�^�̺`�Y��Ĵ��D,$�Z)��.̥y��\�g�@(7�@�R�����>��&ޭ���Q'��|�`���j�'�V�£ş\���'>�YA�*H��`�חv�"%.D��р�7�.i�0gԗR�Y̣<���CRXD�GI<}��)ɞ+G�0b7a�&��dZ� K	!�J��Ҥyf�s�΀ b�S wX����0��+dF�y����ɌN]F�;#�g�P�2�@0^�������P��d%Ƨ/!�Q�G�$N��] ��	S:�D��}%!���7�J{�&��w�{�E?8Y�O\p�oNE��P2u���OV6��E�0}^���eƁtz]�'+ܤ!ǥ\�|�jq�p�|�()�B�pY�A�*ַ���"�(��	!�,��Ƀ�*fp(WD�<,�B�I�8��9PR"4U�!$R�8�pt���s��U��4F*i��@͢�P&e]y�Zq[� ;{����<W���s�����dZF��2��8kC�
3Z�Н*�J��Xm ���7��8��.�h��۵���S�"X.؈��<A�/ߘ�C@΄n<�I;Q)�97(��B���?uq�62hul�"�4<���;D�t�f�.HE�Ak�;{�,��E��h/���� ��ʨ�'���Z�m�F"(�)A]��]�5��	$LL�Đ�L��KC�	=5�䪧'� V
����F�]�=ʱcK�zun- e �.,7x��%�P�1���7gVB�'�ܰF%ԺP��$t�n	��	�P��09��Oh��iƈ)b�l0:���.�+�:X�.=�eIF"@�P�����0>1����ln2(X���[.<���U��_$ �fh�Tv���F&B*�d(qÐh�ZUͧ>3�u� #��WbA!�l[�&Ѻ�ȓ:Dl��b��S~�,�Q�P%.��G)��iEG�AMb�?Cf�$?QH�B����Q��2O�v�Y�������7ʟ~�������ƋHn<�ps �%b���
ТA����$��0.�
�b��.�
=:���Jh,�0��,r�$�x d�0��r���##K ���3ړO�
QL�3G�ZeÀ�INI�D�tQ,�U��̔,T!*��l��N�*4H�хI�B�zeB�~������C��$z�1�N�23�HHl0"�.\1yz�̈G�ig�I�p�IE�ҍ3f�O�����Fۧ���xd*]9`�����5v($�$�zs�!c��$Bc�.-�8�I*O����M�z�J~�=rA�K�0=�$�*cИafD	#� �DҐJ�p�z���ئ-�b>iZ"IS/Q����#���N�b6h"���)k����J˒j�`X�A�fX�)E���#��ݘtJ�&�d`�QIB�=�����^9/���K�4�0�#	_�;R��ʋ8&�fh�1�B�8����t��%�1d?���+1�6�����>�HO��2dٱ���FOq�V�K���,M�-SČE
q�z�B�|$�g�QD�\0�`'�d. ��g���t�=A���O�M�iC-!��I� �bLY��i�*q���>1�ʵ ��(^h�ҋ[@��}�1b�Ԡ��*CxhŐF�R9b�r���J,�r$��m�<����nF{r
Y
)F�`�P%�_x�YP�C����R$N�Q�$�P��'��4y�i�l�A�B��E�������$H��qQT��. �,��F*d�jİ<Q&��!�L���РaI��#c�Z�koR!)T
�
��I�sרXs�:O\@H���"�܍mJ�4���͟P\ �<y��@)��(S���"`��\IF�n�O��HB��&n��1�И�Ƅ�"�'��]�A����Q *����r���F<f逖������\��y�#ikL��=E���=|al8����"S��U�w,\�&����Ǹb,^�|��=y��hO&���ϱ-ڦ�� �Ѩyhat�'��	�Ed�
$��hA,�JB�I��(D/���p��Q�<�oǾb�ؑQHۑr�f	��N�q�'��Ѡ��_�W�Q>�z�%�[�XE��G�<HJ0 (D�H���ڑc�f?P Q��rq���Q�;�a�{���)��$y�"U'f"H�����7�B�I�<��D�$��"4�&Tht�^�|�.B�)� l����
���AX�E=���bv"O����	7&K,}�p�IGt2�*�"O��C��K.�@Ǌ�m 2�"O�"GE(�e2�Z*TF�!�"O�pF	|L����6f��س"O�$���+�B��b��4hn
�"O�H��4�TP�&ĩELؽA"O�T)��Hx�o�#<0j�kQ"O��FH�u�|A�J�J#�;F"O �5�<$�%B#m�&{�$:�"O���˒.e��Hv��.b����"O��)��G&f~PceJ��.6����"O�8��C8<r�$�j1W*j�Yt"O�u��V�4�0���j�E"Orh{�@Ф^4t����Ǐ;i��"O�P!`��%7u~����Ʌ`4����"OaA�Oߩ_|,d�7�ӈ��"OXekEh=��̀��ͯ)��t�u"O��P���k��IQ�� G��i1"Ot��5·.����)��(�pТ�"Ol����`�����6_�&9�"OV�2k `���_ҴTg"ON\� ��h�n�H�[�-���"O�MZ�̅;f����nȗ��e��"O����M��[�,둃�g����"On��`$�F���hN�B���"O�m`$F  p�r���$���4"O�A�1JQ(4�r4��J�r}PE"O���
Ξ,!��)�,��&s"O�y��¼CWTD��i�? I��"O���t��,Dh�ڱ�ϟp�+�"O��!m�"�g0%/lp*d"Oh����Z.�Ve���
�"O���'�K~,�R����zS"O��*F��v�D�'�Q� 搊f"O��#�L'$D���$*�Z�Ӣ"O��8�/.@�`��:6�8p7"OH��ł.��V�\�)6�Pcg"O��S�È	:�l��a"�<fr4�Xa"Ot����v���Cv$J��b"O��A��x�Ju�ݕ'��5J�"O�=�B���dX�!Cq��"O�-5��"H��@�6��d.D��"O<�h�
5/4��	!+�0�G"O�}��*����(��ζ ��W"O`aD��{��	�KK�x��h�"O|<�ܛ ���+g���R��i��"O�4H�;Or�B�	�ݚݰ�"Onu�S��=��ģ�� �:cڵ��"O\� e��^L���glz�"O&��aa�i�*�0(p(��W"O�ݱ2��;ț��ԮB
N�X|��"O��ز`դaQdĹ��;Ό�i"O*Q��L˳4m ȱSIŋV�ܜ�"Oh�R%�[:���P�۾i���ca"O0�s�]X(@<J#a�73a<M�"O�m�#_�^)b�{��S�{j��)T"O|1�p�r�d̉Ao�|}p��"O6hZ���hE`T��(Q�tI	"O����24���� ��9n��`D"O��"`���g�J���V�bP�8a�"O�E�3��3G ��R�JO�a��"OH+"���qzx�
��*1
D"O��y&`��BG�Q3w�8$�n���"O� \!E�,�.u�s�Łr��x�t"O�-��&k"��g�t��k�"O*a��H0
z�(3&P��p�r'"O���¡Y�����N�r<{�"O���oϥ(r������
k��L��"O`��V��i�JQ���Ϲ'����"OJ�W�b��i�W�χ]{0H
A"Oj	8 �"e�`a��6UZ��"O:ɱ�J�E��⤓>4��P"OD����ʳf�xk���>s��:�"O�(�Q�~���A����8s��iR!���
06IR6�ʻ�(<��폽,#!�$K1��K�Aӵ�:7mMs�!��hk4�H�g���{d��/]�!�ė2��q���Y��\�{ Z�b!�$Ԕ���B�b����{�� �l!�$	7���A���]v�x�-��"o!�&f�Z{��P_�X��ȟnI!�4�@2팷V���A��6!��W�0��+#DV���(��K��*�!��43�d��
�y�R��u8l�!�d� ����PL�2Qũ�'V!�d�_V�,�R�� ����x�!�D%4ӊ��¾`���g��!򄙓" N(���4	ug���!�,���mS
�4j�i��!�D�R�}y�!�MZSM<6y!��R]pJ1D{�z��4iT'!�@��0y��M��hD�X!�W�*�*%�+T)84�Qh��:7!�䌸\�� bq�-?����$����"O�)3GtH�a$[�1�D��"O�|��� ]�����:7�:���"OX��f��xN^HЗ)�M��Pp�"O.(Ic�Y�+�D��hF�>����"O�P{@K��y\�YK��Q�Н��"O �Z�&P9@>D2��P�<ޘ	k�"O�u9kK�9q��RP���-2P"O�9�d����8��Q�_y���"O��R���=
�+f�)Kc�@��"O�I��.�v� �Fy[��H6"O�Ͱ��F�R7�|3)I���"O���샴RL]���H������"OpՃ���r�t۶�H�a����p"Oġ���α[�t��K�90�Z9���'�^1��\ʦ�C�˃�3[`�����G�`�9� D��3�
�r҆`�RU�N!�Y�� �f��Y Ϲ�(����+��DܴP!dJ�{,�\��"O���B��#y�;#m�/f���R���.�d	���2��S��?Q�S!M���3I�m�0�##q�<�5�U�Z���k&O�6O�q%��s?Y�^1| ,�Ib�(LOr����-'vI��ʂ:\RJ1�'�'�zUyH�����r��;��*D��5�Q�UC�\�<	�`ô����s,�1-�ٳ���Z�'�d�Yp�·���G�䊁�N���r�	�����E��y��^�P�!8Չ�Dh`��(�2u��U����H�"~��F+�I��EB!p��"De�rC�I<G� ]��+�.h���2�AK�o�t���]Wdi��0XazR�΅h��XC#R�m��#��2�p>Q`/��|�>��Sڗ`��Z�l�#wLh!��ٖLdC�I�~&L�c,C�zS�� �,bV"=y�"	�=.�9��Ɋ<��͑.�|j2��'FX23�!�$��zzP�X�f�aX�"�o;u�V���G��$n"��|�ܡӵ�$�'�y7jR�j��P�v�2�: � %�y
� ��+0
O(2]d���`p�J� ����ѢS������#���(Od��5�5ߺ��FČ>p��Hh��'`���<-�m�&������t�p(	1��g�|a�(�0j�x�O�R�P��d�gH�}��OQ�BȠ9�'��!fV��Rg��&)��>F	��$9���kă/�f]���´*>��"��2�yb�<v6�Lˣ�q���+��_t��/g��ѓ�Mr�"��8O��}��}�!�u�ܵ�ŉ�Ly8z0���!�-!V��h`,^}yL5Ra�;b���B҅���������#�t�v���#Q���ɖj���  ��5/��:6$�9Yb������=)���YY�=Z�(A������5fX����Nɢ]�<Cp)�8-t�Es�WM���A�}�x��B�3-͎�=a� ��c͔܈�(ھO^�7  �IY6Lh>��c"��b`���ceB]��(D���Q�G���)'�9��,�l�±��hCֹ2 PyR��A��-��O�`�̻?��є�^0^YL���`�b���3p���a��= ��G"�#	ENaSg�;�\�s z#6ꐤ�Ǻ�΄�(O0��4Ɯ�z���eҖz�
R�'^"e���� �:���� .�d��#��+�8��f�1�2�F�o8�����[��P�*��U?�M��D' 4�?a���	�Bݐv	:�I��<�Ji ��;A��"D��$!�L�P���ZWf�6u��.�  ��	�P���Ad F�I�S�O�>p�UfS��V�p`���vG�Dr�'8����!�(wܣ��j.�p��|�h+�`���y��J�Fi��`� ����q� �Pxr��#42���>4�jm�E�Lt�V0�`c�I<��^)��N"����ɝ���*D65b�f���`�/��y�ȓEƄ"�l�M�( �$dV�SY���ȓ|�dM��[�{b��+���x���NY����Ӽ老as,�Sz1��v�%"%mBn؈�p	�y�@���:4�q �"�|I��_�o8�P�	�$%" �'�.1
�&ߏ1�$t�!��= ���.7�M�� ��~"�P�]X:�a��U����h�b�1�y���s �4��2��@:S�7��'w$��3c�n@��G��&V4b��-@����LM�ub�)�yb�ߧ:>.��	H.x �e�H�U�c#���	�:*Q>˓_�J�)q
���=f�ӡiW����ɝO��U��2Od�! b��y�a��'��CJ0��B�� '2��W�=xa|����$�R�B�#
Zv:\�C�Oy���I>'K��ɔ��D��L�8
�L7	���95�:UH �A�tx4��'���!�KP.7�������cǆI����a�
�ZSo�O�,��r���1���>�t����V8?0�`�O׮i����@�'W�I0�㞞g_V��bM7R-��$	�|��ir%��,��Dcu��sJ���X���"��5V%��!�D)�DDEW���C�@%.(z�bj���=a"�#)�@ȩ���9��P%'n6�ó2I	���6�%YM5>�88;��Q�IV$Y� '5�\�K�8X�F!�S�N!��h$cM�~��]�qJ� �6D2�kJɾp�,6¡u�؊������T.߄�.���5�a�S�����D�x�%`U�+|h3-O�z�mVV⠒�qO�D��b���±�`�NSVA�É�/'~H�N�b@�de�p;�@ͧ�Α%�<��%�z{b!JvA���ro�<��Y�g�g��򤞻rh5�Pώ�qF.9����8��ۥa�	�,�4&[^�A�Ý�{�0��c�HJ��r6�	�W���� �lj��+�'3���z������484�O�1����5�i���J��P��ԭ��txQ�It�n�[S�L J���0�&���q���:2�ДQ��]��?Y%�ͻnG�]:��7<��qt�ئ�Q��	�M��Ȧ�'���1��̚v�Q>�ػp`ɤ�O�C�~Ec�B�7\��C�G�M��j�V�E�8��?�=���E؞0���hÄ��ƣB+�49I��I"(ٶ�Ƚ�y�OM��I� �����#HFִ8���
G�CR�� ��R"̉fA�P��'A�=�E��Ȇ,K�LN#� Cc��p$�a/|�(Gx"�`ŀ��Ңğgo��G΄p���U;�0U9���$sC<�{�#O�hO�}P��,NW"|��MP:�Z�����;w7B0�/Ĭ	���`.T��['�D�<�@�F��K�L���H<r��뵂ĨF`�Γ
j�̓g9�)�'ZGf�۵	%�B];�+��O+�e�'��)2lU�g�Z�ꔢ@`F{bj��:����mH;���w"�p>�6�^�rG�N��:����,or}C�R
%�B�ɹ;4��2A�7"�V{&��'�"=)@f��t
l���� ��3��أw��)����ǰ]�V"OdUj��1�4в����R����'�s�Cm�S�O�@C�@�M�����A�l�R��"O��z��͠C���g��XF"OJ 
��E2@60�5	��Zq��c"O�XA�VY��@3I��$�4"O�}��� �56�Q���,����"Ol�8�۳\�*qb!�{�I�"O�h#�%�)f�pEY��;,�6`��"O�����&�h�� \)U��<��"O��!$�P�֩x��7h�*䐠"OV�y�iP<q�꽻��[�a�(���"O�ѱ�`��r���o�9}8ja�"O�`+�h
<mݮM"A��:E�p�K"O4Q��Y����Ic��}SP���"O8i3�O��Ca� �� V�)M$�Y�"Of	[�GH<M:F<���.z2��t"O�0�2$y0���4Z�$�$�S"O�0�� ��.0\�ʷ��>���"OiK�BW6be(y"��Y�Cׄ��"O~m���Еh��8kA�Ə$�bL�"O�Uq����yia�
�"��Iz�"O 4��凡Jؤi��X�(� 岥"O$a��a��48�����G�Mr���"Or��dU������z{^�T"O���@�fP<%��8���ZB"O����ܲ1�.Ę���/G+͐b�<�B�`qSŘ%�)��]�<1ѪL��Xyp��$`(Q�C�U�<9���n,ʉ�2-�#�x0� P�<i�(�Q�dȂ�� g�p�5"�N�<A����!����6K�	 ���H�<!�H�D��y����>~*��gUD�<ɕA��y�h�#��K�7 �YC3�DF�<���Q�i��� o��Q�W|�<�#�͞���,M��F�3���<��#��#C1{�
	db䃃)�v�����Z��� ��;Px5JaD��@	&�R�)#D��i�l�*�.���,�}���a�>D�x��� �9$���딪'���O<D�� �ޚ~,T�'��8.�hC�(D��K )I�G'&�#�F����`!'D�p�WO[�pW�1)�3,E~��1�&D��G_&Hr�PJ@+��|��C�	�2��%"�*�5P>.��,�2��C�	��h�go��a�8����Y7�C�ɻa�nѫ�NH�d�6`�RE*f���r�yN���B�^ P��,.�~!l�6�Z��' �K�)�m��;��������L�T��F��>c^�t��yR�O�����ݚn��Tc�GʰS>t��pO�o�S?v���'NLC'.Ȯ!�x������4U$����(�"�6QD�����gښ?��b�T2?���3L��~�P��]�a��m���C�>���X�o�P-3@��8��p0�C�Py�Dف2����I�(	Lk%P����Ƶ0��OȴP��OF(���'��TZ�fcaAc��Ē'LR8Ù'l�9fq�(q�T��}R�)ڪtzp��F�!�0�0�Ϝ���Bw��O�Z����	51lIX�`�A6е��dQ,�T��D�EF���1n�}��Rs  �,�ee��(򫐃{@.Q8/O��Y2��/B�b>%�,M�I3�T�o��^�D!@RyBm ?u�xEQ�����@���O�v�ߢ�
XB��_o���JR�v6�)�����t������ ;�&�cg�~�)�)�'�0��䃶��ytD˾3�py"aLӟl�MQ�?1�YB���Q�2��ԋZ.u��͠`AN�t��O*\��O�r��Bc�a�A*�o�'JD��'��E�cG�r���GB�*!}��:��� �8b��~�zQ�b�L$f>�q8�"Oyb$�����q��D�D �kb"O�����Й��(���ܲ(.�1"O)S�˞�q�Uт�$=6>!��"O��S"�N6G���;C�3�Y�c"OB<k��������-�@��aÇ"O̅KT!��A*�īZ8v+�"O6Y�����i�D\�:rNi��"O$�&�P^�X�7%U�m��"O�Q�C��a)���'EFh���"O����)�p(ر
ڱS4 ��"O0��wʈ�7{TH�F��0{�\r�"O�h�A�(}�n�cg+G <�t��"O�(H��?A�H5p�*�"X�TӲ"O<�)c��9+�(�7H�.u���"O<��2`T�|A֭��ȣ.�6�R�"O(x�fG6AlyڵmX��x�1u"O�:��	>�@,�+U _.���"O�H����C�R@��k� ��K�"O"0
�i��]o��)_d��;"OQ�
ݚ/U�h�w�H�UV��	�"O� x����
|��SV�<AX0K�*O2p��#V��$l�a��c~<	�'�m�b���B��S/]U�!��'\vS0M}}�$ʃB�+X���	�'O�yQ�R5\tx��Q�����'�`�[���y��:���!��h+�'z�� �/C<^p��
��A�q#�'�tıe)U�@�2�4c!C��X�'�6�aef���%
̦B����nT�<!a!���U���	 m�	���P�<�sÜ%4��,����	`��X(4IO�<��kX�s�](#�0n��s@D�s�<�1�!6� h2 �c�d�X"`u�<�1噢UD�Qn��"�I8�b�W�<Y�@ (c�ڄ���F�"����V�<�q�K�8�����(�~�c�˛T�<��	���!;��:@�����GT�< ��2#u,���V"�^D[��L�<� ݧ�9 U��zF��b��a�<Qsϓ�q2��"��r���۷)�B�<Yf�B��&��#�n��\���x�<٧,ʦyΈ�j��C�K��!Nu�<�B-�%��:V�@3[��B�B�|�<�4�ĒG�XtX�iQ�� `�N~�<y�S_��U��J���X8rO[C�<�PO�E��
'��:�6Yc7#M~�<��� �WdB��#$C���t�_}�<� �?@QP1p��P�oJeo�c�<�5��2|��S�-^�$$�a�E�<aע�q������Ҋf-*|�6- A�<�R�Öl���z$�Ų$V���e�W�<ݫYp��鶧AUnz	�'�o�<�4��\��SW��.P��"G�D�<Qc��
a��P[��5MHA!t�\A�<��ʅ^5.!H��

\���b�UX�<�D��.�����d�'�V�+E��U�<���ć��{�Vv,��B�w�<����'
��T`�:.�R�J�j�q�<�R*���%z��3+���j�i�<�� ��|AΡ"ЄE�Q pA�F�J�<�� }y�(���%7*x�A�M^�<��ˍ*gx�xD�Δ2R�y�4�J[�<ɢBP?I'�k2�	D)�"�FX�<� 6�gh͎x����@����"O�|Z4�	�j��[� 
&%��<(e"O��"o�6a@)3c �7k��!2"O&�rTl���V�t��fx� "OZ0SF#�T�t(H���|�|���"Ol(���*`��@���`��"ONѣ�+J
>�� ʥ�%�@��"O���Ӧ�<��xڀ�ң�
$�"OD���Ə 3�D���?{f"OlpɁA�3u) �4�H�t���F"O�Тl����%d�C��"OR� 4jYK�DX�u�	F��D� "O��xՆ�	+���K����W
��"OR�
3χ�(l��a�N_73h��sp"Oؠr�\�ˆP�tM�72t���F"O��e��n��| T��.XKP���"O�H�#�0�b��@H:��&"O�!+�UOu�W(q"O�TE?@�e��.A:y)���t"O`�!� ^��f�A���R(Tj#"O�Xa��K��9����>�
�`�"OL�ڂϨz�q肨�(:��H0�"O�Q:�dP>P���b]�Y�3���Pyb�B#|����4	� B��L�<Yă�>%2�*���t�$%��+�G�<Q5��-���-��:�f��`M�@�<qR��:6�� @�����+�g�<�����>���Ⱦ&��`CoVY�<y�ə�>�F�ڦ��4$<�9�H�\�<g������򌇶r�\q��iTt�<��8\�H���핈UF��F�o�<�5C�&и}�U&A��^���A�A�<Q���UO��!�^&$R��Da�h�<���U�0�Ccǉ�W�5Ba�H�<�����	\h��fD�!P�r��Tz�<@Viݜ ��d�ty��R�EN�<����)ʅ��B�=$p���K]F�<��ۏQ�n�&�E!JZ�`R����<����-b�,��Iʵ}>�b�iEU�<id��\$*���zu���gf�Y�<��e�cժ���$�c��E�U�<�0���vp��K G^� u��D̈Y�<��dO�p�zQ6��\�`��,|�<1���)PJ�	��
� ��m fKz�<	�;D�n�x$ƛ�7�m��v�<A ��
	 y ��$�����o�<y"痣�D��5��l��F�T�<y���k:8��dQ�`8�r���k�<٠�E+���Q���<P�J���GQ�<!Ĉۼ%l4�º2H�<���r�<Y�Y+LH�ۅǋ�lj��3rD�n�<�I�vfȍ��+��k��ŋĈh�<b�Z}���#�x0)��m�<�NN(8m�!b}	�9)2��j�<�A�����4�%A��yX��^�<��*���mҶ�V%~��q�b�D�<9w�WM�N]S#)�*�|哓D�<)��\�g/6t�ѝdZ
�;w̅�<I��V
	B<d�A�J�v1�Ӆ
d�<��Ҵ/�Y;W�}X0c�"L�<����a���+�$��$�:կ�Q�<�'�!�v��&,�.�z ��X�<�eI�'iy�=QF!U9gXP��F��|�<Y4aE�p`K�+�	t$�ee^~�<� ���Br��gY1B��""O�9xqhA^�
�jC�lۦA�T"O&в.�G�\x�򀄡cɈT��"O��ze�		=�<y	r@��ޙi�"O� �cP�.F`��@��	�z5A�"O���D"ɝw��x�+��"��"O�AFER�M�r����K�\�f@r�"O¤�QI5+8�!"P[�D�w"O��X#�%H�B��C��f�"O�h��B�C� �#�&]�nu�"O�.�`񸰇İ"�&�XG萕7!�D�`�.��%�>2�F$0A!Z'^!�D�~����F�G�h�Y6�M9�!�D�$�P1���8���JV�>�!�Ē\�
�;W�ǯt��A�ЮU:�!�S��ʘc+Ր<b��p�n�t�!�<_L����1p�]�FM͍U�!�C)c
0�)K8>�
���N	!�m���r
/�<
��Z;�!��\Z0�����w����R,!�Ę >�8Q�l�G
���F�O/!�$�:�ѺweQB���*�
!��		�9�̘�������
���~����`8`����Q�LW���di�ZƄ�.�Br�#VU`1�ȓji����E��ݩ�(��&{H1�ȓ)���0��&��D���[�c!.$����$+G2.b�h�&.-�&"O���W)�<>&�����Y,���"Oh�r4���q:�⟙/�H<��"OF�R�B��D�"�pH��q�(���"Ox� #`�V��'��?H��:�"O�|�T ؿ|���3F@�8�4J@"O�iF�ߙ^�@�k�!D��r@"O�җ��MR��F�Db����"ONY���*D��
�.E=�R��r"O��Ȅ�*Z@J|JV��#f��r�"O8 c��Z%O��y��U�E�\a)�"O��(@�Y�923LR�k[bT"OZ��Q�	dY(���D�3XX�a��"O���0�l�$=V��t�G"O.Ѹ`-[6pr���$��#-���˴"O��ѡ�ۓ.���i�'M5!�^,1�"OX�S�,V��5�7fR��>�g"O 5(� ��l y���J�N���"OXH�E��.&���0-�`�'"O�q�)�Y3�P&�ӻo��"O�`��D&h��	\8Ze���p"O���R.m���;s�P,0`�1"O��AFmY�]��4�Da�D�Lp�"Ov����
���9b�0��kv"O���B!�\<@Q)R��+�*@Pw"Or0Y5�K�0��a��L�.��-��"O���0"6C�a!�*أJ���b�"Of)� I�
[��)pCD���-Ca"O�8{eF<_� 3��C(=��"O�
�I�9Z(dZ� �{*N��"OL�T�PwH|����
o9�*"O�ı�ßg��T1��?/�8+&"O����)�m8Ĉ"@�B-vt�4	�"O!����8o/2����R���3"O��B���0�e�5�7B��0�"O�Ũ�fP�<'�mQ��596��"O��C�.�.���1�F5H�q"O� |@ؗH�%4v�
�d��k2Ҹ��"Ov �Ƃ��LҢ�^͖�R�"ORp��
   ��     G  �  �  r*  56  �A  �M  GY  �d  Pp   |  ��  �  \�  I�  ح  4�  ��  ��  �  U�  ��  �  ��  *�  ��  "�  x�  � *	 x � � �" �) 0 j8 �@ �G aO lV ] d Mj �p �q  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbE�X���Ț��<��FU0ݰM��E2<P���4��v(<a���%>Cd�e��O[ �E�D�yp���C
Or%��J�H/�L�%h֨k�� ��'2X#<��'vJf��u�� ��9b�w�<�+8��uȧㅕ!Q�$H��K�<�R�H��T H�|�1R�	GE�<!F
D��&0S��*X��QӅ�h�<�3+��~U���Ó2^����b�<�TE���ؚJб�l��C�R�<g ,�dZu�M $Ւ���Q�<�ծ�'�8��'^7z��$c���K�<ЀQ�1��M���B.<@��΁E�<)��K����1�[�P ���C�<�� �+@�`�UGB�X�>`���W�<Y�.7E��4�P.��~wh`:�Pn�<��'S)"��%ʚ�6,�2 �l�<	aN��8��끇ݳFM���a�j�<���B�5ܜ����;q���Sk�h�<t���ER3Κ�Ua 9a�\f�<��%�4AZ���&Nc��ʚa�<���� �F�+�Y0:<����JF[�<�R����� &g��!�D�QgZ`�<��,9h�2�F���I����\�<�peJ81-@<�A&[a[�D�<���q�"���`�8�U�q�B�<���\�%еi_�vI� dPc�<y�)"b��@Q/C8�d�B�i�<y k�$<�B=��j��?�$Ei�b�\�<��υ�#]�A�)T":����b^r�<�SjԲA�c6�<�,va�m�<I����a�>?h`W@�q�<���{��8�Q��.�SEc�o�<��蟿{��X���B#p���Q�INR�<i�
C��JD��M�]���\N�<�@a\Yq��R�v��@��DTH�<QB��6�.�bb�űEU�A��DZI�<��b�F��2�슯�F�p��@�<Y 8v�l��Ü/l��DK�|�<�$��
I���{��D*���Ҷ�]D�<)�C�]0�� &o�����c~�<�#ԫ�2�$$H�f��=B��L~�<��KZ5z�8)kd�E,U�������v�<�3�ϡk�z0D(R�~f<zWm�h�<q���0e:<�S��άI,��qd�g�<���f7�01B��(Y,U��Fg�<qPGG�JM:yd	�A�Sq
�H�<��fH#.�"y�"o���Cݘ�y`�"`�x��S7�p�ч-��yρؖ�9���ã(��Yb�ė��y�CE3r��lZW�8X�nD3����y2a�S��帑���Aj�I���y��oxD�׎C�R�~)�F*���y���c���ud&~�n0����y�����h`"��q*hD�#�V8�y�ʬ*4�P��֚;VQ
ώ�y��ۡB{���N�2,�5Rb��	�y���/#A2$+"$��'�����Y�y�lԠ:�
�вH�q~Y�i;�yR��&6U�h U�Ôn͔D��F۟�y��K:�|K�a@�e�\0��yr�M�>PA�_;sy ��/5�y
� �(X��	7����V䋣{�ԭq1"O���E��T�nb �H�o.D��)��ʏDfda��2�ES�i,D��k�F$+\�� ��Q�r�J��+D� P7�E����KE��YW^�ْ�Oh��Or�D�O��$�O����OJ�D�Ot�h�Í)-��yz]�|��1h\�?����?Q��?���?����?���?�c/�?m?2�ck�ZDp�Se��?)���?y��?���?���?I��?Y�!��khr1:�(�.Z��@�@�?A���?���?Y���?���?���?1Vh�Y�֠����%i���K'�I�?i��?I��?���?��?��?���si�)��^�T�X\�p����?����?����?���?1��?y���?��@|��X5� ^�&1Bf4�?9��?9���?Y��?���?��?I����
I�����!R�� �����?Q��?���?����?���?����?��������W!Ǳc�d8�3�ߛ�?���?9��?����?���?����?���4X�#� ��,�p�S��?����?Y���?����?���?���?��D�����/
��'$P��?���?��?I���?9��?y��?�&�[�6b���T�*ܼ Q�ۏ�?���?����?����?���?q���?a�	�YIZ�R����d!!2H
	�?a���?����?)���?��O��F�'c��R�e�l��E�*V�B�Q��3.˓�?)O1��	��M��I�c:��w�0H,����!�(@�'Ξ6-&�i>���̑7��$�@,�'E�<�� @E��̟�	�'!��lZh~�8��M�Sc��1-�=Bf��FD��P�\�1OF���<1����
G�l��E�=1.`au�G4{�Ҥm�f�jb�x��d��y7b(xJ��A0"�*D1���.Yc��'6��>�|B7���M��'="��잦(������.�*���'��D؟�2��i>����Kp����5��I#�E^_3�	@y2�|bc|�|a��V�.�*�喾z�+�䜮`j�$�O����O���o}"���6!3)�[���ˉ8����O�[���q�1��S�q���$ǦX �0�R�jyTa��d�pʓ��D�O?��if�B���tҺI�`�)���I&�MsWw~Үz�0��^%Hy �e�,���J�5R�x�ן��	��H���Zʦ��'����?� %�E�:��TI��_��;�Ǫ\ў�S`yB��t䋻2a0E�,�Y��u�B�������)�v+�Ip��C��(�����U07���KG���d�O�g��&>=�	؟�����CVdܳ@� �V$
��Р/���9t��>iQ�mӸ��b�'V��'�t�'2��@-M +������-�>��5�'��^y"�|�Dl�dȺg;O@t�P-GDFh� #�R�0O�L��<O.�lZM��|��?)���?Q�j8 ,���  d��H��E/�ߴ�yҠ̐���O�?E���"���/u|kl�>*(�6�ʣmwd�2�bA�]���O�����S�;�2�����a�
�(�&Ǹ9Vc�8۴! ƨ�'ƈ7 �dK�!Ŋ��@��� R�	�db�-l���X}"�'Nb�'ւ}�i��d�O���^
����t�;nn�ȕ�F�ZT����I�\�=�'���ORi�$O�!�D{��#���ɶ3O��O��lZ�{��c�\��?m��ʚ�P��x����?t���"&?!�\�����<���'�?Y���;j|�G_4[��	��k��?yf���C}�]�'$�����p�|�'�!W&Fɹ#�� F���u��YJ2�'S"�'���W�4Y�4K\��dX���53wb��>~0%�@M
�?��  �����I}"kf���j��ۈ!��9:��({l@�����E���TJ�nZ�<��k#p$��h����'-2�z�Ԭ�^4�97F~��'��I����	Ο�����D��T��!�'Vv���/��~�*co�[,�6�Q�S��D�O���#�	�O��lz�Q�4��4 �� �^��Hh����M�2�iɧ�O֭�P�i:�W�t�(4RuI�m��(�#� ��C�h�����	>0�O���|r��Q�=Fmݘ�:mЈ��X,:��?���?�)O�Ynڲf�4��	͟<�I+T��9d�D�֬����3;��?	V���4A����|�?cT��8��\���(�@�����9=��*�% s1�ؐJ��h���u�HIQ�Q�]�ѧb�t���D�Oh���O@��+�'�?aI��>����1�G��Ɉ���?i��im:����'2"�rӖ��5��}���S!*��!3�E��r�ɧ�M+0�i	��G�s������������_�4��QT��r�r��J��a�l�%�������'T��''��'��5#� ��Hde��!*,ܡ��[����4��ey���?����'�?��Î�C�j�S7 �u�<`SH �[8����M[T�iaɧ�O�Qpc�G�?h��k�A��2cؙ�u�B�%�~8��OҰ� ��?ɕ+-��<)�Ė�L����O
`���k��X�?9���?���?�'��$��9�"��ٟ��-�  $D H���z���Q���:�4��' �r��"dӞim4�:��ѧB�~�Fm��� .-zX��ƦM�'�����?�������� �i��닖�`�;����;�BD�A0O���O��$�O����OV�?��tHY�cs�ԓ���x���(�o^����I��p��4�p�ϧ�?�R�i�'V`X
�N�-5�@�
(mZe��e&�dn�~�n�?��ᦝϓ6��y���9,�L;�'W����&3��a+���O@%�J<��V�D��Ο��	՟�R7!̑8'�d �戝B���4�����Ay��{Ӝ����O�D�Ol�';% �a�M�!^�&e@eY�H�X�'D�X�f�d�u'��Mm��[�uYf�y�L���DH��K�F_�D8�EE��y�ȅĺCBoӖ�?�Q�1}Zc�Jq#Fd@-?<�ŢUƘ����	�'_b�'D���O^�	��M����*`g�b�D8+.]�A�ņ	����?�Ʋi:�O���'�7�M�\м�����+d �H�j�bb�m���Mӷ���Mk�O��K�̗����j�<鄉&� ���E�kȲy���@�<a(O����O���O����O�'1�J�a\X��% ��N�mb!�	*�ƠϨ���'N�����'�"6=�D���Q
qp�۲���!���A�C����S�4����O����v�i��$M���0��:A�ۥ�ׂ�~�/��=�9��(��'�	��T�I�Xxa�Rv72,:#���Dd����؟������'T�7�R�9h���O��d�bw��bs��
`��N)���-Ot�do�l&�`[�JW$Hrs�
^a�IP@�2?1���;F������'B��Δ�?�u�V d¬����!&��C͵�?���?���?	����O��r�Jv

���%\$%�XX1�O�lZ97��	ҟ�8ߴ���yG	ڶJx)1rNЕz�[7����y�w��n��M�����M��O6̡��I�V�69�i`#k��=��"
xy2�O���?1���?����?y�f�`�{1�ٍ�n�I6,V
B���.O
0oZ�P�I�����N����Xх��4"�0J��m��sp 
&����ڦ1��4r���OZ
����	���+dF��V�Գ4���&Ȟ4
�_�Dy��R�BB)�o�IsyR
I�**!�b��&��Pr�F4���'�B�'��O剠�M�w/E�?W�S�y�$l�P�P���?�2�i��O�і'�i�7�o.2="Em�$TZ��<L�1�Bu�$� �4�d��zQ�I~B�;Ӹ|��f�%�6��\�n�1��?���?!��?I����O��ђ�/\#3��rf(_';��-��X���ɬ�M#A���|���N@��|2�޲&�
ե�=[��8�/A��O~�m��M�'`� iK�4���X�iL��p4�Ê�~)!L�C��;u��?!��?��<���?A��?�*ʲD:X�$f�7Vz���bX!�?�����$ۦ1SAǟ,�	ɟX�O_T���W��깈�����Zȉ�O���'T\6�_ʦ%�M<�O�̺`J�'w��12���1��*��� \z�i>H'�'�	%��"1"���2���;��i�$��ߟ0��ş����b>u�'r�6��."�L�V!!SΰU(�Gڰ9�H��0B�O �D�ĦQ�?�VQ����4I �(��H��a�l��h��%�D�i�7�BB��6Mv�H�G�.G��tk��O|�@��?1�V��h� ���e��\�Bb�O���'u��'"�'���'�.(nHȵ%�Y{�1��	�;��9��49{>�����?A����?Q��y�Y��yG��3r���`M�1�7�K��q�N<ͧ��' d��9ߴ�y��
��xU/Q�omB�)B���y���W���I�"u�'��	ݟ4�I)6n�0�sD�:A���S�Ɖ2����I̟���ϟ��'h6��b�z�$�Oj���!7���V�>��(�ۧ&N��D �Df}"fmӠioځ��Q���*[6JFDĲ!��c���ϓ�?)eD,K�T�����D�� �2��p6�d_�_�Z�Rt��*�����cӒa.���O���OX��<ڧ�?����p�δJ�æ�(��ф�?���i�&i�$�'`��kӮ��_��A���q@>��%����	��M��i�z7�] �6m%?1�KK9��	R;c�`%ے�I<ᄔ)N�L�;L>i(O�d�O���O
���O��@��OB0j��0�3(h�s�
�<�i��Hq�'��'��O�R&ɍ[=p=°�	�+��9K���H˜�M�&�~�(%�b>��sfY*�ҍ�`���nD�S�^�Tl��"��hybO/{�Z��ɾ��'��	3�(�O�::f�3���Y���Iɟ�����H�i>�'�H6MԜb���!Bƚ1��K"K����*X�����Ҧ��?	�T��ߴPa�֤pӒ����փ��59��>R@�d�/:�7�/?qѹ+�&���.�䧠�k#b��=kh%���8C�¸h�n�<���?����?���?i��4�,g��)qA�da��"���5rP"�'Rq�4��T>���$�æ]%�4ـEK V���iV�wOP���.E�ēr�V�g��i�� ]t7�.?Q�ȖVkθ��ߎ����*��D�h���f�O��K>�-O����O(��O:)1�`�x�N��7� <�p�x��O����<q0�iP	x��'8��'<�S�G�ЅȦŎ`ԉb��y��j�	#�M�ĸi)�O�'`�"�;Ǩ!N������=R1�l�	��~ d宏��i>����'�B�'���b�)9ꥳƢ5	��������I�����Οb>��'�66�0'��pB"�	a�|�k�_x�	P���O��d榝�?i�Y��3�4L����y ��ϙ)_�d�q�i�|7-�&^<6,?��A�v��)��� �q�8c��D
A-�Yr:�6O���?���?����?)���	�"^�Isl��9ۨ��ߨT���K޴8�Z���?Q��䧪?A��y瀆m׎PA�/��^"�a#"��2�n6�ѦٓM<�|�Pi���M�'a�B��y����w��XB�'���'A��D{7�|2Q���I֟�y�C�Dr2��'��\�ԽI��џT��ş��Sy2by�Dir���O����O ({��j��1���	;�hbf"��������4|$�'��Y�Ԇr��\�� �_��yӟ'�H](7�N*K�z���\4��X?Yw#M5�u��O�Q
p×�Q$����G߁W�l�!`�O����O\���O�}��d��؊�N���t(r�^?c���������AB�'f�7�$�i���〚#
�x�l��?t�	1fo��ٴK�V�o��H�@pӂ�I�p�Ch��u����LY�{���:[����^�~.�$���';b�'m�'���'��ٷ&R#e�8  ��2s�f!�R��ڴ_x�����?9����'�?�F��R�����BLX 
�ké�8c�I>�M� �ie<O����)Q yؙi�D�$!r}{P���X��<���L��	�Y$�'��'���'r�p�e�|�X�e�(�̡��'B�'�����U���ߴ#���������f%�h�!��(�'n���?Q�6��U}��q�T}l��MÇ��j����e�Iؐ=bA#.$��5�ܴ�y��'ht����?Uy�O$����V��L��S�)�Ǯ$	�.A�:O����O���O���OH�?B�a�Yk�o��c�"}�`��������(ܴw�"X�'�?���i�'�����U��]rb�D[�II$�!�\ڦm���|2���=�MC�O>=p*��0��p�F
I�+�@��r�F�t��Y��g���O���|:���?y�XKޠ� ��	�͏�uG�t����?�)O�lZ�3R��͟L��x��)���1@dD^�pt���II>��]}}��i�4Tm�1�?�O|z��H<xs�$ θ�2�݅Yp�<Q�d���r+�����d쟶����'8����`�%X�0}aM��2��E���'!�'�b���O���MB9?,��ʎ � eaģ�+�#?9w�i��O� �'N^6��	hx���'ӿh� �b��\C
�m�M�#��M��'O⃝�?��u��+$剛'd���AA3MG���'
�&��	hyb�'�R�'�r�'q�_>I��ÑGˎ蚥+� P\��E��M���<	��?�J~ΓF���wےH�0oP�`U:� Y;	�س�Ai�f�l,�?I�O������IH-w�6n��8h��	V̪�&Ǿ-"���s��H@Oż8b����<i��?y�IU7y��2+E	Vn�dsa�A��?���?Y����dP����V�d����0(Re�"~�x`@0"Љ9���ņA�t���*�M���i,����>���I<x��"�g�T0+�.��<���~,8��	����+O���&�?��'�h\���U�Y+Ʊ �
�b�DB��'���'�B�'��>1�I�o	N��ɯv,�y��gK"� ��3�M�3�w~�{Ӗ��ݳE]��3w怀z㮡����-��.�M��i�(7��G`7-p���:J���3�O~�� ��̢2����HZ.KDp���8��[y2�'���'w2�'+�/G1L8�a"�[���[��	��Mkq��<���?!I~�8�J�RRF/nU�P�;��-8����M�f�i|��;�'!����N F�MJ����t|X��͍*��)O��2k�7�?��{R^�����.b�n��aS�d1{
�Ɵ���Ο������iy��iӜ��8O�L	��<붨�%IM	*�����6O�o�T��R��Iȟ�nZ��MK7�/���E�0�V�Շ.C� �۴���V�`e^����V��މ��I!��2��ր9u���� a�μ͓�?I��?���?����O_~�kX�P����V*t����'���'(�7M�~���M[I>yG-�J�Z(�N_�U��<{� F#r��[���ܴ'��O	�%zбi���9jtZ��͟�G$�,Lc�\�pՠ�"0��� ��Xy��'�b�'D�,�=3��wg�
7耫�C�M���'X�	�M{� י�?���?�)�b1�У�N�椳D�U�<��]�×�ts�OLnZ�M�0�'ﱟ��&�T�+�i��oY,I��y1f�� C�L#$E�69��|�cM�O(�PN>!�rSj�u䈊O?������?����?���?�|b,O�xm���3.�v��a���C)�0k��M@y�mi���a*O�6-͈��B�S�>��}`w�^�iҜ�I�)z����'Ja����?��[�|ppj�mL�=p둃~��k�p�'��'#B�'3r�'�哿Q�4���'E�.��h"�]v� ߴ��H��?!���'�?	ջ�yW��85��X�(*<�H���cϱ*E�7�R���&�b>�R�HݦMΓ
�&Ի�J�a ��D%͓H;����D�OX	K>�(O��D�O�t���ɥ4�$݀�DO5�qx���O����O:��<yS�i�PX��'���'��E ���?���T�J�i�c�ċby�'K��x�	��;��$F��8Q�D�^�y��'<���C��.@���`]���S�0��������3z�.-*��Ȳw��) G䟜�I럈�I؟|F��w;���w��6[�^Q 2��3r�Sg�'W.7MF-A��$�O*AoZT�ӼK�]�'LP��ר��1l���m^�<y��i�7-�ۦ��P��=�'i��0�/[�?�K
� p��[Vy�  ����:��>���<����?����?���?y6�	%e�"�У�R�v�R{'S��	��s��Ryr�'x�xJ�Ǟ�7]HE��m�Q̄���E�a}B�b�&�m0�?1��X%2#ᰃ� �8��ΠS�<�:ӏ	4���<��y��+�O�kM>�)O�T�Ta�2<K8��/�/{�z����O����Ot���O�ɸ<aԿi����w�'��T��+A-x$��Bw�'/r	b��'6-$�	���D�Ox7�Yݦ�+6*��[T =��hŴ0yH�P"H��zI^�m�Q~2C�7Ђ���@C�O���ػi�X�	��
�$��G%B4In���ݟ��	��(�I����	A�'.�R=�A�A�G"�F�������?y�kf�ƀť��D�'-`7�:��U/�B��q���uf�C:�\+��xb�~��lz>!�NE¦��'�zr��M-Cd��U��e�x�D��w��|�	�\4�'��i>i���t���$��=�P�P������i���������' 7�Ь~����O��D�|��@��;��	�E�o��;a�[~�h�>9D�i�6�AN�)Z6O�Z��X��!�`E��
g#�Ukȗ?!D$�����H6�|LS.rJ����g��\�2/�'���'���'���dX���޴9�@�B���+6tkd�ӛg�iZ����?�������$�a}��cӪ�0�kݠ~����6l*ni���Hɦiܴl�=��4�yR�'�%t,��?yp�O����$|pnL�t���~l,!�$<O���?i���?A���?����	S�bxQAڿo��0s�E�1"�\�mZ"R]�M�I؟X�	d��؟�����V�^�H/�E{�b�A\�8R����iٴ-�����O�D�@,��6:Oj��		YB2�G�.-1LZ�4O��1�� �?q�!��<�'�?tc�
kg�W�x�� �̉�zD��������I�(�'�J6�ӧ}c��Ov�$����@���6^v�(pD#br�[�OPlZ�M���'��I u5̤�eկF���b�b5�z���j��%f*QQ�o@y��OՐI��v?��	�?A�|�HH�e�Xa���?����?���?����OP��#��*��L��X�rT��!�O�IoZVٜ9��ΟJ�4���yGE����L9���۱<���Q��O6M�Ӧ�3޴"��iش�yb�'،�4N�C���QoX�����˷ ��9˄�H��䓢��O.���O�d�O���[5n �pp��(-`B!�����}���=����ˏ] ��'pҔ��'��ba�̦&��!C�J�TC�u ���>��i4�6�{�i>����?�*��,�#Bӽ}��d�2�@�<u��0	��I�'Ҭ���P?�L>A.O�qa�^�5D @���jd@����O��O���O�	�<���i�`��'�>E����@9���I�R����'�67�8�	��$�ӦIH�4N��&�W=36M`��Hb#��K�"Ï\ôTS��iJ�I��r-��ӟb�����B����"�in-�V*ɷ:��D�O���O ���Of�D?��G9굂硜�{�dQ��*�U��	�L��8�M[�E�|r�z�&�|ҫ˾C��hiQM	YK����K���O��h��̶nu7�.?��%�!!_.�:cK��f���Ҥ$E6�`���e��&�l�'���'-��'�=��ӶCG�����^<̓c�'bV����4����+On��|�D�U�d-z�Y�OL�( aE,�@~R �>aS�iW�6MK�)j���n �� ��0DP�(x���$ު])wGș�M3 \��>;F�$1��T5��,صb�2�Y��BC/a��d�O��D�Op��<�4�i3d�����7$��	I�M��҈q��?X�'z�6�:�	5���l��1j��|5�(��@!F��牜���۴l�
��ڴ��W�50��O����l��� DT����8Y�V��Wy��'��'�'�\>y2�+Z�^&x�81�ϭr&PX��*�M��.I�?����?�����u��Ƅ\�b�9&�=%
P��҉�/x�HlZ�M�w�x����ޏQ;�6=O�!�D㜜#�F�[� �x��� �6O�ɩ$���~��|�S�$�������K  v�m����*�4-�'"ǟ �Iߟ��I{ybGh��`�w��T�ɚm�jP�VL�������"im8��?)Q]�Ј�4."�6��O��!�X���m�<�jI� kk 	͓�?alL/.Sf���f�����8\���~�D��?�D`���]�P`���J��']2�'m�Sӟ��'���s�& ��ә1M����ڟ�)�4|�8|�'��7�/�iށI��R�5��)%g�+������ym�֙n)�M��Q��M��OZ��T)2�RTI�EJ���Ʊ �R�b���1O^ʓ�?����?���?9��g7��ؠi���-�7)�"���	/O@�nگ~��	��H��G�s� S%IE!;ab�J5�S�&�aȈ���D��eq�4%�铿?�D�����i%�\�SG��=i�\���F0:ɠ��'�P�smɟ��=�.O|���(BH�ak H�l`���!a�O����O���O�I�<�g�i,$���'O����E�x(|E+��@Z�jȟ'�^6�%����������4"ʛ�i�!N�����-�&��F�w�,`Ըi��	d�ys��O
n('?yR[cP ؅Ł7ڝ�1靤Z�~�')��'�2�'r�'S��	 �C�3�0tY����u�?O4�$�O�mZ�Y��[Z�&�|R�P�Ih�M��,�?���غq����>���i��7����@Ғ�uӖ����#D2� ��3�#J�)� �CEW�@&����8�?��{b[�8������꟔��a�#��#�(��b�xճ�DٟL��oy2�j�@�"4O~�d�O�˧>������^�ĒG'�).�'��6��A}�(l��x�S�?y��� Wkx��;J���� ��:s<��4d�(����'*�d��ӟ��=i�fʵAm���L�"�6�ꗤ�?	��?a��?�|z(O��lZ�L�|�˗n&i?���e-�l��$���'?9��iL�OR��'��7MS�X���G�6�Fp�6T1YKr�2�lZ�,NmZ�<��;��!�$��-Oީq"cż���p�!�G��L�3OZ��?����?����?�����ֻ|N,��Xwe�8"�R��E	Ժi�=��'B��'���y��~��nQ: �9"H�1 �l�����W��m��M��'Z�i>=��?5�S��ަm̓&�PY�Ӄ��u؞p�Q���x<N�9=��@�m�O^➴�'�B�'��2�B1:�)H ���u��7�'���'S�0�ڴ&� ���?���Ȁ'�K-����'d�?Io\(;���> �i�
7�P�1f���\� ��9�FHT�3C��tA�����rg���|jQ��O����NZL�CI��&��;�F��3������?����?���h�F��H2��!�bŪm��R$��2��$���͂�J�����	:�M���w(����pTJ�z�Z�4�D��'Nj6��ɦM�޴G����4��Ě�vi4��'¶}p�AS��J�T˅2`��dD;���<ͧ�?���?���?I��V�F�d� JO�q�pla���&����-��D����I��|$?��	�#@�a&����-�Ф�52)�(On��bӼ�$����p�$�R'��D��;+�8Uq��[/��u" ��d���߰
T_�qy��@X8 ��%/p�p �'�N�3A��'d��'��OF�I.�M��H��?���7kʒ%��
�b[&<�fD�?�Ӽi��O�)�'�6mLۦi��4<00I�܉7��H[c��w*T��%����M�O֩�T+������w���3��ʢT6�d�5�(��	!�'��'XR�'�2�'�ؕٶN�!SY�ıH�)MIN�@���Or�$�OЕo�;b6��Ο��4�?y/O�Ӌ�>B�A������Z�h�y≗�M�7�i3�t�:���:O~��N�j��<#��
H#(����&w��i'a�2�?!4�2�Ĭ<ͧ�?i���?� YF��T3�F��(���?����ަ����X�I���Ok`@�Š�d)�����' ��O
��'�6m�̦�iI<�Oܘ�I�������&��𖍙��NIˠh���4�t����X�OM����p�d��V�)4�bM���O,���O��d�O1��˓[ћcF��C��	S.��#�Ϝ N� �'���k�㟌�*OB7�)�ڙ�fi.D�X�Ǫ�%_�:�nڻ�M+JҼ�MS�OΕBDi/�B�*�<9t�_3jXPɘ��^�[%�H��j��<�.Ol�D�O,�D�O�d�O�ʧ=��	��Ђ6����u��(��5j�i��8S��'���'~�O���~��n��N��9z��_�F1@̚�IN�i��Mn��M�'�'��i>����?�j�]Ǧ͓,{�4{C��GF����#N<Y̓3TF�� ��O�9�N>�(O����OVH@�] d�|�8�&[������O��D�O��$�<mx�t�J��O��D�O�}R�$�G'n�a%�#z]¶ =�		��$�̦]J۴!�Y��b�S�(T$�f"
�N�VH��g�6�i̠���
~tRH��T��S�5&����l��H�
�vq���=h��@r�]ݟ���̟���ʟ8E��w�82��Ä ���4[�:hC��'d�7m4G>(˓Tp���4�&�	���7G�����ۂY��)�P=O�oډ�Mㆰi����%�i��	5�8�s��O�4(·-M��J���BO�<O�q�j�q�	Dyb�'l��']��'���b�Ĵ
1��,~b���J�/J�I��M��D��?y���?	L~j��V����'�-al��!eV�},��Q���4P�6�/��i�3>��qH��bl�vȗ�s$��WaV/A��.�� ���' ��%�,�'l h�!G�:�8��BR,^��7�'-b�'2��TP���޴k���C��O[���$X4�
��`	�+�*��Otm�N�JB�I��M�F�i��6�)��Q��b��%��8O�Μ��T�p�����;���?
\����e�S��5�cY.o�GH z��["�yr�'J�1��G��F%x��'�ƙD�$tq��'z��'��6-�	O�Ӣ�M�M>k�(BmGä*��!� �@��R�ԙ�4"��O�>�*��iU���XG`�	t+E�c�F���g]9I���a��B��oj�IWy��'���'xbLN�<n��3��J�m�:�*c�	7 ���' �	�M[ n��?	��?9(��A�LH73>�h�F��Da
����,�Oʐl��M��'ܱ��D`���}5�0�@Ÿb��qg�Lh���ʔ�#^����|�b��OD1[I>�)׹i��G�/",�l�d�Ԁ�?A��?����?�|(Ojxo��-V����O8J*�ã�`7@
"	������M���,�>11�iM���@NN�` %��*^'q��$���y���m�@�F�mI~�N�`9 �Sb��V��䈥('H�&�I�mW#B��D�<���?����?���?�,���j��2D�L2���Z{^(�����}�B�џ@��ȟ�%?I�I��MϻD|r�kAA�ZJ��Ц� J2J��i�"6�Vҟ�է�O����C�iG�� ,xPǫ�#ch�� �ȥ5��<�1<O:9��:�?�S ���<	���?I.�&W��j #�
}�~I��S(�?q��?�����KŦ��IE�� ��۟ذ����fsH�$ma�~hb�L�zE��'�M�D�iB����>�U'ʜ+8bm�w��u�m�E~���;쐔-f�
E�O~:�d�O6E���pd�1����F����A�[>��B���?)��?����h����M�|(�R� �1m;ġ�r�K+����񦥘BI���|�	0�M��w�HXҠ��gv�@�;�\�p�'��7��Ϧ�޴.�v0C�4���	7X����'D���t�����)� T�eV�]CR�2�d�<����?I���?���?�J�(G��q���n.A��I���ĈڦQ�2)˟,�I��%?�ɷT��ث螁f�D�q���$A8��q-O��D�O�O�O��H*PE2EԵ�jL�h�C�ݷ;/�qc2U��a� u����F�	`y¯ۀo���N�5�j���N׆2�2�'���'��O��ɻ�M����?���AI}���� �NX�c`��<���i!�O2��'��7-����o��8(�솆d+�����ie6��E��ϓ�?I0����	�����<�n��.�L��e�jM:��l��d$�D�O��d�O����OH��?���X��☁L�8 �%-����	۟4���M��`P������	Dy��Ƙf�Ts ����["�=4(lO�mZ��M��' cy�۴�y"�'.jL�;n�|�yӢk1��'ˢ|	���'0	'��'�"�'�"�'JdS���v�^I���:M4�:��'�_����4's������?�����'c�m�p`z��AGaL�\|�1�'Z���f��OO����y`�B�����)nrP+'��_DTa��?7����1E�O��M>(�)Bh9�a�%A9F��"
��?Y���?���?�|-O�	oZ�8���C7�B�I�X�ɡOրU9;�jO}y��g���ɩO��l/�by���ނe��#��
N5�u��4k7��C�3���6O���5�*4�'
��ʓS���0ѯ¯H�4�Y���l��4ϓ��D�O��$�Oh���O���|��D�H?Hd�.�4n�ݫ����u���^��'�����'[\7=�:�C� g=P��̕	��ݠ�����4(�����Oa��+6u���2O�\�"i�/F�L�b�!C�{D�M�0O,���W/�?G�;��<ͧ�?6˜-�t�õ�ܛ���(`9�?���?I�������H��MCyr�'�" ʱ`�]t\I;���,4��Q��DSX}��n�h�n�?�O�Y(@��h���w��vҵ�R7OZ�d�UU�mX�$M#�6˓����O�̲��,b����8XF�����C`��b��?)��?I��h���D_�Q"���ɹ3/����!�*d����Ѧ���QyB�e�N��
'��x��,8!���
��	?�M�õiN6����V7�s���	�0t����O9��i�▮p��Ek��$;AR-�r'�K�Idy��'���'�"�':�EJ�G�r��PE+�m�� p���M[�R$�?���?1K~��O:y��g����u7̟9���Q�T#�4�g�O6�v�i�����U"MJH�`�h6(^�	X$"�-�<IP R np2�DS6����DLa��˵�A/@��s�撈t�����O��D�O��4���:����'la�I={G�a8��I�c����K�!`�R�{���,��O�Qo'�M��iXт�����k��9"�����O,<����ĳ��C�C���I��*D���_�}����s
��V�l(�;O��$�O����On���O��?"4���P�Q��!l�kG�U�����ӟ�	ش,� �Χ�?Yײir�'�H�2�D<e�(�S �������$��������?�A�O����'�H@1�cAx���&8b������F"����/U�'$�	՟��՟l��8�~xâDB7B����f��BC���I��T�'D�7m��a>��O��D�|�$���siF!:G�7���V��g~�d�>�a�iy"7��ڟ��~z5�Ld��U�6�TX�R�F#S3� ��Gu�k+O�į�?1�{��U�D�G�ϣ`�
�Z�M�J8��'d�'����Y�8)��7���A�w��a�C�"io0��n(?��i��O���'6mЋI�Xp�R�0l�R����J�M�ưl�	�M��ײ�M��O\x1ElI1�����<�l�>k,|P���co|������<�(O��D�O����O����O�ʧ�(�K�'� 3�L����=y��Z�i�$T�'1��';��y��o��.
�g����U�2a4m��'15"W��śF��O4�S�'��Ѱݴ�y�O(�b�j��+x��y�]0�y2(v����I���$�O:�d�3[wH�[@M�t�����b�T�$�O����O�ʓ[�����)mK��ɟd[����w�b�[0q��b��Vu������M3G�i7��D�>�v�1g�91E(^3$d����F]~�P�gW����I�Y��O|���ɍY�2.L(�tU"�:1�d+�$!�b�'6R�'��������5D���a�K�y��u��I ܟ�S�4�@q���?�&�i��O��9Z��@�*M�N�&�p�Q���Ȧ�8ܴH�&�����f��d`�B�P7��
��s�D-��"Ȋ��ܓ~�|'��'���'���'v��'2��`+�$Hl`%LDDP��7R����4-�f� ���?�����<�!�=o�d#c� �{_$�z�c��	��M���i-z��"�'o���� v�;�J� 5�X2"�?{����R-ֺ,8ʓO�Tm����O�|�J>�/O����մ{�t�H���+r���s��O|�d�O���O�ɰ<�վi�P��6�'s��K�H��������m����'-z6M2�� ����¦��ߴ8���s&.�J� �1���i7@	_�xzԺi���%LxAb��O��%?�J[cuz��%S<+�l��I3�|1˘'X��'���'M��'��V�zAͩ$�t��Ī��*3�,x���O����Oj�l4L!�۟P�۴��.���IlO�6H�B�c�4��2�'���6�M3"���h��F��T�7��e�bPaY�eS�݉�"ÛP��p&�'�A%���'QB�'R2�'����`�_-r@�� �i��M�'�R�'z�	;�M������?����?�.�d ���9K����4쐚7r�]�b����O�Xn���M#q�xʟ��' ���Ć�=N� �g�M�@ITB~�TQ����k
a?�J>ٵg�#w�Ve2˃0d�:�p�/��?���?��?�|�.O�lZ� K��r�P)q��>04�c�qy�.}���q�O�m�4U�k3�L%9�,%�ᄂ'o�RyJ۴bl�V�U�UG�&�� c��9��ɺ<qD�ĉ&��pS��H,�ı&��<I*ON���Oj�D�O����O˧[�tP�
-G��$Đ�~D 4�iWnDK��'�B�'��O�2�`��n��?�8Ѫ�>��8a%�,�6�o��M#t�x��܌F>7mk�����R(,�f/�[+L���Do��A��k��%��<I���?�#��,� MK�m,�z�ᨒ�?���?)�����-s�*V���IП�£'�6{�,���B�'b�=R�h�������M{��i��O"�
��J+�v�pE�P"X$4*`���h��T0i�dn���'n���	��Y�&�:'�2EKpa^d6HaF�ٟ\�I����ş8E��'7��k���6�6E�WB�q�B�`��'܌7�3_�B���O2im�w�Ӽ�g�T�p�(�gl�K��X�M��<	E�i��7������ڦM�'�hٲF �O�u�T;!�v`��J�j�8+Ѭ%����d�O*�D�O���OH�ɛC�­P����S4N��q�O2�ʓY ���P+~b�'����t�'���E
�ʬ�@�^�#"Ȥ�S��>p�i$�7M�Y�)�S{�M8�������5b �9˞�jC�M�Sr�s�<���O�ZN>-O`u�(FGH1R�n��-�4qr���O���O����O�)�<Yǲi� �B�'[�e�C��ɚ��ƴx�MB��?9�i��OR�'�@6���m9ߴ)�|��߫o:t}�@��u'I�MK�O(d��b���j2�	J��"CU�0T��+~��h�֪�<���?���?����?���dg����`&fT(��4[���:~r"�'o��e�ڹ#�O�tӴ�O�k1�ˊf�� �+�v*���u�Y��'�7����S�I�el^~R�X�p>�0�E��>7�"$y�M�,hX3Q��П�sß|bQ������I�J��asd�Rb��
zN��5a��� ��~y2���h���O����O�˧DX�%rfE�'����%e�u����'�D�E����kӄ���h�'r�����7�2�@�E%5b�`G��N~���� ���4�l�����8�O���0��"�R`�0mȇc�R����O.���O,�D�O1��ʓ9����</^0xj"�tP Pɔ�r&�Kî���d�䦁�?iPY�$Bߴn�2�#���>*:y�ӫ#�Bq�!�i`b7��`��7M)?A�*.&�i#��DF4�p���/%�@�c3gA%&�<	���?���?���?1*�$����@F�D����_2�;��ۦi�D�H۟\�	şT$?U��-�M�;L�<E�sdV:���5�ǊQ�Ұ�`�i��6�����ק�OL�x�C�i��d	�NI�A�q�KQ����A-:F��40e�0`��T.�O���?��M@�h��ۘaL-pWL��1�(J���?a��?i*O.�l:����ӟ �IO�f�R⎇8b��MH#���,P�?IR�LZ�4aś-��"D)25�W�c��5� ŜG�I��0��]�O~�p@����ɳTcTP1�1$�x��dB|C䉪���Aeѹ@�ȤSf�fZv���&�M;q�\��?q����4�^�!�a[#3��#�傸|QL���O��|�(�oZ�a���mw~a܊(?�m�'B~�OC1wќٰBc�:Ef�9jN>�*O��?��e[�7� ������܈B��_~"�o�F9Qd��O �D�O~�?}��dI�AP�0�Cğ�bh.D��,Q����ܦ9޴)�R�S�W'&`(�lUa`@���[�_M����.N�2��Ĕ'Q~E�!_��4k×|�Q�D��JF{T(���ڹW$�(KSk����I���I��SKy"�}�RL&L�O�0k$����Ȣ,��G
2Lp��O4�o�W���I�M��iN�7�X'�=�F*[�H���St�^�_�����d���y��3EF����>���=b(Չ�*�0�*���Cr���	ݟ���ş��	����	E����aIYq��L*& ������?Y�}@��Fۨ������'���_(W�v��bț8y���YVl��?y-O���y��ݝNf7#?���F?��t�A	�����	�C�,�S�OZ�ȕ'��'�r�'�H�9U
D�EJ��1�T�*�����'��W�h+�4]�L����?q����)N-R��I���=*����i�M#��9��dV��ł�4o���� ���G+� Ȋ���z:�Z���U~���A���G:���|Ӈ�O"�H>�d��fP�䫜
G����	���?9���?���?�|�.O�(l��5�d�A����K���c��L5�F��WoVXydqӾ㟸c�O��oZ^-�x����z�8 4oޫ/vu��4.��vI�� ��V��P���x���n�xy���t��+V�E%�����*��y�Y������X������t�O����V( v msA��rS�ع�jfӢ�xD�OL���O*���_ئ�TLj����S���IP���7�hi���M�R�'�)��K._�Z7�r��+3��Ya��a2HH&"h�5��|�\����$�bp��Uy�'�N85�5h3�)O�b��$ͭs�r�'{b�'v�I0�M;1'�'���O  r�
F	O��!�DC����, �I��Ȧ��46RP�� V�݈jВA:rəIl8�� ?�td�`�L��S���'u��P0�?ʹQ����BF�����F���?����?����?Ɏ�)�OpT�ax�	���hUX֨ �1�f�D^���{��lybIb����Gz� �TDZ	D,[g'���	 �M�d�'�F��t𛖘�4Cg(�����q�����l܅�ҷ6���7��$���'/B�'0�']��'{�$9�m��~�p�H�mQ�A&���U���۴	��?������<�͞?%@$*�L�f�2��gll��I��MkѼi����:�'Z�ܢFˋ*�Z�ae� � ����4����(O� �&%�?�B�*�D�<��	���N���τ42��	$-���?q��?Q���?�'��ܦ�2��ݟ�)v �B�2P0�� A��d�m�|�4��'�
�P���o��o��踹���	<q���È&c���*��!�'���rb��?�q��Kf���S�Y�4w���E��P	��A&}�@��I�7�T��!��:yN���L邅�I韈����M{��p�Td`�0�O(1�BQ/S��������Rc≇�M+����$��'N�f��Dbͅ�Fs�i�%�ˑ1Q��S�;U�L�bt�O�On˓��'_ܼSd���g�%��*�	L�@Dь�ئ��j�����	韀�O8H�g#�	�4�P��Ce�,��O�t�'%�6O�ѐ���O���2!\�Vݲ��G�ܔ�ɠ��+�"�Jf&s��i>Q���'b��'�l�ve̐hnP�3'��4��XRHS�p����L�	ɟb>)�'�,7�|u�wǬ bd��3.x���E�Ot�$R����?�a_�T	ݴ5��+���<�R���$�8v�[��i�6mZFX(7�0?y�'H<�N�����d�5D��@«A�7$ 5ó�Y9 ���<����?���?���?�.������'6���@�g9��KDj_��	Y ����	ҟ<'?��:�Mϻ���%�w�|uN�>]p@���i|�6�]䟘ק�O��cױiV��
6|i�9�C�K0*��/�$HU���F�0p���O�ʓ�?Y��xb���%ܗs �:���^Ű���?9��?�,Ohil�D�Vy�	�p�	Qe��+�(%JKD���.��~����?�_�t �4:��N�O��?@���V�y0�TjE� ��8u�'�`h���V�G�*	�0��DE�ڟp���'�51�'���HB��n�"}1��'B�'��'��>��I3`�XQd��#Y qPԬK	�`�	�M���@`~�/l����݅*0�-t�G�D� p��>���ɺ�M�R�i7M�^;|7�!?���_8�i²wp^�s�gO5s�F�"d��
A%,�`y��'���'�b�'�f�#̈́)�qk��`֞$�5��I�I��MS�B�<Q��?�M~Γ1Bmz!c�<0E$]�R͎�K	�5k�Q��I��qZ���H��E2t.ET@LIc�(f��ҰO��/��Yd�<��>��5�	Cy�97Mr݈���0��j�]�R�'�2�'��O�I��M��e��<�C�͹X �t��l��n��\
�d��<�p�iq�Op�']H7-�Ӧ��4w���dK�B:�PeO�d��&��M;�OZ { U���L ��]�k7 C��0Lh$D�$�2U�쳟��I�L������ߟX�
EhZ��s���=�����o�J��O,����Uc�M^hy2�b���O�yд��F���v 3 艘R�\G�	�M�c�24��'�M�O�yP�Mٍ:2�X¢�#o�ܴY�@�Ԭ�,�M�$���<)���?����?	5&�)X��=�QiZ�b��ŃӮ�?����$�ߦE�Q����������O�|���?�dͳ2���\��%8�O���'Ϛ7��$��'(F(X���$&�j��w��,$ׂ�b��%V8\i'+����4�`����Zf�O�yҕc3q��I`G�ږE��@$��O��$�O�D�O1�*˓aܛ���-n_<����	)#0��X4AS��@��U�T
�4��';��x����G� '��X�`H!@��K��z��oӌ��tdw�4��-�Pd��q�/O����qI��S�@�v�Y�>Onʓ�?���?����?9�����5 䄸Q�F�S�=C�C��o�Tn�2�Ҹ����	]�S�����Sǖ!W� ��7(���H�M\s��D�O^O1�Vyɤ�l��I�YM�ax���'�漓�$3��片g;(�J��'�(d'���'���'�9!�� V�\�s��xߺ1x��'T��'2\��!ڴ!{ځ����?!���ycʃ�Ui��� q�����ĵ>y'�i����=�� �U�P�� ip����
,~*�u���%&I*���8�*Pm�,��+��\��Ӫ
��e���BL���qV
�����I̟���ן4G��'в�	Ê �\\�4 c�//Xz��'��6��/=e����O�xo�f�Ӽ��/����ɜ-r:��vF?!��M��i��a0�i���8��!�"�O�X�Q�Q�*sfq��\��"!��]�Yy�O��'\r�'L��tЭbb�ګ水.a5�\r.O�Un��p�I�4��w�s����E���g �^1��!І���զ��ٴcP��S�%Y,Q2 � Y�FpIы��"� ��N>% �'���{����=�+O�X ��X�E\ ����Y���O����O��$�O��<��i�rD���'av�7��%9�ʸ��E(�!`#�'�f7M?����$�ʦ51�408�%T:��$��gN()����A��M�p{��iv�	?�z�)��OW`�$?M]c�Hz��L2XH�Y"H�.e��+�':�'���' 2�'Y�:(H�hM3m>yP�E�!�l � �O��D�O&LmZ>D���۟���4��2,��$��(D��h !��l$nY2�'#�	��M����T"� f<�Ɲ����U�o�bhY���Ve��oQ��Bោz��|�R� �I���ğP�&f� >������x`-0E������Hy҃|�D,a���O@���O�'[y�R䥋T�0�
V0aG��'�AA�f�o�u��a�'Ga�p:QᎦR���6�)S��t1�'N�������4�`�S��E8��O�M��eE��"��bӂ[�V��O�EnZ#W.`r֦D�3�2��Bk�/�4���<���MC�Ү�>i��i�D$O�լ�)E.�5���	��i���n��c�Imk~Bo��̮��'���Ȉn���E<p���a�W�)�D�<1�b�������$���լM��� �i���1��'}"�'&�j�oz�iC��L�*Pj�nϙ/2�����M���i�XO1����VHk��I.H�B�)��8<�� �K�6lHz�ɜ��ہ�O$�O�˓��D	bH���KЌ/C �I� ��:ax"	dӄ��!��O&�d�O��`�b=49���o��]�!�(������O�7mPu�ɍS@B�жI�� �p����^�������ӈ۶�M����$F^�S��$Z�j ꈓ����C!��y�ƒ5^rxLC�"�3o>�H�ա��9ZD�C��?B8�hS&⋳W	�h9cÙ#r*�,�G$�)[^��J��-�Q�Ɖ1�0q�p�#9b�\ UJ�/�>< ��5ΰj��΂]����شE���cRd��9�!�Ժ���FQ�eb��P��F2z!: .��GRl��g�����p�d"���X�dDT�I:�����rZ��{c(G+`+�0�3�]�r�L��UlU8}�*���.��(K�RdJw��;_*� ��U���B�GO:L�TiZvg$Q�v�4cAi[lyӊP�{ĐDn���b�=���?��������/ӌ<��A�������S'�u��?��������	ޟ�����q"ŀ>���EE�	d�듢�9= �I��$�	���	T�I����8F�>ȐP抑xՓ��K�EF.	���F�v�P��?����?9��?�g�%�?a�N�.��t�T�A�>jޗ�/dQ��4�?���?YI>����?��Q�u�Jm(%��L��V�H��0
�U	~H듖?	��?���?�$��I�O��f�,r%�*Fj�"D�8�$j��	�	v���ɨMmѪsG(�!w��!Ҡ{.�S �ԮUL���'W2�'B �@R�'6�	�?I�sπ3Y��l��)�1���[#�	��ē�?���l=fI���Fg�S�d �u�P=`��9BmL�y�����M���?Y���)�?Q��?Y����+Okl��!��P�q'��&�[v�F�,��&�'5��]�D40,3�y��tN���%�f��X��jՓ�M[�۲�?�����d���˓��D�k�����yw�D�peT�W���mZ+:q �`� 1�)�'�?Q���t�nh� nT�WE��ӓޕ8w���'��'bٳ��.����`����Af��G������-4}�>1��R[̓�?A���?	G�^4>���z�h��
(�t�.���'����/�>�*O<��;���@X�P$Ѝ4���5��n��t�R^�dH����',R�'�BT�0[� ����3k��e���ekU	^� �OV��?YO>����?���
�	��BJ�
j]���@�~ƒوI>A���?����O*ϧ~���m�&q��8v͟&��ElSy��'��'���'��j��O($yg�˃_'������6��RrR�<�	Пt��Ry�&E��맧?qg-D�b� c�Md���i�(O�O���'G�'���'V���'�A��Ų��L�!��X���NT:l������Xy�/�W2d맳?�����KH"���q��),��(Xg���'Y��'������'�'0���7�@q;GM��;B`�pd�tÛ�V�\��+[-�M���?1����sT�����c̊j5���mG�}n7��O���'-�����}j�&�C����U/Ι8v@�¦���!��M���?Y����cX���'x.�q'/�,V�����ǸB~����z�r\@É4�I|���?Y���2:oJ�ɰH�I0�1����4��&�'"�'R�TY*�>�(O��D���7�
�#Q��F��8����9��Fq�}&��IƟ���*�0�a3�īU��g��kU6�޴�?��3���py��'/���X�#�R!��c�L�����dזs����b2��k���I�8�'zN� ���P� h�H�
�kQ	j��m�/n��	yy2�'��'�"�',:h;����LI y�U"I�(�Zb�V�)x�'�b�'G�T����C����tA��$��͋T.�*8�D9qP$A�M�+OT��-�D�OV��܆*/|�	;>��a��dňT��b T��듈?y���?�,O� ���Q���'���֬�;����(����iӘ��0�$�O��DV�CF�㞰R�nˣt��H�F��T
�y�UOeӖ�$�O�ʓ
$h,;�U?����ӳ-5�$��+�x��
Tq��I<9���?�dné��',�i^�T���&+�*Y��LB�cG�0 ��Z�lX@���M�R?u���?���O���X(��4b�J׆0�:L�F�i�!X�4�	<�ħ����bN����PC��>�l+�JqӞ��Èۦe��������?�jK<ͧs�|a{��8d�����O*W}���i�>�pD�'��Z��%?��������\g69�L5���J�M��M���?��!��Z��x�O��O����r����r�L��F�i�B^��H�*�>��9O����O��D؊i����a̒3�$�j�J	��m�,�ࣜ����|Z����Ӻ����@ ��C�T]@���b�R}R��<U4�P����ڟt��By�L��<�j�RA���+�S�M�F���³�6��O��+���<&ˍRl����hȏW�`� A� �M4�H�����?)-O\���9�4��?N���w�3�P����
��7��O��D0�	ܟ�I*�
��`l�Vl��ɐ%ov^��t�Y�i"`���x��'��	�8)ւ_e���'�6��E�2S<8�0�!�'\�*����a�
㟴�	�4�P�8;a�O���T
Ҽ8K>JT�2(pn-�0�i�T�D��!XD~\�O�2�'V�\cr��T�@�Q��`� M�B 6̲O<	��?�u�F�+lT��<�ORXc�Ɨ�^T�A�W��<1~a"�O&��cYZ��O����O����<�;ɼ!00�ܦ@�ZR^7��o�����I,s�<P49�)��_����aoM�4��H": r�6�1��D�O���O �ɸ<�O��娡e�:;ݺ|��O�t�)94�t�zB�F�(
1O>I�	��S2vK��	7H�.s0�+W~�2�D�O���1_��'��S�x��9%��Ar��Z��i���M7��o�ߟ�'�,J��'T�	��������~�fx�Ђ�*i��� v��Ja�7��O�)�7�BP�i>�IE�	�~�H;��Hs��Yq1�@�=��K�O�`2��O�ʓ�?I���?�*O�dPS�Ǳ!e4�(Qn�^�ܘ�����'������T'���'G|���c�&��1VmD�3�@)��P;'2X�x��ןl��`yB��/��S�	�\��CgN����ڱ(�86����?y��䓻�ep�D�T'�<� �ȑ�%�X�@5C���>1���?������]�V'>�y�&�i�� �a	Xf̀�t�Ҏ�Mk��?))Ot���O>ԋC�O�'7'z<q·��T�L��	������'��Y��EƉ���'�?q��fe�&?�6� �&`�x����p�IVy�I�=��Tܟ(\8��R�2�؍��G�8\1"e�׸i&�	���M�X?��	�?���O�e��_*lߞk�iD66/v��p�is��,Ox�	�	���'����ɶ� qY�1R�	Q(3���4�sӤ@�6n��=��̟����?�9O<�'}���F�P�����/8��6�i������'P�U� '?�	��"��l�D(ЏH�8�h�"ə�MC���?���$yĝx�OF��O�� ��>=�h� AQ�H�2�u�i	�W� � �����9O.�$�O���Dl��� 8Ȩ!X�"	�=}��oZß|�"����|�������!�޿BB�0vM�R	X��_�$����� �'�2�'��X���TCT e&d��\��@�k}`F�I�O�ʓ�?Q+O��D�O��D�&����\�i�������#A�	����H�I���IƟ��'��]{� `>��eE� �(a���T�K54I��bӮ��?1)O����O�$ߴx�DʊwW��G�ԜIa��q��L�*�o�ԟt���,�	ey¯�10 ��'�?�)b8R�Z�lG\��P!�NߛV�'��IƟt�	韠��H�t�OҴ!wc�+� 9.%}(CY(�C۴�?9����l��O�R�'��D�Ʋk�*`I!��(�`��2(�}����?���?��Y�<���?������KH�]�\u W�A�������>�M#/O@\��φ̦��	��p�	�?9��O�nN�_`	ؑCS�~!z��̍ho���':���yR�'��Mܧ:z�LYրQ��4��P�>~tm�����4�?i��?A��|�Iay�dʙ"X����fV�['LpG-A�7Mфc ��O�ʓ��Ox�&]+�z�gȈ),<	�p$G;6M�O����O���@\A}�W�x�I|?i&.��\І���I�x�X��`�����PyRk%�yʟ��d�O���8�*�*��I"~��-Z��X�j�&�o�ܹ�j��d�<�����D�Ok��@���#P=&N8Ւ�QF��	��Iݟ8�I������Е'���:��@K�,v�C�!��,B	;c�
����O��?����?!��> 

!��*_�`xa�U�l�������O����ON�#��a9�ވj���>�4�"P�B�[D�#��i��Iٟ��'���'d	��yZc��Tq��7߶��2M���0��4�?i��?!����YEZy�O�Z� 8���!d��Q$�0)�h�R�i�U����ן���!g���|nZ�(������X�a�`Nߘ6m�O��ľ<�%�`�����4���?��K_�x
���
�Ԁ�2�Y"����OT�$�O�騵1O6��<Q�O�h��.�7^R!��DQ�5��5Q�4��$ ���m�؟���ܟD�ө����~��aL͝$rd�0�K7M�x����i=��'�}�'2��<)���	�.jH3� �t� �R`��M���4%�F�'�b�'��ɤ>i-O�����g����Q��	��5��aR��y�%i{������8��b�'�?�f+�7�8)��ֶq���Dc�l
��'�"�'���S"�>�-O��d��<#�ɚrji�R�Ӹ.	H�� kӺ�d�<���<�Ol��'�	�l��0�0�T�TB�14@7��Ov��Y��	Oy��'��Iϟ�)�.�K6f��&�6ݢs/I�
�p�G��̓�?Y��?����?�/Oޥ�s-���><���B p�t�Ѡ� ,�҅�'�	ٟ�'��'er�fRv�8��� =��X�BL�_4�ٞ';��'��'F�S��� ����B�)#��9!�
1�*Hq#Nՙ�M{-O��$�<q���?�C�<�TFN9)%�VM���c0*�E�Pq%�i�2�'-��'��0aґ��N�Ĕ�,�0X�i�$����S�%M���l�ş��'���'�U��y�Z>7mW5	��=C&E�!$����߭����'��R��	掚>��i�O�����:��Kv U8�KŦuC ,��F}r�'+�'Ԟaj�'��s���'
�2��AC��[zn�����Z�unFy"�E/��6MXg���'���g)?��Y�>.�l�3�H"�E(%*���%��ݟL�4n�X'��}Z�k��j���S疛z�ԋ!GY����U���M����?Y��Z�䜌g]<U9�IF�SA��Ҵ�uڶ�o�&+3��\��g�'�?�V�I5s���� �씢BH͂v���']�'t(PPA<�Iş��U�j�y�i��T�U��+���n�M�	 w��)����?i�w�	¦�7�}�p˛lz ����i@��#o��b�|���i�)I���	[
���`��?4.mXsa�>��m�U��?���?�)Ori�T���7��-j��GX���c�~�j��>����?���ܹ�IҘ������]f���
O�?I(O~���OD��<ч�� -��i�U�̉p�,	�uX�QKuE����'��[�����,���jml�V��M"��׫@���RS��4�:��'���'g�Y��N��'k����
��v��'��R/4)��i�|B�'����y�>�@fV-zF$$Y2ƎK��������џܕ'U��)��6��O��iT��"��ʈ�y	��[�B� &�������P�.r�%����h�t�&�r�n�E�?AZm�NyG�r��7�Q�d�'����??�@S5@ۼ����7k@�5N�m������Wob��%���}�r�Q#;��ɢ�E� p�С*Z�%��!�+�M����?������x�'���&cA2l�1�G̀`<B]��r�@�#�O��Of�?��	�*�P�g�OW����=��\cܴ�?1��?��Μ���Ol�ħ����:B�K$��o:.�0�Od�h�O�U��7O�ݟ��	��*�)����nŘX���� 	#�M���g��$���O�Ok,�Mj<��ĭ�74��A��2/��:̪�IMy��'��'4�8���w�PA�M����Ь�z �u�>a�����?i��<Y>�9��6��;�e�%a��II���<y+O����O�ĭ<���ݔ@>�iۍ;�� JS�	O�8@wG�-.�������I~�����ɇ3K��I�2�5��S��\�H�(9�vD۫O��$�O���<a��Y�=�O|Dj�ԶE�p$��D2V�m���x�4��5�d�O6��X�W�X��*}�b.]%�I���7_r�h�7l�MK��?�.O6�s!
Jn��Ɵ�*]�� ���"��|��0j��i�L<����?ѲN��?�J>��O�z� � RK?��ఠۛq터��4��D^�~�@�o�?��i�O��	�x~Rl��s�hl�  ��3y�e#�K���D�OpiD��O���<�~
�&�+
��[f�N�-_��BDIѦ]ZJ���M���?A�����x�Ov�h)�	D�Q�M���=3KLQ	gӐ	8���O"�O>���.�vȀ��2�^�a�]*�d*ٴ�?Y��?)��^�8&���D�>��d�"K�l�x��Y�gM`�@�)������My�g�cc� ���O��D�"n5̑H##֓#���j0�ӞFn���d�v����p�I
��	�O��OΑ8��� J� 4�M����H+`�U}�d��?����?A��?��o�
[�@]���nn\+g���b�� -O���OH��6�$�OJ�ďH�(��`�u<�5���)VKq�&�T�1����<�I����'xK�1��i
�-�ve-+@1��o�$k�	�����؟��?)�
F}�D�I�J����׾}ۂ��Ǌ��D�Oz�$�Or���O�1�+�Ob���OnTr�nT)vM���p��?�u#��Ϧ	��[������w���%��ؽT�)�,Q�H��!A,�,�V�'�Y���"�^���	�OJ��r�����N��A�G�?"X]�2�Va}��'��'2髎���?�,\76O:�b��A)uل��wCpӀ�4p���in��'N�O���Ӻ� ��Ʉ��?w��X��K>,��Y�i���'U���'M�Y�t�}*�fٿ�H�A1r#�ن���[��M����?����"wT�З'��Q#c�O�qT�X��V1gj>!�Nt���s6O��d�<���t�''���S�]��A���R�>&42�v�����O:���l�.��'���ߟ���`��S���^q����<\���>�pM�Y�����?���^#8�����Y�tI��E�82��'B~m�A�>a+OF�D�<i���)+���[FMѼ]?|�x�e[�G�IrgF���4�	۟ ������'N�UC���;Vw��;�J����!��^�d�����d�O���?q��?aF'�'&����BNy�x�k�O@�q�����O����O2ʓ
��p �?�}���-���6�ѿ8Jxu���ix�	�'y�'�R�W�����)A,L�v�RЂ��qc:ne�I�����ٟt�'���*�d�~���Ab䈄�Y�^i�)�d��� B�be�i��Z��I����\���������{��a���4���	iܹH;N�l����xyR��(Kl���?����fǾa�PRfE��_e��A"Mʠ;�����IҟlB�a0�-O��Ӭۦ�G�B K�2�X"]��7M�<�q"ڱǛ�'�R�'B���>�;lBZ��m�?Qe��j�-ۆr���l˟��ɫ`������9O��>q $�z���2��a�b�B��Q��)�Iǟ��I�?Y�O*�<Q�ؚ�j�J��89A�D�"����iXY	�' BT������P�H�Ӱ�ݰT� �Ҥ�~�AH�i@�']R@������O��I
�p�I	�c�.��.��$�~6�6�T;"(�?1������	-\pb��v��� " �T�8hn�i�4�?�Q�N���	_y��'
�Iߟ�X4=�<��!+�^c�p1��2NAX7-�O�x*u?O@��O��D�Or�$�<�r�䕙�&�# _�=s�jHV�:��\� �'��P�$����0�IO�]Z�g
/����*�un`��u���'S2�'��R�Ƞ�����t�Ծ����v���s��I�F��-�M�/O��$�<���?���z���'�M!c�;L�I����:���O����O��D�<�eΒ#���ܟH!�*)h��*EI�*AH��*����M+����O����Olԛ?Oh��y�gD�8߲Qr�`X�����s����O�˓��s�W?��I֟���=�� p���mHH�B`\�-(�O��d�O�����+b�+��?ݢ�a��'�I��˲c���D.n�:ʓp"<���i�R�'���O��Ӻ�seܒXV)ZM�v�v��V�M���ꟼ�ƈs���	xy���Gll}�BQ�6��= �5S���
�8/�F6��O���O��	H}"P��bs �X��o��re�+�M����<���?����O�r!�9u��x1d�Y$u�B�2��r�7��O���O�)"aB�{}bP���If?��߼w$���T�d�,lsEU��'����dz��'�?����?�7oG(=�yy���"Bp�C��2��'��hY�g�>q)O,��<y���%`	 P�C�ǕF9RbpE�d}@��yҒ�8��G�ϖ�$��Q��
��͓B		�"�t)1eb�<Q��A,5J��`��	�X�P�Nw�'@�Jㄋ	9�p.Ԉr��8��B�)zVXq�i�=h1شp4C+�Q��}��m�WOM/��Qr! "�8�l�+DY1�E{z��b㌆_Ƃx�&R�v5G�^�n�$���wx��q�U�[n\��l�8�0�#�ٔ#Ӵ��vᚒp��)@�	�,p��sƍ�VMBli���(J�H��G�ѿ�?����?!�iYH�}�u��l,��ֵ֥v���A�z��%i Ja�Ds,� `��<��G�v�:7C֒,���E�ط{.��`O�)��cg��6C��w��w�!���?$ ��'�� 1b��vV�(8�����,�@=O6�����g����S���V�V(R^a|B� ��.d*�)�NLa#J�`Z��5���'|�]>��U�ş`�����f�����5�^\�6ً�@y��3rJb�v!��h&�?�O71�bc��x-@��Ɂz�:e�
:6Vt*D�
�V��eh����O�I���]�M��$ydnǨ��V^
����O�S�SM�I:.)h��$��7Mٸ�
R���rB��80�b��f�G �F8"Dl�(IQ#<���)B�B�$z��P��͒g�V\�1����?i�N�F�P�ۥ�?	��?a�e[���Ob�$\�8����w�ݚz	��e�
��IJ�ؔ��L~Z	p2֟ўL�X\�v��kQ9DTi4+J/�?AG�$�V)rgB�	v�p�3ړ%|>��H +������Dl��kD���ҟ�F{�[��J@\����S(yE,5� &D���6G�.��C�i�ha�lH%�HO��|yr�!n�6mS�f?��[���<b�A@�i��5���O��d�Ovy�VC�O��Dq>9�NZ_��iwG�'"	C@�t��@��22�N� ��Ix� �U��)�uc@M2y�r��&����ȧ�E���4�ʦ/����>E��'��GH�(��x/ך��,b ��H�'�BI*�E�:�L+�ϖvs�IQ�'�0\tb�t�l��!�7l�dHX�'�X듂�ף{����'<Z>� NEI�WF����� �0(�x���ב/�v���O�����;ͬ���ZGZ8��k��0G ��OjC2�N�^��Hc�K���R���2k��B�gBx�$�bcG&��Xkw&J9^v��ĭ�<X:1��П|���q�Zb�&c�X������ZU����M���ƭ�*�I���<�	������%���J�h�dz�<�O��$��(A�ԄE��hr&��h���$�{�H������M����?�)����Q��O^���O�@	@��	86(�[�h5��ɀ4�J��@�T�Z�b9��/�i
��'���<)�Cԏ}Qy�JW�79�HǢɘbk�AIT�ŊD���Q��D^�9�eXS�Ͽ+�N`1�"%��q>"�I�� �^ÎA7�[۟x�I-�MS����i=�9O��Da\�QxA#P/q��`�'��'�!�@��%&�cC��bqr����)y�4���*��f�)�4b��&	ryi����wT����'���s��A�-z�1�@�w�8��	�'0�`r���/�ȱ���	�u�۲
�'h�4�u�
v�",�D���o�<�2
�'���r"	4c4��8cꆚY�L9	�'�����"�*��)`�E��!t8�q�'�0c���0~(p#��/�<�X	��Uq�T�
��:�*�
A�t<���$D�tId���-�f�c�,��l4i#c"D��(`�ƾa�FAV�O%� �0�$D�d�q��)1İP�h�7E�����$D����$���^#0 JPF("(B��' �uQ�)O�Xր�� ɈpH	�'�ƠѠ#�%ܼ)B�[�q����'���`��M� �� �cW&�|И�'�*-�g�մ+�Mju	�+ �~��'�v�!wH�,.��PE�ǁ
��(y�'����'��e�dYJ�%�6��,�
�'�9;���
�� �SIƧ&
>�!	�'�ŉ�E�7[���@�K�-"���(	�'"��C��6�V�I�EK$��	�'nN��P�߬
xp���
։g��ɺ�'j^q�n_
t�vU�Ѐ�\b:IR�'$>��7M˥Pv����a��X��y
�'�N!�"��Q��ɰBߠN[*L�	�'���6蓪o<�Qb���81��2
�'P���A&��8�k�,
ƠI	�'R� H�J��d=���AME�'�Mk�'$Z�m�*�l��5b���X�"O���&GL�75ZE�3�[�Z��v"O8��Gރ\}~�#%R�tm�p"O��#jS0
����ԫ�� "OB,bR�/S�h�X��U,T*r"Op��SK[�Amΐf�e�� �"O�HQ�#��t	�كQ&�-_� ��"O���(�8S���6�չ�iXR�'�$iVmǲ@Rx �eϘfA08�@���������S�)�s?�-#�$�B>�5�5K	h��F|��F�a,�������v�cɟv���Κ8D�<H��H��SQ"O�|�w��K����T�"�v���8O|�����iIP�j�o֮H�a�$O1A�d���T#;@�K�Q��yr�ȩB��tCg�:c<��F�׃_��j�'������B�<Yȟ��4v��I�EW� 0AٍC?�1���O���䍏#����&�UQ:�SR�ӜTЎ�CN-}��b+��'�rq��ɶs��;���
�p8� O)-S�#>��n]�|/`�SԡC
��O[t�K�aH2Ɍq\?F��X`��0��a�L&�Ya�NV=U��scLN��|��2�t�5�=3��d����X��'h�ZE�f��B���C���R
}�ȓ�h�C��V�r?�ƤĻ�n0	ю��<iw#PhDZ�)�'���A4Or� @��6xH\@u.�kr$��5�'\��#�����EFX3��7�٦>dT�X�'l�epK>�	݈O�Y�g�G(a�^��CMϸUm���b�I3/���H��ѩp��Y7�,�D�6�δJ&KU2Y�IŚ�0)�Mi��� Xh���*��]*��� Mb�H�<O����ڧf�H-��F�0���~ʟ6xa��πԩ���H�!TȠ�"O�䋀E]�uLL=q�gB�beTl�`�I�P���Cr6$i��Y��1����A�a�E�2�F�"5�İ��7�O�Q�@+�}���98�%xₘn�X��0O:\��|R@ٵF����GF>5 �i� ��c����=�V���'�5I�Ҡb�s�4/[�g��P I1w�|	0u�U��yR�0?�G����C��V1>�X�����<��P> �~5�3���;�!��ә"�e�����9sT]J��ɒ����c��`5ۺJ�$��PĖ,l��q��<�K�)M|��B��]���d�B@��˂����}(�bą�!�DYT�e���J�2�rE��!�R"�*c��V넨�C�K�)r!�D
U`d�b��'�Ҥ8��>T`!�Ĉ���J�J��f���G8E�B��z��1��(�cP�(a.�4s���$�6{�,�\#���X�@�9rԉ&D\�Mo��
O�4#4��F�$ ��Bɫc�R%B��I4:�����8H.��|ʇG��|�� J+�[e�@v�<!"+K�O[��s�]:<@Ȩ�Q��ן��4e :�̅����xy���Ήv^@�Ѭʿp\��Wj��8��B�I"�hH3�Q1��$O�&���C�p$b�8e��b
Ó?}@1�H�,¤����5�R��	�1�B0�S' �	��Z��_6o���!��Ò_�(���Ni<�vQ�
>��R��f��E�c[�'d������D������J��h.��A��,8�0�]��y�b�@�@1��,�3W�=�6�D��y�1=�2b�"~zBA����
��R2M�"�z��_�<a��=��b�G�,Y
������[�<1�/O2�ԍ����(O����kBa�<y4�@�
.�Ԫ� #��(qf@�W�<)�$��F@qan�ȰD��\�<�+Zp�x��ǜ����m�[�<IgOX,r;�p b�
!Ԫ\Z�O�T�<�p�D9V��� ���/j$�5-�H�<	1@[�S�^4#㔞J�f��-�H�<�H!;|dX�@����c�G�<ys �H�IGB�X!J�rѾ�y"d�k��1 F�^�0%p�1u����y�C!�q��P%'�$��7�y2*B"v�� AD.Lo0�4���y"F->l8&�FX��	A"X��yg�*,]�mzp�$8B�T ���y�B�,� i#�I� ���3l2�y�)��,����P���큕�
��yBˏ,�,�R��<̌]rkR��y�+_7nV$�K�'8�L �K��y�
�&�<a!�>/��9BA��3�y,�60��q`K:9��1��^0�y�O��tX��B��YYda/W��y�A�5\��O?ac4F�1�!.�5J���8V,+D� #�&zp��"+�J���o)?WIN&Oa{�͓R��0�K\�A�v�0�����>�g(]��xl�=�4����d�aQ�Ʊ
�PB�ɵ�"�գ߾&z�X��.�&�"=1G��24Q��D�4M~������Ȕ5 B�Q� ��y�n����t�F��~qfh�p��:�M�2Oʧn��<E�ܴ4_wꃗZR����κO�^���H�@�_O�P�� �C�	�'��&k1lO��2�ⅰ5��P��<���Q�'�j����))H�ULQ%5_N�ؤ
Į]���ƓID\��1'UN7$DȀ
]�~��ɾ=!�Q�?)���6�F	2���BU %l�x�<��"҄V�E���UT���ՊΠz�"L�I4=Cʤ��
�-�7����� 0h�ןQ�t��.�`cM��"Ot��D�jg���K�T��`A�JG�<�r.H�� �	�$&h�Ώ3IP��t�KZ�y8E�)�x���)�+-lO"pG�uE𤪰�Iӊ����?}��5Rb	
:y���2��-�^���'BΨ9Tn80��}�q�Ӛ��$Џ}�.�{��;��H� @9����9.��7]?��� ~�
!��'..����6K�!��&SX-���h*����k\ �b6�łOZ`�@��y ٺı�O��ع�=�а��	
 ��`�t��qOl$ŭ��t*��Љ?"�L9�NU*q���dQ�b/���%֤3(Ԥ����?����X��F���C%�+ ������5,O���B��L���E��t�V�CQ]�D�Pi����_[���-t�P�I� ����>I��@E4��h�1/ʠ1���l�ɾ#ޔ@1fN��)Tk���'A���:�����\�lA9�vj�\g�Ai���y�l8�a�T]�U�B\"u'N��P�˂�+5P�Y#�5r7�%��t��}y���1d^�GIٙ%C(��pF.��x�a�	`��h����'�ԑ�gi�k񨨑���&;�y�E	V�L���z�'����5+����oF;&�H��
�*��,�3�Ϭ6�z��� [� I#��=���ӬƥC���P��d��|�����#��^��SV��M�'=�,����	-�@�_z���S�1yj�\��$��F�Rщ� Me�C�I�hpV����J� ��\k4*�oT~t�o�LL�	ԅޕ�?�B�7�ӈ 4�I:��]��y?��r���C�pC�	�<}��rR.����!��ׁ2>$��ԇ�geB��e�?"�~*�KҪ	�џ�(��;ܐ�5&�w�Y0��=,Ov�#�c\*6o�<�dhWXź��� E�u*d�Q�W2������.?�R5���~k����BKplh���<�&����@�-j�y0��S�|�4�D*=P���ɤ@xB�	�k �����<O��cv&�).��*	j�I6P�R]��O�4I�o�P�|�"$-E&R����"O�]sG �76��[�N�_��`�aN�7�2ya7A!�O�u��U(Y�L�Z�-	 �LȂ�'.m�@�h~↖4T�t�� ʰ�^�P�@N��y�b����"�kJ�>0@���yB�ΰk��D ��`�bb���yB�F�8��4�N�(zb��sB���y2��S`�Fm������M.�y�#_	H
n�2����a�����yr�ق!-���LZ?4 �㖣ۮ�y�7\`IkB#�r�� 1�S�y"b�tp�e���-�@�����?)�b�px�A1ĩ["NH��i=��0�G���ab��e�����	�p�L�9���=Q"��jMW�� �?q5�	4g�T����H6Y	*��D)�%S�zy����%�xrE�v"q��'��P��ՅY���k��0*p0-Ov��ǯ�<^�����U� *��(����"ph��P�~�XD��WJ.C�ɧ]��R4#�~�xĪP�.kN]
P�X.A;�젇�F�}`��fD0��d&,0hT�� Z&@�C�Ɂ'g!�d$(8�4�毟5L�6A�Q͕�QU*Im��y��n&�|���'���ʀoA	t&� �${����d�<E��X�f�����]8�	*t�L�<5n�:�X(�GO蜰aC'TD�<�W���(�\0�b�)��!hs}�<�4"�n���]�k �)�G��{�<ɢi��_*P��O�ari��u�<�� �x\�� &��c���*�n�<�ĩ� h�z�ch{��z�,k�<aq�Gm��B�	<n��x���N�<���,!b����X.\ذ�mI�<1���|tL!v�Ȃ�0�p�gZ�<��@����������5P-pDA@L�<Y��
`��C���l���5�OH�<�5���f�<���OMA�uC�G�D�<�1�$&�t�AEO�(��܁��v�<���	'���I'��
*�Д�ao�<� 0d1�@R�zz!�EB�`L��"O,��a�*ߜ�s�M�(O����"ONMc��@-+���Lsg\ �b"O�E;�	Σ'�p�V:Sh�ܸ"O���F'���z���-D�<�*�"OL�q��*E��u���_�@��њ"Or�P�ˎmش��F��TKV"OIb�L�< �:!k�#�D�#"O��� �<�F���:T݀��e"O 0hrȄ�SQ4A:��@�3ɴ�E"O*4���"<�dh8�O�<?��E�g"O65�£F�C�dB�n�/�.\t"O�����~ږTyt�bR��r"OB�t�M}�l5ʕ"Аm�Tj�"O� Qd�@�$7�H��@E>.iH���"O�M��	 �,�*`@W41R4aBf"OVY�A�A�B�BA��H��pC"O�#�A�&y:UDF4{��rP"OjhQa瞂GJh�`$Θ%��Tc"O8ј�"�:��4Z�W� ̚#�"OX]��KB0Z2	{��
�Y��"OQ1�О�4=�lڥB&�+w"O�]��c،a�:���J�R���"O�8�L�#aK>�cף�	*D*�"O���ɖ!uA@Ta��Ƀ"O����)]bTq�X�9�Z�"O\�)�g����;��M�ΈA� "O�!"u�T�_�.9�`�N��X�˃"Oh��H Y���
���v�J�"O���|G�kr�Q;���G"O��R���Hb�^)q�<ͳ3"O:5p��;̨����U�b~�ر"O����F%C.4i��;a�e�E"O$y��嗴J,�X���F.J0��ѥ"O����(dz�t�`�K
[����"OL�	E[�)���i�8m� �5"O�
@NEL2�h�)R6d01�"O��x� fJ��è�(G��q"�"O�Ia�ā<^���B��D�.�5"O$y�P]k=B�K�M�����"O��F+�<	���\�(��d"O��k�(�b\����[=���&"O$�+�'4m�Q"۾7��|�u"OB0Y�F^�#^�@'I� A�"O}��-qHYAp�ݓg>}+b"O
I�J8�h�CG%k\T� "OX�b׹9HqA��K�Ns�"ON�b�N7��" %Q -j�az�'�t,�1s��1j%��[�֠b�'��=0�bD�yhٴ-��S$Ψ[�'�^�	 �Rˊ����0E�>�c�'�欉��\�CI�H�#C�+PB�DX�'!�Y��MI�2�@l���ƣ~,`��' �t����bO�pc^�qX���'Z��CЇ�R/r1�%X�f��l �'�����/[69r@r���Y��yR��0}0��T	
}�B1�!d�;�y��/j����B�m-@�X�gD	�yr#P�?|�k�
H7hZ2��� ���yNF�~�2Y��EO�ڽK�N0�ў"~�Akje#�bÁ{�4
a��.KX��ȓt�V$X�
ˉ4�Hx;!KV������z���i�4�Bq;�<T��ȓ4�F k7e�lZ�����2����?����~� )�"�I�ذXJ6�����"O�kD��2$]��pD�R>&�R�"Op�����/�����C��'O��"O�ܸA��t.L�pq�i�� �\��y���� N48QnAJ��I2�n�y�h�&\!A��3I��v@B�y���+k�\�R���S]������PyB�A� �4��Η�D��� OY�<��LˤH2���>��p�NQ�<!�g��r=�xH�F������M�<�� �(o~�����#l<R���O�<��BU8j�4�2Aa��M��Dv�<��/�%��3�`�άc	�p�<�3)����qDț�x42���l�<�7ꞹh6�ҀjY�G����i�<-�@� �)�v�`TJG�_ʊB�	h���i�F�A[ZD�R*�M�|B�	�}��\*���`�F�k��T�U�B�	/d	�Ukv�ѕmdDX��
��B�ɀ d�(�$��=�`�4F̖ �B�I+2f��'�-����w�J�CbC��.D�luY�/��
8�x���5K�C�I6b��"C�>�hf�:m�B��%Xz>H;d'T"� ���烽^�C�HZ�)1��!X����9N��C��HU��	ڼf�J�p�N�>�C��0�0��!�E�s�[�y'zC�Ik��:S`�2=F2u��GƠA_DC䉐VV���A��q�4��j�'Z�pC�IW~��W.�D2�s�ܟ@�2C�I0&�����
 Ϫe��"�0K��B�	k��H̍�fx����X�Y3�C�	�"8B�i�gLCv� ��ʎM��C䉄8̼T�U%�{�i@&T(7B�I�y��+V5j)4�JQ�3��C�I,r4���$�c1��M��C䉑N���EJ���"�ɉ�-=�B�A"x]��%Y�)s��x�)HJ#�C�	Q'Z���,�������ǢR�FC�I��ibRȇ�~�Z4;E/�+w`jB�	K�mɢ�5g�24�'��i�
B�=w�H���<.tX}�1h��C�	A��ɂ�!x:�
���O����3?c�E�ݖ�]��@�"���m�<���/꼈���?2CF�J"dc�<Q��JQ�ͺ�%N:� ����H�<����(`�Q��T 8aJq.�D�<iE����`���I0Nx��@{�<)�
p�T�Pg���pU���A�<q����-�"���M��!�CFc�<�ag��J�\��,ݛ����-�C�<y���,i����ǝp��= F��}�<�Tf��W��qʱ%�!"�Ό�0nCx�<#H/<�(�EX�Ic�i���p�<����
e�x�y��e4�J��wX��Dy҉K����4��+|l�A�+��y�A� {6�S�oP�{�����ٟ�y�ťZc���M=H���6L���y����U����";�*��aG�y�o�9C+�u��΍�7�<˵�*�yr臨8h`A�d�%m�)�#��9�ybF۲!]hȀ�өq�0��[��y�L��VR�!��
]��j��A!�y"�F`c������Ia /S��y
� l�ٶ�@5A�D1a�]	�`e��"O�m��G��*,2S���j*��"O�l SeJ[��<���m���
�"O�ɲ�⍙i��a)ㅅ��� [&"Ori��ќp|JA��N���oׂ�yB80����r؂���-���y�
U8u%b�ȕ阔h������yB�����T���ǚiW���Ц 9�yҩJ�M|�����0@4=�'�H9�yb�X39� �b4�Ku4ȳ�B0�y�k��8[�K 
uR�LF{+TI��O��=E�cR:m��5��%�64Ƣ|�$�y"�( 樹y�o��|��\[�k�	�yRoP.0����C�g`��[ņF��y�D��������:X��rd%���y2�ҦwBޔ��&��?(J)H䂁��y���)4� t�OnRX5�sl�*�y"���U�\��P��;_SfZs	��y���# ^��уպa�������y�C`�8qɶ�T�6A��W�y����|�J���	U�`��#���y��/�I�'dG8�
1I���y�GC,dm\�ٔ��41mt�z��Ԧ�yrM� ��i�� 89���S���yBDE+~���gA�d���3�+��y�\WP���F:5:�y�V�)��T���9�t�`tG��yBjX;:1^�C��6�v-I�+���yB��C�T�� �5����Q��y2�J�G�S"9��I+��yr�O�_<h�F	�b�����yr@�&�V����^\��@�U��y�O)&4��EhL�i�vP-҉�y.�7"���rD�0Z=|q�'@���y"^��$,2�ߣh���(��W��yb���f�����3N�PŁ��+�yB@Z�drF110G�����*ɑ�y���Eb�ӁGY;����G���yB��na�a�B�>A4QbG-M��y���^��r�ѵ:xF��穜��y"C�Sک"l�v�=�����y�덅�x����"h5A�����O&"�Skڂ1䖩*f+�6e�����ZB�<ī��>L��F�<��C�g�<�k
:Jjh0stG�"����"�J�<���M�a�|P���a�=���C�<!�'G�o�X�#F�1(�V,�@Oj�<�&Ꮈ+�D�h�**,유��m	A�<�J�<B����ˢ� �� fX|�<)T��qN�#���xL1���\�<!c�X�K�l��)�q˃�LY�<���S{��D_�I�\�k�� A�<)�fL�F����@�&&M�b��|�<�"�/#8�L1��\�Nq(��O�<����Q��]q�,M	H�D�#�u�<9d�V�'f��At�H�I��p1� l�<�U��d�l���C�'�)���|�<��Ɩ�JJ�$@�!r(v����N�<���.��@�S�H)�0� D}�<��ᇑN! 3dm��qg �s�-�x�<i7A
J�dp�Ѓ��K\��C[|�<A��V�0g�	S"M#eJ����@�t�<1�_/MBL;aں!�z%H�u�<A6�=�H�S��3t�l�� �t�<� H� q��'G�5�)8��Zb"O"�2�݋>�p��VH�	Wk���g"O��&�3zy�`Z��[+@.���"O�\�$�L&9� ��eH,Y-H	�"O@�����OvJ��9	ڍ�c"O�ɠ%��l>����X��J%"O��	���-�OX�9C."�"O�5x��a:��@��CMdeJ�"O*��hU�I�MZ�z�XX�U"O����Ǯ��T*�LȀ&��dQ`"O��PF�5`3n�3� �Ws����"Oԡ��%O#$$��lRT9Z�"O�@:5Ɓ(����q.#B yjP"O�Ԩ����.�5���b.����"O�}�5�2|�X�$��P.���"O��g�O+Q�V�0��X@�U��"O�uR�ώf���@�8����"O��``��k2�����K���6"O�5٤;?�����)�KoH�k3"O}���JA<| Ň� cj��b"O��{�cP"uE��`�ty��"O
�3�aA�͸0�}��H��G8D�Ae%1�:�� N� 3����`G5D�̘�ŀ�I�xy�)�-S2��0d5D�4:�"�h�	��W;:��B�)D���d����axR#@�r�N�Q�,:D�h�`�K3Hv���p�/5��L2��9D����*7U��P��҂(��Ȳ��7D���P�S�lq�AACP�v���i D��Y�́h��1S!BZE�̰��=D�@�'EV#M�P�@��"h���[/)D�|�����3�d��v��<| "`(D�txBK�'V��e��$x���PSc$D�����3��LѲ��D�j���#D��s�B�7r{��K�B��+8$qu� D��:L�2z��ɠ�T�T�Fܹ��;D����"�xx!��R;,���,%D�tjG���U� ]Z���:�\�(�.D�\z�o�$w$D|�@��<��7D������(B����;f�
8�k4D��ʶF�c2�Qt�BX
2٘�3D��lS�A��2�`ԎUV\ղ$�2D��!�oJ;?�,� "S�>t��y`N4D�,�&���"�Tx�!Z�zd���1D���%e�|�x�Rgl�h��ǁ"D���#��V�$���:z<,T��>D�0�'�B3_S���dOMh�>�M=D��P6h>'�^u���K�=�t`V�6D�d� �H�M��0�B˹(3ZĪ��4D�4�V�Ӡ>�:��V�-p�̛��1D�x�"^H)�%Sc���	����B�"D�8��3�n��u#��%z���?D�H+��p�v�t.r�5���<D�X�2+�
69�׏N��X�� ;D�0 -Z�%¶�x3"²c�:D�X�WhU,n�*)���Lxb� �6D�i��� ��ɀ4a
*p�6�{�5D����'��Sِ|R7��!"�Lt۠�4D�ܘ�Ĩ/l�87�R�@@�C'I.D�P����'|���U��T9�a�
�'��@w*m{Q��bI�B�B��'g�y�J;O��	��·Q/�I��'{Z�{"�ĀIrP����G����'���faI./���a�+��`i��� N�cwmѽh�60�U�مF�\�"OȘB�B�Z��u���9`ݙ�"O	��hE�6�(2PK�;/���Q"O֕Jv	���)�u���Bڂ�p"O& �pi-A�t��J�ȴm��"O�L�M[���yh���:$��#4"O��ä���9�
����TP���D"O$Pk�*V���DمXx�J�S&"O$��S,!L�L�ӳ ����$��"O.��I �!p�[�V�%#�"O~��G���4	��(\� n���"ORȑ"��J,ʣ�q9�R�"OJd���ԉ�۰EG�(n�y�
ҹ�8��<*�e١���y��!��k &!�������y"i��_y:� ���M�v9`�mN��y�,�50�<�*P����a"�ǅ�y���l����a`<i��
� ��y���6���H��@6�T�0-�1�y��E�(�f����PZ@�YP��y�!8�b�CD�NF\��0��7�y�N�֑[+T
K��\ �	D�y�̖�г�B�!�J�8A@X��y�͜V�:�p��݊8n���C�&�y���3Rz6 I�NH�0 ��$���Pyr�P�r:l�8��Ϫv��R�N�j�<	JՑ
6zɃ��"%,QYU	_�<!@E�w>)8$oN�U���EY�<� ��*�2����A�O�(��iFU�<�sA:.��X�B� m�e��m�<�'F���� �ڽ���Kf�<	�1>Y X�C��=и��HOd�<�%�ǡ=�1�$郟|�ҭXe�^�<!׶`��0��LW'�(��A˚]�<���T�P�,���@�FM�4'^Y�<��m����c��?8m<`�A�<IRN����C`�A=P���#�c]B�<G&B:��E1��=��ۓ��w�<�0T�k>�[a �iz��2v Vs�<h֦+ۂ(�h�'Y��XV�6D�����	6(�(5)�~����A�5D�pإ�>;��S���#dZ	�C�'D� �0�_�v�,]y�hʀq�\�`�$D�4�Ǌ��R��52���P�ǆ!�$˄\�t�����Y�j1��$v�!�d�y3~蘃-�26�]3S�7t�!�^�&  C�E
�Y&JAbg����!�+>m�,e �$�< C��t�!��QaZqcCE$.����E���Nz!��B)'��=)*�9wZ�	�&@��PyB�
dxqp2��t�ȉ�� �y��~�ˢ��n_~��  �y�n (��l��,�T�bT
�G�2�y2��e9�t�¦8��u��yb��J��a�.�_��dB��y�I�A��Mp4��!l#���N���y�4(R~ �3fE?��8�F
�y�o��s��E�ѧ�6E*����(�y�`fikfaS������:O0$�ȓ�#�+\<Jܘ�[F�V�m��Q�ȓ$+l�S�Z�)�:hSR!�s+(��M	��"�СwW$S 
G�y��(ܰ��T�����MU11ƀ�	6"O@p��.7~�2���/��G"O� v��&�΁z�up�e_�#�NeZ�"O�4h���6K�h��B}��;�"Ot��!��.l�@!a��sn.�°"O��Ơ����Ʈ1��ʡ"O�$��%w �HQqH�,N���3A"O�-��f��l)�8�ǁ�C�9k"O� q�'Lm�lT��&��n��"O���pEڢ'��`���6��l1Q"O���B�1R��1�1��)��9iC"O�e���I�X;��?�t�c5"Ob��F�=llH�!ƭ
W�&���"O�<� �'Ȏ��֡�)f�L ��"O�Cŋ�V5H!��Y�^,�wO��q�!����A%fX�`��-<O��3�1D�!�w�ہY��YQF�"�B�	&s&n�{Μ�c*qx�� M��B�I�"R�K�(1`}���#%�B䉆Nxv�3Վ�--*@��f��A@C�ɴ�t�����)n����%��H� C��;+������7�
��Ђ�_ C�I�T%��+�� �9�~�	4T�2F��E{�|b�)���!k���\h�����D;FE!�\^�e1A.QKP�9T��,T?!�ѩ���{�m��X.B��u�B�C!��[�^�rd��9CHq�!��2�.�rF	V�^�����ʖp�!�D�j����橖�'���0d�� �!�Ğ�\x`�i�k��!v��3��75�!�D�=3C�3�j.||�3�*��!���}A4�"I��{�,�a2�^��!�D׊�t��\$^(����葫7�!�$�1Ab�ԯ�r�0m�`gD�(%!�D^"E*j���$�4�֡�S�+!�䑙3��Tym�S��%р�Ú���$(����a�>����
PB�I:�ȐR��F~&�R�$մ
�zB�I7��(R��ϗ|�}r�.��"�B�	)!��ձb��pJ�l�G��QC
B䉮��qq#�)a��8���O���C�;xҮ�B�woV ��c��e��C䉇\ � {���$&z��v-̌l�C䉾7�0��M�6d�b��ɱ���d$�Ĩ<I��d�w�����V�XZ8U�D)�q�dC�ɰ<�m1���0��@�=#�<C�=H�Z-X5A�8}e����D�F�$C�-��Ɂ�ŭE��py1���4�>C�	<����c��6�Ԭ ���%,6>�=�çX�lH���ȥ3�HA� n2�'����ן���""���We�lȢ0�į�uǺ��8�Ş��dL�D�|`�w���]3F�ҵ�^�!�$:	8pW.�`���[g'���!�$�F�<�Q]y�����ul!��G/#�f����l�J��+g�!��� �Ɓ��G�C���0��|�!���$���RBf�sZp�S���S��O@�=���L�S)Iv�ŁfI�
�д��"O����A� 7Z���È76��A-D!���CӼ,����q,`B��C�!�$D��:Wɉ8�����!\!�D�����JPހT�����1�!�{����H�a��Y[�U�c�!�ē�� �����:��1(4�1��'�ў�>�8�%�,rj"�%D��{zْ�"7<O8"<�r��3=~q+'-��C{�B�Řn�<� :8R ��� 
�HsI³4�^�R�"O�8�,��QQfePf�X�r��t"O6x���,�k&E�a�(�yq"OfA����=F�:�����/e�Tݹf"O��a��[:I���ʂ���!@"O��2��\]SpY�a�	��gr�<a���&o*�����6X�4)���kx�T�'{8L-ϛ7�NYH���C�\���'t<��J��H�B��e�ǧ=���'#��nٖ�BP8V���=�;	�'�01����-�y�O35z�xZ�'�<d���]+JD2���DF�1UxȘ��$(�'T�R�3��	SșKî�);� ���vL0s��B���E+W�_�@z�܅�hִ*�-�B�PMx�m����3���J#k	J���C��@u(vC�	�u! ĴV�Ű�N+Y{0C�ɢ1QN�U�8خ�A�G�f�dC�ɸs��@ɳ��LO��ȼBc�C䉱x�X� Uk[��|�b�X$A�r�=����?Y���?���?�e�f�"�"���:�VCU5�?����������"�Ġ\����+>"N��@#D����ξ~���`�յ*�<u��!D�,���^�]L��QO?<.թC�?D�� ��H��	��!����-#D�<:�a�p1z}���'0#b�K#D����m�L��x$�����0WO.ړ�?)���?���?A�TH(�Pj�e���ӯ��&O������?Ɋ��i¨3�h� 6h��z��h�����pC䉋m�4����6^^���c� MjC�	�&���H�
c^�tR7$� 4PC��(6,���"T������*
�B�I�$�t*�k�*49� �B�ۂB�	�h\ �a H܅x�z���I�v�=����?���?���?�!B�//�Ġ`g�-��	a��]����hOq�~��ԬF�0�cO�l-����"O,#��.'z ����N�i��MzT"Oج�RÆ>C���#$��Z�q�"O��Qg���hiK��A5X���P�"O�S�3 ��h��}v����-����G�	h�:ݑfö\oh��06�}���R
/x�E
B�N�����@��I
�2R���ڜ'�ԅȓG���_�7�P3E�� ��p$0� ƶqf�0uj�,v��� s.T��5B>��'���<�Ɠ��8*�e:=Kxart�՞[r^a���x���+�&�(��=��r��P��y�'?ؼ�@�G-��`�G�$�y�)��6Il��T�m��Xc؄�y���<sȉɦ,��/�8�څm1�y"�X:^�.(��Ī:�P�(bE\;�y����)��D����<��ɡo���x��
b��š5���A��5!�d�B� Ek�,M��ҁ�4�џ(G��ə	�~䲡�H�i�2A;��ٷ�y�*� �0a�P�or}!�c���yR�\N�P� 0�ڊ3A$��a��*�y2�D7'څ� KI�T���g����y�	!`6�5���N8inŪ׌T��y�ʀ?�va��c^$m���I��y���9a�-���ޔ�f(��a
��y�F^�u��q�i�x#P�A�O��yҥ��.����H�]% �B�A��y
� ��5�D�~S
��A �,G�q��"O�{4jC�+y��SH�))��H"O(��p��*vR�P2�V+$��,b�"O�V�E��,cd�Y�.�,I�G��j�<�Ud޷r:��� W$14��AwfGp�<Q�@�V5n��.��tAă�A��ݟpD{J?�:R�>y;R(��B(�l8�*D�|0@�=P�
�pR��k�01�3D�l����!�i������+S�/D� ��a�!���v�P(D��t
�I/D�@��GQ���Tq���k�g2D����kR,E�t!+a�"*��C�1D�8*��V�(�X��@>!��=)Ê3���x��S�=���i"�V�N�ح�f�Y*7�C�ɖq�~!*�JQ�`4���MEj��B�ɠ+p�Q���se2���-ȃ8�B�ɞ<��([����%b�	j̢B�	(U\�����X5����B+w���ţ|�FDX�o�i���@��I�r@!�dW��R)2����	������1d_!�!�`���	\\���W�^O!�$�5������^�}�Z���l��;!�d̻ �
 �qJ�#Az��!��j'!�d��{��9J#��$]T,)e"
_!��2d�Ω�G�c6P5c���%+�!�$���h@1&bT�o&�2�~C!�F�/S"�P-�^��M#Ό� =!�L�cJt��`�<��3 B�(�J���r�A�D��z�!��y	�Q@5�7D����j��cW�!H��Q�jn�bek:D���T�A�fdd5��+7r����!�<����S�C���3�o_�sx�=��c��hFC�Ʌ&ɘT*ъM�K������E�nbC�� 1��𬏪$~Μ�e��l��C䉨^H*��� 4�����/Q3]��˓�0?1e�����UDӳ!��ȹ6`�_�<�F	�@����"���&\���N�[�<���;.ʲi��W0e���a@�o�<�`�I�p��4s��^�z�mZ��ny��)ʧ7V�$��Ɉ$]�A�&9MԖh��-�1eK�'d�<�PB��.+2��ȓ%�%���ޤ)-\=��o�J$����	%T"(��G� W����J�q�B䉫H�d��ӌ܍r]����28C�I�5��lpq���O�^�T��f4JB�Ic��k��ǔukJ��'$�:��5��o�O^��� 2�$���?}�D�b�"Oҩ	&mK�hѨ�*�3%��Uڠ"O矠)�8Z&ʖ'H��	�"O��Y��R�yRCei `ya"OZ��4lQ+o�0���Ƒ-Q&�'"O�!��(�Z�=S *3F4�QU���IX�S�OϾeА�
/(ruUk^�9 �-�)O����O���>�@� #c���av%��@	�k 	$D�p;AN6(�4J���Y�p-�Ө"ړ�0|Z@��]U~8񅮌HjȢDBk�<ل�3����	b�0���k�<�ԅߖJ��iꆥL6'U}!E�\�<�L��N��%t&�19xAС>?Q����<`�̙����^�N�@��{&L�<�I`�T�Ɉ�~���y����9��|��C�	`L]��7�-����J6��\D{J?͉�G0lN����P:�hd0�,5D���O��(�� ,��+�2$h�
9D�� <� 1OF�b�8w�8,��b"O�1�Ǐ`����φ�h�a"O ypg�æ)E��`a.�� Ъ<��'Oў0E{b��Ny����T�Ŝ�j0��5�!���:HX���A���Mj4�P�]ў����+WVuµ�T&�Q�/�9�̓O��D[��*LrƮ�o�{���G�!�ǿR
њs�K7@ȂVN�Y�!�Y(d��qb0�5���!򄏯�b�hf��,m0@MS,��DP�����+�V�˵%�yO �R��F�$4�Ich�6�hO����&ZJ��r��!���J�V�SK!��W�7e|�Y�m�4<��h�`҅w�!��̙Yk��fjӮg��0	Ɔ�"4�!�iv�����+xn\�d�ĭS!�DC�IS��IҢ�j�xd�@*U;n!��n�,�R��<N0�ҥG��=!�$R�t�tl��;zA"�a ��!��C~�L2CZ,- ��Y7j8\S!��Q]ҰZ�)Y�z�N��4<�!�dV��8#��K("mta�O"#�!�ʡ1F�%�2��,S\Q�a���!�R1*9 AHխ�
#۠1�`GkU!�D�'B��0�T�C��Iz� @T2!��ĕl�.)��,�5?P�$�鞠U!���؛oU�[2)��B"|�ޅ0WVC䉘oH���f�5(T§���pVC�ɫ:[��"-"bi�B(��F�<C�	�F'��x��S�'.y�`��0�JC�S����u$�q�(�A����0?q��G�c7��T��&�>�3�XX�<�����$�g�r!\l�#S��$�Itw��x�.�4O�L�f��P�|�����Ӏ.2�����d� $�pT��46L��ّMJ��ܘ+h���ȓ'� �A�J!No���/Y�L ��Ho&���� ?4LptZ��A�؅ȓF]
	�6�)ɒ@�fծ;s���l��1��N�Vu6�;T�ÕX9$܆ȓbf��r�*.w�<#�b�P>��ȓ}ð<�'�;X���C�$]�H`�ȓ+Z)@޾d�Z�c�Aנ+g�]��,���� �4?�KS�["S̈́P�ȓe�L���Q���s��L����M�^ s�ۂ~"q�b�M�4#%�ȓ{�V< �@֊}ݎ�r��O�
Շ�	E�'R��4H ��nʙ34����'��`�)]��|:dɜ� �Z1��')���M�, y��c��=ӘH�	�'��X�1��^��qp��	�G[����'�<5X�A�CJ�9��Q?�`�M>���I��n�-�$JY(E���h@���{�!�Dȵ5�JUꅠV#	�| г�P�F�џ��IM�O�Ped��>)����j��`�'�\Y�"�#Md�)�d�X�yu����'gl�"AN��!R(�0F-F̴��']��c�  �lHL�O����	�'�����Q�HN��KI'>Jd�r�'a���"���/��9�E�0B�(�c	�'���  ���|iKSHC�8ͮ��ߓ��'�=�a�ÜO�n5�s �,%�Z���')�����Xc
�{F����e�'��ҷ#�z{�	���9i^@�
��� �0{���CK2- �2@m��٠"O�1E��'L%�ܰ�(�-o�"E	�"O��P� �$`mT�pqe
��Ԣ%"Op�����."� 8�D�v�1q�"Od ����+`��q��C�j=��"O �h2A3|V����ߣ��9Z�"O��K��5��{1�6�ҍ��"OPZQ	�ZR<�+�E�<����"OZ�ӣ��;m�P��oG*E��$�"O i�I�5|����-�/2x��kv"Oz��&�hŎ]r -��8<�+r"O ��%�S!Yf�)33���
n�9E"O���b h�t[��	
�d"O�-p ,\!WK��0��X���"Ot��J=t���ٸ�5R�"O�-��؟b�&H)�E	S�,�ʁ"O�Px�Ϝ�q��0��͋���	u"O.��2�o9č`,�"U�����"O�e*F�U��z������Z���"O<l�t$эmL8�?���5"O���U#y�H|���5	�,��"OP�s�!�� �ct�]/���(u"OR-�f�2���6Q�"�xRV�!�΄\A"xZa�lFLQ�'�i!� z��)��Mu���u�E!@f!�D��JbӆS1Z�={w�1
�$�4E{���MԈ+M��c�h��i6^�s�b
7�y�NS�1�N`����"c�fXbG��y��p7*�q9Y���Kt�K6��>��O��j��بr愽 �	;��d� �D�O>����#���j�Q���̀�y�!�G?¥���ו�$eIR+��-�!�d��@aC@CO�	���ˠ��?0������?E��[3R�-�4@�Un�"�C�yr(��i�6���+W�Pj|%�4�G��yB돣a�����a�	P��M�����hO���<M1|�	�	�-�h�i�Xg��`y�'�?qcÊ�u���7����h�AB-D�0馊B��>Y3�FI	R��@�0D�\��/� ���p@��3�(��.��1�Sܧ=�17��CҤ,@�HD�Y�����n�	�)�(k�T�3�	�/T��Wˀ����K����J�C������r~��2q���,n4�#��)�y�/�i���4�ǰ= �DI�nљ�yr`ǈS[
a�!ʰ#�li�s�F��y"cA%?,y��I9!��m� э�y2.ҏ=��ѥZ����@X��yO!`��e��8)��5P��$�y2��"����8Ì@�RL��?������'�7O�X���H7u��93�\!p? �iS"O����2�=�p�RS�<�2"O�1 �m٠T�B���(YnE���"O��e�	P����VED�>��P`"OԌ)���l�}����&N��d�b"O�UB��
Y�P9H��	\����"O��ԣ�k@6܈F〉 ��X�[��$�4��C���'C��]�B,$�@�^(d��`̞@�jC�LB��	nV�F�`تM�Qj�B䉅%�8�ԅ�9B�&hC@�S�LǊB�	/�D�P�޿9��S̱�XB�ɍ�*H��D������p�	v�B�I"YK@��	ٽ}�v���Q#5�B�I!o"d�']3tL����52x@�$�O:�"~�� �@�VoA�H`�@@��6�C�"O�("�>i��i@��;p���`"O���)65��1C�8�P�Q�"O���a�$�@K�õ%�*`c"O i2&��tl.�����R�a��"O�2KV�9�]k�^�dPj��"Or��Վ��Ԅ��v2�U�'�ў"~j'D	�gef�k#n'�[R���yrnͽq�ȁ�/�v����F��y��F�NY� ��� 0bM�ď)d��br���V艐�R�ER��=D�|Q2j�*O<�0¯_�TFB1�6D����牗G�t䱐(��9�����2D��i棗�@�y�W�M�PY���&2D����HG���Ɋ�>C�X���-D���E�^��LE2ǧC�Ir^�7�-D����A�Tr�K���B�2��R�*D� �1�ީXaP�qF��)+��ĩ�(D�D�2MƝ�������?2㎀�&:D�����37��/�5X��E�$�9D�,�4�	:�ab�6P"<�
#�6D�t%'ߐ
���C����0�Py���2D��1VEF�uvD��n�@!
Y�/D��R�$�<��ᦌ�Z���cb�.D�`���:ofdyХ�{m��1�h-D�|PQd�&��hE�7��0c1D���AIM�p{Hhؚ[��l1D� �V��Ib~=��
W�vFŘ�/4��HC��u�%[�Ma�tBpe۟���J4�	@��v񺌚d $`����M̓�qB���[����'V�<��2��TzGE�$|ҝ��#�=b�A�ȓ���p�]NVe�q���\�H�ȓ6�F=��]�j�`�A¾W@����Qg��U��8r�n8F�0��)Ζ�:4c�84>V��`�cJ�(�������I,%����d�KyR�b��/�C�IwsΨ���{�0�8u�'v$lC�U�rA�f �8=s���lH ��ȓ�����D�61*$��/͖]lp��b�zl�B
�#v����+a`Z`��2�E*V��.2İ�a�E�||pY�ȓBF@���+۴gE��2�O_w�|��>J6$��n�bV s�8Đ((D��)U���3��ݸ���8$&D C�%D�@`0d��~%��1��0!74���"D�Ĉ���B��)(�̅.����3D� Y�KI�\���(��W"���B1D���SlT!J��4(B/�a�0D� Y�([�8�A(	۠%<��[TJ+D�8�� ަch�i�F"/9PP��6D�� k�B`�<�E��FD���#�3D�@��KO2缌Z�MF��(�&D���Q��+Hqo^<��HʅZ!!�d�
6.*,��Ȁ�W�X��B+Z/!��C��:��lD>X���)[��!��#��4��c�8�t��F"E�!�dX�"ndz��T����R ��!��˂jG��z�'��`'�U�-ا��yቀv��\�5�Y�4:�PK�ذ+�~C�	,E� 3h�Q.�䲱�X�Y2�B�	 �hD��J'�|��$,�@�B�	���xV��*$l��V U�;�B�	��Be�6/^
(�R��Q,S�@� C�)� ���ğG�*c��� iu�x�P"O�a#��r�m� L�G|�xx�"O�Y�U�R3"��i`��s����"O�]��YS�L����N��@)v"Oޕ��Ȓ[�+NU�I�YQ�"O$��щ
)T.�c��08���#�"Oܠ�l�+Vj��6�ɹF.���"OX<�T'#!%����Ҋ1��\Hc"O`h�4i����mh���%vꬬ��"O<|Ƀ��D2�t�!��f��x1"OP�6"Z<['zԹ��LE�q�"Oj����,쭢��&B��I�"O����(7��]@����\s"OT���%*u���J�"�
R�<��"O.���)W�1���V�	�l���"O�������2Tda�O��B�Z��d"Oȉ�v��.����/ED�}X�'��xjvS��1�#�ǚ'>N���'!�钣��/U�H��v�R*�B8�'$|��J��H�� �%�D����~h<�c	��<�L�z��Y#YL<,���E��y�%]��R�0C�@jR����y2m�HK��kA���ZȪs�]����O���#LO��q�N�)F����ƞ
ƴ�0"O,��Uă��2�9RD�\�X|B�"O���2�_�E�*�a��y�hDP�"O���c(�3Z�<\r� Q�,ʹɫ�"OP)āF� �LR/V�w��Ph$"Ob����ZU,��l������S"O��i�C�*�Ը۴,J�/�t5�"O�̨��E�ޜ��e]*)�F\0"O�%��야(����e�o�4@9�"O��%��L���˧/f(1�"O4A�����6�x@��H�f���"OZ�9��|}�<���ҹ|�H�'���'�ڔHE�їR�"�-����'ML��C��X�B�0�a�#y��9�',����$Ҟ�S��v۪-�'/��9��4_&x�xDe�mA�X��'o�025͆W��-���['m��)Y�'%�8!�I��]{� d�M�
�'�´��IC5͂�����6H���?��
&X�gO0)��}�ŏ=���ȓWh�QHE���}1�	]=xCH��ȓ8v�U�_,k����BL�I�x���V��!�'����Ǎs\�H��j�j�_�7p�8$�]� �fY��x�0��㝌Q@8`�L{�n���M̓$TLu9gJ9;F�x�χ ��q��I<!`��|��`�E�ˆ=92	�)^�<ѧK(�l$�$lB�{�B,��N�X�<	���G��U�ul�>@�Ҁ�`-�R�<�*X%��ͫ�����@�f�<т��$U�����E�f���0�͙^�<�7���^1�
�`�U���\�'^�h�OhqX�Lϒ$��	�!D�8�-�
�'��x5V��#f�P�'j�@	�'ڬ����1Cp�|{u�#��Q���)�4K_�� ��bJ�
I��2d^��y�ؘB"�	�P� �P�u���9�'�$!BY�kaq��
u=�A��'4x�O�2V
[@�O�VS�����$6�'O�Jm���I�I~bT��!�x�vH�ȓD>"�Y�͗	�fl��Ώ�h��S�? ���2L�,��ș ;�Պ4"O���k���\���\�'X��w"O�a9�cĘ���&oU�>�2P"OR��$(�>4�h�vO���J�F"O��ۦ$֦&��Aq�B�z��E)�"O��q�T6/h��;�ެ6J<��"Ó�B�F�`�+k���P"O��8�D_�<nnI�U�L��Ч"O���@W�;���2u�O i�0��$"O���3���bQ�]I��4���:�"O"�#�ݠR� X���]5:�����"O�QB��S�!�������Ee��2�"O\���� �p�na"1# U
�qd"Op�!�̟Zh$�P�A�xE����"Ox=�`G �B@�2!ąC0��5"O�-uG���՘�2X%`ՙ�"Op���^(�P����T��j��"Ode�r��G�θh��[�M͠$�'"O�3P�υ.(���nO�����"O~}��5*\����ʎ{�F�X�"O(���P�0������,t�1�e"OR�#�Ί�?�����/.W�"Onp2H��o�T��8,LЬ��IQ>U����^P 8���>�Da�@6D���`.]�K��y��ȝ�!��z�5D��"�+��u���C��^���i4D��3�W�B��P�JM��b�a�%1D�8��p���1O	�tYT�RÎ,D�B�o�!Z>t� j	�>�2�tn?D�<kW��HL�a�l
)����H �O��	�xۂp�&[��Ndⳁˀr��C�	{�PpZ!�Li.TC��}?xC䉷R�ଲ#��h����5*0�B�I�qҩ֥@f��i�橃}�*C��-3#����F�Sx�����ޢ�:C䉶����ʠM�5C���,C�I+p>�y�nZ)�T!�r@�"F����:?f(w
f,�6� �~�J����IW�<��#�<��"R#4�6�C�NCP�<1'G��2 �R��8S�A3ǫ�J�<A@a�M�u00�C5���î|�<iEAP�O���@��}���I���u�<��IQ�'pd��u�O�iFC�s�<�P	�o�9�$Μ	x����͕o�<q���&7��hXd)�"�LT��IGm�<q͚#����7J��k{���g�l�<Y!� �P�&h�v�)�ν�P'�}�<�a߹�9;�	�~`�u�5o�<	�T�r��4�� ։xc@b�<�R�u���G晩Y�4�3GX�<�u��-L��)�eI�.�R���g�N�<�`��V Dȸ!�³_�6@��b_�<9%������ �	&�Q���R\�<	D�_0� �HU��?:�*��&@EV�<!6/
�ܢ�E��B� c�5��N��h�@h�7.�(DƝ�w7���ȓa��8�o�+t�U��F��B��(�ȓj�R9��مT>��A'�=NrT��[�Ą��0ƭPSi�^� ����l��h@�+�$t��·�1����ȓ�ty�̽'v����d�Ȍ��0��kT/&�<q1��^�Bt��ȓ�V�k6K۷��5��JuJ��ȓoў٠��0���Ǣ=��ф�S�? �-�fȁkl�T���Z�p�`k"Ol��)ޤWt�ਖ"Q�m}�%"O"�S#��"2��� E�'\<}Q�"O��I�,%:�@����U�"Of��g���P�ջ�(P�ƴ��"O��1����D�ԬsB.L�d���p"O���O,|,(�a��*��
�"Or��cB��`]�KE�eԐ��"OX�ic�>d: 
�i߽&e<��"O|,�%�K�LB�xgk-rc�� "O����/��M##��aK�y$"O�\3�"�4ঀs�JN�Bv���"O��@J ��#"I#t�,�A�"O�a�� ؾi܂���ؘ�V�X�"O�%�:�"Ż���9}h�3�"Or����A�Er |R4瘊bz���"O�(G+��0�X���=M��I:"Oz�rr㊿L�0x�^�<���"O����� 1k��
�Cѩ&/���"OްJ@�2{��]Iw�8*8�"O��	jU2�>��#�Ű!�.Y��Y��E{��IĔQx�zpN*S/��a�ŀ6yb�)�'<��p�c�OP��a[�
�	���'��h� F�S�����r�z�J
�'�~����^8٤��@�	z�`	�'!8�[sԩ<��L���;��Q��'�V��IN	618��6(('�:D��'�&���
W.�X��!�^	��'i�4x��0j����A�D���'��S��\f�P���
�$g���'��Q)��>0�F��Pc��'s$Q�'�L��b�� ��%�O�N�����'��12vKF�L#��4��A�s�'��鷅�^_ΑS1�F�4(%��'
�Z������i�c�H�'��2�+�>5G���eJăW�Z@2
�'sb����;3L���%+�!z���''�A%���(h���K���8�'c�yȅm�1��ei�n��Hw�B�'�r��d���*E��;� �'D>(H�'�0t+�	� �ܫ�☜5T�-��':�H�*P�x|�JA�Βd�]R�'D�9�Mv��(b�_�����'e�(A?V�Q�a��	��D�'H�y�WfOQS
�:!�0�: �'p�t F�����D����6_(B�'\۷D8���'��v�D9
�'ը��C��O� qjGd�%7b��	�'����=:"�*�ϫM���	�']4` Q!�A�
����UE�E�	�'��͹!�si����j��2 4p�'�&Q���"~��3��&�0-�
�'X�a����:�����F�d�
�'�H�CηMx���O�1|�z
�'���QO�_9A�a � ����'���ȑ9X0��U|N� ��'9���� �2�����so���'��-;��� ҆�:r.J�,A��'3�	[a���K@�L�80�d��'@`�{bH� �UH�ۭ)D�z�'Ӡ�۰�(O�h	x��$V�|9��'r�x� �լW�.Z�A�Cb|8�'YJ9c&g	K�D,�s��?�ִb�'�
���DS�v���I��_6x�=��� l��m�rnt`�!��a��#@"O\�C�X�}�~9"T�ȿ"XPU:�"O���,J��$B ���\�c�*O�!c�E�Qd4���J�b�d���'����єS���(͓Ѐ4D� ��
J.?\�	�� (<����7D��B���?���!�!�(	�t�4D�<��M�!1Y��iԠQ�;���"�6D�p0-�==C,� �Q�о9���.D����-
[)�6e�*;���pL+D�0["��4B�l���d��\0uC&D�H�4mܞ6���kC�L�(ҖXYB�6D����B% HХy�nֽ%�Jِ��5D��1"�Qf�SW��%�F�Z�(D���Ǣ^^�20��M�kl�]��('D����搨6��"gL֦V�89Ug#D�I��Ѽd�ڸaRO��1��Srn;D����$~����7��!$ԁ�C8D��ɧ�C�O(�@aO�a3�@u�2D�P��cP�,6����9�����<D��c�L�)):�g
:d(�*�C5D�ĸ���,����cH&j�0A���=D�0���@3�vq�e�²Y�aC�&)D�l0B%�VZ�{�e����%(D��ʆ_4#Ρ�'#7z"��'3D�,	4�ʪL��9C�F�\��w�+D���Cگ"���:�L�&/'`�T <D���w ��M<tZ2bW3o����&.D��aB��9ZA2�'�q-굸$�-D�(��(Ǐ����F덗C��9p��!D��(�!ǠK �2m�(��I[� D��ar�D+L�\j��=V�A�G>D�8�dJ0I2<zp�w�p�%k<D�4��د9���%^/�b]{�9D�D�
4����N�(U:��*D� ��Z�=&�h��V8Z��$��*D�b�(90	�W"Z1i����c(D�x�cc�zlH��e�p�*1D��H�-��mG�]�*,Y@D;`A!D�L� b �!�,�⅀Ffʈ�,D�8f�F�[�r��`C�$|���� *D��j���0gf
i�Q
7>Ђ�a 	<D�X�S�_4�nq0L�%�Xt�=D�D���4�J�X&��q�:D� �6�X�w���@���?,RD[Ƥ#D�@PM2-S&��ѫ=q�s��#D�`��)F�F�U�S�&6 3�!/D�X���?)�&C�H��Ib6�'D�H�Å�j!p�x#�UJ�-iu�&D��y�X,[���S.A02����%H1D�К5�ւ���(�J,^9�� Tj*D��;�GWyU4�{"gó1��!�&D���BT�S�n���+{D�X�Cj$D�T�0DȞIy�!�&I�`S� l,D�xp�O��X��a��+N-�nx�C+D����l� j�>�hȆ�lx�R�4D�LhU�H�P�d	EM
�\>9��G1D��ʔ�ʰ 8"e����$(�����"D�<1#�&��	�b��0n�����m+D����� �j��D��(��$D�,�gT8T�G�]�	����e�!D�p��2��9��B��e\f��� D��@1�ۙ	!�h7��Q`�ҕE*D����פER
��#V3k�:-z��(D�� f$�B
�rN��!��& ��D;�"O<���I�tS ����Һp�(�Ru*O��Q�M~M�Sp�G?(���' ԙkЫ�_������)=���;�'fft�5�ϑ@�&��N�l|�		�'6X�D^�G�Vq�Ė+e(@�
�'z�}p��i��xA�-U1q��d1�'�� �\�Z�����U����'|�����%F�8��U�yUn�3�'\����1T��xХ��[�|=�'�H��w(��o��<!�ŮOl�]�	�'�Ȳ���^� `���G"T��'8��(�#�.���uz��`�'� <��aٹov�)�@�Bޡ��'��H26��
/r0t
�e���4��'�.��-Ҹ3w�����T��*���7�����H��|�6��w�S�3ӎ��WĘ8���\���k�C����!�E2�m9#l8�t�3|���ȓ��}�$�O/I���!!5H���ȓV�l��T C+&��V+�'"Bl|�ȓIlၕ�Č5��y(�#1(e��R�x@36ņ'Op����Ƙc�rY��;�<1D�X0�Ψ�5��`h���xg��2��`��#��F���ȓ/�R :�#e&i8�߀��P��J|ҔrA�[&OD�h�@!&���>��� ��wW��5�V�K>��ȓE0�q�ż" �q��B��'�Y��j����b�@b�r􆉄�i���P�1R��Bc�O�0)��'P��B�݀dD�$�b���u�j2�'�.�17�I/g6�Z��J}�:���'ޜ~5ZEB�W�\gJ��'��y����Y��D�;"�ɨ�
�y�.�8�.��5�_���z� �y"�Q�r(j�۵�2e�f�`�����y�[�恻�H�,\�xY:uL��y2��X���@4m�6[��(�*��yB�U7X���!!�0`�rl�%g���y� Wn��b��B�[�>�a�+��y���X�/T>J�A�Ԅ�'�y�͉Q�X���=5�Ke�Z��y2hM�¸�a@�CED��)��y�C��B���IVBƄ:�B��̒
�y���. �\�YIt�a�H�K�fC�I�4��$�:F~��b��@�m�FC䉓^Z�1��B�E��t�U��(J��C�I"(ڼBD�[�Q����%�V3
C䉪9Ț�H���$e7��s�X�C��T��u���Y�����iƛH�B䉢&���`v'�] 2,�d��x��B�ɽ^��Ʌ,�Q����1m��(G!�� ��T���9���3K��v4!��U.X��ȣ�� Lаs��A�!�ɫC	z�r"�q&&�#G�E�!�ćTԈLk�M�|��2�f֔D�!򤛕$���r�L� ����EC!7!�d�Z��A�Dj�O]�X�f��i!�ĕ�y�0iж`!>%��h�E�V�!�>ȄP9t�[�LXd� JM3,�!�Ą {�dYx��O-��T��I�{
!���sbp��_�-ޚ@��g�n�!��F��-�a&O�*�H��6IQ1W�!�� *��� ��hŹr�"y�D	*"OV�f�&1c�����þ#l��bc"O\	1��8b��A�I��]k���"O|�rG��u�@���Ŷ	W|����,LO|�ѕ.V�,c�`����):��� ��'��m'�d�1L�+>`���F�Ιat+j'�yZ>��q��J���5#b�1���>�B@��]ǲ����t��?\J6����G�@���`$"O��Q6K4\�rl�#'�2��i�6a!�y�	/�g}�L3VbQ3AQ
N|��@�	��y2ɒ�d��Ѡ$�!ܰ �����	pX�L��7���Ui�h	�"&)�O�q���%.F&��=��
V�h�|�Dzr�'���y�G�#J�]����xײ���'L�;2�]�r���7〼k�"ɺ���6<OVm ����H!���t�|��v�d5�S�	�]w�h4�4><�Y%�X�{�!�֠3�2\QC��;�h#d�ڙ�!��,.
��c�+)u�荒��	�qs!��B�wLRX �
��e�j���ς�i���b��H���Ӡ��vri���- �P�v"OT��&j�<I���R��7�¹3p"O�%�*n���9��F;t�	0�"O�� q�G�����pgE����)U�iJ��D�9/]@աu��?)u�pO�,l!�J�0�(�ʎ�D������
�pP!� ]�tT@bK�-�Tѐ� �O�!�$�s}`��2.�&�r���2�!���!x��Z��B��$m�)�'�Q�x��	"��17�GheYRr�R	F>r#<i
�S�hˢ��Jd���B�*؆�c��l2�^1� uq�j؜rA=��6����C��d7R��/�?|�r�ȓ0H`�����T8�˺.GD���Z\���L�<]*tK�1!���ȓv�ab܎:
|�)cB�`����aȃ��-���b�?RŪ(��%?��Ji
@"�H��^iU�Ia<	$ h�es�M�#b1BUJT��a�<�$UH�Vy!�,�^�H��m�V�<�0�	�k� �����|3�q�d�L�<٦�I%Sn0	��G���%�TI�'�#:��fT��� ��1���:aɗG�<��c =َ���]� �����!�*=�S��M�T��N\�p���xPtQ� ��h�<Y��8qM^	!'+��T\��
�b�<)%���'�9X#	Ւi�� z��d�<�*�8RZ�����&���u��E�<!�ǕS�F���N@f��% �L�<A0��!)�䃶	\�*��x��B�'��yb�;i� -"��>Q���)�OR7�yB�EΜ�	�$��O^�-#RI\�ē�p>�!C�M�`�@�CP�wRH�H�g�z��hO�2S{ba�}���"��+��5A��U��?Y�'�2e(��O0����V**~� c��ޢ=)!�K53�����f�� ��,��<9�{b�'eB� CG�$4-�Wi�$z��'p�IRS�xF{J?%����4��`!^�
2LD��j4�Ih��ħ|�(�b��N�l7 �{��+��G{��'�r�q5,#	�֬1�%�^yћ'�qOf聉�i�?�т��Q��P�2�:R2	���0D�xB0振&v��dQ���s��c� ������x��s�� o(��fH3b��ʐ"One𠣊�xZ&�y�̑H�T��"O� ��9�ꕇ]8��3ƠN�?�~��"O��R#,�V�T����=bg�q��"O$��o��	���$X3(�\Q���V�'��ӵnUPe� ��5B��ӳ��{���U؟P�4��C�@�*t�T|�	�a D���<]��<�2�ε/	���S�<D��+Ӌ�����|'�H���A3n}�C�IhDV�'r�(� ��:h��hO�O	�� +r���q�ܭ
)p�Xu�G�Y�!�Ķ|6U��t�ĩ�#��|�x��˒ � $��y�����ybc��BY��	�Լ�3+.�y�K;uj�w��	0�H���n��yR�j�p�I�5hA�cB�y��H�Z�<����zOM�xA$��|�������ca�U����0M��m��X�"O�,���	��dcCb�gtPbA�	y�O��*�"�j\����74n~�
�'l�|�)�V9.�� ��y�p��'�ў"~�0�WXی�:�Ã&ɰȋ,IY�<!�CQ�Zؤ���ϔy�4ȳp�\�<�/)�"���V�x1ʥ;�c�V�<�ň,v��V�ż ~8��$�O�<w���!�zyf
���|��J�I�<1�ٛ>Щ�$�F*{�����+�E�<�4
7�t�k� �,u��P���j�<9pj	a�t�t���AM,�h1�[~�<��f�<QX��V�9s�Ҍ�U�<Af� �^��g���\!XDp`.DP�<�X/$�ZTa�K�(&���B��U�<A���.��$��9Ԓ�kTG�P�<�0FV�:���ڑ-C:�}DmPA�<���F>X�ɐ�C���e͑w�<є���,*�����>R"���r�<�SGM�{��9��ۼ	�BCfpy�'j� ��#V�"��fF�0G�b�{��>Q���'Dn��1��+U"�)�kE�'u�#�*��0�%�P?O��Dw�|bV�"~�rW\Az��ό���b���<}��
�L��`ʬ	2�]�[�D��'N�}�@��4r �g�JU�A+0϶��x��ڹa�(��A,g����NZ�kC���)��=�� Z� ���4�N4/���#�),O�T$�x��w����5�St��|����.����'��~�mZ8L��y1W�*k����d�(O>�q���J��4��0o�X��U+=D�l#� @bU4���C�5@u[֨:����������o��2��
aX����Iiy���MI�<s�!C�\�H�JaGm�듵��C��S��>����m� X����A� ������3��s�LC��"lD�!��I�X�� Z�,ړ�0<)�톯ag,���"Ok��)CS)MG�<y�Q2h
\��a�.[`-h���C؟\��Fh����
�+4�<�c��;\\��G{җ|���/rj�C�@�/5������!���>d��k�������ָ}�2�O��I}~��	ܖq�u�c,Z1<�1�!���#=�	ÓZ4�q���y��*�U���ӏ�D5O6�ڵE�~/D�A�OJTA�&�iʡ�ǚr/]0��=.�2qsTD�+k!��6���W��^�hpW��9iZ!�L<�nq{�a�)=���9��+�'Oўb?U��Z�ժD��S��c�Ǡ�l�O^ҧ�g��!zN��@*Y����ֈ�WS!��'7z� �hr�@U�K����(O�	PP0�4Ou�Չ�0O����I�	:Qr��=G'&�;$K̅Zp���	�M��%'�4e��q���l}��R%�׊"!���1$(t��㓈P��ߖd�O��3R��qyH4(���\�<���� ��`)s�^4!���U�\@�l��F~F��F��|�!���U ��/S?��:�e.Y.!��8t�@:�iνB�5�R�!��8�0�Y�Q2��Y�.ׅJ[!�X-jy���pDD9-ub�i�@ڐ#E!�d��Q`$�Ad�_xQ��90�!�DΗjԀ	�N1O�Lq� �J!��И)�a�4A���W�T�i!��a���+� s�,��y�!��ެg*���#S�P����E�!򤄦kG\�1��(gڶel\#KoJB�I�a�R���e�EP��#�d�7<B�84�$�� KHI�"A�#
� C�I+Wfl�ȴ�ߓ0�8���'N��C�����@�KɁK��"0���C�l�`	 &������(���ȓ��LI��F� M��q���+%b�U��ݦ��I�xH
��d��f�Մ���V��+��Y���C�c@TzD"O��!�J�f��;CN�.=�Y"O�tB��R/IF���D�+�mA��yj^/ K�鐣F[�5�b�  @��y"��0
�l1⋚�5	h@Q�C�0�y���I�y�X���*�O��y�o�!�pݙ*�>Q��Ia(�1�y ]6{���f��K��i��ֵ�yR .}Vq�Wf
$Y>r��G���yr��22�ehEkHz�<����A=�y���P[R!k��.lR��Rb��
�y҅�u^`A�.�(>ɱ	ɓ�y��Œ[FJ��B�;��Q�G��yB�U�l�pTK����:�����W3�y�&?�<��d�#��yHяF��y�G�4^�~h��I@ μQCBF	�y�?���EF��7`�!�J� ~@ŉ�A٬�0?���OF�ਘ�Qb��yI�(�x�<���|����
��,q�H�M�<u"�<^Q��f�)�d�h�q�<Y�����ű#i��&`�Y�adBQ�<��� Qg�1�`�Ιns�t ��K�<���F�F��DJ��r\����c�<	�Y'
�E��0�:�6�\�<��O�N��d`����3�Z�H"�^�<�F�F�P�;A�K9:2�9�US�<�6�Śl�^�����/D x���@�<GF�<��)���1[i\�3��VT�<��\)`s�ܲF�U;=�9�5�Q�<�阥<P�ӆ*���F"AI�<�$��![�L�
�[-�
y7Ň~�<���юXh�HC��P�:�[�<yFŖ��4%D ѻ.͚|BeN�{�<�ea�K<������g�&����Fs�<) ,S����Ó7/�Lq�ae
m�<Y�R�[����d�1��5�w�@U�<17k�'_,������Hi��C��[�<�����tڴ��bᰑ@T.V�<����25�F���%���ޤ�!#Q�<A�N���q�Y�Zv`�:��H�<���2���i���	+"8�7�O�<� V�S��t�űr��6v�mr�"O䵢���g��i��[WL�P��"O�I�UO��_xDh��ѻx8kb"O|Pb%,V=;� ��>�������xSڄ��'T':��T#=�0�I�$�:(k�=��)���:�.F-jHR@٠g��}����-ߩ��|��E��Oh��3�g����O�Y��H"O���JG�H=�$R1@[�6������ěc�b��t�#��>�v-�+Y|�=Z��XoD<sV��@x�0b���jRKfP��*! [�|1�XH��9u5X�%�?D���FC� Ĭ�R���$�v��3�:�d�1!�`���⛚�ȟL]Ya(�.䖌[�"�#d=h���"O�0 ��0���X���;v�*���́ED>�O�I �,�3}r��s�(��U ��*4I+��xBb�S��a� üi�$�v��2 ��hJ��H>���I+�����I.5�����(�N���	�6������N���DQ]�y���5,O�<�m�(z!�dƺ�%KsN��@@EB��M�1O�L`uE�O�b�*2/�74O��Z��ժ۴��c��n�<1�ʆE2(x���):���u��i�<Y�a��fB����R'W��#�M�<�נ��ƀ�t�W2%_�y3�*8D�8��i�>�:��ӝfS�ő1$3D��y��F�~���)@�xO@�!��=D��J��ݬ[`�����;_��ѣf@;D��!�	�(L�`��A�����9D��rD��^��uFP��؁C��7,O TB�,�ɯ,hڐ�狆3;�
=��nG�.C�I�k�`2�HT�𪶉�#��'����%͓I�S�'�\�3a�ǔM����Ɉ�I ���h��e`��)ǘL��/h�������Ó/��Ubs����LD�K�\ߘ��F�<��Bn�=��t�o) �a��	Z�)�~C�	�O�d��$�Ejx����K{���D�MW���yr�� ��h0`�B@3�뇧ߣ�y^ f����NܘAc��W-U���	83���;���i��5�sCO�=Kg8�j�MW*~�!�d ���*@>k,˰
Y�WױO6�b��5O�����	*~r,�K�K׀6�<Y�"OQy4Lm���#I�h(�xQ"O���вS\$�#���y"���P"O<A��셉kc�<8���� �"O�E�V�k����6,Q�%�J,�"O�t��(9)dP\r�lZ5OI�4�"O��0�b�"*�K�%�DmpŰ��>����	����?��f`Ʀ1�"5q��S��J.D���w�\_�\��GD�xq`�+e�k�I�yuj�%�.�3�	�I����ʌ0*����$ާX������*2���3,O�$�ˇ7��r�'C���8ņ^�{�~`@�)���?QM=hL��#�
R_�`-S1K�W~R�%4�J�J�R�أ��=W�0��%����JT�]y"��%٦ �T�8�y��F�G�����J\-Ld
��"J��i�hi�	X�*�������+�1�N?���� SPJ5�'�B�k�`BSQ���kF�x[N�
�-%�T9u�ܙ}|�C�Ցl�|`E�R �D壧@A&=�R	�6 N�Tc<%y�
��x���Yv�ڃ���B�d �@��dI��1�t�q,���"%��C��|a�43̚i��h8k�Ԭ[Vm�V~
D������V�'����-o϶I;0�M�3�6Y�aL\�S��V,��Ɯs/������O���V?��> ��C��Qe��X���A|8C��h���vHѕJVv�DhT\ƤA��k�I��֌M�T����쟲���I\n����U���E"f
TA��L<	6d��^>>[�{���'T��ͳsED!c����͋��ia��
f�������{ۨ�p�mQ�4ۨ�@1���-i��?1B
�Z\��``B��Fк���^^��3Z�髣��-����� �Z��E�1g��)%�ʕb��iZu$YH=�B�+�T9�9�(0".�^�QA����O��X�w@ك �
�@E�Q0m��+��z�	 bn1��� �Кq��+0 �[�A��_�b���*O��1��"�x@��]�sN�ڤȋ�നA�
�O���Ğ*��a���O��vMK��M�u��s����'0q`�GI��� �V�� �}��Ka��Y�`�U�tu��!���}�L�)�"�bCD�z�hB�H|=@��?A��)2TX]�����?٤���5�x�{���B�?)W�詃��D+�!�ȓ&&��&�0@B���� o lx`��*iz L>E��'��H�	R��Z�&�>Q��'�f,30�@�d�kg�7��4��'��[� �	�c��sCJM�l���C�#�O2(�)]�'N"��J�j[���V��0s
�',�Mh�ԀQd��א%��t��d[��F � !�O��icSH�.}-��C�����'���2��ݠZ�V��đ@HFi��������,eJ�D��"~2��=!$|`y�JC�&����0�yR�9v��С`����@b�}VĜ�Ie��9�;!��ȯ���8�)Q�y�jH�+J��S�L?�O��#�&?D�,9z�(ǷR�lxIF#���(4�G�D�xl��&�O̅���٧K
6�C�v�<�jC�ɬ7�đ���إO"f��w��S)0���%�B�c�V8
B䉊'��m{�ԇ/2����d�ҩh�	��$ZY��CX/D9aVj=��dQ���.]jja(a�
Z6Ruy��4D�,��%�'r�:�#��Mk(�"�CU3ZXFy2�ÿj8P���S�6Z��g�'e,�����,Cx ,Y!���=����D��I&FW7�HLʧ������� K��h��)ZyP\|`a��=��>9�6(t�h�K��+��蹅��H�'�6�3&ǋi\��
$P��b[>ѐC��1ɠ��B�Βb�A�wG"D��qb�;7gB=h���/���^�&�P�3�FՀQ�����hT�E��w
�HRg��i������<e$u
�'G�Tc�6�ތ�0��7�R��_�@5�yK!�L
?�CND���D�	8w8+��2U���2��-ٺ��dW	e�d��vm�����\i2���dK�8j��bA R
'�2� tcʽ��>i�P"4�bȓV��A�X`rT��N�'�n���	"@bh�ȇ��)>����X>5P�*I�v�l|�7G�c:
�҇�$D�@�U�2
����7/U�?�LP�4[F5��ύy�FA�SDh�4�~���.m��D5fd�"��D}��C�	�R�x1�1̈�	X<�q����P3����x�pa�1�:УQ��?�=�N�b�� �π����ErX�!pBˊg�ε{��21TI�Ǧ[��əg�YI�=3�!�t���qJ
 y�����-��B~�9�,+�f[��u��=R���ᦠӡ���;U��0�F��M!�q�wBL�9f�B�I�N%�yA	C#���"H�a���^��6T�q�ظY"����B)�0q�0a���7"��q�%D�8kr`K�;2��BnU(m�c#}��\*Q3(�$O�F8��8�����q�*Y�]��ɸP�'�H�0�(T^e��T_?$�*��ũ/�@a��JZ�)�"��/]#2�(po٠p���ȓ(4-3���-�ܤ ��P�y	zE��V�(���0z�	՟{M`�ȓ�������k؀�)Ej��R�D�ȓxi����KE!\>)�굆�eŤ�PR(Vc����y�4�ȓ��hʖ_ҡ�ԇ̟?�Յ��	"$쓌-h���(�A�����z�Ĵ���Ǫ�L�cvL'p|�ȓ6+6�i&�=�*��e쎕���ȓ\򴃒��&A����4���
� ��J��3���|�L5��I}���ȓ��ثTeZ���KD��mޡ�ȓ|����۶a�w�Vu�O��eǅ���䌩�Jt���BS�<��#�'�a~���kbF���!p��q��69�2�a�3_���=�T�GL>�( �'��E{�'O%<�뷀�g1� t	����^�ٺq�P5zo�X��"O� ڸ�%nBcΔ��E�K*��2��'�>9`���;NT�0��R�"~�BZ�9�^�$��!L�z4� ���y�-N61����.F��s`'W2��d�;?>  cO _������%Ag�K9�UF�a������ f��D
�ܸ������&�Q�H֌Dm-b�ik<�0�Ϝ���q�Õ����
�Z�'h2Ы�'�$>�t��P��zx��hR<QKR� ��G4z!��O��:4Dԑ=U�Hq�N3+X��GIP5��%e�)�F�� �GB�\����¥?U3
�'1 ږ ]�n�<kǥ��2є�k*Op���L�P�\{�)O�m�qt ���ҍXG��9��'X��ϓ�>��Dg��̀VK %;�! V�^(<�Ҋŵz������3W��aJ��SI�'�\T��I�/P��^qy',�pV,�jcAG�S�\L�E"O�<�@M41:��3��E*,C��h@"O<�ύx/8�� ,D��h0"O��Z���.�#@� �l5�p"O���hB�>3�F�!pm�Q"O����<=v���e�7u��C4"OP�@CO�i,H��b�cf�V"Of4P2m�5Xd(��1"�
���"O��@��9$�Ȑ%a��
�]ȗ"O�ѣ�bX�N |�����X��&"Oq)'�%�
�;���4S|X��3"O�`�		.k(0`���*{8�"O������K^T�
V�\]l`�C"O�xtǏTBK�j�)��'-�y��0�Jf
�f�vQA�O���y�ƅN���S�ݝC���:�B��y��G)���_FD0��Ǐ�yra�fA�a�%aON�\aq H��y��̞/��D��&�@2��AO��y�ο-�tٗ�߄Mv�(��^��y�⏞%:B]���)C~8˔$���yR,��b
��X`��(S`�*�3�y2�x�ҕ�fVB�Pe��&���y�A�uYސ�P���*�`�cƷ�y2l��V�ըM2�5(c��y�h�p{���a&	+�.�
�yrH�:'��)JR�� �!"�@��yr��3K��!ӓ��4O� ���Ű�y�N[�-R����
�	*%�-�/(�yR�՗3�)I��Q�Pvʈ� �#�y�i�>ȶ��Őgi��r���y� JZR��$� Y2�Tzu��y�B�2O�y�WdL�!���eH��yb�T�=�Y"7(��\��Z��y�D�����-3�ݰ�DS.�yF�"h�(�(�����ӵ蕐�y�KS&D���( ���,s�Ï?�yR(@�Z��w�E���������Py��j����8o�������g�<�K�*�.�bfD��_�Ja���U�<��O����1a^y�6%j�CW�<ADˋ".���������Q_Q�<y�䍜�Dh�r@���u�<�Dl�4^'���	�.�)_T�<V��`�>�¨� jӌ`�f��Q�<y�!��Ā��R�p�H���`�A�<u�,"�z+��@�"�H�a^K�<tO�0�� �6."
k<Ex@��I�<QW����*��"r��d�ŞK�<��
�3Z>����4���f�[_�<Y�Өf�H`���V�j�$���l�<� �q�����]5�a�D%̀cP� "OʘQ��9%)�e7w�0�r"O�����;�DK��+IPb�) "OԈrC��4����4�ͨC� ��"O��8�'Z*K&����ױ\��8u"O��� E�L!�؁0n���3�"O����K4`�Έ87L�����x�"OFL��`���AC�K/����C��O�p���1
çIm�`jA�3ڠ�#[7t���ȓr(�J�G'`�š����T�g`ҩ���Z�D��Od\����&��|�'V-A�8���O>�ô*\4:�����_�|�a���O��m�qA�˰>�F�48W����摱EӨ���Awx���E�P2@ܾ�:�[�DSF)�2OhΙ��ǅ�sT5���9D���ā�1�\8�k�Q�2��� ���8T�$��vk�=�ȟ���5b��W�L�k6��7v�8jr"O�HJC�A,M��Da�>D�53��N&3?d�O��3�$(�3}�M��\DХ*b��y%��0a��"��x�k��t2\� $8���R�I��@��C,&D��	�p�I�	��
X��˞�"o,��D���L��+ވ���.}���HE	V�);����)!�� �Ur�處,�$p���#ߔ<1O���$c�>
��G&No �m8�J4N�.� �_w�<�W�X/!������M�� cF�K�<�2;V��a��:C�����A�<�r+э�V��@F69�*u��~�<Qj	������iO�̖�,�C�I�0 ��<|Ռ�$t?�B�I�(1P�&�1'_r�Ao��n��B�	$]j�;F������X��� P"O��٠� y����+5A���t"O�C��O9a6�$-]^�=��"O&Y�����?\���ҭ��,^�1JG"O�P���V��d�u!��Pm���C"O��!sO�D*��k�Q�H�"O�Xw�K��v�adE�m[t�S"O>�a@8�~Q�����^��"O��b�45>PS�dT�y��3�"O��$��X� ��g��=
��T��"O~�&o�g��[��E�3��9"O~	�B�n�����DF�sԅp�"O�EK勝�i��9�g˵2>�!q"O�̛�iʈF������ J"O) ��F�i&q��L[%j�j��D"O��С�
�&͜0���l����"OV����"li
\Z+X�T����"Ojq��d�J�:��
:F�<�"O�ิ�H3P�h���o�(|2n�A"O4p���V�e�Y�G�ǀ0����>��ώ� c���?թG��n0вL>?�f�B�+-D�<'��,^hX`���vKR�i�ΊC�wOX�AՎ*�3托e82�z��!,l��Dd�5<M���ĕ�;����-O��q��C#o7��$��j�&�`��J�C̐(�cѮΰ?y�>*��o�D�j-���Y������	��z�k�>�G��~6}p��6�)��'�؅i2����#����O!�$U�1􂽣uYqf��*FH-V	co�;ZŚP�F\�d�����~" ���\�5��OUs&�U�F ���d>}�r��T�'8�I�gh�1 ��%�ֆI��xYю��AR%� ]�dy�Jϗ�Ơx�eѐK4#?Q`R�%��$�9�"��'Pf�'|mB0ϒ&�-���	:�,���i�i*Pf\�&�Du�@�X�A���Fi�-QR4�OΰH#��f¦\�\�����*"Kf\�9��1dY:|�"���M�6	��FEp����<��sޅC��+W�����]�� ��1D��!�(�8N� QF��47P��	N$�x��T�d���#�/���	V�L�.i�a�2=H!��O�|� P�mb���aNB�/���r�'�,��RhI�.ˎLI@� �T�g��N ��AmP5M�I7��|"h��AÊ�]�Ĉ�r��?9`c͸���2�l�XDdQ�ˑZ�K8l2�@G�w����Y�Y����t��"4n�	G���w�HI�IR�j
@��t卶S�� q�'�49x�H'e�^[�I��1��e�$��a�Y��D�f��(ބI��9�S�{ŏ�]ݬ�q���a�soF`�<�#V�Z�Z��3��Q��pƈ�>l�5�D�=�J (�O�f�|���X�N�Dx���Tmj1��y*1�C�����=��g�8N���b��b!) �4Z��;�ܸiQ>w�����Z�X�������e���K%I:
,������p�O�|9u.��:�N=�j�OPPa˗�����l��Q	�F��x����瘀X�!��X�]|��5�A�Wф�3�F?��=����!_��O?�I��Hi�`��|;��2E͈�w�ZC�ICe�\󃬞� xƵs� ������e�8�#�'w��o��Q=Ĺ�v���)d����'B������ 6�$���B2� <��'*�mabC�3P�A���B5�j	��'?�[�����(L� `�-u4%��'���*�[,m����RW�j�'�y�NDB H��wß=@�N͉�'�D*�hn�YWM�*l�l�
�'�@�ӂZ�'��Ԋ�Y�vD�`�
�'I����@ԝK$�mǀԠ5���J	�'ƌ��u�G���ѓ�[,���;�'�~�q����](�IQ!��1k�9�'�H���@%?�vp��@	�|k�E �'�pٲD��5�q A�u����'z��APO�!ׂpp&Ř�h���'%(²@V��!
P�o�3
�'� T�WH �-
�87F�K�n��p��JMށ$�:Ȱ��!M�8A��5�`Q�+$�#CC�����ȓD�<��/G.��(*7��Z�ȓY�=P5��|Ǆh�a��e X�ȓ?%е+�喃5���{ Ɖ��n�ȓf���&�
48^��H �x��/yA�P�t���Z��aʙ�ȓg]�J���pe�!Kg$��isf<�ȓE���bnFQ����%O�Lr��ȓ���5
����="�	:`�d�ȓ'Q��RABb>f幒���X� \��1�� oJ?!DʔQCoOg�f!��'���h�(<�4���+i2�K�'�Z[��1 �>��'��4	=�%��'u{$T�Z���8�N"<�����'2�j�b�&E��%I�
o�mj�'eƭ)�
Zx(e�����(�|��'�NX�JŹeװY�v��J�+;D���E��~�b�:���: |�y�7D�S&JT8�^�J$�N��d�d�&D�胇%ޛ�h#�<��8$J$D�����\�9�|xF앁��e���$D�H)5���}�$�����J�2>D�\����6k�]�2��.NJ�Ir��=D��z"+��k�
�8s��6|�"v6D�$&��
5���%�7ִM�Sh7D��z��-��P��
F�)�
/D�\��%CL��9!�q�f� �B/D�H!��ڛq��-
�ݧ\��t*O��K2'��GV���u��L�k"O%3qG�&+���(2�K�	�݉g"Ov��럴kj��&�Y����R"O����L�Fz�4H�`��^�L���"O��"U(��|y&T8�oyll��"O�)��B8/7p���7�����>钣Ol4	�	�S�? ����M�I�[3��*��]K �'Ӫ5�g�߆m�X˗B>[�$�Xv,ɔ�5Q��u(<)�
��H����ը2��8�Ću�'����Ƨn�)k%�I�u�����JP����EI '!��Y<�Й����,���f�I�⣋�p>x9!ȓ�-i�)�'�����$�"�0J��J���m[�')&���E5`����GM%qV&�S+O���G�67��q��-O���a"�5&�����8x��4��'��(@0E|��∦X�Y8��Ǻ4+P�Jӽ Ԛt��O⍸����o�y3�Ă�ED,����	6z$z$n��jن4�|rp��B�r̙�j�������.�q�<��F,{����(��0�@	j4
��Ȓ���H��aIӎ`y��	V�_���c&��>[Cl40B�N�<[^C䉥-���a���tn�)�ȏ�-^&˓^6���GԢ< �p��_0�1p��w(1!�j�oؔ���7mN���-AL@Pd����8jظ�1d���
OR���˃�H�p�!eDU"M��8��	:-�8ИTK]�'�\����)6����$荅ȓK��|��x�h�iů[�\��e���`�.��V �ͣ��Ӏ����g�" �Q�D
n�X����A�5��3�ȼ�GjïQ�Љs���%}mp���YxTd�we[�<J�),)
�X��3D��Br�¹�P(@$���*��ر�I<D�x��C	CP�4I��5k�*�c!D�|
B��.dlzEqA��� p��8D��Ұ��^H5öo�5 (��v�8D��ygG��q�ԧ�?�.H�0�7D�8�n�-8k�0��г6�
\[b4D���` H�8�FX��7�>-X@�5D�xӮ�
��j��K8���9D����	�!Ƞl'%��~y��b�	5D�d����:���ӢU�o���.6D� zw��c��h�%Q7B��A�V�4D��k`ݟjm�x( C�~��!� (D� ���Իc�QkW+�.�jukg�(D��q�Ϛ)J�P�1�R�~�,��'D��áD�"WL�7/Q�@����O>D���j�x����͑'����=D�j��0J��p���+�
�q�6D��Y`��6
IEp�e�=��P�0T�,��H��6)v�ZE���6��"O*U;q	�LZ�������a搑��"Od�P!	���ȱ�ޕ'��lj�"O�pK���2�cJ�&O&J�"O�!���8����5�U�"O��"k�Jd�Q
۳!��	�"O�|QQ$��V .4���:"�0��S�
�J�u��'?���ŌQ7&�f�
TM�%�����'j����O���`h�4�H�M���S�'�	yև�O�:\
�f �-|�=c�'׊��g�A�(+Fea�o�&$�}�
�'A�u�¥]�|<7#οI��
�'u�4C i[�h�l�`��3�UK�'W�I ��Im�Q���8�0m�
�'ԙ!��0g�� ze-�(?B��)�'�X�[��m�����<�P��'J�C#�wS^mp��4$@��'8X�:!��⽑�D�*�$U�'.���C��W���eY�(�2${���5OJ��RE�$�v�r�&H�p�P�$D�(O1��ap�f��I�
�ڷ��=�Y�V�x#�K?�S�O"zx��/�$����I%{Ǌ��'�b)Dy��4��7m�4����$���)J�}lӎ8(E�P�OL�X�ΓP>� ��CB͒�QǪU�2&Aٲ����ν$�.�I1آ��5�0|
�n1�Єa�,{�RqZ����~r(���d�ˆ��
,�)ҧNV6�Ʌ�[Vv%�C�ڡjP�do��4�rtc�j�.dwjX秨�(h��%3Vb4��K�ut��KV�¦@XX:sc��:��1@a��:MFF�H��R?l(`	da:�I�,�.��	��6�l�v��M�fm���5@�!��`XB	IP�ث��C!H߫.�!�_�9̌�#�4|Hш'Cp�!򄌏 H4�Q	S�k2P��D���P!�D�.(���0l�E���*���d;!򤗔U��P��[ d@��GE�"(!�d��v6d9bB#@R	2����'!򤔬Q����l(��a��'!�$����h �J�5
���ݖ�!�D :��X"�08��0J�%��}�!�$�lT����\;7��A�ꋰ%l!��:Z�� U��8.����Iߺ&p!�$�+ecpٹ��V:EC0XDC� ]z!�D\�zrb���Mo������5\!�d�&7��I#�!S��!���5=!��QUft����u|`�x�oS�$%!�DS�|W2!*E��Z]�U����8P!�d��u0����k�X��ر̆Q!��ӝS�����L'���jG�M!�R@����vF Kש[r�!��Q��ب Z��F�"y��	j�'rܨz�
Y�y�h����n�f���' �H�s"��q�@82b&�.+�9��'� a�sBt�Rcd���Ys�t��'���d�Y	N�Ã�ёE��iȠ"OƠRQAT�y�h�N1��"OV��ڛZG ��t��.�����"O�0	��K@X��$A>7��p�"O~@{�O�),�k����R�"O�W��dh���:�Cƭ�@�<!��Fɹ0O���A�%/B~�<�V�H>��jek]������v�<Qd�[;y��%�b՝s>00ˀ�t�<��D��p�6�#��&��w^J�<�Q<������$ HA%,@E�<ᆧ��8th���ϵ�J �f�<i�k�$lz�	)Q-ϵfʶ}I�Ε}�<���0]M���&�uI5�1�\y�<�ă�>C�T�b1\�d�0t��y�<)��]�S�vL k�!@��|3@�r�<����;3=�����p�t@W)�o�<��eޓV�"�A5���g^8����U�<!��|+�x���o�nP�.IH�<)��̎3��a*�����*]z�mUH�<aï�:ym���3,N���)���D�<�C�����3�eĭ"qX�Y%��X�<�V�/��h�搿	隀i�FW�<�p%�z�p��AP�)�UI0O�Q�<a�'O�[� �{ǧ�$/�D��RC�<!�C�G�p�B��k�PjW�i�<٤d	u�� ��j.%:Wc�i�<)�@�(\��s�?�]Ӗ��M�<��l�1_W8h"+-:��3�I�<B�]+�|�a�(@$l�GE�C�<y7C�&;50��n,oJ�p�%GI�<9�� M���µM^$e �0!G�<9���#ڽ�D�ݸr-6���@y�<Y�L&Lt��b�'�K����)^�<�1��8��D!��f��8���[Z�<� hz�؄<ꂥ�%�>]��ܚ&"O���ՂJp>$�P��]ߔ̨�"O�9�J&�΀�堙n+@��"Ope�6�ŕE�u`JF=U��Pg"O��;D	�>��ËA��a�"Ov��Gi"AY�3��V+h��eb�"O��d��`m�e� �0�X��%"O:���燽d7n�;P���ڪ�� "O4������_& h!�̢Y��"O�t ��׺q����L� ж0[$"O�a��Z�ay��Q�����q"O$�8qJ��~,8x�4E_�"��q�"O��r���FG�YC
���h�"O�-Y�EN�d �1ܧ7�n���"Od��k�1����)Q�:¾Q	"O� �5䖾4l�c�c�7����"O⩛'e�p��itHW<n��8 �"O(���/!�ah���n�6,��"O�\1 �`��sW)C:��"O�Hwݲa�Ń5p<T�"OaH�"�2hS���>R����"O���6CE�h���I���&Tc�PB�"Oހ;'$����0@�e��z�"O>@���lonib��W�.�l%��"OP����EPh��J�EIZĳu"O�eҳN�-[�PX��� �
�9"Ojq�Q��Hܩ�*�[|d]�`"O6a�/'q_z����/[G���2"O(싦�FAaİ�F�h2 ��'"O8�x�'w\�Mb7䖟b�:e(3"O�`�AS"r
>���#����Xʧ*O��Pނ����J���K
�' �á� ����;� I��'���EԦ�� ��׊$S���	�'� �`�.)`D#f�Ȃ����'�h�sᑐ@&l�JŬ@�\&��'����t�"|EO�t���'��qD�P\t�Y!�	�H�	�'NIZ�g� �4�������'DЄ�Ѭˁe�X�pF�g|ɘ�'�P �l\�5r�d[���-r8p
�'®�� Ć>�4�`��4�pL)�'>=Aǎ\�}I8mB5��}bH�
�'��8�2o�/+�
`�&�?y�a��'u�U�h�ܦ ��jÑ[��{�"Oh�۷�W#�i��	N�<���t"O��[��ռ{Ƙ+ G�{#�Ī
�'d���gL��8ʥ�ٽ���	�'mh���B�>l�ȁ?d�Y��'X��z�$�	� X��*w��3	�'`�cet��`	"�jp,��'��y�A�m��l�1Ȋ0i�H�'&�ʆbU�uB %jq��'u�B��
�'�T�c��&%ң@��kr�Q��'f��DU�8�`h$�9��8i�'�ʹ�2��!,�z��Ç��86
]#�'@Fىe'O�8��
�M�*����'g6��eӚX���ğ#)H��8�'`2P����rN������D٣
�'����i�6�$E;� �>���C�'�̱/֕<4:\{���r� 5�
�'�e@DO��T���'C�s&J��	�'�����C?~(�Y�i�f�0Q��'�� �A�7�M�k_ �4R��� (uB���~%�����T�ʰI�"Ot�+�#�K�`����^�]�@�
T"O��sk7b�9ӀIπٺ"O�x��"֗�	(��S�L�y3"O.�8D�_�\;0�;'�<7���"O�	Z��U���H�D�*��L$"O(UK%�U!Ft楁�c����12"O��*�摭{�>� �D��"�"Or���	F�m���a����"O��W� ��%	QJW.���[0"O K�e�*x�8�D'�1�p� "O��B��ĥ�&�*�C�D�	�e"O����/Q5u,�وUlv�~��"O�t�����6O8��AH�&���t"O�a�e�Rs5$��"��9)�>�@S"O�E�!�܍t-�	{���}z��3�"O�]Q�o�2_�~�
�%�a�ҥ@$"O��9R(�6�ؕpx���`"O(����]��T��S>i�ZD@�"Of���Rd�����+�"OYʤ�D)�.mӓ'�
����"O`��@	x1Y�&T�kv��3B"OʉP*ʝ>���%q^�"�"O��@�U�t���V�S�T���"O���4C�`�ݓ�I�\?N�"O�5����!dZ"5z��d"O|x���S%B�;!b�>]4���G"O��₆N/jlx1kt�ɽ1)�<�"O樀��Nj q�$$E��}*�"Oh��2 ?�Aӑ��,C@�F"O�0���]j��&ȔR�"�b"Oxt�ǁG!;�̌J�/8����W"Ot�	�@	6FҩH��>"��R�"O��
��w�!��L�$���"Or�x��K�B�a5	�P��"O����mM�R�\�0�j�H�|��"O\ԡ��
4;�j�)ޚ���"O���\�O,^��aȆ�\>��"O���4L ;�4FeHdq6"O�4q�f̱Ǵ�#掆��+n]q�<�Ǐ��RG�%{ � �������Lv�<QS��2�9�T�
�xK"��Q�r�<1�-��9]}�儉-7Kr�x���U�<��M�29\�r�ݫ�H����S�<��(Y�.|�cG
&Y�d�;!�IJ�<��̅�"�"�h �6C��%��C�D�<AYM���(B0kq0����?�!�D��l�
P�q@#
c��ҳl�4�!�\�)��B�$�9\H5���!���\�$ ���,�XU���Ѳ#�!�D�'J�"���ں{(�X�	҂�!��D�|��urcj��-��}��H��'�!���8N�|�s�䆦Q"��%�4�!�D��&�N- B��s�<hv�B+oQ!�����c<|4��ヒ�!�$T�W���H�"mF�Q��J�|�!�dDL�,�!Kcd�DH��!�DQ5=!���)��
.tع�#F{!�d�!���3J�q��$U;A�!��ݚ3h� �v�F�"��9gA*V�!�d�(�hUQ�-0	�j�˜zX!��U>X߾��Ɖ�"���QL׹`�!�$J`R��+?l�s7��"l1!��"�D� ;p#t0��I��:�!�� [��ſI�q���f�&�"Od0���7����aU2"w~H��"OB�ҏ�Z�A�I2��l�"OH�Ӱ���$�@�� d
�0s��cD"O�y�)՘i5��hFj�:�"O���ؠ&��Ȫv�O:��`pv"Or��n�+���Հ�0�"OL���?X��	+��+S"O��z!�P*e����j��݂��c"O�A�
�7h�@Ptj�2(�D �"O(�A��B:Kɨ,�eM�X����"O��ȁJ�|x�2ph��^E2#"O}0@@U�*�;EW�"
h3"O0��   ��   �  C  �  �  #+  <7  ;C  MO  [  Kg  *s  �~  
�  ��  ݟ  g�  �  Ѷ  �  j�  ��  ��  6�  ��  ��  ��  �  ��  G�  � @
 � �  �# �* ~2 �A �O (W �e t v{ �� �� �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+��6!\�	�<4�d5h��'�B�'���'	�'/�'�B�'�~p9�nƫ^wh��Ϳ�ţΊ�?���?����?��?	���?����?�'��C�����FV.E�\R��	��?����?9���?���?A��?���?�5���V�H��re��G�0��%�?���?����?I���?9���?A��?�A�+�~�%��T`p@�����?A��?-�M���?i���?���?I�\< ˢC��G�������t+�=���?���?a��?���?����?��$�h ҡ^���"Z�o|����?���?����?���?����?Q��:�&PR�Ħ}���"'Z�{ւ�����?1���?���?����?����?���-��hUjޞ���y �[v��\���?��?I��?����?���?��.���{�ۢFߊ�*�-шS	|Y���?���?���?����?����?��O�jȲ�@�m�dR��+A��U
���?����?9��?a���?���?Y���R�Z���(�`Q��W9]ø����?����?���?����?���?��#艣��N<�N�����rT0���?���?����?q��?y�i�r�'��)7�)~��u �ψ;$O���K�<��������4-MQ��GJ �H�r���T~�|�\��s���ɰHz���@
�}#�<����6V���ɟtw��M�'+�	��?!���ay0-��_{P���%Z�wT�4x���O���h�`���$���åI�8O��4R�%���>�Il��?���wk�db�,X7��]���2��9 h�O�dr�\ק�Oy���2�i��dW�7-8Ւ7M�	Qp<��:w�r���^@B�=�'�?)U���
���`或�"� r+��<�(O��Ohdn�W�fc�� V��(`XVev�0��NO��g�	�X�I�<�O0pg��n��n�#U$�{����	/u�`���+��u��KƟ�agfD�TD֨���[=$p�j��[y�V���)��<�Aݼ�p�2p�1V^θ8�[�<a`�i�L�)�O.ElZC��|(����X��-a4 �U`��<q���?���b�u��4��d{>�',7��/n�|�p��J:9��.�D�<ͧ�?���?����?A��t��
#����0R�����$���-s�ǅ -s$�	����O���'�� �h\&%�8�d�:��5;�U����4`�6~Ӿ�%>����?��6
�Z�j��7�Ŷ?8"C���-}��p������#R3tr�hBW&�˺��>��<��D�;A�����E]8j�$�'�X?�?��?Q��?ͧ��D�ܦ���_՟0�"$X�3	0IWƟ$y�Q����$�٦Y�?AtV�Ȳ�4+��k�D<q)�d���By����4c���7mu�@��/-�bh��Oƌ���?��7)���ɶ�H�)�D��"DU�t%p���	ɟ,�����ß<�BGl�,�d�@���v�|��C�?���?a�iP,A�O\HsӚ�O�ܙ!d�8,��p��;pht98Ec
]��?�MS��i��N?i�&4O4��˝@-E��+��b3㖈�)i��?A"�9��<y���?����?!�b.ƙ�rɕ0x��K��J �?����$	ݦ�p�/ş��I����O�]���=W�B��ŁJ�q�^MR�O���'T7MJ�!��S�S�?�A�CX&|�x1��@p޲S
te�Y)�#MN�'(��H�48��|R��w�8郗dSAb����I�s���'m2�'���4T�Tb޴"�����.�#d��,����6�K\ ,\��I�Lh�4��':������=z.��r擌D�`�9b�z�6��]C�d�㦩̓�?�Ci�"�z��̑��d^���`��G�M����Rd݆6I�<���?����?����?i-�(���W�\x�T�*�Ɲ#e#�����v�Jџ����� �SW�2�M�;x3:�)�(��I/�y����V��w�'��v�%��O����Ov`A�iF��©c�$���+tJ�(��c&�D�+n�:�J�Ol��?���W&�0xӂ�Mt(��Ĕ:8�ƝH���?Q���?�)O��l�zi����͟��I�,�d�����X~V0�DD2*\�?)3R����4����3���d^R "�G "&DY���,y���O�P �/��1B��<I�'i�f��?�%��4�Qy��<�h���Z
�?���?����?�����O��3��X$Xh$\����p�Ĵ0���O�!n��ԑ��؟,��4���yg��h��L���?i�&�K�J_4�~��i�6-�E�6�̦�Γ�?���"E�����j��(7��  q�3W"�=_���K>9/O��$�O��d�Ox�D�O�"��[�T� =��*�2k�<2C�<e�i�~�P�'32�'��D���E�xMP�8�O�@e,��bQJ}�ne�pn�$���|��'��r���M�̙��
sX@ih�&�.B���f`��򤐛<�D�C��:$�ON�RHv�+�)Հ�������	�������?9��?���|�)O��oZ�Kkt��IcL��!�ߪF��a��Ӭ��牔�MS��G�>���i@6MG�m��+�j�0$��ϟ
y��a�%N���mZ�<�1/;m�`A�G��ba(���^w�<�� &�j�@ĕs��1$�#H�NQ�T;OF��O���Oz�D�O��?E�c͍~��u��;H�qjD����	��<K�4$�x�Χ�?�'�i��'?�0��i<X�p��0|��a �#+��DĦI���|j�L���M��'�( ������:�DY��Y�%<�@��.�O�A�O�,�6Q��������	ʟLc7N�+��A�t&�E�UXq������^yRCfӤ�[���O��$�O.�������$�؍U�R�
p/�	��)� P�O�m� �M+F�xʟİA�@ĉgD��j�茰�l�(�b-d�+���+1�V��|�ԏ�Oڌ3K>I�F�f~,-yW⍵T+XA�?���?y��?ͧ�?y�R
��$Q֦�1���#�8�8�aX$ ����-4{1��ȟd��ɟؖ��X�Xc۴YY�L�n]� 9ڗ�4�8!�ֵi��7MG�}�d7-2?٦���I� ��0���EQ��T�0��=d�2WE�'�yBX� �Iܟ��	蟨�	ɟp�O
�<Y2 �"�A�SM�!7�!�bo�F`���<���(��������]������O!�Ј���Ŗt܅����M�'�)����,'"6mp�h�v-�:dƵO�$%^���|��s�J�'>�b'�K��gy�O��I�A�Lp��! ���CP���jZ��'3r�'�剷�Mfk���?q��?1��Y�td�Mц�Eq��Cp��<�?AO>	a]���4M���H.��29���e+�/  r%�A�j��I2Xw�{�ܑ*��Y$?ES��'��Y��p�e��E�F����&(�m�	˟�	����C�Soy��'Т90W��3*�ݪ3@Ь`b��'S�7Mĺvt�$�O���*�d�O��\��-�՛N�Bl��e@5\&���`�47����$��f9O���#\TpC�'S�P�2e��^D��Kv�o��`Yq` ���<�'�?Q���?Q���?�s׹XG|�Q ş8Jb
!Cu�P���DEҦ�@/�꟨�I�$?���bB��@ǘ<~jx�*���9���(�Od�o�MӜ'ƉO����'�M�1HF�H2�cq�N&�2T"�#v�dT��O
e�RJA/�?�c')�d�<I�`��O-Ĝz���		.0�Nص�?!��?���?�'��DĦ�����0�M֦�ꭀ�&�;��8��e\��"�4�?qO>�TP����̦%�شF} �"S��o~���,�G�Qr#
?�M�'F��^)k��|�S�����?1��'��T*��B�$��WF�՜�	������	����v��R��9�$��xY*Ͱ�����:-O�����	x�w>U�I6�M�����B�I�j-�!DؾJ�\�0b�; '�8Qٴ웞O�T��иi��	�b��]��N#:��ؒ�'����L�(�rn�X�	]y"�'8��'[r�Bmp@鵫��?9T�i��+`2��'�剏�MS���6�?y���?�(����႘�����Xӆ,H盟؋/O�DdӀ�%��	����qR�D�b�@p��NX1=�$q��3��I��� ��ɷ&�n�1���?�`h8}ZcA8y�n1����.����1P��'���'����O��I��M��{��Q�WlPf9�OM�\ ~����?IǱi�O�u�'�H6-Ly������RR���J"%_�n�l���M3b@(�M{�'��̥4�����1��	7�0h���Ż9l���H(���fyR�'p����l��`��Z��NI�����'ݼN��Bp�щ#ʦ6MѽQ��$�O��d<�	�O�4nz��׬�(U؈0��,���飷�K��M�i�rO�)�����6�P7-f����g߇oZ���w�Ȅm��1�jj�\�&�3|�c��sy��'����r��x�Ŭ��dm �����'�R�'�BU�۴F�F�8��?���$T�	��\I ��p$�h0�d��/�>	��i26mQ�*|Dz���4��/�0w���	���Aj��B�Ar���zy��O  ���$���1 s�4��M9�Ptz��ד=i��'YR�'���՟��BV�e@�`0းQCt��D���޴}�� ��?���i��O�,a����!Ӳ���1��6�d�	A޴&���G���v8O��ā	���I�'n�l���lˏn��u��w� �:��.���<����?1���?����?I`��`�u�f�%���Ч�	���ܦ���`����I�&?��ɲK()�ǌ�!�A'"<	'����Omڶ�M��x�O/�4�O���Z�\ �tÝ!8�^���J�qŮMY[�{A쏜(��dI|��\y�L��N|pp#IV�-+-��[�b��'�"�'d�O(剌�M��F��?��HzK��jN�I�)�-E6�?���iJ�O�-�'66�P��ijܴb8�0r�� Մ�X&ɋ:��i�U�M��O�@J��\��"!(����x�1�IŔ[���9��fy��1OV���O����O����O,����D-p�N�xS��d��D0ŪR$���d�O���¦qr#A������ޟd�Igy2mܥX�Hk�L(l��x���O���7-�P}�Om���mZ�?���F����?�6.�G�D�D�e���a��ޠ�xUc�dNLt��Y������O��?m�	۟`��}P�{��+S�����R�#\t&�J(�����>��
�.Z�31R���h��%�M��;-�|h�-@9s�΀XF@R���ly����4S	0}s�'�°i�D��p�~�!�Ow�d)	b2�)���>��;44P��1�c��dG@��OJ�I�8�?q!�OD�$8|,+��_0k�i����uLV����?���?i��|*��?	*OЄl�aArл�	±e�����L,,;fhi�����	ҟ�&��]y�/}�8;C�I�_F"����ES�ĠV`��)��4Z�P:�4�y�kXBJp%#�C��?Q�'�� d�c�[�F���+Z,/;"�3Q�iw�)�	ȟ@������쟜����`��Ο��%K��W��-���ڻX~���*A�(M�����|���Iޟ\B�4��7ͦ<�īW�xyP� �$
0of�q��ݿq����o��<m�7L;Fd���?���?�J3f�ЦI��RrdZ�dXp�,N�軂a|��H��S�b��~�Oy�Oc����j�.��RfJ.Vm2�[s$D�oFr�'KR�'k��-�M�S��?Q���?i�E���#�*H�a�&q�Ҟ��%���w}�Dp��nZ0�?�O�L����V�n���rc�<z��A�'%��:.vZ�Y�b��I�?iA��'s�E���P�N ��X�*��Pз�����������Ο��In�O�C��.^�q��Ջz�4z���<2�}�r-K@O�O���Ц��?ͻt��T�N�"��P��D�!&���1�V*v�%n:u>�n^~(ў!kD��S�
�~��������ݠ�/����������OX��O����O\���wD(�JІ�(e(wK	�A��^�Ff�0[N��'��)	+jb �G�#t��7LE�?����'�7-�Ϧ���S�O��Ƽ9�йcKܵp����e�P�K�h��pX����@�2σr�[y�b]M��zR�:f㸝(��5Er�'eb�'Z�O�剽�M�wH�"�?��D)���`�L�T��:�bL��?�#�i)�O�L�'��ia�7����׌y,U��C[��N��3,e�@�I�������/|�įbyb�O���sb 8��N���37L�GV�I����I�����ß�����"���s'�DL��d Ê��.u���?��!�����;��)��%�����4�&��!��(+�$�2����?I�ODLm��M�'Ke.��ߴ�����I�
(�	�&,�0t!ǍzԲ])�ŀ�?12�*���<����?���?a�l��1_D�Yb��40B�X��>�?����$R�ik�n�͟��IڟȖO����+�DJ� �iB���k�O���'�6��Ѧ�J<ͧ��pc"{��w��6������ �7B)2���A4��+OD��X��?�d+&���*XB8��cF7��U�۫I
t���O8�$�O��4���0l��H3�ʓ7�ż	o�)�a@�Z�T	+�e]2e�����'r�'[ɧ�4��l=(��ېE H7b�ز/�rX��ڴa�& H�F@�F1O��$��/*Pe:��ry���>�ąP`aH�HN�	6�N�Y`��ȟ���۟(�IğH��ןt��ӟXT�CP�ؗ)��`u��D�ˬb~c'�
�.*n��h����	��MG���<��f��|2��)Pn�Q��D�|��}�l]� ��4�MSӿi�����@�$J?�o����m�<Q�H�n��`�ma�L��<Ʉ ;m���ݖ����4�����?Z&���	/�<����/X;$���O��dN���O���l�W����'��Iٓ��� Ǐ��M�l�)QA����'�rP����4(�&�v���'�F髥
�Eq@�B���=V�<b�O��R���1|$j���3�?yd�O�X!<�|����1
y�d�O�D�O��$�O��}r��9�y[���U�8���,Uv!��AB������'Z�7m�OB�O��;h��Yd�]YW(� F��*��dܦu�ٴ!*���=sS�<OZ��
c�,��'g��P3�e˭z.�Xs��Τz�F|a�#�Į<����?���?���?��R�Фp�	�}���*������ĝ�C�i�����I�'?���>9��&�Y�IDHC+֪V�&�Oҝl���Mk�'~�O����'͢��&cB1zH.Q�M4a�!k%,�KW&���O�X#�j^;�?)�))��<9!��N��A�Fb�T\�����?���?����?ͧ��OӦ�GaMɟ�pP��*l�r��砊&\�*As�C�̟8��4��'�����Gy�h�d�%U�0DZ�h�54c��+i{�<!q�o����|p�AOH��4h1?��'�k�;!�x[���Uj�H@#��<%s��O:��Ob�d�Oj�d3���Pq���2�`Ķ�x�΅)8�� �������Msa��|���1��&�|r�G$RSZ�i�o��0�=�����5a�ĵ>q��i� 6m�OH�˃�s���ꟼ�ѥ�
ph!� W¶�*נ���
Չ��'9�$�ؕ��D�'���'I��A�����1���]0X����'�"[�@���N
ҹ��ퟔ��L��K[1mT>�j�křo�Y�\�T1�'�T�[��'{Ӥ�IJ��?�7"�?�Z,8p���V���a��z�ЮɘO����B��O�@L>y��L�p�\�idB����M#4��?���?����?�|)O^�n	����"Tr�@ ���kSZ�(3'��(�I��Mk�B�>!�i�JU�$$yGЈz�ֈ�ҹ�%t�.��K?�7Mo�����h\��y��O.�|�$�kg�[�0�by�V���I�<,���d�O~�d�O��D�O���|J��߈<�nL��'�G�|9``�ӻt �Ɉ��?Q��?)N~Z��g��woȀR橖$/x��@pc��x���"�"lӼ�n��<��O�I��D�$��{��7-u�X��L�\I�Yx�
 n����l�D�U�ډ51b͛n�	Iy�O;�@��}���`�+E�$:Xr%J+\�'�r�'��I<�M����?���?�2J�v0���i��Q^�`ˋ���';n�&�ƭs�J�	m}�#CV�вi�y���0Q���y��'�&@�ǈ�>*�I�O�����?ْ��O����PB��4h�k�:\�lpQ��O����OL�d�O8�}Z�PRR��F<4����0mT\ma�x�&��V���'��6M'�i�Ua ���8n͚G X!c�hyj��g�8�۴5����'��!#��i��d�O�S����B�� f�"t͖�&N����I�4A�@I&��<ͧ�?Q���?���?i �֤Q7�q��'��)�R8�'��)���ٟ����OB�D�O���@�DٱH� 1�4#� c$��RD͹-���'�7Mߦ�!O<�'����t! D�������wn����'R>�h*OH�)C��?�` ��<��C��p�&(H5D~l�s���?���?���?ͧ��$�Ǧ!p�������> 2|4rjH�yR��ʟt�4��'��b����m�^�lZF�\��J/Z>��sDLc_��ó!KΦ���?Ic������$�P��\�sv��2"��!3�h�D��z�D�O����O*���O��$.��u�,@��.�F�!�,|������I��M����|����v�|Ҭ�&�ڕ�bg��j �x��O��m��Mk��pC$���4�y��'���p�<I�+]2���kY�e����I�m=�'��	ϟ��	�� �Ʌ�$��'I܁tؚ=1�F	zЎa�IΟ �'�7�zz�$�O��$�|�e
	d��VC�7f��{��Mq~���>y�i9�6����^��P�A�j��	�8Ȥ�10/ГlٞE���J <�P�{Sʣ<9�'>���$N���G���y�@�(vR��ŌW�~��P[���?A���?��Ş������s�V2����!��45��d�]w hM�����B�4��'���|��3ppX0ԏBS<�XH'�ހm��7��O��c@�i��������г	C��#=?� ��p����&�'|Ȯ�W(��</O��d�Or�D�O0�d�O�˧6$1��^�P�����E1}��Xh"�i�ܙb5�'�b�'d񟦙nz��Ǭ�!�	�u�<l���d��!�?��4C�ɧ�1X��޴�y-�)Z�҄�r(}�\�2��#�y*M+�����.��'��I㟀���}ZH	g�[".�$���-�l��؟���͟ܔ'C�7��:ZCh���O��$�PZ��W��0�5��-��$K�Oڡn�;�M�x��J�^�F :6��(N��`
��C	�y2�'=�,�$��6-Z<옐Y����L�RbB�����
*�`Ǉ�!b�I�ן0�	Ɵ��՟(E���'9@��ݎd�G�"&�b�R�'c6��?%�l���O �l�Z�Ӽ�׋I�#k$�(W�B;J�!��R�<9��iE�6�Φ�#wK��1�'6p4"s���?I	C��%�P�I3���,.H��Sz��'+�I���ğ�������69R�a�HBS��*<y�a�'Yn6-��:H��?������<�qEʇH�� w(_��x��ױV�	��M�iL�O1�иq�FŹ(�@$�ԁ�ryB Ǚ�����<i�I��e|�$ʫ����d��/�U��'A�6[(�� Җkx�d�OZ���Oj�4�B˓?���?y�'�B4�u�V�}8�/�<1�i��O^@�'��i$6-�=W�щ�"�4<"�pH�o��^Dl�3Etӌ�S��E�����I~���q~���f,�V�p���;U���̓�?����?���?�nZP�ӈ@�`@Քy��x����@���32獸Y��\�����4hR���?Q���?�)OЅ��D�!y�xkת��[ж������ڪO*=m�MC�'<%F���4�y��'��-{"Z�v9
�J�Q���.�4.�����J��'�i>5�	韐�ɁS1����.d�4�'�
e]� ����̗'
�7Q�5p���OV��埐��R���W�Q�|�)�d�I%�D�O`��?�۴F���)�)��ֽ���)�� S]`a�q�ݟ���˖c�E����OV�i��?Q��3��S<}�2�Љޥ��G̜�F�D�O����Oj�4�����O�ʓ^�6G$��CE�=V� ��kx��yH`�'���'��'��_�LH޴ .��CL\.s��"�&S�u��i��7��� �6�>?q�Үz���+��O��de H��s���0�^� �?O���?���?����?1����� �M�t���A�_I����H$�ަI�-�Cy�'�O��r��.�(j5	�%�V����C�}�9l�3�M�վiJz��|Z���
�#���M��'�B��g	�#% ���䎍&qX}(�'� �C��	�N����'��	�aj��%��=8U�K�y�ԱV$��B�h���D�fȓ��?���?Qư�x�hAg�O6���Oh�q���J�o�V�
4n�OH��?�����yR�'����j�hͮ;�?	�ӻ[���#�O;J�d�`�Mq~�*3w`�R��TԘOK���T��LX��6bh֜%��N T���'�'�r���xa�A�/m�صA4��+���
p��ԟL�4R�d<���?�Ӱi�R�|�w�m���� �z�A�3 �j9�'śvh`Ӿ�$NF}�6c�P�����E�O3�j�N
�\�ʄFG�w^�ТO�h�ly�OSb�'���'�"D#�NI��H�&�Iz�aտEg剃�M�j���?���?a����)�O�8C#�^�0�R���`@�)h.��-�s}�foӆ�lZ�<a��)
{j�B�m_+y�@I�NV�~g^x�q�,@����b1�`�f�'�b�'�t�'�sdA�;��1��Ǜq��E�'2�')���DT�$8޴K|��
��/���f�	#xUT\z�!�X����}W�6�'��'Ҭ���LsӺPl1X�d���V5(g�%����[�(�٦iϓ�?)t@�s����έ�����R>ᩖjB5{p*�Z� �T]���O��d�O����O���+�����������<p�7_]�D�Iޟ�	��M������D���$��akU,
���ʆ��/k��2���ēO���k�l����wB�7mh���I��R� ���@@K�C������o����f�ݨ�?Ad-&�D�<���?���?�-O,rV���
�>��ѩ��Ų�?�������������	ݟܖO�������I3�L�viE�9Pv���O4��'�r7m���u(L<�'��I�}����Û'�����O��}�<<�1�І<?��(O���B�?�6�)��^y�X[ҭ�=
GR	ԧR�(L�$�O���O����<�Ʊi���0t)�0�|���·?�vy!���C��	�M���>qW�'��Y�Un�&+��q��fK�l[nH��i��7���<'07`�P��.s2��OT�T�'�Y�@�P�,4Kr� 4[&��
�'��ş$�IΟ�������@��%�T�J��vJW=/v ��#�&4{�7��>�J���O���+��>�Mϻ2���7J�"���E��:�R�*P�i�L7Mh�ק���O��̾���=OB�r#���"��᠆�4�H��8O��w(ԙ�?9A�*�d�<�'�?�iՑD���S��X�~IK�K��?��?��H������[�*��?���������2\�Y��Z:O��;�9�I[y��'��I؟<lڹ�M�gW� Q���}�+�J�E��8��q� �I�"ߠ�Q���C����j��O�K��H��	`"@#ʔ�RXz�UJ�����ß��I韨F�T�'ɢ����YC�v����$o�nYa��'��7mB������O�Am�f�Ӽ��a�b;D��(�g\S%��<!�i�
7�٦�{��ܦ]��?I`�O�A�>����Dzn��%J.�(ar��D/Q��BL>Q.O��O��$�O�D�O.�"u�ԎO�r���;]���Ӣ��<�Աi�q
��'1��'��O3�OGlZp#$D\#;��M�e��v��?��4)����O��6�$n��A���CB�JT|���D���.9�X�$��O,=RH>�,O��eDj���G���r��ai��Ol���O���O�I�<i��i�v�Yv�'��̡Q��>�X))�gO��tZ��'�68�	�������	�۴e�V�/C���ք^ՔYjT��'(eͱS�i��D�OhY&��"�:',�<���0�k�R�jlT0H��MN1p�gK,v+�d�OX�$�O��d�O>��'��?B�mpsɢY����IK�(���ǟ���M�Rā�|��Q��F�|raE����D�ӡ^:�i��"��$�<��4>���O��}�6�i��d�O>�!����JU�@ĮoE��i�J	-YJM8�FޒO@��?���?	�{A�,M*,2���Ч0�8����	Cy�vӴ�K%D�<�����	�~{�]cG�\y�����H֥S�	3���O�7-u��J��#X��q��C�>*�i���1P^1WkJ�`���b�<1�'9��[wv��<!��*g���*�qV�xk��?���?Y���?�f�?���Q%�?��2���Ɣe�<��b� d�\�- ��$8ԝ�Bs�����'���'��a� (�ǂ4*׮ ?1����V�����4'�c�4�y�'��$)��P�?���OE��8#��p��dx���#m��d�<���?i��?����?�,��pAGC�7���i >dU���BOѦ��� ]ß�I՟`%?�I�M�;S”2��yҶ �w�F<�.�0`�i�6-^��Xէ�D�O������4Ozi��) �$à��t��bNT4ʶ0O���?���,��<1���?)�H�[R֍P��\-��u8'	��?!��?�����Ҧ���ş��	ڟ9F,*W�t(:W(T/t�
a��S�O �	
�MS0�i%T�T>��lA�61�Va�<C��8��w���I4mI"l�≯3W�ٕ'��tk�ɟ$���'%`���W�[y0\!�k�6&�=@F�'���'�"�'�>��^�Z����^8��4�R%ov�	��M���D�?���0��f�4���q�Ӻ�,H 0��=1wlt�:O��o��MSW�i�Bm;��iz���On��Q�C�zq���>h��@{.�)�u��u�ƒO���?Y��?	��?����DB�B�0z�{Pg��V��	�+O��	-[^�$�O��-�	�Of��c̲V��|+�3�\���PS���޴2ЛF3Ol�^���O6�Sr�̂�0��E
5u��Q#�\k�-�P��(�ю4��XF��Fy�տ� ]��78ZX؅��&�"�'���'�O���M�7ML��?e�ܦ;��a��Qd�.�����?���iG�O�`�'h�7�N�I�(��r��;8�X���f܍�$A���ZΦ���?Y�Ǥg
D�		G~2�O���3V�Yx�h�!hp�'�[m���ş����<�	����{��sL��Չ�"�����j[2$�f *���?I��K��A����d�'l�7�3��O:;R��e�?=�T��wR�+k��IA}��t�%l�̟���ަ���?��N�0�5Ԍ��qA�H��T�+Xִ�R@�O(���D�<ͧ�?���?	��^KV�3�n؅l�9bO@ �?!F�J�������13Ԋ��?����� �Ohl����Z�.�����#���X�'{BW�(�4T��F�t��X$>��S�w�XC�C�)�p8���H��yW�՘G��d�Ҫ*?i��$���dV��?A.O\���7{�;�IԐ9Z��d�O`���Ot�d�O��۷H��h�v�<qd�iy�	
�$� r����s�#1f�`�6PJ���$�L��qy{�BUx�P��`5Ȍ�@��ѓ"HĦ	��4���ߴ��dYkҴ������4$5��S��[
���$�ǜ*f�	xyB�'E��'��'��U>%����j��	3P�lxA/ƩQiL6̌c�|���O��$�2t�D��<Y�Ӽ���,�jR�[�i4�<x7m�zo�f�cӄPn�����i��b�6�y�� �Q ��� mn��4���d� 7O� ���S��?���/��<ͧ�?����д�Ah	Y�PI10IJ��?���?������J�遡���|�I���H �.�*�
sB�/��;�&~��m��	7�M{ �i�O���gI9q�Q��B7(��0O�iި��Ci��k�a�R�X��-K�҅�ڟ��_،0zP�K!�px��`���4���p�	ǟ�G��w��<����k���)�7;��
�'d�6-\X>�D�O�mZ[�Ӽ;v��e�DA�fG�L8�v��<Y��i�6���e��l�Ԧ���?���z��	�~Y� ��nFޕ*�j��d��<�J>	)O��?�6LW�F��ˢO��)�����$P~�g|�Fq��c�O���O��?�8���0O����M�M���ǩ����Hަ���4Y�J~B�����#C�4�$j�Ie8|S��Ű�������D��ij^ ���0�OT�
�t�#��kcX�[A�[t���ɂ�M��/��?�E��	:� �����h-�g/��<�2�i9�O��'�l7����:ش���س$,���B�!Q�.�\�uL��M3�'1�!}$�����5���?�]�,1l�Q�mB�u�r\�� K�'B��I\���ϽԖy����V�AǇZџ���ğ���4P��T�O7f7$��M�-'t���K��2��x�+��M.����O}�+f��l��?3��\�}͓�?)��@	��i������Sh�.y˚Р�OԸ�K>�(O�⟔SA�H$�a��FX)o
�#<1�i̘��'Y��'��S�l�؁�	ȷu0f���örg��{��Ɏ�Mӽit����t�Og��y���xuNT`���[S����#��f�N	{��Ă Q��?1��'�p$�p�s.�1A���b�DD�R<y�6�2��"۴Z��"�
,-$�`a�=o�&�i�C)����}�?)a\����4|���q"K�L�X�0����
�<�y5�ib7Mҋiz>6�s�`�	�X���"W�Os�e�'�xl26 T4v)�e����]n�{�' �I�� �������̟��	]��н dԱV΍��`�1t�R�~�:7����˓�?L~��W���w˂0�gF�QxL��wBP4;�L���h���l��<	�O���V�$��j>7Mz��E�%*�	��A	P�"�$�p�p��ؼH�-Bj�	|y�O2mB ���,U��k�-�5i���'�"�'��	��Mӗ�����Oʨ:V��[�Zm[��=jz�bb�-��;���	ߦ���4�yRX�� p탠%2�H�A�1y�:�t���I�t�ơD(�S����b��OB%����P���I�+�N�� 
Z�|��z��?����?����h�����Dp򩙥)F�'���4j54���$�ܦEh�ß����	��Mˎ�w`@����"5��D�JT@��ț'.r6N�m�	���o��<9�WJ��D��)�.$8��=r�,�J�HI����%����4�����O`��OF�@�D8R`,)t�uFټ<�4�H���I�43��˟�&?m�I�5��q����2��[�O�=R!S�OάlZ'�M{�'i�O���'�ة+�LRW��)�@��(Px���*DS$)�O���1`�>�?IS�*��<����h���EN$��KE�&�?��?���?�'��FϦI��,�ş [q�R�]�N횡 T�E�~a5k\�0�ݴ��'�v���fuӎ�����|%���Z�60&a�dK�̬4��d���	���ѯ��F;�tM1?y��o�k�4C�X�%+ݦA�[�CA�7��d�O��$�OX��O���>�S�Y�\��)��T~�ٱF�R��'*��i�@��=�x���Y�Ihy򀒂/i�]A7˝�}�V$�_	��>���i�87�O�h)��e�,�I���d̋5*r��h'ֶV����"
�*�z����'Xbi'�������'�2�'r2|�"ȋ  ����Npk�a���'�]�,I�4'y\D9-O��ĭ|E��#Kp��pA7�r4�o�P~Rä>�R�ib@7r��$>���;�&d���lN�Cd-R�^B�G��.�T(@D9?���Y�������1r��;S �#'T�"��!=^�[���?1��?1�Ş��d�ڦ�@�� y�z���*�\U��N)��蟔�ڴ�?�H>aRU��j�43E��H�*wz��!�f��8�i��ș���V3O���Q"S�l����X���\Cfd��t������0&���Iuy�'���'��'0^>e*���n�&���Z/fd� HR.�M�!�-������?��'����?)�ӼS�����9�`TO�	�J�
U]�vb`�P!l�'��4���	��^1���kӌ�I�A��[Umݦ6�JT��b_9L%��	�U���*���*5���	@y2��uWӟ���ǽB�b�q���Fkl,��ݺ3���£X$��a>��d�O���;��!�'�?���;b��:!oΆ;Y,��Ϗ$�� �K>�¿i���)�M�׵i�̩{q"DΔe7N���^�hH�`��V?�yb�'��m���sl�K�O�����?�n�Ox��F�Ґ� ��f�;��0r��Ob�D�O��$�O0��&@��n�O~�d_%_��<�a.�}cr��b�R9T���d�Ŧ�qJ��T�i�M�K>��Ӽ�"ëOKz4�b_�z�Ԑ�dɜ�<��iT�7���aPL	֦	ϓ�?�����^�����+$&T~�Є�v��,k�]��L��䓭�4�����O�$�O2�D��[��'EʘI��x���ݍ:X��9z��ވ^�):��'R��O ���'XBKJ�@x��lYV `�d$<L����nZ�M�0����O��O�+�� �D�J�3�\�A����DK�!^$���!p]�ɖ�' �m$���'���b�G�?6}FUcq"��u�����'��'v��'k~%��R�X��4+HZyH�'T�4m�`��<���fj
��ϓ�?�����$�Oʓ=���Io�LMnڕ�$�`���M��Y�A{9�ᮞo���1OR�Ď�'��x���0w���?Q�Xc�:<��� 1}�	��LHP�'A��'�r�'��'Y�O�R�ɨJ���̕:}O6��hbqQS�'�F`��!s��Oh�d�O��$�<��� 0P�FT���B��T�QnC�L}�ʼ>�d�i��7����a�o����|�G��Br�Ib�g�dd��oX�UI� j$�'c�$������'x2�'�ĕ�R�G2g���-T�8qV��6P$�T��+ܴV��x1��?�����;k'��hGJ�/R|�b�ϱ[�y��?-O�El�%�MW�i��&��
,���T~��U��HC  �"K*Svt����ӜP��/���l�'X4(��b�Hyɓ���3���'��'������!ʥ��]���ش�h�DJ�j�ܩ#*�D�D��S"��?���?a������O�ʓ*!�M�m�@[QE�-2�j���/�i��7�TӦ	ۡ��Ӧm͓�?��T
>�N�	�M~�� I�x��/Ւ>�P�ч���y��'�R�'���'��'���'|�Q�b7����>,cn��֊��\�����Eڣ5A"�'��
n��-�6Of�d�OP�j��8C�Z:O����D�:��m��M���z˸��|
��O|����X��f?O$P� �N-�,�u���zc2O��a�i� �?�W+;�$�<�'�?�GŁ��z� 	)y��� �s����OJɳ��Odʓ&̛�aĄR��'�є,��Y �V,T8�J���u�':�V�(0�4@��V�~����'�"Ă�F5~I8]e(�x�HĚ�O�p
���V�x�����?����O<�	�ʘ%$G��1u�Z�b��e��O����O��Oj����ZR"�O:�Ĕ!(�HPP��!\�b���o�l�d@æ9J�����ҟ��cy��y���)��pq/]?#>t�����y�n��o�M;�K!�M��OxX��/��7��umF�f��B' �l�1 �*�O��|���?����?)����jf�ȘLJDx�"�3p�
]�(O"Tmڥ ���Р�ǟt�	�?��ȟx���>�48��)�����٦(��X�'$�6M���Q�ڴK8�O��d�O���9�IS�"�2�� ��P�f��%d�	c14}B�O��*�k�*�?	��9�D�<1T�l��p@ m&)�h�����?��?���?ͧ��d������i�ȟp��D֌;3x��mP G�����R��X�۴�?H>�qW��QܴlF��Mk�n�,���A\;;t�*���y�
�QFAz���	ݟ�q�-���*�hy2�O6W�&n|x2�̖:x�(H��y��'���'���'H�I/,Ft�F�V��bD��*�`���O�����5���t>���:�MS���DK�gWʑ�CΉF��q�C�	56��H&���شQЛv�O���;�i���O�D:W���(�bU�&qB�wc\3o�Z����O,֓OX��?9��?Q��������2(%�Х.H@�����?�*O`em�?8����ןh��e�$��'{"I��L9$��Eo����U}B�pӤ�n���|��' ��=��LE:��H���|��EԚԱ��/QA�Д'N�te͟|�C�|���j������3��,33�^�B�'���'���$Y�pHٴi���ie�|9��!��͜s^ޜP��՞�?���8���'K�'rʓ�Mk�ƬNZI��.V�q/�	I�V�i��A:c�s�
�IßhR���
��T�Xy�e��"t�: ��!V��ӁjA�y�Q�\�	㟀��Ο���ܟT�O���Z�C�e��h0��;��D��
{Ӷ踢l�O@���O��B�d�ަ�4&\	Z�Z�LѺ�[�H�{)<���4qϛ�B3��	L  ��6m~�̲�ƴ���7(�38���@�Kp�l+��ܹ�2N]_�yy��'�bɁ�P!JT	B�dg����hƵ��'�b�'��	�M��2���O&i�� NS���R��'��9�`3�ɼ��^ۦ1��4Nщ'���bfɑ�
���g�dEh�؜'����K���@d��{���?����'0�=�I;]6ʧ��0j���@g���<����ğ���t�O��*-�J����(x�����%�B�w��YzE�O��$ަ��?�;46>�����,�K�N+���̓����pӠ�oZ�W�&po��<���r���C����:��J@)z�$��%��xQ�aK�������OL���O����O@�Ě���0G�L��0�i��*)���"����&U��'EҖ���'�~��4�cW�5�G	GnN���Χ>� �i�x6Mi�i>���?�!E�pf�(��ni�.)�E�6A�����by"�\�������'��ɧr��P@��#�Ș"��y�V���Ο��IƟt�i>�'9�6���R*:���WE�h.}����:| � �'^67-;����$���q�شZm�6�s�dUq�L/#d��3M�?v�����i���O�)��ި�Z�.�<q�'��o��^B(A�	6^Jdq�Ձ��<���?���?���?����G׮w�FT��o�&��5e����'�B�hӶ�)F2���d���$��D��&��#`-�w��}��BP��ēC���n��I	&��6�,?i#�áB"ܠ*�����J�e9�9u"�Oơ�J>1-O���O����O��*�D�H?�%a0@��X��x���O���<�i& �Z"�'���'��S�*)N]2MW2S��ո����i����;�O��mZ��M�T�xʟ� �M�G-��'ƔU˰�Nv�Р1��h�x�
TKN��h��|����O2��K>���p�~��ƀ�2cƐ��?	��?a���?�|j(O��nZ+89��9�5:X萁��%��B�ƍߟT�I��M����>)��ip���&��i���B��bI(M~ӌ�n�I��lj~���h������b]�I�MUxe�`�».�@ƃ� x:�	fy�'&��'���'�"T>Eh�o(D�M�@\��H�Q�M�ʶ�?y���?�H~r�蛞w��سA��`L�-� eݭn�~��#i�(�n��Ş>�R�4�y"���D��7DC�	�-1���y�J�za>�Ic��'`���L��>@���;"�G"�`�-,v���	��,��Пȗ'��6m�G�����Oh�DZ,[;�Ո�l��ań�а���;�㟼p�Oh�l��M3ƒx"C�4 V����Ϟ	m�
��!���ܟ)|\����L�撟8H���C�f�DR�X7"�y��H����R��l�d�O�$�O8�:�'�?a`�
>(}|<	 F��1�[��4�?�C�iѰ%Z�'*R�r�����p4�����=���r� ��g�>�� �Mc��i�7m�	V�71?��H��d���IE�F	�H���c��A+Ҽ ��EhN>I-O����O�d�O���O��Q��7/���τ5߈�#T��<��ipT��f�'	��'��O¤Α& �LzD$R�c�,s�\�ue��r���Br�F�'���?y�Sq<:���Y���)�A�L5�@E�)RJ�'!2up2��ڟ0)��|"R�血ė��
%���1(H~�hD`�ןd��⟀��۟��Fy,iӌԸ��O^q	��Z2��ЦHH�{/r�����O��l�\��l5����M�v�i��6M����"�ΉB��ڧbP�d��-}��П��@�R{��DMy��O��\�g����͏;B⚄��#B��yB�'��'��'���)?k�0V�ƨ1l�@0��6&��d�Ot�d	Ǧ��Ac>	���MkJ>Q4$�r.=� ZB�dL�äIG@�'�"7-Ҧ��S}e��m�<��AC�Z�C�&�F��B�N�hƠ�$�V=���������O�$�O���Z:Ed�ܢɈ�,u�#w�ۚ � ���O�r�f�2)�'�]>I��g�K
QbŊ�4�R�q�l����DӦI�ݴl�����_,�x�1���&xW�U�$� >Q��sA$�f�j�Q��F:���U�ɖJ.���R�z�9"mS'�� �I�����ڟ4�)��Ky��q���YE�s�T��B�B����1z�]��'^Rt�8�O���]h}��x��u�eB��	x� ��F$��=I��	���I�4K�Źߴ�y��'8R=�S� �?��UY�,�B)���(IU� t���oj�(�'-"�'���'��'B哜L'�(V�1#�A�ת_��I�4}�F���?�����?��y�B̫��$$V�k@T��ND�b��6M��������4���I�(��e�P�	�wZąbG
�I��m�FC�$9x�I*v�4�d�'*�x'� �'�B�'8 l�whņ�(��`�_�7jX��'���'��T�̓ٴ
�0U.O��D+d:$�Ԃ.��D����ޓO����^}|�N<l��ē�R�ԂA
0ɆM��@�s��Γ�?ّ,R$&l�-)��۰��D�ָ��h�\�$�C�ⱑf�Y�=d.a҃D�\�����O8�$�O���)��+��(�ȓ��H�q�&�$�?�@�i�ԤC�'��oo�(�O��4���Ш\06�x�A&T&%7`���=OJo���M��i�\Z׻i���*Mj`"��O墥
^�G5��&gЂZhh��c}��CyR�'��'\��'��/ש����a	��2�^X��dC�d�剭�M+��?���?�L~�����
��əSX!l��nMb�Rp_��۴aś���O�O&���O͒Mr��o`
���e+�a��W�zXs3R�LV�L��̍[�ILyB$T	"G�T;e��x��0�b�JR�'���' �O��>�M�&K
%�?yw��p0w��*ڊ���� �֛�!n���O�� \}R�{Ӿam�;�MV�<x�dN6Q����c@"zP`�4�yb�'�`|Y�.��?Ex0T���S0�56�(X�	�
�g&L��%R�y��'�R�'~2�'	�����:S�M��K��"�S��0����?y!�i�D��O�2ik�Z�O���C ). �y���)������j��'E��Ao����:2I�6�h�h�ɖy�xT3/B)�V��&c��5�,��Pk9q��i\��yy�O��'�Oی7[�`P�n�)���p���7a���'��	�M�K����O��'O��鰦͢���!I�$rF��'&��dw��Ab�6�y�'o���J���HJ�y4��/��x���;*��i>��'|:�%�N�8A!xY�u�ՓP�� ��Jȟ��	���	�b>��'#�7@�$����ai n��Y�%W�@E@���J�O���ئ��?�"V��m�N\�À�O��Y0%��p��Y�ܴ�?-�ܱ��4���I�~�X(�����A䅘g�ֱ8�L��&L�Hy"�'���'b�'r]>��c��dP!@TH\	
��pH�,#�M[�B*���OH��H��ڦ�z��`��L:}���� IS�	�ߴoț�>O��S�'5��-P޴�yrH�k�>=qPY�_�Q�"c��y�Ӡ���	?(3�'��i>����@�L�XKD� Z���F�C ����ǟ@�	џ$�'>d6F�3��ʓ�?y�$/�H鑧���q��a�A���'����&�{���	Z}
� �����L'P�3���c´����ҧ��l9�j��.�n32�N� �!P�R�!G�K0������|�I؟L����E�t�'s&M!V�]���d22���3J褪��'I�7M�tGB�d�O�HnZQ�Ӽ&�V�`d,y� ��	�^5�$ ��<	�i�6��O|(���a�����0U@�<U�bLԥA�l�e�ݍ_Wb7l�?gU�'��i>��I��t��ӟ��I�`�0����ۮ�@� �wZhy�'&D6�
<8���?	H~��y��Ms�b_m龝���M`+0���X��cߴZ��f<O#}b�JS��J����"6:��hЊ�q����Qr~R������I�d\�'��	40�h���̑F�"��΁�j��������	ן��i>�'|�6�C-~����ۤm�!�4�\+l����-�����^⦵�?�X��8ߴ@ꛆ�'�h�ӕ�͕��H%0dzԐ��ʰ]��F���Q��C�Y�����U2LƲ���d�-�P��$�:|�tې���QR��y�P5&g���M���y�df�1� �2'�.T�ԛ���}
ͨ�XJ����d��"Ӝ�;Dҋ'����'_:r�sN�2W|n%`1�ޕP��	eB�4��7M��/� ��H�|)����]4�Mr�	Nd��Q�O�Vf|y`�+9��4@�O��� �ŐI��2#E"<ت��+J�#Gȕ�<"j���k��t(��K3d�4�ib!���x�V�%V7�d��ː�(
:9��o̼Yh�4`�!t�nD��]�Х�a(��D�O���D?^?���>)��~R����CjIE�=)pm*��' ���y��'*��'-tD��<5 �*sA��8�qr$���)xd��%����'�8"1��/���`��&��R� P<����;{�1O��D�O��D�<HS� �$�ɗ�͗=�Pa��NP�ޡHE�x��'���|�U�X���D�$��	0f�:F�Ru�*c����џd�	byb�C�J����js�ȡ�%��D}Q4g��W�듭?Q�����Ԍ~��I.k�z��7Á)\�� 3�'�H듌?����?�/OFE��kEb��^ L��D��o��I��J:*j��ܴ�?9N>I-Ofu��IW�j��2�癕��1��c�K)�v�'j�S�����I��ħ�?���a�ZQ���R�S<D���#�C�gy�@�����Ӻ
^�pib��wx)Ctkͷq.6�<a6�W�	h���~��ڷ���c#R�eW`Y!����P�}�b�9o����i4��i4�A����z�~�"�)QIdX�ߴm���f�i�B�'���O:�O�i	�hر'�Ïq[���A��:||o�0V���&�9O(�d��)C��ą^���d��I&r��nZɟ��	۟�:�����|R���~��ڬ𲠮T�P��Td1����<�r#_Q��?��?�" Ɛj�,����[��Pr�	5�v�'�@I�!�4����+��Z6`wD�� WB��Ҕ`ې}����'���p�y��'���'�剌VA�A��	w���uo�
��SF���?1���䓔���%�L��Ӥ_����F��4VZ�Z����O����O<�Z;8\)6;�<��ߓ4`	�a3�)�5Z������$���'�j��O�y�@�)��J& ^�1����Y���I�����dy"��$A!�(��� �T]����FL�L�����`�y��D���O��X�63�iQ��� �4�?����З3�X�'>��I�?�X����f�*7��}*Fa�^��OF�"�1D�̱۟��I�L�ҫ�m`z���]�L��V����I�,�I�|��{yZw��q	Eˏ6	���p�A	�g��O��$��)>�D������a&/�`lł!cK�th�6!��5�2�'9��'k��_����(@� 3���ώ3$�P� À�M{`�D�'�$�<E���'�l����!8�xA��JDn܊�i����O���]�}�z��|*���?i�'�be Qa���꒶0/��U�/�I��=�J|����?��'����I�Z��`b�p=i�O�mr�g�<1��?�����'���.D3?�Z�����u��eI�O@�
u�ۂ8��I���Ipy��'���d��F)͂�H�4U���Iq]�I�X�	��4�?���F��F��^x\4!�+ˠ2�\M��'��=�'J��'�Iٟ�y$N�V�4eFd�x�)��)���
��������	{��?YlF�_?ذn�6�����ŀv����L�.8%���?�����D�O��x®�|b��Cz�hYB�
�,�cC���ԁ�4�i*�d�OԁJ�hҢ[=�'�DC6K��=u)�@�A�(�`�4�?�+O��Ą�"L�˧�?���
���{��kc�87t@�Q�&��O�ӈ%� ���T?�Jbg��l:�0z�eZ=H��(��>��_�rEB��?���?������MQ�k޸-n,�El��^]�A`�_�h�I?�	e�=�)��\���N"���;3��X��7MW�'\r�D�O�D�O$�	�<�'�?�3Mgz<��O+`�6}�r�W3)3�CH�	���y����O��1�c-�6����;Ffx���Q�5��䟘�	�u>d�����'���Oz�r�m%9�:�X�J�����H�V��+��\�����s?���Ưl��Z����q�����i#|��IH�Б�'Er�'tB�Dݔ
)���Q�{����mǭ�����( s#9?���?)O���A�? X�6�Ҋ/�⸸a%&����W
�����O����O��t�i	��G�K�g��u�Qj�0]�FEn�,>��?y����O����L�?]�3C�#�0��M-c�V��w#r�t���OR��9�	jy����M{���( :��&��[B��ReHd}�'��T�p�	��<�OK�i�=C�M!a°W�jЧ-�71P7��O⟴�'9��+H<��@�	��e!��[�wV	 �������Iry��'��ey0_>Y�I����8'���h��v�3Ec��t��Ɏ}��'��y��ʘ����0�͘F���Q�n�;v���џ�����ҟ`��ɟ���?i��u�KS �T��j�*%@.ܪmS�����OX�[A�
d1O����)���,a4N�C&�V��6�ir���'���'���O��i>M��?HT�q�ɔ,����ɉa�hܴn��9aeJ�a�S�O5"ŉ-N�h�։@	"��c��	M��6�O(��O|qY�i�<ͧ�?����~�C�e=xd���G�:Ζ���kW�"�c���b���'�?Y��~�̀*���:��)	1��A'��M+�o��-O�D�O~��4�	C�*}(�/�<%rH\;f̓�V���nmN�i�N~��'��[���I;B�;�K�P��,����4[XD�-�uy"�'�b�'��ON��F,gf�hR�,����u�5a(��Hr�V�J1������`y��'��(JAן���vņ�hZPQ ���MͤM��i�2�'�����O�Ɋ�M��Л���D���H�Ɣ�$���p�C�����O��Ķ<��e�N�z*�(�O"3T�G��/�N(�`��L���l�ҟ��?Q�����V+]z�	6OF� $���eT��J	/46��O���?IF�ҧ���OT�$� �8G�ԽG`�u
�#�"�`��)�M쓫?���-�|�<�O��$s���xM[&HZ%��>1���Mc��?���?������ƨy�뇐<Y��LԹT�Hh�@[���	�l48Y)��<�)�S�D���(� �-�|���.0.7�6>��D�O��d�Ol�I�<ͧ�?���
�Mx���׏À^��\��H�~���ݗ��y��i�OZ��ahLc�T���d W�4p3��Ŧ���hy2��)��i>	��П��A��;�C?C�"�QŌO�TM|�����:�I$>��	֟��4�@�E�Wr7�%9#��<swl�oZޟc��|y��'B�'�qO�X�%��	jI��{rK-Oծ H�T��+�,$u���?A����O�;p�Q�t�P���6��\ِ�ڳ%��˓�?y���?�B�'�h�;�h�&�49k@�Łk�Xq#�W�iw腚�O��Ovʓ�?��������ܫ:�4���Df�z
0�M3���?Y���'*��X�?����4Y���nвG���NR"&l��'�b�'��Пl�V�HU���'K�ptf[� vjt���M5{i�<qHr���,�����p��L�I*O��GY��rlp�c�-a�!��i��T�l�IW�l�O��I�?)�cJ��]�Iz�xFk��uG��s�}��'� ���,�.����)�l��U�TMš#��Α0$D�����^ԟ`�I��P�	�?��u燊�`���*��:�4�
����D�O��ېE�+�1O����ǂ�y�<�� ��>Ϊ%T�i�z@+G�'�B�'���O��i>�I7/�,����W[P 1'ω�N����4b��9���u�S�O�!�Y�%��jY-���T�ʫv��7��OL���O����<�'�?���~B)@
J���w Z�`��GÎ�jk�c�l�#I��'�?I���~bJ�W8�Ap�	��2)��ȍ�M��o&V<i)O|�$�O~��'�	�y�ta��$�'V� �W#Ԉ_�d�K����2��C~��'��P����:��8t��8 � �+W#;]4����gyr�'A��'��O4�D�U�TEX�m/	ν:����B\q��;:%�	�$�	Cyb�'u�e� ҟ�x$Y�&����� w�᧷i&��'x��$�O�33f@!Cڛ�ִ6���L\$/�Pt���I����Ot���O��r�.���U?��������`�����K�c�J�z �4�?�(Ot�$�O��Ҳ%�O����A�$:���	PjN�p��i_��'��ɳ`	�uڨ�r�$�O����t&$��D�ݍ4!.�O�1'AI�'�b�'�¡��y�^>�	c�᫊�wf(RgM7�� +Dc�ئQ�'��D)thx����Od�D�� קu�E�tb�ʥ�g�L�bEI&�M[���?�GC��<��U?��|�'O�<��&�ՔK7(�b�U�d�oڿ+����ڴ�?9���?9�'LS��kyb�_#o�I;FK�>g4d�rG�E�p��6ML:7��D����{�N��mB	[�쉵hX� �P�it��'�"�H2�z���d�O���.�$eǏJ!���TiS:�^6M�O�˓M�j��S�d�'�"�'�$���J��F�x*�Ì�?r=��bi�^���cd���'"���H�'#ZcbƼp�n҃ r�0�E��]�`8k�O�����0��ş����x�'����䡊�`f��Yf��j����N����d�O�˓�?���?� h�i��B�L*&�F���G�.�u�'MR�'u��'i�	!f(Ւ�O���kaĕ"���em�14 ���4��D�O�˓�?����?�ӥ	�<��b��s^�P@ھ8�a�W��	���ݟ\�	���'�Z-җ�~Z�s� ��Sb��!����g�*c,"�
B�i�U��	П��	�p���p���:eQ�I��cr��"�����'b\�Ļ�툽����O��$���%@�JJVd���S�"x8�Û{}��'���'Ҥ��'(�'������9��ZK�.�)B�6ϛfS��i���MK��?1����CQ���.=4P���}�r�����j7��O���G$#���Zm��'�q���tȘ����W�b���8b��MS$R�]7���'+��'2�4��>)O���Q,��M2TDK
������� z�7O�ʓ�?����'�8�Ek�$��� �E�\�r���y�����O���K~7�,�'��	ϟ������W��[�
,E&Rq�dl����'_��������O��D�O�Ѳ�K9lШ���'K�:�S7�W��u�	� �܁��Oj˓�?�/Oh����@k�����a�� �|���\�����d���'���'_�_�T	�����\�u$�)�����m/H�X8�O\˓�?�.O^���O����bf�ǍY#u���H�G?g�6(�s7O�˓�?����?Q.O�Q�Dn^�|ځ␓(n�����c�K�ަ=�'�r]�8��퟼��?w;R�	#'���tB�r�j3��֊;h쳫O����O�D�<9�$���������ʎ(��2bf٪v]����M������O:�d�O2$���?}���4� Fύ22^Qx�$V.q���m�ݟH��ky"���p��'�?���
Ҩ±�h`���[#*A`AU�k�	���I(�`x�Ȗ�y"ӟ�m��g�9p���Q�$�һi;�I�&�"�kش�?����?	�� �i݉("o��A�9�śs����h�����O^X:O��$�<Ɋ����"!��MD"T��xY�,ۃ�M3p��"{���'U��'v���>�*O. ��_�zװ��FH"V2��3%�O��`㞟l�'����DZ|L!R�ŝ)\�ȕ����
 lZ៘�I��|AW�S���Ľ<���~�� �`Ѻ�ぺJ�kUN��M����?���!>���S�4�'l"�'z�DaVmX.# ��ag^�\r�Ȋt�eӨ�d�:3��'����t�'�Zcs���>�<}��f�$E�-y�O¨p�=O���?���?�+O~� �灆�x�D���Z���w���n}�e�'�	埐�'�'�2.8R��)�$ٛ)�p�Y�;,d(�'J�Iʟt��ܟ,�'����Ca>����IN��7gIۚtR��z����?A.O����O&��ԋ�do��0��D����@S�5���n�ܟh��ϟL��Vy�]X��ꧨ?��6G��!��tv�l���R	�mZɟx�'���'$��E���Y�Գ�mޠu��!"cnӶx�Ӈs�*���O��N4Xݺ_?��	����ӳy��8C7�M�M!���c��M�|˯O���O��Dӻd��|����
�-�v�ڠ��?W&�J���
�M�-O<��H�ʦ��������?�K�O�.O�����1Hx�� ��/ ���'PR�['�yr�~z����O't0�b�,z��a��wB4)޴v�>��p�i���'LR�O������d!�����a=F��r��0M�<mZ;����<��ٟ����rH���c�W 'o~��F�0Qyp$R��io��'�"�H�D�pb�L��h?Q �Q�#��1Q�.�l����tn�Ǧ)&�d��{��'�?����?iԪ�wm&ܙ�c
��P�1�׹*(���'c��2.4�����'�֘�~r��ףQ=�$�l�|�U�D��<���?I����D�>[B85��H�A��TQr&X#Ot^8{"��c�	�8�I]�I�<�	<m}��4#�<���"!E�?���îJϟ0�'��'�T��2�1�����:6�(�`b_7z,���G����?�K>Y���?�&�E�<�PG=t�� �w�Z�%�4���]	X����D�IΟL�'���6�"�9��J�GM�4x굫��~Em��'���'�E�6�y�>�Ƀ0��9P`$!����ZӦ1�I����'%�d�d/8�)�Oj�Ɂ��
�$@�|����~B�m%�L�	ϟTC%�:��T/J�3t0Y���J�}��sT���M�)O���K�y��������L9�'=I§�5=�+�O�,G�U
�4�?i�c����R�iY�/nn�SU&B�+|��t��-<O��	��r]�6���f�'y��O��b�`q��� 4����� ��D-~�q��>�MS���<L>����'��4����Y�@8z-��{��A��{���O����
�t�>i��~2���5��2��/uPQ�$
���'�4��'+�	���	Tj��h��C��z���[!F����I�Ibȩ�}��'cɧ5�b�?lJ�xQc�90ݒ�1w���'��aS�'a�I��x�	럀�'?�H��� f4ʬ`�L�}k֩�ǞQ��b���	t�ڟ����h\(0c�-Hܮ�S� �f(��2��9�$�O6�D�OB�@�!pf2��#
�,N�-c��>6a`u��_�p�I��%�t�	��I4�t��Ue�;q�H�Kb�8����w�����OL�d�OR�W6Py�4���N�9z��E�E��m�8i����7�4��?)d
ΐ�?	���~�(L�$���QR�O)i*(���4�Ms���?A���?9
��?����?���ʒ��,Uj` ����@��(�Q��'B�'��h��?u�"À�BN�5�5N�?!?j��G�s�f���O���5��Oj���O��D����� �(0�M�xPl�W�8���W�ig�'9P53��K ߘ��O8�h�s.�w���ԯ�.ӀD��4_6��Pľi;��']b�OB����Ʉ�^/�8�ɝ�W���5��	EN0�l�CBf��?	�����?��H�8wS]���	p�����B���'��'�:�t�'��_>���a?�A\r캈��憕��mq# @
�1Otu�q�u�ϟ`��񟌋Ê2�9�T���8�B, ̓�M[�����?Q@S?}�	r�I29h�9�*7E���$HD�a�v��O�H��a�>���П���ʟ �'������Q�4L�2E�Kc�-�T
�X�`��؟h�����?���m�P�qŀ[1w2B̢��Du&��N>���?�Ŧ�����{n�bRV��*B�T׭uW�00�Q֦��I�d��_�	�`�	be��1UCg�����B�r��)FU�0�	ğ(�'�r`B/SA��'����) �Q3-<���ܶM�7��O��O,���O<�q�FZA��'��A�A�7�nQS���|FV��4�?�������q�p$>����?�&O7{ �:0�� ���+�_)���?����Dx��bBF�)c��Eb�#���[ƹi��ɫd�.�{�4D����|�S���[v�p+Zw�h��E��3����'������O��>գU�ӡr6^0��"�h.Ԍ� nx����S�˦���˟��	�?�yI<	��4�JQ����1`K��⧫ٯM2 I�i�э��#�����`��kO�uZ�+k�$�����M+��?y�m$j��+O8˧�?q�'�`�6υxx��r��j~f{�}­T��'���9���x$�V:;�F�!2�֤�J�1D���lF�tr�q(Z�YdH�`@m.\On�&�V>t˳
�~@�h�,��w A�֭�4�0�$�҆\�
X���)r�"��`��EF(.��c(�!CT��"0�౹��ߜh� �a��E�j��2�!ՙ"�42��,�&TH7�H&i.
-I�k{�P-!b�@�~��ĐV���NX�#����#�Ţ9Q���"&_�:�@8K1�'�JՒ,j��'��	�:
Ȓ�Yp@��:킈�,�<�hh�T��!^�Ex��,�J� �im�'�l���(F?7�X`iE�I{<hݫK,6��Y!PI�c�l�%��+�0E{��1�L��|b���'�^1��.Z-)�|��w��&���'���f���@y��FEQY�'E�6m�2x�J�բD�fδ�pVc<PP�<�0C�sp�Iៀ�O��t�2�'�Ht1T ڣr�����+_��pӖ�'eKR�TY��D)�Kؔ�0���O��~��hɘr`0�A4�ɲ]1�1%���	Rϰ�za��)<ܕP���OY2q��E.�*Yド[�6��)K�H����O��d-ڧ�?��e�,h�2TQ��LH�!���W�<�����/��@ia�)MDpi�Lm��Z��$ߖ-
��B		F����(~����~���|S�d��J������x�i�)�!��Hz���bj�+^�@mA�	c>"��g!U�?a����'��,�|&�� �G]Ȑi�չZ�~Qjs/Ic!� �槁�?)�iY?���>�O���ES
@�4����0p�v����OP�b�4m�i>eF{R�Ǐ]�q�p�l^�(+�l�y��C.M��G�/���+�C���Py���)�<y�`ߌS��0�`��z���U�
�t��#�?���?)�Q��O��$e>	��dP�@1�M��	�ǖ-���ĉi/�9{�S�к%��[x�xT�M0K/����J�0C#�u�dԏ?| ۤ�?�>�R�d��(�E��+|Q���� ܡ�6��D��F1Ty�.=\���$�O>�=�����d��p잓�n�ʖ���y�bE�J�"t��F�V�R刦�)�'|����d��(��X�'hrL�s�0I�3R�� I�d
�E7��'� � u�'_r5����Q��B��!����8�4jE�����r^4eZ�*jJ��	�1Š��T�L<b�I�N��|5ܡ��cI�"�Ǉ1<�j@c#�22���r2�@�����OʓJ
Hܺ3�O8+S� ��OPV
���<�ߓ�ti�aK��N�"���h���oZ�FI�
Q@ʐ����Q�JbƋY/�y�U��C��].����OF�'RZ��#�[6M����8�"�S����!3��?	�Ϗ�1�ܑ���X�ci��S��Q>��fL�0,���TF0�C9}�ȑ�X�P��B�X!f�N�~�e�EW.X{��2/ڴ�I@�j��ey��'��>��	�i��pa��1Ӑ�ఊ�E�0C��?_X�РE�͘4������)18^��d�R�'j���f�D3Nr�UХ��9{�O����ү*�z�k2h�8�^�Rr��
z!��I(��AAI��ѩT��`�!��8j�X�D��<���A�@�!�D�o:�$��Ɨaez��@E�$�!�Y7��ə��ӡhK����9�!�� ���0�<R*�+M�![��ː"OB5�r�Bj^�*��H4585ȁ"O� ��dӕ6c*P��#�>4��"O$ؘ�`]�%�� ��;5XXu��"Oԍ��e�Q�XT�F��=L�aB"O��!�������;#X$�T"Oޙ��H�1ھ\���~m� "O,��$��+*d�.��y�a"OѨ���T5�2�D
U�N�j"O�X�$�9d�@Q� ���s"O�T��-�2\�h��FY�9ʅ�"O��q���U�n�� �-y��1�"O�Pa,߿Q��Ȕ�A�k�BaKQ"O���m@,
N�	x셔 ��t��"O���c<NQp6ҷ�u�w"O�y�"o�q۬5Q����N�2�"O ��dj��F��ʶnT�{	f=ZQ"OČ�`�;�B���K7>����"O@����H� �P�sM��y���"ON`8�/]�0"���,hk�Q�"O��q�R?B[ʰ���(��|�"O��P�Ϝ6_2���&���`�)�"OX��%��2>q1����O�9�"O���&Ϙ�萉�
�x�"O^�rA
�h�������P���"O<a��m��S�囐�ֻc^\-�R"OVY��ѠH����`�C�֌	q"O�$�C.�*�:=)b�3��"O���`��R�DiǎV�H�<�""Of9X���">^;��2w.����k�8Z���b�^9��2R���4��k������Sn��7o�Lk0"O���g@B�oMdԘ5�K�1
B�HE�X�;Ƥu��H^�9���,\�4��c�s���ce�%�t/M
h��9�7D�Ȱ�"	�UCB��:5��3���<ko�)o�
(�W�޳0�2��'��PDxªM�c�= �%G'($
U8�C�0>!U�ҹ,ײY!Ӫ@<p+���a�3;�MR�gT�U�Ќ�T��QN�y0�'x���	Π
�b0���7B�h���-�s�
�%�:�#�A�k��re	�GP�\ҥc4J���y"/XW�V�i�"O a��7���U�b���;� J�P��d �4���i�g��W�A�`�5	�1���>J|g��{0 �7�
|�!��V�@��9+�-GtE�fg�(z��HD�����tHN4�V��;��8)�	-I�1OT `�k�fg�@0��݉1�A�&�'nN�z3�M���A�:[� B�� ��!A�.��`6�
 P8�A� �0=�S�Ј|��I`る�>80��C{�'FZxj��Ƒq9��:���5w��]0ଔ�rr�=Z��ۻc X`��kّ���IcL���y��¹N��!�?���{sM�]h,��B%��{º��e��WtИ�ûJ�(����w~�K7★(���ŋɰ22�A�'�4Q��J�A#"�i�_�M�t�E�]$T�Y�.[�Rp��2@����B�㢥j�y2�&*�l� bT���3rA�0>��叱k��a�fO�aƎB�Z!<�CEb׉אi����8���B?P,f���ɏ>�tKS��:2����@"#<I���_�4�3����*N~�a�N��$�^�_0��#b%Iu̓[8��c���)_�=��vI�<H�`�ߏk��D�'��Wd���L<&1���s����O�5Qv�c���'t���Ƭ����'��+���2c��S$Q
TBۋy�����lWߟ|2�I� ������-/��F���,�8��J�:&����Oם:����!�*,OLQyae��{�d�ѣ>ti1 �3^Q�6M!eU���k1��<�he9��x��	~���l�̌� K��Oda+5�c���W�9YX`���@BEH^!����6���������>�|��ʑq��!����=�=�UkVA��� 	��n��/O?�I��!Cp)ɒp0���U�zGJ�k�}�ߓ���I�P�0DP��L�~�*�� ^S�I$:ʅ��?�
���!���N�e$(8K�㙒X~��Q���.��<q���e1�5{�OV���q$A�*x��oX >��� 4ثO<� t�:㌒+Lj����>s5�!1!�	2S�t�8焂K�O�8p��"��Ds������y򠑭��b�b>�Dˁ�,��G
�_;N����'D���'�Н]ͶPr��\�d<���-��'G��1�𙟸�������rE��6+N`j�4D��KE��`in�P�� �8'.P8�钽P\X<A���XW�Ҟf��t:�B��&t���I�{T*=(I<��J��M�5J�&C���IBY�<9�F�|�x�� �bI��a�X�<a��P�U��	��(, ����P�<��8i�$)���ѻfh�dB�	�	K��С��6�*��d�VB�	��&@2��=|�	�2��f^<B䉯��i��H
R���'ғ,���D��@�t�q*Gb�.q��f!�"O����R�&Ɠ�Es��3�"O�xx����oژi#��X9G~$� "Oz�E�#<��}·�r�]B$"O`x� �0/u�y �$Օ:@"�8�"O����:{����bQ,�*���"O�!����#@(�AŁ�Vg�YKg"O��f�Y/M���A.��hM`��"O��P�1+��=�D�Kۜ�(�"O���ȘV�1���o��	�"O ����ϙs�V�c'�ԕ"�*h�%���
GN�k��|�\�^K��ӄԨ���q��(�O����Od<�qK�?nh:��#o��"OLM����7�Z��U��{�N����9�!F���=~C�Ũ�S�f���ƕ��0=��^�^�#cJG�<Qw�ο@��肤�/���c��<��DK������,S��^�9�h�A�gߒZ�n�H�dސ^�~��K�01�?防W��"�x��@.�����)6?Qq,����=$���~���yu����R�q
�?E������__~r�����	 8���Ӳ$�y�b�@1݅=C�ɐQ��q���|I4! �#R�-Y�A�c���D"�O��H�[w<z����
!�`t�W�'�F��
��e8���'l���(�u�\�;�j�X����'�=l���S���Ӈ�3 �蒌y�1$��҄oہ���:�B�H�.L&��ROIe<x�0"O�Q� ]5,�N�?r3N�t����S������1�g~�"Fa�4��ˇ$r��P�@C��y	�O����#N�WS�H��x(˄˥s�nm��'�i�`
��O�@S2`�`�#x��:2�!LO d����;^F=�U0Oxy�6��,	�b�"�.�<U�\B"O�}�U�==��� �@�16D��A�5>T�B��ٕX]?�k���0Z�ۆ�"�"R��?D���S�P���\ 1��>tx�<��^8M��`n-?9�-����F��ڽ��f�;N��s���W�zdۑ�܉k`a~bjťy�tā�L��!��p�F|�GOF<äЁ��4�<�{��0c����}k3+�� k@l��?D�0FB�=3�!E� $��a��>�	  ��!u�?�"8 +�ZP��(�v��0"Oxl�#'�YQz���:��|��Ƥ>z1O�\[�3?�QkЦW�z���F g�=q���K�<� F�L�� ѵ@7&���Y��p��(
P��|3&_*p���KB�d=X�J�	"LO�C���$��-���acX)J�f��� �&B�I�R�V�)���w�>E�mF:���?�Bڎp���<�}���1@x9�g�J�� RN>D�K�Z&ad����3 ��4�����@��c��p�'�g~Rᙍ�H3f�# **8a��yRb�_�L�	c�4&�ᡇ�v-��5���0?1���t^B	���@�zۀ�k��~��H1� G�i�������fΛm�0����C60=���S�? n@s�B��k48���^�sX�*�"O��G��
�X�cT���5�
�q�"OP�j�?�V=����=r��"O��Pk\�2� �YD�[*_NU�B�q����'\��ꂅ1�3�R#>�@�W��i��"PǞ-�!��*FD�D
3P��M3��S���"��K�4�[P�'� �2!�/WŠ4��^�A	�Z��a)+>�>t�'��`�+ �i��iu#
J9<�I�'��0�$+דm"��d�^�2tЊL<9S�U�@m(���iU�O�0QB-ʅ������VL(h�'vr��3 ��u���B�-
',�L���'V>��JPĹ0���xS[��# �V�pJ� �.G��x��W0��0�'i��c~��`F@�Y��$���!}��z�2m�U�G��>{��u�P"��I�y�����$<
�"�*�5H\1n,rl#GF�m��ȓ��(+3f��y;��I�oѻn7��%�XS�ޠs�~<K�#2�$E�YPs_�b�jeف���`Ԓ��ȓ7:
`�CC�x������^��ą�0���Y�H��=�L8�Ǘ/�d��ȓF3�8
��g���J#ْX���ȓ���઀�f�@�Ā��W�Ƙ�ȓ?+�<Q2,ܡMv�M�5�� |>��ȓ=�&q 򨉺݀%㣋޻�4ɇȓbπ1���]ސ�҃�H�Pćȓ	� ��M�4w���k'�9B^��ȓ>��L�e��fB�6`dq�5�ȓ�(�:UAֲ.���2�<V��ȓi�Q����~�p����r� �ȓ5%��� �Q�4[& �2�J���>����Ci��VM���AO_���X�ȓQ}.D��G�c\�2#��Bx���ȓX/��/5C�$���UO�dh�ģ&D�����Ɔ6W�<�dB��$��2�)D��т�_)d��7�6)el{��&D�����)&��٢B)<,8"U�%D���"�X,)�((���-)���#�"D���#k���1;�@H�x�l1�f D�L)��.}��j�E
&l$UHԫ=D�Ce!#.Z�#���ɑ�I:D���GK�f� ��S�]�4l��	�,D�(��i��[e$a��o`��`�5,+D�TA�J_R���"�\�6����b)D��*V��i�d`I��Y���D�܆�yR]� ~�ӀK�Q�^D�F���y2����8���^�Q�ڕ�B��y�5'F4�(��=����D�
�yb��%(��Q*P�/�>�qCL��y2-�3�Z�����'�B��%�_��yrj�9Q��0G*ϼÄ�j�㏋�y��
f�Ҩbp�ջsHL򃏘��y�(�(y+րp�e-*�h�
� �y"E 8�Tb�ռo��m�
�
�yrAJ�+vX����a-
1�E��y��#�����d�Wd��ť�y��*(�8:6C
9E�h�$��y���\-���ԈX�'����@W��yR��� N�����\����z/ �yB��B��<��cJ'M@��q�
��y���Y�����>U��t��;�ybj��N��q���ĔG�"x(`& ��yb��0��pk�A8>H�y���&�y��-H� 9Q�n�C�q eC��y�=A�������j�X� ��ybD �mJd�H��Y�W���a@D*�y
� ���Ѥʀ
�q3E�	{�{�"O^��N�?vGt�Sa'4}D\�W"ObUyV�@�RKv��Vȑ�
$�)2"OLr�'�9��̋���z���0&"Od��O�jf�BO�+lJ�"O�Qbd�������.b�2%"OΨ�WNO>*'�,T�9v�����"O��3��D8� ��$.	q0�B�"Ol��ǀ43�e�4c0H �"O��B�^2d�U��\�f�~�X4"O8�
�G��Z���T�U�T`8q"O�`�Ѫ�V����e+B�{eйY�"O� ��d��)Ĝ��3醍W+�5�U"O�P� �[�xI�d�˧,*��ذ"O�1(�d�B T�x#�Q�R!�YF"OK���Wy ܣg�)336(Ҧ"Ou�bi��:�D�M.���"O\�t&�X{�� ��5+^��Q"O��	B, J���,g,8�'"O*�`�eG�J��}�d�,�d�C�"O��s�iR#,`X�ZF�Is����'"O�來�TOB��
I�Ѭ��g!�],v���������̍Q�!�@1>qM��I�[����FjO�q0!�M?;���{�O<q�T�	��!�M�X H��ԉ�0f�ƀ!6��*�!��ݚv�@�p���%�zAaԦ��<�!�dĄ�����Jw-�� ��éx!���2�:et��&H�ԡD��1�!��X2��o^)L�,hH��2!�J� �x�Z�5Ѐ)iG�1'!�DB�}�H�� Ƈ4�pU{͛
!�D�ch�k� Y�S��{0�/�!�Ā�	g$���g�.��-��Q#!�$)=R,aP�-̀P������!���1���r���l�HiQ���!�$��R��%y�ʍ,-���*Gk�>$�!�dA;�2�QS���l9У�M�z�!�d�	��Q�c�8݈�P'�Q��!򄐌6���'eT5'2t��혜^�!�$Z�/��9�G��ZsReӑm֑F0!�B��\���蚦)Z�d��ŕ&3!�d��%���)a !��U��Ŏ2J!�d�A�<YK��-�f�fG��T�!�	 ^�0#B[��9"5$�/|X!�䙊B�f1��j��]}%�fA�I!�F. �@0cT v�у�A�[/!��N�r�A b�i�8��l݆-!�d�(xu�׮Ov���-X�!�J�?��]*��\�r�gT!Ux!�$Բ|���`�=w�<,(�e�*�!���Tꆍ�TC��n��� e=\!򤘿G�ŋ��_�VK�x� o��O!�_6���ꄊ��U:���c.F�
�!򄏫"1�B!�/r�<=��,��4X!� H�P��Ah�pn���K�&nW!�D�@ 怪�wXhZFT]k!��	K��1Qwaȫp�� B�67N!���Msp�S6U�����*~�!�ĉ�H_��`c��%�N%�R��=4�!���Tl�y`�B�}�.a��}!��#�@�����x��lh���B`!��S:QWba�����McU�=hK!�"`��[��7X�HA�W��'>!�� ܭ1��Z#AV@@
�9C$��g"O.x��̓/;A�
�HA>y,,p�"O���� jI���ӜV]��"O�D��cS'8d4����ݻ53��D"O(!�O�7-�C�C'y+\�ْ"O*��
XM��M���X8p�#�"O�}�%�FLiv �w�;���"OV%�B��	QA+#���{&mP"Ov ��ִp p�M6'�会7"O��sff�jP�����1c��"O����P�>w����-��Jh�!�"OF���֦+߬��7��1 9ry8�"OZ���I�t�.Ua�,ʵs�4��0"O����䛍G0\����/@.F�#�"O�Ɋ��X.Tb�}��e�X�x� F"OX��Ċ�t|n�Q��%)ϮY7�'Oў ��h��eF�CQ�N;\Lv�h�J4D���K��<�H!B�R��DI[G	1D��*0 +{Ԇ�{�%Oi��y�@*D�<Qk;(�<��%�5����B/-��p<y iKv4M���K!y�80�&\W�<YF�=��pA�	�c>X@�V��H�<�q��j��C٣����+[`�<Y�������!֣O���G/u�<�U�R���+	�qC��¤�Rw�<A�Ί+
�$%��̄�8qZ��t�<��[�����zn>�+��u�<��F!%�Ҍ�w�M�D`����y�<97c�$�2�ja�;Ev��CI�|�<�b�G�rM �� b.�ⵘe��z�<Q��1^>V����Z�VC`�8�Ɣ]�<a�k�U��y�>=D�S��	B�'7ў�'Wʖ���%8��ˡ
�<o|���ȓC�>�S��X.4l񄅻T~Э��;���y�I�<��ā�.iŅ�Ic�%5�(�%G�-{��3�I�(3��E��R�1��޸�l��b�I�L>���ȓ0V��ړNH�e�����W0>	��-�0��ΎQjK�lZ�/	(��'������" Q�x{�͂��\��L����LQ� ��m���5:�X��ȓ�&m�nSQ:N���AB�i���ȓa@ب ���}�V�1�U5.��A��($0�C��ͤ_�Da���d$���j�r�82��|�4tp&ӣb����8"Ds���u�)�(������&��8A+�.q�b���͚N�lM�ȓi|�y��^���"`і:"��ȓ����KJ'_j��p����5���u�������'tЄ�M����$�ڸ	�^1-��5@�g�1����q�����M��W/�)o�q��z��"E�T.]��G�(�
�ȓq*�eH͏7xD�s�� ^Q��ȓ[�8Mi"�3){��SV�;C<���+�����8tr�	�clO˂#�[��hO1��Q��o4pur��ŤN��� �"OT�A���l6*���h�,��a"O6M3�kޢ]�*� 1G��X\�"O$�p�(k�"�¤�8���!p"OB�T�ح�క�+�P�	R"O�(�#n�1;�T��Jݛ>�6���"Ob�i"m�8��s�E�p"O��#S7\� �L!�6I)�"O� 8Y�6�Űh�֌r�%W)4�¶"O�e�"U&������^1;�$��"O�0"�,���x��M� b�P�S$"O&yBU'�/eP�8�˛�M}<5s�"Oti�̐	vs�\�d��/�x��"O�%s�Z?u�&�qedˁ5��Q�"O�b�^�MÏ�X���"Oz�t�LG�@e ��]�(+��2@"O*QK�h�_���;� Ӽ)&�q"OR���7 �]�ab�1dh\�"O@� N��.����M�,8�"On��B�37\���#�<{����"O��
Um]�j���!�����Br"O�h�l���6K�T;�!��"On�K��^ 9��� 4��/���0"OzW��5!3j�	���1#\�3"O&͚ �P=$�%i�mL�Hڭy�"O��0D��- ����	��ȁ"OFĹ���rK�LP@K��f�u "O��xPK�+X�F�T�C10�5�"O ԫ�>lԩA�̎Kv	
�"O��ȁٓ&�j0�b��
#; =��"O�}��%�)���)��O� x�@�"O��%�W�D����$��(�	���'o����� �Q�|8�A�!��U(�B�I$O�B	�B�z���HwFɢlJ�B�ɸd<i �f��C���jQM�1�B�	�D��m�,�p�{�%��?TlB�	�UT���Fe	%+��A��[&�6B�I�RSh�{ׁ�5P���S兜�6Q:B�	1V���gЕ2x"�!Y�j��B�	<)m��%I�6vp<�3d�+Z4�B�ɬ?�j�KC� �ib�15nC�	>Ұh�e#/5�t���>4~LC�	h�NňF�>���K��+�DC�	7L���f H�Kc�HȄ-�;pC�	�	�|�*�6E�|@�a�p�B�1]|h)w�B�*��!
�5BʰB�ɪYg� �7�pm����S����`��<����fur�E�?\ub��ȓ1z�}�Vl
=	# ��!L8h&�-�ȓ`��-�C��	%��L�t�M)5�Q�ȓd ����Y�b�j
02�Y�ȓf��Չ3n��fB����	��e�0��ȓz����)H.* ΍!S�W�i�����رj�#��>���Q5CT�ȓh1"	h�I�b' �&�ڳ%N�U�ȓfn�p!�H�r���(Wb �cL����D{��Œ!�]iD2/-�-����He	BN���Q'�ij���ȓXiN���T/z�ltS�φ�R�~��ȓE~x �K�B<x�� �W>n͸����|�Gׁ9M��j��C�`Lh�ȓO��ŲGL�*p�r�J�b Q�	������'�Ę>$��RB��G`P��� �"�@�%%@ܜ�p�H�~����ȓ58Ƹ��\�1�ƭr�&�Q���&�P�i�ibH�:��G/��I�ȓ���k�(��I�~ȡv��T���ȓB����P2�>����f_�͇ȓZ��J2#N3T4p���ͩ6�D�ȓ��h0�̛2]R*�c[�k�Є��d4�`-�0 {~i�� .1]��$cr����H=c)b��D.�m0܇�S�? *��.�Y�	��`'\�Z���"O���B�:h
,k���@D��"O*��`�\(#��j&o��@��"O&�:c��2qb5� @6�t�"OH�  L���D*GÞ/N$�5��"O
50��ʑt ���, �M��� "O�={��ZCb�Dr�,��H�̕P"O Ii��"a����Y�nDyW"OV<! ��R��樌	�&��"O��c�̀ �4T����0W����"O����`�5 � !lH�)�JQyG�8D� ��3iE���$��[:E9��5D���G��3u}��Pw��3>X.Ma5D�Hc��A�8/��q
֊Xg��4D��[�KM#I4\II�ԫ`#�e�EH0D�`���L:��0#���+G`	:�-D�l�1o޺6s����Ϙ�&�||���)D��A�&�9|�{��C&';DXpR�<D���$�"����R��<d&2T"9D��U�UđbǊ\V�U��$7D� ;s�>V���q��m�g�5D����Ҕs7�x���X+|-���3D��RE��AB�Dsa�	3H�,�W�=D�P�$���ty"���F(N��� D6D��B-�:%��P��ŽkrҴʧ7D�p郇�$@6P�5�4����+7D����j��ִ��ر^��9ӠH"D�``�"��-�r�y�$��H��-�-D�dB�/�3�6�kH*df���C>D�X���5B�p$�!F�~���=D����eɐH�]�B��Rv��<D�Գ�@�e**q bb����Q�b:D�$ ���@���+����y�Z�Z �"D�09"kԢFC�T�wg�'�\�꣮5D��a+�&x�4������[0���M4D�4ca�P�L��,c񁅚S�K2�6D���S-�'�N�����"o��\:Bn!D�$���[v��P6J%{UҰ�S�=D�
��X�E0�sD�]�`�ڶ&D��"e�J�ME�Z�-֏o�b�p��"D���f̌Z��Q�s���T�@��!D��/	?�0Q@s�\<UD�$?D��A	U<��ds�-�aVB���n*D�(��c���t�7��;]6�³c5D�����P ?��E 3��8�hI�K D���D�&R�<�f��?Y)B�[��>D�8�1i�-s�(Q�wǫyw���?D�L�"�շ~|e{���,�
�H��<D��h��0T�x�G A( ��t@�'9D�,���g�V(�f�C�W�>4iC�!D�$��/��hPR���Tn,�`I2D��*��G�-����kug:D�l3�G�O���Q�[�0Z�8�%4D�d0�b��w�9�*Ү��V#3D�l{Ԯ� E5�BC�L�4�S�I%D��1��L=��xRw�۱y�N-[��-D���$%,_�j��G{9TTr �6D���(^�;�Ƞ��ڨo�2�@�c6D��c�_�O��s)�3&���F,3D���dҭJ/PQj51Tu�
4�$D��+�̖M� !�A��'��8�.$D�X�i�<����"G^�:j�\��#0D�8x���^�h�ia*iܤ<��!D�"ҏדo&��! ܕ	�b��wf+D�� h�5�Вjqd���ζP"B*�"Ov,q��@�{�Q�d���>,y� "O��#R��Hl��FJ'$�A�"O�Y8�+Sprxhٳ��V�%V"O��{b�V^�
و�g�Ic8�"O����9Ii�A�FT�%xx���"O�|�̗�#�n}�҅M3)eD@" "Ob�Q�D�4W�0x���]^^���"Of9M2��A��/�n�V6n?D� ��GD�I��B�O$�u�� =D�Ш�W8S����̓'3`��':D�8#E`��d�k�'�W�AQ��+D�P���ߎa/P�S��;�@���6D�t[�̔��Y�F��"Uܱ0��8D������TZ���D�?3��u�q�:D��hC���D���F�K�;�Tc��>D��زDzB�#��G,rN�A��<D����(q�H[�BF�����ń:D���/C�}?��0�B�pD,E.4D�sQ�*V�x}p��߲<m�ab"4D��Z&��$Qmx���/V���%�3D�@)�M�8��=�B�%:�vX���6D�0��)��N$���.�3^�`��b4D����.}�d1@�%�"�k��1D�Tѥ`�:?0�Fj>X�V��3D�<�h\���\k�
A9vk`A��A/D�B!I�a������s	�.L!�dV��"�!'�\afH ;!��C$=f- ��۩ D�6g�}�!��9J�`s� �6R'\Ȣ0÷m�!��;f���`l�\PŪޔ"�!�$�	l*�q�,� "�H��e	J�K�!����� �)*-^�iI�!�Ĕ�5*$���zh�ѓJ��!�C�L(Ӭ-/J��r���H !���hb���w�
�p�����i�!�æI���+5h �2��s�����!�$�4Z�l�)�i�� <#!�T�l`ZB��g2΁��@�!�D]8G�3i�:M~��"��3q�!�+	b���C?eV9��OJ�!�䍑T�kA��a"�����E�!�$��(k�PY."���.9�!����ꕁVh:t�b�֣�8B�!�$A� �h���3#�ģ�%� Vl!�E&/�H�&̤0�<��$�V�RO!�d�7w8��$hJ�A��YB�զ2!򄟋(���!f�IY���p�O62�!�$4RG����G��j�xv�٧[M!���Z�nICF�S Xr�b�5:�!�Ĉ�7c�Jv-ܘ����R!��n�X���:�p�v͡o!��]�T�T�P&K�I��D�o!�$[y͂�����c�V�Kq��R�!���[?����,�~�v
�k�5&�!�d	=B���bƊz�n�#���H�!�DU�LmT��"iU1B�^�)��ͷ) !��$?�ޡӓJFh��G»V�!�DK��]8��э	n�Jc��7!�ձ[Mz}ڷC�(V�h�7�7D!�$πCZ����Q�>R�]Iv�##2!�dQU2 P0j	</A����
"!�9k=�e
A�]�-H�R�.��Y !�DN�,�`Ycmޠ|�M*�#�1T!�� v����?X��+ʘ-v�$"O��ڐ���U�.��#+��:����"O|�
����~���&)�1#�~`�4"Ov-��#��
�*��D��½#�"OҬ�E-
#K�� �T�-�~
�"Ol�ӧ�m@"Q�a$������"O�]@���$��J��T(�D�Z#"O@����T8:h���Н�.�a"OT��WF�6M|���b�$����"O|%���[��0����ݮB�:��q"OP񩖇'c&��G��5t�@9b"OD�!u���)e4��O�PIyw"O$�3��!w�z���*�V䩠"OR�0�Ɲ�tU�=Ф#�dA	5"O\��}Kd�BQ�	:�<��"O�4��D�O\�Õ��.���C"O��cIV�����`B�p�Ҭ� "OT�&��gnT�@̑?�b�"O��Z�@0�F��RV"�bT�<1���#d���n��]�yCǙg�<a�`�r��@�t��s3�M1���e�<����f=x�J'!��-Li#�M�<a��V�p�X�qC"�G�\DIb��E�<)�a��
�p� AL0�XW�<Q��C0 0 �A�u��QeE�S�<A��A�S���`@�ϋ�r��N�<1�M7-�>�y�&C�~gHaj�h�d�<Yl�0=D �W��8�L�@�΋a�<Q'B�i��=�2�+<�r%N�f�<�&��>@mR�#�&]��i� �h�<�a""���EE!<�u�"B�k�<� ��Z8qf�ğJ~,��!�b�<Q����b������@C&�[�<Y���s,.)�#�_�<`̥A��q�<U�I�O{|YR�C'g��U�n�<�%�7�\�B�!¤y�����)Gh�<��fO�W��!���)h
��7��e�<��
3=��s͉�F�ၧ��L�<��o�8
1h�p Ļs[�0S��P�<��d�?Y�|�P������L�<�fCQ��3��9)����f�D�<��kA%T+��c�lۏFr ���~�<�` ;|�iȀ+ր���R�|�<����e9����GQ�:(�pb��u�<��40 ���*X�Q��X�䭇u�<ѥ�� 0H�1�T�6��|a�o�<����n��Qц�UWr@	�˜m�<!���X��
��|0��HR�<� M{)��|	@��ao)#�~B�I�1:�@�N�5���e#A%&�bB�I�?��X@��@�_��C�ɧ|��I���onX�ZE�BE�C䉌2G2 �wNH�,T��N��&4`C�	,G�uk�"c04��BIP�6ÄB��/ R�փr��U�fL?j~\B�	���C։@�d$��Js�,	�"B�I��&4ۂe=Qx���AQ�T��C�	S�4p0V狔]j��)PNLM�C�Is�B|0�(Q,"3�̑Sk d���?��?����$$@F�ϬR�M�D(�
�y��.�j�'A�O3䨨n�6�yrm�U�②�d�/�B��v!��y�6 h�yj5%��R�+&����y2�N"X�f��E)�\��Z�0�y
� ԝ��&��@��f�˳i�8���"O`yaDE�^�p��7�^�j=�t�A�ILyR���X)��g��$�PbC�Ke!��O0o' Y8U�I� � �*g�ǀ~T!�dS	���Њ�<!�8Q��GC!��	�[ލ��ϖ�h�����,'!��#���¬N�\ϲp1'KX�!�dX+dA�xb��Q�y�d��jP�r!��Ӗ8.Xy�ri^�*�"���FAQџ$������|�B6�T�{P����D:pM�P�<i�C� ��I��M���Ź���J�<i# ��W��Dr���B���S3�G�<IP�I�4�:���ƃ�4����ĨJo�<	RF�2�6@+��D�0�;Ьu�<�SJ�6t�����c0�	��@�m�<B�+ .p���ܢI�2��b��l�<���R8���Is�US4jEs��'T��
Ս΍kf���1A8s#`٫U2D��+U�}R.ðj���8k�J0D�|�e��4�j��^�q��Q��/D�p���u�ƨ�p	��YC�]��/D����-j����4�וhx)�4�,D��q�[U4$:��Ŷh�4*D�6��B��k���V�X�b��NL�<a�DRCR�ڲ��9u�x�9 ��D�<�Rg�<�:x9��R�����VE��<94C�x��
'Hҽ+�D���V^��%k1D����h����G�#iI�=�D%D��yg�Q9\�.(@��ً��-)�A"D��� �@)�J ؿ
���*Q�!D� :���{X@��A%���A�	-D�h�j�q�����D��l�8�)D��rV���~����kK�hsׄ�<�+O����#��)�A��&��c$.��q�!�ĉ�FA��㳧��#�0��G�#�!�dѾ>�FaʳxhXl�#��wt!�ڿOzRd�!�(� TsD��
b!�D�>\4a�����A�f�ZsU!�D�o¼�K �C��!�~H!�r{F�!����h�d�ʸk!������rr�ʑԐЄ.l_!�d�[�I� �L�Ftb�ퟋ,�!��Dm@��! ,	�*"Ԡ����W�!��X�ıb�R"	���p/F�E�!�4c`�(�jӬ	��xQ�ěOg!�d��a&�!ye���^b���.�.D�!�D\���[�I�|��bpm�)|D!�䐿f�@�0��)��(�k�|�!�� S�z(���WkUd24EܒQ!���r���(+7�r��Tj�$C!���	A���ED�<��3t�)!�$ľA�\�A��R nJ5Q�Iў,��I,9lK�.�0u�0�TJ�3�B��e��p`0zībkK�,���'�S�OR�e���+phf�R�[�	>4�+#"O�2���*fm�I�G,lPJ�"Ov����{����P B�]`��"O�P�������J0"�&��"O�,��fX	Fl�h��"9�L4k�"O���ʓy��V��-����d�|�)�G�"Q1��"e���Af)@6���?�S�O���S�Ɔ�|���:�c�
)�F��1"O��pa����`���Eu����q"OB]�PC�*L�u��)\#��Q�"O� �!�(=��(S�^��<M9�"O"	��Ɏ�Vk�d�C�Y�)OL�X$�|��'���>����0HI$��d%��{ c�<	w���p��y��H0z��M�c
�4��|��|��D��
´;��+�H�b�m�<2�!��5��d�(�����pOF�s�!�ϱei�D�c�Aw{`4�$�"!�d��� gM�Ye��"��L
�!�$E�������� D��!���'�|����3WW"I�U,�8���Ȳ�4�vC�	*Q#*�˃̒����z��U:���d�C7�"~��bC�����'����k9�܄ȓET�ຄ�,^$��B��Tk�E�ȓw��C
ٿuo0e���%�Vd�ȓ1�0��e�U �Ar*̞W����ȓv�2��W`C�ΜMQ�l��l7:��?����~b�%[9(��j��
�`�`���YB���hO�'
8�9�DA�.q�HU��'o�6�[wl����<E��'�0i
�(��?��=[0B�\�b10�'�Xܳѥ|��GH4M�>���'�yxЯ��n�"�����?�4P��'sDt�Q�ݘ8���C�31�t��
�'�l�@��ؙ@e���@	��W��1���hO?!Cg��b���4`}��5�h�<	c˂�Mhek�ծ=((�BT!�⟐F{��ɚ;;���2
F�M!lUcD��)FB�I�'^fܒ�%E�c����C� t$B�	�?/���m��P;�]�Sn����C� S&��\ %K���C řS�^B��dM�$�Y��a�jX�˚���;?y&%�rh=33��K6t��ey�<y&I
<��qӁo��e���&�Q��`E{��)�h(i9u�P�n���jX�4�|C��-$)E�R�)���� .�.x�C�I=!��q��/͗ Z�M��C�7��x�a�<$��Y�GB���C�I�E���w'�*ފ�CIڔrӲ����O��ɮ;���y7*
����B���0�zC�Ɇp (��Yn8�@�V��.,�T��/�S�O��Ic#I�tډrCL����v"OL����Ӓa��u�4��+H�:�;�"O0�Pr�M2d�,�R�� 8DV*e"O���q��)F=�HDn�$��W�'���"G��$��J?T��w!�?qbHC��<	��z`n�T��`��-�#�nC�&�*���ؐk�h|�Q��1˞��Oj��{�'�v x�@�YI��Aqc�g+�'�f�؄��7Y�dq�	��� ��',5��D��4aES{.�L��'2�0�ԂXH�AP\�o� y�'���+�g#$�\ P�,P`��8��OP� f@D��Y'��r��"OL�:�e�]&V�Q��&x���#�')ў"~����)
0d��L4Z�đ��P��y��H�>��£OB-Pm��9t���y�)+G���c��	<I&��/I��y�A4�z���K�lp@���K֕�yBd�F�ڒ�!e�����%�y
��Nm,���X3gG&!q&B7�y�hC�<~�c��\��BA��y�A�|��ԤV�\� :���yBd@�Xc�|(�B�Lx� q�ė��y��?>X,�`K�G���U�Z(�y�h��
hIрǭG�"\p�I[��y
� h�c�"�.��)���c�J�{%�	\�'8�hCF��v��:��
�`�+V�'�ў"~"��W'7��k��O�y*ѳÜ��y��>.�	��_ o�
�R�H��y��=C��z��e��X���y��ٟV�^l����[ P�1
��y�cܐyҔ `���L4$��)_ �y"i�'.��(�"U�w�|!!M���O,��?a���T�UB�P�������$P����yR-�V}H%Q�ʊV�|�nS(�yb�
�7��iy�D��N�\17`�<�yBHݲ4��5��,G��5	4�Q�yRUd(P9RӤP�:;@�s&��y���?.T�i��o�<1�M��g �y���38�]��#4y��t0�����O���.§4�d����L�s:��d�א8%聇ȓ���� b��MU����&��v�z��*�.�D�Y,��f.��[�TD�ȓi�A@$å��8ۅ5"��1�ȓJ� i1�@@�~S�bƯ'^�����@�ۍ7j�D&^"�6��ȓK%��q��T(Rٺ�@,�,�F{2�'W?��/�3¨H���:@s֙x�N4D� �Ao�5!���4R�Sg��2f�,D���D,��A�������A�%D��j���8Ch��z�$0D�� 2'�h�TԢ�,R�1%���7�8D����δ;g��� #���8U.8D�,��	J�~�z��O��v� �<D�X��ȬTDZjpKLI�J4���:D�p:��Q�]0�PA�--$��ah9D� @�nÅu�bXɞ�3�ꝑ�<D�@��E]�IX�0��m��bd��b	:T�02fF��4��cQ*u��`�W"O0X Џ��"J�:C�
��-C�"OP|ۀ担q�N����J�n��Tc "O~-+�^��p RT�U�]u*�d"O���j��|j0��/8y���"O��À�M�E���FN���F�y�"O:5�W�g~�5���ϙZ��YA�"O��0��5�~��2Iމ;�%��"O�8�` ȡ^^��g�"���2"O��J�gV�oh�:UȂ|�@��"O�C����M�ȍ�1�S�K��l+�"ODi�D�0�"��䝩5�x���"O����>l��*��C�Dn��hF"O`���F"^�A���3GLL���"O&��j�V���[����d�0@"O���%&9^�F䡤oM�[�d��"O�<�hu*,m*g�A�4��"Ob����F1	}�H��Q�&���k"O^��C�����H)f��E�x��F"O��c��#�LxP�NRV����f"ON�@3ژ1�H�$�;z��r"O�%b��3D�M�#/�N�����"O~�)�+8(Ҩ#�.��'���6��Y�ȳ��i��}�����nPS�+�D�O^��� "Y]D��ކ4��3d"l'!�Ĝ�JT��|����#�
e!�	V�T�3�N {^X���aW�%�!�$�0?/hC���z8|� ��
4�!��лz�|�Q�똨%&��z�V�1W!�;c�nd �Fk�8�"\;�!�$%�Ԥ�v�4A��ҁNC������Iz��� ^�J��E#p5f��$��2ȂuYW"O� ���;��a���W,���	g"O0�+�5-�B����MB�X%�"O�z�
S6�hL`�Iʜ�Di"�"O���f26z��5N�%TD��"O
��F��5f��r�,_Op�"O�Y q��+X�5,���	H%	E�m��Q�H�S��I�{a~@� ܋K��� �ϝY@�C䉋A8���СZdJ`�4�K�1/�C�I A������3��١'ʕ�(C�ɹScT(����!p�!ܕX�FB�	��H	��ϙ/�ڹH! �6tB䉺b��2'd��<h�xP��;:$:B�	�L$re��G9�,l�c��	v��C�#Q_����L2Yn4؁@iԉ�jC�I�_�F̱�J�����w(Q"�dC�	�k�&H��FS�	[ȉ��,	��4C�I�Gz҉���Wy����"!(�C�� Ӗ��W�V.|�k��Z�Y1�B�I*����`D� f�6K�%c��B�&3�J��2�ۓ-��@�ǓNFB��o�ٛ!�	9L���d�+Q�C�	����G"A� ���ƍ�Da�C�I/���!"-ҋ[��*��L�Q��C�("*�����	��8à�
�uaxC�I!<Š�R���b�\��cE��pC�IVT�(���hGv��򤈡z�t��>��|���
�jw�u`��]lGƙ e��8�!�� y��y
Q�Z Q8��wc�8H!�dџW��Y���%wN��RGiM+!�Dч�Hy�$���K2.�)�I��!�U/0�3��_�z��Xy��R�!��ؠ|��Ĉ��;�l��%��<�!�dEP�!�E�$A��vH0�џ�IO�O�B4!��Q�N����A�D��'�Ĥd
�Q���Q�:	�
���{�J����`K�+��u�!�d�&<�&���d\>V��ѤjαXD!�J������\�EE~Ux@i�N!��ؘ�����M�f��E�ah
��!�D����f��%7i�Y�ӆ��'aa|�
9¶�ӄ��`B���y"��(̜� A"�����2�ۗ�y�Dޛ"�0�Kd��b�D�B�Y��yn�8�����j��T��\�y�����#�9ic�k�cF��yr��$e�-iv�(u&za,��y®��\��5!�2jʪ���g���'aў�Ov�
� �1-Ju*��ڤG����'�d]�
^��J��S2"A��	�'��ӷ'�
�a`�#t}��'n��Q�M4$H�����	�z���'��=PP��(p��3�k�#�<��'R�l��L?~씋&
ӡd�V��	�'e"ećX@���EW)Y�X�A���?����������K�� 0V
ŀ�K��һ B��m��$�*F�7i@�f�.�C�ɨ+�0l�sD���	H�Ş�k�C�IT� E����8Rj��OپC�3	Y����C��	�̀	dٮC�	{E�m1 "�̨�d�W�B�	�3�ni��� ~�t��A	����E{�O��d��TT�(A��f*��B^	_3�)�'*
&�
���-h�@��Y�\��LX	��� >h�4E�"6���ffI�II"Ox���bE�E����Dȴl��њ"O޴�ƣ�(4�zfe�(��=�"O�I9�Ja�b�"A.��.���"ODW�h|H���Xj�����P�I���OC�� ��aqD�%@_)K����,O �D1��p�'� �c=&�(e���ݴI�$��'�n䢥��WHTh�"l��Cs|L!�'	ɘ3��uVH��ʞ�?���3
�'�nѐ��C+|���e��>hZ� 
�'��ӧ��� -���5�K�2>�h��'(Y�h�jؠ& (�̂��D*�`�I��B;� ���R����'�ў"~r��Ϳ4�v����(Cff$x��yRH�j"��Y�`K:wz<P�Î�?���S5X�|��͓~}fe�Q�Y�^�B���a�8ѸrG�) zN(�D-�J��ȓ&z̅ I��S���(w�U<z1L���F0��Pq��F���S��R7Zj^��Io�IVy���G�(&�p��+[��E2�n�(��C�ɸ9��UK@�ΏU��Y�a��e�B�ɖ
W��dd���	aFA]�wp�B�g�(�rC�ɒA�H�h�ۏ ǸB��5JN��¤�V  m����^#�B�Iie�)*��Nh�TiiA�A4��B�I(#�����!M��y��ԏh�|ʓ��$��)w����MA38$e*a�"�R��A%D� ��S�(���1�dةF" D��kp�Z-_�T̛v#�"�h��ad?�Il����	 Pp��#i�2Eֆ��adV�LvB�I�fH<�g㍊)����a��#�dB�I�M�����K^d�Ԏ��38B�Iuʘ�zv�0*�L�/�:C�I3_zpuHs��wmn�ɉ23�B�ɝGw��rE-�fi���H
��B�	�K�IH3Ɛ��P=.")����?	����S�O ���rAX��Jq�RaNd��'��*@��#�R0/�=X�&�P�'zv@� �R���'E%A�*m �'��	GI��V��9�3���8���)�t�������'�59��x����䓺0>�5��	
��\)s��V��v�<�`G3F𱒇� {����b��y���hO�'��,!̟F@n\��VD�ȓb]�qG(F.8�az�J���LɆȓ��d�3*D�����e�)Br<�ȓ,�Z���)�*�
q����1:�2��?Y���?	��IL�c�
Ա���� �sp�,(V!��4	�!�e�߹&�j�al�  Q!��(W�[ԉ�(z&a`5���Iğ��IS�)ʧl[���%Z$&{p�Q� �N����c�� �S�NUjM���X5:D�ȓʖ)k2Ϙ�EP$iQI��y��1�ȓ8��"�G6�j����(�G{B�O��1��i;I���Ë�f�ՂM>y���?�t���?�b�ձ��Os��H��<J�Ju���Z�B�H
�'�0:4�
>z�mX���.>�^I�'Nv$2�I��ܽ��� "=e>�I�'����8\�Z8�J�9#&��'<�ɣW���kN��# ��>'�zY@�'�&���́	�dç�ėLR�9�'Q�aÐ�@�C����W+�t���S�<dExb�'���xp`ۀm���#Aٚ�y��G�}�(i�6,o��\�@���y
� �0+��L�s�� Q�^�~�|�c"O8Mj�'�i����C�09��i��"OR%��m��T�f�h�m�"V<:02"O�tу�'���C�TY��T�'�'�O^��!?�);���ᢘ?{@f�E��P�<1f��6N���J�	�:Zl3���h�<a�$ό�@�!L�cDݺ��{�<i��X�lRX��	��z�e�\�<Ѱ�{�0ZB�f���u
FX�<�QÕ�=��PL�|�9p��V�<a@�K0�ҴB��Jz�(]` �V���hO�R^&�a5�$�Q�cLn��x�ȓH.���J��U�F8�-�Zo���	_~B됪W�J�R3`ʴY�h(�t�^��yrf� h��[��Y�"��GE��y�'ՠjƔ�Q䜛W�� a�)�y�[�M��9��P\"�fٵ�y2�ΫN��@2��[M6�kl߅�yRn��3U�T�'S�E�ȹ@5%C5�y�N�5gs CI�P�h��DGۆ�yrd�2ڢ�(�ʜBt�X�êT�y�Hٍyr���@ϻ?�Q�")��yB�лz��Q��F�<�t	{�$���y2IK#M�A�#M!6��U�a�X5�yҬ�df�#�
)3��	X��y�Ƃ�v:���ֳ1�$�Q��*�yҢѨR����������B��.�yBL��z�2�A���a��oE��y��L�!>9Ġ�*>�Q����y��έ%��S�I9N�QF虑�y⢅)Gtz9��#�4�ڴ���yR�؀EX���%ɕ@r�����y�!ߓU�ܠ���t���aumM��y��)P��Cr��>���t�P��y��[w�D��46�&�s����䓒hOq�n5��0��)�F�i`���p"O�)��"��\q�n��r��"O��j�b��QrT�Ĉ�"O��1��E��Z踄J�?��p�"O��(��\8"�Ĕ�E�PN���B�"O���a�R�`  	f���_ƶ�QU"O$eB0�F�q��oS�f����&���O
��&�Q]~G�FS�D�F�Z��	 	9#��Q���5aC9A����K���Q*		N���b��o^9�Ɠg3�"Q��6om�c�oT�KҮ0�'���v�K����Β�<5J���'\�ppU# X(�Aē�/�ȹC(O�$/�O,��M�
�z�j�G&EL5�5"OZ�r&�O�����:5t�"O�(9��_5�
]k��?Q�=z�"O��� ܕ0���񁯄4D��iy�"OJ���h�
^$��R��U�:�(��'R�|��اdע �� �4��9sdF>D���&V� ��ȡ�G<<	����I!D��� �_�p�p��--�n�H��,D�l0�
3R�`�ǫ�s�`��4�,D�X!'��7;��A��=U���H�*D���'�ْ�ĵ2Q�Z�	,%��(D�p�!j�$�NE	ŮĴj�V�{u"�<�I>���O��k��i ����ƙ40�tB""O��Z���U��\r#��z���1"O@����L��
Ɓ�AR�3"O�`��C�&!n�� �;H����"O� D�`��W*ty�$��&]��ku"O�4iVhJ�*�z�#��̑VV6��"O�\``E��U8D�B:!Gd��a�'��|"�)q�ƿQY�]����6�x�B�5D�����i�z���D .e�f��$�1D����  �Uӳ�\��N�K��/��B�����c�n�SS���.�}+VD1�C��	f� �@/θ!wzy��Mr�tC�I�A���� �.ٞ���+L;H�~B��xON�x�n�[ll���G,:B�%BĺI���Ww7ZD��K��+А�	H<�'$�k�P�h�b���|k����<AQ����g����#��� �q�`��J֦㟔�	>!sU�'qd����~{�~-���5D����@�� �۔k�`���!D��
���Uy���]�\�2�C��;D� �����]�$X��nێ5޼ᨦ�8D�8:#�X����*""M~ VPS��O���8�O~Xg��O_�	#R��*o&����'!��$.�Р��˹C� ���aéL���r��`b1�+:AL�͏�_ɬԅȓ5�@��h�8���i��z���m��c�9�Lиb�\F��E�ȓf��Tҵkɐ����ǗU�Ṙ�Yq�\Q&���
A�,y�$`�'�a~�n��`M�H�NLي%HS4�y2A�M�89Q��w��52���
���hOq���x�6�
i��	8�����"O �0ǃ�����P̏ ^f��A�"O6��cË29��"�=6=5j!"O2	;���>d'�KP��o?�MZ�"O�<����\�HФ
� Cx�3"O��)�G	$M�V�P$�ۮ%�n�(�"O$� ᄆ-x����f��X���q"O����c�#��41�U�]P$"O�e�� (-��8cJ�1U��c"O�i!b���}�w� w�,�"O ��a�4��	�#(R!Mn��w"O@� �� �Bݨ@�ӌ9 �(�"OZ��d�8=��J�>a"0PB�"Ot�hN
`D x$�_$%��d��"On��r��!4���dH�e�1;�"O6� teπT� ��Ħ��D��"O�̙¢�:����H�'Ά�{�"O�:�@U�+Ɣ��N�&g��1	D"OX`���4+Cv�k0�_��΅�w"O�tk�N�>e�*�Fѽ��c�_� ��g�S�O.-��	�z��Ր@�+���'����:"�ڹP�ˠym2�C�'�,,ɲ&Q�����A3�,("OJ��Qn�6L�P-�ƯӚ$L�)��"O��� V-%v�Ń%�I�FMd��"ON-�S��R#Z�(wMĂC�(�;�"O�=���(���ap,�v��FV�xG{��酴^��H���G���B��~T!��A%-u�y .���0y@`�S!�d�?BZP�) B:z��$��[�!�N!p�؅�� ÄZR�W��1N�!��>mܪD�%N��$Y�)@W�!�݊J��E��)�;o�:�'+֕k�!���K��E�ʹ
�XسhY?c�!��HZ{�Y �p��uS�4u�!�$-/�u�aϙ8���IW���S!�D��*ފ8p ���ꨲri��%�!�� �c�Αg��t�Eg�8%
]0e"O��Y��7ZT3G��2��Z "O
!�*Әg���Ae�U� � �"O�,�"J�iX�	@ �N�B�b�ʰ"O��0d�#F��l�s���fc ��$"O�D�AE؀F�81#Q�\pd�0"O(��"�X��tR"��r��	�""O�5��E	=�ޡ�� ��y�6,"OhQK�%����G�*��A"O(<0���Д�T�I�N�p�{�"O��{�瓥%� Ba�F���"O�H2�ȊdP #�.�=)^�D	�"O�2b`
YL��! ؒW�"Or w�Фw��I�P�Z�l���"O����ѕ?�|�ޒ"�u��"O�a �"A+Qתm�UHT�
�P`yA"Ob{ǚ�-�f�RF M�.� V"O��@��4b�Rb��}�$��"O�0�Zi͆�r�A�=��G"O��4�l����L~q
�"O�qB��f@�:%�=#X*d��"O���pc��2B��Ʌ�V3#U���Q"O� 
�gO#� ��ᐚR8�U�"Ol�Itg�e���J��/l�U�"O�ei�Âg�<�5莝����"O��9׀�`�,��጖�pw�(��"O�,��l�6IY�I{Em��|�c�"O�X�h[�M����l_� ��A�"O�!��9R�\|�6ҹc�j�z&"O�Y;���CrE��
�"�B"O�$�f�5g� 9xK<jp�)p�"O��*&k��a��U@qj�o~�-�p"OĀB%O�.FP����!z�%x�"OP�XP
�O��QE�\֞�S4"O� Iw��:*}pXk�N�+a:H�@"O*)9���Y����`�Q�l��C�"OTM�R�
����v(U0n�x�h
�'������*�LLq�6Nq�
�'?�E��Q�l� `�*Cz8(!�'C�A�
�!	���0�W�@�fi2
�'o\�+GBU#R1 ���`�	�'*`��EʣLf���GF�t��'a.@�똚�R�B��T79��Uz�'���	�/�*%�%��$578`�'�R�
��9 � ��C1R1�' \y�G��0C���*�T�Y	�'�d���%�Cp��Z�F�+´l��'3<����D)W����V6X��qx�'Vt���b�$2|S�#ҞI.�h�'�pᠴ�ʌ���[whG�P�e��'clh��`	�I�q��?W�z���'�Ԭ�&怫t�@0�ը�?z����'�
�a�S&�5�HO�k�\���' ���7H��uޤ �,�h�(���'����.�Fȱ:�� *h�=��',xA;�ϥ}�j���SR&	�yIS,�HrQ@j�};�k
<�yr�Ċ�d�+h��f��HX��ȅ�y�a�6�2�j����h���tGܼ�yF�N�J��W��]�� ��NZ��y"e��A��툱c���i%�Ü�y29�ر��`^Wx�sSeٛ�y�N�h�f���AI&#����R�S?�yX�;�s��L
���
r�*�y
� �h)c�W�"
�y��Pn$�e�!"OpĢ�B�nc� Wcm ��&"O捩F$K�`��P�mO�0R,�Z�"O�!���V�V�:u��_��x�"O��	�&g8Hx�3.�	e|2� "O���c�<��1�l�-n�F"OVB�a 0&���1Vl�r���"O�/��[��s���df����!D�Ԁ�M.7W0�qbD��oj� �=D���G�.SXY�1A�O�����!=D�p���>_�(��u���w։���/D��K L��2)��-P�D,D��0u`_(#^a�a�KV���rr'D�ܻf�N�`R�QC@�ǒA��y�&D�r'ew֥[�ؑIp�sB�$D� �IYjoJi�����V�@�g>D�l����v�$dQ��B��
�7D���Ҏ��g��ٹ�L�*�@��ŋ D�(�@j�8�1��B)hTF���<D��H�d��d mJ���-#̥B�:D�D[�F,M�L��N^���	�:D��J�W?H.*���o�SY�6�4D� �t�	 mq1C\�)u�4D��c!ξa͆Dy�@ 0�A9Ѡ'D��c�o�x�2���
Q��$�g�:D��p��]l��j֫S"r �H�6D�p����F�X�	c��O[*��4�2D�,Pa���<`�g.�0��|��%D�(��tFΌ�꘬b�T��-D�h�%�ۺV�ɐ�B�Ls�|��	.D�H�n�-|��+%�Q�'f��2P')D��
pȀB���ۓK
 *�����%D�0� ��5yl���e	�8B�a�!D�Ț0+��XP��
v/�(a6~\s�N>D�$Y�O�*Z*��bt$1M�����<D�4�\�#*!⒩���z�"M D� S��t�:���/aO,���3D��u��<�{�,�5
�m�C1D�HY�'�, ���+�̍�.C,�.;D��	G�b�r�bŊ]�
�@�7D�Ġ���L��=�0`ɔ�YZ�!D�@�U��>A>%��-_� =��<D�P�f$P:Z&Jȹv��Z(�Pd�<D� �b�<4�I� �	����g�/D�|���d{HA9��0��0"�I1T��If��yn����ˇ�k7!�4"OhEBs�6F��㇊�-Mh���"O�0i�#�9+/İJ���	Y9*X��"O"��-~��ڢ�߳Z4��w"O�!8W�E!�zq����7�x�%"O�YG#�1wh�2S��1� �"O����
2"������"!Ҁ"O<< qKZ�JT"wV;E�Đc�"O0LhO*6H��2���;\d[�"O�� l�4T��b�CBSG���"O$=��d�YgX�cĉN����yb�>M����sfD��<Yچc� �y��k��}C�A�y�80ƧC��y�ܓg��sՌ�-��0�բ��yr+	���LS�rh�%���y�F�Kl~���膗k
$���ᚶ�yr+T�3��웄�NZ.�Ce!ߍ�y��1!`D0�� \�6��TrQh���y��7f(8�k�� �X��f�]!�y
� 4u��%D�^�$���IY7���"OhYrh�%M�&9��̎���"O"q)Îԁpl3Qf$��k6"Op����/b�0|���&"� 1"O�d`�f��o�*�H6Mܫ9� ""O�9�"b�-z�Ġ-Ʊopv09"Op��.�;a�<����54T�y��"On�s��
}�N�a�ٟG�e0�"O�T�D�،OV`BQ&Øb=����"O�H6�ѣ�M�7eL3}04"O�\9��62kg�Cev�[q"Ob�&#&:��!e�<Z{^��S"O��`�i� �6Ku��k��B#"OfD��E3!$��d!ւa�.t�S"O*K.��;L\`@�C߆�y"O��3caF�gqR<xP@�r����q"OMxT�5_,�M)`	о{�"1�g"O�5� �"N.d`�F�W昐;�"O4�@��~���s�%��9"O��HE�-`!���	k�>�3�'�Pl�p$��:���ч<u�l{�'$�жcR�\ AKW�dI�	�'u�İa���V�H�p�j�}f�*	�'��4KlXazu�ǅj٠|��'䲌`𥗥  �뤈��dq���
�'�ʰ�4��+	 r��dH�c�@@	�'d��sf�| ������_6����'�	��`ۆF�`@��Q%�z���'�Y��b�-,��@fE�4#Α��'ښ	��Ā$����G�&�y��'|��QjH Kz�ɷdB)S�e��'�>��V*HA�������0�=j�'Ҳ"���.(zK7@������'V6ra���豙����U
L��'tv+���}�HE���R�	q����'%�2E@ѧeW�tF�{[^aP	�'�u0���7�U��O�8s��t��'��a���g��avi7q���'�p����4@���z`*	�'�=W% �5��2ix(��!D�: b8p�i��!���a;D���Ƌ_����bI$���)9D�0�C�ߍ#�ڬIe G6d>��[e8D���R�.���G��D�5���5D���NxI�#�,!
�@aa@?D� s��R8T��@�RE(qi�i�C?D��8Q*A"#YhaI��";uxhɷ�)D��Y7���8b�Q3�m�\@>���&D�tKU�!")H�pB���4�g�"D��sv�M�1����5�@�`�٨��5D�ȓvĜ���b��K�l̾)C��2D��s�I�{
^ �,��Z=V�ra�/D��B M�j�zl!��@��hP�2D�������4�F�O��h��*2�O<}�O��S����K���gj��~��̋A�2D�|�5lF�K%���?g F�2D����G�d�8�'቙H� E��O>D�T��'�+u�aX��=@�(Z�#>D��	'kN�e�� �&E�j�d?D�l�Ƣ&\�
���G�Q�XX*��9D�p�̏�/�$Hjbf"k\��M7D�pҕM�.��@#b#���j�0��*D���Bg׷sfN`�p�P�te.��T�(D���Vh�1g���mK�a|ހ�si%D�� `��#Źd�� 	���rM$S�3O����]�Ԍ�ĂW�#�蹱#dS�n>!�$�2�ji����;$�ݳDҡ�v����X�r���efF��@�o,��hO���+���ڂe�m�a8���y�x">��I@�<SܙB@�%����n 1!�ǘRG��r��۽Q�����)!�dЎ
dȜ�whU:Ǻ)����F��O����5b�B���w�ΰ�f�2��7�O��#�)O1�*�R�����}�"O�X
cj��o4���eȯV��	��'��D�t�>Q�4��z����I�tn��*��DRn��yrI�o��q�+�@^�鲤)L	�0=y���W:5fHhAgKٶj�bĬԮ�(Oi�� ڹ�voW���p��hV�vn�%��E{��T!�
B�$z�߄���KU��y�`�!��Ѻ%��ީ9����'?az����T�؉�W!6�^���'J��p>i�>q1B�5��Pj\��i RƎßLΓ�~r�'b?��O�N4+�
�>��f%Yۦq;��ɧ#ĢZ�#��!U�	%��W��{��n�<��!CI�$�����&dS�ٕX!��Ey��)�OvXrf�ɞvW4���E��9��Q2U�@��	p�p1�W��;r���y���Ysh�	�a~2	�G�t1��p�a������>���<��d�Hx��Q.��YGXix��	D}��'�icfg�N�[�,�R�1�'A¸# ��6�p,Yf�J!H���'��M3�ǵ5�d���H�@-v�.ON�=Ys�Ę�.�@w�7��]�QmR73��	a���;��DC��	���/��q�%�7�r�L+5�O�`崽��)!����(6D��y��;=�HHS�+ {b���#�uӈ��m̓e�Q?!���ȍ"L|�ad̚Ίɑ`O>D�(2S&7� sSO?dXEԥ<D�ܸT皣J�fM��K�4%8�$:D�h��Ȇ�n�P�[��	n���o7D�pRb`�Tl��@#�C؅Af5D�,�pFۿ-Z���hHH̚%C5�1D���a�
�/�R �¢�(4d=��;D��pb�W�%���|rdX4�%D�h8��$��
��Q��H�T�#D� Y �"3,�i)�`�' �@g�5�O�II�F��T!r֪}	1��+?"�B��HM&E��Z�[,@�F��0��B��)�L�K"K�*�@� 蕭-E���$�/U���<ad*J!h,�"q(�{��}�؞D!�Q�`jqJ�G�e��I� ƀq'!�P�/R� ��i	*�d��c�!�D��7�VL����a�B��S�HD���D��,T#Ԧm`G�H�\�����!10!����B��E26.���P����9+!�#0�@ԲLG\8��C�ߗp!�$׳xsT��Ś� u\h��b��P!�$��x����C�)6���8���)�OpHP�{�����&�Qwo�1IGh�!BL�:ǒC�Ʉ2X�ar�B�&V<���g�mfC�Iڟ���G�F6er�AE�Z(��
��2D���1�]�/�
[d�C�X��;f`%D��ȡlB+'@�5b��η��d"��"D�4��ߋT%�T�G?V�N�6͟jy��)�'I?���!ʗ�8��T�����K�jчȓ'�
pH7�� ,��@���Z~��� D1A2�]�%<z`#���BD��'2��z�S�π ��[��a��䭟7M�R�"�i���o8�Djs�Ϧsf��Y�'6h1�2�(}�)�ӫU`P�A 2^p���һߖC�	%m.t�f�\��z�#�Q5#%���&������?8|���Av���(lO�Lyb�'oX�%K����!Y0����	�'4Xt	�B������2fp{�'L"�I�`l8��,B>UX�bO&�y2/�W�B�*��F�Ѭ��1c���=��y�X?x�`L��BK&I���!��N��y�L�{
C�	J�"�qAk܌���;��&�'a���0�ǉv���`��Q�;�L�ȓQ���!��6h�L؄�Ѽw��<Fz�g2O^���'�#[��8ũ̻b �%J�በD��Ix����Hȕ@g��P��A9E�p��"O P�G�B�enp`��^0X�QA��'f1O�PL��6�Xc��W$V�bհR"O���Q�D�a�����F����W��;��)�'M��2�C���([�"�M�rl�ēR�J�P���
� a��Y�"�8��>I�`+�OH�wj��p���C�ɋB0H��"Ov�eH���R�P��V����xb�'B�0rA�I�{g�"&48��x{�'�h$�7�
��>U�� �(��p)�'�LEӕ���8LXǈL�I"ы}��)񩇘N����kFƄ�ZAMA�2�!�d�;w��5`#"��`�0E���["=�!�$�O���Eɐ�̚Ē�K�ay��'[qO8��4��%W�A��툐A��ȥ"O��a�FгA�9�r�P-N^��"O��� �ϟ2�����q�.���"O�����,� ���3>B�0:���3�(O�c>�j�&�
�� ��%X8H�����$?�S�S�k�u�s�W@� ��b�tB�	n���bR0Ն�q�C�;�^��d�<a��+W4Aq�JE"(��+�W|!�E:6)r�҇a�'o�PH�-�/o!�c ��x���;��S�?$o��XF�d�K:SR�ܘm��4 P���D/�S�Of�!@֏�y��0�S	�2#�TT	�'�hI1*�7k��p�+p�h�'G`�A�#�3Z1�8��%?����B�)��<�hT9�, "t���Z��&F����'�a}�J4x�4ȗ(��~8
YzBJ�y�� &~�XƦ�eGɹt� :��?A�'����G�Q�m1&�_a��
��'�>E0�iq]��c'#�2;[�����5���2��3�޾4$p
	�T�(Їȓt�<Q�G%O��!1@� �d�dH�ȓ4O,|&��6q�z̐��&*M�)��x�.���.�� 2̤���l�D�������9��m�2J�ݚl��{���*'��L���bko�D�ȓA莌H�郭iR6H*w�g���ȓn��4[�L��,.�`Z���[R���ȓC��@[��ˣU�|˕�A
xt���'4���AC�h�8DB��d��B��a�r'�8lET�qҭ�i��Y��
L�)�B�Y=!A���[T���W���؁Ŏ�D�ũ�FA�u���ȓ]�*�䚔Jæ$z���c�V]�ȓ}c��G���Ň�7)���"O�U�G�(I��!�\x����ʡ�y���*$�����)�g,Ξ�y
� ^l���TPґ�jL�+L���@"O��� D�<:N�TKR��j,ne)�"Oz����5�̨��T�(�T��"O���`�Qܰ�Yu��n�ف&"O2ܺ�O���
V��?R+x3f"Oh�k5σ�:H�|���˖u�v�9G"O�-�f#��5������K��� �"O��ң�k��2�"�f��EJ�"O����G�\�&�BV�N��j�@�"O�a� % ���E�3m��3֔p�"O���Uj4sy�L�k��'��"OJ=� Z���ēd���3j`���"Olt��%�@�iႦʂ h��2""O�P����8 vdR��R�n3h !*O������p#�רc6x�"�':�!��Z%o�VT ��<
�:���'����&�&I��� 3��i��'����B	�{�y���ܒ^~���'۰a0VKD�j�
 ����L���q�'���ZTk7$5|4@Ņ�6TR0��'����$G]��9�U�^�'�>4�'X���cf�\�2Tݞ	����'oL��K]#�D��&C���)�&�2��	j��U<k=9�$�Ш@��=�d��h �92͆ȓUD��F(J1=��u�f��E?�؆�2��|pCV�J��0J�^�V�r��,���杸>ݪŉUD�8XNv��ȓ\���6�ǄBN ��m��r|��ȓe�TY��~Pec�*DZXx��tq� Y1�T�W��b�*�0���\�x�҄O�
z?��z�̉�X6� �ȓ<Xข1��0��7C!.�椆�k�(�I�BF(m	����5���ȓo�T`Icm C7�0��]�5�>d��2d�H���!��`a�JM�M�"���H1�̀���#��I��ވL�d�ȓZ�s(�U�Y���" �P���;%�� 2�U�|0�a����񢕄ȓo��% ֨M��� ��bZ�a���ȓJ[L ��(�$q�(Y3�^�*��m�ȓ0�x�J֣�a����t�>`����Z�>�;b��6�N�bd���p ��ȓYU>)��U�04;T�ҲQQ���9,����|B��.\v:W#\O��e ��\���
��T
�o �db�,�)T=��ȓ�Ni� )�,YP����?^�'�����׎>X��1��f�O�(͈B�v���A���z�0���'LԥA!�Io�t{Q@�1O�6А���v�с��O�q��!�u�g�	�?TU�I�Yf�l� z�B�������\�`7+J	v���`�/c�$��Et�����r�p5�T��:���F��U9b�?��h�9,��h+P�O5nX����|�)�g�2d�<�J��2?��pF�0D��� A�+(*�1����	����f��DYq�Q��&l�w��7z�l�pE���(��4J�h�Q ��ހ@Uzd�u"O&e:��I�&A!qL �%o �"���$u�� ��Q�4r�Q)W�&a2ׯ�&I9�{�C�3�����9(�(��'�0��<����)�$��G�1=�${��@'n,q�h!RhZ|��U�X�"Q�y�"0��Eg��Lj"왑A�3C�T��.�3�*<�@)Q=�I�7*U9HN�)�#�6dl�rE����9KN�=kA�k������J�z܊��Yy�'���&Ko�O8�ч���vu�CM��B���)�a�,��Pk;�MY�n^�g,����J���!r��ϻ"Z䘉��\�HM�F�I�;�%NYʽᐞ>!����u'f#]��V�,^���ŉ.�bB���1K!f=�ℍ
W�䰢��"U�9�t����'��\�� �*���ř0 N�d��4Z����5�0N�(8��.Gb D1�I? ,B��
�S�(�C�5�F�Aʓj�0X%�Q�g3`��<��Oƈ*E�ĨL]�=
� �ǀ ��ys̏5Xu��+5�[c������P)��5��Q`-^�2h����ϖu�PT�����)[wR&<�%K:®����E%K���[%BP�ʓ�$�f/���]�!�t�_��B�'�԰��N� .�T<ZF�V2')�0¨�o�5��jĠdp+�&���S/�����D�߹X1���d#��.,�@J��5��õ#�<L0��I�U�tM�'n9Y2���D�Yy��9~�����wN��X���-#, �Z�o�U��L1wDڎ!3\�Z"��/`�xE(MsE��0bc�/''��'�޴x�g�;x���R�$E<`\��4r���ǭ�%MtTJ�S�����?5� ��iP�Q��33����;D班UQ\�2Ǭ�^����Gr��J��q���еX����s�4X����]Opz�:�lI�}{�t;a�f�����-VԐ	�ƭ<y�f]�2��L�6g�h_�c�����Y,SҘ�O��<5#�i��k�GW�/O����΁T;\ ��a�'yv�D���Xݴ�>��JK��ͼ� �մ㨰����?��8Ѣ�I�	}He�A.��)�S�M�*ւ�� ���矙$R���A�*kǒPاE�Hh����M[��R���l�~]^`��FJ�Kٲ�K���
��t�EĔMa����]��ល7l8	��&ݕHD�ܙ�̂ �#�#(g�}�N:�<� ���3f.=�"��OK���Ӭ�"�3&R�>Y�`AM�
|Ҝ��b޹Rxc�#�����`̻*���'_:` ���5�~�����T�0 �RA��{�'�*GԌQ7 ��dE9Vx�����sj}�ǠA�RC��#gY	/MĨ�@֖{ t ���&�r&O�"�&)�6H�m��	�@�Q�m�	ݒ��C�%P���X��$�˧s��T{��T3���(�l�0b��@��1sZ�qc�މ��%6k�w��HK����|:��_1f�����aB�B�P8�����) �(��0i]�'.8�ß�"���:�H"�S�}�Fi4AFH��9"�ě#1֐0���уI�`%��B��bN�-B��H����1]#�zFdڠ7ۆ�7�x��t?D��Ò�p���I�z2��i���:=$U*���B����M+`�N�|Q�R+2�v�sF+p��RA��FD������!Q�P��GY.�(d;Ԅ�*Y�8b�`+��X�X�>��'}��W�;rEP�C$L�'161
m�	x����:E�,lj�C��uڬ�����tHF��� <,R�mJ�z�� �;4Lqa'�ǝO8���I�EܓI�����"��<z2��g�>C�@�<�&)F � !�@����s/�a�:B͇�J�l@!>�*i�0��Y���ہ%Ev 
��P��̩��'r���7ǎl@t�B�"͡5E�e�#��6GJ�)����/�4�D�>o�D3Ԥ0oGz�P��"3N���8�P�h��p�C��<y���F�2�B ]��
�;L,��G�]h�6�P��46�4��6g$N����>V��`[jR)i�h�t��K�������mv���DA�sV2L�2A��D�O�my�eB�(� � ��h{���A�p^ d��-@����FD"�U��J��tF�����Y�BB�	�vT ��ω3�|� �q$��G�+������9� ��M;�D4l��A5"�l�;XȬ�P�I��e��4!e��?�i���
qܺ��mG�;L�a勇Wo�����g��Z�#D [�D 5�/��AHo"0X(�K�Sf���J<i'+/"�Ic�H�}u�(�����'�b���d�o�Y""Ofd=�.׊Z� ���@ՙv̡Aaˌ�d�.��Ы*N��@���p`��2,O�3��u!��˦"�����Oa���U�GȬD��	W��8֭O��@�T�
�(��� E�g�����XT�(�܇R����R
�*�E}�e�c|�u8����^�(���Z�,i��_���+E"շ,$����4��=*1. 8V(RE��B��3�^#��%"��'<��XJk�����#4.��S`�"�t�|Cv��6�E|	꼻�˻".*��'D��~>��`˺'%:ĺ�&RVÆ�㡌��8�x�dm��j$�!��	>�(��!�%KѦ�� &��Tƈȳ,�.�ēp�ݻ'N�V��,��S6�!�-�<y�2�JU
��>�4	A���p�͋WN+R�� �㋓�0�%i'͑�$�����R�V�f��c�˓�KMZsf���鞩O����E�
�(O����/ǑYth0�2�
�3h�c���M+X{%P�/�����1&nԍۤ �4P1��H5f��'���h@�@T��s�FFQ@d�5��%6�ƐB��N�'�����GBYPD����'2�֌r���>�4�� ��y0p���6�8���'R�] 8\�w�Bk�m;a���Hp4��Š�z>d�K���2���G�+\����H»w:����LM�:��ӂ�i8YP�Nv��y��tP䰫��Іr�` q7��q�(���8|=A�T���S�9+��1��A�Ms(tHq@X�5�b���2*�L�dG� ��{co�x�I�"�꽋��X�=V�0K���G��q��_9��	�#��UZ��	d�M�&�����)ز?_�5��@�����.{����j�"vQ�U���r����Z�����\�J"=)g�΋T��a�So���t #��R���;���F���	ǳT�P*\�Ul(�@�Ę�r0oZ��F����A�DL�(SC��t ��Y��O �9"B5'`4#=��;Y��1$�
 ��(s�!4��{�U1 �x�rl	?+{,��F�X��B=C2L�( ����炩i
�}kphT3%�p�2�,�=-p8��& �6��$̏�.�Fm1·�3}�1q�3:y��%�)n*��x��� C81��NUС���]4o�8[bd�<)W��Pg��Ӵ)�3'ln8�N�_��x�L�!3b��E���OЈO��Zv�MK����k�����ʨc,� i�ߝ_3�A���>"���"�b̐O�����Xm���[��
)c(���gl�f�f�PF�W�L>8!���y�X�y��'�lX2���GLW�&6&x���*������PpjaybCB.v|��iʛg5�qg� 4&|m�yX<EIc��O���r���5�D��zŉ�ӅO�D0@��DQ�7�J����[..�D�3�F�
K�q���pc���+
�'�|�t �HT\ȡ�8��l��bL�O�$����dكkK�!�p�OI��zp���v	h��٬>�d3�'f����Wی����L5v��Z F��zH��-=�Lc�.�.b8�q��1?i�M��+݋|�Zl[Q�S�F*�&ܥm���ꄴ�0�y��ɗ���"����H�3�ӈ*��MI ɚ)�����$:54��,ߕ���B�
���\�c�
-��a����.��Y�I����� �'|/�i�@* ?�a{��Ż,@]�tC�I�&���dU�Y�0�� ��M>�}�4�ӹ[IX��eHS�p<���c�N��fK)�SdZ��� ���gD'37�Д�	�h:H�������X��}$b� h ��A����+�AA�,���c�F�5�|�2 �ő0wϺ�6HK�;2���7�C_{��k>�ئ� ����� �n��<��$�\@�R�Q� ���O�^�I�'��d�:.�
4v�X9�!3��Yq*D�a�ҭXS'L�cdm(��X��F,FN�?])��J�HeP=�� �	d��"��
6����D�>�c%f��L���Q�P邙#|�f�ŚIU�P
#Os=�IZ<xL�q���
���ć
�2��ѫ�
�zRn��Y���V(��	�l��t)!a�kJ	��E�� {�t�΍�Aˆ���R"+�'I�o��h��Ӧ(����N�<:�h�qNK���x�i
0�U��ޓe�ް �ߌKX8��I6p?�	!֭�����d�ýX˄H��^g�ʜh�I�NP6��5L�6r�"�
�*��f��*��1N�Q��Xpb�e�)K�	�� N��8r]%��ik��!\���!N�Bq��j�5 ? )�EGɲ*=�d(U��yC���#Yu�'�V���B�8K9�l
e�S�/����H�X�T
@�Wb5K'�]qx@�B�)ƔN�
t��%�uҁ���1ᤘh6�6B��Trs�A4C��"�.�c��Ms�
̤5D����&_�Lpf��%4��E@اG�t1RE�Bj�5�㏫^�QT�A�#R�x(�f�� ?�� ��F�@I�e3k�:U�Q���b�vɻD�3�E�'�M����P4�}�tƍC�lܫrnѫR�Dk��7Jb��0���=)����%6P0�Y����F�z���NЩ�E��*!� �3���!jĹ�bő�p�
̇�	�=1 � �n\�-�~��� _�Gԉ�A
� OnA�� YxT���Z�-rD�i��ٱ�F�O3����ꑡJ`a�v�^�	YiT�ʒbB 4�	jw���.��k (Stn[�P�eÀ+�UTLxh ���C���@E�7�ƌ:0A4^�Q�G�o3�Qwg��!!C�ܗ{��U�V�߅��<a@%\;s���Ϊd������ Y؁k� ͌_b�����	8H6�"�E�u���uFO�`�����R�Qʽt�C�*�(����[�Z�88�r�ϯ��?DÈ#w>���gMYB���)�-c�TIR�B}֬�e���:�"�M�#v:�0�\K��HQ�/f�DQz⧂7 &	K�LY�v�X�`mݨ/����	�g�8�{Tb�1m�RYIDl���Mx3��qutY	�*�ZDZM��z�$g�D�*����H4�i8C&�spzyY�"�9~"iA� S�&\���a�R�G��'O�Py�ߧF��sW�%) 
@jW�
�p1�Ej$�	9u)�`� ��I��� D�� ����/�1("U�t�Y�Bqb�2l=\O�{���+^D�	��!f�\��^;4M̉���#��="j"q��3D /TR�aB��#c�^2����c�Թ&^@!���R&.5�!��~�'���!U��W�O��yKc&�&���"vf�[��
�(�52k�1qB�	�eg]��,�!P�zas���$����f�_��,ReHW�6c��)��Q�-M����[K�@R�dIR�y��$j�ҧ��P$j����$�%Q@��yu��+n@ʈs�.[,`p�H@J
�N����V��s���`�W���\VHEk�&9�(O�5k���9O�: piJ�B^`m�:OΕ�D� �� 9�e&?��;Fb��K�($p�I�GTrq�S�ݲb&����08DH��x����X����V���G��L�q�7�C�����g�-R��U3p�� Wٺ�A�)ΟG�P��$�@�?J�
�"���)��KyܫáA�Uܴ�"��A�D��t��?>r��6fg��l"<Zne��( ��'T��Ki��83AX`�dg�����BFnI�t�j�$�al���P�պb�μ��.ǩuK��b&�����;`�ޔ�dΆ�sA��λ 6���FR=�¥!����c�e*0C�j0��g��Z6�o�����?�@�"߳:�,1�aG^N��ts�CS11���07�ܐVF�DJ4r2"-cCkȎp[�!�dK��XW�34���$����L��P��d$	�#���!��8|�T e`݃NJ�pRA��F��wL�V��$��!���d9~�@m24	�3���i�tXL�rf�N�Fφ�rY`��i�;.�|�P�� �W��mۣ��1"mz�s�Q8l�=W����0BUҠI���E������9ch03t���u
�mH�,N9]�%�&G�B&Q3��̘��8
�bY�4��UzCB0�� 5��u*��Ѷu�ܬa��
#1-�ps�$5 Y;��wm:A3Q��'= *�/7$z8�)w��6F�}ړa���\t[�grd.U;$�%9<����yw ��{/<EU��f�(�����(�H�Gb�VaR��=.t��� �$x)4I�O��a�F o8ɛܒ��P��B'){h���f�?N���IQ�ը�?��&�Hb<ͻ�n��D����P�yo�'�H�14MP�uO�9��nW�}V�4B&�ŜG�qS'䚱N�d��7�	�g�@�4-4sF���NW�z[�<Jh��G��%g$�_����
6v6X�uʝvJ����K	=0�|KW�!�		<4�`�� 'Y��H�fՔB��r�  �0�2�
F�_kPY��\.sdSC���g*��զ�@��z����2�*�J��ÌZa@E1t��7Nd�8ӵA޷g�N�����I��D@��A%��Qb��/�!;Պ�c�`b0oۧX�F5�ȲP^l��I%�p�����m�� Sq�$E2�|RM�8\�P��PB����"�O(,����9�R�\9O������'%P,t��k3+!��=}�uJR%B%��Ò�]�L��'>�ϻLr�q��Z_�^&>&�H�)�=�.� Ȓ/-�4}�"ދq�Fd�S���>����S��ēM���M�H�L �W�N�,9q��a��y ���ʄ�yq�lۢ���|���M-J�F0�7�N6-;e� ��61N�Y���1M�Xl�օ��b0^1(�ㅚ�T=����4o[�D;��D��i�f�z`fG�5�6Hj�C
Hl�X���|��q)gå2v��q d��gZ�(��Ä'3_�3qkO�PǶ�ǁR�L����3��4R�;�Z�h��pÌ��[�_����46Z���۹m��P��K�x�؁oD�����L ?��X*�<�W�71��b")�z���/k�O>��J*�h���I>M��y�{�D����{p)Q,XE�ԧ�1^�D�ڣj�ZN�[1g��j~.�%*�+<��eo��y)� �f��|b�սy����E�Z�93�)�Vţ���X�^h��'�AE��O�0�O�6+�b8ʵ�W-X�,�b�B�`h�B�]�|ц� 憊'I(��'F�k�:7�И��D�t�>������J
!'a^�`����]!��=�`IF?*��s�~�  c`�\̈��e�"u����T"O�  �X�dG%PѤ�@�oK�fq�PkD�I5F&�P���(:JU� �*m��� ��ˉl�.B�ɚ*v�0l��&�u��KU��tB䉈?ph�p����Y~N}����7'�`B��.524����+&��+�*�	!
�C�əI#n�"CE�$���P�L�C�	�,/� �,�2*�,r�l��:<FB�I.��Ũ�M��Q�����K�yBB�I�M$Ԥ�G��26�Q3�ˈx �B�	x ٣M� ���U��L'*B�,��h�l�
�0A��H>Y�B��%#ê�YG���Kn�K"S
�C�.l�ؓ�A�ђ<r׫�7[�C��2��)��!r@�[1��n �C�I��2 ��Kn쐒�'łB�	��y��LW�:�L�D�ȟ-7�C�	�Cr�!bw�l�$hb�H� mSbC�I5/����	g)�hH#�$�.B��8<�(�,��:Z��i���q�B䉌j�n�3�Z�n"�1��P\��C�?��ĹU�Q�g�h�� �Ca�C��X���ª��c�^I��L��C�	�ḫ�PN̂	uDBQ�Q�"�C�<
��y���*2��3/�B�	o*%��eͿv��xak�/qRC�	�d�PHy�M���#+��B�	�p�!�B�W��KeG�<��C䉽����!"�;Zz<��̂�i�tC䉻	Q�1�7M	((} �5A�2xۼC���ЗCP�n�:��r� 'b�B䉜"��a��*@Etbu��c�xB䉧!Fu���	*![��ѱ��>�DB�I�:���0"��a1��I®�!
.B�	"n(x��Y+��#D��zd�B�	8���r�ߢ�|�x$üe�C䉜`q�̀�a9�.��4%�2BC�I�7����"A"NJ�[7�
&(�B�	�iG4y�t�0,�^�Ҩ�,��B�I4V�=�Q�
�ewʀQjĥ_�TC�ɲ*��cT
��K��b�C�� �B�l7~+&@��xln�[֯ndB�I7qF�,ɳڌ
��"g��K�C�I�<j��d��<Hį-5l�C�ɺ`Z�K�G���5���	 '
�C䉣a���	�n���#�mNB�I�sA(�vΙ!;G��5@V*^��C�ɦV���XC�Ҕf�N5ӆ"�(ƸC�I dXz ,_ �\=���F&Jΰ��$C(Vͺx����>Aa�[̸豒 	$#j��1IUO�<YDH�(� �A�G�#��)���8�O)��/A�C| 2�a4��Е�bG�L�@���������ȓ 4.�A�L�!G�rm�R��r���#C��6�z�'�ܙ�4�>�3��H�X�c`�B(AN�]�vm�<���d�$z�,P0�cL&J�x ᨏ�[D����l��P>�x�DO��������?��H,�?z���jCnD�x�B	�7a�l���ǩ	&�yſi#̘Bģ�)@DWG%}�T$��'��\�W����ř�A��"�p�Or��cc��sO�%���h�ˏ�i�	O������� L48��c�K!�d�V�LE"r+>#b1����w%.) ɕ�&���0֣k�,i �bS V�HM*b;�1O����c��E�B]��ˆ�xxF�'�FU��F6zl�^tXs!P����Q� ÞDyFn��0Q��]^5�'�t1�%.�2C����e���RE�L<Y���j"f��)�&��Is�US�2��Bרl���r��P�!�@���e�	��RR�X]�Q�p�e��3!�?�
j�I��xs�ՆWd��aM�,S�|@�$
	�12TM ��]3�p�Z��GĦ�'Wf���f�� \�S)Ct4�[��r���k��Ŏ:�4Ygc�p�$#���]�7W"\iSk�8bx�5"�fU�m\X(���7�V�;��أBk\m���D�4P2|)�kT9a|��c1i� v��-�Jmqp��Ea�$��S3�JY��.}H'd	���GZXyv�QP̅%>/�D��ؘ{��<�&�&-�L��&m�����h�n��m�>�ț�s���ZP	.���0Q��U`��Uh�:^��u8�l0?9#P��ܺ�)���0��c�Ѱq�R�� �١$����e^L4��H&�@�:��C�w��K��Sy��:w�U;0oXId ����w��-ʂ\�z~���n��l��u����)P�������M���FJ_I��=Ң%�~ZힷQ��T��^= ��A8a��92fe1y��uCQ�U��3v�X��?�7@�_?�%Ɂ�`��=2.Oz�0���)"�Q��A��{�	!�� *{t�j�X�F���g���x���G+$��e�Q!D�{y��+ )||�D��v~�r�҈][� j��f7FB7��)R�2��%%�!T��˓Z�B��$B�*�F�26'��M`	�%C�^���L}�"�Z�mR���Q*䏕o������-f�(y�!�$C�Z7�C?�lm�eL�'	18u�d��@�b�������1�'R�p�Q"XE @L:���&��ϧ!�M��E���)��ݲ|ـe�G���cG��� ���KQ-
�\��y�Z<uw�(��ݾכ�aK�|����I��]B�xh�H�.[�@�c�0+���I ��R��I�o4-�B�;�3?�c��b$��0A��rr�T47�N=� ҟB6��N)$�NU[�K�j6�A����E��R*O4��D�C˾�9 �NW�Qb��҃7PL�al�����Y5I0�DJ��	���'0�>8ce�Dƴ��aŋ>]z��V�"�-��S����be+��`��k�>h��ɕx8��:���8�qc!���|���6���P��4X��UC�>?a�*m��m�VNH?
�.�x�F3ޙ��o���@h�s����V.�Jr ��"����;�O� 4�E5	.�߈�f�w��u}����Բhf}#��G~�WG߃O�R#0��7 +v0�t�2ovUC02�`���.I�h�T �ՅGmv�I�=�(��O,4r��̫����D�<���Â8b���UD/i��A�=?+��c�F��YN0��&��8'��"[�o�Ԉ��xRg��m�|��w%P�7�^�,K�@��7 �7H;DٓR�]�۸'��]d�L/R6�0���CЁ��>&�	�I�{˔l�D
�h.ȨP!�S�vÆ4�l�K���<�7,�H���Ƣ�>)����r}�1�V�B~2��G��hy�mF�X فt��U��\"f`�5Y�v�����J`��yE
̧f`Y��o۠^T�oY�1a����,\��4�ç1/2Q�3o�%AҰu��lٲ+�yI3��?�nmj��Z5̌��Ж7%"M�/���}��̙�(�Yͻ[�
�xf�̠Q���H���C4�����f]�c�� �<����[4��Rq�B�A8.�mp2i�	^�r���	�dp(f�^"�h�����)f���r�D�����өE-Q��z�i��*/Xj�ə�*�:bF*`�ܙ	�@�6H��It��**�bh���\�T`D�7�۝@�Ҥ�B�'��ћt�Dj�x��)b3�z�'�Ԁ�1�Ǎ2�Z�b��ڢr����̻Ld�8��E+g:�JG�޽H�NdB�1T�"D!@h�$�O��Òm�#��<pW��:r��=(�&�`�΁pJ�<���G	(C��oB�a�nH�$,�p�i�5��Q7,)p`YU�^=Fu��)�O>H�𤐂��ɀ�

�mtn��҂�,n�8�YÝ+�����G�(#䪖jә!;���"
�ns`أr�n�ɜ;D=���@_sf$ �R�|�#>���G�C��(�3�O� �J@J���?�b�J��֮ND��q��\�ց� ��P|Ŋ��	1A���U�]	
cay�Ϛ�!�a�|�Z9��Ƙ�y�!X�r�,��T�	�n�v�[��BG��y�@� ��f��ը!A
r��x#��Y�t��@)�)³_P�>)w�7#��=Z����S� <�A�
s�P�r ����A�vn͏^�nD�D�խ����]�j������ƕM�L����:��U��NL[�xl��+u�+M�?��`��RrZT!����� �V��˒j�놝���_ Zr�he9������X+l0�,��GX/b�|��h�$�����-�2K}��bv��<I���2�ɈKր�d��`�l�D��\�I�p �bt1:+]y3"���arP��,D$�	��B�7%<�#!��s(�Z���3? Qq3BS���E�'�3/�$!*$��kl�`{�D�Fs��b��FK<��vFO�s�F8`��D�Gw��MR��X�O@��(4��dmd`aO
�'��h �(ЌB�n$qֆF7���0"�IF��ȱ18���G�N˂j�=+�zӑm�W: ���K�'9���l�?/�j(�m�S2�#���:�|퐕!J�lm�K��F+��BV���[���f3R|��i�"K.e|��U�J8oj�c�ڙD.��j�Z� �q$J)n��
!Sْ�n_0�M�Q�
�m��Z�Lқ42��[��
�O������+�8�9�c?cg�4�A�@GТ"��a�%:��V=Ga�AD�ʠpu�@�Y�X����L?��M!dn�! ��'�l��ϓ��tJ�˻/�N �FK�~�*��@��$2\����LE m�L�wϒ8�ljJ9*�\�֡
�<�ЮY>��e�H��)8��ɑ��� `�[ӊ<�D�=�c� �P�	�s�����!�&	�0E
#M�䝈��~�u��J�$7�^��d/_�+���A��e�曫���s�#�?�,P��;3�ޘ���-�d�;�A$�!�h��n�`b��8$WP?�5���[�H�� C=t�:Y�S�߈a�h�$ ��6X�3���%8B���AT��`Å<p�.u��Ğ�e�b�	�O7��{��X�U�8�H�Cٸ��٘�i�|s3*�%js�׿��Cw�V32���F���-�-Otyc@��]��agEv"�aq.��4���v&x�����BaC@1�9�h��P!5�t��癷@x�� �N�c�=*��>@{�MCD�N
4�6�Q 5�`�S$g�5Gv��P�N��H��Ź��4� Ŝ���9@�a��zUZ����9H+	3@B y+%�ڭH���Ã�;�v�A��RC���I
70���m��GM;%�z�,MqFƖ9~Ҹ ��
6�����' �GD�q���,w�ўX�A�40`�Y ��n��1B�$<�,#�Gu¤�R`�XMP1�!�!f�|Pa�[���y�����I�wĴ��k�H˂H�m>U�v�@;s�v��[H!��(J<L[T��9q?t��e��i�����4a Ё3�Ǟ_N1��(>IQ@|{6 ]�"����A��[L(`GJ�S�.���O(���%�|��p�B�#��#>� �)A�yvJ��"BT�`�2ԓ�2m���''
*#D�8�B?\z1Æ)��zrN��b�
b�"�ӵ��O����f�u��G��3^i
��^kmN�Aۓ ���s#m��]��$���U*�5�H�Vڬ0�0�O*I�H�c�a��[!�(y��ʳ	T���ܴ|��'�"\�s,�n�HM���H!��	hfڡ��O��2M� �pkG �i��V�[4LjNx��Q_��3��#��A�ܴO]�!��T�#��"��I۴��'.���u�
� }�)Bz>�jaD�8�\fA�?G21�#8���{�pJT�ưҘO|�tRtG2V%ܜ`D%��P�e����$L�FI:!�B3DRRl�1���	,.A�d
T$1*<SE�?a���d�b.�[�O'�����g�M�ҥ16�>)����ݘf:��F&���m�"6�"�s̀-
���Y���0r1�l�p��Dj*ղ��ڜ'o�GC�zb(	����d�PH4ˑ)�8M�ŠpJ��ҵ�O* ���ФA�&A�dT@�g]&y��b�)�N�q��Ƅ_)D�BDɞ:~��}j�
M -�ēQ��ي��G5{Bޭ��ѣB<�+6��{lz\���]�=�j$�N0dH�����5xG΅�3� G6�Ę,zh(��W� ���I*��{��'�2H�X�A��,��p��)���ã�Ⱦb$�9��0x�IJ�H98R�ػ���v�~!Ч�%���Ӄe�?j6�iO>�f ��^=ll�d�L�T^2�"7
Q`��Z���Dh�n�D��� F�(���顪�Q�T	R䭁���2D�4����X9p��c�@�@�>i�l�v���'Yz%�p���l���.B�r|��3�֐�����+�6(��9Qn	��	^�|7�\�2���'�.&rp�1��=t6��フ[�hx 'e'�Ot|�Qg�2(*��w���TT��SX�K� �b�+{!��` �*9���
��3++�����P@���K�M�����1.@�Q�c��R��2
�')�ax"�ͫ�`�0@b�W�*i��k���*�pfd
q ��!Q�5I< s�bN:�x��/�
��p�>�H6R�r(�<�|�"_�+Dܐ�㨜%Œ�s��X:�����M�A7F�2s�N�+�ɘUw�����ph*=7C^��*��V����4��]A�`&l[�$E�:�LZhq�%�;<O4!��ꑫ^
%�F#�DQ����R�n���@��h9��!%]?H�$	�vJ�(T��#ۛB\���ĬSj��Be$��vU�80� ]%9O�*6�:�O�jdKF��{����V�T`�t@�6'cuɤ��w�LI�ŖN@Ts�fPJJ��g̀�R�@L�� �4#ee���(4X�q��ֱe��%r��y�axҪ�"��	#wo)2��k�-�w�]Cb74y��`UNH�Yk�A��' �|SSg�P�H�%F��~~�A{w�mX�И' "�c�_%l�~ɋ�JI't�	N��W�U;"�^Ȑ���ap\����-}�D�SB��8�hz�G�2��%�R	$���c���p����/�zU�񈉯�p=�7��uNd��SM�|%t0
�)�"{4$<j��*9B�t��BF!&��$�����pDv��y.` ����y2k��zݤ���B�,}x�����v�ўp+$�޷)�>������"�Ѕ/��)���D[�g���ӻI"n��,ʀ��-�Ve�ywv����?K¶<P�ߑh]�e�WG�|��5a�FK�:2AU�ޫm?pq��H��'i���3}�����C�P�⡚fC��y���Z1�ܶf�r�i \#oN8���G)�U#��t�)�f�R(�j�2�!�c�Q��e��/����V�1,����)��<	�eR��`p��J�[���(����VV29a�G�'"�����
t��C��H,v̳���?DE���M�=��TbF������	��Uء�NE��``�P�KC�U�QW	 \P��e� � u�d�^d�h�ĝZl�LYMHK�yȁ��%T^��U�� �e��%w|zD�D��?C����.���̉$�O����	ҿ?0��Ճ=�Tm�#	k�4�;A9�B	�s(Ն>7ޕ�ƨ�>:<��ӈT�;�JY��c�m���3�r�H�ӽiuڤ��(��(�1	��A�.��'͊�M�4;�jh�OoT�9�K��fy����G[�J:����f� ������4z���d�)d�-!�(4&d#ڞO1�ͩ&��'R��S��=�hP���5��{e��8��������j��>dZ����-M=�n 0(M# <��Kv�_�=��b��K�gH*q��/�@�V�#��ϫc���;��{�ޑ����}�X "g�^"btN��=ak,M+�F��;�>��4O�?�D�3vF7%c̸�̂;H���s�E<bj(yK2��>�,���X!;�F�+��vypB �0i�[���$�֜ˌy2��0'�¬��+�>"�����1G s���8M�*��)3L�u���:��`���]�ְjs���n�h���m5�j4�O�+6I�a�v�>��x��gޑ+�D_�Q9�:s�|��E81@�Q����&�.�+OǮi*F�k�ߒR�ӹx=rE#�b�'�h b�딚M;̬��(�U��8EgǡP�F�ᤣ�Oޕu��	Uy`4Z5��H1ތ����y��Zg�����?l.�l�h�یP����Z�ɳfB�l�z���-Xc��a%��k$�d��V�َX��A�P���R�F 8������0���E�=+�t0�)�j^t��yihYd�Iî
<X���d�/Y"�L��=-@��+c���!L��ʵ�:|ɨ��˘<1���3���,^ ���wl���C��	�%K��;�BC�~������D1C�pW��X�X>��k7BB7}������5^˒-�5#�:q.2�)#���l㖕2É/lU2Ȣ M�0�\��0�>Њ�eB��X�I��̶h圙2�ɂ/mT0̲0�����wD�I��*ע��ga@pCJ�y�`L&�6�j!͚�{�p�DE��%>	̻<U,�p���� d�; ��܃ÅS(N�e��Q)D�K�N�<T(�@��~��P�xAN0�����yi���"GP��ÀGIQ����i�& b4%J�|zuL ��Jĉ�.��FR���`�ș2���*k|	��C�$xp��h�/�_��i�2Ɩ�x:L@���d	I��x���߸��dyAȄ��d!vc�D���!���^�ypHΔf?
�X�Z��p���@u�(��G#T��ĸ���
WF����ДUEB|�HZ�M�%z����,qh�T)��G�m{"a[Ր&�Av�2`�u[� ���T)��<I��n�8�%Ėj��	Z�LXd�O��X�'�I��@�"aю0 p-h�{�G��Hg�>�nDF���7Lϖ ����ap�%��!Co��A�0�MKLN8%�4�>�O�d���4&q��äUk�Y��'l6\SB��<M��Z��(���G�? ���)�n��3$�(Uf��g%9q�0%yq�ֺ?B���$غx{�qBR�hOb�eR:D0�/9LM@!HSm��#��z�aD=<$����kJ�AXT���&�>��=���m���Ad�|-(q,B��yc��Q/y#~�1"O؍C�(״aA(-�Q�Ɓ`d�c�	�:t܅K��z��r-Ҍ8*�|#�B�=`�C�ɟQ��I��X&��凒<X��C�If���S��W*���uÑ7}�C䉩x��a�)͛;��x;�g	
�C�D��0a�]@zd�`�D8&��B�4!k��y�*�--��#A��U��B�ɊQ�TP7��+-���E.��wN�C�I<k;�����V8L�@A��	3�6B�V��;ei�.ņ��$���=�C�	U������J�d��|T���'|�B�I
���3�)S�}ٸ����(o�LB��5ZF��q�M#}�TP��"�<F��B��2�f�_'|��P'/ֲV��B�ɰM�n�#�/SK���O�1K�jB�	&[�Z��u�٥.o�h:�Jؐ
όB�I�8�e1�OO@I���򮝹j?�B�]o�2�d���5�T#A�~B䉆J8�1�\�H�p�Z��
C�I�F� �b��1�R��GB�^^XC�I
kT"����ór�b�K����C�I�.���b���-�xX�G§\��B�ɾz���cab��^�EJs�W`pRB�ɒ0�t��S0����#0�VB�ɢ]D��w�	K�!�HN�`B���ܤ����FiР+� FhB�I�}J�# j�ؼ���#.�^��W����Ha�gb�>���ŚzD� 'U�(Q@D*˧[MR�r���8�tZ-Ol1A1��0|�R�!�@DZFBJ�%B�! ��R(M��I�)��!��&K�Q?��K�Y]�jɄ�0��!��n�T���H'��q�,�l�)�'F��ak6��"s'4�)E �:�6ec�	]6fRh):gb3���:�~2��߈R~���THg]���˗�SY�'ϸH��s���h�e���h�K��y-�EO6�$��Nľ�b>��!N�X�$QJ��u\���7}�ȵH����y��^�JZ��s@%�!z�ȩ�Ҡ��<i���ȓ!Tf�j�VF	������d��g_���d��2�-"�M�e4�݇�J^�a"hL�bU�C�[^�(�ȓ=�8q�e��i��i�7/��;��U��`XP��cNƏ&}�-� �Z5(
�Ԇȓ設S ���.4a�-E����ȓ5�F��+�:��q&�Χ?�\�ȓD톄0�G�p�sF)F!q"����1��Ɉ�ɘ�Y�лi�8�x��E��ˢ-N;P/p)�e��=^6��ȓyN���D"�2:�dA���=x�h���g�L��ՅN'��5���*�1�ȓrXz� �A�J-@i`�*_�,`��_�");���Nئ\����:�8X�ȓI��:R�F�P<�䋑��#k��ąȓ^6%	M�?a�%��A��)��cd����ۃQ�@X���Y9�2��ȓn��K%���
����(*x�ȓY.\��$R�%y��ʀ���xPb��
ޝ
��}kj�
}�I��{�M��K�JL�R����Z���v�%��.�81B4��J̤oY�D�ȓg;z��� 7f&�J�I���Ї�s�����L�s�����W��݄�Ll`;E	�-�����Wb�U��S�? 6��f�5W�Z�{� Z+4(4ؙ "ODq����24�-t�W�K���H�"O�(��_�&��X0�´`����q"Op�K����P����a�����"O��(���k�8`�� h����@"O����2��q�f�ȝ)����"O2�K�G�D�9���έJs<P""O�|R#�ܬO�F-�.8e\m�3"O"���$��B��4���"O�� W�m�6 pn
�TЂ�"OP�2��>0�|�d _o}2Uɐ"O
zDХBi�� ő�4c��"O-#2�'e�Z8���	�yct��"O�q��AW�cU�� �o@PKV�С"OҠ3h��'�`���$]�d/܀��"O��J���&�h�s䂌x�X#3"O@�u�� [@I����>��U��"O�suoL���$�橗g��yU"O�s7aA�Z'R�A4K��3���p"O4]�.�/w�+I��7n�10�"OR�3F��1&IP�b��@�[WY�w"O��Q���0W�qpG�^"!���b�"OT�q�@ԙf�0�kkZ��"O,+P�ڝS 
��4-%&6]Q"O\�2�Q5H�P�Q"x0�"O�԰��G�R#.��fL�_ܪ��"O��B@-K�/���q��'3��9"O�A��J7O>.�Z��J=��u+V"O }0⥙2<cd<���Wm�diu"O%�fZ�K5P�t�̍b�����"O$�@�B0[R4�q��/h�>��"O��BU�дkY�@�E�ٙ8Ҹ$!�"O.���dՒIj��a
�D"O��vF��.�1�c%tq�$:0"ONĲ�	�L"���b�1J7�h�"O��ۑB)�ژr�a�( ,`�"O = ��D�!9p��d���8R͐R"O�y
 n�2&�{��X�f�qAS"Or(�$ѪY��`1A"��z!�M��"O��X�ț�M�\�$�
/lh"O4�s!I+	:��!�AH�0��{�"O�$(��_ >��݊�S'�X�r%"ONY�d�&c���k��oF�2�"O�8��)�1t�\x�5%H�M^�W"O�ք(��rǦT�`!0k%"Ov�S%�p�M���4#h��"O$���^�)���P�A��"O}{��m�z���ؾv�P5	7"O
���E9j���&�) n�p"O �s�Qd�f��P$D	�	!"O�]Sv�9�������-Ԑ�Y�"OD���VM V��q�C4�n�I4"O-0DIF�n�����=,���{�"O"����0	0v'<@�Hr"O4{e���t��=bW���@��j�"On0�PLθ!٤�X�'�/zr�+"OP�@�ؠ"f��TH�Z��"O�p8#�ٛ3�  ��o"�`I2B"O�9��vC&�{��E
#��ٚ "O�Lq����M��`���9|�[�"O�Z��?Jx���O�����`�h�{��N#G�����E��
�H��my����1z������$%�Ć�|�*�p�	��,t��f�]q" ��S�? ���<}&59���1�xHi�"Oz!��ܤK�v���m�?�B$�V"OXu��b���b�+R�U_�q1d"O��Xb)סr��pza��
vE\@��"O,� (T>u$t�A�bI��9"O(�� H�m�P=0�A�946d3�"O6y۳�G�}�@����v(�D��"O���@�d���Kb��#��"O�d�����<P�pvK�D��2"Oh�h��\:/���W�?�}��"Ot����:7t����B /ٸ��"O�ݪ!������*� k@͙@"OH�YR�:"_��5ώ�G
�4#"O:�#@�=�H��0�C)g�eXG"O�@��*m�]c��(��H�"O�d@��������dB������"O�����8�xH�'�E�JK���"O�!"�m�4LS�4�wl��"G�4Kb"O謁s&H�?]"���76J��T"O����Q)Y�Rhk���G2���F"OT�˧,ӴX�� #�X q0��K&"O\X�*�A%�X9��!l�y2"OZi�j�!&���kЄP�^�t&"O�I��N��d�S$Ӽk���"O���A�?_�2H#��ػ�*�2�"OD�3�I���Y���-_pr<��"O"и��éQv�E�E�Ik$a1"OphY�G_�w�J�+��� Xr��h�"O��k2�8��laS�""^�aI"O�㑈�""B��豊 YBRmS�"O�����	]`�E��,�"OR�X��b>~	;��C=Ny�ar"O��$�Na���� �  !T�]��"O4�1$M�޼x�a�-V:	�G"OH��u�Ue�^�8Fc^�L�ʦ"O0(����4(sD��8>;T��"O2��q"�'�����f��7�$�"O���6l.@��1�$�1/ -Qq"OyX�.ޓq��t�P�G�	zI��"OJ,�g�.%��QV
�%�"Oh;��ɳ]���F�Q�0�0�"O�(����s�8��� }�d9�"OPD��mX�c ���ƈ?�v���"Oz��j�%0���*�����%"OVSDؿrP<e:�Z%q�"O֐!4m�9Y��xb&bK"�.��"ON��go+T�4�6`����&"O��J̞n��`��!�06�~!�"O��AP&�ua3��,%�V"O"�p7�@���΃4q�p���"O6�j�GT1tĨ7�+D���p"Oht��M9T<n�XW�8{]d�"O���"��R��U�D0Z>�D"O6���g��]bZMr�"؅EG�i�"O~�VJ�����ͪJՄ��"O�� ����@�9Ҁūe���!"O�Zb�Y�~�8�CF�����v"OxA�5�ϦM�`�W[?~�
s"Ol]���=qJ�I���p��q�"OTU��сr��5�e�,|�8s"O~h�փ��s������N$�R"ONl{҃��}Q�N���1��"O���4+M0y� M�O�{ꄁ"On�H3bå_�@5�Fg�&�zI�s"O� ���a T>�(]F�F-Lg�DЂ"O�mucR�N3���dD�3ZL@"OR��.ӑ,���B��/�Nt��"O0���,@ ���k<��	V"OZ��T]�2(J1�°I��b�"Ot���N�I]̠�"��/��4P"O�Ya�䝡%�p+���
Ni�YQ"O��T�I#@�q2�6dd�)F"O]0%*̑A�9�aE�B��8(2"O.�{5�Z��T��fĠY�4�:g"O�|1�jv�[�&^�P��u+s"O&��E
��'"��`��&_���r"O��k&'BO�v�$���e"O*�h �R�E��q��!%��,U"O�5��Ϛ3�VL�� d�����"O�囒�Fv�@Sj����"O���4bٺ1��@_'��B"O�H��Ppy�`bC&2�ڠ-�y� �d��š��م!�s�n�r�'}�+ƎS����5�̠�(��'�ȸ)'%��Z�����M��i��,#�'��9� �&Sະ{�N4a��Q{�'�"yǥ	2����C�\����']]����V�����%� V���R�'�� ���ѲQ�� �C�:~���'۸x'��<�L�ccE�/Jn���'���!m�v���N�(��s�'��U�(��FpVE�R�Ѷv*N �
�'Qb�9��|t�"�ى���
�'��D3��Üxld�u┨d:Z�S�'t(8W��2ڴ$�3rN,��'զ�G��KgBd;/�!*�pA �'^�ؕOE[5���cܭ!�ؕ��'(DB��[c�hZfB�/M�<`��'�ʝ"�̋�E(j���P�����'�@$�!L�!&4���w��3	��2�':���$��?(zL������R�'AH
 ӤMS �9f$��|���'�zF��lt�0�Ą��t�����'Ɋ�C��1'Q�9�D��l]6e�'�4�s���=~J�C��$HZ�'~(�)s��%ErP[c���`��c�'x2�Q� �"�I�O�<[�����'p�Pd�5-�T��u#�(M��U!�'�$eكK�} ���᧐�p�u��'�"�J�)�WˎU��D��HX��'ְ���n�/2�.��"�W>/���'9l�S�@���)U�Ђ�L���'~�P�R��\uڥ�Ɖ��6�@�'���B�dI0s���;w䙽�(��'������B*D���E+O��q��'��0����<�����Aiz�"�'贡�H�j�����8&�$�	�'J21��]�.e� �s�W�.0��	�'>��J�A�Ug䀊 	Љ �>���'�{ע�z���;�O�nY��'jv`HSI������`�T���'iph���Ք5B68s׍��U��89�'f���Eߍ @0�Ɔ��9��Y�'�� ��Ǭ\��p���ҐG�:Y
�'��i�  ���   �  �  �  '  j*  �5  0A  �L  "X  hc  �m  6t  '  ��  ֍  2�  t�  ��  ��  t�  �  T�  ��  �  V�  ��  ��  )�  l�  ��  ��  =�  �  �	 F : ]! ^)  1 n7 �= �C �D  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr�	p>!��L�>P^�x�#\`yq�~�tD{���O(dG6â�ߘ<����F�N�B6��~�'.>I��]�(��d_�R>`��	&D��3$l��� ��'y��T"`/"�	�|az�H?X̴Y��ǘ^�B| �e �x�@�?	hlHG �*&���ɵ@�<A&��H�'�T)r��u����`��/T�i�'�S�č��F�P�+ 8x20��ĺ�y��Y8#N�P��1�P	�BL��'�)�s�Y�1~"AۇlX<�XAL<��8h�B��.z��s��N�@�}�'fvM$��E�d^� jSG�>l%��ρY7H03�,D�������b�]S�lZ�r�̹�'i��1�	��~=Xc@ѯMb����ėL��Մ��?�Ox��W���`�~�p�B��>eBV��H�Yw�^�]�*�x� �nN}��/!D�����^����b��WL����O�B���J�l�٧�QM�H�R�ϘB)&��$:��«z��u;!L��;-�Eaș!��5z�y���6G!���.Q��G{*��\�Ǭʓ��-W��S�ə�"O^���.ONA+F��6[� j���%|O0`� �B�v�ڍq�ڂ�x��i�ўʧ`.Z��y��V�k����=y����&j$�y���^9la��&^r�8Ql����)�O�yA�B��6-�Kd�+�j���yrj�8tE�Q���T�*�2����y� G�g�j)"q� �O>&ݚg��,�yb�D�#ˌa�E��^02}RgN���'|z#=%?�j�a�/>o��rw���b��}�S� D�DjF��$o�`t
�H��,�n��1�>��p<�R�� ��x�h�&RI�$��`�<)Ǡ]�S���C�g]wh(x�ԟ4*	�)�d�p篆%%Æa��*`��H��Es��:u��n+���ᑧ y���A�^89�`�<�0��%kwL1��9MV���&̟f��CƸǬ5�ȓ��q:��Ϭc����U�� ���԰�&]/+�d<sF��4�.��ȓ׀)��[�A���Ȕ!d�(U���Ҡ؄�P��3�ǶnO�B�I�'F!�6�@��$ZB*�!Q��B��7s���$�p��� !+ց?��B�IWL����C��sT� q� Եa�B�	�23���BK�8Uzuq1�S���C�)� j��Q/�9�1u�M�I��Xq4"O�����	_��K�	��7���"O��L kމ����-u��Z`�'A�p�<iڒA�Z��N@W���H�n�<�`kÌf(����B�"�j`�"��<Q왻Z���z�䛫b(h9`�@�v�<��4W�̅RQiQ2Ć�k��Ui�<yW!R#b�H%B�̟�`�.��M�<!@�s��@�B���$����L�<A�}��D���^F?�5�p�RK�<�3��-6�&�i&+��
��XGjAD�<��F�a�<:�B!|��aE��i�<��c]!ؼ,��&�06�ݱ��i�<10m���(C�I��8�	w/{�<�3n�'�$={a��;�\��3�	B�<a���zsҥ��F]5g��(i���v�<����~9zBd��W�.��!�o�<�擰a���N?W�t�e��f�<!4)��%9g��7iC���W�Z^�<Q7�'+�𛅏�6?:P��V�<Qt�t�T<Jb��Xd,�3"�k�<��a�?pY��Ht
�*T���Kt�Q�<Yv�H6�\xa P**�Hh#�n@T�<1�
ס�ΡS���)
ֆ�I�!�z�<AE���)4�1χ(U���p$_z�<iա@6��$�9V$0�q"�r�<Qt�]%L�4�2RF�]�jq�M�m�<�Se��\gX0���r�T$�6��p�<ɓ蝟Wp��2T�a��F�<ٖgE��(
@\��2G\�<ī�}ߖ�I�E�l�`�[PK�}�<�%��{�\t� ��>D��� w�<�c!H�Kھ|&�Up�!B�q%�C��CWx� �i���-���
�B�Lu�u�4�R�i��#Q.p�zB䉾^5k�)�T�p1�3L��>^B�	�U��a���=n(��3��i&B䉺k�����Īsx`y%o�'x��B䉦*I�ӁRZt��rD�<U5�B�I�Y�ș��#|�(
�� l�hB�	'���+ρ!AVy�N9}rhB�I5���۳Vm*�b�E~�B�I����U'Ѐh�^��-�B��_�Di:rcʸs�6DY�+T�O�C�ɩNQ$|2g��E��P�a�im�B�ɭQq����S�)���sE�9SzB�*�ع#́����;��â�NB�	&��
nLo��LXg�I2^B�	;����#�����e�KO�B�;i����55�R�Sd���xB�I�E+`�A��Z��h�'��C�I�q�Ґ����/~�Da#֬��0�rC�I-�H�(�ѾSJ�ҤJɂ$XrC�I	���w@�4�>0�BL�\�TC�ɚ@�B�� �� 1�I�K�)� B��T�@-�4OW?;7�ơCI�C䉄Bq�Abe"P�'&�	���	=fC�	3/&)9��]� (���Q�G�B�I;p�i�OӤ-�&��c��q�
C�I�4(��];y`�M`�/�8�B�I�o���3 �X�-"��G��C䉷s.`�B�S٦	9TΎ�8\B�Ie�θbu��:P0��'F7u�ZB䉃>Tb�"�ɏ%�P�āc6B�)� |��V'�4�H�P��-]�(U��"O^�3���h2j5�F��o�6hp"OL,�2��9<ct�AބM��A	�"O${)�+3�y��*��U�D8�"OJy���C�H�쨰1�
U��-��'���'�B�'��'���'���'�~�����|���ZW��tZ �'�R�'�R�'���'���'���'�jp�5*��I�x!�b�7<��'���'��'��'���'=B�'�xt �j	Amtp��@ИS8���'���'[��'��'3��'|��'���Eb֖_�x�b��ڠ-�b-Y�'[r�'TR�'���'��'���'UZ��)���pi�f�0,���'���'��'���'���'��'�\���A�SJ
hbB��,l��U�#�']��'�"�'���'b�'�2�'(�����{�f��D�;��'��'I��'��'���' ��'1�����^�p�l-X���}�Ty��'�"�' R�'fB�'y��'���'����F��
�1RN͏@�"+3�'pr�'���'TR�'2�'���'~&Y������ֿ�K"d'�'�b�'��'��'���'-��Y2c@6����P�y��tkS;5��'�b�'�"�'Z��'���'?�<�\-qD�ѕoSb�"&M3<W"�'���'��'���'�`6M�O,�J+"�I�F�]��9��L�I�*��'��T�b>�z����5H2�9+0�˩g%���R���J����O|0oy��|Γ�?)�&�$�<!ⱉíURȕ��Җ�?���{j���4��$j>a������<�N�IV၆"r-Q��F�.]�b�(�	ry��	p���w$̳+OH�����(3�@`�4^�,��<)��4�k��Ƒ:�.����®���Pg�ҡQh����O��I}���!�0��V<O� Y���>�<�2�%��B�� �5O��I��?!T@:��|J�{%> ��G(ƅZ3ƐC������D-����z!4扨-yx���'�[�p�h@�H�x�̍�?q�_����ޟ����D�2�T��#�	+!gZ���a��O^���!H����O9�?��g�O��È�^�	�#(��@t�pç�<Y,Ov��s����I�.|RL�<N��tb"Er���ݴGc(��'�b7�.�i>]�w�3iy��$jݵ=�����~�8�����	$vv�]o�D~�<�"!���_ۤ0 ��ʍ%.�aXW� O��8���'�T!��'6�i>��ǟ�����\�	�<�B�IԿ	����&З;��A�'�~6�F����$�OR�d�|���?9�B�,��òm,-h��VD�7M-�	Ɵ���w�i>��	��\8vƛ(J,p8�g�.�@���9��oZe~b�W5,"�h���?!6*��<	)O��*��{_�i�I��O�����O���O����O��D�<���i�V���'��鱓*	�{�N��':���kq�'��6�<���OD%�'�r�'�2�����f�:�f��Cd�_؉�B�i��O��M���s����߹K�S>�y��ʷYA�q���t�t�I����ԟ��ğ����Ń6A�䄃�eH�P݈I�UF��?9���?��i� ���_�,�ڴ��56��b�*ԴZ�I���0
w��AK>���?ͧ�(�ߴ������g$W�o��i��#g�1X$挞sD|�	�����O����O���^�L-��3��-t���� �O�V�1#E�l5�ʓN��ƈ@:��T�'���O�'��E��0��H	�hqDq@1	J�y��'��ꓙ?���OUR�Q#'�i2B��B���2�0Z�L�pFS#]���?1	f�'�t��I�4�	YW�MkoP#J="yx��m���h�	ßL�i>����8�'<7-.����	O�lu�EZ�{=���H�<����?),O��d�<)�Z�@��V"R� (��jW�N�����?�ԩ���M��'�����M���d	zo`��%śg.(�䭆KD�Ķ<��?Q���?���?a)��="#CU���D����\�T�C��I3��ߟ4��ɟ'?�I��Mϻd��ԩC�7v��Yxc�3[U<�J���?!O>�|*6Γ<�M��'o$�j4	E���(�pFV�tb-ڝ'�P�Q.�ӟ��P�|^��Sܟd8�nȉ@K����,ִ�,ږ�ß���ݟ4�	fyҠu���+�O8���O:d1�׿��Qb���	]��y*Ç"�������O����@���x����FBњ#l;?�4 �f���7瘝��'d��D��?1fO\�$�^���B��\H�c���?����?!��?َ�Ix>1C�
��7��}0��4C)V�J@+�O�n�}S�����<�4���y7d 7|-R��6oL�S���E�ɺ�y��'��'H��豰iU�i���	�?YÇK���HS�Ř|<��&�C��'x�	����I��t�I˟T��;4.X���']�:� W�ʳ":�'�,7���BT��$�O����b���<�'hԔ3<�"����Gla@�-��	�|�?�'�?���$z�M�m��U:FP�2�[�)M�Q���Dڜ�/O�4�dL��?Y6O�ON� !?O��M�R��m�4ga�x�3Naj����?���?���9q�=K*O<o�-y�d�S��� /N<'��}�B�eQ����M�O>���3��ן��	ߟ�!C%�L�� ]<>��� �e�	�el��<	�� ��JS�*��' �t��� ���g�#<Q(L3���=z�s8O|�D�O �d�O���O`�?Q�䬉�{D^Qk�f�8�R�9�䟤�I��|C�4���'�?y&�i��']�H����=?T:�	p�N�HR�|r�'��OQ��c�i��i�!�GI�!,⍹$@q������I�K�'��d����l���P]��07.ZU��uq��@�	ȟD�'C�7uD���O"���|27Cz5�8������@&&�T~¯�>A��?�O>�O�b�I�ˈ06�LRr�G5�İr�)�D~��p�@���4��89��I�L�Oz=����>���C�J�?P8��@��Ol�$�O����O1��˓D��v��m��QҦ���Ti����"�F��y�F�'���y�T⟐	�O���\��FTۥ�X�q�U��(��n��$�O�5�4�q�F�Ӻ�%����(�<ᷥK�
ͫ��A�]� ��FM�<�)Ot���O����O����O��'V�t�d��"�=�p��M�"ೡ�i��X;f�'b�'�Enzީ�uMS%'��Tcϯz��ɀ"�ڟT�	b�)�Ӣv_~�m�<�'��+cW�� d� N�ջD%�<9ve�
A>��P=�䓉�4���$��.���H�zc aQ������D�O����O���E.Q6:��8�I����8R� ؗ���K*�����	"��=�?�T����ߟ�$��x�g^1K�*���Y�r,"'�>)3�&VǞY F�x̧RƖ�D�8�?�!�����q%d��r�KlϦy���� ������D�O9ǂ�U95�5�;���2���\}�`uӦ�Yq��Od�DMƦ5�?�;���qJ��B�ͱVϗ ����?)��?q��1�M{�O��S���1�*"fҋX���P���8�$��f��)�$�O,��|���?	��?!�6�� 2� I��ƈS��6�\�*O~(n�Fmj���֟4�	@��.A>�a�c�����"�@́��80�T�d�	i��|����?)4�X�{ծG��>W���SFC 1pz|0UM����O�����k���O�ʓN�^8D!�, >��H��1p��?����?����|�.O*�n��u�d�I�y��@TM�z��9��J�7d���ܟD��sy��',��ӟ��iޡ��)"��5ȱ@��E����Yf@�B�iM��O����������<��'��R'pdF�&��|0t9���<	���?)���?����?�����V�P�pta˴V#t	��%�T�2�'2�r�$���:����զ]$������0��U9���f��7�4�	����'ߜ�e�iY����z����t~D�s�g���կ&���V�oy����#�Fpr��_2�ܭ�-N�u����4\�$(:��?���i[�=J0z�C�@Ж$���:��� ���O6��$��?A9��
?p������+N�a���#����0a�3\6�����Jş�h��|rE��-B��`B�%H��4đ�)��'oR�'Y���[��1۴?�N����3;R�Â�W.O��!��N�?���'�����
n}r�'Q�is+��t��ܸV�ŧP�,��'�ҏ;Y`�Ɛ��ʣ'�12�T�~
eY�zl�S�Y� ������<�/Od���O�$�O��d�Ot˧��X)��N�&��E�W�L-wٲ�(`�i}6�ۂV���	�?��HK۟���)�M�;Bs8$��ۃH��X��͑!v`L ��?�L>�'�?I�i����4�yb�32�9��Ȝ�@�<X�b����y������������O����3"P4Q�hĶ����B>�T�d�O\��O ʓa��b�b��'!M�^ަ���V"H��5/&��O�y�'^��'@�'f�f� [�� z�`��D!��O�q��E�{	6M/��	j����O4)x��\�V�TX�A�3R �"OTa�爑SBQ�PK3�zM@ ��O��	�0Ժ���Ob]o�\�Ӽ@�S�S��d#ׇ0	��q[���<9��?���#�� �4��$�2]��)��O�����iV�=��%C�Q<tJB�'d��y\�����?]�	���	��;�b\�h,M�0�ڏ`�&q�5�nyrBg�~a�&)�<�����I�Op��Y	�.g#�;�x�x���crʓ�?������|B��?�,ǵk��m[��#T�]��P%1�h9q�4���W�U����'*�'m�	
I�JQ�E���o��\@CҊ/�����Ɵ���џ��i>	�'r�6E�gAX��M�$	ri�T*�8[�^19G�T^��$U����?��]���IYy2� (} Y�r`�
RT*i�-,U�!��i��I��$)P�OS�<%?�]K������nb��i�:7"4�	^��  �g�63NQ�w�2y�V�;A�M����	Ɵ����'�����|BhW�M:���Óed�Ԋ��/6��'����4(ş}��v����h�w?��s2�&+�|��AY��x��O�O��?���?i��L�>�ʣ͔:bZ�av ҃G��1��?�)Ov)n��@A�	͟ �	b��5\	ئ�.+�>A�t�5��$x}r�'��|ʟX���Q�b�N��gT(Y����u�E����:wi߸}��i>�%�'�6�&����{� ��Sa�-\"��,W�t�I͟���b>m�'հ6��o�
10w�X2=HI��a�V�\c���O��$SǦ��?$Q���ɧ�M��CK�Z��,#���//� ���şpV&���'���҉��?���� �=)��A�72��#�O�����G8Oʓ�?���?��?�����	I?$=&����	/�MS���)��DoڣPF�a�'U����'C�6=��g
+/ 0Q"��2ު!薇�O0�D ��IލU��6�z�x g�+m5H��C�zV�9c��i������O����a�Qyb�'��]������~������>HFr�'���%���0�M�������?!��
{���%�?�|����?�/O���Y}r�'�O����� .�����3fϲ�1s<O6����V�F�ԌQ�Z���S<Y bFM���!宊�x%���E�ڵ��;��^Οp��ɟ����E���'��[��/�.5�aیr�AR�'uF7��+|�4�Y����4�h� +{�!BK�q�x�1OR���O��$?O�6�#?���Z;��)�� 
LH(V�M�A���b�J�,!�H�H>y-O���O8���O��D�O�����e`n]�q�]:�H���'�<��i�f��t�'d��'��Oerb�Y���҅K��O�<h�o�2<X��?�����ŞF�h�r���+�� �R�>!�Z������MS�O����^��~r�|_��re�N<�.py������N�����ӟ�	��Hy2�d�`�Ѵ��O,��gbQ�_zxh�γ1}H�aŢ�O6�n�M�@��	���'e��PR�ڗbȴ�bP�8� ���A0=�Ƙ�@ ,ϛo ��%�J���-��CJ�pb�����L<Se9[X�	ş(������Iğ���y��6�x6#ǯ�j$�@�˙�N��(O,����M�g>9����M{I>iR!�&y�
J�d��!޵�䓫?��|�Q�,�M#�O�T��玺�
��0gK� #�L�Q��D���#�'Z�'x�i>M�	�L�I���0PC�K� ��3d�y�a�	ǟ �'B����-�	ڟЕO� ���h�R]�����Б:�O� �'���'�ɧ���(w�2���F�.?����𯑷5�^�r����!$B7�Bgy�OU����P@Ԁ��/*c�i���'{��y��?����?��|���?�)O(�m�K��3/&u>��*f,Ђ
8���gf�ٟD����MH>��Y��	����)O?__�T���L3�ʌˤ�ٟ,���S�@o�<Q��>�	�?��'^~ V�Y;����q#I��9�'��͟��Iџ��I�	���Z{�a	�;I��(��']�7m;)1$���Ol�-�9O@�oz���n�f0�@�����x��k�ޟp��d�)�)%n��l��<�P��fcЅ��/1�[6��<q6FV�ZK���@8����d�O^�$���|�����^a"Q��,
�R�$��OX���O��^��)K<0���'b5S��� z_���E莕;b�O>��'c��'W�'	t2�%�^H�7�p8�]������ !7�|�rc>�	r�O�D�5-_$�3bo�,�:�z1�F�z!��ڠ<��X��ݰ@���+ɾDb����ş��7��O������?ͻ#�X����'?�xU�äz,�Γ�?���?1�cC-�M��OB�2)���d�<C���>V���AK֚B/�'��K�'R�ɋՂ� $\e��`�a��O �I�� ��OB�D$�ӝ�^h���Z�<��*ۭɶ���O~���Oj�O1��m��e��G��J��V�(�ޠ�0Јs��7�ky�ŕi�D�������$Ī���F���t��t-��@�`���O�d�Ond�3�r|�ʓ��i^�^%��>j���/��p��[��[1^b�m���D�<���Lg����0�'Ed8���Z�9ve�9J��(�7È$��f;O��$����X��<$����)���IF�s.�x%O�Q�r`��?I��?a��?a���O����F5["99s�ʇd	$�B�'���'��D߼��)��$��ѩO�c���8�d�W�Xɣ%��@�	�H�i>1�0��ѦY�' lt���B����O�c����d��g*���䓲�d�O��D�O��$J��������y!�G�=F ����OZ�Sڛ�Tl���'�rY>�Յݾ�©��֤b��)X*?��W�(�IΟ�'��  �|9�ӽ{�(�����dǂ� �ė�.�����A~�O,I�	��b���yR��M�=ZjI=vA.]��Z
96��'��'�ʟ��R0��<�"�i�M�EJ t,�Z(O΀���]��"�M;N>��'y�	Ο�Ò��p:pq��̊ �L���������Iw�vm��<a��|�Xt��?��'�j\���o�����Ə`���'��I����P�I��$��P����$1̵��� �����!2�7�� |Q�#���O��D�����O2��J��wΔz6O֖#���$ˊy��	��'sқ|�O��'h�P�5�i�����\�p�荒+x���PN��x��E
�� ���֓O���?��.��#�퍻O�=��D� A��?Y���?�,O0�oڈC����'Djȝ2 �����!�BT[�M �"��O�5�'@��'��'�Ʊ{���A�����K�O"���!�7�Ta�S�	F���O��FL�84��,��2��굉�O.�D�O�d�O��}���^dT�t�5���j֧�8!Y셊�W���\�Z��'��6�4�iޥ ���傑J +2h����q� �I����;M>nZt~2Ȋ<�i�g�? ��cr���.�� Jti�/$A� ��2�D�<����?����?���?�Ef֮:޾8y��%>V\I��\	��d즱���J۟��	ޟ0'?��I�w�`��EV+$@�`��
�,�O����O��O1��$;`�0/F�9�'�>��b�/F�Q�̈Q#h�<���>�H�� �䓒�䛣4�VD:�Ԭit��l�p{���?����?�'��D�릭R�J���c��E2���ʞ{`qP�e��0 ܴ��'듍?���?ٰh_1�hJ�C�	#-����eJ�um Q�ش��dK�>i((�	����:o"��*��ݳ�zX2w5O��D�O��D�O���O��?)"!� lt9��t+��; 'Kџ ��՟p �4^x`ͧ�?1��i�'ČuI��5j�y�V��
((|R�'��O�����iu�I1cs�9�͵J=��r�N�auJ8�a�ɠAc��6�$�<ͧ�?���?qQ�ڸ0�x�r�)M�9�6���?����$����agH�ԟ���\�O�h��$H���j����a�����ӭOn�D�O�O���yNp�@�_(bj�Q��^�DA��䄞mTU#� 3?ͧ5
��� &��e��ث��� $m���T�
�Ii�<����?����?)�Ş��ğ��q��$��"��ӑɌ��y�D�8 -�'�$6)�������OX�!��
2?Rx[f�S�l} ��ъ�OT��ƌ$f6:?Y��ďߞ�ryB�\q����܇#��۔u��d�<q���?���?Q���?�)�xM*�"���*�H� 5`���g�����$�埀�	۟�&?��ɞ�M�;P���a���QN�A�@��8~:���?9M>�|�5IE��M�'��m`F�8gL���
E�q�'ƈ�r����hQd�|�P��Ꟁ��"�j�f���B	I�:�Б��۟�����jC\Xy2,��`�aA���D�O�̐V䈅���o�`Z�W*�O���?	c\�����%�d��MȊ��x�g^����@Je���ɓ'%�jE ލ
�E�'M�������:��'v�!(���	�#�n	 ;�4A��'4�'�R�'c�>��I�p�NI`�C �x_T�14hRሐ��
�McQA�*��D�����?�;���?j}rd�7WI��̓�?q��?1f&��M��O�7]K��� =A�@<[S�	n���Xpkx�n�XN>Q(O��D�O��d�O��d�O]��lԵq������#��6�<1��id�\���'���'��O�үB+s�Ir%\RI�v��|�4��?I����Ş5<Dej��� rRPh�ca���x��f�8z�(�`-O
�2���?��<�d�<�(�3K�เ�E�͌ ��Ş��?���?���?�'���F���Qh�����D���r��C��|�Ta34N�̟`cش��'���?���?i��(2�!��i	���2M�>��)��4���������Ol�O��Fܷcr��礂�9���ӳ#A�y2�'|��'	��'A���U�y���ea̸��Ē���w�T���O��$O��h�Iv>9�	�M�K>)tEϵ:):�P�H��%~M��ia̓�?�*O��Z�yӮ�BW�\c�T�LX�B��.���l
�4D@�$լ�����O����O��d�)2� �E�I��<�f���*�����O�ʓF�v������'lBR>�h>z����b([4˪}D<?�wU�|�I��'������S�A<S��@�#IE�n��Y�q�+@�B��F�H/��4�*=3��&��Ox4uh��G�\Mi�̗�P��e9W.�OH�d�O�d�O1�F����ڪW�DqT�Z(0�(�s�ɭnl�s��'�Ҩ`ӄ�XR�OB�$�K�|@gK�pFN@Q��V�R���O�`��GkӦ�Ӻ�e��7��Ͽ<�$A��Mè��w�܄��u����<�,Ot�d�OH�d�O����O�˧>b�J���6x��:V�\� �iyj�ˀ�'V�')�OUr�q���<i�z��P�U�,�(�T��u�j���O\�O1�Dٺ�}��扨'9� ���ߐ),����ꖵ�l�I��Y���O>�O���?Y�0g��(��Q+\�J�V�����?	��?)OplZ}{|��ɟ���C��r�/PJ �b�)��.�ȴ�?i#U���	ʟ�&���F�4U�āѷ��q¨��B<?�/�`}���"G���'j��œ�?�3D�n��18�@	�J��S����?a��?q���?aI~�B[�|���$Z���'B����#�a>2M��Vg���T�>��'tb�'��I���7�ְ�AeX F���QI^0Di�	㟸�	��\����ϓ���L^5En�mM-+^! M4��U#���y*2�'�P�'�b�'=��'w2�'�b��\>zZ�j��QXT�KR��1�4=ތ����?����'�?!q��;Vn �R�;!?�)�v�ˏh������t�)�[Ov�p��� g%��*�[&kL�q�gP+7�"(�'C��0чޟ,�0�|�W��c�a!RO��B枥�������	������hyrhg�.��f�O~�dĜ9P.�Um�&f�*9�&7O�o�g��v�����T��ퟐ�r�XJ0����6d���{VnL3+�^%nZM~�ٲ1+�PF��w^\=�#μ3�Ԙ����JkBlj������(�	���	ğ���덺q�|�
���5�	ӱh)�?1���?��i�a(�O���h� �O���A�3;Iƌ������<(���*���O��4��Q�7&y�j�+��P� ��v���aWhUb��N�A�lp�͊��~ҟ|RU���	П���؟�*�&]	:C���3Ö�p�� �g��H��Ly�z�8��.�<�����^m�hjW��m���rW&Ǟq�ɸ��$�O���/��?��%搟b������iu/J�ZL��v �	��FA?	M>g/ �(�QDY�R�D|C��
��?���?q��?�|j,O�io�(c������4D�����BJ<�┥ΟH�I8�M���o�>���a$6��	��D����6�
H��?����M��Ond�Ǉ¼��O>�Y3���aT� �˟�V�
�'�������ܟ�IƟ�����ӽS|��oD6�Z�P��2J��4$j� ��?	����i�Ol�D�O�n�7�6C��5|�L�*rM�[A��d�O
�O�i�O��d�"R��7�}���# �2 ���C���(u�j�
b-g�,����$���6��<�'�?A"aG���%���ͣ|���A���?��?������������T��ٟ�"f M.h��W���J̾��j�o�\�I��	J��I�I+r�$�:�O
�n�j�V�I
U#S�M�d��4�Fg?�����<ː�\�����p\�	r���?����?��?�O5b�9E�'�K�2*v���q+��,�����z��$��yچ�<��iB�'(�w&&��dd@�D�0	�&ڳ�@j�'�R�'Y���]���3Ox�M�}	���'r�"44�H�ʩA�CX%v(ͣ�"���<ͧ�?y���?���?��̸E;� ��Dʆ١b��z����M;�eH�����O�"|�$�*M�0I �D�c��L�����D�O��i�ɧ�O1�9�BO'}��y�%i~���� �2}�\��O��(���?�t%2���<�Ջ"-�	�%H�i��\�(A��?q��?q���?ͧ��DW�+�V�@8`��"PN@��P@�}+2.�ğtz�4��'�@��?����?�"���;֦PQmB'?F�`,�:!��}8޴�����M��؟Ғ�����]�5{�-6�����!s���O4}����OH���O����O1�p����	 b� *p�T�S��MY�(�O����O.Uo92^I��П��Id�I/i���r�ߐTd��F�F�v��&���	������+C5o��<��^�8I9T�ڂY�r��C8��\xs,R�F��d:�����9O8�X&���[D4��c-��?u�M��ɿ�?��kП`�I��4�O$6 �U�� 4Flc6�ʞ8��O^��'wB�'7ɧ��UV�r�в�T�_�)p�Z# N^�`)Ίc46�Wly�O`T���k�܀��U�EF��UeF���EX��?����?Y�Ş��d���� E�r��jT�P$����%f8!�D���J�4��'�L��?y��4�����u���a.��?��X�F�!ڴ��dưPC<��Ot�	9�<Lb��ʬ+6�T�⡒=bz�,��L>턼Z�BJ %
iCg��/0��#�Ϧ?̴2c��3~BČ�SN�{��fC�x����4�z�@sA��v�$�ė<�P1Ѣ�A#:�#>i�O�5�P�a�h�"| 8�%ɏ:.M�X���8�~xbW��(J��xC�狊!� P!j�,`9p��ʈ0:e���G���G��iC����`�£Lh���T���8;��� Jr�jťːS)�)¢���\��ũX@�\a�b&dS�M�!zF0����T�j%�Ħ��ɟ���?՛�OD��Vc�	M�Zy`��F�:z�@�i<2�(`�'��'�3?��	�TH���@��]H��A�@պi�R�'��`\���d�O��	�\H���Ǣh%eHDJ�� ��}b��',I�')��'w�'Z�z�3�1-WK--��y�i��*[�-��ꓣ��Ox�Ok��lV� dED�l]t�)�@��	��3`t�l'���I����	qy"J�} &���	��$������m��M؇�>(O��d9���O��$�#ٖ��U/OZ؀��T<R� �[���O����O��ǂ�'>�^��h��M�Bu��c��$��(1C�i��柨%�h��柠��A�Y?�0��b �p'��yTtc�BG}�'JR�'�	
�f�#��"��-����-G|}��@&�	g8��n�ßh$����ß��$�R�	��a �T�a�,x��i���n�Ɵ���Ey��p��꧉?���bS�g�D�^�n9^IG [W���3�x�'��`E3{���|bן��hrI��W䩳gOƀ("�([�iL�`Wh
ٴ�?A��?1�')"�i��f��|&e�[�t�&��@eӮ�D�O�l
0�OȒO&�>�V�*X�AP�#T���(a�d�:�k6�����	���I�?Ѡ�O
�R������.�8�Qb	�+R ��i�x`z6�D(���Hh��>����ͅ�; ���'hٌ�M���?Y��c��)��]��'F��O���e�9���Ӆ=��ar�d���P�O����Ol�Ė�X�rh o��D���� ��{���mΟl��N����<�������p@߅T�nH�T
�pt�U���G}hʠCT�'�R�'uR]�	GZ��3K�7p�=��g%|6`��O�ʓ�?�O>q��?)"g� ��`�+�<Y,Ih��>�B�H>����?�����x��u�'"XK�=)�P���l�61-�~����?�H>����?�B� B}�A�C@�ِT��-�"q�p�ø����O���O��G�`���R?��I�CJ��;^�(�H0*�%�
�U�۴�?�J>���?1N�ĸ�� qe�T�d��K70�6@jǷi��'��ɹȈ�K|�����N��>����NЮQS��%�,�'\��'}��yZw$dYb��ĒC�ܸ 0���d��|۴���D�>4�(o���I�O��ITr~R%Ï|~$�CbL\$i���(�M�)O����Oa%>m%?7��Lz���Ŝ7v��0�*3��F�ü��6m�ON���O���NV�i>�`2MC|��8�"��U� ��P=�M����?�����S��'�b�7f��ш5��@�H����DE�6��O����O,���_�i>Y��k?q4D'2<�s�ؙT펙��iSڦ-�	F�ɭ�������a?Y��D=���Z;�]��$�ڦ}���{�T]�'��꧉�'�0�b�%b�@�㇛�p�p]�m'�$Ј$1Op�$�<��S�hm�SbN�e����c+״@:½���ɶ��$�O
��+�	�p���Z#팅y��l���T02�@lZ�'�Zb�l��Cy"�'*a��֟б��ǐ�	�(��"Ϛ��!�b�iir�'�O,�d�<a�����q�s�0w�dx���%�<�"�D�O���?y�����i�OZؙ!o�=�5�Ŋ��hJ������Ħi�?�����dP��'�Nx���(,`L`�v�1epvt�ش�?�����䚒u&lt&>���?��:'��1�ߦq���`���J�rO�˓�?1����<��*�������TRd�c҆!U���'�r+ܚ�R�'���'G�4Z��	��EKS$��y�|�Qb�5bY*6��O��oDR�DxJ|�s̖2gR�P�l�˨�z�,������,��ӟ����?՗��閲~���q��:yt��k�HE�3�x�'�(4X���I�On��7���<�>	�ã�Y�,����������8��t\�CO<�'�?���2θչ�"�=p�Z�Br�ƼT%d�k��i��'I�I ��)�|����~� �A�>�,Li�R%��۴�?IP,�����X�������ЊJwYD}3��ȁc$x�'�t�� ?)���?����䑎?��ݓ��^�/�j�c��:x���
}�	����H�IqyZw&^�BO7tC�-c��Ԇlm@�4�?�/O2���O���<��hD���i�#�`����> ����H�Q���韄�	����'�V>5�ɚK����U���dvb�#g���XUF�j�O~���O���?y�Q�����O�����V��8y�oڸi�Z�Qǫ
Ȧe�?����U�'���z���3!ײ��a�Ι�8��4�?�����kĈ��O�b�'��땧PX��UM��X�t@I��Ĩv���?	���?aa��<�N>��OVBB�޷ ����a՗�>�ڴ��ţ=���lZ� ������Ӂ����i* ��G�̸��D'�0ꢽi��'�ڔQ�'^�'�q���q@H ,�r$zJ�-�����i�X�
��q�d�d�O����0�'[�B��M��ۧa���Ǩ~!F��M��(��<�����:��ߟhE�����v�!x�$�A!��M+��?)��x�����X�ȕ'���O�8�1*�> n�(+O�m�`���i?�W�<peeo��'�?!����4`D�� T�r$�VpD�`�g�3�M���6�<�Y�Z��'�Y�S�w��a隭CW�J )�:e\	�'*@�'���'8B�'��X�dS���D�R��/;n4�R�G�l�  �Oh��?�(Oj���O���
�%��P�b��*,��N��)=��xw>O���?q���?�+O�S��E�|jUÄ�l�@Jք�`�d�'G����'��V����ԟ��ɰ����
e��������7,�� �ҍ�ߴ�?����?����ެc�X��O*"�Ǵ)1��ZFXҵ��^�d$�7�O�ʓ�?)���?-�����ܴ?��(���-O�(�l�;�oןL��By�&��b�v꧁?���C3m����GÆ�C�@�[�IƟ<�I��PZ�)s�x�Icy�Пle�V÷v�)��Iϝ��r�i���5#��Z�4�?���?y��"�i�U��"E�Dv�P��_C\H �d�R���O�2f<O����yb����J�@�C�/�5z��{���,s�F�K>z��7��O��$�O��	~}�T�����.d� Cݒ5�\�a���3�M{pJ��<a�����-����`�� )9�,H0e��;1���R��6�M#��?y����Z�H�'e�O$ͫ�@�#��℃ Q���i}�I͟D�%�~��'�?9���?��OȺ}�� v���6X�HӒ�B�^��F�'|^�9Vi�>�-O:�İ<����"�5��4��ˊ��T!���U[}"䗃�y�Z���ݟ���kyB����Ba��j�0��C������>Y(OX�D�<Q��?i�����f^ry�pk��z���Ҥ��</O����O<�$�<i!S�]N��ƀ)��-aP��8v�n$��	�yI��U�4�	Dy��'��'x8�R�'Y<A*
�7M!�qPr�P(W���r�{�B��O����OL˓|_�,yUX?��i��r���n��Hb�ju�
�Ѧ`tӸ��<����?���4͓��i�dQ�0��2)����ߗ7� ���4�?�����$K�_��]�Og��'��D���kj>��V�X\��yW��Hc�>!���?���
C����9O����o� ���ɃLa��QЬDn7�<��'�2~��'���';�ĩ�>��;�T�[�H�5`�h1�CϛV2�m�����u�l�	矤�'rq�� �A;�@��
��gG�CfD�
1�ifLͨG�pӄ���O@������'���/�f�e��0K]^�c8&�a�ܴo�&�ϓ�?/O�?��	�XF\� �^���K�-H�C* 8��4�?����?��bNz�	Ny��'%��̗�:(�L]�R��Т�*ߍPX��'���'~$�������Ot���O0�k�'�(s�n��U�J��KЦA���6��mɨO�ʓ�?A*O�������*�*�h��@���h��R�0��B}���	ܟ�	���Nyb���@X
.�C�><���BB�qg�>�,O����<���?)��k]{M(s��`%.�3n'��"��<)/O���Ov���<!����U����&<�(��cA�h���a�*��FQ����lyR�'��'a  ��'x$�R��E�����92$���`Ӯ���O��D�O�k zu �Z?��5$��	�+q�
Q�m3**��4�?�-O���O����_��$�|n�?r 8�F3h>*�Zw#Ly��6�O���<��L�M��͟��	�?�� ��7f��xE["�D�pB��)����O�$�Or=8�<OT��<!�O�`�Q�\�<!f9�gZtW��X�4���U�7�ޭoZ����	�\������t�w�����P�� �'�L`���i�B�'�R=c�'>�_���}�Ul�f��Փ�/Y�{$�A�R̦�X���M����?����zV_�ȗ'�01a	\<��%;E,�U��*a�!#W5O��ĥ<���t�'����+82L,��T<M��mr���p�D�O��DBa/F��'2��ܟ���j���H�+y��E�O�:P mnZ� �	���㒨l��'�?I��?)��k!ܽ��0k�.�ApDPk��v�'�I ��>�.OR���<����l�we�ݣ$,��P����a}BcW��y��'���'c"�'���(E��� M:��c� ����&� ��ē�?9�����?1�Kd@5�.)&�S$�V�3}< ("Y@��?����?�*O^}Y����|�d�uR)ISP�c�����n}��'�2�|��'�B�1u�D\>��͈�hܖ`F8a���-��	������'YX�Ғ�(�	��
��@3tPg%��~���irӘ�D$�d�O���F�i���5}�j�6��q	��S#kϔhP"���MK���?a,OT��[�ǟ��6L���,ĥ_9Vy�U�lw�II<����?ylN�<�L>��Ocbp8g��	V�9k�.�9��ش��d��^Ȍ�m������OV���\~A�,JD����L�>��p�[�M���?1獄�?AH>A���Ɯl���rLlR��C���M󵯚�OP���'���'�tf*�ɝlR���)o��}�&]�N#|���4F�Șϓ����O��@=�h��Q��'[��%`@D�=��6m�OH���O�q:�gY�I���\?)vM�/�H�(e�(Ʀha�.[Ҧ�$��X��x��?���?�1�I!Za��
���_��͸U�#u3��'�Ęp�4��O���*���Fp���06V�@aL�6���k�Q�X���g���'s��'�O�̥��C�*��ƈ��)"$@_5N�D�H<y��?�H>q���?�V剁ri�A��ܦ745�w� -}P �����O*���OT�����7���b̑ (�0 ��Ɉc(���W�T���X'�P���h��w�� �']��]!�����6�Z=��L�'P��'��U�|+���ħ�V�)�˜�t.u!J�_@�a�i��|��'��J0v!қ>��(շ��5H_�s]Z�ٴL��M����?)O)��(w�Sٟ�s�� eI�=0��D�AB�c0]0d�3��Fy��'��O뮜#6bAᘳ]< �0�	
��v�')"k�6��'B��'��DR���{���ӗ)�jl~ِ��|<:7��O0�K��DxJ|�%d[KFT���u�hbƞ�=9T@	8�M���?����BQU�(�O�z0Q���-!���ɓ�K��H�Gq���d7��䓺?�BK�#Y���zd̆�K�rtK4�P!��v�'��I:JѸ@�'��	� �<��ak��I�+�m���U:�I�ħ�?����?9�-� Ҡ��ě!I�N%�1- �{K�V�'��):X��[��6�2�$&Ύ��so��05���䇜,/b�'���f&0?���?������B�)[��b��-C��a ��)H-j�ӣ�Wn��T�I��?���k ,|��d@�d���1��I���<�<9��?	��?A�O
6pH�O3��ϸ�	��ҧ6i�[۴�?	��?yL>�����%f���L�o&E�T�CW�(�R�Y	��$�Od���OH�>jM|��oN�B��Α,|��<
3jZ?U��F�'Q�'�R�'ɾ-��}Rܔ$\��ZR��,axn�Y1Z��MC���?��O"��K)��O��iH#��e0oׄ8��HR�	�&��Iӟ����>���FU	Qߐ���b�lޙ7N��M#�O"1pG%|�е�O6��O���O��Ӆ��� ��c���] ޔm�������G�\#<���'IJ�Ur�B˳J�X���?р�߉�M����?������x�' (�3����xq1�
A.*����+hӚt;q�)�'�?	�A�#wMX�bq�A3��E*3����F�'-R�'E���1���OH����x���h*�DAb�X�M���o$�I�|�c�X�����I΀ ��T*�9R��'��&�hp��i�2�[�~�c���IG�i���=����Qm��:�u���>!�aWP̓�?����?��O��h�n<�<�Cv�Y�3�h�K]6�c�`�IA��ğd�I4}�l�ڧ�?
�}ӵ�W���%xf�8�I^���b�˚#F^�E�to���Xs1�^�()��"(ͱ�y�`�>S�&%H � �@�k�����'���S��ێ[汪����wW&( Ek�>������.͎$H�	��'�(�8�
@9l��mJ��ȹ����	!�a�DX%:�^�	2����i�S|Q�%BkGkH���wq(����'dc0�gV�m�A�Wй=��25i��=�m(S���P�e�3E�_��Z��7H��Ct�
 K6��rWʉ- ������?1d��C�@XrÌ	?&z�k���wYJ�S@���ۘLl"L�ԥKۈ�*�����	<|�d��V��'���شr>`�V��^���`��uĆ�l���P%1�>q���'��iIs�'h2��џ,Q�7r���!�
ʐNN袃 5D�����"�D��c��)m7 "3.O��FzB�n3DAb!jôOB<܃3��?���'E��'yb$8B-N��"�'~���y7�M�&�cuʚIhDc�T 3-�X��IN�bYn���/|y��3"�|�o�y�*}��2�y�q*�3y��l��ޜ���dR�#������L>ņ�x֢Kb�	O>L�'b��?�Or� ���4퉖=J���;8�AR�_>�\B�ɼ#�J� L��4"��4GJ�%đ��'����0��j��M�,
�d�Ʈ.Ey<Q+��+H�����OF���O��;�?!����DH��(��t����)F���pfʹ]����1F?>�\�k'�'lOF}I�/D�YgM��`�,jf4d��꒔,������܌?m:I��I>������jZ����*�$��O|�d9ړ��'�N !�,2{��`<S�<��	�'/��fͯ7���f��0��y��>�)O��
��]}��'[�А�πRZ��Q& R�	��!��'j"�!e��'a�	�h+N�S��^#/����F �h2�쉯GA2(�2�ý+����I&�̹��.F%�l,j�'@�9��F�C� ��kZ�n����Ǔ2Q���t�'��1n�� w�LP�D�$6UZ�ҋy��'
$�˳�d�fxa�0�*��'��7�K�u1 ���OSS堬�"�>V�$�<I�M��A5���'��\>�R��
ԟ�*���13G�p��o��z�ퟜ�I�  �9��4������#��WՂ�s"�͏��)�N!}� ��(y ��A�-]��s�-�D �e�J~��&mY��P��2�Y��B��Իecb�'�7m�O&�?$k�+�c���/1����kd��'��V����C�p8��M�'��9*�����p����޴�?���i��k[4<�óC_�?���у ��듌?q�IR ���?����?�׿k����5tV����E�直Q��S�A�>�5��

��1�|&�|�l�nຐ"t�^�:����,"���X���#���W�q��'�$���c�VY�E�R��p�U�'"�ɭq�N�4�,�=їm� �T���N;b� ���m�<�F�E�?�i@W`[�$��\hQ �h~rA?�S�$V��3U&X�K��AX�G�	/����i0���j`��ǟ��I��@�	:�u'�'0�;���2���6KK��k	_�GT:�jC+��U� �FB5�O�L�5��^���m�?#$-Â*ƠKq����&'�O���7Q!e��T�͕+��q�Vt�"�'���'��I����?B����\���F鼹P!nO�<�"�_!]ߘ5�e��
x�X@���P̓��uy'G�:ꓥ?a��\�a�b�1�}H$ʴ�?A�Z�9����?��O^�|�&��*W�I���>A�mZ#4�G')$ l�S�#O�1q7���l�\�h�u?QѭʳTS�����s�[�N�I8�P9���Ob�$�<�c��bъ��'(�����p~̓��=��HS�}�v��a盺u�����	v<�i��`���48�H�����3YT��*�'��	,ƞY�O����|"�I��?IgH^��8�-ڈ@(���-�?��y�dE!� �.�S���*���'y��Ce�_)І�_�ft�@�O���S�\�^�$����I�#}�ꎗN�xs�m]3W�(1CQc��f��'��>U�	�h�
	��	�~�R�ԧ���0�Ɠ�% ��E`�Q!�T������HO� 1�����Y%W�V5�)�ĦU���<�I�kgbAUm��I����	��u��*
Lر*O�7t]Y�S1O��8��'��,*G, ZF�T�S 4��{�-����<���XO$��e-�C[�����<ܘ'\����S�g�'����AI� ���\��C�)� P���C�ܠP�l��������Z����n}P�&�N����8���x-�$8��?v�h�Iݟ�IƟ�^wV��'"�H�gG�x(Wܢ���R	C�̂#OD��4�Q�J�t��TC�u�� V�	�0!�тJ�:��hۑC,�40g� ���y:��'&�';��'*�O�a�.	-��q���s�B�"O�@+W.H ��Ӂ�Ra�P`D�d�x}��i>y;�ϩ!�B J���7�VqZd/:D����Y��5ؑ�ӑH~l {�6D��x�@V�S<d�K��̄1�^�(1g:D��Y�	+
�]k�I�*@ST,9D�4c�oV$ @���C�h�ay��8D��0`�_(v~<5pA�6lܙ�s 6D�Hڔ	Z�4��0aߑ
��A��6D����,`<��I] `��!��(D������>g	 I�)��t��IU 'D�ț���4����Y�d�($D�\���G����9��\�����"D�\"��1$Iu2uDC"lD��b�l%D��!��M��Xi�'p�Y@V� D� 0Eb�>s 51#�*�$Y�d�9D�@a����#�|���T�l�H-���)D�p`��>�`�; m�U���[��2D�X�U�C�Dp�Q��M�f��͐��2D��ᄅƷ|�>��D�K� ]��Zrh6D�4 ��N�}�2	�H2��H�3D� *��h�Xd{���1Ί9u*2D�� ���;Z�Y����~U���0D��1��L�g�@] �IŤgXI�4�"D��ꅨI�M QTK�.Dm�Պ�"4D�l�sdōjnBa���o|,��k0D�,BQ�
r*��(���-����,D�|��
�/o4����`��� e*D�HK�)�T ]sF�R��إ�)D��t�Q�v�ֈA��D6.��e��&D� ����r��P�G����Ub�2D���IN[Ґ)�sJ�\�8`/D�(�0��E��#'�F���,x�(D��iӭ�=��3s��i~�4�4D����C1`($aE)"l�|Xx�#3D�(�do��B/����^.��3p�$D����N�;py�-��a��h��ms!�!D���u��!n����O� z��)SQ	 D�`
��V��a�p�!m"��;1E>D�D���Ä.jRģVc�'`v�ӧ=D����bB�4S��q�EL.1n��$?D����Yp�x��y���i�e
$�y' 7�yp��Q:p�����`C��y"�ӊ1�x�9����U��D��S?�y7 Q4�� �O�n�QR`��yB���N�n��S%�Tx<%����yR��#㮉*3�ղҽ32�U��yR��6Gnޭ���v6^���C��y2`̝W2�p�U�@"Œ� 啱�ybl<,!�,B�ۊk� �˵n�"�yB�E	1cx�� ��c���2&"ʅ�yBgQ�4�(�`�&ۑ\�]ؕ'K;�yҠ�.FJ|Z�M�O�\U	_��y(M�?l�t"���@�ɹ�(G��y�(Y&��9be��Ѝ$+��yr�R5 :��FA�C���x��G�y�b�&T�{�DĮ?dP�Wϣ�yb��o��aI��	�I�&e�!��;�yN$F�3�U#F� �R��y
� ���3�O�g�<k��G12@��"O~E:d$FZ���K�O� ��H�"O��Iah�����w�@41�HD��"O�(H�A�D!"��e��O��tQ`"O�X�W/�./$=����k�t��t"O��)�P5>�$T�O�7���q"O�1Ru�W(��!�md|e�"O����#�!��,�TcvPA�"O��(�J�U[XQ��D�z@��[�>A"l�D��Ho9��i�?��rv�<#�L�|�T���ϊuj�����-����s�OM�L����|h�b�\��4AԌۄ	�N�"~nZ*�D4@C'�p� 5��3��>1�HE�<$@1��4Ě�S��B�jU��:��)����+yrߓI�dX�K0P��� ��Y��`��[���Z�+��S��$�a�G�-�Y·���L��l(]"��yǬ=D�xK����p����@����zRF;}�@�L=2]qu��/�v5�FP����~�����
T�<���8�H�h��ҵ*ߑCXa�s�ص$�ک��-���U�ֈ�}/�|	f��_��,O��z�-(�s����V�\PU*¬V�r������	�f�(��Sb=:����A�E�A�=�X��Bم+r�X��ÊŗPJ.]�D�S8�xkR�
e�t5��-�;��{�A��&��aSrGGc?�OԱ�?��t��k��4jj��C�J&C R!����frh�������O J�$�#+˘ȣ%>�Zu��Ò	��5��Z����\�~����H3A�V���Sސ�g�$-�}�%�
?p�2�i[`�� kPcO���'h�!iTk_�J������S�4�S�O�8c%��j<�qe��Ǝ��F��!r�Ȍ��g'���:��QCn~+8�1�`-#��D��=��y#'k ��1�#�_$��g22�Ce� ��9��FB�0V�lt`d_ 	��H1]w �	:!��F1�2'�W5��h�'����a3m�RHrQ��V��8���U 2 "F�Ƅ)'T����1l$���)Ψ���)B�Ȱ+ L�H���VD�>Do6�8�H�h@ "�Ȏ<!ń�A�n#ړM��!!J%PH)�;<x|�f�J�+�F@;���?&���O�Af.D���C�p��c
A�g?�5�>|�z�#☗rH1jQ�i�$0Q�3�ɦ)u$1 U���}��x�%��V�.�C�� �Fϖ}@���H�(r�f�I��<,tlؕL̴�#�OX�ڴ#�t��hCb�,��C�'m v+��8,͉�Eɕv�ny���! 7���Ǌ��xޔ]kK<Q��Y�<)���=�~r`��F��k�'r��4��c��~rHM!xY����A�^��	9�J@���4�:�7&��2��C�Oֶ�	�E2>�NO,m�
ЛD<Н��@:�{�p�d-4�p��3��6�teH��VBA�
֝9k��<�ƽy��iAG漫n�';}� Y�$!�9Yp(T�
��y�I>Yr,\H�OK��I�������&��a#\!a�.,:�yb+L!.-8` �*�`@�`�И'�v	�f��&�L!�� -Εp�4!���ێ}2C�gl��ja�-h��i�t���';�MH��IC��(à��}Y�P�rظT,�52�g�Lz ۓmU��p7G�7J�	Ӗ@��?�t�JrF��pp�@��@B��;��G�sR��'��hI����<k4٩��%qaj0ZT#E��yb��'jgX�B�A�&����rE�%,6�|�r�E	$���!�+��'��#�k�\��w&�y�Vhγp�L����а5X�q��7���c�
�B5(�V"oX9��a�~��c�8��i�'>��*P�B hd"��%扶o�acA�� ��L3w��"'`,�>�B�
Rl�B� �3�,p΂�/��T���	,�v�V�(���ӧO(:����a�^p`�V�,LO�"׭��F3D�1Ea���;�']�9+�K?�v�*ufK�sM� ӭ���D�3A��_7Uj ���)��X���@���-d!��C�8�A�)#z��ʣe���na2@��:T�P�r"�ά8R1OP�p&�ތx�&yx�4�):��[+����X� �P��'�D��"��,�@���X�\�:�٤'�X�x��<٠/�5Ux��tT�j͎t�q��̓>ER-2��>A�|�wfA5U⼄D|үY�A�vԙ#�̵/{�-��B��P���Xd	��TҒ1�࣋{y�i;!jݕt�XI!%	#I��鳓/���?I�������x��) ��9�>hI$��s}���b� Vxx��'瓶2�@9��O��C�|̓�޹j�mY�/@@�ɖ��G��q���fX�T�?E���D5�H���@Q�2rHIVC�A�NUAE��)��)��i>咖���e�杞dG<{���.O1���C-Q|���[;<�B���� H����c��d���T�'�hi
�*6�'44�p��Dh�j-K�$"<�AS>�DU�8�h��Cl(�zT�a�?�T����D�Q�C��8LЎ���-҈��i� X����hD�0�GefI!��!L$����9`����̧^�� �L�0�L��V�{H�}��?��?�����Q��=`�g�n̪��DdD��@ 6ҼD��@y���1��� Ԕ}KR�{�� �7_i���<@b@L��)� �,I�dC&w�v�a�A��,�5@D�ɴe��m����0鑗��F�M�����6�U���csÂ�ÈB䉲F��ɰ��Y#L�0X`D��z�d��-vL`@��R�(�)#KI�)rd�}Zt�R�t�0t�g��Y�$I�v��}�<9���|Zd ����r�lX��ώ�1ʣM����H��		���fhSp�n��D��J���T�C.J�"��-�.Ȉ���v�h�H�D�O�f��6ᒬH��9c��Fi��t�e�5S�rlZ�/_4f2�ʀ� �\����6犉#�6�ۓ':s�Td��:X��]cTe���	�)d~��"O�aL;8�:ɘs�ўD6F8�`�i���b۠��s�/��Q�(�Af�(�k�\�����	lD�x�"��N!�5B�DEI�mҶTO��K��Li�
X!pGD��lI�,��4Ε�BT?��2�d;����G��҈Z���(�z��קt"0���Yl�Z�,N�tP��̊Z��#�.C�u��P��L^'%�έ�ߓF�q�ś0�^��
L�8���<��\�?��ݹe�
�}pP�7�P��O����J�/P�9sU��]@8XS�'6�d��%c�\p�uc��S�si�6�X0R���ȈL�����)�<���ǡ�)\T9��l�<3��4�s"O��6GU8[;@��t�3 � )�PG�9m{D��1ݙW�8T�L���2OE��㟼���S���qT�J�3���C�*LO�9�u-ù�⍣D�M�g]\�)#ɦmm�����[#n�+�����M�R.�<:7���ɺr�Hag��j[^�#%�b��+\��X%�ݠT��)���,.�p�� ȸ�u���=\tw��6!D�124%�+�y��G��X�%� [L������P�r�M_�5�I�͔�n�,�B�C䒟<�Z�w[�`6F��
�x�)a� �1��'?�dB�/�+�Bt��˛�/��"pI7�9�!%���͘%���<���Ѝ\A���ԓWo9�$�@��$!��ͫg�N1�'���	��W%+@Z ��������'f2 ����K>:���#ɂ9z���y�/Ѳx����a*@�OU�(�̈́_J˖C,���A�'t4�&��}��7M	/ Z�� PM^1���O4���3?i��]�J9.$Ar,؏d�� 0��v�<ၤ9f������ʀ̊�Ѧ~��� �`A�i>.���I�j��g���)�KX(eF�ի�n>&�P,� C���Z/�!���:"�����6B�5H�`�!�ս!�^=B�Ɣ3 Kb�<A�ʍD��Y���0v�E�	�.m��C�0B�B�	�,'1I#��.Ű�cr�EI�8����	�Tr�fR�PG��OPK`gԷG8�����E�,)�5�Q"O,䊒F��
o���+R�\+T�[Q�Z�H�t٩��U�p>ѳ������V����#C�j���k'�0.�~��vS����l�3jv�d�>W�!�S"O,ݳv�D���<0U!M!2�av�$U6A�bp�����&��a�B9Otҥ2���?R	��"O6Ti����v��'�
�s�:<(�g[�&�h%�<+��<�R�Άv�X\ '�O(P_�1�TFe�<�hQ�T�� ��K�!SU�5���i�<qp搼�yq�@�
%��w(Bi�<)B&[OP��O��$^<B�J�I�<)�N�S� "Ąu
(3e�z�<aeI�4��q�E߂=�0��*�o�<�5�ώ	�VM3�CQ�6)PX�g�\i�<��(P����B�:a��jš P�<�6*J�t@<��%�H�0�atv�<ٖ@!�29����1T���c	o�<�$�Y�9���c�,1%�q���`�<��#cI�1)�D�'=�r���)XY�<��Γ$�n��ώ�4���K&�S`�<ar�P��vd�� [�
�� 4�B�<	�M� kO��(��H�
�svc�@�<ѣ�P($�b��"aғD ���{�<9E�̑
�px�-Г6`�	!�,T^�<9��s~�/Y�:!��̈́��B䉝V����Ч)>�l��H�a��B�)� ��#`���Q��9�� @/%輪W"OF�S!@�FnJ�f�Ɔl��"O����e-�K�'�]��"Ob�2A�Y�]6z�
h��S���t"O����G^�C�,�tǍ wXR��`"O�@zj
j���¤8C�T��"O��Ұٟ2�Ƚ��C�;=�"O��!C�Wm6aR3C[<= ����"OdQ��-�'���qL��7/b�b�"O��Ђ�]�6,���E��bs
�J�"O�H����hQ2(Sԅ�䖪)�f"O�zҌԉ'����+-v�6��D"OB�S�$@�nH4��+�Z[��;#"O�����;n\%jĈQ�uf���"O`�D� ��ɣ�0K~|��`"O�R��09zBe8�G�S�*xj�"O���O&}�%�FeX()R���"O�����>T? ք�,
�v\�t"O��A��6��a"%�$����"OR�c�Se�,I��T�V�ll��"Oxp�kQ?^��Pp]}ڼ�y�"Or ;��U�e�%�߬|�\tP�"O"D0��eP��2��YƠ�S"Oݳe����<��o���z���"O�QC����
�x���D$f{�!�t"O|�5&��\W�!p#d��;��Ua"O��[�#n�~����:��lCe"O�P�J�d��P�R�_�\ �"O*�xX���*R<y&~ �"O�����W�쩃�hD�m>
��"O4�p�P2>]��3�}��I�"OR�!�lY�$۬�6��:�� �"O��񅫎�6~�i�!�D�6>q@B"OF��ń]�J���ɤ�J�&�܅��"O�hA���r_*��@ Px�� F"ORD�G/�<P>��� hZɛ�"OXHy� дHaO�4F�h�"O<�p %�$%ʹȑ�d\F�-��"O 偅���D�95��-�Up�'�!9�Q�W��!V�e�\x�'��\+��V�\І�VY	0���'7�5��FZ`�_.Tj|@
�'Q����e=3�H{PN�\�C
�'1L��5��r~�H`FB�[�����'N]P$た\�
0Ii�P��b�'��Ñ�F2|1gН1<�|�+O6���J�!�:�`��<dKUꛐR�!�A_��Ԉ�.�.������6,�!�$]�ty88��N;|����ʧ�!�d�4wYhIaD[7?>����3�!���L�d��4�C( �H�ek�]�!�dB�M� �
S<�Ы�* !���I��	�J��)+�(p�I�F=!��<R��u� H�l�=(3h�J!����q�6+#m�� ؠ䙏x!�$F"*�D�b����N�\i���Y2�!��bI8�IeL��N�l�Z�� �!��9��@0C)F�:� o�!�$��:�@�P"�_~5" ���O�!򤑂J�b��&+	�q�nP��Щ�!��R���!e�c�88JdGQ!M!���G@^M������(�H�*g�!�DD�E"��	�nzLtP�(�Y'!�D�P��5��ŉ�bg�Ⱥ��L!�� 0�ui�"z !��Ε�{>EI�"O�P�0���;3&H3V��.xul���"O�Ds��M�4�Z٨�N��ogT|��"OȘ��.H��|���,Ua:���"OLy����k01�`���DU�q��"O,-��"F<c��܈�d�>'�J�R"O����
)�1�c-R�9� H�@"O�]�k��i�~�ƍ��W�����"O�XQ���������R����"O8����J8t��
X�xz��D"O`��bO	S�t@U'"rfV�R"O��S�aL� 2�E�.xF�e�"O0`�Ǐ�.q]�rC
SH`=B�"O�\#0 ��:�*����E�>4���L���X�ue��jp&#��H����!�!�䗱8ɪ�c�.\p���1 	9!�$
�B&9���N�R�� �0e)!��;N=}���8@n2%R��O5U!�$O@y���(Z-_�arUa�8^��φ �|��ߩ~S�K��1�B��>ctY�흊4��M��"ȩ'Y�B䉒_>�[��P5%���@s(�q	�B�	%Q���F��	H�-��%-/�B䉣P��LEa��Kל%sՊ�q+dB�3;V�S4&��*LA$��PaC�ɳ$R��? �н�V�R�	��B�&P,K`�ťM(�!kŔ�x�B�	�c%`b%�=`z��rER�Qk�B�I�D�b0�@�T�2tȲ�L�{��B�	�
��xQ�l��"�
��J���HB�I5h�n����2r�AZ��_,r�C�ɻ�B��w��>,K�qQA�&�B�	�#���q�Ħo!���v�T6	�fB�4i��}0e�N7/�NI2��p1C�IMF� t/�W@:��4��,�B䉒(���C@ͨj��0z�_5w<>C�	�j���0~�Ĩ���mp�C�i�j"�C�B���a����"Ї�O�&�3Ɗ;}�@���"�'}�ȓ�LBT�ڽ\��c�(��(fLB�ɏ<��U"�o��{���b!Ϗ�!-lB�I9GN̬8td]�h�	é41��B䉨�f���Y�+�1q@�B$GT�=�
Ó&�m��nПK̸t
�ʌ�vR0�ȓE_p��4�d	�*%�C�	�g� �r+��n��T��nl��8�I ep���ԽbW����#7��B�d��b�K�"m���P-7`.B䉲����w�ɝ>��"�� �Pa���E{J?�C�m�w��*4�]���%3��&D�8���G�mʠ�'�6y�)Q�M%D�,h���(��E@pJ׌:1~MV�&D�@�U* ������2!�09�+�>.O"�=%>�bc%���)I�酴J�8��Ĥ �O��|�,e��[�m���H��L l4��9oT5�W�1c��Z�U"u4݅�2���tI�q-�8(ק��( 9�ȓF���{��+���i_�h��чȓ�x-AAH��YK���.U�s�z-��U}֘)"��?@��Af��%y����H� 	 �,�-9}L�k&*��	F8��s������a��\s �./
���	I��!0�
={��58 !��X�C�ɺ$Ӣ�r�D�|Ҭ<��n��!�� �l��K!uG�T(�+эZ�l-��"O�j扂�qZ���L�_�2�K'"Oh�a�ʨpP�)�K��_Z1yf"O �p���%b`�,0*R��ku"O�@��ŕW�laz�!�0(ЈC"O֌��ѓ^퀍K�Fղ"� �"O��Xq�# w���ħ�Ȕh"O�)!�.��0��`PC#�� �"O�`��h�J@��
#-��w�L���"OV,�v���|1�L��&!a6"O�1`"���Mf�H P,��9���۰"O�0K�N�9`�v����!p�X�x�"O
�)�`�Ahi@lB>5��S"Oz�p&9��tJ%�YS���X"OL1���/ I�%Y��Y�B���"O�A�g�m0<���dt�|��"O��* MЂ�>�!@� 9쥢�"O�hXS�D1rO���S��a�x�b"O�
P؛��c#��T����"O��٠�"̬Y����R�F��'_^���`;&Uh�L �xҪ��
�'�����ϗ5��� ��2~�p��
�'�0��e@ MP-����tj��	�'��ɹ�A#�`���h9����':�%*�!�g.�:�@�6�q�O����T����j�	q����C��h!�3�TE#'LH4	���a�;ng!��_�/|���.ې<��]�&��:0!�Dӡp}[a��NHtay��L4K!�T=LMYԏ��<H�	kE�O�!�^�0�8e#K,N<�M2d���!�$�:�����k�H�0�07�B�K�!�d�<됉p0I4���R��ĸ��yR�]� ��r�C�}��%��ğl�<�v �	��ɐ��?.��a)�H�`�<)�C]M6�Z0'�$Jy�Q���N_�<��!l��V샫c���0Q)_Z�<��ș#T��q�b�}`b��]U�<!W�t�ZAAg��&e��|ȅ��V�<�%�\�m�"M�@�K�g^���'�U�<qs��#k��#(G�W�&5b��]�<�RK��"�^A�QB�n�V$jD�[�<�5��q�X��5���?�X��M�<F�J�!4 �G�H St0a�GEH�<Q� 7��@�wc��T��Q o�@�<�7�$���ǙQ����a@�hF�C䉸K�����W�>�v(R�S��y��+&���M(l��(�y���K3�(���J�XI��c�.�y���������$�=R�4��	=�y� �0#�
�as�ة����T��y�K[�YL�"�<L�谦)Y�y��b��ܪ����U0F���y�gZ&�=�惚�D���c/�y&�-j��z��z�L8!��В�yR�аh�Z�������^2�y"��LR��ǎ��<���c�V��y.�9Q�7K�:.�^�[F�ҹ�y2�������a���"�Ҹ��G��y"�Ľ&�H��$lC��zE2aHS�y�f��/H�`���M�ژ ġ.�y�I�/FZ �w�N$\ږ%Rd"�y�	�l��S��_f�֌C�y�L\��"���WZ*�+�$N/�y
� rPaա�=X���z�
?�Ҁ"�"Oҭ�4,ƞ8����C�l�.�"O(-��Z�l��+6��G+�XiC"O�h#��~�:V�S�<x�`�"O�Y�qmQ�,=B@�IY�fe|U�"O��!@+�2.�)�I�ad�{u"OP�(g�]!P1`u*C@&<8=Ȕ"OT� !��S�p� s"ȵNr�("Ob��+ۋ&٨E��+�$]騬��"O| ��BCw��@�N2	����"O��Qi�)�h;���y;>���"OΩX�P�;�8R�M0�U��"O�u�BQ7a�u�K"U�*b"O��B�[��}�R �-Z Z�"Ovu)�K��E�j@a�m!(l�у"O&��f"��L�LH�ČNx��"�"OL���,� Z]<�1�lG�E�5"O|1�ۆv��R�$����"O��&c�>%��s�_�p�(F"O`H8�ʖ]j1��D^�J�� "Oz-h���u�ISf�IR����"O���f�+[6�x��n���9C�"O�B��E8^��<x��r"OLH	�DN/R�&��ӂ�G��@�"OT1h��"�0) �݅�^�x"O�TRp��j�3�I��2iCs"O��+gh^8���f� k���s�"Ob	(��Ce�\I��\/ v �"OU�CN�W�^� ��/v��}�@"O��dhS�4?��h��F<�|��"O\���Zt`,rWв;�F��"O,�a�g��D�����p�dc�"OT��ǚ1&7��p �Ńtq��"O.�#��+�6��"�9{s��"ObH#`��!��x�!�ƢD�6 ��"OPb�
"9��p�������"O����i%��!��hԣ ���R"O|Ջj�0�aG˓~ �Z�"O�,��j	!Hx� �E�!{��\٧"O~��� ��0=�P��	)p���s"O.9�W��?�H��Ղбi U�$"O�db���+S��Yu�ȋa��Q�"O�L��GZ�O���R���MG�`��"OJ�v�U�!����#"K�U�j�"O���V��;1�[B"�2TLݚc"O ��$��8��|k4�$0J�y{�"O���Ԭ̋4v|P����uF�5P"O�Q�FM�5
h�m$!9���"OTY�:3r�#�
�k�D�0f"Oج�f��;��Q�Z	G�lq0"O*Q�rdW�dT*��@w���"O
��!�[���䆗*,j���"O���j�l��I5#�6U^\��"O�d�W�[�k��H1p���X|� Cg"O����g��B�0`ӏQOez���"O�h�$bJ8`��y ���-^�4b"O$���l&`��l]�Ma��{D"O���ŀi��tx6ldS`���"O���� UC	~j5��;4��R'"OZ�K!J	y_�dQ�I�T��I[v"OpĚɋ=^�j��%���~����"O@�"�Z��lr͜�c��%[�"O� 3��ޒ\`�E� l^]��9p�"OE� ��5X !�Qʒ�6�z�R@"O� T]�a�k�^-��&\�8���V"O�X�h�$S朒5�?�\��"OL�[ǀ7in��ac�Oh�k�"OtT��˝�|o|��U�U� ��"O:���Pr�&B�X�&��v"OZ�XΒ�?f�*�+s����"Ol�{eρ�)˺�sF�ϔS�2!��"O���Z�p�d�؁oWX�>x��"Opi�F#�|�\x�dP�F�T�s�"O|(JdaV+Y��0��)g||��"O�Y�R��JUp']�4ZZ|K�"O`:We@�b�ec�-d3r�u"O|�j�W�QR(]�R�f0YP�"O.���c�;Ld�9�d�O�]���"O�`�̿^I��hD-�p��Ȋ�"O� �W�5a�"}c�*ۭ�*$�v"O$b@�ڨb[��q���U����t"OP$�c&O</X1�'W�${�d#�"O\��t!W� ߄)i5,�4&מ��G"O �#J�we�����
�#$=z�"Ob�����3t�|Bi��@��D �"O�x��\0"e���+���"O�|J���$zҔћҡF<i<D"Od$�7 ʴE�rx�^pR2l"Oz��΄F�]zv/�@���� "O�D{0�87[>8CT���p�0��"O� ���ߢzN��P�W1P��"O�P3�Ο>oB)�E�ʺ@�@<P"O�0fh�5�JC��P��>�b"OTeK�Z���)����jt`�"O]��ݒ�fr�-ɪM�Y��"O���a��?�6�X�L�J�>��s"Ovmh�OC�SV��U�Z�A��%�y�լ9�±��hģN�X�Q�߬�y�\�+΅�C(N�|�n2e��'��i�r��%�<��O�#Y"j��
�'���9���+x�@D#�*@��Ѩ�'���ݓeS���Z?+Hԉ�'i�U�c�ܢZ���
�h�;\,���'���VE	�S���E`��8O� @�'�*h��� 6�����5*^ѐ�'f�M"��������w/M�XR��i�'3,���-�2~
LhDŐ]I���'���BQ�����H.QY���I�'0�e��I!y L�S�\�O��'H��V
ގ���@Ǟ�u�0���'ݠXC�$O;:5Ps!ȋ�8��e��' �����UʆdS4fЫY�|(9�'|���b�Ows�,��Y�M���q
�'�R�BE	�)�TJ!L��m�1S
�'0�Cc�%Q�ع@)V��M �'������G��ቀ/O�NYX���'$~y����k8�s��A��ih�'�d����r�hx��3>�}��'�FTCd�/ZV�jG�M(-n���'�<`J���i�>xA+�*z
�!�'<LQ���?{:�Ѩ����$wL��'����%�/�0�
�H!�hm��'�:h��L6\���ɡ�Q�?��� �'����ٶ71�b��<�T�
�'�B*�@aX���7� ��
�'o
p�E(��|�5OT8'���	�'K� #4NL $�l|���-�F]��'n� A�Ӊd��ݛ�%?_�l����� 𙡂�0��Da��R�r@q�"O��;�䇁��� �#���vDk6"O�t���g�@ �ԃ�!��a�e"O�`#E�$̙3���;���"OLa��Ie��� � �3k�4�ٴ"O.���^�MJKQ:j�XbE�4�yλ��#�� ]���)��� �y����m�G�D�N���%�؊�y��,O�t�bg	�L���,�2�y���g1�0	�ȑ�7���1CM�;�y§�=|���SJ�3{O��ӣOſ�y���T�d�U���W�i�ᐲ�y"��p�TX���%q-�)kfZ/�yQ%Vv8�1��N�dZ|a;����y"�%_ ��R��k����vfF��y�,�$��VJj.� V�Y�y���2bz�VgH\�)UFץ�y�� �q���`��hBDoŷ�y��_�u,F�@��G�Y/���
1�y�lU�2����0U$Ԁ�	��y"�;wq�����S8E�`�9�G�-�y�_
2�ր��댁l�D��!���hO\��3Q��@���8����F:џ�F���0R\Z����R��� �����hOq�ܘs�b��S#�d��[F �j�"Ola�W*|�=HE��)g�6I��"O.P&K�-�$��Ą˙s�j���"O�Ġ�m!�^��EiOYpTi�"Ot�@C�7U�:U[(�ak�y�U�'��Ⱥ����[nx��Ve	�ܬ��p�)D�x"@���6@+㣈�)u�б�-D��0�b�NdNi�Ҫ�'��xk�)ړ�0<!J���d�������!z�R�<1P �;*:���E L���qd�P�<��LȊV�����l8�9��P�<d��i����UM�I�fe�t�I�<�-8tC.0Q0Bԁ+����G�<1 �K�j��9A���;sL�+�j�p�'�ax��.OoD��Ƀ$o�8!:�#����<���G�>R��� ��6��0�ΚZ!����V0xbK�8� -�v����!��$:AD�� �h:�k�"�!m!�䗴v ��jSoB�s��!��X�Z��'�ў�>��1pw�x�H\9`��@�Q#9��7�SܧhL ��ԧ�l56ZF���g�H#��͟d��5Q�ϛ%��=E{��OȂy� �;e32�ڞ��y0M>�,c��`�Ӎ-��-�gO�V~Іȓ`X��'6��}���"?~!�ȓF�r��%�"jO� S��ڟj�
D��S��xĸP,��6��D2�k����C��$��y��;j�B�j����x��C�I#n���Y����|v̈1����?����) ?��+b[�KED���I�<����;��Y�4�{r�mS��K�<Y`O��X `�YЦ$SPnũQ�F�<�2��{KNA����0I  �m�~�<OխC�*���[�K׀�#3��}�<��UvF��$�^ AmH;C��A��0=A`� �JlB�9# _�O/���U�V{�<��q��x�l�9jv��P��z�����O0�$��N���
�nU�����'���S�%�g�p���<�(��' RYl��;<��B�Ԟ.k�%���� <��b׎ }(�(�Ý�F��q�S������|�&��CO��P+|��"A�-6�C�IN)&��P��6"��5�t�O��x����x�'�d�D��l�Q�S+�x ���x�
��z�u �R9 5r"F
�y��Ăr��9�M��*����'���y��]�wRIaf!�r�0DF2�y�i-�`jDjq�e�R��y�ƅ;Y�|������ 3��8��'Gaz� 	y��%���4 ��KAn��y�A�� :�&Ʈ) y��!9�y$�"���5���'Bz�#P썋�y2m@�B*J�C�3{x��4��yr-C T�Xӱ�Ψ�����y�g��)����e�_>o�0pbC���y�J:�0�3��LQ����T����0>1nR38���ѣݥ?N��R-]d�Ik�'����<aD��Isuj�!A8���[a�<�V��v������on`AkA�x�<�T�1|�
8�T�:K�R\�C��?J\�YB$��Q����E՟B]�C����b3C�:Dp�eC��Q� �C��/pu���!��*�q�^1Tn૎"�)��lN֎�"���#WX^B&�Y��y򏀰<�j�S�lQ#Kn<U���D0�y⏇=}�
����Ќ>� �����%�y�E��ZĴ�#me� ��װ�y���eH��t �"U}��hQ*���hOr���@+[���kakŭ(��TK�
��x~!�U,v���%	/+��hC�nF�)�!��I#�J����@����#��2O{!�DǕp	�£K�El�}�`�MI!��kH����٘Kh��Ӕ�Z!a�!�ċ'@�<}R$J3�,������!��_z��Tb�
|8�:3*���!��W�b����I�p|-Q�
��!��\C,�|yvN�U���cB�7��O����xg*Uh��:E���O�${!�đa[J�;��@�%#TJ���S!��@6��tI.��[p|:��"C�!�64�jL[��I�h�1ɖ�!���)�`Pg�_�"9H�'O�!��5I��x���v�8�c��r�'Vў�>��>Y�a��6UʚT�§8�$*�S�'�Ƒ��L��^A �Θ�o �t��	b~R�.���.��җ\ @�J��
�'��#G�� p��f0��	�'k��ImQ�=�aS��D�2<��x	�'E���/Xǂ,s��#�����'�`�0����У H#ZBQ�I>������1?v�k� K�vXF@Ƃ��+2!�G+x��z���
{AȘ�C A�,!�D�!z$�5�ƤKV���<L�!�J!�����%��DK���A�
|q!��U`�d��@j�?\B�P���!�Đ7v^T�WJ՘!Br�h�/G�!�I�Qi�焦j�lhq歁$.!����4@���V��)YWBƍ<!��L��1��Ց:{䍑�Ւh�!�C�0���t/X�Wu ��Y�!�DĚN���nmb�SO	�!�$	�gy���g��`�`���z!��Ta $��OE�p�N�BUI@��!�$Q�e�p1�g�����a�`)ȣXo!�� "�ʎM`h��lDj��@�"O��Y�LN90#Z(Ɂ,�)���Is"OZ����IUR�È�;?�d �b"O��Z�fQ�3�j�����k����B"O�
6���1����0�W8�T�p�"O\��3C/w�dʄ-·v�>�1�"O����.��P��A��'��'��6B׆��􆛜_��@�ȪB�!�Ĉ�G]�rdB�
����흄*�!��)g��I��D�������&�.�!�� �)f`�i�m�>w��mC�LO�!�G3� L�g��J����i�N�!�K2F���-�0�Rq�o��T�'�a|�E�'�<���'X92 �j�P��?�(OL���P� ��`i�iA�X
��6d�o!򄘔V3��hs���y
F��6B��3|!��D_�\J��Fz^�����Mx!�d��Y��u�vJJ�
����!��SPnm�En�0��-�6P:�!��j�$D����6�r R�횎b�џ�F��M��2��p-�<O��v�B:�y"��>��ip�+��E$4k%@՘�y'ԹBo���g��<�P�)�
ŷ�yB-Ln�R�C��A-k��TnK��y2#����!c(  ��<�'
��y"f�2-|����$�Pˆo���y�e���҉�1�Ѽ"�As����y�	ՇjR��#�#=�ƍ��ɨ��<���D4�\@���#�V�X��ǚ*F!�DV*L��0��RF�0S��,[+�y��	� JmX�&�WHf��*]*"B�I4�e�����iX(H���+'B�C��6q��qm�c����va~C��1R@��A�����p��OE��h�=��'���eZ�u|�[��Zܰ�ȓYa�S��>�h�c�FIa�Zȅȓt�>9su�B�m���5� �r�4���鶨��F�A]]��,��F��ȓ_ЮL��	\t0ؖ��'𮹆ȓc�l��3,����[@�A�Ky�!�ȓ7=��IE	j���EdF�%�0}�ȓ��-�rd�(�X��s��=�DX�ȓ���h�G����cs�<i�x����T�f�F�T�����6<N��d&^���#�����*s����ȓaP���2��9���7����qզt���c �#6NM�Q`v���$����m��镎�3����ȓT%��`�8r2s��W��%$��G{���M�v"8�;�\�>-��b�X�y���V���<x��T���y"F�T��z�㌮~�t	�$�E��y�&S�#( ���B���tɇ)�y�j]���
��;����AG(j�)��#%|LR#�϶5n��&K��j�|��ȓ!������Ի)�: ��q,XY�<�ǌ�0���@P��y�ҋ�T�<1��S�F ^�䁛�FsМ3b��w�<���߄mP��1�.F������p�I}���Oܚ���ɗ?��´�:�pQ
�'<z���Ƃ�Ϯ�Aw�^���$�
�'��5R��8.+���(� �ک�	�'|` ҖGр�,֯.�d�I>y�z^�I�V žDz��RfEI:l�p���S�? ���
 9�FPk��l3����"O�������#]t=�w�]"D!}��"O��&֞�(���Μ6n�ű�"O��Ђ���v��(����c\D�""O�Qc
$T^|X)w ��E�x���"O& Z�/߹')SRA�"6T�p�"OU��+L�oB�(���Q��"O�ɓ�%��(���!�0|����G�'����ʱ�iY�}����Y7T\B�ɵG�J�(���4����[	2B��7
�`��E�$O�q�%n�����0?��Iו6�z�pUbY1|�:�*����<a@KZ!�&���
.O�Z��v��~�<�Uo��B�(t�"��	��[cN�}�<"'V3{Ĕ�J�/=M�Лg�a�<�5�& ��l:�l͹}�l����`�<��Ŗ��!��H=�2��І�R�<9G[0)���ql�UmyfKAP�<�Ч��@r���	�B@��NZK�<!�@���䀐��	Yj�@D%�]�<!G�	y'���BgQ:�F!�*�n�<QBF,�.�el����C &�l�<AA*�,�j�`�/c�l�K2�l�<�aF#����G�"{�.���͈k�<a���@��"6���+�0����j�<��ܤ[P�J@����D��e�<�#L��M�����DЬ7�� ���`�<�BE!l���#Q�Lޒ����Y�<a���3h��c�G�-Z郔'�Y�<y��3M�!�c� OA����U�<���*��p���oV���N�<��˝9_C�ة�X�nI�y9%�M�<i�@�s�^�I�*��9$�MG�<�o[�r�,�@d�d�T@Q�Hn�<9�.��E���i0 Ô~V}	$�Rm�<��F]�S��H�sĜ;E ��*&̚k��hO�':�!J���;l��g�eI�ȓ�M`Ʀ�)�(@T��!�r	��K��|��k�h�I��Ɇ�D ؠ�ȓDI�E�J�ʅJ
��!��|�<�V�ι\�p���7�ؔYâv�<�w#�;Jz1��.4ROd�I�]r�<�+ۊ`"�=化�Rg�:3I�F�<I0b�8.�1!���N�����E�<���Ő՘��D���:p��DC�	�F��-b��ڢ,v�UkEOW�(L�B䉘?������i<����V;,e*C��	h�P�7��D~UkQđ�N@ C�'��哳���/*�T8���2:w���d$?��-^�	E�l��}��	���t�<�K�
vŎ�cal@���Pƨq�<�&��?>w�t�삁W��`�)o�<���M�w�l��Ũ(?�J֮]A�<��K�z���xg" 9JV� R�<a���v�He�!
9ȼi⧛K�<1؛x���᪛!X��a���k�<�m���(	 ���!�Fi�<) �¿�\���--�xi��Ky�<��0pkH	�*D���bNL@�<iEK�� 6<8��R#p��J�I�d�<�R�P�V�~�4�� 8_��R-a�<)ck�X}h(�6�0��X
VT�<��a20�mb��:�
�.�S�<90�3eD���U5t�����Ux�`Fx
� �)�W�ϓ{?D��`�݅)ٸHW"Oj���L6_&� WC��*�vtI"Obe���y�� ����q��jC"O�Y����Аj�D~�t���.�S�)�b�6{�Ԯ8���G[�{=!��-v'��i�� ���1%��5O!�dߟH�
�A����[fEL2!�$� �$0�ƃ�:�t��d�!��Ob�=���ukƢڨQ�>Ts"��4_\V<�"O,=k-�T��d!	A�W�!k3"O��C�B��E�g�;@�~���"O�����H����MJ�"�SC"O�)%���W��|�7FE#��RD"O��D��[��� ���k��@�F�z>)��`R�r�
P�r�_�i'����Ĺ<�+O ��7�&�J�bOC L@a��p�8��"O`1ƃJ�E��x°�U�<n�b"OJ���DD$���&�/Hk�,��"O����
��\�-����f��KG"OBI
�7v �M�񯙿
c�mb�"OTP%��
�����JK�h1"O� qwjİ&r�Vj_��
�����Oأ=�'X�x�0ԉʌb��Ԛ%H�6d�L��Pa~U��J�?��zχ2M���ȓ%��e��'��Y��P�߮3f8؆�?�\��bʄhGN'G�D�ȓ\~��$$:�y�Q�D>\`�ȓu�@P�"h	�{���3�J���l�ȓ�T�a�׏S�TY�んu. �ȓ��M+3 �-/��MC�ꀕ;���ȓ/�2��������sEm�i�✄ȓM�e�T朅1D,AS �%v����ȓ4�4�����0q�+��!=X�لȓՂW\�!��=�� �<O�x�P"OLa@ ������`ƅS? D��"O$�@�HZ�0+��-(��"O�qb�/$�vD�&����D8�"OX��U	��E�.���
�����"O&�KtC��u��(q���z>��E"O`�{�����ʅk��g�P�"O1��M�c�N����7-hL<�'"O)@r%LY��p2 'ϖM]���q"Ov���C��O�D�[��P+LS�dI2"O�|�!� ]s��y"*�%�>��"OJ�Y�S~�X�`@#G]��0��'��	�6�����Q+bp�$L�4C�	:�v�bi[�W������FdC�I4_��@����)hX��.O�DB�	1#_�ѩ����J� �B?H�8B��*.��eR�b�r����f��(�"B�	+Xk q���ڷo!�B�ɚ}o`ȊW��(�İ�$�\RivB�	A<z����	 '��d,��O�C�	O�8����՛D[�FF�`��C���%���{%�8�|��"O��O��a@FXaB�P��p= �"O:�r�Г:8�z�M�;��ʲ"OL���k���Z���S�;�HH t"O`�cb,U{JQ1��h~@QQ�"O�� 4ĝ[�q�L�k��c"O�mj�̕
N�ՠ�JH�,�J�Jd"O6��s�]�|�:��ށ�tt`�"O�@�TH�02�IuGK�N�z�"OT@hb!�4'��M*�-�Qj�H�"O�  �r@�P=�|��5Ɯ�S{��a�"OH��古P�,�4@]�A�da"O>�HD�c�u��Wx����"O�iX&@��	�غ%,C�Bd�'"O��(�Œ.�@����1+���Z�"O`P闇 ��/�/�TY�"O��X���E��̈:�.Q�"Oȵ�0C�7�6AF��l.��(C"O��!g(�M�6��!h��H�1"O8QѓҒy�L ���Һe�Җ0�y�ŝ�b�B82gb�	@hZ������y2�I�o��EI�ď.Mdc���y�%Od�}Ycˈ%��DQ0���y"E��5�0=hu#�O	�tSd$���y�۴>w�M�F�E�vh�S.״�y��?w'�4:�i��:��8��)^�yB�,{�`	�$̎�1��$��f��yRG�#��L��$�te�ä�����!�OL�H�%��T�Z�:�`G2pq^���"O����K:�$�QW�Ę`"%p1"OB���u��X:�-E�NL�$��"O~\h@�4F�t��FT� V5�"O"�@��%%T�Eo
�U��'|�cF�D�[ ��k�	�R����'5d``��uQ� ǂЌF��)�'v��JU����&Ը���'�R��
�' <��SF���(֫P�1B�
�'.��7�(O~T�ȥ��*+�L8)	�'���*pȉ�.��Aش`� p�h�	�'? [��,I�f��qX�� @	�'�l�эNL����AĠt���'�He��C@q�3Kքp�R���'�H�3�/�-,�}�[�lY�-y
�'�X�h� ø�����Nxr	p��y�@��<ҕ�C�=*���[aDI��?��'���F����,���Ƙ
L�0��'�Z����K�_~�XYQ���|Q0b�'S��)Y�?��e��,=�NA�'�p8�I14������*�T���'qx�Q�Um��H@�E��� u0�':���eV�Xࠨ�b	�(1��'(f�2��FĂ5zu��*R|f44"O�����;tV�z�HL�I��"OH��!IK0��	S�N0.<:�I�"O�(Y	ͭO\�3��G�rz���"O�|���ÆcZV<2�D%\�H���"O�y��@M?u�]�t�+}.�˂"O�2��R�"�X��vbI�s��Z�"O���5�������DBk��R���D6�O �;�Eu;B\�g��G��a�1"O��y�HW�dU�e�4%�����'�p�e*W*��B�D�V�9�'^~d���<�=�1FN�B�y�L�edPi�A�;�ވ:��P
�y�	T�M�
����N�:c���Q&�y��?��!�i��+��I"�4��'Jaz�(P�}� ��eω#�xs����y���Z�B�D�i��lZ�(G+�yr.�.p�v #W$װY�R�3c�O��y� Ҥ1��q�P�Ь(ب�r�c6�yB�S�efACǉ�P�l(����y���B��4Q�HH�H�ƭK��ݫ�yjkh�� ^u�x�0J�y�U;��%�2g��ӇF���y
� �U)��-wy���T����"O\
E�6*���I�*�>[e�U��"O�X!6LЁJ�&������{"Ov	�Fg~F����A;;�����"O"�[��?S����&I�]'��"O�hI�R����bfF�l� Bd"OP�C�\�&q�h�#U�z�Q"O�5z�/�0{f���fc�<-�ꍂ"Op�
�G% nd�#T85[��4"Or(��ʓ@� ,٠a@I����r"O����#�;Q��x�31-����S"O(��Aa�q��mT����o"O���#סK�^`�&cD9%�� $"O\�(wI�2J�xl���O�b�C"O��B"-u#J�
u�L�L���1W"OL�[�O9�lڒA�C��0��"O���.L1SنB ��y�D�Ä"O�E+���.n�T �a^��b@#"O���M��z$�����8q�D���"O�!�DL�}���R�-
�>���˦"O�@1VeE�7(j�����/;��"O>���l�Τ�����$<h7"OM�ӊ��25��:�U5��D��"OH	�rlF+g�x���?Qڌ��""O"p�Eꑍo�P%��aײX]d���"O�V���/�Ea��@X�B�"O��R㩋� � 8�).,-��5"O� �d��0r 1�Ph�$^$L�"O��p�I�&�v$�I��`��E��"O��*1�\�
���*y�z�cU"O��fF�i9�ybP���2����"O�����e�4�+�^����c�"O� 1�Ō
<�P��DUx��+"O��bV�DrB�1��)�9y҂ �"O�̪uk���I���&#f�dp"OL(��nS<j@+d'�4����"O2�93��o���p�����5;�"OnT �L�d���W#���W��_�<�HS�"�9<�E �-�S�<��=>҈4���܃DЮ9Xc'Q�<9�n�$w�$@�T�CV`3�^d�<YS�bj��1��.:��T��G_�<)��X+[�ro�)-����!�B�<���+�e{�ʋ#}�KUHOi�<�`�?30Kd�
�xt��(i�<yf�Q<`�ѧ�P(~7td��K�<g#�?b�H������ � �-�]x�8�'���"c��5�
1�`׳[�|��
�'ۮ��D�'L��r@M�6F1
��	�'s�p���Y75��h�į@�8z�z
�'M��D`�+c,�aHܧ4h
�'6R亳e0$����\t����';>�$S�Y��A��.<u�BP��'|<)�e'J5g�n�2�Q�j[b 

�'�*������֠��D���&��
�'��*�c����K���c%Д3
�'����g�,-�QfGA7' *
�'2�!pV<H��9���	v;	�'\�9k�A�6�.y{5�W&����'���A�?&�$49�ۚ���'�(��������;���'���	eU�f������-��"O��3F�V$dn�ȦCΫ\n�#q"OZx��'�z"�?\�@�"O� �x��S�Mt�R(��j��D2"O����Ι.w;Z	���(~V4�W"OB)r�gM}�FQY��S� VR�X�"Ob�xŇ��b�����D�Dd@*�O`�T��G�6A1U��,^�:�xT��OPB���&��PփRA��m^�C��4x2%RP_�'�����2�JC�IQO*xQ��:����d�~4ZB�I�k�(��o"$i�AӦ!��R�<B��&E�|pb��T�m�&a2A�+ �&B�ɋw����^� 
%�U�$-0B�I�~�RA�P��%Rl.��ՊJ��<�&�D{���+�����g�Z�1��,�C���yo�����j�"�p�3�Q)�y��?nb�hEc�#h���B�W��y�삽R�� &B�;a�~�9�bݘ�y���ff��W���*�x��T�1�y"!͔S� )�G6kE��Th���y�	 G�T0R��j^�i�5.��y�'�:m쨱�h�N�KD���y�J�Z��U��@����)3ɘ�y"Ϛ+B*,�bT���%�r,
��y"�X�q;������� ť�y��V�c~����Q1l�(BPKC��yU@�*y�1G�Z�x�����y���H�����d�e����5�y�l�(bX`9�'V4��('#�-�y��8B�0�K�R���B��y��3�0-����*\��	��y���gk�E����k��g<�y���2K��x�'ò�f� �AǼ�y���D?hqG�U\�,H��G2�yB�@�+9 �cd��a�تvBօ�y�WM�ޜɴ��_�xI!q���y��ŎI��˷h�?DCN�Y�j��y���S�t vd�$�b��+�y�����$-��~�#��^��y��͚��c�>	&�C"KW)�y��H� ���FQ�hR	0"�̉�y�j]�6J�x°�X6���y����y���1]�o�$�t� ��	#�y2��;^��}�Fď3<�6D����y��;�.9�e?.6huP0	�y�!	BnF6�0aEH����Yi�!��\h�=��l�[)�]�"�	b�!��>g�v�d/3.�Xa��&�'|!���e���x2���n�`�"�p!�Ǳņ��J�W���	v��Wb!���f��iЕ�N]S�b�a:wU!�D x��8jV� J�1c�`[�H!���7�F�;V�G=jE��)s��:�!�d�t���z����  n��F�W5�!�$A�\5�=�pƻN���m�js!򤁲0K�� !��c�#j�	=�!�����`��DM�N�Rw��	!��.�p�EY�z��8w*B�	�:E�9���"Df�� ��:L�B�	$@ P�I�<}�l)��1�C�I�b�0b#�+�8��A��F�C�>'Bi�a�@)%t|S�$'z!��D�F�BMCDS�	3�A�����&�!� s�\���(��1���®+�!�D�g��bV�!l �.��O:!��'6�J�hքS2*B�a��.H�!�� �d��.0w�\�{�Ù[$Hã"O��[�Nߝ2��`З�W�A$�'"Oe��.��K�"e��Ce� )�"O�p��ߔf~@$���֨K��}��"O�"�k�qRΥb���O����"O�!�1�X-N�ȡ�4k�(�"O�R�`ڪY��m�q�F%�"Oz�z_)n�KBb�H�r�+��t�<aPa�3r~j��1�3d}V��[�<	v�ɓ��e�%"�1�`I����<i3�����2fB�!��d��Jq�<�&@N�~sfQ�#� ~�J���/�C�<@�R�l�Sw땢U��9�uz�<�S\����ǝ���Ш_�<�"惲8D���h�p2\����Ea�<1sL\&J@�B`/D �!�/�s�<Q�֖dz$13'�'3����.Ll�<�+�4�4Pb�c҉cAE�#Ym�<iw-�2��͠3+[�`b�#2�~�<�d�;'D�D"܀W���Ox�<�� ���q��LQ| �"�MHt�<��@M�d"}� _y81�VCBo�<��G�{�N(AC� �D0���i�<���[��d]	n"tBE�l�<a��Zx�1!���w��l�eÆs�<Y� :R�ְbE�/c�Ƞ� �q�<I�C	��1 �%�?;�����DMo�<�A톽nh{T��#|���
�g�<	Q.�<b'�)�	�&TD�y��	d�<�UfL�A��	���C#��@U�<���Ӏ,3p0�A�ӥ#��հ4N�R�<97��f�:T�֋ӇG����f(�Q�<���|�<Qѡē�t}f�%�S�<IEɃ/9V�02b�0u:�z��R�<A�iD�НX��Q(K� �@CTE�<I�o�O���;�&P ㎜H#�w�<	d��@G:l���E�l�Cchv�<�#V�4&&�22�R"�"�"!��q�<!�(��%��\A��/m �)�b��l�<�t["6��њ �@)Z �]�4�\M�<I���Ӿ���K�	/�+C%�J�<�BMM:>�tA���"������]�<�W�#��j0�&^|r9Z`O�X�<9��Q"
�VD`Q��$G�F��o�L�<a���@��h�U���QP� F�<QVe�-���#�Q F:�P�A�<afk��,��:�AB�U�v鐵`�y�<)��ȍG߾�;Mɶ<U�]���q�<�� -	��R�F\��J`�U$Jq�<9\N���c����`ĂF��!�$�2c_Lx�$�����у*�!��Ro��	���+�-х���p�!�DG�F�(�dS�8	�}1�=�!���N�Mj��90��i ���!�D�sN^$yB�Z4Z~e#D�:�!��W�jp�"�(O���+��Z�>~!�$�;<�Bȥ.��"g豢T�N/A�!��?d��j C[�d�颴"�V�!��ϋ���r'�`F*t�c���!�=
.�1b98�ؘ����lu!�DO'p�� ��mߝF�E��Q�pg!�d��h%�Ԙ=a ���AO!��R�
������xARX)�/!��ث_:$9��a�;0X��ĕ�j!�� L5;�cW/|�C���>0�P"O0R���-aӦ)��e:�:"O��@T,��e�J	Xp&��d�RQڠ"O�����VÒ�S�n÷�"r$"O��� �����l��,�*�"O��ԥônL�A{�m�	f��H�"O��7�p �ݸ��_�Ph�:�"O�SF��bąH� ��[I��8�"O6�b$�:]� Y�͂�$2����"O85 ���%��h�`L_4_,���"O��	D��fHW�IjJ�)�*O.�I�k]���eO��)�'.�hǆ�7����
���B�'~��t"-?0��B�H$
2�Q�'2B�@1'��B�:���d$��
�'frY�v�G�$d�X$';Vg��A�'�68H��KK.���]�H���
�'��BǂӌP���Ίt�؅R
�'6(X�#��-T�a�#Ѵo���
�'��ՑtmOr��ˀ,Ѓ\��H
�'��tZ�h�R�Cp��"(
.<b	�'>0��d߅$Y�t;!�~t���'ͤ�Ӳ(����Yj#��͛�'�\<rEL�? Yk���@xd�'��azЎ^�d��,X"_�� �'Kp�A`�E�8��ɸĒ�
�'�0Y�d
G!������ݳo��k�'_ Ax�B��t� �&�Ǥ7/�m3�';H�����;W���o�_�9z�'|=���A�F�
�8�=�	�'�R-Jt�5�
ȹ��p@�:�'�^����6O���)�Z���'1��{���-�`�SR��!R!��'ᄄ
��Dmnv���dS�'h�8�'������% K�6d	2�0��'�!PA�Π;���,��r-~dY�'��y��&M�2!D�[ŧ�=v9����'h�x#7��(<�|h�΋#n2z�*	�'���rSN�'�������e ���'z��"���k���(��ʊd����'���Z�)܂V��<���6c�jA��'eB`��)�Z�|�r��֊�x�'䔽j�NR�M�z�3��/���y�'���hQ.Y@�Ӳ�͑,�8�'��@p�������+Y1V���i
�'��5�⬜S��5֍P:b	��'�P1�\l��[�,W�Eb��',��V�S�wM�LJ�bǝD��I��'�6��cZ�s"��NΥ<�q*�'����%a��psL%���G�=ޚAQ�'* ڇޣgz(p���B&3����'�݀�B]�:V\��4�@�0P�0�'�@`���6Y�&�"[f����'��$��K�c�Z�Y3��)T^�$C�'C�b��� >ڍ�bV?,����'�x��#��Q+��+b�&0�j���'լ��b�IS��x�Vi�#� $��'B�(\u�:@I��٪"�hi��'N8�R2��]X(���$F�`�'ȡ���.��w˓ HT:�'��1�Ǌn��!k��N:z��q��'
��gIL2%������@�"a$%��'9N\�RBV.q���g��p�'O�`h�S�M�hp�v� e��b��� 	�g)�&���N/��q�"O�5J�b�%#���E�D/m�J���"O8�� #EM�~�kT��8O�N�۷"Oh4�GrrcŪ�1�|C�"O��3��pbԩ 1�L�]�X�H�"O
`�C�&J��6�5�8���"O�ݨ`�s�T˷�ݥQW�Mr"O�Țp��;���3,`�@�"O�y� '?�h�щ��R&ى�"O-��� �8���@Q(_5�^��"Oĸ��a߿x){��]-H}�"O�PQ����;�
���Y =����"O:	i�j��x��!���RR�v�P&"O`hHܪM@��r��h�"OL$8�æ}L��2�@�_�m�#"O֝���I."(��E�A8sY.��"O�,{@/��ձE��
V��z�"O0u�R�-BC�aI�� 9Q�e"Oց;`#W.����%W��;B"O�����s�ԕX�H�B<d �"O֩���� )����M<*�p�G"O�Yɰ膩 �@���G�$Dыp"O��eGۂDĐ������>\���"O�if��f�z4���w�`�"Ojx�B	%(I���h�
 g"O˶&>d��[����E)I�y� Ͽ
���[5��Y,F�h����y�T,<]l�sg�7F�(Ŕ/�y"�	�)�	�	T� �g햩�y�m�#x::��(�`��c�O\��yA�_F��@����T�ʭb�Ɂ�y2c�	�N���!��\�CfFP&�y*�=�� ����?~��pɅAƼ�y�IUr�0C�m�Ic���܏�y⃂ �Bd���u�`$�`��y���!��d���q�ؘ0�.���Py�� �|p�D�X�~~R�;�EK\�<�E�T�H�p�cVs7�ȈY�<�F̛�3�,�#�J��2C!�\�<AK��V�H\@�H��o�RA�@��[�<��I��2���.K'\G��c'�Zl�<��C��(�ʌ��CO$Bye�q�<�ь�6I�!ie$,���y��B�<p�Q��R�D�I^֝��E͹!�!��>��"k�,u.���'�^$<�!�䍖?��Q�ɜs!"��"�P1!�� �̉`�B&�8���!�4c�!�dD�Y��1���̫����*�#>O!�d\#X�$(��v�X/�	0!�P�-��L	TC#V�M�!��P@!�$ޙiY܉i�7 Fv�bw)s!�$.?D��2Ŕ!4
x`����!��2.<�w�S�@��1��A<�!�$��hb�����N�lά��C'�!�$��5U7ʃ�s,ۂk:�!��J�o+���6!Ƨt�q�#ߢ�!�d��K��Uj�Ybl��@�8x!��,1YG��p'��'�N!�$�0B�dDq��3�ts@j��^�!�G	����&3r[�(T,!򤜀Y��#PHV�Jyn�8�s!��ݜab�4����m�^` ��S!��0%D����"$Up!�R��H!��>�(���C�+���b��>]!�� �	�G��R/���3jX�;(N�9e"O�\3�(�TlC�� ���(��i+ў"~n�	:"]
�g�=�Ȝ� K��?_F�OP����(b�lJp�[�$k�d2�,¯���^�� )0#C0�X@�I9uD�8��5�.�S�'T;�L��h�!�P�u� gBԅ�e�L5H䩞�6ǜQS�+t��Q�On���ˇK����93�\��"O�2��ec(c��ƨX0��`"O�q/�R�J�W��	?(֍k��'��	6 �"D���
-|����YqB�I�&>Lб�^�*�(+�O�g�BC䉔� |�DL�b%���'杗V��B�	�eP3 ��	���!�+?
�dB�I�)-^���)��drs�KR��G{J?%�2c�/�@%�ͼ+yH��g�j�=E�ܴ��@��S/(p�qw��X���D{��'3�ؓdO��QAn
?/�a+�O�����X"��mݹ`H=����	W+�	�<�J�ЦOq�j��"
�2 Ҩ9@�.��J��7�'i�!��؇dl<��{@�V$�D�MH�	Ex��)T�r�R���� ���P�DY�=�a}>iC�C�Q�p�ްf'��(Ɇs�g��rD�C[���iƲ����f���'h֐G�tcv��yu�P4���L��!�p�A�4D� *H#	�Z̲���-}$�P���T;�4��SF{@�;fIؑxR ۟<f�|*�c ��y��{��ѹ��U
j 
��3���y"�'=0A �O$PcPd2�I8*4p%q�'mڌ�R�*��k���*�����'m�(�P��=\�&��f�O�"�li��'>%���N+�!�ך.6�)P�'���a�/�<ƙ��O�z���L<�r�"|OU)� d`�L ����DH���Q�O�U"�c;S_�	�e�]-u�  	�'B���g� x�B�L5����O���D�4D)�6����	!#<!+A�C��y�"$�z��G�$l��D��yB"�3�����gdv��Ə��x��'�IZ�N�2-�&��Lʂޜ���'�a��ȩm�)���.춨���N��y2iLO�2h8@���<MA����yb��/�� c��	"��wI���y�nΥ#����FT�O;&�/W���'�az�n��`J�9�, BV+�N���<��k�*#��<C�Ӱ�*l�$��@
�B�ɣ.Ԥ,Z�hf�=5st�@!LO�X�>`�Wr���Z��Y�q�� 3',��<���&"˪EksLP`�jYZ4��y�<�U���(���a���Ф�V��t�<���2f�(����4H�9	ap�<��c[�C�,��W��0������k̓�MKS��>IO|J˟�m�!�����D#��?���q2������'cʽѥO��D)fx0��2Z9P�6&2�S��?�&j��c�! �N]D��"'ȅX�<�(ΕkT�E9��؃�|yz�	�?���'���`cT�Y�uNU�͟�L��� � 9��ۋR!����F�"���ȓyl��2�J0Q��Tj��ٰ�B����O�'�Z`3�K\����j1�$Xz�N��3��'����E
�i��\`U%I�O�K�t�Ik�����>�6�ϡU^VP)�'Q�:�ّ��o�<�!�4�0!*���<��ᱠ�7؈OH����(D��ɲ��ԕ5@`'%M1!�� p}z�C:*��p� ٦sH���%"O&i��U�I*(-c�\kB�����Oe���i�Of���@Cn� � ի߰w%ȥx��x�We�����̅Q��Ӑ�|��Z��-� �=���'o�S��?K&"U���Ucb��@h?+.�C�	���r�G5^��)�-�% �P�,�S<��}�pd
�M՘@��D��Z�xQ����Q�<9%��I[�x�HȦIx�����c�<YU��*k���AɞyM"I���J̓J̑��'�H� ��R�B���l�"ap�q�+"�Dܖ�0<a���MVB=��� eߑ��J�͙�<�L>!*O?%���1����BK�_-�x᳥=D�����.Z4���bLK��J��0?��O�Ósl$rG�M$r��"�ߑR��p�ȓ*����G!4Q�4C��H�<�;�4s��oDC����q�:�M��y��X�]��!�#&�8:�R����e��D�>��!1���fV������az��=	\\��?)V��d̮F�!��1�g��z/�9��$ma��"O��Чm��*�R��R0̔�"O���
®�@�{��V�t�5He"O�u��HGWwd�qw&^(g ��6"O,��[M<���� w�(��"O`�t�r�:Q�r��vO���0"O��b2�-e�pm�*]>�H�"O0(��H��L�&	���	~=0P�"O��r�;�8���E
�:-4�"O�Y��1FL�<I+E0E���"O���B�Ƹ4�b� H�`����"OFU�A�V���dȚ(���P�"Op,��. �q�$��1	�L�c�"O0�2
G�z(`��0�����"Ox����m�`4���  �^E�!"OD Ys�ԗF��5:�A,Z�ne�7"O���� J�;��4����*�z��'Nў"~ZЏ�y�ɢ��

k�O-�y�Y�">�b��S!_lTS��@�ybDPn>�+���eϚ���"���0>iM>�dn��-J��q6��/i��H��^�<1���?)d@`Ri�)`���@֨K��hO�1E{��Y*T�kbg��k�Z1��+����m6Uis��5!���W���{� ���$;�O:�PCg]DRڅc�,̏e�t�(�O���&_^����f�3e;d�"D���,�R��R$�t�S`�!D���W���!Y� �wj��/�ȱ2	�''�܁��� C��!���$�C��hO?���5v��S#��5@\� ��<��ضT�<�t�O�,�	��NV{�<y�UC��<1�BJ$��u��5T�X��ث٢a��-&�|���:D�`���{�������Tlf��i&D�����\(2�`

Z�t���8D��S� �@߼�I��l�BV�:D����A�;pZ��dȉ�C������7D���%�N����wd޹rD�4D���q�G�b#~���N߹}��1��M(D�`� nO�`�d��-�{�l�� '&D�̐�!<e.hb"V
U�h��4�6D��1�"�:b3�AT�y��\*g�(D�l`�`ӧ��|eb�m�R,S�*O�]I��0y����Ǒ�Ȣ@�"Ob��RL��NVi�էK�1�\@YP"O� Z�2޴bz������o�^鈲�'��/���9�G҅@Y8�$ �27N��ȓn������ ��5�C!��l�$�ȓfy���rJ#"��F�$|MB%�ȓM��`W�;4��kš�
��1\L)zr�\+J~�y��!E�cȶQ�ȓN9.Qq�Ƶ�d�W �#|(X�ȓx�蕸���3�2����$4t�t�ȓu�x|�'Ý n?�h`w$7�i��yGj<3���.vH��v	ʞ?+�ԇȓF�F�SݺV®u�� +�1���T��u@�(r�͕�[�]�ȓL���@��s�I˓��
j��ŇȓC�Z�J@a[*�J��� Uin4��l��Au�$<�-�@F�{�rU�ȓ	���@U4O���%G3�ȓ0��pQ��2y��U��l۾�m��F���(Q"��(��=��l+�h��p��|��)Eh��:�l[$��@��v�d�##���X0�D*��Ԣ3}Ω��V.8 NJ�������Q�i�ȓ9�.D�s�FZ�4�F!��jk`������ʦ�Ė{8�A�D/[�4U���Y���g�n�Vcؠd:\9�ȓY�Ju��cٓ-���B�����b�(0����!A�H�p��1�K�<D��9�F���K�/�$��C��J�<�T�>Vf��ad�*�<�k�A�`�<�&,8'����.	��ࠀ��^�<A���%*2�#r�� �)X�V�jąȓ������KL*�!���L1�`�ȓ%�ֽp���$Nvyat%�,{�*�ȓ:�D���d� �Q�mơ�ȓN,�KE�H�<�0�"*�|�ȓ�α&ߟh�t�p�@ԟ!8Ҡ�鉷M�~��
�fNH�n#�Z]�i?Pn8C6ဗj�FC�	�xT
��􏛑<�D�X �ŗ,kC���`6�V�I(�C����B�Id�Z�`�#d ��^���C�I	�!B)�6&&أ��<<2B�	1$�T�����\��̂�e��C䉕/��iuH_� $�1��>	�C�I9Pv�:�U�I(x����0DzC�I�=�"Vܪbep�K֣�a�B�I��T��X[��2fiԅ:��C�	��F��M�>E��:�cH�'��C�	��lX$H� �)$�ʬj�zB�ɐ z�hp���=Ghd���F
nDB��-�&"`F��l0�3��+ �ZB�0�$��H��p�����i�n|C�ɹ.w������0p>��Q��V�8[NC�I�h�Ѣ�=Y<��!AmT�UZZC�3=�5��F?�F���s�6C�	�!���[�g�8���[Q�Ԥ	�C�	�&u��*�E�H���x����b#�B��1�A�0�V9X��d�%e]=x�B�	�]V=J��ѕ�p �M،L��B�	!Pu�yP���f�ba`t��U�pB�I{��� +�M�z9�U�̞$;<B�"���g�P	�2AK1o7�C�	+.�3�nD�>Q*�@��8��C�	#txص��=%'��Xr��
]'�C�� ��YH%N�8,r��C��C�I�v�^I:���bU�]p�	y74B�)�  {�!J/)B|�!�XTR�0w"O�XTG͋#7d�HR�+]^�G"OhAP�.�7 uz�H!� ���%"O.��
Q��e�1) Y�f�z�"O&��7��0a�9xC��ɪ��c"Oij�D @��[�!�'I�8P�"O6�(�K�!?�ě��]-���5"O�����6%&�����i�P+�"O��oͮ2��q���K�GX0�F"O���<w����Ɓ	*p^b�QW"O"\Pw(ͦJ�Q�� �Qd�S�"OؽFk�4�恊��W�'F A��"O\�"�f�2��I���$$��"O�!a5��$k{�$��Z�O�Qz"O$����*"h��qԎW����I�"O@ XG�Ø�0���+����"O�P����ݶe*d�Ӧp��h�"Oz�C�.M��;Q��('0HI��"O�h�� Z�:bb�Q���X� �u"OJ��/��h�`��E����E�"O&-�4���0��4����.i�>�sQ"OBTx�c_�>8PZ��ګxd�Q�"OHd�u�ܗc�4��Ao�B�� �6"Op��Q�۸1O
���N�1��}ʔ"O�*�N���r�{��ʬ�Z��'"O �����]�H�cю�}�<ms"ONX����h͚��*L$�!��I�8|���%��TT-9��]�oq҇�X�[U�|���<��U��JȕD%ƥ0�6'�B䉦#W ��-~8:�f�+z�On�x��`�(4A��d�#f&����K�i�x	�G��<F�|2�_4{)��H�!5���`�;9�v�H�b�on� B�[�J���	��䨲�qD@@xP��).V�<A�������rM�pGFL``�
���i��]����F�ή�˵N� !�d#o��!I��K���@�왿�9�&��"f�X�t�f̖��	��o�Q>�����II�邬Y��Eʆ�E�Lf!�1(ƮI�ж�YzT�#LВHp,X�aӦx@�#L�A��T�Ʌ������'����b�.`���#3h�@�r=*
�i�5(�5z���+]k����$u���h�-�-C�ܩ�V�]�O�xͅ�	�E�z95,C�um~y�0�Z.?h�<�C�@�n)i���venY�Nڟ,;n�R\ws�D� -�_@ĩ�Mnf�M��'WNcB��� �zWʌ����wń2 �ӑ耮t������|PB(S8���$�!U�P @t��6J50)�"O�%�3N»>��<C�+f�-RT���9�4�Ӄ�"r4��R&�� @>��vd��=9掐�H�<2�A���"mx���6bۭa�Yc��P�]�<�DLW���*ƮY�B�ջU.I�I,� -Wz�z���qh��tnκ-�,� Ř���O���+��vx��A�,Ϊ	[B���K���@�:f�\���aR}t���Iu~d�s����Js��h���wI|y �j<bb`<�'���c�˂�Sg�-cÃا=ML `��{�'e@��V�։I�8PR��C�2��'�J\��f����zB�B*F�l C�W!O��1�faH� :6�:���1�r	�d�߲m�,rb�ª���P'r��y�����FLU�Y��z�ʊ�9��D(j���?y�ثk��8�q.�3�5Iv��>��Iq���%B��[�`�>�c�MP�!�8����}�'{��� �0H�O� ��Wj�g��(���ɇC�dj�H�=W8�ӕ�Q��Q���#j_���"�9%V��#��ĸ-�v%��)}�sB�<��Z�r*�Tx��.扯_�T	X6/�<KK��A���Qʓ]� �G�1MlR0��/S���e��dr����zם�t�,��Ã��z4H5{��ѽi���ɟj�ہ��W�az�ě1@������I Zj�Z#pD�9;4�J6�,�� ��2+�h!D�C����-�V�!�9#ن	�c�3���B*�������t��@;�#����]�q�Bpo;2c�P����]�uA��(��s����z8j ��L�q
�r�O����CA/b�N=��]�T�#2E	5�d���ɤtJFu:��	�'�f��E��	P�(P����$09������1m̥��Bo�mJ#�I*}Ҁ1�V��P�,RCF��&�(�"�p�ɓ(�R|)��3A{`ʓUKDQ�� �������r�4Z��Vl�	1Dsl8�Yw�51��lB(V�d�a��<��I�'�z}h����<� |!r�V'&n���F.AV؄mא#lqA�F�J�d�����K�r"���$	ƮG�S�<qt��0t�T�[���n?�� ��%F�~b)Q c�L�LU�0y6��s&B �۠nϞ��0�BPy2��U�V*�D��|[�lZ;]��a�?kT����M�Y�џ4,36�����ͫ�ħ_�l8���I�|�����
�'���%/�$�����M��?�`�f�cG�s���ə'^�����)����Q�*�<i�/�<���1}��)�'S�j�Þ�(�I�gD_*d��Эu0��A~A���剷J,�:��W|x���N�pq�L���2Ǧ+���&?���G�sKZ&
��q&���y:�0H��,�Չ�[��|��V|Nm�ǃC(x���bG�X;e�U'x�'F�H��%	r,���)_�Zv�+��J0�AsaE1v-џ�	�	�\�>q�p����;?�|���*��C�M%�M{��׎!0�Lh�^~���isf�1 �)Z�ؠ93b��0h�)Olq[#f�;X�H��|�2"��$;P�%iG-Wk.%�0�r~2�X��LZp�'s�1�1惭8>U�`�\��@Bc'=}�aܸ)�5�����O`j'���:0��Y#V�}*��X8�p�
�/�6!`�g��l���͉4��a9�cC�Hr����� �OV�Xd��`D�<���&Y,�t��ɭFm�邤�R��O�b�i0�V?��4�&��{$�	�'��ZA"G�G\�[���>����O�$��lY+O~�O>�+A%ȵa��Uc�ԁ,.F�g(D����u��(W��9l�ᓤ�&�I6b��A�Q�'�*�p�&�GL\�9�͞>	΀�	�'@Zt)!eѶO$����bD�� �'{�Ǭ�v�L0���?��M�'bP��,F9
.4���V�e��d�'a�1�0o_2�s�KW�X����'����
.H�@�d�78Ɗ��	�'-���E�P"D�.�af+1欀�	�'���h"��\��@�s�$ �"O�8��R*���`�,P��"O�m���6R��˄�ƥqֺ��"O���A�8VXT ���!<S|�Y�"O*�:u�Z)%L��T�Āy3"O���7��+D�\� `�-P���"OF=�)D��H��V�9�>H��"O��kP��MC��� c�8چ��#"OX ���,Bp�"�".�R1G"O�D��H04f6a��)qs��@�"ON):2#�3@n<���݌SP�d�"O�u�6��*a��5{�-ٯp^p�"O����oA�1'F��@^*D�P!P"O>�H��^�S,H=����>Ա�4"O~$����/~"��fƂ�E�< �"O��SaI�K,°ڄX�I��(ܾ�6��i��Y�\c�H�6�� �P�H���	4�-D�k�OַV�k�F.��5��ͱ7�bqsH�g��|��]�tʷ�GI����V��<	�/O;�d-1e��!����>s�r7�i����'�~�!��D�X��QٕzI�]Ys�Y/C��)��(��F 2\���('�ߵ�H���H��Q�0�z�Z�E)oj�<�"O��!���u6�e�I,gL��1�Q���{'����j��A9�q��'J*��%�@�
��%�"#@�+�d	p�'K.���R<=3��fE�����a"K��"ٓ�C�mA\��1+�h��|*�*��R7��Qǆ7H��`E�>O���-�>?�i"'��*)�6[� Ǆ'��[e�=�x"3PwE!򤖏I0�R.\�T'P)3 \��	�q^X�xńM�qwf]�e����G�$O�)8�� "qO�f����W��y��
�}�&��è��A0S����gOC9:�B@���[�"mI~��y"��c"���@�Ӗ�>��FG��?�^'`>$L��Q�o�,�p
 �6�`6��FAɀ��A	ӓ/0��7�E�Cs��A��3Wj�G§ށ���"��a�t��Ċ|j5Ȥ*Q'L�Q��Al(�Z�"O8��Sb҂
�fx��$���<��^�p���ړx�\��ʸ������g�π ��a
�>DΖ=q�$�h��Tx�"O����J��߬l�5��N�ĳ�
މ�0��m�'Y#��`>.��O"1OB�I1AWb�ۄ![v����'{F�aQ�Y-�����ȍ+y�Ȱ��C!dy����J�=�Ș�)̻i<az2i�&��}�r�7|˒D���-�0<Ivo�� ߬�V�˽#`�����g�,���I��2LD�һw�I���`��#͆�+�u#ӏ2P+H��'V��f�`�N�0A Uz��D��l��7�~�K!���ty��D��y҃U9f�P��!�){fV���?
5L����$+ �D�RK�ᓈ�L>)���j�����ʹ)f���H�F(<�ō��p�i��J��=����Pg�|�	��[��=�D�P`GL��w��?r��K�OCX��j��}��5r�(�����+��b eJ�ju2Y�*ݾ�y� u�"EA�=>���D� ��'<:���$��
DD�dD��r�	."\R�-_��y��V'[s�P�Cl������Dt�%���\ܓ:Α>�^�`��2���q�:�ӱ�\�|z ��\w����͇F����c,�:_�L��ȓN\���2 ԋ��5�ɘ}����m�T٪��؞cAq�h��������!I��эlǮܰgj�}5
���ڜ��w���]�6T �J�<�j��ȓM������M�=pL�&��݆�XH8!s�#�$-h�(��A$) ��\8��0�&L�}�)emU� ����IN�{!GG=#��Y�HI�3HB����bգ�!�%�����: ����)�9�� Ͼ82��7C�h��V^he�U��1	P�Q"r�W��Xd�ȓ!��	��G��!$'L%iż9�ȓ� ��Y�;��6�T�OV2\��'V�=�`)�54�j���i3C�J�X�'a<� ʎ���
 �
���'���3�X��u�
����!�'I�\�Ձ]�MC``4\+��[�'�c��Ho����	j��
	�'f\e�X����̎xe����'�,{s�U
K5	a��вogQ�	�'��!2ֿ1�~�c�lۨc�.���'��tjP ��X�.�!3�ޫ^��8@�'�v���M�*ffNt�CN�Snd��'�B��e�>Ev�sl����I�'Q|p��4$k`9���X�F5����'�ruq�`[
�h�Q�.��7j�y��'\��i�ρz�^8s#V))U*�'���s��]<,� j'�·$g�Ԣ�'�� �d��>����6��WC���'��q���Iv��LiX�'S�@Ys�!y!�U#]"D� 4
�'.V��,�氱�4l��Nk����'��҉��L���H�6�Th�'#���dזj�R�J���7��U��'�v�ʇ�Km`|S�iH�g�`�'� @F�1�d
�(�Mk �a�'�t���ֶwn��@�ν,��p�'�8���H�'D�@g��v�#
�'YlE{0��>. 0d��3
!�`
�'@p��
�H�T��4a�� �8��'�4Q�0%T�k�Аrԋ[.�Z9��'���DN�-F.�+VfU�J�'Ԛ� 	�Am΁��k9�	`�'��nJ;���C0�J�<��ݘ�'���Ǭ;�Pp[C��2����'�r<s��j��`�"��2�
��� �A�
�qIZ��G
��'AL���"O�����MR\5�P;
Nh��"O<�����/MƬոdF�J)d�h"O�t[bgʀ I"��`�-+�x�"OX-xP) � _�X�@dU�7@�w"O��	�2�yh��W;�@��"Oޘ��e�>&��c��F+*��`�F"O��)g�3�ne��%�Hc^�8�"O���E�*����'��9q"O�5 _iW��q����P��jP~�<a��˦cX�$�2��mqo�t�<� �	/%U���g����#�_q�<)�
�5/�;Ą�f��)P�/G�<�G�I�\y�́a�4�cA�<Y�Ɖ#2��I &䝴0:Q:��|�<iA"̫}�A���7��l�΀x�<�'�čn���z`/�@S��	e�|�<���RK�,:(��� �D�<����T�\[�H?�\� �B�<Y�*@�sI����ǻjr� p��U�<!B�ObA�֨_�F���h��L�<y�!	Р�hх��l�v�<7��0�,�J,ax�3�n�<I0��*�|lsnD_���{#Dr�<9c�"����+/hRT��L@n�<��O��?v8 �4d-ǀ[��So�<���\1F�Ll�k��x�ıå�HA�<��X�u�gd�*u�D ӑF�C�<�&W�V�87&mv�c�&�S�<!̉�pT�H��n��2�l���J�<y$�Ϧzr&�����N0�ݠ�Z|�<I'��`����C9�t)�� ����ppH��9J:�$�"~F�6鬉a����X����=�yr�y*��Z$�*?Z4��L����T�"�^MЁ"A���<�1' 	d�����l+#�U2�o�t8���	>^�`�9bC)H��ɱ�MȘdta��H�1�2��ēAd�YC2��*O}�9���"�b�Fy��En�q��+M��vd9s٫5s2�8��#x��C�"O�DMԌ ��`�7DZ���Jġ�c�P�h�O�zD�-����2�W&t��M�r�I"LvxvmI�y�a��z(8*�Ń�r����P�~ba��+��PP#�.�ayѦA���0�$�%fC���#_'�p>a��H�z��u ��*�]bUdL�T��ԯ4l~��	�'H}��ϛ]�pp1�A)1o>a���M@U�AΙ^�tb?ɐ!�ھ���C
��`b��3D�tiS]�E�- �\ �C��<M�u� R�T�
*O?�d������Д=�T�H�l	�Z !���N��d@���z���+~9�O�-��4�j���` *W�h�ɠ�`Ϳ:�@ܳd�'�DԣDM��K�4�H���(�L	X���z�<Ћ�"Oh�������{4n��mK�Qk �'�H����37�V����$x�T.�
ynD�I�;B�XX���5��k���`��U����,*��F|�&qYC�&�(��O���ia�	_�BըeL�Q�r�ON��D
,a����$�r��Ac`�T�h���H���]5�{��F�,��!�h��s��O��	��D覽��#�8�x`� ��c�G,��ڳ��"w�J�҆��E�\K�"���<J�JĪo�~�j�@�A"�x�񮊡p�Z���4���f�9Z��D/2Z\���?%B6i��Ǵƣ?aQ��H���p�E.� @xKv�	3CL�"������ �
�{6GQ�3;��pbI��y�Dp��8�C�j��c�ЂŔ�mMr��PE�>�{��<ف�Bt��pk4�ݾ. �HQ����$TGk�@���� kݑC�T��b���8��������Ҡ��c�d�Y��'7X:��Y0�#���8D��A�"�E��]q�#��`Z�3d-,;@,���?�ݠl�,`鱂P�($Z�8��Z�0� �5�[i��
*#N�T�.X?h37
�'�S�g Dn���×�s�P�(BAO9fzZ)84�K�^;`WZ�4�4Js�7� f�@��4�I)�!��$|@�W�	��d���*H��A��(Z?�m�2�o����<Ǌ�1
�(G���F�ќTE���W\�L��6T��B�>�%-��2f' I�`�w�ބ<˓`(I�ߟxZ6��D�x�3�l���E�O�%
`����6)�҉O�:�2<���*���6O� �c� mS.�b��!<O4��DE,�<JR�ݐM7E��%���"1�A�%V�����J_(��l��.���u�Ij��넭G�nk�-�S�E,/4p#�lF>�p?��o����MYw�O0h�|m���@k�$@Y�tG���X�d� $A�bU�!����#�ħBʲ�#s5D�@#�F M�u���U�'�V!�X>�&>*wi�pW]q�gA'z\��"�N�!p�Rc��Q0q`��O�	\�AU��Qȟ�d�>��y�AƝN�~��L�6.��uH(}�Մ�2��S�O7� �C�_�,�J}h����pX2�'��-���U���� H',O���.�Ew٩���7faR��k��C5h
���`/��4m֝�;AF�1�柄d+X�q�z|�Y�b/2j�����}����+T�D^xQh�&'���1�S�,�N�[L>��/�Z�dE���O��a5�
<�H�Cf{e��e�'�WƎ��c��2a���<1�e�O��p��g�#q'B��ig������u�Ds�O?7R�<�ʽ9�+�>i���Gg�?��I/n+�f�KH�S�O��!׾�E(��1�Z����g~B �.g`�p�'.NPPn�8i��ı�K%_<�1��$}BmǖO�`����O�Ģ�� ��S��"CPv	��Q�]dZ(�
��+�1���D$\rDȱd��.$T��[d�Q�'2\d�e$�O�9Y �V��A�!eT�1jB2��� Z`�EXw)ƕP�O�d�,0�P��U�V��tMi�'u��1��+<���*��:7pX�O����v&l�O>հ J)`�҉�J��gr�d�;D��p)F9S�&a��)Ȱ7  ��+7�Mȅ�'��y���Pw:)��� ��p�'�Vt���5��L $qZ�l��'dv���KT%?H0Bѣ�_�hQ(�'�J�;P)
c�|l��GD�~�P�'���� ���1|���Dƭ�%%�W�<��
�(X�}iSL#0��iS$��y�<A�^�>4c4,����a�I�x�<��섚\\��YS�Ԗj���Jh�<6"�H|��a!��in�E8���N�<���:�,�����<�D��`A�<)Qըh����`���.��D�B�<1��ܫ/|�9�!�5oSfx�q�x�<�F��LZ��E�D/�6��AL�{�<�WξA����Ɨy�f���"�}�<)���C ��K���E��{@�y�<!�C9E�xr��[u���f�r�<��($�:Y�_�EZ�j{�<��;,� ��;"4%J���X�<1�O�>������A�:4H1"�	Y�<I�� 
r����l�z`=Z�gNW�<�&F�rd��h��:y�b�Q,�S�<1�i	�F�Se��4}�����@O�<�t'J�:]x�ǰd�DuɄ�P�<At���fN�+��׭Dp�l�ƫ�k�<Ib��B�(���+31p����x�<�&bH���"ή:��MB&�B�<y��_3v`n�t��.iL��z�H[x�<f�#y"&�B!L9��|�<���ޭX�%3����l4z�y�<Q�%]�Ɣ v)R���\����v�<Q�]>ob��GG�x�.�ǃ
q�<A��J�z�3����N����7kXi�<��ٶ�����$2��(A��i�<Q� �[����Z�j� _r�<��'��ҹi��!#P1����m�<�F�3ڹ�6�հvA4XK��d�<0/44��`3�
p�z��A��f�<���4�b ��&�vD����J�<� ��
G��!ip Y�s8�'e���N�KX�h�b씎!���0�L��;�d��F�$lO���%�ԭp�*��#k�dḊR{�=��@V�$�NB�����sI�
8���	�#T���� �A�_�h��V�o[<� �L3�4x5��1J�C�-��D��-�39Fx� 瓝𚨀R�M6j�6�'�-E�,O�P��1H��U�䃁�wt��0"OȌj���j:Ȝ�g�ѭC���C�L(tx�|�f��}�a|"!��c��M��+>k�0��T�G��p=�/�6
�*=؁�x�9t#F&x�N�B@�Yu�Z�� a%D�T{��Z�5<~��х�X�ٱG-��ܸc��F�?�#2�U5Q��8!�u��� 4g.D�@��+�ʂ�����2�x���6
��y�l(}b�B���`:z� 0DX�v`x�B�Q	S�!��z!Y�P鱴��9���A�_b��U��JZa|�̜�K�l��L��Uʳ���=)�)�4H|޵�'Q���5hKz1dL��g�"�¥�	�'��a���-�%��-O�^�q���\+7, �G�d���'\���bƖ4�|3!��!�y�H�������* �M�y�*߅H�!��A�v��Bc�L�<ٰ
�4=������O��qI���}�<����+9�R���,G�S��а�]z�<�D��!"�\��L�[��0Ɔr�<a��>l�	j��ޥ5[��P�)�s�<ycOZ�[	�e����)?��p���g�<�TmG�~���CρAɮ|HN�k�<)��&v,�AV�@�G�j�c&�	{�<a�JR>lTU2i(Φ)��oPq�<�R�
�V=�bGDROĔ���g�<���`�j0Q' �#"R��t`�E�<i��D����J& �D]��NAA�<I�	�l��-y`��&�����d�x�<	"�X9*1A� :Z8�Q+Ʃ�o�<Q嬘�/LdY�alL5~yڭ��N�h�<IW�`op4����7���D�R�<A�&	~�
�`G-�0 ���T,�u�<y�s���;��Ev�s�<�A`_�v�B�i0�P:(��Ӧ&
`�<qď�5G�j�q4��8N6np�`.�G�<���O5�B�PA��ED�פA�<9ue�9�@d�ҫ�4��ax��U�<�u�$�j���*���"�Q��4!0��G�L�f�-T">I���6i�	�k�W�  ׄ'D�T�!��x\�uc@ꐳ9)���Dg)D��i�!:��	[���/�-"sH#D�أ��˷%�
��c�x]F���g4D��A�F�(g.���d�(iZBIS!.5D�B��=�V��5�V�Q�EY�5D���D���;�p��%o�`���>q@��W��H�<EcC�T�M��hBg��X�,��imJ���R��@(O���T��DI�W��7m�(h
���'%U�]�M����z6����oӦ�"�����ԧ���	-vm"u�AF���q��e{r瑦R�"~*2��I۴����R�@:6휖"B\�Ey��	ƻ"���AI�1�@��_�zTQ�P�W�O���3!$��B<���gQ�7^-X�{��[���'C�b�'���b�!��U.1�O��ڋ��i>a>V4��g�)|l�u2'�����5�hOq�����r$|��E��t�A��1U�b�>�O'dc>a0 ����)���=}O8A*��4?�CO#{��t�D�/}�𩈣s.Y`g�ϟ'���hL:5��f�������$P: ��)�p���8t�\&c<�y0��S�L�G�^C&�a:6�s��8u�{>U��O��~4�۱�̥mE�3Q�X�&��W3O�X�F������	[�@���mI-1^z)�o��s߲a��hJh���kY�������� |�bR���Q���]�Ƶ�3�'Čĉ�.�_�S�O]�\�ə|���1���,!(N�����5>���|���.u�`m�<Z��hC����(����{���Ipa�DL?,�ر`�`O'h|�z�̉���i~�r��)�)k�.��R'�L9@�)`D�9�PB�I\M�x�!GB X`�l��FCBB�ɫ8^�:)��pW�m��^�lB�	=�P�B~�������b)B�I�aqrk�G�>[N|��T/�)P��C�	!�F���l��0�'��_G�C�I�e�$�¨�<����É5JjB�	�C�Ҕc�g�>��t`�R�B�	}���'ŏ)��5�ņ��c`B�	�{ǘ�ٵ.J%B��1���\~*B�I:m���W��O�h���_,PC�I�%֨ɐ��D�<@(s#'�3/"C�	kB`��H;,�$��	cUC�	~<���r�E
?�P�aQA�|N�B�I%N�<\@C�O=p�zm���=e0xB�	:p� 5SgNӥ/��<�q�Z'{�0C�_��}Ad
iF��w�Y�?8*C�ɣ*H����*�J�8�&>@5�C�I�_TQ`Gȓ�Z���Rӂg��B�	T���e���,���,]�OtC�I9~���h��C����T0DC��zJԉWΑ�H���b�;J�@C�I>#D���H[��"Se��e�RC��T!<�5K�^����vՆB�?{�9�� �4r0��*U��B�	��0�"c�|��A'J�&VrB䉒F�I3K�I�j�jpe@0sddB�	���躅	3~�L�q���}S�B䉫wY�Hr*߉k�6d�m�1ѴB�I"g��K���"u��{b�Z:6<hC�I����n"��]�1�vfC��t{���W�ʎ$`�QqE��,4C䉯F�P�Q���pi�p��?�LC��&-�` �Mϊ1�4٘���y�.C䉟^-6�@�įq;u #��dIC�ɍY(��0�9O� J�ˋ��B䉪]_T�p�� Wm���q�(B�	�H�S!��[��a�4o�(B�	� �x	���	i�0 ��6q��C�	�0�<�+�J��7��� 1j0fB�0�t� ��5R{�ݫ��P.}MC�-"�B�)[�ta��b&.��B䉺4Q��Z>1�R���[�|N�B�	�@=�@+���1XH%����?wj�B�	3�ޑ��N�J����/��B�I�\�B0�<P����g��B�	%�l���ɾ �n<����1O��B�RE��A��T�mJh�4�̬w�bB䉘E��e���_�6�"tÅ@L�C��2\��Aq��>Zjf�o�|C�I�L
"�jq#8���)c̪	KFC��''BF,IǠͼ'�z!��\g-C�<G��9�$Q�v.��� \��B䉸*�����X5� P��M[�_q�C�	�H�T1�H�@�� xT���d��B�ɪJ����%e;aoL�rW. �y`B�I�ӡIW  ��P��X|�C�	�d�0��c� �g�`���ͣM{B��sHI;�J1�T�*���qi B�	2a�^���/�!7H* �u�yC�)� �yR0�/d�ܥÂ�m �!�V"O��R"_j�&���'Șz�%؂"O�P����S�"���f��.e)A"O����g41t�I�rE�h�nTAp"O T$JӦ9�2���#��X��"O���H>u2� N�T�T�[�"O:��d�^�!X:�Yf�ɀ9�P� �"O ١����%2�����r-R�r�"O�yB����N��#hԴ^����G"O��Sm&`:�b����H�"OXMW�E",�sg̉�U��@��"O6%�%e�(^,��`
K�H���%"OV�IPB��@�4lkd��1����"Ox���K(2�`�ڕ��JV�`�g"O���󈄫#r��gk],n��5"O��#�in<X˂���*���H�"O�I��_=<��aJ��G>@���"O�LYrI[�#޸�qe��71��98�"O�<��%�[�D��eЖ? z�"On�#r�F�hH�Y��^34<��"O(к�lZ]�Xq���Ĉ�6��s"OԬ`W��0 tH�BE�J�F"O�8����%<�z���12jļ�q"O@À�ƤiU�.�1,2� �"O����ѯ%m�BV5I�y��"O�	��c�/f_����8A��z�"O�H����*"+�9P�"���t �"O.�����E
�9bF"I� Y�V"O���*@�LƖ��!��zW(�{�"O��x��c~�����0c�l5�"O ����v����C�X,�1"O���Q�)I8�X��-5�4Ń@"O���5G�o�ųe�u�j�"ONXv�״_K��;��D�:h��Y�"OB8�6 ȷ)s��"�(�iN�j"OV�Y�S�I")e�̉o\mC�"O��� �0\���T���:8�/�!��B� vЁ#��(����!��a�tp��O�0�ά����8�!�T��:,˂L��	R�I�!�$���<���@%h�HDФ(װz�!��*��)��̐Z��cQ�ё@'!��Ê|��L*Ā�7b֌�Q����/!���)~�ˀ�Q�0k�>!!�x�����C�I�RA"P/F!�zKnl"�}$ъ6����!�$�14#��X�!'8b	ru�P/C!�$=
T�x;j�6Q0|��ߩB�!�߱��90��.}��|A�4�Py�E���x1�N��=z�z@Ԝ�y҃
9\����ǎ�1Ҧ}�m��yr� 3J���fލ&�%����*�y�+,� \�%�$�:q؅�
�yRQ��	�L1~Ezu ��yb+ػ�2��T@�p��4�I�y2�P1m�P*�G�r�YBT���y�I ,?����8Yu�@�C+�y"�@ �U�"�$XZE����Py"��,lF�#�E�Y�������S�<�d�N#!BH�EK�5��e��@�M�<9���]��β��X��K�<Ɇ���W�Fux�l@+6����O�~�<�DNY.`��ő�f	�K�z��I�y�<gH�B��9�,:j��YrH�L�<� �����((°b���#Z7�I6"O>=h��
Y�!3WjY 1>�x�"O���E��:�4�G�!Z'$e5"O���φa�&E���!�m	�*OF|�n�T��%)���K�\X�'A�ʧJ�%)8Ȱ�Ƒ&4~��'�����W�`|������Q�'��x;�@�l����g'�	
��d�	�'�l��ЃZ�V��4'�6���S�'bh�!�ț`x�I6+Q�0�����'�q�+Ee�� z]V(;�'����J'5���lo	���'�`%��X�ڔ��Ya�����'����`j������
T��� �'< yk���:	#DD"�K�0��
�'0�u��$�K�H��B�M(�o@M�<�wb�	Z�dd!��6]�*��T��H�<�4��B)��g�	;Zk5�Ec�|�<��B�T��P�s�C8�Z���Q�<��$KA:�Ȓ֊~�X\	���N�<����p�=*�Q���|� *VL�<�7ˉ�9`�S���Q�O�<a%)�'r�
�aٛa�r�E�<a�搐)x�1J^�%V�II7̀Z�<)�I�k4>`3%�Tp��� d��R�<A"�M��x'��R]B@iqiBY�<�p��9W��a#���|&�}�s�U�<�c�AD�%�b
�+�� �MT�<A"��*��#���#9�l�k �.T��K(k��X�ժЛ_G�Aڶ�(D��p������ӑ˜p�]I��%D��Z�`E�~ia;��=R����Q�#D��ZcfY���;�!�	v���s�"D��S�* <K����JM2�hj�#D�hy�g�u8xͰ��	+u��e�?D�����."�&��B$ǔ�y2�=D��!g@G�Eon!�׻2�PH&����yrG�0��D(f�ը~������yB��c����'
�R�)��X��y��˟��� ���L�}aa���y�`T�b�*$sR�Ĥ"yִ
1���y��4:��h+���I��I��J��ybnH�¥
�;E��ݪGƑ��y�#Q0�S

�{@p���0�yc0%ṑL8_����i��y��uE4*ޔ�s����y� �*`��d��-HLQ$%�.�yRk_wk��S2b�̄�ق���yB�:�xd���򈫂�y"#�i�`$��O9|����&R��ybܺ6�Ќ����,��X��喷�yRi��R�p��8n5L��r���yR�I�q,�$��Q3p�@��J��y��8x��dyV�ȝ<(��Ф��y��Ʉb �BRiH�58������y"i�����k��0�q�/A��y�G>�͐��[(�5���E�y�ㄧs�:I�v��Od���ʟ�y2��-�D��@��I���(�*��y��"^b����؁luĠ�	��yg�D���C�ǘa��!:�	T:�y�f&|�@A�F�Mz�ލ�y��+eR�m�.� $y"dT�y�%�|��Õ8Q؄�q�!�y
� ���/�F�b�2�ʃ�O�a"Oj�Bb�!M��$��k.pֱc�"O���,�%F�`1�� �Rk��"O��N6al��S'�Rbj����"Or���B+K%H��BFU:�j#"O\`QA�3k@q���!oҔ�"O�m"���p/�]iZ5V�!"OX�j"C����E7H�
���"O�b�	   �