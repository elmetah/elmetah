MPQ    (>    h�  h                                                                                 H�I=��
�`0j����nş����1��!ON���c��f�;��,�>����]�0��<�I=������$��K#�()��G�Gu�ӯ���b�ڬab7-8_�]6�@H�<J���f��6��������L�����=�N ~+-5�Uۿ���D��q'G�xӴ"0��s�r��	�儣m�*�	/��l��S��.kw���/c�*��������̣Z�$�¦��|ټm��tHP��_>�����8O���ϩ��� �-��*ϸ2>�q�>�]H�E�\�����_�n����Ȅt);-����f�3i��W���~~��ͱ3X�ƔP\g6HZ��r�(�dU���
�T�Wҫ�-��>shVpj�&=r��Ҝ���?hF���ްwq��BS2o��s>���|���ԋr�V�oӉ�p� ��4��52�~JG���&#:�[�����	hq��@C��Be�'���󑰯d����W+_���~x���높~G�Hq�-T-ys�|�.̳5a96�}� ��9�
T9"z|�dx��Wl��3��a�@+�X8�����<�i��Cx*�����P��|��c�i&�S7�,kͻ�u�o��9��:U쏐�=���	����<�+/���}wZH6L�\�4b,�T2��QA��PӍJ���%fU�(�~q�(_v�Xg9�>[K�n@\v����_A�-^�m�����"��������q|27���p�9\��,��}�}�zV�(�.����>�X �cs���P���1�����4�S�jK����ع;�����+]!�B\��Q���v�S�o5�
.�Ȉr�F(���nUP��w� =e�~v�w� ���FK�3��P�v,gִT�,�\�K�K����Y�l\8j��҂�9k��L�� ���_�,g�b��x[^�z��%-����}�^���VR�X�A���9�Z#W=�X�N/����䨀fA&�Szõ��)D!�KB�<SZ�2���<�Pܑk�ĺ3�:xD�Px��R<�A1���P���H.69�Ơ�R�s�#���kWh�&:�cd�e���Z>��2q
�f�u=��K�2S��ts��g�m�CJ�B��P.��(�h@*�'��h0�y�`���}O"�Ȟ�`��o�H�9/�ra�L�t<�����J��TI��e�'��$�h�
�ٝL9��?Jm��9�jYxP( /� �lIı�+��Q�{Q`p�e�6�vvR�8�LT�������g/�Ǘl#!��J�!�#�=��̟���2w��0�A$I��r�R�Bx� c��:ړF���!�)僻8Q	�߻N�rQ$/�Z�����������y$�D\�ƞd)�^+[P���d����g��������c������@�N�;k��k~/e�T�v:<�oN&l�V�ĥ[�b3��㖆�kX��������F
�5/(�9%|qc�z:}g�.~�Ժ�:���m��#��qj�%WB���ǊK�3=�#��H�b�*-�f!~���ƥ3��3�/Ŝ^�s�����净v^0�EF��
Tfl�Rʤ�j��r��:?����{n�e�� �7њ`�Q/b37��&ϱ���#t�>5��ց���v�d1��go6#8it#��6F�Nʸ3�����]r,c�*b��BL����J8wF�S2q�C�`QTS8"8�:#�x�q�j�����$��Qy��p�K`���>?�0fP�L�羅z
&>x�Y�uR��h��5'�.H\���O���+�� z�[8sx���X�d(AaX]p-d��t�#����Hb ^����L�T�$g�C|�����1��M$��t��ک�-��!4��'�R���pR�No������w���_W�9pf�H>=�Ơ��^^�� �uk�O;��^ȍ��+�)1TY���=�	���%�K<��Ԫ�Y��4�����p"nۭ�)*0A����P���"m<ub�Ήy W̏��6���mD�k�{Ǿ`�^����X,��~��������ߒ~���5��~������9�ܳ��j�=������U��2��Mm	\�3Z��w�Dv�c�_��TCጩ�&L�n�� ����Cȗ�]|
��/��Rd˴�b��wz������\�
�ϋ}P���h+�J3"pB��rJj{%�����olРl�NT�V悐f��L����w�"�F,~n�N����2 ^�6��\��#�<���:��>Re�R��,�㕃cqu�d,�p�d0H�PwJj�����bc�ѭ�&�ԾI᐀;�&��O|�O\���L�$6��2i+�^���0-])i��*0��l�&C_�};m����H��E T�8"�S�ս��q��"�
a��Q��X��&�w��'���Q4���ݱ�I�iAR�q]�X��ix��@1��KD�;7���qD�bZ�" @���@���̭�]9I>\XK
��O�sn�B.0�Lp�d�N�#Μ#k�BYdv����p���5��Į�$� �?��,xSt����|:��[��~dЅ�.���}�!�W	0�U����F΃�Q�{Y��ץ�E�'��䵘�<	p��������l��4���������ޟ疹pÐp
F���*��9p�]V���>�k�~Ɔ �D[��=SVrï=�(~��)������b�|e,������HtPNr�{���T��֕���YN������}��è���:5�Cm����=�^�����G��}�+[B	�ݰ(VU�#��+(�p�gnH��=̽�CL���J�z�b�2��$2ŗ�@sЖG¥y��Y�X���Z���򨩂r����q6�4Κ���%h�T_���.�-�l��o�)�FV�y�"w�8�R$��"�e:�B|zK�o��{K�\�L<XyZF0IL2)F�6&ށ0�����n��w~h���|�~75#T���D�����?f��Q�zmjP��~f�����z/T�y�Gʽ|#0�r��c0�j��
��潑u�Y�Jhx��k�~�(�@j���������U�b��?t�@p���)BgE�r����>�z��,,>U(��k��J��������*=��1\��x�1���@�:���V�QT3����8笡D�����L�����;����Ȭp[��uU¹r>�u��4*ӯ�g"qH�.�Ը�q��`SQm_�P	j�`r�d�NG�.ƊO�E��c��t�����޾N$]�`��+�����/R`���O�?k͚�,��!s��D�7��+�7�q���-��� ����E����7������n��kL�?�S; %��D��f�}���r�=�~�j����́?\�8�Zg�-r��&���{�}�̓Oy�Ȁ�zt#hq]�jX��M�ݹ8�ȋB�F�?��J�A�]+�o�b>q�|2�	�&�sV��i��p���}4�!2���J"r�%e.��[��ɪ�K�h,ss@^2B�)��nv��k;�$�R�ն:��xK���+�G���L+�Th@����.�5a���}=���]
��"Us�d���W�k3܂��B@�Z#S�p�d�Z��i�̩x�o��`�q�P]�����i�.��,��\��-��_9#63U���Xۙ��^���w<I��/X]{+�Z����À�O������푅A��.PnS���l�f�`�(w"�Czm�����u�w�\�}��\���-����V�e���V�!��g��2��B�qE!�TM�ʧ��}�!Q�ul(5ঝ�p>�q� �\�s�����/Z�2��9�4`��y�X�o��f�����?�VZ����̻j�S
�[��Cx�a�k�O�`U+%P��K ج�~q�F����WK�&���v�ߴ�C`+��F�~���'�lw��j�z��p4��:nH�z>+��0��W����xv�bz��6-�4�ɸ��ؘR�VMQ��Ԛ��o#r�&�,�N
����|��Ct)fz�љ��۵��JD<6�B^��Z�./�𳎏�::kz�x��3ux�P�P�ʉR��<�誡���a��.16I��U��.�n���W��&�dSc$�d'�>���qe�֍0ϥ	�D�*f2.�et�.�gd�Cݎ���OP�&�(�]I*w���C؛y��2��:��bׯ`po$�cf�/�Uk�'�<��������}I$F�e�-���U�5��
�׊Ltv_?�M#�-�j���(�V �"R?+���Q�?5`H����v��m8�����1�[�B��7��l�ך�E{o!��3=l��̺c�ʭ����$B#n���MEXB��E ՝����������) i�8�x��NH:�/P�u+�Bk��e���D�zƙO4��K��󤟱U�-�������=��x����R�C���n�V�i��e���N[�	����&�K��ep�[
�̷rjT�����:�(8�v����ѐ�3��o�|�q�z�N�	����Ǘ�٣�)�(hM������A���=�cك����;Vf`��M�����3�t���,|^�����I��vY���o��Ł��T�;�REW�j�����wV�8|�{i&A�_�J��34`��b�4b���b]����>0�P��&��1�&L}�g�I�6���t^;B�� �N�ƽ�V�K�Cַ,~��*�BB'��ɨ�w�ʻS-J,����`Xw8=��:�Ƭ�L��0f��9L®s @p�ڽ��7N?2ZA�|L�|��*vE&9�mYE��u���M}��2\�6VO��+�,,z�Ԗ8.����[6�?��aU�p�5��o�z�BH0���<���C拮�$�+'|��F��֟1<�oMߠ]܏���$#Y�d�4��-'K���f�R4I�X���ߒꕋh�:O9�'H�O�ƛ�A^�#� �F��j#��ٳr��7��O��T�"�8-3	;�m%�� �����G���\��i�xۨ�p*��g����k�z�Fu=��	V* �Z���'6h][�(�@k/�,�9-��9��0�,e�D�ĂO�A�����������������������س�?��9Y��"
��Ԉ��MH���nGD�>�v���3кC������kn�6Ьõ`�Ǳ�Xod�Pc�Մ�d�	�bL�8z}�����=��ыx��P�1�\�p]6>rŭ~%[o)��}N�;BNO5���8֨T ��w�EF������^s�^�)�g�/�vb%<��:�R@G�8��~A�cl�<��*�pO.�H�QcJ�9G�u�R�j�lġ&��c��
��
Y�rOO��4ze�\W�-��$ 6�m�i�)A�p}]H4��h�*�Il*l�__��;hi��6��H�1� o�"Y�՘��q���\*����s�-X��Y˒�h'	Au��j4-uٌxtBD�
A��5]r�����̌޽`DX%�7H�l%~b��' ������<���-IV��X梁�J�?nJno0R�֣V���I��w���Rd��������5|����kڸ8���Z9v��w`u:<x�\+_Р�~�t�օ�ǁ!��0//Ԯ���F)0���{tg� �?�J��5�<�ML���O����g�OC���6���L�ˆc�1i�Ë���i��Q�E�ت�o]18'�ya����u�r���_�Sqb��Ө~�S���q<[�w��Qv��c�tk�rs�%��b�_}�2J������a1z�8	J��ł�s�5t����J��y�^�`����ĸ���+v�X�!V097��
����nCLա��S�ɳ�L�5�Jk�RbyA�_b�;�zs���� ~�����X�y�ZLZ������gS�9h�6
���ՙ�i@N�V�_ JM.Ӓ�lҘ���FQ y�|���<�$-�"ky:t�|�VoL6SK�"�����X4��0dK�2�c$�ᅁk&9���B�<,��'�hC�,ۗ#�7��~��Dس������D�Q>��m%�������rÜw�oT��Geq#+��rV�0��)�
(ƽl1`Y!�]h���]�~�Y�@%E᳴��hl��0'��tN���ֿ�)��	E_Z9��I҂<	�&k,y�I��R�fn�JD�Pq������k?/��5�1�j@�w���JV
�1!��[�'����Gc���ULjN��Y����������R����9��iKӪ¯"� ���庸��Q��Am:�H	�pP�C�I�>.!�X� .�c�������a��CU$��7�����r
���{4�����R��@��\���VB��U������{��Fk�S�ME����r3J�un�@ ���Ӂ;;\����fy��?����#+~�J	���<
�\�ZZZ�Y/r��T�ڕl�ZԃJ�V�a��5�h�jKj�g2(kT�H���&e�F����f���ux#o��=>Lq�|mF���m�V����hK��a�42�2�RJ�*�`6�Y�[����8�Vh�i�@y cB[�<��/��&HƠ�UtM����<�x{����Gw��'�,T�'I��u�.��0a�� }�3�a{
JGq"0��d�{�W��3
z��o@���n�j�Y8�5�i�#x`��LN��&RP��	8�_\Y�	�i,�1��ӣ���9~�kUb���s@t����j�<���/�ׂv��Z�0Yc��j�b��8��T)A�KP	9���cf�(2�:�^�l�N����0'��\�����h�U-�
� �0�Ѡ�ҭ�"VL#?��2�U�,��o^��"ؙ}c���(�[y��~.>R�8 T��s����F�*��e�ti�4��J��"�_RNy��ի)�!���o=��e߬|ݻe5�
������v�|������U���M� sT~lN`�u��}լK ��Fu�v�&9�ʮ����Aƍ�Z��ϥ�l�hjy&��KO��u丷|���!���g����x�d-zz�S-�����s3�3��VH���,���'#��NnnN�@!�(	��އnfu/��	'��Y+0DW�B�5�Z�J9�+K܏��:ku���ďx�P��R2��d��������.,S�V����/TW^2�&���d����{>���q��f��2$�kA�r2	��t��xg��jC	�����P���(�r*�x���y�шͲ��o���`+X=�~f�/vYa��q<�\-�(V���I��e��r��ګ��
t�L�O�?�N_�A@j-(�g  ����[��d�Q5$�`��V�Զv,��8u@��X��{���.r��lY���@%�!F֫='�����(����Է$},	ք�H�B.� �=��4I�ډC���{)[n�8�Bx�?
N�y��Y����߽0��@Q���$�D��ƔZ���;ћ���¢����a0��R���������U�=ؑ���q��a�e�C�=�p� ���&"6� <q[%�m���k7��u���8�����������|��1z0@���0H��2W}��`�~�������AJ�=Z�پ)�`jefb����b��<3�x��%��^�A��!���svT�`���J�<ڡT�*�R�)�jo��Ձ�Ӏ�{d��ʺ������`�bb)R9=�8���C�Y3�>+Jr�7����,gB�ge��6��t����l��N��#���w��na,�Wt*X��B�'�w|YS(Cr����`�{8XNI:���'qZ�B���Z�{GႮ�cp^�����?��4"�L7��ő�&4vDY�E�u������=2�V�\�ոO-��+�z@n	8����x;���\a���pc'��j�M�m@H���ȃ����f(�$��|&V5���Y1��gM�{Sܪ��ڟ�0�?~4�y�'����!,R�c�����u�L���m9��Ht� Ɩ|�^i$ Z7+��+g�T�C�������@T����3~C	�M�%t#������O�o����������ۣ��*�(.�D�|��sU��}u�DB� ��\�ʰx6�#���GgkJM%ǴƖYn�@'�, ib��4)��$�U����?q��"��!��x�o+M����EV�~�Z��s�(�6M#���T����v�?z�x�uIC�j�Ǳnw�Ϭ��Oy烆S�z��՟�?��d�b�
�zX���!s�@���s��ګ�����2px��r@n%6B�����7NJޏ�8ƨ���^�w�_�F�Y��A����^����壭1�<.��:��R-�?|ʇ�cg�ǲI�p
H�r�J`~��PSę��E���&�P��S���o��~4O{�U�\����Ɠ6�B�i�#�+}�c+C_C2*��le��_��;c	w��>=H\�n ���"�~�sX�q��@ԫ�����^�X[��˭x�'�����4h�
�W�?�A�Y]-z�����6�Z���D��7�&�g&cb�� �)����������I�@�X�[R�Ew'n��P0�ᣚ�����R�F[ d�F��~�7f�57P���_;�1ړd�ɢ����r�3:����=лT7��ў�!�N0�(���uF��m�8�{�Zcכ�Ŧ��d�+�<M�����P�m�:I���1�>��Z��v��O[��8�Æu�&/�Ё�ۨ`	��/��]���4��>��k�=��XoS�r/�3�~p֖�P�����r�ɬ���b�t���r���a���LH��Zƛ�׈�Ԉ��-�p
�w�5O���R�<�s��^�O��Y��R��+�Ė��yfV��
�즥�n>&��ֻ���-L���J��bTp��&��-sƀ��[�9�m��X� %Z��B��t��|���$q6k�P%G�${���)_{^.�l�s�_4%FlEyB�Ǖ��$Hac"�5Y:OL�|��}o��K�S�0�X��H0��2���컝��\L�=�����O��h��۲v�7+p�Y~�D��� �L��dQ���m����ª��ČR�_TN��G E�#&Dr��0ywvD�
t�G�Y\ٍh�.�oy~V��@�����~�6���!V�t�s��ќ�)�?Eb��)������\X�,�!6�a�Jh�����l���Q1�j@'�����IVeִ�Nɋ�0��rŶ��X�6t�L�T�ν��_��\����y��:�o��"ra�I�dӥ��"'IR�%���VP�md�	�	��N:�D�.|��c!�P�jTY���h�T�$�+G��I��͈D���̄+�J�5�$��t�ܗ���z��9���V�FP��²�ζME������0�fn������ȵ3�;V��:A�fTq��zGb�s��~�J�D�����\��_Z]��r�$��f���1��E��Ҽ���?Ph���jN8_K���{����F�K������9�;Fo�>'��|�,��\mV�2��Ñ��Q�N4M�2�U�J�`�'��#[�ŏ���mh���@���B�l�����aD�ZْH�w���x�$�׽|G�#dT�.r�Md�.���aJڠ}�F��%
Ŏ�"��d)��W=\T3ׂr�@\���O�f���jiG�x�����؎'~'P���$҃�9���}�,�:�F���9��U�^���#y�E��<�1M/�r�q��ZY�oU���R���N���7=A5O�P�>*�Ǿ�ff�(���yt��B��Ϥzb�X\G����D<p�-�|μ;��L�o҈M�]���,����2H�(���Ȋ��ʝ,�}>��+#(U�j���H>�� F�s����Ng��/6ܯӅ4P�z��H��4	�Ȕ𲾒���ө0����G���`�P
?�Rȹ�/���[�EIU��A�(�r ��~g�n�O��8�EK;kڧ��v���:�a�d�<y���o݊VZl�0�j��Y�&��İz����!��2T�=����K<x� z��|-����.����cVC�e�Rk]�j��#�����N����c�Z�y��fp�ܙd�L�}�Dr(�BT�<Z���f��!X�kp��Dv�xu�bPɒ�R���?�n�<�8���-.'�mƱ�Y��p��W�t�&�1d��ݼ���>���q�����?2;�%+2�6�t$��g���Cc��S�P_Y(*mQ�����yR��h�V�r�`�`�ә��/�|C��#�<7K&��*�/�I�6`e@5^��	�+T�
O3L�H5?o��ujj2(Q+ ��5~ӵ�MQp(`A?#��v���80ꔫ9�����z��Ul��B�;�!��=��v���:ʣ ��[$�77�7��COQB�@` K���O l��e���)��8"���N��I�����=��8���n�*U�D-T�Ə�~�o@$�q��ի��#�U�<pJ��#�4�+���L�Lh��s��ܐ�eZ�ă���R&}�e��'�[@,�h��F�Sİ!Wn�u�능�F�+�==�|��z�Q������k����:Y���w�޴S�V�S������C=5�����5����f���`��=^3ݜ�[^y�O�>����T�vO�E�%�����uT�9R;�jJ�G�QR��n��{_v��K@�hY�`�xb�����7S^���>&�O֒˃���v�')g�:E6���t�A��ֱN�Bf����'o,�'9*���B�]�?� wv�S#\��T�$`��K8s	�:��8�_*�}bm����B�_�)ǒpXe�.d�?(����Lr��`�c&/%WY��u�v"�OVs�x�"\5��O�D�+� �z�'\8��j����:6����a�Vp�8��e����wH�����xj��A$�*|�һ��֯1�MUvm��I�.��Kt43Zw'��7��#RꝈ�&�4:!�,���9!�lH��Ƒ"�^o�� H!��S��� ��M�ū�T*~�.�O	��"%/�u�ڭ�����o9���A<�۞�R*A������qXQ�u�N� ('��ŷ6
����Qke6f�/&$����{>�,�gخ�_����騌����>��xh��F#`�
�9��Yc����9���3ܚ�A�M�~9��`�H�Uv\��5��0�C2+ǟ���nRP��9s'�N�L�h�����d3bBCz3B�\W���K\�n���A_�{�p�-r��I%5Q�R�n�qM3NE�&��5���l��w.+F��u����ܔT�^�Б����?�<IF[:
�MR�u?�zে��xcb2��u�Zp�!5H�J���+GU��O���Q�&�1��Z�؀lj�㪁O*�0�X\͔��6�7�i<2���~B�=.*�R0l�V�_�3;^ɑ����Hg9 ���"�.�NM�qF]��k����)I�X���e�'�Ah���U4�����Y�:;�Ac��]�:�캠��c�3�D�Q�7~��bGDbk<� qu��9},�2�5�y��I��WX4;�@c+n %�0�p����s����-�c�bdGa���5E���5������ě�n�Nj�o�@�mDN:������ ���W�j�̅��5!Zn�0eB���:�F��E��|{����"ئ�m��f�x<�6;����Ƚz�ɜL��y���Qa��A7��g(CÁX��qo�<M�{N����]����'5�.���.�,?�Cq�S��A��m~Ky��TN.�r2�mp������t��[ri�d�<�1̇Q�h����o��7��F��(vw����5*αэ����^�^z��� �K�+��ɇN��V�`ΔJ)$�A��n9�ҡN��?yL�́Ja9Eb/�&��Px�qtWs�%=¶�ƀ(i-X��ZB�+u�r�3���o�6 ��Ϋ���� ��_�.��blH�C��{�F�&y��Еi��$c��"av:*��|+�;o�{�K�њ]��X�L`0�;�2�Z��Ƕ%��Ӑ�/������Mh�������7�F�4$DNV���y��\�Q�nm��%�� ��h�- T�^{G�8�#!o:r\m04��_	.
��h�"	ZY�P�hIl���x~��@�^$��:�^�#��/�\�t�=E�̙f)S�EՉ��D���x!{�7�,���C��\��Jò�ƶ��+��a�ٕ��1U#�@h��V�������&<����w��q�LU_θ���-�۬��2����JB] ���4vӠ�3"����_m� s���~�m�a�	��C/I�?��.ׄK�v�5c<CĿ��C�d��̏�~$.w�����('��`/)�F$4��XB�e���Ҁ:��_��IK�H���EU��>8�IƹEc����Ǳ����n�2S����p��;q*����f/��,��8~�j����7Ͳ�'\��Z؄6r�yA�PV�N)
�@vF�G�����h��j�(X�J2���r�\
�F�\���r�a�sro��>��|�2�����V���2���}4h�2�WJ�����8��\Z[����M$h]�7@��hBQ>�`��`���|�CǢ�K	6x|�p��aGm����kTVo��r�.�{�a�� }n�
�
@�Y"��dd��W��|3 ���<�@���Fឃ���i�$Tx���������P�Q5�?��U7=�*�,W.x��R��Z<94��U؆+�j��k8� 5�<�� /)-�l��Z�����E��9�x��~:�Ap��P?d���f���(�������D!�ƪRU�S�\� ����+�~-J7�V}����6�c�K�:��R��m�2�2��2�ȥ�����}��f�<(����Ҿ>~� ��s�L/�<������]\4�t"����i�ĸ���ے�મ4�=%.���ǻ[��
�i��tH���Ϣ�r?U���cnT �C�~bd9WJ���@#KVh`�<�dv�fܴ@���扎7r@��#�E'�l��jo�	����0��KW���c����N�+x���zp�-g���i�X�i�XV>����.�%h�#�uDQ�N��|������fk�<��S����FD��	BϮ�Z\⽜���Dkk���Gex0�P�&�R(�-���wcð2�."�9�뱈_�h�7]WT��&�ʕd�ؼ5�,>��6qv��a��Z��7ӏ2���t_��g5��C�UI��YP�(	�*�I.�ԏ�y��U�h���s�`���Ӵ��/l����.<rY��^�8��I5�ze����.p���
*��L%b~?����j��(ju 6]�Ww��V7Q�L`��'��v��8�2�9:^����>����l���6��!�<=�K���"�u�r�$�q6?���>B�� �)�jן�p�b�w)��_8��?���NYX'=�����߳:���b�e�?DȫnƊн���LGg��X�"��&��~z��`��Ꝃd�������W,Ye5�S����2�35&���3M[[�ȷ�Ն!�r��L	J��6�ѡ���|�[Rz&�'��ARԦ �h>m��.�9w���9`�7#�=���4$�'�fƚ�^�-���c3�௏#�^T��y%�Q.GvJ����6PŲ)NT�h�R�.�j%_�����	�{ZN|�p"�#�`9�6b��b�r����r1>!p����Q�b7�,�g[�6�W?t��̢�lN����g��t �,��*N�2B��Ąz��w��{S��A*`=#�8��:"���l���+Ϙ���=�X��J�p�F��I*m?��	�s!L��٤�(G&*��YV�9u>�`� d��mS�`\pt�Oc+��z� �8_���LZX�У8aADp�j��`ih�#�HN'��q���q�|�$S�J|\o����1M�M����ڕ������4nZj'�����RE������O���-���֛9\�H�G�ƌ��^�S �x{�����J6��o�� � T�[s�)�X	L�=%�z�����E��ʠm�t�W�܄&ۙC�*����^������3ouΝ*�zu ��	����6y��Y� k�?�ǪRΖʰ}Զu�,6�������R���E�M���w�SϨ�e<ץ��}Y��`��y�1R�Mِ����㻋v��0�c��UCM�˟�An-_�t^���P�I۹aյ�+d7Ɂb��Dzm���ٯv�i��a��6��p���r68%�G��h���?N@�����%���]"U�w��F����:9�/��^�FΑx,l����<d��:���R��C��d9�O;c]������p�KH3�JVgT�[���x�=�y&�{<��F�'�H���6O��B�\/C��i�6�L�i��腡���y}UX�*���l���_0�!;Y�H�G�BH�1( ��h"~)��)b5q��؀v#���=E��S'X�o���r�'z���J�4�Fj�I|�5�A���]���՘}�,_�o�@D	�7"f]�!bƜ7 ,��T`���q�T�hI�~X�,<�;oKn[��0�g��`%����g���wd�İ��C�y5�3���r��R�I�?Q~
��h��:M�F�����|����i���w!�`d0 |ծ��F:�=HV{�X�ב�v��/.��}<��q���&�#����0�g]-���b�,���|?��8��|["��R���6���P�%��]���*;�Q���!�����1S��;�)n�~&<ļ�l�,X��h	��b?���N�t�2�r�5�L��zz�ܞ��q�r{��i�߀C��m�5�(���<�L�^�2�����$+��D����V�$R��h ���gn4�ۡ�),����LʝJܸ�b
.2����s��1�KT��XgX�ΌZ�Y�P���n��
��6�jz�$��P��l�_q*�.d��l�YHĕ�F�y�K�$�9$~�\"��}:s|f8NoN�K�4+���vXe��0��2H���)ϐsU��M��=ht�v��|$7!=���D��~�V"���QO>�mV+������'�~PT���G6L�#�lrg��0ﺒzr$
um,��$�Y��jh���
��~��@V����ْ}����z=t''�Ƕ�)��E��;�_���C���,*J&W���W�NJ���)�F���'��`,�1��@]V辞�|V�P@��*;x��v�|?4���EL��;γs&���x��ܛӪ���%~#����ӛ=p"��\�ᅸ^|�Ĺm��	V���/p�:��.25�1�QcW`�`gZ�?\��ʏ�$�����Cك���I�a�e�+=��@<n�p�ϰzr�����y���YՐ�꺒���E>���#�S�f�nާ\Q�+�+S%;����04f
囤�1����"~�������m*x\�bZSJ<rc����fw��@9�;�X�r�M�f��h�QyjD9�j�������_F����w"p�-��ˆohW>�q)|Y�Ԓ�FV�T��y�ڥ�d04�"2���J�,��j*��[�}ƪI9{hl@�*(B�/��;2b�ל���@x>�	���x7���ЎG��_��CTT�@����.�}�a =A}) ` E
�}p"���d��Wso3��(��@�yv��\q��ƥ>i��
x1�?�����݌2PI���Zf��T1��@,���|�Vǽ�9��U��<��/��������x<5�/��g#TZ���f�𻒁��-�Y]�A�+XPکBν�!f�(c�Ǜ�&����ƅ ���M\}�C��7&R-�C�q��B*�>�Ӳ%�����2���]l���Quʓ5�}���2*(��U��,�>c� ���s�Ϸ�$�x���%'4�fB����L�;�&!����.��}G�xڰ�}2��V��
�Xx�/#����;��U����.j D�~]��d�خ�DKq����Vvvs6&�{�v���2���k8� 0l� j�襂�_��&÷����ڴ��Xʠ	#�x�ݽz�E�-B1ɤ�I��eV9������n*#�SM���NvS���m�䯂�ff�ؙ����xD��mBJ��Z7^8��н�W�Lkf���8 x��P��R�� ���eB��$t.j��g
����R�-W�Y�&��
d?���9>�>q�׍ڱu&����2��t��Jg��yC�h��	��P�]�($r>*cb�ݯ�'y�����	�ܞΌ�`\����&�/�#����5<��t���?�a�I��e����I\��!�3
�L`�[?Q��=j ��(��r Q;+QG�rQ��`w�d��0�v=�e8����T[��֮�#Nl*�J�1�"!WRT=X���&�rʙW�w�q$.�)�Z8�9�:B?	{ ��e؅�[��JO�=�)>�8X����N��$��=�����.Ay��o���Dc#�ƅ;��%��}c�&���F��OS��6�jC����JfY���1_�������e�:pxA�k��3e&3F�Q_�[vR��^�Æ�X!�&$��՞����g��(|��z�ԅ�u�z��L�b������Z��_4�������=���o���1��f(����c���M3Eӏ�
3^/fy���/��'evEу����m�*T�_R1a�j �&�Ǭ|��N�{UF�������`T4�b�j���?���/�*B>3?�H�_����Q�g֫�6j/�tJ�,�=+ N�>��<�/��,�'{*��iB�Cބ�a wM�S�,�
��`��08��:����z��Ř+�L8�m���ep�U��d?@��LcL�V���b&%�0Y�P"u��c�ѹi�}.�o\�s�O���+�TrzQ��8�jM���ūҎaAK`p4�N�[~�H	/d��n_���U�$��~|�+���V01�3M����M������4�4�z�'�ؕ�HR�r/Dr��j��ML���9��HE�GƇ��^%�� ��9��H�š?�J��;��T`Y��$1]	�^�%�V۴4+��a�{���z�w�۔��*��B�u�#����4*u��E��� ^����%�6�6���sk�h��%�Ė��=���x,��̮�
��i����9�-W�xMĢ.V����@�z�x��Vk���e�LP����M���Z<��~�Yv���d	Ц��Ch�x���n��UJK�D{%����p��dR��b86z��2��=�H�dF?ڼ��>:p�v�r���%�z9���_Ч�CN;�H�I��@�= 
w�*AFs�K�u�G�ʵw^�����b��<R�: N4R�g�����/5cXPҲ+dp;��HN��J�����>�Ш�^�&��<�����cTOu��� �\C釴Sk�6��&i�˅\<:��fВ�*wFWl��_���;T������H�; ��"��s���q��������*��}�X�������'��`*�4"����0G(A6]^���,�zLJ)DD�T7���X��b!= �lj�oc��(}��/+�IB�9XREU�6��n�[�0>~ڣ�N��|O���G���Ad}H���}H��5h�:�5�z�U�$�CzX2�pR�c��:��q�H3�A��`s�b�!�r�0��p��4F�!���3{���'��n����<����O��~L[z����� �o�ɲ[6��g{�g��w~a7Vvв�ʨ�8^����]�WS�en��CH�m�|gb�)S�b����~�ʪ��]@�c��ɽS�2�t׍8r_�ӊ�ٌ��á��L������~u�$��^�ɂ��5�P�?K�D(�^z�&�j�<��O+���D�V�������wDn/�@��4���L4�!JWX�b�-�K_���s�Ϣ�l�သh�X֌Z8D�+Ԟ��|p��e6���a��U��^�_�_�.?f�l�ـ�0k�F}yS&����$���"WW�:��G|�ôo�@"K�za��uX ��0Ыg2����}��W�>���z���`)�h/��0b7�S���nD�xҜ��[��RQ���m�P�=T�^�e�QT���G�T#��r�H40�G��b
�<��`�Y�h���e�~g_2@��� �T�Cޜݙ�<_t�0���� )	uEK9��zk��n���,e��p�R�hJy�g<|��a]��W�4�;i�1˳�@�5 ����Vv��gZ�Ep|���W'���L��:ήpP�������\���}� u�ܐ���Ӗ��"8����t|�6iE��;lm���	���yP��5#.�˾���cr$�� ��E&��x$dnŦ������^��b.�|�߂�Ab����H��Kqݫ⽂�����w�9����?E�E�s�^���q
n�<��1d��d;�x����!f��<�+W`�D��~�
ұUg��(u�\	#`Z�/�r>��Ɩ8��x �6�&��;�!a�h��j�i���P�4 ]Ȓ/�F��5���)��}��C�o���>�\$|Y�9�-�V���ҵ��Pg4�i62�H�Ji�p�L��-/[�	��DrhӄD@�xBGAx�sU����+$?9U��V�x��V�(	GcQ|���T����.��xa[�a}䌌;2
6%�"�%�dڄPW)63�m�5%@��U�B�c�͡��i���x��Y��k �8DhPw��u`K���u��,���R��@�9�a�UN����u\��D�<p�c/_�bq�Zj��O��b��niW�4�A��DPu�θ��fw:�(5�����:>�`���\���ݐ_��&-������j���I���g��QG�ի(2Y/#��������}�4.���(&6O����>��� @�Bs'%j�2�S�H�`��4!xڶ(��1�:xz�A���<	�dk쳯G���Q�_
Ph;��2��4���}0Ur=��� ��~X����i,�K��ħ27TvN&����N2l\�-�c��l�ݻ(1l�H;je.���*�a����X��%f�N��ľ�x��zf�@-R-�߸�؟݊V4=p�c=����s#�Q�:�NQD��z*�J�fa���u ��E2nDÃBŧ�Z����[���ka�c�UJ�x�@�P��R>@�
�퇵�h�K.G��Cb��g$�mk�WJ�J&\��dz�k�>���q,���,��Й-�]2u�It��gk�C��ǒd#�P�;.(?0*ޚ�݊��y*�9�Q��)J'`;��ꦦ/b�r�n��<��ɔ��>�*�I�0eq�9�d�T�_w
ଝL���?�@��Ij{i(�G l���jC�MȅQ!�5`������v���8a���o���Mo։>^��l�H��,�!��L=U��A +���R��$iFu�4��B�� |��ؠ��uE���)G�*8�4h��~�N�B�D���Pߩ�d��d��ۥ�D���ƀ�p���^��)�&E��#q�����>�G�F��)��n��}�p�ݛɲM�ve�5$u���Ɏ�T�&�M���9[�D��꽆�N`�a��?ۨ���=�W���na�|�zF�PcS�y9Ǟ�=��|�������J�"L݊-| =�
�٪�}��df�	�Dy�nr3.�^�/^
]���K�A�v@ݩ6�U�(�
T'OR���jۂ�����?��{P^��&1���Q`o��b��M�����1�>Q֣2���2�Ӗ�gQ��6E't����؅kN��U�����,X�*D�Bn�g��_�w�fSgc�eR�`�J�8��L:�e����.O���31��:��pJ�/��?�	��EUL#���1@�& ��Y?�u�C*
�W���	&N\撌O���+�.jz��8�4�!)"���ņ!�a|upp�-d�V�s��W H����4��	M��O�$���|�����Z1��M�&�� �ڋ�G��w4��'R Y�MtR���W�腱����Ý�V
9�ILH���Ƃԕ^��� F:\���@-��%���vN�T�v5�^	O�%`RT�+�ò;8��V�C�o0�vۏ[y*R։�0LN��+R�Vu�03, ������6/}��Ϊk���Ǡ�����,D,l#K��<)��%�A_،HPɊ�}�	�W��I��ۑϳs����j�Ƙg0֚�M���ɡ��v�SJ�+��aT.C��͟=�n�殬�n���?,�߂�+��dm�wb���zĜ��ᐯ���_���9���p�V�r,�d%�������BN@N6���b���b�X�-wxY�FN����f��e�q^��.�|J<�:{��R�]�+�x��{gcSN���p��Hi79JL������y]��sm&�o��k������4��O����\~����6��iM����{�G�K�j*R�lQ��_fy;OɊ����HH'r �i�"tT����wq��l�������ʖ:�cXG{V���'p�O�;*+4T�!�+�At��]=�����"��%�[DP7O�%Sj�b|�� �����a���
�aI}ňX�}��1��n'0��u�]�� $ξH�2�d������+5#���P�������Sv��@��^��:�|�k��'%*��u�=:�!�J06O����F�m���{�ׇ֥�W�I8�(�<������m����5bk������ܲ����C�8���r�\����m�����3�C)]x�&������P�{��4��t{�S���u�~�!��	�b���^���.�N6�t��r�ҝ�͇��8-]�9�כ����(��ߒ"�yH��c5�x'�>���#�^uKW��{�>8W+�H���sVwʔ�F���xn*.�_��p��LO"J�\b�k�����B��s�ԏ��so�Y��X.�Z�N..ͩ�j�@W�6��Eμ�=��k
q�_g�Z.k�l�y����F�3y� k��Y�$��v"���:�Kl|�nooSS2K��s�n�X�^�0�%2�Q�Xg^��u"��0Vu񥦻y�h�\���7����uD�9����;��/Qm��\� ����
��T:c�Gl��#d�r�70e~����
k旽��iYHv�hH�� ��~�0�@��7�;�ϡu�w�utUZS��P8)dqE��ԕ�y���@��_�,�����M�J�������|Ǳ��bd���1�u@�5����V�_���`�H玔X�2/P�"��L&?Ω����"H�s��ͪ*���6���U{ӑ/�"�*h��(��Q��B�bm��	̮���0_b.���'vc�%�V���Mp�@�$������9����,ׄ�ǡ�!fd���+܃��懠�ݧ��Y���2ぐ.������E�T2�t���n�����ȡ�;�OZ�&k�f���f�2�߂�~��J���p��߄\$�ZI5Lr8��-�п�1���(洐�V�h��j:�o
X�o{P�-�DF��l�-�C���2��go�~Z>�g�|���V����/��=\"4��R2y/:JDx���,�`ƽ[��m��o	h��@ �B�ru�����Mu
��'>4̌�\�`x����Cb�G���n�cTʋ_��^�.��pa�b}�9�Vv)
���"w�YdW��3�z����R@H�8�K�Rv��|ISi3��xg+��C���P�9�Ðz7���P��,�h�����9EdGU	+��r��?���Y<�>/�P]�JZ�Ӌ
����R���\m��A!��P�;γ�7fҒn(٘������|1�;FNO�\��7�ؔ��8�-{wI��o]�8���pqI;S���z�2�����?\���ʉ�j}���с(����@J>�� ���sB�#ϭ��.��ܛ��4�������z5����\d���o�?ў���߳K�L�
��ȥ8{���13+UM�f�2 z�X~S�h�z�$�SK����7�v)6���z��	�(d��!��vY�l�Fj�_����(Ĝ�����ж�⩙ՠzx$�z�R�-�������:&�V/�V�d�V�`#pQ��vN,U.�O�����f\�ę�0� (DތB@�HZ��RΏ�gk\�@��{6xa��P5��R����q7�(���.ć�����O���JgWžG&7�$d�RB��>�!q������	���2Pj�t`�gkC��գPK9�(Z��*Y��eg�y>w���g����'�`�×�Ge/�J�I��<#D��/"6�tIF��e,�5�R��N�
�j�L�m�?�1����j�?�(=�Y ��!�k�(1�Q\yR`������v�F�8Ѥ����ъ�d���l`���'W�!E%=�	��\LKʏ�>�-OI$����]�/�B�Q� 7<�ػl��_i��fj)�h�8��`��^�Nj��n���$����y^�V�D�r��{q��۩Gx4�A ���g�����yP��h�۟o�H�8������Ⱦ�eƠ���?w{ ��&�&��v[���T1Ć�d/Ĝ���Ӕ����Ѳ^��)X@|.f0z��ƒ+$��WU��9	���S2�J�a�BC%�=��X�=�v���m��g3�f�K��o%o�)�3ImR��9�^�sc�*�[�"{	v;���������T#��R'&'j�DF�=����wn{K�4ʁh��T$�`�bb������#���`A�>���<���H��9g̜p6 ?it���s �N���x���J�, �]*�W�BI�a�+~w�L�S ���
;`n&8�5":����nV�iGm�a=�.�쮕��p�e�<�?�c^�L^�l���A&!�YgM4uo�%�=_����\!�O4c+�(�zMh8���<%�xxG�a�a��tpj���QX��4�XH��O��dԌ�i$K#|-���V!1^2!MA�>�1����{�.4|'����\RV���]9�n��w��\ƹ9��H{_�}�:^ۣ� ��4��.� �����WT�����Z	]_�%nQ�F:d��.u�1_U%�z���ۊi*�q��������$u_��k� ������6��/�� �k�;����[�-�g�k,�!�����cl���[�c���nܡ����2��v{��n#�i�%�+��o䚏�Mj�B��v���Y�v�;A��'�C�˟��$n���%'	�eh�:��r���Bd��b.e}z�dd�H�j�G6��Z"�rv;�g�3p�V�r���%}@��>s!���4N1[�������Is�Yw�F)�a��?!� ��^�"p���I��zq<�ޅ:�`�Rb�q�f�&� ��cN�����p��JH���JǴ��V���L���j&}R�ƢπX�=�O��Ok(��>�\�����6zKSi�Ñ��[�����g�*-��l��_&�;J	�X;�HR� �"�iպ`aq2���G
����'��2bX1"�4Z='����J�4�8���1&��A�@�]�}��&AC�5 �D�*�7�yN�b�}� ]�a������k����I��kX����,STnl0���!�+�r�Ιi�mH�d��u��Q���$5�x��k�b�}�?��y��ۭ��Y�Q:^ h�����B)��V�Ʌ��!F��0������FKڦn��{�J����$5��R�<T��_{�4[���>��� �e�����K�-@��&�m$�}�(ľ��Ѫ��]S'J��4�"�1����2"�/DS����(~�DѼ@����.�Y���s(��	Z�t�5rU�s��U(�s���ԍ��k!��3��A:��μ��L�5���yG��z?�^p��� �y��q#+�f�: 5VR0��6��n%�����+p�Lj~bJM�;b�:���9��z�s����"8���-XID%Z.yG���w�۳U6�ڕ����ˀw%�<_�*�.���l4:��fڏF��y	;t�U��$ϲ/"M��:��|:~o�K�fb��J�X�O�0��2�ȸ�3⦁�Kz�DΨpBL��h��e�9��7����D:6�'�3�)Q`�m���;ٍ�T����bTuO.GG�#Kmrx��0 ��m�
��?��8Y�m�h�&����~"@�\�VK�J��RtH!t�����)��E�hc԰���dk��18,��(V��H>qJ/~�����Q<�M0@��B1A�z@.U����LV,�q��{:��	�{�W��]�*L���Τ�t&k��ì-\'�|��¶�hI��PKmӌ�"���K���l�ﺽxem\��	���u�+ӽ.C���b�~c�[$����vj�{�B$��ܦ�D�ٔ�0�LD��諂�����WBܾ�ρ���ر*���e��W��I���5D�E�����p��7�%n��ab���\��;�F���E�f�����z�s~�*_��͞jA\?�SZ�ZVr�\�<WW��G�,b�҃�Ȑ�lhh.Y�j�*5J���������{F{�ވ���^���4oy:�>n�j|ϋF�c_RV��������a4ԏw2�5�JN��½��~d[���Z�@hI��@uVB=Ğ��TL��ΠaKu/c���"�xh%M�^��GYj�I��T3��T�.�C�a�B}Z�qڷ
,�<"R�dP��WD��3�Ƃ9��@! �^ͨ��W��inY�x�V��;���4Pz0ë�Am�+�,C�v�Mт��V9�� U�}�?��k�.���B<�/�W�Xm�Z !���p�c��dpo��2A\fzP�:�ή;�f-�(��� ��0�`�Ja�8\N���Ӹ7�O-6�B��Ux�����I��/!�(��i�2�����i�e���E}��R��(\�J�z�0>t�� ��Xs]}E�(L�	�Z���?4W�r��L��Y����w���1b����)���N��G5v
�!�`s�91���U('��O/� "O~N��s��ߗAKI�(Xtvf�,��hq��#J��|���1�_l4�9j[��m����Iⷷ� ��g	�j�:Vx3w�z\	 -�=��U��ՎV*Y���C�#/�0��N�t���䀝�fW��+-�����D��IB� 
Zȑ���v�(QxkW�y�͑xUPP�2RM��A�c,x���b.�D�x�KW���I�W@��&��d𿍼��>���q�h�M2vƄ!#��2+G�tK��g��C�a6���PWf(u�k*�kW�@�yy�N�oR�K��$+`�l	� /X��$��<^�Д�w%�NI���e������Y�\#
�H�Ll?"���Y�j1��(��C ���������Q�#`H�k��pvN��8�S��~�xv��?N&��yl�U��"��!h��=�ޒ�w���
s��.�$ߚ���$�*�BP&$ �2��s��k�H���0)�-F8)���^�Nŕ�)�*�2H_ߟq?�b��Q&�D4Jq�v<�6�p3~��\M����*������+e�;����5�w�7�������C�De�+���Q)o����&D.�肢6[��߷ϗֆ����ח�u옞�&0�

��nB|ITuz���ԒQ/�ԌJ�򥤅���ÈX�z�#UP=|0� u'�"�f����&E��c3d1���k^����e�_��ԏv6��'\ŞH�T>e�R��j�&�x�,�u<�{F�T�ܿ׈gY`���b�N_��^����p�><��Y�N��	��gG��6�vt�����N������a�`��,;�*:˗B$�˄f��wRcS
�Ģ�@`)��8���:�[k�I䫉������)V��Sp�A@㵂?���>�IL�*�g�&p:Y�{]u*@l�Xv��{\\1oO�e*+�Bnzb�8KWA���<2a�)mpq��L=o��@�H:�2�j�g߾X戣U$?��|�!F���1���M�;�Lęځ�[�a�4Z�?'��#R��
u���K3��n�7V�9H@�HR(�x@�^6�~ �{͓'�Q�6����3���ZRT1��T	���%֩Ҵa��1E4�E�`�Y�H�`ۅ�t*m�覹��(H����cu:!��k� /����L6�i�ERek��ǖDp�6�]Ԣ��,�@P�� ��������~���2�����m�6���iJ	g���X����z�
NNME��D��O�Tv�Cx�����C�]p��7sn�@��`�0E��5�m��#�ա��d�ݍb�=�zzLu������~�U�E����"��pw�r"i%X�^�ya0�x�!N,t��ZS�qjK���wn=F�Ą&9�ܛ��^�Vޑ�9~���<<�Դ:q�R=�6������rtcI���<�pl2:H�ٺJB���r�[��[Ш���&x�f�!�}�ܬ�jgO�w�w}�\���$0$6u�#i�t���SAP*��l��X_��G;Ei=����H��L ,�"j��Օ�zqm�Ѐ�A���)A��X�2�O�G'f�;��4�s��F�!ɅA*�]�މ�A�����ۉ7D�p�7���I�ob2^N У��,X��p׭���I�G�X#O1�'��n��0o���<�}��#0�t����dN�'�Ԩ�Y��5�z�Ć�B��R'ڵL+.Gv��T�8:��3�yd-�]M�Ѥ��G�!�i0l����F�f)��{1�w�}�i��v��[<����%����6�Ӆ�������h�p�n�Y�h��H�a�����7�4�].����l�������/����gS.s6���~��`�{%��.��T�Y��`d�ĝ�t(_�r��U��CN̮_��o^q��O���H�U���t�Y��5q��Ѵ���{s^k�l�{8��˳+3K���BV-t��q�Z�H��n ��O���TOL��J���bv)���`�x�5s�>��}���WxXd��Z����AZ�Z���v0�6���r����{�@�k_]��.���loc�� F���ydu��Ec$��"ȘX:q�|R%�o���K�-�$��XQ`�0!�Y2��}_�BF�ߋ�k��qz�h`th�T	L7W�{A4DuF��D�H>Q�k�mBa�V�f��m�t�sT�[]G���#R�rӛ0����V�
a�3�iԄY��hP%���z�~x3d@BNd�q��0�-R��C}t�`��j�)�E|0���Hy��,�~#�,?f�*�C�_J�w9m���n��ȕ�ߠ1|��@ɔ��ٴV�d�,�P���9��j�螬��'�L\tIΟ���(��[x�H�h���
�g���`WӇ�:"I�s��x��JѺ8Gtm77�	BAJr��&g5.���+cñ`�Ln���̶`6$5�<���P��:� u��)��M��K)��l��/����_	��쾐d�֒��+E�r��d��U�nʻ[���9;�]0�@3fvL��܆���~���fE��Y"\Z�IZ?�r�۴w紧U�&�'���ޚ�R�9hIF�j0�*%*W��3�c׊Fvoo�㷗�`5l�o�>Iݵ|
2���̛V����3G���$4�R�2o\�J�C���n@�W#[�m���&h��@6#�B�5����O���E����* ��=x#�n�ytG�&�$
�T@�ά��.��ual�}�j�^�
��"-��d��hW�Q3��j����@��+
�H�S�2m�i�6�x�9��S�I*�P5�����
��k,~w�������9���U*�0�P����g�{<!o/0�$S�Z{���	��'���ߣ]��(�A�d�PF Ω�>f��O(O����J��Y����A)\�Ӌ�����T-�߼�[��.��ҪB��C���Z��x�2j���I�;�,V���l}`����)(��L�u�s>ϼ( q�sxY�ϣ����(����4�ls��Z�0��k�Q��}g�~����6�d������B��
aVE��y�9��'�$U̙�o� �i�~IK4�ؚ}sK�9�����vߵn�g�$�P��\J���lO�j�VO�H�t���R�H��8U�_Z��Q�xN�z��q-��ɐ|��p�V%�w�t/����'#J����N��j��^O��ufR`���s��v�D��B6�Z��C���.�ï�kR��f>�x׶�Pk�R��a�<���ǰ9��.	�}�Ӹk�\��h�W���&�#d+M�<L�>�tq=zٍ������2Dzt�p<g<��C��u�kP��h(���*O����y��_�
]8��͞:B�`H5��;�/�����4�<����e��E$I��e�K��������
qF7LL��?�Ҧ�Mxj�g(��� �S<w@��b$Q��`�$���l7v�c_8��ū�K�:���R�0l�}�K�!÷v=D�D̒D�ʅ����,�$u�F!d�%m�B�� �����������)��8�z��~�N �\�m�M���/�=��aD�A��q' �����w������^�&��&r�������n�خ���.����e|�%&�������w�&���=N{[���J��h�}���%���r��h�ퟥ�|db�z�Z������m8�o0��ax� �i���&�s�5��qj=W���[�:�0sf��b�%H�����3r���^����W�XN�v1�ѩGt��Y �TY4NRk�jl(�����!V{Af�77#���`�\�b��,:����$D����>�ִ��	��$&�g�O6��t6UY̩U�N���.�.��,V��*�^B������w�w�S��v��`��+8�:v: �$�܉��e��>
$�ۮK��p{о���m?
&"�KLԞS��&ߵY�Fu�0[V�UͶ���\���Oj�I+�|zz��8�r}�n�X��Ha-�Yp�Bu�GB�����H�-����ZZɰ�c��$zU|c^]��ւ1��M����g����N��<�,4�;7'#����aR�~0����H��m�	9�� H�d#�s�^�Έ wL�B�zﱏξ����'�T̏�5I	�D%�ش|����{���J)�S����+ۀ�*c��a���C��uz�uғ�7 �<����B6@�� ��kM����<^��i�,=�֮��0���r������d�/���g䨐�׬���d�k������M����<M ʧ�F1���b�v�ky�A�В,�C�ǽ�y�mnt������Df�0���(v��\^Td�2�b$6�zUTּ���}�@�P~U�(Q��!�p5��r�I�%3�K��o��oN'�]��W�,����w��F�J��aRK�6��^̪h�?S�Nث<��:��R˫��ٞ�VOcD*���Pp'��H���J��\�M�͙*�x�D�n&s�׾|���0 �S�Oa�<Rܾ\/$����6p�pi^LX�H�X m]���*�fl�_7�M;@� �Hy� GP+"��p��q�Q�}�Y��t�KgXx���j�'�Dd����4Ϙ�P	��A���]J_��\Q��(����D0��7 �	D�9b�^T ��i�ۯ��WO��BI.��X���"��n"I�0* �WG��hU��O�� sd�����"W5T�2ġ/k�s�Zڐ�f�Kk��O�{:��4I�x���Llх���!��J0|����FX��{L-���Ħ��?�ȟ�<�򒾋�j���fJR��[I�s�!��H��	fS�cJ����О?è�e��ܐ]	w��Q{�X�{��d��\*॥�SIc�����~m�_����3���O�-�)����tC:SrK.D�^Q��(�
O�S#�9�r��U��:P��?�5LC���ύ��,^fXQ�־��oE+N��0��V����{��s&n�n�p(��Y�L��CJC@bQ8}�7�0s��?�� ����X2�Z$.������ϸͦ6�
��Ї�A��[gC_�u�.�9{l�lĜ�)F��y��F���$M�"C��:L�|�0�o$KsK��Ӛ53X�#0<�2|?K��7��CX��zi6fD���*ph0��o<�7���V��D�=�]MlˤoQG9m�LY�q�g�JO�O�4T�@G=�&#y�r.��0���`.
�t�D��Y��h�Cp��l~�d�@��P��;@������ot&����'g)u&!E7=��'��Z���Y5�,Q�(^�>.�J��(�>���I�C+����V1�T!@d�0��,�V�9�Ջ��^��=&����ӊ�L�>�Κ�J�yy䐬c|��r�k�l���)���9ӂ�c"�������պ��5�m�J	}�����!�.��&�أ{c�'ſ�Fa��(o����$��Ԧ�"��J}��Ij�芘���3��_��4�eϷ����%C�j茸c���'b�+� E�1�J���m7!n���CF��Q�;�g��ZQfQ�a�,"���~��\��$���&\u��Z�or�����F���"���9����NhdShj�k� �N� M#���qFq�:�>�Ѡ�@�Pd�ooJ>$Hq|E�#ԙZ�V�Y�@�"�n?l4
6�2ꢉJ�Y��8@}1P�[~y;���h��@Q�=B3�u������q���%�moLx�T�-�GO��u�T{�Ĭ�j�.�g�a�c�}��'�
"7"�QdƍWzOJ3�a����@y0�F���m��/ki�3�x8��������a�P�A�ሣ7����i,�.���8���9V+3U:���K�k�a�r�B�<\/�,SN�Z��;B_�B��Z�7���A҂�P��uΤM�f�[�(
��6��&����H�j�\�$Z��`��-�!���&��l�҅[��wM$������2Ũ��m��Gg9����};���.<(���p�>*�� ,g�s�U��+㞿�-�L;j4����{��j&w���d�����о��Dl߄�ɻ=5�
����H/�T�R��$Uސ{���� K�c~D�gyȖ�U��K�����v�%I������"�v��2B?ݧ�lj)�jQ��#���M���舓�)��j'��m�xi}�zR��-���������V m���j:��p#e�&��N�G� ��䶤{fM�i���{�19�D/h�B�qZ~�Μ��^.�kM ����x�s�P�?UR
�v<f'��P��tZ.�2�.uĈ����٧:W6Ɔ&ȕDdf�`�נ�>�g�q�aj�÷���I�
2�`�t�(�g�I�C᧕�Ь/P|�(���*ʼ4��^�y�`Ĉ��5�'p���`�V�/N�E�ڧ�<�N�� ��͎�IWq�e]�B�г���
Ld5L��[?Xӣ}aj癦(n� �)���+dQ��`~����K:v"�8M����Rn���OJ��l1�e���!��=���̭�� �D�K$Uo8�b� �~B/@ h�����ao���d�)3�8_'ڶ߾�N{���/Ӄh,ߕ�ʮx��&DjY��l2��숃��뤒J����9���*B��q����-7�i5��I<�9q�eW�a��H���&�����D[�a�����Cf��M�3�}��ޒ�����Z�2|�wzL�&�����
����u�[��s�M���8���=2z�ٖ�!�8_Cf��8�����Ze<3����oX^vxK��2D���v,����b��Tt#^R�=�jGJn��>���%�{<�iʒΎ��L�`�6vb���c�Ԍ��10">���|h�ĩ�?��g=vp6�Fdtq�v�D0�N��I���[�ִ�,qX�*0SBڱ�ܘ_wT�'S �����`��80��:�8���_���@�2�5�}���gp6���n�?�o��h�L3U���5&nmYx8�u�j�vǠ�aCu��\�O�OS�+���z�"8���ٮ���Oah^:p;4k�Bg[�E�H�}ѻ�<����>w$�
�|�����1o��Mr�܂��w� ��s4��b'�~��y~Rg�2�.��e���ϙ��ը9���HL���n,S^�� 2=ϓ]��,� ��	��b�Tg-[��:	nP`%L�a���v�'����p��4��~��{�*�����a�^����gu�$ e�T��ht6��;��U0k"ǌ�	��.�a�30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�*ڜ47{^�6H�?�q����|�emHW'wNn�㣔��Ld]�m�fh?���D�����xо[����9�nL�/l�Z~��p �G��)P�A�U{q7^���h�j����%$�59�����w���׏c� ����h���u�xW�kE�V�Q�bͬ�)b� d[%�G��'kf���Z�Z�;�H��^u�Ĕ��S�l�ҧ;��(�6�Z���?��l���gtǴ�'���t���s������=8��m��GB��2��6�YOf�F�V�%�����Zo)ξ�p
�ƃ�=SX�����[��\�KOq<d�'� �@/?+�h��	-�'[��G��[8���	l	o�5rv�v���h#Lz��-��`Y�~��)�gDg5uH{���Z^9��]����5�,�'�Bo�(�s��Kw�=Y�T���h�a���/�,�^o�Բ�Iӽ��u�&ka�a��Ҷ���\,�'&�m}㾃Q�aV���H��ÿ�Y/�>�w���Jߕ��x��`�j����k(h���۷*���E�;Z����Xb�X%	�0�v��Ko[��:�3�e�r6?{�j�X: nN�$�F_�r�io�~�0�*w`^�w:8\��B@�L�nl�!p�|J�O\��_]�Sf=� W��1a *)"�V��[9���&E��Pz���YO옟a�-��~<|3��ɲ�~;��<7��7���8w) ����dH����?��;V�$� R�����L�#�Q�jVV��H:DFm�(گ_�9*t�s�σ�=�4n=ڹ���P��ӭ�p�U���8aK�Ǩ}S$���逑����4�ɥ�Ad���RI���?�y/G�ÕX�F�c�v:�m�]�V�9^���-�4���i�N9o�7̣�N)�}�[VK��;�Q�h<�ч/k}�[� Q�?(�W�[(O�����ƴ�}ư��x&#��l���^B�a�'i�
W�p���}���B��yO��xNW]�:��?�
_�oC��l��ad)+p�8�}Wbg\��@��!�r��1���S��d�3	[����X�|��R�-���1J&<v�L�^����?P\4Cھ� N���
�9�#���S�㹘Wj�����W�]�{��ϧ��w&B~��q=������	�W�r�sxS�E��^x��>�
�o/-���H��Q=@Y��r������X]#yE~�����ȿ�����;P6���Z��̂Y�q��&^)��=��|&^`����`���׌k�����"sI�MtZq&��
�?8�0W�߀�~�!�s������;��?}��Mӎu>�؍8��B��]q����mp�ۣM��J)���/���'P=a�7D��EB�?���	�K��4��U�Ku'%?J,̀�y�����.����X�94�k���9dƪ���i�Z��w������DFh:��̭tR�;�۲�]��!�%�s��۠���~�m�B��������`z�{-"q���i�����_���}��.z����
��B�J�#��g�I�z�N�NE����6�qZ���Ba-姌6�T}.���+��J|�]��.{��> ��$� t�i3(�*���sA80�.�]�����ļ�WF�i*r��z;,�3��"C��UD�����.�.���'y��P�ې�峴C��v�h�C�ݯ�T�5���^b�8P�Dxu�:y➷fA���D����G6g�*�M�y�e|��s�I�xD�٪�>� ���W�[@B��[%Jx�������j�IE�b�T�5� ���F�Q�jk��ўu��^ ϡ������������"�?���`�m؇^<]�C�arp�����ǒ����Y����A&0�����������I&ƴ���f��@�J��4�'l:X^�<_)����J�ِW�0rV�"._���r&��k�w�E�$�)��b=�l�d��k�_�W�d��ʱ(���9~��'�5l@�Q���Η��f���N�'G�_9E)|~��;����!��5T���ɫ� �ؼd����� ����B��ݘ�we�� $�^��W�.w�& v�'E=�A��'z�I�[-���ò2�/��F�����ueH�zS�T��F��E\+��Z�պ��rr��7��F�D|�Xe��K��b�>-�� y(
fOE�5.'ܫ��/���R�Q��s꿥��{��|���.,|�@Z��_���O��)#O�{��� �[�ͯ�x�gU<o�������	���5;��yS����Íp�U_��M�'L�&7�/W=ܰEl�.` G�$�2K����b<%k�]�,�/�9�4=�ρ?������	���ʌ^0<?�g�)�T�����adA��D�N�	 ��N$�m�	��Z��t�Q���p�h��o�{|�Ϩg������Vx�_��"�h�:j5+�w����10/�K���s��Mb��$rᚍ,J2g�+^�)�<m���qЏ#Ӥ������,�C�Jz._��Z=\�ٮ�i�������[:T��������r�(65|q6�2����aI�s�6�
�"����_��xq����f6�C�)u�'1�K[|lL�d��p����B�fe/��X�;a�{�K��РX����\Pʫ%�:�f^�jXD��}Ҳa�}3^I�w������/�%��+��H��j�F�/���i��a��5
����-��cL�\�-x;���!�z��Q�F���S�e���#��ű�^v�t]}n��fy�ǈ 'ٺ�2�{����*np��VT�M��f�K��x�/?��������aP	��u�$8/V�rB��e��l.���X2���˾R�c^���I���N�4�G!�R<�p_"�K^�-8g���>�a���\�,�˞bFt����g�G�l���)M��fA���*�t��)7Mbvr�=+�ti/�b�A08L�;��)�p ��d�D� +	��&�/���,�(�ɔ�bG��-�<m=_�,Q����x6�~�(SБM�7ĺ�U�ٱ��?�co�3�t�Һ-�I���蓟�<7hP�{w��i��ؔ���3a�����`� ���9d�vS�!��n`�����O�j��$�|2�߃n���M;��6�G�ɠ;�1��Ͱ9{��5�<�i�P|��6T$�H��tgB��ԩ^1IA<�����o��x�8����]gR��5�y���W�|"��ՁT� �����]�u"az%/��.m]n7N1����.!OL?�m�5CDB�em3�73�<�{w��-��EL��Ұ��D���o����hB�IV��E��ZWknV��(�6�
byY��ஹ�����[ �$�:�m��ޗ��i�m®�9��pz��=$a;�ZŌq�!	�d���C���zR��D3 ���L�/Ɨ�8R�a*�Ϝ� ��&R�$��̬dc�6��1�|�IB%����3��@0�Ly)ؤ:;:H���zQ4m�>:��Q#�cg�.�y0S�B»K�0��%$�S�PTGsKo 뮵董7Q��`�3��S[^q�Ȇ��?�d�"-"�MnJ}	`��d����L��QQ1Ặ�ݛp�-�:��E��_zG�Ś���Į�n�BI)���x�kHf�UN5�d!vny:��Y�Y�(���v���5���¹h����o��l�n�)i���e�&%�Գ%�:2B���P��Ʋn� 7S�{�ş/���8zi�ɻ�+@�A�˘�̒���'����:ȰW��̪�Z�*}��W�"*}yQ����Z�N�gGQ�f�N1o"H1�R�b"�J�E4�I���Q�|`���R:	o��[t���� لI4FR
�i�|�<!	�Q^�G���O=7���Is�w1ņÚ�3�#���$d����
�?Y��@V"�0R���zZ�#� ����Zu�8t4�%q��l>��0 ��U)p¯C9!�׊v�k����矔��� Ϟ]���G���XQ#|��,�I����	;���䟲c'�xJ?ܖ� )��h��9�a�GrzlD��r��!,�v���U�`>��F���'� ;E�9��ԩJ˸�f���b
>��#0
�P�vEo j�I�9_��_LIT5k�1��Ӡe�Ḧ�nݘ�������*	���s��`��a�_e��*e��7f?=6� [?59��������W�u�'��jLO��m��?���D���O�Љ"���O��6KLy��񥲆޿-#�!����$�9��^l�`�S�Fj7��_^��@�G�x�c��ٸ�����h ��V��;8�@)kxb��E�����נW�T O�%2�O�ҙ�xZ$�c;�A�����O��������>���;(��Z|@�
�1l�t-��Q�n%d�'0�;�B�������h8�R����Bh����rY�<�FA��%ВTo��ށ�����mSC ���D[ɥ�\׻�ܭ6�`� ۸c?��Ph��;	x��[�W��E�X��lԨK5��v&z|h67��T��Y����W�ϣ2�5��8���GEL@�pߐ����'���S+Ps4j���=��E�_�DXa�'���}�����T�M��i��2�)���v�.��Lk�� L,.!)���s9:`��ânk�ݟ�v�A[��[�(����yd����q���Sw�HϾt����u���[��39�=�����b��D�ǀY*��_C`���bt�jo\%�nP��w�u�����*#�'��S<Y���*��������w��x|�h�����۔ QwV�D���A�)����[��|�{�V�?��Q��얣��#r�ܢO�+�X�,T�����Q������
Ҧ8�9W�P�F+�(K�-��}?��<��'x��F[�,8���]�ޅ���)dx�[s���K��ʮ`=�㜯��ߚ�`��6��=��/���T@C	���lJ����ߧ	�䦛D1�6�p+�ڹ��zN���6k��/;~e8g]{�F"o�M�ӹ1u�����
P
I5Ǔ���:�F�4�+r&�XAw�Qڠ���Ae�Y�&�����ڒ3���m�<j�+���+Ń �2XWΑ����۳$�mH2c2Y��?�	�>��Gu��ws*��Y�_��'�뫛��TLL�u�2$G�L-~��2j$��'!�H��ȹ�T�i���(����E�]����!ё�f�(>�`n�r�m���������1��Ȯ���M�.��F助����7��:)M��w��=P�lk�-�5*�Q7��8�b�|mCj%յ#��s���B��hW��0��xbe����t	�5��_��S5��#���#���O@�����J�P�5�a��NXf�-�S	�w�Ή����ʗ�[��?��{�ch dW�^]L[�5�(��)G�G�pMk��1tc��%���ڵa�t�|�=C{~� �p[���̾����a�j.���ѫ�Z=�.�]�D��?:E���ʰ6�/�i;���n{ؽ$[ OE�h7�O��Fi))稼"B�\��$�gFɄ��y�I���~$D�ߖ%=�O6����iBn�q��̍;,~`$�cs��;�������yB˪`P�[M՟�VS�m����غ&��[Xj��)ɇK�2��;%������j���waQQv�Q� �� ��02l�z��s�D�������U����/܄`�Z���p�bY��ؔ����J1��ZZ��o毐_G�ZY��Ş��{+z��Z��3��
44\k��Y�S�E�(B��[�@��i�J�3��⾅�[aD�Co-N���@���eժ5��+�1�{L��!�{վ���b�<�Ԓޚ+c�1ŞhQ���I����%��1�KE;�)�@Klb��l��bA9��3xMn%�7^�����{;���ن.�e�;N�j�����3���~3r�w.�ԔӜJ�NN��K3���`��+� �>I[[���= �V��sOg�W�u���yQx�����Ne:�4ՙ���>���qku�':=~�G@l�F��;O�����3��g�:v��� �\9'�}Gk�OPK,T]��c�6�=�|)5���v�\s������}�͡W��r��J)�·nt}��]R~z�r�.�b�kȶ
]�d[%�S��2���Y��eiO��4U�P� ;�=���E�yx�5������;K�j�؝K�Pa�hض��B��׹��3�%���8^/`j>���7�|D?	:��ĸ�\�=��Ikm��1	W�?H�g����IR������i6��V_�F5�ʑ�F��ґA<N�v!c�v�� k�^�lǚ��j*�!p0�z:O��x��4�k�%0��<-�Z��|�pEc�^��1@x��q���
Z
.i*e�i�ೆ��Ev
Bn6�\�(͋f�۠Wҹ�b7�n��9tƃ��
,��:M����l�$`�q��հn���ie�a�,�9����D�����.���=���t�?!>�|A�l@7Jl"��0��-�
�V�k5s0�> �w�ੑL��#����X/��%v���>��8I��x�'ʺ'lrc`�7��:m����rl��V��~�t��W,}++:���O��L��	�����W���S����� >Qٍ(?��a�
�"\����c�9/@�&rl�ϕ���%O�T�a<k?��/%3�O���1;�.*<gx��E�� \�B߾H��p���;�Ӣ�����oL�Y���V�o�H'��m�o��e)9��ˢ�� ��0D����|��=#<�`_6�q�p�� 4�Z�tZbSq}#��Qi���ՓD��k�A���_sYɊ^��'��5���͎��Nm{��V$�i������`w�[�;D�������JD�V�D�;�8<h�w��|I.�H��QA剣��(�*��[O���}s֜��@���k�oA�Bƕ��"q
ħk�'��}>4B��O��iN�-W��طvu
��OoP�@�K�c�]d���I�W��x\}�����g�c�1��W�_dظ|	�0�DtX�I�ܾ� M���1��Wv�HK��\�}��;����|����&�k@F��%k��Fc����]h ����XC�&XTv� =<��G�	{��r�S��)ʪ���\�¶Y��ːv@&Qrc��� B�ofL#�O��G�a�׿�����4���sPh�U�NZ��'�o#Mql��^V��=� &�X���ə|(/��k�]e�}�sv�:t'�&/) �8TU�WA�9���J!z4�s�:5�����Cr9�"��M��e�Z,!��.r�xd���qq+\�ڿ���MI��v8��m�~��'}���W�ڲ��?���J���q�4�ʾUn��'R��,�fy;J�f-cN�¥w�4w�<�`�����ͥ6���FL��C�r:F��ӹ��RZ���ߐܽ8���Ǉs�y�1b��4�~�W�>�^�(�f`G�.-�Q���Wq�syr����6%#�z"����F�BH�#��W���wz��n�;1�-��SB�G~���?T*����q��t�ƽꞩ�[��л�>\� ���i��*�'2�A��.ɲvU���1�WS��iו��ǭh;�D��LC���D��e��'ͩ��'�|RP�;x�r�C궵�5�d�J>�T�f��^�41P�A�uA���ˣ$A��.��M��`U�,�p��R����b�/�x�ܪYΞ��p�/�U[���t�%׌=�Ԟ�v�fI���aw��0�j9�㔩��)�*U'u�·^��W�`ZѬ��J���\}"cΞ��N�:>/^�|BC�n�p<p��0L�}�YeI��0����u�Ǽ��8�NU&�\��SSP��SJ�|��˅�p�I�˅�&tJ�W�W�x�V�h�_1�j�?�U��w��'$���ï�2l��_�3�f_�+pd� n��8���9+<��t[l-d��F/��H���<�X��'TG9�~<$�(��_��3!X��\�b�����iA/�
C� ���+|��xh�b�oe�3$��!�c�*.�� c�SEʓɲn3��u~zHQ#[:ו�5|�F���<*�o��Ǣ?�Hސ#z�#����݌�9c+B?@��M��b��:(��'�B�Xrt���(Lb�����9y�Uif=.ZEP�.�:����T�����s׌��+��{姯|w�.��x��@�
_Uֈ<Rl)���{�C	 �*��3�U��s������6��h�yю��;��Ú�MU�3�ܣ'9��&�1/�������2�G����lq�D�<��]<�d/�i!4
G�������	6o��ٲ�<,��ᶇ���.Ė?#���	�a2Nq�v��,Z8��~���=�#���{��P��'��C/���t�O�BhO�5�����������1��(������P�g��J�ʬ+k{N��_I�$�m�%뎈�ŗ�2Ok�=J�&����\�)X��2Ӥѯ���[��p>�߯�(C�3q�y24跤�e�IK}�6M[}�:�ZYi_��qb�d��u�C�R�´wcK���Lt���H_���@��/:TX�L���KAΒ�m�䝃�I\]L�%D��f�#�X1}_s�In�m�r���o��N��A�"�����RL���m�m�?J�CD�����<j�1�'�P��l�DL!��M��g���٥�<97��&N�)^�_��j�N�Q����G� #m�8�	���� Y~�[�I��C�x
�E��Đ����\U �$%�Z��z�q�2@#Z�la;:c�͚A���я�E7P�_�̧��A(F�~Z$�����lf�`�4���q�����>�[x��,��82�Ł�pTB'��(�rYBB�F�u%x����o�k7�CVPƶ{SS��һ
"[q�9\�r������ ��g?Mt�h0$	 %[:b���� ��l|��5E�v�mDh�����ҩ��I�Y�Ti��j��*�5H�d�Q��c��K�ʞ��}��?��';�(���sܭ���=L��큃��a0�5��Of�1j�Q��.���_���zY����v�#������
.ɼ�J|8:ڽ�JAOą�?vW/d[Iw�І��G5^�w�qT�c��qHw���ԤO�zjްh��c���=[b]��o�!*�,7�%�eR�b�vo�n�:'wA���R%�*�FU�3}�<J�ێ^���Vͥ8��wf�|80Vɣ]���Q����ڄ�b){��<���$������?���Q~�ʖK#���\s+��,��`ޚ����Q������}�8/Z}���0+-|����}綗<=h �gF�b8��]/<�v�,)��?��hsk�����V\@׋�l���B'�`�l��s8��I?�v��C��8��+����Ol��NS�1��p�(ٹ|i�z��i��+ԑ�R~�X]#��F�C���-�����=%n�Y��
�2��M�	���HFN1�+�X��/w��VŵA�v���{���傷֤E|#m5+i���>��+n�2 Zt�lnu�9b��[.m�H2�[?�j�>Q�]G������1�_t�}\F�C��T�Գua�6G�S<L�%���jؓ� !J��p��T�v�s�1�N�1ő׮����X!y �f����G�r���v���8�*�q���I��X�u��$���z�� ��߉��"uM����+Jպ�e�]'�>-�s	������5b-��C�;;�]*ΚӋ��\̦��ͯ��]0.Yb�5Ǽ�t��UF���C�ݝ���r\��Gc�g�@�/U��N�J[|��~�a��fN �-p����Bw�,���:��r�n[(�ڙY�c��d�q�)2���o(f�*G���p�[c�7�ca�����	!�t�3=�l~���p���t��c�(a)��ʐݫ��=;%��)S~j���D9��>j�X��/uS��v�7{�˪$i�EJ�/�&X2YUiѥƨd4�4���*�$��c�,f۶!R��jN~����>_7�3�N6��÷>�B�^�S�5e~�2co���x}��i��l��y���RƔP��%�ɩ���X��J�b��b/���x�j<��/s�2d���H,����j�g�w	�Gv�����6 �C2.闝MD�'����2K&�f�UR%����ta�ud�YRr�����'�11x:��O�|��W%�G7-Y9K0�g2+�":�N�3�4T4�#��{s��B����\V�k@Tȸ�/�3��K�=ҷ�P@xD����N/8�@2�Ne}�҅�1��n��.{}`F���
-r���}�Ba��ٯ�h�s�?~��5��Q0�K�^�������n�Nʭ9�:-x�_J�߄l��}�#�����h�e�S�NS�ɯ�6���B���&̳_%��|�ݜ�C�N_9y3L`.2w`LӨ��I1{��� <6��$+��{u0"��!���q�ͩK�:?�_����[;���us�x:��G�|8FW�O{�Q��+���g>�bg������\�_ }�O�M�Tj��Ѭ��Ƽ)��+�db�\&��F"�%>1�I�ζ��x�)�Tn����$z+6�;�y���������T;���s
k�����㖈��kUW���A��OJ���!Q]5F���hA��B>j~��K.�}��c�/�ͯ�M���z���8OQj榦϶�s|�����`һ�[{>��]9�+y]	���HF9��J��R�wĂ5�i�B�VŎ5X:���Z�{���j��%YcU�C�g�7k��lo2�v��=C�09��O��Gx���]kx�h���r���|�%EG��V�-x@�	�R�6
��i���m��.l�Ei
��p�MT��SS���7�a�D7����B<��s:,P
_M8�H[O�$�qb�%�WR�'`s�	��,ZzѢ"s�X����ǆ�݀�x����]o>�pS���J�������@���ұk݄��F;���Q"/�p�әn�Xמ�%�`�Hxꭠ����ς��9�r���߯�:�b�qŭ��r{�բ~4js��ֶ��:M��LG��떮t���ൄ���4���e��5E�W��au�"}?���Z9ׅ�&g���O�.a�y֦s�3D�&�0�q;�Qx<�ފ�L+���O V��Hin��t��;+���@9��y'LA����VK�]Hσ=m�Z�ڄ�w9��袈�փ���Iڮ׮���O�E��`#pa����W��2�	JS�~J�A���}V3�>��Ay-�E�2ܽ�n���X$�{��Km#�7V�

�9�Sɉ_�ƭۛ���~���4���V`�;n*Fh��ч$E{���Q�j�,?�(ā]���Ӵ���}%U�m%�>Jr��Bn�����l
lT���>�}�B��O=G2NM�W2���_V�
t�Xo�$dbꮻd���mGTW7�\%��,���'��1`�P�H)qd���	�V���N$�� $�gEzBO�1��`v��n������%1�HZ���Σ^ΡЎ���ΦO����w�q��b�]u��� �& �vl=��Ǚ,	#�5r���S�F�峏�3�]�p�Ed�s�@��,r�'�נzP��%#nlZ�m ~�	�J�`c��{,�P��P� j��=�Z�Z��$�q�^���=0!�&smP��xf�$a޺Hzkr���%)0stt�T�&�e��}�8�[sW�T�O��!"��sU��pb����7�ʈ�MVȏ�0��m�� �/�\�q��ڂL���9M��d<�&�H'%4����Zc�?�+r�<�}�@Ŭ4��Ub�'��,B�Iy�&O��ש���M�!4ԋ����|�������"s���	F]���a۷R)ۇ�"�ep��:�s�س����s �&5���6��Њd`�A�-7�|�A���E�t� �,~K͠�z�����B���#a��;3~q=�{�4|6�C'�d�l�|v���}(�)�G�1sp쌯]��c��'������t�y�=�ߌ~�91p�惕K#���a����i����=r:a����cAR�j�C.���m�/̄�ܭD{Ϯ$��.E!�c����iH+����k�2��4�$|E>�R��ظ��U�~Cهߕ^��j�"6�pî�8B���Ѐ�����~h�crն��W�����c"�y���	�PFyRl�g�U�֥L������Y����`j�r)�ƥ�2ۄX$}q����j�Xw �vu�_4� 2|2�:+���D�-�㱾�)���=}����z^�����f�Y�f���@���~1�Jj�j�77��?�G���Yp�B�~*�+��B�ي3Jt4s������R���m��@KM��S�3k=G��G'��h�DV"@NF�j@)A�eT�*�<TI1=����{���}P%�!��߷���S���h�˰������������K�q�Ȭ�ʢ��%s���4e9���xL̆�|6��[�M�|M��k#WeBe�N�3���	C������t�6�-�3y����tN�@3��8`e�wxk����IھΛ<� ӕ�ve�V�ug8*�h��̀��:���#���B���u�Z:���G�9�F.J�O2�g�^�fR|mg�c�����d�\�#�}���O��WT��M�����<��)k��{*�\�(ap?�ܢ����ݶ5Un�XA)��n3�����z!��g��޶)���c1��2����މj㛱�� ~�a�A�UΑ������-���1�5�բ�Qz3j���K�DE�GL�F2;�v�g���ѷCa�8��pj]1����|#"��:��W�l�2(���ݼ·�	v֧H�y����R����y* i���V��~5��D�#�� �)�5�acL�g�>)�kVwl�����Q�0p�<O��Gx����k/-u�0�yZ?|~�EBg��m�[x7���)5�
� �i@�-҈����H�EU��
8~^Q���})�K�a��s�7�K���5���i,G"}M�)A����l���h�EXC���YȰ���̥[Zƅ����"*�UQ����[Z���gG�f�I�o"�u�Rd2"�e��|�4�$��ʌ�|`L��R5yo�V�t��.�(� �� I4!�
���|���!�������j�7�%0IN`�wlb�!v��.�#�.�$dg�˒�?��蒶;V](0R.
�zUX#�{���VVu�S�4��G���>W0 reU)¯�T!I^���k����z���4�Ϟ�������"aXQލ��u�Io��~;�/+�Mg^Y�x��ܖ��)�
:h�8�a~�rz����ǉ!'�v�1�U�;�>��e��*� ��97r��D˳݋fSj��>�7�#0�P�QBo X�I~#9_���_�;T��1!����e��`������V�����*	9=��.Z�`'v�apCe���*e�s7fڲ6���?5����w����W����*$LO�m{z?�U�D�f���jkЉ�N�t���qLy!)�E޿���!uh��?M�����^l90�S��j7%�_���@B<�x������e���B �cx��6��@�_xbiHE�	��{�S9 OA�%2�o���.�c�Z$��;������p�Oၟ�1���9���](��Z|[^�
("l�O-�M�n���'+��;���K����8��3���B� ���@Y�7JFAQW%�M�.wo�Le��b:�SC�'�ؐ[� �\�v���D�`A� ۓd?��lh�~�	x��[�����a�XĹl�#h5��Bv&��h�E��O��r�Y�L�W���2�15�����"zE��L;��+�숭�'�-��SRs4��q�=�jEZ����a�#��h{鉮���ܜ��c��dٮ2+̍�e�v�I��L��� '�.!d���:`��â�8��ZZv�-�[�@�({�������n�q����S��H�yx�M���~��63�n��=���ʈb�Ph��;�*���C������bt+�o\��nP�Xw��B��@�*#�x��Ί<Yƪ��ey��H|���w���|�#(������Qw1�D����ܩ)�����^�|]��V3�?��Q��F���#r��J�+쳟,T����ϛ�Q+�廙
G8����P��+��E�-Q�}?�~<��xr�F[�8�`]�����0-)I�'Cs�e�K��ʮ����7-��JߚGa`ٗ��
��*��/FC	���l���ߧdf�V+1�Q\p+b\��;zN��6�*~e�]{�5F"�ƧM+������ꋱ�
I0Y��_U�:�	F�Ok+r��X�Gw䌼��O$Ae���&f���{�ڭ���=~m��f��젿Ń�2X�����!��02۳��mH�2Y�?ۤ�>��G��w.���t�_�b ����TL�<u�-�G\SL-9��2�d���j!�#�����T������a���j��]����!�l1f�cW�`	
r�	���l���cή�LƓC����V�.ԥF�6����7�:��M������P�2l�-�0�Qu`����b��YC�յ�\�s2��B�a��c��	o0��Xbe�����t	?�4����!��h��t��#k~��@�Ɖ��mJ��0�5yma��NX�z-��H	 7w^���6���[�R��v�ch{�dWE�]g���X(��4G�EpM��,Uc�?&���a7t���=1~�;]p[10�̹.��a�%����?���G=�	n��'��r?����ʰQ/���Τz{E$[��E�cyO����i)D+���	�{�J�$� Ʉ��yR��v6~$_�ߖ�O�*o6�L�!�Bn��q+�̍��~`?�cs��;��9��ā;yB�˪vbP��M��Vθ�m���
�غ��V�j�?Wɇ�2��+%����aj��wa��v�L* J �2lV���D����H����F��� ��_�`=I��7�ݎY��@��`��A�1��f���*�毫G�~.Y��)��[+��Z�|3��44p��t��Sle�(���r@����E3_
���N��v�D mCJ�N���@�W"eեe�݆�1�6g��<${�9���f�b�<�o�ޚ&^�1 �hQ�%��d��T&���KEv�)e�Kg(���`�r9��{xM�p�79d����{֖��j��pe�N������v�u�+�~κ�r���ﮜJG�N��i3���`��<�;E���I[V&�ݘ ���sjp�W��u�^;�y���ɒ��IW:����VN�Y�����u�l:=��G@BF���O�_����3~g��8���;=\9º}GfOP��T]� �c� �=`�)5��꼱F\s`H��L�}n�͡����Ќ�)�nt��]�Hz�m�.D@�&Q�
x��d���Sɩ�2�X��G��N�W��HU�k# ��=��܀/yK5�ߥ���';�j��K�˚�h���}��T��3Ĥ��p8^�j>����@|D:76ĸD��8D�I������	W��H��u��\R�M���i6��V_�5����a���A��v\�c����k��vl�UV΅L���0�UOOܯx��4��kЀ:�����Z�|:!Ec���l�x�y���	
Zeci�E�i�س�u�Ev��
B����W(��f�;���ҹ�E7����9O܃�
�,��3M�~��ǈ$�q����n��D&�a1�,��������Z�.x.�=���ЈP��>�(�l�Jl7�0���-t�q1k5�W�>��w�,���T��nX/�i%ve䠹}�����u�'e_'gDrcr��7��:m D��Э�`rlܱV��~�o��W��+��:�+�O��L��!��Uє:ҵ��!��J�� ��ٍC����a��t"\�����9/;&rǊ�Y���`O�χa<F���jN3��ᲈ�;ډ<"�����Ek� \��B�H��,����;�.���[ύ �L�����V���H'v"m�i���b9ް0����׫��d����=���`Z���<p��ޢ O��$�t5|Sq�x���e��+������&JA�U�_�nɊ�"��N��������(��2	m{[�V$�&��r��;�Ǜ;�o���#�J�WV�_�;Ƴ�h�R��|���H:QA�z��_(�F��v�+�}s�b��<���L�o<�B��#���
����'x*}>���tμ1����
�}�� we��?�W�1)��5h��g��3r�\��Bkt��0�vOkU��I>jU�����A8��z�ƃ5s`L���P�ۻl>f�/#1�P��oAo���}y9���� ���饜���e� ˦�q3�`'ͽvpj*��~�U/��A@��b�ue��U*�@7�{�6��?�
���T�PW�÷�hv�`T�L��m�9?C�D��J��%jЊ�$ l��M�L�d��&]a�`(S��.�uK�w�o�^��+봡jj��4� j����Y^�����}�[7� I�4����EVx#_E�i�|l��%��A ��2%�J��sǙ�K�HZ�/;��7�V��������8����z�(_(uZ]�E�t�l�(3l����ը�P�����t�E�e��8���-�B��=��Y��F�V$%�%��o�z(��Pc�O��S��DҔM[j�\�a��*�a�c ��?�F�h�I}	��.[3�6�}
�9X l�3�5�ԝvg�`hom��_xK����Y���8�\�3�5�2������T>�ߐ���xS6'���t8�su�_��=%�����ai�Q�����ql��Y���`f�Ӗ���E�v�!��M���!{O.b<7���:���CF�ĞkTv�V[����I`���=��0 �q-����_oH��S�S����1��<�I��О([�{��bV����E*ܥ�D����b�Jo�Sn�_+w:�m�k�%*���f�<z^��'8�^m�v�w_��|Q�l��(���Q�Z�
ڄ@�F)Tw5��=cU�7��?u�Q��ؖ���#�M����+���,�N���R�R��PK��8�kt��E
+&w~��E} ��<�u��N}F�~/8>�J]N��o5�)Ϸ����s�2�l���C�Dq�En��;]'`�a��������-pCJ�����9nF��H���gQ>1���p,��\z�XE����q�~�d]< tF.ʧNK�<,M���R
�h�F�6��F�D�+s2�X4��w%b9��;A�˽�ǿ�������?m�Y�^���M�*�6�2�n�����r�o۴qmi�2�J�?<��>* �G�K��8��j\�_�FP�F���}T��u:*vG��fL�Y<�����T�!���	��T_Ƥ�L�5�G��Ū�o�>x=���!��f9�2���Nrf��ok�Q�֮�'ߓz�����o�����j�����ڀ�q.M������3n�����:r-q��E�����bffC�0��7|�������3�~����0G��bFz�� �t*I��BQ���O�v�P�kg����@�N� .�J�J��� 8aq�4N�Č-�8��o�w�����C\[�ʪ�r�yc	��d�>(���P(�S(G*��p�O�_�cZe��m��BI�t�E�=),\~3�p�KW�M 9\P#aB0��^?��3=���?�{ʨC�7����Տʑ�/�o���{QG�$�WgE#�Z���K�Hi
I.��>m�<�N/[$>����v����	~�ߗ�@�|�6No��p�B�A$����N��~A�cty�\�`�T���%�y�2/�KAPȨY.�T�W�g��36�E�����b�j5���H7�2�FB&w���-j9��w½�vwJF��� ��2M������D%���3���/��?��NI��!��ѭ�\�$rY���1�U��1
����e������G�6�Y��� ӟ+pY`��[�3���4�K���T���If��L@��� 3�P,�Vî��TMD �md$�N�h@�=�eVX5�~��1����ku{�D+�V�ң���y&���t��3�hs�x��������UK��k�������g���g�'9���xN�w�X�H�S�i��/ә~�1���(e�h�N��Y�����',�#����f8黛u6�b�N��3�ʱ`�E���O�d�Iܽ"�~� U]\�T.��X��u������5�*_͂�:8�9�����n�����u��t:~�G���F0�Ot�E��d	xag�׈��i�H�\�0�}Ƞ�O�0�T�|�DV��>�X)V�M��\ԟ�c�>�
��b"۶��ѐ�)"n�������z�~��%�g��Ф�eK7�t���s�8,������l���U�^���^B@�P�ř5�ʢa�����j��FK�"-݉���Ș��8ث������P	8�;j���z�|e�K{>����4p�궞�D�m	8@�H���õ�R���;�i���V �5q��Oz�̑b�ַ�%c��@޳k��l��������;0��xO^�xcM��V�kq���˽;�|��E������[x��+��
���i­�J����rE�:�
��@a	�]�9�Ͷ�Қ_7�W8�Z}	���,	�dMT�$�E.q�'��o��������4,���{?O�QU�����x���؅�'jl>*��ͷ�J텦��iM�� �╎k6�Y�_�U����
ڼ�Ix`Ӓ��X�g�%W���,����1�������Nr�����:N���-�d�r�C���2~���2p��~:�C��P�L�aq�/n�hZW�]K�-׌�I��n���a�
#"�Ō�Z�P9�Xg&����٭�O�Ŷa]����3��5�	!a;{h[<������F�� }A,�E*H"I�M�t;$@��?<��[�L��Kf�V䆌H��Hm��\�}��9�š����������GDp��>��;��Y��pz���L�F㴕/S����7�b���v,�W��A�n@�`�ɫk�>��vf�T�-�Df�m<�V�߷���XG_�*���G�O���hN��#V�P�;��h
 k���@���1Qp�%��(ݶ;�ݸx��}�?��������BgW����
�U��(g�}_�;BR��O�<N&�W+��x��
��0oQ�Aۆ:��6dw1��F��W0ݏ\>���e�耯�1�ŉ����d9R	i����h��
Z�����R*1�v!���傒�
ª��z������@�gm��@͹��}�]_�{mC]ICwۀ��y�[&�n�׸�=�0E��n�	<Ur���S�$��,9\�̻۷�[�ڧ��l��@�S�r�G����^���#Ώ�&�_��^�Y
aĔ�z�+�Pq�v�Z,E���a�q��.^�<�=I��&��݇2�����S��k+m�����s�t���&��%8u��W����c2!� �sx����f�$��#��M�~����^�&�`��Au���q2m�ڻ9r���Mj'�r ������'Iר���ړy?	��Q��\4F~U�CJ'�8�,[�}yf������2���4����_�x�1���׎'����L��c�F�2���bRۏ/ۀ���~>��s��s��R�*�3��ߺ7��s7��bQ`v-p`���Ba���_��`�嬢���zá�٘��B�A#��ъzQ݇��M���v�?� �HB�����kTK3��	���k������?�^� ��7i�*겜O�;AFj�.j�{�l�d�WTC�i�$G�!$;zhn�'L�CZ��D�?��F��(�x��\'�iP'�s��I�C��M��M�+3�Tm��3�^�	�P��u����l��Ao=���Ë�b>536������Y����|�x�s��:eS�i��P[��y� �%X��uW�7�2I��Q�b����l���g	7�a�������u��^n
������c�&֣Ia"����^(���<^��C�43p]�_�q�Ըފ=Y�C���-0UBi�V�W���Åol�BW.���$�N�J�Z���X��>�J���ΗJ�W;��V)_�pw� �m6_Vw��$�(5��PlD�(���P__�dN��v��i9Lu��,l�:_����;�ݢ�O�9'UB�9V~}��y��V]���ϕ�=C{���؊-#�K�� C��� ^�ǘ#��e�$�sp�U.<� �3EK	Q�Y8lO�z)c�[;%��C޲���2WH����Cv�H���z��7�ӷ ����+��.�#9�����Ǹ�O��8�� Xs���Y b0�3�Uv�y�!fކE7.u?�����a,����s8��5�{��|8�.a���@(�T_��j����)1!{o�� b���;����U
���7XZ�C�Э���	�)y������Û�SU-2����'���&E> /%-ް�.��|{]GH� rt���x<s}_]��W/�t4�d$����\	W��M<�'�7vWΏc��� ��/	N�_�W�Z�/����������{��#�5d�P�Z�s��%ED��`�h��5y�^�褽���K"�2>��aw�r�)�(��J���+l��
:��e��qU�	Nl�v5�,A[J������\Ɣ���P�2g&�i����n��1�"��/=(D�Xq�N2uh,�4��I�{6�q�>|��;*M_���q�����{C競�5�K)�L5l��ir�����~/{6�X,����K���.�d�L\^b%e�{f��X�\}����K]WI/۸�Sg�����%X� �_�8��U�=�w�7/J�s���M��Z���ec�ԗb�h-����d''qQd�X�T���!�n�?�TLj��7�BQ�}�M?f�3�ǖ	�و����)���*"N���8��۩�fk\K�F%x�H��1��z�a^ǳCz�8�}�=��&�D�:5��n9C�a����R�!���(+�cf�\3;��R�5h_p5^�Mgi���xd��j��t,����,��t��h�g~�2lNn��w^;��A�b�zt�;6E�D�~�*����ʶ/��A��ӆ�3KV�w�~��������NLD�+3����R�s ([�ɢ�1y����m��S,_�G�F6as!(�V{Mɇ޺N�u�e��J=�c}C��B*����dǗ������
w�PG�ǂJ������u~3� ��E��D*�=��;^!���`��٩���j$�I����)��n� M�ov6.����t��:�[]�{5/��J�Ѓ�YĄx�W6�ف�j�H��(g����"V&1Ww��V�S*a��Ƭy�%]5����w�P��e��"x�c��1K�m����]���"�0�//u�.{��7ָ���U-�O5	�;���!�+D�ue{�7�<+w���0�%���c�>��D2_��}��֖����Z�	!����9��V^�4ㄐ�b�u��L{�n?�e����ͰxEτMj�Y$��{���p�^=r���W�Z�-����o��rS�wy�-R	�3��������6UU�o�u�� 4��R�ٷ���d103�
����W��jXΤ��QA�0�?y�d�:�`A�	�QBo�>�}cVIU Ag؇my��I�Ж�KD�z�3TCS� �T�z�L��<����7�%�`Ge0S)~h�V�p���Jd��-��Knح�`��S��<���Q��˺;!�~�P-k������*C��T���R$���%W:W̖�k���s�5�L{DXȽY%�Q�6��D4��ȼQX��v������D>�n-� ,?�3#P&��L�s�2P&"��=��E�n<rS����̟�����3i!�����@o�x�̠Oh��iH֊^��-J��J�Z��W��3�"xʃ_v�X��ZnA�g��}f��o��?��2C"Շ&n4l��X�|�c��`6:o�y�t>4�h6{ ��WI�(
.�P|5�!3�ۼ��,L�;�7�+�I�~�.9%�܋=#�-�$�?s�O��M���`lS��60���ш��#�h�C�u��4	��j�1>�4k0nA�U7̝�}y!�}B�[Whk��{���x u��5���Ƿ���X��l��S0�W-3���^;K������s'�F\A�$Be)��h%��/�yrϿ�/'�/j�v|֕Uqz�>��k��&��qb����"̐�$ �4����	`>ӵ�#>�P^�[o��D��s�9mC��-(a�~���MeP�զ?ۜ�M�c�a�*ק�"w0��o�e��*�77���6���?�R�Mn���W �`gE���]L���m)�M?p�-D{ڑ?��З���v��R��L��M� ލ�ƽ������t�K^�"�롨ijE��-�|��B!��u�����C�ר�� �칡�����(x�4E[<}*��ͥG�B�U �84%@��������CZr�;�t����������H㧴�"(,�{Zʷ"�rl��y��.�����5hw�	揬A��Ҳ�8��ׁ�:�B�����cY���FP%^��^f�o���i�HƜ^S�J��!q%[���\e��*oF�n� �i?3��h֛�	�s�[`[]�n$����l���5k$Kv��h\\��D���xY��¥.��@`25nߩ�7*���iZ^�O4�z�����'�'��!B�s�Z�L٫=�_/�Fx�aց���~�W�&�7@
F�}��-� ���|�7vI
�Z<U��>(.�u(��Q�:nd�p��k��v�gG[��,�����-tq� vq��B�!�H]Pxb�H�
�Ν�*yޖۦЋŭ��^b�{��U�d*I��Qw9��ؓbGo�M�n^��wg��8sl*qQ&����<'���t/��KDϥ�*�w���|�I���KQE�9�4��-F�)�h�b�&�
�qޤ��?#e@Q��x�1�#�^e�*�+��>,���@�~�_�J�Ui��	8��^��+STɰ�;�}��9<���F�F��8+�]���ʜ�)����\�ds�Y�<���1Y���S��h��`g���l"'�����CC��+�t}�h4�u���4K�1-��p9����z�p��ؑ%��~3�]	wJFp~o�[�g��K��#&����
W��s�#���F���+�MX�#�wrt���(�As�ݓ�ʽ��o�(~&��lm[3Ů��s�:�őL�2&D�R~:��n`���vmw2�VR?)Zc>�sDG������� p_ژl��ū)��T�
�uǺVGϊYL�A�������c[!p	��V�gTL���ټ0�t~�w!T��v���!�@ff��&��r����w��ȅ�Cj���~��߼�x��h����������M45$�L��u�ގ����-�u��\~�x��b�i�C""Ճ����9���0��į��50�b��g�"�]t�
�,:W�������7����D�@*���L�JA?���a��=N&r�-V��W�w�����X4�[�����sc6�d彨�����b(�,yGw�p�}�W&c���v����/Lt�G=�a~���p��<������a�Y�6bo��d=a;�h���$�}��F��%5/�B�ܜ��{�,o$��*E��ҥ���iw�ɨ�)p�Z�K���$+��ɒ��G����T~r�ߤZP�Y&�6�Nd�]H�B|(��?^����~�]>c�p�	���\a�cyPV��x��P��O�|�d�ץ;��������&�}jbN����2
�O3VW���mj�fw�]�v���@ �EJ2�l��a�Dҧ��v!��l&��d�{u���;��q�}$Yx_�f�ތB��1���ٍ��b����G�L2Y_W��M��+]Ф�h��3�� 4·E�!'(�ah%����<�!@��1�$�q3�и#�ʅ���D-J7��N��@��e�&2ҫ)=1�3X�M�4 ���ԁ����>j����ط�y�o�]}PG�P�)=���f�y/ح#J�k��jG�+ɚ2/!������"j�9nwT��vI����+ �2��Y�ȣ�D7CJ�~�}u���`;��s��?����Yݏ�k軌�ld1�f��h���T �"Gby,Y��R�+�몭��3���4G���F�!�&�N�[��Au@�C?�i03�^����iD�`�v�N��@}K�e(7ҐC�1�^�r�{����ɋ��`���o��;�����hd9��
ݮ�`ۂ��m�K�����}�B�y���6�9S4x ���j킥'��n��P^��Nfe��N�;��d��9uluy�q�(
q������]&<N*i�3w�q`��uKl����I��ʛ�dU �S����
�*��u�ˈ�����*�T�e:J^ݙ���&����"Qu��:Я�G3�sF�cO�1��2����gi����\,�S}���O{�Tp8���lT��W)h�)�Onb\f��5�I�0FOʹ୶�@�+L)�nX��Piz�=���Wy�}�ϛ7��Ȇź��J��Ɉ�b^�ҡ!�9NU"��Ӛ��p�o�6l+?5���sځN�2jI�hKYӊݛ����ʯޮ�}*��TP8qDcj�I�����|w���b�ī����˷��i����	�SHq0)��d%Rj\���`Qi��uV��5åJe�u�m.�t�'�	Nc�5d��`k��Nl��+Ak�h00�c�O���x�����k�pA���g���)|���E�4��A$;x�#˝��'
X�i.���i�YO�E��I
�Cx��F{S�陠i��,�7����l�Ӄo��,��mM�-f�$-*�q-���A0S��^�����,�G!�M�B�c�[�A�N��X��U�9�:>|���_��J�������@IƆt�kT�q��
>v��%�6�Ӥp�XB�Y%�P\�sB\�+�������z!rw��J.�:���6H�&�zr���I~��ڇ
�
>�d:�)�"�_L�v�%����޵/�Ƈ?U͌3Zp� �A�{�a �"ﮠ���9��&%�<0NM�k:�O��|ao�D�^ �3�2"��X�;��<I{���� �,_Ւ�H����M;6B6� ���t̙Ll/I1CEV6�HD�mf$#ڏ�M9�~�S�(��)A֑ڙ���0�)泉��k��p��s���,`���+S���@��!������AD5�2��ɽ(�YS4��5�&G)�VRm�q�V��|�dY������.�h�ߣ�F��]x=V+�;��h�͇O��;W�Q��i�7��(/���o�ȴ�WY}�xZ�X거���hByB��
7�4����}q>>B�i�O�đN�)@W=���ӕ
?�{o#����G��E�d	+��WB��\�H����	�Rt�1�$t�3d�|P	;sX�� -�\�B�2�wm�t1*n9vs�_>��dA�0�$w����٣�C��Z�,3���x���(��k<]���[���&�E�iz$=�$�����	�KHr��'S��,�>`�Ų�O�Ѷ�My�~)y@9��rz����࿄� �#Y	≮Z���k\��F�JgP�aƙ��hZ~���by�q�S^	�y=�v&>p���z��� ޥ[k����Тs)#�t:�s&��Ԕ8���W�}��^�!͎Xs�ߕ��-JŶV��ڍM�_����M���ax��Jq���M ��M|��	����?є�'0Ux�X��%�!?�sT����+�A4�oPU��f'7k,�t�y�0߸�;��t�8�4j�Qٳ��Ɗr��I����ǩ����zFH��Ӭ��R�w�ے�2��b��4es��doL�^0P�qb,�����6`Zo�-�A�u給Q��_�>�w�Fx�z�g���6�B�:�#��+�)P�zc�V�.%�e�͏Q�WfYVBA�L�l�T]vK�m0�g
	�=�2�����qC��w T?�iP�*c�����A�.|uth�x��LnW&>@i
zs�Z�;J��_Cl�ED׏�������t���'Y�P�;S���C�P�H�X���8T����l~^BeTP��u�v��~o
A�3Ϊ$�j��s�G^��-���E0��i~���x$Zڪ�Qe,l�b߷[ �)g�3%*t���p����uI%���4oh� |L��X���E��)�u�9[^ ����۴���{�I�۫}"��������Mz^�C��po騏��;�p��Yj5���Y�0��>��+�n}���QdƔ���F(�� ��J�x�`�8�����ԥ�Jh��W͐CV�~+_�q�R��Ȼw͑�$����Bl�O����_qZd�Z������J9^���Jvl k1����/����9��^O''�C9%��~�2�܊���om�4xr������؜����4� ����~�pe�up�e���$w*�햟�.W� VQ�E��!#v�[�z���[�����6�����; �U2�H��z3�>ߥ���M�+�وԵ:z�R����/3�&��\q�XEq�+�pb�"�����y��f�&�Ec٧.,y��	��ں��1s#s��W�~��{��]|�s.�[�\7@:I�_�D�/c)k�{�B� ��%͏���raU�e��7-�՟�����1y����ɷ�m\�U?a-�',�w&��/7�����6�05G��������<+C]��/�q�4 �K��u�%	i��l�7<GS�	��Ρ��Ax��������Y	 ��N����1�Z�C"�1�@�P�d���#{\-��G�cǢ�Y�6wg���^��ahb�5����ɽ���+W��ĳ�f�K��܂�zATJ��+>���o����'���I�~��JZ>��f�\�a��Iqt�����;6���tK��k��R�(!�qjV2�	,�ƹ�I�O�6�i��v;��n�_p��q�ʖ�FzhCy�=��pK;�dL���� ��̎�Ŏv/�;�X��[�[��K�� Ѐl��"�\0V�%wB&f>��X$- }�.��]+�I�kE��ɓ~��%j�P�,Y�J�D��W�I�*�l5��Z���F�Z�c,p���q-Xw��vهZe{Q�6��&���3U��X���G��z<�T��}NtFfY$��hXٚ����x��*�i���g�-jf���K���x���gb����Va0�9�U�8��R���0.�Lv����!���n��R��%���N)��.L?�'ITR��_UU^��ug{&��R�A#(g�$,���~ft�\��K�g�?�l��m�	����~A�yr��te_7�V�V�|��Tg�/ѮXA ��_��h�PZ��ʨD{���ZE�������q�~(�/�t�'eC�g�mo{,1'_��36�i(3дM�3G�`���M��/#cO���T	�����)�_��o����P��N��9T�o�Ӕ�F3A�ܢ�G��SD�G��V�;!��r`�~;��w�jv̸�\����z�n� �M�6����,��8�#{�p`�^��GF�ʣ64�7�w"Hݕ7g�%���	{1)��h��|C�X�A����]G$�����9ӵ7�2"�`S�4F5��2����B]�b�"AQ/�;.My7.�7��K9��=�O�WN�M{ߛs�DD"�eM/�7��<}�W�����,�9Ґ1�D�ڱ�O��֨�]�)�������%�K[2V�!v�~ bY��������
������k��[�냑�M^���ApZ�m=�����c�lʶ�t����D�#�b��m7R�S�3�"n���]���Ș}�A����tM �gRcϼ��OdCY�Vy�?z�)~ʟ|�E�g���oh0�@�y	�J:ޢ��*Q�e>��������_g�:`y��"F�K�0;� S�F�T'�+_~뎡B��\71r`����S;�[ب�ʥV�dz��-�`n*��`�]i��l��,+Q1e���1��P��-}b��%��?~��6��1t����N��)�P̨�-k(jSqՖ5v�yVf��Y�w��C��V�!�rc�+��H�������@rn�y���
��E��&�h�)G2"������yEn�0 S�������T�E��{9�FN|�ܵ�z�"�z���J˥
�]x�@"�T/�y�.�_7��&�� ��HO��X��:����D(!e�E7�|%<�l͉�+AȽp���@���^Dʓf�j1�.�$�o5�����rQ�@�V����HbU��F��eg��|��yg����-�񈳙-���p�=
	��������e.�-�4
���y��@��R��3��qŅMъA[���$��7�5 �b�Ri3���/d���\�&�6���U|��2�YH|��y�0���y�#�:a򤬡�nQ��=>�ȼ���pgp�y����h@�K�s����S�cjTm0�1���T��N�7w�`������S��s��m�%Rd@k-��Bnp��`��&�����^Qwަ���X��{-��k���EOE�ke'�܈�!}�T�L����.�kn��w��5<l�`�vY�e���y��Q��[�`鬩��צA����k^n�ϘL�ˉ�&K e�P�2�%/�)	�C�3n�j�Se"րk�`�A�Ȱ%�i�8/�R�A@��r����8sY�� ^�"o&Ȗ��rzZ,���Z"���L��gZ��g-Jf@d�o���x�^"�Fb��y�4�����i|F0q����o%̽t֭o� �+ CI��Q
�i�|�n!��)s'%�:�?��W71��Iq��������t�#C��$����=Ż�We��z�|�08�g� �d#T!���9u�L94������>E.�0n5Uϋ��,!4����kGk?�MKX�Zτzb΄�'�Y��Xw�0�{$x��u�IU�;����U�%ca��>�ܼw�)���h� ��Z�r��Ǜ҉�qvѲU	Ȃ>oﱟ9:����*�_f���X�qD����T�@o�>kε#��gP�9-o&MJ�/j9{���R�z��>��y�we�H��df��v^���%*oꡉ�U�F���pne�g*�H]7L��69^�?�K�����uW�c����EqwL5�;m�#�?lD�����/)�eu���~2L_ӭ�K�`�%L:�G���zt�`��2^���9�pj�@��ł��f8v�^�h�6�x�crS�@�7 �! �Y��S�x�%�E��{�oq�=�uڲ/ 5�Q%؈z�8ʑ��@Z
�3;8`��X�k�u������]@��LrZ(��Zb�����l$nUy�Tp��wz������Y��j��80���r�~B�T`�f`�Y@�ZF�8z%�!7���o��*����4�xS)�Oҹ��[/�0\�W§d��� A��?� fhn` 	�[������>)�lz%�5��vL�h�8����$�qk�Y�$�=����۫5�R���+���n�b�u��}�~'9�HԹH&sZ4e���=J�&�_2�van��<����I��1�������7��6�ލv����� �ful.G󻈎):4�������v�0�[G�ψ�ŕеt   8   Ĵ���	��Z�tI�*�� 3��H��R�
O�ظ2�>���& �H�O�QS�� y��]1��S�x%�D+QlW���K�4;B�^�?�vR���'�V7O�`����4y��Y�t�B.3	*���ņ�S�B���4A�qO����D���M�`��DO�꧇�=rF8��ʋ^y�?l��pS��(��$֊wo(Q�&č5o��I�	*��e�Sg|� 4l����	��'�'Y����O�牚!̀��t萧��ʓ%ӎ9��J]�f.v�h�џl���O	��07��hy�E�{)"�ҵ)u~2�ݠ0�T ��ݺ��
��rE���NHb2`SQ�j� H��(��|�(���5A��<�`ԑ��Q��y�.Zu�'�ֹDx�U�Y��''7�̀�f�W�+ђ"<�q�%�!2P�o������?�����ݶlD�x�O��Ӊ��ْ��'e^����$M��(B�Ӝ`D Rݴ��#<�Ҁ'�MP��h�)@=H�h��U�}�iɥk�\�;Z�"<yc�4?��.Pᢁ���_=�x��aSoy�JT�'.>��?9�KL%�����>������)L�:#<ɂ�(�|Y�����+����∕g �����?�1O��r��$���w�|0����]�v量[E�'ƐMEx���M�'A)²
�A��m��/�sUÏ��W]�'|�i�;c���ˆƳ}�{�JJ#.�qOp������I�8���F	x��Hf�ݿB��JJ#<yP�6�V ��l� &I�4	5$�Rq�ȓ	Ĵ   @�?�_]H��O�#�(�ñ�3D��u�   �                                                                                                                                                                                                                                                                                                                                                                                                                                                      T   �
  �  !  �   �(  �1  �8  �>  )E  K  �Q  X  Y^  �d  �j  %q  hw  �}  s�  ;�   `� u�	����Zv)C�'ll\�0"Ez+�'J�Dlӎ���4Om���'Ԙ�5`EK� yw�:u_R����՗��HH�h��$�^�ׅD��\�DHc�!aӇ��?q��d��?��Jپ	N��$oǶmEqq�D�����`H�2�B"�e�d����u�$@�d�']�|a�^�8~�:�jZ�S�"� b�ݥf��8ë�O�X���T�]&���ƏΦ	����ٟ���֟��Iҟ��rT?��Qc�/a�J�GDF㟘��K�^��4���O>L������$s����L��N�T���/��:&��Op������I՟���R��x�����?���:��iѸf4�p�Eؚ�HO�">��4!t|ı�
]Nհ�
�3���wZ��F|B��K�b�'�L*��#N:d5�$Y
"@<ܑ���Ov���O��d�O��OV��|b�w)"�"�#m{9Y�)7gN����.��Im�Vn��Mk�H:��h�^Mn��M[��J}��1D�?|Vл�Tg�ƹI���ȟ���o��d �4c�KM�X�y��.Z�k�A��M�V���mq�NHo�1�M���Rk���t����g�E#
��!`�$5�(�MƵrn�n�K3���Q�]q�) 7oΏB��9T��Ź�4y�vEq��z1�R)1$<�e�N�&�yJ�ʏ�r*e���ԬP�Hnں�M���i}�����u�1�;d,뎁κ��X�V�x�*��<#�@��~ٌ���Ψ�ٴI�6���׋ڃgf4Q�Q �>��=Qf,��~$����O��:I�ud8+��n�4=��^!%���b�GE��
h��c�g�����X�Z(�T�&a�h����1j�Zh� �i�$6M�Od�����j7���e���p��O���%�M"c�C�R�j�*TH�O��$m>&���O�ӗxf�P��g�R��%Kǎ�]�1�S���	�2� �!��V8yBm�8��O��	V�	/h6���^�iՏ�	~�P%2r@�`҅�6��;�F �U�'�����?��OİsS��06҂q���:i�y`�'�b�'��OQ>�zׄ�Qt|�I#怑�)Vl��8Y���.RvtN�P��K�w�`��m�3��E��9��|.��F����U�
T�}�s"Oҩ�6�7�0��wǇ9X���ٱ"O�9q�X!J�ԚW��?	� |��"OrDS�M`� ��s�T���d`4"O`��!j��R�&.�C��{�"O�H���ڔ[�+��:�}��	ğJ�
)�S�Oy���>n\"���·)�<�(�v�<AG
A�u���Pe��U,��RjPv�<1��\ % ��lF*E�f)�/�i�<��]�0)�U �̣3�Ƥ�գe�<!୞�HOm�E� 56bؗ�_y�<��.ȁ��)���B5�X�ӢMP~yR��8�p>�c�4��\CQ%�"��K��x�<�.ԗ�X%�%@�,À s�Ϗp�<�J�8dN��`FK%J��0�X�<��a	�.�`wmӝUp\��(�U�<��Dh)X%H&8��T3��Ox��b��M���?��M�O�v;�j].Um�@f��?y��:����?��O᦬����f2��F\�>��ĳ�e��!�b��(v���6,�6�"?aR�T
Ŗ���ȑ�X�����@�|�����2+�Ԁ��!C�*�L�$�N�\ˑ��R�n�O0�$�O"��.M��h@��˼�{� T�m����?1����U���+ 	�+ ����h7X{�BH�O"��v��U|t�
[nX����'5�	�c���Aٴ��'�����?1�j!O|j��qC-G]�
S�.�?��u�\+c��0����"��Y�AR!�%f24P��H�P�G���gi��g[H+!nF�����
�n�U�Є[�lQccF��uw�J#fL�O�LZ��%>HY�@� ����O~����'=2����Ȟh������9���V ãf@�'�R�'��� �&z_���V'��@����|�OR~�M�1m�e	G�K�e"H�g�i���'���Q6P�%3��'��'?��1��g�6�JnS:"uVس��/ 4�9�_�N�p�+`ؘ�1��1&��	
��}FȰ����D��G܏y�>��A�Im�\p�+ֳ`�c>���ڳ����=j�e�E�Z 6`Y)�&�9Z;L7��|y2�J��?������?���$�,ɡF�z�Z�"� !��'JDXv��D8t+7�1<���H)O�Gz�O�2T��3� �)�n	JB�^�i���pw�� M�24�����\��ğL�I��u��'�"7��y��d��u�6A��������s�Q}!��O�C��D���C2�����i�uZ�|�RO�T���>�(���_:r�9�j��AY�O�L�"�чR��� �N��"O�%�a��7+0̽@�@Ÿ) ��q�|"�z�B�OQR�^����������"�6 ���`g�%zmd��KP�,�ɄR�f�I���ϧ)���I
�9Bm�mݢ/Z�� X]�*�&{���kĈQ,z΀�agXn�'���gc��v�b�Zj��r��/��8q�pG偒C�v	�6�J��.8�'"ғ:�����0�'��`*�\
�� yӈd\������?�����(��,�Qm߻t�,ь�X��a��'�n���5,Z)�2W�R��ιh��Q�0��٭�M#��?)�"8�m�Ox�CĊ3/3Z���֘?��"��Ol��׵<.�=�2�B4R�ZMs�K*/G����Ot�ӯ�R�/!d��!E3u2�OnL�SŇ�)��6�ۚeG$�B�b�� ^��$>q����>#�И$�4���3?�I�ܟ��I`�Ķ$G Uq�h
)]^�`�sl�
&�%�0�	d��ȉ���8D��D��T4Ш/����>�3ĩ�Y��cPm�:vʺ�j5��y}r�'""#֖jӲ��D�''2�'"27��TP��Ήd{RL�fǓ�kj0rW��w�� U��QD�"�!�^b1��i'��i��ʉ)I�B��O�g]�c�Ą~�T��9d(D+�@�8�b>�Z���8���v���	�_x6���
�HA��'��G�]���Y�����E�=r,�'�~��4�7�܄�H��hतk��l9W�R;(�t5�'�R"=Q�'�?�,O����a��A#��v��<�����`_�Bάo�ԟ��	���O���k� �<��A��Fj4$1'�םy��!h�-�I	>HՅsհM����(O�X�O�&��-��ϝ�J�� $�4�����MԺD�6d��j�'�ݢPmB��(O(8i��l����*� ����*�y�R�'���d9�'6�4RG�-�����X�??�Ȇ�2��=؇��U�։�Lݠ��%�tY�O0ʓ'�Ph���i���2A�AV�
>�c�
U;����<q��?љO@i ��/N$@�bO���d�yH��P� ^CQ�u�7�Lj-N|���PcQ�H����S>n��$n �[-�����j� rcID�6Ɏb��U�>"���C�9�Q�� ��O��D�M��E]V����:0��*�/,|zɗ'b�4�zc�ȹɖ.4���R�$|:����:�OP�m���v���dK!c�Zu��p��Dc�4��D޷_d�o���ȗ'\����KfݵQ�֙�cώN��|���������2`@w
=D�c����b��E� �
����n@�r��+�N��"�ғ_�<B���б� �7��L����yYT�H6��	#p@���~b��<k[�4S3"B�gS%�z~�FD�?��-�&�'��O��	�-�<a��]�a9�i᧤4b��'5��T~�-@.møMQ�����p7N���OJXo��MS��T�S����%�#5*��U��?q�n�1������䄦d�	�h�,0��hE�,=�!�D)u+|�3��a+0,!�����!�R1BP����C0'��"��]�r�!�P��@�z�>���a�Q�!�dB����[+�N�@����!�d�z̮p���&٘��$`�d��ɰ;?d�����P>i�(
�EϜH:�D�]�!��I�2�Ȣ�我l��,aE����!��]�q!s*�&W��9Yca��;�!�$���$����G�� 		���3n�!�W�G��X�E�Φ*�i��E)x��}R���~BÉ�VAl����ش<]U(�i�8�y�(,��v�`��ΗIp�(5�,D�<J&HFahH �s�+T\�Z��*D�PI%��a��e���FF1)�M'D������2�T��D�f��\x''D��s�Ɖ���\��Oߩ?��st.%�k�\F�4B�Dx,1J��ְq��L�����y��>a�4�0Ȁ<A �l�'�B��y�сM�f���5?M���rfQ�y����4B��G����iW��y��N !�P,� =�����!�yB`
,�Z�kT��,>hI 7eȑ�?9uE�E�����LZ�lE:T���&	� e�Qsvl8D����a (]xO^�o`�8R�1D��z��Z�1<���k\*"��Q�c�$D���u�#~=�Iy3BV�K��Ч�"D���w	Oc�2N��N�i��+<D�`��[�N2��JU�Őiu,,�t��<ATĊB8��Z��D�_��bB��+zF
����7D�� ,��G$(�v]��I�_ �%�"O�])�hҤfĹ"槔�F���u"O�yaQ.R�*shi�RL�,l<$��"OZ��mԤIT8�Rk(\+�	v�'�,���'��9�C��9�*��ò��
�'`��A'.gN���KE�2�#	�'=�"v!RzZ���B��
H��Փ�'������d$ �AJ��T�;�'XV���� P*���"�8z�vD��'�F�H��َG ����ŝ td"�����]n�Q?%y�c~G��� 醤[<���n*D��CBl�2WA<4����0\�zu�F<D�d�n�$51RA��*���S��4D�$c�D��m!��ӥ���3h>D����� w�iyf	�9|�`9q�(D��8�@�/7[h)�C��t�7��O*�D�)�'5M,UX����Wxf �DC��`�a	�'��:���'>mjm[h�����8�yOA24�켫��)�����W��y2*�E�vǍ �$��Ǌ��y�N�
)H��r%�yL�CB�;�y���D�:,x2OF�p1�����f��|�a
/Dۖ�Q� ��	���y/
�M�2\���D)��B�nS5�y�֫4nL����� DX�ٰ��yR��1���o��N��Ę�I��y�)G7&x�<�&C-J|�s O;��>9�ϐD?	D�Ց/�d�U���u< U[@H�|�<�2͊� ���3��S���Fi~�<����DNޕ��dK�>�iDz�<1s�7.{�Ա�ǝ�GvV=@�m�<	��.s��}�ՋAuNAp�aj�<	��ÓA�fI�4�ƥkV��;���A�'�����ąq�ƈ�u툄c2�:.�@�!��s`4H�aJmҦܚ� �Y;!�Bb��Pp��q�:i����{-!�8m�p9d�'���%�J�m!�Ö���c7�^�DfE[!ʅ�  !���̖�Y�r�(�/R8%
���Of�D�)�'f��3�R�gB0c�NC���a�'�� cN�8��-p���3q�̫�'�l1�:A� p�d�&eO6�+�'��p�c�R��(�IZ�Q��!R�'���4L��`�N�`�HXC��8+�'�ޱaT�ǂD_`��%A4S�y�.O�z��'/�Q�׮Yu�4�c�^2(�x���'�T���E%��℘��Ek�'����MI�7(&0�&f�)~A��p�'D�a��Our�s�*G�61�'�8��e�l0���ŭ�j���n�9���<%�M�~�	(T+?���>��HR
�N�"(أ����%g=D�����B���E�,,��č9D���R�ثS:�A�)ː�����F�<��❗5Ը@QS�K�{o5�z�<)wl�<�����D=ws�U�˞z�'4�`���U�3��R1�������EN]&�!��X�!/�Բ�'�@Վ=�$�1�!��
a*�a��*t��`��,ߌI�!�Ċ�F�1�g�ք�N�i2C��!��@L���WOP�Z��]X�i�3�!��ͦ:��p�#-����p�� �Re�8�O?�"�	�/}��	�	E"�ry��^�<�gB��$�LZФ��,���Y�<� DD`��ۙG��k��;c[� �"O��#���CCd�A&��`]Ԍ��"O��zPE=����C,px"O�����D�x���0Z.qڗ\�-(�O����m��rT��p4��5K��"Ov��ԁǌk̠��H�6Jς��"O�q�B��c��
bH��L�����"OȽ�� \A�q���v�.�hQ"O� ATQ�<4^�:q�L��ഓg�'Ih�'����1m�{���؂̒2p)�eR�'[�y�q�M2w��鱂)WZHL��'묌d�[pL �b����|mh�'�^��fG=o���a�o}9���'�葠w!0�����J�vc*���'��p���d��CEmZ�n>�uی��L�;�Q?�Qi��� i�͇D���pF.,D��c�Т:�0�h«)e�Z%���)D�|���õY�H�����IZ�H&5D�\iD�6x%niS�A�N�t}y�-D��s�'K� 
�apaý_���Rn1D��;�n��-��e��� �f��i��E�O��#5�)�]$��@�0�d}�7�L w��|q
�'@bd2���~�2���t�h�p
�'�f�G
��oJ�p4�+kE0}a
�'�� �6@[s����$M���1�'�`��%�½vEة���]+(�T9
�'�BYW(	�Ycf�C  I� ��)X*O�pbB�'}�- �����cԄ9��+
�'�R@p�"�2r�)*t#,b��P�	�'�>%�3���g'�Ty@���Uh�1B�'�R !�6-c�Уh�Q����'�
L�ơǡXU*eo�2GxN|��8�����Zq�11�E�&�iƥ�s�$���%{QbV�(6p�ҩ�3����xU���*�5[\=!�P&�d��.�Tr"B_/Xs����B�I9"x��Y���A%�+)�P5ң*��58xq��'`N��JD�^�(���
�$J���E{�(�'�����`���R\�a�-���@�"OXq�B	�D`�(� �R;�l�"Ov ӄ�6c�h�XH�I4&�"O^�;���m�hY�f�>O+�@)"O������F�T飇I�%$ƈ��"O�`#PH�"kxЗ��#8�)��'z
�э��S�1��۱�ǌ $����És7���ȓx�	���=i�, ���-%T<��S�(�
e�]�[vܐ@�K-K0��;�*8��26����oҨd���ȓ/4��V# n��Y8�cOlɆ�F������&k�T� ��Y�F�'gRL�
�[���!}_��!A�<���ȓD+6 ���7*i��s��ԮH��L�ȓ>�:%Ӈ`F�?b4,���܅wla��c��娄��SĞ�y��R�2)�ȓL02U�v
[$'r�G��;n�����	�Ad�I0�]���� �ȱ���v> C�Ʉ+���XG"�@'��q�/�8$�C�I(���Z��ZRK( ��m%p��B�I8|p^a�0H�$k25�W���Z�C��$XI�`s��,ʶ�8V@O<OW@B�I �nx�q�\n���N��P�ʣ=��/ZI�O&�����B	�9c )��ۘ=��'���A-�!j��@I@�آ`w<!Y�'Z#��_\] ���LlA3��� ��s� qU�80o��1���4"O�E#qG�AĤ���Я)�Th��"O>�qq텑:��,ݗ�N�[d�'(��R���ӵx���A!c��A7���B��`"���6�$�z'�O�~9�`Eҽ�:Ɇ�s�y�"�S	zh��R:
��ȓe5c��C�&Q�L��e�b� M��G���X6�'2}֬���[�%�\���^�J`bI�v�l�[�AH��1�'�&�H�7���JԿ >&m�X<�A��*�Fu u��7@� 0ఇ]�p�d���*�����Ht�P���S�F�؄�lczm�R��$�4���NI.Ѳ���vζ�x�*���@T�1%�%[\`��I�Z�����:lDd�d�P��s��	^B�ɤi��"�A,�����uvC��4p�0��F�V!�A{KN�L�,B���}u��5o�ȝ�uI�+��C䉤"����-�P
�M*�h޺:
�C�	�;,St�\� �B�*�L�b?ў ��1�j����9X��ڣ� 2Vw�a�ȓPE @�sf%I����� �����me���mED��/B @��=�ȓS$��;�T=!��л�NA;sN �ȓ~~����H���ik�Dؼ[�Xфȓg�bHj&��M1�}��	D:c[v��I�f"<E�$ɟs��-iE�X�rX��mW!�ʒsLAg��#e���F��K!�kf|��ׯ��6}��C#B�!��
�(x��d�e6&A�b�+�!�צ^���y�	�:+�(�gbO,u!��[ݛ����]��*��Ŭ'Zџ|��h���M��j�.�?��O"�����(�`��� ^�tM"�Qt�2��?��q<Ph��� 4� 8�)�Y��O�$�k�D��8sHX�bP��BQ0���[<@NX������D�|�Aՠ�R��7!���c�+�A�'�6���?)����Ώ�X{0a��I�ظ��N��D�O��$I���+�ǉ�h[�Ʉn�� �'�I�J�9���(q~Ԑ�fgO��e��a��B��	�.O��'���v��hկЪ[l�I`�)+!d����^��}�6@���R�����p��S�E��2���ڸ"�
w$�'"�\�Q`�X��y"ğ7D(�Z�ρ�5HNU(���"(�)���z�'^��ug�M�~���8��	�l��Γs5���I���'���Ԇ�d�	U���j�P6쑸�!�[-J�q���ׂj��x�*X�$�ўH��i��g������>�z4�TΒ�q�4����O��� p��� �����O(���P��ث_��kp([�i-q�JBW̶�O2��D}8
��?#<)�oV�tҺݛȈ(I�������� w2���sm�Gp��g�'ڄpB-_<Fm�{�t��O�x��'6b�	�<�'ظ(̅��	1��	y���Q�<1���eĴh�-�b
8)�o�ПT
��4�X�$�<�s��5N�s���8vɠ=�Ł����R�˸p�@p0��?�������?Q�O�NhA�&�0Om�h��Ԁ �|��B3u�d�`��΅AÌ���S#E�l���ft=�we?;J�C�-ԯY�Q4��[؞��5��O�������p����BĻ%S��"C��Ob�=���$�N��Ki�'*d�x��ֺZ�!�D���"@�$=�T���LT-~��I��M����'c�H*M?��8K'�,��
�HG�0CG�?D���bZ�G��!�c�:]v��%�<D�\JAcD<�ꁺ�Mݿ{�Hܡ�C?D��k`�\��d\۲nF��8���0D�ر4�V1!@0�A��<B���� $D��ZUMM4}��)
8Z]Pa#��t��#<��Z 1�+���@a��AS-Fˈ��F"OD� �W	p�J��ʗ 	�L��"OZ�pae�%\E��V�v�+"O� $�a�D&'���	��S�
�Ip"Or�z'	$x1:؇�ќ`ɶ� "O^)@wK�M4>q92j�9(&}��J��O,�}��#G"K.I��t� �Y��Շȓ>��B�dR*���k��M,����E��C0d�����۪���}T�M 6�O>I���¢j��dx�ȓ	��$��N�YĤ�8v!����m���[�$3{�t�I�3\����	J�,��d�R�l�yS�
�Ob�d� 3#:!�� 5�dp��)��Yn  ��<2!���\o�����Y�;�)����X!�$�r��mZ'�/����0J��.-!��w,��[��Y� �4�p5*>dџ\(sd��M����?��O���+ �\�2�IR/�Cv�@����"�"��?1��1�|
������!��8��׾}��U��ۈO�X�x�Ord@�c��>(��?P�P���΂�ᓯ�
X��'H���qt��=h�6C��18��p�4�	)_�Y�BM̵p�"���Jy��X�GD�a)��){ ����eH�����O��D%��?��'��3ŋjW��H����yZÓ�hO�\s�j�1"����a��%�&��`�BO��҈��"J���鰔��#ތ�Q�*ـ��I{?�
�T>�ɢP$��%(S�"��x�ۿM[��K��Ia~&>}�H� ��	���'�	W��"X�ҝ�C>$�ء��/}r*���E��'�EP��U�s�Me��(�6��57� ԥO�P�O�ꃑ>)�V?y�ȗ���g'R�0��+C��dS�[�pE�t 	VS�	���1@&�)�� .�B�ܰ��Ƀ��ɻ3���'	�7M��>�S!߭u�r�$��o�ɇy�(ҧE��1g��`�Ā��+��k�	�t��4�'�Z\	H���<9���r~�'��J����"�⡱��]�dTj��$[��㗦ǟ ��-��>%��U�~�
{��\'2�p�"���OX-��'�&�A�O�s�܊Ub�����ED��ə7a�80��Q0��OT��aoJ\�����^?\��r�<S������.�)���<}0��G�N;�R�lZ埀$��@���I_�ܴ1����Hw6���"ϡF���'E�'�ў��;��:�W�u�:\(4�@���y'�xD{���a޶w�X��q'Z�Qr8�����yrE�p\.m�bD�N��8@���yb�T�e/�p�2�W���"7�y"-��d��`���m�2�yRl��It�KR �Q�lRv��y�߀keFBG�4��-��D��y��_���&A�WC0� G٫�y��)�T!҅-	�P�����yr�Bm�Ěd����P��ʢ�yrL�f�A@��$�%l8�Ox9��O�{�'O<k(h�@` I@��	�'��Mh�l@6A>l]��`��'�aӉ}�HE�z�~�2��H1���u  �|�lD(m�\�$LO�W��H�j%*n�34�¾_����������g#u��<Z�JB�c���m;k�`��Ϥk�Ę#'_�iJe
*�R̌���M�/f�u�Q'W����0���)�:�i!Ӻ<��3�V�ga4��Hݛ�M��遰;~���Y)>	$���
�=�r�'����%�i�An��+:�H��HU0.K�)r�Z?�"����Pu���d#��g�}3ҥ.�D�fX���bG�uq�Q����u�DQ�V�'肉�U�9���x�e���le%�@3��O����O��?��L��TR�HK/Yb*�ؤiR4v�,�	mX��DJ��\��T�U�S5n��?O��Gy�gۯ@���`��SA��i��'h��n����ȟxC�Ϻ&��\������ğ�N��Q�v���N\&%�x1v�܄[�0|+v��7M��Q[�Kp�l��6��w̧B�,ٹ�I�O���t@��a� p��ѕA��A�{'�}{5/H�'%�]v�R+�$�>�Dk@��y��&]����0-ø�^�!�?xj��d:?9c*�ٟ�>�D�O�6��(g�~�S3˗0yL�s���;6�*��ē6���P�Ե$�,p�R�W�i�O��Gz�O�V�sˆ�R^r�;��4VK�P��۱)V��۷�	��?���?��QZ�.�O&��w>U(�!����x�lD�\o�ǉWJ����ꂐ7����X�P�&G�?�Q�H�� R� egE�tʚ	R㒂 ���#�Pt��z�n�=]nC�cӪd���B�'�4�Q��G�$I�)����$���u�C�?1�����h�r���-3���Ջ�7bY��*Z��y�:/6�����!q&P ����)и'��6��O�˓'��I��W?�n��qe�޿B�j�av$�5�(!���?頭��?1����T�R#9�BMq"����yAMϰX*��L�1M館�Q�S�;X�"C���@����ˤ^��0v�Ɩs��CM�I�H�%dߒT]��1���f�'w �����?�OR�F@V���m��	�!�r��1���O���$�`>�)�w.ضF𴬁`DE-�����LT,���1M�����C*o^����d�O*�5��QR�i!B�';����l�m���ё�9 ��QiÉd������?����?I�y*��I�ʩ#%ϦC��U��i�O�����)�ӧ[����T�����|�j;s�Ov%�P�'1O��R�p7���]�S���?Cp�)�3"O�}#��(M��Q���*"B�HRG�'\ʢ<��K;�`r�,�.5� �o�@?�	�(�t� �O�4�XPB��A�Z��%�ȓ�Y0�ks�i	f�$3ZP4�ȓ"F�ɡ���	����"&*R�9�ȓA ���ɒR�R�E�B����h�b��ўQ=��Pǩ
 Z4��2�e҆���{��03��)C� �ȓ/ �}��,ڮR�^uH���Fڍ�ȓ?ځ����-B<h�M���T%��5������l<�P˓�(�����\��1
���'�4l읽I�C�ɧZ"\2��7x�z��ޅGbDC�44�HL@3��.i��Y`a[��B�ɓj_��#�ř)��8�Χ#�B�ɪ�k�ز#/
�e�Q�Z��B�	=SG`p�򌊲Q�M��j�X}�B�3V����,`T�}ɒ��a��B�	qK~e:��)��h��M�jB��"\��lA��@,&Ѽ���H��	"B�	,\�5����k3�X�OV�4�B䉴
Ȝzb�_i&��R#�� �B䉙`�sc��U!T)�`ՕGo�B�I�=�L�2��xP�8��O%z!vB�ɱ42�0�"��7@8-0RL� �,B�I�L!�tI+�9���y��!v��B�I�[/\H�3k�j�ʑ���@+	6&B�ɑ2�~���W�&ݴ���J�>��B�IFY��ha擿}���I8X�B��x{�Ih�.?\e�葻~jhB�I�5͞���!81�>��`�ӣbp�B�7ɮ%s���MCV�ɔ.ͅ�fB䉸`{>�+���bA��D��ئC��U)S��͸\&���b�ίd�PB䉄J��|��d�6h&��S�ha<B�I�AE�1�0�Z)r;\��'Ə�2YB�ɩP���@ ����<� �#�M�B�I.�@�f�&h��͝5q�B�ɨL.4�(NL8� :�$K	w�hB�	
J� |K��y:f��GFA %�!���J�4��!��S��	ʔ���!�DH*"�-�6ŖT̓3�I�3�!�d�Ǣ�0�5F�}J�җ�!�ė"��4Z� �K��2g�}�!�D�|򖘣���=�ցJb#�}G!�%
�4���#a�T�W��)E!�>Y�H������1d�F�y2!�ę��Jy�OO�I����85&!��A�WJq;k�:X+zT:5 ��!��c0�@�g%f��S$!�� 6QK�,ݖ`��!��M�n%ѣ"O���C[eĎ �E�#3�F%!�"Oΰ�A��&�Zt�tdXa���˂"ODu�dE��3�h\��c�61VY�"ObtX0L�m����3���%#�4�T"Or���G�I��X��w��	�"O��h���>��^$#Ԏ�q7"Ovq�!�N�,��K��X�A&\u��"O�Z��J�"�.T:5K�z
�@"O��@�:X�v|�͙2���"O(�p���_QZa:���e���HV"O�Pb��ʶ?���(V2D^,F"O<�9�Bˣd�����`2�:'"O� �t
Ә�|�PB��0����R"O�q뤩]^`Da�2o��QsFYC�"O�-h�mƀ! �$k1�#/{�}�g"OAʥ��	T߾mZ'M@�l����"O�E�.E>����ʠ+���"�"O��@�*B%sK|(��AN,(��,i�"O��5fڲN�L��сW�=�5��"OxaH���@z��`��,0P<{G"O�"qb��gК�(��O�"��"O��P�#H_�0�"�R'n�֝h�"O�$hP�D�w=��*TMW2<�Tl�"Oa�f�1JE"��Uj#C���"O�����ǫe|:J�cכ]�B�["O��!�#��XTi�%��B���a�"O�P  dS�Sx�ݡU�B;}*YI�"OD=�5)L�����n�x�M�""OȈ�)O�y��ȩUk�;A��{w"O
�(!#<�Dȧ녘Wr9��"O��*�'���V�P���
8`&"O<q���Gn<MU%��y���j&"O���V�L4E�]ƤV8$-["O I+ ����h1�ƌ�m+���"O~�C#�D+.
�!Z��\�a"O�Y��D�n��UΔf��0"O"d��(
��4΀�)���P"OZ9a��C��E��j	S��y�"O2mZ���0B��<�t�,��5"Or�8��E>bV��PWH��V(�!�r"O@E0��L�4�����>4�A@�"Oz�cA�xl��bE
C!�� "OL��T��r�,	��n���7"O�)�F�,H����P�Q>\�a"O٪�`�uD(���BH9��T"O&�b����0��Ƶ(��,�"O.i�ECؚ����p̘(l��q"Ol ��g"���� ߂,;�՘�"O��0�l�P��]�����-!�$��M~FMa�˙	%�Î�n!��V2�ar"\�&��8����1T!�D�*2�}�5�U7hx�M�̐,Y1!���5tc�ٻ�,�TYp�)p��<"!�����
 IL�xޞ�� O�82N"B�I?&p��R��1U2(�>[B�	5o�\�i�����'Zz��C䉎SGz���ҏV/2��4oٲ%�C�I*RX|5�F-'7}a"�)גt�C��o$�M)C�]�O�"Z����p�C䉪48���gmE�)�ȵ w�G�K�>B䉙3hTqe��'���c��УB� B�I6$��uk���+��pd.�`�B�	7b��|�D%ZM,�EabB��;�B�)� �2��:��i���	S64��B"O����P�RA�@ a�,x�5a�"O�l*D�e��%"����"O|T���S-Ud�q�*D�B���"OЉ1S�͢�*���A�e@�"O1P���j	�D��)sl�i�"O��S2,�@���^�-��iX7"O2�K&D
��Uj&眱2���@�"O TXp@�#i}2h���s+��Z	�'A�ST�ܡq��C�A��(��	�'��`c!F�1E,�x��̦6'���'��dď�!�zg�� 4KR�1�'6u��K��z��V�2
F���'ԡ{R���=�FF��$��1��'�0|s�c�)sdMn�W�yq�'���>V�b�2GjJ~�8
�'��	��H;qs�[�W]ƼP	�'�R�*�N����%a�>:H���'��,��=:� �����u"���'��t�<_���P�!���r�'���ړ-�-g�ҝ: !��%o�QP�'�jрw����:P�ґl��'�z��ˈjB|����lM
%��'��8�"JC�T9��LM�k��A��'E�s©ڦu��EzpC�l�DmZ�':���(['t��O�*Y�l��'G`��QhQ�G���ϘP���q�'>��֮�P���0'@ў�ȹ��'��xkb��9D��iF�\����s
�'�ȣ��C�0��� �6K�'��]q�-ߍ���T�ђ{&I��'��x+��k����T�])H5�8��'�,<�j�=z�	$�߸/�μY�'� \�ցͪ�.�:�!��c�'�\��3
JX�=�Ao
<o���'|���#/�0�t�p���L3��B�'�u�Ռ�1j��X8!�H!W��I�'q<��_0�쵐gL
�O��i�'%�P�p��:\����=:0�
�'�葘ԏ��\e����OV�l,H�	�'&��@�$�,Z�χ�2$͐
�',��b$9L��lPf��%,�����'Ʉ��0��FQ�͋u��\�N��
�'"�}U�V��H�4D��B8���'�\Uj1`	܂"�k;|?:ec�'���[�f�%��鹓��kf:���'���y�!��#I��hCd �h��5��'��)���J$��cf�N�Z����'�>�ICfW!f�VL�E �W�*�'�(d9G�ޡG�	"E��I� ���'�$�17섁�$��O��IW,}�'[,����|�H�*��8:`$A�'1>�	�'w�tp���(L��'��M�'a�l���2���w���	�'��Pv�ܬlu�-#R�Z
!�����'\��#�JN�<�Ȱ����'��u���[�/��$
��P>�
T��'yΩ��@p� 9A�Ū
l(�Q�'��b�)�*}�	V%�8��'{������5���{"�9OB���'>:��dϙ�JE����@�ص��'O,�����V�1�1-��Q��'�Hd#��U�B�$0��)ό#�.m3�'�1S�I�,��Ѣ�+$:��	��� �4+*t�|���7D� t�"O��	�bH5q]�u�2�X�U���i"Ona$^�J�Qw ��>�x骤"O`X���5
.U�F Y<���f"O����7.&="�	�C�X��"OX�s�L�l����d.Q�N�����"O ����˧b��80��$4���"Oxd�fV.�n��B��3|x�I�"Oz���ԧv��y�Dj�+b�֭�"O��)Pǂ�\3T��	�"z��<��"O�œ��
�6N��ͽ}�V�"O���"�	��܉K_;"�ʑ�"OΨ!ӣ��R=����=)XP�e"Od�P�P_���f�h�$	�c"O�%"w�P	������6vvycb"OFM�n�"<P�b�e��fp���"O6��&D��*\a���Pcv�"OTY �"A�"-�I)6F,!i�X�"O4�`b���b�8[&cƧz�^��S"O����� )��haA׽G�x��"O���a�,�N��O{�PXSs"O��B�����MY�g~M)%��E��!qE�AC��{�߄r��y�_�KB)�!�͝�`Q4����y��#c���b#�U9đQRhS
�y�C�zQ��[3Aޟ!�ʔ�E���y")��<|��1�1B�źG*ƍ�yR���L?�Y�7�#m йإ� �y�O�Wi����[�E@š=�yr��Mv���mU�Q@L�k�
�y"�F7�=�S�(�`a$E�#�y���!�$5�w�̠6�D<j#�0�y�ŉΥxb�:-�L�gT`�<� �:K�H1bg�YwHTZ���P�<��!��#�QR��KP�#RCAd�<���	�Қy�s"��(��C��a�<	��N����R D���h��a�<1#�ITX*�@�ep�N�}�<�h/[(�p�i{��sw�Rv�<��'��\�<|�DkU���8�&�y�<y��J�zs�T�c �"pg@[�<�׎>S�9��섍.��*ӏ�W�<1�	أb���o֮ɸ
T�P�<�4��,pB�E�1��mt��[�͙S�<i�E��ѣ@��B�9*U�l�<Y��f�� hy���b�D_g�<ِ���x��	�n��B�*Ca�<!4 ��k`��Qg[�0-��+��@z�<�DA^kβ�+S�Ȏz�X�p'̓y�<�`8P����Uo�\4j\�C'�_�<���~����t��~�LI#��\�<1��Z!y�>a���J�M�(Xh�%�Z�<��c�.5ZH(j�D�~C����m�<�vς�Z(|���R�fX���i�<�# \�2.p�a��	J< ��I	l�<1�GD�=����@�C Yt��[�p�<�'��x�BD*�	В8C.A�ŀf�<��Fߏ~��PBb�U�|�����Ox�<�eɂD�@���^�_�T�Cd�v�<��&�q��!�C�
�j��#.�n�<��
e�D��pB_y�l����A�<��G� z��cAA� ��Kw
g�<Y0͎,O��ꓢ�
) Re�k�<ᑄI)-�����a߹8��� e�<ـ��ق���D�XC������<� 襡ǧ,�1b�Ú`��f"O�q�Rb��Na���-E	X�����"O*��͟U�"�M��FL��C"OBl� r�>�@�#�"u�I��"O4Pa��%!O mѡ�K"����"O���mH!H���ن~mx<�@"O Ej5D *���*K'R|8i�"O��:AD]�I:5IU��	u"O��CR	�{Xd�V�$̦�hV"O�襂��B0A� �۵g6�-c�"O��JTN���$�� /Hk�"O  a (���.IH��,"�X�s"O��*p�]F�Q���^ls�"O�ɓ��9=B�9��F�,`0��f"O��HՅy�(��D��!;V"O���c_�%5�[��e�� #"O�a4c�\�z0
�O�flΈ+b"O(|�7��G�椺�A�Hɒt�"O�uJ�"�nXgkʋS���聬)D�t9$��(I	+�!^	�R��u�:D�\�œ4��MP�䉼2
T����8D��q�%Z,D1x�fLȄ2PTq�%D��u�ܷY�0Q�&�K~�|0��5D�i��%Zӊ�����a�0�&4D��b6aT��B��hé��(�vO'D��JU��7����"�-9�L�E)T�T���ul�E�	S��(�"OP���ڱj��#���W>����"Or��m�tH�����"2~@�"O�I���#N�6����ӶuZe��"O"�B�i�&O�PDpQe��j���"OZ�	􄎝Wi.d�����~�[W"Oν�c�� ���Ά�`X[�"O���S�
0/����k�4v�b"O�p�ޞ^x�D�C �|�kS"O��%�_���pg��^��J$"Oz�p�FS�@�$�G��6c��2a"O"�3B��9�\���D;Q"O����[hs�,�V���7�H�""O*�Ï�%�aj_�DPȂ"OV�(f�U,9z�; N4>�^m�"OJő&*@�9�����ԓu��$�p"O��fo�!q��%@�dV�4�X�ȧ"O��ؔk�Au���a�%&w�Y�"O���F
?%���4s1L�>!���ŅۆX��$*WH�>8D���"O*q
A(�'�Q)��5���"O9`�LV(&D�h�Ȝ�w��"O�1�(�L�����AQ�X�"OH���y��U�7G۬`VF{�"O�q��`��x�E���@�T�1�"O�īF�-|<�Q4�څH�����"O�!sc�Ք |�q��
`���"OԬ� U2$���k�@�]԰P*!"OHi�E�^�i��[^�p���"O��#Go�u�ؚ��j=�Eا"Oʈ�F�;Ĭi�a�M(���"O���ŘqyLh�"+՛0���"ORDɕj�K*�d3wC�Ll �"O���.Z;�LI�emH��KD.�y�$��q�|���'�gU�A��Ą�yR@���{���"���ɟ	�yTjv	" )�R��F���yF	)R�	s ħTZ�!	]��y
� dȢPnD���J!��#3�<9"OD�P\ �ā(§��x=��҄"OvaYu�?[j �A蚙N5��"O�ٻ�M̮Gx���Y�	\��"O``���<���%cm$���"O�����+8Rt����>lo��9�"O��0�J�_�mq�/�KkFh��"O
U���"|?���bɶb��w"O ]���Di�m Ќ�P�±y"O
D"�C*�t��S���i��"Op5�4� uJ1��,÷&4�f"O��b�C�'XߢYj�閪/3$�@�"O�=���%���c�WT�D���"O�,k�bH6�qs&B΁�(�"O����K��.Z�����E�Y�:Q��"O����OH9�P4�`�+4�\�s�"O�-H��)=Q�K��?*g�u10"O�y���ߺ{w�p�3���5����w"OT�
��K�
��1�)@�ٙ1"Ofy�6 �(aCv��3x�L1"O���iL�lƤ� Æ�klA1�"O�]��@RWR����5;���"Oh�A$��)�<�s���
uqT"OĻ6�U#m)j����ܘXXHȩ�"O걩�eAbx`�5��Xu�eB�"O$��5�D5���a��@�%�h K"OD`�Z- ��I�v$�3e�xS"O68+��*$�,`A$�<?�4Pq�"O�%�G�9�*MM	Mۢ�3�"OԐ(�܍|��0��n^0.�
���"O�|����,R�E���єg�<�3"O0���V?T�PM��)"Is��X�"O6p@VA$Y0��2)�Rj���"OJ��Q�é?.I�)wNt�Q�"O��#��,�"�@�2O$���"O:q��0W��A��Ym�rd��"O�}9A����T��+��F���V"Oj�ѕ#t�6YxqA_(��|�&"O��ؓl�x�^��� �����"O x��ϋ�7�:�ص&àM�F�I�"O�ii���.3�z,���V�� ��U"O�q6$�0. X�W����`:r"O��Ag �4F㦉J�n%jQg"O����ϑK��0�7�8f2�qr"O���1  4@(L���6n�r"O�� �d�=+ѲmÐ�R?3����"O��[l��� g�!b�j� "O�QS�ŉW7T��tF��[R��h�"O���'D�+"�1v�<#L��[B"O��Hb�H�huz��E)H$\dHq"O�x�V�_�'��#"�U|:�3�"O���	51$�s��7wJ��1v"ORaӱ*�K]�!�	�2v�l�'"Ox	��K�8)�� �(Ͻ�<H�"O�98�Ra��Pqf�"W���
�"O�I��N��{�f�+e{ldj�"OU"��E�4z���+�lk�"O��ɰI���j���
^
6k�7�%D�|��7|��� �V'n����F)D��qaH��>�R�j�?=jJ�bU+)D�xsl��1�V��gG8_J@��D*D���a�;Sd�㖋��r�(t���%D�Hf�\�-���W�8:JI��h D�\����oj�5��JٻRBF�!3D�� \���h��E�X	ѷ�/(h��{c"OX���A%v^(���`�M��4"O���q��B��`P��O�%��ٚ�"O���2�L8N�|d��V,�ƅ�7"O�<����f�]�í�X�h���"O��[��0x�D�W�j��"O�Q�ÐF��B⍝B�T�S�"O8$A5�Z��D� w���T���A"O���bȑ=vî�3�L\���IS"O�x�rKO	\c�	R7n0jdP�"O�����e�	�6-<Z��$��"O���2���z%/,� HgB"�y����-Tv�8����D�*� �y�L��H�Pm�9cZ�2o���y���5(��Ug¥0蝲g�6�y�ܦ��@y� [�r���W��y��B>$�t��#a\�DN,
f�(�y2�˸H�,��� ߺ}朽ł��y2��>hA���RB��c@L!1!��y�.��S5�}A������jG�-�y"��{��p��S�*}�̔��yb�׏�Zmb2n�5aK8ԩV����ybkO�>rK��G�N���hűnW̄ȓ���g�K;'�^%qXX@��"D� ��-��V�N1�R� zT ��F>D�4����^D ���_oV��`oR#;n�����M2Ϟ��b�hx�4*�AG�6DbU��ʅ/5��� UF#D����+� tl�vbB76H�(�F6D�T���Ɔ�Ը�U/$D�lhG�?D��!�艁k#�e�4 Ųw0;�F9D�|)���	v����V3��Ebg�*D�hPm�Ns`a�5+��b��{RE>D���[y�{����2)�UWO:D�H�E���@��ɢ��C�Jnɢ7�5D����Ǆl���P�OBT�PqPL.D��k�(E�e�e��!T&�F�P��-D��y�iZ;����$��z����ӧ+D��a��U4h�{��A*n@�Sm'D�I�bN�T�< "B�:��A&D�,x�j��]hؠ�]#K�]0��7D�yE�Όb@��D�(��0D�px�� Z�<��d�Ox�(2'/D��C5�Z�;BV�A��I%]ν �D:D�Hc�N�b�ȸA���,ƑY�$D�\�5A��nd"��(��y�#e"D�Q�w#~���.�7Q@ف��!D���.�2��"cO�0����<D���!�?77H��@$]8��%�:D��@w3�:;���=F*ఢ $D�������a��)�B����'D��X�4�\z��#o1a��I2D�\���.��!����ek2@b>D�LI�D
`<lQ�c�,�J�(��<D�h�1Ə,�8�طf	>��J` %D�|��˨@�j:Ae���p��%D�v��u@cdN�P91f��$* 0B�	#0iy��/K'p0	�j�	L6&B�I"0����f��Wm��H���C�I�v8�
W��.� ]1F)w��C�	�M|h�7��0f��H�u� �nPTB�	+��$kG-�ia�*�M�7BB�I3%��A&dN���ʳ�_.0�\C�	<L�`��Q^K��y�i]�[WC䉣`0q���7#���Y%��2��B�)� ��x�Ʉ5m�xm dj��Z"O��ؤ�Kkt��W#�&<K��;p"Oh�J�	�A��3�C^�/"ly"O} u��:Ů	Dl�+%*L�1�"OҔZ������k �^�#PXX'"O\x�e��-~I< 0퓜d\���"O�8@�DK
���LN!?�b��7"O�ȕ(WIΑ�Q���"����"O��񬓑�H�v���}���"O詪 F)�L��D��n|.���"Ol�� ؈{��z%�C�V��6"O��[��(6@�:����!}��!"O�;0J+S:�k�.��RH� � "O��R`"��Ⱥ�
@F�s�"O
5z�׻i�0횳NZ*�赠�"O � �- 4��s��9�J8k�"O���.[�Q X�:3%�{c(�H�"O�58d��*�R%�"�	Q���sE"O�$2Q�Y�(�X��`͢UYx�"OZ��r��`v4x�NSD��ze"O���r7(M �#7�L�}	�)��"O,�Ie�-�F�j���s�E"O2��#JÞ#��H�6	C�Mˁ"OD�!�&؎~�zݩ��߃7E�jf"O�$0�K<K���j"�i�V�
!"OZ#d�;Q>0hS��*�2�� "O|��)��z��`G� �$�;�"O�d�С[)�^�� )�<C"O�c�0��w�>P����"O���$��	%"�q��ߴ���"O��x��Eªy���g� IY�"Ov���MX�v����Q ��<p"On�+q��F�&��0�Ag�8�8u"O��x��Ԑ{�d��v�9"O��sgR��ݹ��gr0ԸW"Oll����^���8�#��g���"OB�1-����kS�^�^ �"O40`�.s�.1�de�=
�A�"Oh�a'
�a���a�$\��"O�u �'��@R�eBǆ� �^x"O����
��X\s&��~~��3"O�,r�R�%�MA3�3/y�ԱV"OH�9.].6f�F�M(99���"O��AV�]�;�u��+0���"Ot�F���Ub@u�.	%C�Sw"O\i���-'�h���Cy?�
�"O|��@#�x,)�QM�)2"Of�ᅠB0j�"�)I�IA�"O�D[F��'p:���A���P�"O���p��;] ��� ��F0����"O�ԩAI�-U��5��·@��p��"O�}3�O�-�r}���R5���u"O��M� 4vF}� 3sn�q�"O��S���*�|�FdGQZ00"O.i�@��A��x�a>)E�9��"O�q�0���.�D��uoF_?��y�"O
@�$샨L�L��6Y+tF"O�U2���mҨ�Z���-#tL c"O��K" Du���FH�1���&"O���� C X�����.p�9�"O�0�Gܫ� ����5S����"O ��e_8��תS+Q��w"Ol@A� /2, �n�'1��M3�7D�d"A�����A���9g���D�4D�� 2� �)��00Q�Ŕ�`(��"Ol��e RW�1���jd*"O��S��U$�T�R
�xs�a�Q"O6M@Ҏ�+�� q�NQ��D"O��ҋ��D��6nS:e6����"O ���9��s��Yh3HQ�a"O�|Y����>���
(d+jT�3"OH�F�ȇ6d�1a�~#ܙQ�"Oz ��ɨh���1���7��Dp "O<[FF�)�|}T��#I�����"OʵRb�לK$��!@�Ĥc'�5p�"O��֊�t���0���.\� ,;"OJ�%��_�~`�hW�f��"O" �'HB<g�0Y��	a:X��"O��`"Z diɲ�B�s[^�R�"OP�ssCP
i��yq�%�@I Lȶ"OPU ���G��0�dM�R����"O`��w��R��B�U�h��0"O�t��*Hl�x��+^!}OйВ"OB�Pҏ�� at��엂3���"O�УsDڐ5�0����	*f0�O����N���Ճ{gู�����!���^`�𠫇L�U���}�!���C�J���.�8@�\R��ЎY�!�$�8#�jI�֏@���!��<H�!�d8H(���e��[ՆH���^�9'!�$��#����f�7�� 3�@�,�!��L 3I�P�T�O�OF* ���_��!�D�3j���wm�5 5����G�s�!��M�F{�%����9NfI;v��%F!�D�� ���õ��2(1�Ń��P"7�!�$E�L��ْ��T~�a�
�*�!�G�<h��SB��Z�hq���G�!��R)�T��-�:S�|	y@�:�!�d�T(|���Y�*i�'�Ϳ^�!�@47h�驦�T!\�
Q��ԙ+!�dg� ��ퟛA���3NIE!��!&� �)��B�y�\��@k�w�!�d�<S���@�A��l˪�.�20J3"O���	�P�]y�D$��	�"O${5L�\��)d셕c��1P"O~"��^�1���9��a�Da�"Ov����Gd�$���D�8����"O��8U��t���;ր^�+д���"O*�b��Y�d\0pi2�|��"Od�x�A�%� }�WȆ'K��	"O
aB���tm,�J�%)7M ��!"O�8�#,Y�*z�2&�,6���"O �P �h�vl����� �F"O�d[�.���e�4ԑ=�BIC"O���ˮ%��<H� R=A���0�"O֔����E���+&��5;m2��"O�A���Kso��RG�->�,qps"O�x��jA=w7�!��#.�j�b�"OBlP����d�ݺ�nR�|NH��"O0,IQ��^�<�C�	O��,�"O�UJC$@/a.�mc��ѣ{h��"O��p�ڵq�nLف�S�_��:�"O^ ��}�^�K�b![���"O`��D+�D�&t[� �)2��i1�"O�Ű�H[�^ڴ`��Ӯt0���t"O�TR��͘rI^(R]a7"OB�W�ߠ,��y�)��i�"OeT��g���h$H��a��"O� �P���.=@ ,��_D����"O�Y�2Lõ5>�y�p�O�`��UZ"OZ��`E0F7M[��X�C�$պ*O�=!��ϢAL�#cAƪd��l`�'=�s#�_�l߸��i�L�J!�'��  �O,b����]�I���'�4@��G9@tL���&��0��'yr���O��ȄBc�A�!oR���'*~<A��V� Ύ���M��!�'�!j��!���J4�P��'�]�eiQ(H������H�|�)�'"��"f9;�<��G��>x-z��'xr����\�g��g���oh�P3	�'�5)�N�#�E{Q�CV��D	�'�du3Ez.\�Q@��F�,L��'{ (V�ffi��i
<p��'t pSN�.u�:�iQ��/!21"�'2 ��]�0����$>���'9��"�˗L��8����	g�����'���H�����+�.�7N���'��}#&@�_1�%��C�4AU���'���j ��J�RY36�G4=�h�'P)�G��-R����e��J@]s�':�(��LT�th��� $u����'7污Di�[&0Rr�]�:1�m��'��Y*��7*L1���#1�,���'u`$��z����)�1����'��`��Á;F	L8y���s"J��
�'Ū����x�����.@�Y8���'�2P�
�$`�ܴ�/ֻW?��`�'� Y9C�
���*4n�K�:��'��+D�
-]Y@���"=zv|��'��{S�͸e���)큁F�!��'%� ��?���j��	5D护��'�ޜ���D+׀Xb�H9*����
�'�0\*#�
�rOf�����53.��'�����̉���+c�DaH(ph�'Ѣ �G� cɦ��É�7���'��+ G�0�ޱ2S�Չy��AY�'Y"}Df] Q���{bΒ�j@�8�'G �"�H�+�U�1�Y>y�(Ũ	�'�V�8M��Y� "&5al�8�'mTqq�]�D��pV/`��L��'���pcF�90A��\��yA�'�"y*4���mh���SM)Ðq��'sp<Ȧ��T���b&GJ#ɸ���'6f���`P3n�¡� �ѕپ=B	�'Q$9T`��͈��s�m��'�H�h��.Cv"DX� �0a����'HJ�w*Ͷu��j�J(}+<	�';B-[P���1�*K(�*([�'Z�i�H�܄���I�s���'V��:��{B�<"G�7g�*`��'t5�����͎թ�O��\Q����'i,�rD������A\��,p�'WL�1�O��9�����#[{��{�'��1���0�b)a�ٹD'�h�	�'G��`�
;\���"4h�5@E��'1�uY�G�3Ach�cn�%+��@;�'~��8���4�}����L���`
�'C�M���~�������2K����'X������(b|��!�I�Js�'�V9링3)<���4�ȿ3�R��'���p/?`5*��Í��+@��+��� �080��2#���x��?:N-0b"O��
���&{��(���˩"����"O�����Ƅm��"%W�pc"O�]�qI)V9@Ļ��U�����"OT��`aB�sI��@D �%��(�"O� G�6� ȁQc��YЀ�a�"O�����2~�<��GѩE���J�"OF5�421
��1	�Z��؛�"O �B�%�JA�r͙6v���R"OB�R�ʤ9�0@b������}3�"OTyr�#@�����e�B��"O�,�4F�-��Cu.�8{�p}Y�"Odp%�R=��m޿}W��"O�̂.�9S�:0:%Z�Z@���2"Ol�E��,*�P�k�&��"O��r���3��|AG��Ao��#�"Om�n��������(dJ	�a"Oܰ�dJ_!>�S�JR�:�"On5+a�&qEiI$��# �����"Oh��q�ٵ,'*��� .Q�č��"O���@�,R�P1'@��}�0��"O~�h�,B��0(�ŅP�	��9"O~\`�	�3.APJ20����"O�����>Е�fķM���+�"O�iy�N}�H�5⃶c�&5˲"O|!��f�fi�%� $դi 0"O���pe��o�rI�u�U=wL�"O�ct#�r�XX�BX�+�R�)"Ov��Q`��'7>$a��A8Y��Q�"O.�N�C��d�qoXl�V��"O
59�bNJ�`e�G@�_�t���"OV��L�,1��A��4��L�"O�$	K�\s�cD��-w谙�"O�	�m��-D�i` �tmN9�"OT�	�F̱v�XtB��; AW"O��֌A#O�ʅ+�(�+`x�"O"����p��|��!Qb�}�"OV�(���XXD�.�V �"OB!��o=���(U�{�8�`"O���-�6˂�SwMW�[�J(��"Ot��r�Y�u�6�ر@z��G"O�ī���T��2��17f�@h�"O0`#�S�3���ڧ�W�[R~izr"Oxs��Z�<U����]��sw"On���(�%M�IP���wR�"O̙�¬ѽT:� "ʎ�!��{�"OXıU/� ��p�r���{
p`e"O�����Q�S�rpr��#��"O^�!QGU�6c(�#"�����:r"O��zaE\�Є�`���8ό!�"OvD��<e��5
"�d��	V"O2��'�*k��y��Gۺy�|�1"O�����s�prRF�
c���:!*OҁɁO�k�(̪wm"L�\��'�6�3�NɻR�0(�c�KY6�j�'��l���0@�x��;��z�'�
	���C��I��:�(
�'n�A���NI��Lƥkb��	�'ؠ��B�8���F!.�`�A	�';t�Ҧ�P�
�Iy�JҹV<�,b	�'����S��6�p��c_�I=�1Q	�'0�Y�U	1 �񗥊T�<a��'��H���4��})w��P	�y��'c���[��\Lᶋ�t~����� $�i%��)l(�{Fb�&��A�"O\��C&�2����L�A�Ł�"OTp�bO�y��]��I�/kU�Q"O`���^A!�4�ՠ2��E�"O���E&�9h�@�g�g�P �"Oܐ(AC�Wh:�RU�Q;?\,A�"O���!iF�q�~����'Q��˖"OFqpF�7dH
}���::/$�"O� ���25�̓6툉8���"O�  �j��m��ۃF���	�"O��R��7'�ɋ#K��W�0y�4"O$������O��\g�:*\�;�"O��CH�#r�1���8b����"O�Xx��I U��`�j�VK�<�$"O�H�נ	xc�iPi�
*D<]�D�d���<�2��*�hu�2�Ԟp������[�<)��:x�|zm#0I��(3�]���x�K�	hgDM�r�L�,!Roޘ�y��ǂ)>"���Ϛ+m��)��R��y2�S|,�-��ca4xt	v�y@� R���T(��O!DA��C�y���$?:��!&\E���ٖ	\>�yrE�11���N�D`�y F	"�y�BQ�S��9�.A::=�Id�ߣ�yr#ӏt�L�yP�I�8� t���)�PxR�iC(j4�j<S&g�3���r�'�8�;�lB
m����u*H!h\Q���HO��#j�		�N4�w���z)ܡ�s"O�hS!,��U)Y���!?kJ�A�"O�5Y�ċ�.d������4�( "O`��%qT�ɒ�p|b�	�"O�=��S�"1�%!���t�4h�&"O��iŒ2���Ս˭/a$H�t"O� �w���`�P���}�Ԍ3"O�E�GM�!�P�9�@æt���g"O�b B;y���bg��xj�-YT"O$�3B$tbրX�b�2�"Oڔ�ԈD7z�t����BO ��r"O|<�ŗ�,(l�q�iζI
�s"Ov���ץ0�hd���@�0^�W"Ol-�$�Á,t�#����>�S"OJʑbVt/� j��ݫG�b��"O���@��
K�Y�2��@��y�"OB��#�ʛ0�"H槂l����"O�-:`GQ�s|��˳��j%,iK�"O޼A"K��ha�S�C�F�"O��P�bԿC������z@�#G"O���Õ���!�գ;?.��"O����܏x�Lٙ�ǉ�SXx11"O���v�̜jdI�QS�=�.���"O$1��
:_T � S�;�"O4���׏}�$���kY�D�&"O,�ᄎ�p�F�h��5R����"OE��-$2��0��`� $��"O<��C�\�Z41rLSP�>Q�`"O2���ȵc���P3��5����V"O���'I���Z��\~���"O��6ǀ�Ls�����al��`"O�Xc7
V�j]�L#pB�3\�1Y2"OD��dgJ�I�Ľ�UJ�0/�p�V"O깰+^&<똅B�+�:�)��']�Xʓ���u����g6*�	H
�'\D)��O �o�� �m�S��
�'�A���d�6�z#hF�Lu���� �U�!�Y�O[t���ڕiq�8
"O$�Q F �fw�9H�Ɩ^j@@�U"O�� �@z�FmR1��lV6p�"O��a_�s�2���N�%T0I��"O\�S&A�2��r�>)��"O���aާ=�Ƭ���/|P1�"Od0��/ :EAH\: IZc��B"O�)�$�7F�г��B2B"O
���k�8*��e�Ӫ2���"OV �*�"�
%:���t"O����Û]��Ze%?�z4:$"O���P��e�PT�E�K�o���R�"O���mL�Lp	�R�h)+�"Oy 7�R=4��PÒ��*����"O��؄Q�I�jDcM�t�X� p"OTQ'P@&E���@2HnyF"O�y�Y�sr�jLV�FUh�c"O��i��X2\��=�� ^����y2�_�3�8H+��"~vR����ɣ�y2#�kRHR���,``�%2 %I'�ybN�S��c�,תW�d�Q��P!�y�*%#�`����P��q�K̥�yhR�m8v�;F F�I������y�f[�pI����C�:�FS!C[��y" I�}4z�Q&��,�B1O\�y�(Z�N�������)$j��yrꌽH�5�P�
zV5aD�?�y�'
�y�bQ#��H9tB��B����y���<�*��U�*�0�#�V�y"�W�L�A(�#��$k}����y2�P-LГ2�G�P+���b���yb��-�N�1w�_�B������y��S�:�4��e�#5 �0AT@���y�[ڜ䒠Á�0x�����u�͘�|$Hn�}��9O������"��R�L##���-��R���b�D�0
4bш��w�
Y����'eJ2S�ݣW��6"�pd9W���MS�L��k�&=SC�����ɇ�^��H���Ƣ���*�P���c��&5��F�i�BQh��?��i�R�sӒ��"����h�$��1XC�9H��O���9|OX7X)�����i�����ae��dZQ�P�ߴ�?�M>��'�M�] ^9��A�
�6��A��O�ɀig<X�۴�<Y�[%4F�WXbo>�e�Ջ~Eb����Û@��}! �	uC�iY�O5�DxBk��B�fX�M@�L+��&eھh 7M˚5^<��j���~���Ȁ��{̓ ���	ھw��[U`�B����'��s��?�$�x��'V�X��9���p�Dpz*��gA�Y��K���G{��ɍ�:���'!T����i��^���S�4LZ�f�|�O%��[�Ȫ�˽>>�D���T˓9`D�XP��Y]�>�����\86�ׇi��3E
 Y�%�RiG�_��h�3��)%'fh �b��������9f��ARE"K�7Ȁ�/��G��3m\�Y�4D�����-K��&鉜	m"�D�4DTte{����*�z5��V�3y�GŐ��1��my�'��O���pӔ���,�6��6B��jNt�KbLYϟ���	xب�`w��]�x-i�Mڊ>��I�M�v�i�I^��X �4�?�����!��P4h]�q����DM����ȟ��	����VB��F0.Y)�Q�D����-ѓs#�)���9H�N� [���`H��L�a��Ph��F�C�R��u�0Y�1 ��KT�{�#�V�(K�@��HO�w�'r�~Ӹ���~���&���Va�>$��Y��+\zp���O��2b� ff�8FZ� I�����A���OzN6n:#�<w��S���<7R����VP?��D�\כF�'m�i>���T��"0a�aE��Od�� 7m�n[p,*A$ڦ�1O��3�r�1��F�M���}���ߝ�6b�O5�|8�9V,�� &f��D�/�.��!�#e�f~�@���I3�j��~��)�=+��J*i?��e��)�p�mZ�f"��O`H��Z��i��ɆC\�/���Q4�İ~6�!����O���+�$>�u`M;&]�SB<��S��?"���Gy��gӀ8n�]���u���K�`��|^f�S���=�~b�'QLT"CA
�_���'�'���]�xoZ�o6���&Aҧ>�J�����<mf�M؅E�&_>&�k��Z�"��Ū�Y���?�S�? ̸I)!r�bT���O�D����  �<ZFn�&n�� y��	o��S+b^��r�B�D/Pp��vAX��vt��	�f�T���j���I�M���~�'h�_��{���<b�d�5y�PF"\���O^"=�g��/��RViT�.Ɔ�������Emڱ�M��ƛ��'_���'��'�5E_�` |  �   8   Ĵ���	��Z�tI�*�� 3��H��R�
O�ظ2�>���& �H�O�QS�� y��]1��S�x%�D+QlW���K�4;B�^�?�vR���'�V7O�`����4y��Y�t�B.3	*���ņ�S�B���4A�qO����D���M�`��DO�꧇�=rF8��ʋ^y�?l��pS��(��$֊wo(Q�&č5o��I�	*��e�Sg|� 4l����	��'�'Y����O�牚!̀��t萧��ʓ%ӎ9��J]�f.v�h�џl���O	��07��hy�E�{)"�ҵ)u~2�ݠ0�T ��ݺ��
��rE���NHb2`SQ�j� H��(��|�(���5A��<�`ԑ��Q��y�.Zu�'�ֹDx�U�Y��''7�̀�f�W�+ђ"<�q�%�!2P�o������?�����ݶlD�x�O��Ӊ��ْ��'e^����$M��(B�Ӝ`D Rݴ��#<�Ҁ'�MP��h�)@=H�h��U�}�iɥk�\�;Z�"<yc�4?��.Pᢁ���_=�x��aSoy�JT�'.>��?9�KL%�����>������)L�:#<ɂ�(�|Y�����+����∕g �����?�1O��r��$���w�|0����]�v量[E�'ƐMEx���M�'A)²
�A��m��/�sUÏ��W]�'|�i�;c���ˆƳ}�{�JJ#.�qOp������I�8���F	x��Hf�ݿB��JJ#<yP�6�V ��l� &I�4	5$�Rq�ȓ	Ĵ   @�?��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �T   �
  ~    �   �(  �1  �8  �>  BE  �K  �Q  X  s^  �d  �j  <q  ~w  �}  }�  C�   `� u�	����Zv)C�'ll\�0"Ez+�'J�DlӤ�;�5O���'�hA$cŨOo��b.@�`u� p�v.Đ1eʉ%��Hj���%��¯lݱ��.��?����?�YA�)Qf�)��gU"%�E��:2�⁃tC�*N����*�M��ү �u��Ⱥ+����'�6�p�a�+f��i��eX.~�Q�`Йn�J剒��Oz���
u��`�Aަ�*�$�ݟ��͟p�����Q��S2 �\�#�Kľd[��	��M��f�����O��⟀���O,����3Bv4@�B��r..X{�/�O��d�O^�d�OD���O�"��i�X�����ѿR�}����9������Z�'=��mګ@��ɱDU�=�ll�D��J��O2�	g�=�xlyV�5��3��@j�"J�N\�%2c
@�O2�'8B�'�"�'�R�'E�SӼV��7�$IriO5�}kNߟ�����M�7�'~�f�'��6�ia�G�ئU�ڴ�?Y�!�`v��c���r|�k�+�hO2d@��	Y�\a���c��Z��]	0#�a��u���j���U�� k&6͊��eq۴�*�����7���bZsտ9����؀.�^m[֣�aèU.na�!��
�%v?x�x���{�X�#�f��M{3�iM 7H�#�����&/��!�g�Y�"���R�_�"^��q����գ�4V$�v�/�b,Y�L������H�;)ϒ����q�J���!G�/q���f,�Ft��`ӫT��M��iɺ7*4��%	E���8��$˛j��ѰՇ����'²8��x;���ΦQ�V����$��R#�2t��ǟ�?A aŲ}J=��.�	%n�����?%D(�Q�#�6Gd�h���6����ɑ�b5���d�$p��S0�C��,��P�t����<1���?��"��� i��t` ��&�<n���PHM�р<����G%!�Q��Y�';R]�S�����Ф!4r��Ďا hZ���(f�f<;W�	�@�r X`�'�����?A�O�h����>���h%˘�f���a��'���'��OQ>}����zni��H�k#p�E:�OZ��I@��*5�L�6�h�A��yC�$9�	$G�"|z�w��]�-�(X	05FE&�1�
�'|vd�����$PCDkD��
�'
d�PA�+�0� 
R�8P�ِ	�'ZM�CF�� %ۻ~Tjh;	�'w��Ӏ�*|�k�f׸v�4� 	�'YpQ�s�6�Q�&�U��,<���@H��Fx���O��Fy�֦�f���5À�:$B�I:	$$�S�N(����h#BB�5L���"V�5�X$����a�lC�ɺ<:}�[n8X &�R=��B�	.P��f̋n2T+��	V��C�:J4�Q2)�1c.���i�+�p�S9rD��I�����˧C��I�g��'�C䉆,�M����>����#]+��B�I�+��T/)Rr� �E1R�B�ɭd��h@�;��!�O�O��C�Ɇ8����g$r�Tkɺ#̎���m{�l�R~���ߒYqD'i|)5O2�?�)O����OX��&T��� ��Ń�uڃL��fF�P�AU�c���Fb�,�"����Q�1��Yu�e��01E�Q5o��-����X�ن!8$�]�'cZ"<.,R'�N�_8�<"�剣o����OV���O�HJ���3s��"�E٨]H�j�H�<�����(�N52�-�J�]t��|��:��'���D �L��I�#L@#z]��� ,��	e2]�5\�unZX�W���'� II��%l��+���~�HTk��'���"6z�KH=`I��Hvn%.@e*�ၣ��S+(��0�&�3C��,QgV�(,�F�̕8w���q�����5_Hx&�rN�Oyx�e�O����1i	�(j,��O�=YS�'Ob��D��=>���B�-�J�*h��\Bt�'���'�l=��H 7hܐlBfC�.s��Í�D�\�O�h���*f��L{E%�Mv�1�$�i�X�(٠{>I���<��Vy��5hqJ����� ��LR$�)}���aY3|12Q����5bL5���	�, ���'�P��� ��u{uf<b�6��rmE&)�(��-f$L�WH�	��O$�
���T?�,Ӎ,^���P�ò3�E�+_ҟ��'d�}�����?9���?١��"`�1牞_ȴ��SC�5�y��&f��9�!	��B�|�Ӄ�X���dY[���D�'L�I� WYбa��V�d{f�A�&�(Uct���M��e8p�1@A�*S���'��776^�f�Dt<	���c�N8�bmC�]e�ғC[7P�Ȇ�`�N(����[W,�$�sXbQS���ӟL���:�٪��Q�E�
e 1Jڳ[����(����V	^�K�VZ���Q�5�$�ަ'�8{��b�<�'��$)#ǖ�<s�b�a�1Y[�taÓ�z-8��=�BI���;@v� ��C ˟(�:��#/�W�V�jP	'�"9c��D����Yja��d��$kaH?-�����R2����0.�J��U��Ԧ:�������ng��o��`X�	�WYx�,�~�`�7�Eß�������ayʟZb���dj��}�&��G��%������ �O�a��B����Da�	m輨��ʒh�<���<���T+_�V��O>�	 fy@�@��ҿ;�J��qJ�a8�V�]9䁞����z�*�$)6��4��NR��O܆����]�`��v6��HUɉ���d�%^�hӍ
H[f����ܣA�zij�&�%���7r���ь'wxY�A��4K#�O1�D�ɳ�MĽi�����O���u.�SB	�Ē8�n��W���	֟��	�XS�5*2�����H��?� 퓙O\�U�s��M�1☜��Py#�i�2^�0K��b��G|bJH�Hq�'ȜsD��&\�H̋�A�Q�18R��y!��b��B	�XN.%�����^��`P�R�\��C��&}�Xݡ���nR�e�)�ģ\6�mj���L����/���C��/$��9S1"7�S�)�	^5H\�I�?���|������j}`��ԥa���ic�M�%�V��ᒄbLW9��=�H��`�'�#=)��iN�V��y�)Xe0bJ�<M$Hc�[��@�
�� ӟ�I͟��I��u�'HR5���&�Һ���kX�f�^1�!�n`�`x���{�eC%j[)fay�'٣����ǘ4,�`U�)��֎d)��R�m��[�����$�*-0�����WJ�X��N�, �ae�'{��'��O\"|�����&8��ſ\��Q	'&o�<�SiB����ہ�I?ve�))�c�t򉀉M[���$�	.< HlP���+0Ѫ�9ՃՁ/ܜ=������?�+O����O�瓠�%aD�D/T):�	!DҀd�Hk��V� �j�X��_�]�e'ڭ���j�I���Y�+?il��f��5'�.=ؐ�'Yd�Q#��a�U�*ۃ?���6�ɼos��$�O&Po���"A�G���aFa��(>�ם�Z��ߟ �?ͧ��'���)R�L��s'���d¢X)�}��VK�S%� �,@��֨g&�9G��6��<bǑ$2`�f�''�	{��'&@̈�c� B�z����2Me�XS��'Y˝�&�K�,fϞT��a�{װy�3	�)���W �5�vM:j�A�6�ثD��� ������G�<պ��)6�<,�A	��.�OD�=@u�У	��8��ډl�d���O੡�'�b�h�T�$!��u>)�s/θ'˘}�׮�tLj�h3-7�$�O\�=a�O��#��U�-~��4.�?�&y(#�	��M��i�1�|��Q�(CĈu`���g�	b��'�@}�c�4�Q���4LI�)>�cpcR�>�̠�.D����Cߴ�~ա�,�7�pʴ?D�Dنm�0p� \y��<eBJEQ�9D����L�b͒49��M�H$�5oq�<uf�e�R�JG]�f��y�b�n�<1�"�._Z��g���L"�.�iy��@��p>�v&�p�TYh�K�����g�<�J��P�<*3��\��ѱ���_�<i�!ڸC ��gg�Aw��T�	]�<��G�ji����/�&,���PO�<D�'<�f��/�$[frHyt�Nx���������2}�<�r�"KHh��H0D����σ�N0d�y�AZ�j���� 3D��+A��m�N�`�a ����6D�\sÕ(����ĥY�s9D�Ʀ3D��X %��E�v���Ĉ^%,a��1D�HP�LB�=�@Tke杤
!���a0�>��D��ő���e��Q&�JHu��y�m� �\���M�*HJdi���y2�ٙ��\
#�!=�(�S��y"` 0��A���ل~5ȹs��y�H�T:Z%�FD3 S\Mʢ'6�y����2�,`r#��c��P�e���?��#�Y������4.��?.�P �.���.�r�<D�|`���:��5Q��2�,��1�-D�L�F�P�3�lM��L��[N�� �*D����U -�d�H5��^�����J#D��5�T�p���Ҁ`˰+���@�!D� ��OF�n�$�"fʎ$�8x��΢<i�eGV8����E�C)���E�KE�$����>D�� ����
j�
!AB	+��{2"O  )�a9{�����:;�yQ0"O��y�?��Q�C-�=���"O�P��c]�7L͸r��(8� H ��'-����'7J��BNבj�pA��.�}1�'\�9����*���{ ��+^G�l��'�����i	�fh!��T1�m��'��L"p�ܥ��#�%��H%�a�'Z�ŧ�/��%CDќD�(��'��	 �Ǆ7KДS댷@�����D �Q?Y��
̈́P����ӥ�1)�6�:D������7K&\�Td�{�q�'�4D�@�� T�j ǌk���
0D��5jQ1O<��5):-�¥#�D;D�t��ˠ
�Np�
�5��)p!-D�P�E��,G@�T�	M�Q�|Ԁ�O�0���)�_?����T�@�T�bwl
�' DX���.�< `B�X�4��';� ��M(M�,�:��ȣ�nU�'ڴ@���(7��ұd�*���'��ؑ	͋|�u�t�v�t"	�'1�*@($�b��d� �,BAyb�U�p>�tH=�AH�=�^Y�ԏ�C�<)c�*Si:��Ћ��-P0���}�<�M�Z)r��d	X��IR��	~�<� 
Z#`�mcS·��\�5�]c�<9�È��*("��aCP�i"N[`x�x�ա���*��9^w�i���G�B�T�e�+D��cD�'j�yq脎Y�t�VN*D����^�h� ,�F�H�.��xP,D�H�暘1x	�v�Q�fn<hU"+D�t�͐|1�� _״\A��(D�x�0A4�����.N�X�L��(ړ_!�1E�$ȗ)�`<Y�Y/�x�`.Z��yP-D=�qH�-S�1�g��y�Eh�:�#�1�L�P����y"`S p`���7 ��q�Z��A�?�yү��� T�ۧu�$%؆.��y�Z�@�2�� �"�!�ҫ�?��+�^����xx�U��^���G��J��-D�d�2)��6}��RB�J[����*D�Z1��)Q�.�J��N��ga��y�Hl��@��Ǉ*��4Cco��y��T��Z�:T��M0��O=�y���&6��r�ٗuкD� /��$����|����/hzћP�nq�p�$�yb"�#F����"�.��Q@���yGE�CNPE��+�@���Ŝ�y�ŽTY�OҘvҼ°[��y"LJ�-��a���'��$���\��>Iwj�o?��J��U��}9�d+r�]��B�\�<�C��#�h��X?BH��0���s�<�R�UY����y����t�f�<1��Z�\��aLU�Fw�}�p�f�<�v��[�H(�6���+ON�e�!�D���l�K^?L��H@�<Oў�*� �Nk}��"�0�,���G�L�Ʉȓ5�8�'�]�2��Z��ȓt�iRꐌA��50%΄9U������(�!��؈�F�s6�׽>N��M���9`�9͔$����tJ6�ȓjT����i��d����N�N|���ɣfx#<E�g
��00���3�V�"u!�D� ��)3dS�F�p� ΍2_�!�� B=+��+V����jG1q�Y:&"O��i�b	5!���t	ɼO1UIU"O�E)�&��o��8:��ɂXtd�"Ov��I�8�Ga� }	Z$W�d� �O��1@�ߕ��y
��;��؛�"Oh�'!D�3�@e�2Ň�p43e"Or�jS��W3p	�$O�^�<`��"O5�&	?	�Д���ȳ~]�q
E"O�m\/�2�[�tp�����'�hDA�'l������4cL��p1AybIZ�'ڔ�S�I�eQX�ˠ/�ug����'w(�ZD=Ir48 
R?t�]K�'��Q�m�+Q㪵(�I]�!N�-	�';$�3��9�̰Θ	E���'�0�֪اnR�)jQM�}��)����x�Q?)���WYL,�QF��7j�&$�g.D�0���V-���R���53��1D�Ĉ�nN 6H�5�Aᖗ#��!�3D�(�3 I4YIH�
�Ĉ�B^p Y��2D�t���j�N9���� <���<D�����Č(��!O$��(Ä�OB��)�'/#��v��@ȣD�,�$�r
�'qth�q`((F�U"#��3 i�i�	�'�X`�� V?&��yX���tt��'δh���[_�����[>@�x�'𤽠f���"���X3ਛ
�' �}�2IC�lj�S�kċYhp:)O�MRB�'�F�!�a��"B	�e�0��x�'Ot@aPjTY`f$��T���`�'�h��1ܼU��&��_RL��'/ <�V�Ĕk@�P�$ [�� S�'"Xz���,�����ěN	5r�1����p�>�Bǝ�e�&	��È$z9
Յȓ���y��(i�P�96 U���i��9���`b܈.�YWh�4oPՇ�J5>��
��������z0��ȓ)&ʜ��#ǖ,�H�]�]�܆�9��l�B�uHE��@ד|[6�D{R��¨�H�R!N�	\�$y6��MM�({�"O�p��~N���eÙg(8��t"O#a*��$����ꁹR�[�0�!� ;X$hRo*��� #��*l7!�� J�X���&VTt�B��`5!��3A�t�R�Ll��!�9R�k�8�O?QV��G�U�&�G�.Ƽ*c��I�<�UE�%l��S�R����]I�<�"G�&q�%�
=N�P��E�<1����/B�@���G;O@�]*'��C�<A�f�x��H�fD7M>��5���<�K�D�T�j��%��S0��yyBD�p>)���_vLE� ��t��<�HY&{�<�Ҁ�Q�\��%[�+�T�<a�U�j�ZոT��8ZK��b�T�<�@��<S>R�˵�^625{%�l�<A����I�QNO�����\|x�lBi��4�4�]ސm�'�?Z�.�(C�&D�,p!΋�`���R�wS P�	8D�\����8��٩t�.R��T�8D�xI����}[���#��B4l�K@C8D������6p�!�'.E��!D�8�����)�2Ę6̇��D�ɣ� ړ}���G�T��48"<�D�̋"6��![�y�95�z�y��L�n�DtKG���y�l\�y��A:Uh݋gu,��6����y
� j�0h́	Z}�n��F��"O2,����Ab������QB"O�Q[�
ס/*���6�۸)���D�'V�����S*p�0H�B�/�J5"�oQ�[��ф�	t�p��,��t�
��$�,y��,���#�	5�|Eۆf�B	��ȓf+J��a]�w(�"/�Y����Ĝ�Q�&ޯ�� ��L?D�`���Q��1!�;Lh�BkN�']65�'��Z�)$2t��Má<�8���c�0FȨ��R��ui&ӫT覵�h�)a��ȓW�J!T)KM'FT��Ό��t��ȓ:��E é\�@��%fȐ��zs��^/>��ŢN�����7l��I3MF��K���R_	$0Ĵ{�#7D����;�<���������5D�,��l"X�P�h�)�p��O9D�㲡߷K4l[�ߍx��9QS6D��Cu�_��!��\�f0�
��!D���a��m����Z�"b)ӵ/ ���E����|�d�2D�fBhx�d �yR'��]F-i�N�.b��l�&�y+��i�t�oY$Ҵ�1�C�y��Gxp|K	ȉp��D:D!�:�y�nÕ#vz���T5��8��'Ş�y"��2se�)���E�(ڰ�@����?ɠIFM��������G�[ȪuՅ��s�|�&�)D�`b�%��S�.yz�ę�)Fv��w&D���Nd4�Blͭ3����ҁ"D�����>M�!�Ԣ����k!!D��ѐ��t���e���~КW);D��ѓ�W&��%�"\�_&^8��7��$>�Y������a�B��BH�r�xd�rg��˓�?����?�>g�� �X9,8|xh��B�}�N���_�N�R����6.�	�$�G	\'$EyB'�yϊ%�u�Ԥe~��W��m'������(t��M)}F���֥1`�`�Dy"k�?q��O��Ls�
[�0�И� ΁�S�d��(O��$"�O@]Y&��_�b 6�>���'�ʓO�"-G&J��$ؗ��Z�dI�'v`����'?RP���O/B�'�pɛd��uT����ϋ�*��;��'V�q��C֤o�p��D��C2��#�edEZ��4�̓e7�Ih E�v|�1��K��yr�2�D�!\�:Զ�AōT7&�x�Haܧ6NE�%��&m�T��;o��Γ[����������'����i�R��V�U�,�9�+L�!�ItL�q�đ
}φ}��o�,tў,Z���Ρ[{D��E@��x� <�C�>�����O:��q6Pl�OV�D�O��d_�����]��Q����0�c�h�7N֖�e ��M	�EĬ2���k�)����?ᨥ@�	Аin، u�;m�M,3� Mॡ e�����b7Fx"g:wxn���Y�w���Ŝ���������F{�:O�QB� �o ��j��3�@c"Oh��!˝k���[�/Q�L�̝:`�'�L#=�'�?y-O���3�C	�0��2K�-V}� �M4	{��c��^�QL@���O��$�����O��S�>p)���� �j&&U�8���qS���e�P�	3D�7ְ=�D�V��4�6��|��Y �%�'q���hD�_3Fź���E?���ቢ[0.�d��j���N=8r��Ŋ���,�$0ړÈO�� ���y-��#t�O-pH�+�"OB�# MT>�����MW�080R�x�۴�?q.O:��D��ܦ́�(
��p�'h���B�څ|F�d J,G!���	+Y���ݟD��@�p��q��O?�`�&�wO��'8��+�@
f��$�u�Z:yx�E|�U��ș�j�	>�V�#5��{��"��Hy�"#N�	~�
$�W�'^\�	�l�|rqi9Qέ#e	"'g hJ�CKy��'���2�'\�h&RUC��B	����=��I��B���_� �a�O�X^� �@������H�5��ꙡN" 9���ȇȓc|���
I;��� ׍�6Cn��ȓz����M�$��)H�nЈ�����S�? r��G�8c�q1�aO�6�5H3"O�Q�����5:�W�,��m��"OZd��-��~����� 7@=�dJ��O��}�@׼̘`�C�X�$E)V�^�~̅ȓS�dL���*u����A[sh�� *�QB���&�
ő�N�$Y���dٌ�CVɗ�\5�𡑮��c�"=�ȓq,ja
�g�i�,s@^�1 "�ȓNE��Vm�>40g����"��	 *���dE�ED���e��h�������z�!�$7b�xq�V�ۜ>˚��c4@!�$D�,�����W�n�(xҵO�g4!�P?�t�����!�N�����k!���w�����'٢$�z\��O֯(�џ�A��Mˌ�d�������n�H��չ�W��O�(�u�өe�lj�p&��r��&�4">G��L�OA�ɒ0L����#3$7w��K���5Y����2Ȑ���4UХ�v��
c�C�	�:HI{�u�h]x���_��� wyҎДT���B$�#/r��`"]0��$�O��D#��?A�'������?b�`4��Kہy��1�Ó�hOv��D��?3atd�G Kcպ}���Z7/�'걟������ѱ���ME#������'ˈE�J���<iW��6� `S�!P�P���[FJ��e��T��O���Oxq�p�>9��tf���|�U� -WS%�5ȒLc&��O�x��h��.R"䠀��v�Tq�#��4E�(�*�>�f�>����M��Zm�d��'Ř�E&�!P
X��.�?Y"��S��]��?=��[�IE�y�ǡ��sE��I�/F�H�TD&}J"}�-^���M+�HP�-d�}�EN�G�ТIdyR�W����3�ȟ*%��WI���j���_��4��I?�tĕ\�T>�I.Y|�<��q��*Y��Х��-FcT���!}���1��D��H��uR���	*� +bh��H�KD�'��0�@bm��9O�ڇ�O��c��$�)�&�%�T�C�'�0T��� H���B��H�Xy���%2ظB�I"� �!��X�W`�i�bȝ�}�6-�OؓO(���D�|n:z���闌ȗܦ����Y�:��hO��<q�i��n�VX��_��As�{�	~���O���Ӂ�30�	�UΏg)FIh�'�x�2� D�D���ʓO���A�'���[��b����]����!��}�<�çηZܔ�`*\_�~t�e�{�<!@c�>,�AC��UG� k&N�w�<Y@nڍ>�\��e.ËG��rR�Cq�<�lB�ڤ������SDn�<��JS�@uJd��k��n���#Sn�_�<i�Ț Wl��e�=I2|��l�Y�<	f�R{>�R�\
[�s�Q|�'�l�S�'UE:$:�VOܕk@M�*#$����>�����:D����()J��>9
ʄ��)��*�Y�,���4���q����ڨ�3l��=���x靂~�z)�4#��3�I:cJH���y��-�9wGj�ڰj��	�ld��Bˊɓ�%���V  �)�e��q�c&�z�"h�� Z�����
6r*E����Y�|�o��W�tс�`]L����e��Ԧ-�s���ܸ��/�$i�� ����?������e�*g��	� b!�.6]>��Oꬠk!��=6�rIXR��*`��N<	���	8��!�o��FC�܋T�S� �!H�L
i�(]zt��4w�RO�]���'�R�զE"�$O P���ݰ@%�UQC'T��x�"M��HG`��&%��V��p<���'^S&D��OW7�6�@2�Y׸��%�i���'R�O$�����'L��'���<��0�
�4+BЅ ^�3�����&��'�j�a�ߦ�2W�!.yb>O�{RU 9���;�$H1]�Dj��J�5�@�F�@1��N^�Db?O�ɔ�^���*��F�m�8 zW�Zȟ��'��q��|"����'g�p���n��Q�TgUp��'Ir9�1d�?Dv�!b��R_` J�T���4�*�$�>��@f����M��O�6���jT��h�H^��' B�'�ם����	�|z ��r���$%���qj*q��x����:	�S��S�/�T9��\A� f������&�L��1A�.L�	�5/H#=d:�XQ익-}�M��'}�4s!�I�2���gF����4���Z��?	���?�"��^����R�_�FFdx�b#S�!�$�1}z�4��숕w�d�+�T1qO:�oџ|�'��-��'O�ihJ���T_�5���
�23�f�Oj�DJˀ���O��k��@����9�h������Y���)���`3,�q�mP���#�,��Q��+�ja��4��a׮߆�,��i��7P��*�H+� ��󧅫I�d@��$�D��a�۴�M+�� ,ҍr�ގ2O��ĭБb<B�'�'��)�J<Y2C,��,��L��]z�-J(<�u��/yn�e�QE�=z������/_������$UF�xQoZ���	i�䩊�_����<=1��_�0���"ȭi����O ň6��O�b��gy�ع2���0dm��U:օ!FP�ē
Ĭ<Fx��4�?B��x�g͆z+��T�����Vt�Ir�S��:m�­�JMԹCb���o��Շ�������A+괣`fߎC�@��I��(O�P���_q�� `7��b)<��c�O0���I;�i�P�׽��4���]��!�$*
,CCb�όT�N�;O!�Ğ�gi8i�RFՏ$O2̀�Õ�u*!�D���`О<Z�1U#Ѻ2!�d_�R�₣�2�i�+�����'D��"@O�>#KT#�i���T�<٠ [֒��6��c��`aGMS�<q$��7��� g�M;�d���J�L�<��B<y���lӳ]����C�E�<�S�#7���SfӲ
���["NX�<���@6#5B�P墝�ͬ8��E�S�<9�IZ�@kv�B �V#9�E���N�<��fu�q�d�#t*Q3�`B�IP:!��UT��Hb��ʹ}dC�	�\��B�B��J��4� I�Pv�B�	��=�,V S��@ t`9R�0C�ɹ�J!��S�]�p��M-��B�	�S�}���ʫ�d�I R�`C��$��aD��z*t�yg�HT�"C�	a����*A�o�(S%��D�B䉥':f��j�
E���*�-����B�I�H�65��	�Y���cKJ�KEvB�*a�T�7�G)9D~��*S�`B�I�:�@�ꔪՐ`^r�i��O�5�6B�%x��AS���9$��q$A8�dB䉟tmԕ�(P�86:�&i˫F��C��0hV4q F�ӓ"3"���^�C��C�I&��
�T;NB���j@^��C䉨�DŨS*Xl�"
�'�f��C�%X��a�MȰB���%J��C�I6���k 	Q�����N�C�I/[�ܩ	�Ņ�5�Ja�$A k�rC�I�)@ەl�r� 	*���Y#~B�I0b:(Bt�JhB�� ���ovB��-ik�)k��ڬG��`pƆ߹4lHB�	�_�z�a�F�T��Kb��i�LC�	=W�h�a�C�G�KH�^�L V"O� ����@��b�,���� �"O��#��K�"��q靈�nT
t"O\+��6t���%y\T,{2"O*p�N�5It��`,G[�d�"O>�	2�K$$�2ab��z��j�"O6�"��عew�]K�/@6M6	3�"O�H%gJ����P�V/d��"O���(
3C1�L�A@��4c"Ol�g�Uՠ<�  ԎB���"O��G��-	��I�$��/�Q�*Oi*A!0Y���r �Ƿ>vD`��� �}�EΆ�c4p��/B�e ���&"O(0�b�R�-����S�?T�9�4"O���g�i�u9�ƙ�u9�8��"O�e!�h��k!�i���>��첃"O|A�eė�g��̢RřM�	�C"O­Kq��>��]�&Í �n�H�"O�y
���S|��I6b��,*s"Oĸ���4�@|!� �<����"O���䁙�J�½�`�1���$"Ot��kR�EL\i�Q%6m4q��"O}�Qk�g���r���w����"O�i�����\9!뙼-�!���0�����݁l��k��z:!��Л0tع󆋠��Y ���4�!��Yղy����H�a��3J��D F�U��σ/k!�A�`E�y�X�W=�p��J'q<p�U��y"^����ɡ@�����ϔ �y�+#F��S
�6��Zw����yg�_:vPK0J/`�XY��]�yr�֨q�0'��#�>{�ȋ��yB���T(��r���M�\��N���y��ɏOǤ��#.�����y�$N�`���dM�4�TI�-�y�i
�'
���À{�"����:�yh]�@� �7F܊@.8�T	!�yr��3����A���?�H��Ҫ�y���J�{��9�����;�y���A��҄@E�Du�]�%�8�y" ��&� x�*L�9�q�J���y��VxQ��H�"�D������y�l�=P�4z��(81��	%���yR��#R�L��b�M�.���%E��y�DӔ�` S�ՁY�)X�� �y�)H�{��s%�B�R��4��=�y�T�[�P
,MBHթ�(٠�yǒ=����f(1������T%�yb��.��Y�GG7�nI��y"��
*�J���AT�M�F��y����n]K0m<.�TH����y2��4t�ڀ�XR��R��y"�	o��=x'*��PI@�RR���yT�`�&l0���I5�U)�'�+�y�l�'j4&�0D��k<HyjDD��y�E(�8 Ѥcם^N�%त���y���k�b ��Y�W���p���yB���rIIbn�9[\����yb.���c��L�\P�*��y���zrpP@r��9S���(�X��y�m·k�p���Ô~��y�2H]��yң#]HL�����7p3v�Q���y�D�	-��S4e�4p�E�0�yBΕ7+�T@��JzZ�ճ���y�@�0銸�PeөxG����(��y���9J(Lqz��+R��yt���yr�+]�l�a��+V��)C�<�y"���.�*�C_��B�ۂ��y��4;_�<�C�A�ZN���S�y�NQ>�� fɘ�bxTe˚�y"A� ��0� �\h����	�y�T�J����r��X��͓ulH'�y�g� ��I��L�<Ke��ĩ��y2KJ������>k�y`�	��y∓�2:�"`V�c�00�b	�y
� �h���?m�̘ҷٍ�8�kF"O���6iR��Ѐ��b�2}�"O��;��3K`�P̖S�25�0"O��c�o�.yX����(0ӄ���"O)1�Ӯ�l���	�)v�P�"O��Rg�M�opj�g��4�$�F"O�Гb��8��e�sPI� ((�"O�puѡ.W"M�"d>\�IW"O�E���[G�h�'�S%9;N!�q"O� ��*�}�����@5�xt"OL�X��]�]X^y��g|ʨ�5"OH��Ř~��Q䌽0��h �"OIJ��@w_�h��I5K��݊�"OnXy��}&xt��@��9%"Oh�)4���kz6�{Q�ܚo�81"O�i�f&V�V�*Ոa��%ӐU`�"Oh�����,����G�%�&t"O�B��B�râ(���7R
b���"OB��Rh�a�a��F��+RdJ�"O"Agf�9g�� �Ơ-F�,�4"OH��c!Θ8&x����\:K�-�@"O�pi�E�X֚����=AnuY�"O:E�&��
ܨ�R���B��p��"O�2��G4n�ڜxpeN5 &,Q�"O�a:��%w�8�CK!&�~��"Oԛ��x~ɣS���I�-"O��[�'C�j� A����7Y�-0�!�݌+v�r���F�j$��y�!��t@H�h_5��@�uQ<o�!��_C@h ��ˏ&Xt�g��|�!�$T丩R�j�,nР+��%O!�dT�ax��Pԥ2Bt.M22#F�Qp!�d�{�Ii��ťX:H2q��0t�!�D�.��e�SI�>Z/�#1�Q�[�!�H:8��I7(,,���Uq�!�$G	?F�	a���A>�����!�d��.f��r�nM'4d�ə&Cr!�dӜ/��욁��B2���A�w!�$�	j�>؈��ę���E ãnS!�$Ƴz�f��E�N-	Ui���hB!�Q������P���&,�5M�!��f��kS`�9:l-!f�Q7/S!��ɱwO����Fdoʵ��If'!���gQ���决i���:�W)7�!��>A֣X�\٬!�/؟`�!�d��� ����Ie�0��-d�!�$֪S�^l8�l��TN8X�ꅺh�!�C�TF�3��x:Ag>/�!��K�,�0��)�� L0�0F�"h!�D9y&�0ǈ�o�T�Y�E* *!�R$$�(Ƞu������2E�<F/!�D��G� d
 ��K6��k���!y!�$ʂbWx�Q�"� �f�yeʴY!�D��dH��D�G*L���I�Ȑ�!�$��m�r-��pS$eQS�(w!��M'wA�)���:{;Ji���!��[�'&�Xeꍟ'И�C��V�!�$���(�B#A���2�R5
�!�D�/W$*��F��:���i��G�V�!��Щ��p���l�L��v$W�}�!�DC�"��bf`<pH!�0�
�@0!�d�5a%41�Z6���g��
�!�d�
C�6����☁�p�Хf�!� !)�j���y��u���@Q�!�� ؄�p�H�"��X�rB�AYtuAU"Ol�`�x�됡^g��h��"O�1(�@˥}���bE`9��Z�"O��k�$�;4��+G(��e� :�"O��j�#��!��] 	Ӫ(��"OV�����5fI���dҦ"O��{��ε	n0��^��["O ��1���T�
�Q#K:h]"[t"Oژ3���
%}x��&tF��h�"O��/̇h���CcնA+�;'"O�h���' QiӔ���!Z���"OLL�uY�W�ԁ.&Vs����"OȨY�jލB����/�DfT���"O���+��s�� �mN)K]lY�1"O���DL�8=����4!�N0��"Oj ��.K�TP����<�4�B`"O ���[�?�X���N�>�<�b�"O�;3K�%a�� .��%��͑�"O��c 
(t��/Y%P�
,R�"OН���T�*�#���6��e�"O
PC�LY2l����N{�ABq"O���*ߎ�BM�5�C-(nD`1�B,�r�i�)ܤ|�ԃ�B,<O@��Rd�8,<���Ҧ��Y[5"Ol=�Vn��0��|��g�E�L}��"O|��/�����/R��^��"O��1/+v*� �P�W��|B�"O�H����	6 �"�N��B"O^�M��7­�%-:�� j�"Ox��@�53��#�ݒ6�n[�"O���n�?0�����Bc�	[v"O:(#�#D�U��L8&ʟ:Ak�X�7"O>���Ƞ<YZ�[�
�eH �t"OƘ�"�>L
4
��V|� v"O���7C������$D�q��"O�!���X7G�3Ǎ�\����"O���7��4��q�ƒ�����*O:�a _�>��\y#aѣP�*	�'��h$,ڢ*ȱ R	Q8<r�A	�'�\�q0i��Q h Ұ?����'�R�(V�B��`Jfe@�]��'��{��O�O2�XX�͐S���r�'��I�0�J*7�� ��>�`��
�'U���@������ 2$t���'�8 "��y���WR���'J�ԁUn֢c�vA�Rl�%.�M��'�2�h��J�$<�C�6(W(D��'�����iy�@"R�ܟZ�z]*�'Ϥ@���$a�>D��j��Q䌉�	�'ĀX�Ӌń�\sCEG�[�\�	�'Sf��p�,:��bT�Ν<�J��	�' L`�$%V�p��M�%���x	�'�=Y�@�3"�s�">��	�'S�|�2�Z�7�|��RMƭ.f�]��'��Q��+C� ���P%G�%�X���'0\�"��)Xd^���U3 ����'�
#����4���D-Rh��z�'VD��OBL����L�At���'/��y���j��%�� �.�����'�p�a�L	L&T�O��1�]�	�'�^UӁ�������"�*t���'K��C��
�s�.�S�/4Ӛ���'(�y$�C�?Q�(��,�5*����	�'D��;�!b���#UfPA�\1�'8�{ś�5R �S4뒒{3���� �Q�N��*���3� ~� -j#"ON��oU�(�6����	qD��@"O"�(�O�4���z�EKe�\��"OʔYb�L�j
^h�ꙴpM�m�"OL��1�G2R����ӥ���"Olh�V�g�6-D�ĬE"q�"O&/>Ԉ�Mȝo��y1 �/n�!�D�".x>�	���� A��
���<�!�D�8/�4�&M�.:Bv��w�ږ^�!��L.����eũf��-�Gʄ7~�!�ӝh���nW��9B����7!�d��q6-h@���;����b�q�!�$�'����R���¯]X�!�dȐE�4T���-b�D)x���<�!�$#��sFg�#T�"�*�e%�!�dNA���IM�L�L��$&@�!�܃#��U����Y��Ū���{�!�D
 ��y��ǃ踀`�_U!�Ӹ-�F��,�|X�H�B	!�N�zg�ɑw"H�m�*� ��w�!�D��
�P9�IP2Ǌ5R�a�/�!�O&ḁq�s���qoN"!�$/SZ����O P7�({s�
�G�!�dP=I�S��K:/����	�!�䙧|�	HT�=&��2�V-v;!��
����B)N�@E4�#�Jܬ6.!�H32v(�
�O�Q�f����.!��8�PL')�7m0����+��m	!�٥~&�!WcE8.,n@��̦_!��I:���E���~�x�ˤ��ai!�-}4�ҥ�U�x�Dh�A"��oZ!�DԺ9�4k�`�J4�EF�	}�!�$Հ.~�� ���(?�� ���o�!� �T�D�-��Ӏ'� yz!��X��0��hF��_|��Z�'��ܨ2�D�#��a�Fɭ�rUq
�'*P�֣�3��\��Q
l�\r�'��e؃�#$t0&��1Z�'���*I�mfb��-I��Jy�'�\�wNY<?�Ĥ
�%� u$�'����礜�3���#0'hjH���''�e���	�`�{#�H���Q�'��)��M;:-���#s|��	�',E��?D��(���,7]	�'`�Y�B��;["v0��9��HA�'����GJ
�x&x�!Åa��c�'�~P�F�5&n5���$6��'�` �-��|^Q0kD�3@��
�'��x ��<$\�F	Z+� �
�'�raC���-+T�Bӎ_ c��@
�'x�(H1EZ�X��u�b���`�J�'��Uʔ�ɻT NdX�	�=�fT��';�0S!b��M������9:����
�''��@�
L��$:/
2�Z X�'&`9Ȥ �1a:��D�(ϢAH�'�~�X��֔gF�AqTLM�%�ʴ;�'��M�wDT���5�t��5xT%��'
����@����5ä�ي�l��'����&�aQ:��jZu�LC�'����c���w��2i�Q*�'%b�/Ś+�p]��v��'�L��3V�b� ���\ ����'��| 
��b5c��°(N���'�FH�Nݖ|Զ��R�N�XU, ���� \�HV\��
��y�f<� "O���_|�Bh��iC�,U��"OL��u'�I	Mi�E�w�XD�e"O��QG�:�X��E�.�V=qA"Ot���Y1TQ	�ր�0�c�"O��6�\5W��y��V02X�4�"OB�`��ڠξ�P��G�l���"O^� E�?*[dy��*����M��"Oji���.���)2jr�zuJF"Oj�YŊ�ue2���
<�4��"O`ps�FT������.��#�"Oni�� ^�.�K���8����e"O�5�ٰ��m�9s��l+ "O�mCjʟ�֨��LQ��2�"�"O"�b���7g�6�C ��/G0<��"O��A����pRB�E(j�A"ON�[bo8T�!�M\�,��"O�`���B���V���3�|���"O�� ��́[|�z��(G�-:b"O��A+ĹD�P�sF׸O� ""O�ؘ�%�Є�f�rGи:�"O*@�E��G����̆?Fv��0"O`����n���ڗ�<L�tx�"O��Jc�S8F����
���"Ox�0lR����d��.$� Iv"O�h�#�0'0f!C��4a����"O����� "��"�'c�V$�1"OB�I���*+b�E��M�@����"O&@@`ŏW���]"I@0��"O�U���	(�ٰrC�<��	a�"O�h���T��Qs��4�Ш�W"Ojx{D�0y<hY����R����"O��	�^J` �efM�o|��PP"O��s��ْ5�a A�+<i{C"OvA
$��*W�x��bċ"&�<��"OX��D(N�Q�j����A	"O�H	cȍ
r(x���֪{� y��"O�Lٗ��� qIR�Y'~�\���"O�,y�T�%.�A9� �(di���"On0�/ϑF�~U��$C-T�4�!"O�u`� I�x8��$��\Ш�5"Of�z�)�.@�PĆQH��A�"O��u�ȳuV�QpDkS �2��%"O�A��-���ғ�ʁ)�(���"OL8�q!��-�8�1	���p+P"O�k����M\X}�r����"O�m�G���{&��#&����2��"O(ɐ&-��+�t��C��܄��@"O:|r�ˊ_h�U��eD.D��\8�"O���i�'z��Acqe�3|��ȁ"On��F��XS|0�p�Y}޾�Y�"O�Xa� �ty�`j� afj�D"O��!��H�WK���F�5QH�k�"O������xM,	A!C�4I��M��"Or���ҳ+�z$�s"��z�~Փ�"O�tpVO�k����CgO��b���"OF=1�)ֻMm�EK��>J����r"O��cGOƥ���s%��8>�g"O��iɋq�tњGDX�NdЊ4"Op<RG�|����3F�A1"O8��A�����ˊ���T�"Oh�9��ߝDlX�БHj��IX3"O��:'��_��DKU��(���"�"OH���K��R��Q��ٲf�@@�"O� :e	u��h���b
��܈"O�la6� !ZXV�@�;V޲�Ʌ"O�ehE*݅R�!�3)���a��"O�M{�ł,X<��(��B�i�C"Opp�C"�]OL���<٤К�"O���1FY�fL�(���&H����"Ox�{�N�n�����u���aR"O옰��K'^߾Dv�?T�ڍr"O�2Ӏ�(lZ�1R5B<>�ґ"O�݀��E6N���l�* ,Z�"O��I�+C���L��!W�i�11A"O�ABw%A�R�@A��G�,mx�4"O��(po��!��pA�F(S�<!�"O$�ڗ(V&%��8� j�V8NL�e"O��s.�kk:��r���HF��Z�"O8��� Hn���'�]D�k�"O\�U�U~�L�G,XUହT"O�h# Ô1cF5����=B�l��"OPl��+ĮW���Q6x�6�)�"O�H*�-�SL����s�(,9"O�L1�bو#�H�ے�R�Q��U�"O����DD'&&���\b�a	�7�Py�L��Dn�;"e�|F�R�}�<��F�$Kt����F���ТRz�<!����a%KƢ�u�D��@�<1Q ��W�АB!ʂf�{G��3E��{�)	T",��e���<ɕO�e�Vu{�II��*T����O�<�V�螵9  U4�X��l�A�<�1�-w.�Q�G/�L��0� T�<��&�PII��Y.ް�b6�v�<	�d��.�&%`pM�)hH�c W�<s�өG��q�i"�
Q�LW�<�W�6P>�!�A�P�D��Ra�S�<�#`�,c4�@�-~o�LSs��P�<Y׊�&uM�I��J|�p �5�]K�<��LK+A{��ӡ�9.z�tOXD�<��bɆ�8)�&�/;X�5Q�LRB�<��C8l���E�
#��<��a��0���c�~�#a]x�<�i3�h�#!�"��ERF�v�<1���,�k�M�4�e� -Rv�<�A����V���3������Ss�<i���:H�-���)0HN@+��
m�<	Qج@���u"N'�R-k��@a�<9eDĈG�vԲ��%A6bt`5��u�<�Q�-Z�0�k��$1 ���PZ�<��I�k��DR`+��$*&Ģ�C�X�<)Ì�K����2�y�.Ͱ��z�<�c'݃z�W�)Ru,�(3�Rp�<sAV'	�X݂&Q&:>%�7��m�<��*\G����@*]�^bd��k@�<Y��:=�P����M"�� /Mx�<��\�z�����C�f僱*t�<� �Ě_P��b�>���3��h�<Q�	��t:*�5��[��Ma�<qƘ�-�������#��@8� Z�<w���\N��pc��=���!%�W�<Yw�*$#l�b�1
�X���Io�<�%]17J*���N�Ŗ$�� i�<y��=2@H�ᄁ3V������J�<鵈D�d;�ʃf�q��1G�a�<�3
��TH�ԥ�Ɖ9pN_V�<��ў1h��!"-W�3a���T�<�f+�7�R�Yt ^2{�pK�M�I�<� Z��be͒A�X=��d�0"O\��)�)n)��
Ai��t�
T"O��x�F�0�ε��M�g܎���"O�]�C� N�̺�ၙ�8I�"O��8ċ�'(�"�Z�4(�hL�v"O�|�S��H"좶�خa8b!��"OH��	^�K�DXQ�-�$�б"O����S�!	|DӔDPe���"OH� Wg��)Bv͊�8X�4"O��Q�@�3WJ��ɔ-.U�LQu"O�q�bF�%�P]�+�7%V��"OZyt�v���I�~p�-r�"O�����]�F3�Г���s`|3D"Ob�8�y�`$��fD�H�zYD"O|�a/�v�/C_� 9�"O̸{�,�B�0ę���P[����"O����@�b�M��ęV�bt�"O� ��H�8	��P0jJ=<�h�y "O�h�f�j���kq���&ضX[�"O�hX檟; �U��G�1%xde��"OD �
)!�0�*%�)Bi��!"OHI��ʍAò��&_�=]P��c"Ov��KΛG\�T�Y��T#��yr�-[����u%�lB�S����y��9��U�aCҖ'�YE��yȅ�\o:�he�=�^��w��	�yRN�АA��"�X�h��:�y��U�e�&͙'��~VV��!�C��y¦��j��DbT*1�0����yB#� s﮼��M�/��p$-��y���'v��h����]@S�Ȉ�y�����h��
ג}��r*H��yB�Sb�p��gH4r�0QC��yb���#��i�RE�F�1P��)�yr@� ��-C3����r11�8�y���[��p�W��$ِ���y�c��s8pR��E'D;"<�l���y�;v��Y0 ��S�V��V�
�y�5����'e�HB�P�'!Q*�yb-(G� p��	AIX��l�*�y�AXL��j�JG�9�0�+e���y2e�0/���1|Z�����yrC]�O/lA�rl�?D$�P�m���y��љ(F��C�o�/:��ɣ1n��y�'F@�"�aӅ�4��{"a��y�⃗*��S(�/;�A��ݱ�y�ő+<�Hs�U�Z�􍺡��	�y"!�%S�-��hM {�~y�q�I��y���$F�̓"-Y=*L��c֌���y&V-Bd�E��`�'�#��_��yB	B\J����mStu�u-�	�yE[��,M#1��{u������yB����Sw挏@�BhBԃ�y����?<,YI�ȏj���fi��y�o�/r4P`r�M24	<H�@��y��s5�` �рY[±{���yB�Y3'��j���5&(��@�H��y��)@{�u�G���NQ��Q��yR�ڷ@�\,��lS��rЩް�y�ٞm���ǮȬ-b�a ���y�E�' e@�K*�$8 
]�yJ�k h�B?�,Z'Fϲ�y��H�Ix"�qG����q(��Y�y�+:���`�}�z��C�y
� ��&.]6�
�cUoJ��65�3"Oԥ�⧖�$�v��A�^�7H��"O��P!�-M�NQ
���tt "Or��cA�'���e�:8~�i��"OKU�H��&C,wgaRr���y2j49�J�`w/շh<�#"�Ҽ�yB@A
R�. ���#]
tY�ś�yҥ	&g8��:�cU:R���bW郎�y���/F�1ɤ]�!8d y��S7�y­̀�q&�[��|
�jM��y�!N�z��1�	j {ԭ���y�hՁ|u��jd-��x�i�ś	�y��8_�x�����b�@BE���y2��0�D��Ks�l���˒��y�kٙ\�("$�n��9����2�y��ևU�Z���l�#Q��FK��y���qў� q�T�1�g[��y��`Ҵ��f���:��l���4�y��^��*a@�#� LK���yr����-"r*�!k�؊���<�yJP9n��Q��l���	��K��x�'j����nƟ~/��A쌞n8Y��'�\�:I���h��n�g�ܰ��'�Z�7�"P
�kZ����Qd<D�h!k^�j��S��,&R�IL:D��r�V�S���Ӆ!�1P��q
8D�D�T�X�,�f����ϵL�E��o4D�P�R(�CX�0 ��J���1�/D�liEJ֖3S�T�QE��
��j�9D�02�2%�2e+GX�=d�$�)D��#������kץ�:�	P�:D�����$�yr��4q�Y8�9D� V@E�HP}��oS���F%D�<���0X%.}Ra�ҳ<�.��Э#D����n�f��CV�E�IIV�r�N"D�Ο]:L z��޺i	b�� �2D�8�bCH�%����)��z`Z3$>D��w ��{l��Rƛ�Lظl �;D�lk"�9s���[U�Z�Z����P&=D�d��B[\@XЋ�@�ֈ�"#;D��C��J)Pjz�c"Q6g v܃4F-D���b�(�2��B�xC�mJ!�D�2*������)�!��\�.B䉋B�,�r�ۏ>l�p�M2PB�I/(�p�h�h��o�+�Ά'��B�	Q��ʲ��`tv�ST�CD��B�I��,�a��%M�<��¯��,G�B�ɶY�Ӥ��*xW���q͉#z�C�	Re��0,�4?ڛ%�K��*M��N�D���Q)!��bu�0cJ��ȓ ����#��;�,��+A�l��Wm���RGz�X(�aQ�m�b܇�5h��h��F��LX�C!oA��ȓw�D�SC��:�T��rdH)�ȓW>�cahV�a�f��C(���P�ȓ6|�;�nH�0�&���V�I�ȓ6$�(��̡e�ĹQÏ*l�����U�`Yd��Z��5	�ѡkLe�ȓ��3��l��r�W�i܆�W����'����h� �?!�D��B��u(!ò>E ���f������O�Ep@"/9x��Rb'��Q�l��ȓ� Eyd�W�4?iʄ��!�f���,P����8.mf�XQ��;?%��S�? 8���X�z�.ѓ�!�:O��[b"O`�K�%��+�z�86&˒o+bE b"O������* �.����tȉ"O\Ec�^X�ҩK��D�r�@��"O �Rp��#|	\�g� .Eq�y� "O�;n�7r܎�����"b���"O(�J1xv�C�ʅr���"O�\c��]#��({��G$5Դg"O\��v���WՄ0��O�Iz91�"O��1���'~��U[t�%��<�"Od0��e�
^PE�W��򂤹R"ORd3W	S�<M�̣�m�W�f�"�"Onu[��(x�d�m�:[���p"OڐQ�ν}Ȁ\�T�B� KW"OlȐD��7=��Bd�� ���Rd"O���⩑����!�#��Bt��"O���(�'G��]Id�-+N�""O����+Du:az�+�F���"O^���i�!3Ȝ *O�4�"O��p�F�wNn���k]�B��u��"O�+�ˣKYn��a���v"O���.�:Fo������,5wD�'"O����*�r�V]2��.�yҩ�OP �DH/������y�K�qFM{4�D#����� R<�y&�{�z��e �e���*A!�y2�(~��p�&K�U��A�yBJw���"4HA�
l�M�C�[��yB�!5L� 	"�@ᅀ�y�b�Hv�y&C�Sj�Bn@��yb�:))d�e�ڰxzQ���ʏ�y��&� �R�]>N�U*6���y� �&6�,1c�i�]��3ԧ^+�yR�^�Qh
؁6��^������P��y���C�\�c�9Xڱ�����y2bO#K�|��aN�23��-�*��yR���o��iQ��ðf����L�y��3%����/k�Z�ۧƮ�y�+��v��s��M�z�&�N�y2������\,	����!b���y�(F���I�2�+p)�C&D�2	�'�ՉT��3yn�A��C6C�Q��'������,o�܃�J	=5�v���'����ą	LН+F�.Ѭ�z�'�
U"�M�����;�(P{�'_��
�|̲t��Ȗ5CRQ(�'W��/�CTU+�H[�0�����'�	���2��˄���$�mi�'���12	˂f��PS.��|;
�'��AgB@6�e���R� +�'��e�AE�3W���R��}��ܻ	�'�29�VKO�o.02"��|��A��'SV���h }Kv9Qh7JE�=k�'�m�è�1k,>�cAǁ<=�x�'�&���ܒ(��݂0C�*:T\L9�'�,ZqeP� ��T8p�ͫe���a�'���i�ղr�l�vfٕP�z��'�NtH�C�#2�H����Iq�H�
�'�H�U�K��(1JVW;G��1
�'�j��b��L��U�E>>#p2
�' �8�����ո���+़�'I)Aq(ڷe��-z�)�#V�`�	�' ��2�	 *���F�/��		�'�@���eV1(��	�'�u�`���� �q����.c�Ƚ���(L�p"O�e1��'xL���D=N01"O") ���O2<��#/҆� "O�����*�(�a��͚]T��C&"O&p��Wwx����;@04"Of�9�!�8�Ⱥ�gJ
Lq�"O��ҳ��c7d	�"F�2��H(�"O�9:�JÇ8�j��֥
�S���
p"O`��"�DyJF�	���je"O.qJ"��p�h}�@�WNڌ���"O>9�OT�?�2zQj�(ؐ]K'"O6��g��P���8�)ߙ,��p�"O@\���B�n(�| VN�/��56"OV�1�dɜ�HPJ1o^�,�	z$"O��)�*�s`�a�Ô� ;vݙs"O��J�)��ܥZ��	�]$6�w"O�L�7C�N��yp3��k���X�"Oh]˵�/xeZ�����	M�L�Q'"O� Е�� 2U2�z7��)w��Q"OT�jW�t��蛐n�UN���&"O>lF���h1���b�O�\�fx��"Ohl�5�@�pu
٫NM�J�v���"O�!֮E�J�n���,B(H&��b0"O΁�@���tӕ래'�#1"Ov0���ߴ-��{��T9%�Di�"Ov ���'K�!��_)Z�@�e"O�§�V�/
Nȡ��W."��H�"O���#f�)�p�-�S�,�"OH\�0��q�� �ȣRt"�q�"O����� "����eUN9��"O������~�̍3�,�>��P��"OPh�U�U5M�L<���S����"O�}��R�BV�s�j]���Qu"O�]�@.ZW��{ CU��%��"Ovx�mW��ƥ����N�*\��"O �z3Ν5:r�0�P���j��!�"O昪�!�4P��#-��ޝ"�"O�)�4�D��!���zs"O�Hp���Щ����lcU"O���SK!�����Y;�� ʷ"O��pUŏ�\嬁�V�
�K���E"O6�8�}׶<�
�Z�\Ʌ�=�v� ��_���rg��7���z��p���ql��ȝ�)ϔq

�'`�L�痔T�Pl����"(K��
�'>���i�\�Ui��wX ���'�B��u�1���%��p�����'6��ran��f�Nt��� m��{�'��|B�nY�%�8AY�
�x?��0�'�d�Ċ��%Q,t��m�k��h��'͞r%`�7V<�l`b��"I:�'��=�7O94R��8�_����'����k�E�z$ʶ�� w,f1��'0�9B1_�@ $��,Y/]O�=b�'�@q���0Q_nQ�W��RԀ��'e�q�fH�.�ha�艣NҤ�
�'�q���R�D�aF� �Ig6}�	�'�Lz!���n�δQw�TA��U�	�'9�BB	�X"TD�,4=B���'o:pJ�J�~'~p�b'

p\�'����NO
hŮmh��Rb���'�Vqp��!p��m(��V���'�tչb�*Y�H���L)w���'Rq��!X%��;Q�Ҝh`����� �����K&6�3]�R�2��"O����h��)z�q#Pk�>+ ���"O$mzu�]�K4-��I�2`X�"O��� +�	�-zt�U6.f��;�"O8�۲�qj@���E!
y�A9"Oh�؀��6d�Eё���{Z�ts"O�Q�.�)���w.Q~evU�"OR��a���8�bqjgO�'.^��#"O�`��(�N�|ء���	X|��"O��cj£��\�f���iRΙ�7"O�A���E�nM{���dQ�!;5"O<aSk�*T����㎿=�v"O���Rg��UGW�O�PL���l�<�!):w����O���\PDk�<	��C.oRu��&ͥ\��A�a"j�<9����_���bkּ$�{d(�e�<�Ecú}�Ҥ���N=Y5D��`�K�<!U��:B��L`"i��=�2��ep�<y��jK��V��<dN�k�<�SK̪.2U����$ �l� rϖ\�<!f�I;f!`�:���: ���"V~�<�C�;H*p b�}9�|@��^�<ubP�[Խ@��@aRE��^�<9�~� ���r4�`Pw�s]!��=9��P����,�H�8Vǀ�<G!���O��Y��J�T����6��%[�!򤄢,���KD���Y� ����-5f!�Z7��TRa�R �b5*C�_#>F!�D^,��9�A-�q�� G&Ч!�dA#=0���-�*���ҍ!�䑫uP�SeA7x��A ��B�8�!�$�4Y�L�*��%~���W�qY!�D�(P���{g*�=�~��E/� e�!��(��sF�V=v�.�G�x�!��F��Ae�
4^yr�c�2d!�ܤb�~a�AǇ	��Q�#dמ9I!��2qy>�cBG9_����!"!��D� �TԨq�ڄoST�I1o[?!���>	$b�.1AH��P���Q�D���D,���@H�U���`bm.�!��� ��	+�䔆�Z)p��ڝ c�	Y��H�*�K��I"YO>u����; ���s"OT]�0��D#PYӧ�<�։y2�>AA�'����A��*p�\�Y��'�h(C��>$�r������j/�|2�'�ʆ*��%xƀ#�[
k^:@��'n\�(@ U,3�u�ˆG���'<ִ��j�o4�dR��ޫ1�(8�'��X	�F�/_�񙵇�5x!�|��'y��3W�ȝ����e�2f/�1J�'Htг��$s�P�	�F�X����'�8lb��&ъH�g�$O7���'�0�t��²`�w s�Ÿ�'�<���%�(��GG��A�3�'{z���jH�f`I#V����6�'D �s����E�y�Zd��'W�4�1��!�=���$�c�"�c�<	��N�S�M�3m%cX�,C��Sa�<�����,�4x���*L�|����_F�<p-�JG�Б��''8��v�@�<y���|xf甚j4�ɐEB�}�<I5/�#R{�0r��#�N�C�w�<�v��# ti�%LL�*S
����s�<�C�n��R���W�n���r�<� �(Т� �G�� hI4�@���"OL��&��7R�Z;_�YI "O<p �G�iL�K��|�(�P"O���g��}0��`&��_y�92"O�T��݇}w801Q=Ds�e�!"O�I�a��}���bD�D�;�x��"OT�%�o>�x�"��r�@�P�"O�0ce�
�H��%�DlP>�޼S�"O�Ғ�ӚT�P����9�re"OL`Bi�&E���IU��/xYD�K�"Ovtˢ͖�G&��
W措P����"O�$�gR����@f�0Ie2i��"O|@�r�׻SpA�0Ñ���x�"O�	 ��vr���$'��5#�"O�Y�eƛ:$�x�eO���"O�{� {�2���NU.J�A$"O:X�1M�
��0��_xa#"O�0�
S2.�j����]F�4a�"O^ʂG�'�p���j�EYQ�"O�U�E��~�%C����y��Z�$���v���EJ��yreP/$� ��I��")�Ժ�d��yBmE$*��ʒ(�����Ϯ�yRJM�8U�%����5���iG��yL��}�(em\<'2|A�j� �yC�	T08Qs�U����X��S�yB!��oB�U)�+�%'b�,
4�V�y��T��,\�BȑQdx D���yrOˏ�\�D��/+��X \��yҭ#&�^����1!tPoּ�y�̌mO��3�"����h��D��y��]'��H����\��b���y�� ��99��Y�N��r'�3�y��gOb$�F�̶z^θ)s"�6��ޔ��LoX}��9O(h3����$h��'�A�(�*� ���z�,H;jz�@M�eP��������L?nbD@�!�.cHh�h�g��Ms�
B?T`H�f͖,���t�Ԅ~�� ��,�s�x�LN�^�<��+�5����uӚ��b�'���<��o�D�~nZ7{�u� �I~pH#F��fbt3��?�L>q����=�^�0u�\ _/��@���.Q���۴�?���:���R>�m7���"AZ�p8|A��$^�X"P�*O�0�!
VЦ9��I!'��Y�@��9"7H��
S�Y���S�-�(:��z�%Ȣo�ԥ�iA���`#�rI��;�Q�h;N�{���7@
}B�Ѻ���s;.A�g�L<��i[\^�-zJ>� (�pTry���̢gu�t��+}}��Ӭ�?Y��_؉':��'���v>�����L���r�T� ���h����O��ل�Jm�z��c��z�<��l�&�Mk�����|"���䝐9��L�䣆���H��h����#`Ga>b��D�O���p'Kqm�ԉ�-��g�Dl�b�@�O?��Ar���X�� ҥ�H-��Ȉ���	avx�&޳P���hua��b��E�TAG�#���,j���5�яMw�$���
�X��i� ��ǎ.���"�C�Xw|�q� �O���<Q�����4LvD0���C:�Qj�	5���hO����%A�k�IP�"Z�y�V9���OP�o����'H����j|Ӹ�d8�II1x��j��ƇVƘS iDE�qO���C2|:@�#�H��^S>��C�xW蔻�O��
,J�_h!�T��(=i��$ �m�H90'����C�ؕ$Z�[k]yDdx��#��i�mM���1��PC�R�'��OG��h�Wƌ��0A�'d�3.����-�)�����%#"���4����A �q�'����}J6�i¿iK�h`�@R�#"Ҡ�I�Y���*�'��l2��qӔ�D�<�OL�'ق��AـU�0�*�l�8`ٖؤ?~^X�靵�&�Y�]�P�����Ͽ��I?p8�V�ފy3N����殮�����N��eJbiBԦ(iLS~$̳D���Hm�aj8:��`"A�y-rh���i0HmJ��?�B_���<��5:�Kń<;nI�qa@�)�\#��@#�?	����D�O��'���5H@�lv��A�>~DT������I��,�ߴ��}�:1֠�G' p��ك5ז���Smy2b�l	�6�8,Oڈj!J	�k�������0�����i��!�|PXW�ŕZ ؘ"�
�^�ڌ�SB��� LU��� L�Y�"��,X(�kv��k��	�`X�e'*Ȉу�$S��S�1Î�Z�|�"@�)�P��
HSp�H�j�G)�$�x���O*(z���͟4�'��*��U�_�6D0�[UD�($��<���?	�S��R"ذ��Bŀ\>_�:P �N�8%|`oڜ�MO>�'��L>��4GpM � @�?   N   Ĵ���	��Z�JvI�*�� 3��H��R�
O�ظ2�>��j& ���OP�se��c�T|h�L���$�6���ْش�/�Oe�'������͓oO�:�W8K8��s-��]�ڠ���N�P��6��{�/�#<���g��A�Ƽ/�"$�!�π(��-5_�H��gP�=E@�#�`�<qdi��gߒ A�F}R��z
��C�X0`�����`��G����%���u��Ӿ�yB�X��4�S�`�l�I^�"ɣ���xӊ-8��&X�j���<&��NY��~��αN���� V|~�3	� m�w!@�˧�YJ���[�K�-�!z���A�I��tJҝ|�c�9���.��!�
1Æ���yb#t�'�l8Dxr��r����� dK�� n�1m��#<���)�8J���Ċ�ab�x�YV[	�O:�	��G'ȸ' �۲.J�q����3ț=}�\�ݴ[("<y�4w�ܑ�3�1P�����zi�ة� 
f�KvT#<�d)1?�g��k�6h"�"~�~	�C�DbyR�L�'��l�?���֒c�IF�ԞU�)݈g�"<���"��`���*��P��,8Z6%���ө�1O�$P����<orѪq�L7�49waAu���,g�#<Q�3�D��%�b}�����t m�>�W�
�Hھc��!U��H���"v&v����Y��x̰�������%!CN	������	6?��`S�O>R�n�!F�,�L�]}"<��K0�n���I��x��]�򠗬�\@��TS~	  @�?8���5�͕
��lARC$�x�U�<���	�O�``гm�2�f%Q#�"�[.9bN�zrF�
*���{Ȝ�"V�"�B�Pj��
�'��|���T8kɔ���2��=����5\����?p�ê�":��`�@ U;nΞ��O�N�E��m�f.�*pC�f�9e�a��&��}i��RCN����pԸ�pNB�2�&�8�Ũ,�8(G��F�&�ɈA@���O �bL��:���H����/ ܽ�B�?�A�hz`NY�$�*p!�N�`�dh���?��<�R@B�lJ���<\�<�ci�O")D�''>2���S�? �ș!IӾwt�͂��XB��ۦ^���S/�*ɖ�PF_6tk�Ę��_�9�hY�r蟛���8=�d�j�%[�D��D�F�8�ΓcH<�c
����D%�~
zQ���    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  ��   �  E  �  �  �)  35  {@  �K  NW  ~_  
g  .q  pw  �}  �  H�  ��  �  }�  ߣ  7�  ��  �  #�  f�  ��  ��  1�  ��  h�  ��   �  ��  6  z 0 � U �# �) �,  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B�Ż9�`��Ɇ*���S\�@���%A���ƭ��U��qKe|B��$/}"�M���a�$M�$i�F=�fj �y�H�,�.�Y���b�2��Un���y�5*�6��h�KC�����S�y2D�P�ơ����n���!��2�y��� ���G�U��i�@.9�y�M�8t�X�{6�_B���b�&S%�y�LǪ��y;𡎯L+�L�e�/Ӱ>�K�(3a�J�E
M!e�[�$ H(D�T(g���c�X@t�'-Ԛ՘s�!ړ�0|�'d�R(��( ,�#$���2��~�<QkȐYK�Q�U�B�4a�թG}�<yt肸{+ �p��t�5a��n�':ўʧ5z�9��'�����sEʒ6t`(�'��~��T�,U
5EG��
L(S(�&�yB]�S���J�/8Nƽ#C���y�íu��P�Հ���2�]��hO���IV:\��U�rf�"i��X��L�-�!��6zH4�R)��(0�4��γ�!�� q+ �	�# ���ǲS���"O�,�u�L5R����S*~� (8T����	�^e%�gƋ<0��tY��xL����)�&&����߂M}���V�	:�"��M�vQ��j�f;��� � �t�`��԰?��"����Cpd�l���`G�A}�<)7g��*^�Y��ȂY��H�	\u�<�q�~�@�qKO�VR�u0#s�<IH�v'��It�"4,d!�qΖJ�<g����(DZ�pCp-���C�'9ў�'�b4�𠌉R�n
�m:JU�ȓk������{n��Q�FM������IV��~�hJZA�ݏ(��-1#N���xҌV�b�䠣�J)t@H�/s�H��:.~�%BA�ĴР��Ĳc�ƁD}�R����I%��Pj5(ʋ3�q���)(!��2S�&H�t�@:}Ȕ�a"��!�D�;5�J��4@l��q V��!�ʀQ�ȼIW��$T�lM�X�hH�+O�����_oX�Z�
$��Rz!��=}Q:��7Ç-UpN��1cLu!��L�C�숥:fd��G��;!�;ed�G�(��$#E�Μ`!�\ �P����t�J�{5��- !�d̷}��1�e�������C$
�&�!�Me,q�n
Z�F5���آ46!�D�D߲(��&p�F�4�͝/x!�$Ŗ"F>�r��E<��@ EI�&$�!��3r^A�@�˰H�(����!���42� �)�	�n��*"!�ĐR�I��/vI�ڂg*D!�dO7	��
�k6#G6i"O�5���؅lkJ���;B)HI"O���H�?h~��k��Q
!(�y�"O�M�v	�'k�J=�ch�#f���"Otyb�	S�|�VhJ��h��7"OʡF��*#���!g��J���"O>�Ƞ���,�P�Ra�D�q��	��"O����BM�nLf����� m�R��"Ox��N]TƬ�S�@1n��q��"O�`R�/j�H@���j����u"O*�B��c�x�����t�(�"�"O4Xz���^�H�[�
�
ܼ���"O��I��ʌxh��aC��0��Z�"O2@{�)$�X ���4X��#�"Of�1�Z8O�6��d�R��aa"OF����R���X�G�>Et��"O~�{�cH)�
LZ�@���G�J�<Y���oHL�aP�.n(����D�<��@���%�iپ%�^uXW×B�<Nۆj� ����:?����Vw�<�'k�>eQ���"3OG^�3Wg	p�<JT��$�����+L��MS�Vv�<�� D�/~1�g��c�@D[���u�<��F"Bq�_����Pai�<��T�c�P(��7v�����d�`�<i�F�-�΍:SK�3Jy�g��v�<	�L�6A B� T��7��SBWK�<YV+��T��������!u��^�<1t�	�Tf~�J���e�J���e�<Iw�@?5� ����?>j��8��_�<�%�J;�l�a�1C9<}0��[F�<��CJ�e�P;�Bײ(y`��3K�<���Φ*��X��~������A�<� �Q��ŉ&B��@�i�!��E"Oz<@����`P�ѥ��U4h1'"O2Q����0;�Mj�����R"O��BII�/b�JB�4��D�""Ob�hDD�!�Ё)�L���Y{4�'"�'��'�R�'���'�2�'�Tҵ#K�
�R���ؒW�V5��'$��'���'��'���'���'*�}BBMXM�Tl���R�x�T�'�2�'ur�'���'���'X��'�v��Y���1(�k��(f�����'�2�'�2�',2�'�R�'lR�'�|aP�P�$dI�kQj����'G��'���'���'���'vb�'0�k�)ϐ:��|��9E��q�'��'Y��'�2�'���'"�'����Nt:��$݃n$d��D�'�b�'�'�R�'=b�'.��'Ϊ����U!{o��M�4jB�$��'"�'�r�'�r�'y��'H2�'>��eOB�`B�#;��<��'	R�'��'6��'�"�'���'���I��.�p�&��T��uiR�'���'	��'�"�'�B�'���'�P�r �ҴF��XI&�Obj<�F�'R�'�r�'S��'�B�'h��'�%Җ�2ib6�rD �[���B4�'���'��'�2�'t"�'���'�JL�E��6GO�Xy�,7m�D��A�'�"�'���'���'�"cӲ���O�(�eRbĢJ�nA f~�ܙ��ry"�' �)�3?���ijT5� ��2R�L���ڶu��� ��������E�?��<���Y.�3(�)k?�ԫ�O6`�Ě���?�N�>�M;�O����M?Y�4��"�fxS�ۑX�ʈ��k9�џ��'1�>� G˫R�����%�lB^Q���M�w�RV���O��6=�l�Jp��"[<�;q��I�>�����OZ�dq��ԧ�O"�����i��O���1��Y4p�a��,Zf��~�x�����=ͧ�?�ц>g��0��uR
$��<y.O8�O4Mo��	;�b� bɈ�u-Z|�S�G�;&:� ��H`�Rl���|�	�<q�ON�"RkT�e��	��BZ,�zj��H�IE$�2��%�S�E�΅ɟ�`�(W�)%!��j��L~L�I7��Oy�\���)��<���"91R�� A�Z�윀��\�<11�iN ]��O�n�I��|����I��@M�/�İrf��<���?1�0� ۴��De>�Q��Ktb��`G�1؜$�A��Lu6�d�<ͧ�?���?��?��eP�&R�i�Eg��w������ĝѦ]Rv�ퟴ�IП�&?�I=�� z��#(�e�E�Q=R!���O\�$�O�O1��Y���	uX�:e�a�k�jgޙ6�	p'�I(���;A�'�N &��'�H[![+TR HXe��'X|�8��'.2�'�����V���ش>mԘ���Oti
���?r@�Xr��]���:��D�F}��'Yr�'#Pd@FX�F�z��#e��j�q���lt�&��`��b�Q>��ݳ*��|��NI?<}�| � �9@��ן�	џ��	埈��i��� �1��,��$zvG�,[�|�{�k�џ������#�4c/v	���?i��i�r\�l�����i�J��dx&`�Zv�2�	����	՟ (�����ϓ�?�@e߃A��H)��Gb��h9b b�n�OZa�H>I,O4�d�O��$�O�,�&e]
6�@�RΝ�0�Y��'�OF���<)D�i�r�'?2�'���9tO�e��-�uҒ�bE�B�����	���F�)
vONB����Q��^!���c��a�P�Hb�)��M�/O�	�?�6�7�DX��m�F/�dö���`�{ �$�O(��O���<���i)L��FS'r��ضnK(0��υ�xe��'x�6� �������O61'��$&_�p��	�P C�d�O.��M�6�6?�;_0�H�'��ʓ�Fy1U�S[�ʕBՄC,�͓��$�Ol���O.���O:��|b���3��  �ƿSF �"�.���f�_��R�'���I���睥z������0x��q�� ȥK�X�I��'�b>�Q�����̓Gh������>z�Q@	�F��hzl�y���OD�hK>I+O����O���Do�aa�;@�2[%��{U"�OT�$�O&�Ĭ<���iI�P	`�'bR�'��]"$�z�	�e���ا�$�b}"�'�2�|�@�q������~��*����G�X�zAy��%?�P��O�܄`�Fa{"N�%|�d�"W�>�V���O�d�O���?ڧ�?���, Dh��j�2Z�:�:�  ��?�#�i��P�'���f����4���k����6�ʸ�Q)R�;�
�	ƟX�'{����i��;�"M��O��zr��/�8��qB�iAa[�#r��Dy��'���'+2�'��� �Q�:M�Q��+�.xA�Ϫ?��	�MS5@F��?��?�K~�zO���c꒺{}"�;g$Z�y/@�Q3T�\��џ�'�b>%(v��>")�ԏC�x7�1�+ע-����!�=?q�C]�NZ��������D5Q�2���;�r���4x'����Oz�d�Oj�4�n�v��L�)�b�@>P2�3����r��eCĀ��yr�i�����O����O���V�bî�b��֞�8� (�t���li�F�L �E�8�'ؿ� �J��=d�,0�	�Gzb!�'5O����O��d�O.�d�O��?Ay�_>6��8AjB���TQm�ԟ��	˟�ش
1��*O|�ls�	9Tqҙ)a>c����g���'���	؟�S,;b��oZ]~RU�tl���ީ`\����V+\{8�
q��П�
֕|Q��S͟,�	˟d�&k_�<EL�N4)FF�@%�@ڟp��|y�Fs�R�	�/�O����Oz�'`ެh�Ŕ�=��P{3nP(f��Y�'�F��?����S��2"y(�� �b�Љ�t�C�U�� "�E��+�����<ͧ&3��	{�	6$ ��fMջ6�hMKU��'c��	��X����)�S{y�Hoӈh��;sҔ-ړhJ�.X8�;6�3;���O�eo�f�,��	��YW��~&�{�N���1�����	,(��oZd~r�u�\M�}
�N��xw@�����3Qn]�<�/O0���O����O<�d�Ov�'!�rq#��ȸ-���`��м!hl����i� \�U�<��Q�۟t#����A�L��0�3�B�U����į��?����S�'(�b�޴�yr!t�^�8�@ 	�`�"���y��łs ���)r�'�i>�������Ge�TT2�˗:
��l��ܟ������'&�7�V(��d�O���A�QԎ�NŌz�d�#��#CF⟀�O��D�O��O�側�9#%<����PuF�Ԓ�<x "۳i���IJb��h�rI
�\�O�?a�.�C3*�GH~i���ޟ�����(��ݟ4E�$�'8X� ��v����%�t	�5�'��7m�5���S ���4��у�4�|$K�0:>D��:Oh�$�<)'�4�M�O6�c�����#��;6�DB �ˬe�$D)S�3�@�O(˓�?����?a��?���v���r�Ϲy��1C�G!�P\�/OL�l�)oO��	��@���s�Xy��B�aB}J�dP�{��4��-�����O���1��iO[|��qS��;9��BC,�8<09'�~�ԕ�'0����`�x?aM>a(Oh��)C�?�4ܹ��0V:�x����O"�D�O��d�O�i�<�i���`�'����� 5�,�r�E��H�,���'6m:�I���d�OV�d�O��t�!Wq�I�Ǆ���F����L��Ms�O�)�����"����wm��)b�=h�8\Ɂjƅ =a��'��'�B�'��'���E0 ������8M�(lY@��O���O�Io�)%J��\Z޴��D�̠*��W�.�<�Rᝩ
:�XL>Q���?�'+��4��4����x���A�=pe��)(s�Z�%	��dQ�䓇�d�O��D�Op�DO�:T|Z"-�2f�f*\1����O��_��6�I�'�^>M�	K�>��j��x?�\��#?��\�����d%��x�|@р@P8�q(fz��՛g�+(U���X~�O&TD���1��'4䬒�m�4�NM"��2��%jW�'���'7b���O�I�M�f&B�H��7+�I<b��G@�/$���BY����4��'0b��?�f�=E�"�;Dˇ�o<�t&C�?A���]��4��$Q�(�&���O���.Jb��Q�P9D�%ȴmZ�`=>�I|y��'��'���'&b[>	���Q)W�"}E���e��*�a��Mk�k��?���?H~�ɛ�w*��5�\�1�4ibs��%#��Pk��'��|����*
��&9Oj����Y�
�t���;?F�x�q8O��+B`��?�c�*�D�<�'�?1F�k3ppqk�4$Y�

��?9���?����DZ���uoJ؟x����CD-T�ob�YQ�5!����*�s�|��I��H�	t�2*����ǋ !��8Qᣐj��5B֡Y7�R����|�'E�O
�X�&�8�"���xT�O=8������O��D�O��d�O��}�;K�z��@l�$3�<�;d��b�����4&ڤq��?A��iN�O�_�XS*0q��-�D�U�I�7��O�D�OX,�ADz�X�����d�?����U����ᝓ<�X�[�O�K�Ry��'��'��'wR��K�UЧ�Nk�ά���Ȋ,���M��!���?I���?�K~Γ*�l\�$(��)�ܡScN��ER:�X�Z����&�b>��vK��QX�p���l����΃�7%2�x�e*?����znB�$ʔ�����L�R4@drWb�}t����J�}����O���O �4�.ʓV�dG�e���v�tU����2�"0cQ@V��"�v�
��ӭO
���OB�d�A����3od�^�e���X�����x���
�cS����>����<��)'�<^]�Pb��Lm��I]��L8���X4\��[2e6E�r��ş��Iß(�ڴ8W2��O��6)��/;}H9�Ea4�()I��^,$��O����O��:(.6M4?�;}b��G�x�\��u�4Up�p��j�.�?ٷ�<���<1��?q���?A4��$�*d��5a��I$��*�?������@�@�ǟ����(�O8D�5 ϩy��,�V���BNH]��OD��'.��'ɧ�iQ;����+� J����������T�~�>6�Vqy�O������v�B ��P�}B������?���?��Ş���Ȧs5@��f�aA����WaS.]ov��'�t6�,����$�O�K�k�$�8�0t��[�&j�O��Yi!F7�$?i�#�*7�I �� <��LK#e%�u@��HwzB��0O�ʓ�?���?���?1��򩅆*:��D߂l'��	�F�t��lZ4t����՟$�	J�s�p �����Ě5yF���@.W+H����ȑ��?����Sܧ/��4mZ�<��O�}��+r�ͮ+���x!��<��'K�'����K�RyʟJ(�I�>_��d"6�Z�/Fe ��''�7�K$u���$�OP�DL�`]�<�'"A�v�i��(z��⟌c�O�$�Or�Op0�S�_�n`VF@�w~F��5�����@
HNr4Cы\�SIIr�OΟ��w��rf�6JޫasLLs$�����	�����PG���'��YR� I�5]B�ӖK�X��i�E�'T�6���S�T�+����43�B��x�<���w�r5j9O����O��$�&P��6m*?��G0[�����9Q��R,�?v�!3㋭)6�0�K>)+O�)�O�D�O����O�,;7@>[�nE��䅠}w.	`n�<7�io,]�S�'e��'���yB`�6��58���A�֖"r��tQ� ����%�b>���h	�0��8����Z.�dh��#D�"?��ϑ/-L�d�����Ĕ�n,"h*A�^]`�4�QB�nk"���Ol��O��4�@ʓ��6�^,5���\��l�;�O�+���BE��y�BwӴ�Ĳ�O���O��]�0�\RwE�D@Y8D�ڀL�V����g�P�k��ڇ����>���BY*M�d�Y8"�¹�a
��>� �ğ<��˟0�Iޟ��	h�'f�����b_�R���bw&-�r�q��?I�Y��&�U�4����M�M>Y�Q�T�1Ѥ��t�S������?Q��|b�*���M{�OR�V�J3�5s��E7L� e.�MU��9�2/��O���|���?��Ak������UӘ�@�f��;�65��?a,OD�n� h|L%��⟐�	_�d$�4��H��&��6��l�V�T���^k}R�'2�|ʟ@�r� �{�Hi��8�B�2-*���s�f��x���D.�^?�H>)aB	% N�	�������L��ɟ\�IƟd�)�Jy�b�Ĺ� �T�?�p=�3B��\��(�E57aD�d�O�yn_�/���؟Pw�Ԍ@ q���ofq���\џ��I�~��l~~#P@�0�'��P��u��(�B��R!�Ir�<i��?A���?���?i)�މx#i�9o����
��U��LĦM�'���P�	�'?牕�M�;UӲ��abE�x����d/\�n��R��?�O>�|:ժǩ�Mk�'����SfM(W�܅��J
un*C�'g��s%�韈P��|]��S[����y(0Ey���(Il�������џH�I[y�#x�f�{���O��d�O��S��Y�U&�a�$��#"����?������Of�<���֓}I����'Ȱ{m$�`�g;?a%IW�h|�����P�b�D)�?)�a]��H��81�~\������?���?����?�����ON�e�C�bЄ�\,0��$�#O�O�oZ�����	֟�X�4���y��M�&,VߚS`!����y2�'���'j��JD�i��i�y ����?��hT�㎃�|ڂ@�ͬt�'��IƟ��	��	����	2}���bj�;2��c�6mM���'��6��5n����ON��=�I�O�����6JA��"	S�/��Р'C}��'�B�|��D�=WLa1dg�-g�4Dã�Ӳ�Pf���d]�)�)*�,��O����P�Ѓ�i�\
�Ǎ�	�L���?���?���|:(OP%m� v$��I�}��A�GF��@��E�����ɐ�M���m�>���?!��@q����f�'A\s]d qc�Mc�O�uA�Ć��2*����d1��iJ2��y�F�@bgّ�<O����O.���O@���O��?��A�%�N�%�l��$������H��ҟ�Qߴ|k���'�?��ig�'��L�@��
L�@I�f�
:�����|��'w�O�h���i��	�7��t[��͇|���6� {����A�3n��/�$�<����?���?�R'�
|�1���ސ}",� F	�?	�����̦����Hɟ�����H�O���dÚ0W��M8��x�H9��Op��'h��'4ɧ��W7F&2\0% �i�*�x��̄/G|u�f��T�=����<ͧhA:�D�*��D���#CU2V�ّJ�,�y���?��?i�Ş��[���s�\�h��U����5�K�gYn��rN�O��$�٦I�?9�V���	8D`�t
�.̘� 8P�n��3i���I埠aJC̦�'���Fqܧ2cd�$W�K�x���Y4*�9����O����OX���O���|�D��+%ޥ�CL�<�* �t��*c֛6I�:4q��'������'V7=�*=�'�4_�r��"��^] �R���O�b>��I����ΓD����ɋDu�)@0댉z$r�͓/�И	t��OĘ�M>,Oz���O ���
�����ٶ[��I7��O �$�O��<)"�ie�a���'���'r�-2�@�\F���W-eа��d_C}��'��O4�I�bŏ?BP�4nH�sh������dj�7w���u`�T��6r"`�Ɵ�AA�Ơ-��(��g�-�
��0�^՟h�	۟���ß�E�D�'!H`�$��V�rV�Z� �����'�7��bπ���O~�l�G�Ӽ��≁��Z2�D��dZ�<���?��M��I�ڴ�����5��π H�xDjۄ	Ln|`�'Uad�8#�-���<a���?!��?	��?q�<Z����)�'.C��������L�1��������	��$?�	���l��Ѓ ���i�'N |�O^���O(�O1�r$��G�)�%#��	2W�|ˢء}�Ҙ�@�����FW2C��a��sy��̤n�~M�SE�(&���@	�N,��'l��'��O��	2�M�3�I��?	�EO 2�&����2�`�����<��i�O��'%B�'�+Չs*��ɖAbU2gj� :��p�i��ɩY��B5ҟ���r�.ձW�Ĝ9A�դE>]p�m��I
�d�O$�$�OL���O��$0�)'��a�'L)x���賆�UXH��'��i�@EXQ�?��ߴ��X� s&��� �.�k�dC�?-�H�M>i���?ͧ5�bA �4�����:��u�P�d/<hJ���$3�tl���9�~r�|�P�X�Iޟ��	ן,��IM��"�0�F2kb�	�(������Ky�bnӞ���F�OZ���O�ʧH��a�,)v�� q���/TΕ�'����?�����S���0MC�X2͕L_��Q�� ]�M҄�^18�\�9�O��=�?�s�+��Ǉ�X*�M� .�����؛y����O����O���<YӲi�E���5db��+\*�]��)H�|~b�'�27$�������O��	���^�<�#G�}���<y�L�MC�O��[d�O3��wK�<��߇jP��ռ_.n���@�<�.O|���O��d�O��$�OʧyZ|����;8r� r�
��2��i��D�@�'B��'���y�hs��l �x�`[9@1< X࡛#���$�O��O1�agw���I2fg���ݳ.�^쀁�F #����/��}�R�'l $�l���t�'��h�t
Y�l�� b�f�`B�'�"�'B[�0��4��Q�(O0��\�9�6��cH�D��	�L�F%����O��d�O��OJhs%��s���J��[�J�����@3b���=f��s��&��=br�ɟp�H�3�\�r�T
�i��^��|������ٟ�G���'[�e� ��4J���dHY�;v�1��'V�6�M�i�
˓b�v�4��A`dO�>��|D��U�8��6O���OX�DT)h@J7-'?i���(���K�,��G�RY�����T�٤�$�����'"��' 2�'�y��F2[�@$��M�Q�!^���شA� l����?�����<9��V.{z���B5E�@��#��,t��ן(�?�|��!4n�!�a�^ݢ�� /��!�D������H���Ewj�O�ʓdʽ�w#"����$m���?!���?���|-O�tm��1�4)�	dm�0�'GܷU��-��k��&�P牧�M��>Y��?���`�%�f�A�:��i"ȝ�_K&:g�O�Ms�O|-9Eș��*��T�w������ ��ЉA���P3� a�']b�'�b�'���'���q'�\Ar&��rg] A��C��<���_�v�����t�'�f6�7�D�?=>�B��'S�(��"ݲ:T�O��$�O�ɖ)�|7�%?�ωG����$��K�4�s�L�S�����O樲L>	,O�i�O4���OP���@�7w��z�
ۯS#@�s�F�OV�d�<�ǽir �`��'�B�'��"Y��0'��R6Հ�f"z��j��	����	b�)AeJ�aÌ\�+\����	�p0���ܩ���ȟ�Sc�|2e��P[�|a�lY8'��7�^�$f��'�r�'���t]���4�a�Y�Q,@� ���6=��͐�A��?	��	t�v��^}"�'�!"��Ya8�]`a�Ҙ.Z��@f�'l�Dօ)�&����a,�A�S�.�>,Ѯ��1 *lK4��IF����ly"�':�'�"�'��S>]��֮@ͺ!U��-��c�Å��M�U)��?��?�H~�4`��wl�1ce��0
��'C �'�����'��|���h �0ʛ�<O��{�˲N��5��nM8�}(1O�,k����?��=���<�'�?�� `�T[�#�3w
���k��?���?�����ͦ����������$�!�I�a]�Hf.�2w�HkfE
r�&��IΟ��?YDUadB�	񩑂=LȽ�!+�M~��.ڒ\�aF1$��OіH�I0$���ٻ܁�D������S�*a"�'��'k"��˟0�� ��.<*Y�W.�~�2F����z۴Jxx��-O$uo�m�Ӽ�2DB�b!��6�R��U��<!��?�YEkش��DD�<�Tѐ�'$x%S5dN	$&D��M�!��j4�7��<�'�?���?I���?���$�ȜcV���*��J�/��$�������\�I͟('?�	2�, �b(D 8���M�G�XѩO ���O��O1��%�6��!k;T5Z��'t�M��ES.0��FD�<�7�͗E����������#J4�yW�߆xkpy��f�?�&���O��d�Ol�4�^�o�����q$Mį1�P�ZC�����
	5�dI���M3��>a��?�;P��i�lO�3�:��g�8��|�e#Ł�MS�OT���ք��S�%�����L�!ɡj��j���w��]j8O��d�O����O��$�O��?!����U�h���킬X�%��byB�'�n6-�8]F�	�O�tl�y�	�m�L:ա	���+E ֿ}L`�%�����擎�0l�B~g�4�� �U@ƞ(w	 4�rf���J���?!�  ���<�|Γ��e&�1�:�H��̾ho�0DxB�k�N�c���O����O�˧r,1$Ƈ�
�T��f[�h_F��'�0��?)���S�@0\�!Ae:?�x�	��ѕc$��c��,9���Z�擊P�. x�II��;pI�$F�=r���N1f��	�|������)�qy�a���h�=ow) �+F�(�����.L���Ol�nZQ�T��I�+�",d��m����bJq����	�R�Tl�S~��/c� ���i�i�JJ¤S� O5p���>^�Mٙ'b����I��<��ӟ|�	Z�$����6�RD4���,�*7�HA�.�$�On��6�I�ODnz����vg�,��y�������8�?�|R�����M�'��`H�o?e�N ��mL�n\�j�'��)S֬D�鶕|�\�h����t���5=�۳�-$��A��`�����xy�(k���V	�O����O�$�DƞB",�wg�-0|}�`+�	�����O���r�d�J0X´�NT���L0?��OO2AY?��'Ji�����V�g�p\�e�X�e�F�#�$ZX$��B�O���7�7p�% ��ĝ/��Z��_�qɜzbW�kx�d8`�le���7``��*��M>����.Pw��|�����y�U[��4rJD�5 �#8�^%����R�A�#A)B7��b�lR�eV�K$�n):�´�),�E85��~Vr� U%L�X��舑"�)j����G/�V.���4M��JhB7H�g��
$ �D��H� �#~�6����l"�/5Y�l8��O3F)�զ�L�r���4�?a���(��I{y��'!ɧ5�*C�#����T��!U$V�/w�(�'�Ɛ�S�|�'���'��IeFp֏�w�z���K�H 
�3DD���d�<����?�	�A�� �m&���	 �P� �����?	���?�(O<�sP$��|��i��?t��8p�4iAn=�ʐΦ��'1B�|�'0�l�w���@�E�p�B�Ci�(zehRj���ן|���T�'��S�F�~��E�A
���=Y&$b�e�
���Խi@��|��'A���T�qO�i���qI~uȶ�֛*�@� �i���'��	�X��ѭ�����OH��U�[er��d��*�I��P4�='� �I����+�N����Nġ,�F���]&1\s�ͳ�M3,OB�"O������I�?�r�OkA:"���ɥ!M�x��� �Ē��V�'��O�4�O��>�I��ۭGg��Xn��ts2e��ow���������ݟ����?�a�O�ʓ5�HЁVn��3\BE�c鈆��|{��i����G�d:����*W�˻F�
�(��8C��u��;�M���?��*n���X���'��O$i@�✂0��Ѧޛ1�i���Lc��O���O��$I[�&�z���7�*��F�0G��m����"Y�����<�����c�V8<u���IF�t�B��A�W}��Fޘ'���'*R���Ƈ�,����Tfҡo���"s*�%M~XѪO˓�?�K>A��?�a`�Qgt�� ���{�BŜI!l�P�����O����O�ʓsL��#2�~`Óߺ#eb�*@�����4�i}�Iß($��	ß8�s��e?�p��	���I��- Z���,�}"�'�R�'剚	OB�a������0�"��3ʌ;p�5Q�Δ7*�ioğ%�|�Iğl8���c�Wr��̘'D������e��|n������Vy+Q��'�?���ʔOZ�w@h�z'J]=:T"�.�J��'ur�'Nܤ1���?mpԇa<�<��� ���Թ�8�+O���������|�D���'-B�#���_��K���(3��Iܴ����O��Mb�{�$�O�yBb[&|�q���+ko@�+��i�h`(�dӚ���O����$���)v�Ġ]��ɷ�ӥ4�Tt�ܴ�?y��?�L>�����0Wn���gʁ�8��aCn*ymZ��$��ßLJ�� eyʟ��'��Ѧ�H�Z��d��iq�5I�#k>#<���)�O��I�T�\H 4I!Ftv���&4��7M�O6X�֨�<�5]?i�?��bȰ?g�Lȱ��&n���K���'��!щyR�'��	���Z")�
{2��aLB1s�p�3MA`�0��'�R�'�O��$��pu�L5g���y(��.d��ه%v��`R��O�ʓ�?au$����Tl��E��} �b�e��).�M����?I�"�'H�ɑ]:7-Q�x1��ږ� w���%�.,�'��^���Ʉ
���OFR.F�k*m�����,�ґ)�n<6m-��ǟ��'I�L)N<Y�����
BŠ]�}�S�~	���'��R�t�)J�ħ�?����b����@b Q�!���%����u�'�"�'�"�'Z��yZcC�AjM	1�Hk�A���=1�O��DC�$��d�O���O$�I�<�� ���)��
:(y�� �Pp�YmZ��X�'��}y���TA�(|,Dt[�'��E��bP�G�MSC-��?���?����,O��(|N��"��ߤC�ɸVKK�~� �O�����)�S��#%ˈ<u���E'R�wM����F���M���?Q�	�l�p�x�OS��'�ԑ��R#1�n-�&&�v��١S�oӶ��O�ʓT�3?A��?�Ci��" 8�c�k^�EOƥB7�Ê��f�'�V�"3�)�4���$�O��" � �tB���/:a#�bN�Z�fR�iI�	�x�'q�'��Y���&�߭��1r4I�a a� �8&��=1�O���?�*O����O����)����R@��F�R���x	�i�59Oʓ�?I���?i(O�����C�|�f����1[b�%��a���V��Q�'2_�T���<�ɒvV���lT��U��:��G�NȈ�O����O
�d�<���F8/���Οh���� ��;u��4�`�@4��M�������O��D�O��ɐ6Ot�䯟 Ga�|PHxq�dL1!H�-��Jn�V���O��(F��X?�Iҟ���EI,���kC!]��𡍜m(� �O���Of�d_�J��<i���4�\05�M�@��K]�����M.O�5�h����	�H���?M��O�³�\h���by�!
�\S���'vrnЋ�y|r����^�h ��3S<z��aA6w����"6��O����O����D}T�$8��'a�����!�"k3F��7 ��M����<iL>��T�'Ԅ�`�)$�&)��Y.f�Z)�R#v� ���O��ĽT_���'��IПx�(>�E��O���UC	q�(�n�����'h�U����)�O^���O�E�`̈́D��S&�I�0wbe�rK�æ��I>�&�r�O��?!-O���� y�*�0�������6uh`A��^�p�J���'V��'�^�\�'�؅𚔈�o{I^,:�LHጽèO8��?�/O:�D�O��$��mFz�K�杽�b�!Vʍ�e�H@�6O�˓�?����?A/O�qB��	�|��9l�r����I�M�az�c�����'/�Y���	�������s3F��0�˰FL�Ѩ��"E�VQ{ٴ�?����?�����dϵ���O��n@f�(�1!��R��6!�	EJ6��O ��?!��?)�E�<�(��,)UHҴ9!dP#�ԝ-A�,���¦���ٟ��'��#��~J��?a�'A��([�G��$��pl�04*բsP�������I-̎����?�;�M�4�b$0�#�*�����l`���\Ӓ���i�r�'��O���Ӻ�"	�p�N�Rcg�J>R�
a��������0�m������4�S�����Ƌ�g��!�!��j7M"r�zumZ�P������S����<$�[��a�G#*�#�e��9��V*T��y�'��	�'�?)�ᚇ ����JO>� �����F�'Y��'��|Z�̴>�*OL�D���2���� �1�&ȸl��E��tӔ�d�<y���<�Oh��'�	 �.�Ѫ�#'����W��'��q�$��O���<��'��hB����搜a� ����`}�o�#�BQ���	�D�IEy£L6s�
��F��x�n�sqh?R��H:��0�D�O�#�d�O
�Uc
r��d��laF�@���31杛��O ˓�?y��?�,O��Ja`�|��a�[s��s7m��+w$|��M�O�̟$�$��̟ܘ�}�$q����96���)�>����p$A�����O��$�O�˓pĴ�y����i�O	�vÈ��JB�26��O��O���O����=OT�'��Q���<	�Jd�$>��Aa�4�?)���AV�6%'>��I�?�Q�a��\���Ck |e���ݳ�ē�?)��l��9������4h/L����"�;vā��M��M�-OfEb2�ߦ�ۨ�d�d���'>��u �zDpu
`���51�1�4�?���XQ��z����θO@�[9KRy�g�܋c_����s��yh�g�����ן<���?MH�}2j�%Y�8���ڱ	)T�AJȚB&7mވO�P��%�+�ğ��W���ȁ�ĊO4��COA&�M����?��9:-�xr�']�O�е�25b(��I[V@�׼i��'PLLJ�����O����Ov-2��V<2��I�S�ˡ/��x�@����	�kh�"L<����?�M>��(��*W�O�v��L��l��<��'�thڜ'��I�����ן�'ۈ���;f��"Μ&ao*�{��Ի@Gxc����U�۟��I;T��{�J{&4�a����H��	7�џ����t�'pԘ��+s>m��`�~":��ǫ| Lq ��>9���?�I>1��?A�LN�<I0�L�Q�D�󍋙` ��N-���ޟP��Ο��'L4�8� ��T�2:�X��מ)��m���7SD��m���&���I������P��H�O��x�aӦR�[%H s�����i B�'��I*n��H|������5"�"��`��"U��z,^.RC�'D��'��z�'��'��IQ KР��䘵[��A��J�:Z�vY��*B�M�U?��	�?�z�ONu
c ^��L
V��1w:�0Źi`��'�Z}��'��'�q��lzp HLl��
ۛ$�A��i$-��baӞ��Of�ퟨ!$���I��|�X���߈y�G��
 e:�4Gr�M��䓓�O��c� n>`���^qI�:�$��4
7��O��d�O�AH��a�i>��O� �uF
Dr�(�� ޺��u��i��O<'>5������I�3L��[q�O�"���g�E4nfh#�4�?�E��W����I2WV I��僶)� [��D`<O6�d=?�������'��=����'v���s"��bw�-CA"O^����Ng���c�cAH�ڧ��Z�j���Y;��P�d+uhx��)Q�dl�}��@~�h"tO�5LjE��݌wp���Ɖ!L��Ӏ%T�H4�D �td�c�I�+;4��+� ���AO�&/����_��(F���ؒ�)Q?���!�h0�B��ZFA��d�md�1a���1��ȩ���9��Bբ�7<*��å]�ApJ�D�O����(�je�)�~�#FdU7H���O���7�L���όsJ@2���?�J|2���RrÌE��3RJI!1�Bi�F��j���� �ֈ~E���D��k���'��p�to�� <L���_Lҍ��<O���$��Hh�X �
7#�ʈ�Î���a|��;��D�2hy�83���1EC؊ ���\�8��'��Z>5�ቒП(�I���	�m\zF`HF�U�c ���vjל8�.��Ba��WD��KT�ʧ���?��k�jh�#F�&T@�{�n�1i���u �X+�#�>E���T����5!ީ��k@6%�ƀ�1�1�?�������4�|"�Q��P��m8k��c�¯�y�H�#�D���;���ʩ�OޤFzʟ�em��Ќ��˘_M$E{%��O4���j^��8�D�O�d�O����������?���гFtL
3�D�7ԕ���_?�P�>J����j�xLGNu����L��4��|��A2�~bH	�S}�$���G�?�R��D
�>)@@�v��DDJ�á��w����cr�'�ў��'x��3쏗zv�����8N���'mJ�3�-ǌc��Љ1�F�{%I;�S��P�d���MSV
A>	���#�3������*�?9���?��x�6��'�?�3�8P�Nޱ�?!�q0� @B[7e`p��^8���3럨&Xn��&�����E��wH���k�!>&��f��(+��1ģ� �Q�*`��O��$ݓ=����!F�1n|�A�1/*mZ���'yP���bmĚ�r���	G��-�u'C�<��	Jt���ԚY'���GwrX���>��ob�4��ݦ5�G(���M����?��Ӽ�c��3*\����C�lX�ƨA-#8=���?1��a��h�Q�W#vɧ�i�2g� P �XUl�����!A�Q�PS�-�"%�E�Do�_���Qb�>`�H��E��(O^ ("�'�"�'aRQ>Q� _���f�E2'v����E�ӟx�?E��'h2�����
Nؾ-�s 	-k��I��|��'5l`P�+�7�2��ȴe��Ï�#<O��a�K��%�nl����^`�W"O�l���D�Ҹ�f"��k��Q�"O���bG47��yiQ$�$^���	�"O���	?���ڔ%
�a����"O�I���T�a�X�FF��E#!A"O�T�Rgؔ]��d�k/�1h$"Opy�AC0w���c�2>!��"Ov ص*�e�]�Vh�fb�G"O.����'\�9�g!�C���"Otm9s:,MF,�%�K�.��0"O�M���R0g��A	4��b��e�A"O���t_ k����C'ۘN�.��"O��X&41�5���>�J)
U"O���"�G(� RL-[.$��"O��'nZ5w~�Hˠj�dr\��"O���1L� SyZH9�,Y{���"O4q�煒r�b����޺j�
0A"O&���Q&Z,�	�)�x��#"OF�{��F�z<��(�(��-�"O���TW�v����\�\��V"OJ1�5͓+�������(@��)"OJٻɏ�h���6�_0��"O�X�J|+Vix&K40)��9�"OH��dgM�L������X��"Ox����Y�4=aeJ��H�(@�"O��iA�����ȓ�K�� �(Q��"O�1h��V+���ɧ#�^��`"O���<�m��o])Y�<�yE"O��s�1R��3���c@��a"O�abgDG�d������EF�1"O��Yv$�=s����b9y(��w"O���F]�Lߢ)�t�k&L["O�@+ ��>c���B�օEjF"OBtU�0���B�?&�1�"O� 
d��O�lq�(ʢ��:3LB�"O��C3�D�P�b4�VFJ�.*BhH�*Oh�J�aQ�n~�	���]P��	�'KFR��[1Ş��g����P�<�3��1@|���u�? W.  UiVG�<�`�ˇ2�py�ȠSZ��+0*{�<)P
A�u~bH�E�fN�u��]m�<�r���A�[dBxcJ�g�<a�vV���I�c���3�.�f�<��A~Z0����C�;i���\Z�<QRCZ$Q�@`V�ͻs���b�V�<��ͅ#����Q5h�VabNk�<�O�0 ,� �[.#Ƣ A��r�<�׆.7~�� ��D+\�d�f��u�<�B/�!{Cj�ڗ�)$���)��FI�<���O�*��yX�OC�3dA�]Z�<	�F��y�l�oe=�=�d��X�<)���5�ir�k
9����IT�<9�n�,U0@9�$��1`dxg�Y�<i6
=�2Q�K�~��F��Vh<�gB#�"��J�zX-�p��$p6tp�)ӽm��}��{~�k��Ĕ���C�����<)"�Ŗ���U�,�%%��N�D�R��=��8	#D�<ga�>^��A�bW)4�5��f!�dV-<��Pf�a�OFB��v�u(�58	p����
�'�4������yA��b��\�5H�x���'�bu���>q �10��L���0o*htCB�<��03F��7þx9N�����UǠ-�c�*y�a}r�9�XIq��%����'��y"g �\��+a�F;I���`.��y2�W�^��(o��������y"�2B�j�挚!�`{6A��y��ۅ[��͛)E�!F�q�K�y��+I<����2�Z�2��L�y�&@<�Tu!�����m8�&D�yb��W�쒄� ���c쉒�y�hτ`�^�i�a�
�@�5�֫��Ox��=§�n�˳�
�5kJ�r�Ȥ{�ʬ�ȓ0��9��ǒ�?�W�yq�q#��OvY�؉2`H�O�>��b
��M�:-��H�!��C䉹[k�%{g�)�|A����*s �2������S�5&���I�OvZeٕ��%~4�qs�J�|�
���J��R}��FR�Q㜨)�鋵g�h��$B�7��3OJP�.�-\_B��e�ZH��c�I`�Rd���S�< �H|�F���!QшP�
�2�C�<����Bn(��Ɠ�$Z, Μ�<y&螒���K���` �)�RH|�է�'P!l1j�(�D�ȓj�2Т�*�.�����q� }��"����A��85����#Fx�w�D�pK�>M��E@����0?�F@Z�uNl��ӢJ�(�
hR�FW�)�Hܓ��O_�*u�4�8�O�XZHݓ"��d�`�|����w�	#+뒈8Ԉ��,��-���~ڦ�� HD�� �*T�������a�<�#�(�:J�BV�������<���[���ɖD�-L:P��S1�CP͟u���2���C�I���kb�� �J=Pg(�1(��7�O(s��'A@�?#<!(q V�E��+7�(�����K���xV�#"��jGJ�NவI�j�u0B��D�dd���'�j!Pf�@=v����E��>�3���@d�0�A�F�[}H�!N?uI�W0��lޕU�t]8W��v�<���R!s�*������P�<1ѠZ/ꀬ��M�0~�����ӁM�$��bm[�Z1+���~rNC��#%�U3଒�al�8��,�	��<Q��O<`���9�� �?#<ф��8ؚ@�x�x�@q f���;�,�u��!�A�TTS�ٟG� c��P����" .�0`a�=Y�D=�b&�.z����0���:��M@yr�1klȡ!�$S��Х��� �#J?t��@4E��Q��y��"O���U��{Nx��n�n�;g6O�����ٰg��D�ל3f1��B�|�B��8�\,i�H��X4�E[������ʱq�H}�G��#{��cf�8"�[7��g?�e @/s�Dr֫����O��UƄ.+ZΈ�G�1o�5a��	�r�dx��ND*n��2u J�xU��3lD��p�.iT���ϓ����HiS�y�Ns��m��I�m��ɻ4b���!d��X��I�a�R�!f���5͠ biC3���ˤ��"-;!��I�Kf�,"�VoJ8Y�)I$T�˓��DC����H�+�l!}O��a��f	ڵv|�d*�.Ǣذ?Y#�8A���M�"*��S�A5�E�АA���GU�K�G$O�lr��8��P� o��h:��ɰc�؁���nU|�'�66Mˮr�|̋'�Mr���#�nʯr���(�'���I����RI�Dě'bH��۫Op�z�Bb^<A.O�<�S�'7��9R�/ĢQp|�,��'�������r�9%���2r�F�9��h-O����R�hD�J|j���9��-��1�ҋN���v%ٶK1|Hى�$�k=��'��풶�K����f�k�}��ω�j�%
�~��"�i���;u�Nm8��t^,�$P��& 
���>a�,��6o4�����Y� R��З�~�*� aj(����v*uh���k*��%؊ɒ�e��0��lȅ�\4E�6��ئY�U� �0B���dS|g�(�O�X��*�C��8�Ջv�,���<R�:bA8}�H
u�4[��̨cF#vd��������Ĝ
l��O���8�oV}���	�:������uT)'�_@���Hz�a4=��I�J d��޴^���V�e@,z��ؕ|�@��!�Έn�`�ZBԂ'��\�c4O��a`᝶½����.���P�R�l���=��v�,��*OFq�х���y2��O�p�3�܍q�P��
)?��͆N���0��T"��u!�	ut��Q_8�-O��*��c�������2-�hd81��%̖��e�ü`����4�'��tj�
Oop��$H�<��c��>:ܨ���p˂UʗF�;�!�˝j�g~r�ȥ7Y�|�d~Dr�Ӌ���O.���e�(�!�+��^��A�S�i���xu���gj档��V�z��)�'ۭXx�nz9lD�S �~8��
��ܢ%Zb}@@ Мmݾ|��I�>��"B�m��탵�z��ff�r�'�"hk�O[|�����C�*<J|c�"�V(<y���1h�3�� �j���"
æG��X'�3,Q� �R�a"0m�;fn��+��u�b��*0Zg���ɿ@���:wd�'v���F
My�Y��B����$�<��J��s�&�{f/�(T�AҐO�E��ֵw;� ����_��p��싽6;���٥�'D������˴&���u�j��Y
/<+���a�@H�0�!��0p���
�<�M3 >��<��Bs" h$ĕ:"��b �}}	Pa.��u�#HO�ԃs�������.̯,�h�bښ%��Xi��y"��Pzpm!1�Űob���ЮZLrX!
��6R�^c��!_���M�B��\I,,h2F�I��h��iʐf2a�D֙xX��FD� �pKa���I��2���OD�(�Tv]�P!�39:���	2;�P9�wg�,�4C��Ύv�<"?!���{Pekd�	�m�v�a�	���](��	D�i��L�)q��X����R�ʑB��'��##��;P,���Q䎜de&���Oހ,��*vO^�r��Ik4�9Y��S�i�,\�ْ ��(X�a��j4!��t��=��aڞ/�4̉�mޡH���K�ͳ�����O���fh�G˜��P�!�╠W�,�D$�rD�SX!��@�a
�L*���1I��X�NZ�U�6D�a�'�����%m��[�aSXV�M(����S|��,�9oMnE��@K)Dў{ ��G�b8Ie�K��<1��M���J�LF�(q��!�g��a2�KK�DJ��c �'�dP��F[��NTR�� �J��4
1�i	U*˩
�*�Q�I�c�V��=��5�gѵp/����*w��ɀGǑ�ybk���P��#��Q��`bqJ�W6�h�c%��-���V\�� 2����z܆TQ��K\� �g,n���� V���1F�˰0�Q3�*����!k��تP �7�
c/bK�gYرz�3
P����'R0DGz�)ʓllX<k
�9E���rO�s�to;6�Y��l�8Y�������y鈀3��,�Jd�胃�=�Mt�øE��BD��A�p����s�X��A� �4�BǮ�<v0RD"Or���jP&x}�x�Q�F�2��e!)�y�Ϝ�WI�j@'C���3�S�? XѢI[ H��p��� U,�jR"OBx;6O�a-�Yp*Ec�����"O�Yڦ��b�*�#u☝G���W"OR�S���� \��AT0k��{T*O��c�k��J�m�Ǣǟ,ux0�'��D ���8ZP AY"�)VH(	�'�@�gŊ+z5���M�#wI�Ȱ�'z��CK�19�(��ÌhoH-��'{�D�IY�w>�+%aĳS�n!��'MH����ݾx�L��U����Y�'f���Ff��9�X�;b&_��K�'��8R.@�j�DS������'��и�GJ 4���Z3G�h0�'�d!@g`��I
&H�5c� J�Ҙx�'�����]8z�z �ţW�?12�H�'�nQ��
1	�:����jL8	�'n�eZ��M���قZ.y���{�'�
� 6����س⅂�H/����'�4!CbB�,��x12�Bu�j���'4��
cɶQ����]��b�'�Ƒ��BMs6	�-N'|w��'�����ټV�����tD�9�'�
\�a���Q'�d�P�s�`=��'6�@�҈ *'�����n 1����'�V���=[_�����yԍ�
�'�pl�k]�7 `IbW��g�v

�'���1%AU�fےP���_�J2�98	�'�HĒ�l�.\U�#�W ����'�T�0Mӟe�B")P����J�' :�OZ����H��ހc	�':��ل�ǽ0��5�G�YW-P	�'�a!��7|4nuhp�F�SXF+	�'���#�I�/1\aGN��G��	�'sf�!���,j&Â�D7mc�'� ti��lJh� O+5�LC�'�t!@�Ț���ظƇD�w�&Ey�'��ek!�KMfrfS�mR�@�'Ǿ���ĎO�l�2a�0��x�'����%Ox��ԋU�V� ��'�6]h�bO�\[й��o .$C�L��'�$ՠ���1�X3�@��F���'� �P�ȟ@������2�N���'l�҈� ��uS�#�0%M �{�'���J�{���2���2�"O��	g�Kj0�P'H�w�pq%"OF$�6���N�Ag�v���ۡ"Oh��V��#Tmb��W�}2\��"O��0�Cž�$yx��ۆ`i�B�"O����΋_��mXp��F\�� "O����d�5`h� �&{7����"Odm$LX6fC�	� �"y���٤"O���!�Y�FcV�ڣ�_Xܼ�3"O��1�JN305d���M�z5�ei�"OL��L�[�`��n��[���b�"O\���N�:+;���$�-R��EZ3"Oz��w�hI�E��|��`9"O^Dk4@G*i*�m��I�WHѹ�"O�HqrL,Pp���U=�hT��"ONuS� ˼4�N��.Y��%��y˂�ƨ!kǖ[��9�c0�y�͖�f�<�LܼS��st$	��y��P}�U06���\�R(JgKâ�y��'a��� U��	LS��D��y���Y~������#<�tI�斉�y
� j���[6��틴e�""ֹ�r"O��c#�	,M�إb�#Ω)0�'"Od�hG�E�/X�tMØWZ壢"Oa�R�Q�st��BE��^��)��"O�H��I�'�%����t� ��7"O��1oė�zK���\�"=�"O�ٰċ�8*��q'-�K� ,v"OV�i���T�6�9���~�R�[S"O�k�#(���f�ӂA��}h"Oҵ�*>���h�AԽi��bfl�<y�,��|��b���$󕈘i�<1@
4;Ȋ�I!�u4)SK]e�<�@曳b��lq�oE�Qz��8!�J�<qׁ�Q��E.��%2y�T��Q�<Q3mq�ur�)\$eȈd��Bx�<��B�d����hL:.������s�<9@���pߤ`k6�Ьp�n�;Pu�<I&/ע'�v͚��˥��9�e�LY�<A���>h�������Q~B!��K�<!���  L�|��,ZI��=�#�n�<�e�-QolM�g���]4�=��l�j�<�Q�L�F���/*&G2��T�[�<�פ���,1e�L"/����l�^�<Q��6@�����)�
�^����MW�<a�k�(�Zx���-4�@p!��Wx�<�T䉚@GZ��T�,��ܡЦ�x��|�?a�n�	%���7�iז��J�M�<i Bݡ>��Qb)��)�C���B�	f�8����,�@�ôi�&�bC� �d`J�>t�8I�M\}RC�	���ݓ d�DM�*>>]C�Yz\Pq1��ry6��3.YD�B��y����Ш�>	+Z�P�'>�*C�	�<���G���	�F�)7M^CPC�@ve��cĵ�D[4�H
t��B�I�9��`�d�%3��2���xC�>M��锩�"���	3��.�hC�8g���Ad%��b��(��lW�I��B�	&�r�������]��$��B�ɫ]ʉ"���Z�,Ikf���b�(C�v�!* ��AV�C�1��C�	}�����CнH'���lC�u�C�ɸ9�j��uR1F��ĐkebB�=D� h8���&�h���Ȁ�NB��9���!H�$������r("=i�9�,�	�Hj0Q�ԏ�8�t�ȓ`�0��&c	$�ݣ��L�BC�\�<Y�e�GEDYRG�6f���-Z�<	�j�)J��0s�I�:%�a���o�<���ɓ8�:��f[������k�<���-Sj��S-�m��8���Ti�<A�(Ɔ��G��a��h��e�<iA��[��WQ[�\����	!�@:%Ѯec��
5{}ƕGb�7P!�ē�����:{C�a �Z>!�	��}��b����p���6O��|��x�� 	Tv�|���)rJ�02$�)�yBb]LA0�2`�9|j-hqJє�y�)�/l�pSh�s~n�Z��W�y"ȿ>�^Ā�{\�9U	�y�Ǉ��U2��I��h B��9�yrI�t�����Z0vK�l��Ꝫ�y2�\�\y��y���|Y��8���y"��Lwpقt�.mQ≹ MΆ�y
� �`;��3s"�`+Z�}���"O��Ԍ�;ff09�xd*���"O� �qč�3_��ƒ�`sā�"O�M�6��ccN�H��UEld]a@"O���v�M�H���"�5X�8U"O2Ahǹ�[����� a��XC"Ol�Jf�
$L����oҁs[����"OTL�@T=Px�Nֹ2B�7"O�ECBBd�la�>e#f��F"O|�
T(L�b��5D 2��M�h!�
r��%C�mԙ]=�Q�gղ�!�P�TK^x�R&]�C=�ᒣ�Q'�!�S�������W���_�!�$S(h+5K֥��=�Tm��×=�!�պQS8�CO֬^��t喇0!���;0ZEP����b5���p&C R#!�߫1ި���&H�E��L�c�3p�!�T,>|�8��$دi��]����,c�!��Оu:gn��h�(����R�!�$*Gw���5S�Y)���Œ#ra~rY�,hA��d�fA�E�Z:�hq��,D��w�	��(SJ]�C+6�q��.D��1�-�v~�8�bn��F�'�*D��q��Y�܌:$�C�C�& D�.D�p�ËT|}�%)���+0%�AH-D�D1��+��8k�G$�Bd(d�5D��`r'�� ��;5
L�f&D�\x����{��[�.X�%v&%D�d�t�J�3��K����U�#D��:� G�6��s�D�*-�yЃG D����-��X�:�DQ$}4R5:��=D�\�ael�`��ҁC���'=D����BS1G�������O���v�<D�TZ1��K���{�J->f]鑀9D��8�'2;�`����>"l����;D����]�&.�;R��G��Pj�-D��3L@2.��Dʙ����c..D���$N%�ug�.!��G�1D�����+[4Ru+��2zDp,[�%4D�0�Ԩ��~GFM�1��P�h躒�&D����cU�]�t�)K�l��Y�e� D�́�"ԜY]��W3oʍ*a�3D���A�+>H��p��	|��p�h0D��b����d��83�V2]��X�*D� !�*N=gW���Q��8I��]��B)D�D�Q��`��-`T#a���1D�\`��hӨ)��P=!e
�u�.D��*6�>8�T�6g�Ld��T�,D�����'ptҲ���Fo�m@��.D��{�@�u����a�?i��%�R�-D�(�c�ðu����rG�	�t���)D�<e� �젓�)� ^Ht�3)��<�S�':�$�5խ4�������N���uY}YA�=V�d`����?s\���ϔ�� ��?\����B��pPE�ȓ=U,�[��S���{/~��� ��Ĺfʀn��x�3aI!+�"i�� p�%X�ZJ(b�ze��BXPl�ȓ+�i�/��	!�\�s�
J�y���d����R�c�j�bL��)����ȓYm$��w ��mp؃5�\� �܇�@":����I m��uqb�:t��?;6��p�S;�f)��1p�Va��f���@D��O����W&����S�? X�G�b$�Y��چzN�Z�"O�`2�OK�dl�Պ�NUIw>��$"O������%�^૦�̶1�l��f"O�5ٖ�ĵ'8�M��Å�aD�BG"Of�"BI�R=
�'�S�MC�9�"Oh��g���v�c�ء(%Z� �"O�Aqb�B.&�.	�4�d"O�5@�-�b��h0`����R"O�=�EJP�a�<t$��(���T"O@c�̱t���IS#�1���s"Ob ��&'~�鳢�?eb�K�"O��C�Ņ%��$�uHC�� ��"OðF Q�RH�ǒ�����"O�H@�ډ=/.�"q%R�(C��z�"O�����<����RBH��6"O:L0fO�'/�A �ѓ�T�4"O�e���2S��]�ra_�Gܡ�W"OڭzJS�x�L�[Cҟ9��QP�"OzJV���R�m����x` �"O}B2*FM����ݱx�d��"O����*�����x��(1"OH;1��1��m�U+��p��"O�M	'�{�dP����;m�`�"O"��U!�^j ӵ蒣<��e2"O�q���3K��7(��_�X�9�"O���(��7��P�H��2A@�"OJA��D�k��H�fE9V�*e�%"Oh�{�ʕ���	���e"O䨈SMX�T`�˥�L�'����r"O�a��E�k�@ ���-}z�pC"O��g�L�"�H����x|�H0"O(�2bI:�v�*�
__:���"O��!Cm�� �8�Cv�ʄf����"O��s�C�X�0��ìL����"O܉�2n�(��̩p�5+�a�"OHkPY�r�>	��"́]�՚p"On� �쓨C�d��/���R��"O~�Ӄ �2��	�b. ;$�N8U"O���
!Yal ��$j�"O���Qo�+8��U�j����9!N!� �y<��Y��ι�~A:&ևH!�ċ<4�YR�'�(���Fި*O!��Ы/�#�D|���:�4~��C䉾fgE�ɉy@���B�7shB�ɉD��e���\�{��I��՚�FB䉃#���6��(M:�����^ZFB�IIæᵀ�_Yjy �f6��B�I�2H�-!X�Vu�Т2cC�B�I+Y0�������,A\@B�Ɂ�V@a�fO�K�Dx�C�)�>B�	�	�  CfĖ)9���;0%�C䉲�*!R&H̍
��y���C��/eKt�H!��/=��pVIn�4B��<"n`P�3,E�e�L�� ٞ'� B䉏/����]*}u F�X!%eNC�I�fv8[�	��W4�ዑ;Y�vC�I PX�[֪_�t� ���ڥ]�C�	>�$�ӊ%��:�d��p<�C䉽5�t���eW-��	I҈� �C��-YJ-��HͰN�v	{0 0G��C�IU4��ק]�F�d&ו(VC�I~$���Ȟ�&3`�ã�=b B�� ��q�f��
;hXsl�	`c�C�Iav�c퀐"E�y�呹L&C�)� �8�b��C��,7NK�w�=!�"O�D��GO�)Ԍ�w��hE<5��"O�j�O�W����J_�I(��h�"O��qQt�Uq�`G'jr�"O֍і�߁4C|���_�����q"O,�L5���C�#9{"|��"O\�)I�r�
���Ռ5N�\�"O��x�$�q�^�bkYh��"O��hTNZ�7[V+Lcf�4�"O�i�,�2O�İä�݉WDPۀ"O�4Xw��g>8Y��Y^A�w"O������9+�=X"���6�^���"O��xpk^�W�p�$��c}>8�"O��K�aY�U��t��ro���W"O  �c.�'V�:5����RM��"O
 �����]�A�,�:���"OԬ�DM�9N��+Qb<*$"O�� ���y�!ㆪ�d0e@R"O��U 8]-Tt"�D�c h�"O���G�|�$U��i�Gz��"O���a��/ ��a��)��{�l�1g"O�$��G�}�5��W�(�Ӓ"Ov�a�K,B��#���@p&"O��1�ʁ(%��	�!�-���"O�csL�o����U�4/�FHp�"ODr��ɇnѦ����W���	xE"OtuZB@�=%���
"�O,�NI��"Oz�Xa�9%^Ԥyq#x�5�'��H�g���\p}!f���P����'v�ɒ#�νG|.$�u��N
���'��`���=,�X{�T�Ezl�Z�'��+Q�ڊ8!�����8_�q�'¢��хيL>ՠƂ�7�F4+�'�� @�=;#�+�Cã.��L8�'u���G�	����Uc0#	(�P	�'�T�E%�Q�,�u"�� W����'��9�j��I�����	H(P���'����oǴ`A�H+!/���F���'YhV�\/��芠N�3%��X�'�I�vb���;�Dp�j�
�'�V���9=|�X�G$HUZ�S�'��])�.D�"�t����L�pE��'�(��C�T�|��w'�->�9z�'��hPF�P�Y����aӂ�K�y�H8 �@���ʑ�8���S�N"�y��ؑe���c"D��2�Fmسj���y�.Z����ą��$�P�/Щ�y�ު1������g���G��y����p: &şWSNy)����y"�\�W�εI�I=Ě��cfO��y2 _�X����K�DpkS��y������E��J���J���7�y�Jְ;�6�`ä?!�t�H��yBB\(���LV7?�0���y����J�D��A�;3�na���&�yRH�	$�����fJ�8��8�g! �y�ҽj�-Y��X�?(���	��y��1���D:`��KT��!�y���T�*�� �?+7�D�� ��y��=�i��iN9dؠ�C���y��c��CAET��L:d��;�yb�N�`�� &ܱU�7�y���(��q�%i�P��lyGA�;�y�m_;a�����B�J7&p�G7�y
�  b�Aό)G� ط'�
C'���"O@��#O 1�JHك'	�$���"O�"�^-6M���a�ܤ%��HZ"O�쪦�	!^| �E�9��5�"O�s���Rq��r��E'�N�"q"O��)uE���0A5��!���	�"O�aa�%���Y�L5,�v�G"O�H���\viP0# � z����b"O�ec��_�{�9�3�+~�� +�"O���d��R1B��l<
�0v"O�1��kM�&�I��_�4U�h�2"OIc��H�ZMfL���\b�I"O�a��[�A�\�P7��=>(Ĳ�"O.黅 ݪEɒ,�elJ�v�43c"OPEp���6~TLj�J58�*ə�"O��aɓ/�.�GjO��4��"O�ɫRk�/��LӴi �1�6�� "O� S�3�b�xw�ˊW��<�U"OP��AB�t�>��O�X��ܨE"O(��%J�_�*@�"�_�l���0"O���V�E�r�d���I��bMt�%"O����7�ip	H�y#� g"OT�BW�Z� C�Y�0�j,��"O���AI[���Y�E8v��sd"O܍P,C-�%ڃJ��Yo0d��"O���'�Y�Q*P@�	�5"e�X�S"O��JEZ�d�@ă@��8N�q:�"Oh���o�X'����W�@S�"ON�SRO�+=���v�5C؀��"O����K[��]���*[O����"OXa�[�*H�l��J�k��]3��|��'H�mvɎ:ǎ8�7�;=����	�'v�@��b�:N�@��3�(	�'i lRC�=vv20"��@��(#�'��u����T��ā�tM��:�'���4C���	1Yn�J��'U4�����P4�̸�B;^�r=���O*���ӑ;τ�%�:^L>$x�"O���gC52���%N�*i0|`�3OB�$��\7�� F��T���1D�y@����\h�Ob�� �/D��i"b�!'�*<C�і(q�5Xv�,D��ˆeܘtA�u��샷g����b&)D����摶>%�Ի�̟�o�0��$(|O�c�P�ѩ�2�<�rk6nK���+'D��#o��b��4h�	:J�5(ň%D��;6�Ge@w'R�4�"��Ӏ$D��!E�5��z㧑"^�ӵ� D��q �D&����P:����H2D� ��;oX�!a�I�SR��3t!4D�Գw%U�6!�|Q���
9\�pa3<O�"<1���"@��d���/9	T;GK�b�<Iׁ@�H����P&�l<rڵ΄_�<�bGB�]^���%���	�@�<�7O��*����D���/!������S�<���+0���8�a���Pc�Wi�<g�А�L��g�Gu�"��(k�<	E�
~ZE�!��r�\0��he�<���V�,�R�$�È-.��I�+�l�<�BbI'+�h{լ��g�2�Y&m�b��xΓ�q�wn���	p�a[�S|Z�&��D{����ݕ2�"]���/{���[C����hOq���: l�)0�P�P����T�"O �R��D3dpyb��W�^�2Ai"O� �!)��t:<t����B�X9��"OT��tN[�h�4��
E�z\�1�"O�8��R.8����ln6�TU��D{��IE�Mf*U��nH�{����f�-N!���R�JFlN��s�K�# ���
�'��=� �C�P�$���
ޤ:���'�p=�B,x8z��W��\��'��Ls��А]��ٵ��#4����'+䝙�� +��%��2�z��	�'��̚�+.!/�IXEKȅ+�r���x�Ř;k�Dī�^�A�"����=q�y��́[�N���n &Tq�A����yr���W4E��f��x���t+�.�y�*O/e�H�A�D[4\f $�$���yb�C*-���J&a��}޴���b��yOR8NL����L#b������y��
�8�̨q!)[rS��(�$�yB-Xd8��d��D���JL��hO����N
-�nl30hp�#FoN _�!��H�]��h4ϐ�_~m؄��&�!��fwr�;=��:ᆯG�!���FϦ�"qf�45L�21��|!�$Ē{����C�j�6	�D�M:"��{R�|�(�'xÄ��>9�Z�c ��8�!�dQy�N�۠��}�ę�!�D��L"��`�HĄSܠ���=JbOph�$�˰S�Jq��G�
����"OB����G�|�*d2�pq�b"O�p��	�
��Bk�
���"O��:�*��{��`0gӈN�
�c"P���I�Fx=!.�>�%#�*� TnГO>�Ol�=�U��Y2 ��[�L�i�ѯF-�?��'[��*���4t���θ! 
�'�DdLT�(v&i�D�C�"�'W�̠�gC�
��q�"j�9n��X
�'��$`S�]�j��ЉS��Z�t�:�'XBA��A�4�d+�f�R��j���hO?a��+��^�#�*�\�:l2d����?Q���O
�+c�G`6<���*�6,x�"O�(c`�^�1�6H�jA�(p��)"O�qS�v��L�HX��"O�U��g�q�$�p�<P�.1:�"O��� ��4ۢ �@���+��<Q�"O6°�l�!z�j�5i �uX2"O0���(�1bؘZ�H�3�x9S�d<�S���:w��!�.���KAoL�gb�'�ў�y�K�֎��r�A���j4i����'��'�O�Ҡ�$X��J��ݪk�lsȧe!�d@���ٛ�m�R����4J͢+�!���|��2�[�M�{�)U�=D!�̢��I�r�[���������N��p
s���BPS�����YW�<��0|��F1�d��8^80�V�t�<A.ɱ!TD)j$i˶T�=� Eix��Fx2n8���(���3f.��c�y��7=p�q��.��B�a"�yR���ՊH�� ր���K�yr�Vmh�Q�M*D�b�N.�y�i�W$�x�$r�#bo��yR� 
oZ��� ��Mk�+��<I�� *	��ӷB��;Ri�#I�-�I^��T�'eǺeBR�H�j� L�(�U�(�d=�O�0S@"�+~J�eN[6A���ɥ"O� I�(�1Tźu�u����`�W"O� ��cdы9x�U�4�G�G�
�"O�3'���1p^��AM�q}�h�"O��H��!z&B��,ǫxT�b'"OZ(�$EZ$lzg*��!@qF"O�4���=z�`P$��E�b8��"O�Q�Η)70�K�B�|2̙3"OXϦ"�&X��o�oBM��"O�����aX	��8���1Q"OlD"�A�Gм}��#R� ��a�"O�|��E#.E ��S��$�H�k#"O5`��U#I�j}	���2u4���"O��+�}��D"��Y�~�婓"Oxd�퐚�Bź1JR�$��`�"O�q3�(�cz� 
1�[�
P�""Ohda3+��1-�A��Ȕ*~;F=�"O���B͛4�t�٥�8~v����'��IA~£�!�����`�-:���ኆ�yB�^H�Ń@mΡ5>x��(׍�?��'���"�%q{\���T,�jh�.O����\�pzD�Y�� 
(���!⒄�!�9]v�˂���k��th���
73!�\�[�Jr �w�䠩W`� !�$Z:gvJhTj��s}���G�<2�{2���:�&�Z�'�m^��2���	!�D�8����¨4����n҄$!�'?�R��2���Ę#$�F�"�!�DYY8L+0�ғG	J�`�E�P�!�$ť`yfH9�E�/fM#�� #�!��t��Cd�M Y��b�I��?�!򤓕x�`���aUM�Й��3�џ�F��hI%xp�D)\�C��Y��ۜ�y�፩3�9����i�0��� ���6�OHU9�	�E��4�a�E(��"OD��$����@FgF�����a"O��cBL�Ʃ��F��8�f-H'"O�|�	ק�
�Ig%D1C���"O~�٤*_�!n�ű��M�g5�P"OP���-��(�-ח&�d�G"Oݻ��Hm���P�,�m;X�3��D.LO�X:/�;T�e����V�u�"O�I��Q-aI�y�@!&9��"OJ|p*W�~*�q2BW�L�8�bD"O>� ���P &L��RM��"O����:Qr���c$��{7�`��O����]�z�����E!zה�зe#D�(�,IS)�oS*9iC�+D�p�B�u��5`�4��@�߹e�!�;zx� B�b��.�.$1�j��d�!�'� .�Kdh#ਙ)D�!�DE	R��Wl�&f��]��H��!�d�5p�)�w A,h*��ꬒ�0�OB�I����)3$ ic�z�⍌v_�B䉂�V(�tN�>*x�3�NM��|㟌��	�`��J�l��:qn�;4��"oBC䉿LTYWI��=�x\[uA�2cZC�	��H��S�SU&JH���&/#�C�	�I2$��)4W�8���gP�.�C�	%,x�p���ǃt���v)����g�D�6��Q`��X�ꞏL��T)��-�IT��|Qe���4ʌkH�+��M�T�+D�t�!�H(�4%���5]h>չPo$D�p��
�l	y����)09�'	$D���p(\�"V^x��h�����>D��8bB�,F<l��!�uR��9��?D�� ��b�e�19dnłc9�0��-�S���<R�,}�k�bԞ]�a� ��!�$�+�lt��R�J� ���ʋ8/�!�d̕J��(���T4ny��
�t?!�$F�n�1����>���OR
-!�5�L���K�6e�mr�Z�o�!�S
%����,�����(��`�!�$�@��1��kߟ�Rغ�*��b�!�ĉ_?�-yS�ˇ��5����?}!�$��i�X����&9�6�R�.F���	S���iBlN�P�z}���`$�a�G�-D��+�	7�bD�r׆H��p�b/D������� XM�g#��	�D�(�A-D�`1A�'8����/ݚ(��
.D��B e�M�ȸ�'Q4d����H-�O��&�
0[b%ԩl����&K"I,�ՇȓX���0��Z���Y���	���ȓ^��}kT�=z�졉�����t��]�&@k��'^�^ј]<�d�ȓp<\x�k�
k����'�\��܇ȓI^\ѧ�^�q�t%z2%��
��݅ȓ3������8����2��;�&؅�p�L��7.��PT� ��Y�+���ȓ'�tI�$�N#����R�8�l�ȓ+(hW�ޥ"��10) >�R�����Ű�hͻ4�B�(�jЅ#�R,��Xu��3�#�:Mx�K��UL4d�ȓQJ��􋄁ߎ�R��L0nd,�ȓ�^��g³m�؈���V�d���ȓ|��0I�>�����/�9����q�.-�Se�.�6S���
^r݆ȓCJɘ3mA;�=Z��� !�ȓ{&P�u��.΂�)��	":�-���~�@���1j����ǂ�%nنȓ� ��dS	9�*�QH�Bz� �ȓa(�`���0=Y��FRK�ņ�&�A9����5�v=��A�&VⅆȓQ�(L�$�ݕ.}���r��/G���M_}��/�*81@�a-ג��m��(�x���C��a+��
pbi�ȓ+�
Xr%F�	ie��7��a��̇ȓ������`q@GCצȇ�}k��Z��b�Z�*���"M��H2�����izq"��<�������'�ءy�`�X��������#�'I`�1֌�c.���&� "���'�\U9�#���(����
�ryJ�"O:��t��^�Hm��W�P�^�Ġ�ȓs�@R�%^��$Y����U2�ԇȓK�����HQ4��4P���FCD��ȓ~��A�E�Y�j�Fu��F�6$脇ȓp��AGP�: 9�l�7K�^��ȓ	,�����)�}�tg�
�����t�x�aT?'E���O���(-�ȓ{�f8�M���9��^�̄�V��=�tb�rG�tӠ	6N����J��
Q�ߌ3������8L΄A����<I5ƅ�H4�⁕�g���0��U��0=Q��JJ�ȍ
���k�\��H�Y�<a��@�$���Ζ=�,��>T�X;)
W��Ѫr��>$�ܳ��?D��+v�_�Y��0�Q�C9�`�w�>D� H�45��|�7"�!ޘ�aF�&D���@-3x���$dX�g�/|O8c�� jp�P�w� $Q��4x���"Oȩ!���&W�p�э:��  "ObUdM�..+�p�'3q�9�"Oq�$!�w�y³励G	2��"O�*3'�S�6�e�UIBd�"O�YB���)s-�rH�)�F���7@!�J�P���`�B>9 &�Й*!�D�K}���+F�g7�Hz5��
s!��ve������_�6�Q�$���!��$U�%�vOR'Ξ��y�!�ā�d�����A	\�P�`a�B#d�!�Č�8��E�A�d���Sw�7�!�9��rU�V|FU{fM�.3�!�䗧zk$�p$�zb�(���_�!�dҢ�&h��Ζ�W�Ir+�!{!��ًbAt��B�|F腒�O�;!�䐩5�\�����C:v����1	!��,(�� ��Q8�\���T�Ib!�$A�7��r���<&b���	�tZ!��"W�@�Z ���,���� 8!򤜧I|�	��T�E\���ņ<!��߁B# �e�7'���;�\�'�ў���4# �a���lU�;�n����C�ɷ[�6�3w-�4��qrC�S�B��iE��#玅F3�@3���2�HB��>"�lݑ/�X~`���ճ%E�B�	�+vP8�U��bLZ���ȩGVRB�	�n���"��E����[�4B䉶T8.H�*�.���1�#�.*�B�IN���7�J(pH|i�q�#3�C�I��0(��
[�\5����95W�C䉅K����a��)�]�e��	[�C�	�C����f��$LƭHTD6��B�I�*e��S��ΪU1�γ_��B�I�!��Z@�D�U`�l0�ƅ;D��⟐%�XDxX5������ ,��3��1�y���sr\�Eo�&O�YX�1�yfS��!�V��L&�@���y�T*'�t�k�)���Э���y �Q�~
�9-c��x�����y�mBu�ؙ�'Z�o�2�:�
-�y�
�ʒc�͚hz�!ХK*�`C��$�2�i�k]�Zl�p+%i4|F,�O�=�}���+x�Z�*]��!�NG�<Q��ޞyE0��N�GEj��#mRk�<��+^R��G$�\�b8� �<T�k5e� a�u�R@R/�Ե��2D�@[!���q�v|���*-�Y�$�4D��{�%�u�d����F�pݳ1k-D���`׶���[�פC��)s�)D�̸�Gה[��jv쉸9����G�&D���D�:�F �5	1�l�� �)D�XH�D\=Dp��b��"`!r"�(D��d��"#~��4�:q�1�4�&D�H1��q��PاAޝ2�Nu��H1D�\���t��)0`Z�G*�9�$%��v����~�8�[Ӭ�[�~�B�%Y>{TC�I�!7��KtA�>y��5���V�9��B�	�S|"m)���w>����\!�B䉸J���� +��E�ca�R�q��B�I�PH���/<�|�R%��_>�C�ɳR�8��F�n=bH��O,O�hB�	<V�^���.ބU*�R4M�J�O��=�}���\�)R]�ԏ5ͬ�ڂ�Z�<� ʑ!�I�!V��T����)�"O�� 2. #V�tI��[;6�V�Z�"O.��aBRn�UH%h��J� F"O6��&@�������|wf,X�"O��@E [�y ��4#Q=Z2�0`"O|x'-��d�13 ��wSd ���'����t��y����*���ǣ�8n!򤅷��pF�M,����tBޫ"Y!�P8]�J�ecϭ/�ܡ���	ag!�DQJ���%Ig"���J��jS!�D�XԠ����7;k>Y#�	� Y!�De��|b�/T�^Y&4��J��^R!�D[)dӲ�����JM��Q�R�0#!�dK0oܘ9�H�_N���sM�m!�
 ��7��PIj���
P(�!�!H���H�
�"=��!)x�!��P?T�i3���ڭ*ҨĻR�!�D��Ty�{ �9(Сi�!�$�8y��,��A!F���sD�
�!��G�g�`��+�=:�г�3'~�Or��$Ɯ4I0=��$<`2$�5�G4Qb!�DR������! %�((����^T!���:}�s�.z N$J��Å
�!�� q�	���X��y�A |!�dU�h:�*4�H�OD�*�o�;{o!�@mS���q/X�2F|��Q�td!���P�y�Nފ���,�;!��ʌ�1b���:�d�送�$/!�d�*TU�-sn��Bܺ|���Į!!�ٚC���Z�d�~Ţ� � �!�«Kf�pvJ�&y ��� �/M!�d�&���i�a�	"�����5!��>r������ T**��Ȣk!�DՃ���Z5�K�&VxX�ڛS!�DM��Uy��]�P�ɀ�ïT�!��8dȥ��b�;v �t�qȒ*v�!�X�|'���6�T���-�!���NdRh�QHG.?�m{�!���!�XX^!�*@�ԉ��V�Y�!�$�6#�^DfV�(�xI��;�!�$C�<��#TP(�Q�+
(�!�9��7�,k��pj�T!��K>/�E��!�����j�+i!�$͇nVl�Y�F.H�b)k�*Ů'J!�d�*/
P	 ���g�9��+BZ!�$��CE�[��㵁�!:=!�d��VP��ԅ�b@yUgŸL8!�<j"]B��%.(���V�r�O|��&�	F~��$Z�}[TG?�CTN��yB� /gxV��Ԋ��قź�M��yr"�T���� �=4$`#Gԓ�y�B&`�^	�ɔ+mh|� ƨ�y©I7-�4��2�J>e�p�eO_��y�'�T)�ܒ!g8n�P�Uʌ��y��7X?�I�q#��`:�m���y2�޶Kth1B4#��R���1��&�yҫ֊g��yD�QL���͒��y2K�9,��90�'ʲO �ش/���y�	�e�Ɯ����A��̡g��$�yR�W/dY��r�f'+���h����ybς-W�X�!�
���&
W'�y2�͌Y�8R�E;Kh��%AJ�y�-X�)	�,��pd	)�D �y�#��1�|��/d�D�s΋��y
� ڝ{B�'Z����!4uj� c"Ot�0�hO�D�����*sp�X�"O�0��j��!D`#��Ζ7\��A�"O�}����n�q�b�)"�P�s"O���1�[6w�t�j�k��N_`z "O��KQe̲�X�#�)�,{�I�r"O��"�JGL���)(}cХ"O�4 ���@J�!�v(]�U�Xi�W"O�%A��ԧ^G�P#�GQ�nE"O�tZd/��8{�:Dq��˓"O�834�U>v����(SD�S"OIz�ˀ������,=څ�w"O2���,{��0�Ǚ% e��"O��b�E��q�v�֮R�B$yq"O��!��%��I���X�[�4��"OF� цܲTk�y���1��}��"O %�6mE�O>�d��fR�Q����"O<���2E���F�U�.�1"O����.�IK����/Yk�1;V"OR��%�:&tHgA;MnTp�"O��IDn�%2��� @�!n��y�"O����7,�F���4'��M� "O�}�g�M�$�9b�o�K�,U*�"Oq�p�o�Ya��>lx��w"O�p�ԧ1���z��r�#�"O*L�� ja� ��L����1u�!���/@18����(*�B�v�!�[�*�d=Cs(L) �|�##��7F!�D +u�#�Ǆ���}�C+�)�!�d��?d���u!��we�%��ǜh�!�.@��'�̐:U�a�C(]�N !�D��"%�K������0�cm���!�w 4�0	
X��$)�.ӀB�!�Ęnhr`Q*�A�H�k0�"�'�T��>�L}j�D�;k�,0��'�Y���1[��Q$@�[�ੑ�'!�t��Su�H��`i�"ծ��
�'��qKF�m%t�p����Դ�+
�'G��c�KB gL^ɁU��$_ˊ 
�'O�[�ݏ'$�,c�Rd��	�'���a�g�e�"Ms�"�$J�2	�'4�t��;i��i�C��2^0e@�'����/��|Yr�®'����'��80�Ƣ=:�iAF�q$�� �'�>���G� �q��E����'�\�猄3N� ��� jϪ�X�'2�$�vG֫D� ك�ܵ9}�Q��'\�Z��)S��=Y��Xh�:��'��T9p/U1�Tl����c�x��
�'�lȪ��J�`%$`���V�4 �'���bQ�Fmw���ν#J�$��'B�21(�T2������,�s�'������N��ÓM^�n]�)	�'�~�q�J�'R��hʒ#�T�����'����䭜�v�,y�
J�}Qy��'�B�(6Qx�f	9p-�'ڄ�"�ᕔ*��tI�X2����'�Ɛ����;����H�^�jȆ�UG�	1�Γc�9X��ާ5�,5��m��U�<M0.�P֩�:G�ʤ�ȓ��;�ƙ#��!�g�J�pF<%�ȓY{�1���]�_��e��H�D����j�ꖥ�B�@ЙR�E PI����)�g��.��ͩ��g�\y��S�? ��#���#��	a��/I�Th#"O�-��Ô#j �1�IFz�"O� 9fχ;k������i<LA��"O��bgL�_�n8����w�Z�!3"O���ޜ[����eC5�^�@�"O����M�Jl�cf%: &��!"O���b+B�U	,Hp7e�:���!�"O
de )j�NLb���rŸ��"O���ˌ4P�3͞5r[\�G"OH�IӃI�]C��U�s�J�"�"O���*�{�vcqjE��
��"O�1��.��Ȫ���A��TYY�"O2ՁgD�m����s�Nv���)"O0�#��So�T#��I$�>*"O�M�T@ϲc�JT  Η1�p��"O�5�QL����B��&�� �2"Op�X�N-��+��ĢI�i�"O����^<1�YxҪJ�d)À"O�Y�w���� ��dQ�	��"O���_(���̍a��8Ղ��I�!��G+
5$�B!#�X�P0%��gQ!�d@� k�	��b�a��h)�U�r;!򄌥	B ��QeX�l��x!L��8!���F�&=b�*��$c���ǚd0!���)�0Y���#Wzt�¢H~~!�DȺ$HP��
�h.�
�'\�	!���0J2TpC��U+ddȰ��\7�!�$	� L02�6���1 �;�!�dA�4h��9�YLt�z%I¶Y�!򄌿C�D��ɗ+ԌE�@GDf�!�Ę@vfX�I(C�޴YQd�E�!���G`�(3@������qʡu�!�L:W�V��qǓ2'�,���7#|!�DږT�^qTL��L���#O�{!��1�X$+��
J*a�3E�=q!�d[�pJ.)iWnٖW.Dh�K�jb!�d�3*�uQ�G]?@P�7�k��B�ɏZl�c@��nr8�M9�B�I=H�ʐbl�?4��QEP4ۘB䉟/��KF�ɾfix�B)�/=�hB�	l�H0���JY�7 �,OiC�
�֐Ѣ�C7Q�Z%�iN�&G�C䉎 �� DA�J[*�
���/�PC� Z���f���!:��h�@̇>C䉛[P�آ%'-c��Q��K�XC�	>�dS"�N�f�!v��9[XC�	�x�� Qh�*a^3� �)T�C�	�sN�珂> �<ձ�cɆU�XB�	�i��K%�<j�r�J6U�:B�	5v
:��C�&EaJ�A�ΗMsB�ɆNL�aE�oU^1��E�0��C�	<fH8ɀ�gO�g��}
w)
("$C�	�t<QAkS+H�(�����B�I:T,�2��>
�1c!͹_�2C�	�6��-i���7�n�
UC��#8B�	�th�t�6�-^��k��-��C䉈-�RW�R1(��+��;es�B䉼��xX(Z� ����"I%-DB�I�Y�Lx��
ʂ��e��=�B�I�~:�xu��=z�^����� PB�	�[
�@�%h��E�����#��r�PC�ɖ�,���K�-��9����}�LC䉩������s��3��a 4C�	X��s�C�kвd3˗:A,C�)� 8l�A�0iB�:W��N�N-�V"O���f��(C�1Q�̔�>�.| �"Od���Y8q��D���ٷu��"O�Q�ɖ� �"%a'/+$t`�"O��qD"[ wH�mr1@Ё�lP4"O��Ku���~�l���� 0���"O��V��n�܀JQ��HYv9�"O ���ʒ�<D�e9#A�{X^��"OZa0E�:S�Ny�GAҢ3U���"ON�����u�
dψ�Jp`�f�<�&�݃;D�)�v.��:5N���w�<i`ʋ-��t��"´c�Z�b"�r�<!&F��`�H4"��=R �@i�<QE�F�W� ����%�.* "�c�<i�l� ��<�!�U�'�D�h<D���s��/�,B��R�.V`qB�.D��@M�).%�'-݅6p�*ҍ,D�,s�hE�0�܌�a��X>x��G�&D��+��E�E�@�a��G��YҠ!D�P+�	ծ:�L��rCS�
[�qb�i+D�����Z4ͦ���ϴ�֩���(D��D��~�2P "B�/yU��+w�%D�����
3-~\,R!iɰ)�xm�#D��Zv'J�x�"��H3g�P͛�-D�\¶�Z/j��YDc��P�u�,D�X���ͲN8�4�����^FiZC�+D��2L�vࠈ��'�/x��A (D�ԛ� Z�r�~5ه��"G��ܙ�I&D���U��+��q�e���j^�Ȩr,1D���rϟ�Ҵ���#cG���H;D����Φ1Vf1���T�U��iyt�,D�Pk��֎4^�J!��_J����b*D�DzcMB3SD�%�� q��Y�d(D���@�D)o�$0B�Ν.tp��!D����L.0�ݛ�cM~�rf=D��f@�>A��;��Xdڞ�;��<D����C["�Py�Ē>$I�D`;D���@�A$���zG��$1}*����9D�0a���t|����?�-�pM4��-�O�|�4��ʙr$��]�,H)6"Or��í�t[�ՑbG��;q�m��"O�p`�cĀh�zw�P	X�0r�"Oh!�',T�5'�(Sv�V�XTpͨ�"O.�)�Mِ>y3��!N���"OإJA��:Mz���R\7"�R���"Op����Z/ f�aqC�"�By��"O9����z���"Ӻ&�VP�"O������s�hIq��K�a�1"O��ɳ��j�ا �9��U��"O^|B.�:�����QM�&"O��틢��ez��ѿH�}a�"OJjGG��S�⤟$L�@@�"O��$`�x��-R�A�1b�АU"Op9��U�8�P�1-�xYc"OD��v��!@�E2�>��a��"O~%���X�c���mU���`8�"O�C`̄�$����%	�g�4���"Ot��ȟ=XF����dJ[��8�"O���ƕc�v88!�cҒ0`�"O>�ku�y���6�:���+2"O68"�H�����!K=\�N�c"OFh�qI:2Ti�q�B�K���H�"O���*�>z�>MI���E�.�ۃ"O~��F^(
���A��y���"O� ��K�"G�lE� �x�Y!'"OH��"K2q�*��2IL�$�� "OF	��M0A�!KUh�[�0��c"Ot�J^�L~�� \�4/PR2"O���dO����c&֝1��H��"O���L�W�i��^�(�� �U"O<�Xt�>oŐ��B 3jȐīS"O^5�r��g���@2���.@u"O8��F
�8��.̵4�:0H�"O�Qj3��[h�r�U���8K�"O)s�D� AD�`m�y���"Obʣ,�*\)F-�D�[�:jRL��"O������i0�#g!�>FB�ä"O4�c@i��f>@�� ��"���Y�"O���F%ǧYŦ��I�X�8�x�"O�E��yFx������`�T��"OLA�`D�D�N�Q�/�����؇"O<�Sˋ�Fi��/^�ؠ�"O@j��>Q���Z��5v��Ā�"O�R�/V(]/�������^�ɂ"Oz�Rw�T�v�2ȉ�_x���`"O�Q�5,ַSZݑ��Usq�(S�"O$C�ҏ��TsA&�tZ�-�"O�m�����r�k3fR�xQ��ac"OvpX��]+����ӑm6p��"O �e��c$�a�@�V�-`U"Oک��D��)�t͚��ZE	�U)"O6K��C�����:&��1c"O@��H�ஸ��ǿ� �S�"O����P%y��ˆ,QY^��@"OD$0Fc�2;�<�T�өYY��8`"O221�]�T�i���-�^���"O�0��� ��sb*K�A�l� "O�dF7��y�t�ߥE�n���"O$���/Xe��)��1n� �C"On\��M�[SH�ۣIM�p�t���"O��8d�M�1�4	�3�\؎��"O��oJ�[-�$��h�,|�~� "O��Ǯ����y�!׌:�Pt0�"O��hF˛4�~�!�� .=m�MBw"O"��.�;/�L��K�7g8P��"OP�x`��ٔ��`[02��@"Oh��앚@CIiA
��aO�x0"O��Zr���sc�EK�i�� �|���"O���)9u2�� i�'`��@!"OHpq2� 88g�`.�l�<���"O6��,G�0�-A���.+"��"O�`��Y%�<򷏃�1�<U�!"Ox����M����P�XD�"OT�#��	�h��hwE)0���n�<����#��7%P�F�I��%Ig�<�����C��\rC,X�MZ�x� �Ja�<�BE��nRt�C6,��$�JZ�<�A���sX�K�AY[y<x��ɏK�<�A�/5h0�  �8e< &A�F�<!��E�8}���\�{�z-�@�x�<ɔ�|�(i�7,6^��K ��q�<A�c�%`�r�lԍ;��ţu��F�<�Si�Y��Q�'��r�0��D�<��J�G+�@"%�U�
Or��B�Wl�<�1��+^���$�
.P�&�p�̆Q�<���ո>��).t�1�3��]ٞ,�ȓ�b��F�[̌
S����Q�ȓA���@�	5;��*��^�%4��S�? r`JF�-MݠEc%���]��(�"O���s#�'�~�لk (g��U��"O����̞j${rK7]�vؤ"OxL3��P;'p�(�j׿���!"O8� A�)N���IFu�K�"O�$��Όh}6��xR���'"O�y�tOܒ{�l(aq�I14�pq�"O��@7�T2܅��W�$R�	�"O0����m��L�4��nxl×"O�Uqm��
�4]J�5q���z%"O��T�U iVpԒ��_�9���""Ob���.Ħ,�����N0v��!E"O�Q"��!BU�Y�2��
o��!s"O^a��_5c����C�kAj�j�"OΗ>Y �,"�W���ya��R�y�$��\����hk�aQ��
��y����4�+�%,�d}��J�y��Z�K����vÝ=.|@�B1n��yR]������ԥ\)\�%��y�%V�"�B��'��`�K�&
.�y�Q��~m��,�mZ�Arpd�*�y�FP9�#R�M ;-p���>�y�C�<��(��D3�|=If���y	S��������~~�PEoX��yB�ɣR�(L��CG�H��0Ơ�$�yŞ�D8�Q���̯J�6�1%�'�y��D���hTv n��W���y2�R71x�j���:Y�i:�g��y����rA�)Z�E߲PN(
���-�y2-�2�4Ź��U���ж�ˬ�y�,~I|�hc�}O,��3��yb��C�t�V�ܗ�\���[�yr	��-������](����-vh��'��5�v,H��1��)ǻW���'�|�)'�K�>��KSȀ4!�':��8���n�`�²�I!o�x��'�h�zT(|���H�o͋B�����'�d��e��_Z�a��3�6DH�'�4�v�LP�h��'�J���'��� �Mׂ.��|���x���'��H0��XB	r��Rfβ�ب��'~�7�2#� Y�gM� ���'��`�#��"	5�<R���c!�I��'|2�yԌ� f�T��kRUL$�P
�'�"�{��˯X���I׏["����'�ԥQd\�5�i[�GVQ���'�f p�(�)5���+Ԫ�c�` ��'�FT�S"�O���Ӄ܎	��ɉ�'mΔ�p�$.y̽�$G1�tb�'M
�{t�F�\����d�E�0$PK�'�.�x#��x5Rp0QL��M�'`H�M�~�!F*�����
�'�Zi��ٶW��Iˠ�S��ܸ	�'r��X�g>0���Ǫ�yx �I
�'��i��%Ԧ�@$��)��Y�	�'Jlx��OA�jF&@�"M�ֵ�	�'�8ѐMK�&��#^�����'��$���y-��E�
���'BXed�
!����OFmL�!	�'���LV��S�o��L���'#z� ��M�);0�Z�+&p3�'���'}�]I�nB<���a
�'B&����@�e�d`�$b�)z�fy�
�'~I��aQ�y��|��d���
��
��� �=8S��(Piv1XfH?m�<e�"O:a�F��!J�B�q�]ٺab�"O$R�`��bd^���\�z�iq"OДp�A�-��T3�gB��a�E�y�D�!$rV�Z�׍<�D�`�=�yI��_v!���67��Aeغ�yr�5!�Zq"��A*Q�$�d���yҤW�,�I��Ʌ,'���b�A/�y��2Hv��tK��%{@Y����y��#:����%�3mi�����yBE�O��YwI�')�=e�O�y��ެnt89'��&4����ԅ�yrl�����ϗ�h��!'"���yrZ�Q�*�kac��][��i.;�yb/�=vJ@�nO�f��\�`B��yb��38�A�bN׺d�P|�� �/�y2"�63�jAO��Y `��GK��y�J�7��Ћ�%��Ln�{ ���=��ycӾz�Ƅ၌E?FTܝ@���y�(�Aw����@*=˃����yb*C�����k4f��,!`�C��y���eE2 q"cڱ
T%K�/��0>H>	`意O��i��	=` e��V�<��&�7�V��� �3l4�:��N�<)5���j��s�����f�<�Tő��� �N~;ڤ0&B�m�<�J�<ExV�0��*.ې�����b�<F'��c��>p�L0)k�=��O���Q��?;(iye�RJO����{�����6m�+w�8e$���Y ����վ���g��TdA��`�����;?yK<�|J��+d��5v�	Th���_�0>�H>!�郯)Q�)˒%�)Nj�7JEU���_Y�c��� 6'���j#)o�&��@�&D���O8 �R$�1��AadK?�IQ���2��(0�[8)2�U{2�ӽU���>��d9}2I=w �I�6��\�4M(Ҩ�7�]�?�¸�����kɪ��t��_F���R�ɏ8���O��V��A�B�K��K�'4���� X{H�� ��#KP��
���O��'��K�J+r��� Q8w����'���DN�P@ �WH�"uU�y�,O6Մ���d���;!-CW��X����Q�<�=i�:b�0���]�~lp� ��+&�ćȓ2��䃑��P��(�I +*nn����V��o�EE��WO�CC���]�q��\*:1ʁb�NA�I栈�ȓ,�a�c��`�%k�������D~"D�p��VK��)�eDZ)�y2�)N�@ɵ)ԍU�hB��8��=�{�Í��r ���_+3njP�Dy��'J��$j?�eQ0fن]P K듴�I<urR�� ���FP�e��5�lB�I5^�����,���E��jB�	5%�^�0�,UU�ܴ�$a	�4C�	�;9��&�M㶜�w�#Ox���F{J~rg���d95&�1�#oOU�<�@9/�I���p~��H�W�<A��y&�0����aTx�R��Ux�<�Ʃ.2P�Ɗˉ ���Rlo�<�t�;d)t�j�	�x���ğV�<�@ ����3o��XB�T�<��I%t&l��>t� �;� G�d1�S�'R�d���6|�s��Q��$-��S�? ��#A�-_T��X��˦Yj̩s7�<lO�]�%K������~7��A"O�M�R�ܷP�6Y�` �V����"O8��&oP�F�֨c�G�L��#�'����D�C�B��Ѕ�6��S�+�9�!򤜔y�v��b�O)�Hz�	��o�!��ѬeL�3dO1йyֆ�8!�DN5�x�`�(�$J�R���:�=E��'۰��C���10�h�)�5Pu��'���iQ�Ӟ)�z����qڐ��'�5 ���?�d��K��m���@�yr�'��TDǶy��X��]��N��մ(�@��d��6KCp=11�ʿX!�dأ�xA� ������X�"��F��!udE�Fh	�vM��pL^3�yr���9{`&DX=�����'�yrJ:2��)�D�Ǎ]��l9�ʽ�M#�'�0C���h)lQ�sM��8�O��>y�{b(Xel�uU�{+�P[�m�(�y�L�]�% q
 bi��RE _��y́3 ����r��X˦A��D+��<i���'�b���nJ�L��`Q2<�n�I��D4O:�0�B��J�	:�A<^\6�@r���4�'$��s�¡�� ��G�����dpE��(t]!�*6ql�3�XT��}@�-Eay��I
�ʩ�5M�B ����6 h�C�0�J|:`	��0r�(ِ�nC�I�y)pP��L$b��A:3�ۘN����d!�kANp�%�#��Q�*��?���?�	ӓ��Y;G#*(di����'�dx�ȓ[���X���;�,aQǀՙS0��ȓs��-"%C�k�E)��o0��ȓ'm���'O�u5F�XF4ꂀ��\b`�����ԈCM-.�r!����K��7�(�а���E�l�"�[�<��+Y�UغH6���S��L�M�<i�f�2XW̠�gi��wtv����F�<	!WQ�`���I��G�C�<aS��pH5gH�)aW�ͣe�Ng�<)��=��YX��+F��!��,�f�<��hǌбLE�c��|�D��b�<A�P�9�{�<��;�"`�<�-S2|oސk�߆}T��CB��[�<�$ޠiB�qg��܃�KSx��Gx"+H�e�����zVx�q���yR��Ya��J���sY�Ӏ)H����O 7M2�)�'_��͓�&ȶLC���)��]��?���:��B8-�h����)�伇ȓX"��R��'A�@�G��:���ȓr�����H�i��irЁ�]�h�ȓT�2��тP9@�v:��Ia��l�ȓ�q���2��A�)X���)�����'m�s����@^��nU�>��s������� h��:����9��ȓ[e�e��� �`ΘHxK�'f�8u�Ȯ%3�*�@S�Rn
e�'��B4��$X��ʄ��Bj�< �O���dFS �M\{����'Q2	c��l��ħ�~b%C�l �;��7f��cOU��yr��-��� 6�MP�y���)�y2`ҷ�P�b�uo��;���y�ӭJoP�� (����d&A���O����n�n *K�W�J\ۢK��d�!�7ZQ�x �?C�H�Ag��x!�� �`�'�_�^	��WJ=;��p�u"O��`|BPSC�Q� ��t��"On����U2�n\��X�Y�J���"O�y�I�>[
3�#ߊh��\20"O��1��c����fm��I���cT"OzI�C)'Iz��5L��"��H`"O.�`��2\+H<4� �䌣5"O6�i,�� [��rp,�'q��}��$?�S�'nΌ㣭��<�T�bKW�v�T��ȓ9����%i�3;|�� o�1�X��>�����;�ʖ&�%��N�� ��P��y�h��"E����G�إc�/�qH<Ʉ!�\��b�^�Cg@����^yx��c"���  Q������@�Z�B!�d^��L�D�� ���a,W6t@!��U�7�j��6˞�e�1Ҵ+�|4!�Ǖ 7���'%D5"��؊��(	�!�d:��칖KQ3	���f��H�!���?y^`�`�@�NLD�S�b��u�!�R�%�� b3,A
c+�PI«O�T�!�D�=*p��$����#��+g�!�dU�O+Za['.��s�D(��ۍeE!���C�8}�u�T�Jߎ��D�7!�d��8㺍�$nԣC�$U8�j�%�!��R�T&U���E Jn�2�̉�+B!�D��OF�Ӧ.�6wY^a��L�4!��N�^��Es6��{V�ZgN��@�!��u{*���N�a��e�bN1/�!��9�.!�F��C2����T�2%!򤁤S}$p�u&E�U��.�"T��"O��c֊R�������0�(��G"O�us��Ii&����D�hYJ�"OJq���j~ B�O�L�P�ҷ"O������,]w�\�V5W��Yt"O2]P���	>H5�G���X�&��"O6�hq�K�b��'�3P�� �"Ox�"�@Y�J��q�>�\8�F"O�h#�U��\����#P��X��"Ol���b�N|X���=jr�U �"OH��4j�'wz�Qf�0y[NAp&"O�8�w&ei��J���8hZ�"O��"`�,��qxp �qپ|2"OH Q5��}�TՐ���y�Ɛ@V"Ot�{�(�%dڍC�!�6Pz�9��"O|�Җ�B�y`��aW��JUH,A"O ��$mʦ]�ˠ�K*#�Ҥ`�"Oh����>?���C�.W��e"O�Sc1ut�|�I�2�R\"O*��JO�v6�)�GY=Ȋ�Z"O���A%����lS�K��z��#"O&�)E%� �4�J�_�d�HP"O�� ��Y���'��)���z�"O�Ȁ���+ 4X�Q�L��\�C"O�!��DY�x:�<]���"O"��b H�{<j��dCң?;b�hr"O�ׯ.`_l���E$�9#�"O a+�\� >([F+A<.�� "OL�x����,�Fjw��M�:O��P0�i���	��w�R� F�	9nl,@�e� W]��❯T�6C�I�r X�	���,4K�i0f4BB�I�	�x���A�3P P�7d�-oQDB���uZ%�I-�JXd�& ��C��VV��!��Ⱦa� +3�ӳ�tC�I�<�E�����D ؀%�< ���� Pa�c��Ҳ���� �6�4���*Oh�xeA�G����œ1� }
�'~xl��'�5,upAbN�?N`e��'%���cۉ$��*`R����'n���ed֬Nx *P���w�� �
�'<ŀ��� 4i�a���Ul��M�	�'�� �ҵT�FTvoUH���'��3�
�SuV �U��
}����'n��,υUA���%ñlbq�	�',�U�gɳW-�[���"�f�0�'��=�լ �+lv��	¡$�,��'�60`��Q� �͚��@��'����fә%�H1��&�(S�q��'���yƆ�<fĩ1$�D b`1�'Fx"*��3uj�+2�hY!
�'%���_uFhyb��<��5�'ؾH�$*B�\�P��67�l���'t����
�N@x	�_�~>�	�'��� ��`������*s��-��'�4�q�FL�0�����C
EH
�'��xQ��Ӈ@���*�I��N"v�!�'�2B�P�Y�"i�d�´GB��s�'̰L1�
@��&`Jĭ8��]��'1��f�@�69��݈7��Z�'Ӧ���AY��9�FO]�(���'���P
�6�^rA�:
T��'�8y[P�
'����0�םg�Ђ
�'Jl1��7RL4)�R���"
�'c�)�F�6l��Y3�A�p,!�'	�a�%�;�� �fK�2Xh
�'�
��`��&|����ۆ	f }{
�'�$J���e�Јc3�Ez�����y���0~��Pc��Q��1h�yR�ŏ.V�"���N^<q�Ǩ�;�y���'��};��)�l�3w���yRĘ,�P%J�ϔ�+�f�B2���y�ۅ]�<Y��K T�R�耚�y�H�7�T��H�-Hp�f���y��G�Rvz���lN�\� �h̄�y��i ip��"�T ��&�yB���1?�����E qK5`��y�a�1L�$��� 1�z%Q�����yR��7An>��E��%ӄQ�ÅB��yb�I,qۺ��i':��9�(Ϙ�y*Y�"�9��* �Z�b  2�yB%�k���#�Q8�flQ֎��y�̖3��,�R(�	$;���c΁�y�L�d��
� 7k�P%�֫�ynB�4(��A:c���E#�y+أu����!t�,�D��y�#�3h���B��%�ְ2$�+�y���nTX,9W���'�`��D����y��i�4�$��3���d�܂�yrB_�T�n�c
 ��h�`@��y/)&�*"F��h4� �a��yr�\�v�5��b.��d�X�y"�
-�DC�B�j �u{dW�yi7)>� ��L�ge���S�0�y ɕ~�b�e^�\� ���y�(�<N�^HbE�E'Jv�}m��!�dP�!���V�w����@��
	�!��R����Q�Z�޸���
 �!�d��V A&o�!a�`ӆ��=a�~2ϘDH>�aU��p;��CW�K�F�l���[WL���S�? �U)��ATE�u�p��P�$Y���ɽ+�)��
�>j'?E���W+Ătb��_.�HѣJ"D� �d��3�T��F%�~���1f*�O�����lRL�ٷ��b� ��7,ǿP�nh
�	����́�Z��y"� ��ν+V�F�tJ�pcCʎ�cw0�gꜻcQd$d53��������K�	�9�,\�Ӂ� ���5F���1E�Z�EqO�L���Jcl^;DD�Ct��_v������_Âł�;A�2��5G�zX��(�zc�a��fЎZVZ�R�"?�fC�!����]k`�Z2��4Ь� È�.-)f��O	xġ���7��S�P��[	���c�`ǝH����Q�,T�>8��%O�|�~�*�j
�0`�"Ej�	P���Gl�/��"}Z�iW��[�`X$eV�b%�4!��È�D�?�H��G���OH���I��l$�$g�ŉ^�p�8���&bH u�L�ȱ��
���) �gH�M9BE�>V�Q��aB�.�p�d]!Sس�ڴJ�)�$>T*��E�!�DIt��Q�l��6c��N�6 �@}�8zE.V�>�Q	A�/)Jau,�Y�E��F�<�"ԐT������2Zf��I�)'Z!�lH�[�A+���ô�1uv|�Ȇb�(
r� �')r�B��>����� �L���ȅC\�4"as�ZX�~���L]Y4�}"��5�Y�5��|�O�x�o*=�6�Q`%N�hQ"�'+(���LCe�Qp�E��˝:*��T3�bVb��QĠV"s>�@�F�4A(R IU�ݟ@ vB'���kC��%�M5N���n�k`��R5D�[�(��$�՘\�u�v�+TB��'�IU�#�h���Aƥ��i�%^��Q�cԬQ`&��%��.Eµh>�O�c&�4�1�'ٜ7�⌈��'2lM1⬂vx��Y�n�	z��)K�C�%�>�!�'�4���'-��pcшT��r����Z?~d��	�]�x�5���/��t2O �E��C �8�͋�,�!�n�� ߦl0H���Y=��HE�45O4]Xf���Pk�X0'$�#�ʰy#�d_5gp@�0H �H����!�&�6�#���=T�5q$H	��A���<����e�D����7i�<����R!z�d��̍�Xe�u�f+�
X�"�O���|�0K��S�Ĕ���l�l�A�M�wQʈk��r���H�&�'����D݌u��Hp�HL>Z��dX�<�e%�@�ăe��#�Ý�v��\h6�h��xQ��iƕbs��뢤L̈͐r
��p>)J)Uz\�ɣol$��άv.\� ��
g�#on((�A�-	s$H�0���?E���J�Hhq�X<�l9��*�:wy��c��E"��Q�b�BJ�0:��t:�'���S��Rގ�	G��q�'��ܘ��!T�T8#s)� ��u���U��
����Ƹ6�q����(;�RY���:�ܛ�+�L���J*0I٦l4�P�\1gE:��)6<���ɞ�W�x) �(�%e�*C�I�!\��	�L�N?2����O%�"C�	*(`9B2	�^�$�!��^B�	�;P��ɸ����h���C�	�y9.\(�� B��K���&/���Ē @��CK<�Q���UDn���b�6T�t�aSB�]�<�F+̯�@�d�.	J�#��Y�MY�2��s�)��*v��DC�+1����H*��C�6`L�1�&|�d��%�_s�q�!�$}2E� ���}&�����]�\q|!�ũ��/��=�pC���'�&���D�N�^�q�ւ7�n�!j�]=a~���00y�AÉ�;+��J҄U��p<��%>�p�k)?���RmҐ��9u �ãk	T�<�!٣u����f�;>:nukƮi�č�tvl��vl �0|�/��P��r瀵5���0J�f�<�5c��C��ay����;�p��/�\4��*�[� ���_�Bvq��'`�pAE�#0]<�h5fĵQ(���'w���E?*�ib$�� .���45V�����'D ����%V��i�1Ȉ;s�2�S"M��x���! �V�a,
岁�v���G^%�x)PU��|�z��Eh2D�́�c����f

HZ�K�o-�L���7f^�=x�G�D�F�s̀�%���
H������y"�O�j�V����*��M�W/�,����������޽yb��?�'�-s�MZ!/�*�2eF��~��
�'SN�n�.}���I���y"2�N��촁�	���0>DA��	���+Pj����]���L���2Q,ƺ~vy�%3OB�@E&�-
�P��@$l����"O�,��O"�8"��p��$����^9u`��*�	����� �u戗;���:S�ˏ<֜�xF"O~c�"W�8I�� ��a�/13Af5b��>�H?�gyME�,�La+W��8�%�Q�ybB�^%ɶ�#1=����@U��Mc�@K"&ܾ�p�Y�tA��ڧJJ��:���v�$�Xj(xGP�TQ .�a��a��W<*C��[\!���0Y�0�ҵ�T"w���׉�K�!��B ����"c���b�EȞL�!�d�`���A��>c2����E�'�!� 	^���Sm�t���Û�t�!��F�PD��Q�ǒ'����DI�!��8 L�Pc�"|��a��N7�!��EqD��F�$~4rD�V�!�����YoI�>��r�+c�!�K�u��h�Ќ|�q���L}!���c�d[M��|S�)6!�^�u[�bT�+\�`�2"�j*!�d (Jz��ْ�T= `xM��L8x-!�Dʏe�.�)TFë6	,�s [0!�ĉ&XDf�{s!�'9�(<@)Y�L}!��K�y�d<�T�Q=|��ˣi�{!�D��	g&a�/��U����(Y[J!���$=m���7���j�a/o�!��K�lf���&� $�=x��_�Z�!��p˞ �$k�l���q��� �!�մ_�꼛㣍m�x��E�&�!��h ���F��x�x����V�>!�dN�C3>��É�h��dq�dw!�$	u!��q��z/�9��"�.�!���_q� A�'�D#Ea�FZ�R�!�D�70 ��h���?)6��[sD!�dX�$��A�Ɔ��s���+.2!���:v��%i͐�H��#<A=!�U���p7�_8G8	!d1M?!�M�	�f�9�l̈B����
��z�!��Z'8�!o�\�21r�H��T�!�B�`�\90�'K&��	��B�j�!�d����-��nʄ����Y &G!���<0�b�pa�9W� ���%^�h?!�d|��}`t�C�4�T5ɀ��A@!�d����PPT��)|&�z���h�!��I�w{����U�\l��\<�!�$J6��}H��UT�t�!�B۝E&!�$�$h|r��D0Fm��')]�!��/A���'�̎F/�P�Gʺf�!��@:�A�jػ@~�lp�R��!�d�/��z"�V N�<��1�֫F�!��-<Z��A�[�*��!�@��#b!�d\�)�ʘBB)F�f��P���P�:h!�D�ou���#�u����#_�yA!�$��P.���`���V����C��K�!򤓂9�.|�%�-N��ss(N�p�!�$�,_pZ	䉊�l�}��h��!�D�I���+ҢZ�j�.U׆�;t�!�ǅX�3�lȍ&����T�v!�J6=LaE� �&�4mp�o��D!�D�(yh�����<��=x�臭,!��\�����+	�w����F��+d�!򤎼:�A�PbZ=B�v�ZE�
0!�D�o��R�r��IFe?!�dП�| �OF�iunq�f��'m)!�G���@��H�,H�Y�bA'M!�	&V{L�9֏�:C:�����!�D�
@�ҎʈVG�6BW'F�!�� .M9p����޵hH¬-Ϡ�Д"O�m!Ň+LȐ��n3t��4	C"O
9 b�*v �#�+W�y*���"O,���&���`�9Z���"O����89��L�v)ǎ7�(��"O��t�L(��3%��RVKr"O&I;P��\���$��!��av"OL}xb�*A��s㘅tp|�"O�IR խw����5ቺs���0"O��3d��m��ѓ�� o��5"O�R��˭p4��#i˸s����"O��zG�άDϺ�r��J�e��T�"O��s�ϥ`�< f��UΤ��A"O���Tf����T�T�E�u�d��"O<$�Z;u��y���)�4���"Od}��M�^d��_�r`�@JD"O�a�g� p�Jܣ�,O*��z�"O�\2Bڞj��z��ܑ@�|k3"O~h
���U����<a�:�"O�����}���S5�P�^��B"OB4�M:}[>��L���l
R"O}���>�K!k6_�����"O��[2
.OÈ�����l��TK�"O�Q ��!�"����ʿZ'j��"OF-(QI�G�`5MH/#�5�"Oܨ�4F� )�=�1��C���#"O��j�9nD����.j��E�1"O�8��]52�z]�`��;�~�h"O��(�/h�=���N�:-y�"O���"Q�6����@�K�TES"O!�Ɖ�i�����jB�!r���"O2�3��W�9�삐�Ȇn��iZ�"O�y���N��$Ȃ�� �N��-j�"O\���&� J�Hi�᧞��iQ"O��7$
�.�N�($�!�pta�"O��0�O�w�(�D�ϣ	\rM��"O�5��	@P�tjٗC�:]�s"O��s�̭'���K�# G�E�E"Ot�+��p��A���?=32Y�C"O\M�%�w����lĊe5r`I�"Ojps������W,�.����"O��� �XM���KҰ�YV"O@�q��k@�h#@����C"O@̢cʀ�\k�t��J�&!�0�"O y�֣Y�P�t�[ �A8Rw��"Ov��@�(YQ�y�H�{j^%W"O�����p��q�F�CN��"OB���H/H�%£&E%z#¡�"O@���m�u�4����Q�B��2"O�˦'	R��Y1&���"Of�����%4�L�f��,\j��T"O�@3��˸r�������TJf��"O�)
���O��@TC2�=�"O:��q�,A�0��N	�!27"O�����S�8RU ��z�j-�5"O"���鍌bݴ�� %M���r"O�$h���+"�B�,x�C�"OpբbJ�?���㇩ʢo�x"OV���@5�T;ANZ�g�����"O��S��o�����'h���j�"OD�k�7Ll��T���[�X���"O.�+�k�&~E��9�B[e����"O���@�#G�a�'���Bv���"O�|�#�=Vx$��$OR�j�����"O� ��S��W?k`��v�4�����"O���0��%�����%_&Z��i�3"O�M�%M�u��d�ģ�=<}�Qy1�'UZă!�7��1B� �DD��/ly�ii�J�]<���Зa��CU��E�&��d*Fy�'v	�b,�0{�������N�+��,����n�th�d��y�Ə�I�]��f�.b	8�@�)�?��Q$j8��`ӊ6�fX��i�42:�11H�%g�d��P-�)}�"C䉈^!�ѩA�@��H�9�G�K
Μ�U"_ݦ(S��+1̀ȸ�I@X���d��?<�PG���}�BC $!���;�-�{J|b����O��9Ф�6,�hy�iS�m@���X��C$P�/�faرI3�O"�h�mz((A��J�(B��՘�T@��YPU�l�#
6NXy��D�ۢ����$a>����*_�<�xu*0�k�������i��P*��ζi�x8{0史$�bI*$�,܀d����2Y�+���J�!�b�7訟x0)��V�e�%K �׸pP� 2ړIH�A�u%Ex�b?�y�����Q�w#F���iU S�qg~���m�|?v|@@쌟S*�g�'G T�q�"E�$9kP��!%"Q�s$���2t�1L�S�!'(I����*�0"�Ԁc��	'ƕ"���	%�V%af-�O|LaWƍ��ݸ�*��
Kxyw9O�00���\h��$�������;5T��tAIo�t� �;���x����$aė���=�a�!Ar��H�58���K�$��|�!� Ѷy�*�O6@Q��N�`:�g��u�#�U ��`�A	I r�*�[��[p��}��X[fk�^	�b�2��0�����áv����Zޞ))[��'hhS��ԩdf]�G�����٨&�|��įIl�%�I�z��b�'��>�ɮ>��8 ��JXH��s!ɶ�"��c����"�0ɛ /��/��!3���+���S���)��i[3!x���)��,5�ĔA&�PCBO�c��{BB�4!�,h`6J�)��P��F#Oc.�Ă�:1���"O��c$GÝ��ѻ�n�>�>4�B��چ%S!G����H��0�d!�*4���B�,~��c2"O��� ϖZ��u���� L`��_��bՑuKg��-�g?�թ .yR���{{�2�_�<��@�Rv-��˺w�>\hbd��<!E'�\���s�i��bcl�*1]� ��)h�����I����R7Of���	�|�@a��I��U��q�"O��⤦E�
$�W�P>�Y"��y��
�g�:d��'�@4H1��m�-�y2+ʆ ��P��8��M��ȓ�Ny�._�L�$�yA���̘��r�f�`A�mZ��Q�ۂ0q���
lhc��M�ta!�@ɾFM���|�� �] i����(�>,��y��HI��ِ���uT�a Y�/D@��ȓ'�"��rlR��t)@Ƈi����ȓl����5�Ϟ8C��hBa��h8�牞9A��xR�x�+� #h�iR����ȃ��yr/�+~A Fl�$z�v���
�ēI�����K����S�z�J����g#�}�B��p؁�ȓʜ���1�T%�4��v�.\9��I�DP��A���L>�Uw��"��1]]Tu�_}(<���H�a&~1�0'��%�L�J1�$D��IƢ�w���ݯf���jE(�.���[1ܗ,s�x�ՠ	z�<��ED~�#��y��rPcP1���!���y�ե9>(*��І]���FT3��I!�$Z��L)dna�4NQ<d*H��K){�&�T��?�yb��%T�$���	�i����CV�@\HR�h�<q¯�_�>�O�D�geMC�����H�ABPz�
O&ტ��o�ȝ1񀐶Z�<�)�$�Arh���L��m��ɝn��ؐOӑm�$e	c�i���DþOA�}���L$}^�ɛ'x����)�1Ө`���ij�yH�'����w�^0B,��� V+j� 0�J<9��A-T��)06��;8�?!��_"���ht�v�I5,,D�hQ��@�FQ����({t|h���2u9T/�<���	�����	n�ٲ3�	!�i�B�NޘB�)� $�A@���*��c�57i�тvE0�	��S>�a|�CӂG�<�8��՜s.l��7i��p=ie	��e"T�k�|1 )��8Wt�K��Q�\)�Q;�(&D��A��8^謈&��!t{���D�+?�p`�S�#g�?���ÐX�p���ͻ��E�+<D��1t꜔�je��%\��H�bٚ@��QA��6}��s���d�f�D�R��z0�aY��Պu�!�d�RԢ��ň� =��A�d��V�Z2���'yޝZTj
�~�с�(����Zߓ8���8���>9_(&U�C�5@ oC%Lĝ��D�z=��lG��\A� �=�V�ȓ(��Bc�=qA�@��O�a�����:�ˉ>	�H��H�*q ���&�aT��y�*u��/�%@F�1��x��%q�OP�/�Y�� ��ȓTA���f)��
8�I�W��W�4���)q ���I�4�Μ��	ݭ)2�Ćȓ	pF��f��"Yf��{��M$"'���ȓX�~������8����Y�\,6$��MR��0"ȼA�����(NɄ�I��4{Bm�d�T�3��ՓO谄ȓv��\i"E�F�ԸK�G�kD���ȓ]q��S�障=��%�*EPf݄�o�8thoL�*`*iP�B��������À�YN�H��.�Q>�=��qǶ�ȓ��%�9�'EÕb1���Y@��eʫG���J��_ɨ݅�B����ʴft�qF��\9��P�޽�C(ZXzA�L �E]�8�ȓY�d��E�!�R���U/#,Y�ȓar\�1!�M �:3�ѷZ&���ob��Cɚ8p@��b	�BB���ȓN����]�8xC��֠2V8m�ȓ~�*9������kA�\�j��`���>�Z�-8v�
C �/�����4Y��N����T:�#N�����M���f�r��wx�Ņ�Hm�%�Hq���ZG�ϛ �DQ�ȓL6)J4� �uO���W�ܫ���ȓ\6�HXe���Xc%���"���ȓGĆ�;�kK�:��a�CǶ!���l ��
YT�P83��מ]h��ȓX�j�j&���Jv��7B�q{Z�ȓ-<�x�/��	zLu����o��a��T_��A`H�&.�7�_�#�f)��O�v����V��jb���I����ȓ_א�Ked�	V����	�(n��L��o��m�`�=$�*T�>a���ȓw����1�A*y��i�7�B��p��ȓ?�r�����os���-]W8��ȓy����Eܨ|"x9  �3Ip�Ȇȓ%�֨9�^'A�j���#_�c�dцȓ0�4)HAi�$tX�cQ�Pn����;&�� ��-$r�Q+�~��{�h���M�N]j��!��'��U�ȓl�Ȩ���ٓv�6�Ӗ�Q;G����Hy�[�J�qI�L3*��ȓQ<�Y��#z�P�Bt�E�ug(`�ȓ_�p -��	lH���c����g@,�b�����(�h��1�ji�ȓ\���
FN�W|�ũ�+�?3<ąȓZj@ah%n�*��M�Ub����ȓY��pa� 	f��pM׷6G��ȓu'��� ��vmx$���;�t���S�? tx[4)� B���!�=O���+"OP��)7Ha������d�be�R<O�L��F�+lt�3&ʗ�*�l�r�	p����5+��#�,1A�%)��B�I	��R3��@���Ưm0B��0NE]�4�ٮcm��F�D�&Y B䉷#��� tO����Yy�m���C䉆s��rR�S�Qn��r �� C�I)n��h��,�X%�$c��g��B�	i�h�`��lN4"��.tKdB��;!gHTy��GF�:�XA�Vw���	jx��?E�T�wJX��j6lk����*@V(8q���Hܓ��I#ʧ/f��5N�nޜy0�Y�y���r��^�	 y����ӂ� 5I��$�����TAI>y��G
�PI	ç]���"�J�+ P��@�Q���'%�H�bK� ���Ո��=91����[Cb¬w��T����r| �A;5%��7�0|ze�xf\="p��E?X�ƍ+wQt��w�c?����5o�����4��32"����	¹�NB3K2��6�  ��i�]��^>M#�i�t���[�Dn�\XƑ���I��^u�Ԅ�0��ަ�yçK�\�����
��q�����I:Ψ��ρۦ]�2�iza�4��<@*Wh��7'�]��`�9�~���#!�M{���>+>�1�O���J�F�(# m����z�����)�Mu$� � ��e"�a���z���b�P��U�Pl
��M[R�=5Y���J�;J�I���s�:��;"i���hT�ra:Ն�Ty�*�f_�x�4%HW�<I��Pm�J��	��5�3 ٚ�������"]� ��8�7��"4~tY��d>���.Bl�T���h�����fR�l�06��J����߷1��HF�,OHi��l�2���$F�i��P��i��i�B��"�ƌ�O?7I,
��͡$EޤC��rK��c!򤟋=�d��Go^0yȖ�$וUI!�D#`�L�5
�FP�<�Dc�0ld!�&[�(yX��[�GhTD9�#S�bc!�Y&�8���+�)ZX��p�^�Z^!��
���р�ѫe4x��䏭iY!�L9>���V�x`�)��i�!�D[�6^b4 �瓗YLX�`$� �!��Cǐ�#v,G`�:�]7g!�%�"�*ë�"��#�/͑�!�dE�zۖ�����b��$MpN!�$%L��Ѡ�Ŗf�I�Tnҁu]!��ű>Ң,!rd�!X}ꠊ�DJ!�տ1� �+�U�q�fI��hB!�$B�V���1���BЎ��­ǐ>-!�$I
Q���q�/�/��$��M#w�!��T��,ф*� ����-��u�!�&�ic��L�p�dC�{�!�d]1*�>M�ՍumFdɥ$ǻ�Py"cN��)8�eW�2'���j�y�@Q6P���,�z�P�gÅ�y⡒8��F0p���W��y��	�x|�"ٶ���
��yr$�-? 2� '��, ��B����yBAǫ�Rc
��t��Y������y�c��n�h�*��]�j^�Ɂ'�y�K�DR%DN��������>�y��1V1��i׈���@�Ѷ���y�BZ/1Y��A�Z�^�P�/P��y�䞫N@y�#�OS��q`u�
��y�\�r�ΔA�� ���gJ��yr�W�0rθ���зcC�]�&攢�yb�V�IX��۵%�[~	ӕ��y��^$@\ (����C�4�B�Ⱦ�y�_�8�isdPH�|��(��y�儀p�DA���38�`��1�(�y��4\<Q��̰)��s�⛠�y"	ݎ������0����p�F��y
� �LB�cŤbg~!rFSA
j�z�"ON����3!"�ř��nh�6"O8�P�Qf�b����0R�EKW"O�� +J�s\Lm`�-ȷZ@���"ORu�6M>O�a�+֯A?Ɛ[�"O�m�"/�?#v4��Q�M�M'n�C"ON��w@F�b�Reb��˷��hW"OD�� ���z�j��v�\Z���"O�����](i�* ���E\�)��"O8P�CJ�2�XdS���>��%s"O
�j@�A�X ��#�R>,�2	�G"Ou3�D_����ȍ8�2�x�"O�9�u�*LN�ي���42�(e��"O����<*ќ���ċ��V��"ORM����O(^���0�NI2�"O�[Q%�r����R���^�����"Op!x �qn���T�d��%�3"O
UK /J$V6b���	#�y�"O �b)F�0:
-*�Ú�F��� "O2�HQIG&?~q�2 �>�S�"O����+P�^�`������z �c"OJ`���#�"�n���0x�3�=D�c��U������z�P�'D����dT>G�q�P��)�0�G1D�Ly�(��dR��
�-=�=��E-D�L�C���H���bGY19r���j7D�$��.L�\	Ir�
��qW@yZv0D���� t�yP� [�,�q6@3D�8hC&��}��}�v�˽{����o/D��9E(F�cdF�j��
��`�&0D�L13Ϛ9Vp:X���C&U�j�b6�-D�`��N��k�T�e��oyp��(D��0%�R����6K �It��U	 D�i��I�(�
l!RÑ��3�0D�� s�s��ĩ�B_��9�/D�TJ�bͻ4��`�ebP�|�XaE*O��!@��5
�9�(�R��q!v"Oȁ�u���3
�@tFJ4�T�s2"OF�b�E)SnY;��ڂ;�R�A�"Oz �� �.Ql���n.S� xh�"O��bp,W�6�1Ѝ�:Wͮ5*�"OZ�(tȁ'N푆"�(�>�KW"OH��'@�5h���'�g`�{"On�i2Ă�7䙹�l�����@"O�l��,�K���c��ԋ:�a��"O< ��dֺ'�H�+S�҇��s�"O�R�IZ�t�z��ȣp<����"OR�z�)�۶�&��}8�� �"O��v�aC*�r!,��Z���"OH���c�|r�t���Z,B���"Of���]�}� ���iO�y�� ��"O�n��l��ĵA�(T��"O�}�6k �8�]�G�V
A��"O��Ӓj��[��xW�A�����"O������SԚ�i� ҔZK�!�"OPi��䄉<H���`́\Ԟm@�"O 0Ѕ�0*���6L�	z�-Ie"O�3V₀A�����M�D����"O�A�£�~պգ��A$@|5p0"Or�v�5h:�	У!�0Uj�]��"O<�`$���vzj��!�ʜ��QE"O<@��eD:%}��1QO������"O60rdHQ=2���0h�>$�f"OV�薇]2c��p����9��"O� ��%�����e)c+ԍv�$5�"Odr⡈8
g��1j��s�pi�"OẂ�xe���h�t��"O����@�$��K�R0���"O:���.�y��qq4DýV�9Q"O(\���%=�}y��Û	����"O��q��C�ɸo۞|���'�t)Db�i�Xq��(L7n
4a;�'Ӷ%�bE��W�q��(�lO╈�'�BXШ�2	�a�P�Y]=f0��'�)*ծG�G^�,5�K�[����'�d��ʜ�bpeЄQ�T@$�`�'9`+!ϑ�tEb��9T�r�c�'�� :b'W_����@�x��h�'����
&�����<0� ��'	r�3� ��#s��@F��:e��')�����
�eq�&ۥH�*qr�'](*���>	CMX��ݛ-B��
�'����&S�0�ct��-;I���
�'���¤H��T+l��S�:�x"�'���z�@8D�J��3���]��:�'�a��[?�fl@S&i�Pi[�';�J��5a�m8�)�,�Q��'���F�i%���3��+$�:�'�$ [�aG�W���Tb5*�Ƙr�'�Ni��+T#]�qATȐ�Y�lQ�'����n��C��0VmA�'Ǵ�˲��0aFp�Ue��)(�'b��놭$w�	��I/
^H@{�'�H�s�\�JvN���!A��I�'�8}���jMl}s4O<�ԍ��':}�C�����9c��
u��'*8�O�x�dpү�<3�����'�P�+2���f]AE���t����'���{��5	A��IՃD�dz\���'3�T�0�B
M���i��P�X�����'{��P��BN��]:sG�0�'�Lx�/�W� �HuE۳"w��@�'����R(�a��`B ��i:�'Z�8`A��$�.Y���,��'l��h\�V���Ӷ艠l�A��'*��
\�~��&�H�U��'\t �ɟ���(��F
��L�A�'ҤY�̄�:� C%Nӛ{�L
�'28���΀L�Xj�
�4z�"S�'�Мd�J"��!�ז��i��'!��u�ɫg�Ɓ���$��'ٖa�����B�|$���y�'n�`�녤#/�]0UL�76!��'d��T�^`k�&�}:%1�'�|���L�+��"sI�r=Fs�'C&���!�������E)_�i�'Xj��3Ñ�:	#q�S!J���'�r} ��I2���)�$E�;�*P��';>��p���ZL��(��4���	�''p��OV#Xq��j$&N
;;��#�'�t]�!��@���9�e؁72�'�x�B�D��HbPHč),�*�'9�j$GI	W�
��d�ݎ �d���'�ҁ�C�O�3(�D�T���6"5��'�	�W�"��VF�=�0l�׈"D��c�*��u��H�&?:т� D�t�dN��(����r�M�d�F"4D�����za)�d�v�F# ��y
� ���J�Q�vԻS�L�;fH�t"O��b���:rIJ�OA����"O� gցv�0���'O�(���`�"Otɳ�Θ`
'ԉ^�p�V"O�P���ՊeE�@��B�̸��"O��3�̄�q�x�,P$��A��"ORTpd�K*��ɳ�(^���"OP1�s�l��)�%�1_�:Y�"O��)!�W�!V��5
Qu� �y�"O�)��jB_#�)*�I_9ՂI�"OL ���-�:hs�R�o눸 "O,M���S@2D;R M=8y�˲"O���!aI�'ö,���s4�Y�"O ih���~r��#@�|zj�I"OV����$+�0x�LJ�.Aj��6"OXL+SJU�ʍ��kϽH7�a�a"OR���gWt�Z�W����R5"O�T�2h��iR]��H8ߊa��"OZ�H�'��]`R!PC���	vZd�A"O���GӃ^�|�FT�;�p�s"O�p ��d�.Q�v��Sc.�1"Oz)A��<p�B�X���A<|)+�"ON���-I��z��9tjTç"O�#ҡ�+�Ƞ��O�
���"O���'�R0�g��7�r$"O���+2@�"@���@O2!�A�!-�| �)��O�����M-.;!򤏁��M�q�Y7H~���Z��!��WCi�*��{k���4�;!�DAܴ�لF�Gcr���댝`�!�$����Ư W�]Ybi�7f!򄈈'� `  ��     P  �  �  j*  6  oA  �L  KX  �c  �n  iz  ��  0�  E�  ��  =�  D�  ��  ��  &�  k�  ��  ��  X�  ��  >�  ��  L�  � (
 � � % f# K* h1 �7 1@ OK �Q Z d �j �q �w +~ �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&��E����8�8��͜"U�^�p"�ߓS�!�d߅X����%.ͼ2�EO	n!�� D���f��Ik���!ڨ$I����
O�6�L)n4\Tb���>5����� M�!���r��� �� �6<r&��/C�ax�� ғV�1q-i����
"�F̅�xl�X`��+D�ez��%� ��\uj�0��R>ܲ%`��T�ȓ%z�d��� �l���;�.N:d�!��_}��i�铬�O$�����%�tm�P��3�<�9p�'$
��,������/"��( @_�EZ��p?y��g0�@җ�L�Xw2)��@�'P�}�uBC�ai}1.I^Ȓ���&�v�<لBޥ9�����d�U��0�cLLy"�)ʧD~R�W-M�|E���P�ÁST2؄�?�V-���d�����=f�05�ȓ`�ꕉa. N�И���,eL��Q��=(#�UX��|��.ýN�Q�ȓ1���vh�9��R7C�7���ȓ0��	�kS\58�qr��*����y�nU9��ٷ%@�g�j�� �ȓy0��&�C�cja*�ɜ-w�
���W}V��K�:�qi�X-+����ȓx6Н"tLt�r4� �_!S���%��!��	�_Pq�'���x⥇�z�`���F$m�,�:�!�(T�ȓ+d�a��ڀ�XQZ"L$$}�ȓ[�P�Q@�>�fM�h�c��h�������ɓjfD��3�??���b�L�e�
*��@���1&�Y�ȓu�\i��K�c,���ɏ>��̆ȓmv=Z�'��CWx�1�����5�ȓK'�� P�yN��WɉQmj݄ȓb�ƥ2ڟg�a񃊑+y����E��B�X�`��i��h]>�ԅȓm��́��:("ĉ�gvͅ�e2�q�
*Y�P+t�&�Nلȓ�F˖�]6AI�,[@� =o*Ȅ�b��|�1�р]���:CCS.TRT�ȓ�GϘ�1 ����l�(LjB��ȓ9�^��&"�$|.)��J�wN��:M��vHP&%z��b@%g���-z�!�7;L��7�����ȓ^��x��iI[�4	7o���x��i�!sA"� F^<�R$��	�q��0�yb� �Qi(P��	)j����jR� �uk�$�$�����j�p�ȓ=g�`7˛D�`��+ɨD*��ȓ�p�R�]�
>^������h�ȓ"�������\gـ�kQ�@T��De
��t�@$�� �,�e��=�r�3BΏ{ DIHF�ԌM�^ąȓg>x��e�hF<�m�`Mz�ȓkڸ�iӇN�R��@���yF5��"���ł!n&5�KՆ��ȓ�����G�1Y<�r4�Ŀ	'��������p/҄"� ��Z�< ��ȓ�Q�IWL���2чF8�Z��q���K�	J}�܋�ɓ	A����u����wP�|>h�#�G��x|�̄ȓL�̠�Ve�]��l��K&cD��ȓB�v��nӝd����ҡTh��ȓp"�Y3�Ϲ7�``���5����ȓH&�%H2�@�f�@ (Vc�:o���ȓYj��p�،=��-�%AƭJ�l��ȓNH0�
��"[~�x5*M4NB4��S�? ���09�45p!�Ђ�=��"OV͓&��!]>�j3��E���S"O�q� f�1&aL�Xb*͹	���H�"OH|P0ßb �9q�dhʤ�"O��S����@��B��:�f�'�b�'���'B�'���'XB�'�xH7H�3'HZ����N�0̺����'�R�'���'���'^��'�b�'������&@�1�aDA�V�#�'G��'}�'�"�'v�'���'IXݣ`�;48~�Hg�i�eq�'�R�'"�'���'.�'���'��	t��w�(��B�+b9�W�'HR�'���'���'~��'!��'F��Q�˥R�\��F�H����v�'�b�'���'P"�'�b�'���'�L:�#L����MB:p�0���'�r�'�R�'���'���'*��'`��r֥�Q�r��φc�d�t�'B�'z2�'�r�'�r�'�r�'�����uM���C&K�_�����'v�'�b�'�2�'�"�'�r�'x�<��B$1��Y���%a�|��!�'22�'���'���'b�'I��'�&8���<�.���eϫO*���s�'��'XB�'��'��'�r�'�<DR��9��h�� �����'�2�'�B�'��'��'���'�P�rr�;�MZBn^�y}Ju�4��O����O��O����Ol��	㦕�I˟hz�	̍Y�LP���l�h�W	��d�O4�S�g~Ҭz���!7�R�f f<Bl�/#4�a����BB�I��M���y��'= x�O^�M�����U<D���'�"�������'1r�D�~�%T�zP�!1u�h܎��b�\{��?�*O�}ڐ1�\$��LA*z�h�%U�,��6��Ę'�|mz��J.A^e�DC�"��p��ó���D�	�<�O1���ZT(Ӝ扆��JBH�M�F����ކ!�d�I�<�4�'K�iD{�O� É�JS�藲P3h51wHɌ�yr\��$�Z�4mOV��<���R�c�P�E���H2A��'c(��?���ybQ�$c)S�J�6=" �ҷ$P)hD�&?��A�\œШģA�^��'�?D�O�Z���ʁ$RFxsE%�
���<y�S��y򢗯Iu����a�E���3��۪�yb�sӘ�۰���ݴ����DNˑ<�1* a�F.�h���y��'R2�'�()�ѿi����|Z`�OF��Yd��9���B&M����1�ݟ�'W�i>}������	П@�		)���GIR/O�d�U�f&P��'s 6-�j�����O���矲�	�O���N1�DM�s>�|�D�߼VL��'
J7͗צ���)�H����1�S��a�6@�6L ��F���`Ա����eM͠	�Kr�I`y�L��U4ǎ�6���Aj�(>tu������	����i>��'��6���h��'�hA)��N< �`��#� ��85�'��6�<�	5����O�$�OBE�'��1N���je�+��[�(�,l46-$?��oբZ����K�������lף<e� ��"ΐ�6��`�p�8�IşH������D�b2EM�a���	�h�0�2dl �?����?�D�i�(	�O?r�s�$�OV���(�H�22��v�f��$%���Of�4�z
��c����h4� �����a�㭍�63D�Ivl����N�ICy��'<��'\�k�NX�<��7*����L!$���'X�I&�M+�AM'�?���?�.��-h��Zq��i�$ǱBq	�P��|ѫO�$�Ox�O��N:�h���H��bK�J�꤇N>x��o���4�����'��'��+�ᑠ5ά� s�ף*ؾ��'W��'HB���O�	,�M��GP8 �� OL��iQ�I;W�d�#���?���i��O*��'.7�	:<w&4�g3�]��ㄛ���oZ$�M�u���M��O*	X2D������<��.�9B>p(7k�4T�6&Q�<,O����O*�d�O\�D�O:�'K��d�0��Y�A�eO�)� t�v�i""�)s[�x�	e��<���w9��kG͔�{���q��i��1�KmӨ�nZ��Ş`�rݴ�yBhFv���2����P���_�y���s6��I/e�'2�	ٟp�I>��1Y���8�@H8!>lx�	՟,��՟��'J7팰G}����O��D<�X"�_E�D}HD�!7r�ګO�Qlڟ�M�x���Ff��T�:Q(�W�Y���$�st��xQ�3r�"����0��p�����Q?h�2I�^dPȂ&Z8j���d�O6���O��'�'�?7�����8�	�n�Ƀ� G�?	2�i�РP��'���vӒ��aQ��Sva�#���F,�.e4T͓oț��W؊7��Ch�7-*?�V,�!f&��
�E��!�V��O)�(��A��K�H�N>�/O����O����O����O�M�2�Ҫ90Dpiáh��f	�<��i��`V�`�II��,"G�n�JT���ԕ�܍xS"O����Z��]bشn���O��T���R�05��A��^� ��J�g(�C�W����,%RM�	ly�" �k���Y��X� 	�\
V.a8��'��'��O���M37İ�?y�#�>z�T̉�̑&U�Ȱ22i�+�?���i��O���'�7�@�9�ٴL���1JBF	���"6�rg$��M��O�����%�:F�9�	��� �=�4/؅	I<Y牬"�i�4:O����O��D�O��d�OJ�?��gJЙ:1��2)̊n���ܟ���럘�ڴ(� ��+O*�lZZ�ɞg��I˃)Lq����!��~���t~��'%��Owd��зi����g���8 �G��(���Ĝi��ܩ���b��b��Fy�O_��'7�B��K鲝�B� ����5�&bR�'l�I �M������?Q���?Q*�x	3S�سU*��t��k�L��!��x)�O̵n�M[��/���N�"��Ǌf�(A��M�LuAT,Y@U�b�����i>�t�' �'��X��ĭE0X �������*K�����ȟ����b>I�'vJ7Y�"Ξ4J�fã"�]Ivk� %\p1�<��io�O�]�'��6��
��1�5���8�yHf��!�ةl�;�Ms����M{�O�9z1jU&�bfĤ<Iw,�M�.I�����u� \p��K�<�,O��d�O��D�OB���O�˧R�`��7(pڝ�gF�>{�Hm;��i���C�'���'���yx��nݼ3^����(J�Sbn��������oZ�M���x�O����Oh�d趱i	�ĉ"CD���j͍,b�qz3
S�a���D�I��Ѐ�5���O���?��=�A���:=���SeU&a�X���?����?,O$Inڐa���'7B��.q �K��L�}�Ҥd��$(�O8)�'�7M�٦�BK<��f�5g��Xa4D�e�\���m~�h�`Z6�d/����OE4�����"L�	�b�����,j=JsLђ0���'z��'���S��婛�*w^�F�I�:���
�$�x�ش^D�4y,O�nu�Ӽ�Q�:��o�&B܀��B�+�yb�`Ӣo����H7O�Ǧ͓�?A�ƞ�R���z➹��P�rPБ�����bY��O>�)O�i�On��O.�D�O�9��/ʐB������5���btI�<�`�i��5���'���'Q��y�H^+Wt�bS�`S�m3G�Y����r^�6|�9'�b>�6m�#c32A�T鎱!at�����y��2f�vyBo�#�!����'&�	���D֝w�d����+]ˎ	�I�������i>�'I�6��v�\�$����=N",�LSM���'F�6M)�	�����	޴]��F�j���s��paj�=_vN�e�i���Hn|骵�O���'?����h�a�o�Z8���	����Ɵ���ԟ��Iǟ@��_�'_!t�JG��5(y�x�e�Ў2�t��-O��dަu �f'��i��'W���p�ߨ#ƹ��C��1E*���O�6=�*1�F�aӸ�)S.|���$FV�� ��6T����	W���
����4�����O���tx��� ̾y����Q���p���O��i���*J��y��'��Y>� ��t��!{d�_ Y��ċ4?�X�0��ӟ�'��~�V헱_ez���,�8J>�2A � h��D�ܴ��4����'8�'[�=���@
J��q�
�!������'���'�����O��I�M+tH�U[�Z2Cҥ{���h5�^�.8�'��7�5�������O�(����r[G�ģa�B��gG�O��d�,{�6-(?�%K4���>=h��2i��@�!�5,��8�)l� �'%b�'_��'x��'o��8FЫ���BR9C��Mwݪ�"�4.g|��,O(�$=���Of�oz�=��Θd�<a�]��(�$�ȣ�M��iںO1�fP�e�|��牎P_�Xa�g�/��,��K�5CX�F��8��'��y%�(�'_�'���c�y����"[k|�P��'r�'�R�H)ܴ� �y���?��}����F��fI���T�J�2(�>	��i�7m�R�Ɋ6wȘ9�)��b�6�g�� j���oŘl�DIT�������'@�V�$��?Q�/UV��;��V�wwUu�ʕ�?���?����?э���O���!e��@x�ħ%0j�(���O^1m�6��$��͟�ݴ���y7�T�D�l����ւD��A@�(Z9�yB�f�^�nZ.�M�MH�M�Oz9Æb�4�B��L�+�摢�Ύ�tv,���&Z }X�O&˓�?����?���?�q��t@�)ߟ#���j�! )8�-O��mZ�T	����IN�s���@dȞ�>}"���JYr� ���Ц��4jC���Ox9�NM�I�T�)�/�|J��Df�Ԡ�aX�8y@�G�tW�NGs�	Uy%	aVX�dቭKbV���Ԑl��'B��'-�OH�Ƀ�Mkf�6�?9�ϔ9$T�"bI�~<6��K�<q3�i��O�P�'�z6�����ߴ8����_+A5�H���C:3�¥��a$�M#�O�4ۓ��:���
9����r�� [��>�Iw��>1u"u�36O���O���O����O��?}х�KV ��`�laS֮Oן���ɟ(p�4z���*O�n�@�ɮO"uɶI��8�{����*&���L<�i��6���89@Fl�j������+�1��y��M�?=�������� s�'�t�&��'���'���'����vaۤ8��z��)~jιa��':�[��Hݴgu�p�)Ox��|���̉|C�q1!/�7W'<�a�J~ �>�u�i�z7��O��~J�""1afm\6��D�f@rj7���gMu~�O=h���8jm�'��)YF�P=���eo�2ATX;0�'�2�'�R���O��	/�M��G�(߀���!F�4U� `K�x�r��*Ol�n�D�N���͋P�of\�j���! ���c��<�M���+̪!�4��Ċ78�9�����3� ��g�};d��rL#�jt`�;O�ʓ�?Y��?����?����IK�8E�B�.��cJ&�F�UL0nڈ�������	T�s��[���k��Ք9i�Mp��Ju:���H�6	m��ġ<�|�DK0�M[�'�ڰ6NJ?9 �u��&Q6��'椬�s��֟ő|2P����@��ȟ��L���C @YHD��Lß��Iȟ4�	xygiӊ���!�O���O.̀�!�x���H�&Ìu��	���3�����$Ʀ�ٴ2�'p�(����n�`�ʢ%�(�V���'���,���ymEo8�	�?���'h���	�`3R}�,{T�k�mI����	۟����� ��t�O��EO��6"�Ԕ84؊`V��cӞ̀% �O��$Nߦ�?ͻ6(�LX@�$BJ�I*�˚�5vu͓EE�F`iӎ�nZ0�Pm�n~2,�35l��Ӟ	�\���&0W����Wol���|RR�D�I����Iڟl�I��dJ���(��%�2��P�v��C�jy�$cӎL)���OZ�$�O���$��(�\���b�\f���f�'5�6���]JK<�|�0K	�Z�s��82}<���/_���i�� E���Ͽ5P����Q��OV�a���U��&$Y8dǜ�;T�t[��?���?��|�/O�l��9��I���ԡV�ڳn�:B��:�ɔ�Mc����>	`�it�7��¦9��S&j�8���_�����[�N}�%�i����;CA���O~q��.��0����f�H���g�P�=��D�O����O2���O��$:�5�����1ڞ���!J�~�Y�I̟<����M� ��?��$٦�%����.6�R�c];�ޭ�ݿ�䓺?���|��Eٴ�M�O�	��:(�<0t��Zհ���ah����IG^�O���|2���?i�w@�J6kS5Im0��ۃB{:�	���?�-O��lZ�p|U�I�t�Ib����7ut@�J�,S�VΉ#� ��s�O�m���M���xʟ�qQ���^��i$G>�,y��@+,6a�[�L��i>ʠ�'���&�(H���d#��*r�1�FB^ş�������b>5�'HN7mOD3��*C���$��T�̔<&��&#�<���if�O<��'�z6mڡ
b�A N�/�x*�I8�nZ��Mӱ�)�M��ObxD����H?��RJ��܊�aP�)�T�@Ug�@�'8��'r�'���'哒/D��Ñ�4☳��D9(�N ��4,�<����?A���OϮ6=�q��IZ�FJ@9�¤�;BY;2������4Q���Or����iZ�dH9K�<�0��ԩ.C�|�eMV�T��DSWkz���Z���Op��?9��?ܜ!S� L�;�RD,�z����J��?q���?�����EЦ��� �ǟD�Iן��A��k��II��PD8r BY��@��� m����JY�����.C�.����L��by�'�J5b�+�1R�Ѻ��4J�ĺW�'>�@#��@gJ}ÃV1�@1'�'=��'R�'�>����Ezr�Q�{��r+ıe�}�	��M3���W~q���+�.�Z���k	����_�`V�ڟ��ҟ4rG&������?�c�??�>�S�:�0 ��3ɒT(&�`��S�IDy�O�'C�'�fP�mJ�g�X���8NR�I��MS�ς��?����?�����V����bmK�6byk�c~�`�Z�fv�x('�b>q`2LC�g��TkG���	v�ڝ@�My
]gy�&طkm��I)t��'i剜}�d��O
�U>i��˛�~f>��	����Iҟ��i>=�'�6�+����H�b�@�mt~UIRBI#�t��BȦ��?�aR�|��4���kr�l��-�,k��;���*~x��9n��E�t6�o� �	�=O�q���OӮ%�'��d�wI��8���1E�`!Jۜ(8�%k�'_b�'���'t��'x�9еM�X��pȓH��#<PTKu��O��d�O�qo����ڟ���4��]~��gK��Z&��QF��!�����x��fӄ�oz>}�$,Q���'���զ�H�ÕM��y�|bC��S�VI��9\��'��I䟔�	ϟ`�I�iTP�^4�20jM
wE��ԟ�'�6�	��d�O���|�#L(�)�m�N��z��O_~��>y��i6�6MSJ�)���/�>XB�[i�a"b�]^z��쑖D���,O�I�0�?��n�O���1k#o[�`�rP�#��DO�m	���?��?9�S��'\�	��M�F	z��Ņ�+(x�BS+�a|�`�������I��M�I>ͧXh�	�M����+�}���N�~��aa�эj���'��Az��i��Iv�<u��O��o�("���}ʗ��M�������O~���O����O����|D)��u츓�cE�
��{�J�`ڛVA��wb�'�����'�R7=��yu	�k�rlʶ�_���8b-	ߟ�lZ���?Y�S�?��dm�����b5���gN�&{���&���Γy�<hr7��O��hJ>A/O�i�O|�H��R�I��`�E�ݨV *Hb E�Ob��O��Ħ<���iL��*�'12�'f�̡q/�e��}��)�4�=C2��c}r�'FB�|�DŴؐA�Ǎ�<�D�0
�����y�L2�f}Ӟb>ݑ�O���J�h�����ej��q��)S.����O��$�O\�$.ڧ�?����?b@<@(s��d��3�IX��?!�ih恫�O��l�៤%��*i^�	� ˏ[� q��J�D�	��I��ȓ�/I��Γ�?��%Q�.���3� �@�����fD��� '
�{��dZ�k.�d�<ͧ�?y���?���?ٔ�S�Ht�uyF��i��趃֫��ڦ�JI ��8�I�8'?1��>qx8P��78�8ER4��!N�BE˩O��$�O
�O1�TTpr�WT>z��F�-m�
M�WN�+_��7�R]yBh®rl\������Ē�<��f*��c��L:6N(ro��d�O����O��4���;ݛ&	^-7���T J
q8�ASQ*~�P��<=��Fp�0�)�O����Or�D�H���Ⴌ5�l< d��y�y0f�a�r�7$f0f��?}%?]�];oP0�)ug�!5-��J⌃`;�I؟���0������	g��Z�b7ǌ=("Ԉ��v�`�s�'#��'�6��ޯ8��	
�ML>����59{� �၀�C�*����A�}��'�F�s�l�i�2;�6�y���I�_t�UQ&�ʟH^�=��O�G�CsF˓d%��q��RyR�'v��'�k9h�T	���Q�-�R*ŮX�r�'>�ɹ�M��Z��?���?-��=0���#Q��xĈ�A�,�`Й����O�lڣ�M���x�O��$(�Մ��T��97�(�oׇX��1�a��G�jt��W�H���*S�E�M�	�>���Y�8[�^D�&��b�<�	ҟ��I���)�wy"df��B*ƕ2���jEAЖC=�LÒ�I�l�h���OHqm�_�G[���(a��Zb�l�T�C�6���a
����ɩ䞜m�Y~򇖈?�$��'��D��.����˝�o�0�#��m��D�<����?���?���?�/� �Z�+�?$M�u�  D��(�ېI
���`�������	Ɵl$?�����M�;v�jM(���1��H�ԀM�6��a���?	K>ͧ�?���l��8ٴ�y
Qn*\�Q�Ѻ}���j���y�µs����䓸�D�O���ϨM�DI��N|�D�+��c����O��d�Ol˓��eG*|vB�'H����0~�� Kwv��3#��O2��'��'�'��@t��W�⼙&b�=E�P�a�O��y1Mǡ>��7�\z�SCy��O�X����/Yj�Ӟ�V����O0�D�OT��O��}B��l�Aw�DB�,�y���7E(`H9��P��F��1:��I��M��w���#��P�<�L�ڣb��XNaa�'�7��ɦ�Pڴ貄�ܴ��D�c����'~��者� gmN$3#f��7�`Ԫ�� ��<ͧ�?����?9���?�u�3W���[E�U�^H�N���$�Ǧ���g���蟴$?��]���afL	]��`��#�����-Or�Drӄ1$�����ۀO�2^���Hw�1��Q1V�5!�(C5��,�ci*|c�k_�kyb��U����*/Y �Rh�v,B�'�2�'��O�I�Ms��H�<��E۵gqZy��%U04�@��<ag�i��O���'��'�b�2-"�c'/�2s��b�j
�0�v�@�iE���O�M1��/��s�����]T�Z�	{< �&-Ay@��`�j��������러��ݟ����d)31K�-�X"(��L�<Y��?�Ƕi�v���OFxo�|�	f).���lD�*��g(L.@,%���	�@�� T: m�<i��!̞\Zwa׻/��-K B�$����;gz�	Z�	ry�O��'��a̘v%>Ȉ�jM� �rxi��׷e%��'��	��MKq��<���?A*��I;TO��+�ظ���K֜$Q��ĉ�O����O�O�S�IT��+�# 8j��l�S @�$c�n�Xhog~�Oh�q���*��\0F"�p���A��0WϨ�J��?���?�S�'��Ă��ձ�a�'Hn�M{�IM��A;�GU7R(�h�I����4��'�
�N����Չs~�����2����V`�+<~X7�O�#�F�����'x
9�S���?���T���w`߮ZR�RF�_�"%����di���'x��'�'�b�'���V��E���"z:t�%hV�qRdߴ8
\�p���?!����<���yw�����q��wU�U�#d�9��7���U�L<�|����M۞'D��0S�5g�	wR	��=0�'t0�Z����0���|�W����۟H��c�*������s�cJ�� �Iϟ���gy"�lӪ�H���O8�d�O\�Y������e �&8�11fM%�I��������شy�'H�%���x4ؠrHJ*z*���O`8PD�1ڼT"��B1�?����O�h�p*�'aP�*�&ԆI�dɛ �O��d�O��$�O*�}���j�ԓ䯚�'����g�(#�!���j����Q"�����A�?�;K�b���n،Sv&���@�)�VU��?9���?��/���M��O(�
�
N���ḋ(g��Ű"c�.�2�ZU`�!u��'��i>��Iߟ��ҟ��ɇ�<��j�%����hR)I+H�'

6�ȿE���O��D)�9O 8h�^?��1�qEK%P�r��"@EB}��'�"�|���n�c��l馡Ө�8��˜hM6�s@�it��.s���D�O6�O�ʓJ�Z�
V'�]��T�W5Ԭ<����?Q���?I��|J/O.�nZXS�I�:��AJ�*��o[2��Qe�	�Z��,�M���)�>��?���r`A�v��,!��Q�NQ& "���%"�M��O�X%�X�(���.l�xjC�A�ݲQySbY���Oj�D�O��D�Oz��"�Ӧ��191�L�.��1��C='��e�Iӟ��	�M+�f����֦$�,���>%��yF��$qT�V�Ƴ��㛖%z���B�Qr6�<?y�k�]�? Hh(��"C����d	�,� ���ǆ�?�	(�D�<�'�?����?A㇖3r8��9p�"��v�W�?�����R��ck���I��h�Om@��ڀ��{cG�l'�U��O���'G��'zɧ���'S$`򰇇�W=D���I"
qJÃ-�
l���:�����&�Y�O�P�ޔ{PFޱi�,h�jD��I������b>!�'�7�V�/��p��� z"�2�~�"��%?��iU�O=�'c�.��5ateΩ�@)�
�#�'��gFwG�V��Hc��9�q�����T�g
*���*K�R�*Q8OL��?��?���?����i	?I����H޾C���񃓶YX�n�#?�����0��Q�s������k�BW�	�	r'i�7o�NU�Fċ�&+�6�b����<�|�L�M;�'^f�Id��zL�ӧ/ V��A:�'3>8�ǆN��db�|�V��џ��$��2�R���n��LAjH�BӟL�I矸��iy	o�ZD�%��ON�$�Oָ
�H�\�F��-���|�2 ,�I��D�Ѧ��۴*2�'�*lA%F�^-��P�Ru`���''r&eP����V���d쟚d;��v^�E8	�$U/M���QJ@5��@��'���'��'�>��I�2�|���Y (..I�I��_��	�MqǏ%��d�ئu�?ͻ�f�c��%g��+��_�Q�|h�Vۛ��lӂ�lZ9���m�T~RDE�r�����)}��,���G��������o�~�Z��|�S�����	ޟx�I�4i��1u�"@bV�U!����m	Uy"MpӲ�BU��O��$�O,���$	�M�P�
D�R��I�PkЉ:ƌ�'c�i�L�O�O�T�aQ���l�E�vL�I#Șfq�轀�[��P�o?Z��}�	~y�b2b��fݹ:9<1�6�loR�'z��'9�OJ�	�M+�J6�?�3���>��E���� kA���<���i��O4��'��7�����شٔ%B��6]�x�� ��	��AQ�oZ��M��'LR�(/��S4l��I�?��?;�
IX1G���fX�`CKN���ğ,�	������,�IK��TP�
dRw]�D��"ś���Z-O��dB٦5��d6"��i�'�&�
E��%
�5���	`���Au)2�$ۦm�۴�zq���MK�'�i�P�((K�"]�~j�-bW��^> �)d�B���|rY���	����쟈�B��	",	��Y�-DB��I��,�'�6��r�����O^�d�H�I��`hB��-<���z#�W�D�O�ɖ'i2�i=�ʧk^d�jٗgv<�ygfڮG��慔�}�� �c�s~�O�V���'f��'���1�^!rx�݃ea �QR`p@�'A��'���O �ɭ�M�v�G*a�0�Ȇ,�/Y�)��5rz�.O$xmZN�Y�	��M�DDK��� �%<"�SC��/iF���'��	���iC�	��l���O�']BU��%���,9�ƀi(m�����OX�$�O��O��ħ|�2G#F5S6�ې17�ճ�@��楓(f���l��u��y�lX�?T�a�� 'e�&���G�<x��7��ꦁ��ny���#�4w��5O���ɑ�B1�'�X�*�T�I'<O�	���3�?ao5�D�<�'�?!��q�2ap˅�,"�����X��?A��?����D���Q(��şh��۟0���ٞ5e��iSa�&?�^,5�R��0��ɖ�MK�i��ON]0�Ǖ%k�R��vNRwbV�x���R��\�}�X{�,�{�S|��,��4"$a�*^ʘ�dN[�&�HK4C����	ʟ�	�`F���'����LػQ����f#�4_j�!�'�7�%��I��Ms��w�L:өHf�8���Vo$r�'=r�'B�Ħ��期D �������5f�b�E'!�>e��j��}3*�O2��|���?����?���: i#Ȓ��l8�*�fh+O�nZ�Z���؟���K�s�dKD�R1Pب��b��4���R֣�<��D�O���7����}��L�%�4X�0�cs�Z��fNd�v�@ �Cī��T$�8�'⅑p�ˑU�@�HO)k���g�'2�'�b����P���4m����F�P	N�K�lE8a��3�ZA̓4���dd}r�'���'����f�:��Z�h¤9zT�BAݠp��=O��dn�Kx|��y�O�7�,l&0�	�+�� ����/��yr�'�B�'��'w��I�h��ꂣM�6��l�/ ]p���O6��[¦qp��Ny�#qӲ�Ol� ��8xhL5��MxɴĈЃFp≖�M��ig��)ZʛF7O��D�0E�zPp�˟ �)�흮v���(ą�?)��8�d�<!��?��?���B�u��
_2���{�'
��?9���Y̦��U���\��Ο�O4\P v�֒x���	!8%�x��OH�'EB�'�ɧ��ޠMp؅�smH�y���a�fF�qG���G�f�\6�Ay�O*p$����<"~����&�dA�<o �5����?y���?��S�'��Dۦ�I��.|r�@��()�	�S���*i�	˟Zٴ��'�X꓃?�5����Y�B��txdxPRoT0�?9��'��8ܴ��Ā%"o����O�In�$�֊��E�ē�F²Z��Ky�'���'n��'��^>e"�A��H�fY�5'�xb��1��6�M�7̝��?���?�L~�m0��w���H��J�m���0��j�����'K��|���n�P��&=O� ��ŬS�+CC�4q�r�[V=OR�z3e��~�|W����۟`�F�N5��Y��Y�|;�E�5"�ȟ ��֟���Zy�Dz�ֵ�Ƭ�O����O�@㵍̷���iU���#�b��a,��&��������۴�'kȹ�W���
y�Ԍ
}��K�O��)N�pN�����?IF�Oְ��!��O�\|Y�I�5�ݱF�O ���O��$�O��}j���"�8RcX�J�4|�J��m4�5i�� {��%�o��ɂ�M+��w������ʬfr0��ʙ��d$��'��6M�Ʀ�z޴-�:�ߴ���3#���'9���+vL�D���p�%J�r�;!+�$�<�'�?Q���?���?�kB�c��P���/:�Պ�<����c�� ?q���Og�`2Ё�6Q�Z�{�[O���S�$�>I��?IM>�|b�,��\	���VL}��k�-O�X���4���Z��~yR�'��'�削������G�Kp4B��W�-�r�����h��䟈�i>�'��6MMw8^�^/ �$CB�&0}�L*PJզn)��d��9�?��X�������� �^��+[�:�T�d�M�;��sRZ���'T�|9b��w
M~�;)���哅@��N�d�̓�?	���?���?�����O!B���� 2j00j��|Pf̐C�'�b�'�7H1s���O�l�x�ɵj������I�O��z�tU'���ϟ��spm�I~b�Z�2����4�l@����e-���2Il?aN>�,O�t��D�Ob�$Vͦ<8En���Q��K�uQ\�d�O\�@`��!M?fv�	��O���厈H�D�"�3%��=z�ODD�'�R�'Rɧ�	�=\`M����1���3c\##F"���E��b�07�fy�O�6��������4%һ���A�`�Ö�?���?���?ͧ*��@����D���=�&�K?���ŏ��4�3�n�.������ �ٴ���|"�S���ڴ3za �iR3�h�P���#[Ფ�iKr�;��f��8�T��s����~�ǦY�0ZƁ{a�U�]�fvCn���D�Ob�D�O��$�O>�D�|�+�&`[�xoُB/��#J2Q�o�/b2�'t�^>��	���2���ǡCD�x�b�D�T���`Q� ��f}�@��<�|�2L���Mc�'�V��&�@�R���@
��q*6��'�
�!��QܟL��'��zy�O�¦���a�)�0v����m�-2R�D�OH��^$B� ��ei�(������5S�LqW�\$c*P�����k��x$���	���d����:޴�?�*O��kёF����n˶P64A@��(��ݭ߬�j�3�S%����؟p�4�Đ �J��%Z��R�g^�������IȟpG���'!@����;@��ek]�.Hh�'��7O<A�h˓��6�4�V�Y�A�gځK��9@8鱇8O�AmZ��MS�ta�Q��4���9K	|��'Y����G"Y<Zcҵ3�*��]�6�z�;��<�'�?���?��?�Wک��Hۆ��#�;U� ��$�ɦ]���|������L'?�I+q�;�h�3fr����ř��*�O����OؒO1���QL9��+b�('��e�V�ܑ,446�&?�WaF��IB��qy�Ҡb�ܘ�d) �Q�(�Q �N?
?��'���'�O��	3�M;q�ܱ�ɚGE$�R���R���^����ɫ�M��RH�>g�i�T6-M�I�����,�=�b("P��1�"�X�n�X~���+����Se��O��.�cn��� j�L4�֏�6�y��'�2�'���'~r���$4٘�%J�'��2�l\�T�
�$�O������q���ay��s� �O�qQPDS�:T��,2)ØE1�MXW�I2�Mc3���4Ś+"֛f���b��<6źy[��ݶ�>X��Nغ��k��'��i'�����D�'���'���bf��.%*(ȋ�NāmM��G�'DQ�<��4_�53��?	���i +8Nzicg�
+&2���I�������pݴ\ۉ��i�ny\Xb���b��eq�Ǵ8�N��'�?y� �����S3�R�t�ɀ}�����`�S���R	vd�����	�\�)�Sfy�v��yj�5T?<a3R�I5�F�JUC�#h�|���O�HoZi� ���ܟ�k�	�8XC �*�Id*���	��HlO~2$Ζ������Xp��p'h�_eX�+����(?��<i��?����?��?!*����1-^=sǦ�\v���S��ݦ#�fٟ�	�x'?��8�M�;Q4���&.F�@��b�IR�����?1I>�|�g���MS�'ǲ0xS�$ad\
�۸-�X]��'T�@&a�d?�L>�(O6�d�OʽQ�e J���'c\�_��5���O����O~��<��ip����'���'����!
QpDD:"��(�$�<�	���D�O��$��ߣD��s��ݝs4jsA"�:uX�ɻ;�h�#oM�ţM~JǾ���Iy�<�C��44z���;:�j��I��D�Iğ��	R��y��B*���i��ŉ.�:�JW�g�r�`�=�����ش���y���fZ�31O�)�fq�Sg���yb�'3��'�i����Y��Xфן|�(��,X�`8��@eY(��2�'�D�<�'�?!��?���?��e�-}��@�B ܋.\���c! ��D�Ҧ��a�e�P����@%?牓=��	�� 
�X(xZ��F+7ܐ�O����OL�O1�*��� �xs�N/�rQ�R@x'L����|���D,��%��'b.WhG�i_B�AV-�;��@�4�'���'�����T\�X;ڴy�`Γ���u�w����@LE�6bX�͓@����d�m}��'�b�'W�9�F�T;�ar�kT7-�D �_�Xכ����{ry�Q>U�]:.]E�5���V�<�B(�� ��	ğ$��՟��I���u�'�Hg�/ BH��D`i���?��K���K�����'uN6�3��ҙE�2��V"͌|. ����<!�.�O���O��FT�7�0?�tf�W�N�E 0�6�k�M��µh���$��'(��'��'9Zx��l��|���-�8mN����'�"R�0`ܴtA���?����i�.K�,�@eӬ:�jdr�m���I,����Op7MB�|�B�B(rT��/G*AV9˅a+TP�`3��#K�Z���G�ϟ� U�|���<\lHAMďr\^��U	��y��'�B�'����T����4Rb �� �&-�%;�gS�aKh��Wب��$�ߦ�?Y�W�p!�4DhL����8{����BL˂MD��B��i>�7-.��7M4?��l�8t����)�MN'Y,�#���SQ"���o�;�y�R�@�������Ο��Iџ@�O����̐@]n�Pt�P�#�ە�p� � ��O$���O����DFզ��<���{�),.�R�Ǒ�#�V�����MC��|J~چ`F��M�'� |b�4	$t��O��:A���'N`��`aB�����|Q�������W�\ό��b�n�4Zǆ�럤�����Idy��~���b5O ���O0<�B�)O�����B�4M:!E"�ɭ���O���#���s���Q�~$���' �}��	�8�HĐ�	I�9�|�0볟��ɏ �*٨F,�0�r�>C$�p��۟L����l��Y�O>�)�9*QrD�##�>z��
Bg��b�nӔ�QUo�<!�i�O�.N#Z�J8Q��
�)�F̰@�L!���O��$�OJe�q�"�3������?��R��\�lx`i�\h(P6	�\�	Vy2�' ��'|��'W�5��f�19]�x�$��F�Ɉ�M��ၨ�?���?)��d��1rAK��W�6\�!nY>I���"\�<�	՟@&�b>��A��c��<Cd�W5�]��E��� o�����J���\h�'��'N�`J��sg"Χ��)�j�F�������ßH�i>��'M�7�@��$����G�F\��r1*��V�,%�ls���D]}��'m��'"d�fh��5�����}�2p	$��:g����ʠ#P�Q>U�]�`�4d9�!�f
<��+����	֟x��ПL������IT��;�M�e�ԃ M�D�%J�.R�����?i���D�3w���M�O>�SN��d~̩� ��4�j"(P�>�'��7����XAnpnZf~ҧ�{��<R�.��1���A&h�T�,�ái��H3�|�Y���0���p�� 葯�zF=Rk����JyҌaӦ�8f��O^��O�']�݃�d��B4�����P(a�e�'�f�1��k��<%��6�Jui�I��6��XR" !D�\Hc/CE�$� w��O~�O��i�ɚ��'���p�*O	qh����2�`��W�'���'5b���Ow�I��M�F�����'��=_��yIt�ϳ!���(O0nb�Y��ɀ�M�`�Ɣ&��t�SKT:P�TYǘ�-t��D{ӐT3�w���&ڊusCK����O���)'��L�����Є$<lp�'�	Пx�	�l����h�	S��%�a
�ƃm1T��f�Na� 6�_9d���d�O��3�9O��mz���ER�ur&N%p�8���M�c�i��O1�*��q��	&"��1W��Ք���h֍6��s�H�y��'�f�$�����4�'^�葔i.'�XT�U�"L�.m��'�2�'�X� �޴
��b��?������S8I��xz��K�_�T�ۈR��>�1�i2�7m�W��*���b횇FzmZ#۵H������e��#���|:u��O�s��1-�����uv�mh ���*�!����?���?9��h����T�����3���dV$2��$U�!��A՟����M[��wL��b���Rin�YD�@6䀐�'�7-I�Y�ݴnc�H��4��DZ, �P�I�'~U.�*��۠
����a�Kj{�Y��+�d�<����?���?i��?!%`��FO��cԋ��/�ݱ�1�������ώ䟠�	��&?����C�<%G��R�8��P�ٛ|�60�O��n)�Mk��x���oRs�<�4������^)X�SC*����	k�z�x�'Ov�'�ܔ'��T(���7I�,܉s�ʄZ��]�A�'���'�B����^���(pvT�IqPD2Di��Ȳ��
=r�ɭ�M���ɰ>)��i��6�����dD�*�A{����|���	G�gT��lZK~�� s"�/B��Oh7O�-c\�pk�H� �F�PŭB �y��'�r�'��'���A�jT�óM�I�VD#&����?Q�i�X��ȟ�=oZZ��?A�ͣ��Jk�9B��� '��L<q��iP 6=���P1&sӤ�}�$���ŗIg0��←�W�|����P���/������O��$�O��d<[� =9�f#}�l�zu�ۤA�����O�ʓN�$R��?Q��?�.�L��
�)�6}��m.I��:�����(O~�D}ӤQ%��g�? � 3�H\>;󞈱cT ���B'2� �"H��9����|� ��O�|M>�w̏�,~҅��㕶r�����t<���i!�0Z���,�L�fD(��xy�*��I�M��rf�>���i㒹a��٫���`Eb2Tpq06y�~0oZ��p�nZs~��Y�����S2�I5,g�}�䢁 b5$)��%��D�8��vy��'�\��t�ЏcW��(#�P�\o���Al�.�y`l�O��D�O��?Y����ŢOè��5�
:l�0JP��.��!x�v�%�b>�獑禝�,��X@�2an�aK6]�m�5�6!�(��f�O�őL>�.O&˓nh��6#O$a�Qc�6\ą��I��M�T5��$�O�A�Qf�j>b ̘79j-B;�I+��dEݦE"�4b܉'@�8y�!]�#��q�@��|����OZ�3Pa�;� �A!�)��?�!�O�;r'��YY0f\Y�)��@�!��8�4��rFl	� hbfƄ/E����ߦ���ܟ���;�MÊ�wkļD�qV��B�Ɯp�d��<���i�6���S�������'���:o��?����@�z���+�|��Ē�c�'��X�'?�D$���Fi⇭�&��lI�O��o�~���'H�i=w�����/��1��:��,�'�6��7�OG�)��\%6�:�
_�n�����-D���:�Ϛ����'�MP�� �����|�[���SNC�`0��`��jj��tK���T�Iʟp�I۟��ay�oӺ�94��O�� �ĩ|��8����νR��Ol�n�a�����8�O(ml��M�W�i�\�F- 1HR(�aj��Aj�pbBߘdO������C�ɠ���F��ߍ��46��J�y�g/|�H������I���I�L��' �,~�����G+�.�	D&H��?����?�i��!�O�"Fo�(�OL��� »BH䰑�C��n�E3Ն�X≊�M�����G��F��� ���H�E��p�b!���3H�I���E�Jyb�'$"�'2�� ��}I�.&<~PA1���#(B�'��I�M��T
�?���?�+���
�b���hJ\.��Ib9O6��ZH}�loӰoZ&��S�4�R�CI���HĊB̢����CHG.9�j,D�`aX��S-l���Es�I#*(�1�ǃz�.�ȆA�d�BT��ܟ��˟��)�Oy�Lc��rE�%6�~Ҷ�\�l�$AA�!�V~��O��n�e��Ο�+�O���­ :���P�L�7�Iʔ�ޒ8����O��˅GnӠ�&��ԓC$�?��'��)��n1gl2�Rq��$`���'����`�	���	ޟ���F���-����@�"���K�%oM�7�/G����Ol�� ���OB�lz�)�DFA�	�xLi���8Vhx0e��?�ش(�ɧ�b�",	ܴ�y�81wuдOݏh��r����y2��!M�����-F�'���џ���2���k dׇkW��D�I{W�|�	��,�	�D�'��6m�!�*���O���N� ��0dBCF`�q�s���Ov���N}�'���|�i�-���D���ژ����?	4���"/j��]'?eѥ�O<�d�$��Y2��&9"\)	Z�^]���?A��?a���h��.׃:�j�J"���D(a�WȜ �j�d�������C�<��(�M�O>!�Ӽ���L������V�p�_�<����?I���ڴ���5+���O\v|���0F�&a3H�$|}:T�|2R�P�Iџ���Ο��Iß��f� 8�n�B"�*M�pa�q~yr�a����K�O����O����D]����	gO�!ݼ����@�y�'zd6̓ͦ��I<�|2�
�7ఱ���4��.=�P$h�YQ~�iZ�]f@��	�"��'d��;�<X�5�	Q
*���	O���Đ֦�s��Ɵ��(&�Y9j�940)�b�ΟZڴ��'����?Q��?᧥#�zz��
>��P�ҥ�#Ml�(�4���K�&��m	�O��O�g�֦0wt�z֙C�-Qu 
��yb�'/R�[�6��yZ�ϛ���ҥ�'�b�'� 7�L�h��,�M�M>q�Dl���x�� 4'�h�ğ.���?i��|"u�R��MK�O9�򣚈B<ܑ�d��S�O<���'y�'��	^��E��I�3b����#g�!4H�Fx��`�vŘ6	�O���O�ʧ���ZS.ױHk����]��'���m�ve�Ґ'��u��Ӎ�%;�nHA�ڥ8���kP'	k��u�IƮ��4�������@�O�w◆9.��M;?h�����O<��O���O1�Jʓ%���]9rDB��`gV<}��,�u�
^�t�*�'rb�m��⟰J�O��Dܗ'xZ���4{���{���*A����O�ܙ�k��v��aM�?��'�^��U�Ѱj� �b�
G1�9�'���\�	��@����0��E���*���Z�� �E�N��"#��¶6�K�p
����O|�1�9O0Xmz޹�Ӊ�*i�bl2KC�{�� �$J���MS3�i��O1��I	��l���2`[�T�F� 6�X��@�s��I_��xhS�'�'�t�����'�|X@�h�n5�pIшDfniXG�'q2�'��T��Hܴu��P����?A�5H�5�"���U���^v����b,�<���M㗐x
� �H���,�D�B�ۈc�Y
�����E�C/b!(��T�(�S�b)�����Mn\V͛#B@� E���֎*D�8Y��N�t�����ƃ�8�x��d�П`8�4�t|����?!òi�O��/��	�c
+hTД��'E2�D�Op�d�O�Ł�'k����%��ɱ?�xV��XX����
_ �t!S0�PY�IayB��0|�@�pc��9X z���TAj��R��F�6Sm�' "�i��E��!��^�r'Pi��	�;�5�'��7ͅզ5)L<�|�qMR�R�j��C^fu��A
S�Huz �����MTx�j��d,�Op�yO>\A����쭲� �n�����?!���?���|R,O"mڈz�\����6��<*�nݮY<��� ��z,: �	*�M�"��>I��i��7Mۦ�*�.1�Z)�#ɕ�2�m�v�U���mA~��W�L����V��O��K��"�*���-O�.�bE��y�'���'R�'�B��ܛ&X��W�#c������]'��d�O��¦���d>!�I��McN>Iইom�`�DO	(�6,�SIֈo�'�r���4��1���4pSO΅G����ٓk�ތ�@d�Y�h%�wmF0El�	�j�75�����s�Nt�@�Z����Nt��y��o�|�X�J%*GZ0�X_�"D�6H�]@�u*Q��<d�|ӤO_��zE�X�������,&a�$Q�M�Ih\x���
�J	��b��j���'��i�.��p蔰O+2(�F�ӭp�Ph16i��fY[t���y�V����}����E�^�;dD9eB�&8���"�b� ` o��I�������X}8u��@��d~tC���8^�~V
� �#D��>lvPpA�K�y�H���K٠zְ=j��	�+H$s�l2�����O���d���� �r�J$#C�o����/LC�i&�t�	��+����/v�c�������*�T�d����*ߠ<n�� �I!Y U�	��8���<�����i��b���oit�	��a-Rm�)o���O�X��J�r�1O���}3���8yz� /ŝq����F�iqg�'Ab�'���O��x��76*`���YF6�=��b:/�&6-M !Y�6���<�PE�jr�a6�F�n&j!����M����?q�'�4�,O��'�?1�'gpY�$�CVU�E�	&�:!��(�ɤEPz��O|*��?���k�I�RP�B+@(�G�>�*����iZ���e������O��Ok삝9�ܥCg��7|���
QiF�a@��*U
���Ihy2�'�B�'���>Q�j=!�	�wm��D!��)�)�֡��$�<Y����?Q��ty�<����0�T��ӡ��l���srH7���?���?+O��j���|�.�i[V-j䀒 ;�$�� F�є'|��'���;4��Ֆ6l��#��v�@�"�I���ҟ<�	ڟH�'�I�P �~��6�-c����t�Xk�l����YG�i���|��'�2��)d*qO @�h��w�� ɢNXe�IW�ip��'X�&������$�O��IO�vN�z f��q�0�C�E�Y"�$�d���x�� �I�����\�H��"p��F*�6ɘ�Mc+OԽsAI��m�	ڟ����?�ۮOklvvlV�z}�,��Le���ش�?����8���i��S8����PF�A�ƊC2Y��a����7M�O��d�O.���~}�]�X�a��1cw6���z80)�)�MK�GY��?�I>).�����3V�KnH&����҈�������M���?�\�0\X4]�Ȕ'9��Op!�!MI'a���u�܆3�I�0���!Z_(�O"�d�O^���42\�GK��^�k�(��v�:�n�˟H1���9���<�������Ěs��x�UA�I;xA�#�}��	�'R�'�[��B���Q�"Pyq�^�T�����I���O�˓�?yL>Q��?q���'qޙ�,�~��	!�Пe�0�H>����?�����$U<Q~F�ϧD8̙�e� 9d����H!=0|o�xy��'��'��'�����O����$��Et1�`JJZ��S�Z�(��џ4��ry2���F���9�VFD4 �>>֠�����IH�qy�O���~� EO8|�~�Bf�\��@�u�����ɟ��'l��"I<���OH���Dh@Ԡ> �"l�0�Ţ{k��j@�x�Q�8�	韬$?�i�-�Bͺh���`Ėh+P���B�f�D��i��맀?!�'��I�����Ѐ��f��ʘ%G"6͵<9���?Q��t���4a<| `U%H'mH���rA�!��4l--����ܴ�?���?��'������8I%D�W��Y&>h��N
��7��O��D�OޓO��<���;�\�Iժo���Z=��C�ia��'�b-T^��O���O4��,pl �F�NyhR�AQ���7-�OڒO^���y��'5��'-p; g 
D!��;���3\�4`���$�"Xf��&��S�'���%=_D8�D,U/r�+�-��L�,O��d�<����?������o�4��3�O�u�"m�A�,��XK^J�	�8�I|�IlyZw� ����u�t����9��T��4�?)*O��$�O����<qfߞ~�	X� ,`X��)wo
h����ȟ���l��Hy�O���b���Ι8���PG� \]���?)���?�*O�p�5CK�+b�J�{:pĊu�A"تz�08�ܴ�?YO>y.O�i�O�O(虚�.��p�\�r�ڀl�zH�ܴ�?�����0>���%>�	�?�8� ^��ƃ�Ha�C�"ҸXd�xRW� �	���&?�i�1��
��8�=!1������i�>���a=��H���?�-O&�	�<��Fh5��aV����/LaZ-l�ȟP���<R�r�3�)�ӷ��)���#I�Q�X��6M�7f2l���O����O���<�O��i�%ڤ$�,R&eZ�&�T!�e�j�đ�S�� :51O?���e�7h@(�!��	byv#����Ms���B$/��S��>�Ԯ@O�"��r��"gBDeЀ�$71ONLc@`[짌?��'��`��P�*Âa����f��5��4�?������
U��d�u�\i{��8�ٰ�g�,,����'����A"Y�Ø'��Q�����w�~p�e��x�ܠR�J
�|���Ggy��'/����O���W� td��N�4yĮ߹>�������p�����@���ܕ'uj� ��>��m8���0�y��s��>����?AL>�/O�yC ��O�m2��Y3�J3e��,Yn\`W��A}r�'}"�'�r=�,�I|���&{z��@V`�+RO��I4!�%4�f�'��'i�
f��!��h�	�6Ti���ԠVJ�:���E�+����'�RY�t��d��'�?������X�&rB�bF�»y��#LC}�'剷W�r��	C�X���"C�BcF�jp��ŠR@}��'�hL���'���'�Ol�iݡiu�A6.f���L�2�&����,���Ot�����Io1O���`y���r�8�J��R�s�)8`�i�>���Ev�H���O���f�&��s����n������S34º�Z�Ao�V�RQ��O��d�O2������g~�k�(o�H�:A�;,�c�C� ��6��O �$�O�<�DOX�i>y�I^?��o�)��=�ni������	Pye�+�`��<���?	��LX���� �<R�T@���T-�|s"�i�B��
P�ꓢ��O���?�1R`�IP�P��L=Kq����y�'B^|��'���'��'�"]�|��F�iW���@CV85���
�kU"�n���O���?�+O����O��dO.m����6C�.ܐ�v/��,F>O4�$�O��D�O��d�<	�O"vH�@9]x�ѡWɖ'*�0�"��:қ&[����Sy2�'�B�'�1{��5Ƈ�X��@�O>_P� �M��M���?����?*O��'Bo����5V�	TА#sb�U:���N��M3����$�Or���O`4��3ON�d����O�(	^
X��O���)�Ct�l���O�ʓ��\��Z?%�inZ�?�S�ò#QB� !lW�,X��v�	5����Op�$�O�t"'4Onʓ�?��OGȸ�sNG�.r���c�*[�*]�ܴ��D�9��n�埜�	՟��=����}�u�I�<Ud�/T����v�i���'�R-��'��'�q����r�:G��U�C�@y^��6�iR4�{ �h���$�O��D��T�'��ɘU&q���ҟ1��9�l�(8��hJ�4���ϓ�?	-O��?��I}�\ �'�2Z:�h�kզz?fLJݴ�?	��?YAO��5���ry��'x�D�8�5��)��Q�	�0�ȼm�ğ��	�� x��p��'�?����?ٰ�3\�Fȳ��@�O�i�Fj�fc���'F�-ap��>!.ON���<)����i|	���<pr��zF��n}�%���y��'oR�'2�'��	�%-����B�m6����&����BP�0�
�'v����X�'wb�'�r�Tb'.  ^�H��MS X�ı�	R�<�(O���O"�� �r����|���4�H�,�U"Ĺ�dP��'"P��I�d�I�7���0r��dM��$����<-O���On�$�O����<�1mЄ7��Sӟ�䮖�*F�@����;'�@2���M�����$�O��D�O6T{16O&�'��l��AH��I��,9~>�r�4�?y����$ָFYf��OR�'���L�2K�Ԁ�)@�/?@l�	F$^����?���?����<�,��d�?`D��*�( �u!��z����`ӊ�$HH�i��'���O�z�Ӻ�`�ـNk�L;�㏀K�����E�=��П��m~�����/�Ӻx��!Q�����`ԡH��6�]o��)nZ�����|�������<�A�׾��͋�d[�}C��zu��s��F�͵�y��'��	C�'�?1a� �$�6I��o�>Bx-ڑH�(F���'���'�藪�>�-O��D������=I��D�9"B1�f����<!4���<�OB�'���e�$(��h]!7��G��5n�R6��O�K�f}r_���	zyb��5f���f5����u4A!�Aú�M3�c�~}Γ��d�O����O��y��[t⎕b� ,`�O�#Ft�D�ձ9$�	yyb�'`�I�������9�&D)��X�%	M��:��$- �d�8�	şl��柨���T�'�hy By>��&薨
����oðrpl �v���?+O�d�O:���� �ѭ2�����Y�A����E�WI�ƕn������՟��xy�9G�r��?�1_v��soH�,�"������p�n��@�'���'���(�y"�'��ąG�~5CWF7)NH*bT�˛��'�2U�P0'悙��i�O����<!2��J�~b������X�P�Br}��'_r�'�@��'M�U�����6�զ��"�&�csL��9. 4m�Fy��cI�7�O$���O��)�u}Zwx�!�`F�-R<蓧��9���B�4�?��^�������O.`Ȋp���Rsp	S׀�'.j�yٴ]<��"b�i�r�'��O�J���DQD�? r��g� D�f��a�	�B�(�iwX%؛'<"P����hby`���; F�IѮR�=L`0��iP�'-� H��0OP�D�O^�	*s*�AЎ�2^� �CuNf6m%��ݏ+Þ�$>��I��,��6 |�x��޶)T���!K2�j�l��<3��
��ē�?q�����Cc�7Oښhg�#�ŀaA}R��y�\�T��ן��Iry�L��;�<pTB�7D>��7A���S1�,���O��D:���O��d
�;����N�!V�I��!��.������O���?����?�.O�}��j�|�D#N� �ذ"E�hR���� _}R�'HҞ|B�'I"������T ��ST�3� %�ŉ�#i���ݟ����L����٣��'Tle���S!J�h� H٧\�ܭ0�iRX�����@���}m<��o��� r|�RU�� l�@����H����'�T�0��@���'�?��'(r����m�?��D
E�*L�������?���1r�iϓ�䓽�$	�*�b�9Pŕl������8�M�/Ov�"V���}Ӭ���d��je�'���cתl�l8IE$]�D�HHܴ�?Q��,y"���䓧�i���Y��PfΑb�I%*PJ��n�j�������	ɟ �I�?9O<i�v��`S�·CU�@Ia�F\��a��i�
�;�'-�'m���N5 ���EK�2���Ʀ��ʥm�ҟl��ޟӐP���?!��~
(qXHp
�J:	�����' ӈyb�'V��'�0(Aum�9��P�F��iq"�'�Ӧ�d��^�0%$�X����$&���1Ndy�`dǆ"�*q�� �;���JS�N>A��?1������=jyv�#�ɂF�ҡ�6����2��a��ON�D:�d�OL��Bl�P�W� �԰;�
M�[�r���c�Op��?A���?�-O���.�|
����N0G��4o�1;�H~}"�'g��|2�'f�CX�Xh2��f1z<چ�ڴR҅Q\�[E��>���?Q�����Gt�'>���	�
u�pA���6L| ��ӊ�MS�����?Y�ĸ͓��ɍB�:�"��;@��ZP-քm�6��O����<��h!$��O���O�:���������F���a0��#F%��O"�d�]�`�D1�d�?��u��!C��dA�Za�dJSo`���=-��Rƶi�꧉?��'o��9)��!떬1a0E�b_<�>����O2��^��6+տoT �JgB�"oڥh7�i�*���jӄ���O����"Q%��S�Yb�7a�.����}�,�ѨOz��9�)�џ@��#C7%y��0�
<V��e��R��Ms��?���LD�f�x�O���&4�䦘>K��;ţ����LoH��ӉO�b�'"��)(�#W�J'ø�^�FȰ6M�O
���d�w�i>Gy£܋�ⱙ@�Ȅm�04�WM ���?�+O2�d�O��.Z0���T|*�(Q���_�X��� 3���QM<���hO�I�>�}�gF�'/ARC �[,=�6�O\ʓ�?Q�����O���7�?!��b�F�p�HSv��PEm�L���O��$ ���O��U�����[�V�I��@�Y,����&���O��D�O4�v*��Ē�T��9
��!��o�`�ȁӓ�6��OޓO8��:�C���G�g��a��:-ptm�џ��yҧ\�W������쟂Q�a!h�P��w[5SBًp$�^�I�����R��"<Q�Os.���]]����й$���:�4��DH6p�0(m����)�O��	\R~,U=LG~4��
+;D���f[��M���?���_i�'3q����V>@�R��'#���%�i7���Jc�*���Ob��쟲d�'N剁}Nr}8 �S�=W�
"���=��4q�~]��?�/O8�?��	�yv0�6�]t�	��)�`
�qڴ�?I���?!���FM�IHyR�'���Ý)H YJ�B ���2������'k"�'�������O����O� �&Eģ(]�5p҅0+�<t�fF榍��.�0�Odʓ�?�,Of���,�h�
A'Ɛ৥�;c�F��BZ��U�l��I՟��I՟p�	py��ïu8@�b�o�â4�d!�1�iSl�>9.O��d�<1���?��]�؊T*ŪC���*EC��v�@�<y,OT�d�Ob�ı<�țe}�I�#�:�k�f�n&t��NOb��T���	iy��'���'�Z�O� ��!�"JT'ͣD �a�i ��'���'��ɜ]�����n���*�X�/@r����0g	�[夤c�i*r_����؟����\�Im�ܴk���
J�: �5��H5KP�lZƟ��Iy"������'�?	���23�[�jS�\~Yb�fȿ:%��ҟ��I���j��d�����]�@&��G�,��$�t�Q����A�'�j�Z��j����O.����Qէu�t#H=�h6	�b`��̮�M���?Q1j_�<�M>َ���X~��1	f���z@Ƽa�F��M��{6�'d��'�� �>y+O����Շq"���GĆ�w�t�C��T����soa���	ny����O}p)$�T�4=6 9�dݦ��@y2n|-���i�O�ӥ_��(��?K��y��K'.	@��yr�[!������O���S�v��qz!�R,�v�0R��:n$F�mZ� ѣ�0���<)���$�Ok� &T������];R�ʒNގA�@T�؃z�d�'�"�'l�Y��q�٥d$L�A�]6x^�ـ�̊�+���Q�O�˓�?�+O����O|�d�<gO���ga�i�]c�A��q\IQT0OT���O��O��d�<	��U#Q�ɓ1=�i�3�ع\'
�[F�!N�&W�`�	Ny2�'}��'cl�p�'v��٢Α!Q|D��c�!���铯g�����O����O��&���qGQ?��I:Gn�QuH�/	��@P
�7�8�ٴ�?a-O����O���J<�O`���|��-�7��"��)�iPR�'��	�~|�k����$�Ox���3ú,ـi]�:�*u���J����'�B�'W�����y�^>�Ic��iݤ��Y�ǍO�)���Q��ަ��'u8}�o�p�D�O����P�էu'F�z���rK�IU�e �/��MK��?��k�<����?a���O�^(`�D��`xµh����q��ŋ۴A�I#�i "�'�2�O�����D�&uؙ�ڤ":��	$��\P�8��8;O��Oʓ��Ov��6u͜�\85*aB�u(�q�b |���d�ON��:H\���'��IƟ���&2��Ӷ%���8Tl�>:4LoƟt�'�M˘��)�Oh���?9B��&��qP���0Ӗ�C5Cwӈ�Iu��ʓ��S��(%� ���'���ۤ�Q:p2�9C�� ���U�'�2�'U�T���0G>Ԕ����'W����7'ƄZ*� �O<1���?�����'R��R�KҚ��К���S���Z�%���'���'���'+��O�%_�KR�g�Ҥ�e������ ��6��O����O"�O���<�O̦�锉E��8�^2N+����f�>y��?y������>��'>ib�d�T�r���{�F�I1���M3�����?9��~+΅�>qA ���`4M5&۴�L��a�IƟ��'\z�) �!�)�O��	��i��ha��2zX��jZ/TFʡ'�������c��6�����L�{�qk�+�]>j��eF��Mc.O�Ck�]�������6��'��)��Fٻ^��\PbJQ3ޙ@ܴ�?q�z#��ExB�)���I��h]�T34�IѪ�v���	�7��O���O>�I�b�Ο��k�>-���B�Y&�q���MSV��G��������s8N-���*�q0�nV-GP�l�������<A����M�$�'��d)R�ƅip���t	��M/>�lEx�,8���O���OJ���ǜ%1���	6��?�B�Sȑ����I�����O<ͧ�?1���In~��P�74�x��`-~�VqjQ�<���?���?a�j 2�Ƀ�@)�y�e�<xճ�l �?���?����?!K>���~r-L�z7�5�5��;�:��V(׀�M� �F~��'[��'��Ʌ2�p���O.���R��V(CCK������O��d�O��O��D�O�̃�Y�|C� �E�^��&�J�G&��B�>��?����ץ5��T%>5HTm�7������("�� p5C4�M�����?���|�$�>�3蕉V�*9��c�
DA�ٚ%NU٦��	����	��,�hP�P��ߟ���?�2�$�!6����ca/d��ًBH�6�ē�?�/O�L�S�i���抜� ^��*��.{�pa�bg�^�G��۱�iav�'�?��a8�I	*38�)
�V (���D�J�O��j�c3���?O��B��?Q-�B/ �$�}ɶ�ic�A�g�'	b�'���O��@�$�N�,K䀀���=� ��G(�m�>�{Fx����'_`��%�*%������5Oc��P�e�$�$�O��d��Z�$�8��Ɵ���:�����(/TD	R`IE�{K���>a�N�]��?���?V�@�
q��Y8�`�z�n��&9�6�'J�'N2�$�OV�D>��ư�a�BG�[�̥j�NӔD�RP�R\�PEg1�	��I�� �'�,!J��פ}{���'�-c�!zU��0t�zc��	|�؟��\� ��冘aCR�#�d�F�u�&��ԟ��	џ��'k,Yu(t>�c��W���uK&�Eo�*$YƋ3�d�OȓO��D�O�]��X����'
s����e�e�T��a�>���?������Ѷ�`A$>鉢	�)���3�IH�	)� ��M������?���� �>�����g��ˀ�T<>�w�_��a��Ƛ�'Ɗ�J`&+���O��ɓ�*r<HD��{�hH2P�
)G�>&���	՟�@��,����e� W\����Tt��t�w	���M,O�@Q��L��Qy��b�$�>��'�6a#�
%(��wEHP<�cڴ�?����4�Ex����=Q�t� �ڹC�L����>�M�1LC�6���'���' �T	#�I�=� J�L�)�����BC>�M��ɜh�'����$[c�}�DM�^5l4J�FK�=8�m�|�I�<A��fy�]>���b?a�B�K�BU���ٛ �>;v, �I����J|���?y��EK�(�7��	@j���c��J��]Z�i��b W]t�Q����	e�[5L��y���81����%/E�'}�'���',�'_���.��5��@�e��G��DIbp�'�r�'��'��'��O��XN��$���+�:��P"�i4>��N��5%�X���
�Z�@cb��4� �gm*����@#ˮ�b�L�y
� �-ᤤ[p�be��Ót&��1��M:�z�(�lH% ֊���+Y���-T�<Ү�CԀ ��q�R�#���AK/*l](A��kep��(� �Fٚ,HT����]�7[Hi+�L5u��i����zɐT��<f }yB�1$��p)�G)r�`#ʚ�+�l��q��<��]�7��	��Q��B�e�d)��ԍk^ <�����B�'��au�O�MA�|XS+�e��d�sYVr)�����CE����]	>QPkő>9ӈ�!%��(�(A�zq��T9,�p%*��~������T�W�:�J���B�D��XR��'��>}���	?�|��\4% �K�E�3��C�	�5�.�h�NT9SА�%h�����d�'�$���W�j�)�D.XiK�>!���?Y�QA�����?I���?ͻ �����G
$���b�B����{cH"��SxJ �'	@�g��)"���է�$�hl���m��!�# �!h�ɀ��4��|�-�B?��	#h����V�Ґ��S1�O�)'�@w*b�N�K�=�b��=9�U�ȓx�#g$�4PGnU(�0��'�"=�OI割dp�:��N�)�Т��k1�@)�%�>�4�����	П:]wr�'P󩎍F� ��/� /Eh̀T$,"������ ���� �ʗ|+|���E1M���,B�I�+ք6T�@�Q9�Mb��oެ��d�9�Z��~��ȹ@��A� q��'h��Ic�Lܸ��.,Th1�m�- ��ȓ��	1��߇ #N(��!S�?]PT�<yA^���'�xа�l�����O�1dƏ_;�c��[1Nq@���OF��/����O,�hW��$7��Tosd����	�yΒm����	�x�
��,���*��}��)��ց+�2e��$YuT���+��=k����	^;uOz�Ey�$�?)L>��b�-h�6�YEA�!qq��AD)�Z�<%_�����G�]�7�Z��I�z<��i�� ��I�-'�T�"�=hM�Qىy�+�6FI�6-�O��d�|j�d��?&.R3K0�ԃ���m��Ȕ"�?1��Iz�����蘧򙟜�f��MLPT��-�6���u�0}B�V1�O��(
U���<���C��&ԥBV�>Iqc�����<�@h�:]���C�ςq�(<��h�i�<���c��:���/?�=�P�Ld����$
�t�ɢ�K3@H$!�����)瘟nZ̟ ���<i�	S<T����I՟���ן��!����ف{N|lcd�@ =Ҹ�<Y�'MHx���Ы�/p�����g�9�n�B/�I�p[J��$^���S*S�8vz-ʴ�Kw�c�0괅�Oq��'���toʉ%�n$ ŝ/_�q�	�'�4	�Q啃.jU��m)	>�y�O*�Ez��)&#�*`/�tm�"�H%U}`�aU-y�P���Op��Oլ��?����T�Bش=p�BPv� ��7/�dl��	�M_�pZ�}�R0P����O
d�e���\��!`��
I�}��	{�Ļ�	��!+��d(�.u�����?�!��e�r}�O݄�f�R��CF�<�󅋭7�����F,d�t²��C̓S��O��b�ƦM��ٟ8��ɐ\�\�2��]0tNhЪ�E�̟X�	%,�)���Lͧ�����r�ɬ��Y�7wלu[�i��R����;v0�Oba�u�^�)�����É[8$٪A�'�2�����r�&����	0��D��'�1_��ȓ?<�� ��#Y����u��,E�P��@Û�h�}�tQ���P�,��po԰Ԙ'r�UO�>����)��0�ğu�l�F�*f�*TOZ)i�����O��E˳u�x������T>M�O%^-�6\��j3��<l�
J�� �A˂N�ڑ9ŀH0����p ����m���ؔƋ����6�>��)Mޟ��	R�O|ҧ	/c��}��O��H���'D�@B�ɹ݈��⮋�@3VL[R�"����[i�'�B���A=b��)��C �Yd�����OB�Žk�(� �E�O[nן��i�E�T��ND�jR����2�c��d�&����ɼN�R1�G�9$`$@y �F�qz� 锥?<OD��s$	@�Jh�մOE`��)5�	�ME���|R&�2Hs��ڑj�
3�1i�&��yR"�=0�F)�N�`�B숥Eט���CC���ر���@�R�,,"���?���p�&2vSD����OF��O�D ������?�O��86��yt�ӤO�6@B���xBg��ڼ��E�D�R͋�G��q
�'�Ҽ����ش���CZ,�ȡdGD�?i	�S�? Z�0�A��@ѴT1t�wl
��f"O,��s�K?�,�VBݻ]zJ�)q�D�f�A��i��'"t�&/�r4�(�PꝒKN�Y��'��
�2�'?�I\�H �q���3�dɇv?���s�[�nڀPɂSt�x2X�^�` �x��V�b�H�I�MŹ(4����+���p<�&�៴�	iy�� -J*1!��o�ZY��I��y��'���ᓿ[����P�/�>�0������C�I �M#p�π+��Er�*�_T�9R�S�<1+O"��d�=��ӟH�Og*�i��'��چf�*08qx�N_f�h ��'bۜ�r�T>�vg�S�W6�p�2
*��9�O^��Q�)�J'�1��)�Rgx�u���N�'���0��˘��O�^�I�j��-[.�S��G1�8j�'..u��c� u�AJ1H�)#Ó[�ĳ@�J��Rýe�l�˖N5D��iqLM�N1�Y��vf���(D�!5<)VP8p%A�iUyZň%D�����o&�q���C�5]R|��'D��J��_+^����ÿ7s6ȸBB%D��	#HĦ}F���wA������ D��6��f�\!ЃN��8
8-1�=D�ī�=�@8�.F�F>��7D���C/%�rd8$'�-H�i��0D���զƤ�fM��j�!{bD����"D�pYH<����ơ(�"�;�D5D�А3k�z����,H0[��	`�=D��� �Z�!�rUy��K�![����-D����k�!0�й�򋋘�� �-D�
3�XnbiN*(||�f8D�J�)�ZGbtK3b�<`�X����7D�,J�m��'�p���5| :ѩ6D��FiQ�	N�Z7Ȇ�����2D�p��.�UZM9c�y4��+q�1D�� �#�袱��ݾo�5��n1D��JG��+;��9[����B�OlF�B�*���k��4X��S#M�B�I'u�̓S�
�f�&iK�>L C�	�h��];�ɃQߎe�Zp�p�&-D�<��fJ/j9\8dX�#� �$,D�l��3����E[�W%�<yW�7D�T��
	�=�q���C|���5D���VKM�#@@���2#h@�5D�!7�{o��H�Dҽ
���@s`-D�,�u��q���ӇI�.\�z�3 �,D�<;C��0TQ��	Ho���ܳ7�� P���Ot�V	װ<B��B��$u`<�A"O\HHd�R%��%YE(^���O:� �.�(�0>	�iǌ]�e���741 ��}8������W��d��hD��p����׀д<�!�䍄}� <��M��/�ɉd�ǘQ���`ጆ����=�eGś.?����U�}U�$a�"Opa!��.XTS��R
����V&蜭��y����c�X�@E�7c�r��
�4D��8W�Z�i� ��P	�|	;���O��ن�f�|Ҁ����E*���F��p�t ����=)�O���"ƜeJ�"\�C�T*�U�!��p�ȓ<���{��Q�A�0X��bߦ
z��?�4@@�Pq�qG���y��ɹ7�K�l��QK�.��y��\�����W:��q�cCX7P �U��{��h���X�A�H�h�Ǎ�<?ڈxp��!��q���%F��"��p.юR�	\jh��:��hт�z9���M��(㤑��51޲���'����d�		1�ׂhF�!#�' H�Qǅ�,r�"��uE�J6<1Fy��!w(X�~�cmS&7$����1�X�$�c�<� j��کd�p8��5~͈b��<(��
�}���'�&��g��I����(g�@	�'mXyp�-H=�[r�I*3�����'I:ȡ�g<�Ov��b�l�.���DZ���T#��'���Ɔx�020��0fcd���(�Qg�"<O��#��h�NA�$���F�NRܹ��<�>B䉞4�}i���$\b)PTO�0(�x�Or	�O�2����O*�-ɱi=V��do�9��0)
�'8�m[��R�.���H���2�b��<R����Ol���ʄTTZ�	P
�	H�M��OJ�9 �� �RP)��4T��1C/]�G	"XJ��+��
�A,mz4J�E&�옇�	�25
�N<IqaG%E�<"� Z�
��EQ���y�<yg�_*=� ���*E�E���@#d�m�<ɦjBBh��@2ዽQ������A~�<�u'ݞR�X�Q`�Z�֎4�um�p�<��E�s&Q��A@4x�'E�<iV�L I�,�!`,<Dxd��eGD�<�B�$?;�q �&��q����`�3CP��>�萛w��y����L9�5��e	{����cZ��$,���z��R	I��I��D�=�!�6`�A5*<b�L�K���=��O`�g�I�O�D�;EZo�4���C4Ee�|�
�'�J�p'��PՠU;!�\,>d%�ѯ�
#y�Oz�}�JHI9�O�X<�hX Mۢ�^	��_�������'Y�(3ng
m�f��0�O���h�m�S�i��(��E�X"W��8�
�r�!���| q���ܛ.��xADB�6ܞ1*@1�	u��~Ba��.��͂��&��9Ra�=�y���ǒ�rdI�@H闂�?��,.C��}��P�R,��kq�ʖD�JX�B���=	T��7% �	�u����uJ6E��x��
����B�I�b?���
=?!�[T�]�h"<I O>�2kF#��0� ��G
j<(c�#D�D@�bJ�qۈՠ��ާ8G��b!D��s��.4i���X �sEn2D��Q��Y����`�+K�X:m�g%<D� ���zV~�!"��"q�� >D�ܩ���Z�uRҎ0%�Z�g)D�D�#��"�X�Ǻ8�+� )D�(�Pe�D�xkbeK���щDC%D���d&َ8�VQC��G(hޖ� AC$D�  '5���ae��T`��5D�`�w�_ u*RKC7a>��	 D�h� :T@�h�#`|
l��H1D�����09R� �p�P5��u2�-3D�L��S�h�洺�,���A ��,D�<��*�8��\���ݒg�BaDA*D�Ac�D�N�����⚾Q�$���F)D��b���aТ��UA�,5�성�(=D��
���2y>�D���	�&���`��9D���t�&l��Łc挵C�,L�'�9D��7�O�Qi>\�h ��,B$B6D�� �Η��|8GeÎ��( !D�,��/\�6�6���M� ��I�=4��3V�?{��e���JU[�Ə1gmч���]�ć&q������-+�����$u���<�g�����:��H;6����B$Po�<�f�!",����5tBx0��m�7pJh�?�}z��DZP�Ö.T�r���#�@f�<9�%K�t���ڇ!O���e�th�J��h�	Ó5N�Q�o^�puzL	`�S�4�Ɠ=���)�D�bHxbd�31ߪ�q�:�xb	D�?9r���JI*,���y
� 2�a![�as�Ż�g��Ӥ"Ot��A!�@h��)T��e�i�e"O�qj��4�i�0!<v��A�����L��	2���a�B�2H�Ѓb��$�"���2#D�>���hV��'���5I��ژ(�wn�55;H��ϓ҈��n�7���/>i��c��G\�8�O�D�1O\�:�G�����O^���	�?Qj�i�㟪`6 M2K>)A㞨d>mrçizP3U��:`�R��s��צٙ�7�ɣ+S�#|�'zp�E�Q��T*�!�bfX d����fvx`��ܴ]�8��!F�Q��ڕ�L�;�ܩ0VK��$T��O�I�5��8/�9k�H
# z��x#H�e�te�t���B�yrʋ�B�@�ϙ�w$�rFFtb��R=R^P�h#C� ���ax�p�6h!G� �'.��H1J50�"T��ae�@Л'#�AS�_U	R�$y���
��iہ,�r$�䎐1�!sQ�+m�=�2+�<�D�*��E�T6O���C6 *�Hf�^�{Yʵ� 9,EA&�Q�$��D�/��K�3�ŀ�y��m�DP��oݹU�
����c��ِϓ
��T��9����U<������	�l �7 �0>�^t�g!�s�'�������|�I2�l�K��3`�|]�4��-4�#>�EΈ�3I�bD��k�����|�T�/H���i��f��4�Lwܓo��,Z��ڦ~�h#~
���#"V&Z��҈���"A��?!fm�,,�
�H��5I��a̧D#�;T���a��] '��,ȳaq]�-%�N"�%�O����
[?�C�ùc�$m:W��;�Ձ�o�x�*�:rAä3�\�WJ=X~6��ãҋ�Fx��[-}����!̊�>t	�ϓ<ެ��W�ѽҌ��O�X�!�ƃ;�8�[�CΧn��x��?O�qZ+��*L���ҩ�q1��0�FL��k�Q���Ǝӫ�Qq@6O��?+Z�#�Ą�?��̘U���<���b�L鸕@׾=��\c�ɿ �v����m>�0��#o hxRD�.D�Щ�,�	 z��C�F݂=�?E��?��r�  �H�vhP��\�A_�A�&��yrn�Q�LeYvɥ~B[�3���0�2�0�p��,;�b��W6u�@tB# ���x��?ҧ��s��Ђn|5��$��/®��ť2L����N�o��]�$�*�M���e��it1�Ӫ[�P	D��%��G)��1���8F�!�� ��I�p�ѐ}� -��TY�U���?h��22��b
%[�/(X��D.2���P	[��������I��I�*���aܗe�IY��%m�u��B+je[qi 22ȝ�Y�f�0T��1����Q��Z�<1v��	(��9	�) �h�tЖ�������F��P� 9�P5	���&>o�F�4�*�:OM8U��6b��m�p,�9��)`Q�'�
-�v��h�P�*B�߁/Ff�:�ԝVì}��B4|�flV�S����% �">����X�,C��*H���:�l�u�'��x[� �Kj��)��ؓ-V"-;E �Z_�+�	�(/����/��!�$�m+��+�K
 �b���f��I�T���CS�C3X����e�2EQ>yX�_�6�V�9Ш�Q@���4D����.U�c����R��0�^��g� ,KlR�:Ҁ��?	��E����>�O�*�&��CA�'	��
�,��!��,ke�����@	o���7+��!�d�%��ȓ�
�l�*Qc��-�!�ĉ�MW�QYD�D)n�y��bՆ*�!�$GH�6|iP�ë�(����J-g!�ˍԌ}S��)o�d��뇡Va!��@f6в0'ڱf�J�7+$D!�D^!�ܐ�B�138U3SjR@!�ȧ)V�L��Z����r�У%S!���9�	��:hrz�h�옃e�!�W��3��הS( J�iۈj�!�C�_�<��TaH@�Ԫ�;'�!�
y�!;u��f02E�@N$y�!�d3p
s�9&PB�ڤm�!��L�pG��q�ņ���9�ʖ�!��ӕd�0�XAG�B�)�԰;�!��
i�	�%��U�6c	e!�Ą<�m��C�/$�@y��g/!�(��c�.9�=F�	gy!�$ҏI>K6iA3��ck�Ar!��N ;��xgn�;|�В�J\?@T!�$Ǔ�ZDc����<�&�!*�D�!�؝ �����J�E�}s�&z�!�� 6�J��C2~�&�j"F0B�D#�"O����D�\�vA�#e�(O�f@��"O���Ѯ�'*%���D
��f}ɗ"O��c�#�:m�t��$�9�(�"O|Q:@�D� _��jUcI�n���+�"O����È�.Y�J@S�9*�:W"O����	�<����e	�bҔ�r "O���&Q�HW0�3&�J4V�����"O:��˒k��m����p��8"O�L����-���a���,9"O�t�\�g�he(�������"OF�8�f_�~����0�ĕ��"O �y�N%v��3�,S@�HL�0"OhڇC,��$Kǈi3���E"O�iq�H]���J���	o$lB"O�x���]!�<�sW��CB(�F"Oj4�G��9F8�A+Öv;r�("O�A1'��~o0;��3%�ū""Oq ��l�q"C��(�"O�ИLD�]����q�Gp���x�"O�fLK��8�6��F��8�G"OHqbt��>rqL�RF�?*f��I�"Of��`O,A�U�Vbԥ$n�x�"O6����ܒ`�R]�^�%I�"OȬ����/g�=1�FQ��0"O��wS)^崤�f�%��q�f"Ol)���F��䫃�}�N�Q�"OD��hC�
�ڤb4�Hlj\{"O\\�GOؠ-5>Q�B4e.M��"O��s̐,Gt����R5-��V"Oz� U�D(v��mX#�_�1r�"O�MH托Z����̡O��$"O�E�A��wv�i�E�A�M�µ�D"O�}�'�iRNp�SH?H����"O�����;D��Ԁ�I�z�T���"OZ�J�E�w���HM2M�x���"O�|b��i<��i�<�3f"O|٨�/dS��d�4\�Ih�"O�Ah��z�ڑ1��>jhv]�D"Ot�Q+�,��4s��W�
�
&"Of 0���<��,[�%	<)�����'À��4'�S��jbJ��X�P�	�'n����/�(v�0|I"e�,O�RR�'����piD!9�0qrT��{����'*���4�V	1߾�:�H�@��'�8�'��jF�T�@��N�4B�'1꽁�J�*�(�#��A�ii�'s���bI�u�ѪWBW5�fQ��'�H�Btj��h �9�!�&4	+
�'ڞD�M%k�F���R�;8�!�'CV5��V$��a
�@>r��i�'�.�xь�7X��|!kJ�s�F!��'�܀R.�K|�A�Ō���H}��'���Ej="�* 5��
����'��X��=4�q�R9-)@��	�'�MYTf�.*�tI���=<�6�#�'̠����L�[6BI�Ul��J���8�'7�I�ć�$&�� թC�BI�'�<( �_�lBL�g ��9r��s�'�4�Q��#|�mkw�4�b��'OTLA`)�q`x���!B$-��)��'Q����Nݡ0\��ID�0�@Ѳ�'z�ғꊩ=�`0�yby�	�'Q���#�ԙl��J g��oǬ$s	��� �,[�"�*pQ�-Q�!m����'�'����'�D9	�D �t�$����7i/2�(�'&�=h��*��a
��֚0�T5��[<&(#za`Ф��,X��V�Q�(�7'J~�<)�\l|�'�ò6`j�h��"�b�ȋ���O@��� ٩`�H��@+=0���"O�T# .ڣG�����J�& F"O�m��Q�<`��
�@�?v��Yf"O�I G��:@ʄ���Q���S"O�M���G��� ���I#o�|��"O��c#��&
���ऀ1?T09��"O���2"B�P{a![�g�0���"O�|���.�
X�e�-��J3"O|`�bNިJ�m��-ۈ[�؅!���6�S��OE���R=�i��+Qk�!�$.6��$��*�bU��R�A��!�J�2e���݄DO2		w
Q�b�!��A�FɚM�$)(G<�R�� !�䘿.����H�H.T�� ��v_!��"9M&-Qör$�\@/"!�ȹeը�Б��7*
 ��$&�/5�!��čoL�[���$3���G�!���1E�J�I�鄱V�rQ˔ �!��e���+`m�RP��膊�)T!�d��YA풍+7����D�UQ!�$�=;.fy!�eM9q(*F�dH!�d�1~�T)2oE��j��P�@�!�$�$��"AY]��13w`D>�!�$	�F�b�A�VoYҝ+!�"V�!�$�'u�(��3	@*�=3��/�!��I���i�	�&&v��w ��6!�D/��8��C\�C�U�樌#=!򤇬S�"H�"@�&\t��?�!�G�{#@��@I�=B<A���5u!�D^!~s q
��΀qk���Ɲ�g!�P�l"�Yf&��A.\C�%��n�!��fyر�FKV�4(W��b�!�D��;]�� d���s��$�rcQ�!���c��jǊ�:+���D�E�b}!��!6%���w-�+n��t	�LQd!��ۓp��Z���a�v���(R�!��6r��������	ǘ=�!��\JX�t��8��=&8!�5�Z9��� L�P�M !򤙁_�i�.O�X���:$�ޭ0G!��O���зcʦy#��ˆ&�-I*!���o�N�d�Y�%7`}s�	�g�!�$G>��@�s�[�o����C���!�dA�mo���FX�z��z'B[� r!�#9$<�����+g��y�@ ��!�D�=|��E1W�SA��3�!�x�+$,J<ar��PX��	]�O�8�1�� -1��W�.�j�':���	�5*Բ7k�B���i�' �Ԩ���.-RV���)͒
J���'9b�� G�6;��SB�.� \a�'�Z�+�H�L\�m
�ϟ�"��D�
�'w�e����f�v5K�fH�e6����'C�,c�+bc`�W%_aq��I�'�r��d�E�}�1���҅Y��+�'ib�Q4#����kߒdMظ�
�'�jT��B�:_3��i�e�5c��D[
�'g��b/϶MH����䛃[<���'� q�!iD*H��B�c�N����� ��j��ڮ�0�Kv@�*�(��"O.�P,��%�S�NW�\�eYb"O���E[i�@��QM�<��"O���%CaR �+VSv���"Od�hd�X!���b� Ui� �r"O�<�E��=2����j�TL��%"O��`N�t2-(��ئ'�Ô"Ox�#��әA�(���;V��x��"O��d'K2������p�&q�"OA�SF�>3�D���N���h�*g"O�!i�C){ǈ���Vl���A"O��*�F�P#��.��8F*:�!򤎏*�T%�u�Տ�B��Ei�E�!�d b¸��3��"M���fF!�B
I��yQS�Y$0�0h��NȻG9!��>��� �藱h�<�I�-��D!��ŏ.Em��M�"��,I@g_,!�ĕ(�N=��ԾTè4��e\�!��:���D�7��bd�!W!�d�K���rf�r�6���LW�K!�dR�A�4�ط��j��hе�g=!�$Y�H |�,H K���*��#(!�;m96U�V��#Cr%�R־e�!�E�t�t��6�˹J�2�q���!���M� ��bw��
��!�dB1zpP���)
q�T &�-�!�d���Z�f�R4�`�[�?���ȓ0P&Rס�<�<�[tkĘSZH��W\"Th���-LX����"��'���PZ�!x��U�A�U=,c������q�wDƍW��ېߺS��C�r�^�Z��7��Ja&�!R:D���N%a�.U���kH�%��N9��L���11J-U.~1��K��Ry�Ms&a1D����o��!�x��o�Q��J1D���Td *3챐���,���f(=D��2�?1T�}�� *vِr:D�� u�Lp��Ӥ"�
�dI�K8D�� �@_'TT���^������2D�����Y�hѐ�![ ��m��J2D��`K4�|��s��/v2����.D���'�[d��m����� >����� D��3ܷ"��`"eG�v5�u">D�x{�-�Һ��U�.Q`^��>D�����%�D@C�	$p�<�	QJ6D�����ͬ�����N�4�0��1D�4;�
�{d(�h���"����j.D��)0�;&�0�y��:Z��VE:D���梜�)T�P�Q�V�"��rK6D���!��Nh0s*ă �
Fm9D�|�0�ـ)��)) 0�]��!;D��J`H�9�L�z�ݭY���VO7D�Drvf����(6����2�� �4D���tn�U��84��"(�5H.D�����:O��(�Mϱ,�:u�V@+D�X�&ʀ�V��Q fJ�x�H�g�,D��0���B?��B��A�H��!i6D�(rgk+8a�3,΃T�� 0�i/D�<�'��NY��� )�`�g�'D��aJ<y իf�J({��y�#D�lӒ��	�p�;�j�� Ġ-�d?D��
щ�,�dL��瓣�:�	��1D�<�"+)K�0+Ta:$�(m�b	:D�L�CFf]PѮa����#c6D�� ���B��6���3E^%9��df"O.�ʃ��`{� `
�$�""Obd�p� i*�jFB� �60h5"O(�AA�Q�7��X��A�;��|�"O��(W�@,�B ��$`#�%=�Py���E*�8�FΊIւ��F��\�<�fK�&&���M�;����p.�t�<�Rl��n�\�� �Y�9�OOK�<�#ĩ�Ԙ�h/�
yՍ�D�<���
6:�܃�حT���ơG�<���]�u��lhw��)������B�<��;̤l��*�I�a�[G�<i��>>%���U�ڈcP1%l�C�<dƍt�n��w�T!�ҭ#Nf�<�d�B$+��E�"W�$
�<�+�[�<�%�@��)��j�Z��ƉY�<��T	�yZ��΄^�`�0�	K�<q��)q�B2bF�l������J�<����%i���k�Ȕ4ٚ����C�<�@ͤ@}Z|�ï�'�jU�Q��G�<I�͝5�:T0����(�i��GL�<�FеJ_�hC���vW2�Bo�N�<a���FF�a���H1o(:�i�K�<�f�Db�����Z�!_�\��iB�<it醧N*\��eZ#�>��FPv�<�Cg~����Y�:�,�!�p�<�AI	�
��ĩ�9���`A�o�<�7�čh98p!� @�~�B��C�<cF��喙*#��w��=��o�@�<9%`@�|�"`�V��:@t��NJ�<Q��QR�Ţg.��O`��PuMQz�<9��ʎ��	R	ւn,Nu�z�<.�0g��Ɔ6vh��K��^�<ytϟBƂ!� 0ZEpţ�O�<��cW�M��h#�2%�ʈ�1�M�<��Y�?��j�W�+.�{R.b�<�bkԀ��,xW��	�N=A�_�<A .�U�nhz�ސ.4��b`h[�<�a������kQ2��I��U�<�(����Y	��Y-I�z�1���M�<�f�\��$�ņ.E��J�@�<i/ʍd�L1I�h�-T
Q@'ÈR�<Ѣ�����kH)�}@���K�<Q�B�	7�Y�'�"<K�ab�n�<1���$�6����LE��]��lk�<!1eM#<�V���D@+g�Q� l�<1jC�-��� ���H�&��R̈~�<�q� �X0L�Ign������@���<I��Q�5�X,�r���E�XAa��{�<�.u��̨���:Y�`�֍�w�<)�-[� ,�u�E�š	�U3«k�<ybǔ���Dj� �2j'�s���h�<Y�(�"��XH,�%���ら[�<YVM��l�4T+�@�;s��`x�X�<�歜�x'����iB7�N��#MWk�<q�,:u���ۑCǅ.Ў}CV��j�<qA	Ps�:���?(���E��~�<9�N�**���Є;~��,)!a�P�<��A��^kb��&U�&�$�&��A�<	բN
X�)�OV2=e��x�l�B�<��l����LQ�"�Z=pu+��_@�<��M*!>�j1˚�Lm��3�&�{�<`�:7�pwAT @ 	�_�<�gm��A�1�0k��v��d;g�^�<� �T�jR'�ֈ:�kO�\��� "O0�ن�B*,2�tcԋ
>� XY'"O�9�vd�gk`|;�dMZ�P�!�"OFt*�e[�L���F��p ޑ�"O)*�_�~���'&5n�S�"Oj�{A�*|��sG�hk��3"O�]#3ᙉCFȉ�)�>|>�E��"O�h���!>�jQi�hɀI�D��G"O���%�E�4
��1�Z�G��Y�"O�pH�ɚ#|W�٪�̟��(� "OV%bìŜD��zc���u��	"�"O@�RQ�A�w>�J�I��9��"O���@�oW���ݶ^��|K2"Oh%��=-���GN��}K&��b"O��{���8%)�c��E�g;4��"Od�b�Qy(X���` 0dQg"O�E���Z( Zp��s-QtLq"O� �oZ+
վ8
��S�q{����"O���#	�K�]�r!�gB\�"O��s�M� �(9���G#�ѣ�"OB�`���*0�\QrE��ui��C�"O($�ѫ��]���,߄Wr�R"O���!`ُ�b� �O�lh("O �	�d�2ː�h��t,H�<-L����o۬� at(�I�x���F����8��X���ny�ȓ?,�:����o�Z���L��L�N���5F�0 5*]P���{Z�y�I�ȓq(��0��A�*���I���(E�t���r�RqQ".S&{I�A@��~�0�ȓRVu�q͇)J��3U��?R֐�ȓY���	�2/l�+a��_ސ�ȓF�ؘ{�GE"{������7c�x��O�5�5b��r���c�䑺dUh�ȓG) ,���4EZB�K㢓�;� ܆�s���穋$����hT&2܆�n6���F\�D�qdP3L ��J� � ����Gf���2J�6��}���AԁL�^Ej��DF
�1�ȓI���� J�p���K���fxb<�ȓ!
@u�.��P�u�'��>�RI�ȓ��'�W�XDY��F�,� �ȓgI�$�b!�\�Z�0f+�&k����ȓc�����	�=���S�B��ȓTŘ���F�/m̽c�K>Fΰل�!����ծXF���`�S
U�u��z�����*�%;�y���ȓʀSaD։�P(�d���BD��LS�Ъ��U�F=Li���[3Z:p��x"� ��Cw܌1P�'Kj��ȓ�^,��@�7a(�]��$�u�ȓH�H��c闚m;��f��3��H��0dr�#C���X#Q#�?LdI�ȓU��aB�D�!D�i3�
$it��i�h�Ԏ� |���cb�q ��',\�[1fƢeM��;��TM�.܆�s����焩��-�sBL�U�ȓ:��	���-.�� �@�uEb�ȓtO4@��d��W�����H��
܆�Zʑj���`̒����@�Z��ȓK��x���P���n��R�\���N1{5����LY���8���ȓs�.yk@�3)�i��)�[�
t�ȓm��RFc��,�a!�m3M @݆�S�? ��U�طI���ě��.�[G"O~��T�� )��BC߁Ē���"O��KgF�݂9Ģ��O��x�"O0����Sbˀ��a�6���F"O 8��Û7z���)e�I ���I�"O��	�� >�}�mT�(��R"O.d��bV�w��@��+=J �"O��j�eI�0$.�V��_
f�C`"O 8�!Bh�.�` J��K��K�"O0�yaH�l�P�( @���R"O^Y{��Fb��u��M�9ڍBe"Or\��ő�+���
�'X�AߦHS"O,��Sw�^��$e�;p�n]h�"OQ��<+|����?J����w"O�2�� F�b��I6Pp|Z�"ON�аCK�GY�\3���g�9��"O�j��ʰQ&���#%�2&W
x�"O�p���M�����%\�*��W"O�m����nL��z��Srz�
"O�!�%�1
�@�2�̌S�	:�"Ot|����G,��%鄝,xb�z��	ҟ���F�'aŀ��܀Lb2��A�~fJ��ȓJ0���˸�Z�A%�;����_6ؤ9���#�	"eD޲\K­�ȓi����@�h���Y3��.*�6�F{��'!��Hn��Lb�B�m�$Tn��	�'6r"GM���1�`�>nH�	�'~L�SEe)8$e�D&��9�\,�ߓ��'��}Y�:K��IST�ǉ?����'s��ّ.�X�4�QGj�b���'F�}끧�sH�a����YkJ�"�'��ty��u�� !��� F�x8�'�\���W��ء�HQ� �4H�'�\U���u��}�A	�B�>qb�')b�AIAo0��`َ3�� S��D�O��$.��]�R�� M�&oa
4�F�X�WS<B�	�S�X�x�%W����n���C�I�Do��ڦ�B�d�,�PE���C�	�OَL��4{�U1���qp2C�ɹj� Ī���N�Qj�o^,L��C�	4Jx���hN$wڄ��b��C�I�3$tP��bt����0/��B�	>`���L�}�MC��	j��B�I23(�ɚc�W��M�Ҭ��#���=�
ç:0RůRu?�F�+ 숼�ȓlJ�����,}�\0��M�=��d$�`��I�(��]�+ܔ�iGu!B�I(��Usuk�b��9��|�PB��lr��Q2�ٻɎ\H4����C��B�@�[D?pX��.^.�B�	9K/H�0%�ކdl��M��|��B�	�M��l�V�S#=��p*��MEnB䉭Ui�P�w�ЛzJ,���-y�0��?�\��M�@�U�A8ȸ���q����ȓ��)�,c�dtҕ(�M��ȓQ���A���qTq ��D�"]��V�^m�AG�8>*����OR��H�ȓgTy���� h0<��F�nD�ȓ(���"@�	'�Xa�����h,L����<I���� N�$H���a�d�Q�'�T�<��R�a�2�!Ҫ� r���oZO�<��E�3���!J8���H �f�<"��~���D<JX(�@���b�<�D�)S��!�`�8j�$�� '�\�<� ~�0槃�q�xq�&H3%Aۡ"O��bgε&�D��w��?
<X�O�()�"��v�h�#��0CYB�#�(D��8U���n¨� Ԡ �l���u�'D��*4#Ӊ[�(ѫBʵ���B`$D�pА �]����1J�#Q?��+G�!D�<�`K4f��KE9sC2���;D��	w��C����O��L���:ړ�0|"e��;+�vX�Mɖ*l�qiV}�<I.A�T��x�KS7>{��ㆧQv�<�bn�����E���;w�\pQ+�J�<	�'�)\�a90�Q�\�6=(� H�<���!R�����I4'+p�&�C�<y�$��N��EX��T�6�����I?D�`���ܒ]����I�7x��݁AN;D�`����"C&jeQ�Ӱ,�}�a�<����(�����N�	J��˵=H�EZT"O�Q#!�ʨz�8�E�h9���"O���1e��%��9� ��j0bp�f"O���i�i��O1Y'N�cG"OF�p���=�蕛CF�`�hk�"O|1[Ĭ��e�Z���e�0��AbO��E	[U���ǬϜl��  �K'�&�S�'c��Y�'C��6K0�i1N�sH<�ȓY�&��u��u(��6�H<q���ȓo��Zf� R�8�d̆�g�F�ȓ��]q�jвn��,�vH�7HZ���
i�oU=EFq�7E�Q�ȓ�vx�c*�v��e�9L���ȓQ�>���,��@A���<5N��ȓ-�n��R@�&OS(RSeS�9<|��0�͉����dņ�!2
�$$�Z8��m�<�ز,+B������!E�� �ȓ~0D�P�)R{>ܰvGR<#2-��	a~�D�lN6�6��Fxn ���ς��'�ў�M�LqC��K%ĜQ���1t�`�;�'������Ǿ�@�r[�~HK`l�Rh<!�C��z�t�r�`_�ddѐ�����yBB[�v���S\\;�F��y��78�B!��k��D"����� �y�d��.Ar��F+�:�а*���yb��1[#��a�O)�q�0�!�y��R[��- �� �Z K�0�y"��&5�8�Bo��;����V��y��G:�Y�� �!4�P\"��yҍE�1�JɒĒ�6 �]J�>�yn�3��ە쓾��]Y%�F5�y�ڍ_<@�p$x x���i̩�y��K]xi)���dg�hqP�5�hO���� <����
H���
�`�)r!�@ A���D����!�µBf!�O�c�zI�a��iP�xL�@H!�d܏=�>uاe��(ՋѢN�B/!�D�,R���NS*\b@ G����!�䌌]��Hh�bS
;֐�3�|!�d0mde�U�ˑJ�`��f]�Jw!�G�-���a0O�!+޲�R$ƗDs!������Į�i5�`;r@�J��yb�ɥm�rѢ��ӑ 8H�#���9M#$B䉥-w�H1�H>��\Z�cB�I���řG�S��x����.P�C�I $&��R	_�T����y�C䉱(�|�b$�2%F��6�,�C�Iq��<� i��ݲ���?F}�C�)� 1
c$F(w�H�bMU*{Teaq�'*ў"~2�Ŕ0-q����-e�-�6����'OazI���8d�@*(�8�S&ҳ�y�&G�>A���-	��q!�J��yR*�6���Z�M�1�����E��y"�C�BC�%3���y�D�{�� �yb�I�O�����j��U� f�?q����'��=��J��vv���3׃YZ��G{��I�<qt�P�8���k� �O���kf��Z�<��!��I�e���
1�L�"��HS!�
�W4�����K!���.�=D!�D�R4���V��#h� �F/�!��L]����n�D-
�,Φ]�!�M�1A�%�=J�����B,+���)�'F�
�k�%R:G2�t0�A�.Y�*����hO?��F��.JP�Y#��
-#���G��e�<�'�� w���5�v�~u��_�<1Vg=��9-@�H� ��B�`�<��ɵ�(h���>$�ʄ����^�<9��\.���k���6"̀�[� �Zx� Gx��~R(��2��|��������y�O@�K�� :�N)u� I�j!J>����)&
����0���UKO�9�!�$�7G�b`H�Q�hP)Jտn!���*�N����9F@���(�@b!�,G�5��1V���gĻ-V!����9ۢ��� ���!�LFFџ0F���I�`�f`c5�ԇ-��������y"�$A�%	��P8+��� ���?�S�O���6�R�p���-�]�
�J�'2�5r�f�
Ci�<BR��W����'D+$�Z�Veb���њK�����'���@ש|��9�mL�Q���B�'l$��O��5��u�;YdH��'��Ӈ�Y5su��ҕᅩe����'���jH�@5AĂM�Z�DI����hO��̓x��� �T&�>�!s�.J��5�ȓx�F̐0�H�?Vy��Y�3<H�ȓD��`.�D�p�ȖD�"���ȓ+�,��_
i��9�/̟�(����<�cɖ�#2΁�! �)v���o�N�'�?E��ɞId��J���7��S�l*D�x�/�$4(��[�(h��P�G�'4�(�A��g��Q�.tgrQqD��J�<�b���0Lr�)�jm
q SD�<2i��]O,�SŞ�t�Ĥ��,E�<)d��]�ŠC�:Lzp���C�<iV�òER�����*��lz�Їȓ@�8��EO�W�z��0g���^)�ȓF�n�*��Z ���W$�YM�D���}Y����7.�7f�.L�6B�ɧ#7�-2֮ڽ$��ԙ�DF/fB��<G�ֈ"��K�-�0	��aZB�	1w�����L�i��:ƍ��|@B�ɓ�8=ȗ�θWitB���Y
�=��'6>�qP`8'D����A��5��1˂��-�C��� 4k(/!N���^�t�Ռ͸[Ͱ4ʆM�:Z��؅�]ސ)�b	�A.Q���<2��ȓ_�xE�V6�;��ڸge&؄ȓ[m�՚��\@�x�W�Q8�U�ȓd����1IZ$f�&��'ֿ<��ć�:�꜁&���'�FU9g�I�u� ���؍�S��q�$�өU�m�tA��S�?  �zB�4jX������t	6�q"O��k�kC�`,�	Hp�X�$�Ne8�"Oh���OX;Uj�Q��o�F�N�Qb"O\q	bjπ d�c��ڂgd
T�B"O P�2�֖s�!�f�x��"O���g�ٻv��cc@80zBE��"O�ȓ!�Q+��j��Pbxj��a�	L>��L՘=��	�u�t� �bh7D����Fֵx�Fy�!��X�4!���6D����+�@��@�P,|v�lR��2D�`�!�ח"�Z`I�
�'o0�p:��/D����!G&�@��,ũ2�H�۔�8D�t�#�	yK@|��E�n@hȠ�(,�$(�S�'�����`׌bMb���P�RuEB�%|�LC#�5�� �cℎ:�fB�	�6�<sA�D�n���c3���C䉤{��i�TH]5F�m�.#]� B�	";�:}Ӓ͋�0ѺpI �ҊR���=YL>����b��gw�� ,�5"{r���i�y��k���5!�5L�����yb�;x�`� �釔�Hbeh��y�f�@Z��ǁ'kf4��Uᙘ�yr�-)�i0eh��q�e�C��?
�'�#���4����%V�:I�	�'۰���l�>@[jL��P=nf�ۉ�$)�n�W)�d���*5�J<2C���e�'��П���Oj�ɪC?$���d��E�b7N_#snC��0p!�Ihb��e@Y[��� N˓�0?Q%��*Md�ػ�IR={IP�R�Th�<!u��6�`�rS۴�2Oe�<�A�6~L���DF�D��4��j�<5N��iB4 J0�?ɖ%��g�<ٕ�!�R�)C���X���J�`y�'��|��������+�;!��aKF+A��B��>d��A�v��P�X�*����O����D�=�8 ��;��D�&�٠R0�)�c�ܥ���C+��C&��$�f��'����WgVl�P����_�����'�T(��ƃ�r�d`���\@���'�A{1A �Q0�ͲfiA�X���+�'?�=�5�>Yi5A�"ӆRU���
�'���'#]�&�<DrV`ٗ~����	�'��IS��Q����	�"+'�Z���'��� ���(���!?�Ҥ L!�Č�D����1ӚMX����1!�Dٳj����h�z��}
pK�
/!��^���r����NT�״d���'�(�@�Y�6Q0t��'+��}��'���T �ˈ�CZA�!9���C�'�a�ԡ]�(���-�&3�%HA:��>����?ّa�2C��C���h��g����y�f@!} FM��σ� �݀�Fˤ�yrٰ[BH�J���T��ȶ�2�y2b(o4LʧS�@r1CJ��y�BD/vW�5����69� �Ѵ�ٟ�yB�^�\/�y	��ԯG*�e�g�F����?I���� 
xN��3A$�8�0r�`�1�?��'y2l3�^�iw.�2C���/�?i
�'�����4r��y�c
P��Ih	�'^��x�K�m=���B��HR������hO?=�b�F�F��yU~`ޡ9�F�<�%h�!P�,�!��2�����S@�<�Q!L�;6č2coӉP���s_t�<!�ɔ�$F����ވ	�´��K՟H��S�? ����ےR�]+"�%Jmpѫd"O4��2�K�e�&��G���>�����"Oࢆ̵�2�	�φ���=�1�'�������
�&�h+�1��<��q�œ�m������!��\(��ȓ�<]�Њ�����5 8�>]�ȓg�0\ؕ���9Kf���
j���L<�Ā:D���$L�$Av=!s�F�<��'O�`@�AK�Μz���^K�<irF57������-"Ԝl�d̚I����<2l^�:�hB�A�$;I�`�p�G�Il��$�Uݬ� 玬o.Pt���!D���b�Ȇ6<b�!'& �x����I;�OZ�o�*R���;%��C%A�'9X���ȓ#�`e*U�Ymb�0v��� Y�ȓL}��X��X:+�r	Q.o��ȓ@t���uMɿb�HUP���Ow���(d<��HzH9U�X*�����'�����ך]jDI�����h?PA��'?ı��J_!5�0���e��= �'Z�,¤!��Z&�T�b�L�V�ΤK�'�"YR%�$�hb�,�b ^a��'�>X����T��)c�!�	��d�	�'�5�/
�"���ܲ����hO?y���7S#���6�*YRL�� x�<����==*����2iZ��{�@�}�<��j��/j��t���~�.MѲ/y�<��l׿}3Аy�c
|�� Ф��s���0=��M�/E�0p�&�
`�p� � r�<YC�$��<�f�;V.i��H�<�# E8�*�Ab�H>{<�a&Hy"�)�'l~p��� ��KG��0D̰�ȓ.�<�䄁::��k�-�%����n���E&Tvo�[F�ޢ.p2}�����'�fx���l�6�,A�p�����'��>��$@�Ļ�dJ�O) =H1��� �I�ȓ]^�P 5�;E-�P�r��6��4�ȓ�^�q�'��+8�8��c�F@������R��#g���1N��P���U0�� �o�8u�Q�0*�ұ�ȓ�\9�Ft�,�뇨�<��q��=��K��=f���D�R�c܆,��i��	@KZ����ӄH=H�pІȓri��-c�	:�aI,Wَ�Õ"ON�Za��L T�t��Q�����IG�Op~]cg��-Nj� @��X�4y�
�' ���C�5~X�w��P�j;	�'����%R�B�^S"C�G�`���'�f,�p�&yg���g[�>� ��'!�Œ�d �E{-*ᄙ�9����'U���`��i�X�r �G��j���'&L`�I?�!�4�^MY�q�'���ӕ�س%���H�m�t.�K�'˼����!]TdӠ_�q�� �'���	P�ʇ*��)RU��j��1����?qpφL[��ӎ��J�����y"#_�T[�g��Q��]���y2c�]�r��bK�H^��O^��yB��!
9��e�E;9��������yB�ɭ'����ČfﶝH2��6�ybC��S�	��nBV�Ġ�Ѩٞ�y�&Â(=j��snԮO��)ԉ���x��y�L�Oǳ?���5Օ��Op��2&M�pZ=�e�ٶ*_��"O� ����"�@p�RG�ޭ^�#�"Oh5���D�uH҅��`@�_h�i �"OJ��@H�;�t5�A/K�neZ�"s"O����KmH$(3u�ބL��a"O���n������D ѿ':���S"O�q�6ş�=?`%3c	�<4f�p'�|��)n��1 �,I�w�yeŇ,�C䉹<�����8[�0"2�XC�ɊM��i@���9�� X�J�n��B䉋K��d�ԺJ���C��~��B��x��ʃ�&7�F�a�]�h,C䉫P�>�:Q 6�$+�㐉#.(C䉒'�
�@7��4,P���C�\�R��?A��OI1O��	�� 	<�a+%`ȇx�=��"O��`"��t�XU�¬ưn�Qڠ"O�0��1N3 �x� ��2w�xhp"O��� NFR�f�#g"�>uk��k�"O~ݩ4c��;u�l!ōvV�0$"O�yYqK�K�>��/P*EP�U�"O.�1c%�t����-ɃOG���'z!�Ĉ��C�B<%�TQ�ABQ����!�'�A��LP�j���l"b ��'~ҭ��.��X��|�(�Q��)��$4��dF��/ojYD$A�"�i2"O��!��E ?\�吃�S�'����W"O�8�S-1�=:e��T#B	�"Oʽ�3�=4T� �T5dn�m�E"OB�� �1Z��Ĳ�&!iv�R"O�݊�[�Kv������VZj}z"O(���C#c8#�U2=XN�q�|��)�B.qD@�=p=�b�Ų"b�C䉍La.HBd��*"�������4p��B�	�
�<J�ycŏ��n�xC�	�u�F��Ħ��B0ΔaU�W�/�FC�	z:Jl�S`�NN�d�R䖁�>C�Iy��٩�@��p\$ u��	iC�
����3�Nvw���K,Y`�B�I5���ʕ��)��7�ɸ_h�B�	�wiY�	0p���8�'�2*=�B䉳Ob�M����x|�D���X��B�I�d�*Ѹ1c@�&s� ��:6ٖB��b��)��NW�5V�b����6�C�I�%�������7%>�9�d�o���Ɩ7h�0�')ɶ#�LuH�l݀d�!�d'��tr�A
L���`�3`yў�����R��Q�܌[�*�y��U�!��B�/BIJ��KS�����ZF�B�T�&���&��l�ܠ1�Y:>[�C�	#`Vi!֥ 3'�
�|��C��
u�$�O�'��ҧb�I1�C�	%�Ơ��ʓ6��A��">�(C��Kz��R�٬Y��͹!N9'�=i�'p8X��U�Hzzcw��	Lp�ȓ3���.<}F��
u���oq�Ʌ�)���*bӟac 5�7㍸&r�Ņȓ4,�����1\+��Ġ�2k�|�ȓ$���0OÀq����L�FL��ȓ}?R��%Ċc^1��.q-�ȓI���5Ν���k(I.L*�D{��O�r=�I�HQ��[����^Ƙ��'�,q1+E��5�a/MA�p��'g�a��m�|V�A��%�C+ �S�'|X��u☛W@z%�0��0J�)�'������.p��=J�f�-#_I�
��� z�J&k�:"����F����� "O�"�ݐ����d�P{�|���	]>I��������dHe�� 9��<D�@��(��N���bӌ�M�� Q,9D��r0F3"�Pq��
)#Fq!G�9D�Q�)@�\��Sq��Cp}i�#,D�0{�(��"��	�r�z�w,D���B��	ᐱ���Ԑq�LQ	%�.�O����@_����	wH(�{��W`"�=y�'gf^��0��y���f�\�M��C�~�c���8�2pа��!n���WR�\i�F*Hj4��m4'�i�ȓ q���V;��L� jZ2 �d���[7�T"�@Q�y����1�Q�ȓ�Ĥ���Z��j�cd*}�X��I�<�r�L�Fj�H�����̑ђ%RV�<�/� g0���@��橕y�<���#+v��D\��>r��~�<b� F�6Y��ɐ�Q�8�	C��@�<�������d��j���i���z�<��dίU��) �b��(Nh�0j�z�<�fτED�]9jћ2��� "��w�<qT@�5~T�Y�3�]f�0�Eb_L�<!QKp�8@���E��x��'N�<����I��30)�o����gH�F�<��K}����!ڬO0hU��[�<)QG�)K�5pg�=8'��ba�_�<!Q���)��i
�ϋ��8PA��C�<����Moͳ�ꎚp��p���Cx��Ex�n��h�E�^1��۵Đ��y���o�����O3Y��5����y���yZ@�3���:�5�tF�yb��2't��"�܄��}�$���yR�W�5�0H��n�����ʣ�E�y�L[�qCjp��B��,��� �ybEA;��NX�
|}��']����hOq�����n�*H�m��W.(�T��"Od���/�;@���9a�x�9���'�!��
����E�}��L�aoߴ-b!�$E�X�z��ChӺZ���c�,DH!��0$lq����^����]/@!���&]��p�Lͪ9��|(���U-!�#UI\�x�HD(;��I�B^.K�'4ў�>-�Q��X�L�A↔�Z��h;P�+�����B���c<!��jB��\�<9�Ϥ]�dp����+W$��a��b�<�Dٳ�\��ĎN��ܡ{1�N]�<���Es  ����8`?N���+V\�<a��Hyj�Qb˶`~�d@& �T�< 	��D��cG=�x�F��xy2�)ʧ�.9Ç��4Ndy�$����<��t�,�Bw�S7"W5#0g�6�a��/\�t��N�(y"\B/�"9���r$�`���60N$m��?u� ���
���G�Ki�E7���*@��ȓ?�D���N,,���i��2By���JA�B�&h_�=�`�	1*ƾ,E{��Ou����ޚM@>�"ǜ�kP r�b�'Q�>��f}��w�Mx�X:4)�:Y�",��]�h�p//)��Ղ0+ҵBUh0��xI�1(`��2s]�<Z���af0�ȓ"���w)X6�v����ƭo���:��q�"��OX�ٖaM}=���X���h�C]蕰��'�����b���	0�)� �䈖�_�Uo6ћ�@ЌM�~I30���O�=1�'��|�7/M)*�	��&ùE�H���'W��59}�v1t�T��
�'�Ti�`H�.on�œ��_h�B�I�P`�P���"����qMݯ>�B�	�(��p��pO8��S��6|�.C��(9�P�X�㍳f,AᝇS"C�I:;F*�[a��<|ʴ�PKN��>���<I/7�D�@�C\;$xDCCJ#�y��F
 H��j��͆ߪ���y�"K�E�.���
	x��)�1�y�DD!]�m� ի8� ��G��yr��uDd�` 2:K�\��Q��yr�GR �I�6��!�q��@_��y2%�k�@�K��2%
���?a�H|P�SU��j/�zU@�;3��z�'��Mp�D�&�ru�d�Z_|��'�^��a�U�<�VmۤHѵ��4 ���<�̈�	>=G�T���LP �"Ov�� �D�"{��d��V�J�*!"O0�(�Y*�]s�A�%Q\Q+!"O"�P҄VOg���v)���!�"O�@�l�62&
c�����ɨ��|�'�azb/�|6n̊�"�=�"AB��-�y2��9^��7-W�.}.�kf�O��yb��*f�}q�*])�څ0���y2�R(p�)�v,O���Η�yB�B���Bs/B���i�R �y2-XT�hh�0v������yK�7y����H[� ���MK���'�azR��b���ш�}h����
��y�F�zc�SU�خ"�B�&���?��������FM�03�2�JFN�.��@��I~�<��&H�p_V�1�ރUd��C)\v�<��M�3pv�(ہ�RX����4Br�<I�Q�54q ��?��1����c�<�P��+BҌ�VT�4���j�mZe���0=iA#W�YDh<H�J͍ \Z,
�k�<y�nO�}ѲmPt/�f�b}!��h�<Y�o��$0�0J��@"`�$�b�<��'Қi���d��D��! �[�<��+�p�~�dd�e�,"�J�C�<��)I���u�M��T�<�u�T=^x�0��,,�K֋N�IF�@��Ǆ-@ٵ��6X(��Y��&D����l����a���ޒ,V��{u$D�4�3�_�_b�*���~�T�� �?D�4Z�dR��[�ےx� ,�'�=D���vB
3\N��r m�;fN�{&�:D��
��L.c% �Q�@��V�>�`7D��Zuf�$��ĊU�A��X���5D�hN̓pd6	�a
�U�4��a7D�4�#̷+�F�(��&z�Q�
4D����@%�~Y��H1��	�2D���Af��v7�����-���p�!$D�ȱ��7r��q� d@&d��УB�-D� ��A��%��<)I<>�V��D-��W���ӊ,�X;�ØR����6㗥HB䉞I��X+t��M_�]C�'$~�B�	)�Zh"�G�X���W�BR�B䉍Ta��{�� �{����B�I*`���->	�(5�a.��B�I�s�( PbI)oQ:���N��B�I�8���9��x�@9��&�e�f�O��G�� �
�H�+|�4y�g]�"��y5"O��{�MC#���(!l^��ax "O(�
�ꑶT�|q��Ӯ?{��q�"O��PSd��Y��%qpiգ=c���"OV���b�u�Z��0�N!I���0"O^�d����1��&c84��"OL�:�f�1j�x����
(ݐ�"O �������Nr��v"O¸  ÁK��� td2���"Oް� �W,@��G@b-\D�Q"OB�k� (Jo���ce;u���"O2�����6/�>YC���6V�`��"O����,O5"�pu���w�����"O �x�)�*
+4d�P��c��q��"Ol�SU$#y��2"_u��%��V�d��	�>���mN  8����v�B�IFAz�iR�ÿ]�@$㒠�0�,B�I�4>Hԛt��mE�C�6O@B�I�0m�ps�T�C�^ J`��/;jB�	4��IS��aJH* ����C䉧	���u��:Aj&h��g��,C�ɣo�ƈ����'��*�*`oZB�I$ ߂�a�5��1�bt�.B�	����홸~w���W(��B�.UDl3ԡ�n~�YP$�$�B������ODr����JU8B�ɭs��)#-�& ����p"�i��B�6�`UH���G�\)�H�]ȊB�	�gT2�¤J�z|��\�@LB�	�a��A�AA�,\&� ���>��B�I�+}LؕG� ?�Z��6�B���j]0����1°�V>?�B䉱b��%���CV>j=�rg��=D�@�g��z�lɩ���E�Ja!.D�x гh�Ƭ�7K�)�p��SM+D����ǁq�D¹�yt�:��B�I�!r��b��?m�0I��N}�xB�I�O�0$J�J�4�4D�f�U�"B�IeL��WH�!(��1�c��C�	6Ȥ��s���OX!6E��|�B�I�y�d���D�X��Ő��^�*C�I�Z`�4AS9�z�ȃ(Y��C�	�JdF<H�(ю ��az��R n<�B�I�5��ᖦ*r����p��C�I�2ƀlyh�HfrD��ꚙ7�HB�I/3��KI	]r2�X�5��B�ɩKET���1���`�|B�I���`�! ���"�Z!Y
�B�I�l��9)�FM7�8@�L�b�B�%fn��B�.�u�D��
DC�ɞ(�xQ��]�b�t�s7�ZL]<C�	U|&\I�ㄺF39ҦMԏ`�0C䉲: Ѡ��ԙ<�����'# �C�I9z4yAB�B�]+�hҺ]�C�	7\�֐��EJ?IY��VD��>�tB�I(Y*�e�Q���6�V\%���D�B䉘)� T��b�*&��dl��[�C�ɤ�b5�Е�F�b��ww�C䉅��mP5�D2e10jVd�	 �C��&aG��@��^/������ l�C�ɶ$s�!��$&(r��Ў,UHC�	�|w������=�ĺ�P�2~B��e?,]ѧ��B��H �W��B�I+�pʒ��Q��qb��( ApB�)� L`����5^(�� �J�QS
@"O�����M�v���B�����b"O���� ��S�2�@�䔱Rq"Oh�q�@�&B��"QE��Z�n�Z�"O�X�F`���6���C�x�]Ц"O�E���]`+��!"u�1�c"OF�gJ�i>�H1�ǅ�m扲p"O�eR6���F{<a���e��e �"O  �� J?;�vl;ԯ=?�����"O�q���=@�5�g���T�q"O��h�턍� ����7x1� �E"O�)`�=���ԥ2:Α�B"O�DG�g�D���K��`,� "O6|�⏝T@�S��`�R��"Oi��䔸#��E�0�Q�<�NU�"OTma�kO.f�p�s�ʄQ���X'"OB͛w!_7"1��[���"O�P��f$(҈�F�G;J(.ű�"O�A `*�.9��k �C/&�|�p�"O���QE�@�$u�s,� kC��"O|�;�a^3����O�:S���T"O~,Xtf�/ JJuYc���]5��1�"O���C�R�L�\��&�@�3zia�"O�}�� � X��K�aUl�"O"!��̫�b0˓#"�"O��ˆ�1dz�X�+r% �"O��8 �`�rL�D�c}M���S�<��J��>��<�cT [�Y�L�<	����(�����!>)yHp�E�c�<��	�2��|b�ܱh�>��ե�a�<1�X�[6>�B)J�v�ҤQ#D \�<9C%����jp��&���A���Q�<�ÀN� !���_�q9hYqc#SO�<qg��,|�Lp�V��=�}�u,KV�<Q1 �!�v��q`��<��P��N�<�`GȖ#_�8 ���
8�L��k�U�<I6��Z���w�}�����gU�<��N\�R�Aψ'��A�I
y�<�q��8~�TE1�m�5�@����x�<���R��J	@w�T�B��E��F�t�<�V�S� �e؅-� v�l�s��[�<��>Wvz�I�E��p^^Qq)JY�<���1dLlM�t޻r��6E�R�<�'�J��j#���=5��x�<��Q�d���GFWҨ���t�<��	E@� ��hƖ �L�CQ%�r�<�0	C�M�(�"���<YY����h�g�<�e��4d�,�ZdF�&���\k�<aa�1Yp �fC�%���V�SQ�<I�G˪��T�E��y�P&Dt�<��A7'����U�M�����3�!�$�	Oo��ɤ���UU�y����4�!�D�1в�`��� 9�u�Pl
:�!��W�Q�L ǚ�2�\(�ʼ".!���uc�p7��$0�����E!��&(6�C �'����g
�.Z!�$Ǣ��K�;pn�I ��B!�DW7`�s�( Q0z�e� 8!�DH=-y��`�U1������]�!��noR�	�<�&����ׄ0�!��V�v���c�b`J�!`���Q�!�# U����uXt5��mZ�x�!�U8���� �_C�и�L\�Z�!�$-�٣�B$vZ�P�
��3!�� L$RUC�6V�(�*g&Щ~\1Jf"O���ұq�0����ksHѠU"OL5J��];�d�c_=rࠐ�"O%qvL y���aײn@�ըd"OT���b%[���:�V�8n���"O�e�p��ba� ��NƎt��,K�"O���χJ��qz ��Y���Ib"OBQ�0��Sf��eA9?�$�Q"Ol���I�.I�i[��\I��ӳ"O�:�-�e�ĸ�c>|�"O��id�ȸN����Ϙ�YS�ЋT"OF��׮�~�4��h��FS8D"Od=!��\�qq��E)�LJ�x�S"O0�t�ur$Yc6�]� �$�"O�1v�˝>�ZXe*���x�U"OX�k%��J�k��j	#���?�y�茵*��T!ˆ�Vb��°����y2��@A�H§��U�<�����y�L��h�J�z��I�I�"�Щ�y�`K26�<�DH-CO.��b�چ�y2m�9�������@Lj 	R�$�yrFM�\�D����͎��{anދ�y�� H6+�VPh8�U,�yR�N+\� HW� �I6�0�a�'�y�,HS�D�� �Ev�@�'^��y�Ė%M�M�s	˞|���Sv���y⦈:�h@�QI�$;©���խ�y��~H!ȵ'S�d����쀀�y�.^�V�"=d
��}J��;�y2E\��\RF��46�@I���̪�yҡ�d���7A�a��#&C�	�y���457�xZ��^��pYd���y⨔� ��xv��y����L�:�y�i ���gA�Bю���/«�yRD͈\{8 �d��&&��Q�ݒ�y��Ѷ@Hd���ݭ醔1�Df�y��2>��]ɴ�	��&ᘷ�yB�<
K\ڰ$ƫ@je8���;�y�
��tĀJ��^�&�"b晌�y�'�xJju�c��jp���"�M��y��� v�svJ\9a"��	�풗�ybW*�-��@_-p�B�zTH��y��*3jUc5j�;bK6i�SeǗ�y�# �YO�iQʋ T��M����y��Rvx�i�'K4�j�־�y��LN�yb�E18�yy�h���yg��8�*��+�-� 	��y��6�&��c�1y0��c�yO������2z� �A`O�0���ȓ�e@�(��)H�`	0��1W\�4��Q���ƮS[X�ct���Mָ��q�=a��-G����b�*X��h�ȓ}Tn�i��D�Fp`�b[$,ez��/d� 
��
=[d��f��%�Jp��5�Lj��)VQb��ٺ��ȓ|=@�S�4TBhcU���C��X��6XD��ˡ*��z�dۓZ��8��i��K��#�f�:@&D�>(5�ȓ�8���A�,I���2`]�t@\��ʓ?K����F"�
Q{�KJ�}�C�	����ۈy��8��	�T��C��$\@ApSj���81��MjG�C��g���Q�_�e���fL�G�tC�I�2��9� �[4t0B���2�ZC�)� ��3B��9t�H#�M:=f Q�"O�(�C$C7wRE�F��Vl�Љ�"On�j�hT6���0�� ^�eC�"Oj�p��qoRa��0��S��'�ў"~�&��*]�K�D};6�9PRL��Ua%�7�_Y��lCUj�:{T|�ȓx8��	��ɻ|x�!�m6Ȇ�I��DO?GƤڷ'[�na9��#�!�A�,�n5B6j˂i�Й!�!�!�Dŵo�fe!gB\�Lެ	  �U�ўl��ɥ����4�T�z���H-��|>��:�S�O��zǄ$N8�
��.�"OBy��
�H2w�K�Y����"O��u�H+8��;��ڴ�d��Q�MCH<�2@էB����٘t�y@�O}�<A���-�����)p3����d�<�F��8��܉s�ߪ�����J�<ɧIY'"�� �c�&��C�j\k}�)ҧb2P9�k؂��IZ��I6'k���'��~��:L�H���dW�F�$J��6��:�O4k����KR��H��$�4 ��"O�\A�F�_f`lcC%Y�]l�Y��'D�'uհ�-M��ha{�aJ�W�.���'i�d�_�z��d���� H�h-)��
6�S�T��K��x�窑6ċ�G�!�y"�g�\đ5����������y"��J�l-�E�D'Č�Ғ����=�y�cp
���h�,C���I [pzC�I� d>|���5��x%��h����ĝR���u��3dƅ��N���Մ�[*�qDO�#�84�S ���zT��~����S�ORn�"�A��hPqC��--" ��'�D3`Ō�(4��^r7��N���'Y����	T����m3.ʨ��G�KS�C�Tk��H�@�H����ب!J�C�	�;	����[�m;��0A�Ҵm	JB䉘��ӱjB�/�� �p Ҕ�6�?)����!���1��"l���q�]�!��:8��1zV�z㊽BM/May2�
X�\h�#��	ĮY*6� B�I�~(X	�	�� ʾ�¡�/�:���'�O?��W�D����<�c�^� �!�U�Dl����+]�ȕjJQ8/��'�ў�=��	C���u��hzj� $�`��'��`���"r,��/C'J�N���!-D�$9�%ǆ�z�H��Z	x�6�5����	������2�M�1��hzB�	�{dBAX�N�;�t���m�
6�h�=�~�N|��O�$R^{��D���"�<Q��ʛ[���A3��}JƼ�ծz��e��=�'e�H�)�%^��:�'�"�za�'$~!�=9]�\�� ��WjE�W�= �
Q�#�x9O�}��W�:<k�Cj��E�է��jJ������YB�X���`��I�����	"�a�Ƅ�q3�r,*}����Ă�7��O�23艓F�z���h�<a�\ ���I�P8����L��tZPq)c$=��"��$�ƨ�vl���z@|����A!^&��D"O��Г�˚p��P�W�=M���<Ov�'��z�Y�h�� ��^�jw��FE���O>i����?����u�1(���5�1��B�	\�ƹ�F�]�Q`l�s F7 �ꓔM���ᓟq�*�J���I`���f{�F|!
���'�4���\d|QK䢓���+ٴ�hO�,�S�? X)�a^�hF̋�B��1�P|�p"O*��`�3��UbsB�|�j	��"OX}:��KD?{��˾"���0�D8�S��vlV3U�¬Tv(M#��T�L��a�����x��+�?#���b�1��9��	h8�<hreH/����PJ�.A�&ZWX�x�'꾙�u�ҼYԠP&�2:S��'�ax��d/>�hHY��-�0D`��V� Tў���~��ɟ[��0�"�XXt�� �DD�O�=%>�t��d����O�'\��1VM(�	a��ħ��y��WG�C��7u8d�=��'H�x�JCqp)�mC�e	ܨ��	�OZk+OR�<�$�3zԒ���_6ܝq���_���=����A���Y�@�4*j��C�¦�������X��Ӛ}�!��Xo���3Q�"�,@#~j�Γ	Z�r<:'GJ-<
��h`�v̓�?���|"�B��6ݳ�Ѿ_nxlq�ؔ�y��2j�@-J��������'#-e���^ �`�B֤��(N�X�Ŏ�2+�!�D Z$B��t���U�
Q�1
Ҹ1����P��s�E��sJ �C��	���'���D��,�C��8a����j��YZ!f���yRF��L_�Ȣ��6\[�UI�GΚ���hOD㞨&F�z�4��ǣU�
L�� �9D��3��ѨG_�q��ϒ#pP�����8����0=q&Z�j������	T�L��3#�py��|�?�JC��;��}���T(*��5D�,i�W�d���-7,J�����K$��d=CL���U�O�~�HlB"k��H�a|ғ|2׍5�pl)����u���Y2�y��'@NQ�bGI��sE��F�0��I<	������Oh�䙱�L"�>�;�g$��!	�'�}!6�c����D��
�N�3���i�"~� �&��wlBc=����^�A̲,�ȓ@���p�;N`Y$-J��P���s� �Ń� &�L��㜺
����#��0|z�͎�P�"�Y���m�B�K�<aK>A�4�O�S
RŌ��J��:�B�S�MW"�T�X��)�e�	�,��I�P�U\��{�MʔB����:�S�OÆ�Xq�/{*b$څ��	|AHbr"OĽj4c������M.^��A�<)Ó?�D�'�=�T���mV�e�B� :���	�'��ph��B����sj�-/d쳋}��Od����",.�������i��Y�'��?��ׅ��v�Y�����ԁy�j��W�)��<�CT5!�L4Rb�"� T�^��G{���iQ��A� ͱ`n�p��*Bb@�ܴ�~��'��y��"ĵ� 4crNT��T��OV��$^*F�Lg�?:�ԩF#N �!��=��Q#�KO3U4�ȗ$���!�$�%BR�� ��2Hj���:�Q�,F{*�4�&�̠\'��BA�22�h3"Ofp��*�Y`\��U��a�(OL�D��ORE�r�.�ʖʏ�*�Ѱ�"O�ɻvd�Ą�X0�B�]�&�"O��9�	�}*8��%a�?�v 1&�Iw�O>���BO�� �H@���7[S>e:
�'�U"���z˞���[W���ə'qў"~�MX�*��ͣq̑i��rug�F8���~��*edzH����5y��9�T�1�y��	���%�ٸvO.�p����HO|7m&�R� �'��"9S��z�6��������ቯ]%�i#�)ݾ^�标��4"##	W)�E+�h
�7�f���S�? �,@�E�}"<`��M�Q�����"O�\B��@�Z�ҹ4��*� X��"O~�p�Y��zq0�'�Z�ȩ�"O^H��S>����N'KV5�"O�r�nēC�`��.Y<cb$�w"O��
q��an�S�+V(	J�0"OrMkf�k�yb笏(9�-��"O����L�Q`�������W"O���̍cX���P��W���G"O�$�'�
f� X�D B� �Aa"Ob���*ԑ$�<H�4m]�E�z�;�"O�x��c��Bfn<��V�B�U�"Oj�b�(2#��̹�d�B� ��"O�	�'����е ���"O�D׭
a�d,	bk��t;�"O���p��7�X���ٽt�9�"O6��f��?;�0	w��}�&�p�"Op�9U(c"����29��	8V"O��j��M�,�	#`D��|[�"O���q�i3
8�b��;jH�Z"O>����_�Q{w�L� bL�"O��ɷᝄK�[3s H +R��A"O�q��\z�(��H�;@f�:"O�ɛD�@?[*�)9��
�W#N�a0"OvP�H�=G�l�� �i��MJ$"O�l�MR\. RQ� �H��"O�8��f)p4�3��-�"u��"O�S�cĔVf��Xg��G��u��"O�B�,9��[����U"O:1�Tf݃#
1� F׷$-z$"O�)A`ԽN/ y%C�3���y6*OV�Y3�+g�8ly�+�=r��
�'!��ئ��/^l܉�F�?Si蜺	�'b4irbP&K��U
Da�R�[	�'f����
#qQ��ό�;�`a��'�F��D&����z��w�����h�<���I��T-* )�:_��YJpPc�<)�NE/#Y���&�ڰạ���^�<	!�B|z�o�a%�<CፓO�<�t�מ6Qb=�Pj�)H�AQ �Q�<�c3���Ú|�1I��K�<�A�:�V��#'��8�Z���f���� �D�:}L���M�M���;qM��4� �b��wj�ԛE�&D�8��.[?	b<��Ӭ$��<�a'D��0����-���p��E��V�"�E%D�l[�+�5	�l��Z�a��/D��+�FS�F��I��v�,D�$�*D�� P�m.�r��S�N�FԁF#(D�$r���S��!b�G�q��D f)D�<���u%��{����dAA&D���d38b�ѾR���i�)D���5��@Q�5xUF@�Y�p�c1D��!���"x����)I���I;D����"��hR��A͎8�6M��"8D�`1T遂|+4�!}�
�ۆ 8D���7�_,!SX�+H'V�6D�PJ�<��(��ǩ7븐�n D�T`�,͎@F�,aG+ŘB�����%D�x��	�)2	�)2�B�LpZ��B D�l8�U�C�@|��a�:%-L��G�2D��00�H�@��#����M�T�Ī2D�L����$G݊@rD b��]��N"D�|��A5�� ��~���:�K!D�L#G3Wt�hɰ�	8���H�M:D�� 
�f��4/���(�ܔBr��u"Oh!լD�d� ��EW"O��s�"O��󢎑P�
ĺ��͏BH(�2w9O����,�p>���0
�j|ӳ�?r�ƨ�5�]���3���XW���.�h��4Dq�2�2U�V�/ؘh�ȓJ�d�i�m� m�L*�K��B&��>�FJh$!��-ڧ1d���' �xlj�.hn�A�ȓ��=ql�c����3\�h��|i�\b�j�(N��ي�Y���"�C#r�����!d��4��.)D�D�צY]�ҸCݴwx���T�{�� S+^q".���/PNlB���i~ �c�5蘇�u+��9��ǜq\���,��L��m��b�@����y��B)s��Չ���3P
��!ᭈ��'rBd{�G�)��aF�T�ۗr|]��iȇ�������y#��AUF�R�KF�n� V .7��H�e�+w��?X�>�p��� �8��+`��S�ظ�ȓ?~�w��;,^<��R][���o #��H��uY�{"Q/;�֙Z��/w���IƯF6��=y��f�bl�'�f�P�cJ2���b��J"Z�'}lՠ�G��ڬ0�e*۰L8V� ��$G
��Т��I� @��G��W4R�0i��{�!�DL�(���G(��.!lQS�����!���RwPy�5T�V�0����/{!��"����ʵ ��A�wkB�M}!��ԮM1���d
��"$�[�WR!�DS�	�mx2"]�K㈄aԉK�|L���Z+����w�Ͼu� ���%��y�.tZU"���E��E��+K��y�c�%%g`� �����ӑ�Ɔ�y'\6�X�{Vhq \��F��y�ƚ7xh(�
��~D(
6���y��I�z���BiI�h�ҹ�����yb!==������D-c�Zh��:�yR�ƯlV��3��͊ieJ���y�D�!�b�q�>lz�,���y�+N��)5Z�XE��"%K_�y�NQ�D4��A�I�:\�\d�C���yR뎩&a������Bk��3F�Q;!�D�_��/{��M�dk��=�!�DJ,6��g�V}��ivK/D��AY|L��
�������'$'����1Lx~��I����್Xf~
�U���RcNL .���QM�~�<1'g�,}*����ڠr�✳P`Q�s� �>rs�?y����Hex!�VA] ��=�u�=D�`ZE�A�raֱ����	����Vˈ�P�48O�l1�S�g��ȺR�u�)��s�p�!6}
��J�RW��`0 >3JNe�d+@-P��aեO 	��#����?3HJm�L<i1�R�6��� ��o �	�g��@x��(a�)h��GZ���	��-WMQ W,=�$�'<�$��$]p�iBo6��iM�X�c#mٔ*��y����;��'��e�&e�8���&?}�ƥK;��)�>^k�0;g^����DG���ϟ/��I�M1|����|����L9��Y"2���&� $^ ����C?}B�P N�d�	'񉚡�l)��㓫z�.YP���v���'�GZ��w�Ӓq�����c5��
c.�*Q����&Xf�'V�d#�'L��  l��\d�����5&��h�'[@1hA��65z4] �e�:v.�ӓ=�&��b�;��$U$�X�R��Q2y��Y��-��
,PM�p/U*w���'}�~����>��ҵI��� Aџ8��qW:?�6�G�������a䈅r*O�e��N�*��S�
�V2 �xrB�"hY2=b%��Д���g��& B�'0�5C1��JJ�D|�I͑xex��BL��b�|��[���c�\S`�ڿ"��4���ƙ*��8N?�r�԰�8ِ��ʃ=B��Tl[Z%���K�a~�"Ҁ^+q���C�D��'�*&':%�u�%
3"t0���>~G���O�<Y���Bc����'9�=��t�LU9�˕r/�h+
�':x�{T-�+K;�[؝c�m�!r�+���(N1 �Y#o�;cӊR�x�ޫuì��O�5��m̈3Q�41�( �v����'S�(a���+%�x���_��� �q�I �v���&�)b��D+c#�5��'��L;Cc_X�'cJ����F.,
��Y�#9*��I>�!Y�&3>��a��-z�r@bP ��O��@��pǒ�����%�Y�	�'��|�D$K��`pI�q�0(L�J�j�a�����e�1���O=�ɵ3������Va��'샋m+rC�	�&s�-��¤p���'^106�yr���"�,H��/hz�s�'�2雃"_Z\x��W(�oݎ�ד������O�	ۄ/N�K�t�!	�	`�ؕ��D,�l��'�vܡe�\, �,(�h^�c��:��Ď-A�h�E� �ӫ:��9`�!Y�S%&X�wDٞf��C�I��TmG	"���Js(�"B���ɧk>F�E��BX�S�O�J4C*5�=��"�|D��'�4H��sM���%�"j'9�M�lC�KE-@�^ R��'��:�ʑ.X������ۈcl�	+
��zǄ<`j�;?*�ڑ	�/���@�*2t�˓�2�D�i�W���Q����rvႧf$��1�/X�fJ�c>́"�W�}/�`d�ߞu�<�ku�%D��qg�O�NWĤJ�o�
=���s7��|�RfT�x�B��ԗ>E�䣊<M���P�şh(D,�sM�9�yRh�5r\H��^(o,R(�Ӯ����	�R�H� ��q�ax�C9�D�3���owl���Ν�p?�S��~�j����	6�D({�e3���b���;[bC�I']�4����V�B����A�y�|�M>�����{�֝!Lg�}���BB�i��W�?�����! �{�G$��J�)��|8a�2!0=����OX���N͆�n(s1BS3ɸ�(����G$;Bj�ӣ��n� Xi5�I�]�Q������O]��c�Fؐ	hX�e��9՚#�'�t�+Ʈ	}�\�!Jk+O�IC��6y><mPp�-����L�Tf����ˈ��g"O|�V/^'|���`�'"� (����.c��� ���b`�|�3�I�h=,�:�~�8׋��X�A�����p`
�!ưl�6-�#	L5�q쉓w��$B��'�O@4����Ś<���� ���_��$����	Z���=��KA,�ά�4GXT�����o��kHt��e�ϳJC��*)u����x"�*VV�$z#�	���TS�0R�w�n���,�P��ӥ�DX��2O1+^��� �E	;W~��A/���(ȥŞ�aQZua&�)CҰ�Y��@�|����%Ud���
-�>q����/��<e��iرO@ݡ���{Ȑ�����9!��0hT��J�0܀��I�xZ��;��E�DՉ��y̘���I8"��(X�'��)��
L�c���fm��0�[�F��H�4a�:5/�b�D��NL	>��� �C�nk��|��aq�^�%���שb�:u�Wi��VR�sR�^����1}��O�*+��a���=�D��O���P�HU4M޽����Ce̒Oک�0C�Ei�t�	��PM��]��ħ�a�oV1 �D ��"p����qa	�d�dD�)��J'-ϭ�u��O#�Y�VƑ9oup��-��A*��,f>y�eI�S�X�bq��&+�˓$ @���ܴP�F�*�͜7RU� �88��y���?4�Q1�U$�����*ѝ%�|����?Bu�@��y�Q�
�! ��i
�țb/hH��N���� Ͻ��	 >��c-��~[�]����hT���  �%�2�+G��+G�=��� 
8lҺt�B��"�>�I�n� �W ̈́�������7�5�I� ��0�r�x!��jSLѦ
i�P�+���؇"�.4�U&�6�|���L%���J"]<���-�q%���R��.�m!�B�O���7�Zz�EX�I�2{{
��!/��}u�5�G���D���g'�;����O�Up�I�0~p���w�`�K��N�#o���$�/g��5p���96���O��K�����[���N��*��F��� �ݨ64x��E���X�-��	�̑�`��R���j���'����Тk�V5ѥ�B5Ul�q�
�0n�%�vM5��4c�j9�m)!��q�&j�,=kV]+�m�2/��4��J0���x�,I#fY��WȜn�b���S�.���:%n�(����$�Ă�����bG�UBt��b�(�8/z�h�!���#ˆj��ф'Й؋A h~��ȓW4H�� G=L�2�;�͈����"�Uu����ӻuچ�@,U6�S&f�Ѕ��t�n��WO �bj�$�թ�A�T��$܎+	L�:� ��DptQx%�F���P		����Bķ�N��"�?o�0HBƼq����	�$���s`�^��pvoQ���$�@]J�y����>�:0�a^#�?���X�-Y*=Z��? �l8C�O$g�`��R%Ӡ3F��;!�'�tP�aW/n��9��A�*��G�wx��6��"�aY��Ρr�rX�!W.m��Q B�B��w��P�d��&^*�{��F2m	����'5p���
I�xqK!o���6×��ލ�t�V5#Jq��AJ�n7r�갌�Ȧٺ6����0Ty��ƛ��W+lU��6 8΀I�fC��=�v`�5��@�e�]�8-<�ZBX�)@��hSoԗEZ�zӵi�LCseH�lb�H*Zj�l���q��� �!r1eQ��,�K�> 0���s�d�5�찻v�D/B��$C-c���#۟��JC��O��=�#�!2�tp;�۩5vȵ�d�?�O�)�ǩ߷J���e,�4:��( Se�{��Q�4�PX�@��L2Q�>���'��)��:)^V�� ��.gfM;	�'��9�#��tD�M����) �љR<��yஇ�rݛ�!ѷ������ C
��g�
&a2�3�c�U
a|���8�v�B�'��3�bϓN�\:#���U|� 
�'������M��,q��˦&�& ��'�~���ɂyk8�,�����'���zf��m'�l!M��l��'7܌���>G7c4G^� e���'ޮ|{���?<�1@c�	�|���'O�(�#�C$$d>]j3�ҹw�,�A�'ǌ!�t�J&
�T��Ӫ�/Q����'0d�a욘W�A#��DB�
�'��1@hw��E�V��̴�
�'�z�R��"�4��kK��l
�'����c"�O��8[fG�(¡��'�� �&�)q�^4%=�4��'��� ��kMl��l�& ,��
�'Κ����ʑ,c��D�:|��$�	�'`�-+�e]�h��HC&�Y�T 	�'G&�1��?sw�����E�U�<�	�'��ũM+n�>�"!D����'���v��Ö�ҐA� -h���'�ވȄ�	�d���GkB�K)0�@�'[f�b�ö3�d(�w�œC�����'ӺP�ө�!�ȳ�#B>,�@�'L� �#c+Ь�bvO��<���
�'"�z����=E�D�&��DS�i	�'0h��.�J�r�:ņ�#Kk�s	�'���KA �%dk���W-M��Q��';��H���r�.͓�@րM!na[�'\��[��92P�zgeW�v&���'���iv�qj�QswIٞ&��P�
�'(d ��[��+��P�aO�yr��zE�䋂�	LPa!�?�y`N�ʹ�Гx#�0��yb�	?^�u ���hv�a�"���y2!H�~�1H$ː��J�	A��ybɂ�{��%��挵 ��\Cნ��y�AW?�и�%�֭t��س�%�y��X�J�h11�&N1`s��c�8�y���<l%" 5G�dn�d�b��yb`B�	�0E�Sf�4)���'�H��y��	-��(�c�=K���6����y�=u�Y�㔡I��0�0 Ə�y2�P5=��#�C�q�Fy  *Q��y���VM����턬j�L�W-̹�y2�<Ubx��I:]�20C�j�=�y��A*�s0��WϢ%F���y�GK���SS�W/bX�eI��yb�-Hz)p�.�D�ɘdn_��yR� @s�]�$��)�9"wE��yB�I�H���5���,�]u�=�y��'�M�r���T(V�D
�yr,ĵ,�X8*��d�*L�T+���y�JK�t��@m�e�NAJ�&�&�yb�-uN,u��	�K�RXQ����y"%�/�M	2/�Lc�oI?�y���8O�pT�WN��(:�9�Q��4�yB��g��SŅ�tz�`-O	�yr�#7�`���O�l���!��y2j�*Jڐ<�
�u�^!�����y
� ҜZ�H�<Y�I�
/MP8�w"O���FW�2���ꎉ l�R"O��G�e���3I�1I
��"O�I �ζOn*�@���,V
&Ia�"O�H9C��+Y/V�k"�V�@x
�"Ob�� E/GR��2ȅ4"��@��"O���A�sʆ�k�C+=�� �0O�(�,?�p>A�����pYA 	J���C&ǂ���(�l�fv(�ϓ{�M�j��+��T8��
�\T��DxT����
 he�CL�9&օ�>3�v&�yU�*ڧ �UXR� u:�3���h/6��-���q�1$��AD7���,"�d	#I�����Y�jP�M#fl)�� ǁu����� D��3pcS�7 ���@��q
��I��m�jxRP����<���jl�A��L�y�M�K�>9��<5h��.@�aZ��'��V�^�Q� +§r�@	�'T��+v�ܒP.`Qu.�$Q�L�Y�}�8V{�a�wXE�O�yp@՟�`�[eDW�^�Xբ
�'���h��Ѵq:�<˓,�U�a��
�3PU;��>a��>)���;"G�d��G�_�\]� *�N�<��(^�>�C�aK ]��!Y��;& �u�<x��'�r�@�c�70T0�B1;��<�ߓ3�( ��HM��yR֓l��UB�)U�2>"�
�lߝ�y�Nӷ ����̆Z�����A��O�(, �a��I��Mlz����1D\D��eńi`!�db�vEy��4?1�X����T!�$_5��۵압	6�E��YY!򤐩J�=��)��/q�)����x�!�r�(l��0on�|���T�%�!�Ч��}A	Lu�(;���8�!�ϩ�yP5&E�#�dŪ�.�*M�!��Z���Ώnܨ���#J�!�T�1ܐP�ek�"�$J0�O�r�!�d� e��g@�x)��q��H�8p!�ħI�
x	B��S%n���E!���-�,�Ӈ%=b.Eٶ�<@!���I�:6�Ҥ?�h�rЉÙH(!���Lh��s������c��!�D8l�� 1���C�P�����q�!��"�,�A|���[ы�?F�!�dPsW��6K	��a��A7��d��L�d��eQ@��4G�	�yR-�Y �Ⱥ�@�v\��S��
�y��;}-��� �����K�,�!H<����
��0?qQ��b����6�^�D�<�Q��b��|��X�ؔ'��a��
b�E�c�0p(�=��'�X��eG�?F�ai3.�5{�,��L>a�
�x�"��$�%�'�Y��3-D���E��N����ȓrhi�c�O�Ɗ��䄻SE�q{��'?��v���G�L�kB�J�z7�m
3��+g�pY{�;4�PIs�W:�u��)J�M� �Qd�66`�(e�Xi��d6NS�dzM<���2�BXP$
f5��qx�PxTJ�j))�U��b�S������GBz�bAD(���*��(���Pq��($)�,&X��� V)�'$R���S.�$?��'�`��2���Z���Ev��eT�0!��d��0ȢYV�"�3���#�ub�C�'p �D�E1(xIyr��g��L�`N��2dPb��(���eȡ	5he�7qd�q(g��KF�E��cЃR`y���lt�8��!ޑT@���]4U��X�O�����O�ա�-N�p4�+�"�l���O����MȈIW�M!��ұq�'�"��V��^�剕}��& Ʋ'���Jg�ֲ`��]ɷ��k
t;�JX)pLx#��>}RU�W��z6��?"$Ω^	8� BXA0H�%�=�I�! ��^� 0 ,���P���C��݉4F�/{2��c��?*�\�҈��Naz�OP|�b%Y������.'�h&@�=/�A*X	M��'�YC�j�H�TP�"��c����~Ҁ%D\J	!V(ҹ���F��O��a�a�&��� 
��&U<+z��3 ��C�Z(�)�+mJ��҇X:N���	�G��	�?��(/M!���V?6��X!�]�KR��A��G2==����%��"�^5�4y��M3x� D��!�!}!樺Ń�c���I 񤇑#��9v/�����béj�P�����ND�@d�!<OT�۷��HN�\:A�8 .d����Rn\�0��7��0�VhI�)8�O�8�v(���O&��/R�0D��%ثrQ�d(f�|"�X�v[�Lh��2�[A�,R1��)k!�I-k^�ҷ��q�v�*�"Oh|c�@Ɲc�|� �U�w�hh�k6E`�)� 	6�Vjg����N�?u�0� ��e_J-�*@L��ȓ(�*���!� lmt���aX b5��B)�<: ��f�)|�vc,O:uӠ)�7=��I�JX�d.� ���'��6c�˟���&T� I��'!�mRՆ� �~�QO�I�bђ2��H)&�T1�d��	������
qܧt�n���Q<@,�=� �Q�����ȓ��B�D�J�)���_�P%��'x"M�E���2d�ҧh�z�Ν$pE��zE�4=~H�"O6�!aC\5;8|*C)�9C�>��8FC�J(O���''?�")�3h�f.<��W�'��I�7���<�VLZ�IZ$��l��1�d�AoCA<�%vw���5j[�B8j�HS MX�'S(\0�'8\��m�|���U,�%:,hw)�V�<is�ڍ'T����L���)�I?i�F%h�P�-0}���݂w�h�+'���|wVx1�Ψ!�d��*��n�~~FX�%D� ��K��RLJ�kE���$ͤS`8����ʰvy2���d��=��~r%ϻ7�@���.*k<e����H���@��N<y�F����FƢ��L3�p���{uFtzt�|�	zwB|�;(v��)����Ӻ"I<�$�F䈾-���k)�k<�S���(�F-E�nD�GlD�b�t21��h�P�qQ��4{�qOQ>=�nv��z����=i�9��-�EVB�ْًY����ϟ�,�F@X8�옲�KT��8�"O�pb�����2#O^
�s�T�$8V�K�9(Qi�N�R>� W!
�Y܁iB�U�J�BB$#D�$ ��l�d�����$gŀsD\��H8 �����g�2	�Hɖ��1�,�����>x����ɀ0�x�ר5I|�3���%�^�;qn}�Ta�aW|�'�$�Kr�U��T�	(�I����"B)��J�?����x�@@CL�Di@��h��$��
XT��l 6)���K��`rJߝ+~b�p2�
.t��&@3�'b/�eI��<HS�)��l3�r 	��L��T%i���y�.�S�Og��h�'��Y�1k�C[��H�5?�!h^$���(�U��a���M�g~"�%��D,L�<��up�ֺ~B��p�� K����3�in��W��&�ўHK#�� -"�D`�T���"A�6�%����&�D�}��.U�.�k�$o��X��H��g�� ;D��_.H3��z�~�R���0ÈO�� a�o*D�S&OP��趁��
��L�An�J��H@�/�$��I��x �m�x��lL���L|JD��,<�L,��`�r�Y�Ɉ.��PٲњB��i1����0DI��
�5������0��!M�]剌'\���O85�So$?m��K5J�
>D �`R�=�>hʃ��>�q�H������S�*�b&��^z���8O_)�)�.`�9���'|O6U �m]�hȬP(gA�hq(L�"NC���F,�w.8�>��!]����AG��y�d�>"F&���NJ�y(��D�=��<����;z <̒P_�=I"�w��%"�c�z�x�kJ���p�@���:-'yr��	R�~�T)P'H�c�H����Z=A_�'�L���$Z?DU4�ۗ	5�'5m"�1�h��I�l
ÅI4κ1y���a�4�'i�eK���!�GN�}�F! ��Ey�pL]}�(�'-TB?�S�Xaﱟ�'�\� �d C�`����H�=��%c�1LR T-6|Ok�L��YI$�X�Z����0\.|�A�XG�J%��%�O��!K�6 ��0 B�V^er��'�L��*BJai�齟���� �\���F?<�����#D�d{��.���ge��4�(�2�>}�o
de�a��l<nm�?mc���*��q�a��7+[0��ש?D�� W�Y�Yqt����H#�X1�F�t/�a�-O0�[e������|��X�W9a��Q��"mi���?Q��͙98�(��ᓟ%4xQ�� ɓG~~�B��A�yB��&�)�G�NX�P�u�Z{�٣v�ʩL����ʴYPD�ŧ�<���T����?o����t�ϫ��� j�J�H��Q�����qZ0��"O�=�r�ÄT�<,�BVg�Y��iW@P�0�T`�N̊���Xʤs.O��Q�.�^?Y8�cA�2>�0@Ç��,0ea{�gфo��<���ͼ�MSf��u���F_��I9 i�g��XO���2�������Ia���BA��/J2E�Wa����>�UB�F42�9���E�O��U���"˜m��#��<KXL�5�J�0��'�ȭR�ŒV	�S������(@�J�1%1?���>����B�V9�ď�r�&�"/}�<�$ϡtC�,��ƚ^Q�%��E���bGd�[j�M��w<�C�ׁ)��Aa�OZ�_�����~֌�5}�RU�Z�B������w��E�F-:D��7��<%��=B���[1N-)uN5D�@�$C!�}����I����?D�tPW�#90��ۤcגŁ�(=D� )�N˳â��n�<*D�ũ9D�0�`\4e��% ̭rg�ڣK8D��bR��+v���0u(��aH�d 2D��跮4K��q{�˳$��,2h=D���sh� �Q�gӶd�2M���,D���t�	�@�$uٷ���"�x�IRM$D��)��ѕ6LP�{rbY�8�HU��g$D�dSQ�Z'O�t�pu��	� AI6�%D����(�qׂ	�_���c$D���F�]O2i�1(�+��,hwM6D����U
^���TMԡ�Bd���5D�L"�]:p����6J���?D�xK�b��}��qwoB�XHl[�;D��9�T8P�Z�t��*��4vB�	H�u3�I=W�%xq��:~�4B䉗H�ֽrpm	3+fi+g�ԜG6RC�	�.��@m�,}Z��v�ӂk�
C�ɣn���K�-��]�:X�-���B䉷�8ŰG��~��CE��j�B�;U�p��v	!�ՁT�T�`B��%�p$)Ӣ��.{ڀ�$� *Q�C�I�ZU�<(��b���Ӱ�̙w��C䉢O��YH#��c�)xt�K��C�	�{�F]���Q�#N��[c�[u�rC�Ii|u���2L��8�$L:dn>B�I�A��h�	�9)��c�,Px��C���n�	p� 3�X�2�3|��C�	 �\mP���|J\h��˒�7�B��_�`q���:m��}�3�E�-��B�IM�\��#��V2�M	�oC�r6NB�	����[�.��"㬽v	.C����,6����q+V5'e-&G��$"OB�S` ��4ގ ie� L�	 5"O�lx�I�!l�Z���:;�ձG"O&��]$#�R]���Q$���ӕ"OԼie����҉�U�ʭ� �Q9���AY�(�V� ��'��!B���,l\���[�d�6Ł
�'�xU�0,�0eR����Q��	�'H8%���9,�p��#ڊ:��,��'0��q�G�{֕XSOM�.q�Y��'^:�`��8n��ū����'����3��0�BjF)���z�'sޔ���T�;t)k�81�,�r�'HXġ�A
�B���cI  &E�Ի�'��ճ�Ќf�0 �X�r���Y�'a2�J � �]%���Ͽ`_�Y�'���J�OɊ�.�XV�ёU�4�h�'ʜ<KRNT�T��� ��q��
�'�����ߟD�,2����,Y��'i��1$A�<c2L�
���
���
��� =[F��(b!�p���ڎv.F���"OBtҡ�ްg5�8���E���q�'��	sF�>9���M3�ӎM�l����5B3ּ��B�z��iS_<��'�����O*(MIW�T�Z<T�z���=k�(Ტ2}�{�"<Yҕ?�X�����o�kv'��N�����~(,��v`8fv ���ʔ�]OB��S
j�W��b��U���� 8��H���n�V�(�pT�F�a~����0|2b�_�mzٓ+S�7� e
p�@�#W�1�'n&E�����On�OO�I8�D���`�9S�N?c^�:H�Ġc�Vĸ�e�O,�P�7�D~�jר	�*`�4��O
$�3`;FLQ%� Fx�/@ЂB԰W0^a3ÃK��y�Ɛ9�:9R�::b�`��y"�4���	��"-	N9{����y��=������%��DX��V��yB��8���S�ȍ"�:Y���_��y҉^}�,�ě�FCS��y҈)�⍻������W�y�N��+MӃZ�����Ɉ�y"��@���b?H�rTzp��y"�#K�������8��`�t�֨�y��� ��,qd.�")28���ĸ�y�=:�$]����4�{�뎌�y�S�Ɛ�e>��=Q���y҈��/X����Y��,�Hm��y(�8//J�Ѧ� �@t�#�yB��Pe�p1�[�s3������y2"��p`���
K�A��)i��݅�y%O�ZK�tl�#lDcc���yR���	�R�Kp�T(�fX�yrJ�2Uީ��EE�ZMD�yB$<W����W�QLx�C�ء�yr�Uu*��FH8�XS���y¯��H֬�SOH+=��$8�O^��y�`����GN�9O~����Q��yb!^8��@˃�3/|�eR�M)�y�D��ѶN�(��dQX=�yb�?d���ŵf(@PeQ��y�h�p����P������y"-��p������7G@�՚����y�]�=���s��(CkT{��X��y2�7dj�i�,ǚ	��Z�j�4�y�ŗl�5i��ƕO{��귈���y��9��3���}���2h��ybnľR늴�&Q8?� qQC)�y��X�|��]��m	�0w d��S��yB�ʱp�em�X� �*�&�yR BU����wBM���w���yr��r��h�q�3}u(d�QK�4�yr�Ĳ� hD/��	��� �c��y.��eR��˝��ɹ�IZ��y�I��[HbL��
�*���q�ݫ�y�� ���"(�,���)'`ƴ�y�� iP�!��B�&�̬����+�y��B3Bs����FL!l����)�y���6�`�U��-���a*Ϋ�y��ɧiV将;*�>a� �E<�y�M�?�AX�̚�
�<9�-��y�����f芻M����Eԏ�y"m��?:�M*4*�F�`�7M9�y�ɓ��z$���H�>����W)V��y�n��llHQ��H�7�H�`���y(�,M�`§df	
���6�y��H-u�}U�ϳj�pk��B��y�'W.~����N�h��p�T�+�y���*\д�"�Wp"���;�y
� ʸa.ճ��Y�)ܫ#����"O�H�ĸ`E�`&��(*q8%�"O�\r��� �b���V�"O�3Gg�?p[ �pth�A'�e[�"O�t�P�	`un�zHȊ �Q�t"O��" {���2���~�V��"O@�6�\�FɒQ��GW8q�M�c"O�1D�W�-4z�j�K�B�ٲQ�!�Ę71wd\�3��F��#���{�!�"f:�P�ߩ�X�!�V�b�!�D@!116�a⑘(�\�VbP�o�!�dT>-�Ե�d�](b&�Q�#՛m�!�䟣2%u��-ِ=��k�@��T]!��l�,A�kӖe�1�Y�V!�D��K�J�`��� A�^Z�-��X#!����x���Z��\ȡM�!�Dߍ"V��0O�a��г����Y�!���2��h�2��O�x��Y�x�!�ČvX���0f�PR��H_!�D��!xr�sū1���Nʍ[A!�dߢm�D$��AH�m�t�`���:!�/'�4�΢ZzQ� "�<!�$��T��(�Z��81�6"^�^ !�G=T0(ѮS.h��)�G!X8N!�D�-;:Q�H�u���	��!�Dʐv4j9Ӓb�8|d�6�8 !� 3k6m�c/�H�1!�^�dN!��$a�bE�	�]���J�gN;.M!�d]�u��E�%U�j	�A۟rZ!��>iP�
�@ث8�abGG!���Np��f�ƹ� 
�wW!�D,7�&e�m�?/y�u�tE��!�d��H���;t�N�(N�䂦D��,�!򤊴��H��ץB���(!D��/!��Q'mJ���J��8��}��җp-!�K0bb�s@�z�VI�+K|!�䂢'����Dvݖ�#��W$
a!�d̿K��ɀ�%�/*��0؀e�4 !�d�6*��a{���8�r<I��̫<�!��f<�+�{�vCtiK�4�!�d�=%��;a�D�zMx�����!�DU�;½���(�J��î@�z�!�̃6�$���B�	�Ų�E��!��#PN�Ԁ��Tk΁S��Hu!��#X�J��ĕg^�V<x�!�ф5�Q��]A%�h��i°^!!�G�@/��뒁�6p2�)�1��R
!�ڭL��t�"��<G��s%C�L*!���TX���`�$2^��(/#!�;B��P��L"t��6���Q!�Ć:N
J1,�cd�,!3�$(�!�?�
p��^xTH���!��Y3*̔��j�@?�{���T�!� -�I�4�%<2���މ:�!��9>ѐKe)@�d�VA*���o!�D�X�|H�pA�?k�b���.�
!��]h�)�A�o������5!�B8i���1�ʝ'"[�ŉ�i�%!�$�Qz$�b�
��E���8"!�d~���0�%U>������D\��'!��JR��{�l͠V�X�:���r�'2���Z��t#6LϷ6A�Ș�'"��ځc�=���o�"����'\�}�����x>�c?�֘H	��� �H�kڀH���S��.5L\��"O�i �L+}���	�i�g���b"O
d���Q%t���qH����I�$"O
]S�-C)Q^�ِ�Pl2�y�"Or�lވ(z��ּs:��� "O�)7F�1(�p��C�RO�2s"O�I���	�F=�8r�K�$`�y� "O�E�2�׆�+�j�7}#��z�"O2����6{��:c�	
�� �"O����X�./�qq�Ƌ6�t�b�"O�0��V:?�&�Y�*.(����"OJ�A n^=Ic��l��}��"O�8�3f"Sr��x��$:�켱�"O�0�D������FR����ge/D����O�d�Hnت>0�q/D��E�����*V�T�{�H�$�.D��a�CO�3�̭�t����eB�+D����k�D�H��kQ2J�a �(D���1+����rf���X�AI!�'D�4����_Az��!Z�ԙ��+!D�<�$`�)t�\-`B熇Ϛ�9�#D��ÀA@�;�5�_�un!�q�5D����@�-yh�*4�ɥ:�09k�N0D��z@��\�va�a��7i��
@0D�l�0��+2}N}��D@4U*>�ȵ�#D�<pqC3u����_j�RyPC%D��*�ꏐU�Rew.�^ak�o5D�p���[�${l�;�&A�]�(��� D��(�I��J@V�)��ԄJ�D$3!A>D�(I�"չ}�~}���ϔR�@ i�<D��YwA�9b��u�RɊ��~��-:D�Pc!�ؓl�=�kP^���7D�H�0M�/I:����ܻut<�#�7D�H���Ϗ0�|:Q+��%��\��e4D���2�Q�kحHab�r���"3�3D�T��/S�����&12d�94�#D���v*̑�`��5�� %�Eh�&D� "é�; |�Mk�C%?N}[ņ0D�������c@UZ��m��̭��y��,\F	��_�GO�����^��yB�]�[�Va ENU�v����B��%�y�+*�<�cЉe��� "��yz7�l���-_@K!��3�<C�	W�H0�BZ���o�R?C��-Lo|����@��)��N��C䉔]9��"C��v���0xέ�"O�؃R��1x�P���c�$�`)�"O,��R�Ȑ)�X�Ã��:�2h�"O�qCg\�.��x�[�\ϐ%hF"OT�Ä_�Z�����n;�L��"O���@��:3�:�Éײ8����3"Oh]�	E!|t�Rp�&�֨{6"O�����q@�PR��O�1��ea�"O�Z����u#�P�G+*m<<9��"OjXғ@�_zj�J�(�7'��b�"O�Qq�ٜ-u@iQS���W��x�"O&�&�G�Qߌ�e�E'S�l=r�"O>����>b!Z�j��D,�8h�""O
�� ��<]A6H�����"O��!r��G�r)��&f�$��"O$���I��GV�r3(�$4je"O�[�閆z����d&O�3�4P�V"O�b�*�}@���R����"O���7+˃{��8���=]��4�1"O� ܀9��H�B����;Q��C"Of4�7	R�q,!�ʛA5���"Oz�*6�˿��̢�\LRhq�G"O�l����g���8d�H�z�(H��"O�)��!��j�}��CLkf�"O�!�C���:�v�Cq�&$WBa3"O�j"A�g�}�GQ��^��d"O$4:��������7��}4"Oةi�.��>�`���I���"O�;0��	�Q�I��y�c"O���p#C�p�~��HE�mP�1�"O�t!x���F�'=6�]*"O^�	"f�-"ek�T҄� "O�z$oݰ4.�#Љ�b��(�"O��g�*9>�]� ���C<h��"O*�8�   ��     r  �  �  )*  j5  �@  SL  �U  '^  �g  �o  7v  �|  ł  �  J�  ʕ  +�  ��  ٨  2�  ~�  ��  ��  B�  ��  ��  ��  *�  m�  Q�  ��  5�  9 n ] � �" �(  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��l���_�a�)�Y�!��-�	W<)���&M���#� Z�kY��3���p�<ɒ�`H���p�ݎNLJ��m�l�<)C+��5���k��n�d<V�o�<�Aa]�K|-���J�ș:C�t�<��E<�	��I�����n�<��K�
Z6ͣR��3�&�Y��T�<	�F��l<�p뒔g�zhz��˓Pn!��AbM�#& W"C&)ӧ�ܡn�!��;
L���WQ%�=k*�,�!�DǨ0�4���jR�[ �&�Wa{2�dF)�bUY�C�,_+�	i�E�xH!�$,&Ttx"���C��yuk�'[�Ȣ=E��'����BAA�9��m�F��o�@��'ζ��1Ǘ����E��^��N����2 UkW�^	&J��*pjѳw@��=����y�ÆF`R�ʵ��%Pq@DJͷ���0�Oh8�ugL	Vm�E@�M*Kx�[�'#��P����'?����*m@�X`!�;D�$�j�Sľ��"�R47�����8}�[��'��?�+W^^-V�уI��zG*2"1D�� �`�ckۧ%�>����B��$�R��iQ�'��)��|"�	(KHA�gMկ��R�\��Px��iDH�ş�`����#��Db�'.�QS�$+4D��I�<;���D�h�`�n�;�����`��U�!�֛�J]��eE7E�l���	)4�!�d�v�Z蹠k�Ck�)�����O!�䈫T0��c�j�? E�4��	^�c�!�$*n��\����5�uQBbJ03!��P┨��$vd� ��o�!���d $���A��IpoC�y!�DD+���A���3"� u�3l�".�!�DO�*��؀B�:�|�q!V"l�!��,<xСY����oI4�!��F'��!��F�f��#�n95�!��ztX)���>7v��`K�U!��w�N!�b(U3/����Ȕ�[�!��*Gb��Uo]�L"&��L��!�D�7+�2<�6*_N���I�!�6�(9���Q�lL�3goݥ?�!��N�dx��XU0�y��9Q�!�� ��8�O�7\�xM[�b!��<�"�)�XF�C�!�D��/�z��	Y6=���P�F01�!�dI�U�}�C>Y�(gۚ0�!�$ťH~�%T�qZ҅G��!�D(=Ŗ��̏Wg|I���Ǒ?
!�DǏq�Z\q��&nH��K�.�!!�DR,Z~���4g�R�XSn!��;%��0&���@��8�4�'4!�d����I�jE:�\�f�D�T!�;`����s�W=EF8�!��`j!��#���U�M-�T��a�@�!���nJ��`u|�BN�"�!�Ĉ�^�
u�E҆9b�-�b!���D�x�T�N��e�D��/=p!���g�]Ʉo
4_�Α#���G�!�d��Q7 �����)L9Q�!��,
�,T�����mڔ*%��3�!�K9
�X�V�e�T��,�	�!�$�\���S�/Q���Y{!�d(��a#�]K2���K�<�!�d�6]��z��8���s�]<�!�D�[Mj�ifFR9l�<���@�Wu!�$�/$�p��v��=nT���b�M� E��^��H���8e��2S	
4+�n�3U�$�O&�'�`��T���y?�3���e^Tb�'C���6�ďy����6��?bȦ@p�'Ҥ\+�cZ6���� B�6X^`��'#>��0��H�`���~�TR�'NB �� �-������v��i�'Z�Y��C:e�sQKª����'vL�b�MňE
���H�������IR��EJT�V� d���.H��B�	#"��+�`սt�^�"7�У=y�'$�P�ՠT?9�P��@�Zd�N���O&������H�^���J�>���ȓv�lt�s�J37�.`� �Յ~ �EyB�|�d�?� �v��<nF�(6��b}B�'����j��9y�	��߲|�'�<H��g%Qx�dڂJX�]�x�'�bQ�l�� d���ۆ����D(��Y�ӎ��E�Bi��!4Ph h�"O�#�-[�h��U���C��Q�"O� n�0 ��c�6 9�n���T���"O�"�&�!bB�%
Z?��*��Gy}�'I^hP��V)
+�Dc$�Z$0�~|3	��hOf|��.Z#_Dv$!w�δ#�����"O`�q��!�(Պ��U�n���O��D�@�Y:�L�G@©�F���|!�$��#򬺀jHf&ν E���!�ҠY���K\�-�a���r���"O��ٖ��cVf@S������"OvA�&!_ ������"�b��Iz���I�#y����	;f����'W&�!��K�l(S�M�=��"�$%�0�Fy2���0��(�p�w�Μ�$=$�\#�#5 yY���!��1V���j١�ҡrP���7O*
�y��>�Q��'y<=�|��c�=� �J� �$�z��Z�<�2DM)q(l�����TUx 1�c�U�<�W�FfTY���%��$�rDS�<��M״Q�&8  )�91��Ny2�'��R�K�_���b��IG�`	�'#ك�+1EJ=a�(,����'�쉫3iy&����-�����'L-�W'�&��$�ێ�l���'o|�1t/C3Y������C+{�58
�'
�8u�$Q�l��R��n���x�'r�$�Dl��a��8@3M�+l�b�a�'�p�ì��.: r��c ��r�'���$��>�Ωp�EH�ո�'Qvj�e�5iz��;�U �:`�'�b���d۠)�9�CLƔ�����'�Bሰ�W4[����E2s,�Q�'ɂQ����==�0KC�q����'~ ���K>\@�5C��:��-��'d��Á<����v��.6�r���'�h���e��?���V�ֹ^�>�	�'Ѽd9��
9�d1FA܇ I�\S�'�y���(PY��;�(ղe'J���'D�R�Y�y��i�PY�88P�'v:�HFD��bJ%�B��4Nm�d	�'�܈Q�"{�y���z�& ��'*��{�d��J�YCT=jr,��'�Ze8��B&/=����c)�LZ�'±3E�0*���C�[�`-�y�'ِlx��N�<|�tJ4.^��@�'���1�!i{j��<A�H��y∟�DUy��L�3���9��0�y�\#G�eр���I�Aq"�I��yr�D>�:�HV�ن>%h�Ӕ+,�y"玪7M��u�L>&6�P�"�2�y����o_�mP��Ņ,�.�b��ǎ�yR�<�6*T�Uy�%K/�y����
����6Lt� W'݈�y�M@�[�<9�Fn�( �*6/$�y����y�r��0j���H��\<�yBʋn�	�g�5>P�iU�I'�y2j�J��ѣh֔+Wd�2r ��y�lǨXc�4s���	��Y�fb��y���2.<94 ��b��%�1���y��Z�t?�C�@�.?�|���y2�C�4 �&D��aE��K��P��y� B�:(j&ř$�ܵ�Шׁ�y�HT�i8>�	!�)� Ԉ���y�)W��� ���ݢ6������y�YB�X��]�;P���I��y
� ����b�z��`��M7���!"O�)��B4$wP,�E
g4��C�"O�H؄��#@���P�\~(�ȣV"O��0��M�2�˱MQ�Dh��d"Ot�ѐK�(#5�d ���/3��Ȱ�'���'���'�b�' ��'X��'�^H�nrR��Cb0I�\i��'�r�'m��'��'D�'��'�n�	d�V�,�� #��V�ڢ�U�'T��'���'�r�'���'���''x}��+̑B����B��&*�B�cf�'���'�2�'�B�'���'�R�'�DeB��_)Y�e�F^�7�.%[��'�2�'���'���'r�'���'����T/ÍZ��,�X�PA�w�'���'���'���'���'��'�R�릯�7WH��2D�V� E��'�2�'��'72�'(��'���'�Ʃq �H�N�*�S���BĔ����'"�'#�'L��'���'��'�*���2TZ�a��ÖR%�康�'gr�'��'|"�'���'/�'i~Es��20��Xqg�@�W!8+S�'��'�B�'b��'��'+��'q��5,�	�}(&�� �y�'���'�R�'g��'�B�'
��'� 8`�ZU�v$8q*�F�R����')��'���'��'��'�2�''"�Ң[�$%hRo �}�ZS�'�R�'���'���'v�D`Ӽ�$�O��R(R O�N�S��%d�F̲�DNy"�'��)�3?��i�N�j���.5w�d)4$̫Z�����4��d�ܦm�?��<���C1Ҩ1V�Y�j9��Q�ś�;���?�a���M��O����N?ٹqE�9ZT�I{���(yT|���%��x�'��>�x�M�0cWص2�h�ܒ�o��M�d�F{̓��O/�7=��թM ��^����Գ2f���k�O��Dw�4ק�O!4XzӲi�B�T�t���L%��"��C�R���f��Y��2K8�=�'�?�6b���!)J5f�U����<�)O��O�nZ�(۪c�t���K�e�٠d�4���3.G�{i�I۟���<Y�OF-�d�*k
|1�'	� �����$���Y~y�5o.�*Y"o��H�"jK?a���;E�$dt�)��TyR_���)��<�R
�0M��!�6� @m����f��<��i�&%�O��nw��|�1m˂ho�|H��D1���#T�<����?���↩��4��do>� �'-H�©E�:\)	E	�)C�4�d�<�'�?���?����?��	�0~8~T`'��<�,�σ���DޟPp�D�O���Oܓ��QB02qRL�� 4�P!�$6�(��'���'�ɧ�O�}��;C��!���X(|>X8EM>h�+�Ox�� J@��?qW�1��<yՍ���Vu� 	 3+&M��	�$�?y��?Y��?ͧ��AĦA`�A럸ZGcI��u���1(&��6��H�ٴ��'
^��?����?)D��C،����E�%ϹM2؅�/V�M�'�6q`��LI�O�G%$I�R9�2KY,Vty3��V��y�'���'���'�����'!b,B�#�>\�tD ������'���'p6m��WV���'2�ɜ㖤1�
2x�(q`F�� �>b��������&x�r�o��<��9-�-���	�v�a���:R&��$gу)���D������O����O��	�Xbj��T�ǡ[���`o��3T|���OHʓf<�fJ��1"�'�bX>�X%�E:c�����ܜu�m��#?i�R����՟�'��Qd��*!H
�T>�)1���:� �	E©� �Y�_:��4�`�:�{��Op q%��i�&P�M]S��[B��O����O����O�)�OʭS��<�#�i>�=$옂HZ�ͫc]�4�0�s���"A��ɽ�M�O>�����Ο�P�LP�\�����]���0�- ٟ��ɴT��mZ�<��43P@}sa#��?	�'V��Y`���.�Z�`��O-*�H���<�*O:���O"���O��$�O6�'`3��
ϐ!V�fp�c� �6��3��iq�:�Z���	s��V%��w����r#Ϫg�H`y�I��xQ\Pv�'��|��ԣ
Ow��6O�9�v듦 mD�Cwf��l�hL��0O:i���F��?���/�Ħ<���?Y��@F�ѻ��T�C%@5;����?����?����$���u�c���t�I���`�JTx�J��Ҩ#ŬD%�J��$�������ON�O�E��C^<�D�A,�0��"��4B7�ƨX�@��%>�-X�b%��I���jL\����
0�`�Ο��	ԟ�������r���?�dÛE�Y�&蟅5m�ɢ�,�,�?I�iJ:���'��f�O,�4��T��k�0d��-r?�C�:O��$�O�8W�6m~���ɉ[�~ ���O9��I��>��ͬ���§��oF&�$���'#�'���''��'�b�sUܒ5�m�F鑙j�̩�[����4�lPS���?������<�5�ϹB����n��o
Xt���	����	a�)�Sp����_�3����ꖸHL��J�N[�y5��p�8����O~xaM>�-O1&離1@0	4*˺*2��#L�O����O����O��<�i�U��'��Svj�PJ@�
w !��'4P7M*�	���$�O����O��8`NRA���kQß�5�0����$ ɔ7m'?����g8�|"�{�?  �P�悟
�nY�,�x���t8O,���OZ�$�O���OV�?���W 	!�"]$,��Xy��^yB�'��6��[�	�O �n�u�I4C��iI@��>N�5�#��.�,d'�4�����S#F�UlP~�P"}��0��*@�<$�� .�P�y��ҟ���|�[��ß4����X1A%	�v��Y��ߒ!�����ٟ4��]yb�p��0���O����O��'b�\��g�J��,j��A ��q�'��?!���S�4"S-|�bw+����t��f"2�3��ճl��ƈ�<�'$����� �'48P[0���a!�@@��+��'Vr�'�R���O���MK��W:"T`9vHӠ6�R1p�Y�0?��;*O��o�A�3��I��8���v�ֵ3�R�*�̑�0��@���,�oZQ~���u�NM�}�������xAO�%�K�� �<	)O�D�O��D�Od�$�O(�'w����0���
�M
x#Qi���M��e���?Q��?yO~�f>��w#��b%I��~�~t8T'�B�z�b6�'2Ҝ|���Y�L���6O���N-vl���

�b�8�;O��A�"�6�?�
&���<�'�?�" 6uȔ19�;4��J��,�?���?�����$���)�u�]֟��I矠@` ��l�p��
@���(�ccTK�in�������h��-a��҆c��=����-��Z���~{��
��q����O~����O����g�H�c�h�
��e#�KŬmҦM��?���?���h����	���M���f�J�KKl֎�DU�I؆,Y�`�	��MC��w`��#E��h0ɐ��1K�t1��'�P� Ib�Ʀm�'>ų�
W�?���Э)qzIq�}�h� �.�qF�'���џ$��ܟ���������b�L5��M���!��ΉL���'!<6��LwD�D�O��-�i�O��Y����w��-���̫[d��2�]}��''��|�����93)����I�U'�`��E�&��L���i�L˓(r4i梟�'�0�'u��"dP6z����dԠ#i��B��'Jr�'������W���ܴXo�%���jZ�����k��X"f�ˊ=��̓;���~}B�'�'�����ǅ}'R�Y4�:^Ɛ�Sk��J"����pCKίm�������]S3�`p�,b��V�[��d��4O*���OH�$�O����O��?Qrd'�F�́b�Y ������ߟx@�4hG�e�,O�nE�I�s���T�á3�x��&�T�*��]&�,�I��S�h&h�n�g~Zw����C�X�z���Ks�C)���i<SR�o��Ky��'I2�'2�ŊS��u�����;���#�A��'��	%�Mc!녩�?����?�.��+w�
�(�h�;���:mo^Ñ����O^��0�)�h ����A�U;	"p����
�jp	ԯ�1DT9�*O��?�?y�d"����<�;��)?�	�I�>�
�$�O����O���i�<Ľi��iQ`�3�D�0���M6��2�M�� �'W�7�'��3����O�`���H:݄ UVp�,Y�pA�O����/4
7m%?)�NO7+	J��wy�F� XS@H�1�� db�]�$��y"U����ٟ��	ߟ��IӟH�OW�t��)WlZ�ˏ5&x�ȢAi�\|#���O~���O�����ܦ�ݷ]=��Ph�.D��Q!FCƷYj����ҟ�&�b>qʅ L���͓}�"MA�
FN�`[��R"Z���U���I���O>�(J>A,O�I�O�`�oä�4���V)Y*�O��d�O���<a��i{��x6�'���'����F���H��,y�ڐ�e�$�_}��'���|��ң	��3ǫ! }��r'������Wj@����H/1�����~��	��QQ��e:D�`'DO��d�O���O��$.�'�?I��(NW
)��D��=���?�ֶi����@P�D��4���y���_�dzF#׉{n��#̝�y��'T��'d(��p�i�I��|� #�Ox|R�eS��=���Ȓgt᪁a��Sy�O���'qR�'��dM�d�n4@eL̾�Rl3�D|x�	 �Mc%�ȡ�?���?a��Ԉ߂;��T��B��#��#ckK$C�듵?���S�';��}X�+�%2`�B�#��6X�P�%�>��'l���kD�� ��'���ny�h�J�S��dj1���E�<���'�"�'�O��	��M�v*��?iB�j@����'��L�ҙ0�i�<2�i��O��'�b�'E�L���)#LB>@�,5!��[�'�P�҂�i���n5�
��O�q��nY*x��px1 �5��Z�ሱ6�D,�O&����VX	i��H��<!��@&�v���)Ŧ&��P�m�{�HUd'�_��;P�O�����i>����ۦ)�uw��r��b�8g#x�6�Y�n�^�2pf����s��|"V���?�G��)r���1/+0�S��R�'2^6-X�tF�ʓ�?�+��]#6&F>V��lZ�G�����[���C�O�D�Of�O�S^�P��Ǌ<_ږ=H�E�2�UV$��Qy�O$P��64�'C��s�P�A���s�
	��z��'B�'I����Oh�I�M�p��b�"���!Pz���	x$:.O��oZZ�|���ܟ��G`�%}g֑#�A[�Yi�س���H�I�O��lj~Iߍu��x��X�� D���N�T,�2��@�>�X�I�1O�ʓ�?Q���?����?1����̬#�b@ �&�'m%R�8Q��33@$nZ�@���	˟8�	X�S˟t�����-�::� 3�W:R�ZY�d"���?����Sܧw�2�nZ�<!$n�H~u��+�#����`��<�$R�/���IF�Vyʟ�b�@�@}�V�R Tq8|�p�'v�7��w�&��?-8����`�Hْ�j��~��4�R�>���?yJ>��aR�<z��I򌈢%V� ���Z~��E��-2ÉUd7�O��1��d~�Ȏj�zhi�==���C�Z���'D�'���쟸�5Ꮥox�tqSN��+���3M���L(ߴJ���?1�;���4�V#��Ͳ���TFL1�e<O��$�OZ�Đ&x�7�2?aU@��T�r�i[�4�(S�Ӧ_>��QT@Ԉ{p qBK>Y,O��OH���O����O��ȧ��6��90hIH#�� �i�<�D�i�� A�'��'���yrG̃�ъ���<;����pO�L����?�����S�'[����L��B�'l[w�X�cG	�[��]�'���@��ӟȻd�|RV���AP<#�&	ps%N�0�YҁĈџ��П������py�e�>t�pd�O���1���b�7��E&�@[6O`m�l��MK�	����	��.׹BK&���J'L{N<��dJ����nl~�ȗ�)�B��SP�'Կ[F/Q�9�np�C+*uz5��O�<���?���?Q��?���$Dǿ?��]9�mX��T�h���*@B�'���O��"T���4��s�f, C_:�AZV���U@D<�d�O:�4��l�p`m�f�r��,Hp̍ U@!��P!m�D�p�N�%���D��䓎�4�����OR�$�ei��iv���l\7}.���H�O����<)2�iF 9C��'���'�ӛX�����
�j�فJ2/����	ʟ<�?�O�����N�vR�Q�F��5���X-F�`)�"]?��i>))��'T��'��ABA�n����+z*���n]՟p��㟤��şb>i�'%�7�`�R5��A+w�b�C� p�:9$��O��T����?�_�t�ɠ��uH�L�F�"%�����C�X��ǟp�`Ӧ�'0RE�t�,O�(y�L��JXd�*���*d�:5��1O�˓�?A���?���?����U91���/�>h�v���	�h�}o�1d�m���P��j�s� ����cq��L� qެ&
�U�9�?���Ş:Q�ěߴ�yR��>rK�/WZ�c5��4�yb�C!�����9V��'��i>��	e�Ty�сY52KB v@�T1DI��۟�	͟��'(6톾'�`��O���=*��9zP.�c|��zf(�!� ⟄��O��$!�	�j�p�hÌU���ق�Q7������Q`"
 M$
�!L~*@��O �i�w�x4Kp�hGDC�w��!���?����?���h�>�D��=��Px�i����+S�Ǵ94~��˦�y��������M[��w�Y�EL�r�8�Z�=i`�Q�'��'I�N%n��F���ݏ=}d���[�V	A�I�"�t=:U�#;�r�0ӛ|Q���I����ɟ���⟬Z�'W�
:�LI�,�$:)��G`yRab�����O�$�O����d�+J��"O�U"x8��A��\�'8��' ɧ�Oh�����6\���rm��΁[A��Yyx�q�O2������?��+�d�<I��܄O����I������hٳ�?����?!���?�'��D�঍���YßDAE�Ӡ^kvS^�j�+�K՟I���Ă�)�?q�[����ڟH�ɋ7�Z4ⱭE�L���pAa�r�2A3�#��9�'=��ʴ�M�?Ekњ���w�$�F�F�E�H	#���G�4=�'5��';��'��'���mR,��#F���LR�M,P��s*�O���O�]o�g6L�S՟�Y�4��h)�5��/[:{���*r�EHR ��N>)��?ͧY ���4��$Z
HM�5I�ř)O@~ب��� �Q�o��~b�|b^���	ПD�����	��4R<x;d��2� �(Qԟ���{y�h�
]�PB�O����O��'k���Җbҽd���D����� 0?��Z�4��՟`'��'d(��oz�=�O�+�� ��%�8���;��4����B�ƓO�YR�m^<jI$\�pK�s����T��O���O~�d�O1�T˓M��fN�9�����˥
Q�4
�b֖	JP^�p��4��'��?y�Үu����#U�h�$2Sh���?��Z˞m��4��D\��b�P����x��	�h�0, �"����yRY��������韈��ǟĖO�HP	���.���0 �԰#!.��`�cӚ���a�O�D�OJ��
�$��睽*���� E�H(7�����Im�ŞT�@ʦ�Γv4%𵤟�2���C	^���ϓ_K��c�h�O2��O>y+O����O@2��'1Ĭ�G��gv k1��OT���Ov�d�<ac�iY����'.��'� iP�H�mx<r7��/:�d)W�D�V}�'��OR�Ҁ��,��� V�P89�҅A���!�����e*L;i��O����	:i�BH�:��� e�h־<Cue�����'t��'q�������@��J�|�r�����
�؟(zݴ_�n�����?�G�i��O�N��O"Ĩ��W'�Lm*�-�"��$�O����Oʁ�Ja�J�R�Jm��?� |�@,F$Ӱ��T'2�YT�.�d�<����?Y���?���?1��L"�0�-��O((���.E,��P���!�����I�4'?��	�
��x����N:6O��Y(�0ҩO�d�O̒O1�f�#ծ�
DfL�jgӯFu܀ʇ
N�] جT����U����i��_y�ň+8�B�Q�@�8��&�vn2�'2��'Y�O�割�MˣOE��?1d �*�akuׁ:	
�����?	F�i��O���'5��'�fD�6r@�Q��T����ݎ{���:�i)��2w{��ڟ쓟����59��;�BX~����Í�1��O����O���O���=���- POU�8��9�.�e�t����I��M�6f@��c�v�OzT��J�7k���7ķh6p��'�d�O��4�꽐S�u� �Uf�#V��<E�CF��H�����iT�	m�	tyR�'���'�r�ϰbk��C�ץR�v��g�D�uQb�'|�	(�M��1�?���?9/�Dq�!�2Z�<	��^�Tߎ��g��T�O��D$�)���3,�~Y	���By�[�5~-�1�3�˅]j�j.O�	O��?���0�$=Q넨�!hJ�U�N��C w�p��O����Ot��<y�i�,l9� �Yy��AA8h��v��1#
�	��M���>9�/�Fku�]�:=�)��
V�����?�6�Ɨ�MS�OH�˖O���M?���g
�%2�l�eL�)}�rx��nt���'��'���'���'�S�9ټ�%���رxT�Ėd�Hڴ5�D�R��?������<���y�!�q����E�pv��@�ԪD�2�'Zɧ�O�	��i*�dM ���)���lע�E���$��D��
ZR�]8���B�G?s�ܫA�a3j��A��&�P���e�6?�0p�b� =����s����N��Q�,zLYK�,���y�R�M���O,-/wP�%���B�G���� B���$�
��{�k�
8Km*��R�� ��Ҿy�� �%ԭt5F�ѥ+;u�0����'4NK J�S����k�\"�@�dK�:܌y�&-%I���ie��\��
�L��
M�S��v`fΌ� ���+��1�Rq0Q�JV�,�������� �Z,mhL���M��?Um�	ClXH�[刌�dϐ*>�&�'h�'U2�'j�l(T����l����J��'��ѱ�l�!#���'��T��"�C���I�On�d���I�TƱ;%RT8��B�Fޙ1�U\�Iş����+>6��?i�Om<�#4��m�ܝAI�$�x�ߴ���ۺ[cn-m˟��I�\�����Ƥe�WLY�W؍�e�St��R�i���'���p��7��~�4܊��O��C�/��7�E�H��mZ��@�������0����<!��/FT��
e�Ȉb� �$���I囆c�F��O�?���,*er��`��!d��Ճ��\ۆ i�4�?���?���D��Iwy2�'���Ƽ{���i�J��m��Z��O�=[��6��Oj���O�E��.�ff���/6a"����A��.-��1�O���?yO>��e��kӊ�C�$�� � ̤}�'+��Jw�|��'�'剴HIԥa�.T68^>�`-F>VΊ���f]����<y����?q�y\�U˅a��%��i���(���#���?���?(O9��|�螮�R��W`�B����� զɗ'�b�|��'�B�Im��C-Mx4�e��%d�¤��P
4H�����	՟��'3��b�~j��-Mp��̝	<���h�Q�t{,��i~��|B�'�ʃ��'�x!��\~At��!��m�Njڴ�?�����u	l�O2�'7�䇐|�^٠F`)��C%I�e}0OP�d�O~�%��On�O����g>��!�!DDK��Y�/R"6�<AL�2͛f�';�'���ʹ>��ּ�Z�׿R��aV�I�.~J(l�����	p_� �?Y��D�0��QZ���U��M;6@��(�v�'���'��4n�>1.O��Q�@�2�D���ƚ5Q������y���i����O����9�� ���<9K�ݪ�EË�7-�O�D�O��I�bJb}�X�H�	\?2�[!Ҹ�g�L_���C��E� u�}�I>����?9�sp�i��P
Je�7�)>jv(a"�i���:L�O��O>ʓ�?�%��'����Ϫ{��1t$6A��'��Z�8��ޟ���jyr��JF��""]24�e�E-�FoI�D4���O\���OF��?y�O�R��5&��OG�YY�hH>#4\#�4�?i,O��da��'W�������N_5&��)ޜo�<j�.��y�F�'�����O>�n��o�B,�W�Dfp�<�Pe&!r�OP�$�<���b|(4�+����
-�]J3�I��p��mXؾ6M9�I��,�'sT�BK<qg윔R��hd�P�zڹ2S�NҦ��	Yy��'�&�:f^>y�I����s���GDg�0��g�25oA�NC�'|�U��6(&�Ӻ�s�Ҹp#ҹ���Ө[�dAʴ͗O}��'>�;v�'���'���O��i��V��I>C�D�<>��SVmg�H��<�
GM��ħQ%�)��2< ݂妉�6��ulZ'��	�\�	����hyʟ�)�q���VЕѤ�ȧ[8�1�E�E}rAS��O1���$ʻ[<���$�/jl�����DD��1lɟ��I�0za,����|j��?)�� !2�%�
F�HS��[�aI<I���'�Y��r���˧�?�燎 �� A�K+y�
�sd·(	�|pb�i7"��t��	��i*�I	"3�@C�*a~\IH�D��1|)O<igVW̓�?9-O����>�,�i����C�~E{�M��h��"�<)���?ى��':��צ\PU���5�-�@lF�]��fn����O����O<ʓx����28�µ2A&�2C�ޑۧO]+T���Q�������}yB�'����4 K4�V̸Q���r������?�����D[�=tt�'>M�]�'ez���c&[����Y��MC��?�,Op�$�|�����B8�k��Zp�l��)ޗ8��6��OB��<	��]!hf���l�I�?�(��E�"f�i�Ś[5`��S^�����O��d�O���4OԒO��ӳ �I �gכ$"��ˍ��7-�<aȞ3m���')��'{��ɭ>�;rz�pn
ml�1 @j͘Jc4%oϟ(�I�<���If�~�')Ŧ1��*��ے��r��n��C#�@;ܴ�?���?Q�'��	Vy���
o$ � =R��=C�˃�*�7-6C�d�Ov���O�2E p.)�J�Aו@�dqd�o�����O ��Q�i����'�����4��)��A)��!��J&����>�mZUy�'�,5������O �d�O��qQFi���0fy\i��E��M��Q����OJ��?+OH�������˘p<X{v�,d&LJ]���{�Ԕ'���'�BS���q�ؿ���c�&�4"Α�b� �O ˓�?�(O"�D�O|���Q� ��]�b��(܈sG� ���<����?������J�=^̧?�B�Ԧ�-YE&i�`���\nZjy"�'��	�P�����x# v��:���;gHH���z�������Ms��?I��?i+OD����G�d��5V��:.Qb�r���0�������M[���$�O$�D�O2�0�=Oj�'�i d�*k:���2���F��u�ڴ�?����÷IDZ9�O�2�'D�T�����
Q �R��$"�DΩjp���?9���?).��<H>��O���kg�_, xQ�@��(n�ɐ�4���K�LӨHm�ٟ��	����������G� ~��)�*Z�;<♁�i���'��yb�'��a�'Y�~�y��K�Ii`Aj��� ۰n��r�۴�?����?1��<a��]yr�-$��ӗcQ�d�����o�6-�, ���O���ON�?Y�I)q�#���#4�|j3mZ� ��Hݴ�?���?��V�o��	Ty��'����l��Q#A�Y!sN�q!�L
-����'&剧H��)����?a�O���剙]�B�..рl8�LN����1��^y��'P��ޟ֘k��,Q�T�`~4Sd�D�&�p�Jq���?����?i��?,O��a�S%-J��P�
\k�)X2�P)Vg�X�'����Е'�2�'��E�+����A<��h�
@<S�R�(�'���'��'��X�HZD�������6�>q�B`ܴM��
�̓�M3-Od�D�<9���?��TE���Or���۵.=�j�-Şq�N���4�?���?a����U9;���'>�'+�#5(��QbKo��lG�L�Ms���D�O����O��F��O��'c4yz��M�@��W�ڙyVu��4�?���;��0%>��	�?9z�MH��"l�<��a����ē�?��Gh� ��䓟�mU,*��1���K��Yq����M�-OƸ@�Hʦ�*����d��'(ڔ���김�i�17R|�۴�?���`͓�䓗�O����iۿb�T����(>���۴��ika�i�"�'9R�OՊOx��L	�%J3�х~ƞ�	�eZ�C{fl�@H`�	r��v�'�?a�HX*L�3wY��\8a�����F�'�"�'T��z�>�I͟���>��U+�/(��X3Ș� ���=�$�k�������Od�]��������i�ɂ�(_
T,Ho���[�� ���'��|Zc��|�4��:J���$�,Un��O�ks��Of��?y��?�-O΀`� �3:���0�E�;u��̠�Ь3P5�>	�����?��	��,�ɗl^|q�U�s2�Ӗ ��?�.O��d�O��Ļ<��9
�)\4��]�aE�V�z�#$ǅ�t���Ο4�Ie�Ο0��0���ɛg��		���y[�Y����	^�.5��O��D�O����<1rK6?��OF�թ4뉾A�Z��2%�z���s��rӤ��9���O����=hO�$3}��׺0��))d�&�(��d�ˁ�M����?�*Ob��k�X�Sٟ��Ӿ0���8p�ƈS^��ʁ'-Eq֙�L<9���?風�F�'��Ɋ\c|�R��d͞��'F3 ���[��Cd
���MC�X?9���?y�O@�iC��=�4���Sbvȳ�il��'�R���'z�'q�Taf%Un���㳇�1HT(�b�i�& #r'p�p�$�O��D��	&�4��2+Ya��$��,��0�S��x�ڴ��d������O�b��'4��%ϝ�&�҄h G>7M�O��D�O�8���g�����{?����S�h���/����AÏ��%�re�x��'�?���?��W-IT�$��� 65��i�+q��6�'��H�o"�	���'���| ��)Ti�;kJ!�O��_ˈ�A�����O����O��T^�|s��+{i�h`�7Js����7k�'���'��'���'o����V������P�Ĕ�yrY���	��x��ey��V�%�F�3� ��"�!1ͨ\cS���cbZ�B�W���IK�',����@DC2�FГ�'�Y�!�T���$�O6���O��>n� �V�����@s>�g�;8+NaUe^2.7M&ړ��$�O��'-�$1�ńM���d�pmn�I�Í����<����O��&�ҕ$��H��M$�3�"O�y��
��!��(N�1㥘&cv�� ��T�.�j@�9J�Ҧ�ٍ
�"A)�jǡ\5L�pb��,w^i�p�SS#HTH��I�s�N\Z����2s����K�n=tZTjɠ����^gK�4��B�_���P♁&[&Ɋ�5i\ zbk��X6�1����@�:u'���`�$QF���a�O���O2�����wd>#�9�䠛�V1R��<K!� � d�i����I�jHˏ�t�(}���:`܌�H�(ۈmz(����H��,C��p�|�x5aա�65���D,�A�r��Y���i�f1���l��y�g��O����E�i>�E{Zȉ*Fe��R}<%��C_�P2�'h���*A�5Z�0K�E���*� �OJ�Fzʟ.�??mɰ��( 8��%gFz<8,G�],����?9���?����p�d�ON�ӵn[J,f��)(�J�2�
�H]XD�ʯq�p@��	�E�NP�'�F�l!���Z��	2��%9<��	�%9��2e��r���k��Le���f/�O����O��D�<i���'ۀT�0G��R��X�F'�b�Vb�'�(u���J�$��Ma�ͩYu()�y�o�>�+OL%"���D}b�'qČ�TA̎^�Z=�0E�"Z` <� �'2�ϭB�'@�I�d�"d���٪|ܸ�Pm8��ԯ_:��X� Å�i[h��I+Ia:d�`���dը�'�z�Xu� `�� 7eF�H浑Ǔu�]�I؟Ĕ'jP ���R��� �m].,��y��'F\EH�j�y�y��M�6jƊD��'��6͙u$��R!b�$'�d�*UN��E��Ĭ<A���!l����'g�Z>IK���x��aW�"o�Y��\�v5�]��b��D�I�8)*��N�	U�dU��+�� ��]a�䕦x̮���5}�0z�R��u�׷A�*ᆓ%�Ll�k��k�Ũ%hB 	wn� ���X�'�����?�c�i5��I�1~������0`�@B-��Gr�D�<�����d(�L�]�v�҄&T�U��/����ۦ�Jش�?!��i�r�O�Dc�)�c�$�ҵłX�6�O����O����'O?S�����O��$�O��n�R����7� `i	��;CZX*��҄�����*Q�i#�|�蕖'�8ݙ7+�}�$���LR�7���O�E}R�U��<�}&�<2��-L������/UH�t�Cb�,QH��)�3�Ɵ`jX�se ;�V�8 C�O
!���r5�t�-;���6���;��ɼ�HO>�A�&ˑOr=As��*f:���цhUP��PH�ӟ��I��,���uW�'��9�,� �#�g�.%���!�X��7J�I]!��Q�`�K#��+�j�+��x�X���xrk_R�H,�V䐦?���%�ĳ"J�T ���?9ʵl�py���:<B����G�<A�o��2y��p���#�Lx�HZC�sܱO� Ǝ\����ϟxT�	`榝c��[ `]Dm��Rџ���16��)�I���̧C�~�b#�S}����OfԨ���+s�؅�bcMl�
�ʁ�'�C��#�#������c:��ц�Y��9O����'�'������Kb�mqMK��$ �'�(� �b7�6�AB�|�p1�'.�6M9^r�a"�ȣ=����n�6L1O��N�˦��Iߟp�O+\mb�'wH�!�+�:6'�0��H��fK� J��'�r�¸}���T>����&�;D�I����JI�Y�Ot�w�)���Il��u�/3-�C��9\F�'aR8�������Ovh�Ie�S�.�rSG�88~�H�'�J4b�CƧGo2=Ks��?��HYÓ`͑���7�a������I�`��Cwh_(�M���?Y��D{CǏZ��?����?��Ӽ�A��F�%�ceޏ(M���"J[���'hQQq�'���4&(`%���D,�).h,=ʌ{���ay�~�Pi�EҴ?��qd��=���'Y��G���,O����
S�Dj7ßfx��k�V�Y��C�ɂ��	�$8ҪA
�&U�n��7����O��#nV���Ƙqg.HPc�QY�B�	�x	��`oXy$��F\I��B�	�h?X����1,�����VV�B�I�\c�(d��>Rv�ґ�Q�#��B�8lk��#�ېh5��8�D";�B�)� �๓j�b%ʈ�`�>8P��"O<����*�B��Wdh �"OH�Ä����QQ"�'|�!�"Ovy����b!�ܻU�_^h剕"Oj	ӥځ�h���m@1ZNn	�!"Oll�����3�~i�`�ذ&���"Of���
G	C'V�qD, 5���:�"O�p��D�P�JŃ�dN&�SG"O���НG��ص"F�c�-��"Oz%u-)c؈��S��M��q"Oz�`�V��Dd[Ǯ�F�&���"Or�B�;�pC�����q"O�H{猓'��-�l?���b"O`P��
<L˦-c�Č�B�ظ��"O�9��eҖ4�Ζ:���d#��y�J�'�r-Z�*]�^�y�ǚ2�yR�D1.�: �aƑ��dt���y2�ƂN|MUL��;"�@�N��yI*f�P�J&p�QbSEQ�y�W �n��ī�>4C�Ԅ�y�
�;<_���j�@:9k���'�yd
}w�	ʤ��KJ&�rªI,�yr��e%�Ł�@eH�aEՖ�yb�	S��aAsσ3�]�
��y�IC,Q<!I��Ϋ��y a����ybF�#~Z0횰�Q	EbΨ��դ�y� ��bx����?�x陑Cȍ�y"�^<{���d�K:U�� ϱ�y�d�5��P#7
�c �ز�y��Ԣ�Ωa�^%"ЃR#���y¤�j \��P�I�uQ��y2IU'Q��p��D֮v����iM1�yb�0$�HM�V��;j�0��%��yBkCO���0�]�|���G��y"*�8$���#�"TF�A ���y���;�dڷ��6 �� P͎��y���4g�^]Ckx<�pS�B'�?qB��$0�d5� uЖ���`X�]qE��.Hy�.��L��9�f�c ױY��xJCJV��H�7a�.�M;2#G0�H�H�h
	��d'�$⮰���XF���j��#��]��I�9(�Y8v��%db�����5=�5RkX'��h�"lH�[��@R��Me0�t@�iY�l��a�2�Li�������>���SB��d���q�X�0�)�Wy��BO�!�#M�A0�pW,��%A�\���.���m�b㰘ۂ��/���"��	^��+2��m�L��N<%>q�3�Hp�7E<Z���������"O.���D>pg�X�Ξ�]��-z��|�Ǝ���,x�ᒟ=�@�sN����'N&9z�kT�D�,�����S���ϓt,�����6%���l��Wrn�3�D�<
�q�&�&z\ɲ'�Cϴ�q��	�:�Ri��I�$��1f�O� ���G�A��O ���O�c�UHv�M�&�!#�;*��YVG�:���c�x�E{҆K-g���Q "��t0$�,,�;�b��G���bUHX'Қ��޴!�Z�'��OJԹ�w'Ψ
f*̥Y+bP; �Hȵ���d��|�5"�w��������h�%群��o�|o��2�c�8��ɲcx���a��̺k0㐲3���ۋ{Zuk*{�퀮>�~I���<�&ʓ�ꈻ�!��r�qO��ДIT<�
LBFf]�=^��u�=P���@mΙH�P9����p�a�Y�HT�#>y��(��3
y��$�!Q��� �ǜ/T� b���ό+ ��]"Z���f�<��]mҤ����:Lݸu����F�4#>�0�L�p�y�I��q��Ѳ����FP�0�ݜ���K�`�y�dIC�̗��O���݆ng�9�˲�j�R˖�#�C�	'G�M�.�+t9�7k�\�qp(OT����όY�2q�[w;L�&�~��c������4�z4��+�"_�4\��I�f�xZ�Î�kGTsQ�7�pơB�d��-Z&l�$�p���!�*�J��'��h�TkR���l���Y�\Y�r�}+G6#\��aB�	��`�I�6���O\� )���-aź-q!j_T��|���� 8U�E��;�pU�P���P��C����i� �{5"Uy���+t����k�p��Hc�]4a��\P)4D�P&��4I�Ս�5��A�� ���IW`��W����)'tb�@@�g�]��sG��SEvػ�"�O�\����j��Ii�!�\�$�8�T�b&��\`�T��r���r���x�B���<�`0���|џ��w��+}�� ���N��,B���v�Fq�dW�0�������V����65�\P��s�x!�D�( �)�<!�T�h��(bW+�%�Т|�s��� �w`P�"�X��Ee�i�<yU��^���j󁜍��TE���*��q�
�v���I�j�4#|�'�4Qy�B�3T��0:��֪|�����'��tA"��7"\xh�-{�b��[7dr�Ir'ʕ�v_�@��	
HZ����_�v]5���U=����V�n	�{�^AP�B�B�\
��9��Al���!��H�!�dB�o$0�T
�&\|�X�F�� �1O|�Z�N��@&��B*��(�YA���P��P �m�,]F��"O��p���EF���DU��rQm/3���S`,L��~B.�����I'~v̭aP͜�M�J�+�0F�bB�	,�|�c6M�m,��끏�o�B����"[D��ª��^x�zB`�3-C�
�ʷx�����^-�0=q�K8k�(�b�Bc�hadJ�=P�r�[�	�7{f�0 �g�<A�L�<�x��I[�$��.�`̓	ۮ�g&�$n�yɰ�#ʧHH���G�h�E��<c�$��ȓK~��"u�	�`�BU�%�;m
H�`�����	�&��hQtH+�g~�/L��*A��wl�|�gGE7�y��>nMT�I$�%,� XQVß!vH����Lż�,Q�6�u����#��x�vM���9�|! �#7LO�L��<:>�ٕ�X鸅"��vޒ�c�N�J�b�s�"O��k&��#Q�5�0�"B�j�����h�Y�&��8���M�&�L���És0����o�~�!��X2��}Ip�˦\)l�yq�T0q��$�U�ε@��m��'&���O���pU>�\6�Y�����9 �
��0l��	�P�F�'}HH4
�|jzp�	9���[׏�4��<�zr�ʞi���x�P00���,�=c �\X3a;�	�O�M���@?��$�#��]Z7i���u7χ���D 0MN�ـ�Ȧ�Py���VZ������U�1�"g׻hP (�i����$���e���i�ۼsugI'�0P'։0�I�0��|�<	�)W�$kb�C����2F�)&�߁ ��0"�PK
�(-O�.O�@��<��#Z�'*�i�ύ)%9��y��z؞�2�(��\/8}B��'�|@@��ԅD��	��� ����'�L\J@E�@8��2��R;�`ؘAn�t���
�$:�I~�$����*��	�4���ܟ�%8�HM��D� M>L4�� �"O8�$���C�g+�Q��!�j�������<�E�R/N�8�?U�wFv�zR�@p���ШP�^�J�[
�'���Sn�98n
wē�Uچ�xv%�*�6����iݩ�Ub�q�'~d@�p��D��;�C����
�����G��=|�D �(�v-��Ň� i$ܛ��Y�X�dǒ(�|y�P�&�%D�>�4�����UV�g�`��I�ek��!Ɣaq���/eӦ6mъK+��ݘ4 Z�7��y��9���#3��B�	D��}� L��Lt��ߤ]	�yB��߮S7�3�M���B��!����$!��ʧ�
x��{^�p���/f`u��c�8y�@Q��'�|� /�sy�˽3o�����C �x�	WA��y�"���<0d�W�0uz�۝s�R�FyB�%�M���:��͂�-yy�>�OKL����ѫ�V����,�����c.�S:D\����RM�t,<}f�2	��u�g�~��� a��9��ە�J7���1�n�'���i[hy�7�>�*���}pl͛��Q�7"����"O�A�O�3C�lMї/�b!F,�^py2MO�8누�'}�91@æ|��[�C�G\�^��e����)�x�#!��G<a{i/8� ��'-���"A���2I�0�����Z��
V̵	j���SDM��Dg!ʓ{ߪ̘3F	���"ұs	��>�p�L"���?�ɗj�>�� A$�����
6K@�%lm�(�V��	d4$|��$E��Չ��6Z[�ACBK҇|�HP� I�x�.`��}R_�ͻ/�P\�� +@߮�b��R�M�I�ȓ��HC����$�� w�ʤ$�T�5��D�(xEJ*0W�MHvB���&� r���.<�HAA��Y�oq8��W�'(�<i�%�{|��20�	�\��B�ϐn��L����Vn��ú��7-B.GlZ�C�U W*��Ey�ȝ<�rl������:=�S��7��'��*�7rȵE�#?�~	�H<�[^`�0���m��,�$���j�����.�.�q�N���E�����E~��&�=Gm��� N$iY�=�{?Y�8��E�ac\;�� D'���H�e"O@�cb/� �<��eCQ��0��Q�X�L�_w��$�ȇ�Z<l)(њ>ID�8$!�S���n� Q�S/A؞p��E J���"���X"&�&�)�T(9�%]F� 3'jR B��0�C��s��$c�C0,O왱�Q# [D��9	���u�D^"b�~\�c�V��m���`��h����oQ�?lDQ��������'6���`�pF	�u��}A�`�ri�)K�vPci� 8��9}J~=���KA�gz�K�jF�_ۀ���"O4�b#͹N&�0�'��N�h���NSQ�D�;D�Ђ��m�A���LS���=�!�#:~��WK��HĹx��`���+�L���^ �%㙳i����Bܴ ��Ũ�#Ә�rgۑz��L	f�@�J��G8���`B朽'��S�3��< g��0����Ō�;�*E)��<��ߊKf��W�>��l��B
�yBG��v�X ����~t�Љ�w�MiӁ",���C�}�S�@tn�.�%��7옽w�nzCYI�!�Ĕ��|(Ռ�4O�q���A�dB�&�p���Q�Q�B��U�ڧMhM�c!�Ƀ��xB�F�{�|�K�>k���򄆭w���� J<V�y4���I �eƦ�	 :I��C�1�r؛ �K!�J�r���]�a{R��{D���%0 ip̊�#���� ����W }m�|f��px��?�ҵE ��a��,\!md@qTF;D�TY�@P�řAb��im�xU|T]�@R�չ���ke	�8�|c?O,)��-z��l���H1\�Oʴ�aO�L�(UY�`C�cV4\J&��XvD����B��6�8bM�E��H�r�a�-z� (�<{��+<O�,x�1h+=y���hW�}k��E�DY��݆ `���� +D���AE������� �XQ2l'D���׃�Mk�d�ӧ�
OEQB*O�e��j�͑!w���X�"O4�Y�L��
d���چ� ��w"O�@�ҭ�=�{�KC�G��,h�"O���L�4��V ��y"O �+��^�y�
H�R��6���#4"O,�1Ѵ�.0�DS-�m�ܐA"O�(� �0���q`޵�ƅ�g"O�Q{�kր'����d�θ%��!�"O�ɪ#زP$­�c��
���R�"O���L%�F���˄�2�l4�"O�p�0�З����k��� �*�"O�Ha7��t��2�
J���3"O��"�͔C<\���_ c�|�ز"Ob\x�. �_�`����1�h��"O�hcѮ^L��G��*-�����"O�̀��ɨ Kr4R�ɉ�^����"O��g�0��}��I8`���"O8qRsg�-n�5A`��F�2d0�"O M!r'�\Ɛ9����0t�UZ"O�)�Pc�	dQɧ��oqRE)P"Ojp8e�S��ęP3-z�Jq�$D�`9�i�<=��	QAS�7 ���e�?D� �5�F:nOV������!%��>D�0;�Kĺ ��,3&BL6dμ:1�<D�`3���x��]t�0�4�=D���Otnr�a%��l��bK/D���j1���5h˰~_0IS+#D��1�TV����A����釉 D�XC"J��!�r(�Fo� 	������?D�$�%���?z�3�n�9I����7D��iD!�,�����:}cz)�A)8D��Ԏ�2��+��i	P��4a9D�� �h&���_\�* ���a��R"O�XR�%k���b�e�2X�v"O���v�)��� �ɐr���%"O��
�+�#~�xq!.VvX��Q"O�`�c)l�n�[�̖�FZF|�"O��$��(^'Y�6���B;�m�"O�Pʴ*��x�����6=��"OT ��jп]�����!�S��g�<饪����!��F�	�f�R�]d�<1�/�� [�Y�g�@�5�p�Rs�X�<�3��M� yHD>�Z�r��S�<	�a$�	@)�9]�HQDS�<	Х�9V*j��2� �B648�dPu�<A�)u��"B�и��*v��n�<��.�,���x$$�26�H$����j�<�P�R�,X�@�I�|GHx6o�g�<)�K�__���,j:�ų�aa�<�f��P�I¦	B��y�0� h�<ACA�oوm9���Y�L�� hc�<AG��$B�h��S�0JJE;��D�<Y@�B!C5�z�'�
�����)Ik�<��+��2��. �z�$��! A�<9���Uz��b��A�a���"���z�<yt�_���*w��ev ���� D�VA�aO��#�� X/f�A$����y�nuU�)� ��7W6����	I
B�	4�q� J
�(�R�8�G���C�	\Hघ',H�A���	"�K�C�ɰlT�#d�G(Y���p�ϦX��C�I�g�F�H�N�u΀Zm��;  C�ɩk�X���^ ]$�[`�:��B�QVj�b�ڬ4���3n���C�I#�ԕ@�͕�E�=&
 )��C�I�Ih��C��-q!,,`#.޻z�C䉭,v�m�s��-\�\*!��C�IG�l9;�)�~#HY`�[8ck�C�	�|Ғ��oμeۄ�(�G�2!!�$� `cL�[3jc�aV3v�!��3I��@6���17�1G�\G�!��ح^N0s�W�wE(���W(w!�]-�¹�qNF<}+0�����Ad!�D�n����q���>�n�C�ŨmK!�d��}��L��߭�ƽQI�rF��!�O��(=KU@i��LH�~2�Q�"O6�t͓�|i\�hA+~u���"O~��f�Ol-���8̸Q0"Ov���sQ��b�N�GN9jq"O��p&�Γ<�z�LP/cd���"O�8�� Cb5�4^'���p"O��QoR�aG�x��é8�	�4"OD� Q*��YA�H�XW��pp"O��`�(�FĀ43CHV� 黣"O��`Q��2���{0�������"Ov��#.��c�ZD���&gE���"Otx�I.Ƽ!��9[#>X0�"O̩�,:,~�s��c����6O��=%>��OX|Ag��A>�r'eX�j�܄97"O")P+O�I�R �hMyg"O���!m�$5���P���'"O�͊c!>2)5�УRZx��t�'�'%��"e��0�+۔�:���B�	����w��(�d/	�0�7"O"�
��@.�.DӀ�#v[��s&"O� �P�F�@�A�6^&�Y���
}����
� 0A�v��%pR��/ۤ?����"Ob�9*[#z��҇싮�`��C"O�Ka�
t�!�+Τ����"O���FE�c1�d߳Q�RYy�"O�����X�{e��<J����b"O��,mk^���k ��"O4M��P�-�$daG!�Z�p���"O���#�����/1OF)�� ]��y�&�q���z���w������yb-�E2d*AUtr�ё#���y"'E�<��p��.l���Ɂ ���yRa�U�4�۪Qp� ����y���:c����'ΣQ���r���y� �?3��As�D* �\�8sO�5�y��2
ƈ"t���r��щ�/�y"J	9Xg p�����\򁐑&B3�y"	K=�J���ˉ�R`���L��y-��x�h8�F�VX֨�ɢg *�yB���D�1q���]Q�ȒBT��y$�pH�d�^�W��%2뇄�y��,��Kh�2\�(�0f���yB�G�RL.0F�<
`V�C�m�9���F���O��QY�h�-N`J)p*K�H5�Y)�'������?�B���YC�-��'aN��w�/P��ˁ<>f]�	�'��Tॅ	��l���,ݲ���'ᔰK%�*n�\�����)EDZ�'�ƌ3��Z�@ ����Gւ(8t�'O��U�z��HY���%
׈�!�'��`��e�P1>��Ӫ&����'^�I����;Dc�-�F�@�}�0U �'�2��0B
&X$%�va��If&�+	�'r��b�C��S��}?<����\�<#�[�����G�~VE*��Z�<A�C���@FN�"� �ۧ%�T�<i筇0#�0�Qu���{&
���M�<90�@-�X)�aˢ-	L��c�YO�<��c�!�0�W�%5�����I�<Q �8o^m�vADD����B�<�G��9�q&F�4����ti}�<Q�iR�KZ��'j��K��RPoy�<i�/�=�v`�gEen�U��.Eq�<q�[�L�� ���-:���d�Un�<9����v$�	i������Ypb�t�<�aU-@R�@k@�ڰtD8��kEp�<�e� ������o~���/	e�<�v��o�E��.Ł7˪��@]�<�u�Wz�NP�D��XV<d���t�<�o�&]p�	�`J�*"b�x�!�o�<�� �2aqnX9��էB�j�JnDT��hO1�H��W��iv�eZȈAy8}��"O�}"���4Dm��'�
#/�J-h�"O8Y�3f�(%����s�!����"O��q	̳N"���gɆVV>�p"Od��F$M�/��+��jO�KB"OU�q#W�u�r��Ӈ�{Cx`�v"O)Z ���E�V0��J|1���q"O�p���ƞ��E���s\ ��"O���"9�L�1�/|\�ica"O1�Dh�*h�`aƥYW�1�"Or��&�4�!�#��lx�"O�١�l͢Mg�tH0�Rz�^pq4"O�����0]�D�zF'*�[�"Op)1��:S^�}S���9�r�i�"O� �� �^;t�������c'.� "O�1�G�˔v��뎱h�R�"O��IA��:���d���P���"ONaB-O�&�A��P�F��(�p"O�y$��:M'���ugz��mb�"ON�*S.ϛY�>���
�$�5"O���t.�	P �D�4)���B���"O�+gJ��_�����"�����"O��34M^�:s� '�ħ�5Ҥ"O��X��bLiEF�JM���5"O�����q#]�R�A�{�)�G"O����/J���t&�&�=�7"O�xb��1t�P]��D,F`d@�"Ov�Q#GLq֩PqX��E�"O41k��Z�IG��(�	�~�l�"Oư�`'	(hx):a �W���&"O���͖8|'�Sq��<R�"O�����T905��f	q�S�x����T�U��y���{�h�'_z!��0J�֬���]++���"�˂�!���<	_�����!1��� $�!�d3qZ��c�m/!��`K.
P{!����N���g��v����l2[�!�D@�%wF��A@�A�\���8�!򤃃>��\����'l��顫W�!�dNk���Aq+MF�@=)T����!�䅐p�Q�#�GlֺH	�آ*}!�$=)��!"H�?B�|0��I-j!�$Z�E�x}z@JO�c����E���"E!���xR�e{diE�Pj�A��'�!�dl���h�>C&�s�P*2!�U�-��pwG�
��)�ï:�!� !>�p�՘@�2dB���2�!�ֻ�RL���6~.���@<"!�S�X�����b|z�|����d!�ӑxٔ�D�dm(̋�&Y�jS!���]�>�+&-�)Q����� 5!�D��h"t蒅^����!(E�2�!��<n�����N7b�J�r ǋ�j�!�$2)#~��Pc�A�Zh�E��&�!�;$�xhE��0��C�'��`2!����*u5�B�P.ZV�|?��ȓU��0���ťU�@��e�S,���ȓ=�"q��:M4a@�h��O�L�ȓy��𠊸v��X��^����W��ò(�����FF�.fRɇ�9�N@@v[�-�h�W G-6�
��LrQ�w��]}N%:d��0,�b�ȓ���k�- z��	�e�4=�ȓFd�1m։ƙ��"تڰ�ȓ��h�s�A�P��S�,=����ex ���T.5�A��d�8z���LXpX8Q �b��*��b�-�Q�<�K�j�5�p ,)3��I�gKN�<q�eF~=��K2�E'y�EQ��J�<����dْ�#7.O$z���p}�<	g�ʀnm�[S��I��Br�<y�o^����1gH��
+��� �y���!~��2��W"U�tY!R͎��y�$ND<��[��Ғ@��>��e�&�c��"s��1+���2#�漆ȓ-���t�̤W�z]Y�M%w�R������Ckԓ(;"���T�.j85��x�n�QF�(�� ���6'�6p��S�? D񵎈8D��s�n}���"O@qH��L�^�X�q��_�>D��"OĘ���E���q���  �D�	G"O�����4YU*,	��{�����"O,�
c2�2�F��<M$�f"Oa{Ճʶ>�-���9��=Y&"O�@e�+"\ q���&���"OxM�DI�"�rx( �-h���"OZH%��OYx��	#j�H�"O~Q���͢�J��ǰ4Wz@x�"O��(b�I�<��Ԑ$�C�Z"O�x
��ƍ'�,يRÙ(E;�\I�"O 0���ŭl�Zd��Z5"21Q�"O$-zd��B�����&�J5"O��r���T��u�C��$bZ��H�"Oj�����(`B��osR�I�"O��u���H�1u"؟F���K�"O4,A%1�j��w��N��}iE"O$:2�\����&	jh&|�7"Oֹ(�"ݩNd`��� �,�C"O���#�f3()3%�/-h� �"O
-�#�X�p����"�p:9�"O~9���L�CV���1���K�8��"Oδ:rfѽs���/��D-FM�"OxXs3��?-����T�85qA"O*i�� 1j���hB�zt��"Ov%�'�b�ԭ���ԟ�֤K�"Oء��],bh (��?��]A�"O����*C1a���;��Z(c�h��"Or\�Q�?m�4ъ��;��\��"O4�Z'��7x���)�ԥ�D"O��;�-	?Ђ��t��wP(�S"O�X��
;-4��b�g?�V�{�<�҇�	j����K@��8�q�w�<�v��{	��ҫ�lNZ* \�<���C={W�����X�z#�=�d�[Y�<��]+yƨX�nUb���1��[�<�$KZ?R������j��I���o�<)��FV-��I�C�!̬��@��o�<	��^�9G��h# ��D�Y	&w�<9"�}����O�"I0��#P�n�<)��ߨ]R4���	dRn`����P�<���ԡ@:��˂ m����&PL�<a��:x�<��튞 p:BŗG�<�P�v��&�]E��qq��A�<���̰[��A�&��w$�]{�Rf�<ᑋ��G�(!�@BH�$�KT�Vd�<�Չ��2w���s��(�V]����_�<���3}n8zW�C;,X��3��g�<)�cV �t�`�2-BiQ�/�{�<Q�L�oZt<!�-	c��$t�<iF���ё��r<�@1�ȓ#"z�Sĩ��N�lX�cfQ�|N܆�@Sl�H�G\ \2�m2T-G*Ȃ���paP10�c�B��*�NM�pr:���~࢘+����l
���,M1dU�ȓ7DJ؀��΢����C�/դ	��=�ͩ��û%.�1`!F�	"�4��b�|��Ӈ�����U�E��ȓ\mZ]Xe���<�~X*�B�T��E�ȓ5�D��əu��
V�R=}����4��Є4P�����e9'��͆ȓ%~uSf`�'VQ*�	 �/Z܄�z8�Q��J�i�B�9���&�<p��S�? 4YJ��
���йS��@sN @�"OX	�׏S/j��a9�}S�4��"OJ��'
�%����*�QPفv"O�@�$LD�~}���e`�;|2"O���%\�H�	d�ɣ���Pq"O�E����@�o Y_����"O��!�"�{p��@�af,A"O.�s'��X�h��5.p��C"O�5���DS�!�F4<&�7"ON\��1|����P�B����"O�`�`� x0����@;[q\P"O"}�e`W�q���Z�e�_t ���"Oj�RC� !!�"�"4i.%��"O �2�l��_�$���N����rc"O���P$k(�D�D�#�l��"O<�R�Æ'�%��CßH��dr"O��ІJ_�-���A@|$�*�"O0 ����:��T)U���;R@I R"O�}�!l#��F/����ru"O��!A�ܷ�Pqtnˌ}~��S�"O�Y	w��
D�x|����!yL�ّ"OV��#�+�J b�$q�<��"O�4��h����W��'j$%"O֨���0B)��`��M|\䑫�"O�س�U�,��8��@\1n\ `��"O���KΖ;�F@Oԋ{;����"OZebd�m�a�&G�
L�"O���P��B��xK���6�Z0�	�'$��Z��W�]�����d�@z�]��'����_I8��%��9V2@Y�'?\��w�e2┐@e;�
q��'�4��^�5�&E�BC_)+�2���'��p���ZuL<����:ZTr�'8Fi�A��98Ԩ�$��_Ҍ��'�"w��[�N����0
(����'t�iC�kݡDp��  W%����'����C�m} �0��d2�'�lB�!>jt���
�%�@H�'C.���C�/n������C /:}��'�>��!E�8��ZPaU���,��'�!`�'�72��-8R��lMĄ��Z�$��H�)�ƕ��?)����VpK��w���"W�� F&��R�`x
�,�*J|��@!�@.$U�ȓi�hc@U�|9�mXJn��ȓ&f�8u�:�m(�$��b�I�ȓ,�+풶|��)���_Yc "O���a���fD�IB�=jx	��"O�:6BNO�aY���:\I[C"O���AՔm�=����3�U�"O.d�1�N<�|4�0�%
�(`P"O�E��&7$p!j��ܠ�@Y�	�'{��[� /�v�S�'td��;�'p,�kv�\�w�z�!O�lg�$�'O�� �c֦� \�<[k����'3<��'!u
9�`�$XWBy��'�<����7Us|�!A��O�����'���&�A�4LD��l#pJ~(��'��܊��z�! f�+:���8�'�`@3��K�(�����9���ߓԘ'u��&�U�G��IS��B����'M�,c�-�)j{��q������	�'��8�T�Y<y�H�پbˤ�	�'�
4xFh��>>�)Q]BP A7�VH�<� �����N�����b 6t�"O*�ipꟀ{�ʀ� S��0"O�뒦[iz��gcz�v����'Fў"~J�n���f�c�	��;�~`Q�f��y�&� "񇇙,=�5S��ً�hO�����&r��CLք=,�hʓ�!!�$W�_�p�3
�r9L��h�;;!�N-}�p81ɇ5#vd��! �4�!�$E�:&z�F�=R+�@xy!�D�,0�x��kB�Up hML�X���b��(�����<o�P�o�8�J�"O,�`Ώ�q&Q��� ô�h�"OD8�0'�n���%D�o�����"OF���T�	!�D#F�P�i���B"O��X��+X����Xqz"��"O�e�T���\x\��tʗ2Uo ��"O�`g��$i�����.в��'�ў"~2f�\�[�N�١���XTΰ u�7�ybK�`k��Z��HF���MO�y�J �E6���8r��4�Ulޖ�y�g���*�i�?^�e���  �y���Iɒ�U�7T�Ը��J|�<I�#L�_R���d��Y�X��SE�<�p���{�9j0C9)Yܕ�d�M[�<)���Fu@��/||(YkǢK]�<��D�����Iu�+E�c��hO�Te��z�DW Q�M�Psr��'Wa~� G��|��O�&K�f�k�I ��8�O��vCǖlp�����͙c����"O>�Ě I��_.\oz���"O@�H�+l"��F�9je�q�"O��WoΌOl�q�N�(Xr"O�N��D��m3�ꞏo�\t���'�!�dRs� �C��9.���p䊞�!�Ώ��.1�x�1��_��@�'3��a�˜�4����p�ʱ6�z��	�'`<��Fw�&��6g�_P�!�'ߎQIU,���x��UǄ�Q�8�(�'
]"$��%�(�bƥؗM�h,Ɏ��6�d"X���G�1��x�+��9�������	ؽKF�-��j�0g7긗'�ў�|��5R��i��e�.�����y�<���ڀ���ތw-�/Lo�<1���4;Rm��
�Rdj�X���i�<a�g{5pmz�
ɊBDZl�ӧg�<���=��y�Ί�)1�T���j�<1��O<.�H�QI?RZ�:W�Qh�<I0+�|X[��F�<��J��m�<���(k�n�H�7�h�[���b�<�pED�sk��pʐ>{V�ؚ�c�b�<	7`l����da�%1��`U`�<����+&��.���Q�!g�q�<1 ⛴�"��d#H7}m�:���ly�|b�O�hb"@�;e~�%�1�]06�x;
�':���WF9&\ވ�a�QQ���
�'.>�r�;,�}!  �A��1�J>ɉ��	�"*~B�	%�J���\h�GY�X!!�)�y!�$7R�Qd�!��$@� �q�V�H�xz��Ęt��yR�Ih6����TiĖы��'����2扔Wc2�0�.� l��`�D�SF~�=����hO2<��.�Ḏ�ޚ4�\�PeA$D��P0���x��X�pW�O�R�x��%D�0Kf��$�B�:'��t���� D�� �xy5��Ovxu� ���`+�<:�"O�m0�/U	SG�1
�G� �p`�O�8��ؿ�,�hl�"8��m�'�;�O����E�J��uؠ��iф�W��B��Q��EB5YH2�@�� lړO��=�}:S)K�O|��O�!�X5��H�x�<A�CT�J!��TEL?6д0�k�s�<)�bE,kR=��^�L�"j�!�D�<1bK	;L�I9"��->�@&�{�<���Ѡ#���Q�(ۀW�>T���Fm�<�rC�K�T�sv.��/��)e�T�I}�x�a!@�6��|�G�]�o�I0%D�`��n��;2�[�W���
�!D�TBciH �:��殘,K�{7�<D�<��,�>"�^q��
 �n�[�j/D�h�$� |�V�أZ�4��N(<O�"<���� ��P�tX�oR���vD�A�<!uB�$b��H��WM���5��|���0=)Q�;�����w����̝M�<��j �>Lj&�FI ,1��@n�<!5�%v3P��w��]de��-�g�<�ы�`W(A �	X�F���I�<�qo�(+��01KX�wî\�p�B]�<�Ɋ;q�>i�c�	�M�B���&�V�<a�,Y���D��-[�a"�SQ�<�Ɓ�%�8 ���0n4nұe�L�<�8S��,�C)ɓ���I�gG�<��Iՙh"tu[�lr���!�Ey�<�ҥŰT�\q�H�<$kT��i�<�C�I%.��%��F��,����Pf�<1���M�AZb��"B�Z�RS$�^�<yӇ��@N�a�{/,D�g�P�<%c�6<d� u��//���P�M�O�<��,��p�N�Jp�!���`�N�<����g�2l�Fk�@Ȣ`r��H�<171�de��XVHђuLHj�<Q��_�@����LEq+�³�g�<��]�0�Kʖ�$�5JGf�<a�k�8Ea�%ܒ_t�5���Re�<�`A��J8�	s	�$H"�zAF�<�q嗉N禍�4���PWڙz�I�g�<���4�4�u�ׅ?��]�$�d�<q��R!m0̩��(�"$@�Ƀ�[�<��-J
+�x�cP�zƽ�d�GV�<�G�SR�ޔ�* 
 ��`1eeCR�<e͗�R�0�*�#�	s�Hq` �֟�F{��I��pP�e�bdڢ�%%׌#=����"OrP��� ~$��&���)Q)�yb�A	hr��ҧ��*����E͗�yBL�
�4��N�N���r(T��y��ڭ+�^T%	
��VA�w���yrnH�Y{�6�Cmz�!"
-D��c���
QזiI@!��\�`6L�<����S�I��D�W��Z�hXh��E�pC�	r���+�.�Xx�r��;�>C�		�R����Ţ�H\�`GE�F��C�I�u���D�(>��@�B�7��C��&�r	���I6n�q��T��C�Ɏ-F�e�4���L�I#��Ɇ��C䉢n�&��'�0FN�$Pt�2�(�=I�Z4�xJ��M�>yHT���kP�̆�`[�1�	V��
�����6 ��9��:�4ړ�BZl�� ��m�<��ȓO��\���� ��y��D8q����S�? �&�F:'�BhJd�ǨiԼ�1B"OʨhǩɺV�����0A�$A�V"Oby���"�	�z�c�"O�U#�/��H���&>��r�"O��Z0h�H��T�F�L�)�p	��"O��[�@�W��P��hM��Iq�"O^1 �fӾ_��i�X31�d(�"O���N##��%�a��?��1;�"O��d����ӖԊ�j�)�"O6�+��'4o�����Q�t�:��	z>��@X4E�����?��C�1rc�Q�6�;0���*�C\�e��C�?m�踠�����:׈[�Jf�C�	w��%#�e��bb�����&C�	<L��t�D��Gn�R&*lC�Ɂb��RFՓ�x����,����4	��r ���]:�U)3J@�\=�O�=��´8 ��]��%���%	���q�"O������n�*����C����V"O��r�L����Ep��4"O��Θ�tٴt��F�7�5['"O��gGJ�J����+�1O�Fp��"O��RagI� ��q�k;9��z�"O^Mq�+pG�4a���82����d/���d[�m�vi .]kn���!�dG�X�`q��? >��� �o�!�d_+c^"d�f!K$�y�#��!w2!�֪,v^H���
e�t��(ѻy!�$��8Q!�gB gx
�[s��+m!�d�6m_�d���O��5��T+_^!��pМ�n["F����j�4�'�a|rf�>m�tus���,�jİ��ɢ�yR�G�jC��ӆ�"]���
3�H��y�U�R�RU��#�DF�;��P	�y�iZ�:�b�k�Nˊ;��8k&��&�yRM�)[� ��2EׂHMrò�ӟ�yb��d^d�s�K�2�4Q��y�M��D�ܓ��Ы9=�0�%���y�-�l���E�d(�p1�j���yR#]�|޸���X�.���]0�y���8.d����� 1����ߛ�y"(
0R�`=H����`ʐZՏO�y�`�K��q��
1e���T�5�y�茍1�āY`��tADis�n�5�y2�w@���i���������hOq�b��v���?I�)6�*0�(+�"O��� 7t�+�J�T�D�ӵ"O>��k)(�jԪ�)�:q�pq��"O�,����;� q��cN !�L���*O��{���	fq�A��DrO��j�'z�L�7j��5����E�Z.y�'��0&��e��|9p�H�l�x3�'��xPD�*TJd�xw,O:R�����'~��F�)Z���F@�T�j;�'�(�`A��k�f���a�?�{�'���o]�H-:�q��
+Daj�'��U�
N�qq��`aj
��Tr
�'���ش.̺��$�p	ˢH�,@
�'s A�2J߸$'�l3!�O�*�e�'��y0���b��,����y��L0�6��Wi�V�� s� M(�yb��2\��3,ɊV}1���y�[����C2��7V���0����yR�%#�}�&#�K�x�(r�5�y
� �H��H^��!�3�!\��(�"O��Y��A>�0řv�c%���"O�s���y<�]�uϨ<0�t"O2�����"���r�B�w�!Ca"O�pv���p#��
���T"OV��5��4y9��:�2C�شa�"Ol����_�\ӂF�{�p�3�"O5 ��#� �֣�6"���#"O	�m�7���@BȷP���C�Iu������h�"�0�-�x�|�g�
�}�!��D-G-�D���@��)h�� �Q�!�_#G�LD[Ef�3b�"�P�o�"jc!��L�����U�g�m2DOͨ?P!�ތ<��3��ԑh�b��&�!��'OV��E�(Z�z�R�I�8H�!�]�ņQdmCX��u��+�6�!�D����ôD9[���Q*�a�!�d�=�ځ�R�-1"��BJ¹�!��I��̤˔)	$<m� h�/A�!�Ě�0Oz�A�M'&缨�B>N!�$�2�>k4*_�E��o�)p!��
��`-��x����+Y����%"Oz�$�;Uwࠒ1-�P�f��>ړ����*�ڙ���Q����kU�݉,�!����sDh�&z�|�j�U�d�!�r+gD�ї)\�x�9����!򤐙,�� �"zP ��Aw!�Z8]�|z���tiހ�a�'<�!�D��m���@�Ij�]b!�YG�!��aS�\j�G�;!�n����Gl�U��(�e�a���;+H�@��M!t}����"O�Lk����cI$tj�h�"OZɀ@S�7��LRvG
�Go�E{�"O��:��,(�.��g��NY4P��"O�ҁ�ݼ~��:���yR&���"OQ1 e�.�41��UQ0D�3"O���3kr�<�*2 x�X"O֨��f  Xn�"`�yp"O2Qh�'C\(��Cl&MT�U"O(9�a(�9;�8���Ou�]�"O
́ Kˀ^z�q�
v�Ĵ� "O�#�1 x�׌]���"Ojqi�D�TZ��X!�ݪ���"O��1�^5=���	B*V$i|6т�"O�5�1�؉���`S(��@UB�"O��zo��A�6Y���k���V"O�9���ڱC�q���L�gir��g"O^�h���	�fD��b��D"O�I2�BQ�b�@��фΎ T�}
"Oʄ�q� ��<\�u�"%@�Z�"O��^�	q&���S'Vx�G�'���7_-h�y3� �8>4T� ��Y�!�d������
�:Q������G�!�!Q���P ʩ\�Q�EFK��!��ף]��B�6e�z�C(ֲQ�!�DN j�ЍAE,]
�l���i�!�XᎸ��R�1k�y!�Y-t\ ���&?:dxZd��> !��U� �Vq�+ߌ未r爌p�!�d�#)�� � ��:�2%�����9/!��,/��Y��K�a��]	D�2H!���Es��V�c�����E*C�!��zqXMô�B�{�X��Ӥ��T!�$@?��v�O�[M����.��$R�}��� �:g�7Ŵ5�� P�Hiʐ�'ў"~�qJL4;�J�J��ӻm��X����y�Ћu�2q ��b���)@�U�y�N��lQH���%P�|��Oƴ�y��
\�؃F�=Qبػ��
�y"�ȣ1Y(�Æ$��H	�@ ��y���N8�T)-_D��$
/�y�l_�WL�=ѥ��ZXb0�e��	�y�`��{�:�)U�ӂCΩ�T�ĥ��7�O����`�&���B'S6e�HZ�"O�I+��H�T�MK���]H�e)&"O2`s��Ɂ-NE�����i��qAP"O�@� ��+3��H�� �n��ps"O �ZŁ׻g�����ݿ`�z�� "Oh◦	�C���4D�;Ix�Y�"O\�34&�:.~$�J��Rd�Bpɥ"O,yChI�:�RM9��Qr��4hW"O�@�䟐��hs وK���hT"O��R;~d�c�IÌ<^X@�p"O=x�(K�X$���ӯX'\�@{�"O�$�*�0j1�@�E ޽i���"Ol"�!�A���R���9�f�z��|��'�x�����,�p���!dZ8��'�����~�F�v��F��	@�'�xQ��oH�����](8�N���'>�����"�z���o͚/"���'� c�+�t���s�&O�c�De��'����En��\���W`��_-��'�ڝ҃�O�"���$����P+O���	���YU�EL>������>�!�R��j���	�`9�����D�!�D�g]؝�s�ˋK)�1K%�B�!���[��(�C�^2���ʲv�!�Ad=�	��e]#:��
��f�!��o��K�A¶-yT j%��;v�!�[���@��V�A��hZ���na�O�=��Z)��'�� wt��n�r�!;0"O~�''�-~��$�\�5Z
JG"O(,9��:=Vj "�@�9V,��"O��1�?A�D@"��8T���"O����IR��1*��ܶg�2գ"O��x���=>z!�d�т5x�3W"OFuBl׽?h��2�2i�(v"O89��B�B��̓+m���"O��
M�N�
U�u��{l�q�G"O�*$�GK���g�B
w`&Dص"Op`��^�+�4�)��-fB��3"O#n	0y6��F�A�2�	�"O����B�b_R��`�����a�'��I�4i~�QnD�+�l��t���7|XB�	���\�lO�.2I��+�( *B�	�L�p*��L� y� �L��C䉀b���Em݂5T$-���rB䉏E��h��Ƀ/��;�+����C�AH��[�	V��cFG�	�C�I e͌�����yA���$"�#aC�k��H�Ȓ=�t2�.��FC�ɊY<.$c4��R��52CgL�u^B�I${YT�yh%S�IrB�+c��[-�.u2��2��T��C�I���ϒ*^���ई�6C�Iw�:0#Pa�N�J!9��"^C䉺v�l�BV��IE��76��B�	�]�ܴIs�.|ۤ�*��'l�B�)� ~�p(ޥU���qR�D)b�ek�"O \[�፨�5�T+	��>Y�0"OyB���b4J�����B��K3"Ot�f(V,<���(��
�����P"O����C�Z�;��ہs%F�xr"O�$ѤʕB�8u�N+i�"O���mI�q��p�'f[�.)F`�@"O�E�S��;Kۖ0Y��+R/�8��"OL�{�Gǡ,=N��������r�"OB����Z�8��/�,����"Op�0&�
�y�j}�/���"O|XEI�C	���`�� �"Oju�3�I"�npi%�
�@�8Du�'�1O֌B'o�K;�=�n�7b�:��B�|r�)`J�i񦅙��R�;cw�C��:�~pR��1G�Š�JЪ+~�C�I�7����E$m��k0�"��C�	YZ�8xb�@�*�Y�h�"�dB��4:�Z �԰Jt{b�P�5+�B�	�C����k�&�8̐��P�~B䉪 mH���B[����eǌ�n)XB�	�Zp�J��o��P�&����VB�I�4�RJ'x��K�+�55�C�	�v\qHS?Q�̋��י2�$C�	�::�r�1������e�C�I!F�sU�/yEn�ɷ�� 9�C��?g��Rd��p�<�SuN���$C�I�\hT��Ũ�`��/A ;��B�I�7��`�#B4��SFd�j�zB�	.,�e����<:¸���.#u3bB�ɯt��ܫt��1m*��z�����"B�ɹ4��%"S�ưl3�艅[-L&,C��#��I�@����C��.b�B�	�*�����M9�ƜB`�Y�O�B䉅5[Nx�u�N�U�<�'��W\�B�	9"�����t[�����@�cI�B�	�0A�%RZ�&"i�RE_	G��B�	�K�&!(�.�c"�D˕��a��C�I�'���14�A�(�����e\���C�I�6� ��]49��}!R%�4aB�I�%98p�B�����@Qf{�C�I�CM�mY����6����Q�c:�C�	�~��$��#E�pu��f��C�ɭ/�@�Ŏ0��c���%��C��46��+��O�Kp���	WJB�	2j���SH�+ ��#��	'B�ɽ5���g�P4 p�0��J�.B�I�#�P50��/�0Dh�DP4#�B�&$rb�s�_�l�R�$��0r� B�1 tr���wE[�-ͬ �$B�ɥ"U�5���	?��Y�#L�L��C�ɇSBV��礕�Ks�$�r�/�C�It�B����	]��z��/;i�C䉿A������T(��dU5f�&B�	7J���1��&;|<�
�g��Yi�C��J�qc�W-m���F��lh4B� [�8������}j���e-Y'u$B�$�ѱ�A�=X�Ț��cddB�	p��0���s��c�
Wb��B�ɜ1 $d�GL�4,�u[r%� QHB䉫d�ɰ,��1�)kWK���$� �[Έ'�Mhg腍i!�ۿf�6X� ��c������>$!����q�=e��)V!3G!�� ���uF�+O�9����e�*���"O��B._	8�%�@��{�ґ9"O乡c�-��۰#R�j���"O�	��ՙd`Δ�$�Q�hu�PC"O���Ӎo� gaV a.�02F*V�y�O�z����fcAX�fH��Q�y���(\`ZI�dH�;�a�I��y��՜;����Wǘ5)8s��9�yBhٻ2�LE$L5/�\�@h���y�Ɓ�*9�@ł(J���^�y�g�E�v�q��\'|�h�&@�yB��h��@��g� 7X}���9�y��3q9�i�qG�% |(��M��y�F�c�6@�AX�ҽI�T��y�Y�,�A�k�u����3�Q(�y�;�Dcԁ�;b�섚��J�y���D&��YeZ�m��a�.ս�y��Q"3h� 䇕n����G���y�O�]��pү�:czl`�'�R��y�b��&�D= �ŗa���Q'�ܻ�y-^Wg�j�'�^���1eٗ�y�ì#wa�4'�U�p��nY��y��9*�V�ئn�Ku�sd�W�y�͚������l��$�H���y��_�da��v�Y;3��#u$C�	 1/�r�]���$"Se�C�I`ծ�yDJ�u�Ʊ�� �KՔC�	�k�\��S��V��%��n�B�C�	.}���J��P�ZR�K7~��B�,N<������]Y֮��z�B�	�.l����S
E��m8N;�B�	�)�܍3͔9P�$4!����B�ɺ���K	������ !#�B䉙,�I�K��H�'ZC��B�-9�b�ZH��ゃ�lC�yQ�b)D����]Kʴ���p!�A��K:D��Qa!Z�h�B��#�ؠ
����9D��R$�3冬�Q��6��a"6D��X�&8F���p� ����)�� D�$��!��M���|��e��� D�0��$�!_�h��-б"\��CA�=D�X;uF��Y��*���[��e
#H=D�l�VŞ�R�2�ǯ%$��i�+!D���R�WQ:��ɔ�I�|�Qa+D�Dw�\=]��a�ȈM�5b��6D���sc�5�3��0K|1с�6D����AN�4Ҽ�  ��h\u���5D�����
�Xز0A�nđ�L4D�����,+Q��w�dc�&�l�!�DţkHv�
ႎ9���o�23�!�Y��ʡ{@��7��(���,]!��2H�n��E��x��8qH��dI!��2}�i�$�9�hT�Y�'D�8��NCq�#�/v�J��7�0D���$N�9@^� �I�V�>�[�./D�DH��
vܤ��Q'TY"y(e-D�Ԃ��^�':�"q���L���?D�`���)����#��(!F�>D���'�Y>Z�q�3���|�n��4#'D�t��P%-��x����`(B*1D��xa)_�Y<��KQ��)f�12��9D�,��!ڋ<�`�� ����K9D�# �/l�H!pъ�0i����Tg1D��#�f��@Ej� ��/(�щ�0D�� &�a�&�3׊�X��8k�L�3"O���gd�OU<	��g@���D"O��P��J�T�b �	i�@� �"O��AQ�U�jnP�q&��5�4]9�"O� [BGC�]��8P�ޤyI��3"O�t���Y� If��
Nd\�c�"O�:t��	&AN�0���CL�y��"O�@��f	�VM­!�L�~� $"O�Rd45BD9��ŤHz���"O�$Ct�$d��ءÇ�A>�Y�"O*pH�eлb䂉{��!�@90#"O���%O��e86�Q�,{��@"Ol�W	&f<t�Q� S$gn�Ӏ"Od��%*�(v�FoE%[�y�"O64��gC#k1ȉ()_����"O{�BS~���H�f$Z�"O:�X4E�m���U%�dN�lA"O<�0�C�35C"D�u�X�AM��Qe"O 8���RV%�Fmi�	���yr$G���0��w���ؒ		��y҆�,�`1c�j�.�т�E��y�ȇ&V\�ފ`�x@BoW:�y���Co`�*�Ɯ�Y�&����Û�yb�˒w��0IĄ�8c�28X�"�y����ȝ��@R�rR�Ywh�2�y��)���c��f���)����y��V1x�n�ӔL�2Y�6i��
�y�"�2,#����׀Xq*�23�y�Ë�!����ȭIl�Lꂫ:�y­U�Z1��qF
�I&�I�k��y2�V�V�<���9��I�0����yҭ̫=p���Ah'~��FS�<���įt��u�,c�2��cSd�<���(Wd�S�d �FLh`K�x�<)��F���e��\�d�p`�|�<���ι�uͲg�5zuN_t�<�wa�;&� �rɑ�Y[v<�'�o�<�G˔�4�UQ4E�����*h�<�n��b¨m�&'�+Gv�[�Go�<!1,ۢqyu�a!���Ne���n�<A��;w�����kܰ`�j��¦�O�<QE��\,���Z�g�e�AL�M�<���έR$�9�d��#���D�S�<�����b�� �le숻�de�<ٵ�UӶm`���c�� �!�Pc�<i�.͡.��
 � n��䊑k�c�<���S�P��\"ٞ�a'��: n'T��`'"O#c��Z4K�`�pK-D�p׬ɛjI���&	�)$��h_�y"$�� ��h��q�Z�3�	��y2 F*q��H�ނ�m�(l���F�yRm";�0�IA�D�N}Hi�a��+�y"�X�u�h��6;A�R�i!hC��y�'�f�@ u����ua���!�y"F��xzy��óUV�����J"�yr�W�c�#��:��<�����y��ؚ��XG	�f��0 ��<�yB�K�7cj����T#�T;�@V��y�-y*T�$Nѝ�JM�5�#�yr t@`P0�%�<}�dH�)�y�-�RB�\I�-MS:�Z���5�y�Y97y�L�� $8& �B����yR*�a���" �3/��U{
M��yz���i�<�n1!B��
_�9��S�? X��֕3=H����M�5�@Ag"Ov-KG�(3���WKW�r��"OJ�&F�p�e�0�^�]���Q�"O���s�e*`����<�(s�'�1O����K���zDK�0�Πh"OFdi#�\t�I@��䆜c�"O�aӥ��KvP��(�ݶQ8"O��0S*.��T�"��{2��`"O��96'Z2�(��a�B�̬<��"O���ʠ.c���@/ɑI�4"O,��iȰPl��R `�%��Y
�"O��'��h?��㡩�3���"O����=A��r%	��l�|��"O�Y�Ģ*S����Az�d|��"O��B����c�<]Õ���E꒥��"O��R�Ұ(O�j���7��!�"ORԲ&F_qd� �#	�$�"O��3���!.�00oÐ
oI�T"O~�{���,:�u�f́k���f"O<���dݛ,r�T0��4iRHa��"O�!�v 
�[����al<��f"O���0
O�@% 8X���}WPU`�"O�\q�Å�R����Itf��"O�l85�
�0e=�φ!U4J�"OD���F�*4쁹���&@ص�"Op��oA�M�1 ��ަB>���g"ON�yq*ׇv�PK!MN A�y"O��P�i�_�j,�1!,4�N�*�"O I��H�=�BH�c�`��%�!"O^}��g�@-B��4�ٶI�=:�"O�mF���f<�DO��xs"O�8YpK�34P���a.�� ØU{�"O��3iB?T��@JAn��1�� �3"O�� C��2\�m�3�Ҍ-zTh�"O=c�T�Rdxi�&�9�p�`�"O8���%"J�`����"OҠ"Q��<�H���g�/7��p�"O��+PS�2�Y�iUl�A�R"Oj�±���n+pXB7�Ç �~�"O ��([y�҅hö^Ţ��"O�h`@��i�hd��2��(a"O�jF�G���1�f��b�N�2�"O���R�B�H�K�3^�t=b�"O��3�(� ZW����5!�BxR�"Oڍ!Ó�tX��ǘ4"O@@�cZ}*%q摉O�$	1�"OTDI0��IW�]���n��l(g"O��� �~A�d���f��X1�"O,�8WHU$H�(9�/=�Ru f"O�<���Y�{.$0G�ͺ��u"O������b%R�[ ��		B"O^���Ԭ|��F#%� �w"On����\�.���Iae_�݌d��"O�I{@�Y�h���Ú�AԖT��"O�1��;]�.�b���5T�pɀ�"O��s�C�m�إ)��g�h� "O؅Y#�F3:D2�Ǧk���"O@i�ߢyo�T��E�C�쨳�"O��8!���0��J'@z���"O
, `���p�P�D\1A#D��v"ORQ�BI &i� �dcJ8i:�M(�"O�
$2D�=�L\�3II�Nb!��)/z1�N6<q��I0�K=uG!�d�9�4C�լSR�YS�E�m>!�� �Z���5�a�sM��NN򴚓"O��2���-F���UY�)�\�"O:�2$�LL� Y�(�8cpV�@�"Opu2�@W7���ڡ�O'r�,�"O�.}�.E�.A=;��h�$ݜ�y�M��+�Dاm�7E&E�Ć��yb�ގ,,A¡�˚B5�aN��y���<~�\�$����s�ƅ�yr	ȫt%�"��MZ�p�j����y�P�!dȰ �κU� �q���yBL=v��U��U)���.���y��]�@�b�K�`�k�c5�yB ˂t�P���y�U�o3�y���E�8���ːz���`����y��7Z�jU8�\n|�P� 1�y�I��m�V�b�lG<e�a놀	�y�9��ܺR��Y�����H��yN�0�P��̈z5�T)!��>�y�*ĊhJH1G�;'�@�e�I;�y���(e{P�)'S�/j�"�Mʰ�y"&��ߠ �u�L"���;�m^��y⏙�t��a'n�%��o���y&�����Q:	F�):b����y�*Ӯ=�\H�lؓ{� ۢ%[�y��7
g�� "ɂ-\�%�	�'���[C��C	�-b��")3\�i�'9�M3
��s��8��� ��S�'�5�o��E5�ܫud�	�le�	�'��
PN׎�$y�!� Y�v���'�l�ϛ{a
����+V2 �'+f̐E&��=��iY��ӘSԤ�q
�'~$�)&�"^�;T�I�6���'�8|j%
T��Dg�9�����'s��R��п@\��he@�+��+
�'"u8uDƽ��1��N�ӆMX	�'�8�3T.�$S��1V����'B�I��ƛV)C�턉,�N		�'Lԕ��	�V����R�ޮm48,�'�ȩ�sd\�H��2b�k�z�Z�'i9���D���rN_78#�%B�'_͊ׄ�y �Q��U�0E�!;�'H����M�H���2���/���'���s�ف_�N1*gC&�� �
�'��\�էQ/4:4pX$$��"9�R
�'���7�$.34�H��e�h�X	�'#|Hhu@ƠR�@+�1*��m��'�&q��0E�BأF��qnT �'$`Y��)�x�YF��)�
�'��欂0#򱘶��3x���'��@��31�a�%L��Z�
�'2��5��[�j�8���;�h�p
�'�N��fM,Ӻ��fl�y��'H�"@�IW|  �ݒ(���'y�i�vfC��+��Y(X��:D����  _��J#Ώ�o�r��8D�pp��"Iq��R�c�6��x�`,D�l�"kܩc�R�ؠ���zWv9s7i*D�T�
K�5�f�X�� ���'D��K�"���\�!h�*
��1�-#D���AG�w���h�v�R�Z�"D�ȀW�A:|��a!w&!x��s��-D��H'	4Q*����
$OX��x��*D�ܐ�L���<I����U���3D�4s)L�nx� �@Ɓ-G@Mڷ(3D�� P ��d�~�Y��*4���cU"Od���U?BuP4`�@�/t����6"O�|␮X�U�l�1���$�*�"O�%"�+ɉ���iCK�+K�ZѐE"O�a���")f<8��*������"O2\!���b�j���ճB�"�0�"O(T��MQ3ԥ�d�V�vz!jc"O�Q;���Yo���#"3�01�R"O���(�d����E���3�ސ �"O���G4#�\��CN?5�r���"O�X"�'�$��	��B$B�
�R!"O�t��ϐS�%�����#BHB�"O��㛨���u�	��)��"O�|�C)K$:����&M?Q��Q�"OJ\b gϸ8�X\��N��X,�y�B1��,�F�F�p^�X�!&��y��]*Rz�9����<E ��p ���y*l7��� �/>굨����y�K!S�`����,/�u"R��y� Q����6�@���e'�yB�[�(�+�W��=�1��y��F�=c^��`��	��A�����y�O��n��	9��l�N<�@��$�yd�	bb轋��c�ir *�yr#�8�.y*޸R21yc/͉	!�D-%w��ENڡ�j��(*!�Ĉ�tx�%��"^�\	-��!�D3$+�e����2�����}�!�Ď 4t��*7�N�^=���ug!�DK�A� �9�h�ٔ� F�U)P!��<	����QbF%a�G�k!�Ý5dRr�$`f�*��UX`!�$ʞj悥�V@��}9���6K�8Q!򤏚�|���-ŐYq�$V$9!򤛽9���05�	5-�<��&�A10!��2%(�2���UG(�K��� !�$��t���Q�5	'He��%�q!�<��(� ��b
��P3EI�*!�$�����_xM0Ĉ�F�!�ա/�p,	6�:yV�� "G�!��XBFI`T�	%��B�@�7�!��o��5B� ��fۤ��6�!��˛T���0`˦7�T��FA�8�!��f�j�1���	���"o�e�!�d �>��91�^(6�޼���^�!�䍒a�<��'\�):|�����(%!�DF�&��|���@=5 �e�t/��0!���9:4��{e��'s*`3ɫ.��_��(�ʔ�D�[<+��9�'�>~S���q"O�Ca���y���d��0<�|@"OP#o�5,��zZȕbJ30k!򄗣6�ԓf��C]�s� ��@Y��~�����Æ&
�>%�	��B1d�� �r"Or��@��#֊𥢃P@`�PR"O���g�S@D4���<���"O$�0�J
�0= N�:;#ԠBu"O@���-O�u0&�
�I��ѫ&�II�O����$�:*Hɸ�Ᏹt� XB�'f4�!�����Ȁ&��=F}��Ob�=E�DO��0y�(��KŢ}8N�*DM��0<1���M�#�>�2�A%zH>5V���=(�e~"�i�ў��Ϊ�r2��V�%���щ;�(��hO�~~� �5zr�c�� h�mChC��?	�A'�S�O��q��"�%�$@Y��Y�j��"O� �1yk��>V���CO��ќ>aÓ��ɇEmd�`�RZ��1�.���J���ɱ"}�?��#O5G���U��D��r�"��hO��W�И�f��Cv � �`
���ay�Z��?c��@�/��m��ZE��s�&ђ�`84�<��Q��N,rӄ�82Jx�c@�0��$�S�O����V*$���P`��nrlp�7��OLdJ�����YK�/�J{��	��'��ĈФ�{Q��=L�0�e��=,�!���"s�����N�2�嚛'!���*Y̚"O��Cv�X�	!򤔑7Qx��Ó5� T�!�R -!��J��� ��f�2��֕1�!�d�x*P�b,
wBlQ�c��6��';ў�>y�3���"����#�F���N6D��'.�>�<(�H�j$(P�`j�>A����dT��Q���!�"�!��2v#<�z``5D�X�s��`�*,����Y�I��/�%�S��v��Օx\
��q͋�|)vu�ȓ�ZEҖ����b��J�Y�.��ȓ�8����V��cĞ�MK��ȓ"@Z]qV�N ���H���8��Ot���͔k��m`��֦.�cS�Њ@!��+��,�P="�@yt�!B�!�D��	�\�+F�Q�T ��,�X�!�M�Z�:i�5�ҍ8�Ly����
"�!�̐v]�0B�(w}�`B�
�a!�X�bl�xc��]�>o�cjEW!�$��G��Y�abJ8 u 9�(	�vT�d"�O��סB�^vP�R��C�����'��'�p�cB�\wWQ�cE1��Ex�'����#�/Y�v(r��={�� ��'D0}y���{�ʜ`D ��)���
�'L �S#��YU|m���[u�AY��������d؍.���A�V�;�6=Z"�CFQ!��(�^���!57帬�mB.3�!�L�-7,9���,�<t�l��an!���O�i�g�"������	f�x�7"O,��%���G:��0�	�lG��"OL�bĔwt ���[�v<���'8�'�F͉����C{�q�SA�b�ء��'
:P����K�@��:����y��)�5C��\б�7>�ukt��c~�C�I�`�ɻw�/G
�(��Q�gP�"<�ϓ7������s$>�Y. �=��������"�K�a�\�@�X�	[�HE~b��8R����Ms��(饊O(?1t�� ���'ْh"�q�4�-��$����hO�>�*!�;O�L�x睐'6�DX��=D��.�3�V� ��'6�PS@):D��a�M���FЀ�! n��Q@�O��d5�)§�y�.��i�>ȉf��d&�0n��xB�'T^ �	?\�UA�fZ89�ı�4���>���T?��J�sӾ@b�T8wd�*ab"D�HY�@Ӵ8ݾD�����	(��StM~��=E��4+�T���)i�N0��:8���ȓN�={rT�6���I7�S���0�ȓp(���V�:1c���Y���l�Z���O���& u� {&�6�^��U!O,�B�+ߖ�*1m^<V$�A,T�k��B�ɵ`�@%�2T���{ �ռ}U�B䉠{�鰠e��*pm���?pB�	Z�B�@)�$�f o�PB�IB�������'A2��FџwE
B�)� ��"��$&ݠ��s�ݝ,]�Đ "O,8���t�d��$f^�CU ¶"Oي�c̗|���`Ǐ�0Q��ؓ"Od�2,����U1�ޖT� �1"O�E�͈#��A�S��\M��%"O4��&����b��4�F�+��@'"O��� ��v��t��Beιy�"O0�$��ic�%��kX(n]�X�"O���c�w
R�	!�>2��2�"OĬ �&��P��yP
�,8�i�C�'�ў"~r�%Ҷ$B�zs7N���kסO>�y2�'+f���DI&*ұ�G�/�?���M��A��d	O����س@I|i�ȓE��EIdG�n]D$3� �/���ȓR(��K�k�"U�$ "�ԅ�� 9��&ֳ"��	cs�
e�4e�ȓ{�8�"׎U<Gr���c�cG���ȓE��H��V(�V�p� �E�ꈅ�����O�B�Hs*��1"ȼ#��Z�J!�d�)�5B�"H�:�@�c!�ҿ
]!��]��PiQ"�fr�`cD�ʚ�!�ĎL�e���=0�` cX��ay�I7c�:�"GO=/�����Ů'��B�I�`
�ɻ�pX��x��31uz�h��(�S�ӑc̄H��^�`F��B?juPC�I�4̆,��ĠH���#H��|�C��4�p��L�p��\+7왥O=8����<�$I�Q9�'Jh�ْ�L�<����>N�>��U�Ԍ .��ׁ�m�<�@ܝG�Ȥ��jG�&��A��Z�<!�@*o�(����w2~���w�<)ѭ�/��L{�(�GCj�8ԩ�G�<y�N��2�:�Sa�\��h�3I�Z�<I��i��,�Bkΐ��`��kA}�<��F����#AM�[���'�^�<)��!�)���=��ً��NW�<��H�<Ad�S��K�{��mS�+
z�<�f=6���j�cB�/��h�$��w~R�'�F��Ù))F�r�b�)T��9����ɝy]$�B�֥6'I���O�#��B�#�U ���s�Dk#�?75x���U0GE�?��5������=x�0T�2D��yo��"��1��18~,d�`��M��)�S�O�$��ǿ#��h�
�Hr$"O�Q��1F��	j���9��Q�"O��1C�"%7��� h	5Ԑh1"O� �n�2!&ݫ���j�h"ODEs�
�������%0�Z�x%"Ob��GF٭X�lDY6'BM�Pd��"One�D�A�@:��'�	���I�"O<�"ĪOU$u��(Ό	���T"O�c4�C�00�b��$L"�c�"O� s�IH(HH �HL�hn��U"Oi����<W/�H��gD�i��§"O� ���!8DLhp�[;3a�x�"O*i�b 	��,!$+��}��"Ov=�C��D��Q(aё7G��i"O��r��D>;/�%�Tͅ$b>��x�"O
}��Ж9����tkH�n&��PB"O��P*�0X�Fi�p������^�!�DØ���$�
�_��e��+J��!�$�؍s��N�s�R!�Jٳ:!���[�.��Q����-��C
!�$��cBh�r���a�[+_!�� �L����w�h��#,�����"On��ȼ��l
��7PcP��"O�(A7
	���IO*4���"Obq1PbҪ?9<�@�S;ND�a�"O����
Z�½V$L�ҡ���yi�"m�\I��"Q�f,�af ��y�+�w7�h�GD L��8f�_��ybGQxG �����4CH�ݸ�l��y�Ǔ�D���RH	)sV�����T	�y�a�FGf�"4""��ɰ���y�	\,]�]�0>@���y��.7��ԋs��lj�G��y��/Рej -S	K�p�6�yrjU<w�|"�f�:*�5� DN1�y�gC&}K���k�})���5�y")I&u�(āǱ_#��a X��y��J�2�9� �֮ uV���%J��y���4? 8k�#/7Pp�V%�y���tܘ�`�	��P�FL[��y�-A�>1:�X�J�0��d�v��y�#G�+GZ�"�0 �,�F.Q��yB���=�HL!��\75�!{e�L��yR��%@��Kf��|!�q+�>�yb/�7m�tU"◇t�@�T��9�y�ťe���u�@�u�Z]"u�U �y��҃Jj��� �a��2���yR��sg*`�Qdx�]��ʃ�y2g	��	�'al���[��yr�Q�G�$��c̆[z�pPC���y��\�C��-yb`U^;�zo�m��')�)�vL�� @��!U*���'�D $�*z� �[����pA��'��k M����8B$�G4�p�'��b��M#�H@����M�yC	�'M�1��厩�N�s(Q%G�z5y�'tܰ��nu�� e�2r`aB
�'�ص�ƒ-�P�P�$��-�����'B��s���E$�8#b⛙!^���'.yڡ���oY������s	����'�9�FaY�:{�)!to��tl��Q�'��t	�hE*I��4�9c�P�'G�!�7$H�4hD-�K��P���
�'�t)�v"�6	��q���ŨT�����'G�Uq�P�%H�r��Ұ 4�
	�'�����D��}�Τ�TA�Y6�pH�'���jSA�8a�R%����$`u�U��'*\�V�S!e��Ę�+7jŸ�(�'jA2UV�`
Z!+��]�;����'�D��k�}0	��l�" `��	�'����1fN?r<�� £*	�'�r-Hac�	J|b!���:N:u��'�n����?$L�P��3�v���'�<��EI�B�`�[�z�`���'�^Tc�i·N{ར�k�M��d��'��ZE엒Z�4Z3��+'R�R�'�H��`b�7�y���I���(	�'�VEp���=z�aaӇ۳a\ri	�'�9I��X4r`�����d��x �'٠9h��Q	+�֨Jr��$gu���
�'U�dg��O�
��A-TX�@a�	�'��1�Q��=�
�q��%Wd.e��'�m�"M�2zgj�sT̍�M	B���'�J��!X�?��� '�'i�$���'������Z��*�dH$p�b1���� �-����$U��M05�ޚ8��r"O<�da�m�nኲ���D۞�H�"OVX�`��z@�I"ċ���F��B"O�l�kW�9ֽ��J��j���{�"O�=��� (��d�$H���D{�"OV-K!AW�]�(��GH�)V��7"Od�BG(�-W�%� ��-+���"OTc�+Қ/��訧&I3F,4-X!"OP�z5���i�UA/��E��"g"Oȁ��̠*N���ư$$�W���y�����I�E'�W���j����y2
��(MI�X�Q���3ʚ �yb�M%o{d�"a�8p�`&;�yb�U!u��|�2�C�a��a2�[6�y��X�lP�y ��	A������yď"y����`IJZhx�#K��yb�@1H�h(�`��V9 ��B,�0�yb��<6���'e�,�<ģ�枤�y&ۉ}LM��ǈ�	��
@��;�y�iF-=Θ�
6�SY���Gχ�y�M�5G�i����L�Z岧-\��y�,TP�0�1����XI'�@2�ybD�6UA�a��R�t(�l�!I5�yR�F�flI��uy��Y�a���y�J
�7	��GF��xs�(�<�y�M��|�:Up�����,��"��y�DSTڼ�"���C���h�	��y�f\�tJ���NU�O�������yG�#<�\u8��?��T���8��'@��r�9�\�O#
��C	I�&���qC$R�^9
	 �'��ᚗ��RF�V�(U<\�egL�{��Br��Qyb�������$s$�0�%ַD(J�၁,�B�ɤdD^�@k��K+����M8,	^�Y$��7�ze�Ģܾ[sڀ�鉠t��y*Cf��Xf���%�	���$��[n�W��oFH�w�],w�Tc7��� �as�"�5��)#bO�,L$<�V$����+ue0T@�@�B3kDB�W[�1ń�A�.(�d�]�kp���3�T�_��p�U�T�R�鉯ft2т��y���2D�"�9ʐ}����S8�	��E�+fi��L�'dP��L� ��"�.n���#�̾�v�zc�5�$L>�x�B �����fA�7��
���%)��r]f�Y�gS})���m��Z��Hw�ƚ԰<�pG_!u����d@S�d�ha*%}�rי>��T ��	]' �������U�$e�O�|�t��Qh��Zpl�Ӳl*P������}�pX3�]<���$�ڎ>�V�q��޴2�����ᎨK����#�E�D��QG����T�(��2n��T�`B
��0<�W` gc�A;��ÄP�ɭ]Q$����@,]�5��D��t��U��:��*PeY��M�֯��?Mp'��X�3?q�HL�&��hf́ �䍁U/�fy���2 `���W�	��(�O`��-�Y�6lΧ.fVi�sC+*�^D�J�}>�$�r&�<5���"(������'	�3w��9LE���TZ��V�4 A?pC��I'X�D�@Wjߣ�3��O8ŲbG�Q�18�ܻc�Θs�X*&��3rg��U%����u��aa/޼����.�mn2a*�����ˑ�j���֡���/�=�蹖.:�D�>z���c��a�t�%�0Dn~P����!���p�ֵ<����yO�0�@��?��p(7jJ�HmT��� �q8���p�����K���3dH(���#�삾v��m�'�n���Ͱ�н2��O�e#<zl�}�WN�8/��"����t(�馁��
.�y2f����H+ĵj;���!ŁgR�Ԧ��b
��+C� �N��ڏC.6X����(�Dk�'H2(��[�A�PX�'��<�4+\�%hr���+w��P��B?3
�1b&�:��jU;ci�pXAh���4i�K�~BK>�D
�(��$��$� ��2OP<����^���=C�4�w-�S�V��A�	�Ny:��Đ}�0h��D�.���'���<�7��;O��25�X2b!�b,�@�DL�e�F  �O�0��+Ԛf�`��I�i��v�:=��fN�E���#�/U��C��4p4|`��J��
�C�����8	"��F0_&���·�/e�Q����KCg�H`၉,�e�Ê��yBG�>&v�P��E�h�Ĝ���Y	?x��g��{Z�)̨[������|
� By��.� mI���I6��:�O@u0���[jV�����!������Ӟj[а��	 �Rߨ|�>���$J�v���$4.��a��<^ax�C�'��Q��mJBr��ɲ��%m,�qs�D�3$qS�ړ?3!	�O�Q���ޛ`�Μs�gK9uo:��ѐ>)�@��q��P�U�@=��[#,>�'Z<��Ɣ8J�4�ѵ��ijA�<�si,)�p]���4&�h�6=����2ɗ�)Y��A� ��4�||�}&�L9��ۊP�pAO�X�� c;$���f��HԨxx�,O�<Śy��҆fRT��$mJ$�� �̉Q��Ģ���}`j"�S� �NzӢ;,O����&
D� �F��[�v�KgⅠA=҈���#?�<c�mXl�<�T�ӡ���Y#�4�0A@-�h�I�4�6M`V�)M_*5z ��^�O�����/0N��KU�8x�Nr�'�>�@p	�!x�������v�~����Î��)��
ɮ�~�\~����3vb�w*ȝ>��Q��"
!��T��d��̛9�Ҙ1�P����&Zɨ�+pnL�Q�azBOW0�"d�@a�q:�8�����p>q�`�)Yw���EG̲V��R���}+1��%c�'9�M�W`Z<i�F�yT��+�������81�e�נ�k�B��}b�,�G�p����t�� u�^�<�2ϟ�qgZ� 1�ŕhÜ�U�
.��=(F�T@�f��P?E��"F�2;,i"���R��0�ȓ*�%(�&�i�8��U�5$zj��'XX��i�w����'O�;�M'T�F�rH�i.�����'/�����ݳ5�J$���LE24�[���:3赚dᅃ�!�d@�HI�A�D�Q���];���Q�,���L��C���I���']����`��#�!�p<�xQ��ͅS��$��	����3��e�!hAA�O�>�b¢YBݒ,B�}o2�2e(D� Z�i�C���aZ.�ҥc�*"}�C�X6����D�,�bR9|���p��7�y��K$�Ox�:�@�	J!���$:��My�*ˉG|V�y2�ğC!���#[�(�1m�a*�	��zG���Ȓ�	4r$�m�}�cC�3��Tp��ԟ��Q���Y�<�ÄF%ѦA��Cܙ ���iJZymNpe��=E��n��}-��F�C��M�c�.�y���{�X��	Q�sm�p+3'�y�mq*�q�'��B�������yr�F1c'�E
rHY6���d�y��ׅYF�8��r�HM	g�݀�y�����y��hM�s�r�C���?�ycM�R�P`�-Ȋu� ����yr���\�h��@��lG$d��.�y�e�$Sfҙ3��Y&0�Ѫ�y��!��c�6T�<��i��y��>9��@k֭eP�T
�)��y�lS�q��TrG �DŸ�M��y���%=�"@����z�pؑ��yR��c@H؃HM.o��l��㘧�yB���t�	����Z��)�3���yB��N�9�1ɓ�,H��q����y�;�IA���]Ya��y"* ����)�"�$��}��lV��yB���	L�2���?F]0s���y�M@* \N,��J�vX��2�Χ�y�A��`�Z�-vzAx����y����h� H��^}X*�x�g�'�y��K�<�|A�S)��Y�}"@�Z��ybJ[5@����\
m�:ĩ֎�y�
0u������?�4)@gFT+�y2bMM�p �b���<@�<�6L���yB�5��Y�nO2��t�fӡ�y�)�WE�Cs�G�6�*%a1��y2���B��򮕁)|�� �_�y
� ���6�ٝs�
�C���
a����"O�yщ�%Eo�)�q�
�T�$ٲ�"O�Um�O7���g��6�`t"Ofl��eٰ@{*E�P�d��В�"O(� � E��ҡ�D��]`�"Od8x�n��"F0�@V�H�`�I�"O@��T�˱x�.��kD��>q�T"O(Uc��0�V3G�X�z�Ū "O�L�����3�\ �/�-?��i�""OPl�"U�z���)PiB�[�"OB=�ʃ,���i�FBE�ܚ2"OHL�BY�4(�!҅`8mHY�"O�����O�Mj��9�o��J�[C"OBT�ªg"n�A�u�q�"O��"��M�:����U��0P�І"Op�ʕL ���u�3�S�a�d��"OJ��5������(�MM���s"O0��)��fh"�R�����P	�"O�y�g	T8fW�0�V�2)��T��"O�����7����X�*Q�"OHљ��7*X���)@* i��;�"OFT0Ce���(7�? X��#"O�P �'
6�Đg��#At��d"O��#��'hJv�� �2<֙��"O�l�qC10�|��F�D-�9��"O�u��jQ�1���b��Cׂ6D���$I�2���9��[<Ĥ��a0D�8SM�/L)qGo�%pa�`�Cn D�ؐ���.�@X��%�3B��s%� D��Z cÓEH�e�`B�$ZBw�?D���n\�y�d�Y�&�;�|�vF/D���'�U�@t�+�K^�o78T3t'.D����fO�����u�^#}�����N+D��Zq��1���D�Q���	Ad$D�������Y��9� �#��Z��'D���GED�(i�q#Vm��0� D��(r��l�R9��Z�
9�1�>D�L�"_�t��	{��C� � \��:D�`b �	�w5�<����#j���9D���/X��xgdI�k��-J�O#D��A�GɃB5fY����,t
b%D����ڨ.g��3T
��B��-@>D��9%M������g�$_���*D�d6��ZO�q(�̇�<��!q��&D��� �J����=+3����'D��sD�� �>I��2	���S��%D��to�!d�)�#IѧyEΩ��'D���f掣f�Ё��mE�/y���%8D����&�#C\�
�,�
>��5C�( D�|�ԿrϤ���G�r���% D�@��E��n��Y[�#�1G˲����$D�\����d܎@ '��㐼pWM?D���#	 >�&9pDl	�$V����?D���I@m;�5p��� � c5�?D��H��Υ��m a��7�$�@�<D��B�֒]��hi�䔒q�4T��6D���B�$F����ӟ_Z:��@$&D���Ṕ	B|�A�ʹ`��=���'D��j�ώ�KP"��a��鲡�Ʃ7D��J���/v��&`ϵq؞��'o?D��R ��e���@�fM�5HY��?D�l�V�Ȟ���2Z1%�%�T�Կ�y��ס�xh24�F�rj��ƒ�y���Q��ɺ�A.�Qh�a�%�y
� ����$4�(�2�H	�|�&"OrL��c��J�\p�wA��	��hau"O���G�eg�PF@S������"O,����%7�����ǳ[p5*�"O$T��g��gvh\�1恦a�5CQ"O�P�a�<���	4o�4Ie�\2V"O��s��n�`�؆H|�q�"O�}�p��.�-;qLW+b����"O�]�� +Ai��`D+�b��"O1wAؓK,D��`�=5VЙʅ"O�}��i�$MF�X�BQ�6$S"O�հ$Ȅ Y��q��׵%^��Q7"O�m�����Vp���0[�t�"O4}+ǒv�ڰ��Ȧ	|H�A�"O�Dn8$!�L-3�`��Q"O�"d�:9��"J��L����V"O ��Q/_Ib� ���QdZѕ"O��ӷJ̧30ї"߀9881{�"O��t!��Zi�4`I�S%�DK�"O5+��sYb���M[!H+�9Y�"O���_�61�tL->���"O��¬�)| �upw�W�T��ʦ"O�����,G�)�c�B&"��
�"O���pX�j����K �1�"O��I�@Ǎ �=C�L�%�+�"O�h[���	*ʂq*����f�a�"OJ��7KA%C_��C ϋx�Q�"O��p��.m��(g� �GB��Z�"O�A�lFy�&���W(=4"��Q"O"��g.~�F�!�� j��"O�Y�g�%%*�qr��0V�as"O�����X����6
0 X�Pu"O�=�c��}(�8�@	�1}�������xrB�c��A�����`K'�E�P^�ҡ��$�<�"c"O����,�l��|27N^t�����ڈI�����Ϩ<Y�n�v����I��H�x1�O6
�>��*��:š�DN`$l�7�ҳnR�*���"R`:��d�~$!�F�#^���O|��� U��08����B�_�yr1<���Y[ ���7��<�А�@ Q
J{�����O�xC�I&Do5��`
��T�I�dJԦгK��D)JO8���O@�Bg!������O�4H��J�4��
ㄒ�2착�M@�Y�ҙ��DFR�t��I�V��"��D�zDA����� �f���(7e�y�g��I�A'��R�B�oH�(����')��'I�<��"&*��D�T�	]&e���K('=�C�䄾%�r��E�S�"��;QMD���	�&b��f��}	���@�;�BY:����+t &��O��M�"$"p#%NA�S���I�̝%H�����jҫ��)m��Q��'�(I�v�S�Y��Y�Ƣ�>)ɘr��k`(�u._�h.�E�âQ*0�Ղ��)�w�&\1�δ��/,M	��'*�0�چPK`�(0)�>��B��_#� Y�Z:7k-(���K(���U��:��NMڦ�Y�)0�g~�H&~C*�b�/S�t�ҝ�4J����>�僚�v�^y����Q�O��L� `��l�4,&� �|�����*L R�ۦ�C#b���׊+,O6P�/�l�X�-]�6ݤ �r-�1�����o���E���g?ɂ�
6O���u�W7����$��BȒ��.۰?�5P�4"�	$��O|�10�P�CR� �ScG0���7���bE8�{��z|�I���t��1Hum_GV2�E2�M�[s��+����c�'TP�$�
G� �!�%CO,����p��p��`YfQ���ǭz�L��'9�yɅ-!���#��O��-�t���j����F�y�6 ��'�|�bCC5<C�a����~�0��b�7}���$I����{"��%I�h���J>X@9�C��?dL�Jw伛FO�ςJ�=!L�g�Kipꤳfo1�O��U��+~����w� .�@�c��'�X�S�l���'@pMi!"¤r3�AQ� 1�l1��'��p�cP-q
Vղ��,/���)N���E��8X_qO�� ��2�9�}!v��+Z$ ��"O�)�f��(PO����Y�l�"Њ�"O�dC���.(CO�n��P��"O�{��Y1:=��
��Z"R�ta�"O ���P���2E���h��"O��Q�B�I&H}G��`��m�w�<��:����@��5(
QC�J��<9�����s�)��Q��Z1@�A�<y�k��Kl���Y?0@Ấ��E�<ydβ�x ���M a�0U*$��h�<'��{	���U&ߜDl�������ڹ[dqO?8��\Qw(L��i`�@�q��{�<�FȒh����r&T
�D3�C�u}�L�1��@��'�T���/��UB�S5��|A�M��R�	G��',1`�J16�B-�*&/�l��6D������W�|��`�JYjlC@1�e�.Z֠�R���!Y3��)D�.�f��d�
4��B��c�T�	���h	~�A�D�� 4!V�řF���Ơ'}���'�J�y�UJ�d2�x�B�r�'"�
���w���SM�%t�(\{�'��eΞmE$���IKeRȠ�B��D���*�pjL��T+WؙQ5'�)��s�m@R���q�z��Y ��?$���6/�Z�t s�B	�!c�隠1ʓ��ۖo�Y�~0c��	B������$X��S��!�$ӭ*�@�C��)D�IB��%=`2ٺb��=��j0��%����O �����#�J�4�Ë[�tQA"O��ô�<0�
ٸw.��d2TU���h��p���3擠�0<�2-���xB�	4(Gf@�GE�yx�D�g�8-�:�!�jNO�M�����l����3G�쬅��`.��WA�,O�9�c�ӇP���F}¢�xJ����Çi|xR2��18�ha4b�=;�4%��G*H��7O�?Oޠ��E�u8>E��xGJ�2��?*ҧh��l��U%K<t䂡#C"y�@��"O��$��@Y�"�B�9"���F�>a��vNdc�,O�	i�CV�,�px�GĸO���Pu�'9PI�VDY�"ᢆ4_8&Y���6?=���n�P<!�%+u��U)�F���1�Im�'�L�C�կK q�����g�����o��Pҗ"O@ĻРK�^">�+t��)���Z����P�wqOQ>i
�!�$��$�A��k�T�؄�3D�Ě"�,M��d�kİi>X+.D�l�B�	�;�x�H$�-`�:D�肶��d��=�'%�0�ujf�-D���C�Uo�S�e�<]hF�Bg�-D��D�O0:�i'D���rK)D�����8hWpxه�M6�����)%D���0-�R���5*��9!�i�r�?D��r�B��lE��Q�';�Q!�n'D�phv��R��e�e�=3tIh�M%D����ŬQ� ��$�["IV]Hw.D�����Y���X��-�JZtp��
-D���$.��(T�K�iv6�; )D����]RlV��
�1�蝈t�%D��8���E0́�FoIf��}�� D��9��Q�yk�d�e�H2l�y���;D��"ƃT�)�0|A`�8[��C��6D��`�FL�1���XAg�8X���"�7D��ZE �S�~�.$�)P�!g�B��ib��rÚ��$�XP*�-LC�I��dC�&Y��A+v�˱Y�$C�ɡ\��	򊉦k����t�ڳl��C�I�Xed`˧/�.	�ܘ���/�B�	_�F��5X���e$��sNC�I��r�Sq�4]��XAlN	L�C�)� �����'Ƚ�!�ը���"OŒW�ӭ7F���A�aB�($"O$�����	��<r�̆'k���f"O�<� ��
b�d$��#Ź@��@�"O愫E�ݤ!oq��!F��"O��R��
<.DA��U*q� 	�"O� �@��T8e$�F=4�$�C"O�mك�\�D���`�T�D�jq"On��D�p2<m:C'ßv�6�("O��	�K�F��(������@�"O LH�Ѱ|�[��P�I~�a�"ODŇ�����K�)`���"O�@����+��	�Æ�no��F"OX!W�Ɲe��ED$l��+"O���� �%s�D٣��J�l`�"O0(²I�o¨�r��ͱ)0�|�U"OށQ�GE���$�	̜f5l�q�"OR� E�O�~��(����3I$<9� "O@01v�æjF*,D�[K㖠�"O���VL���@�"��#�D��"O�l,IFR|܋���x|"���"O����Ίb� ����A% x	"O���MR��B���.�"��d"O��X6�T�.Xpxӭ�i����D"O �����r�B�V��n��eq�"O0l(��*^,
�	��b���`�"OkEIʩq�z�H����p'"O����㐚?����M�,���R"O`E��-�i�vpXק��Q���r"Ox�ӱ���*Bt���\eF�: "O�`�[A��)ã�`n��8�"Ola
��Bj�ȥC"�ųr��Y9"O����H�+Tx�"������'>Q���H��|����V
��`qg:n�F�0�Wk�v�O-��ӯCm��u��5�*���يO���2��
�YF��L�]�Txz�\>�E�'�1`G@��n[36�@Yzâ��q���)�1k�+�%7-��ç5\��C#o�`�׋��\����y�
 ��M8^��
T� ��A��X�|i9�O��
hR��[�J��Y���s����q�O��.�'a����cD(�HhydkA�P�����>�B�!���<5jA_>��P��$1�j�J1*��XY�\رĚdLӏ6?��C�u>��ՏŗAP���c.E8QV����Y�Z�O���"4�����ǋ&H�y0� @�>���hV�|�  >���`F�OeN������"Z�eI�`��vҸ��-O�l��A�ؓOQ>��T�*"nR�{v� 5F�ő#)�Oj�*�U<g
�IQ>ͭ��h��e�O�F�䒿JŎ`+�f]'\G�p��IT]?!f$�4�8���^�V �c�ٹF��M�r/޷$�8�'���&�jӼ!y�'pwn!J�/��*����-B�Z�h���.��?`��A�FK�<%?7�F��MKT���2Z�1R��E�Q�4��Gp�����-��b��覵��iGa�dA�rv~�R�IK�\��D�"�vu wǇ��M�Kp�8��%���S �VT�6#M�_	P݁���J'L�	�Le�d�A�A*;��<JA��I>}s�P�Qt���w�S�-��a)~�� ��3^��u"��#.���S�&����(�6w
6e�փi�qcb��j��m{�@��Mk� Mt>�z�iV}����-��_^ :�F[/W�d����|Ӵ�Z��D��l�� h�� �0�dջ��AG슽	P�vӆ�A�,z6T= �q>�$�wlչPKB�Ef�thdx���M#:hM�I�"ʕa�	O�x��V�^)s~<03�Z/\T��$�G���>!�N-0JFHό�1���
m�<I�C�Kut��Ec�)q~]3CnD�<�"I�:T�����j��ఎ&T���I]�Eb�e�2l��
vC�*z!򄜇}��0@��	�A���c�4c~!��՞tV��@E��\�'-��>m!�$^?p�U�0,K�f=�#l�h!��}�<�2C�G�f�����k��
�!�� ��eH�X-p��E�3 ���h�"OZ��r��!]�i���}t�(2"O�]�vDˤ
�@�`�IIt�<�#"O4�ۣ$�BN��G�2vl��ɵ"O:�" ��w�u��ǚ%XW\���"OX�r֨�Wo.$����+E(�
p"O
���*аߚ���	H<@^~	��"O^@���;�i� ���t"O8(rd�)�&�Q�,m8����"OP��!�T��Aә!x|�"O���CL�(��-SfN��(�E"O�${�B�'t��h���!-����7"O��QS)�J�T�G,�:$�W"O2����M�"/B��%��"�ĩ�'"O��+Ubbx20�ש w��@�"Ob�a��>x���{A�:my���"OX�u��>%�XP&�!el$�2"O�Ph'�1�p4C2���Y��CV"O�-��E�F��j�Μ �Q�G"O�,p0�D�2@pբ�+��B"O��t�NGF^�v��r�����"O6��e#ع
�<J��_�x�<U�"O2Z@iI5tF�H����Mʶ풕"O޵�i�!k��d�$a�i��y�_�<ON�JQ)6M��\�� �>�y��˼D߄�)��C4@���a���yrh	�~��)�C��-B1!��yBHܶXƜ !� �9R���Q�y��<9"`���Ɓ\�0����y��3� b �
.M�	��J�y"�X�i�ƽ�5�^%>'ĩR��-�y����-#�Pp�M�^�n��!B	��y2�J�X"�M��T�L�Ґr��+�y`Y�y�=SA��H�N1(�ʎ6�y���,�r}���.�lR��y�h�
�t�rch֩��	$�y�aݽjjj`cl�+���a�넸�y�È)+��X��\l0懭�y��\(A�rh2��+M%xIb �L��ya�d>q�#�8[#�(�LU��yrOHg��wᗝX5��vD�%�y�M�3&%L���H�&�2IJ��yrA�v��]s���V���H�h��y�O��q����{����镧�y��D"l�j�E�ɣr.&<!��[��yb	wJ����^9mж�@�`D	�y"�ȥHߪ	�w�g��0�ѷ�y� \$��HP' ��	��نc���y�W&z�����E1`,�Rq��y"{�|l��G��.�@��E���G�!�$�%^��	�/	��A�� �!�$�,)>Dҧd÷5�}سƁ=u�!�Z&*��@1��/���$&@�\�!�d��0J>t�5f
�z��	9u�o�!�$ +�vxK�-�t@�O�D\!򤓴i��pC�C^ܘc5NMnJ!�$^�c]α�3@]y��-w�!�D�.s����
� ��Sl�P�!�d�,s�`�t��4	l��z�-Y{�!򤒔fz�ɪ��E�t_puy�!c�!�b,(K$oM=�L䫒�@�)o!��P�)1���'܍s�����*a!�7<tD�A�D�7r���B�0�!�Če�zabt#0��4)�ܧ
	!�� z��tF[>l������"���� "O:��0C�n�re1@��)eI�؁`"O��Ɓ�?)��P���4��"Ox���T
@��88���GT]y�"O�@j4��%l�4���C-=�<�#"O����ŶZ
���q�����	4"O�j�g�]r�dK��ׯlX�x"O�HS��2+>X��b�̩{<j�K�"OB��L��J�9%��+pYh�"O�	��P]�i��݃I��a�"ORy�[�"\L�e��EBc7"O$@6�J-'�Tɗ�K�8T�"O�E�3 IR@.�B�n�.J�T�d"O��A���#yc�0CoI�I�y�v"O^��Z�T઱����$"O 9X���7k�9C�P�P�F"O�Yр�JN���C�� ��"O�\���i_(if��E���:S"O�DS3!S"+)&D�aMX�Z�Dňs"O�0Q��/^���a�lI%"O���R!A-iP��%V�&�H\�"O6���f�IuY�����U�*a�v"O��r��d��i�7n��p�
�8"O^$��D��#�X��L֬��"O$�`�V�pJPp��1����"OF��NN=�&haf���>��"OΙ�QHJ;�6}:��d2lT�"O��*V������7B3�"O1%��:��� S܂E��9w"O�yB���yj%y�oF��@��"OD�I`ܒM���fa\;X)�|x�"O�b �����N�S���#�"O���3̙�M���j#��3�B"O����'Z�[��7��!�`Z%"OZ �,�1,���U��\�21	�"OH�â�TT̍���ʤu�`���"O���ㅞ8F!�1ȤE�^>��0""O��D�H.�Q�
�-A����"O���7LOm�4�V�U0@�Y�"O��4!�;ԶjC�Ax��Qr"O�ta@ �R�ti"�J��u�"O��A(�
_�n��	�{�:��E"O^�"c�<;�{3S��UIu"O�հ"K�tn�`c�ذ{���8�"O����\�*�&G�T�.8\"P"O�%��H�"5 ��DKř�ĉ�@"O
1����t\H�**rF��SR"O���Ё��A�h����6Tr��3"O�p�B��uQ����`ȃ[μ�b"O�xS��@3�f���%�f� }h�"Oj�b$/�!���DT�l�"O�J醃w�(���D<��80�"O|�bRf�{b���3�E ��8""O�00��6=�Ĺ��*�r�
�"O��S�k]�&<���͐K�R �"O���LD�WY�� d�ey~���"O� A��Q�{ �\�2�T�[y��{u"O`���U)"/|��0M�&FN�HH�"O����')�]@�	Լd����"OJ��)O���=�!�4�F���"O$�3�,ۘ&dڜ�֫[���Ļ�"O ��Y�N��� S� +���"O�	�j��a���`��S�C�2�y3"O��Jb� &S����'�<��p��"O� T\pBf	�bN��x�ȭM����"O�}Ҥ瑜�RH��+@I�ru��"OLE��hW+�����S���"O��#l��IB�T↢z�0��"O�i��#˜@��c��K
Vr�|J"OJ�a�e��*]�8P)�:Wd�X��"O��A4ď�I^@���~A�`2�"O�	
E�\Vv�$�V���f.B@C�"O,m��B.S?6{ㅓ%"�\s�"O�p��ʏ�k�q[�B�dH d��"O0���9Z9&��wCJ:=RvM""O$�A�>jr��bu,�y[�"OR���
u��8�J�)��*g"O����z[JI �!X�B���r"Op
�fT�j���� 3o\N�Jt"O���0''8�<��&�+kU�0[7"O���to�J����&�HRx "O(�S��8^TjҥB��`+R"O�,���8z�ވ�QE͏Px>�rB"O�t��NaVt��MWϖ@�"Oȸ	��1:�0@s&����d�"O��* ��S�P%Jx$Iz"O�� �z�J��	�Tw8p+�"O0����M%��k��ͨ?X"��"O�ģ��Ք/g0�� @�M_��[r"O�$��'fb��nF�O$�%X�"O���p�ZP Ss��P��#R"O�����a��pᄬѣ#�ؠq"OĜp��Ih�"eK��=�BL�g"O��D	��=��Iz�e��"O���F �z`����Z#_l\�V"O����w����_2�n4Z2"O�Ȋrݠ)(�������1��a0"Ob0�K8JA��ƪ�p� "OV)�3��*̡֨#�5�@P"O6Q�c�ݨE�P˳�Ѕ,��0"OnXX��ǉF5v<맍Q"<��tys"O�qIBC������r�гjJ�9��"O�9� *��%,W�2He�a"OH!	�� �D�P��:���"Of ۴
@�H;����i�?@�T��"O�B�K�"�R��Q 9$���"Oܡ�"T&f�,X�dn�q��d��"O����o�`�K��c��!C�"O��F%"y�1�5i�c�64��"O
�A��`�>�!r�JKv�df"O8�W�A��H岳�1.]v�	s"O�Y�m�?@��%�].6��H�"O�D���Ƹ)�V���&�}�"O����_�"��X6�?QbQ��"O,HH�����i;�Y=(�:�c"Ob�� ]);�8H#4� �RQ��
0"O��RQ@���͈���'?.mH�"O�Y�cF�>�>|*�j�
G̮Tp"O�a�.? ̎��'_�]�"�@#"O������lhPeg�_��۷"O<�;�ΰ;���"��"��@"O6L�B��a����ǩgǈ��"O���n�� Q�	
(��b""O��D�ګ�v�x��R�n�fA�`"O$X�   �