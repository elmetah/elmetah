MPQ    #    h�  h                                                                                 ��A=���)�r����,��w+AT]�!��`�e_F��ۊ�F]�>�(��TNH���C�����Q�y��}��&0�)�>a��v�����\Mg{��4��c��3�� ��3(*��rfH����b^��� �ߧ�>�x�-�l�IE&����I���3n��Wh�jZXw_S�/��㎤\N@ =Aٱ�M�����>ag^���4����!���gG�<��y�]s�up���l��jۥ�����,����ӆ�J�H�{bz%ݗ/�:����ڏV\��أ:���s%8@p�ᠲ?�h����b΍"�}}��w��s5Ā�H2��D�z�g����;��x٫6�~6�:#lUiQ���p��š//�4����+]��8��u�� fZ�j���:ՁUV��s��[����� ����2"�1�Mi���a.�ڃ�h�V,�q԰�AԴ�^ٗ��3y��&�͈�.zwy��A��M!D��t@B��#~�њ-��K٦�SS��}i��!���}	�cB�A	.�9�H�[W�.*�ꌋ�����o�o	�@Q�K����`|VO�.2�R�%M�rǫM?�V�����q#XZ5[����Х�Z�|(�;�@�l�e'30�M�s��&ˏ��G;�))^�Ӽ
.(8%'-k��k|���cm�Z��s�.q	��]@�����3�G��W��1>��'�� ��:���=ő�D�=8��cɰ�KgcPOu�s�0d�T������T�]���ռ=Fw���'�P>ta��u�I�u��m����"|����y��_Z����`�o���S"%r������?��3�����O�l2�I蜦|� ��5��P� ��O�J����L��ٍ5�變�o�:�EQ�Xa60T�%.Ú�ס�^�ŭX�2�qa�J���y��91*� ���ԝzDRa�����v���}�LX'��zc�����&e����gn��u�l�0j,�T�����y�t�q�f����f���"�cEQ���ﯝ<�R�
�a�zx�ڪՇ�p���]���e�ERl͎�r=-4�[neI��l��j�7�J��cs�J�Q�HtIm�7kл�>�>���:u)���.ҽ�q�a�Rz����p3�_z���_װ5��<hC*�x�f��+�4�3�v�k�� �2��d{���K�w)C�!MYC�.S���z�F����fHW��9�$���UH8�7υ��[�`*/�"�yn'>�`�D�}|4�C�إ�}U� ;ڴT�#��wb�4������8�m�s�ٯ�wD�/x��8H�!  sG��>(m������+�\ �:� ���ܮ��6�Q0}M/���!�����˼����$���xH��~`Ƃt����
�O�L�d�䭎|is9��_�;�$ER�>�?�K_�<�u��8��|X������U�ޠh�Ǒd������ANͩp��kY��RZ}��J�'zTb�c=����HT�Q0� �1��4L�|\��l&7�m�ֵ��ēu$��Le
˃h�-�$8@��<)xA��U����ȣf�^v"H2�oRaj�� Y���ց�V_6,SרSظ����	`m?�����b�?��XYM�|ik��"��{�x��`����S�Iشa��Y$�E{iYpN��P
��Y9O s�ϵ\�o�-q�`qJ�� �oE?�͌��E˞���#�:��yv��%�'OC�Ľ{����@�@�C#0�ޮ+[���9���14�rSt�K&惞��#f�����g��I�����XgG�/�t�_N;���|��N�U�K��e�S��D�jS�/���E~C3�O��+	L��+�C��S�պ��������E��?�x!����Hi0|e���}����,��x��m�&H����'~+��z���R�#�����]����}�k�v�������!p	�}_�5=�)��:،����>����U�:͞��o2�;�g!��|q�㩙��X�)�e��x�t+}��`+�C鹓�K�ĝE�G_�jZk��nߣ7�x�����~V�d@/
�i:G�l�-�I�J�2GYl�i �ֹ0��P�� ��\=�UsP#�L����z���}ƑÌг��[����B�qʰ�u�ǘ��k�<�z�����J��92}}��]�ޑrs������]�2�{�1�T���Uu(/�$1���+GqH:�i�ܷ�"(-^[5���I.�
�Z�Rˁ`|�X*�w_c0W�����U�] ����J��2�K5�5��1S�����MC흫& C(���S�k��|I��A;��c];(6��4ё!� ��w�Zw�Y]����h
<W����-~����U"��^���s�+n��c�(Ş�+�^�~�V�SC��!����&�;����Lʍ���K�f<KO�"�1b*ďE@���/2d�3 tJ�2�D5����W6��K�j*�a#�;&隝��q���}��
4rr��Nlr��O�����4�Q��e�щ,ro]iA'��	op@�7�#H����e����H���;���bs��j��[��|&�u��,��ᕄ�:I��U�!��*��=͝��},zW]��G\���F� �t�9Y��w��O=��յ���W��������v�r�:�^���xPM�?�`�B�\K�}3��O���CØ�1���>RȒ���(c3��k�1����L�/ȥFW�%$%vTS��<�/I�y�V�CYm��^�i��?xS%�+<8��4:d��Ё��jy�����gPnVp2*A�wY-oP�q �Uh"���$_ �`/�;$$�FW2eə��~$Z�]���3�E��c|󗛭����ab�v�9G{�zYr{QbC�sf[F���
1�2ψ���G�i�+�&Dtx#��gYyV�P�=�����2�=�nE9��A;�Qs#���KN�� ^�YSK�)1O��)��K�2����J�5	m�ͧ�b_AOA'�����P�f?�� �N�d���_
4O/F�X��{ ���K�t�����N|�V1�+�d�	4�Z�.#T����Y,�۴��Yj�'?7C{^d���΄n(�A6���u���Zȏ^M�)�g~��T���3#'ޅ���]�H�-Y]���� ((��g����Ν��tr���W��%M��3����� �
s��f�M��o��#�g�H&��d��&H�I�1�����`d]#jp���li��`�^����qgJ�a��6b*đ�u./4҆�^r���i�\����~s�  �%ӯb���?*+͒Y�GΨ�1}��S�RBZ�J��5_[�H-�3D����" )��։	,��X�~q��:��1iL�Ls�t�x/L�J�K4���i�ԟf�S��^Zu�����lj�^զU[xU��hs�T��@��	s �I��ɋ���i/�a�k�����Vg'3o7�A.[߹�J����y��c~���\�~w��C�ܓCMi��_8wBEM3~
�-!C�K�R�������{����c�iA$`9Q�[24..e���'S������o�$6Qit�}��`W&�O
�����R%H������nVǸEy��#3զ[<ջ��(�РA��ט�;���9���<3��Mk�������BM�_GG���)y�m����8Z�'hWp���{Jݟ�E �P�.�ҕ��,5��sd3�>-���N�,�����z=��U����8�?��x:��ɫKhg�l�0^��ψ���we�i��a�]'Gշ�!wl�����Y�Ե@�Y�����mk?���5C|���c7��z�8�x��Jө��E�r�١�s�?%���q0�j�El�@��wy��;��5P����gVO+��|��-ԛ��b��[d��uIXE�#�X\�T��UB���8[�@���;���GJ[~3y�R��Oϻ���mDͥ����F�����?�G�c'�]Nz%�
��e(v���E�C=uZ0 �p,#Ʉ�O�y�k�qA���uf���"<paQ��t�
=��8��|�����M�/���]��x��`Rȁ#��݊=���[I�ɓ�@������J��sQ�BQ*I�}�k��> �?�$�/)��ǉ�Ag��a���$�[p��_�-����5��ח�#*z/of�AL0��3��sk�J-͞UP�_0�x�)K[�>)^��!���C�Z�6�$�^��)��W�cM9��s�\��H��7C���CU;[W�v�d4��>ѯ���W��C���?��3����7#m�����@�i�sXĪ�F٪��w�!/3#~S5���� N�um�����d��]����ݪο��W��|�/N}�ԍ��z������@(����џ�3�Sv,ƹI������.�O6�Y�s�����|�������vwuE���:��_L|y��~��	7��L����0���}U�ųh��d5�(Ө))�\
ة���FN� BZD}���
'�x������<oT4�+�ۅ��JTN9g����7C����.��%u��m�'�˾��-RL�@�U<����K��q��H�A"�v]s�2)AaPF�{����'�q�,��@�.�O��!+��m:7tB�tbk���=MO3�k�Hh�ļ��[,��N�?a.ˀY���{D��N�ۥ
BvX9JGL�*�^�*�tq6̅�[����o��[�'XEư��Hu�:M'v4%�oC�K�{�U��{q�> v�9+-[>��9��41��SO&!�2�b8��Mt�ᩇg�?�I��SL
X��JG>@���� Z�Y�W�7�SN6V���%�@�>S�+J��T	�*�Ġ{3��� ��	Ǒl+bvx��K\�������]����?VM�!أd��'�0WC���}!C8�� {�n�T�(B�&c�"Վ�\���+����#�����d���v�s���A�}*I��C������_gu��{����I�;�S�p��ђU��j͙�o��r�"�����#�^���H,�ef��x�Bt�|���1�����۟�"��/Rj�B��i�\76�{�c*љ��d����D�ϧk-;�L�EmG����$m��H�6lr���I�Y̷=O+Pv`L]f�u�ƀ��>�����9B6-nq��!��S������<C,ٸ�����ٕԵ�}��k�^r.Z
��L]/�{{�����@D�(*՛$����W�qc��iv$���^�^�G�]tI)�����|�{+�ӣ(�RA4kt��t�YU����zJ@$��f��5��lS^���u��8ۓ >K���dkA��I�A���c8s�6,����k!��ȿ�lpw�`�Yx&>�j��h���WYԑ�V-y�Q�X�"Z�i^���Ņ+I/�cr�9`��YpqԱ��C�}O!����/;{�~�S/�(�����jO�1}["�
�B@�x�/O���f�E�k���X�{k?6�#��Ɉ<�+;aSܝBk�}�¬P�-���is��M:��/0�o1���hф�]o��'k�@	�b˜��#v�MC�e�Xa�����ҥ}P��h1�61���(uS����'���?��G	�&�ɥgs�Z�pz�i�"�G���D?���tbP!��B�R�w=Hx���ZWE�/�ז��+��:��9Dt�%7Mls�`��\�H-�8f���ر�P'�s���ӓ�Rc1���f�����&�a��FL'�Ȁ-0�`�^��yg/�`Ђ~��^c�m��ɋD���zE�%��;8��4]A��u`����ym�N�֤�n�H�*�}Y(BX��2��j��SA$��@�;S�v��ᡅe�7t�tZSf��S�EؘcW�=��(����]3���{d�Y��)Qݱ�sA��FW�]8�1�L)��܇�i�C����x���g�}źۺ=��P�y��2��n`�5��;r��s^���D^�����bpS�a1jt$)U[�K�q%�5����	h'���_��aAB��q-�P��Z?������%�p��2
�wF��a�\a��8�Kܤ������x����+�:a	O<��#/Ƒ�����vW��O�)�L7��"��I �(�,���u�����o>|�H����͌4�A#bi��`A�Xvb��d�b���;vc�\���.���쌹�vWX������ls�)� w�n��2Mu=��Eg��������JZ�Ė���%���]���p�z�lg�m���0�б�Y"�<C禾��b�N2��-a/���\�dX\�9�Y�n�[�2%n?�׆�?�Z��p��̀}n�-��Ӆy5�UH(�DN0����-�Z����ϛ�~��:YiG����3sW�e��4;��D�#�����n/u�v��j�-Z�p�UL8\sp�l�#�DSE] ���=/1��<i2�Ia$ ��jйV���
��A�]�V��Uray�h	���7�sw�{��w�/M�^��B �F~%�-���K�셃��}�B�����3�cybA?�.9�S?[y�.�����:���cĜo�oQ'����s�`2�OE�5��9|%C�=�a�o�DV���>#p�[w�н�cЛ���2)c;SX�T�|2^3�-���8�M��~돺�G���)��/� ��85��'�c腡�~�vQ��,-���.����S92�h3-V�����'�Q�9*�5z��pl��3TLk�P޳\6�L�ɦ� g���%�	�5�y�@�B��]��ղ�w�O0ʝQt�𵻿���b���mo��h4|H����ɕd~��P��%��Ɉ�r�ɡ�q�?�O_�,��مjpl(�R�Rl��v��5����0O���7u`�H?f�+1�6㰢�E���XW>T_,��������̻�ގ�	�J�i�y��n���v�ڱ
 �DH
��mvV��L
�݅B��'Mǚzٹȶ%�e�%�����~��Є0���,~]f�
y���q�;.��Xofx/"לQ�@��e�����9����p����t��j��T�4]��K�R����
�k=#5�[$���T�%���O����	s�(Q4��IcY�k�1">;k=����)����2F"�Fa,�����)p��]_����h�5��/���*5�f����3���k2��9�(�Z���!K))y)�!C��Ca�q{�Ұv���k�;W�P�9�S�׮�H7~Sq��n%V����;�=�>��:T2X^C�c��fT�K��
�v#(�5��*ޚDOp�@O��y.٥��w�W�/�hnz���� )nm/S`������ڰ�����������[Z.�}��_���'�I��A����ux�.� ��Rԯ��r�O�v`�0���|_�f�k�:籋zE��U�5�E_�jv�z����(�ra-�_;c�� U4�h�[�d��o�cnS�w�J���!���BJ&Z����t�'0�z�ټ��T���ж�Wp�
��,�7�n�LK���שu�ɓ����Ȼ-퓮@zV<ߌ��1��w�D��ruv���2ĴaV����׷[�
��O�,J��	�V�x�Q$�m5I���b&0�*M�	Sk��=��6��sVȹ6�郿�aI)PY��{��N�G�
�i�9E�aׅ"!���qQ�g�*�d�zo����p*E����:�zv,h�%�v�C`�{���vE�9�7��.[���9��1*�"S*p�&\~���lB�u�<q�gw�	I���Ι�X��^Gy�"�;�UT4���8��NQK��A�A2S#ϣ�G_��%QX���Y3;�q;�3	Bu�+=�h���V�&V-��#���G�?��!�nܴ>V?02A!?p.}�#�����>��� &~`U�	y���E?+A[b� o'�\�j-�X����a�X~��?RC�W���q!_�>��p;��2#���^�o(�mUE�͔\�o蚩�� ���?��>�˨�Gg�zeOx�tᛳ�� �L���*��z'0��
j�:E�d��7���\��Ѵоd6�m�#��fk-��a�@#�G7���!t���ģ{I�۔҆=���P�	L`�?�0�$��D��y��\��C�\B�e�q�(Eh�s��+���<��������oYp}��>��r�6�4��]�K�{Vi ���g�R�(%��$�l����q~�i�ދص)^�y5��I$�;�F�=�ȕ2����NV��-C������U�-�t�nJ������5y�SS9�U��G��*� 9���uxk���I#;,A1��c�&6g6��j&s!����-:�w���Y��\���h���W�2���0%-t�ϳ{3"�w^րni�#+$�!cNۗ����T���yCn�!�EyY�;V4������u�m���OT6�1���ąH�@[|/���i�,@� ����663:d�`��ak;����<ǰxწ�3���������D0�����آ$�����o�$'&D�	�t��-��z���/e" ��^�I�5�`^��MG�`	��`�\�u������ReO�i!�A��� S���b��X�'z�8�SG_���^Ṧ�t݆�𨅝ߍC3=�`%���W�` ��}��S�h����x�O��Mǉ`ذ�\���������W�NX��kR���������u��کL�>��[4������'���R/�\'���y��mx:��5rõ2�%(5�8�4�h⣅���D/y�8R��n�@H*w}GY#5�'�,�˃����a$U�k�ݏ�
f�|�e��fY%Z�����NE�c29S�#���P�X��wj�{�,Y��NQX@_s��F���xH1��<�>dZ��E�i(�����x��gϡ`�U��=��	���2X�/n{����;M�js��Ձ[u����=��S�~1�`�)��qK��$`�ڀz	c���]� _��xA]s����P�`?�%F�6����`�K��
��F�[��f�p�NK�f��C����|�f+k0~	j��Pp�#
&��5�f�<�e����7�\K��0�ě(w7D#/�u�?��q��>+�!h�dc�����#�����ǘS"��㏓���V���������������߹���W�Q���.��ń���� R;�XU�M�ž��gQ+�e���9�ԥ?^K���@�*e�]D��p��l¡����ȹK�n�gl���ͦ�PWbK�8�~0/�`����@�+~�\�LZ�4�ǖ0�%	�o��)�?�'�����ї}w�����,�5�pH#��D�3���f�H�Ɖ��ҫ���~���:���iBD)x����桀`;4|y|����XA�	 �u�z�w��jA�����U��{sK�}�^�l� ��H��X�b�YiMqa���E4wV��2���AB��o/Ηw�y�t�̈�Xw*f]�דMI�!�B�L^~@-��K������N����73c42AZ$�9G	[��H.ۣ9�]Be���o:P�QB�st`&�O��5�#�}%>�mǼ}�=>}V�(oQ�#�*�[��Y���ЖC�̍�|;�oA)�ȋ3��~�&���ڥ���Gl��)���{r-8��'ޏ�<70�qxq�k2�ƈ5.�����e{�C�q3h��(��"���[P��@�`����F���q�矜ɡ�gtT�$nj��;��+�C܊]]pխu�w"״�X�$�r��6�'Ӧ�&nIm�������|�U�� ɰ��n�I� �����r�������?�,���!e٠
�l�g��-�ױmr5��I���O����0�c�8��7�����wE"E�XR�1T�_g��_8��Ι6�Ȼ��a�"�tJ�u�y�0�J�@�1Ϙ�%a,DÎ��H�6�'����=��'�P�z�n��@dKe����DŻ�.���'0���,�H��U/y��qVU���yfH�"r�aQ} ���ۑ�����	w�H-�k�͇��c��_e]��K�vU<R>��%�=��[�D���>^�;���Ll �sǌrQO�MI�TBka�>v1��Z��)���?���TWaG���.p��_+���0a(5��n�M��*��.f�&��3�Y}km�b���8�U�-�.��Kќ�)��T!��+C<�b��Kۑ�M��ƪ�W?]u9䰚�R��H��w7�EU�y��Q��,���D>���w�JCS�ǥu8���e�#�|ᅉ�������H�D��٠��wU��/�^�������m / Om�����+��!�k/+@��MIu��AL�}�)�Ռ.��J������5Sѕ��	2e�/|��E%籼ְO�YU�:�5�|��?�F�0��3E#i5�0�_y3�5�w�c�합�:�e�6@`U���h�U�d�,���a���%�����(�}��ZNGȉ�9�'�!ߔ�%���TT*Q�Б����Ԡ�E���!7��Ҋ����u��ѓ�S��4)-��}@uu<:GX�H7F��˖�������xv�)j2_��a|\�1�u�)e����,��ר��͗@�k��asm0����b�2�*�ME �k����:�TI2bQ�}�1%�zl�ad�GY��v{�K�N1�l
x}�9@5��������Nql~��T��?/o����]�TE�4-��wM:À�vG��%�M�C;�({H:z�/;�4v��0[�
&9�q1��S��&�+����|���X�g2ŀI9�IKX��G����R�P˿���G.Nl`���v���S^�Q���� σ�V��3��tV��	�x@+<���ź��u�l�V��?��!Z\����0_HzI9}W$�����$҅�&�6�Մ���+|?䍻��;v���4@����w���3���zA�����_(�n�����d�1������GgU��2͏��oC�������6�T��˃�W�كe��xx�dt<���K;�gi.��5�U�m��/�j+R��_�7�W���%��=Ud� ���9	��-qqO�;�wGj��b��
�,�V�����=���P��L�����}�����4 G��Ҥ�~+Bl��q��������)?���<9�4�}�ɧ�1�
>}�<��8r��%�O��]�\{15w�5�v�( ��$B ��Mq��il���,�^�j�p�I��?j���쁱���(ʐe��ݪ�CU�����&�J�	���cU5���S�L�C&�n�� 4�>��:k���I> A�ac�B�6��;��!�*���'�wEr{Y�fc�`E�h�EWϰ̵Sv�-o�����"�
^�E��+��c�d��o���Oت�g�C)��!��c��;1��@\�^���X�w'Op�1�)� �!@6�T/ů͍T;.�U����Ժ6N���h��/�;ׇ;�x.&�s����������Co|E��{����z�	on��'��	��ٜ���ٟKã�e����V������jT������)-(�u��X��I���b�$	��\��ɛ^����"���Sz(־���~Gm������ԙMtX��������$�=~iq����W��p�M�e�1��]����-�� M�:�`ӗR\\��ˮi�!K�����)ԭ�Ib=R�������t�^ל�m��Lv,�6[�����G�ō�S�/Zy~���"���om�D��f��?a%��8+54�ѣ@����yc��~�nY!*�CYH�������AȑJ$��b��F���-����e�Ӂ��5Z��ɖ��E_cٛ^�4��~KSe��2�{ڕ�Y��{Q��5s�tmF����1�lϙWx�x��iC�����<x��g
�s��Rz=�
��/Z2�pn� {+<�;(m�s�k������K�վS|�~1�l�)KZbKjO'�E���	^�N��_�_r��Axj��g��P2u?0� �ќ���I��Q�
e�tF#���R��K��KRed�U�j��.��g0t+&F�	��Q���#奘�pk������	��ߧ�7t���WQ�?WQ(Rbs^��u������%_Z�L{��͂B�u�#�kۅ��N��>��K��qrR�R��g��N&��Ek����WȌ~#`��>ބ'{ -.����M�:kŹ�g��#� kr�T򶥺Ezè�L�e]߯p��lnqۑ:��f8���v��&Ħ4b��֑y��/EX�珺I�F��\�&�.�����%������?;24�������v}��:��i ���g50��H�D�f�S��c��z����C~"��:�B�i=�d�����Z���[�4�����q�B���0�u�(�'�j�*P���LUBk�s&>���H�� ����@�3;ihB+a�̓ �V�p@��A	�v��(��˛y��������).wep�խ(pM���pEBv�y~[��-���Kq���?����"��醊c�l�Au�W9�ވ[�b.Ŀ��i�ݱ���Ao��Q]���P`�UZO����>W%9py�#!��V�c꼺#��[�W�R��Б� ��;�����xr�3n�P�¹v��V|�pِG'a�)�1,��s�8�m'���
�l����X��z�.��m�I����3�����$v������S��t��)c�!t�)���I�ɜ��gρ aK?m'���%�~I�]�$}ը\w}~Y�W^�\ ���Ӂ��a�3m<^*��.K|�'��0����a��!���
��?onrSz3��͇?6*��ʪٻ�}l+�������5!%���"lO<,j�����~u�!.g����&��E��XM�jT��Æ����C��S�u��]2J,�6y|���js���@��D>3��#��b��R���8g�'��zOC(�[�'e���_#m���KF�B0�$n,4�)���Ky-Lq���iL�f���"VFQx ���C�>����K�f�D�F�Շ��r�7N]��O���R����@�=�+[�$,���������[Y0s�� Qj�IYpsk<'[>����0/)|X�ǚ����ab������pqJ4_f����y�5��רU�*�f-���:Y3]:
k�ߋ�o���P��܉�PK�>J)��!9��C���i�������!��W���9�tJ��nH��(7�W-�bL�ܯ��e�>"]*�0
[��EC��?�г����_U#�`��<� y��H��$q�߸&ٛ��w�<�/d,
�dɤ� �f"�KTmehg�Ύ�nQ��&��)�ȼD�zf|�`}����E1��"Q���Z�P�5��%��Y�j�f���6��Z�OG]C�_��P�|U�D�!'��'�E�DM�+60_]�����#=�h�q��8�q��Uj9�h�oydF����WT���h�.��ך�����Z��!��F'楓�O�B��T�;g�l�E��I�/��lX7T�ߊ�`��0��u+���8��o��-#�@p��<�!�]ɉ�~�%���q�v�/2�ya±���s���#�¿,������{�:���m+
�S�Ab�nV�EeM�mkc���u@��hL`]� �53�aEgYO�{��MNl��
��9;�@�;�[P�q��]<�P�o1\����E���Y)�:~]vb0�%xEZC�,{���ݬ8��/W0�J`2[orc9�k[1 DS�s�&��h�36wK��_5g�ITa�ĔmX}PG�h�q2=K��h�RhŁN����7O���|S�uS�}�;�m�ı3�3���q��	8��+�Ι�?���\����o��8�?���!)e�4F0���B�}�Dj��<���Y>�&�,3���}���+�C�Vfܠ:>� ����u�����W���ֵP�������_x1�)�������[�����U{]�͊fqo���S`�����S��^yw���e7�:xV`t�:b�L�����Ն�01ۮ3`jƉٙZ��7G�r�҄	��ʳd,1��y?�X�-�6��GŁ��Uî�%Q~��~-�1�f�
?�= �"PYQL�s��i̙J㑯憳[h݆�|_B7Fq� ��Ǆ����\D<� ��X:<�6��� D}�n���Er_�ٮj]��{!��@��Щ(۸$�a˓�q�
:i纵����^G>�P*I}]��˖�>�����xDm�����E��U�}n�*޷Jq����]�5o&S�vs�~��	*, /t��+Lkr˴IY��A'�c��e6�<����!�x9��4�w +sY�6R��nhvW(W
O��۫-j�a�i�"�b ^�#_��+ژ�c�s�
rN�J����h C�!r�o�;F{��B����՗ҵO���1ή�{�@�l/ o�E6�?��Z����N6i�Vh���;RY�@��nKz�aܺ^q���H�񾹖W��� Q��Z���u��o��'��	��\�#������MeX���	��� 0��I	Χ)�V�C�ǠBh�u$,m�������}�w���$�x/�Ζ�zÓ]���G�_!�u�����t�S��^��&g=�յ�.�WV������:/:�^e�ʶ����#M=�`ΞI\��t�i�<4�v��pw��y:R4̀��|ϸ��W,J�c	L��
��[���:܍��/��ՂBua��@�mn_T���i�+m�%^��8
��4n���	y�y��]�g�nB�.*���Y{��݉q�Aݑ1��$K"&�̎�'q��A�e�����Z�@R�,t�E��c��Λ�5�����N.�-�{��VY�g�QN�s��Fv�.Z�1�����j6�3#>i^5|���x�O�gEJ;ŋ>.=�i0ߊJ�2Τun�a!��2;as�Vշ�����>�S7&c1��Q)�	�KE�ֿ,ڶݻ	Y���9_-вA�����+PZ|�?kϝl�:�Pη
 :)F>�G��� &��K�����R���m��+�{�	���Fq�#�E����G�)��N:��7/���/Z��2u(-��[MuUz�����	�y���\��-��P��#X�1k՘I�W��FJ�"x� �͋�B�Ή�ڊ�V.��;�Wi^/9�U�����O zC��×MF�Ŵk�g�8��W�ov�5MÃ�H���]z��p�|lxZ��L�C���C�]�����ʦo��b�|�t�/�on�J�v�a�\�g���z����%?�]���M?�t��E��<}u�ʛ�a��6�5��H��D_���4�~�V��9k�`$L~]��:*Ti8�߈��d����vK4rV���Gq�RK�?a�u��x-�j�Y�����U�4?sx�����$�l ���N�����i�3�a��ȃ�[bVS�ۑ�A֍�%Bҗ��Ty�jjH���x�w��G�H��M=��ˉSB1̙~vu�--�KLzM�z7�x�����D�c��%A�hh9=ԯ[�$.Qzꓱ���̷t3�o���Qx��i�f`å8O�f2�Y�%4va�r�	��V3�eH�#� �[(nȽ��OЌ� �C�0;��(���U3I��W���T�I��n����G���)�f�q�8�f�'TH��r�;�g&��!�4�<��.�6F�������3�[�^�3��x�J�f�W������l�d�ĚLɗ�g*�=�Z�l�� ��S.����]�Y"գ�w�E��	��f4�,H��\���~Rm�����p|Y��Onh�����d�6㶲��zSr��+"?�G��]�T�֪`l�K����'�	5��ȭ�KO�tY�h]ޙ@���\��Ǜ��an�EX�-XH��Tp&��A�W�Q�,�E�yy���qJ��yw�� 	fϧ�a�[�D��P��g��Z.�Y��3�('^��z
8��v\le�܃:"�/�����0�ye,���;5lyH�|q��G�D��f��r"���Qs@�v������}�s�!����%/�]�m�,�vR�%�[R�=���[�$���qa�������s=�2Q�!Iԫ�k�>������)w�����SS�a}���pL�w_��P�f��5�XA�!�*fJfH�_<38;Gk��h�
$�K��䚈KG �)ʴ*!���C�I�"��ҁ�����|͹W��-9Yb�H��HQ�7/����{�GK~��_� e�>=,����QC�̥��ǸS����#Y�tږ��v�����_�(�z7ٖ �w�*/��	^��J� ��tŞ�m #���͇��� <:@��CP �U���N}T����0�Z+�r�s�k)oы���m�ƥ.��{&����GO�����;�kl3|�v��-�b��EY@��&�_������>����^�������U�ph��Yd���Ӕ�*��:����˲I��Z����#R'AJ �
�c� [T F��G-��=�k���<+7�|�}q�K��u��擓=@˪I�-�*E@k��<�������-�.���=��!pvI`I2��la(����ѷ��F�ݧ�,x���^��:}�"=�m&;��K1bW�/�`8 M;Mk>���N�G\YG|���a��Y���{��}N�L
��96�
ז���9q�����6���ol3�͓L�E�86��v:9Z+v}č%�\+C� {��o�Gb��*�f�\4[*��9��1���S�%�&�M���r- �M��g���Io˭�?B<XX��G*a�2lF�,��!@#cN��<��G���1S�x��?R�+o��K3lۦ��	���+΁��z����v��^Ç�?B\!D�t����0��F�[}�� ��K��X7�}�&�B��z���n �+�g���
YB�{���U���1����9��;�(�����_�Z��� � �'�6,����U��ͅ�o�7O�@�ej�J��9��D�e�r�x��t������O��ڃ��x�n�jjaᷙU�7��E�z1�x�d������ϓf-�ֲ�1HG WD��@�!�"D�
Q�E��=���P
:�Lq�ͻauf�2;�*�ҳ6����>B��q��ryV�?7R���</2A�3�^�q
@�}���ONr!R��g�]a{�,��{#u�>�(�$��ʓ�Jq�Nib�C�iz-^�б��I�(�Wxß��l��'��-���W)����U�U����J,ox��w}5�zSʃʋ�VU��y *����k--It�YA���c��}6��;�!����>b�w��Y�&)�V#hQ�{WEص�ac-e�	��$�"Fƺ^'�
��E+���c�־ťb�E�T���C�xF!!8���;��L���ʔ����y��-d�O�C1�_P��e1@�GU/;N�:��1B�4��g��6����ч0�-�;M<k��qL�i���������g�9$�2W��[F���4��p�%o$k'W4	�j����j�I�9�*e����Z{ґ��ǽѪ�ۢ���\u��Y��b�c���J�ђItɑ�7�3��	�z^q����gG#��0n��
�tN��9W�>G�=��Q����W��2���Y�UM��� ^��ǧ� �M؁�`��|\��$텩W=͡�A���+���R��x��n{*�r��
�'W�LEU����L/{}�j�ĭ�/-��\���'m�!���
~�f�y%��*8V4ɞ���	�$C�yYf�B؟n}�o*H<dY���8<t��6�Lhs$�z����[�bԿ�MDe���w�wZ?�>�GE��c�5�ԣ�!ʿI��#H{P�1Y���Qɫs��vFC�%���1�\�O�����biy�4��#�xj�zg�ζ�&J=�����2��>n��!%�;�tsJj��R_��R�NȍS��+1��0)AهK ��Zg�Q�I	T�f�n��_��A���]�P5��?����r�0�\�N
�FY�9�H7W��Kȥ���
���d �%+��m	����!"#��������!e��f���D7��'K�5.�("�!Ju��_S���8�4.���xt��+�#N�h��c �D����N�����HZ�r�ľڊ{�)��FW����/�i��p ���	�aM� ůrgbo-��d������t�^�4���];p�npl�fu�J��6z��c�Ө�ᦪ��b!ܑoME/��x����|�=\�$����?�G�!%ڽ���:?��� ���/��}��&��y��q5f�H��D�{������ {�p��;��~��6:��i3�:A�­�ѱ�4������ ��t��ڱu�F���jr�֦�٢U8�sܐЫ�s7 �����P���Ji�D-a2���V�#iv��A�� ߀{��AEny.���ǘ���w����+�M��&�B컽~�\l-���K'���r��u��"�����ceB�A�:!9��[y�Y.�dh�.l�GԷ���ok�Q��X��5I`�gO1�.��Ò%/�%���Rn��VN�����#zp[c䭽��Ї�<̞��;?��/hL]3$���2f��#�}�&0�G���) ɼ�ֿ8�ױ'��х��b���|b���w.�f�?��Ծ�3��I�J>����!�����x�����ޟ%ܚ��Wɒ�<g��Yׄ�u�9��BH��G��%].�_՞͏w3-ʉ�=��𵧵��7h�6�mr�ŀ�tR|�,��
̂��e��r_�zǶ�Ջr����~��?�7�|b��+lv�w/�bx5W0��┼O��Ȣ#��޴+��뫢���G|E��~XC�0T˹A���]�.'���fƻT����~JbXQyrma[��bl�vDgD4�$�م���I��0��.� '���z�L��e�#�A��j�o|�0���,����Ԑyc5qwe���f��"C��Qn����9���I�0�\9x���v�V�,��FH]�x���4tRo�ώv��=��[�D��@0���n�d�s��Q�yPIO�k�T>'D��+�\)rz��PtXX�a�F���p'K_�㒽y5����^�*!��fc�H��J3\4k8�ͥ��F���?��K�{)�́!/��C�,]؃��~���WpC`95]���HZ�[7jܹ�JB��=̘�\�>Xj�&���nCml�F�s�뿴vn�#F'2����
����!��x�ّ��wf��/�'��κ��� �6 �m����
�$�ڜ��U�$ž��0'2�f�}��W��+��3��-�نİ���;���/����½O���L�2���|KL����3��E�[%�!4_d�f�,�Y���^���
O��jU�&<h��d��M�O���'���Tˍh�.3@Z�=��H�'����;��;`*T�pK�"���C��UȆ��,�7
lY�8�[�f��u��nb���	�-Y�<@fF�<K6��y��Hæ�������cv�+�20��a����B��G�͙���,�%�u�ӗ�4���?m!�u	��bF��{+-M���k�5���(�Bxq����� qa��Yr5{�^]N�8�
Ix�91���{���SUq�yyS�}��',o�*��.+�E������:�v.v�x�%n�hC��{�����n�%1� y6[��9*��1)S��&H�F�imu����Igc��I�U�ܺ�X3*�Geyz��QSA����m� �N�_��-`��7S�S���@�	/�gN3'$��T$	.C�+�T����ʺ�l ��g��?�/�!_��*P}0�x+��}(���Ɨ5L ����&�x������I)+-�����q����ֻ�q?I�+���MX���+ϋ�������|_.�����;������=���U��d̀�.oT����?1�\P���@���S�em�xv+tMY������\�u -��F�� �j�XN�P��7�VX�H��� E�d"����Y��Γ-B�(�,;zG{L;���y�[�����F��4�ۀ+L=VGKP;�L̾�����Mp����*����/�B=��q���Y����Q�Y	<��	�1���9�'�}�|7�Ġr�b����Q]}�r{�X\���!G��(C$S���~�q�li�i=�DQd^�����*I�o�D�43�w:`W���:��p�{dU�M>�ଁJ�Q���5e��S��Q����?� %�I��A|k��I��A[`cj�6S�g��PW!|t&���~wv��Y�6����h,=?W���$-`E����"J�^B��U^+��)c:���@s��@���x�GCZ�!<ye?�;��8��(�/;��h���2zO@��11��qZ�@��/vM��է�,��f-H�"�"6�jv�L�(�\�;�Fq�I��d5a�԰D��vd�-1]�[آ����k,oem'oT	�[���jμt�;e��9��	���*�L�^�,�Lˡ�}�d�I;uZ1��e���:��U�iѭ�&�A7�_��D�z�n���V�G~�*��I��%3dtɠ��ݪ�y��=OC���W���~X��p��T����l�;bFMsU�`��\m�d����rfȡl�ú{���Rj*Ɂ{���;�����Bk	L���Ǐ~���5nq����/k����d��Omd��<�á'$%��"8 �P4$F`�qN�?-�y�.���n�a�*㻈YA������:ӑg=�$A���~&��W�����e�-	Ҏ�Z�q��b�tE|i�c�D�2����D ��Kb{ѐY�4QD�s���F~�d��1�0�Ϫ񒇩�+i�A�}�xEA�g�r���u>=��G�@'�2D�n�CF���;���s����B菼v�qES���1�Px)�ȼK���L����O	O�,��|S_�o�A�%���Pp?�z����A�0����
���Ft��ü9� �Kv��&���/O�xO,+WG�	�ݍ<�#v�{�!�Ͳ}dx���i�G37���@$��I�(㢡�u�������6�����	�v���1���#���g|C�?��O}�	0�����������R������>]��	�W�����Jj����� �q��D��M|�ŪϮg�p�Q�%���Υ+���9���h]�\ p���l.����Ϲ��8�S��Ӄl���b��B�j��/V����"=ɗ&[\x�ؠt,ǂ�%u�+����?LYܒ��<�J&�}k�N�t��Ӭ9�5iH�aD)���T������� ��ʭ~�<:`�i.hY��ڥM��|4h�Ұ�C �Ƚ�u"Ou��m�Ѡj-����U�'�s�ɡ�JZZO: �CY�x�N�xi�ua������Vɂ#��A������V���kyI�^`g
�~vNwO�~��M����r�B���~�c�-�GK�̓���庑x���_��4Qc �\A�,�93[T��.���ɠ���*�o&'�Q����_��`y��Ol]����%*���(��)AKVi��[��#UV�[�z�#zpЂ�T����;�Be�M��b�3�j��ӣp񩊨���CGXU�)�S�g8�8|h\'ʀ΅�E(�]Tk�׋O�..)�ݺW����M3T�G������_� aN܉���pz���������S�ɍ�Ag����*��w�I�Wq�/Q�]�"5ՙ�w�4�D����T�"C��S,m�'��G�|_���I��.��ZKT�lbW��r$�&�yG�?G���ӄ����l�5��
+םfq5��'���^OMe������6ԍ�@�}����@�E��X>�T&mu÷�I��" s�/�P��?J��2ymlt�����:��%D��D��دY�#'U�)e4'�:z��f���-e
s̓�����xd0��,E#Л���y~�uq��j���Df4�"�[�Qi���,��o���$���������[~Y]}���⾱R*����L�=��[k�_�{k����Q�dWl;s�O�Q��vIʂ�k͇�>b������)m;�ǫT��C�a�h����p��_5i���5�P�׹�*�`f~6Z�3��kY�?�@˫�A<�ܚ�8K��:) !!�@|C�~�?ҷUry��2pnW+�v9P���>��H5_�7�Nn����=6��Xp�tP>s*V� ya�C?� ��ݷ������%�#���M�D�����(�թ���ٌfw���/�U���ߤ~;� p�	;�(m6���X��e�WR�p�~�9�;�j@-�}�V��0"�l_���1١�с̈́�u)��ar�������OOX'�l�願�|Ƶ\�������!E�����_n�!I��t��٧���N��"}U;�_h�}.dWR��
������y�?�h��i��Z����̍�'��9߀���VǁT����@~�~i+�D"��<�7e{Ɗ��jƁ2�u����I��� �-���@a!]<�p��4��c �yf�c�v�y2��a�S���~������G,n��Pt�,_�X��m�6dL�b��n��>BM1ok�ܣ&��=���^S�fG�a�߶Y�3�{fO�NEl
��9,�R�Lb.��5q�bO����� o�A��)pE����j� :��v�L�%��C��{46�}p� �G�[�8[�i49EIK1���Sq�A&� T�T�hݞ�6gP�I����5��XǔG���B��<�y&���N������bY�SJ�Q�Nt����#3�i��$	���+�G���@
�-�I��^��?�#O!zF���+0y�f�-}�fu�ט\��_i�Zj&Ϭ�p�+�$r,+h��'�� ���1��,IY�F�ȼ��{�f>��^.���z_�DZ �V�|����I[�3��ULBe�{�Go�@�_[�9s��@�q���7�.qe�x�5�t�Y�}6a�ӱ��E����D�䰯j��K 7XA���M�;2�d��[�f���	/-ݻv�'��G�a���u�vy!��5��uۻ�_=��P \L'����&�h3�� ������j0�B�`�q���/�bǵ���((<%���鼳��bvk�}�3�[�r�Ď��y^]��{�����{n($�Ej�9�q7"iXq��H�^�T�!�I3�1�o����,����t,l�����8U�e��;�J�TĆF5���S���/c�ژ=  ���<�tk��I�T�A�C�cZb�6���q��!w"g���w1�Yg��LSQh�rW�鳵�̺-[�N�z5�"��{^]�����+k"Tcu��ۣ��;(o��RKC��!W${�;���,�C�ʵ���w��� �O���1"���nq@�o�/�lI�p� '�P��F���'c6�F���&�^��;�pk��4S�_ڎ�rIa��o�>��/YK�*0�ѐ
�+�S�f��o�ԏ'���	,�ל���Es���e)&'��DF����oZ����X0n�nu�㺈�k� q�v��9�ɇ�"�:	��9�z��
��'AG�����E$�@�&tDw����ߴ�=�˒�֢&Wg�t�9���鱕�#Գ[I��v�eMI�`�s�\�}˚��������Õ��5*R�q�v���׈�7�]��L��.Ȣ6�����7����1/�*܂s�6� >�m�̋f���ܴ�%/��8���4У,ƶ�Z7yO|z���Cn���*~[eY
���� :�rx���2�$��8�]&A���J�4e���-�9Z�:D�}��E�L�cy�Q�J��W�?I|>��{�$tY/i�Q��	sc��F�A���
1�$C�e1�d_�i������x ��g�6��\��=�F-ߛ�O2��n���F;���s��Ո��F=�;�Sh�i1�')7�]K֊���ڇ��	J<o�$q�_^�(A���Sl�P�k?`��=��P�)
Q�F�g�>b��U^K>fc���I��Z�ә�+�	�*2��#Q�g�\�9��c����K��7`��!x�+�i(�M�J�u&�+�A֏� �;�$��na���:e#��F����:^J��H��f����>����S7�:�����ȹ� �Wz�jj��ec�ٖ �i��qM�6ť�Gg����~���Q��#o�D��Q �]K�=p���l��y�}ٚ�Ҵ�Ψ��^n?� CbR�A�e`/�u��{��ɲ� \���{!IǽYR%='��8I?���vy��e��}�@C�O	5��5�՛H
��Dp�T�?�ؑ� |�f�:���~t�:�[i)A������q�� 4��f�ϟ'����u�n>��j����U.Q�s�"#�����Ju ~��_%a�	�ji��Oa����\V��e�A�#��6N闷nMyd�t�&�Y%�wQ�M���M��"���Bb�~ǊH-~�>K�'��+}��U�����}�U)cۗ.A�>�9�t-[/�U.���dH	�]��o�l_Qɴ���Vr`TU�O�$�*�.%%HBǃ��yV�q�֪�#0�[�0ս����}�h�T+;��I� ^�%3�pR�u�%Y���jG<�)6j�⹨8W�'M�C���X��22��m�x.I��5$_��V�3����/_|�	Nݤ[2~��)�����������/�Ɉ6�g;��Mtd��l����b	��j>�]d��Ք�3w�[-���Ea���n���M�m��A��:J|j�����7����C�Gj7�+��r�d(�t?�_������'zl
y��t����tS5��K�؆�O�(������aύ���XU?�ZdE)HiX9VgT�@I�rYV�d3����K�
�D�I�J��Lyh������ͱ�&�D*����ȯN���=B�$O�'o��z;֘����e�����m��d��_0�84,�w��lt�y��>qm�N�ճ�fo7k"yH�Qd`��M�*�*�9��R$\���ׇ�����"]x��=i/R���=8�[F����g�BI��z����sn��Q։�IEqk��>���a'k)h��U��Oga����n�p�a�_R�ӽ7�5��O�C�*���f����@�3��k�9�����<�C��=�Kx�)`!%�NC����v�R�FtW���W�|q9k�̹{HHO7�����|8L��HQ�>�Y����T��Cz��|"���z�,��#���hȗ�/�f���RתK��ه��w��/P�~�̤��8 K�LvX�m���Ƴ��F��+D���Ŵʻ��̾h��}%ܤ��i�kĹ��Z�ټZL���P7��V*I�L�e����O��<�Z�^|A?��JQ��_E*�ݽ��_ɠ&�����A��T|������]\�U֓�h�#d�+}�Ū�������C�ZU�9���^'R���;;��qNaT�%`���[��^���U��lL7��S���Ɯ�Vu�@�$��[�-��T@\�<ˀ��3�~]��f�>�;v�!�2f�ja����-����. },�.��+/��g���uKm�����b��Ԟ�q_M��2k�q�a�P]u8�X:��!�{a��vY��{A`-NXq�
�s9'��קhq�G��q�kmI��oyz�dHSE�����.F:j�v�@�%dc'C�{�{oE��������;[[Q�9`(V1�USL��&�mu�HceH�^��g���I�ɂܰ
�X��G�	ߥ��I7f¿�؈T�xN��#�i=�1S�B���>��%C��3�a�t	$j�+_Z=�+���ȷj馹���?s75!��U� �0T�}�g}^T��L��r�E��& E�������+��������u���X��r-�a{e�CAOz�֡ͨ������L�_�����qǌ���i�n*oU�#��v��o
���?���T�����.��`����e��2x�gt�@�8E���n�k��ۜ�r�a�j2���F��7�K>�B�V?�d3��A�9�D�U-xޜ�"sG1�M�A��֑q}����������=�BTP���L�_ܻ�XM�����@����`��VBsYq����P��p�=�C�n<����}�"?�ό}�
a`�rKFS��2�]s��{x[�,y�}J`(�>$	'
��4q �?iӘu��^�^3G��P#Iqr�h=J�*D́8u�0%r�O��Pݱ��U��~����J]w �#�&5[S�S[j��j8�u�� �����k^�.IŹ�AL�c5z�6��)�&Z!r���O��w�M;Y5��Ǧ�h�W�еZ�Z-VW�����"w��^x�K{�+F�c���v���6�&�.6�C��!rJ�[�;x� g!�eqn��!�>/�O�p 1:3��g��@}3�/쫺�ՙ"���b����6�Bp�B�]9�;��Y��
�Z�8�ͭCJp��&%��#��D��P���d�a,�o5d�'�DY	G����@ 8N�D�eč�����kJ&� �:�O�Bl0�3��T �u��/�����t�d�˜����C�x��$þ���z/ʉ���G4�4�aa�[9�t�m���H���j�=�tW��^�W�����g�JeQ�6��Z9M�\�`��~\#uU�U"驨��b���p��pxR�r�q�;>"�C_��x�Lwk��}�a����N!獵�/!�3�.ԅ�}7mZ)�A �b�%�P�8�r4��_��C�ua@y�醛���n.�l*�Y�"�I��-�ّ�G�$7D,�8��,pe�	���*Zp#]����ErP�cT
���C��*3:�m��{���YJT�Q:7s>�=F����F1�8��`�o�^�i��N����x���g1b��,/=�%O����2�3n���r�;ops���#�:��_�_$US#��1'�?)�kK��E����"$�	E�-��m_�XA�����<P���?Weҝػ�����mN�
%eF�� ��'���Kyve�\���%!�.=+͒�	��2�#,�������I'�����R07u<Ў���=(���4�u�p��������e�?����뼰c#�!���5�(�49�D��fٹ�c��tO�u�L�l��W�W��:%L��|ׄ�� t�� �M��EŠ�<gs�L��J����<�!���ﺙ��r]�o�p�u6l�K��8�j��N�I{]�9���[�-b��ؑ`��/X�6��ͺ�\n;�V����8%��ڝ��j?�7�1�΀��}a��*��" �57��H�QD�〳�e����X��G�����~I�:�^�i$:�K*��P��"#�4^�F�A��>����cu�2��8�j�T�-�U���sm�T��b"�f� yA���	��!i�7�a����g+�V?�G�A�}�ߑ�[�r3yM�V2�4�iw���մ��M���7�1BKB~�т-��K����f2���*����7��� c�r$A�p<9)�[
�.=El����S���?o��uQ�ѩ�U�`/%�O�����@% Κ��=n�V�ybQ��#,�[�Y�q�xIy̯��;p���3���Cv���aA�R�7�0G�B)QH�][�82��'@9����Sџ��j�(�.d�xݰq�e�3�x��=�� ���#�R�7�-���8�h��P�ۚ�yLɃ��g��`��HҔmj�=����Ku]�k�ՏE�wD�rʺ�1������,���mC���M`|�#a�;�j�R�H�P\��"�g�f�.rZ��o�$?��J�I���Bk�l���O�r���5(�g��/�O��T����ҍ�V�3�A�M��EĨX4�,T�3��-�H�i��P��鎄G�J3[�yc�Nl±ϓi$��G+D�Ii�j����עYt��Y�'�(5z�J���̏e rn��]ƻl�M��0�,�딛'ty���q蔾���
f��;"U�Q_ V�⷟��щTvl�IИ��Ї���M�]sYh��3�R��h���u=��[!d��A���+;��u"�"s)qdQ�A|I��>k���>�v���t�)c��aug?{�a���t p�7&_�7ҽ�Ԣ5��7�o��*Re�f�2���3�~kϬ��v�5�7J��P��K3G)6�7!�YmC^9�n���Rso�蒣W�IP9�)��4cH��7�����3?ޯN��>����ƀ/E#C�Dƥ���r��#E������-A�\�KϪ憩قl�ww�6/F+ށ�t�� &^��+�mlM?�Tc�5�G��#����/�'��O����}��?�����<��^� ��U��wj��+e�Ƒ���-����ONK}i���DV|����h#h�N�QE�n��_$od��\�����pѻ\6��[�Uqz�h��sd%�Ӏ�n�4kҩo+Z�E���Z�P��w['�T�������T��г�I��si&�!����7� �iF�Ʒ6�uw!����˖
�-*	u@W7�<\EI���V��ڿ�o���! v5M�2a��A�S��x-��I��,d���
˗�S��s�m?���bCy���ĄM'gk��أ�F2���3�b�5�����a<_Yw�{�N���
�39"����t��@q���?�a[zoXЪ����E���� �K:%��v�T�%���C]R{���ݳH��h��=[Y�9{'�1�pHS'-�&�ڪ�:]�^���d�g�U@I۳��+80X�`.G�ߥxpY2���/�v!N;��i�I'S��J��)�c��x�z3X���4�	�-�+:�>�f=�c����x��?.k�!�|���0/�� �}��J�� ޗF�� �m&;��fK|��c�+�8��] �������%����|��� UI���|u��;��_?@)С����y����f���(U�%��q/�oe�-�����o3�68x˥��`e>e�x�ot^�H���L�	t��01�w�ЮZ1�j�b�A��7v�y�z�qlFd���� ���-!���9G������֬����ףxuZ�1~�='��P��?L��6�M����~��{��5j���Br;q�������+�)�^��<8k��^ɧ];��R�}�P���r�ۮ�P]�6{S���g� 9�(e�$d(���=�q;��iNೋՕ�^nY�W��I�-��iw�����S$���ѐ*��C���LRDU����R�J���> �5�0xS6���7A��� ����h%k��I�>3A�t�c��6�����!m�|��W�w��'YP'��B0h��*W1F`����-Q��0�"2�M^�^��9�+!Yc�;��e�1�ԉ93C�s!�����#;S"�u�� M\���ʗ�]�OqjY1Ud ����@X/' ����(�wٿ�S�6�^��E��l;9%<�x:�U�^�(2&���A,��%+�~�G[��a��\ܯo�5'C�	bsǜ����%ŧe_*����$�}�]U�����0q���u+�|�������M������}C���^ ��E�z�'��)G����v�v��t:��.��*�= =4��:�W@7��L���u�����K����MD�[`���\~���t��áj��3��K[���͙R;�ʁlv����;���gL�b��X价8x�*V���U/|Ë��;پ6��m�k؋�o�R/�%eś8�z�45����􁐫yEw?���ni�~*��FY Z��E ��SC��|'$���f�N�&�v�e��M�F|Z+,ږ��E�s�c/�.���<���I5�Z�{<,�Ye_6Q��<sKF/�5��1�l�ϻ�N��|^i�ç�yIux֛gl�Œ��=�$��Qb�2u�n8��w�;Jis6��վy�耺��-�S��71BU�)-W�K�����ڽ�2	@Fh�ڹ�_�N�AՏ�I�_P��F?���s�@����ȭ�
�o�Fŋ��4�m_�K�����(���P����%+�h�	'%��#r#E0����N����~?7�aZWH �!\�(t��z�u\~폣I�G��� ��ZzZ�dΎ�F�#:su�8���0V#�`?�:4�g��4�i���ΰo��H���>W0.��M���r� OՒ����MM2�śՍg�4º�����ꏥ�Rr��QF���J]�)!p�bl?�~���>�����m���ݦ�mb���[m�/g����u�贤\�Z�1��3JS%F<F��H?]�Œ�NΛu}�1�� �]�]5Ҫ�H �D&�������\��2	~��:1čiS+�b�F�=ށ4ٮ���ߟyY��F4�u����,j^#��H�0U$,sH46��7+�� t��"r�m�i
ɒa�C&�BohVz`K⒮A��e�젮�-�y�������w�M��O�tM�UEiBغv~�8E-ta�K�;����勧C��9cQm>AÕ9��[�.x%+�����J�;3oWX�Q�U����`
BO�i�`N+%t��9�7ZV����S#��Y[O�̽�R��s���
,4;+��,'�Tf3��d~w��[�{��я�]�G�i�)lF��B8�|'{E��y�/�N	^��ޘ��ĉ.���+��@n<3��e<����5~�)�H����C=ދ�Ú$�8�~P:g���	������N��x]�@FՊ�Hw�
��ug�Lyr����ӣ��W�m������2| �y�����m���˔����綡"�r����j�?X��_��]�hl `[�*���N�s5��{���.O^����T� ލ%��q���E_)�X/^T7G���6ߡ��O�����J=����J�F(y^)� e�Ns?�∧D �m�E���FR��$���'%��z�ߩ����e{!a����V�(�\�0��,V�w��Lyϻhqc����'�f�! "��QZ�p�=w�����ox�H��h���B�,��]n�����R[�#�ⳗ=�8s[�d�,��x.t�}��s�1kQ[I;��k^�>���Y)^>{Ǽ�l��=aRp�w�Op�-:_��d�m��5ʴ;���+*<�f��~�@3�k
iH�6��2�ܫJ�K�)Qr�!�C9�TI5�҈�j;ݟCTW\69���̯j>H��7VeD���Z.�쯩���{�>�K��
�C�!�������# �Z�\6�J<6?����vR�}O�w���/ƞQF#�� V���m���Iڈ<>���Ū���ޟ�}[GҐ�;��!�������p���P������������Oi�8�v��J�|7��C/牭�E`
w���_]b�R���ݝJ�b�7�<��zU��h~� dh>-�;��OG��ꊉ���4��Z�����'`�߱�G����T�Z�Ў�G�/�&�z���,o7viΊ$�p���{u�ޓ�5)��J�-�PM@Rr�<��Q�e�r��wX��ǡ��pTvp��2�ɡa����nJ�3�ҙd�,�%w��S�ݩ��)�7mdu�_b�t,��7�M�=�k��/�ק]�N�.(�QG��{a!�oY�7�{��N�)O
��+9f��]�7���lq)ށ?���<W�o�G�͚�!E���{�0:�)$v��%Z��C8��{�)�NE�e��l*@[р*9�F1s�S/&4h��ՑxY�o�,�gO�I���ܦ�[X�]�GQ�!-l}�����WN)t�����lS�hE�4l�������3�|�	�+���뀺�����*��
?龍!�G��J}0
���}��Y��ɗ�Ye껖�&V�����f��+�$��K>���ܜBun]&"闝��9�>0���L�/����@�_�	l��'�������}�T���UG8�l�{o��eµ~���x9���Mˀ��30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�+ڜ4X{^�wLРr�A�}���Jdq��B�Ϥ!>m�gخ���T����r�2����,����.��km�EZ2�X�?C��>T�Gt�U�����Z_4�ӫ;�T���u!U�Gip�L��C��S��S��!
,/�0
Tf���3�^C�Q�$�Ť�^��!9]�f`ay�ȳkrMX�6Q.��� �1�F�j���xߖ��0�Q�:��澀��MN2�x�^/hĔZԙ^�O���T�J`�%�/�?F�)w4^�> -\5�����ek�#�M��\��T6).f,n����Ψz�f8p]Sh���駛f��ȕ�����wձƌa�P��HiUqXB���|^;8�5����WA��j���K�97ݪ�I�	t~���5c�&�N8�Q5j �d|�j���m�z��嵹���gV��	�XH�����,�&�Mô�F�J��Q�����J��9�-���$����d�O@��#.���i+h���ǯvk'}�PH�55���[��YB�GY�u�;����#�Z�˅ʶn3f��4�di�&�ó�y2ኍ�B�|�n-��S�[`��1����ȉ�i����k�W@�|J
@`̱ޕ&�v�ۓ]�o�;�k��ZE�V��"i�]p�$����Z���g�4f9�Do�1���"	�}�0�'4���ө�|~S���o>�jt���Y!� � �I3f
�|y0�!����X��s>B�,3`7��nI
"y�V�����m�#\��$Ò��@b �^�l5 e0M��L�#mF&�q�u��4ψ���x>�H�0��PU�8e�.x�!mR��L�Wk��X���������]���}5��rdX����#��h�P��6;�?~�^Y���������)��ht�`�rY&�h/���v-8vUB�>Ȁ럲�c�D�%σ��yj�-��h��y�>Ĩ3#O�P��oߴb�w�9�����ˈ����pa���c�e����u㘾�}���)*�l*�����6~ӀgMe��%*D�7%q�62j�?���
���W���le��ӈLzym��?!��DL��0PШ���m�ڣ�sL8V�Dz�>�H���ۦӻ.+��o^K����j�I��(@���M��L-��@ϸ�|}��� p6סRa���x��vEL�;t��!i��� cx%�!}�Q����MZc��;��������.�ٟ\�֞V� �e3(���Z��)�l�G�_��-�a��♧���g0��o8�<���B^VL�?�Y9NF��%/XOO�ok)��D���4�S��Ҳ�d[H��\6p��s�� ��?�t�hG+�	�:[���?JN����l�
5��4v��h�̷�}é��Y�YP_)o+�Q��5� �������L����KO��֯�'�C�R$js�$��=C���_�I�@aǄ��C�[���)���\��eﮱ?��M
`v:z7�k/��b>.  �aF-:��K�!��<�v�,N[�'�'FW�~ߵЎ�GqKO��[H.��S������ѐ�����{r��X�b4���&��*:x�b������bS4�o�n�\w!�	�*b9����~<X>���:���l�/�w=N�|�r��:�d��yQv8�#�U���5)r��%��ۛ ޕ=
?4MZQ�jϖ�"�#1�����+k1q,����1���p,�������8F5^��:-+ ��m�}~E<��Lw&�F:RI8��]&�y�M�o)m*ߒM��s���J��ʍ>Nע6��c�����`8�1�]P���q��oC���+3=����&��@R1g`pJ��.z-f����c��^�~�[�]ڬcFan��l������t���p�=
�e�$7x�F��+���Xunw�베m��A5���L�[>4�0���>m�%ծ�3���*��"�q2קs�#w^�Ё��|mG�*28Px?�}H>H�G��d����Ȕ+_늖�.�z�eT�uXM]G�o2L��x�qtV�
ך!����PT�{}�jP%�%���Hݻ�����!жjf���Ͻr����M�t�����T�!x����������������Z0��4M%|5�r�.�/MS+j�-����u�I3�b�� C3x!մ�{�R	�Z��nۯlh0��b����3�'t�}z�Z�DݔX�I⁴���5�M@;z{����J�@����a�eN�=>-'�{H��w-�F��:RΩ��[?�ڐ�c�#d�@���?�!�1(�	8G��p�g}�nc8�x�G~���m�t��=�:~�=�po��k��:��a����'��A=�Z��	A�k(a���M��cb+��%�/�@ �̈́�{��4$w�EA���#�C~ih��ۨ����P$�-��#>m��(ەu�~c�OߵZR�(�6���ΚB��������~��_c��G�:J��e؃JNy���)kJPf-�� \�u�Q�l�d���y�H��e\jC���y2�ܒD����x�j��w S	v���$� R�2��˗e:D.M���h�ICW�]	H,�t�������Y�������Ft1(z���j�3k=����G�R�Y���n�+�h��V13j\24�F���z�r���')�]�@k5��?�3�����Q��`OD>R�B��Nf%�@IIbetϣ�\��1]D֚>�t{�����Aa!�ׯ�9�簌�h�������𬨠�K$�����D����EC��	69P�xl(��6\X��?l�:�������ebY�N������_�P�=�VXϛS�����N��3Ø`��<��M��U�I�jʛ\AC �ɣ�.�vپu�.p�X\~��^u͠�:G�C������Ku�a�:�xG�!^FN6�OR&u�~M"rt�g�_~�|���\�+)}�WO�{cT�Rˡ����\��)49��b\2������R� �=�U���^)�\nSD����z"m��70�@�IG}����Rd�����K籮���'�a�U�	�5�<Ʈ��8��5==Ȣ?��G�jaLK����gl(�fV.��I���P�c��8��j}���-v�|CbR�w�z�R�ӷ��}��5	���H�U���3�R��ę�i��^V�C�5�1<d7��@}��U�cl�A�^5�kv�l&S�/��m�0�J�O�p�x����kO��?����F|7��Eb'<��p�xW�"�I�z
�Аi`� Ҩ�����Eu��
!�����n��m`�k�v���r7���8񧃻�,g�oM/Tm2QC$yԥq��&���m�~u��@��,qA�љ�*�/�J�� �|X���~�ڂ>�w��+�kJQTӯ��ԌP�@�|kT��=*U�VFp�h7O�g�>�p%:X�0w%�h#�S����ύ���j���r�7�і]:�A��d���*rK�|9�~+0]��[��3:�ߟn��L������N��1��{��.ҌL����0Va�p�";�H��E�9�Y�&��|̰�7��O&�a;`	���-3[���'`�;Y��<cSn��6d�dp� [�!�H�m��kz*;?��L|E�@,�L�����=V���H�m�C��[�"9=����b����d��]���@��4+�7�gp�o�?�7��s��SP�����8���T,	��'A�π~�<ɉŨ�����o�/�r
 �"�m�7MVcYʷ��������N��ۣr���IV���;��yh�Uz�[�:��mQ�v5��({g�;}�� ��}rC�� �UZ-��BEj��S�
�A�F�|}=GB�"OT~+NDW	�
��p
��oob^���B��d����dh�W�\��\��L�螹�1�	��3d�N�	�~^��u�ը���}����1�hv���
����X�J`��z�b�ՠ�������y2���uf����]��u�D��W
�&7�35p�=��{��u�	���rV߶S'��
+�j����Ѷ��y�J΀@���rF�,��ĄnK'#���̄h.� ��7��2��],P/�-�T��Z��	�.�mqV^�=�=�̆&
�6�1��{+Z����k�]��vs��t���&n/G6z%8S�W �m�f��!�sV���'�LłG��A�M��\�9m������Y_h�q�Ú�dɻ7D�MHB�U�2SV�'�AH�c�X��!�?0��쓉��w��4���U�
'�/�,���yz�f�/�bB�46-z��0��Vw���6���/��}Tq�F����x[R��>�^�����ѧ�s�/�0����,�=ܖ���zۧS�`�%�-� ���r�����|�CLD�1�z��R�6yBM�?#��@����z�:��φ�j<���'�B�u��� T)1��*��3���.����/�q�}xq �\i��*�OÜ��XAd�h.H�D��R�p��Wr�,i�L���D�;��E�E�{C8��D#P���{�F��~�+'��P����,Ci��Ȕ�핉�mT"���W^���PsR�u����J��A�r�𥠋���U��yT��
� ,��]�xppZ�����K�.�q[l�#3�y%v��S���Հ�I������̊�IAl���8q���huBh�^̖��:��ѫ�)�ϣ���"����9����T^�C��3p;k��B�<�vY�xQ���0�6%��;����O�M���j�>�l]Jd1کS2��2�h`����J��{W���V*��_�E���X��w��$�<sÎ�Pl�};�Ҏ�_=�Pd�De�������9* �Szl�;�}f�z��@pFƗ��'s�F9�L~����j�.�?;V�z�ƛA��ҡ�h;���|_ d@%�ʩ�<Z����yeP�$�{��b{.��� "��Ei�8��#
v7z�]�[Yk��Mɲ^^뿐P�7=�!?�H=�
z�����;>����+!ƽԁ�L���ǖHz�r��(��X�f���^�bΚ�Գk�y1?�f�K�E���.ӳ^��=��e�}w_s����{d�t|ֽ.��:�D�@ �_4������)O>c{M�  ƾ�[�]�;�U蹀��S���E֭�V��WHy0)��zu�ù�[U0�y��'��M&c�s/�İK�j����G:@���m
�#��<��c]�_�/`�@4i{S������ 	5�ʸB�<��U�e�mݭ�~��~v��3�3	̀�NP�;۵�Z����S��0��R��{����r��H�Y1�C�d��+h�,�5���#�Ľ�6�w����0.�Pm����}Jފ+�CK��+߂����#�'[�T����J&>��_K\��}������Ň����C��-��K(b�"q�M2	���VI�(6��Ļ���
_��cqa���CEg�SĽKuLL�r��UD}�,�թ/\ZXz|��K������"��RC\|#%C�if���X�bc}���)�I�]H��=*��Pz%6����d��+7�[b��Դ���W��y;����3cx4"��>-�~$�B���o�QŐr�����Y�ݨ��;<���� �}�
�f%��Ǵe��f� E]�D,=*@�X���?�y$Cf�*�K��0x~&�����aG}a|�.�!,8[X��X�D�ߍ������)�庾�Rs���C��-�zIÍ��WRhKN_���^ �gGS����8�qG,����r�t_�/�0�6g\x5l��ܹ�$?��A�8���t1Rc��"7����=� �/PA��цg��:����j!��Lά�IA��ې]����(�������5�Y]�m�.x,}���]F6�>(��dM��,6�*Ш����c���� ��BY����.�{y��P��g���绣i��Ad3�Hb�n���,����"Ԣ!t!Y|�`����~Uj¬�(��G��n��XMg�6�Ǹ��ک�KH�� J{�fT�hW����V�6 ��
�H���g8d���1u؇�4^�ȁr�$ሔ%�]EL�aDݐ�G�����"V쁀���F<�+}�]���"�.�/�& .��z7����#��]�O4q�����U�D�3�e��7�XF<��	�L1
�C/��=b��Y�D�)��B�t�h�u�gM��=W<��V��A��Bb�������N7�:���1�"C����ꙙ�L��p�e�=�@1�=/��8=�4A���ގ�c����F�R_�E3,���t��Gku���薍!~�{y �0R/7\�z�d�b:��ݬ��u���H���_����0.;y�w:gNb�g��Q`<�>�����C�@�g��=yܩ�nBK��{�Q_hS�oJTsŠ����ڦz���7}��`_��.��S����|����d�K-Ξ�nv��`]����+��kjQ}�-�bջ���>-I)F�q���?���m~G��?�>`u^`�tS2kt��=�5�O�"�jf �Y�3�Tx}�"��a*`�퐹� ���9M��>jnnA��̘���&Q����52n�j�oy��IMn�S��1���6�G���v2�i2ޜ��d@���w��̾k���	��(�w�\=���EwZr+&�#na"�Xe}��6W^Z�!g�"f�U�o�4v�~+E"v�=��4J����	�|o�~�Gok�htܾ{���� �gI��3
̍�|f��!9��_�@��֙�7�?�I������iqh��~�#���$�r�֭;�kZ�>b�0��Ѧ=#��
���Zur�z4'�F�H�>KD�0�DoUU;P�[�!:,M����k�m�������Q�J�Q�
u�ן<�X}-�AT��u9'����;�4��K�8�^`�$����l�)z+�h%o��z�r�䍤>�M�vZ#DUc>>5���������e ������W�1�F�>10�#\��P<%Fo,�����j9��Ћq��?������e.|#��^����2�!D�*��o������,ӍV�ea��*���7!z6�4?�5���N<�|��WpE���K�{L���mG�?N�UD�
��&е[^�����jL%@ �ѡ �k��M$Ѧ@��8�NRWQ^��t����jcl���l]G�$�^��#'�����F� ]ZO��C����x��E�(�H�̓���� �#�%^ ��~2��V�Z�S�;�*�͞�;�{���I ��������(�/Z(���61ljo1{�{��S;���¬���0�8������B�$״,1�YƳ�F�RB%���J)o �Z�GZ��: �S�-��?�+[u�y\�����_� �w�?�<�h4�u	� >[>�)�qS���l ��5I�`vRz{h�;�
���7^Y���ѣ^�5LM���S����xg��|R�p��C�#'�������s`B=���=Ц:���Sa4�"�&7��5BQ������*i%�޴��%%v���x �鬦�.M�B�N)d:�'_�N?�	�jv[��[�消��Y�˕�{uuq؁,��3�H���V��(�~���4������&Oba����>a*�C_oP�i:~b��=o��n|TJwE
k�֯�*�!����R<�o��䄩L����wj�|���ɧ��f5Q#M�pNʄ��?)�a*@�<���K�`�?A�jQ����ɡ#*��HB<+���,�A�ޞ�L�}Y���6v�83c��|&9+1m��Yp�}�c<��M$R�F��,8���]����z�):����s�k��`,��ܰ׏����D\�F	�`�$������z��C5�S�8����S��ҹ'1��pW@���q�zz�2��D��C>~--]��HF�>3�yu��Ǜ=��q�]��
u��Q噔f��FR��+�W�X�qow~ӠZfA��N���K(/��:k��_Hm9*�IÂ���ůs�2����=�R��-�m�`�2��?���>���G��ȣ���5٭_�\a`"S��B-T���u�],G���LY$N�����fi!NOl����T��������R�(�®�	+]"�
!}��f$q���Pr��zzv��&N�uu>�.��\�{�ZMk���Z��.�f��M���B��վ�|����-���Z����b1��C@�@�aڋ��������)�ﯙۻ0��?b�`�@lt�F���ӼGQ(�!�:�v2��O���Ρ@HwQ���VJߴ/���Qa!�Nk�-����ĺw:���6���g}[,���xcOd��9	��.vr(jb�G��p�,�
)�ce���K���nt**�=��z~��pD���!wg�!a�H�ʔ���t�=?m�*r ����j�0)��\� /��1�z�5{<Xj$��EΣ�����Oiդ��Q�8�I�9��$���ɰgG�%���B��~Ы���7RL69��û�sB�/f�I̹�S~x�c��������?�P�p0?yn�-�V�P3���܂�p��W�0�W�f\��DF�j@5�ɳ��2h�Q8饌�;j$H�ws�v"����I Ɛ2՗!�mD����ӌ6 ��c�YXL�����x�����YV��	����Y1���n� R�[�kG���Y=w���+�_Q��+�3��.g�sR��2@��~�%:�A��q��ά���_U^�Z^!RP��&��).�����S�R#a_n�K^��6g������N�S�E,һ�j�t�]���z�g�K�l�(P�u`��C�A-�{���t�#}ª��h�����/���A|e�;�T¬�<�
/�0m��L�4��0��{tJ�]�(Y
��`���u+����m�J�,pH���,6�6�(���M�C�̉kʗR�H�{c;��������AǕ3Fƴz�ψ��P�E��Hm��[s)�43-�T����̊υ[U�B)�!�w�`�K�*��jb��ȇ���n3�4M�B6,cp��%��aOU�{3Ұ��@�c�4����6��r���HIXg�5_� 1X���ѽhip�ļC��)1]��,��ŐN�#��"�$�� ���k�h��l�]^}�"-�*/-rA.9��7�9m����Sy�O� 	��A�_MMD��e9ny7��<i� ������^��a/�|�#D0���;�x��^�����+��&��y�V�!��bE���,[��۞cJj��󫰆����y�W�r�9!�녿�pFn=p����>'��@�Ը��mJx0�y���~����R��;3̧��k"��]�4Ԗ-�ʟ�� r�R�$��ɞd�'>�x�}Xm�� ���d����O_�0��yu��:�ŬޥQ �Y>f�_���S\�g�C�y|-��:�KB�+��SfãT�$����z�4̯7'`�0�έ(S��iؔ���I&dfOe-nb�n�`�&��c���6Qǌ����<N~-�s������T��Y\����P|���1ne�W�kz���5b/�*HuY#o��'���LâB5O��4� �'����&Bn]Ͼ	�
X&�Q�q�O2Ź��ȼ��n:�_S��G�Q�
�����~)iҝa�8��@S����^��s�{�Ș���(�혥QZL��5R"vo Z��z�Z�2mg���ffU�on(���"nq�ݍ�4�oOӖA�|���M-oht|�G�f� �TI���
leu|�M!�'�YI���Ha�9�`7WOzIW��C9��k��^R#)Xt$0��Mw*��q�ޥo"6�0� ��F��#:1�����u�\4��c��a�>���0l�U�Z����!ڳO�YUkm]��3��¶%���:Ϊ4��?��XUs��o	��/�/�;�,G���K�g�����b4�)�hŞ�����rF�H�-0����v��U��9>�FI�_~z�l���L�� �5�+j��ą��F>�+I#�gP܈o�x4����9+(ً��) �V�}��Ye�d�}���Ký�#*U�ɉ`�w�3J�-�eC�*1 �7�,6_�?�����6���W�����ƣ�nL�r�m�"�?��"D�1z�=���UK�K�mڐ�1Lŋ��qa?����K����=�H�ڸ^8��럃%j�K�r��%��=��\S¸I����b� ��'�-���x.X
EY����#��ȭ �O�%��Ԓ�.�V^}ZpO�;^���>]P�bT��˦����2�(jזZ�;���=l
s���ɴ�����z����^���T�8V�Q�XT`BK<s��<Yf3�F��R%�l!\&%o�Nҁ�G�ڷ3S��p���[\���(M\�,O� '[n?q��h�Hx	D��[�?�ଘ����l�=W5�v�q�hZ'���o7�W��Y���£H���S5�p��u��� g�TpI�����E�'__gԟqs z�J�B=pF�����Z%a�ז�Ʀ��ե��u�D�2�ʨ��~�B���vG���0_�L�p.�P~��:,W��ĩ��v��[m�Ոt�N�k����!qxZß��H��r`2���R��t��rЉD1��2Rb�^��ƪ*G���	�b@<Bo��On�w���v�{*o="�WHb<�yq۲��I���\Eew
h9|\�^�G����*Q�pS�Ʉ+2)�an� �H�ޢ�%?��Q"�o#�U�����+8Eh, Iy�>���ɂ�1��MZ8�.z�f�+Ѡ ��}�=v<aó�UF'kU8)G.]S���ڦ)����ZS�s�_�n�z�&�/��֐Ķ��|e`�v�j����l�+�C�b���y�����%��rA�1+�lp�/u� U�zV$삐ڑ��$~���]G�\FnZ̧`�g��ai����
ɓ�8����F�2+>��X_�Ww�����A1���r��Ȗn�&��i/pm�BL���ܠ8ϧ�O�2������l�ݤ����m���2%�m?'_�>u�GXM�CU���t�_�lt &ȫg�BT�-pu�=~GMeqL�k��~*ط�!���┭aTJ��������ŵ�����8�!��f�(M�g�r�1;��w�\�q��ғ�p)������I�jT������X�jM2�r�6D�^9����|-�p�������V|b�S�C�*�����?٧��¦ɯ��9�0R\b��	���@tU
$j)��|V��v.��(���9B�<@��K�+�J�����Aa�`lN���-�GU`�w��ۉB:�Ζ�[��Aڽ��c��d#���S���%�(
cG��9p�8C���c53�2�����t�y�=T�~�`p�歹�A��aM�X�4 I��cq=�P����f)+�*�����P�����/�~H�x{�Oc$�q�EnP�VO;iu`k��CM���˲ْO$)em�Pg��w%��DJ~pi�bR���6�-�[/B:φ˽�6�Y�~�s�c?F���4V�ߙ����y�C����Pӏ9��1�"�ݥ��f��vG��a��%�j���S��2Jj�绥,]dj�_�w�~�v�(�Lg[ ���2�����EDP�����֫����K�k�,H��t<��@Y�d0�`E�@�1UѲW"���A����+G[x�Y�������+[K��&�537�4 :h���r��t��z?@�T���P�3X佸a�r��~�D�1X��4NS��@֥�e����)�:1�q�K�G{�WJ����.}��dI��fJ&�}��hʅ��j�Y~���o�KC��u�����k�rp�9,��xA��(;�ޕ������>��X>�e���N�������R���F��L���� 1���	Nlk3pI�`ҝ��,J�O�eI'�*�)f� `���#�Tu��ǶE�Ψ)�;���z)�f&& H:��*��U�\�*M�'��&Ts/���|6��+}CG���o���݊<���]��\/q`&4���<e
�2��	�-?�iC-<�'�F|�~+���o��ύs����	]��N|ۆ_�Z�$������斣��T/\� "�1w�������?M�� ��*/	��H���>5R�9��v�iR;�V��C5�3�?m4�����֒�LcI]����k�\�l�KNj?C���0-��O9��x��3P��kl���I����|4�(E���l�x4}R�ƀ�
���i�>�糢�E�a
^�{�=D�n*�(�%�U#
7�F��s��®,DH]M��O�$6�qV�9��m��E�}E�,Nl��SؾLܨ�J::�٩W��AU���(>(@�OJ���̻!�I�a��R�kQ��ړ����0�E|#��a�Ӎ3XK$�%��*������B�Ð�C�r����Si�:	�9Xy����r�`���~�j݇��`G�:A�q�k&�L;)�
6�ߵ�.ˇ(�\�<���)�\�eai�"x8�����9K��&��9t��!�O�Pa�J����38���!�;v|�< hS�@���a�` ��;^-H] ���hM;�%�	�ݍ��cL�mV�J�V��KH���m/_��xk�9��]�|���(}6h�"cg����|}��TSSp�Ƣ��4�J��lS��w�r�E�c�qQ���܇Am�I�{���&1�Ⲫ�L�,�וּ�?q1m�m�V�FY��{��}h:ժ�ע�1ҵ��>F�fmVT�;��h�[������NQ]s2� V�(8w/������}�����2�[Ջ+�Bb�8��
`�}�C�;}ڴ�B-�O1y�N�s�W&��ӳ�
h��ol�GV���d�x���W+�H\�!]� {�蛳,1TM��T�dtca	/���5�e�ξ[�}�A=1��v�>'�DՂ-���@B]���0���HЂ�-�B:Zܨw�A!u��D��/�]QA�E���*�&t��,�=X�����	��r�A<S���쒪�����ʶu훿g��@Bl�r�k)�=O��#��a>]�}g�T������D�\P,�m��Z�k��q��^��n=��&gX�.�c���.�kkf��m�sGitC��&��3��8���W]{P�C6!� ss�-���������>tMJ�͎v/��a�1#�k�1̎�&-���&+E�%���}���<UՔ8�F��8��G]Gu0ʎD)Ϊ#��*os��\�$�n�ף5քdN�Z�`���������v���C�)��,�'�!�g�m�fb%1�՗p�]��A�z�:��i����~%�L];�_F��)��k��?�U���q��
	��es���<#FfS�+2yX��bw��5�n3�A%�9��9���D�q��]y�mM�ήݑ���D��C7�2F\���Z�Q���s�+m��2�?�9>i��G�#��7�0�I�{_��t�[�-T�uy�$G�o�L�����ث{!b��`T�����]��f5�ũ����R�!� �f��� ��r�%C�� ~�PoF���?��>2�p=@��K������m����M��ָe�����Z,*�-��՚�U��|bE��C�`>�u�5�3���F�������0F�b%p�����t�2�^`,�[��ݵ:i�����v5�y�@܄o��F6Jsw���!a��UN�-��/�C�w�艶�Ί~�[@v�ڱc(�;dѵk���+(~��G���p�O��Ucy2��l�!��t�3$=�р~�g�p�;��ծ{�OaA1�ʨ�����=S}����B4�r2��V��e<�p��/��܎�9{о�$�Eb�8�b�J	i�G�|��Lo��͵ $��B�D��9&a����~�"J�Vܖ�Kޝ6�R���XB.3��1���M$~ ��c3����0���$�؄�-y���j�|P�t4����-�F�ĵ-�z����jTSi�G�	2|�Z����j�R�w!Иv��(�� ���2,�㗵*UDħ��tK�J1��~��m�� I�ь�,��4Yj1���t���71I�$�����8�o�-GO:�YQ����~+�8�':3�0U4���x���
��.nf@lv��֠�3�23�U鑅h:�D�[���NG\@J�
e��bҝ�1�B���8{�5Y^_��"������Z���s�hO�W�=�M�i@K"����e��0�f�D9���xe��,���(��;����^f��\�e��yNkI���Ӻ���@�WQ�>rBw������
S�Nw+�3d�:`F
`x'ר�<�I2⛝�S T���3�ˬI�uH�v�98Q�������:W�5���_s]2�h�u��~:�$VG ��FotO�3������hgV�{B���f>\�e�}�O:T�Q�##S��[-)���|��\3Ķ����=�B�a�����He)��9n4dl��zC	�W������{�$Rk�����3��؅��FIߗ����HUo/-��H��O=���9�5^������j�w�KF�<�('�Gi������^���8�)j�����m|N��U�xh��s���	��CxW	�H^^�bP�R��Ěc�i�3sVٟ5p��%�8.�� �6�2cm�I�7�k�M�l�a�	�U�v0Q�O��~x��-�~�k�Ԏ��a�^`|���E#���n�xX�H�j�T
y�i�p�)�x�F�E6��
�����#�&�?��A�y��7�%9��$��6,h07MP�%s[$�&�qz(S�..�?�ź!�,r8TѺ�ӾpA��CL����D��MD>�c��,�XJ,��������$��t�k�i���Ϊ�7�z�i���z�ӱBfX��&%6���`�����1�s���;r#r���(:-���o��ԋr,����~LK҇���5:eo���L_��.��]ĵ�sX�L^������MGmo�a���"hF���>9�&2�L��U�O��a������
3\�#�H.;�G<�-3�d]��gH n�H����{;C�"��'k��C�LY����<VcV�H癳m�3ڜ��9�<������'a�����"����&� �p�x�]py�����a�4�`S1�����FY !l�V2�A��a���JT_��:R�pš��]�c��m;'�V�4[�Q.�ɡo;�������6��7��
�"Vxc�;�/�h�FЇ<�N�Q<o�D3�(�����:���f�}3e&��h��V��/X
B�����
�F��s�}�g�B���OU�DNeKWJ���w��
�#o�zZm�#~�d�h4����WOh1\=�V�D���?ZH1x�)�`4kd�7�	�������	�ݾ�nZLW1�Nlv�������r�=������&��vc�Ц�����l E߹�A����z	{](_��d�R�&�o6��=��Ǫߵ	;F�r�3KS�����&�KN��>���˿��@��r�A�׸�ʄ/��#�o�̅���!�]�x�?ē�-h��P������Z���/"�q,�z^��=H�A&��H��h�<7���{k�I�=��s6�t�S/&�GEע�8$�W{�ga!:��s�i������Q��E�Mn(������m{�8{���q1�-ښ^»؎M	�6_�TlZ>�'=Y����`�r�?���TY��XX�4���U.�'��,ZWmy�h޸�\!##�e�47b�� cƗ�����=������2��FuL��y#R�۟���}��Rf]s����h��[��>�^���E��.(`i&-O��욎e�3������Dԯ幢z��ٗ�9B�fA#y�v���uz��&�����҃+�^$r�B�&̧YUIT�&:����4f���0��r�������} A/�i�=�*�Nߜ���A��.�aCg%��o�W˾i��î��0;�K	�f��Cy.�D�Z��%"����?g2'�#�P��o�2hoC�����|�
�TÒ�i�^o�nPt�mu�⋒�An�A�q�N���4�?��Z�[����֟����ix�;��-R-�����[M�<4��%�#E���6�Ir�X�!�э�C�*&��bשY���u��
^M�;����li(
�-����"#�{�¯ά��^iyC��p�����re�=��Y�;1��-�0TF�57�[�dB��B���ݍ�J�	���9��1�	�k�a�J��iW��oVK��_��R��	���w�@�$e~��oFl�3����_~�dM�V�U���q�&9���4E�l�b������ݡ���^�'~�9��>~�
萕�O��|�C����I�����)Y���� eI����u}�[�"��eў�$dM��# �.��� #) 	߈������'�V��B����rrG%�̆��k�Y�ϸy5�/�4�
�VY�ߘ&�P�4<E���A�Ĺf�N���4�=n Z����x�#L�&�-%�c�2@�'��7����jn,��S�Ѱ��/����,���i����g@�Y	�S̐�9��rO�z,F��27���Z�͙�uRI"h�IO��H�Z^X'g���f��_o��+��A�"���4\�S�H�H|�H>�P�o}Z2t.v�X� �RI�ӕ
�X|�	�!��ˍ�V�+��7���I������i���#��N$�5�?r�=��P%�ԣ�0�DY�x3�#���3�wuY34�M�Z3t>��0^�U'C�mk!�<D�K��k������/�h����y���(ױ|X�o������GX䜡�5;;P\��}�}�T�6���f)*	h�?��er�eW��o�}[vlG�Ua	0>�[��1���ڌ��� �1��'��$G���!>�~#.�8PN�o~R�����9]6��y�����oZM��|ne@=�/B��=�W��CP*����q򞾂�_��esRl*���7���6�ɦ?�!V�=�"�ܥW�YW?W����L��*mg�?`�
DkJ[�/��ЇXX��9�B�sL��񣷐�}�m�������2
h�d��^�I&둭�j54������a������T��<�ט�� ��s��|����3x�&�EK)'�͕0�2�� �L%0,Ȓ�ؓ���Zb��;��SͰX���ˠ��k������XQ(ʄZ��I�yrl|��p����X��%˓���8�1�E��o�8�<L���B��𴾀5Y���F��b%N�2NYo�ك�Y�*ƌ�tS�����	[�\\UJ�_�^�8 ��?#F&h�0�	v�s[P��^Ӊ��e�l��L5[��v���hL����g��ɉhYo�����0{�5^X��'���SJq*��N�j6/��zA'�2i��Us��<>s=�b�.{hK�a��Ƞ��Z�G1��'��6���m����lO@v9c �J'5龇.�ܮ���P:^G��`Y��[��v�[�� ��ڧ˧�Uwq�Sj�@�HM��R����m���S*ކ"}�{�L����bs���E��*9[A2ŝ{�b�}mo�b�nN��wW�L�(��*a^����8<��dVy�;Iz����w|�p|#��9�R��Q5��Kք;�)��*R�P����ޔ��?��Q�i�!�6#�Cܢ��+�w,��Y�0{��O>��.��8����N$+C%��*�}}�?<�J�6��Fن
8ن]�YZʌ�k)��W�L� s��:	ļ�,�M�!��¦?�X�
`W�g�\ψ�����<�C������W�e�x�$
�1u�p)�𹒸�z�'��t�4��~#��]�%�F`�KԖ��Ԝ��/���
G(X�cW3����F�.�+phdXќ�wb!��Ac�4��;�z�����"�mK�-����*MEŁO�2f��B�����۱�mpq2�͗?�W>�f�G�a������me_ʃr#B�f�T�O_u��QG�˰L��p����>�!`B��F�T<���ɏ��d�O�gp������s�!�i�fv�{�-�r�\������`ѓ ���n�s߬^���篝��#���[M$��[��~�ε<���-�Ԛ]�h�>b�f�C���s������娦�i;���~0"ab�ٰ�k�t��A��ي���BD�������4�*@|���%�J16��ss5a�>�NC*-Fz�G��wo����,�H�[��G��ֲc&��d՜g���� �T(|�Ggi	p��ܪ�cw}m�f���܌t�D�=�
=~p��p�E��U+y5\a��X�&�E��@=Q�|�4XQ��PR��r�����/�m�܌M�{�ӓ$�k�E�;z�&�\�ig���D��J�����$1:ɂ�x�7U���k~b|�ߔe��I��6��X�M�9Bl+��/�`��~���cqk\�������%�l�y@I��h�@P�RV����T�5�+���B���	����jR�r�N:2�4Z#1�����jv�Lw���v��r�?� q��2����+�D����p���ȑ���'�k������
��8.Yhx�V�B�2��1��ɞ��RL����G���YO`*�=�n+M��XS>3���4����$j�Q���M,�u@��+'3�8��0��D�\��N܉@���eөқ
?1|2��=�2{��\���FY�VIHޘH��h�_��-n��E,�g{KÞT�g��I����$Ut9 �xK����'����!��l}��`#�ʦUe�T�N�
a��Ċ���`�⓼����ț�뼜ȺbN���3�F�`DA>6>|�A+�IY�'��rQ #x�B�U�uF碶�,�C9�� Z:UG`�b������s]u�i7:��G~�F��:O��cН�qwg�ZQ}�B��\w.L}EZ�OQT۸l�����;#)�9�:,x\�*�����;�h����TF��m�)��
n��V���z��O�sONP�H���b�/����~{	{��9���K��j�U��Q����XTZ����5�KŢ~�4�iGj�
K�l�&N�p��.�1Nw��:78��&j|�/�$|�k��S������n/��	�2�H�Y��`��RU|	�~di4��V�F5.Í0O����K���(.c�m���\k��lE1?�P�Oc0Oh�O�Fvx@@2��k�¥�^qV����|�E!���,u�x֑e��)
��i��ҧ�׳�d�E4l�
�O�n�&�$񾠊r���:7��^����ZO�,�`�M��-q�$�n�q�g��l;��=ϕ��X,����A?�n�희i�{�����|�ĂB>g8�˪k�Jj�;�ԫ��?�k3UĘ�!��5/�����wӯ�X��R%��s�>h��8F�n��e��%;�r!�2ѵ^:�[�-w��c�r�6��:�~�a���y�8�:���M�|L]���lN��EBF����JZ�� ��:)�h�a��i"ڒ��7e�9-i)&0��/)�6I%O���a��ۦI�P3ڮ*��^�;�U�<�e���C�C�� u$��(H����g�;A�2�k=��?L���cV!�He�7m /ښH�9\0x�bT�����4ڄ���{���^ ��v2�p7�t�><��2J~S�d��)@��M�2.���AKO�]���H�T�D����8�ѳՎaTRm��Vbz?��#7ɟG�� �y��W��#!���MV�F8;Ă9h�0��
����=Q?���B=#(�B��:����_}1>�Ca(�� `�mxXB��-�rY
fQ�%��}�^�B���O�3`N���WH�B�5�

�6oN_xo=��2adT�]�üWM��\��ѩ�8��}%1v�E��d"�	��.�%��Ǚ�����u�1��v^�^����;�W<�y���BФgf�0�~k��#8[���8��]��������1&�v�pe=:��ݑN	���rUAS�Nj�ɢߪ	Y̷���W�G���@�G�rE����x1�-�&#DXt����_Ď�vǒ�Q��,P�6���Zi�k̭�qj3�^ǋ=~z&	e��c��:<�ސ -kY��{N�s4D�t�'�&m�9^d8G�W�����j!x��s����F��Ł:@� _�Mli?���4����v���q����)�oM@{���҂|�;';���K���2�?��R��u�4#>�Ul_n'�e,�yy,���L!���#T4���^�Qƕ�L��^��^�����0��F3%n����RX�۝��;���e�s�|���?οI輁d�<���T�`�N.-�M������1}��J���� �#v�z�`0�UQ�BL��#�H/���CzN
��yz^����\��Ѯ�B ���^�T�Wr�X)3��zn��-F�b7�N�|rb �&i���*N}ɜ,�$A���.�������o�SWQ��i���E��;W����rCw�DB����F�%�=�'D1P�(�p�PC���ȳ��nTTXg�0^-dPP�`�u?܌≊�A,�5�����Ƕ���>��'���)���=x����N�j���[d�ܼ%��`��A����fI��_�_ы�*�舎�����Րuag!^�y$���j�i�4��&��"aM4�����t ^�ZC�<�p��Џ��f���Y��ٻ�0����<����F����?2�������RJ��s�r>`3>�G��_p�JSٜW*�V�A9_�7�3��w���$c��-�l!��1��_|d�)�Ӷ%�eR9�Au���%lk��[����P�_��Ɩۍ'R�Q9���~��f�R��zv�BAƚ���/�'���<o ��,�)��{�x��u�eOX#$�6�!1a.B�� �q�E�ز,��)��z�GN[8��\�=��{�"B�m8��`lYH\U�z�w����L�H��+��� �n��I��D�̑<W'�Xpn��bbm��2[@y�Df��E���.�Jv��H�e�s�"�s��)�4{�n�|���.�}�*@š�_Ӯ͈z�Y)���{��� W�Za�a�U��͖t\�� b"�4g&�yOi5�y��ØE�U�oƒ'w��&�r]/B��jv(�ٺbGs����Ɠ�d<P#]:�k/��4����p���b�	��Q�Wؕ<jZ|� ά�ƭ���}g���	��{N���4`�Z6;I�<�F�,(�Q;Y{�y��y_Ǎ�����+��-��Y]h�� 5����ǖ���E���/w
����E�J�(+i����E�W�Nr#���������J%k��,\c�p�4n�[h��|���*���|���(A�Nq�P2��3�o�II��6Ν9�+����_�aq Y�1�rCĹ�²��KF�2L��T0��E,P+{/�iVX����;K����뗚����\[�%:�f)קXo3�}]���h��I��Ʋ�5w��Hf%��Z�Э��
.��1e�T������(����Ę�c�p?�`-=���T7�AQ��(�Q��پ]ښ|r.)9(�M�'�_K�}��f$)lǓ���%tZ�U���8�*�%O���	��TRf�^�Kؔ�x=V%�R�E��b�a�/�`>8z7�M��#��׏SΫ���>T��9yR��f�b����Y�0���wR�g_M(^_��g���5V[���r,>�p�i't�:_���Ng��Xl�l�Ԕ����AL�K���t�X�˨aj����S/�.�A�����W3}�����+�/�Ϋ���(������\�(84��32���xV�m�K=,\�\�o�6���(~^MF��k�Ix�����cz���ߟ6����t;(�s~��'s+P5���L�>��S8$3,!��"���f�$n��''!XF�`�吩Iăja�ܧmŁ�knҚ�M��J6� z�ԎƩ����M8{'��݂����5�T6�w���Hh��g�y����1ԗ��s	�	�#X�1�]�w�� ���-&���Hy"��h������L��
C�]}F",�/.�i79Ϡ�B���PO�g�؎"�^>�Dm0e��7q<��KU �"Ӏ�]q�{q�D��vZֳ|o���Ԟf H�jP�$�V���a�/bw���}��+�=��������� �6���:��$�pŒ�=��� ���I���~�L��]b�.Bt�e\rR^�3XŊ���>��BU��Xs���� �PR.&���HKdΎz=B�\`���h�����~�]�a�0�k�y��:�-���Q�Q >���|�M�g�`Uy��,���K!+�ʰc9S <T�]���{���S@C7!`�(���SFJ���ɥ��d�
-���n��`܍��k�_�7�Q���a�0�{�J-_������eo�P���{�N���rTǻ�3��k���;5!(a�U�T�Y���3P'��|� v�.����'����B�nm�2������&��s�Pũ2�CX���6�h�n���Sʪu�p*��L����i�kv��To@�LRvb̝����!��yc��)��W»Z�3��B~�"�l\\d��fjZ���grjf%�#or��"u�d���4	2ӕ@�|�y���o�z�t�,S���~ ��I�B
k�|�ק!�1�����_�.֘��7� {Iv�
�BVX�D)�Y��#�Ȕ$�>6֬�)�J^S��M�!�0}L�9	#��[� I�uq�]4R���>�6�0K��U�Q��q!YV��G�k��o�R��µ�W���iz���XX��@Q��T��N�n;�����\D
S��c+����)y�h{���#rE���*��vev�r�U.��>4H��)Q��ԡ��ԃ�I3V^�QO4�e��>0��#;}XP�J.o�~m�t~�9�k�J^�����>g����e��8�|k_�*Rx���z*������
��<�l�e c�*0$17��6�? �X�
By�{��W��d����!+Lz�em��?�=D8L�����Д�jZ�ڏ�L�W�01ު+�lu��?I���^7g�~t>j�؂�J��]?�#�V����h����¨ �E��>^��+��x���E���'�BJ�� zW%�J3���b�մ1Z�u>;���]���=��	��B7��%�(�<�Z'Qп��l)\���Դ��Aղc|�&Q4��Ҷ�/YW8�S��w�BJؾ��X�Y%�hF,VH%����o��h������Snd�Ҟ�#[��r\"4��/e�k} FQ9?pN�h�B�	�	[}-t�+:���l�:j5��v�h9���i�����YY<{�	j�=��5�O�t�@pX�:��]�7��B��'��rԾt�s��)'�=/i|055)�a3vY����W��t�i#����7����9�hv�T�Wi��k�.���͹�:�ǿÍ��(�tvZv7[�������j�A��Pq7[�>��H������*��=� ���hG�����b����ѵ*�FN��(�rb?n�o�\n���w�#����*Άv���?<Ė�۱C&�(�ĥBiw���|��Tɦ���LQ�<�6��
o�)^��"��C����? ��QAK�n�#�I��|�+�7�,���ޝ���\�K�P=�ջ�8�\R��O�+p�xm}�B`<�t��.�F&h�8�I]�~ʹ*)YV8��GsΛJ����y����)�OL�߅�u`$�=�ɥ&����9b1C�}��^x�Mߒ�*���}1�h�p6N��?;�z ��az���#~P�]�\F�<�X�ǹ����`� ���
Ԅӓ�E��TkFQ\+}C%X~ٓw�݄�ٹ�A�Q֓�GFE�5�����m�5���Qm�C�&�2C��>�<3�۾�8m�f�2$��?�>4zxG��]��"#�4�_ו	w�f/�TwB�uD��G�-�LxH;��}j��0!�⓱T)[�V��]�4���b� �!<w�fûA�Z?rp�������ۨe�t;F�����Ƥq��t���"x��tM��!���}F�s��M-{]m�<3��5o;b0|C_w� ���>[^�m�麗�b�؂�0�:ob���ttu�i�c��+�݀篵��n@��	@'���J�J~꯼`��a{:�NC��-���U�wi��a4Ε̬[���|cS%Kd�,�8���()~�G��px4@i Oc��^�3�+��dt	�j=s ��	�p�����+�By�1�2;�K�w{�Xv��l�.��d���f�j�}^�h���e��YP���&K�n�u,���Q�r1|9,��x O��I	���:��)��ɿކX�|eϞ�N��8���T�R��Q��ʭy�;%� Ң�sNM�3pJ�`Ҿ��m>�OD�I'+3�)� `I=���#�u�I�E�s����)":�-���T����S�uC�:	�G���F{��O�Y���[�gb([��Ӑ{\���}_FO��=T))�tX�	��)��N�4\��������mzѶb����)8��n@&���?zO~�zn]���Ve��0m�ȟ9���A��f��Dkz���$�U����X�݉����R^5j!�<��j"�KRz�ݴ;��S��# x����0?8*��j�>��ls|�.����3�y��� ʼO�	���Hj����WR��_�&c�i%�V��y5|5->����C��B�c����t�kC,ml���a{�0��O��xN�O Hkt�����Z|�$,E�熆z:lx� �vz�
��i͸�ҵ���RluE�mN
�+k�DB�	a�؜���	7��7䅫�����,�+�M\	�iU$��q
"�:���,Ӻ-#A,�����\������ot����眣��R��>���˸�zJ8�B�|�p��w��M�k����G�C!���o����)�=��X��]%���l촭D�(�E�s4�0r�D����:�����C�?y�r8����~X4釣�����:�L5�H�L�q�뺃ʔS!񵨨��4���,����({�a/"(6�Er�9�&�=<��9�D-IO�2wa������3�靲T��;&��<�m������ �B�l�Hi��;ϼ=����MQjLeO*JbJVo�Hs��mߘ�(ێ9��,и��2�-�l�� �ao�,g��s�p�0k�L������!�S=.�"�e�w�!!��b��A��+�r��X�������Yӡ��6����mG��Vpr��]��-@H�H��&#����?n���CVm�;�jh5㺇H���Q��5@(�L?�H���F}������\��$�;��BSɡ��i
�p��F�}���B݊�O�nNq}�W�Q+؃�
��oQ[9�/��db����bW���\I5����KŔ1��l�~d$W|	�����ո�\I�Kf�1C�_v�,U������S��͇*������f~�2]��ײ�����kB���%�]���g�夂&$4!�/s=�ѪkL�	G�Grc�S����W���Wܦ���H�%п"�@���rSw��ľ�����#�I��k�-A��ğ����UP�(~��jZ�O̻	^q8�^���=T�x&�i�ބ��ȗ����k���I�s¶�t���&{���m8�PyW9��!F��s#�����1ŏ�3��\ M� �&�N��M�D8�5gjq="-�&�����M��B�x��UJ�{'Ƀ̨�Ye��
<?�ǵ���4�d�G41mU:p�'��l,fy�2-��WI�yJ�q�4��,���#����������A��F����}�R&�e�+]�܉_N���Es� ��}]����B��:u�
�$�t��`�-�݀�m��H6������*�>�znCN٣��BZ`�#��g�BP�z��������T����Q_B�t�e�
Tv*�B���ν�Ү������Aኌ) M��i,b�*�z�:�A�S�.�p!C�}�bW��i#������;e���rP�C��D�����K���n�#�'�qrPʖ�>ixC6��lʕ��T�9���^{5/P \Au9e���Azx����}���;`���f}��P!��8��{{�x�G�����^lڼ{�[Y�'�3�%��� ���Bu�I�C�-����x�6��"���eC&�vִu�y�^��J�����!��s�4��"/b\�Nξ���^��C�Ep�C���������Y��g�0`������ga����H�ͤg����ݙ�vJ1����C���8��wJ��QW&gMVW p_}QJ�ޜ�dw�G�$�f��{�l/oʍ�� _
ibdY秱��j�}�?9w?�@��lyj �&�G�ݭ/ƤK�' 59>8~��td��[��ٮ�V�ƨ���}ص\���ǭ ��<��c�	ZZ�.��e]$#$p���8�.�� ���E��?����w�@z�A([�8��h~�K�C�s��;����8�H���z��ߞ������+��B��n��c�E���5K}X>���Dtb�Yz�@�y^m
f�?E\.�β����w��j�s#g����{1E�|CH�.���U=@S�_!������)|&�{m~ mmD�hA���BU5ƴ���U�.�>�
��y�����f�UX9�f��'��&�y�/�� ��h#����G�03�+t_���<^�]ߒ/-74�yY���N�n�	�xʥ��<x�����:�����������M�	��N=��BO,Z,�ʲ��	i�_{{U�Ө`�
��;���ݽ�p����h�A5��7��<��*���d��c\�#����3^�J�J�+7n�5#Z��斏\�9�T+�!�h7��J3�ǯ�~�\�xm��k���Ŵ�~�fp~�<�D�+H�("�q/�_2 -Y�D�I%�6\�I�I��}Q_i��q���ƽCҼ<+JK��eL@Y&�b���a���/�TX����U�K���9���è\)7%�}�fw��X}�}+?���J=I:~\��kw@%��K������!��`����%�ȇ��&�ce`�M�_-�YZ����Q�2
�a��L�h��q�7"���|���}��f2��alSٳo�2�r��O�*m1�M+�渕f�LxK�Dzx���������a�����W8�	J+iQ��b�e�V��0<�L�����R@�F������'g��@��RU��_[��^-�}g�t `�,̞˷LGt�	�]��g)�0lY�=��:���k^A�Kt�U��j���5#�-�[/ʄ�A)��T��A�`�Ʉ�7D2�'�ι�����(X@��1�(F����w�g��Ƽ:m�{X,*�����m6�1(���M0[��X��L肵�cH��m��/Dǂ��A��ϵ�PRw_���y�hL����3z�2��c�Y"�ϲ�{���!f �`�ᇩ�9Zj�ѩܵ~�t��n`'�M��6�b��x��F����{ f����C������F�6�5���H�i�g%}~�H$1�����5�L�1������]`�B�N@��;���E�"#"]��:w�ؾ4����]I�"zǀ/�_.�T�7�Ҹ������O�G��fj_����D{'�e�s77�cQ<66v�Y#��b�E�_��,eD=6��=��A���}�t�����d\�V�E��o)
b�+��Y�@�y�b�к��qt�3���PY�DxY��ݐ��p!�=�i���y�Ņݤ!�H�ZƑ������X:Rl�[3ٟ��֊4���!m��׆�H�7 ?�>R<�I��~}d\~�O٬j�͢8=���̣ �C�0���y"��:T����0%Q���>�d�a�a�]qg�r�y)>�[`_K/��~��S�b�T�z������9�7jJ`�s[��S�Z��aޥ��fds��--"nc-p`�P��9����XQ�E�o)C�I��-����^�A��V<��<:貈]L�'OM"����ۧka(�Z5�������Y���7�o.�NY�<�r���ʦT��O�n{̇�˸��^I�&>�m�^@�2� ,�<Z����Yn�L�S�>g��7�42��Ii_6��ey�@ C��i�k� �	��B�� ��%{Z?Q����"��*������Z�=Vg�#�f�g�o�����|�"��V��!4�"��I�|��d���o8��tI-����Z �k0I-
�j�|�8v!f�5�g��,u֦��7dZI��;��Ӗ�'(�#VS�$��ֺ�û�:�oQo5�0�	r�ӗ�#g	Z�N��u#�4�g����i>8��0Yv-U����(�.\� r7:;yh+u6����<~\B;b�އ{̚��~k�c�)B�(�M��at���y����PPK�x{ܣl`�Z'D�o����*��R~j�ɔj_2i�"r����Ҩj���w���v���m�3  д2Gz�B��D���(���^�����[H�mL�y��s�Y���e썌!�v1VQMx�������\��G��Y~�A�Lpn+<��'|�3X'24Ao�Θˠ�����;-Y@��T���3y�������U-DDl�?0`N�@���e���J��1	7��P�{"������̐�E�p�g��瞁�h^��D�F�����\K����VdkL��3F�i�9��Ix�l��$&܂�Gi������dl�y$�e�NX� �D?��Mo�������Q�A�d�WNd/o3�xM`s��E@��0onI(�D�Jn ���� O%��Euu"���H�����!G:���`�`�Bd|u�c4:�7�GmW�F|�O@o��,��సg�)���r���9\f�N}95O��Tj������Ѻ)")��I�X\�j�����hͮ�����|�!)�Ռn�����zP:���1�Zo��-���AD�@���:\�����4��GK���U\~M+�*ei0�� 5k�/�-��H��j�c K�0�U��j���j� ;�Q.r8kU�j�y��[�|1�F�`������������	ͳH�A�����Rd��� i0V���5�j���1eYw�.��� Fc�&����kd�wl��y{i���i0~�nO���x/x��Dk=���Vz�[�|e�lEP�Ԇ;�ux�HR�w��
ǳ�i~�I��ȥEcZ�
���T��^�^����f��7D:��&���i��,��M]-� P�$'��qg����]�l;n��>,�:*���i��n�;˶��Xf��9��>vɍ˙J9�&ӝ���:�����Pk�5Y�+F�f}��L ��D�^N�X<wH%#����C����}{��Tb��	�r�n��D�:�D����Mr����j�~Y�}�Ġ8�:RT0��;3L��`�{[�4��tY�����-��:�a��a���"�>��&�L9�T�&��*K�� OF$a)�ЦX��3�[ݲU��;G��<���QQӒ�l I����H����;����鍮��L���	V0�lHT�,m�(��Ik�9먧���r�$��ζړ��jƲ�-h��%��p�u���9e�f�a�S�+��Ҳfo�B������A~Ӻ����w3ĊS�R��`ޡ�٢�4�m���V���ޘ���+��͛h~3��`B�W�Ve�,;׾h��_�	�Ѱu��Q✣�d()V���A��NK_}`��R��å��<��B3I��D�
q�
�t�p}+��B�}~O�WNr$W�؏��T�
yd)o�PN��޻�%dCX����W���\�#��1�����1�ժ�     i  �  �  [*  �5  A  WL  X  c  �n  �y  =�  M�  ߖ  0�  y�  ĩ  �  J�  ��  ��  B�  ��  �  w�  ��  G�  ��  ��  8�  � �	 J � t  �' ?. 
7 �> �F �L 7S 2V  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�=A!L&�S�ӰS�����<l༛L��5_�C�I
/y$Ցr�C	ʔ3d�O��"<yϓ|���q"��L��aрFF�1����`�^h�Q��hPN�}�d�ȓ!��x!D�<Tt
iz��ޭL�e��~��TbԀ�.͒��G+/���ȓr�]2)��ԭ��
�Vلȓz�<���!�P��fͬ3���(�����w���t,\�H���K�D��`���58�Y"���)A��=�����v}��B"���sΝ���l�{��ı;X�C���zC:T��'�J�x5��+s(T���	ف����ȓE��G���V󨤢�.�=x�i�ȓ�P��dC)'�l1�c��
Ѱ����`��C�
iv�@1
N ��Xpz��)k�<Bd
�>r���ȓ��
�h��l�R�ѻ�����)�J�0���Rn
顂�T/��A��L���S�)	�T\J�c��>�r��ȓ|6`IV�5^���Y4��E�P�ȓ�b�෠�3%�`��/@�J���NQ
\K�HJ'�]	��Fp/��� ���b�BA�;�:��L��K��@��}vMc��O'�=���4��9�ȓX,,����W�Δ[���L�&���T���'-JH
��ZT��,Z
�'	�p3Bl�v�`CRCς\Z�'��$B���q�(����"M����'���Z�Cq��%��K	=d���'�~�:�K
�gM+t"ݚ8�4����� �����H	��hT	�&`M�jY��HO?���<���K��ˉ�a�ʇ�<�!�.
��9����"�!�D��?�!�$ݨR)Ҙ��F�3\}� �)�i�!�d�%�����d�	�� ���/!�,��e�J���H�G��Y!�D��� 	҇��Q��U�Ɓ��B�!�
Xۄ0��݁�L5b��ՙ%�!��!��)�wI��'��L	"'_�z!�X�`�┥�6>��pQ#DG�!��͉să��w�e��ˤJ�!���6L\I*��n�����'JB!�ۂ�|�b�RS9��JC�s8Q��D�t���I��D�&�S EN	��n��ybh6S���HO#<����gR��~"�)ڧ
�~m��%��>��%�\\m��!�L��Yq����6ō��R��ȓ2�|�0s��+vS򹫑!<6J��ȓx�<y��'C9Y�D�3`Ν0{$�ȓs��MXIE=)�����*oHd��]�hX�Se�;�̵qEg��l��C�����8��1�e�^�F�dQ�ȓIȐ���C�k� 1ӱ�2(����u����呼	vzQ�jTl���ȓ>ܒ���!}[� �0�V�fxh4�ȓiw�0����)��0�%*D�|��ȓ*������J����\k<��ȓ1JX��i�,*����C�Ϩ���<2��(��6Q�6|�Gl,^�hx�ȓ�z�yqC�i�Eˡ��+���ȓ"�qy&��k������Q����[g(�(c�\�j�a��_6�M��A�Z���/t"@�A� 
�%�ȓN=�)�����jF.��+<@�ȓmTY�D)@)X�HARd��e��X�ȓ��u��%J�=��eb�K�N��Ćȓ������Ƅm�`�V� �Ƹ����i���Bvu`"Ԧ͖��X���ޱ0��:)VE�RR,HЅȓN��ra���R��hg�-n`(��F�D F�'`�,����G$�]��|�J�:���(��	>� �� ��"���*k56�MC��G{r�'��A��� W��9��J|HYY
�'F�z�*�*`Q9�%ARC6������x�,8/�V���L� W���c#%Ư�p=a5 9扡{�*`l�q��Ff�4��B�I�q�|���	,}�x�NU�b�E{J|juG�7`��H�G_�N(p�VL�<)Clə	d��)H�hlT�#��^�<���9)�����j4R��;֬v�<�ǒ���@R	��5�(�Cd�L�<�G���;��@��"ƪx�Z ��AF�<�0�X�%jFL��r��	p��B�<9�˙9[�$8dOH'��X!����<���)4���� �;j�ny�g�x�<���\0(}�1K�-�<�*�LWq�'@axb�H��H�2$�k��\�j�<�y"�.m��A6. ]�P�s"���y�N�61��#c�V�AB��y�Ά5xr�A��W�Trt����y����0h�J��R�P�^�21�ʂ�y��ۨ1*��I�I����ע�y�n��P9,]P��4Bfh��ɣ�y���� ؍��C�W�rAWF,|��Q
��'ԉ'W���\;����R��7x�Z�Q�'V����y�e�"�J=��
�{2��L����$��f����`�ѰZ���"O|�P���9Ct���
'� D����O�㟐&�L�,�GG��#�kA/(Ѭ�*7g)4���`��.f�Q�&)V/\=��h]n%!�$P~�i��M3LWF��4�Y0w-�y��I 
��A���`)�ep�!P�mښC�ɛ9(R(ɰ��S!~��M
�dC�ɏ"��Y�h��:�(兌!K��C�	�}!H�K�G���&���L�L�*B�0g2H5����h�6h{$B�&c�B�	�:X����3V��=�a̳.�DB䉜_��V�pU^@�vE�1�.B��(8�U �"��21\���N��r���d*�Ĺ�
�-�������SVν	bi:\Odc�@���*�`��7O�v��"�%D�����
囗b�4�M��N�40Q��>��ŌÊ)j�G�4.:%o%D���D�R����+�e��6���)s�!D���N�1:����}]��D�%D�p�ǡ��Ez�����]�1D�H�Ç���L���'o�����k"D���CĘN�p�kD�%~�Ci?D�t -��H�t��"��]U��aE�)D�|�Ѓ�.�qIW��TeU�2D��Ņ_���1�M�-�)�Af/D���4eտ;���r�g�Si(�K4�:D��s��/a��I��zl��m9D���榇�2͒�
1�P�C��<D�l��d�f h�hN�FI,m�Q*O:,P3�>0���(��'��x"O�倎+@ܨ�pE�9Hz�c"OD��,ܲ?�:� �$Q�o�1`!"O �����*mL��m�=M#w"O�����ӽCE�����/$쭙�"O�+�DN)ܦ����1Չ�"O`H��/ZF�� hb��2��u�3"O8�A�7q !fe�
pt�0IQ"O�����+A��:	�Y��"O���� L�Q����cT6�i"O��'�Y2!����߼GN��{�"O�H9�74�X
3kT�#N�Q"O.��ckN-E�|��WI�'?��9"O2��K��z��!)R�v�|@�"O��A�lM�/��������B�X�
 "O"Ԉ��?EE�`��.;� �8�"O�}�J,Զ�avj�#w�� �"O>�[WLPj���A)��v��� "O�1� ��b|f9�?�JM#%"OZQA�C�'8x�p"��a��`:"O h��P+x�lJ��,*���a4"O\���],|�>�I��Y=f��0�"O�G �(rޙ#��Ʋk�	�Q"O �RvfB�v�,�zF�:)�^�+!"Oĝ�@��pH|�P6�[h�*�"O@�G,�(v{&A�����^ѸG"O�8�r.V�p�
w'���r�"O8r��V�NeaElU$u�ڢ"O��ƑR]*=��k�*W�0}A�"O��p���DE��+�/d�|"OZtk3�S	�D�KS/i�u��"O��!�%z�^�9K�3s�*u0�"O� �- R����W�D�<оy��"O���ǙR.±r�
��L!�"O�E�a��4+�ֱ�B� >6	2��1"O��f *~��;d�Ԓ@�j�ȗ"O���f!�`�J�*�^�>��xs��'|�'�2�'��'E��'#�'�I+�A^$ܴ��P��E[6�{��'�B�'���'+�'_2�'Qb�'�{`�˾RO��A���'|�x JT�'���'~��'���'<��'���'�R'�X*J��l1� 84���'���'�R�'���'F2�'�'�P�._�Bi4q���H@�h��'FB�'�R�'j�'r�'}��'W��s&�y��E#uÏ�#���(&�'M��',��'Z��'���'��'oh�Ȕ�F�O�͛r��|��l���'m"�'o��'��'L�'���'���8�͙\E
%���D�4�v��@�'���']2�']��'=�'���'���p�� -��)���1`�'O2�'���'s��'��'��'�V8Ir�ߘH�2%B%*Y�`��=�G�'��'���'�R�'���'�2�'�b�fҲC�`�ZU%����q9�'B�'�2�'v��'��'���'��3C��xz�A3���k�e��',r�'x��'��'lR�'a"�'"8@�"$N�I�mY�	��N��g�'=��'�B�'A��'lr"`Ӣ���O��ac"�>1T����
y��*Q�Xy�'
�)�3?y�i�8p�aa��0f�'`�~4́���$�ڦ��?��<��4>عR�Q�gjH��'
�(*�K��?i��ʡ�Mk�O��S��
H?	P��ǡ`ʄ�����%�>Q���4�T�'��>���f�-$��(�6n�U�Τ�Іܹ�M;���Z���OV6=��|K爎�A<N-��K��6���L�Oh�Dv�`ק�O[�ysr�i"�� <�0ň��'f�z�����'6��r�tj�{+̢=�'�?���$C�`X��8�� �G�<9,O��O�qoږqwRc�xX6B�"�&��ݹ{�6�a��G��="�������<�ON���b+�N��Z��s������U^̡�3)�+U_"�韬��$Q�}�<쑦a��?�$YŌ�Zy�W� �)��<�j
:zⰅ���£G�6mY�$V�<��i+�9q�O��n�n��|�RN�%1�
�'Kغhi��AC�<��?!�na@���4��y>m����(���CB���E��*i�0�2�$�<�'�?����?���?��l�Z������ܰoon����O!��Ď����0/�]y��'2�����̇�ln$���.��ݹ��I_}"Iu�<�m�9��Ş��,�.\0A�u����,��,G�n�	2�u]҉�pMУ�j4�^w��O��'� �ppj�=�شΆ L[hĻ��'���'�����X�"�4|�@Y��_oB�O�b`}2�9'g�d̓�&�Q}b$j����'+`��ރ ��8���]\^X��߿X���>O�pC�˫4B�J��\?J���]�2��`Z��܏�":	Y��I�D����`�	����Y��5����$��4�A���p��{+O�������%|>}�I��M�K>QSOA gNT��D7T(���k�4�'�$6�R��v��$n�L~⦞�@�>�CPh�0~����e+��=B�����w�|�_���?G�Y�1����)ҳy�&<���	L�'06mN>s�����O���|�n�:}0��"��9���hT�U`~B��>i@�iz�7_L�)b��.�ڸ�C�dB,�7�%4�p��@#H1^<,O��H��?Q�9���u0��1A׺����� b���D�O(���O���<���i�v��NZ�b8xR%��"{�M�D������'��6�/�4�>�'��/T��Ф��&9��d�	�9r�'����i1�i������?M�]�T���������w~}s�}�Ȕ'Ur�'>��'���'����X���Ҁ��@c��5Y���j�4�zX�(O��$��.���OB�d��6��*��L�_ ��ꔖH9�pi��M;Ǜ|�'�r�'p{���4�y�$ŗhh�qcq�A}��P���-�y�:x0�IE��Iڟ��'���'A��c���%��iR�?~��'���'��U�kܴB4@,O����;���h�69�lm�&�>ƪ�Oz���y}��'S�|b��AKP}�R
Ի���0��Y����Z'��K���ɼ����s���.�DX)sxq���6:�Ի�G��3�!�DD�J2�!�B���,�w�U�uv^��ަ�	!�Qڟ��I'�Mی�wT��`�'㨘x�) �0P�8�'��6mDզqشHafߴ�� <a��9��[D̓�@NԴ#"d�,5a�i�'d-�ĥ<Q��?��?)��?�m�=��*���P$L��Nġ��dU���0Ilyr�'��O�R&��Hd��'D�%���x�aAR�l��?���S�'%DJ<{Pቓ%e�1	gAύ]�-pToM'i��(Orq�� �=�?yJ)�D�<Iw��A���n�cg.t�6i���?Q��?���?�'��Wզa�hP��L�bş�b�:t��O'E|��×A֟L��4���|Q\�p@ܴ>�����q�V��P�ɲ@�2[����_ ��qog~RD^�~���S�9&�O� �p@
J��y���4t!�!8OB��O����O\���O��?E���'#�ȕ($mǕ)>ӗMUy��'�6-C3&i��O*inZF�	�:�����e�]a�d(1 wX�h&���	͟�S0�nZm~Zw��P�#W�+6��#�.[�$���A�:7£�m�	Pyr�'�2�'[2'~69h�(�+ )��@�rZ"�'���M6$F?�?)��?9*���!�
E<.
�sc���Ұ������O��d/�)�K?]I@��udL1N����I!��+!.^pG̨�.O�8�?��3�D�S����+_�z������@6 ��D�O����O^��<�&�i��{3j
�'����d�¨
��Y{#@�+7���'r66�I3��D�O��S�-!b>Yc#�6	�p�4�<1j���ic����EGL%ji��&�Oy���K�R�Iԧ�������y^����ݟ(�I��p���(�O� �E
��2���h�3y��Y��m�r�3O���O���d����)f�t����/9��4c@l��5�f��	���&��ן�I�6�l�<�7G�Qz�V#"���6K��<�g/x4.�Iw�I}yʟ�A�ц�=T�(��+lp���'��6T�[o����O��բ,�����ȴ-9h�*FGI���RϨ>���?�M>� AD�@��`$��c�AJ~�*�>T��(R�Vc��OE����c��/Li�j��B�I-�I)�E�4g���'�r�'q��S��|&o�&������l��yā����۴F�PC��?��i<�O�N�5I��)) ���i���>:d�d�O��$�O�=	�l���ӺC����´@�@l��##̓�'�ŢALD9d�O��?���?I��?)� /�r��({�ܸ�1i�iv���(Op�oU4X��ğ��}�ğJ3�*��5a���0��%^����O�$/��I�`��b��"4`��j�$>憱
��A/cN�˓@�L�����O�9�M>�.O���AAW�D�x���%�"!8�m�O����O����O�i�<�a�i�b�ʖ�'H��iWA9N�8E*a�`��cKr�u�D�`��OL���O����%V�H "F�M��5�>`�h�S��b���ޟ���	ԊM��D�nyB�O:��C�GYb$���O*2�P�4"�#�y��'��'��'v��)z���`2��W�X�s���C�����O������� �Rvy2�a�P���<Q��O�B #��N `0���V����?I���?�҈ȫ�M��'5��.kK�шUʔ����pf���QZ�9���OX�K>.O��d�O����OY�IЀd_NP���E1E�d�c�O^�d�<���i��´�'g�'U��*b�5�eX�P)x�e숯!�J�}���ߟ���S�i>M�	�h�,t娂�W����gT�����¼=���{5�@oy��O��4�I"��'U�2���qaA⴪ʧ}� 0��'���'�"���O����M��&@�-�XŪ㒇@�0�{t�>cݠ����?���i��O�'f"�ِ2ԞD�R��_��8'G��	���'�����i�D�O�=9�����qN�<�Œ�Xiʄ���D�6�U+&G�<�-O�$�O����O����O�ʧ`9��9�uy˵M�
,-pE�vmۣ�M[�-$�?A��?QN~�Ǜ�w� �� 폠:t�l �&�GR�ؖ�'2�O���O���D�.��6�f����N9k9
q[S�Z1N����Ix������4"�b�uy��'Z���& ^(���KD>@�!�S�U2�'��'(�I��M�Ca�%�?q��?1V D�d��pʴ�"#���@4��>��'7�ꓤ?ɈB�C(W9�� O��!����)����$�R'��;wIX�g�ؒ����e�J�D��_�)�3��15��HV� ���O���O�$5�'�?��'��S�� ��	��X#AH^��?��ihB�2��'%�`l����ݲ1MD`:��[z2��E��i��	ޟt�'���HW�i����^�8�V�OHD�j�`�3Chʉ���P�L��z��Vy���X�Laq`�M�(]z���0�,�c�v@�r:f��O��?Y����d���kJ4m�0ت4�R:���CΦ���4Z����O�fa����q?� ��g��j�i`aύ�xapW�����<>��O�	ByҨ��Q��x+e/��,җ���0>at�i�Zd���'J��B�\ x��Hk��k��:��'��7�4����$�榽Yܴ%ϛ�j��-H#��.ܤj&������Q�i����7Pv̂�OR�%?��� V�d���M?,	�.��`3O����Od�$�O�d�O��?Iȱ���[)(� �?vtrC�ş���ϟ��شL�8ļ�?i��ir�'9��� Z�1�na��>;t�᷃)�G֦m���|�r�˃�M��Oz4i2��NR^��C�*���"��*W@��8��O��?1��?���r�M�D-̅� ����$�u����?)OPo�n���'m2T>���U�͆x����&TO4�q�%?	%R����4)Z�6'�?ɩ�]�I�EI��p7�H"�蘝z):�I�#�\�JȖ��TG�̟P*��|�o�BKqCQ�=\�dX�3^�"�'�B�'&���P�Ȋ�4&B�KT@��z�ܤJQ�K�5�5KA���d��y�	m�	������8jWl{W*J�O[�I>�������ٴm0��4�y��'mr�����?HrU�� �@rk\�b
D�r7A�i���=O�˓�?����?a��?A����0Jtt�F��<'TIA`疟.DIm�f���	���	y�s� ���c���/N:!�4��!��i��	�?1����Ş� <Hܴ�y�P
�w�H.0���!�b���yR� 4qp�������4���dH �̩
��� v#��9a� ����O��$�O��A�����<��?ac� ~Bvđ�y����$k�O$!�'\"�'��'H�j���vVՒ���	��O ��&/�8~?�7M?�S�q���O�K4O
�n�A����(�Zp"O޹�a����.ś2�ډc��huB�O|�m�.x�I����@��4���yW(ڲ4�@ �-+��t�U�y2@dӸ	o���M�c
��M3�O��k$(�+�r�揃t���3��,NZd&�עs�l�OPʓ�?���?����?!�I�tUض�3=F��b��	zm��*-Oh�m��L��I�X��]�s�,� JU4}�a*Q�M�5m8����OR��!����<�&��3�K��l� �L�@���>L,ʓ3MJ�5b�O�0�J>�-O�����D�s��re	%/dN�Pw��O���O����O�)�<Qa�io �e�'h���gH�g�3(���iR�'6� �4�dq�'v�7���1pشr�p�r���>��D���%U=�(�@�E2�M��O\���d_��ڲ�(�)���d�&�Y	�<��la��>O����O��d�OL���O��?5( `A�)��Y��MܑJY�<�	8?����vl���$M�%$���Df\/LqX� ��[�@U�2@h�����i>��1,�����'�"	7��d�
)�t@ӓp+z�	NT*B^Y�����4�6�D�O`��5������O�̱��I����$�O>˓ۛ��ȗB�����0�O���S�[�B��!���!B��p��'.�>1���?aI>�OM��yFE��S�*�p �U9j�2t���
�g�E95���p��i>�"d�'<��&��ڲ,��%%�9�!$���J"l�� �	֟��	��b>�'��6�Ϙ-�*��$ɞ,D�a�ؤjhq�(�O���٦1�?y�W��I�e�m�"a���P�%����I����'� ɦy�u�d�����%by2l�c�z���O�u��X��H^��yBX��I�����@�I�ЖO������,PHǍ<FaC#�k��9*��<�����?�Ż�yW�A�'���S���!#f� !�/UR�4��$�O^� 4�a�b��xƖ��7'ÌW�hl�T�L>"�D�I?}E2�h�'P��&��'�r4�p��\�k��݃6��1HVihp�'�2�'�W���޴n^Eϓ�?q���t��!�Af@O� $
h���k�>���?YJ>y�K�^�9�dd����� ��<�dFJq��Ϟ�M��O��)?�~��'�(D��\��}�ׇߔ��� �'4��'(��'��>�]�M�h�+���µ��B�%tJ���I-�M x~�p�d��]��\1h �?*z�Qc�	hr�	۟���ʟ�Pv�����?i������?mxj��t`B�.�r��ҁ�:KlD�'�������'���'���'b`���$X�J�:
vb j7�h6U��zٴw�jT����?����<�R��*u��T��G��2�����)s��	ǟ��Ie�)擡kn�9 ��#��k�"��cf�y�����8�'���p������s�|�V�8Y�l.9L�q��"�$��U�T�ן��	� �I��jy�`ӂ���G�OT��� ��`d�<h׶�S�&�O��m�C�i>��O �d�OP��Ӎ[�T=��!Pbȉ�G�/_ށ��oӾ�I
|QT��0��J~���UPT
 EQ5^� ���0 ��L���?91�ǌ'���weO3
���4�ܗ�?a���?�r�i\�͟� m�V�	!6Rd��T�P�"\Ȑ���w�v�I<���i��7=�*�,}���@<����]+T�b4�o�n{F 2N,����F3�䓮�$�O��$�O��G!��� ���;ĝ�p/�BN ���O�ʓc�F��PR��'��X>�[5�˝`h����K^���z3l=?�`P����ڟ�%���Z h"�**P�p0o�;ľq��� K2�ѧB�4��4� e��T��ObLtЀ9���xPm��2��(����O���O��$�O��
?FK�<��iO||#�
�]/��YVi�U���v���B��I2�M�J>a�O���ݟ���7��������U�8A1h���I:USlDn�<a��oT	�թ񟠜1(O������I���s�0��W;O�˓�?9��?)���?�����V�cv�s��v�B��fk
�F��m�F�RI�	�`���?A���ş��ɞ�Mϻ4��r�a��P&��r�
&<^(�H�����T�'��o(��=O `'��x{,�@ʟ�p5��h3O��8�'��?!W�4���<!��?Q'I_�����VH� �Rg���?A���?�����Ĝ˦C�������C�#܏;��9�V�̹2ǲ��Èx��ea���8�Iy�#=�dR��5 Ą��JՔg��j�������~�<ВN~� �O(���p0-5c���X��%i!�i����?���?I���h�V��D�dV���+�5uv�2�%p�K��'��6��"t�	&�M���w����gGa4	��(�gn}қ'�r�'�rlށߛv1O���P/1����π ̙*�dún\(������B�<�d�<ͧ�?����?9��?	�_@_�Q%� �ݓb�U����5e͞՟��I㟼&?��S�N�[U)Y"�)*Ş��5B-�>�`�i��7l�)��G#8�p C�w�y����2����A�5z�'�����i�ş��1�|�Y��;`��S���S�*L�S�`� �o��l���(������IyB��O&����' �\����
U3[�M��D�'47�8�ɢ��d�O:�k�(<@d��3���dH�7P{�Ea ��M�'��nO�(ܜE��g@��?U����$)�F 2|��!�d��[ˠ�	ҟp�I���֟p�Ia��}C6�kbǉ51*e�3�ƪ5+.�/O��F���3��h>��,�M�I>���P�~���ʀC+2꒸��
z��'D�7��ަ�S�*=o�P~"ѓ����K	u�a����d�
1������0��|�[�������������5CI��(`Ȓ)nta ̟ϟ���By��gӼ�<O�d�O��'KMX�����	U�82�N�+Y�R8�'���?������|
�`�<�u��r�G�+]��;�c�LlA�4������'��'�9�pD�0>Tz�Z���d����'{��'hR���OS�ɓ�M#���1�%+�G��1|^�KZ',x��'��6�,�����O`�C'�lh���� ?�U����O���W�W�66�e��I8�д{��~�*���H'eŠm� 9CQ+Q������$�Oj��O����Oz���|�Q���u0$9Q�	�F��<x���9ߴN=q.O���&���Oмoz�A�ŌX��`�j�c_��4���H��V�)�S�ve��o�<�v�$4�e��;c��4ۓ�<�1 I�W����J3����d�O����$v���u�ƌt��2L�o����O���O��[��HT��y��'MY'Vt��v��p)	5���|��Ox��'�r�'��'�ŀ���/kl����'�m�����O��!t��/a�x7�>�S_����O$�`"h��|��{�h��C':y �O���O<���O�}��DW�t�Hf�a��!�Ca8��%ӛFj˶,�R�'7�6�)�i�E�E��KQ��1���<6%��h����wy��A)6o�����c#�Ѱ[��̌#J�E�#��Kׂ�zt��<\+'���'�2�'�R�'�B�'��`�B-�$���d�L�p���Z��R�4u����,O���?�)�O���f�ɚ-�@&/ �P���+c��n}B�'��O�)�O��e<~}�"�ϗ=y����'ؠ��Eؗ.Mjʓk�`�"��O�4�K>�*O�t8��J�'��qx�c�9T�����O��d�O���O�)�<�P�i ��C��'fr|8W�	�Q������
R��Zp�'�6m?������O���de��B8~�=�S�S#qi�!��	�M{�Oƥa��ų���6����~�k��3�E�d�N��s�0O���O����O�D�O��?͂���5C
�%�r�P�>�P��H�my"�'��6�G4l��O�m��I"&�8b��B�Q���/�6�c��	Qybg#"ԛf��0 ��$!dL�	��K��������~l�'���%�d�'nb�'�r�'�X�	C��=�r%	�G3QH���'��[�h�ش8�H�q��?�����iC�t�F�('��4��y�i�=n%�	���d�O6���ʟ���\��슆d��DRސ��,�=@���`�O�hM�y�'���Eџ �v�|�o�dB���0b�	�c<�b�'���'���Y�ȊشrR�$�U�÷|�& #�ᓦ5*�5��b~"�`���4٨O��D6 *�ɰ�Er�2a�I��o����O���Oc���Ni�lr C<Cf���a�]��r�D+��V���|yb�'U�'�"�'U�Q>1tNշ��p�-T6[��:,�0�M�$��?���?A����9O�lzމ4��
R��j���6g���!ʜ��,�?ͧ�?i��S��۴�y�o�.+!��KF��!Z��{��ѣ�yB��d�H�I�'�'��	ş���e�]X�%H�DG"�!uf%\���	��D��ܟ`�'Jr6- 	6���?�u�4WFT%��l�=e"��Ȧ����?ISZ��#ڴ̛6l$��0&����� ����9�+�:\Q�	1#���W�6u�|�$?���'�|��	>���w'�+{�!S�QV���IƟ��	����	S�x���'+НÓhՉ���0����@�T���'�27���2'���O��o�q��李���Ӵ�T�\�n��'I�K��	ޟ4�I�,��(�IΓ�?yu���6����U�J&\��K#���XԂɟ2%�(�N>I,O���OZ���O��D�Od���ڞdUfM��"[;��d��Ƞ<��i��y��'��'��OK��.�� �O��Z��Pr�"Z�>j��?���O�r�'f��2��# ��Y��5 �4� -��AT<(ze\�@�ǂ����c�	vy�&B�[NXmٲ�؎{���7��ct�'�2�'u�OU�I��M˥e�1�?	�ć�-���7��&i����2�?y_����?��Z���	Fy�F#Rf�P�!Բ@�|��� �'d��TK��i�����A�O.�M%?���LN�+$o�
`ɘ1_%~X�����	����ܟ���B��	�x��G����ZM�lKΌf~B�'�6-X���$�M�H>��ʝ ]��NbQ:�������?a��?�d"��M�'�%F��� D �a��Xo24Se$G�r�@��~��|P��S����IƟ(�5M_>S��x���j� ��w �ڟ$��Gyr�xӼ�X�?O<�d�O�ʧ|�ޔC�26�����=�F��'�4��?�����S���Z$Ms����@ڝVs���'R�
���Dk�5u��&����$-��D.���Uq���S(C�^�p,A�k ����O�$�OP��<��i���
 �ӥO�H�2͚2c=3��:���L��?�f]�8��&	��в�C	/�ll#@+ɛH h������`Ԧ��'�,aQ��`ܧ>+�z����zP����Jg�e̓��d�O ���O>���O����|"�j@�)���;A����\(`�F���m�&�y�'���'�26=��P��څ^Hn�)U��-̀R���Oh��'��i��o�7�v��:�#Ҿfi�5��.e�0!)D-k����f/X��$)�$�<�Oڲm1�VC.5`��E�D�Q
Ó��&�fT��'���%P����M�Y��x"4���\�OX��'��'��'���IA�I�x�(��(G�����O�Qx�	�jk@S=�)��?!�Oz	����L��l�iA�i�h�rR"O��R�G(���.vHe�F/�O��m3�q���L[ߴ���y�M�/C�Qa�r|f�b@��y�'��'-�1饱ii�i��c FI�?�2�B��&���b)�9<�ʁB�j�ma�'��	X�'޸!����.^�ĂS�Ǫg_bl��O �mZ5H��m�I����V�'J�f9x!�G�J�8B���X?�Za_�T0�4��6�'��ɗYz�$ �n��u�T<�dF���͙�U�b��c�nd�G�O��I>�,Oz��*T�tIЄ+�@��2S*�O���O<��O�<���i\.M!��'��ի&�W���pґb<�vp�1�'�@7�3�ɓ��$�O"�$�Od a Ɓ45{6�aa�)z@��D�H?<7�r�,��yٚ�P��O`�L�'t�t�w�:LQ���-AKx�`@���#�Լ��'I2�'���'��'�2��ƏM�n� ����؂p{7��O����O&alZr�d�S۟���4��N�в���C�R���M�w�Dp�L>����?��?{���ش�y�ԟD�O�#@�P) �]���FT?9����䓻��OP���O���ˑ�0=I������J��=y����O��uśf��P���'C�Z>������_��A�b�J�@�̝��O<?y#T����`$��\����r�C���R�ٸD��|���+i\y��/��4��H��%h��O��RD%�46�t(�^,/>t����O��D�O,���O1���	���ˁw�J��&���)���0aF�[��p�[�48۴��'��ʓ�M��G<h�J��T'g�z�NZ�q��&�r���f�n�"�k���ad�p�K.O��d��?2�@�1Gē)sEz�#0O^ʓ�?Q���?����?A���I�:r�^L�A�_C�m�ࡕ
�x`o�~i`%����	\���H����{��@>Rz@ ��^��lug*��G��j�Ĩ$�b> ��զ�͓<]���1%ɒt�,�&DV�qK�ϓS-����On�SM>�/OV�d�OR���:AK1DZ:8������O��D�O���<��i�����'Y��'P>��F�2����Կms��`��'i�'����?���6Z�@Kr/	�a� X��y��'��x�dZ(dD0u�X���Ӑh��a\�Q1���Nq��)�M� u�y�4�Dܟ��	ڟ������E���'P�a@�)-;���4.��g��8��'**6�0V�����O��o�K�ӼC��	(a` ���%80��(�<����d�(�<79?�c�E�/�h�iщ_Xp9�dI؜G2��b$E�L���O>�*O����O~�$�O���Ol%�ta�@��$!c	P�Pk�4��<���i�~�S#�'���'T�0x�]	%�����)ǛXXM�E�D}��'��O�	�O4�D@"�	[��H:U���"T)�KJ�s�E�0��jt,a�n�O�;J>y-OL<RGm^'o���I��8L����'06�̰yD�DJ4�X����V�y��H�ʶb��ăȦ��?	�S����4{ڛ6d�V ��ŗKP����P�e�j9 �t=�7�7?��U����I��䧔���l���U�*ޗY&t(Ee�<��?y���?Q��?�O~f�I�c�la#�b �\����N� ������?���or��-��s���M�N>�$�?��eԦ7�n�%�Ox̓�?����?Y��&�M��'"D�%+��`��}�=�����|X�,�&����|R� �?YS)�	\tq��k�7+:�Tb�u�'�:6mv,�D�O���|Z�2����5���u>*����q~R��>	�i�D7��)��N�H�|���N�d �\�%��!�6J&B��h,O�)��?��9�$�j~��h��ڰ�KY.y9*��O����O���i�<yV�irzTz��"Y:��]�F��e!� (g���'��7�8�ɐ��D�O"�RE&׷jf�y	u�R|�u�� �Ov��H�6m2?��Gf�q1�'W||˓
j\E��N o2��{Wc�"Ex������O^�d�O��O��Ĩ|�����
=���ʤq$�T�#T�]]�V��
uR�Iޟ��OV�'�d6=����D��l\�r�̈W�5Z�L�O�������I�ҘDm��<� Zp�a��(� 3���I*�r�;O��1s`���?���'��<����?��`��a ��@`eЫ oD�c ���?Y��?I����Ħ)���U˟�����X��!��_���
�L�
�"�L@g����"�M��i)O�EE��1�� f� 4P�	唟dA��T�SN�|
C*TL�1RG*ޟD���h�&��!&fytSDm������ڟT���pE��wR{�D �BŞ��#�T���h���'`6��8'x��d�O�EnZA�i>��;,�h����Qu��6ʽ�6�I�M��i��7��($t6m+?i�m�t>���-O�`�Y�ሃk�(@*���4Bf��N>1.O��d�O����O����O�My�&�x����mC�͘���<9��i_L���'�B�'d�O��a�)6�Aj� :V�p�T�Z����f�`�Ɯ&�b>5w�y8lԚ��o��r�e�0_+����#[yR�]��z��	�l��'�剰]�	��׌D����3D�'l�D�IΟ���؟D�i>ݕ'-�6-H�M����!_g�,�V�ҥb;|e��` �D����զU&��S�����k�4w���"��N�0�g��h�"�!�G��fQ�1�e�i����P��O7��&?����l~�hb
؇W�p����Ѥn���l����\�I�|�	S�'x��؉�-�$�����Yr�����?)��S��l���d�'��7�?��V*Lb��0��/w�Š���(7}j�Op���O���]5�63?�;abHc�O��(P��A!8mH��e��?�q�+��<����L�j����Z�<�(S�X3�O��oZ�x2!�	��I`���T[6� �Od�.ܙ��@����X}��`�ޑn���S� R�9����A.�>ٜ%c�b1"��c(�[�y�Y���&qz�ev�	9��[F��3�ؔ���O�09�����	���)�by��eӞ}ٲ A�4��U
�:{p܁a<8
�q?�F��H}�K~Ӑy �_1#�h���c�Bڧצ�#�4U��M��4��D1v#���,�<�ӥ��,z1�O5{>��do��<�*O����O\�d�O$���O�˧"������PVǬ񚒫��4pXоi�F��'V"�'L�OU�q��.�}zP!9��U�0�eH�?ݲIo
�M���x��d�[v�&3O��If�C�ca�A`��n��<O64x��҆�?10�?�D�<�/OXiP���+'<�r"��],t�A�'{�7�ȣ=�����OB�R�vt�S2
��<����UW�"�(�P�O4��O��O�"m��^��X�$0a��a����CeI�(�x�c�j�ӕ)��\�����K��b�x�/͑]G� Ӳ������؟L�	���'?E"�kt>��I:(�>Ȁ�k�y��L�:E�a+!�'}�7̀1n��R�Ɨ|b��y�!�5"V �(E`�:�"��_'�yb�'���'@�c�i���O��EFJ?��FD-g��tjQ� L�ꥠe��cf�O���?���?���?���2S4P���-7�Q6��
'����*O*l�*i�T�I՟h��V�s����O���S�À�D�cҨJ%���O<��>���I1m���R�&	2!��	�R��	{,\�bD~��;���a��� %�Ԕ'Ɍ�{�B8q��Ve=�<ɐ��'>��'v2����P���ݴI���y�∘��/;����F�_Lل4̓2#�6�DO}��'��'HZU)�`F.tl:��e�V�*��!�iȤ��v���#���VSQ>5�ݲ+	&�q�K�R����.D���Iݟ��	���I����IV����D-S+y�ޥ�#*K������?��<�fM������'MR7M/�D��K�s�\�-�ĉ��̌m���O����O�	Or��6�/?��f�&�B�
=�`�XԨAqb�C5G@��?��)/��<���?Y��?�I[)VK�x�JU�+ 98��^��?I����$��},j����O��D�|:#�0%�1�C��n����jG~�l�>����?�I>�OtptH�\��j`MT-$*�Q���G�0�+���"q��i>1"')�	�4���G�Ue��G�
2�K4�g4�9�Iȶ-��H�@Z�^��������;�L��u���Kl$�PrOŬ�,��bG��,"�9�kՈ�j��fB�8+s��9��p���
u�zAaB�9"P	�iQ��:=��g�� ��>Ŕ�Q�-��%�@骷���C����8Ê��p?�	a@��4�$��(��	ؐI�4�<�B��Ȑ�C�f�
Q"�I
��1gȰDWy��营
���u"�g�|�����W����Ӥ�f`��S���� w/��:�>$�%(:�f� b��r� ��C��'��|�P��KҊ�?vL���G��P8 �#���b���Iϟ4��ny�ɓ�8��~���n�O�X���J�[ .��?	�����d��c���u��az���95��xqP�ՉE2��?����?!*O2�{�&�[�S�e��,{T��,U����&�J��Qܴ�?�L>�+Oj� ��d�0@���A�C)�����C&>N�f�'rP�,��)W��ħ�?��� @�(
�[������F T����a�x�Y�(( ?�S�T�V�_�Y�/�*�"m1�.0�M�,O�)	P٦�3����������'�p�R�ĭf܈PB�����Hٴ��䄱��b?]�#O�'�����+w��e��duӞ!��#٦=����,���?8�}�NX�u]V�Ѥ®W����Td�+h7��'��"|��5�X�[��W"�h�J\3`="�"a�i���'��ַQ�
c���	���� 6�����,8U�2,ρz����@�1O��D�O�����5!`DRgC�?Kbu�J�j���m�̟�CI�ē�?������s���5��l��F�EJ �A -�W}�,���'��'��h{t�Uo
��!��4@��1I��`V̨%�����%���';^�pg ˟@�$l��jƼh�f���յ�'���'12Z�@��+@,���d��f��ԛTJ� VP��f�����?�O>�/Ob�]��SF�{Dy�T�js#囫��$�O@���O^˓]kM귖�tF��#�ʸ� �]]��"�gK&s��6��O��On˓�l��>�5�Ѵ5�)����;�ư0�)�ߦ��I��ܗ'*n�C:�	�O����4u����M�м@ǁ�{.i&����t�X�g*�1YNLpe-Ջ�7ͱ<�WD�(��&�'�r�'��s��X�!���&hP8�촁�딎"p�6��O��K��f��!�$8��"vN�����;�I��I?&�7�^$M�<o�ҟl��ɟ���1��ĳ<�#�~����"5����#��(}�+P���On�?��	�B�:�`��5gjY��d�7' ʉ�۴�?����?���9Uq��uyb�'���ya@D!d)N"J�;��E5Yg��|��U�2_��������i���4
�O[R�*$�ۿS	D0T�n���d�B��x�'����d%���/���e��AwP�òh��J���H4�?�$�O��D�O˓Hg�ə�m�ni@Q[Fi�
n@��`2�ٜ���sy��'8���t�	����B4D�8�:A�M��SG/L��\'�X�I�$��oy�b��U6�S�rł�3P	C�&V��#ɕ4�.7�<������?��v�vs�'+�*�:A���˾M�t�O����O��D�<3�̿h����*���[\�C�'�*k�b�R ���M;����?1��Eΐ�b�{�K��>�j��e�TZ����ˊ�M����?+O&)�4C�_�d�'��O��P�A&~���Ŧ�&V�,A{�M,��O��dѷ+�:�t�'E|� �"S�]����"04LAm�^y��ô���'��'���X��X1[bF08�%D$$���c̄ p%B7m�O�����4A��b?�"ǣ� ����f�3N�u�CGp��C�@�A�����	�?=3�Ol˓���R%�B�SʤXǄ^�#�T�ƶi�8��`�$5�S���ӎ�n����Yz��xc��y���o�ğ���ݟ@s֊�����|���?��킀.�*(ha��b;���ĬJ�sϛ�',r\�${��X�'��i fm�g.���H���,�'e�F�h�O4�)Ub�<�)O��h�פ�:>"B� �Ο�~���0
��ē���<�����$�O�P8f���|�@	bM�Ff�(ia$��?1���'�2�O�|p� ��}���+�����i��8�y2�'���ߟ\;�or�#$�T����H���S��������D�?����dY�ěgQ
D|�s��!9N���o
���?1*OP��PA��'�?������[���t�B��T&\Hڛ6�$�O�ʓA�m%�(����K/>=y!�X#~��;$v���O&��rA�Z4�ħ�?����#�+5�����*}kTl�G+�h�Ky��'/����u7��$/�h���M_V�B�)	�����O�S�
�O���O�����Ӻ�ԚC].�jt�Ɋ-� %�U��̦���Ey��N�O�O��e���PZ	��m_�h��H��4�&9��?���?!�'��?����e��|(�86mX�����MS��Jp�|@�<E��g�/�Y[#ڊ'���Ԫ[�Ur��'+�'mj1Q5W��'��$*"$K�!��n����2���$9��Y�y�+ԩ
�P�d���O��d��a
^���o�Z}���	 y�(5lZ˟lۤ��&���|������O\�z�cWT�P��0b�5l�xMC��D|}�'1;�Y����ʟ��	dy2�S)(	qul؊XݒE@�s���;��2��OD���O�˓�?��E����`[<EF�
SI6J��Y�"���?9M>)��?1-O��u�W�|"2�G�X?�ȃ��=��B��a}r�'���'T�៼�I+X������
x�].4��bg�ߝD�tl�$�ۑ��$�O��$�O�ʓ9l������T)1?������D�D?���M�%z�7m�OԒO��P��}����S yW���1��9A�h���ДZ�V6-�O���<���ۼ_��O\���5&�E>90��3�&��=��J�%��ē��$ί���8���?�����\57D�%��+e���E���h��i�R�'�?��2	��(>7D��"�=l�����#<6ͦ<	W�X��?A�����ܴDg�B6��;`qީ�f��"L�2 lZ j������0�I����{yʟ �$�H��Px�O�"�lh*U�צ	(Gx	�����rL1�����h	-|xy#����M���?���ǁ�'���|����~�̿ta���x=<-�-Z�0�BP�H�6�]���9O����O���_�8��]�#f
M����0Z��m���lBE�	����|�����Ӻ�gϜ"�!��L��3�� ��X}R��hv�U��������	Vy2k��(p�G���(p���oďu��i��"�$�Od�-��<�� ��ҀC̣M{�,(q�ݟM(���d�2�?�-O4�D�O��$�<��H�
N󩟡K���剓9P^6<a��[m�I��K�	nybhU���+7n��DD�h�,b�� �ꓼ?����?�,O����P��'�iʥ����H���p��\B�Fy��d�<a��?Q��#��<Γ�?A�'y�9�G�Qyz�G9�l�۴�?�����ě">�L��O��'����^(S������f� ���N�!���?I���?Y� �<�M>��O�B` �%�!a����+z�۴��$Ļ��Qm��D��ោ��������(V5/v�C��
Ct<m1�i���'�L}x�'��'�q���:e�,�d���N��}+��i>� k��rӊ���O����"X�'���'[U�<I�O��>�ry��0J��u!�4[������Odb!I�y(=S�E*c�j,Ҩ=��6��O��$�Oxi�G@R}�U���ID?顭I$�ek�ȇ�A��d��æ9%�T�Rhn��?q��?aI��u��%�G��\��������'S|1�Ģ>Q)Od�D�<Y���.��y�P�c�(��%�ԄSLUT}����y��'���'i��'h�I�S�<�ˆ �ZnZPR@�	d` ��r�����<������ON���O��鄭�G��)��G8;��Z�c���$�O|���Ov���O�˓~yJ�X�3��@ 䢔�^� �(���5)PH�Y�i��	���'���'���ɴ�y��ŵОɚLF�i 
�g���{{�7-�O���O��D�<	�o�4d��ܟ�X�p-�1bSl�6���D�3UL�6��O�˓�?i���?�Ed
�<a+�f���@t�����9\��,���ͦY����'_�yK�N�~���?��'^��!k �Y䄩0��(fp�(i�R���	ş4��-3c\�'��Ĺ?��QF��3߸|�gD2k�tbc��ʓo]�]K�i>��'���O��Ӻ�&���z���jb��ECrͨ�/ئ���ӟH��m����yy��ɐ�G�Pc��rl��� z�f�D�j��7��O����O���y}r_��RwhփDu����)Il@� ��>�M�&��<�O>a��$�'BI�J͌ڌ|	�팜GF��t��j�D�O���'����'�����p��I�f �y0�my"��%�@!o����'w��r���I�O����O�k1�dct��g��VP����U��0�N��O�˓�?�.O����-������d���MxtQ�d\�Ry�ȗ'J��'�2_�L3R��Z*H�X$�Υ�z�a��G����O>��?�.O<�$�O
�DC Z	��҄
��֑��)Soj��0O�ʓ�?!��?�*O"Aڶ�M�|���ɠ���Jڃ[a��������'�B\��	�������I�AT����<:��Rd��-�V��Oj���ON��<a1LQ����'�4-�I'hd��q���M�����O����Ol��$:Oh�'[N$u�D�S�����&gOrR�i���'��	6=��ѹ��f���O0���u���i!�) ��}���[+O^�'���'�����y�^>�	k�k'B��c���s�`:�h�⦉�'߾5�Shs���D�O�����`֧uMXyμ��O9y*<i"ҏ�M#���?)�"��<�W?��yܧ1BT���;��Yc1��T��em.-��:޴�?���?��'"��	my���+dP�3EO�,H��#¦�\(B6퉜Fh�����2D`b�D�gr��$���Q��iYr�'���
�*�D����O��	&(��u�D(F?u:��Q�jV�IB 6��O�>@V��S�4�'YB�'��E�T�ߙ w�eS#+�-F�B��s�a���䖆{k���'����d�'�Zc���W��,�Z�;P�M9r����4�?��JI�<a/O����O����<���T�0 ���6��R�U6F�y��Z�d�'�2T�`��֟����?��@5�? Mpk0��W��R�y���I��x�I�X�I}y�B��+^�擾(	���b�> ��-ѤA��6M�<����d�O@���O�a @=O�i��E7ʝ�U�A$ r>��qGЦ���ן��Iʟ̖'��Q�tN�~����E.�9{v�(hǢ؝C&ԱB6I�̦���]y��'��'*()��'��I�s�R�>���w`^"7��H{ٴ�?a����d	���$�O���'���JYj��S��	8����J Lf>��?)���?����u~BP���'P���:��y���;�%�1�<Yش��$�:�8�mZ����ioZ�?��O����T�1�ݜ3�TY�D埡!��'9�
��y��'*��'dq�� '��u��Z�Ɏ_-J��$�iz�+rӼ���O2�D���M�'���6	� �w�ܤ[�*X[gZ�EGD͋�4^�JM��?�)O�?)���z|p�r�#�x��j��β,2���4�?!��?Y`I&��	Cy��'���`Ί-9T� 2c���	'�F#<�V�'��	8�2�)����?i�`��ѽA��rA��?��@#0h���M��4��uZ�W���'	�[���i�����8�>Q�8B� �1:(�d��YΓ�?����?����?A(O@�XR$E�@:�`���Z����AE�2D�Y�'���ҟ�'�r�'JB�A+
�V���zb ����%1^X(�'���'&r�'��s��fI6��D���҈s�ߴb5Hf/]��M{*Od�ģ<q���?��a�\Y�$"H��B�g=�m�!��(",< �\���	��D�IQy�F>-�Bꧦ?��"NAX�`��ns|�h3�ȣ_͛6�'���ɟ������:�j���	�
� �Aj�!�j�����^���ixB�'��I)�"�⨟����O����H����cMW�5�|m�����G����'���'�B-Y.�y��'���T�P(
�`��0#��9x�i��cĦA�'.����#s���d�O���蟌i֧u!\p�\�Fh;~�����޼�MC��?�0A�<���?�����O؈H e%T#�n ���*�-�ߴ_�0��W�iO��'�r�O�O���)�6�I����\L��O'j�oڭ`�*�	K�F�'�?�G�b��D�3$'�r���%Q�pқf�'r��'�j��!:���O����|�Ʈ�:W�(��c'�

=^I���w�ГO0k�aUo��ܟ�	⟴+d̉1�8��[�
��%��n�؟ܪ�â��'���|Zc��AC����(�pq�TKR?P��ڬOް���O�ʓ�?�����'<��
Uc�g�(�[GI�	V:�b�٨,6�'��'H�'��'�
�R�E4#�l̘���>@��@���yr^���蟐��yy����F擳az 
�#�+0���1��R��O�D8�$�O�D�Y���A�5В�zs�W�"Θ���زK4���'�r�'�V�\ �����'d��"�jS�hԸ\�@.H��<�y�ie�|��'d�����>aAʋ�,����� J��yk6˂ߦ���ܟ�'�&�)e+5��O��ɉ�.�b۴ė=w�z�)��2C�8}%���	�0�DL̟�&�t��j9���U��Z����L�-g�qm�wyBI�f�h7mW���'���6?9P
C1D��a��eY)��Ś�֦e����`*�e���&�(�}�R�܀	$Z�0@�-r[i�eM֦Aa�Ė�M����?I��%�$� ����`��0^ü���	T*1��o+S��	v�s�'�?�G
�N걑�����%��3қ��'��'H5��):�	؟8�)�8��S*��XH����B(oF�IBb�)R��?	���
�q�e�:z���ک(O4�ӻio�.:2GDc�<��U�i����$�&y �)�(��@�JJe	�>)��έ�?.O��d�O*���	�'L��}���B��\�� ���ǐQ�dd&����ן�$����ן�
Ц��{0�=;�#�`��!����Isy��'X2�'��	;@X !��O�6�3D�m�0����&m����O����O�O����Oz�/�y�ΈT� @ �獯d�tř�$�_	,��?Y���?A(OVt���Gn��4 C��F�L��6���,�d�F���4�?aJ>���?�o��?iK�t�1�J��>��A�9�T}������D�Oʓ<����e��d�'I�4���#����fB�A^�=w����O����O0�� �OܒOz��n�eQR�<����5 ҭH� 7�<A�jL,P��6�~
�������	�xєY4 ��#����%a�<��O���FG�O��O�>�f聽M��桓6h,TH[�!~� A{��^����I˟`�	�?uH<ͧX�����MO�)��וn�ms�X� �If�S�'�?9H��4��4��P�%���E�<;�6�'^��'��D��<�4��'T*�HnG���/��aѲJ��MS�2$8�)�O�D�On$��fр�@���+��N2df��Ԧ)�	4(pE	J<ͧ�(O�hQ&oա9.�Da�$]u��xE�x��'��I���I���'�E8 �Sy�`�sa ��֢�P�KS�8O����O���<����?S��L��a��̐h|����/r��U�<����?�.O|��O�}���$�V�4;C��t1�q7I�H�>�m�۟����`%� ��Ay.��M3J�r��Ju��:ޤ�&K_}r�'w��'X剼h��5�I|�Č��6�Hmt	P(H�i7#D�N���'��'����=. >��coä~�Ryi����F��7m�Oz���<��mUt�O���O>,�m�`R���g �<[|d)%<���O ��'[T�L�'~�Q�R"7�l�A�*�l|o�|y�#U�u�6-�w��'k�Ԉ*?�@�%C�:G윒,��P`�ަ��	����:��O@�DQ䓵_���S2�
�j����4	(x���?y*Od�)�<�OS��b!�;e���Õ䒖3LDܓ���>Q��Q���O��#ۇK 0n��#9�[�06K�O,���ONh�Ɵ@��ß��{?qeU�+�`s𩅡�d�(0	�y؞@�Iǟ����&��9
� Ƹ0#P���a��D2�4�?�5CJ&�'�"�'-ɧ5�̝�D�|��`�;L)&�ÂE���F�G�1OF���Oh�$�<qU�ęF�=���72���E��a���x��'�b�|��'�2��4�j��O��I��l�AG'wb�ۊy��'02�'��	�h�|��O��sK�I:11l%J�j�K�4���O˓�?���?���^T}�.
�Z4��dn.�4��C畇���O@���O>ʓS�	�U?]�I�Z�l
�-���ܙb�
2�F���4�?�)O����O��D��z�$�|2$-3Q�UcEiεX��ؠ͘�����'�[� B�#��	�O4���D�T���]!"���N�h�}�Y�(���|��qo���P��' �IU+��р�舕|�V� �%�4K��vU�,�����Ms��?������U���5^x��T5e�� p�mI�'�&7��O �dM�Q���d��'�q�� ��"���B�l�W�A�= ]�C�i"a�A"|�\���O��������'�	//�N�����-P	�$�sN+Q��K�4� �'��I�'F7>yo� q��!�c�||���"���p`pB�I�>(��W'eӜ4i�A��D*^��Dފjxx��oV��Q �,"vu�0�����`��@�c,z�`c�P�_tl�qm
J#���#�8
&չ��ʝ*�N  �
� ���0F&1f�[v��:�X���MuH
��w�Z�{2�b���D��%C:O*��'�C�-���PrFCK"����'IT�=x�% l��'nB�'��� �'b�0�f�w(}���$F�W�r��*�&� �y���J	�|b�~_��P����������J�F�V4��DQ�r�'��k�h�:h�����f����@�|��'�b��?��C�)�� "��(v*��+gk D��i��ٴt���kQ#2��p02h`����4�?�-O��˅e���'I哙'eB�ˡ�ӝsU�"�ʏm��[�)�����Iݟ��# �%"�%����D`m��S���E�h�UBK�0jL2�X1�G�(O��`CȲxj�rP��(j"��x`�&Q���˘$NT8�Q�I6���Ol�?i�dN�X �lYFB!@��uj��q�(���+m8�`��8NwHc0*����e�	"H.qA ��!S1(yԦ��8t:�Ie|V2�OX���|���� �?��?�HT�.����;	��ы⢗)ښ��,߲vJ��CP�I*�c>�dC0L똝�)I��,��r�6D���{�LLɰiN����)���(�x�|�Â�Z%Ĩ(5&/x�R �I���'��(?�<��4{�BH3%�H�l���ȓHn��6C���1�'�2�~\Fx2�*�S���9&��c��D����E�K��'���fа]W��'Y��'� ��֟�ɚ��j腱1���3���y����pHj�����]!@��Ơ۳����99�B�U�ָ��I�R&��:DA��<(�[�	٩j��	!R����OD�O����OH˓\It8@��>;Kʝ��$�	�� ��-bS��[�N/�8�4 K��+��)R�ʮ�<8id
����A	3�y�XD�ĉ*�iN3��<�$��y2j�w�"���ي�H����y2�I�f[4����fPf�j�c]�y��2$��tyRÐ/XZke,��yB��*p��iK�A(M�d%��y�Ǝ�F_�Yc�m�-�x9!�ґ�y��G
�8ZG���Z�ha*��y���q}`�s�]0^M^��U�G��yb��U=� �șOr�� �'�3�y��TTc\�J��ËE��t0TgO��y�#V�~��1��Í6���-�yR��y�TT�3�.0L�*�ŝ�yR�T�G���6�����i8�fA"�y�	��XgT-�%��O�����[��y2��:94���D�%wfrx+����y�-F
.ߨy(v�G�q��AG��y�k�4T��Q���e�֝�qo׵�y��0d�H��O�R) ���"�y�%�4B�5�s!���k���y�-��>&(�[w옳d�Ѱ��y"��U�q����,Y��P�����y��"�����N-K3�y�h��4�`���ńKf�R��+�y��xx�J琴�j�)A!�:�Py�,f}R��OܹU�h!�U&�[�<AF&�)� �{QfF2):��3%c�T�<A)UFv��7O�4���UR�<��S�%��y��֫P_&�ɦ`�F��(ڦiخ�N}�@fB^�5�Щ"@�4��gH<ɴ�< g�H�I<-��АM.�k��tΘ$1ј�>]�F�[����Ī�ݠ�x�O?D��	"�M.s�Xi+��+T�@�S�M�`���0���v0�H�F�i���G�,OT�Q�8v��	p�*� [d�P&"O��ćdbIЁޟ4�8� �(K����B"��D���Kw��)�p<� ����&:(���&�Y:AG�݀ �'�LY�$��cXnA���7v��T�n�+N䮅�,�6�y�A\e(<����	����Ap����J̓������i���r�I ,�
�>��o�zM����MG�p�X$�5�"D�� n"Gz�=j4�;kI|`i�,`�!p��̓�h����1?�|������.%f�69`,M-5�"��$��b�<��i����#p%	lѮ��c'�@��ZRX�\K��^�A�>��N3?��OB4CJ�o�u IH"TD��'��E�@P%UD9
�Y("�^MK"N�3�j��K�04 &�Ŕdb�2ס��=�Rj�%V�x`	�J�i�VHƪ�H�'�FQ+1�����z�m�+ %a��?��gH�l��(a3I�:E��"e#D���eE��G�:Ⱥ���Pƨq��}ӬI���N'�>���n�<�!�(�k,��,ܙp�pWZ@��U�F�!�؈ ��%1�ע2o��cu��s���
��N�,(��W��:�W?�p��d��"�Q �f1E���K�C��1�a}�D�2[��l��K5'�r�J��,An��nF%i��Qq�"G�D��0��A��L���+/j���3��?E��ҭ;ғ.]&�
P�7u�p�����b�������%!]�|�}r�Ñ1(����p"Ot9kgr��QVCS*�h<#�i��m��J<|JjiH+�'���p�S��5��Wm(E�� �`�j�奋)�yb Șx���mn�j!a��^�����0�R�26�P8��Q?�s����g�D���̡_,*��R��+Ea}��?
ѳ���GU�Xbb,EFh|��o>7�]sP��fFRec`��W���3	�9i��bK��6%cw*ғs��� ꌔERN	��␟�����)S,7/��d��DW��HRw"O֕c��0�nţ�d��2�ű���_�/aV=��@mS\$eM��S�I�2	���*W����Ԉ��תo��C�	  "$��c:��,�E![/;�^�(R(�&�qš�����%§���	�B�� ���.���j�,�BB䉵l*:I �� �؄"U�\9����@2�	pŀ]ΔA�鍕,�Q�8ʑ"K)i��;£ٍHR���E�-LO����Vi��ݠ��A�T��h���P$�Qҡ�{6���N�Fx��2��<�
���p���@V��<q��� �V��W��!_�09X������O�����[@�t9��<O�� 
�'��qR���KXJ����;l���8g��8���D�j<�����ة��'��ѐS�I$\�i������'R(� CU�t�l ˵�ߐ�|�[�L�TtI������×��R)D}�L2U���d�6��Ht�_��0=1S��"[Qn%����l���@�Ğ�Z�09�dT>��d�7�M)��8�A#�O��c�	�v'�1i`�i�Nēq��7)XNőu�M�xv��is��FfJ?�1w �6d �EՆ$e�屡�.D��{�*@�.�������A^�D#��-U�V�(xZ��m�O�"|�BF���2G��C0mJ�҂Db�ii@=D��a���uҲ��q�NR�FD�1x��)���:C�B���a@Lc�'�p-�B%H�s��1V���J�����'K�!�U�Q�P_�lb"@�� � d�%D��I%,�~$�"�G�V�tqs�M;6�`��D��x-�<�N>a��4*3�s��MqU:XA1��c�<	� ����}Hu�ߋ'����e�ɟW��9���鍟]=��c��2U=�dsb$�"q���3�|�N�&�&���r�Y�.	U:�8���!�	��ұ�M@��*D)��tk�Ze�R��dE7:��͓Q.��p�%O#uFFT���i�*��}#��bME�mW��!4H�U��%ԎN`VT��DȄT�:x@wA�)Wdp�*���: t��W���(����5�h)��BO'Oh.�sa����1�|J��1j� �P'�C�N��A�#\�� �O�"�i��B	CL�u�s�
4fԢL��d�/묵3��G}w�AaB%�]��I�4�#��>�jأm�dQ$�ѻN�yR�he�'�@-;4�Z�(�T:�����#�ʨ�4�U�^�~䢠K�+���8��(������_J:��P����Ԍ��)N,��0a��-{6��
�r��D"���S��.�=s�ܱa/��w�T�)A�_�g����H(xĮ���üRd�D���13*��s�<'vࢢd�1��\Q��+�Mc��X\�r MŬK��U!�� �^͂�E�g��ͻ	��c(@�Ԅ`O�s����ɻ]YmP5�	.�(!��J��0.����^*�aƁ)e4�I��P1{��K�
,�8!�TJ����Y��0��<\Đ
ْD���"�)�$Y����R[2�I0WX�3� �P&+��<%4�Jp`�(X��D�p�r��UNK�dǖ��#�X�O7��?�gNM�\s��J�9�$ �<����7SҸ�P�L
�!��?Q��#�bY�% �ÌX>�i1�G�Q�<�{ЇT>{�v�k�kA�V����Q���$�@Ǚ{4�EO<w�՘ ki��x��$D4$<&�<�ϰ$C�z��$��&��NG:� �0��`��	!�N̯3�a~��֛]2��y���<Z��"�E7r�v��� 3"���c�"�Pu!Ca� -q�1%��>����D��S衐�S=}�Z�`Df[)<!�D�Φ�2�j��c�*yZ����1��}Y5j�O��8 ���%�x��ɷ#���$ýߖ�3ɋ����sP"�Dџ|YRn�Ħ������V�.Ib�O�+�bx�g�;�8��	ގl�hCF"��?��" �-,0���.X�=�1kˇ����/}Xt��퉮�.у�� �+uHT�V���`\!�HL���:�z�k���y�Ǟ�"3p�B�Î)m��D 7Y����j��p������Kv[���L|2��εHd�!�'�����A�}0�����F)z֦�����(��X�W�2%Ćb�Ū�fL.̞zu��PMj�O�>��� D�Hb�'��\S�L�&����Ɇf�������$������YE65�`$w�	S�\�p�CE���~��<;&Ŏ�5}ܕ�@�'$H�J�$	nu�b�c̞%"�'�8!Kt�TS�$9R$~$������x����BV)s�<�`Q)�� Y!��vk,�@�*�2���h7bZ�oS�W�����fԔ&_�f�[�V��?���M�UԔȢs���Q
��CX؞Г6B>6V u
'i��L�V��&�4X������9z��}p�fޟL��!_�{2�X%�hP!�ȺYH@B����'�HA@��#U�4Sv�5R����<�$U_��8a�ݵ�x��cA�g�B��4>�&��شa�L`�� C�D@L�`���L"��2�H(O��Mk:���u%8S���TDĊ�O�yYuE�{��b�)	7r��E�����Y�d\�B��џ�@��>�O8�r�� CC�Q���` *5�'ÎP���7 �!(1�C;
}�$'��,C���6�F�xԚ����?�6��+.�l��AȚ��΀,g�(��x]1O�)��
,8� P���Nay��gy��*L����P�'l�q�LE-W�����[�^�{�>:��DI�A��L�q啝����S�qϔ�O1�Л�w����I׭8[��`5˥/�����g�>�اh�~�ٲ+�M^K�`�*LreX �>!�$Ѭ
�ȴ�/�v�����˟�$�Ȑ���Pa�P�E94���9w�:}r�݉v`���<�r�ͩ6ఠkw��Y�\|���ˤP��MrU�O+<i9�d��3	��M��E����4'�qGz⍚1��m�
"y����c��9�j���RU̓y4j���B�l!� ��	,l�湦OB7��c�8��H�� ���"�x@;���|��D��^
�@R��ב]�hhK�N��N��u� �z�ᄖ���	H?�'4��λ�t�	S��3N��T�ï�p�,��.ԎQ2U���@^�0�"�G"�>Q�#�H�d��+�$	�[ ��c�MįbĄ|�rO6}�JFE��!bZ��`QĖ��ɶ VE��}�%�Ѡ��j[>��)�ԍÛ ��<�OåxЦ���ڔ]8�V�ٳ(p4]�eJ���#=iqlK�*��IjG�
e�r!G_�[AD�!�,�ɍ`"��SN"���4��A��%�2�����ƶ	����:�XZ����0NN�E�����gs�m4 	�^:��s
_7&�~9y2�	�-%��''�ta�w�x4AU@G�b���u � z3�1"�'2*�P��&�)�'�p:��]�x�`yc棂=|X�O�����W%W�z7m�a�mi�&.��O�)�'~����ʰD
�>I���1D�O���pA%���:6Xf���D�\�	ۄA�k���ی"P\�ʐCa0ibs�.�2_��G0C�(9��_>U�IK%�\��㞤T&U�	��'��H%���祅�&�YG��1��`�t���5�k�����"§�	�����sV�0���6������ɩk�l��O�p��#�D-	W��p"��w��|"��O����Q�����I��th.���:o&@����0���� 	�͸G�޻I�D��>	`l��������'%�9��"�4u9

 ��J�h��K�4h� ],���hǧ�0�ا�ɛ�2'r���@�*���Iǉ�)�	k�"*����,,O�],y���+g'ā�U%D�8�T�{�L�13���I�}���/θ'���ff� ~�l��kY;F?Tػ�'E������U@��f�8�b�'�>�B�`��4KP��?�}���34$�s��2(� �%fq8�,H����~r���qp�(��m(��&��'�Ҥ#��'��W(��G;BeC5hA|7� ���d���F��/Y &��@*�-
nY��D\u��% �O� L�b7d@�E@\ՂQ�M�X?�x�S�i�,�4)��~2�G_���YS%?D���T`F�h�ȓ'F}��M�,�u(�(�Ext�ȓ9&Aҧ�Y&)d<Ї���tt ���*����y��q���?\|a��,�l��i�nS��Y�`=�P��P{�e�rn�5���dER�3�`�� �!�bF�.�q21n�O
���-��l��kK��l:���N�6��ȓ.��ݫ �wu~���ԏz،d��x:�)�$ܨ_����5E�GT�1�ȓ6nz4��d�3+�<yU��%@�X��43и�G$�	9�*uKBo TTn]�ȓ)$�J�P���b��$S�&���?��P�Ѩ��$��83C�EAm��B$�}a�/��/D|h'�[�ұ�ȓs�(��T�a'�XK�5ɖ5��.w|�ڂ�: .4@��HZ4�pm��d���CU/� `r���SB��z%�ȓ<� T���b���k�AƾC ����a��Z% (Qk-�j�(Q��F^�8s�ʾs B[���N!���ȓ�(��%^�;���B����7�Z���~e<�V���;�n�J�%�:X�ȓV���'�ȵr��)2���4,��ȓL�0��Y<	A6�B`ElE2�2D����.�LK�iS��<G�ѷ�;D���Q���C�ڀ�eE�W�ơ��+<D�����3;��5�&B�)�eؤ7D�xI��W��-Q��]�Zw6��G�4D�(ʳn�D^Vlk����-*���,8D��"��xj��a�ܣvm�Ѩ��0D�,��nL�?�:A��[�<J��)D�TR7G<n��`c��]�
)���;D���eʗ.6�>��@��hŪ`1�O9D�ȳ���	a:*�[ �C�'~H���j8D����
Ц��#w�,-XD��"D��&X,Z�����'.�0tP �2D����Vc�j����M�O�*xؔC2D���#��L��	w�ߒbT2[./D�2�ձ<Bxa��^�&4ԙ�f8D����!f��P��o��h��*D�H�!��,W�Y�w�B�k�A�*D���𧚾�p	s�`��><ƙ�4 'D�I1	T>�f��GȎ�d�����1D�L�Əۇ]���.i\�lz��߅~�!��Ү<d<�wf̛fD���D�4�Py�`M ,�!� �iV����j��yrb%xQ�&���b�B)r!/߽�y2��<x�F�!pJ�"��F��y�J�,>���l�pBʽ8�)��y�L�7)&����,ٽ���y� ��y_�)h�x��'�%�����$¨�yB��tUt��Gڪ
�R=Z�_��y�"Q#�������Ţ�C�yr�(�n�X&��)R�J�I�3�y2��)M����-��"j��BV��yb��:���8)#M������'�������+�OӸ;H�X�'ר���E�,%��-v�:t�N�<Y�"��=!Rpk�m��,�8JGiH�<)�o�Dݸ(��K�}���a���D�<�w	��
� ��dF�缵���E�<YVǜ�%y����m��i�
<A�Z~�<� &�(U�ۦ7 *���훅?W�T�S"O�<����8;�
�R��	NI8aK"Ò�P͞�KCBu���L@�UA�"O,����e�����ǀ@-<9���(|O^}�b��q��a��dP�oFT��"O�1����+|Z0��-��2g���Q"O@=����
���p+N�~lNU8G"OVI��*%�����  /�@8iv"OZ!s��	ƕ�s�D�]Dx��8Oz�=E����/M�L� ��|'L����	�yr��m���$�Z/t��l���W��y��Ʃ.m�y3F�oh�L*���y�I§Y�*��1Kb��x����Pyr&�G vp��G�$�y+2�<Q�].�! �1e�Ts6��`�<a�����B�#��0����E*S[�<	�FF=`��0�ЮЪ���1hT�<�cWf����q ��<�F�{�*�G�<����$h�TH���nU\�0���D�<���(F�h̛b��L�ν됪�G�<�rLN�=��и�CB]NmR�D�<�����f(3�bU����'k	D�<)qh�9���`�A�k�4�� �B�<A @�s/:�x� ]�>�����{�<�i�U�bM8cb���NT���w�<���X�mV u�
0Vh�=ɷƓp�<�毝�[�^P`���s���h#�Ul�<1��_}�4��� jźN�g�<��&v�
i;T�6P\����m�H�<ɲ�
R�􁙤l�4>���Ȓh�A�<�bmS8�(	�I�O������B�<Y*ٳ
�&�!SA޽'� � ��@�<yTB�, ��\�W��7QA�肱!w�<�V�ʨ�ȴ��.'����&��\�<�T쏓)�,�h$�B���HVdY�<1�aW�}r����b2~e����W�<��OC
~�`xiDڛkX�髣dGR�<1�I�	v&��oF�*����ëTv�<!�K��~Ȅ�#q���D �ђ5`K�<qGa>h��D#�f�H$��%\J�<��c�$fh.9�� ��"r��L�<��LT�r�>��t���^L�<&ߦ^�<@�F�Îj�T���K�<��#�1���A�y��Az��]�<�щڞ	]Č��-�By1��@�<yr&H�&z@9S�ǅK���p�UX�<	��U�#sʑZ�lHWo�(��Q@�<�]"3��2p$�7�NȠ��@�<�Ro�<lDÔ+��c�84Zp�[V�<y�aB���� �,�ҭr��T�<���_�z��h��
�i�v�$�L�<�v�[�qixy{p.�}�j9�A�c�<qc�T�`Gt��"&�#i~ A�z�<Ѧj<FX����`��`~��H%�Y[�<y7�\���T�MP�\����Eb�<�+�:$@�!f���iT:| !��t�<��tT�qdHa�L�S��U�<q�ě�5��D׌84]����jW!��qKh`���w�H����	�!�J�B�C�Gє�8D�-b�!�Đ������G�"B'R-Pb�17�!����p�7���	���� �0U|!�ĈT�\�P�͚A
ęx�� [F!�DY/JV��S�V1��6�P�e�2B�)� FE҅�А{�.���F|Ur`�r"Ori��� �\�
���8�^�;e"O�;g��<u��� ��U��Q�"O�� sG�&Da���piS���-Q�"OpLs�5D��m��gT?b�1Z�"O��D�+����DF�x4�4��"O>�p���4�r�Y��[%-�6n7D�<y�Ax�۵ �dd[h7D��@�!C6��(�׭}9>[I#D�\i�%>����N*� �#%?D�� �(	�-A�(�oљm.�c��On�=E��d��H�Rr'�xP�����?z!�d��@D�4���gQ:�!��L�$#���I�D��兜'�!�ڵc��8�K��`��{�N7uZ!򄛐O�r���ω�e�2�{�mOxg!�$^?<�֐��*P��a+T���*�!�D]$<��DI@���,�z�y�(�=�!���߰}��)R�.���aHŰQ!�$^�-����f[�@�D�����
Z@!��O��X�BJ	+-�Vu���Ȋ8!�$�"�D�bjG�N�R��B3�!�D�-\��@f�ƥ1�xL(���?f!��
Q�Dl��Ȁ�0P(5A*Me!�Md�)Ӂ��Q��b޶+G!�^12��%�&o��@���+]N+!��-��q�!��c�n0s����~'!�DQ�gT�A��p�)q�	
�2!��ի7L�eb��͘oY�(��ƒ�b!��V2��l�񥉏g&֭[��ƟSM!�N�H&\l���@u �8Q���d6!�$Z�Vc���a��G�e85$�p!�B^� �� ۷7�����!�D1J�P�� %a�����k�!��Z /���D�:1�P��d�:�!��:YMεe菋��ڇIQ��!�y�R�'nP�Nؼx@�E�LL!�U5Gw�U�ƅ��3�����'+!� "A��5	�ဴ_6���	$�!��]Ƣ���CY-mO^"" ��!�$�p��m��@n��Xp7i�!�D�/��q¡��$%Xv��o�?{�!�d�
?q�P�%�XE,�y���`�!��Zi��	w��;3�LPN��e�!�DFx�<mB6蟇<<��R�0,M!�$�<$��6#[5	�@�E�/!���W\���D1� �rs$]#!��\�X~�P�1��4��"��!�dJ2�Ze3�E�k��͋�"?~�!�DˉN�0��S�M�:Ҿ\p���q!�D�v���@b˙o������2o!�D��k�B�3mI"�8��ǄWj!�d&�\�9q��^pp�c�	 j]!�D�#�t�ǣ�7dc�+/�K!�䙧1T"�GITQTY�T�V;a"�O|�)� �f� fA�X��Yu"O��A	6m�����|����"O�,JN\_o�d��o��|�,�W"O��X��kS"�z��ӆ4{�%�D"O��R.�e���brU�g�Z�6"OƘ�e4"]��"-צc8�PG"O�)R�ʘ�{gY;�l�0w���g"OJ 薭��NY�\�P�M�!�(���"O� ����	��܋@�١�&Q:E"O� ��K&KУ=�8�H�N�tL3�"O���"�6 7ִ��G��p�p;�"O�(Kp�#<���(�_Z`Ÿ�"O��	X�e���R+��g#�iH`"O>�a�#���0���Jt('"O<�b!QL�D�&�k�`T@"Ov�sj!Uj��Y��"��7"On�iD�ُd�X};v�H�=~�5q�"O6�Bp�dB
,��!Y0Pĸ\�s"O���CxbЀA2^�� �q"O��@	Ǽǘ�pmO�F��Z�"O�8�'O�nZ��a�ˋ�w4����"O�Xj��U�|L����w��k�"O�5�	HNf���#T D)��"Op�@g	S�B)Y������	1"O,<Z�UB?칑p��< ���E"OB`H���1�p��
L���"O�a���9W�P0�Ɛq���Ir"Op��$�15t�QT����"O�p{��b��a7�σ)0�8Qu"O����JL��hH:�� ��"O��#�˶'m���Ƿf���V"O,�z��_�\���'�d���"O�%kX=��z�&�
�p=��"O.Q���_ $�D����ۂͨH�$"O�Mڒ�"H\r�x�C��D��5�1"O<�����8�!`#["jP��"O8$KCN�9g���L��y�"O��K�W�-D ����� ���2"O~�
��ʶy� �+�h��X5���@"OHD��A"=^�0@v���(�"O�%�6=��ٲtϊ#h*�B�"OT���.��c\�9�7���A��y�"*O6]��	?v]���H�|���3	�'�P�A�_�6MX�\�+N����'iE�j�U9�l�n���D�J�'6XtUE�fZt�2G�"/���
�'�$���A�7�ᘁ
�������'�Ȃ��B6\c��;DG� ����'v�f���t��t�I�r4��	�'/��"��N�L]��Ԩg]F��'v���$ek*5"��R;�D�'^���mߤ<
��@7����'J�� Q{RT�����0x��' �0��n�)Q�p���ɸH�����'P�`ғ�Еvռ�1)[��B�'���I��Ĉ-��5�qj�]:��	�'a�}AUBf�QF	�iW
H�	�'�.�Q@"\]T�����ȈP��d
�'�lc��_�`*�#V# ��	�'�
���C׆
f�2TR;j����'�E�rb��XUDKc�Z�i��e�'&�����
-?m*h��>]�0��'���*vXyy3�Y�0Ȏ�¥��<)�����Y��fk�H��'[A�<A%���7K�e �K�EÀ�c��<�e`u뚔9P䕐n`|�7�SD�<AbH�v^:�A7�&{."�h�}�<�'D� �8 (1E��{A���/C�<�G��d����ጟit�1��z�<�
Xd�ؤ� M��}a�ՈeXz�<y�K�T�WH޿)��D	��Kv�<A� F��d�
�:��� �.o�<�T����9�3	�(�ʵp�h�<� �݊���<7��YR�?���"O^�;u�5<�A��A�C-Z9�"O2�������^�`�"O��#u׏l�bݱdΔ��|�e"O�`�Ø$%��p��31�P
�"O&��'�ٮ:�����;q<��à"OV`��ȃ�����G��!"OX�f�Q���9�6��_��"Odi۶�Ƶц��t�֝f�Pq"O0�( ��!p*��iP6?~���B"O�����R�����	�eF���"O����l�:�y�FG�OO:`��"OBL�G��kG�`��Gޗ)9(RU"OJ�Xw�N'fB�9�L�4
v���"O���A�ɀ/a,@����9�2<6"O��uI_�9�0�2e%C��Hta3"O���C��_  T�Gk��`�2���"O& � *D/G&)rB�qJ��s�&D��a�ʧe����!B��aOB1�7E(D���ً��tSov6�ǯ$D�,�`��il���ϙ X]+�c/D�x-)ty��/�4Y}�����wI!�$ʒ`��!;�Ȁkv���h�4p�!�D��r���Έ��ͱ0�M�
�!��}�����"C�
�X�Z�C�-�!��8~�z���aܑ��|�F֙�!�dD#,h�p!�V�Q�V]�����!�9msx�k�Zc���T� !�DW0�����c�F���O�S�!򤛎7�����f�6Mn�q5�K�i[!���EϺ�#�e�1uW�B�U�(!�d�+Y����JNB*� f�(!�Di���TG@�h�&N�&�!�V:uT|�Za�W
%��"��!�EyM��o�{���R�Ď.W�!�$��)�
|�Ձ8�2T�DL�u�!�$�<�&�P��b��R�BB.�!�DS7+��c�*��%�E�Z�2�!�$�2�1JT�͹v�$����9!�d6y����9!��r��K!�M6�mq"T�s�,q��0.!���?.��ik̈́W�@�)��޶S@!��/m(�$�M�@I޸���:f!�d��/��B���A<�1����!��e�L�	�OTFJU�[�@�!�$H/i�6�s�L�X7|�	1NݍQ@!�>U�̺V�;>=(����*6!�ؒ��]�dk�]9�e�a�&!�$�+)�i
1�Z���V�V!�Y&i'0�hV#G%
n�5�4$׉=!��M%��H���{Zb��$ʀ}�!�$P�B �Ci��%Ex�Q��-	[!�dQ�y <yI�R#w1\if`O !���,-�� �s@�-#,&�"��	:�!�d��x9�ER).P[�/T1�!�]-7T(;�j��9^����/i�!��<����C�w*fL����&yp!��kv T����wv(�ԍݩsW!�J�<>�;%�T�,�媴�VGZ!��ef�2AG+�P��ỉE@!�d��<8b)� j�6Q���b6!��6��cO�^�r���,��v�!�dɡRD�9���%�v]�􈀸[�!���.1&D�� حR�pmb��܇=�!�� X���H�S��P'.;p�<x�"O�2'G�Qo�cs嚞D[�{p"O���Y��F@hS^�*�"O�����E�(��=8F���<�"OT�� U��)C�#�{唨pV"O����\�+���Bh�+=��}��"O��0.�N���JD����)�$"O�,�"H8+�	��	I2%���#"O��@��D�b z8�r)�7&*��S�"O��P�O7DY���qB\��0�C0"O�!Sk`����a�7��0��"Of�b#��.��8� S�'�=z�"OH8���H����n1h�1�"Ox�3�D� �:`g΢hV��"OY�އ+�歑��II�1�7"Ort���ޢk5��;��Ў3~0p�"O��֢U�=X�ȓ��� �y؆"O�L��N�=��#�����C"O�hy�)��%���G��$B(��"O�	gG�qf&�C`-��B�����"O�pS B�)h�U���X�3���G"Ov��$J�Eg�$��'}l�+�"OF�)�%ȞQ���2 ����g"OF�
�R�E��L�Џ�1l�D|��"O� 	E�y�Eʳ�$(�.��a"O��j֭Q�Ey�U���G9J��p[�"O�BD(M8s?�5�U�Ȼ.J��W"O>1�	�5��y)�(�
HS���"OL���6/Op�J@(ӍAr��"OƔs���p؎8�Sg�#�jUw"O��9e��]�$)r�4y�$��"O\=H�g�%BT&i�0oY�J��'"O ٷc�?Nsv�Pm߷3ȼ� "O�!��73�v�x5G�Y��"O��B�62�H��#�BGHIH�'�hܡ`��b`��-Q�Cv)
�'�|qP��Ĕ:+�D00�Їq�2�`�'�zE�C#˛J�E��+Gq�]c�'��1�C�*hH;q���|�[�'�v�J���N���Z�NĤ`;���'�X�u�M�N�P�A���f�b)�'�)M.B�00 c��<c�'ƠT����~sPk�Ѽ�~e��'O�d*U�u<�c-�$T(r�R�'�F,����;z+6��ɚu��]I�'(�$�a�Ũ1h�+�H�=i���k�'B��p�l� p$��(��iexջ�'�ư�v.���Ȭ��Øh�A	�'D�x���?jd���O�	�<��'w:48���+D����U��u��'A}Y(� �����H����0�'h� �m�9��4h�!�
�'Tf 8#�U�-���X���-����
�'JTd:V �9R$�Z� W�W�,K
�'�zP��#Ԯ���*�R��	�'Se ��E�,�!�c�:B2�!�'Yd�{���I��W*_55^p���'F������6"��@���#�=�	�'$-+T�N$4Z�颶�ձk`4��'��e�2K�b�� �\d�t�+�'�$���N�2���%�`2��'�6�P0�U:}7T�q'
;&��*�'dp���'�u��C� Y!�*��'�� �f�w������b��� �m��C]
�ic��n0L"OlЈ䮋�P�PH��A��8��p"O��¦��+����L�	��5 �"Oz�z���p��]z#�C�\���"ONT�&�<c4�]��C]�z"�!�D�=���1�եX�\(���!�Ċ�4��������!Ԧ�s�!�d�7=��%Qt&�d�1�D�2�!� %�>�K�\Q�.X�)˲j�!���Ua�JG(@X�5ɇc]S,!�B�\t�u���?B&a�C��Uq!���S���թ�� �mb�7iu!�䛄e��p+�>opɖ�ʊs!�$�@	�tHT�	�U�b�@��@]!���|��xY��=g `�j&�F>!!�䂵y�� �G�a��tqV�	&!�dڸr�LՆ]-~�ňD�x!�D�$0bF&C5L�:1{�iQ�!��4
f���GnՒ ���&�ʯb!�ė�zf�`7��q鲩J�J�V�!��I\�[���0W�R�*��Ƹ�!�$��L�� �7n `���:CS!�$��qDS ��,�fX���D	k5!�$X�:N4a�/I� �����Ɛ)3!�Ńh0lE�'�
E�*��f%M2@1!�$�;G�Q�:��LKd��<A!!���?L]���)�Ȝ�F�Q!�ċ>Km2��e��e�����N	~!򄂄i�^�p6J#.��dq�g߸ ��t��(�:\P�F���e	�*a���!"O�H�A�Wh��ДE�W@�т"O���A,ʝ���Y`��E
(�"Oj��oҋD��(�
TS)l��V"OQ����_��b�KI�	r"O�$��Tb���>Q��ڃ"O$�]�=�&�� �v�"`͂ b�)�'b$P�!@l�L���ǉ� I�$�'P�!戄:N�����).#@���'���/���b�I �����'��T3b�?YHn�)����,Z
�'`<��7c��t�`�P�/��Z�'Rz��g�����'B��4�I�'	��%�V�`�9+��$x�@B�'�:��C5+X�83�Ë{+�A�'�^���A6, ##�@�f3�]{�'�T p�AW�E�4�s2]����D4O>���٣f#t�	��I��"O�x�hI�O������E7
�"O<���cN�a�cе�`#�M!�dӓ @J��g��2P6���k�%�!�$sڠ1 �@�FN���+g�bO�X���Ld���S!߄a�:���"O��0������	k�J��^�dX��"O�(�%!f�$ԩ��l;�P�%"O��S��-�(`��`���"OL�� 0Nz�LSZ�8���<�y˘�iE��3T P��8�(�e^���d:�S�Ou(E2�:'�\d���A4V�)���xR��
;9�E�e玣x"�!KF6�yeZ���Ɋ�Hm�Te#���y��K@0	a�>e�6��w,���yB��A4ęw���l��j�ݻ�yR�ҖJ�YK!���vzͳ`Ǒ��yRڏ���� �c�(P�Ε����?Ɋ��� v�!�Q�r[�ԅ(,��%I4"O��@pE�N�,��&�R	i(�{F*O��2��2zr|���Q�߬���''������.[�1�SH�<��,z+O>���ǵo�X�Q�o��G�4� �Dٛ)�!��J�ɳ���uz�9����!�$�
r�=�TLX8cލ�F���3�R�'��O?ɡ��¾T�m����E
`���h�]�<!���s�(A:� �6h���m�2�yR�%/^d��q���.M"�'�"��O4"~�B��5̲���O�F1lm�uK�<�f���ubx�oH e`*�3q���y2�Y�ocV�3��o�4}A �y�c��;Lڬ"Ԫ0o5p�0Ņ��?���,ړ;������C�~Y�����\�j
�'�����D�u�B%�����
�'��0���
9$Z��[p͛�- ���'��Y�W&�"A�`*@'�z�\���'{���b<�98��M�H�a�'�$��sK։<��Y���$j~>��
�'ۂ����R9c�v}�u�+^���
�'��mF�Z�nJ�2I	�1��!�"O�L��`W&�ĠV
V:ieVx
�"ON�D�ҜI`��Ǘ�L<-��"O`tC���k�Ziൄ O-�M)"O���e�٧���z6�+g)�lB�"O�
��|�4�2�Z�8�Q"O����r ,����d�<�Q�"O~m�4KX���``��}�x	!�"O�[��5yF��7K-v��!�"O���Uǚx�)ٴ�D�(Ϻ�0a"O���`���9DH�UN�
W� �6"O�Y���'{h���D�<R��"O���dҫYd]z� �>@�Z"Oj�!�^�[l��-�f,؄36"O0x#�/�1cd���=j%ޡK�"O��Y��� ��2FdݍL����"O�@h#!R9"��-Hq�K�eQ�"O4�@A͠*P��S	H�����"Oz��Z�c8�m����-c����"O�y���b�v1� #v]�:$"O4,(2��	Y�����֬X�T��"O�1��)T�vpp��/�(D����"O��g挀#`U��Z�|8�D�"O �)G�_ Ev�]�K ����"O�*�M�x�b��j#`X:g"O�a��$&=�ȃT�Yg��̨�"O�P���Yg��,T�E�>q��"O�
�닒1?L�)�BC�̀P"O��%Gئ:�:Y�5c]�T0w"O�h����&^x�-��BU
AJ"OB�
GKT�;�d�%�� f/�G�<ѵ"V�X�� S�N�V�&I��+�~�<I�ɛ�b�^��a�A`��,b�
e�<��Y�:f��F�R/|>8�a��k�<i��$M\����O�p)����Q�<A�J/�@�`�<|'�i�/BO�<��'&D�|	tb�>>Q.%���U�<�$��K����%b04��a�Tl�<!`�������[�G���C3a_�<���B1
C����&�v(iR�^Y�<��c?B�q��F�0$�Y�<����@�4�b-Տ
�b��T��N�<!@�Q5[Zhɠ�N"	F`�v�U�<� �U�B�3B�z̩P��j)��{�"O��sJن|��EX5M��`$D�@�"O��a�/#~
D��]N�ʷ"ON�rvL�
Xpx6j� �"O�I�B�F�g�*(�'LN�"��"O���
!zyd��3�z\����V>m�sIߪ��H0��;iBr1A��2D�Ĺ��@�;���)6� ?5r���M1D��X��"��I�i��)�х-D���(4:��Z�#Y-��,�6J&D��Э�-���`�+D�l:�����#D�����@//!��oŨ:_4����"D�Ȉ�j.o|D�T�A,�d�%�.ړ�?��dV�B����&ک�<rF�	�(JB�I�!ؤ9a�J�w�.��̅�CV�C�ɌTPZ�{fFU�e0|��ߪ;�tC�(FЈ v@�!{��Y����t�
C�	��FEq�O�3Z̹���U��B�I�_����CCO���%�xSrB�I��|�ّ�)*�TMC5�;:Y^�?!����*(D%�e�Z�?�2�0,Se�!�$�'i��|HfZ{PT�B�ȸ=v!�$I��~hs�؎_^���G�!f!�Ā�X�	h���=U�١�]���e��(��ܠ"�Ʊr��E0eõ�t(�"O��B���o:I �$!��l��"O��Rnʯ�U';E��؀��'���4��Y��4�d͍*7�4��P�/D��H@b�&,�� A���T���#/D�p	��*"�xȐi�.w&}�,D� [��Ӫ@Xt���4�
%*G�>D�l�R�5��l��Y�v��؂�n7D�� �A�r�| �AY3R�8(f4D���Q���x"9�d�&MU� ���3D�(rb\�;)���S8K�D,�v�3D�`�P�J�06��O�0'>���/D����%̉8�`�;C���M#2pJe�.D��8#	
�#����4��L��� �,D�1�����[��^%z����)D�t���U�#�.��S��^�bY�B"'D�d���*#��0���9yT��'#D��HƊJ�#ʾ�HfPΒ�Ӷ@5D�,١�������-˯�.H
 d0D�@!0�*,.�� ��~d��Z�/D�ԣ�'��x�׬ܟ!���ע/T���'$=X�lB���R~�(�"O�U�@/F�pvj%� �=8N�(�"O0��E�,V$Pr�	�9U,�Uw"O�����M��f����C�_2�a"Ob=�n��9�"i@�	�;�TYg"Ob�M��?m�d
��;#� "O��4�-J��;W	T�g��� �"O�[�i��('�%�e�]7��"Oұ uGٌ+^�K#H[�3Ҫ�S�"O2��O�-1�x��c̣L��p"�|"�'�F��a���*LfPk��ÃP8ja���x�B�##� %(k��\�r�L�y��	��9+S��4��<0��ƾ�y��į@RE��O|O�+���y��4Y����%1p�ʉ��ޟ�y"R�`�����:d<:b0��'�y"�A�	b)AB�\14�@L��B=�y�Vze�X��8 2��-���!���'n�b$� ��	(Ā�i�1#��� $��R�]q�Hiu ''��"OA�'� 7�������(:�V\��"O�X�d͇"ӆ0�������|!�"O:��L-I��0��Et���"�"O&����M(Z���â�Tq�m��"O��b6ADZ����A�8Y��0��'f�ILi,)�B�V�Vg@պ���{fB�ɼ�\(e��:yT�@�Ġ-5PC�ɛ>�V|�J@%&f<��D�þS~DC�M+�-�W�:��#p��'@�B�0nAhmzfb_�,<�uR3�)�B�I�x2�a�1�W�|���PС�{˨��0?�a�O��N��ߪu���S��T�<�ć��.0� :GK�%K��R@�M�<�ÂB�~��0)W/^�XH��qU�I�<�2+�A	�O��Ct�i��H�<yEFF�x���sf�ŇJ<���b�G�<IwM���"�U?b��C�G�< )��>��`Z'ZD�nd�"�l�G�`����7�hIwA���p-y�'D��{�F�4i�`�$��I�l-2�%�D!�O���B̒&k��!��#�R30"O��ZvbPW�(�"���^�6��"ON�r3�F�e8���W"éE�����"O�y�Pf������9P䞑C�"Or�	DX�yb0�R�ȹM;
�*��|B�'_Lɠ6 �/�V��CX� �ݰ�'�r�Y�p�q�C���<���'g�l�Pe�=��a-�7���
�'fH��H�9`��(tj�.���X�'N
t��e�9t\|������
�'�B��Ʈ^Ț��)��6�+
�'ݬ�h��ɹ:��I�,�C�h�a(Of�=E���sZ��%�τ	�`���\��y�%K&C�(�y�L� 4�����<�y2�Ҏ#'��%��JX0O�5�B�.a������+(�ؤ�TĐ�N�@C䉌t��iq!�B"��C��l�LC䉠F=c���^��KʈF�C�)'`^`Q������G�EF�D�O �O��g�':p8��&�$|<�!l	)C2Ѩ�'r�R���qK����� �q��l��'s�Uk��$t�yt�zR4p{�'G�K��;G,Xt���T�'���'wR5�����1!���U&�i�'�f��PbȆQ=�\8�͊%�M�'s&!2����Y�^�۱L�-'x1����d�OF�S��{"Ђ)�dU�$,><(�� @�;�yB��f'F0?L�פˀ�y����jH��EM�)/}�y�v��=�y"�N9$َl�G�Y��	�n��y��w�R�(E*`���L͉�y�����҂��c����Ⱥ�y�i�:�J9��@Ǝ=�Zq�f���'�b�'���A��)��I�3cP�
�ɢ�'���u�X�.�4��gֲ7R�8��'�$՚��H�b!��E�'�v]�E�M������0�Z�'�zm)�M #S�[�%Q84� ��'Ŷ$� !R����B6���']�,yt�E�J����sl��7an���'i�\�TNľFzE�S��5�ft	/O���,Z���)wI�,T_����k��C�ɨ9�	���+h9�\���˓EҦB�)� �8P`�;;=���
�tHF+"Ob���Q�&�sdc�K*��J�"O,�8�=Xꅫ�"K`(>bq"OĕH1M�VDy㢠�,2#��^��D{��)��t|l���� �`ʢ�N�K�ў�������5,V:\�\�`�U��dC䉽�l$Iu�A���4� ��-�`C�	l��E�]��&�A,Q-�tB䉃[�:0٢IC�gD ���D;;�C䉪J�zeõ�
3k(�L�3;ҲC�I ��U ��T"�Wl
t0�C�I9S��I ��(E�0�ĜW:����q�P�'c.�8aGƲp�聁w�A!L���	*љ�" 4���a �uY�9�ȓW�Z��iՋmZ���@��(�ZQ��>e>�DhP=9��	b�(��9��n�2H2�C�A$���G�p�-�ȓJ��nI*3� `a��D-s&h��	@iJEۆ>P�Bē�|
���2�ɠ*�ƀ��MZ�2Q����zJ�B�I�9���!AQ/a��́��Xb��C�IC�N���$wp����O+�C�	�Zm � ��V�c>���$�߄\rB�I0� U
D/@!B}�i��Iû| NB�ɞkpNP3ɕk�J!�Q˅�*b�=I	�'d;޴CS+ַqDFp���#34�!�ȓ*�A�I��T�@�)��%Q&<��ȓs��]��S�K�֠�V�ݠGaH	��D#�Ar�
](�zd��V�q�TلȓD�TѸ�-��K%�%�&�	/\V���ȓk�x�C�K��˰�Y�� ��Q��l��I���պn�b���5o��5��NA��I��V�vڒm��E�<�jy�ȓaC.��G�s.Q�!F�#g(�ȓ}��i�bcJ�p� IG�Dm��U��xm�sa�-tٓ-�,9Ҝ��0��ܒ��:ܼy0���e��ȓM��j�C��lG~X�A�G!S<��}����'r��1�@��'S,X�ȓ��	�+Civ����#[3Fޒ���I͟��<����930�!*��`��b�<AV�S�T&����)�%g�D�c,�V�<�E]&��AA� �n������i�<��(�
*�Ԕpd��W�z�2�c�<م�����s�ʊV+d �roUF�<�'U=�4	�/�+�Z�����C�<	��_#:��K
_)	�v�z��B�<1H��0�{�O�E�Ԍ���c�<��T/iwx��3�]'GpȰB��\_�<Yw� PPN��׃W	^�Ґz��Q�<�pH�d$r�J�k���`��I�<Q�
?�&Qb1�S�W�Fm҇�k�<�A���LA��:=Z��B��m�<y��V8����2$7���3͛l�<����?����ɷ#�H,b��d�<Y�9�44��F�6����"l�b�<���1Z�Rb��*%��	�Ãd�<�A��E�`��I�(x���x�<�㡏�I^2���/j0�h���Z�<��-�r8��u�W$5� aF�Q�<i�F��Q�¨�6���S:T �6	�d�<Q4-�G��aia��/;��k�	H�<��S  TAa�#��XR
�3TK�}�<	�
F�{���=L~���D^�<� Ā�3��. h� w�Ѩc�Ұ[P"O�5�q��X���R�T����7"O|�7ES<NU \��ٱ۠�ss"O����

'\Ē�
G�) ��1"OH��-|�l�Z�(G�,-�1�"O���a�N�E�W�ג}��s�"Ov���D�uv i�@Π8.%"O��&ʢQF�!����t�d�P"O�tlֱb��u��YpK��y�,�.d�S��Z��������y���1j�$�`q�ͳ&��q ��
��yRa�0cL�I������P��ۈ�y�'�?o�@����վٰ�Z �y2�/`� �1akK�|4"�ؒf��y�m��r�v�!%'��m"�AJ�'�
�y�I'4&a�A]>SeZB�iT9�y�"�4��;S��BTv�y����y�ɜ?*�R�!���BeX�k����yf���� �ǝ:'��`��yү�B�QP���|�)��C�y�J��d��DÙs��9%���y2��I���0�҄i���2%�Q��y�+NB�d̢p9K�1
�S �y���+��l@�"�?ɂ0�QdǇ�y�aE�[�@X#��e����P���yҧI�M$e��ꂰXQ$�)��=�y¥�{Є��F�#Uk|B�'�*�y2��+
:�1���J)"�B���yÒ�<��}k�'K�G/��q��E��y��� ��ES C�\���\�y���%\�d0�@n��?v��be-�=�y��H\�ԯ�;��	V"�y��E1r�Ҍk'85^M��a���y�����f.�)�`�{3���yR��`�hi(ǧJ(x�l�.��y���q�x�#i~���"H��Y!��![wv����٧L�LEb5��#-!��;���+�FX/%��@2D��1:!�䉸�NPp�V�q�@��ܮr#!��ަ�N�"Ug�����jp�_�:!�d��.�ɠ0�b���tMO!�dQ<>8�IG��Gˊ�a��R!���f怄�sN��r���V�i�!�$�12�$pר�'9w��T�L�n�!��O7������;˴Y��ɪ(p!��1l�Z#Í<7U�����M�;m��џ��?E�aZ�'�b͘%bS�$�D�D%۬�yrEI#C�0肅�,Ed�"��œ�yߢ#p4� 4\8
�Y¤�5�yB��R�<��K�+�+b��O1�C�I98�ŒC��%r��#��]-g|�C�Ut�l� !�bq���޾��C�� �l�f$ �)RQ�\+b�C�I2�L-D�ܷ-��HI G�(	j�C��}����nC+A���t��O4*C�I�����Ώ�d��B��)8u\B�I�Z�ڸcv�
�Dmҷ#�^	6B�I�n�@�@7�#s8m�t#?��C䉞aFUX!	�i�L]���N�"��d�O��&�O�苦��VpB�眸m"a��"O�J���]�X�6�;}iƀ�"O�<;���L+ ��$+	HX�8��"O��rdl`W��	rM��Tɮ݅ȓl�d(b���-�ƨ!
v��T��S�? &ܩ�FS�G�T����?��ȡ"O��ct �F�S��L�f�g�'t�	C����L�H ��x�# �vM�H˰2D�|�怐j3��K�ΞD�h%2�O��NM�p:�o&8\a�-H�I���ȓc���#B/S� ���� Y�H=X��ȓ g2лt�ʥz�R�X�Ҏ_\��y��k@�X�
��t�g�G�%!6l��b�f���蕅M#d�1F���dz
��'���'��M�f�܅b4W�}>x���'}4)S��^W� ���(s�$�*	�'�ơ���;$,�Y�R1h1(�8�'�ztˬ84�G�C#f�t�'���ᓯT�'K���,Wl<��p�' ��%%ߟu ,l�&�Q�6�	�'�.A˵I�-3�h��Ȇ2�و�'�1��/O�8 ��T�ɑ%&��Q���?Olq2�8Ut%�R�-I��Z�"O6dѦm�� ���@�3i�S"O@����N���T��uT�`"O��iÔa��U�u�ߺG#R ��"Od�A��S�*pAE�rĂ�"O$hsE�1a{^�w��78��4
�"O�9�e�1J9y���e���x��'Jў"~�O�~�|���
�l��L?�y���-7��:�'2vq*+���y���A])�S.� @vܘ��M�&�y��o�Ε�D��n������yr-�*	�e����a�`!i�f�yR	�"��ђᄒ:n>�p�.I7�yRcN��p���iZ��r�N���)�S�O_МB\*r�j�㵬CLc܌c�'���(WML�#�� H6�ۇ=���'���Bc�^0b���f�~�Z���'�n]��y��<X��%�J�Q�'9�d��M��S |��4"�%�n0��'1�dcbZHq���ސx0��'����̘�)R\E�	�(	^|����?���i�60I$,�"LB&;��B̃�f�C��$9A�������-��\�i<j�C�	�s%4����pk�|�� JjC�	+X�bY��L�<U�����W�&9@C�I�{(�)� P��\ңL��4�C��w`�v`�'iv�PQqE�[4�=��'@��hADٝ��n�O�N��IU��Py��� %�@|م�'7T����0u��B�I.5C�+�7V����Y�s3z�O�����ZHr���!{���"O�=!!�Dп}�*	 p'� ��ȵ�B�H!�$X�� ��n�L����*Z!��HX������FPx�ƶK!�D�N���4l�'D��v�[�4��'&�f��~h�cCh�� �a��0b����Of#~��@�/A��I�G�ɋz�.�se�{�<�����'�"l�bھe%�Ы�y�<����\4`kA.�<���y���~�<�'�p�JPzf��'��\��-H|�<��`��i��B'8"�erF �b�<�e�s_*�M�9����`�<�mٰu�xpr�֑\�}��F�<�wi�3\Z��X�Ɗrr@��'J�I�<���>&٠���Kщ���b-Q�'ha����D�!��N�:��  �]��y"a�t$Z�ƌC�8�,԰�i��y
� ���2@U�	�hD����>c,Af"O�}h��
3 �L���eK<(U����"O�A+����O4��
�"WOJLi&��v�	O��A5*����M�/��Ih1�F�y�@)2�S�]~Tq���&�y��B:C��!�K�<�*F���y���'�� ��µ�R:��;�y��1���S L�|^�!�c���yR�[+0�$LcU#��c���5�y��,����lA*X����Q(�y�̝�l��U�шQ�9\r-Qq����y2k�'A���vfې5+&���g�y2�K��Yq��*�t����,�y�f\,
*k�'�
���%ؔ�y"�;k��!VK�o�b��G�ÿ�yR����	3�b��oq:At�]>��=A��?ɚ'�&�`W_i[���v���5Cܨ�'uP�C&.�I�H�犋&1;0�h�'��'cAK����F(.�.�
�'Pz�$�Űj�`�3��P�����'��D�f�/3�~�1�ۖD����'�lɛ����
��5%3D�r��
�'v��j�kT1ss*�ŮVH�ƕ`	����v�����
'�琴h�*�� �8D���T�O�k|�	�F���`��f`6D�ģ��M� Z���ױ`v�4L)D���f���] ϙ�|�n����%D�HP�b�ƕham���b�X`�-D���ď-9ʲ!3��9�R\k�6D������#)��P�%� a����WD:�In�'%�4O&H�ǟ/g�p�"3Y5��"O&�y���(ks��2F�
s:H���|B�)��"J�H�`C[1V��LХ�S<C�	j�F��RȈ�m�쬩�K:~1JB�	1
��\�����!�
�z���x�B䉫$�U(g� �[��U�r$��'� B��+�N 
3c�Y���)D�46��C�ɓL��]#�k�7p���4�
�=�ԓO��=�}�țk�<��f������Ɓ�s�<a�dY�%��сB�Y��ĚcZW�<� ,��t4 )��R�T��DRS�<��$�/v� �U̒wǶ�A獗M�<�Ł10��Pt��B��	�J�L�<���J:.8~��5@PW�h��`L�<����
�ڭr���'!^,QP��Ky�)ʧ3k�xSN�DY���}�h��00"EkR��,��Q�ċ�9R1�ȓ*�2<!0�Н1VP5)��B�-QE��6w�:�Ő�b���x �� �K4D�ۣ����+�#pV2��c�<D����߰x�J��7C�4u8��6D��5�d��c)Q.�EÃ�6D� ����:J�<�R�
�a������9D�L��=bM�@�'[�N\�4D����m_�-�$����,I��N.D�@���Rܤ��cC�V�(X��1D��P�o�%�5q��?*��u�0D��
4��1?.�&ٍG�p���&:D��i�i�cD�����N�J@"��;D��PQl�'xL�Gl[T�:����+D�H� D�?�,�k��ۑ5���T�*D��Q%�	.E��Q�W��;��ղ�A#D�Б�$H&v>� !��W��+EI,D��Ñ� ;Hxf�zR�� �t�"G�(D�� j@뵡߼~g$��!��$ 2��b"O\�Gɖ޼�sP��9�0�$"OC"�'b��K��T	���g"O�L�T	ĔBE�H`+��|"<�2"O�m����63,d(r)�n�,H� "O�ps ��G^J�hP��; t9��"O^��g%͸ ͤ���h�8cSV�)�"O����Z�R0ȣ���$��`ag"O`m���) �P�&�E${\x6"O��"f�� ��!3X>Ax��"O�I�4m��3�ӌD�ڔ�"O��� ��J2D�2)IE�<��"O�U�4�	����۱�Hـ7"OT��en�>=�N�;F_�Z�<�Y�"O���Ń&ZFn]���q�6���"O8�Ƀ��e��#a��[����"O.m1����g;�]C����|�{C"O�K��H�����S-O���Pr"O���)�:m��Ms�`�\�����"O&Q�/�8��@Y⮚�B�Z�YS"OZ�����g�q#�6z����"Ol0s��[S�8��,>'�|L`�"O��{gH66n��4�:\�(�A�"O~`rq�'!�̨Z��S�]�U�r"Oh�a싊HJpA�"�Dn�L��"O�+��K3MOPhQG�g��"O���A�q����f@XМ�v"O��SO�/|ސ�4��\�l%��"O�YUa�2g�Z� #K��&U��"OHL RB���R����g���q"O���T�)g���2�)�_��)�"O|%1 �3�L�h���~�����"O��yb۔B�>��lN��|aV"O4���Φ�|�x�j�j簔�G"O�h��J�g�<�����|��"O��P�o��[�8��H [�A"O��3�'J%?��8�5��1f]�Xqa"O���&ժ'�p@�C�/z~p�'"OzI�`�MZ�Y3P�@�#z�]�
�'�6pq7%� Bt�l����;���'�2��kT?��
WK۟;Q��'�����'�	~�6:��Z�A��� �'�43pd��d��<��-�N�Mi�'�੢�C�6>HXQ�ȷo�t@�
�'��,)�@1L'��PE��:g4*�P�'��uh�U#!iB0����z��'�!ץ����@c⁥a*����'� l��(H6{Ӽ��"m�7%�|���'l��@"#P4A��,B��jD�UZ�'i��T�ҝo�`���*��N,еi�':D�z4��H�C�W��5;�'>��P3b
o�L�AgO>^�%(
�'�)�p#�_�"��PfzE �V)(D����ٓTR�����f}c��&D�\�HH���p����6@� �p�%1D����GN�L$���p�Y�ڙQ0D���QiA4}�@�� _p�ٛ�l:D����K�&r~�hPr��.
���k-D����jݗ��Iq��{4�A���+D�H����dC2��ԋ(+�BІ?D��)(b�����R�
����"=D�`�	_73��yG9c������9D�d)�%�&0 B�"k�z�d���9D��إE�;�p��p�W#g�6�H��7D�� ������� �H��i��S�x5Y�"O�QG/ȸj��g(F���@W"OJ�r�ǔ �8L(J'c갺E"O��qCKD)��8!���Ia2��"O��R���[���$��#cT@hb"O�(���yD�ѡU(R��R"OR�7k��C���s��Ī\�)!"O"1�tE���"$�E�f&��!"O&<�¬�->���$H=[���"O����%!>b�(��v(���'w숈 ��	h~��7��E���'�nm"�	iy��:���(3<�)z�'������_�B*��h�lUY�M���yrb�+#D>ɢ��.
(��B�C��yǇ �z ��A�~bz���^4�yB ��U��	A��>Z D�dX �y��Jb�I��hŌm�ƙ9�O�<�yE�ߪ��@�ݠuz. �K� �y2�������	�Y�ͣbl��y�3�J�㔧��H��ay3Aˈ�y����4�����@L1� ��y�] R|8�F�65ƤH��M��y�oʻv�V� �d�<)D S� ɫ�y���RW������'��Ҵ�7�yR���M޾���*�������y�n)R,�ݱ��M$m���m��y�*��m�"��?	�2���ɛ�y��J,� z�$�)rb�j�"�y�/�^
��@�шh�n(r@@��ybn(�`��R�	�ru� ���yr+ҪJ�<�;i�&~�*�r�M���yR���3���qf�y2 uei#�y���,�0��g�	�z'���Q�y��8)��!�#!|�j�ߕ�y�E2����A��\qr֬���yrϜ�MOF]ɦ*Ƞ��6��y�_�%�<�E���*, ȕ�!�y��ڢqv S���}�
`t���y��=3a,q��O�D��Y3o�:�y�茝f�~� @�=JHx�d��yr� s�2��ԏI�	�(�wE��yңQ
	��st��
2�K��3�y"�8װи!��6i�/�y�ՄXP�ǅ�8wA04�D�2�y��/�F{��ֿt p!��-���y��r��\�Eဨ:e i`�4�y"l�%PBڙ"&!�';BSӊ��yRC�.� %�@%�0.� ��L��y��	% i�1�Q��F�y��I�ک�Ǣˋ&JHyR�y��Q�i_�A%F�u�4��l�y"�7~�l�Q���1�`�K-�y��2j���@�:r���w͏�y��?;�*�ʰɂ2r(lBkH�y���|����\=b��*��^�y2'�v�!�E�go�t�3#S�yb�����I�F�n�	����y��\���u�׫j� q�����yB�F�M�|�(N5jV�p���y��A�'�,�i���1T"je<C�I�/<x#E�]�=j��߸E��B�n�q�3O  6PSwS�B�	�@��A�Ď�6	��p��#[#B�I)lC���ŝO�M�振C\B�)� 4�;C�G�O �ySA�1l.�d�q"O��+��F�/=�Ț��.E<%"Ox�#�ܻWK�%CPĀ�c�	��"O����ʀ[�~dHd�����y
"O�i� �{止� �2s����"O�	둆ʖ�{%jμP��"O�谳j�<Y��)A)����"On�"!b�\����ƈ9��])�"O^R	.�HS �ŀ{5���f"OԜ��D��bP�Ϗ	w����"O�xp�]:@�͐�o!G:qj�"O�S����P�^��h�>x�\���"O�B3��H�xg��pYb��D"OT�@P���)nv$zT&� .J��7"O$0�1aQ�X�e�q=� ��"O �W��G�r12WgɹT��q"O�=�s�Q3���P&�*/� �"ODA�^�@������:�5�+B��y��\ V@��B����$柤�y2�D5f�zb��^����W�a�!��gG��6��xv�y�lR�E�!�D�+>�j���"GF�D�^7�!��Fz��wC�8b/����ʹ0!�$��(�I{U%e�q���T�?s!��t�0�PF�l\�{�hL�mq!�$��\E���Th���PeH�(!���yۨ�@tI����1�){!�Dˀtz����_�D�N01�m֮<h!򤝋0�Hy����9~c���U+Q/99!�D�3l ��2�R4D�i��M�u!��$&3z1��ǺT��R��3�!�$
�@.�x ��c\������!�d�n��Y1�K�xl�p��GO�!�C8d�(�[6�	&UW
հΔ��!�$\��� �CF8r"��i�K]z�!�["��qʃ��"(A�+����'F|;Iֈ:x� �^'a�6͙�'A��p���l�`P�DOͽ['�!��'�&��Q�o��d)���[H���'B�
�"��\'�lb�hٖS�j��'QNhqfW><�D8@�LSF�:=�M��m�W���0���z�;��
y��<�vc5�OP�n��1'ꅛ��x!#ςC��)r��d?�>��	ڂmx��cH�:e�J���d�b �O��N=?)c׍޵0p��%☄�`$x����4�=����O�20��6E��0�Qur� q�"�S��yr���6�7��rlh����y�aGw�"lsp�ԍ �r�k҄�	�y��ԛw=|(��$�mSh��iR��y�aI
�3$e�c4��#��D�y�
N�V4����Mړg,����՘޸'�ў��`k�	�,M����!k�S���:�"OD�� ���l���vI:V�&Ty�"OP�!�-$1�O�1-@���1�S��y��,_i�1�͵Ea���S��y�k�0�����.��)xg��y�@F���+�-9�yr��y��?](pu�7���'?`��E.Z-�HO<�=�O��y+vď�8h>�����7=Wv��	�'W�Y
'.
�BM"� :@�d]�	�'�����*�Y8��ӾdƬ�	�'<x�p���.;G�h�Al	ZP�Q�	��~��/3�I�vDJ?�P��$���y�`آ'kx	�ጟu9u���ך���hOq�� �)-ןԸ,AǊ� k��p"O��bG)�+( �hp���
@~� ��"O5sv�S/ad��qŐ|F`j��|B�'1�t:���<�4z�/�ʞ|I��$,OL0Ƌ�Id]��kO]4PY"Op%q�E�}�d}#���3�~��"OD�Re�	���s�iI0�B�x3R�tn�q���O�~��6ˊ$�������Y�j�'>4�V�s<��H�)UZ* �'�a�&w�:-��c�,W�ѩc)ݚ�y�,�+:]�dܿ"��&��y���l�B.X6����P-�y��"�����e�$���K�����yr��1~m ��m/����)J�M{M<鄧�>%?�O�Lcƿy�Ȕ��.�<��쀳
OT7���p��ubƥ�"1���Ɔ�i�qO�=%?	쏱!�p��DŘ-��02@/"�?�j"}���aV��4���Hu�R�Qz�<Qu���m��0H��DX4��3��y�I�A�Q���yҬ�1'����˺k�A+g����?yp���x�j��J&��г ғ:��!ʅ	>��M?�O>i+O��Bq��sd	�CI\09��#?с�0�u���o ��Dk�am*��&���M��'b�	a!�!��)E �hV<����O�b����$"�*��NqP�-Y��"ĤO����Q�a7Ѐ���,9��8r�����!�Řp�T��e��?v���bT�$�!��Vv��%�a$�{��HV���џ�F���͡�.i1��X�<d��1E����<aM>E���>P��1�B��A���C!C8�y��S5[om�"�reh� �B����-��Z~r-\�T�[җd/yM������8z�'-a|�n��Z[h)�7�S���1 �K��HO��=�Oޖ��w� .ol���i�oY4uh�'{Z�3���@ �� ��(I���7�S���)�x@H�Mv!���yb�&�|`i/�p^�P�1M�>ˡ��:j��&̇`&��13��2z�$)ғAU�&�D�=x�L��o�UL*���B-�'a|��J8�ra��?��ڐ甆��	Z���O�$yZ�+ǠA� !C!	!=�ĩ����'H�<b��pg�ɂ@�5<*���'�@�o؊�F��7��8�9�
�'8M���<�4L�P���
��y�� }�@���� �5��o6ў"~�%T6Dz# 
�^~�g˓&�t���H�-��kV`�ț�.�$�~e̓��?Q�ix��Q���HWz�7O�YB�I��Th�(U(e��X0���&k�BB�ɱv������]p+�	Wd��{��'�S�t�����O?�Z@�f&�	p�C�I�vl.�C�)Щ }���A�0ܠ#=�Ǔi�h}i�đ+_X� +Ҽt�ؘ �'�*Р��1�4�Bsi��j�Q�'�h�2Ǉ�,w��t�'NRq\Xb�'�NE���[V���'�!gG���	�'AШ`��D�Qj�7�}�a�(O�=E���1/�pؔ#F$e�p*T��y�ɺy�����ӇRmp%ɰ����'7ў�O��=��Tb⠨�n�v��8���yB�*�� rK�����DD��y���"��xBg�?b��C�Q���O��~j��՜����&��z^%p�Ok�<94.�(}�	��O=$����jy��)�g�? ���,�^�8�8�k]r6��s"Oؼ0�b��rr�J��uꤓ�"OV%�eOJ�Vd;��:@�(2�:,OE��X,{ʒe㇀&���5�q���'�<сm��<��R0��­ِ�'m�>@���m�: T�{����@���Ӏ��'N&���N9eʐ����@�����D'��>��݉ *C/8��0�a.��6��$�',b�)��	�l�2(@���l┬˝^X��� �	�W$fyk	����x�W��%�P����'x�A�.�&%����+C�D!)�'r�5�v�ͨ!����. c��D�ɦC��D����å���E��Y���~��OT� k��5��ɒ��osp�9�/�$t�5� �'�'m��*BF�=`�HY�&���-�8YT�b�@m�3z��OԒO)�� � :b��3��=��"OT�Y�E\�dPT�&ͯ�Y��74�P�3G^73����� ��R�M)��TӦ�ow?�*O?�I5}�a�/n��!�7#��	d�B�	fX�\caL�ꐋ���8I���~r�)�3����wœ>)
��U/�G�`��$�>���K
38���ҤG)YG�r�� �1�O���$��vb�2%��%�e�$�"w�!�7�(#`ϕ?ʹ;$�Ŵh�!��i�<۲�T�j�g�7!�D�
Zzu�BG�,ѼP!p(U8!��	�P9��Ƈ�(yc��6e�!�$�&G,�w��<y��x��� 7�!�E��D�r���`M�i����(|�!���$1y,�Z4EJ�T�O�]�!��(U�hz��� #�2Y)AoN1!��M�_L��`�CM1)���!�d��	��UZ��׺5Q��O��J�!�$��B0�1�$&1��B¨��$�!��0�HM�'C͐o����e�/�!�$�)I�d��,��u��M�E瀽!�dQ���2#h �b���	e�R�w�!���h'�L��;!�6!I�%čGI!���<H�݉��W�`�J�k�iȏ3C!�0>ND�8.:U;�i��<U!�B�'�$`+�n[�d��fնp.!�j��Q�g��]�s2�V!}1!�S�(y�e���46�xM��d��%$!�$
65�b {T#��	z����j�:7�!�J/C�B�y�$��3e e!ƮI� E!�$�!$݁C Î^L�X��Iq!��&"� ��C��$����	E�!���	а
��s�BT0b$O�!�$�4J���I2��!&�@ �Q=S�!�\fy�D1�ۊ,���"��!0!�D�Vx1Zp�31(|ܚw-�!�ޑ*�L�@DdC/)���!�ސU�<}��Y�����L%;�!����,���)���رfEk>!�DH�
QDaA֊Q�n,��gB�h7!�dN0k:��d��n<ɘR�^:C�!�D��f�8l���a`�������gja~2��2m*3���[5F1-m�V�h��4^pU���e�A�<���X2	Z����z,�%�r��) t��H_{�)��s�>����ҡ�"5�CϘj�E��dQ:Њ����R!ADo�,�8̆ȓ9�*���l�%1 =ᄊ�_��C��L���=[�Z��o�?��a��S�? @���dхp>^1��,�8V���T"O�+�KK�K4t�h@j��x�P�q"Oʨ�qN�$TwR���KϚr���9�"O�A��C�9N4�J�+��5�v"Opqʠ*ԛ5D�q ����.A�"Ot���,������9��@c�"O��1 �Θ�eȂ�w����G"O4�2&��) zL��h�w��bA"OX�HF\�E�Qza%Ž\y�pZ�"O�f��}׎I��$�	q�$)t"O��`�@N�#�0Jb$�4]���"O����. ��E1�d۶l<�p��"O8��g�!�N��pE�52�di�'�v��!ẻ&2cC�nv���'���ش@�&��0���%-�h�S
�'�r�R����##_�?pH��'V
]��ß�7Į�rI�8,��a1�'�H��L�ULzM6�Kq\��	�'�<QH%Q.�4@�@r��*�'{��Z�,@%B���	�Ӆx��b�'C�P�+\#'^���ݔp�u��'.N�{eS��᧩	 %����'��hw�F'h쬳eh���a�'�|�sFK��	�$A�+g�\��'/�a��`KT�����!�[c� k�'���s���?.mʀ�\�H�n���'�ْV,Ϩ&�� �4��(M%HU�'W4Es��]�|t4q�d�<X@M�'d|=�mM:{�(�J�H�$ժ���'�8��ʗel�������.�!��'�PS'�P���K��9Lt��'��P�ï��dR 0�0���j�ش��'��I���kaZ��Gʀ�\�L)�
�'ތd�K������I�6H�N���'��i�A��Ih)����C���C�'nR���A^S;��wR�G���:
�'����$'��������ܸ	�'?�ՓfB�3M~�b����:j��	�'���JGfU%_��ŻS�:G���
�'�pR�_,@_`��C���l��	�'*������6I|�Y�j�C��I�'��!!΃F��ay�җv�]�'��]��k��%��j oTb*$��'X�YUl*�v��_�ԞB�'�䩂N�u���{%-�'
����'�*���A�q2��T�%��``�'{e"�|��#�Q,
�h�!�'H��ů��lϼ���A�3�n��'�8I��c�MY�!�g$�'7v��H
�'��q���i�}#.�{���y2��F�0�@o����(5��y�.˙1�����P=��Y��A֚�y�L_i<��PǦ�	�D@�uk�yB��\�\D@�̟p�i��#��yB��gAyqB�6"7���7���y�@ͧ��u�`�#-��xD$ʔ�y҂ʂ\:X Fj͐��1r�أ�y���oTp�1�aR�?��a@��ξ�y��-	���lB�X�t��ԥ� �yB#O#���EI)Ur��4f��y�K��
���=H8��a����yG��0�65@d�6H�4 K��!�yD��RB� ޗH���$��y�<0��kA��0ހ���
=�y
� �0s )E�z��T ��G�l�BdK��'�P`�w(
EX�`��Ŗ.	�Ja��u�X)˧�/��[� :�-�<�{�l��?�%�Oa�*D���=��:�� 3��� �'��e&	Ε7e��2D)/����O��	�Fְj"Lu!u�O�A� ���1i`�N~��Nd�tx��M�P�l��C�W�<�$��L�(�.�|�@�]*O'$����Op��@�RA�	�б��ҕ����	3{�F	�d̝S�@�0f�>=����O8s��mJe�Ca0�:�ka���F/�)m�0�!&��-P�:�QP��n������	8	�t� 2�ێs#�y���E7���X��1q��X��I��JԳ@+� iv#[�c7���l�/�=�࢚�n�" h�#>��?� -�@��X���^&�h��Ɋ�� kL�8A�U��i,K�����N�B��L�$'���$e�탲OP:Rq�rH��n Ѱ��9D��6@E�7���[�N!sN�8in
H�s�'�0��'P�T���>4���sA`�#yV�t��V��84 ��Ɗ�Q�l��'����B%�0�Jq
�)����R (ā�p(���
	M��eɈ� �Z,`0*��[\���ϓ�:\���H+i�Ty��È�P�v��'D\Yۅ�i>�X����0H҂$��j�@U�ɂV�b�p/%f<@Њ�GM=~� SGFSM�q�C��	ya�	
.k���؄K}��'�S#d����FJˎL�*����H�{."
Vi�,o�����'��'���yw	��1�C2AΙq��IG@ٓ�p?I��'y�HBa ,������)I��¯���x��N�.n��2�$ڑ-�>IR1�*����V�@�M��b�s��pv��6��$h��H�jAY�0�e��Q���@;N����D��&8
�X6>6��!�$��ڸ��P,^
���� \M
չ0�J .$ ��B�?2��#>�E��%V0e�vFR�`֔e �@r?��i�6���������
	L�(�<a���2m�*�0 �'���k�O�EߎX*q"��&J(��W�p�,8a��(�O��r��D�~]����n��GZ�E�D|���ևN���ဠ�L��"t�ŗ
�je�D�?Y��wW�I�eb ���A�%��s����Y����T�VC�U$I���S`͑�8��ކG܎��!�<��ٱ�OB�]��
����M��󄊝\b���!�Vq�$Zj�,y�qO�(�6�iݍ�U��-zfA8�:*	� "aÙp�t*�`[F��2@� w(�Yg�Φ&�ԕA���{�'G�i&,1-ռ���@9΄q�fܓb̬�3g-�Y�&�ݎO $�I�FM�&�>�6,=9ߎ�Г�I~�)�l��lČ̣���J���`��&�ܴQ �A8a�1�P��U�c��� �
�#��"`D�ɑ2&�ؤypKA9`�!��hVHɰ@�,�󕈎(Q�jH��I!n��r�>��c��*��u�U2X�.��j� [9�L��_Z'T=��I��wP>��%��[�"���Z��3�)Y(N�r���#�~�;�!�	��h���4���� �8LV}R���!۠m��V���A�ŕ&G:�����'<�&h�c�P�%�Z1���2�!$/@�6L5��d;�*.X֎�����OZ AQ
��5V/١���੝�C��K���y����J��򣊣1�r����#����tn<�O��Yc�'A�Q3��!M`r�k�"O1bwk�7_��`�֟9���P"O�`��.�7t���t��iu�E#&"O�=��a�� ��8p�g�$|er���"O"�ZpDߙ+��|�4��\RM�"O~܈�Nۤ 48]���J#co0�3"Or0jD�Z���x`� (:!�W"O$��Dm9e�X�W�b����v"O�4�B���p��yD�;A�|A�0"O��qWbS�*n�9���c��2P"On9[��̡^^��aUG�;|���;d"O�:�V7I3"�aE��5�p1"OB�Ռ�[}l�[�ş�F�0"O���rBGt�����Y�?�0��e"O�x ��5^5�@%����,�H"O��� ��eӶ,��j�1_'��2�"O�5�#�2��\�"�[�$ =𓑟ԩ�R�H�z�е��A��[�Mb��
�eT3��>���)UC��ֈ9 T:E��HA����� ��y��B)@x���.E?W0F�B
��HO*��AT�#�D�[���@K�>�θ���]On�������y�	�%L�xё,�:F�6�0��K�M��i*0�b��>}���iofى4�E�<��y�c��^��4��'�F���,xT�9�͙������O�ԛ�LHjĂ�@ϓC`�e�Ս��t�Е��P�$
f$��I!dN �0�H�9�� T��G�LF���2���#Jμl�"
54�DI6�G3]�9�C��QY8%s4�4ғp��{#,H���?5���H*8ؙ�j�	sHH0R�'D�1gb�	b&:4HtmƬzDd�xe,e�H���Ņ��݈M��}:G"�O��R6��)B�uc��n��P��n;�|�sh��g`4���X;6��3 ��>	��ϖ[�ԩ���<9ԬL'<^f	[O>V�ѳG�l�HBc��"���W�qx��K�c9�1eV�xRv�[҇M�DVh�`�ChyB.	5�E�5K��)Jԛ*T�<���ha(�:J�">)�I�{�B�|*�j��␉��d|�&�՟��j�4��O���gܓ�P2!�
z�hb�݊)X@1����h'��"�JH#��"�z��慌p~�b�'m��z���X��Y[��yir�����1�QՀڂ|�����@�y�S�]!sC�
�!��xqg�+A#DB��&f� �"HN�@?�S��V,dB��R�/���1T��?c`�1�"�g?٤���0��8��/��A� գq.G�<�5 O�`;fmB3�N	&����	B=Z�,!փ�7��@�5�0̯{�'� �Sb��v�X�j�!ȋ?�H�X)8$)Q����M1���
�ڽ����7�C�@7i�@@�[؟�� ң:� �b���8Ӡ@1��-�I�*W���S�J��+�+J��OC��L�]{I���*8as�'�5+�<�x0�F�"8~��g.Z0%'D��S�W Rh� �۴0��>�zF�-q�ѫ/�8��L�7�\؇�_�L1��G]�(��=B� ڙI�|o�Dꘋ�E�0EJ�{�{�\�Th];#�(���J���=y'd\ _�p�e�OXd�J�����d��^3���"Ob�(e�I�wO�Y��"ɡ�dCt晰���h��I22��<Be��'���:H��"OƘ(�ȅ�Q�]0���B/&I�'�0�Vx%�|������%ZȪ�e�פJ0:�n,D�xK��J3e�>i����q�څ��y�0C���O�|�^�(��l6&��`��Ǟ(�yD�7����܅؀mr�Ȓ�yr��(�
���δ��i򤟉�y�^Ux�Y�ԢN�����@�E��y��M�������~8�J�'�3�y�����w��P8�7ț(�y2)Гl�q��7�����c2�y"�D9HD�Ҷj��0��t�S��y�!S�<�H E�Bv�*̂#�y�o�i䖱�����4�*��R��y��\:2�0P�@!�SC�͈�ybMO?��4+�A'X�{�i��y�
Z��>��K�4(90q��e�y�'\��y1�/��'���҃�:�y��ή�f�ӵ���V�@�Ŗ��yH�D�L����F��Ω�AgȌ�y ��"��Xc 
_P푃�N��y��hR�� ��4$ b���yr�X�Q2�
��J��l߇�y�hC$�+�m��K��0��yBHTsf ���Eب�d���y�3I���g	Y�Ƞ�Z�U��y����u�:� �kĦ	$��(�m��y2�� tڡpqʆ���T��yB��~��[�,J�)=�=X� ƻ�yr�
O+`}S�A��]�p4��G)�yBoK�a��r&n
�W:^�f%�yb��@��(��լO�ʠ"���yrL��Qk�EǪS�z�y���y��*+��z$MăkN��e���y�\ ���+��Q4�
�1���y���"p�:�����}%���F�Ȱ�y���E�tU�$N4iqĂ�b�1�y
� "Ax֦"K�85���W	z�T��"Ol�Q�C�P�hB��6$2�S"O�)�f�̕������țzN�T"O��ĮN:NЭʢnی��[�"O���	�7MH��1*�6��d�"O��)��ޗMIRH�	
$>�Z�R"O���F�t�ĨvG��"2���"O���/E��l�G g�L��"OV�x3���Q��u'�Lc8|��"OD�H2ə0d��H7�PA�Lx�'�8�k�g MJXx@@����	
�'�hqP�Nǅ@	��"l_��4��	�'D�!2�"���"X3$3
���'1�5k�o�V�ܸ��L֬Kv4)�'��]4@��2@Lp�'�(:����'a�H[d� ��Lȃ�;�
L��'����'Z/�!2K���PK�'RX��/�3_�U����#��9�	�'�����F҅&��i�C�+g�Ւ�'N�<
!��Ѐ�&�� ����'Y��!󨖥N/Pi�&��^����'��xU�Vy�h�F�ra����y®�>���҆�+e���b�gϗ�y��߹��0��%���`���2�ybI_�
,��)@�DU�fx���*�y¨��'�&��p�@O�|��ab��y� �(� �D̳1Qv]��IU�y��.?|�]s����6���9EO��y�%ާYe\Y��O�{��� �f���y� 5��@�㨃q2�@���)�y"�8p.X2%�i�z��5�#�y�A��2� �pHP���֫��y� �Wc��R�p����ŷ�yr`�_��T;�/�i٨l��FJ�Py��J
qצI��*u�'"OV�<�Ӯ�:82�
�,߄"��4va�S�<��Cר�J����)+�Z�pďDK�<AƮ��|�"�"�[�!�� �U/�D�<�gŉ>!X|��A��*jw�A�#o@�<!`���� jI�dJ0 Ðl[�<)d&kI6�f�Yz�gc�_�<qE���/�<M[���D;y��&�W�<�#�	;^�a��)�0e� ��1�P�<��ɏD��yWeZ�:�IT�H�<YU-Y�4��a랭@��4����G�<)'�+l1��)�FA�v��5a�LC�<)"��e!	[U�?x��-@�C�<�tJ<�l9�F�C�MdB��D+t�<�F ����$J�@��<�3Kt�<�@�:_��@��-k|�I�e�Mz�<��Ϟ8�FIB� [�I�]m�<G*E�)���0�ιG�8b��@�<� � '�` .�#Y�켘�T�<���_�P���UHL��h�i�<��L�^4������� MQb�h�<�@
�W�X�;�cT=C�|a��Jh�<��JǯO�����h�60+�yu��g�<ْJT��Re�vײz�>tГ��c�<�q@#d��iC!,{#ܸmPwj!�DX�:�{�R-�^X��ݥRv!�N�Vm*=kq� �v�b}!�4l!���vV�xS1eX9�$z�ǒ@[!��ȅ(��#c"M�@�,YӐ��:D!�$X~�B�0wJ��H��%c�60#!�� ���s�@�f�([Q8��"O�x1�dE<J���Æ�?W�8y��"O��RQ*&cԹKR-P#<��XK�"O��r�P�}pf�����4_��e�T"O,K*�x�� f�M� �є"Ov��#u{lQs&��8���(w��Q��U���h^���)2y�]��NE/L�!���8\?��#�&*j�+wJ�z�I7�Dy��y�)�'��i���>8yѵЎV��ȓ[���u#=�����	�rL�OZi�Ý���ÓJ�z�Ʌk�F\n$Y�`D�;w� ��I$�:����m�-����54��(��a�#� ��O�0('T�$�h�@��"r��d �CLQq �ΪdEZ��ю;�S�i
���&��,m�q��+mt�C��)w3�d{@ԇ �J��2A
3���ZgcH�VJUh)U�+&6M�_��������@��O����m�h�!�$���ɤ��= <�a`��7%ɒ�H��O��+��p#Ll{��'1��跈�	�<�g�����2�N��9� A5y�@��^�C]$�`�?a)��*W���Vz.�
�2�x(�i�\���5h�8*�P�v$A��l�Â�Nnb�����@:�Y!���uR��*:�1"ŏ�7N�͊G'N�3*���c8�O�p���K�L
� wkJC�Mh��M����Ks���9��&x�x��'����" �w>����e�;
����r����z(9�'S��z���
3�<�j�
}�>qsS�X�'��pа#	""�L��g75S��B"�9�(
�*D
|�:y[�'�e9g	�-D A�L�s�T��IԊC⥝7�C�E� �����2/f�(Z��T.�.<�@�^E* �2���tDŒa�á��#>�`m� ]f�	v�*=)��A~��J�P�߄iU
�BP��1p�^�)Q�m?�R`D�fܙ���	���k��c�Rd
v�\({�a~RG@/j|�ѣ�M8I#X|�Cۚ8q����8p̤Ô��-0�����-bp���;O)Vh�Zwj��]�a�2���@4<+:��
�	��B�I�v�!!��W��&G�
Ya<
�U�`� �P9ot��������)1��������	_k
�ɤ[Ȋ�������JA�,ۄ��/ќq�%,�.�Dcu�S*Nv0���M*�j�"��T3S�.��䆑OԴ���-�J#>�(';	*`PW��<"��!1 �L�'0�ZIO�̥8ROC	%j\<(�#�!"�|Mqt'�#�@9�%�h�*Q1%�Dp�(��'�����,�;b�h��/��iBD͹���>�s���$�f��f䔝����q��:c�b�0�o�Z��#��@�!�_�� ��FOƊ !�^�Er�8c��G4�¥��Nͩn��Ht�M�5�pa�]�ބڶP>����+snp�kZ���(�3�����E�^��IQUC(�O���q��G\l�	FA�6z��2$��6m��)�d�b�i�g�I�A�d��g�cu��-4y�L���D}2Y:WL����ǟ�� .Jf��N�8nkXaI��ӄg����C�&�!�dV?.1�te�"�"�Ǐ�2P�!�ě/V��m9 �ǳ�H�۴���!�[��DY���<�N��'�4!�D_K�f� ���i�Ak&���!!�D�t���	R�\j�l�G�ԁg-!�dР
��d���1QH�
���3!�$�8G�R,�t�Ɠ�V�9G�M�;!�d��kA��XE��ce��2t	!�d�>n$��MM�sH�s�
:"�!�$����C��o��X����Q�!�$�6��Ȉ7C��,�Z�iC�O�y	!��:)Ӕ�f�����)�!�,!�V�5� 'X�9<�h��J&!�䙼%�
�h5J؍9F��7��<�!��J�t���!���%�����-&!�ě�$���Z�` ��QfG�.a�!��4o�iߴk����e���!��i����gM�#vE�EW�m#���kE䚖�'�y�CNJ;D�B����ˇ,�\�X	�,�T�pQK�86pĻ�@O�l	j����+a�X�	�'-�9�1��N	�� Vk̍U�i ��d�	ʒȠ� �'��O��6*�&��`�ef�q�Q��� �HR�%/e���C�%D���iȸܠl��d| Q�O?7M�T�e�C/Իc��೦^4�!�䝫��9�㫛/nZEQ�O �����]ڈHjK �y�dX�lX��MC��Ƽy��J���>i��	�^�$��M��~( |xBfF�QBje�g�um�B�I1(&n�H�{#N<y��ϋvߢ"=�FE���$:t�/��ED\�ۑ	-��2���2��C�	�!N���Gb�+/��p���v~6�	7�\�(eE��)�'!L�I�R�d��2�O
p��5@�<"C�	�ˢ̹�,��W����ea�;#[|�d����$L�	i��9���r�
���"�;�УK����y龈��Ix��	��)�y�d�@�8� �"�Т�*y�'����tk�-@���OQ>-+�VR��!��X�)U�2�e�F�c
 ʧW\���'W���SC�(:�,�Q�>��g��T~�iL~�=��'�6��ŚSgB7+Qd����g��t��gՂ����Ѽc@��H%`V*_>���ɮ�a��� y�a��ˎ.���1�C�O|�Ё!��A�5�4'vڐ<�)B�gR�x����	��c�X�$k!�$
�ԊL��Ϣ��M�a��u�� �ȵyB�0��N�7A�[����e��B��X�gg[�'�J�hI2D����&��^ԠA��Fy���yc��R:�,��kڵw� ˓��2�*��{�'&��`dٹ����u��1��ۓ]�b�3�f¡}�>X���eN&�!�\
<���Ӵsx��`�$�I؟xP6
�9J��I�%�C�V+�����/�I�!;d͉#�2�,�*v��1��Oȶ���)U�c��j�8B�'�vm2BCّ0�q�b���L��r*֥$8�q ��.�L9cٴsW�>��"ݘ�%B!5�:���oK�F�5��C��ç�D�h�$;q�+W,Ilx��Hҍ�f%�{RhO+,��@����nረ�/�.��=���P���%��O�U��!_$ѭq���	lV�"O���0n�P�
�Ǖ�	y�m�U�D�x�d�;��B8�h�����i�)��#4�ԳJ`ʄ9"OP��r��>lH�ʙ�	a�<qwD�.��Ӗ|b�����2�vL�FF#%�Y�)D�l��"U6z�渹!HJ0C��Y��g�`�)���|B�Z�b��!��ש*�B\�0"\��y"@o��t��
!�
x�`���yrj�l�dr�O8�BQ���ߛ�y���2���)%Mܟ�bIA���1�y����;��9�ĤJ��PTEK��y2�D."e�A�x  �@"����y���ERD�"s,�x��d"R�9�y�K�E��X��Áx�,%��*�%�y��ԃ+`JH��F�(K��O7�y�I!y�|C��+n��4aΚ�y��"~��C� #$����ĕ#�yB�M=(#^�yũW�jm*Ջ��y�[%yQ�C4�L>'J�R�N)�y�fR�8=��3��;*� {�D���y��C&�lY`C(%4�5��L)�y�̞.8I*�H�&���c�K��y�#� �X|�Tf�L��pV�И�yU 1N�TS��7j���.t�D�
�'F¡�\���6��01u�X
�'��)��㑪6�5C1�)=H>���'�t��Ae-t��P�gnB�0t(���'{4��AEӞ*Fp�	���(.缝 �'P�U�Q�²v�n1B-S)�U;�'-�x�7U(02�vLA "�}��'[�0RE��*(�#v���^̊�'"���G�އ=�^0Xfg��V�I�'�p�Z�!�9U� Ui$k:�
�'
�����.�HE���T4��'H��X2�N�f�a�/ڲ\��2��� ��zc#Zy���SaJ^��H�q��'+�Q�irE�0��FJ5��H�z�(�7}�JN�w� ��A�O:f(R��^}נ���7;�XI;*O�Y��J�P��tj5���Q?�W�޳*e".��R�ʠ)�l�O�9�BF��r�� �LBɆ��)�
P��%�U�VLa�dZLI��#C
�����
)m�)�6���If�A>x�A��ж#/T�`�kd��'H�<YU�OZ8��d'�C����F��e�ذ�S:Jw�42΀�M���B�a�4n��5��{�H�X+�\`%��
�4mPCi�1��Հ.*B��)�kj0 � A�$���*_�U���V�@�$#�+|�T1��SaoN�Z��4V��<�!�UCj�i���qc�+:��4��*e8����Fb���m^�gN�	 qzUa4&��q��O���L�l	�@M�8����F�' �@�� ��T�}��S�O[�$�ތml*��V�=Șd+f
ĖC����&`�I-a��a�$H{ؠI5���<��Y��K���H&�T�`�׈oa���E��U`�O�%y�Q���B���ɲHJ�T�T-G��S��,cdd2V�V�}��|��"��oL�]�"f�c�l�w鎇L,�S�OK��ic]Ȗ�p�� 7.ERq���]f1��ٕL�H}��]�'E�u!*�j���c�;�  ���C��`p�,�~ I�-Ʀҧ'� �0|B�-��:O�ٓ���b]��;��П���$ڽ)�Z!���=S�� ��S�n}�@���w8� -�c�b@���я)��s�K�q��ulL>ɫே.]$�,��)�64��m�7��<
�x��U"�X��lK㋚�rH��	�F��rt@S�Sx$z5M��z�4`��[�G61�7�"W�ֽ����$՟�O��P+��cT��Xh�:�%�O5"nR%:a�P2�>��)1ʧ2��2�J�51������-.���!�'��]�'�n��r-M������O
��Շ"M�p2q�H�D�zU	B"OT��̏ If쨘�i�/9���p"O(YI��Y6yMtj�U�!�zQ!�"O�!wK��~�����O�o5���"Oܰ�(� ,����&0���"O��"��[��Y"CJ�RzE""O�`K���:��P!]�cd.8{0"O���� D20a��� -:Vڄ	D"O*x˳o܄)ݮ��aZ�"n9("Oځ�mp�1Xe��1��E	u�<���]s�-�#�fG���r�<i j_)'�&1J��W�`��@���]l�<iT��Ka���cP(T�<J6�]k�<I7n��~�
	�K<H����ng�<y0�9�*	���4tzݚ5��e�<�c/x�x�QpH�v���g�e�<��B�C��!�-�%G�\2��Mf�<�	P�h8�!����C�@����b�<�AɃVPt�p���,P�nG�<�υ��c� 5ݐ�I�Áj�<�K͋~f�� �ea�}yrJEf�<i�j̦K6�Y���lD�m�dJ�f�<�GoG=��(qdG;
�����\�<��`ǧr>晐F��qz\c�iL\�<���2{�*s�͛��tY7b�[�<i�aثs4��@M��y���4�T�<aWFc����jى(>���dWQ�<i�(�4a(�h�C��=����'K�<m�!^��s�@ʾxk��4���y���� C�!��5�� E�*� B��3f�X]��"Ub�LKr�:u�B䉩l��p)��U��ᅍ�ѺB䉝�*�h�b��4M�]���@�P�B䉏A��'M�&�N�+�-B�6s2C�	4g� ,�⣉5(e҅q�%A�%f$C��)3�|t(h�LՀ�[��2W�,B�	�H�x�{��*]�(�(g$ѩ3X�B�	�mRV��b��,X���gS�B�(6��LN�>�"pZ�&�+>�~B�I��r���nȁ^�բc��4bB�)� �MB�%w���L���d��"O(���`�/�|(ړ+�t�4��"O���C	V�p�0��A�Ə qN,�"O�3	�a5�8q��5Y��b"OV\Y!#[;9���Uś�vGvl0"O����;]�IR�M��r"��Ȅ"O�A���^{��sLI(�Ru8�"O���śU�~9Ise���N��p"O��#��.G�$-�oW� z��@"O�����_:h��*b�BX�B{"Oy�(D�R4H���#G�=�"O�hRV�ð~E��X�AD���"O�<6@�:l�� "�@BY��"OH`k�i��B
��1ԻC/��Kg"Of����� ="��yC3Y* ���"O@�0�>'&}���7E���U"O]R��C2+6`���.�|EY"O��%O+z�N�p��(Æ��S"O��2�JU������TF�[#"O�P��$�*~�8����z�g"O�|���Q�6��#���r��+�"On��v������AT�b�4YQ`"O�d�R@�9��`��b>t�`"O&��F��#|���h�.�UMJ���"O�H��� +G�<0��	;1I���"O��)S��.Znl�ĺI���:�?D���Ȗ�3&�Dh�BFj�9��#D�x0C%>�꼚�"�l�I�D�"D�(�����ZԘ�P�TG�0إ.>D��B����j1�B-N%;^��S->D��jB��/��h��Q�p
�ȇ�:D��F�[q���P�8ơ�v*OI�R)o޽Y�e��P "O6�),��\@���P��-k�"O8����<1����7@H˲�R�"O���AA�f�� 5ŀ�z (��"O
���+t1��C��Ve�pA&"Oh���Q��8�,3+����"O*<@��S }Ak�G)V�+�"O�$P���iZd��� KW���"O��A��� 
��` ����r'"O�ݫ��� PJb6���!����`"O�tv�&�Y�6- �m�"O�\d��A+q������ 05"O>u3���F��<;�A���2Ѫe"OfU����$r]F��j+l��-z�"O��aBL�'��Px�	�d�~tSb"O D�$"ն3I�q E��;>h&|�"OŉFAE�>�������w�bI��"O�q��eܳUJ֙QaHG"VHt��"Ob'd��-`�7�����J"O�HA�^<`hH� ŋsAڬ�"O��1ǩݽv/hP+�AI5t<^�XQ"Oܴ(�W3qV��q7gQZ�1�"OT�k�*Ң,�TQi���)E�	�G"O�]Ң,���^A�YH�Z�D�h�!�X� -�%M"�R�\�x!��U%x2ҔI�j�62@#��Ɓ1!�$];�%�A��d+�!@�X�v�!�$���%�� W�	��`���D�!�d�'4���Hv P�sܥJ��,m7!�Dښn���6C>�ȑja�6E�!��̈r�n�qc�>^�E�زP�!򄆊L;���+C�/W�q�%N�4�!�� � 
'
�_�i� eP�<�Je�"O2� JSO(�Ly�-�r�!�6"O�HcA�J�"����':�A�"O�)���!(,�����X����"Ol���$L	vd��hW�M��uI"O�y �ěrF����
6[���d"O2�BR(M0��Z�)�S�Z�C7"OD �r��[�����ȧ"�z�sb"O�l�Ǩ��c���I�l X��"O���DS
 �0q���QXVi:�"OD-1��"p�Jy�i�5V�IҒ"O�V�?T��0@(׮ut���D"O��Z����48tX#�fOZr`82"O���p��0�y���	U:\�d"O�=+��Q�b���JO�ڶ"O���E�Ek���"w���\�<HU"O 	ig��#U@���T���jU2�ʖ"O�Y�	I�Y&�h��G[�#^�Q)"O����(\P���b�$,ڱa�"Oll{��b���C:7j�"O���e�ͼ{����'=�p y"O�t`�EA:Nh��@Ʈ �J)��"O, ���
�'><ȓ�T$E���f"O� u��I��e�;Q/h��"O&�� ��ܜ����$�}2�"O¥X���z?�̢j͞
�B�"O(4#q�8d���	��P` �1"O��Oυ?Eм"g�s�:���"O~qs&��n"���&�{��ds�"O�ubU{ìys���:!����"Or��#M�J�(ʦ�إt��f"O�0�mN�nQt5p�l�K�֡�"Ou�u�Ι3�*��RIQm����Q"O�mI!�L�Q�䉃w��1��S"O��CFA�"P�QW��<Ӣ%#�"O��j�j��1*́D����P�C�"O�8;�h��z���f�І
{��7"O(X��g
:�,���.��y[8�;�"O<��B��~�h���,��3�N0��"Oh��[&rR.�Q�ʏ�N�x���"O�Ё�L�0<���G�M��	e"O�����9#@�ˤ��E����P"O�����%�����D�@��T��"O~T)r��f	X��C�=yn�8��"OBU`�C�Hz�� !>Z�I��"O48�7���|}�" �O�Oj,���"Oq�3A6
�rM�eO�3A�Ę"OB�qŭݯ#�H��]����sd"O��"���#B�� ���� ~�*0 "O��s�Αq �Uqc�_�Q�;0"O�� 0g�1]�@uiBl�+��9�"OM92g�:���`�d[�E���"O  8��"1����P)V4l2w"O������� ����3.��A"O��0jߺ=�ġ���+N0p��v"ONiq��J���P'�.b0Zٙ�"O�Q�pEQe芰�v�Y)aw ���"O�
b�]E�Lӄ�ϳF]"���"Oʌ�p"��3(��{E�:f["O|$@gk�SH��P���#U	ʴ�yҌ�k�ء�1�T4`��s����ybO��Zh����W$,�|y�I��y��@�VB����6�!�d��ye�2ލK�Ô��4#0&�8�y
� ��*�-�WS�4���>�P��e"O�$�"�1����D�f���"�"O�Y�R.D8n��ɣa�7e��u�"OR�*�	�
��e��3�t�"O���c�G�V��X��/l���"O��s�o��zĸ��;<o�Q�"O�Q�V��'�T�0�	i�iD"OJ�$��]?��� �4M[ڔ��"O�-hP�@�%L���-Ld�C�"O`�
�E�N���c�]�M/~� �"O��s��1F��f^�'���w"O��8���IƜm���4H�z�"O�p;��|.8|����
��e"O6���M�<��{�X�;�dE(�"O~�kE�?�Jt��`҄:�Q�"O���WcD���3�A.+V�2"O�	lʵ� BG�/: ��"O�4�7oC�n~��gG�[2�Rc"O�eӄ�H�@UX$h�G��5R�-�"O��K�cU 52�!��:u�"O��#�
�8<���Q�_�P�ٵ"O��9�g�R@��"�[��F��P"Op`��*������
kD ��"Oh���]	-PH�%@�:X 2��"Ob���`�2�����D�@%��"OP�C E�HY�j"��s�	��"O.D��N��L,�볇�%����"Of�bv�R�O���qD���b~�`�"OT����6�j�2ƇQ�"%��"Oꤳ ��g��嬓�^�^E�"O<��f   �s�VU�߁s����S)D�@@�>@���0�ǭx�hȳ�D$D�p�ոV~��A�E%3R,��/D��hd���\�j}2����8{L���/D�(����Q�!H�M,@p���/D�82L���Хr%C�3C(�8C�/D�dbe��An��Hc��
K����c9D�(���0nb8�S�H�P�}[C$D��)��������#qs��)B�>D�0XU��!4�P80�)Z�bd\aG�=D�Ă���
d:\�AFX�y1nU�W�'D��ȇ����Kq�Kzd$� ��(D�P ��/	�h�情+I)�!��J*D��H�;rQnQs�G�#����,D��JCOQ =�QH���`�$B1�-D�dC'�C���ʰ)��D�0�`-D�<��&�"Z<���.�\��5!)D��1�F>���`�@F�,C*��&�&D�ۦ��!S^>D�$D��� s�6D�h"�?n�X;ŃQ�*��I�Q�5D��*A�%��-K��L�aŠ2D�p��lH�z���.�%eOb���-D�L�
+[E(�Abf,bM8�b$,!D��Y��8Qjx��O���4�� %D�lR���x�C��V#)�
���H$D�X�˖p��7��G-Ƽ�q�'D���H���&�C�%���ꦫ$D�|�,�&3�p��uh�1;��`h=D�Ӈ�]W�钂̅Y�^D�Pa.D�� -E�G��3r�&�,��AJ2D�h�C�qܐ����ֈP @��.D���%kJ>0�S�@6���r`�:D��@��υJ�f���C�%���� ,D��R'�E�
K���㛟u~�(�J'D���6��2^�1ׄ�r�@� ��0D���񆅔4���Pl�?��@8�E0D���堎pRH�0��Sj?��V�-D���J�3�|W�V$:A�l[�h+D�� ��aFz�4-@�
V�[B���"O���J2O�fX��,ՈV�<y��"O`()"aЛ �~@!�+�%�
q��"O��b�?JT{R�ʎ��@�"O�0�2�J�6��(��m��r�p"O̐F���\�� �+~���1W"O��GF��TN��DK�2���f"O M"vM�7�b-�4��m�Ƞb"OpС5'ӟ!`��
�	�$
ג�"Ob(��kH�0�Ե����?���;"O�E���>�^}Q��DQ�tE"OB��@@%:b�8�%�G���A�"O�)j6��N"]��o_�o����"O�i�f(��U]�
2N�1%����"Oj�"��	�������\|ڤ"O�	!�:<���
�On0"O� ׾^ޔ��Wn���	�"O� �c�z�Dhc��?# �Q�"Op���y/>�bk�| ����"ODe��C�v/��!L[���`�d"O�hc�i��۱����"On�񧫃9 ER��e����"O���vM{IZ�jת��}-R��#"O�i[F�-@��x�R �H$慺�"O�����&U��0���8�ā"O�!x�-_�b���0J�}��p
�"O̀��	T�nɡBKV�~oܕ�`"On샢&V��`\+!�Y<a�0��"O`�& vG�(���9DM�u{�"O~1�sd�"mx�Z&�e	)嘞�y�̽Lq�����@1�d�#b���yRȈn[|�Q�@	/���ٔ���y�� O���v��*��a�
�P�<�&ܶEoLl���
;�H�u�K�<IǍ�W�ʉuG��7}�<;F��n�<�צ��Eq��.��|>Y�&�
h�<���΃�֍kê�jƆ��e�`�<YE�s2 �g݁W�ʱ3�#�`�<A��(X&2�J	�5��H{���Z�<����kvX�΁I��ӑ�	X�<9o�,���*Wج!�s��V�<)%��CPڱJ�g��u�	�P�GV�<9�F�P�aWd*)���PcP�<aGc��1�\:0�	-��A:s&�H�<�d�b�|�9VO҉?-�X�b��E�<�@�;n6vX ��˂wy�];�iGD�<��־H�.Re�x�E{4�d�<��-C jJ�x���߶"�t�qCTa�<)χk팤jף���n�MC�ɇE��Q�A��|�d�ѷ`�q��C� 3�.y�"�P�`����K6��B�	�D���#q)l�)�.4*�RB䉟D@�������D� �`G&�3.>B�IVm�T:'���c�DZp]=!�&B�ɰ2��(�fGȶ0|\ٰ`��%�B�"��`I���n�2eH��8�zB�	,0Z@�P�H{_�A��!q�DB�I�%����%��|�urQթ�$B�I���dZAف_��!�!œ*wB�I/�F�'E̡a��B��P�PB�C�	>C>6�Aĉ (�zxs��V&B�Ik�l�#��̓K�)��!=�B�aŖ��A�� >�A�!r:VB�=Z,�X� D�/��ɦ F�Y"pB�)� (a{���[��Z`���.b$�1"O�(����<>�a!�M�^-*Q�"Oڐ���ĨgqL�0!���-���"O�-��U�s�|�0i�;'�5YV"O��K@�Y-s
HYU�ю
*�k�"O�����PrK� h 0Ě�"O�aĄ�6���5�M*l����"O8p��O1���g���.n�H��"Oju���]1/d�jR��"2Pb�� "O!�a
���P8k&,��G9X$��"O4�q�/�F�vz�֫�t�"OF�J�����,�FjϏ_n>9��"O���#@Z�	���Mk�a9�"O�%"�	�  �P   �	  �  =  �  &  ?.  �4  �:  A  _G  �N  VU  �[  �a  !h  cn  �t  �z  ā   `� u�	����Zv)C�'ll\�0Kz+⟈mڃ	g��,Q}~�D�\Kv����0MX)���޺l(nIe�ڐi��q���)�(Yj�J�����/�T\���z�8ł��jHp�RíQ i��@�4������'��k�)/lm��� [ᦥ�׿��� ����D�`�	����N
�u���
J�<����E a�^)��V%�U[&L# ���޴zc����?����?y��2w����IJ%4ȘA���݊��? �ir`���W�,�am���SޟΓh:JR" �)�D���k�����Z�͕'gr�E1m���蜵����	R",�:X�X��v�X���r�!"D��I L�1{�hBg���h���>ɛ'�O�hRB�N#��Z����]�0�D|ك��.&����ǟ\��ӟ���ܟ\��� �Od�Ο>{���N\U
�I���;���O����O>�>�
hӬLn�0�M[��Ld%2���u��@�(ES��̣���J��ȟ谈��@�@�.<���S����P	X�A$K��*
6l8u�z�p	n�M��'a���K�3{�!P���m<��׀�8m�x�ww��l���ĭ=�n �S� �x�Y��?f�H�i�40x��`�D��`���5u�-f�͂e(�0;�\cqX�tj�2��ix7�Y�QZS,Ra�jy�n�"0̆���`��߬eV�������\qJTA�Ƒ,#K��fB��Kb��Qm��M�P��$X@��э�n�H�q@ɒ� 2'N�ҰtBR����a�d��ia(	'f�ԩ��J�0$r���'�r���kYIc��5̝�y`,dI`��/N=lY�4ki�f�o��M#���e���	����S��=�?�ϕ�yf�T�ڕuO���K�yb��9RB��v���;���B�F��y"C&,\2M3")Y,o�̡r�ó�y�a��}Ѱɹa��a����x�|��ȓEBF@#�+�3B�d!0OY%hcb��s���ss�(j�$�w#Z��E{�)CҨ���镬��E�3E[Ry�+"O�K�Ѱm��P(���Ox8���"O���¥O�?v�u����J�Z�V"O�MA�c��Vv���@��B�a"O�u'�ʋ-���he��}fT��"O��A�D��)�\ c�l�;K�5�'���b���S)�p��m�,��gU�l��݇�h��p3�a	�ŎY�擸g��e��s|�c�eW�U��P`�\5jP���ȓY �hW
�8��`�Ï+�"Q��F����p� {}\�X���	7^��ȓY\P̱��sP�Ur�%�e��'�2���Q4fEa����u|@J�c�/JO���ȓs�-�rh�=y�P�� 
�-��ȓp����+��Aޘ���:X�4�ȓU��1�-o�hi��0)�Ʌȓ�\)��٪q�A6��������ɻ�>U	�4�?y�c�D���N�r^t����}o��A���?�E�Z��?����doöi�p��mz��I�B��R7�Ȇ
������=<�R��$^�8(��aF�Έ>��	Q�sb��	<B��VNݡ
�����s*�Hvӌn����I׃]�0��u%�*&�8q[4I_pyR�'��OQ>��0.M,+�a��N9����A�7�O�t�Ɉ�Z%BD��("�t:���o�f�$�<��]�?����'�����)�cCB/fE�d@�^'b�	d�\����ӷ~b�3�,Ώ\M>����>�\�Isj8�)§m�ɨ��>�����VEh��'|�!���?qN~b��'� �Q��1L*T8�'G4���?i������� :ysi[�\�Gb�,ڧEyV,fO,k�ب�ǘ?V�(�z�4�?�-Ol�
3���#>i�bϓSG,�IE.��p��#��#�%Duy�[�V�Az���y2�>�~y����:�d�w�ӥt���@]��� c�0|�c>c�h�ႆl&�b��@*58�#u(�O��Uhp4�IF������$X�.Z�h+�7��{���3�m���y�+�mu�qGo�!hmT��#C�4��$�B����'G�I-$�	�c�d@�a�GI�e�P����~�d���=��0�4*L�!3%iɛ4�J�x�$7�,�Ud&u1,�`���v�<�I	p�(C��'w1$�����`{��qe$�{�tUSg�O\C��!
�pHV2s�0Ё��V��B�ɃG�1�f�A#du�}�r�x*��O\�og�	J�,���G��m�.Y$d0�M�ph>O��y�/]���J�� �������s��Ck�5��@r��'4!�'��c��8�O�,��]�-TL���cV�c��1���'��m���?����?y����LB4E@���p�SKǛ���O.⟢|:��q���0��{�Y�C�H@�����c�8m��Ɲ\�.h�d�F�RA�h��Vy"�!QB7�3�i�����r>ŚqAE7%nl����(A�<A�*�O���T�V"�Q;W��J�4\�"|r�Ϟ�n�9���$��� ���Q~b�A>c=a���\�?U ���.M�܋ӌQB`��N'?�7�Yß���|�a̧T�9a��ö/S`A�Ak�v9'�8��A���
&k�74 M5�ߗDC��8�&+�v��>)h���K�����ʥA�Ɲ�G��O�B#`:�i>�<)fLB5DI���D�#�dQ �R�<��F��Iғ���G�ݺ�J	g�<��+ō>A�����*�ژc�k�<��J
_�^t��E
6���Xw��g�<1egQ�	&�I��EP�1�k5�Xc�<��C�T�ԭ(��+���±G`yBM�p>y��Q߀� @�ڀ!ڔI2�H�d�<'\�tD<��T�#?mN���V�<������̀��� 4-k�C�Q�<��J�m)��rEFN�k1�ө�J�<VG.�����!a���ҩ�Ix�(!%F���M��]�zD�C�?	ޢ�i�#D���\�H�H�!�	Im���A`��yB���]�� �.?���tBV�yB�4��� �
׋9ؔ�����y2��
K04xPɆ�h�ej��y����J�P��D	�:�I�.ҝ�hOX\����L�&��!�#]��Q$��DCtC��(g3�#�e�q�����j�(�B�I�{�L�� @I_"�΁f��C䉆KX�$B���?�:���X�G�C�ɍ?H�L ��$.:�᎖�w�ZB�I�c��!��'ĺ#���6��QF���G��"~�'#+%�L�ɤFH2�.���g3�y��0p4�4I��!,�X�AE���yb�T�\�r5�a������u�^��y�'��s��	�e̝�(�V����I��y��Y�2��Z�[!Td,�P���y����<�&��"�����`�O���UQ��|��IHm\�cFSC�>�!���<�y��F�Nr�8���8=>l��H$�yBhU�.0���T>�>���B�3�y�j�>v<�p2`��Mhb�b$DJ1�yBg�).��h��F��P�	%�A���>��m�o?y��K2nc�YQ��\*�co�u�<qsk��\�D3���tFNMBc��j�<)fM6Gd�Qyt-8�h\��%�b�<��Īwr��Ի��l�E�S�<�Q�V=/��D�@�߸L@v ���Q�<Y���E:�4��̶J�r,I�!P�'�h�X�����#͆@�&޵<h���!F�]�!�E�Z+\L�%2E�;�Jڋ"�!�$�6
��(3p⋓�V���jӲ9!�䕔̬�HFo^�{���U�B�;!�$��MB �Q�*Ed���[Y�%!��_�����k�2<\!I�e��}g熏�O?9ʵ�Ϙ3^�Q㟌^�vI!�X�<!�mN�p�P��>"O� �KY�<	�-ɥw�ސJ���8j���ehY�<��&���u��e��u��PƩ�T�<$J��6�ⵉ�������T�<9��� \�\��A��3�훴+�Ry��л�p>Q�l�;Z$�d�u��H�V'�K�<� . �Ť��-�8 �D��z�N` �"OB��e3M�8�����l��T"O�Er�އw!�����<i���"O�E�FF��r;<����
�h4�6�'���3�'l0�{�)ڶE���Kݬ^�� �'Kp�����;�zP���@��x�'C4�v���@�����#d�'|��FK24
J1ꔈ�+�P���'�d��v����XT�d(U�lP�'adYr&�V�}p�ZdE҂ޠ����$��&iQ?�JG �Qk�)bI�>B.�
�/D�,����?]������l_�-�r�(D��H���c,e�FKD(/FT�C(D������#�(�(��R&-[ �$D�@)�'Y+'�6p����AE���/6D�����;\�-�'*ߞu�����O�@4�)�'<��}	 6R�\����.�(D�'�:���e�)R��h4���-�8A������۬|�8|²-R�JY�������V�q���DL9{�bB���Mն	6p�Y-<���ȓ=;f1{�@J�sR��)�D�[���'�0�:�w� �Nݕ
�T���O�otz�ȓ��"�΂fK�Iw��%#mRĆ�$K�a�n�̰�mL�/���ȓ6�!x����i[rFռvN���ȓ5j���ȟ��<�q
S�C� ���q�h���l�5r�ҋs2T|+�(Y�v>xB�I�B�Hh0�@(a�0h�nû|!nB�ɫ?-�Л� �I�� C�ԛ� B�	�2s����e$P�Ʊ��+Q!
��B�I{Q,�����`3kN�PC�+D�<*u'��a/vqx�I��\Z�l���5ړ)p� F�t �c�< �/TL�؍�2l �yrΜ�

`P��[.T��؁�=�y�GX!��T�#A�EY�xZ���yb���&�N�s!_=�� �*ٖ�y�K�x���@�Aް;�,�q��y�[�j�$�2���r ��&�?�wT�����)�f]+&�l,j@�+Bp�M(D��QV��(1����$�\����;D��x���*h�p܉2�x�>�¡c7D�@�F�+���D23*4�*D���,�H6\Xq�bA
�E�4L*D���N��$�Pk��̀�,0fa�<Q�B�@8�ɴ營c���B̏\B�����#D��Rq

*{����!V~2 h��$D��3D�)>qb���
�`��q��%D���RS��J�xRc�*!� l�¤%D�@�7��+Mz�{���S����#�#�Ozhb��OR���n� zX�yB�Cr����"OXE��h_� ~�P
!iĊQ6ԝ��"O�Q��JñJ!����h�s0~ ��"O�Qu�\'I��x���o���"O|��J�6"�g	�SP����"O�ؐ�BNll(5�����<�����ɰUɚ�~"7��~��䉓7S��u�D�<9��˓/0"Dia%݆g��ؖM�|�<Y��N��vH��O�P��k&Iu�<94K1y�21�D�z4�w'�{�<�"�ѥ^�Р8�e٘�~�e�w�<9a�	L��� ��mlP�d���d;G>�S�O&m�&�3A���ʇ��/"(��6"O�L)F�\�b�lܪG�	0��=�e"O� �8��M��G����S�BM�"O����Z�1+�&�2���"O�x�!H#�>Ő��G���  �"Or�9�gY3�1�żx;�9�\���+/�OF�����S(Ф;�m�_�X`I�"O0�3%)��#8t]z5,���\���"O,����<�6|�rj�&�$`I�"O��k��Ȇ6�b�p��F;�^���"OnY�R��-j�Lt��H��xTT�C0�'��	��'n<�)�h�'"fVUlH,��iV"O���&ҷ-��@W�I��Pb"OhDhbcQ-'{�,PB	 �� hF"O�������@a��C �ٝ%�(]�"O,]�Pȍ�^��Y=2�J8˴"O���0'�*V��ؠK�kQv���/£~���U'2v�y���{�V��%��D�<�iT��"�3��֭pv&��2�x�<��g�a�������%����^�<�̕%d��9P�
?m|4��
a�<)�Oߵ'�Pk�DΪ3=��6W�<	e�	h8Ja��*$�>�'�ɟl{qL+�S�O$ty���:��2�&W�2s�EK�"O�)��hYPRQ� �ß��|�"Or-��T)��,H���}y~8�E"O��C�	A��$	?e����"O����M� �z��7t��Z�"O���4b�\.���"�\`��+�Y�D�-8�O^Ѱ4i�epF�(��(�`<K�"O�a��2s����]- �H!*s"O�l��%ۅD�Щ�r%A�9�P}�s"O0q�tJ[�PQ�@Qqb�Y�t�I"O� ���h���!� E�@ǐ4���'8n�y�'�\��	�&�����a�p���'���Q�nk4����ح���'>��VI���Q5A�+�Dq��' >8`����ni��P�(�95��[�'��BD}��՘Uo���C�4D�[��BT���ehF�P��k��4�-:hF�4\�Z�d �T 7|m��C%P��y�����ˇJY�l0����)���y�V/h9R ��X9�%���y�N�QPl�KD	��P�� ������y�N6}�|P��5x�dJ$���y�H��(��Zba�Ex�<{R�-�?�wmDV����(:�KH�@VE��}�Z�k0�+D�£���Xu~T�F��p�
�Q�+D��إꞢ����v�ƒ���R�>D��p`g�"�\�󶋁'�d!2S9D�d��+�Y��sR�*�@Q���3D��*0�>.��)BEԀH.Z�`�m�<�Q��k8��a�S���3�b{:<x�B3D�(�tNQ��9B��&*�p�g3D����%T� ���$\�T!@MxAl/D��X"�K�oN�S��D}$#&�-D���AIA r@��SE��q��� I/�OB��O� :5n֊n�
���-[T
X�"O��ȣF\�`bHHR���3L�l"Ob���g�^����@�MOX �"O* 1`�Ǚm�����gJ�c2I��"O��X6j�;yȮ8aG�w�x�f"O���b��rb�� Ɖ
W$d� �ɇX�N�~" ��=<�a���GC�U��A	w�<y&G�*?�v�S,qb&ŠR�O�<�B��7�K��سM�tz"��N�<� ��6�
�s^e�w+�pa�@�"Oz;�jżBWpYc4j�s-jt"O@���%�0�QH�;j%�L
4�'���y���SP�V��r��
gjݱ�&Y+x�N���C�~�Y�i��C�(U��f֮���ȓ�`��Q�V�⧆)k����1����c������Ȅ�l ��ȓP���[�#R"5�zi��+;E�I��g���S��-#�6pI�>:y��'Ir�!��5�莏]( ���n};P�"O0��K�2���mזc1�l@�"O����ǘ��R���
H'4J�"ON�)ꇹH�Z�����B�<8"Or���18�t����\-
Y����'�n��'l�y"r��@����X�wǀ(
�'f �AtÕP�8�ɀ��w�L2	�'2��1�KP��j1�W1u���'0�`�c�� �8� �)B�\D��'4����D̰+ɀJ�����)D��3���'x+�lɔ��˪`0O'ړb� F�$AK�R�,��l���R!J��y"���U	
�#3����H���y�)��j����ۑu�����S��y�*I����N1�����*ǆ�y������m� rd�꧎��yBC�6=���9�@P4h9�,�wmL�?)EGb���������j�2�J�%=jP�aC:D�칒iܽ����D-E��k7D�H�7$�a�t �E�m@Abņ3D�$K��D�6�ذ��N��%���0D��2c�� �; ���B��k<4������<n2��	$�ަVI��P��<�Ol�'$�(q�On�'��활T�(k �˸�<�+�Z� �I䟔�	/�m��!�����ʢ�?ͧ���D<�&�en]��t�P�1� )�0�a��r�\9b����I	r��&j��	�hp���[�{���!A�O �1擵L�h�Sn�H}��8l���0?Y�"GQ9vp�1��%31�#���`x��.O��	gb߾b�hhW��wM� �AW��3���0�	[y2V>q�I۟!�	I�`����@�+��G#�џ���ȅN��a��IX`��S�O�Ԝ�f��"C���
dˍC~ḙ'b�{	#w ���#bZ�,��?9�tFN�BL��R�'˞au(���.o��2���O���$?%?]�'W�	�'��lV�"�┸Y�r� �'P�P��ê:f�(��M������k�O�.H�bm�m�T�Pԋ�6T��]��'��	�n�E�I�<�	������$��Z6`܂ �A	h���IP�V�2���'��D��O k�D%BΟ�\P�@�0qd�8x!HO�6u�h#)�Sc��� �&XP�/��g�'�4��̏�a��hh�I�q�O X��'��	�<�&�G6`TD��A-=&����UD�<�f嚹�(�pa�:K8�AqgN��d ��4���d�<�i�1p�r�	��ͽA��hs��ğ�Vܣ���?��?�)O1�D�#2���+I\Q�2���<��RO�4|�����,:K�=*S�Egx�T���T7kX����8dԪ�pG�:	��`��X�>c�"�kQx��x���O���:+Z$��Iδf�f��O��=ъ�$��8�5+�e�M�b��GϜQR!�ĕ�,�6�5M�@��m�5Q�	��Mc���dI.��A�~*�K�#����D�\���&������O|�$�O���O�<C�m��ҵ�?�'N���a�V�O&�БAH�eժUG|r���lUQ�0��6*[�x�Z>ic��K�390�J�"'��H��9�no2x���@�|ҳ��4j������I�P��� �ny"�'	a|���3a�ܱa�4w9��8�n����.O�HC���#G�
����J24��2_�(���Y2�MS�A*��d�|*���?Y�U4_�}@e/�3x���oJ/�?qe*ܚ`����A��A�~tz��,׈����Ư�0j�ѥ��J��4O꭪�F�M5 p�C�X0����ȃ=8.�q&�@�aLj%� C�{+��X?������T��� � #A��#N���j�c8� �"Oj�(���F���sS�\&A̤���I)�ȟ> ��5HpR{��ΥIR�0%e�O���O��P�/R���O����OPԬ;�?�vK��1�a��Y>Vd���@�5i��j �'@5*� C�;�^y�͟��H�Σ)�Te���.�R'�"�4��I!g.Q�r�Ӻ�Ο�xzw�N�er9�3��z3�0�f�1?Ig�t��o�'����+ЦQ:%�B�~Ur����&�!�$E�v<l���O�H�t�䁋�/�2,9��|����'�nXR4��R�a�3ML��
��:��q��I7���B�� v��w���<��C�	a]����O�'C�a�焕R��C�	  �$�g�
>�Qpq&P,��B�	#�H��V>�z��,���XC�I�W�JQW��* `C���n��?Y0���<�����:R(�㋱f
�����7��Oִ��
�(�b�9��?s�8Qk�kD��L�j5�ɜ$(l�D哙1��(��%:j<�"�����">9&���p��F�Ӕ�D`"gQ3ڒ�P�E�u�	��?E��i���h��N=+ ����ş:_~�}*�<ie�'\UI�C�ބYh�P�G�Zy2�'b�'i�Z�E4���B�0i�B�Ð+N&� @��o�'�|�aʲ)D��R�J�������O�,)򥇛�94$�Z��y�����d?1��OZ�T>�ɏt���:s�V.8T-�b/ڌw�^���͌M~R�,}⃌��	;�ħ�<Te�o	h1��iO�7<hع�+<}b)���E��'��h�C/	�`�R�`R�C��a�Bdφ��	��'T|�'�N�'n�$���P4L�B1�0ĝ(�<��	:���'1z}ʉ��68L��З�i�,�EQ�
xB��L�}��N��I�Y�O�qn's�D����l��)`�`O�{iʓG��O,�E�D �=8�؂�.�&o���zGN�~��I?ra�ҧ�9O�i�&���S�*"��P�P�Ԝ1*�0�&č/>��8nT�'�� F��NO:Z�ap� #TE��߲�?AAè� ɰj*?��y��?�~�.87��xb%	�P�a�
��?Y�*�O�賲�B:0J˷��+T�F��*O:�%��7ig����ݜb��`�ܴ�?�����$�O��|�+��J�t���Jd���,)�tq�AJb}�|�T�E�d�	��УI��Pn�4��.-���hO���Y�P�ߛN���!��'�8 4"Ol5r�a������⇆�w��k�"O�ܳ 'S�v�\8��K�N�q��"O4ۥ�ɶˆAA��N:M�ɂV"O�I���H�!D�he�>��H��"ONI�e�ʹMG����$�5kȦ�ɖ"O$ᢴ`MPzx`��k'}�
�'Z����J�d���{�
A?"];�'��Q���Q�<R4��+	��p�'-z�!��:wL	�p-��;
�']1�`D�G6\4HA�]�����	�'����L��h	f��tAӏ�a@.j���C����88$��ƅ	.�B6N]9n,��k����!�ti�P�!΅WP�V�ɟf:���g>,N8�2��5_�d,ȅ'�H�c���/?�	S5��JmPq��A7h���9��ěP��0
���� #�H���|��
>z��� �\��'�:H�§	8	g������ l���'�f��G%� (�4kB�L��'�9�P�ts�x��C�5�
���'� ��<y����n�.)n<"�'#B�I�Ȑ
Z " 
�.�(Y�P��
�'h8�I3g@�Y�$�3q�%p~<
�'�2e���]��	j���j���	�'|��$K5g�������s,�1�'�ʵ*e@���i*G���M�ʓQN0yu��P�����s�V��ȓ!^�T��y+`)$n@�qk85��)^�� �.@�T�n`������y�ȓi۲P�DgRD�\� 
��-����S�? ����;]$�-���X% �r"O��cRmˬ<n���	H�"�"OHxw��o�\���.�;*l��5"O��V��Pr�x��L�x�D��"O`�J�B�V��HI���b��}��"OX���Ƭ.���h��A����1"OVxbP�Xʄ��Nˆw����"O����.�9Z��x&Î9ei�1��"O\�0���<NT���ₔ
Q:���"O�z��Ji�$k�kE<�4a*�"O�I���!9��!�
�!+��U�`"Oj�w+^�0�4Z6i3��yC"OR�#i�'�0�ӧ�=AH43�*O�XJpDA	"{�M"#o�:���'S�P0�"��tѨ�����#_�9*�'G�������]�*��.F<G�.X��'�n�a%ʤ <h��D�=��b�'�zu��͞�
E�A��@R	l�5�'CBh��m� '������F����B�'Z朋�뇿<����1��� A4T�
�'�P� T�:0@��gŤI�.���'�u����2F4�a*C9�D���'���`T:O��L��.P��	�'�x��/N�b�[�&0$1�	�'���T,�����,Mx�	�'N�*&��zRJ��U����`r	�'��a�9yY�=K"m�.*��H	�'$� � � w�ȁ6)�����'H*�R�B�zX��@��}a�1s�'i���WI�@I��#'��*Hh���'BT�Ơ��I� ��&�1D�f�k�'� E2'�;<	�<�� �@�����'8�xൌ['=L��U&�3<����'uH�Q�Q+D��5��4q�
�'�Dۡ#E�i	��'�®Z4�
�'����,R�%sX��/^�|f� 	
�'x��*fhI���yCh�!Xxl��'�.U�� wd�C/G�`����'��J�-O��z�GBQ ����	�'����5�ʠ{��H�6��n_ڴ��'mց��`������cP�e�n�I�'�l$��8�҉��*�2[4D�A�'�ࣦJ!X��4���T�����'���:�)^"D�@j&QDx��!�')H�-Z�I%lAŚB9BQ�'�,t/�=7I���Gȃ90X��'��8��/A���"�/]� \b�'m�3�Φk��}�1�\�����'�B`ڰ�Ȃ=Ht���C-cT@��'N!�K.;n,t ��Y��8A�'�ļ2p�ݲ ��A	��Tzv0`�'E����h�/B<�!K�J�Q�'�j}��&E+U�6��T'��ȶl
�'�t�7�+� �j�I1����'?�dY��E9 ���FV>)��T��'hJض�C�z�E ��
�"tx`�'ֆ�+����e�D��L`�'��d���~�uQAV��n�Y	�'�:�Ib��Ԩ;���"u"Od|�GͪU���H�2=0`��"O\�JfEZ}�{֠
��;�"OD9&ݴQ��	K�hF81�{ "O�)[r�]=0�V��7b����Qe"Ov|`C� ;:d��W�ʙr"O� V��`C׉ؕJ�* _�~��"O�a�/K7 y�l�U�S�r=���C"Opx�a ��o��<��đ�-���s"O�p�w��(j��䘕�T�p|fx3�"O.0�*ܣVDHM{с�$X�"O�Q��2qdL�I��4���"O�2a��i�Hċ��W�-�����"OB�aQj��>��9u�ݖ
���B"Ox	�ej���l�j�k�1D��ݲp"ONٲ�x$Z\I�H�8��{T"O�4��ŶC��xc�I	Iz���G"O�����	�SzM�W"O�`ύ�	~D��G�?{L�
�"O��WÓ�,`,{�F�RK��c�"O��sCL�)=�ج���D�52�"O���c�"2"�|J��j�9:g"O�s���)��TD2
c���"O��qn˕}�	����wK���"O�bAiG�V����"�NJ�1V"OxTh�č�0�:�A�;r���HW"O��!�Ƅ��z���xt�H�"O(p!#2���Y��/	g��J�"Or�A@I3Gl^��R��WWFPv"OY�r��<����e��U��;b"O�	f[�>�ҍʇ"M'(C�7"O\]��)�0u��Iׁ�>-�1#�"O��ʵHUGQ���+�{Tع�"O���E�ؚ7 �a�k�ms!"OA��@!S ��3�]1qL�ɚ "O&Ydk��-M���_�^�r��U�y"�\�}��@�sdܽ:z��gٸ�yR��9�x֍ܶ,c�D�3.�)�yr�
a�Ra�R� '����*��y���>=��ۑ�X�N�t�G'�yR�l�D�W ðM԰H	��'�y2k�!*h0gL�><�j����y2G�"f+��
�&2J�i�m�!��
H�X��T@ٚ_z�:��Z�{�!�DX@%zT��%[ �"āL�!�Rtp~p*'�3CNjP0Î׉}!�dJ�)%v�C�AF @�G��_�!�׮hK(A��2+<��&Z~W!�S�5� ���H9i9N� ��,�!��+s��K��Ԃ	���e�D!�d�O耐:��%{m��/EI!�C$x���o�e �G�
H!�R!�
<�0 gIC�%S.5a!��ΰ$��mБ�ވ55ibv*�MQ!��'V�B�!SmF![* ���$D�!��ǋ�B���  {�(T&pv!�->�j4�'hE�9z@qr���qd!��Rj��$����	x�Sb@U�tN!��!Y���"al�U�"Ĉ0��/[!�DI00�	����!��8��ܷCr!��J'-BY�@���B�*T��T!�$c�����C�n�"�Y�b��!�d�Q�
�q��.-��@��vz!�d\�)�6`��_�N�d�b�]$f!��,
y����L�nX�s�B�DE!�D���)ˠl=W�J؃4��'-!�D��v�d��v��
~_,�2�jC x!�C~Ǡ$2�	�b@8���HU�mn!򄉎\
�P)%��h=�!��{-�ٚ&��>1q�ܒ�(�3 !�� 9��:�ܤ���L�lTJx	"O�@��O1L1f/O�xIp��"O�u�7������4΃<?S
�w"O�1ɶ̒�Y���B�ʞc��D"O�x����c�
�:e�,�a"OݒEgŭmu�T{ċ�;e`q�"O�r��W�)�
\X���1~����"O���w�M3l��[Pj> @��x�"OtA`v��!��=�H�2ɢam"D�����]�AR�%�kЏ:t�$D�@S����mHhPX�'Ͷ3SDq�3�"D��� �F�|�&hc�K�1p��;D���ga�
F܅��,I;[InYXҪ-D��i  ŝb�b����DH�&D���E�=6׬x��(�-;:���j#D��Cg��(��E�6u��WN D�pQ�ǁ9ly�h ��#]Q�tWE;D�0ҭ�+���K��(]p�T���:D��ⶣ��w�T���R�C����b:D���j̕a�ѻW�nپxb��$D�`Bg!�{�5;�D�>���V�#D�X�T-�[���#dD2�v|�TL%D�D��Imo:�C5C��bq2Ic"�!D��b5||�(ac���6���>D������3jJ��c�Ypd�:F�8D�x�b�^�)����B�e�mIb#D�|��E�0S�X՛1JՁsˈ�r�M#D�0�L�5Cf�9ie��"v"�R�"D������MIX��2:
�@�č%D�D����<������-�~Њ�`"D�8b̒@E����+�wH`�T�?D�ԯ��J|��#R������g���y�L�m�b�*�B�	��l�cះ�yR�_,�H�+,�r�K%���y¥%=Q�A���R4'��d��ۯ�y� 0K��d�וo���h2j��y�Z��Q�-�Y��PR�T��y���9���w�$7������yB�ѴR���Ir�K��xQI�J� �y���|�(}�R��\���C���*�y��?L�L�1P1RW~��۰�yr�׷*"R�t�UE/�(�(֫�y���91ET�p��@<<��� ��
�yB����h0B�J�&L����>�yB�ò8��!�i�T}����4�y�#�����΅�>����-N_�<1�&�/0ub0����V<��W�<�����U��#�m��(�ϋV�<�`�=����+���
\h��^�<��L�:9B�rOݤB=���R��p�<a$�G�J%�B���i�8��c��g�<��D�@�!d�˂v�v�`7�W}�<����2t(*���)
�g���Q&�x�<ɣ
�"� �rt��'<���Or�<iqLZ�uine@��Q�u��B�<�w��ZVQрBO�V�V�KC�I�<iL Lj��Qd�D&8����b�C�O6Ip��I#0 �aSA��2se��$�8@���'o�:���ٌqn�ɱ�K7D��#ň'd3H�
�A&.��*�k:D��ᘀ��)k�/˙0"�]
g�2D�8�SĄ3:�^8�CWj���o$D�lJe`В\���	��)z|��!D�\�',�� ��xJt��u�ۂ�!D�h�dB]]��{ӌoN�����;D�� ds�ဨ+��bhÂk��M��"O����Lږ"����%�3�-��'8|�a��P���x�}mn�	�'0z\2��O1h�0�9R���#s�X@�'GT�Z剕�A�H��'�M����'�eZ�-�$^���e�[�DdY�
�'��@��N�R�tMw6�H �'Ͱ���,�t���T�Hn�`��'Y�D�6�U�=nt��J��g!V���'���P��߭$/p��O��nQ��Z
�'7F���f�O�� aC=t���#
�'�Jeɤ���p_t��!A^�n�tz�'Z�0���'8��� 1�M�"�#�'��A �Ωm�V��P�
�*�'��m�eK�'q����$	H����'�p-b�oP� &έc�#n��'�P��]��,���5\��a�'}t(��.�
S5�V��n�\�3&D���2�|ڄ�:RXՑ2/D�h�. D���Z��M�_�V�b��,D��Hg �=3�.�r���X�>M���*D��	(äg9h��@�� ,ɪS�*D� kׂU_�#�41:U�2J7D��S慍">lm9�(��� �:D����A��jL��Aʙz�j4��+D�����#~3�Z@��h@��{�<��`��l�l���R���^t�<yfO>2��7�Q���A��D�<!�^_��(��TG�6�y��Z�<���q��V�\˒٩�X�<��lF�<4� ��fP��9o�K�<����p�9C���^ʈ0�ƅP_�<1�K/0h\��A��bᰔ�W��e�<Y#̽�9W�ٗAx�XD�G�<)�Efx���͛&ˈ�(�A�<9P�Q8�� �W��ԅ�X�<�Q�U�2R��5���X��\T�<� �L7V�zU8-E�iy�@��AS�<y�0Ӏ*�#ӬE�<��ff�<U��2m�؅�&�J�h���a��b�<q�ɒt��rb�%_�]ڲgQ�<a�C��iXг�#"@N�霤IQ!�� >�x�ug҂L�8D�v-�5%!�E�'��m!w�Uzf�.!��fG�a�"*��=�B 
`P=!�^��>Ʌ@��"�zM8GoHDt!������,H2�|���M&o!�қs�l8X���1\ö�j��Dp!��̅8(���Ak�4�) N:AS!򤄊6�ơ�c��<��8"�M5tO!�Dmh�*#�=o v��L�o�!�ص)�����٨a�$:R�R��!�䄆��$
�N�9�^ ;g	q�!���@���PQ��R�X��E���!�$lO�=Ѓ(�g��k�%	)!�dK|F���΄�x7`���ŝ�!�d
�t�Ra�~ƌ�z�KbR!�D׷g�V)A4�Ӭp��DJ �&Q!�'8�����
g��Qǉv!���,c2��%B]:%��Ʌ��!O!򤐁2
8�j��ت4�$dVÔ�6�!�d�V��i�1&�D����� �!�Z�jb�QcQ0^	�P��N9iF!�Ě�=���`U'Z"ȑ�f�+hB!�� �%�a���2��Td��8U�)�B"Ol�p�
@"(`�`�d�]8F-,aj"O�9�f�ܗK���ҏ��R,> ��"O��D+^�����-Ό�>9Y&"O��T.�4���o��HH�	2�"O�QTL��6���q(��hA�Ii�"O����K�R�	�A��.���r"O`|�7�D�rHZ�H�Q��R�"Ov�IտS�29��.ڄ%���Z�"O�8*7�
�:8�Xt�H"1N���"O‡���[|ƵZ��C)Z�����"O`(qAаJ��LYRj�@�ڝ�D"O��b�%�97���$�ȃmN� �"O�!��Ù�m��Aʗ�Q�S��І"OQJE��jc(y��ޞ`�t�A"O��r�F�R$�e��܄�a"O�ly4�A澶��~�"Od�g��
w� Q#�Y$av���!"O���Qb��aZ%䚳dg�U��"O>���'�#kFrc!ި��K4"O����hZ5O�r9
�
1"�̑c"O،8��t���X��o��8�"O�	vK�9W�$��ʔ;��r�"ON,#&�D<->�xs���M0Q"O�p{�%�D�ѱv�� b�Q��"O�b�&��'֎h(a�@�|��أ�"O4D)W�ګ?�h����"�Hp"OL+fLʘ� P;�W�Zt,�S""O��{jτ*�^H	�Y)6i���e"O$dbb+̻D��s�(��p��"O��`$j����1Id`�5�h�.���$w��]0TgG&@��Q���E/[����"O�YIąo����ai�<��4�'���<A&�	K�<�!r�"bʠ8 ��	t�<a�O�jb=����ˎ���F	wy����M[rD]vʸ��#/�$h�9��gKz�������'�V��ȓL ��y���&��L���ͭc�)� ���G�m�ɴh���8���b�3�\�r;�D�=Sz����
�
���KC8����./0n�92�_�+%+�߿r�>�IÃ�[������:|O!ڲ�1I�%�$���C��E��ɶ% �H� �$L��'
7�ɖ�D��,r��B��SU,$�yZ�P���
�hM/=�]�J0�~�G8�z�c��J�z�`aB%W�m�>1��US���Q�C	�-�ʧ�:D��0 Y�X� Ѣ�J=x��TY�A����� J}�ՁC\�E���O�OL<�'`�@Ƙ�#�8T}^d�'���2�ď 	�L]r���0�TZ���Dz|��������Y�EXa{��P�g�9�nO*,&°1���O�tNرk���f*�PîH��`�]�&7R&�*��Ŀ8:�HT�8D���dI:��M���k����#���{�dZ�`}�Y���X�
�j�,}�O0jB� �p�z�6��%�	�'�:,S�]-$m�l9�U�ig��ڐ��U���@�Nʶ3QZԙr.���g�zb��s#�,s: �X�A��Y�4���� t�����RC�d���#M>�$!��"@HZ�(1�Y6m�<<���'N���v�D)I�}�#�M,^���A���ʙS%x%���<v1x؁cq>�zvg�MU8�q+T�p��7l+D���:h8�ݘgJۣwf}` �<�rk�	-�X���8������8e~HҔA�k<(���X�,�!��]�bppg��%\:�W��T����`�F��LIJaaAj�g�I7K
�i�Ƭ�2j�-�`��.`C�E{89���O�yE
x�k�2h����I;���S�'��ʇ�^ ���G-��N�L�`�����C%�����>�X@��m׫
^�ɩ��	&�!�dK5PmB���呹3Q"�r  �X�qOR8@8�)��D<l�����z�ʙW)'Z�!�� ���pgѭ���1p�Y�%�Ҵ2�"Ox}C1a]>]�r]�6d	*u�Dxxb"O�(�0Ή�5�n̛�薂w�x���"O�HҖ�C�c����c٤M�U�`"Oj=�g �����S<����"O�mCT.�� ��p
b+^�"�Хe"O�1�1�S(Z4hD`�Ajx�"O��jN_�\^��b7��\�����"O�]��j�$��̙���_?zY�q"O�$rQ�D�v䃒�q1�|k�"O��1�B<r��8�����P�s"O�mK���d���C,F>+�0�I�"O�UʷBͺ4U� �n�&8�v��"O��n��M�F��-F�	&���"OV�@0a�z�ܩ��̌�(�%"O�}�D)�1-ی�:��7
y0�"O\�òb�-���v��+a�TT"O:�*bF&�\���WYt8�"O����S�.�n�רR!?V��"O�]��h �8���icjK'St���"O�,h1dֈ��Ѻ�cK2T��A"O
(a`뚴A�t�3��?�|�"O���o��N��5��(^5D#l�8"Oy�`��,?L���鄊d�`h�"OXM��)"��%��H� D�t�a"O�(8��
��!��aV {��Xa"OR�D�(;vdaZq�=<��M�"O���v/"x.���E�5\)~�"O��#d�&v��p��#V�p�"O<0q"�J61S����T�y�1C�"O�MBIMj\0�ZE�Љu:H�ja"O��Sf�G���#V�Ȃ+��H�"Or��K�(b,<����yBLyr�"On�۱�ƽxM�����/���r�"O��YA�7�~L�0��J�8A��"O����L��*m��`��71�V ��"O,L"���u�Ѩ��]���PE"O�8X��"5�`�f�C�}���*""O�\h��ܓ~X�8�ة!�,�C"O����W>U��q&g�)��)��"O�����P(���G0+���"O�%��� Ne$��u�*Oj�[PJͼA�f�"b�O48��r
�'��oE*(_
��IC�c�����'���AG!��6��0R$��V@��'�`Sr�J.s%"9#Ȅ&=� ��'ⲝ�bD��8:����(-[:z٩�'�n�Z���$xv�	ѫ�0Me�-��'��H85H�394e�0CΫ�� ��'���[�$�|��|�#���t9	�'lXȂ���4T\�
�#U�5p�'"�L��9#��er��Mxؕ��'�����
�?=�U�BI4kF]�'Z-��	�8EK���jR..Ġ1R�'�r<˧j�?��&�[."����'e.�`t�\)r���D�ۣU��s�'�����Q%��QT�]�N��0
�'	&�����|#�:I���
�'j�4( �@�v!���Зv����'�J8��!�EW�0��P��V�q�'�S�k�&��1Y�h�O8�	�{2M��!�n9�Đ|S40`������&��0A'�F���'��N���jt8��iI�[�B�`��-Pz(���v8hrƓ=�`D�Vf��i�X���S�? �U���Vt��Ǘ�~Ȁ���"O�MR��"p�k���(8bV=#�"O�L�vC���ax�G�3�rE��"O@q��N�L�tH�Ƃ�M�IkA"OP�æ�E1�P[tE�w�H(�"O��`�"P�Y�Z��8�`"O~e2�NzMt�0BJ�9$��f*O�u���m���� ̵8��Mx�'�q��T�P�I���a���$�2D� p�J�H���@f !�R`�W�,D��rצ	uk���t*�SQ XR?D�$���U� @Jl0��N�"�DECׁ0D�dI�g�7~�QJRv���a.D�l�b%�/u���[�V�m�0�?D��b�B::�PL��d�gp��0D�!D��`fm��f�sc�Փ4���C� D��E��Ufp0��/,v�ؒ'�+D�L@C�Wn6�{�ѵ;I�L��+D�,0Cf�G}�2t��:n�ڀ�4D� +0N9c��$�bS�cʲ|*��1D��x�$LK�֥O)8��0U�1D��83�Ń	i�\�>�d�j"�5D�Ĩ�ӠLj��{�,O3D��I(D�(y"&�8b"B5ht"��u�Zd+Dg9D��9C�΃Z�*� IC�y:�c2D�\�)O��ɋ�'2�� o3D�L��.�&Sʸ�dbR)k�,9�!$D��AmN�)�<[b%,� ᣷�&D��A���.hH�N��@�8 ���0D��j�E)tVu�p�H�H�.,#C(/D�ܱ�D�2&�:��R+�`�&�,D�����Y�^���e��R�@I�*D��u�F%`ׄ�� e�zV�q">D�̊�ǈ��4��C["k6��0�<D�0�ޕMP~HY�EV0D�5��;D� z7oO)3��QG�1-4F�Q%=D�,Q'��<N�p=�^L�ҍ*�y��P'~����0D�&�[qMU"�y�2@f"pj#"Dv��`�ĩ�y!Ğ6�\�3E�G=4��q����yү��2����E�d�M�qe���y�1:P�5Xˀ�`Ao���y�bڒbNҕS�݄"xy8��A��y�-<`/�<��Y'�PQNQ��y�K"kUFXF�<#-�ɡ�����y�'���e#@��~��f&�$�y����0:�nԫ  x؂�N��yr�C�!D�H4)�b�-[�Ɠ>�y�M0.:�!�ω1k���sȂ��y2#P:#c�X��k�:�T�X�J
�yr��$k��$�$� C�����@��y�$M�&�Th�U"M,P2(�G�� �y�
4k�M�4�Q9)�M�5@��y���n��1� HY�R	�����yb�2T	y�!���Pq�t9�G��yb���@��@˲!��� ����i��Y;ĉ��@�F��f�P�����ȓM(���	��y���пT�`��fl|\�A�,{H�@�JJ�p�����\h��9 �t�AVH�.d7N|�ȓY5�)�/£Dr޸*7@'p�2��ȓ$S�Hp�Δ/dv��L A�t�<���ܒZ�
A�c�R /C��A5m�n�<9ǯI��A�E�v�mY0�Sj�<� �\z��\�*�`�fF�t���!�"O0����_%*ҕ"4�[�/.���"O��� $�-W]�H���ݠn"��A"O(�3��H~����P�N0M��"O�AC�D��VE�#P(G�|G"Ojx���D'<��B�����1�""O� ����͓7���b89�"O�T�g%ӎdq���#O�3e"OJɸ�8KP���mY�K3"O�]�6*Y�]C���&�E>L�l��S"O�A�3F�?3�UR�@@�.q=Q�"O��g>8uVd�c�O�ZNMA�"O´�ƀ�.�V4;��E�v0�"O��:��&/���񔥓/c��Iu"O����J��+:��գ��v�xa"O,�#%��q��0��H�*d��"OH=�B���?&�=�4Ex|ʆ"O�H��-#D��Q!L�����"O�1�Q+�r������R0P`"O$(`��� ��4�	D��rq"O�uC'��6U�#�a�x�$k�"O�5��L��M��X)9g��k�"O0��tΌ>Av���-� cW"O��f@�гO
�p
h�V"O��jK8bD�r��_��RU��"O�|�'� ���@ �3���x"O,��'�ԃ8�
8;Ј��)A�D"Oj�Y�D�b2�P��Hϰ�%����y�%[o��4���$4,��Ʈ���y"O�1��z�&��9�厹�y��8Dt�+��W	��d��Ɔ�y�*!����F|[>U V���yre�m�>�:�bUokv,RB��	�y�H��.d���\-��RaA6�y�X@��)� Ā�TiJ)�)�yrK��<�*�N�P��	��e��y�0�pp�D�IE�-�aZ��y�\_9~T���m-�U�WM]�yR��/B8b����Īd�2!�B����yB'�9f�ْ��cL�8S�@	�y�-���4�
%28㡌���y��T�F��}� � }�~�:�'��y��'�l(�R��$����n��yr��T d-ԣ��%Y�d��y�Ĕ�Jur����Q���Ś�	M��y2'�/>�@̋��\m @Y6�Z�y��\.7�0x�_Y���j��WL�@B��2*0�fU�vh�V��x`B�ɌU4�����,3��Q1 *��4��B��WN~�C��W3���s,�k� C��	fj����K;�l�1N�k�B䉷{��`D��Q�����K�3`l�B�I�I�dRCg�1��y�B�C$�B�	�"x��q$��af�AI�jI��B䉲<rN���$��k��m3TKX�d��B䉩!�Ե��\7PS$�H�cՐ0k�B�I	1�B��ץӟ�H=8G��

�B�ɨf���फK�t�h�đ>L�΢?Y��)
g>��uL�.�R�`�a!�W�2���#3�1^[��q%'�*M!�A!��X�@���IZ<x�2�NM!�$�E�0�PÏ ;>Pi���Šc@!�DV	E�(1� ˢ��0Ys�_	k5!���K�r�G���3��h4��&!�� �p���	-i ���n�	��e�"O~p�M��h�<���lU��~8;�"O�,H�⑄o�����3�
�*�"O�X�#�59p��N�^�8|:a"O`�J�ˬz0�@�U�\�1j�Y�"O"	�e��Le�$h�K_ 6-�D9b"O2�s%L�-
�#E�̵t"P��"O���M��`_>Yj!ޒgv��"O^%"��4;���!�Evy�"OR�{�g��1�Ѥ{�x �"OB��B���a�V�Y�8J�l[�"O�۠�ŏT9�@����D백��"O�\�!�R7_��c� K0��"O��B䝮]4��ġ�"t�`�C"OZ i�Ȑ�@�������t<���"O"=X���:5t%ꀊ��NǶ�+%"O ��E́
R�:��U�L��"O�iU"�"E2���*
$���"O���O��QԚY`ß�V��J"O*@ ē�h�
-�3���P���"O��1'�X73��ȃ�!Ls�]+"O�@H���4+(�p�DYl�A"Ol�8S�QkQ�a÷��.��l�<q��F4Y����� �.�!*Ї�e�<�Fe��{U�m���P�2��x�a� ]�<�6�4r�I'�״v�L�a�s�<�v ^�Sa ��/��W�(��&
Qr�<��+��#i�ժ��6؜$QG�h�<Q�웻q�P��ǔ�����ƣ�[�<��&E�j��S�JG;~�@�G�@V�<Q���#y��7�Jݣ�L}�<�d�d޶�3��B3Rq�y���t�<y�Á�[�4 Y�#K-I�^�pb�\s�<�Ӈ˲m��`(�*��xl�E�<�6�d}�DE/�#vذ���\�<A��	"uJҽ�S�Y�k�p�q�Y�<�1��-����K�>��x�KL�<�����a���@#�=o�����b�<QP
^�rpY�f�8���E�w�<�4��c�6��0J\�\�"0Wr�<9��K��嚅H�2��JU`�k�<��-6Z��e݂E^<���Qk�<i��L!x⦅J;_������Oe�<�`�3^�J�K�X���e�<!�O�6�F�B5��� ���ZC�y�<�4ᆤW��E��%�?bm�XZM�<��h�;yԡ�$M��!�>���F�<��tk��"�3)��D�"��k�<�`.�'�����/(7x���CA�<��	�3��As��/7���bC�<��b�{��!FM�(�=؀��}�<�B�V(/�4xd���6�Xh d�n�<�&�1p����_|y�p�ƪ�u�<q"�ExA$|�D�هf�@��BkKr�<I7)V�=M����
D��ڳ�q�<q���5�@�w�=m'|rg�Pj�<�EN�/=�Tjco��y/6̡���c�<a�EE=%r�����p��R"�y�<y��L"�l<@�(Z�i�n��1&�t�<AcL��4�P�V��2��h:��Gx�<��� 9���j&�#0 ��y0�T_�<!�n^,	�vHP@���aԮ[Z�<�
�I��TK�J$}�YQ�b�X�<A�/΅zL��lB9V�:�6��R�<� �Q�'։za048�쟣K,&i�f"O<t��b׮};�pa#+S ���a"O@�t.U�kY0���9�h)�"O4�ˆ��,R��A�C�3��1B�"O��vIK&?/�Ղ���	1~�da�"OjY�e�
�RQz���K84t~��"O4@:�d�#,�؈8Ջ�&n ԡ�"OX�Ф���3#��{�m�1g�:9��"OHc�^l�F(�RC�?p��H "O����_(�jF톇ye|�HC"O�XDG(L�����8MV��[C"O��%�.b�����F�BH�%"OԴ Nw�+`%�,+$��"O&��҈Ҭt00hBWk�S2�cd"OB�S!�t��=���φ��xk�"O���3/K�;���@���#���"Oh���j�\}��� (�)r�L�@!"OnE��IJ�
��u"�e!���D"O�d�á�4\�R����ت��(5Z!�$X,#A�\���5\&Vybj\�qC!�d^�z������Z-+ �Iq� �c!�$S���x�ã�&��p#ņ�xT!���$�����)Xn61��G��!���<�"�	5DP(y���b��1c�!�DB�3.�[2FT�T�$d(�(��;�!�d�!FqV��V��IH��HZ$j�!�?_�X��a*�A��UII�6�!��J�Pda��?+{ �K#�ſV�!�䘵W��X�p� pD��/;!���!3���,�ULXvE�p(!�0vέ#��ʬmP�Sg��~�!�d"o�����ơM$���!_=8�!�dX�NB+�/��[��	ӀaI�Ou!�(���j���b����m�Ai!��A�g�x�� 
-!frmY���IT!��`�X�'��bl)H���z�!���$}�%�ł"Y:(z@/���!��R6@���&�A��p��G��)!�̤P,4\�&��.}*u9D��UF!�dׯa[�(��ڛZ�N��dfO7)!�ήRn�����{x�����iB!��Ĳ:�m�W�@5+g������O<!�$�3ʢ��a_�D���&��>\�!��R )���XbL�0@��SF�}�!�4��*��]�y�l "�M5e�!�;b����LaɉS�F?B� p��'6\�������"��
�K�'�@��u�^7�P��+L���!�'>�qБˍ�L0�ڳ�ЇK�<�`�'����qd� ����eB��k�4��'�|�ا��>6��a�P V/]����
�')�Z��ø�6�� �W�bT��'��U���]�i� �B;N��HK�'�(9����X��� G�G<az�'"�Ei�l�I5X)���ˏI�t�0
�'(۱��U�z`���瀲uX���'�T|ɥ/��n<�( �@Q$nJ6ճ	�'2���S�3�b	�'���"�Є1?��� %<.n{	�'�q!�	&��`eO���9Y	�'�{���z78<Ё��D����'X��+?��(�����l)�'F��1"H���f�Q 
�^"��',"-�@,���j���y���J��� 4�!�
+^��6�KL�,)A%"OdE#�J��nC��P��i��y)��<D�t�С1��q�0���O>�y� ;D�p;f�DLr�\:��ެv?F �ӊ;D���A�O$x>���GH�`"R�!T*O ��ӵX�F�Pq_�=�&"O��[�ʉ�k�ẕ7�
gl��
�"O��v��f오`a��&bP �"O�p�7�ΧF8��I7WV���"O�P��d�rFh�i�jK�Mj��	U"O�1QTcD�|����m_��3�"O�Ț�J"1��Y�f@�LW��s"OBp� ��3�X`��Q,I?��0t"O@�� �UU:��A#/�ĩ""O\94�(i�@� L�"�4\��"Ov� �� ]Hظr�ʺ*�cb"O���_���gl]�;��ɀ����y�ߝvZ��W�28��z����y!Xp���Ub� ��=)�'P��y�
X:h��q�~j�\A�	=�y"�W����q-za:6�ֈ�yT�pG���wu�F
\��y�� ����mj4Bq!�����y"i�7-��*#$Ƃc��� 
��y�V,'���Sk�	a>�h$a�ȓ5��&�ˣ��m�E��9���)�\���&ʠy�(i� rk��y�o7i<#�'��5?��!��y�
��V�xrLA�4Z�L��O@��y�&�Vb�@*D��&)�޵J��)�yb�3h�餂P+'nIJa�ף�y��۲'��-	���i��*F�y�_�P9� [ (g�@+W$R5�yB�H�� GGP`�f,�rm�A�!�$��[Ƹu�e둱2�J��İ]�!�E3S�<�c��K! Y"0�P�p�!�Ċ�P�F�b�nI�G�2X�Wٳ]�!��;�h�bo��8}AgAܝ&x!��<# t�U�'Q�ơA�3_k!�T2Q�uK07�
��@o.VN!�zBLeS�%X�s�*���gU�5i!򤇜C4�Ë
A�rak`��#N!�D�xOx���F?k,i��W>u*!���89Z��Ğhj���
��E1!�d��[��uH��Ǉi,��۲N�s�!��?t$���_"�<��!�*z�!��J>A���ր�1#U��k��!�d��7V�ip&M8N��R�T��!���$z�~��ҥ�-k3d=3�F�'�!�X�pRz�qC��g%H�c5�/*$!�d�ʪ�Cd�0�A"�>`�!򄔼W�MZ�EU#V���"#+O�|�!��V��bF��B�4���D�-�!�d�z��)�͇i�|L��[>1{!�t�U�`�c����tذ6Y!�d]�/aH�X�����Y��� p!��76TX�Tk�������	G!��.m�<��s��<r�"��-J�G!�M�.?�� e$��|��`�Q, !HU!��_<^s΄2g+[4�t���G�!�؟
��)��`�"S�4�svE8�!�V@�ܬ�V쑟vv�$�A�A��!�͢j�v�su�_�;a���wb^�V^!�$L�w�ƀX��9L�U���ǲY\!�� 2�!BGa�&pJӭ2+���"O�둆�h�4��#��&!�]Qw"O̘:C�T�M� �]��d1�"O� �'�Z�7'<�QF];�n`��"O��R�	��M������6��q`�"O�:gB�	�PK����p��x�"O����*�LYd�Z�`�ņc�<Y��F=u�Z5�2�>����]�<A� �u��]K�֒�	`�n�<udО50�3Ƌ|�QQ�"�l�<Q�	`l�ȉtA��fE
��Ȁi�<�r��&��	cܮ$���nIJ�<�kV,Ye�����������Vk�<��o��T1���1` aE2T���ꋽ=��TRs�դNk�1�V�3D�DA��L�] 
 6���Vd���0D��Ƭ��G^�M�!mͼI��Iq�0D������&L��s$�*R~ta3 .D�,��O��w���#DK�B)rȨ-+D��0R�ˈ.wX�Ȅ͉�Qs:�Be'D����Ė�!��4J3<�l2��!D�hi���H�u/;,`�E2�#D��Ȅ�B�N+�q*׌�7- �hc� D��B�	h�Q@��X- Bd[��:D�hP'#	$xlA�NC�4��@:D��ye"��.�v�`Q	ǜR�ĕz�m7D�8�6 �6&��%��iAL��fl6D��JQ-_��-J�Lש��ux��4D���S�� JX���V%wb�䒀,5D�D�P%�X UC���oZ��0�D3D��X�L@�#���Qb]�m������.D���1H!<��\����!Ȑ�W�!D���T�̒g��¦3~CX͘�*O:�+��\�RDp�
t�	9bn�5I�"O�R"�P%��B�a�"t4��"O�q�G��vL1 ��C=D�0�"O!3dH�z2H���_,~2��Q�"O��W��s��U!�D_=nn�k%"O`|����n�ܑy��O�]���1"O@l��.�1:x��p�ΗGر�1"O�5��I��U���.K��M�$"OԱ�r)$'i4��mB%G`�3"O�(�O�D���C�R�|���"OJ�Ӓj�o�^1��`Л�0��"O �g��R��<(4i�)Ъ�yRł�,ټ��l߅_6�A7!�D_�>�Q�mO.Q�~�����2!�$Y��`�A0�Rz�X���	�/�!�z؉!��Ӱ����f��F�!�ڪ�n���L.K�,�K��'!�!�W3\"��ZQ���.a�3oM<"�!�D;����,S�|�t���ܯz!��(V����R�ި^꼵�ǃ*	=!�䚌K�l�+P�H�@:�8�(̐LE!�ގ:����F�ȜZ7�|�`�Y�'Z!�D�/f���c����!�TG�S!�dW��zH2G	܃_�� �DO��!��ݞi�ع�C��@t1��
R�!�d�<(
��-��D
&hޭ/!��@�e�z	���E�:;�f�;t!�ǗY�f��-G�N��y���%Co!�DG4\�T��!޼{��l@G"=S!�$Z���VB�Q�n��h�N�!�Msi�8����c��E�!�� ���Ņ%!�r���Ա{T}��"O�,�0�Z�>>T��[b�"O@�Ӆ]�]Z��u��3!Gt�*�"O�Ā6#;M�i���=����"OpI�2(�� �VE�0fVH�%�����*����>I�f�'I��X?1C�Q|���A���,��0�3��T����?���-h�(
�7���R��+����`w>������8ޠr��(�X�`�;ғi�0u�2ʑ=���ǔ�X )�N���M�C$��`t��iT���(!�ft�'/������?�I~*�4��4"Â���!�g�r�y�p�'#�'����'&�b�́6AD�c�i�7Ԭ���'���'����A¤�#U������u/
/�~���'|6M�OB�ħ|��+�1�?a��M����>T�r�iTOT�KPB�u+�J��i�v��f����V�
j�LwYe�/�l��q������EX�bq�X�c+���u�gӲ��
��FZ��±J�)#���ഥN,6�",�~��b*>�B�� '[��Rc�-AAB�l�<B����Op=�����ix� �/&��`�%�WM<�i�'��U�hF{*�(i��>�83cB�j������M�7�it��ݚ&��@�]�ݸ��ԃ�T�����?A�ID�Ux�<X��?���?�7_?�m�*��\�c���[�2t��
{W�)��-ϸ	���F���M3��1U����G�'&i��N�977Hpڴ"4n��{"埆s�di���%nD�kg�%���V,V���<)�0w�j=X+M.����ҧT�2R���%�R�'%N����$�Or�B��x���OxB�
�m������IK�'}��`V�6|�|ًT�Õ'	8�PקC����	o�I=��I�<ѱ#�s0��R!`G�:f4b��4R#~�bM
��?���?���q�V�b���?���R`�dǬ#!d6�&���I�e!�,\#�q��H�R( s�V�6�#?	��ݔpܜ �ιo4,�+3�A M����A�#�0L�\���ǈ�-p��|�#��O87�ծ���8���Z��\���6�Z��I<���?��*��l×��17b�K�Dd���2�\���	�/"�
ͩ��V8p�X)��ʚ`����̦9 �4��d�!��l�P��J�$�8]�uFbS(3���M�8�@�ץ�O,���Ov��nI�C}~źe�Z�h�Bj
���eQ|&4�ƬB !ґdyEz�h��rAv)��Fި9M����O�+ �ة�擭E��5Z�bP=d�&� �gW�"=���V�(����M���	T8w�u���2 ��!c�L@��IRyV�b>�O|����5g&��f�LWdP���'��ƃv�J7EU�N�#���N^b�Q���*�Pj�4pi�TY���I��	t�b������o��pW������\¤p+�n��E� h��մ@(E�&L�# ���{�-�+L8B�n���O�kL=L,���AdƄid@<�4�rE]oڲ-��i!å�<IPջg�Ǡk�:��N����5��V"R9vuY�!V;(X�}�ӁC��MCT*G�,�I��M��߈���o�����cD�U�Bȉc		�~r�'7a}B��re$Q
f��"Iz�����O�~�|�gӰY�~
���u�A1Cq��C�Cv#̥���}>��O����+� 8  �   6   Ĵ���	��Z�Zvi��:+���3��H�ݴ���qe"���@"<A�iB���gC`�����Q�R�y��U�6��7�i�X�����f�TYؔ�.(�r��j�j�ቄ@2�Г�i��̩�+�>8Y�A�Ϭ\?�Y�.O����I_>7r�P�_��Rs.H=_��8�>�@��/H^.Mr��S��
�r㠞�?B�r��r�$�	�< �"{������
���[�$z���SF��F0��&�� �x3D��$oy�M��Li���R��8���4@x�'��Fx��Ba�I9Н�s�a�X�SE&,T��	69x�\��ቱ�PH���>��8[��P�<����ď��O��	�O��ҀK\lQ,��	x�N�i1�>��-tB�� ����^-:�0��I���!�a|���������O�H-�'!y� bf�T��jԋ�st�O����d����� a2�l���S.e�P�Е�	�ai�	9NF�$!7���(]n����@}ƴX��`��G/"�*��Z$�O�@s��;FT�kS����p��J�V�
!�<y��!ϬOF	�e���Y�I�(�n<b��OR�����Z��ē��D�,Nb�(jB�K��P��J�U��x��J�G�\Iml�D�9jE����'X ��j�-߃x�	j0��n�Q,O��p�O�{8�'@ \�gC����axr��S�P�k���U��C�P��s!C~�<CI>�'yQ�x B����W*W�~�.��"E-D�蓇�   �O���?1���d�O�Ȱp��'r�L���X��Ȑf5O���̈́�2e�4�j�~������`��-D4�c�b��\G�q�@��(�`T�I���	����x��yGeKT~���S��骡��X���O�A0�]��ڴ���y�]�Nhڅx�.�t&	��*��y��'M2�'���i��I�IRp����O�:y�4�I=b�J j!M�^��G�`y�O�r�'���'$�a�"G%��rlÔeNh���^U�ɤ�M���?����?)N~���r/�����ڷ��gĻF�LZ(�����O��d3��)Ò3���g���V hF ��ހ��#�~_�	>މ	�'��T'���'�ZMa�"��瘼CWvd����'t��'B����S�XٴS�x�Y	�̉%m�oz���@��8��!��*ۛV�D�t}B�'��I)LҡP�eP   �	  �  A  �   &  K.  �4  �:  )A  kG  O  aU  �[  �a  *h  kn  �t  �z  Ӂ   `� u�	����Zv)C�'ll\�0Kz+⟈mڃ	g��,Q}~�D�\Kv����0MX)���޺l(nIe�ڐi��q���)�(Yj�J�����/�T\���z�8ł��jHp�RíQ i��@�4������'��k�)/lm��� [ᦥ�׿��� ����D�`�	����N
�u���
J�<����E a�^)��V%�U[&L# ���޴zc����?����?y��2w����IJ%4ȘA���݊��? �ir`���W�,�am����ޟ�I#+	r�r$jV��TA5��(jA�I�8]�ԕ'c�"�=c�����D���%*��s �h'�ɋ=����L9D����_��
�a	3\8٠d�>�'J�O�a�Ū�ēd���^_�<<QFg�4S�I��Ɵ��ן��	џH��џ@�OS��]�8�:����_;��X��F�~����O����OH�F
�Vl�p�oڸ�M{�tQP�3�m۪2�B��P��؎�D��ȟ��B�+�I����,͜Q,�l c���TCz��D��-:�E����t��l�?MC[w��Q c�E�T��q�����@����25�)R�ӎ�C������;Q�ŋ5E:@�b냮R9��@o���Kٴ2כ���l��BbC�&z0�cr���h�@0���A�.�FMa"�r�(o���M'�F�
~�0ѥ��C6Ds�/I�M($<;s�ƾʄ�j�_�6�x�
ó;�|�po� ��43כv�u�E��@9`,��'��%^q���7�����Z�>#��4��	���K�U>�Ib#��?Gb.�Á H�?ʴ�3��]cp2�T�f���B"��V�<!3��]�NUa޴(I�F�u�t����G$�l'����O8��g)ߥs	��KCZr�<5h֯1D����L]:�d!�`�ˢ5�t��5D����푈[�6�qĬ	�&�hY�P�?D� �f^8�H���G�_�X!xT@)D�`�4�ɹg��y0�C�w�PA8��'D��H�%)nI�w�^	t'*�x'�%�h�,�E�4H[�`-̴	 ED
!��)4���yRmBpT;q"����:vD8�yr�]������G�	V �u�$�y��>;=p$�ӂD����
����y�G1J6���2!�*_�uz,]��y�D?[���E��,L7��iP��?I��Wg����l��se�����Ul�
�)xS�2D�� i��M��qA��5��	�_�!�d��^�
�0c� -����{{!�J�!�6N2 �2U���4s��5��Ig0��TN_:�v���/�Cf��	<������ ���_1<�H��'/Н��AH!��Ύc����Aǅ�� �ȓ⤸a��- �����ި*.jm�����#lC(p��=�U�S&a�`���:�Z�Cq�,��!v@�$o��h��r�4m��k�>F�~�ke(N�&~<����/\[��cݴ�?q�$�\�QU�O����'I�( l���?AB����?�����@�	}�%�����	
b�h�f��P:1
��čC�axȧ2@A�����d�?\p~�C�cߩB3�9���\0�ax���?��i�7��O��Ł�6r,*|
�,8�-�a�<�����(�Vp瘕,E^��V@[/�D%�T�'����:dp��� �?�6�؆i�.�B_����������Γ�y�h�,1��b�kϼh� �KSgJ���H�r�s�{��	��^��%@�[�9��d�0��.s��&R���s���q�1ѷ�@�j	ұ����!p���.���	ٟ8%?��|Z�Tx������
�q��(�Y������!@5���%(�	fqάk��G
f$֣?A��%�:��A'�9@��s"
�S��1l�Ɵl�'\uId�O�D3�ĮO��8��ބK���B��$ܐ$�'B�����Ϙ'�B��'��]��
'@%|͞D:oʑL��ɜ:�(�RQ�,�3�'_� �A`�gj���n�3L(��8?��͝��p�|�����I�`ah1�'�R+@MH'�qHb�ȓ��`��)��F02�C�z���'5�"=ͧ�?q+O�k2��kߤ��bmZ��@�����$;�OH����$>�:��E�����9��
�!��?´�Ic�\��y���҄L,���O��I#f�*IQ�݂�C�Q��@��@jO�ԫ��_�r2QE���/O��w"O��1v��[���*� �=?�R0�|2�e�|�OV}�S�d:/&���ָ� &�lTaxlJt�v�	5�	h�� �9��m[0���ˈ&vyT1+a�'��<$�C�e)�!�O@��RCΈhG��A*D)=bX}Y4�'sDD;��?����?�1�� 3v�!�C�Eۖ��%տ���O>㟢|���E�n�t��5�*�����}�� `�bzl�F��eJ�bP��>�b���vy��/"�6�<����H��}>ف��B�Q�% �� � Pc�O��$�:"�Y�C�9Xh���B�	���p�&5q`�N]߬�󁒟�qF ��]�4��t�O	��a6��9E�RY�
�S!�E��O.����'n��T��Ш]}PU�H�T)j�j�0
��'7��'a��c爼aZy�`L+ $�"���Qb�O�i@���W4^��cc�#a��c��K�򰣌��(O���v�_8��F(_&,��"O�!�'a�y��&��	
�5P�"OJL����@`J�Bŭ�z�~h�@"O )bG�Й�1�r�?��=��"O�cU��5�A��
 9I�PQٖ"O���©9�,U_|i@ i���Ę�j�|��x��H
D��@1�1���y҅00�6���+Y$o���$%���y�/YJ:~�` �����T�X-�y�i��ɪ�+�;��Dl���yR韊3�|���啈��)8��ҍ��>�dr?��D�w�b���A�����p�<��m�&���̎�n�D@*�NOj�<9(�<�8)���2	uHD�2c�<��d�e|�@�޷WB�0����a�<��@�/�R�BE�@>%K�t���^`�<1��Z4[�� �WEF�k蜂� �R�'�rUC��iýe�PY[AF�pM�.ܓ1!�D7�Z��+��"�&����]#!�Ї�-0TeP�����0'GQv!�$V�W���F�0p�Փ�^&P�!��ɼF�����(\$ػ$���!�Ϡ)?B$ʷ�KZ�͛a��̛�O?����Z�L��%���1#�Ժ�v�<�2�Ɣ:x��fZj!Z�d�r�<	�+�$xt}���wz��mDk�<q�K"�n@����:1:`�n�i�<���2ђ�1�J�+}�ЩP�@�[�<Q��%$]��3!+ &|UHEx���My"![�p>�m��	�t���[	 ��0P�ȝB�<��	IH�&�	Ք�PG%_B�<�`�S:d�
\k�Aڬ,� h賬�t�<��B�3�~e���a��qU�Z�<a�@�Z.������L���!/NLx��P����,���AT�0сG�9[���k#D�t�RK !x�
d�4��:�`6�;D����d_I�$�h�b�M̰xm:D��ar��%L�ز0����֓�yrd۳#$��3!J�W���Tkڷ�yb!��X�К�.�ְE�� �1�hO��3T���8�(r�O:)S\�Y��Z�X��C��('"\PP� <I��VJ�$X?�C�I-S�mB��C������X?$C��#'3���@��l$�[!+�*U�C䉀\�>M٣-�%��r�#�B�	�8;b��1`�.8���0�NPz��ęc��"~n�^}�Y�Ӈ霽�7�F\T!�dlW<���!�J���[^*x�!�$˵Nξi���P)!9��`	�5�!�䃩6u
�������0�$�K��!�K�Lzh���2
:ј0b��!�d����I��8��tb/%�剛:� ���V'[�P���Ѻp���`�R*~!�� �āg�	�bR�yC��ϻ�(�e"O�x)�év�~tA`fW�"���"O���V��i& �� ���#�:�"O"�󄬗&)!��a��A
 0MY��'�����'|�5���3L� a3��#�����'��a1k�UR��ŭL�	�2d��'x�TA�Θ	�5��&Ǫ����'g�93� �D��J����~��s�'���	�FUq=�IK�V�-��X�'!ֽ�A�WS�|�`jS����%o �~"�i�R��\!��jr��O�X�<yq$��<?��Raυ�-��QyAAZ�<	��C<G~��w�O�=f<�_�<I�G^�aNF�۵��z�J�P���b�<QW�� s�ʑ:�拜�,5Ȳ��g�<�([�!ކ�&��8<�'$���h��'�S�Oe��s���,z:^@bF�2٠ԫS"OzLqc��1�\x�GA�Q�0U�C"O�|�a ���	�+����b�"O:�Q��
h"f=��j�p�F�4"O}�&G:EE� +��1,��P"O.L{E�3�,���B�qŎ��@[�4H3�;�O��KeL���\@��&�*�8G"Ov!����x!4%B����nu^PC�"O��H)U� `�Q,&pb�/�!�@�7�r i7�ȶhtVM��:Y!�D��v}�ӢT1lv�I���#P�}�K^)�~�H�����.��f`H�����yB��ot"��=OP��l\�y2�˓X!4ZR��98���,ߦ�y�h_"_���j
)zi�+$AF2�y��
1f�6�-hmcuCǅ:��Є�X3���"*W;{��9[�NU�hD{R�	3Ĩ����e�ڄM�"r��K����"O�i3	%# ,=;�oG;��X��"O� ���5s���2��V�,��"O��ba⍦O%u6�ЏP��@"O,�ƃ<R�p=�$	n�x�*�"OZ���ž<��d��=n���T�'�0����p�}���Y�~X��D�KOl��ȓkB�6F��&����#�u��{�ѓ�b����&Ř�B�`͆ȓY�n5��^�8+H�@��K�b�^ �ȓI(д0snaŘ�PW���k�"���~p���@�0avX��
��Gw,Ȕ'<z$�
�7�B@JR+?`��+��$FT��ȓ+�H9�7��HЃ)�%I)01��=	8�SGm�2P�C��ǅc��=�ȓrh�DjB�5è�A�Iͼ�i�ȓ=����4R�SGJ�@Vh���
?���I�0�z��'�Q$ ��z� �(�B䉌D����k/Z��P�a �;�C�	X����LC�D�Fpx�'��!*B�	 M��lsׅƬb�t�%M@4j��C䉒$���x`�[�@ߐ��s
ܼzYB�Ɋg���+�n��D
~@G�
]�2�=1G�\�O�������)@
��UKR�om�Er�'�b����>R��
e�ׅ�P �'L>uiEnʶy\��A��3
�'|eH��ǉ8�J�Y�T�Y�Ah�'���  O4}��[7V�;����'?�1��l�T�;g��<�i
�o̴Fx��)Ī4+��{0i�o����$S��B�	�I�0��)L3	;�)k� ?4�B�)� �ųW#�?$�i�!��2"Obp��h�m�
�j �*3?B�"O���&�E Nst����3J-��g"O�z��N�~�,`NA)"+���DR���E�?�O<*�.��,,�%!"��?��ԁ�"OP�94���V�`��`/Z���Br"O��i�kW�c���"�nI)c�� ��"Oؕ)�FՎ~�N���gO� p|-�a"O���ŝ,^�d8��ra��/��}�IІ�~���8�����&U���{C�κ�y��}�L��� A�n�Qo�y��Q)	�l�G���>=¬�q��,�y2e�U���ōǏe�.tP�i]��y�e�2{���aܗ_�8�H�,�y�Ț�\Ъi�g��shM@Pg���hO��IQ�S� ��($O)%E ���(�!|C
B�	�d�(�bMG�n�(I���R�a+�C�I<4;�1dЩ���bO0!��C�I1}.! ��F
�bj��6j�C�I�]n���u$���a��;�C�I�ARD�C.�'�puK����Ԛ�Ě;A�"~J!Ձ<�|��!<aVf��C?�yR��K��$�����"h{DF��yb�S!}�r�3P������F��yr���
{�T	�oY4L��,��KU<�y�B�i�\=���H�BQys�N6�y2���aj7��%952ypc�J���DIi�|ᐊG����p)�5�LP3$I��y�
��/@9�0b�uY��"��y�FH�$��ȝ	hV�gX �y�΋% T<���m��M�2] ��Q%�y"
"+�8���7�� 7�J��>���s?�i�C!šP��F�Z=���]Z�<���,a�<-BEn�?D�qK�SA�<�'̀	gtH�3�.Ͷ%K�� M�@�<Q�-�yЦerƙ'{�4��vNWd�<I��p"X!����}�qhL�h�<����L�:$�UDW;*�}����M�'��Î�)�G�	��O^� |2DZ��!y!��0�
� '��� ����gE?-v!���p�,L�E�'@��	��nÌ{z!��s���mGo�~���BQ�2�!�ɵ�CU�ܖYp���E23�!�$�_ ��Bi�_:�1���y��Ϧ�O?}�p�J�`�P��^5O!����a�<Ѷ��3��7d<T�B!s�"�4�y�˴/'�1	ᢞ]��t�B+O��y�O�n��s�-�: ��$1����y�C���)q6��a
(�Q�y� Аs�Fy�uʇ���0d�)���`5�|BhӠc��U� C6(n��E��y��o�D��("1�XG��8�yŋk9���W�i�d��J� �yQ-^v��Cр�d�>)r�^%�y���6��� �e�<cQN�i� ���>�s��a?y��Т6d��9s,�����]]�<I�$�I�.=j�)�+&<�'��}�<��M�a��a�$��&oش�Q��z�<QS-L�Z��5��nH	EP��2kRa�<�G�V�M~|QB���z����f�D�<�e# �5���Ɔ[�;����}�'�$�����t���`@x��d
A˞�h:!��=��q�酥wq0$��	:R4!���X^8��L�sdTE	�!�!�� J[E�H�
^ 3E�] SV"O���'HX� aef�w��	h�*O*�p��%\0H0�,L�9��8�Ex��)�;7S����! 7��Y��k��B�	�b5�4�كfǨ�����5woHB�I:��BRC� �LuS�Z�3>B�ɿt�\��Ǧ�^����I B�	�Y�`�u�kA����n��C�	�hm0�����KW�C��@�F��˓P�Р�� J$���ρ/�M"��D��C�IX��Bd P�E<���Rh� E�C䉳��� ��W�b�`ș NS�s��C�I�4��-1�m�6|.b̢�+;@8�C��,T�����L�(�#qcU�r������=_�䌎�f�u�Dv܈���o��Lf!��T�x�4��Lm�9S�[�,�!�]�0<ܝ�� �M
� X�.T�!�d� �Yz���jL^}��@��]�!����s���(� ??'�D �����!����*p��w�����x�ў��A9�'
I��c�C�O��i�'Ǆb*b��U1�YU���
� ���=��' �A+�j��9�J\	%�V�-�6D�'�|ᰒ��K�1�N '��y�'�rt�P�UT1�Cğ%|h��'����̓8��Ek��F2�X�� "�uDx����A�<��!�A�|%�԰�@���B��%M��Ha���W���p�͊R��B�I�B@!r��U�?���1�˷-��B�	js䕳'KʥPU����Ȣ9@�C�I0Tv0i$(I�ر�4|j�C�I�'���Z�g�p�\����2)M��	R�d:}2�_�@�D:}��A	i��!��M��,DB�cN8J�֟���֟h��T��PP+˷;��ՠ��|"�DJ�H�\V��'a9.�����S�'tB��!�����7���r�Ӌ@�prB��P�YA��:j�>">A!��ȟ���F̧
����Q$ǐ����f� ��'a~RǔK-���b�J$>��z�(!��>�W���!��l�*�x�b��w��-:U�<�a��?����|R���?q�J�):�����@�98Y��A�?!�ׁKb8��c��Hpl�a������4�lKk�XR 	@�Y��i��:Ohe>��T���8�J�&��� �z��ԅݩD
�\S�nC�<1P�՟T�Iy~J~��O�q/M�H/�\�!�Ϋa�dE��"O�`��䄁^r>5i) �	�8 �s�	�ȟ��·	 �	�v%�$F.N����O�O0ʓ=�R����?����?Q+O��@�H�׍�2
�X���-���HWn�OX�2FV�%G�P�P�?#<Q���|O\+C!�=��2!�h���{zy��U�P���Oh�XU��G(�ÅI�*j��P��L���O0��4ړ�yR��Q��``��=�>0 i�y#۵�*=2��\0��h����?a��i>��	^y�#��H�m��x�C�DZ�����D5�"�'u��'��)擶:~<تCE_�4-K�+�d�~$I���U"�{P��+԰Xpϓ}{���\0 (�H�%ϒc�~`�ą,�F��5 � ϓ�F��	�7P`��J��a�G*a���Ij�'�����ׇ6lx��f2{A@�p0�8D����X�Y��h�3.
r�$��%G�<)U�iP�X�,ŭ)��O� ��Q�f.:����JD�`M�R���I����F���=�j �!��?�'R؋�<}&�P�%�7���D|r���L������ �xԜ���T>�ae�Вs�� m-�E�#!�6�,��͟��|�D�� # P�p�X�G����Yy��'a|�C˻B
���ր�05#,	�� ���>�T�ȳ�	ٷf/�ah��|�hI��<Qr��6=����w���|�T�O��*�'5G�T ��Y<Wv
u��۝�r��8�B}r�a\\�`m��	]�W?u�E)ִK���%P�'2�Sp�l��o��qܝ��#3�R��V�S�fߌ��Ѡ�	ւ�h@H0��	�~r�'��)��%?� �m��攏j�8���Ϣ�"��"O��+��$#� �`A)oE>bC��6�ȟTQ�U�\�T��Mep`E����O���O&�P�$R93}^���O��d�Ob@�;�?�,�Kݰ\P�&Yl,���-V�Z����'9L%�5�	/��KΟ��R��λSs��R�Y{m�ȉCƅ6S�0 �I�L��Ԥ�(,��g�'�k�ę^T�n#a�n�;M ?������L�'0�dU	5:��/��$��m��13!�I6>S��&&2���2F�=#ª/��|j��':�i���c�" 4dV7�f0b����Q����02Ijto��T�ޫG�C�I'!"x8��^*)̖ qw�$£"O�AXw�>4(�����YfBh�"OX��� �<uh��W��:N��!�"O�	�G�6>j���L ���I�6����C�')j�d����1���A��}hj�F|�y~=E�dE���A�cг~�Z���$ňO(<Z�G_*�(�8�����0\�ӳh�Ew�-+f�I�����O����K�%71�)�!oQ8/�����O���?�)�8�,�f�M��>P�S�@[}�i��$��	��PA�Ռ�1_%��%M�;
�ʓ�?��?��4��4y���
X�qq#�)�I9��(O��=Q���8|>|9�!�@0;�pB!Og��L(��%��~��1@t䲂#C* kVt�`o�H~r��P�`�=}*���D�XĨD0���C
�!n)A��N,?	��>Q#��X��RⓡS`L,���)#�ʙٱFM�41�2��>��O¢}Γ �Q��A�g5zH)Weӟ�B8R`�b��`���o�Ӽc*>���A^;#O�5bwOFAC��d����� G��)�7����ҰX� 0¦�� P��Y ��7��	OÜ�'xH6��+y��X�%S2J^��S���?��I�I���'��#�a��Y�<��҈��t�`���Ï3�dV�F��S��'M�9��O|����Ĺ|}"y� l	�NQR��@��-��I�����#}��i��8��L�Bb@uX�H:�N� ���On�ˢ����<�&�]?��H]�W���Qa��Mnm�̎��` �'�0A��-V4,C(|��F-l��y�'@\�aeƺGB4x��Pì�zݴ�?I�����O���|�-��9����Q��GZ�:i����Hh}B�|�U��G�d̖�K��U
�M`�`0�����ē�hO���	Z�)J�T$��V+{Dĩ#B"Oh��R�x�Hxz��B-D����"O��{G� 2\�T�u�1��`RR"OmZ2� Mڶ4��%۽OV�q�"O4�Yu*X,ЎܺC�\�2U��h�"O��EJ�;�x�g䑸4F$��"O�)x��JG�ɸ���A<�%ȑ"OJK�<9Cʌc��E	��h"O����@	f���6A�W�
w"O�E3�G�>Cw�+�oÌ���S"Ox��P�VOL�%2%�P�qw��[�"OH8At�r��8:�ǟ�=fLՃ���){tމHȋ�	��	te�Ro���f��*��(sa(�/6����!l���s��9�ʨ�#NL��~�	&!�I��.�5�,$��k
�&u0�B�#5�L@�.�,C�`T飭��8s#(�2�����E�0�b�a"�� �@4��O�r���� ��A�I�PP�c�B����W��(p B�ɭ/x�����/"��*a�f�B䉉~N-��HA�\~` �T� X�B�f}�m[�d*ny:�C@4K$�C�I�u�Jy�$Z�48��[�� �~�B�	9z�ڤCF/�{����H]2�B�?kļ���F#8�X��_�@��C䉳`X���Ɨ4c����`&j�C�I�rSV!��аo��	�.ҮC�I*������:$ZՈ܈t�C��5@A���{���@-ۺC䉳&����f�2l�EG
�8�RB��*	U��!�Z�/���J�½\�B�)� ��:g��/n���{��/�Z�"O�<0i܁jw��Z��"jZ�e�"O�q ��n�� r�=8G� k�"Oxe1���]�M�!iۚQ�|�V"O����b9+�"԰ŧ٠4��f"O��a��O�C���gE�*H��["O
E!"'5�� {��?O@a��"O �����1T����F5=R����"O����.���v���?�u9$"Or�p�E�L�иZ��,���"O^���ON�HR�8 j��$D��p�"OJ�`��/&f�$�U��%'@(Y�"O<-���6�rI�Q��97G���"O���0����%�!jȋe����"O���҆�g0�]��1o�&��6"O��vEB�1�P8��6ޤ�j�"Opйp��D�b�@S��	i��`�"Ot83&ʊi�-X�.�pZx���"OZ-�R!�V3���mKN6i"O�ă!�L:pC�તm��G*�e"O��2`�P��s��+>�M�"O� aB+�[���["̓t�v �U"O��T���h�H��-W�R��t"Oha�&$J�!�報L��]����U"O2p���͢IJ��n��3�X���"Ov���ƁZ���Ä��z�"O D��C�����xd��6�� �A"Oa@�>����7TM&�`G"OP虷ɞ�d�u���%I���6"O,�۴�([5UI� T�"E �ن"O�I�V`��q�������q;��"O�`IZ
V�2Y�C9eG��0u"O`�I
��vTHR�YU���E"O�Z�H�T�)D��
6���"O�K�
Y&>��)���~"TQA�"O(e�p�V�Mf�+_�����۽�yB�/J�0��$�&��kP�R��y�✅q��KdB�iߴ��r&~q�ȓ��e�!.��oh���5F F���`i)��. �t�!�ƌ>Q�ȓ[�ڄ��]#Et`�[�
PӴh�ȓ���HG�I����5��U���f��Ȼe�j����2a!�a��P���
n�=Z�d���������Q�* �Uz1�O�o����Gg��fۣn����GȈF$�؇�fa�T�ņN�N{��F�үCo8͇�E��d%�
H���@6��,"�:���@2�8��Fg:dX��[�-hy�ȓI
.h��~�J���E�T�)�ȓzl0��FH�;y(��`�O� 	M0y��8�P#��������^�Si%D�<�@oA�+&��ص�<Pz
�x��5D�\+�o@65&���ȟT$� �D4D��a'gՔi䑃T�^�q���HC2D�cA�C5#Jδh a=�t�E�1D�4bn�'�PA�q�L%, ~��b�-D�|JG�J lz��U�=]�8��/,D��yv�/l�� iI�gX�$ %F,D� b�QM�V�a��Ȝ�l*D��R�E�85�����?Bv(��(D���cD67�D��$^�?�L���'D������Y$8�Э݌j"FQ!K)D��'�ѕO��1Y��Z�m�T���(D�� �	����(�����ڛ{�L��@"O ��$_f��$1����^���"O��S�nȫF*������k�6ٸ`"O�As�H1���"���}���"O|��J=��q0�ȘF�>�S!"O��b',��8P���qk���>P�u"O�DabM�2,�4�!$ʝ5O�x�"Ob���mӏ5�T��L� ��$
�"OBu3R�����p-0~���G"O^y;Ń��C��ԧZ�ΰ�Q"O�0!�a�'3��)�b�J�d�:���"O�0J",�^\�Q�ѵ�\�r�"O&�Ʉ"��4Ի�*�*���k�"Oj�Ғ�O�&�����4+��,9"O"0��H܂Sؼ�P1&�(���"O^�q0GL� �
h��ʍ�~�b$u"O��1�z������s�X1	!"O~͛VjW%P|��$��5�`��"OV0�!�a� �b� "U�1"O�e�"̐)�j�p �!n�L�C"O���s��CS��A����d|�D!�"OT�@R&Sp�Afn�	t�(`�"O0P�m��a=�;��O�5�Y�"O8L�4���T�e��ލn �8��"Oh�R�Ɔ�.]p�3���g"O��q��خT<Ay�:C>�� "OF�����"<萐��^s!�*E"O<����7]�� {�IF�~�Ys�"O���4+��/���%�L�?�xp:"O�Y���f���Q	 P�$z"O�yq�e��B�<�r�M�:��e��"O�X(MK�Mn ����G�� 1"O�������EЎ�q��tYw"O<�y�E�Z��iH1S�CȄ��"O�m�����~4l����3�V��c"Oz���$LL�k�^U�$Q{�"Ot��Q�N��Y�3nE6*8����"Ó�m�?, (�!��>+)��g�<a�J�
W�P�c�Oyt���y�<�o����8Y �ır}��1V�]u�<�%���[(m�,Ħ1D5��w�<��A�G�Xܻ��O�J��ES�� t�<ab�ߓӨ(b� ����t�<a'F��ҬPÀԙ<�n k��s�<Q惒��%B]'4��)jÇ�)@�C�I1E��� ��V�[@��� �׮C�	�kJU;��۝8��(��ћ(*�C�	�hq�]Y��Z~�@	3@�+:{RC�IG�t:4�L�F�����+	PC�I7�\I�����ea���>@XC䉡6l�@��N֐�ڂ��C�fC�	�|����6}��#@���QC�I#g}.�I����l��X`�� �B�%8�2�rA�G��ѱa��iN�B�l��!�q���j��]�����l� B�I��4�CG�tA�f�W��&C�/J?BYQWc�,U��RAۉ{"C�ɢ �4�S�%U�H�
��E
O��C��	�V��g��*^@<M�%��1��C��>�x��̑Y�2�E�*f��C�I-d=V�!&��M�w�P�n;D�|�SϜ�zf���+�0~���Pb(;D�X���ԁT�`(�e���U�$%.D�,��&C�U�N�;%�7MJ�D#.D�� JI��C��� y�i=(�`�`"Ot	�1ܾ1��l�fȥD����""O�y�����4ۢ	�����R�Zآs"OD�k�*@+n՛�eF�S�j	[d"O2b`(�8;�|���G�f���"OBy	�rH=s��v�©	c"O$�t��)� ���X4sJ�y�"O��B��XR?��	Ī�PRb8+�"O�|�#I�H�p��؆��P�<�#G�K�xbCm�i4�� �kP�<r��
uɖ�(�oT�@��p��N�<16I])������D,�Dt���<Bd��Mj慇 	�,��&��Q�<���o"�7(٦%5<T��H�V�<�%�� ��0H�ˑ&|+D��b)JT�<Q�M�N��R!�V]�fl��VT�<�]��R�N�|S���n�5Y�!��4�(� �Lx<�<�CM�+��$Ϙ!�H�
f�ȹa|�Ѧ剁�y�盍���!F�R�r�l{7��y� �~�����m�)��-8�y"�[�Aͪcb��iZ`x�nB�y�j�%o�U֙u���#K���y"&�0"�T�&'r�6�J3�#�yR�Z0�3'���K~�rcƏ�y��_�@I�5Qu��?\N����Ĺ�y�_6/\�J�EF�W
��SR�ղ�y��6`�J�8d �H�BY��y��i��ḁf��?�n��I���y��ѠN,7�e�:|�@�ܖ�y��,3�Nx�T�b�����$	�yR�� W�	Q�Ŝ�] |8s��y���u<��+��Qp��C����y��N-+]��r�σE���
Rl�;�yB�I/h��4�[%if����y2
	z����t��bp��aE�Ԙ�yB��_֝���K�X/�|��KD�y���B���p�O�U�8� �퐅�y� A$r\ki�6��P�b��yr�O8}��@Ғ����Z-�a �+�y���R�� A��/Ҵ��'�������HH�d�V���1�'�2H(�mW25�l�6!T�ֹx�'��9w�l��EjF #J`ȝ�
�'�D���n��6��孕�Ee�@�	�'���aFܥ��0�5FI-p��	�'�:����M��$����W����'�j}�GN� \��@a�����'
�p'���'c���K�+ָm��'�l��,�	vf��S�B�2��8:�'�`@��ht �#Fފ-F� �'�,̃��N�m�  32����X�
�'��a&�,.�ڱ�ڮ+>�
�'&�T҇���&l�{�K��8��
�'g���ş|�}x�ꌤ?��3	�'�H����Ԛ[P�rwa�	)D�	�'!��cGd.n�U�GIθzը�3�{"cT�Jj��+�pppѨB.��v[ ��#�0~BH��O&)|<��,T�Љ�]=��Vd��8�݄�G����#��b0�=��/[z�d��N�B�"�¨=O��1aiJ�i����ȓzXڀJv F[�hIa=ց��Y�fi��
7&���lV��T$��Mqȩi��ێK�D�é�
\�(��S�? 0GC��Ѻ�S�i-d�"O�M��#B)��q1�͙�16��"O�h��U��P�
M"}mI�"Oe#H�e�-�p���;b��"Ox ㊑�sߖE;��nt��V"OX&���t@Y
��D��"O܂B� W�h ���O�k�zI1T"O��21nB�G�C���8�d\�"O�m��M��E̔�"��5���d"O� :V"����2V��]��M��"O����؆}r�ZA�\)`��yc!�d�:ٚV��c�uRs��vS!�d�4f�`i�4�ݑV����N��R!�E�hy�X`�#E��L����͍wL!�dSC��H�c$a�p�t��D!��י;o�		����T�9@�Nc�!�şg��:�^�9`"y�$ {�!�$�����Ԡ�)-B�1�5�T�_!�DV�F���k��90�
X8㊃�VX!��%/�L�Sâ���`ȺШ�B!�Ĵxt��։Qv/��.�0A!�$�2�DE(#eФB������!�D��+ʹ#',9v b��K�g`!��h�6���DXnI�c]�_V!�D̗h+�l�0	�>K+�{gB#�!�d�V'�$��e� w=* ��*
/89!�d�{�B�ѣ��>v#h䂧�ڝ
!�õAx�ɶ(B /#��!��"O�iJ��;L ВcCN�H�~}!W"O�h;��E�hs���Qb�//���J�"O��`Q��KGb� 灀(?���+#"O�[���r�%�p���B�`��G"O4Q�	Į�&�K����U �"O��a��3��	���fΒui�"OL���ѵ@+�!�!�M�'��l�"O�!9���N4	�G�7�
��R"OdayIB.E<az��I^R�RG"OAK��C�;wp���� ;A��p�"Od�Z�:��m�����6�ޜ��"O��3�Y�L���zu��/:�,A�"O��"�@�AF�:���%}�`E�d"O����KΖu;^�۰gP[�pIP�"O��3e�º>���j�/�0,��H�"O>8� ��2�6��!Qx��p�"O��g�I�#��P:,��a"O�E�R�_�tU��T�LQ��< "OJ�aA%��1 H2(�'/���5"O�T�O.�t��'(�_�hi��"OB��1�t)��Oϭ/��T��"O�HeOG6� ��M���@�k�"O�y�r*C,q	��¶U�_�Z�Za"O��@R���Wf��C�
�$Qb$B�"O�țAb��yߊ�p���C�U�4"O؅:#�
N�>H���A"-�"O`4H�J_�X.�)P��Z�����"O��1�8gT�Yɗ,܂8Т�"O�S7 ��� 9�m%*w�3"O���DƚN��q�l��,�p��"O�I"�A���L݈�cמ����6"O�8�q�Y���b&�M�s���"Oz��&+5��+�AP:H�yw"Od�Y���6%JH�G��P��TA�"O��&���f�N�R��J�n�bI�"OJ����Δk�*=c�Eּ<`st"O� ^�X�M�/��9y�KX|Tɰ"O�X�dR�:R��2V��6}U�*�"OZ�zGC��'ۂ\�A�W=(C�@�P"O�p;VÂ���� �͉G@�T�"O��(�V���z#��.�z�a�"O���ӧÝK�xd���9���!"Ot��d�-w8f�ŀ�!"���/�yҫa
� ��jQ{���o�y"�Q� \xZ�b�.EC��B��/�y���>Et�2B�H{�����!�y�(L,	g=��o'v�'f�y�c	�RFiR�۩f�ؐ"S�Q�y® "@��@8!E9��S�mA2�y�`U%NX<s@�O>R���
�y���f�j�R��93� ��'R��ybc s�V4��BX;~�*阴�	��y�,^n��$Z� P4���y�֊4�v�:�C�� !�)·�yb�Ƶk(2�{�зw������ybm�2{�A�S�."����W�ʌ�yr%R!4-�#�/7]�De�sę��yOɅ@��T���C�Je�;�G�y"HBi�Ҥ
L�D�p:��T��y�'U�1C���>�6�&���y2� �0�\��Պبq�xi�A���yb�I�<�X�+sb*g������y���},�hx"�N��%eK�!Z��eWHT�eR�e�h	�B�OkBȄȓ
*~�p&��9FB�bt,�V����ȓ*����Si�"딕����^̆<��/9����a��@���i�f��N> ��McD�K'17~XsdV�љ�'GU�<��i@H!���)(�x$�Wz8�P"��Ұ*���*y>����3F�!��(Jj���@zЭs�M��I#� 7m��/��������#~
u��Uw�e3��FP40�Z��s�<���L$��em�3P5ڜ8E�
��̕Cv�M��0Q�ݩSĨ�&?�4�E�@�Ng���!EJ�vJ�*w�2�O�\h�!R���	Q�F"S�XͨG�!D��#�M�PEn%01�Ŭ��=i1��'@U�$��+%�Xq���Xz�'���:�J=^(K�GҴ�S98�vi�R��y�Zq`1���C�	(+f���
E+h��p*��n���ɍW�P)XE�����t�B�U3r�D�DCe��SV�L���H�.���y2/!gV@��J��	(��z�$M���k �SIk�HQ
&�O�OR|�T	G�E��Z ���",�Ń��'q`�I�BA	��g�mM�����=�b��X ;�`��Ҭ;P�a{�nߖ>ʸh��أ�x|:V����O�l맄�6+a�<h��ׇ#5�m��foݝ�g��¹c��	F���G�*D����̚v�~�h�*
>����#b������U����@�>Q�|x�rn][�O�ԉi$��\<B�Z�&h�Z���'��s�F����[6�1Y�ⅲ�h�W�h��4�	�%S��a$N��g�7�J��4���	t�8s�1O������1�Ɣ�CnΆ*����Ҋ�P�����Wd�m��i-x�
�'9������3j2���l�H�I���ʶ&vΩ��Β��4"�.e>�(�l b,� �d�%����Ѥ4D��x� ��t���'ڬM4l��&��<с�N�(36в�b���<��^�m=�d�dEA�Ϧ8H�S�!�DV^v��8�D�.'� ��4㉁Cmd��a�>q�a�3C��>�O*q0a.[�V�f���7:RD�a�
O8�2�
�} ��I��S4&�����h�+��q��
��0?��f<�F_�\�pB1�CJx��NO�xq�'��Z��N'Jݜ�+F%��J�"��	�'�n٪A�Y�<6��r��r��x	�{�N���O�O8�1��dR�Cɼ��B`ٱc���Q��� L��G���	�Fp��eV�n,�"O�I�Fmߪ0��`�LT�BQ��"O��v)��m��M��A������"On�×���9X�ࣁ(��,B�"O ��$ވ�๻'Á&����Q"Op!L[.Y0e5A�Z���PF"Oള�"6L[�;���6l�)�"O2�Av+ʫ\�bB���J�\	�`"O�[%�\(rVBͺ�B���P��"O*�p!�Z
C���&����T34"O2�pT+Z.��% �n>t+Jy�B"O@H���۱UH��MH�9�T�"O�� (g�
p#F-dyt��"O��)�B]�>����"zr4=�V"ORa�#c�_���T�G=���p1"O~��U�4l��s��*B���K�"O����(��ղ��f�*䣔"Oj��@�^��[���N�ԅ 3"OtM�u��c��1��Ǟ	���T"O4r%o�U�T�AƜ ���!"OD`b4�¸4rF)����V���*O�l�%��;�n�`�-�e�vq�'ᒼC@	4����E쌳i_j͹	�'9���G:/�u/ڈ4G8�J	�'��(I��_\���i,&�r�']r���U�i�D��L������'�bp)�1\�< �h�����'I��)SKO�<�T���4��pJ�'z޽���M�$Z ���˒y@.�j�'+���
�9r�*p9c��q�
K�'4�!�ǵ$�D���Z$v���r�'���в�)��T�+ݐCpj���'�&mJ���#X��1� ţB�<0��'�h��ڴG�E��lˏ��S
�'�aB�E�TԼ���D�Z%��'�aF�>?��X`C��@�y�'��(%�5o�L:�b^>y��5�
�'��Ř'�h�ܰ����r;ڸ��'��P�C�V�'�޸��)cw���'�	���8�ѫ���'��M��')��:0C.o�Ι���Z�w�Zi��'��@�ʒq�0�s5&[�=�� �'���1���@���g���0~��
�'���T(ȫz��S�l��GǺ�
�';�$�B��;�N��j����
�'?ؔ�)�!j�HB���8�i
�'	�V��<�|$R�*�!���9D�� �� ��	Z.6�-���9D����p�&9"�Nܩ.��1�G9D�d������7)Z��pl���8D�<���<RE�����
M��@2D�x�@A�5B�zQ��	=����:D��"��\�x��af�3<p�(<D�@��W��%�R�K2�8i���8D�\�e�P�H��[�	M�^IIQ�'D��2�hA-Fサ:Т�*\�:Y�"@2D��@��,b�9�'%�57n��e0D�ȉ`�39)6u��!�-b�};6$"D��� �47�ipa&ͽe"p���(.D�tِ�Y�-�����O�k
 �z�B+D�X��\�3��D����EB�(�I@��!��
���Ԅ�0M@�ODx�#�5b@�uG��<v����"Oj�x��ѴaQb�˄��A�"O��@�O 5���V*�D\T"O� x0� ��<L4��k�^����u"O��	��[�%��L�n����"O��b�e�yZ����a�-ꮨ�%"O�a+5.b��AQ���-*T�L��D¨@uZE�&��]~N�YA�)D���/O8~�D5ؐ���A�(L �'&D���ҩ^2��"����	���$D�!EN ;a�9@@oBUB�!8N-D�(c�ں$M"����E�4�FPz�� D�ܘ�˙�3��yz���x�H=���>D��B �Z({̵I�aU/F��TՅ D�D���^�/H��abe�'n�р<D�`+C�$R�k7�R1��@���<D���P	օ�@1x7� �j��:D�d��E��2iN���	��a�%O&D�t���I^^u��ט]�XA�%D�(Tg� �bd�Z'>cz$���(D��R�KJ�1����#ث6���pC�(D�@��B	��z�̨���ϓ��y2��T�JA���Je�9HG�y	N�+�,�R��!Y:��V���y2��Ut\)�s�֑R\9lƧ�y��ŲoW�p���G��ɲ����yB'�?_\T`!��C�V���=�ȓH�p]J���uA�č'����EFU�!�F�5��X�͎7�Z��ȓQ2i�7�`庵HA`�,��Q�h<�FU������sYF��M���pR1s�& HP������ȓ#B�U@d�ДP�na�ƨԃ%z�Ȅȓ0DT���߆Kq��#-
�\L��ȓ4)"�
��H��G"�Q>F-�ȓ]�1����=t��N��6��(�����X�����bf�B|���_0xp$�5�P�ajA�`�ȓ���w��!e� 3d�/ �}�ȓkW��Kn�bpР�u �1۠���;�0���CZT`�R��	�����	���ٳe�j~�e`&���)�b��ȓ��ч��K����G+CI����܎\��jQ=M�Ό$^(X�@�ȓ �
����^WLa���Ѥ�jQ��'A���S�oP�����
J��ȓg9P�@kS9�ZA�w)N�M�i�ȓ!�Ƥ�M)���Qh�}�T���o�D\qp��,{� ��EÀF�x��ȓ<9*g''yԐ�;Үֽ|�FфȓS��a�AQ�3�e���2}���a}���ቔ_�P����03
���f92�;dn@�nZ��yp�Z)���y":���K�I�	���j	��?�̼PDGI� ɎxA��#��܅ȓk9z��i��\.$qg��T�d���B�`H�埛&	�	a@	T�����^M郧�mu:}��E�a�"��ȓE�`�1F m�RDce̝	!�Ї�Q� B&���2�2��d,�>%<VT��b�x�SV�T�-pP�j�'ۼg���8�$�2�Α� ����\�	����aӰ�D�B����#Ph_��ȓ��`�J�,͖�B3�³~^d��q�r�hd��Wu�l:�Q!��m��\�#��B@ '00����tȊ��?
�c��,>���S�? x���!�=����F4�""O4�IR��R��"���c!�a"O�!rBb�,=*������c�c�"O^<C�M]���hP@,~^��S"O=*u%�"h4$���Ku((��"Oj��'�_���сȐ�u\v"O�3����!<�
W�gn.���"O
�B�4d���"�T�Wg6���"OLq��c�(Q�<�C	]#Lbī"O����� K�Գ��ʟc3@�0�"O4��cJ�1�dx�p��\��\RT"O�ᴫϙ{�p#Q��p�p��"O�5Ѷ*��{�\x��bHĸ5"O|��S��U�\���"]�X�p"Oܘ8d@��e��"�d��^Xlh�"OL(�b"�w@�����kO�i�"O���S��&A]�|u��m3bɅ��y��Y
+O ��M�6�<�&����yb�v�tu��@Z>Y36l�(�yB��# �4�)gjC-X��B�)���ybOZ?
�DLj���g���n/�y�BǙF6���;
�fY ���y�DQ;_ʝ0sl$	j�({�S��yroɎ;����@�V�*����?�y�/ �M�YC#/ �V�i���y��XNc�!���,���eH��yRϞ9c��l�4L
|iVɘ�j���y"�E�.`����<�P�3
տ�yR��
,g��kpG D�$�7K���y�$Ӟ`9�	x�9H�ږ����yrl�;�l��%	Z#-ʦ��E�O)�yB
��芤��[�p�ԣ

�y�������@j|M:�K�)�y�O`�ހXq 06��uq�矧�y"
s�[r��4x�X
C���y�E�<���qo��d�V�&[`C䉔tAx%qV�@>a:��iUI� @B�	+wz�	�	^�-��z6IǆE��B�I��Bh�!��U>��VC�/B�	�J����60�4+���y��C�	�=���r/����
矴H��C�I/O��<1��>�ȕ"t�\/_�tB�1�x0F%S>Vb q��YaH�C��1��A��,�hL��G��o�jC�ɓG����a��!B	tiQ�ȻL�B�&tgr���'M�x!61h��B�u�C�I31�иE��T.����^�74�C��dg�p�%OC�|�>%"���*��C�'yJ���G�*N(��Wm�$~p�B䉥2��Ѓ���<�)Zqw4HB�ɣ �8�&�W6R}�:�O٣��C䉍�(@@�I�c�lY�M��B��@U=I�L�xb3��><B�IXŐكԃ�"B8�Uɕ痬(�B䉔�\�%.SI��G�A0v�zB䉣@�.=�P�w��2�J߯j2C�	ej`e`�KA;,Ű`�3�^�|h0C�I�Hu��R �8�)�s�܇�4�?Y��IZ��D�۽�urR'��!�!�$���UsËY�|<�E��~}!�dɹf}V�ڑ�U��.d�g	5{}!�䜶Q#v�(@����yS���p�!�D��A���[�7,��ue�4_�!�	=N4����o_�f ��D�ړ'�!�� t�1�/��>A�$�$�Z.x<e��"O�HC`��L$�'�C�b��S�"O�8[��n����#�F�%����P"Od=��E�6��`���q����"O������p�r�!Sʓ$�0��"O ��@�S\��az�'T<�&"O:!�-���YQX�c�KN"�yr�s�

���;�}�����!D�<3u�j)��s��
;��EǤ#D��Xu�)D<>Tp1�̔K�ųģ'D�(�7E݀A��iR�*;43��Y��'D���r"�=[�	HB�s�`�P('D��I@�
�M���De�b�yrK#D��a"BQ���g��0E�?D�0��&�1A�m`D��$�y�E�.QT����w��w� �y���]YB�(߃m���`����y­-(��K�g �bx�$�._��y"+-~��-
ц�D�l�AӶ�y�%�����JG�OF$���yOX�B4b�ʸI-�Q��ybL+x��Ap���1<�<� ���y��T5B�d[ץ�:30��0�G#�y2aőv���x��»'����w�Ȭ�y�-ѷ���!�Lvx�p�I��y����&tPRNZ|@\)b�C�2�yb�SX�,i�E�8bhp%2A	E�y2E;d�vQE�F�
��`��>�y�	�[Y^���ލ�j��C���y�m��Gx�\�VcG
?j������y�CU����H1�%X�̘�2&���y2NҊ{���ڱ,Tz��ԙb�E�y�&)Mp��`�s�F��0EG8�y�A��[� p��$��	7Ѩ�y��=w����Un���sAU��yr�6 �͢��ӝ@�}�P��y¤�sw�d��f�	<�<R�c���y2N֌M����׮۝8k<�W�ˆ�y��ȷ��U��Nϳ0��������y"%�7���A�)E�M�wş4�y��N�D��)�%�H���M��y�"�x$#��ޜ�A���y�C��t� `��U���h!�Iȸ�y��'B�y�wĞ�w��)�դO"�y2��
�s�hT q`e��*X��yB'��8�#��n`hب􀎒�y��Y)8r�ȃ��T/ݪ�Z��y�CI��p���
F�}�̘�'X�yL�-6(h9PD�{�TI22DL�y�	?}!��A���g���1��yRG�O�Rd!qL+af�y�LN
d,̘��H,l"`����-�ybi_0��@���ə��}x�&��yr��c�)R�n�5/ؔ���l�/�y�
��Q������>,˖9��o���y��V�&�4�3��� 2kd|���X��y�e�� ��=Ro�.Ez`�o��y�ⓠ_�n��g%X U�@4����y���5Xtp`���Z1q�#(�yji���t����8��-��yҬ��2���BW&�3��y�b,���y�vvtt�{ !��K�y2#\��ţU�k7Ve��O��y򅙘4= hI�L�!7ڢ!��+�y
� ��#ԍ�S���&�!=���"O.�1R���֍s��d&py��"O.�@cF��]�jQ��K0b�Y� "O��q�m�1$嘄��j
�B%�dз"OZ���-�\�`5 Y.1�Y�Q"O|�{"&B�j̍�/X5��"O�[�������N��i���Z�"OBȪ4�Z I�����̏X�B���"O�8�!�4�H `o7\��qt"O8� �F�+&xQإ�]�Mk0��B"O�,�QƎW ��K�K\����"O�a GZ@�1�bkP�s��u�s"O�G�һ{J� !WEQ?�>�I1"Of�j���;N�4#���Y�!�"O�kT�\wl)+BA��%o�P�U"O�Y�U�'xƼI@�O3T� "O$��%b�:` �@��Ң~`�i��"O�H��یZ(]PfP]���"O^`0����,W� 9qd�@�<���>x"- CѶ�r��y�<AC��=a+��K;c���;*u�<	�$Ą���Y �D2~ Z�;WlBm�<��H�Fs��CFD�O�N5�͒j�<�WJPLt@l���ZF�ES��\�<��ŋ1
� �Qd/�$�7�PC�<��Y(Y���m� �����H�<yv�"8WB݂aaվB��4�E�G�<�C*
R�vc2�	�A�-��g[�<y���6�I����TݐR�k�<Y���� %`OB���q&Fk�<	R�1�P䙶i�4h��=�/�Pybn"1�6��c��
?� ���Kc�<!������w�Ceh8����Rt�<��Y	a���D�#��)s�s�<�%gS�����L �8ϼ��`�o�<��&J3���&	4a'����_j�<acg�6��@"���0^r����Nk�<�3�[!�Pd��
�/h�2��vm�}�<���O���@g�/@��A1�L}�<!6*�707�PH�A�:���w�<Y�b�m�F�i��]�E\)b� �Z�<YC/�K:�����%@
u8f+O�<�3�Z�G�4(��?������N�<��*T5� ���E9#�����[N�<�4�­M�.�9��E5y��Ii��RL�<A֎�Po~�.GѤu���KR�<��I���1�u���I�ʝ��`�L�<!2�"erY��c�e:R�b�F�<qQ�]u\8�4P�\
��X��@�<��-!b5L����3\s�� �b�<a�C�D�T<��0|� ��2(Ja�<�d�FPz�y`��i����kZ^�<� �T�yzb!*��^C6�/�X�<�cE�/90�q��l��e�"C�[�<IK	�\��Dx��ȻG��Y���\V�<#��=M�dS�H�����k�y�<Q�$L��l����Եu�Lp�/^�<A��O�MH��2@^�1R�Y�<���6����k���|�Z%X�<iao�A����Eo+DRZT�#��y�<��h��'� ����'X�6Ѐ�"�s�<���O/�2Y���]9C�n%�*�k�<�t��&�JsA�/b("3�e�<yvL���E۳�_"U�L�q�IG�<� *l����$vd���aG�*=����"Oj�+#��+C�R��V�׸�{D"OP+�i�>'.�AEQӀ��5"O�q"��k`���l�|�G"OV��Ζ2C�����-�'¼S�"O0�i7�T2N|��Z3MߘC�V�F"O�8��M�:RpPrbX9\��(x�"Oޝ(�N�GQ\���KČF��r"Oh�CK���T�,
4��h2g"O�xWf1��Iv��u�X%�c"O,=1W�M��4rFK&�X�8f"OD�CD8� ǭƽ�� ��"O&�D�&mO���mW&w�R1(�"O��Ak�dH 	cK�d�4a�v"O<���X�o�E�`�	�>�fTq�"O
���B� ���G͎7r\��"Oj]�� M����GI>-]lt�"OI��@�3fU+���)�JI�"O����		�o��VC��l)Hw"O�a�,	|�c��	�u��Ź"O�EJ��x�*�[$���n���E"O�豦��< ����K�e>�˲"O��)���q��`�!�{  ��5"O<Q8�c_�@lkU�.1��aW"OhD�jn�`��K:N ��"O>5�#��>p,��;,�(ra"O�(E#��F�x��C���`3�ݺ�"O�h0D���&�@١���O��3"O2��C�B,x��7P����"O*њ�m_��"����՚%�81�"O΅yD��]
�f#��a�"O���)0w�و2�9g���3�"O����(��4��*UC�e�0� 5"O�i�p�EtG�:0�;",��&"O"��tbZ1VK�D�TBM���q"O�x��m.�5�r(D�8u0�"OJ��bQ8d��Q d��3R��E"O�}�Ӌ�R*rd1�0.�q�"OR�R6J^��P�܍��if"O^bw����"So �#��@�*O�(�6�ݪ1����鼍	.!��+l�@S3ɒ�S�FaEI]�-^!�D�Yd��"M�3I<A��(�	V!�T't�
0f�J�Z0T=*3�GX=!��A=i HlS�IJ�! D�З��&L!�QN��ۥ�����T�S*�Py� �
��\��A	&}�8Ё�I���y��R�|Lj����,uw��N�<�y�c�,e�$�^� �8�ג�y�;0����%oӯ"&�8��V��y"B_]�Q����:��%C]�y�Ƕ`Z�Y�*
�42%���A4�yX�r���Z�&� u��8qhK)�y��)D}/�q�������y2�ӣy)�ũR�`y�u��ߕ�y�嘥Hm�Õ�պDL��PхA*�y�.
^z�0AH��*�JQ����y2�	Nv�@ӢÚ5l|\�&j��y�m�&�JXz���8��P�F���ybeL�T
�"�Bb�����y���*+� � ?�Bᩔc��yCY�;�I��ؐP����/H��yR-�?0��-���2� �{�%��yr%ѶM�n1k�뉸R;��z���y
�  �
B��*>鶉X� *;�����"O؈*3�!b�ba��i�.Y��8��"O.��0-��F���r��Ѵ
�:��"O��)Ԥ�.`��ƅ]�)�ͣ�"O�i�g�ݦD�n�b$C�!A��|Q�"Of! lE$Oz�� ��Ϡ��B"OR<���E�b��s¢߸"ɖ0 a"O�����!��ۓ��3y���"O|���C5T�d� ����w"O�A#$�U��*%�V	F�<�*�"O�������Urަ��D"O �:�]8CV��lD�5��!�r"OY��B%d�
��T���Kg"O��s1���d/[:��TR"O6��������DP�L�DԂ�"OH�
�֞9��vDI1i�<�i�"O���3��/[��む$36�"OIy����u�=�Q��y�l�b&"O�� 7�ȁGT90���|��"@"OZmD����` ����'I�b�ۓ"O���Cb�Wk �I��k���S"O*�+��<^�p �H����a�"O����M�L.�fǆ���'"OJ�aEa�"p>�X�c�[�|��g"O�i�,τg74�)#P&��<1"O�}���ȱ��E7�(��]Qt"O�P�C�rQ��]�D�h��#"O\@J�O�;B(���� rJ\�P"O4h�a�Xu�9i�I�7���Q�"O\!ˑ��<(<t�)�	?2��U��"O ��cS�V��89�o�GC|
�"OV���:n|P��ޖ;�P�b�"Oh��s!��$�d�sI@)M*���yRh��j�<"ĠC���
�膧�yr���%��@
�ܵ�����y��7.�`H��N�g����Y��y2�W�Z�i+G*x�:���L��y��Tk�h��5O�$ph��	΍�yr��%w��a��_"p�B�r��9�y��	*4��j։4XE�F��y���S݈ɣ3nQ$���gd���yB/!|N��5dɤU���G ��yr�+��ie�ȉ"���c� ���y�mF�A;�ab�Y $0JA��y��I������*L�h�6���yr��M�$}�Ƙ�Smx5�5!"�y��W�k�J��F��9`��� ����y���<@�K�D�%�Mb����y�-�$'�� �0�H�K�(�yU�;�@��'�ס�*wL�5�y���17���c�=2�\B�. 
�y�ժqU��YvE��t���j�
[��y�΀�Rܡٵ�K0$�$	f��y2益^��P�dJJ�"mIB#�;�yRf��;�dͨc��G#��"�՗�yBoK�N��d��BJ�[�#'�yaA1{��mr4�F�&+н�Rʞ4�y2OS�rH����B/	�d��b���yHQ�xr��E�}���N�y�-�S]�U8J\?d���9d����y�@.
����ܡV�0!��oþ�yb��5(T<�J��\5;q�ǅ�y�+�m�p�3g����Ejq��4�yR��0��јD�5ur	��/^��y
� �<Ҷ��{��3n�v
���"OX��ŅH�P��Ƀ�/�
�6��"O1��%��4�R=��o֠j�4=1�"Ol��C�,bPiW��|L�AV"Op���9"rӴ��7i���e�	���g��r"�V�'���^?9��	;|�]�c�[0N	�@Zj�����?��xhN� d�R�%�}��\WN��Du>�rc-�E����wg£~|�hum3�B���2b"�v%�:-
|`!��ީ�McƧ�P���Y�Ʒc�*����Lb�'a1;���?QI~��4���j'��B��s����O�����'��'���'�^� Wg� �h���^2z�p�
�y6���'��&�I�26Z�ѐφPHD�Ɋ�~r�:c546��OL���|r�)�?Y���M[ ̴km (���[�m�08�ʌeF�:Ն��{�t��7 d����Ao�.���)b��EP�8���5I�4q�Hh1wi�&�k�P��ٚ�H�������>�5�~��3,l{���	.��Q�1��o�l�"�d�O�p��J��i���K���#����5ď�
�.,��'�2\�LD{*� !0NR���TW�$��剎�Ms�i;��]0$�L��Ĥ,b�l�!�S����?�$�W�5�,@`���?���?��U?�m�[A���ÅDE��-s���5�`�fb	�`R�9�ϔ*�M�5����Q�'���*v��}��e�\�|���d��X�>=h�|) ғ`C���	L�@��y�<�$��+�:̚��H"UV����� �M��)���'�
����D�Op�>)f���
1<0���H�%;N,��Iw�'>�1xDm'l���o[��"0X�G̦-�	M�I5��I�<�� c1�J�,G0�8¶.B�~1���#�?��?����0���?i�^���p�xǄ�	��sμYb�uE���7#��n��d����B#?1�*A7.��Ē�!�����:PN�[�8M��ǄJ�������4�$���,I���X���O�6퇂`R��geM�_p�(d��"v�~N<i��?I�*���:F�D"4΀-Sa��39D����II����Ll��:E��.�.؉ ���Y��DHঁ��4����Y��$nZ����E�DG�ty�Mk4$4������jt�����O|���O|� �!�):Yx��%�G,]����
��!��e��zq�R"Y�d�q&���HO���s��6��=���/Z��(1=��Z�,� I(�	��m�֍[�$�/�HO~-Z��'�rbg�X��~r��\�15�\�T
�XG�ju�~R�4�����G�T��^�%Վ�P��'m|9��I��ݴ�M�!�:�aK�nE�}8��_���6mK2JR���'�b�'9����l��'6GH�p�6��߾
�bTa�$
s��D�"�Q�ʏl:j��r`�����_>A���ہo�W��5jf�9V8����������V��ST��i�F���$���
��\c���&E�Lo|,)X6r��8�4B�\�	񟈨ڴ�?����i�>�2�CZ�t�,�Ё	�C�p\��'�"�'!�m�!�V�_��s�&��B�lB�'��'�z7mDF질b^wfpH�A�m�PԒ�#l�`�ff)�D;lO�(�  �   6   Ĵ���	��Z�Zvi��:+���3��H�ݴ���qe"���@"<A�iB���gC`�����Q�R�y��U�6��7�i�X�����f�TYؔ�.(�r��j�j�ቄ@2�Г�i��̩�+�>8Y�A�Ϭ\?�Y�.O����I_>7r�P�_��Rs.H=_��8�>�@��/H^.Mr��S��
�r㠞�?B�r��r�$�	�< �"{������
���[�$z���SF��F0��&�� �x3D��$oy�M��Li���R��8���4@x�'��Fx��Ba�I9Н�s�a�X�SE&,T��	69x�\��ቱ�PH���>��8[��P�<����ď��O��	�O��ҀK\lQ,��	x�N�i1�>��-tB�� ����^-:�0��I���!�a|���������O�H-�'!y� bf�T��jԋ�st�O����d����� a2�l���S.e�P�Е�	�ai�	9NF�$!7���(]n����@}ƴX��`��G/"�*��Z$�O�@s��;FT�kS����p��J�V�
!�<y��!ϬOF	�e���Y�I�(�n<b��OR�����Z��ē��D�,Nb�(jB�K��P��J�U��x��J�G�\Iml�D�9jE����'X ��j�-߃x�	j0��n�Q,O��p�O�{8�'@ \�gC����axr��S�P�k���U��C�P��s!C~�<CI>�'yQ�x B����W*W�~�.��"E-D�蓇�   ��L�;�) D�(�e���8Z�A��	�5r�Y�b��>і�6@�����;I�U��aʤ	�H��`��ra}�Ɋ���)� l�����?��j���#�.�z�"Oz0�seۅ6#�T�!L^�*�:=R$���z1�wm˥v�>	�$��._)�L�f�W
E���<D�th5�V�p�UұBҗ]����u�Z�h�Z�O]�4\�u��?Zﺓ�4]%��2�z��x�收#����'�O`(���C���ݹ�� �d�H�dD�-N�"[��߿�J���Ɣل�	?4Ƹ�Za�<n���n�T5�3�	�R#�Q�g�L����P� � >�p���D\1�	�`�r�CM��y"�Q6u�hu��9=
�X�ǃSy"Eճ����`�?O�k��V=r�D�?�X�#J�+V� ����$q�p�#D���S�
n&���0�G�7i�	U+N?|Uޡ�    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  ��   �  ?  �  �  �)  5  k@  �K  �V  4b  sm  �x  ��  g�  
�  ��  �  e�  ��  �  +�  }�  �  }�  ��  S�  ��  .�  ��  ��  5�  y   � l 
 �$ �- &4 �= �E zL �R Y �]  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+���6+\�s
�<4�d5h��'�B�'���'	�'/�'�B�'��(#`/�P`b2-��
�v1��'�'�2�'���'�R�'���'�APΚ<�z-�,�Ŧ�@��'�"�'��'���'�r�'�"�'�d=Q�n۶P�r�B�oM� ��+��'��'�r�'	r�'���'�B�'�ҩ�Ƃ��K��Y�RmɂX>����'S��'���'�b�'�2�'B�']t(�t��7���A�k����'(b�'���'���'b�'a��'&:)'Ƈ�S�d��R�k�ܵ�c�']��'U"�'a��'e��'���'S����l�/U$�L�*ĶI�.����'���'���'9"�'2r�'�B�'��l��Ѡ{h�1� �"PN�e)��'nR�'���'(��'�B�'DR�'`\|ؕg�
Ɗ}���sʎ�{�'f��'j��'�2�'�r�'���'hT�	���,8������=�q7�'���'`��'�r�'���'��'� xRP�ڜX0x �S8�D���'
�'���'J��'
b�'2r�'.i�B�{����Y0�ㆀ`8��'���'��'��'ZR6�O��$��x.��2��/_��0��ؼw+���'��R�b>�p��Fɉ�ʊx��j� ��%a��U,h]a�O"l�D��|��?�D�٦����ǯ�/V��4(�@�*�?��^�J�4���e>�#�����y�F��&�"6|�u@�?��b��Iiy"�S�JQB}�sa�!b�-�T6J� �+޴����<!����r��N�a��� BG�w��Mh���}���O��ID}���͈�2�F6Ob�Sel�Fľ$�p�3zZ-�6O~�	��?9��5��|��_�6L1� g��5�֩�TZ�,͓���:�$ Ц��1�	8�J����8xJ�i`��фJ�\��?�EY�����<���d�Y��m%�C&kͅi? ��'b�,Ú<�~�����ڟ �%�'�n8*1��<G*�}P�l�
^]B�:[���'\��9O@m�Uj
2z���B�/L�>��"3O(`nZ�!^�ڛV�4���r���^j�����V����8On�D�O���9W��6� ?)�O���镇=B��
�F@#NYE�J��zL�P�K>�.O��O����Ol���O��CC@�O��gI1
5���d�<	��i��<�q�'��'M��y����{a�8Ѯ�:5��<A�3M�ꓶ?�����S�'ؠZ�	?\�zM�f&	D�Ɂ�K!�d��'�4��+
֟�*��|�[�(�֍��C���XR�G�J�n�E�H��`�Iڟ���̟�uy�x�(�@��O*�IkÆR�09E�W�"�
���OlilW���ߟЖ'�>8��ܐ�l8� VT{ԍP_K�&���X1�ѽ�dd�S���i�g�ZC�Dzp�Y(Ŕ0n�`�������ҟ���ş��J��T�4����^�n�
3�ֱ�?A���?ɔ�i��@3�Ojbca�6�O�5#b'�;sR���ˢY��Eل���O�yw�1�4��$Z39v�lSV��\��8q��R�
�!�iM��?�Uk#�ĭ<����?���?��υ"�����b�����8�?!�����9w`ȟ@�	˟T�O6�-�w��#�yi�O�G9Ld��O
��'�b�'�ɧ�)@5j��c�R�g�X8@����)�D���Y8*捬<ͧ0�h�䙷��1�(mXP�Y�?o�L���ɠG�:����?a��?��S�'��D�-R0fG(7��};���/��X�V&śJt��I��l��4��'����?)�h��8�@ȺҌ�Fx1��/ʆ�?��D�ش�������l��l1�.OV��O3�2 F�z�ْ�;O�ʓ�?	��?���?������G�~���6#XNj83�)�'M���nڠC�d��'������;'3<���ƙf�>����.���	ɟ�%�b>��Q��ҦI��*BQngN��'��(`LĂS?O��D��;�?��$�d�<ͧ�?�&��Q@�
`閲|��"T��?y���?����$�Ԧ]�`o��@�I����`N�d�3����S�J|`|��?�cP�`��ɟ$������uf0�Sa���8MӇ�&?�u�ȤU>���O�Ķ\?�����?Y���@�88c�Һa�txj��?����?���?�����O��bp����x��� X�'d�pf�ON�m-B�I̟d�4���y�j��&7P�ւ݀2R�4�`▬�yr�'m�'��ˢ�iT�I)�(Ȱe۟f�����N�j���'�x��(�C?�D�<����?i���?���y�Νmq�ZfJ�^��gả��ɦ�Am�xy�'��}R��>/��jSގV?��wk�g}��'p2�|���V��T8��!M}z�ӑ��
GeP1˔�i��	�.�I��Ov�O�ʓW�%��aD�Q�R�`u%�!||���?q��?��|�)OHl��[e<���*�LU��/K=i4B
�z�8�ɏ�M���	�>i��?��N@ �M��GR@�	'%�/P�H�ɛ�M��O�D�BR������ �P(�R�7D�-����5A5�:12O(���O8�D�O���O��?�(��
m@1"��G�>F
@��̟����hhٴ0a��ϧ�?QQ�i�'�zeD*iA�Y�$�/^�Iw�|��'��O��d@%�i2��A�^u�1(P�5�����ND�X=N��f_����4�D�<�'�?Q���?���)~�,e3�̂�s�H����9�?)�����٩ ��@�	����OE,��f�:%0���`�E ~�d(��O,y�'�R�'`ɧ�I��b�1!�3��Z��3:�v0)Kn��B�i*�i>ᑳ�O��O��I�Ȇ!f�,`'ǝN�f���m�O�d�O����O1��ʓ!�֎�� PZ���G�]�����V���@�'�"gq��PS�OB��dlH�����
x�ycD��d�����OTA��Ӿ�Ӻ[�/7�*cD�<�@�>��% `� "F$鑭
�<�+O����O��d�O��d�O�ʧV�A���qB��!�M�l�`��b�i2�$x`�':B�'��y�z��n�"�d��.̢@0I���J�`]��$�OƒO1��h!�Hhӈ�_S�R�b�\u�s�T�1'n�	!5s���%�'}J$���'B�'�@�wΖ�*P��3"Q�F����'�r�'_�2ߴg�T���?���62��#c�Ր1ȸA�EϞUL �{�Ҡ�>!���?N>��	1!�f!����_^ K��u~rG9�,a���O�.q�	�gr
�f0�%L�$0�@��Efɸ���'�"�'M��S�������9�M!�2X_>�RQ���۴	�F�Q.OLn�N�Ӽ#�Θ����e�Bx`�����<��?Q�*P*��۴���6�yS�'f��c�6����dl�1M.�P� ޝ����4�X���O���O���V5%�� �nE�M�Bp�ბ�˓69���#�	П����IX�d:�lŏ~�0��p+K=k���ɟt�	G�)�S����p��+| <@[FJ�-X�N����-�h�Z����S��O��pM>�+O�T`�(�'#���x�BQ+y��<W-�O����O8�D�O�<�ֿi�h���'z�q���c�f��֖9�B����'1�6�3�ɥ����O�ʓ}�X`��#����ї)t���cC�M+�O�` .޷����!���שּׂ��)�
U^tx�vEϿqv](a<O��$�O`��O8�d�O��?�c	�E���ֆ+К��L������ҟX9�4$Nȍ�O�~7�+�$�(=iH=��I_����&L϶�v�O��D�O��^��6�1?�;iHx�Bƙ�D5Ba��'2u�h� �(�?T=��<I��?9���?	F�R~�m	�c�__t��S&"�?�����dFͦ�ç.L���	�ĕO�1�w���i�Q���Ǳb�<���Oze�'r���?�1s�A�zD��%��#�a3Q����Gqȭ���K���!'�|BG��y�<��P��o���C�6S�'BR�' ��^����4C-qJ4��ܰ2,�>L�T��+['�?Q�~��D�p}b�'��mq�0"t�!j�*8�����'�r��
%�������CL����~Jh̀4�X09�ǘ����jA�<a+OX�D�O��D�O�D�O��'!x�Q�Ɏ g1���⍑5K��!��i� }��'Qr�'@�OR�Li��A�P�	�bN���򆪂(PcZ���O�O1�P�PEia����*2�;p�!R�̈Z�]���	��D2��'�J$�L�'��'t���1��Z��dеa��[�Lig�'���'(�S���4Z��Z���?��/����C�[2d��*2K��[� �Ҋa�>���?iJ>u(��s�и����+>:$P��F~RÒWh>IP�K���Oe<Y�ɹ �"�0 �N�� B�@��Ӈ�����'P��'�S韐:c��*�8��G���ykꟄ(�4[hJl�.O�m�J�Ӽ��`��#��1�YS� ��nC�<9���?����,��ش��d�#�,����0N@�R��B!7��U�O"1Ȑ1r+4�į<�'�?)��?���?	7�!�(8 D%W�"����N(��D��%����ٟ���ɟ&?����Nz���	ٕ|�l��=b9Rp�O.��.�)��?�� �Ua��y$@*Lū0�݋A`H
X$I�'�����oF��T���|�_��
���L@x'�>QN�}�"G��t�	��$����sy�H~�K1��O�� ����&i
�:!�� ��\W2O|l�c��P�I�����ߟ�Ѐ�1A��ٵ_4Jf2T(&O���o�R~B��1<&60��Rܧ���r�[;R����ᗼXL�w͝�<)��?���?����?���cJ�7�h�!uhR1:j�v�
{2��'�b�|�^aSs�<	!�i|�'����Pm��g:\���ڳTb&����|��'�O"�蹕�i���-68p!у�!*Na��U�g�,���8�TV�	Ry�O�R�'^B+S22`n�	����G��1��Q�b�'��	��M��Q�?��?)��hJwf?R� t���Lt�E�����O���O.�O�S�\d�h��D4ny��z�FL�?::��E#��S�T��6�/?�'4����9��'vة��&q�p3hӏ-kzDp�'���'�b���O�剐�M��, !BHPUb�|���B�!e\$���?��iB�O�y�'�"8"%��������� a�R4r��'�P���i9�	od���O4�g�? �\
�.��C�+@���(�Ti�3Op��?���?y���?����ɓ!r	��8g���Q��+`�~��Yo����I�� ��f��r���w{��!��#<���̐"2�����'��O1�����bӞ�ɦ0xP�Y7':&^�M�lB0^Ҭ�ɛuEs��'�& &���'���'-�0�BD��\w�=`�&]5͘�+u�'Q��'}r]�\�ڴv�D4����?��2)\��ʸ��m�6#A>-�|<:��o�>����?�N>�����/R!�	� ^��L[V+Mf~R�4�B�Ǿi������'��C�,5�n�T�B��*�h�n~�'�2�'�b�Ο<j��\��A�3��L���Cd������40��qP-OR0m�Y�Ӽe��,�d�8�,�*S�R�cGA�<����?�|�HY�4��T�<��y�';c�LRsHUH>�''܍%$ �ȕ�)��<�'�?����?!��?�aK�w*ƀj�hG�������d���MEBM�X����0$?U��=�L�B��.]�`mzW+ɜJ�DY�O��d�O�O1�LpI��ư\�v��&�K�b�PF���<6��\yk�"
��U������E�t�y��R�4�KQ)I�`���OR���O �4�2�<���OT�C��=r��M���ٗG��0�f�nm���$㟰�O����O��$�*'��-�䌒�j�^�')S�E�fT�T|Ӯ�L�~�J�>�>Q��5��MY0��	�t�3֭�>^`�ԟ�������I����t�'W��"���v!b��*:��R��?A�֛F��6P��ɨ�M+H>ID皫ь=��/*��f/C����?���|�ƀA��M+�O뮑+*o��G�pz��6eԘ �!�F�Od$@M>*OR���O ���O,aă�@?��a�k�&�`V��Of���<i��i��l �'���'O��6�h1���a��#j?�IZ�O���'���'Dɧ���o�$x�0���N� i)!lN�mj�X�+��c�8����擸��)_`��A&\��n��P��e�e�H��� �	��d�Iܟ��)�[y�Gz�@��޾sҾ*1��X��ɠ����{�˓{i�V�$
Z}��'��U�w���.>��Ȗb�3I���a�'C��/W����a!���x0�D�~�bE��>*x�3�a˘X~*2�<�+O`�d�O��D�O����O��'��(Pjw�R\�V	��H¶l"�i�2]���'���'
�O�rcx��NYdjd���ĕK.�pf� E���D&�)��L��m��<	�H�k��H��sN�J���<�O��4���Z!����$�O����3�ސcF�ӱf���� Gޜ�2�$�O��O�˓����_*Ql�ğB�h�dֶ|�CP�9����6#X`��I��	П|�?�`R�CA~X
�>^�;�J�n~"*�%5��p���3Q�O��d��2Q_ۛxU����2Ú�ipI�J���'"��'���s���e���
m�<hèJ"�Rq@����D)��r��J՟���M���w����d��AZWbR��5��n�8�Ipy"�Ӵ2��������/��)��DH�V�nu��ې���� �D�nu'��'���'d��'��'����D��::5�ւ�-&�,��X�,i޴d�<5����?1�����<��C _ ��ʠlH0.^�Y@���x<�I����z�)��48�1u�ܱQ���%'�\�0,�S��=�'�s& ��g�|2V�pa'��?$A��U�=�<��sAٟ�����t�	���py�ee�`�S2��OH�`f+��<Y�r�ߛs�>(�=O8ll�f�]���|�	�|B��C�@�ܩ�/�:E�p[��/R-�|n�D~�m��k��F���w1%�2��v�N5`���hZȰ�'B��'�2�'-��'���L��n� s��Y�An�� ��O �d�O��l�?s[�ѕ'y�6m:���K���U\�%J�	���"�h�O���O�)ԍ�5޴��D��c��IЅ� �R��pI�	��"�X�i܄�?y��+�D�<ͧ�?9���?ia��M��=�c�$,�Ѕ��
��?�$���$J�Iє��?���ԟH���?���H
>d��$��*!��%��Go���I���$�Ov�OR�'�?�ig�-8���#9��īf�Q0�
�� ߙI�2Y�)O�����?�di.��<]���bG=W�>=ZR��W��$�OP��O@��	�<11�i�5����p"�0M�i����(�(��'|�6-9��6��D�O��2 ��	�h��g!�=���B�O0���)�6M>?�$�ǻ>��>�Y�S�y�aD�K�����n�ȕ'#2�';r�'b�'���I��؈���,!�Ej�@˿m��i�4+�ذ-O��D;���O�hoz޵K��0h���2�W�XT�U�I㟈��j�)��d�N�o��<1���
D(+Ő# o�@�_�<�@�J�:P�I`�I\y�'~2ǟi�,,���R�B�\�[�E�f��'.r�'I�I'�M�f��?Q��?�a�<,N��g� �@��n���'����?����V*�2�S�3{80��EQ3	*���'e�0aT/N%T���,Y��'�Q�Ƈʴp���i$*L�/0E���'P��'�r�'0�>i�	
;�d���H%I[>��M��:���%�M��ꇧ�?��G���4��%K`	�N������21&�)Q8OP�D�<I����M{�Oh,�b"�b`� $\�`�x���8,�.�Z���i+�d�<����?9���?���?��Pxaɪ@�/W2��R$�7��d
ɦ e*T�$�	��L$?-�	�m��P�NL���p�S�^ӊ�ЮOp���O
�O1�v���c�3-p��A�.��0���)�kb�<����\P�S+��%�x�ky�-N|��Y0@�W4\ �A�b�'��'m���S��@ߴkL�x����Tx����82.��i B�m͓}�����o}��'~��'쀐Xf�=Yr~�#$å+�0�J��MZ�������bԸ 'Q>��%Y�2��&%ʫ6�<�9WhI�z���P�	ݟ�����t�In��)M�-jV睽jizSπ� �N��*O�DD����<
E�i)�')&�놉�,��E��rʔ<X��|B�'��O=�Dk��i��	�I�������&h��K���|��b��ֈN�d7�D�<���?����?��� �M�BA��TD)��S&�?����ꦡ����T�����O��y�6ɓ�r/TMÂ��X��Ya�O��'C���?�Rv�άA}Z���5G,=�d+e�0��]+�0���ԀD��pS�|��ȫg��� �z���ѳę1{��'B�'t���X��ش,Ԥ)��[�3=X�2Úg�.H��j���D�Ȧ�?�2R���I)K�ft�S�Ē0�6���@JՅP�d�	�?@dl�R~��O�_����@�ɒ�jؕLׂ=�6A���-\�Ķ<����?A���?!���?1(�0ոǮ̰���3V)Ai�zAq��[٦�Zb%Uyb�'��6Dmz�k���(m�����
1rr���a	�����}�)�.� mn��<iI�R�"��0LQ��Jfn��<)5�E�d���	r��ry�O���T���02��%g�����,��2�'���'��I��M���3�?Y���?��J�h�H8�/R.F@�a V р��'bꓨ?9���Y�����ʜWK��Z�ݑ ^|)�'���au��>�К�������"�'�ځAF[1��Ʌׁ�������I˟d�	ퟤF���'�6q�����4�EMGpu�(XA�'J�7-�1F������4�]���X�HHkW��Jˤ��t1O����Ob��$7&?�u��2c"6�)M
\H"5��"�V��\�W��`�M>���?ͧ�?����?���?9�b�#I�����cN<���Ŧ�?���`�V�#6�S�?������?q�i���O0 A��A�7�2G��<6=:\���O���O��������u�R}��8��kԊ}J4��L���"�%
*B�Bɺ�@�(��KN�恲��T� �O�˓u,]�F Ke+���Ak�m������?���?��|R/O��o��L$����#Q����GM��N� 颡β$�t��3�M#���>	�����7iX)�o�8sD���Ld�R��}���|^9�-����J~b�����`r@�2r�|q�!�0j]:mϓ�?����?���?����Os0(˔k��?`ȩA"O�'}�H�'���'�d7�� h��c�F�|��R*�i�ŠƑG��|j¨��5��'9���Df]�rO�f��0����L>bA�t-	���1E�ӵ>`��ɴ�'�B%$�����4�'�2�'�`i�&�9)<����&E�0��')P�`��4J���i���?����򩃄$M><���'xj�`�v	
.5�I(���O���m���Y��V�k�*����"m 4��F)O�8-6����+��4������J���O��3�3X�b��T�xp���bh�O���O��$�O1�4�����8�:����3�D�"c[�?�v1�'bKj�`�@��O���v�l��C+�0���˔��>�����ɛ�4���F�"���(�'NI�˓P��4Ҷ�υmy��"ŮMd��(ϓ���O��D�O���Op�d�|zAH�k2�����"%S"�;�-	�tA�vnשu>�	۟�&?!�I0�M�;5|��\�]CU"O�;��A��?�M>�|"���M��')�\�Ԣ�*%�|<�c(����h�',�R�C?�O>�/O�	�O��Pè�#!~,�v�F��L�����OH�D�O��$�<�i�`�22W���I�ZF�H�#	�Rft+e+��8I�1�? W�H�	_�"�ܘ���\�!�b�8QL���R��'B(��`zȱ Ð���_럤 S�'N6a���%~�H$@!��\�n\�3�'��'���'U�>5�	�e���&�A-u�(��Ȓ"m����I��M��\�?A�ʛ&�4�p�B���,�0��G�i�6O �Ŀ<�U�Mk�O���&��B��>I��4�b!ڸqL����ڼN�̒O�ʓ�?	��?���?���~G.�+��Y=W��`�MG6z��-O��nڑt����蟤�Ik��4����V1�Cu@	�P&�xZQG������O`��3���X���m�3a_@�,�GN��AY�X��u�̖'Ӕ���|?�O>I+OX��c"�
@Q^,@SG؂]�^0"��O���O��O�<a��i`l�y��'��u�a�-����)U k�c7�'��71�I���$�O��4�T�B�Ԋz��9�
��֩�����7m,?Q�3_���D��ߩS�`� ƀ�����0�Q0�{��I�x��Ο��I����%T�,0b� �LŖ��(��6�?���?1R�ie�Y�Z�J޴��GL�a�FLm-ҙ)f�A9���RL>)��?�'y	L��ܴ���J� ����	�]U��S��>XX�!����?�UE.�Ĭ<ͧ�?y���?�G>X T�cE�_�v���!�H��?����d��E8(��4�I��ܔO� �P-��5��CFO��N�)�O&��'�"�'�ɧ�IA<<�2H�,Ы\ :�Pu�H�B�c2K
$}���n0?�'/���$W��VxF%��o޲��[�ʆC������?I���?��Ş��Dʦ�;�M�.d��$��&��r�>uS�eX�v�����,"�4��'-�듴?D΄S�Iz�����J���k��?q�>t�C�4���Ճg��$:��4c�.��󢉞I���+�	�y�Z� �I����	����IǟėO�Ll��-�{�\�W��J���n��5�r�L��D�O��i����$�OD�4���".ר]V����B�lt�}8��O2�O��4�����O��K��w���	�G�T�kCO�s�.���'8���ɾ6�+g�'y�$��'��'FN�Å,#M|�7�\ `;�AA�'�r�'��R�Њ޴G������?���@CA��G��J���;C��1C�j���>����?yK>I@m�Pc�i��5:�l���
�y~�Dk�<Y�����O�>I�	�)
�h���̓�-d9��R0
���'�r�'<��� �v/��"��ak�+4�,���G������4a�iY-O\]oN�Ӽ�� �>�0��2���T�����<�����䛦p��7m<?逎i�<I�S}�J�d!�m�<���.˨|y\k�|�^����ӟx��ퟀ��������/3wL�	�K�t�ÅKyB#vӐ}¶��OT�d�O撟�$޳&`��a�KrY\I� C��8�'���'�ɧ�OXX ���n>JK�݃bFm���b\��"�Oƌz%�N%�?�E�'�Į<9&J�/{���RƲYQz�ó�A#�?a���?����?�'��DZ���C��ܫ�$�x��)Aʡd�h�S��m���ߴ��'��듃?9���?��O:6@N麄�EK	E�U�4��!�M��O)�U��?�R����w_�!a�HO��� ��/G�x7��	�'���'���'G2�'��RT�ǟ�t���@�h�R�I�O����O�0l"�<��'�p6�)��4���b�V��K�m��@�O\�d�O�)[�7�)?I!Ĉ*`5BC�3)ֈ@IA"_qbpF���L%�<���T�'�2�'v���m��?������6�� �'�'�"R�T��41��yK��?�����IZ!W[>�[�IH�`�� a@h^*E��	9��d�O$��'X����f�ҋZ�P�	L�F(u�J,r�H��K3��4��i`�-�>�OX�e�ZE�x�#�H/y�)���O����O��$�O1���u���������D�{)0iX��iѤ� p]��ܴ��'%0��?y���:9��f(A��FIQh��?��-m6`q۴���O�q'�j�����B���T��`�\�1�n�U��ly��'V�'�"�'IT>��D��X�N,R*D7v�� SEٛ�M�H���?���?I~���Qe��w<z"���	����J_03G� ���'��O1���#b�R�	�Z�,�$�µP\,	dJ�%��IJ�*x�Q�'���$�t�'"��'���B����}j�|ہ�S�X���V�'u"�'R[�����{�tT�I�x�Ɏ4�|���b�:	ADXb�H�N����?9�Y�D���4$���� �V�Ȕ2Q�O�.= �
,?!eb<���ڴ��O6z\��?�b��M����&���7ٚ�%�?���?���?ً���O$�nʵ�i �پJ�e����O"n� i�%�I���(ش���yG��+0�	 ��@;r�bC��E��y�'��'��0`¶iN�i�mB����?��"�S� �zu@�+n�L ����'����4������۟��	cO(hPʄ53��I��F 5�:��'�l6M�Z7
�D�O"��:��O��+���lڔ`jLC�<�	qK�>������O��2��Ժc��|A+S�"�6��0���<"H��[�`�ԉ�&_/��|�Ify��ߔ7�*J�%�j�r ��(���'�"�'!�O��	��M��n�?ٵ�U,f� Q;��3y�.�4��?	ýi��O�u�'�"�'�����yꁋؑ[Cz�wgII�*��q�i$���%w$���S��)p1��yI����핃j��Qrbc���	�,�	�<�I͟��z�hʇW���A��A%W���E偉��d�O�Aoڜ7kN�럸X�4��/��Ux�H�;j*��v���B�61�<������oOX6-%?�b�Y�L�2�#UZ�>�(d�ٞ���s�n�OX��O>a(O����OD���O\D�w�cB��`רcn�͒ՠ�O
�d�<95�i���e�'
r�'��*"�1�E�L�8��Ee�^���1���� �	q�)�14 ��)�p ��>/$��6��s�A�#ʈ �����g�П��Ǘ|B��9��x��,S>�8yu"���'���'5���\���ڴ.A�h�4�I�8�2�c�&�'9@�+������ڦ��?	�V���	� �M&�R97�� �U�M���I�����B����u��R<6���UVy��2Dt�"fi�4��)�чĀ�yT����ԟ(��۟��㟤�OS��AB������e�w�A�R�a��٘���O��D�O��?E�������\7��P�I��U/Pa8� �;�?q���ŞZ,}�ߴ�y
�  ���	��E���Q#)*��(B=O���FHI��? �3��<����?��n��O�����L�0�p���?����?����_��aG��(�	˟@�3Ł�+F��A������G��u��d�������	_�-{�F�j2�`9 b�>7���dj�!w��#Rn��|Rga�O�����
���IJ�No����Q�Ҩ����?���?A��h�P�d��� s��3	9|�Csg٠�D�-�g�nyү`���ݼ�\}�Ջ##��Is�@ T���ן0�'�4u�5�i��I�4�
,Ru�O�\Aᆤ�% t@���Ì�K�F���YF��Xy��'���'U2�'.R.(kkj��G��,�h��"�e��I�M�EÏ��?���?����
%޾�X�*[n������� �>������O� �����aτ)x��j�p���LѤ(����vX�D���1D��K�s�	qyb�O5 L��@��W�&�2�����';b�'��O�	��M#�d���?����@jXʐ�3,G��('̂��?��i�O8 �'�R�'5Ҍ:}����5��dŬd:Y�m跈9�M{�O�@��AX��(���n�q$����Z�1�҆S:���O����O~�D�O���8�� c֑���ڽ��K0" >6���	���ɨ�MC����$�ɦ�&�ܐ$��'r��'o��U�� �O��p�i>q�E�ئ)�'6$��#n��K�b�z%끾s�B٪���"�Y�I�W��'��i>	�I�����ٜ�*�H�7�P���ˆ'�
��I럸�'ظ6�xOR��OD���|�5/����5�'f%B=QU�A~R�>Q��?YH>�O��R#�2�(� C"!&��hgA��-�L�C���>l�i>9C�'4��$��Z�.0a�������m(E�l��ԟ��	��b>ٕ'�7-p@><���Cg�p�.�1`��Q!d�O���H��!�?�N}��'I���ᩚ W�ܐl�i�Ph��\�L��L �-�'���r%�M�?m��_���C&��� f�Q9l��"�x�l�'�'r2�'�'H��5f��y4�ޤ1b:��G�o�4D��4H�Ѓ���?������?����y'��|IhT�G=x!�Q�X���'mɧ�O��q1�i���	0*�i���E1b+4�.�󄝦_�@K�'Y�'!�i>��ɐ
c���f�0'�������#!�t��ʟ���<�'m6�\taV���O���`�>S.�/b ��LE<"��0ªO��$>���.M"�c/��t���>C��-*�Ћ�|��3L~��+�O��{��IHu�+�<5��!��EW�D(��?���?)��h���*hR����־'��)��]!>���AݦqhCʄ��I��M��w�Q�
�=�d�L�|ș'l�'GR��*1қ6��Y/��_ ��DI'E�PGi��ey$$�ꔸpM�p&� �����'/R�'��'�|�#�m];&|"�p��R�a�޼0Y��ڴ#��	���?�����<
_�Q��5C'" S��73��	ʟ�?�|:�N��a
!u)��	1���EÐX��YS�`���D�C|1+�[J�Ov�d;��7�Z�c�I1g̅(v
i��	(�M�ц�6�?i�Ҕ
tB�OQ�&� �+����?���i*�O,(�'�R��y���BBTl�D���^U+c�H�V����i����A�"�27�O�>�$?��=�*ae�}pܱ8#f�$I2�i��<S���J��C�[�o����qe��0����4{�4j#���OY�6�9���		��(�B�:؞Բ�ĀK,�O^���O�Z)K��6-8?�;$�������}�b
�d $�W@	��?9��7��<��nF'd*i ���bX��@�>�O��m�7���	ΟT��H���AH���!�U.��B�ڡ���j}B�'m�|ʟ�С����'P<!e)J6hO�,�G�D17��W�2��|�0%�OH=�J>YK]�B���H���|���PC�GE<i�i"�Q�2lR!40�Ȼ���:�0�H'
]/�"�'"�6�0�	!��D�O�kf��+f�)��(UB��pT-�O���
� ��7�5?��ǂh�b��GyB��-�(42r��F���R��L��y^�p��	 t�����	ʨ�
u�(�&+�D�ݴT�dE1���?�����O<�6=��x3e�h�(�h�%z�\ո���OF��"��i�.D�7-~�<��M�2Tp*)�`%�4�X���~�(C�҆R��5�ģ<q-O��#�a���`R'
Z$�����'M�7ʠa�����O���M�:%� �K��(%�
��r��⟸[�Oz���O,�O��z!/;�}����sTr���4���%��D$�i��$��$�����`�.I����S.o>�`X�f3D� �6ə'����`ғVm����B\��ش{DHZ���?1c�i!�O�N�m�@����L:z�
Q�0��-���O����O�xH&Jwӊ�Ӻ2dP���ƍ��V�r�&S�2�4����
�z�O>���ON�[S�ʫfQTLJ5o'���	a���޴%_�����?����OP*����[�'�(q�Gp����f��>9���?yL>�|ZR(Ob�? z�xT��V�pȁ��ʶm®1�Y�B̨˓*�	3� �O1�L>.O�*WHD� )��s�*D�	s"�'^F6�X�3����2*����νt�̱S����2���$�٦��?9dV������]+1�\�S!��*Z�*��E0sܘ)%�@٦!�'��1qӁ��?}�&����wf���R/EGҘ`fbKB�BA�'~R�'=�'}��'\�Xx��=!��)f�>SORd+��O`���O��nZ�r����쟨�۴���,�CB�əܖ٩��l��<����Ŏ;�6�-?Ɂ�=#6�n��OV<�3�A��^�(��O���K>1)O����O8�$�O,욦��O��@�t�V/X,T���O���<AR�i�d8Z �'u��'�Ө:�ٛч�pW��1.�9�D�n�������)�E�ŉFx��Z���,�h���K��\��EEU��Mk�O�U��~��|��B;�J�{�D�>�F�6�L;�2�'P�'2��D[��:ڴ+&�ԓZ �*��^ r��1��M�bЋ���?i5�i �O��'�S T��4�'���Z%�4f�9{a2�'���{u�i���(<��5r�����TԜAٔ����l�[�ߓi���<���?����?����?!.� d*S�ĜM�Z�/�)v�P�[��H�Q@�O�՟���ȟ,�r��yG���r����G��ww\CF�ΰC�R��)�//��7�s��j#댇0�ư�Tg��)X@t�k�|i̹Ipb��W�yy��'��
FD��4��J��Kf�����_�"���'���'��	*�M�gB���?���?�5ǌ&%+JT�a!�$�T�VI����U�O��>��&(<=�0c�.\1��"�,I���]���soM�c�PɛN~�S��OZ����{��ĳ1`�'iaFpk�T�2���?!���?	���h����]� sN(ɵ��1�r%�1,�*{���Ʀ�:�doy��n����H��}�KV�P<���mյRh���ߟ��I�����Ҧ��'��iZ5�[Bg�B	L����tS-u�����aޑ�����O����Oj���O��DD�`��,F���P1�4hH�ʓ;a��e�Q�b�' R��$�'�P�(f�<
�2���.B����d'�>)��?�M>�|�^����"E�m��V*W"���B�J��M0W����2R�D'��<�7NA�ʐl���mG>|�V��?i���?y���?ͧ��$�Ŧ��R����L�T�O�v ����f }��܊Vğ\`ߴ��'����?���?Y�oM�1\���� "�\���<��$�ش����3(,~�{�O�O-M�!e�\�fJ�p3čPfDK;�yr�'�"�'�'�r�	I��-@ �W� ���Dɏ#n]��D�O`�$Iئy��k>���MCJ>qҭ�m����ʈ�h��DB�����?A��|�d�J�M;�O�t+@��"є�����Cw�7>ݐ�X��JP?�L>a+O(�$�O>�d�O68Y�k�9s��P�$ 0G�Z	�,�O����<Y'�i���\�4�Ii��f,h� 2LAf�P�ǅ5����B}��'��|ʟ
�1��4e��� ����	3T� C^+�<ks�!�<�'5���	T�!n�z}�h��o�8����2��E�	������4�)�}y�q�e�F�I{����#A����Lոx�D�d�OJ8nZQ��A�����4������B�'�F��4@]�D�	�g�6�m�n~E@�iѢ�����K�{����c� I"�z��آz��$�<���?��?)���?�,�(�d�5�X�q�������L�֦�[1�ʟ$�Iӟ$?-����Mϻ����p1�`C?e�4pj����	@�)�Ӓ!O��l��<Y�K�6!<�)R���t�~a���<q��*�����䓨�d�OL�$.|��8)�ER{�r}j��2~@�d�O����O�ʓ2�6��7p���'-��$P ���$3�d��⇊:)��O�U�'���'��'�l��䃄>w�����Ӣ.2� ��Ot1+�EJ�e ���&1��H�X\lD�u���.D��jR<'`�Y_���Ѝ}�:UL\� �`�Vmx��]�]�� a���>�vyʓ�ۛ) ��f%֭4��+V�	9�}��%E�wd �a0w/�`���>)}qOrPiv�ߕ=.b�s�hѦ4Mt�kV  5gA\��`�޻I�Z�*���|1z���GS���)Ǩ(u$<+�"�}\"n\�Z֮ȷ	�أ#�A�:�<�p����-2���6,.t�
"Ny"�Ȱa��)E�@8c��D�.�l0��,�ZY�w��.L��h�`�_��B��\�?�Ȣ�g��� +yIF��'��	� $��ؠ}�T�CA��=e���VMLG�t�RA	K>���?a����s4��G�X*v$Gꊒx���#G�}�S���I\y��'V��'� ����	�~=�2�VhĄ�[&l��}�B[��������ImyB��.e*�Sq�*B�#׺4�NiR��A�&6��<����䓝?���i�) �'`œ���J�<Ă�+K�{׮qJ�O��D�O���<Q��݇,��S�����ʡ���c� Z�l_�h�2���M3�����?9��'����{BoB�^�,q��A�o��Z2��
�M���?�/OIq%��o��'���O�zU�
���Tr�Fa-zl ��5��OX�dq�p�'	�,��%�	kn����F�<mZy�
��~>^6��O���Or��K}Zc�u�t��T^X���DH��c�4�?	�t�Ʊ����)I�+{T���U8"��p�N1q��v��E46�O&�d�O���QF}bQ���� T��f�Ϸhiպ�,)h��9�Ѽi�:U���'��'���ĝ�^�n��G��>2�(�B�V�|�`�n�x�Iߟ��6J��d�<1���~퍲V0z̊Ǡ� �~�;�
���'�ޡqs�|2�'�B�'�Z�%�N<q�xɳu�^,c�	�v���$�T���'9�	ԟ�&��X�H�dI3��1\7p�'T�$�*�I�H�I>���?������pG�P�k_�YF�9$M��H2���e�WJ}�^����g�������9h
\�'����x������A�Ͼ��'���'�2R�@i�������h�n�c���AT�kfCC5�M�+O���;�$�O��=o��	_�5�2D��b
�1�A�0�Lꓹ?����?�-O�qACL�}���'�9!�-Z�!���@��&J��(��boӶ�D3���O������9}�JϽ�q�J>�d9�����M#��?�(O�1��J��<�s��*�*s�8��J�"8�� +�D�<I���?AM~�Ӻ;��C3��q��!�S�8��U�Kʦu�'�"<�g�lӎ��O���O^���H�t��+3�*��&��a�l�Ayb�']��$��2��i�$L�U�l�5
Y*ܾ(�ش(�����i���'��O7�O�),hk�$+�D�<W�����L�I_��l՟0�I���%���<����Z4�ϫ�j�Q�$�)d�>hcv�i���'(���m$HO�	�ON�	�~t��u�3~D��d�Ҋ0�7m�O�O����D�O��I�\7@ݚ� BRZ6��u�L'<�D6��O�8Pj�<�$R?5�?�
(<�Q�&B�n{�	�[�1�'"!��y"�'�؟Л���&L0p1	�Z6,�d+�eǹN2m�'{"�'��O��䴟����^���fG% Tfq��*�D!0�$�O,˓�?�DI������<j8D��*�f���9&���Mc���?��b�'3�	��7�ֺBA�5N!�Ȕa��ޜz��I�$�	�З'��EU��O1��хӡ}3�y)��`�H]cy�:�&��<ͧ�?9M?}X�?�P�cJ��;R�S�'|����<��_Ƣ(�.�v�D�O|���R$q���nh��
��@u+�����x�'��I[��#<�;Q/��ڦ�*��4!�?"�m�Uy�㏒a>26�_��<O�dM#?Q��$4vҴ��C�	�`�A�զY�'�"�'_��R�����O�FIÔkF)]�邢���Mc�뗨�?i��?9��,O�SO0�Y D'>��	��ۇ+�fm��O��s�)�֟8Y ��%[&=Ҷ�إv�Z�0CL�!�M��?��'TZ�r3�x�Oq��OJ�A�JS�J�0���n�.�r�Ƴi�B�|�~��?����?I�/.,2�q%C�5���LV�k��5O��a3=�4���0��}���R`���
 � +6�'���IK�	ȟД'B��nPx���95��R�� %:����V���Iʟ��?A��~r,Q���ȧ�Ot�
��M	�M��/�K~��'s"�'!�ӌxo�U̧D�n�2��	{���C�M3C��o�oy�'��T�	�#��j��z���L��t�kL�pz��5�
3����O��$�O�˓*]:��'^?�I�L�p�3!.|O�T3�F_�~F )޴�?Y-O���Ox�d�[�$�O���
5p��9Tܭ@v<�)��6!N�n�ɟ���NyZ`و���~���?���0�IIU���p2&��BM�_���X���	ן��	�o�����x�'7�i��QM��EnJ��v\�Q���D'�&Z�j��B#�M{���?�����S[���"U(ФJ6�W�UQP��48�6-�OD��ây��d6�D*��@j6@(�2U�FH ����7mJ2&d��n���	��������$�<��a�)�fh��(_&;�ָ3�����֤I��y2�'a�IT���?�N�6�8�SG�=Yw(Բ��(h���'r2�'^�i��j�>�+O~�d��[�kթL�p\S6��0�|"Эk�f���O��dвi5�?)�I럔���Uؔ!�vT���m�.:���4�?Q�NŊ.���sy��'N�����k�j}���]��Ap�,)P����� ̓�?1��?q���9O(X�6��c��PbAeԹ�c'7~�|`�'��	����'���'���	k� �C��?��
w�O�mM��"�';�ӟ���ԟ��O��h+<�I'��c�.�S���:BT�����i����\�'�b�'����yrN�5�P�H׋��M���1���6��O�D�Ot�d�<�e탦{���֘&nt��+�1K8p����C�7��OZ˓�?��?i4`�d~�O�s�A�O��1H�ƙ��U2t�i���'H�ɯJ�Ѩ�����O���S�L�>q�%���E'������
��`�'���'��Ƚ�yr]>��W�uf1|F�"EbY�N3U������'JܹsE�x�F�D�O�D��קu�G�\��L�Cj�4�z�G�M#��?�F���<Q!]?�F�'b�\(F��T�G-;8<oښb��Y9�4�?����?Y�'W�	Ny���:��k�H^�sG0L���;_5*6���(��2�ß|l��
�(�&&�ܚC�{4�l�ҟ$�I՟��j����$�<����~�dH'>}��)��T$I]>�j���9�M�L>Y���<�O�"�'� n�$��LF@��@k����6��O��j�(�H}�_����~y���5� .��@�>?��m�_�9�l;�P���#�e�������	��IOy�g؃L/,��R U��B9��l:DM�t��>	,O����<���?���w� �Hf�3�i���A!ʝ�����<�)O��$�O��Ħ<A7/�
���P��j�0�L f��q��ԒX��R���I_y�'���'0(ڛ'"�a��E[!�����ԁ-���� O�>���?i����d�b���O��E��TU�FN�B�4M��� <f�6��O�˓�?9��?�P-e~��M#��fx$��D��k�zP$oDʦ�����'�aq᫳~Z��?��'#�U����MD�0  \���I蟜���4Z&�Jy��'�i�Z�¸2�꟪8��ep�'V)P��F[� ��
��M���?9��2�W��J����D�5*ʩ�t��3=�7��Oj�J-D����O^˓��O:Z�����p�B�:�@),l�rڴe���$�i���'���Oc����DYP%���P�[A>!kvmW1��mZ�AZ����'w��䉞;���O�5� 8�g
X:O�B9nZ���I����!,_���į<	��~"ǍcV��B"#���1��0k�4����OHL"�0O��ޟ@�I�l1㋎��I $�)}F&�A֪�M����<��_���'d�T���i����j�!p.-�©G3���CȪ>�1�U~b�'���'��Z��
���?�p*��L�H,6���C�J�O�ʓ�?�,O��d�O,�$�JI鶏Ɉj��@�S�ǆF�Eв6O����O����O����<��,Z%0�	�<s9Vq�0� )g��Ar捵w#��^�|��Vy��'��'�L4S�O>��ňM�s�.l��/�(Iм�i���'�"�'A�ɹ6K��د�����r�#2-?UڞYbWG9#�}���i%�[�<��՟����'�F�B�d�
�\-2Rj����T#Ӌ��'�R�D�S�X���i�O*�$�
�GʘT�<d�щK5,�\��RA}��']��'eFiX�'�s�L��-,��i�c"l8�i
#È�
7֤o�^y�&ߑ�z6��O��D�O�	�O}Zw�h�	D�O���c"�B4)޴�?!��_��͓F��s���}Z�&=��Ez �rC�DÆ���q�@R�M���?9�������^��&LԜHjiX�i�1-��n���c�k���?)��۹d�r,0PF V2��f-��/��6�'��'�t�Xs*2��O<�Ķ��q��T@�pEc�n����{�v�OHU0O�S̟�������T�ۈc�z�z1�8��hsJN��M;��@C���Гx"�'���|Zc�$�c2��90��N�602�p�O�m+�5O���?��?�.Ov��q�%Z����T��m����ԯ>�]�>	����O���O~ ��ǋ8!S
 �b��(H��A@�Lڬ|�D�<����?a����s�t��'�VxS��b��Q�7�X�@-�j�I���&��	���t�d?q�B]�R�j�g��=SM�P�Q^}�'9r�'��I�U���O|ZׁG0U����s��E�zx��-h���'l�'Z��'�ZA���'���ȼ�t���3g>E���:���lZߟ���gy��^�X� �$��輘� !\QE����S�� 3�XO��۟��Ih�0�c��qڀKM1`L`�b̜�T6��
�����'�����fӀM�O�2�O"n�n��Y@f!��Ƥ"�ň1;`�n�����I��P��m��t�'bu6�Ѳ���'�0�FJ:LxmZ_4��ڴ�?����?���KR�O8���j�3s*�@[�)�j(�W�Iצ=0�g �d'��B�_�@"�A2���v��<� 4 &�i���'��8�O���OR�	"��I2D�*P��0J	x6m5�����?a�	ȟ|��+B\hҧ��y�BT�C�"X�ݴ�?ѥ,D>��O���-���D��6�Z��8��6��m�Q��!b�🸕'���'��V�lp�e
����C�Ub��X��Y�9��
�}��'��'6��'�Q`��ڬ_FH��Ųj&r�'bY�kl�U����؟���Vy�\qʐ瓖_�Hك^���ٹE��`˦�7���O"�O@���O~5�q�OƑ����-4z���V2���(��g}��'���'��I�c�ZxQN|�t�[2�J&��'WڄPG�47��V�'��'oB�'�dH��'��L�b8�w��v���F��e:hoZǟH��Yy�Q�x�����k,	v<h�m2)JiCS+2ױOX��?��Zw��@ӱm٤�HB��ۧA���[ߴ���C޶ n����I�O��i�`~��*p�)g���0UQ�G����d�<������'pq6�3M�;��H���ѻ3
�$m��h��a��ߟ,�R��?y,O��� 4�I�����7���\x}���O1���Ē�"t����R�ذ�#)�.{��o՟��	ڟ��3��?���|
��?����*>�ʜ�3��5�X��O�+ƱO
,+��D�O>��O�|�	?4�xѣߪ:���Є�jyr+[��?9����O��O2��v�O�NY���!�X��C�-Yn≃eN���?i��?���?���h�6��dC| �ԉ���'O�-��?���?q��䓪?y�'���+����Ɲ�A狀R�<,�ش�̍�'<"�'0�Q��#��8�����[��3���v���������O���O:⟘�r�~� *],2�(���ϯ5�89wS�����L�����	�,��D��ڟ����[2�G�|�vH��Y6L�b`l���$���I{yB�ݱ�ēR��S5@�?<�&��!I��;�mlZş0��dy%��)�����$������O��hdb!+�+�!L Ӏ�@�	Ƛ���O�#<9�O��l����*s��y��HW$Qo8Da�4��Ę�W�d�nZ��	�O��I�h~�НV�vlz�-S9�^͓��_��M���?I��o���OM��a%Aw7����䇹H��I��4|6�%�վi�r�'��OO�O&�$+�JՀQV�=�8�!���8��mn<h��#<E�$�'�jԡ���8ҢyY��=A>8���q���d�Op�$_�tV�5&���	�X��7}��ئ��6z�)���Ĉ;��(�>)d�P�<q��?��{3��P��I>`��rE�V|���c�i)�d�M��'z매?�J>Y�қ^�D��/ҏk�ٳG�~�'(ډH�O���O*��<i҆Y�E @8q�`�b`U���	m2�3�x��'s�'&�OL�@����'_(�4�N5�­���&U��?���?����?	�L��?9`OK�\�ĀZTǞ�ISf�QoX�`~���'�"�'#�'�2_��TJh�<�scKjڬP�3M��jQh�V�P��ɟ$�	[y� H�J����܀�� d~iR7"*��͎�5��k��ݟ0�	
PDb�d���DR��iC��8b,�od�<��O*ʓ1�|�A��4�'����b.�8��I�P���3�A&?�DO��D�O�`	7�	}j�bߋ5��e��'�1�X��H˦�'���d�`���O��ON�%�H}I��F�C�U9�*ԁ{oZ���	7R�#<�~BrJ�E.u�VJJ��C�Ȃ��!����	�M����?����֕xr�'R�ㄨN�"-�e��#��X��-��){�H���)�'�?�V�T�d���r#@P	*P�mӛ��'�b�'�t�b6:��Op�d���ypM�5k���LǛbNAs� #�ɶD��c�����,��5=](� Ό�di��A�H��6V����4�?�0�	L�O��d1���L���A�JEYɧ� {8�	�R�,"*���l������ΟlCDj^�^�VQ��/�7�$psV��
7R杖'���ҟ�&�t��R?)t@�}TB��P���]n�1c�eRզ��D`5?���?����Ă�l_�Xͧ9�&�0���$$�t�� Q^�'�b�'�����iE��+	�(�� ��1?�>U�h֧Dj&ꓹ?i���?Y���?��!������O QX0�UG.N=�����!3�DQ6.��=��m�	ڟ8�'���bN<�S��4 @����XԵ��������	˟��'�H!�):�i�O\����k�1B���+1LA���Y�[ξ'���I��Yc� ���t�^�>X|Q�cۂU��M�4o���M#(O&� u�U������d埮H�'hB�bc/�F�l���h��AWά�ܴ�?I��}�"�Gx��� [%#$ ��--L���Q��?����,3��c��?lO��9��٪MIL ��E�,�D@�a"O��:���A�q�V V�;���1�l��Y�x����dH��Bh�i���{4��U:��*�Q�'��qn��M�(�VΟ�9��	:3%�6�2�q	�`��I{�J��9G
� ¯���Q��̚�-�����&�*�B1��t��!�!��t������#c0:5�7�� <ЈPn�O��$�O���ĺ����?I�Ot\�q�D�ܙp`���4�X��g��$�l0w�ٚ7���b��	4Ny#?���+
����A�F[P����.�欒�M�"h�\����i<��E֜c{t�BW`�tO��b5�G�wz�!�2{V\�K�F.d�R�'ўt�?I���<B�J �͑��ъ�V�<�c�ϸB�:�S2����b�Ȥ��K�sm�IXyr�|:�^��ɘB�=!1ă%G& ��,B�rs<���ן�R�oB����	�|��Bͱb�f����E�$��!�~��Q�	:��Xr"���x�KJ<oI4�`Qd�(%��	%�����O�.��:�KD�0����Z�>���'��I	76�L�ℍ-��p�i!24bc�h��	�}~|�P��#L�� `fgU4}�<C���M�G= C��R�m�]ǚ���Z�<�(O0%�C�W}R�'��Ӻ}.� ��l��)���U�b�v��c� <A���ڟ4��I5VV���F�[���|(�tL��߁AmX9h���3� A�b�>�"$�9Pt����gٖ~�Q?e��d�����ɆEP,
�ĝ�m-}�m� �?����h�>���!y���26�ݶni,���>m9!��<D�>��V�D!a�0����m ax.0�n�t=����rH�Q1���p�}�&�i��'��S�uL0y��'�b�'��wW��C�	K�a1�BS JFV�f�|"�y2E�%Vcr����/ǄD�t�,��'|͛ϓv1|�w�_�o�<�C��U�qin9�y�@U��?�}&�������P�f����5��+D��V�
X~T��*��:5S��;?QW�)�'Tp�aWC�-E�d{"���'�:���LCQ8�Z���?����?qG�� �d�O�擢:	� ��JӁ��2�!Y�Vf"H�$+#��3�O�x*��J��<{$�{����:�4B���z*pMi���6UA��z�4�҉�O8��䟇gL*f�<>ܸ)Q�ԍ}�!�d� ����b�F5;���v/L!d1O8�>Q��L�O���'���\�A���RB.	2g�b�'$X���'|"7�8$3�'�'nE��џ+��3�����8Ǔdv��?Q�dL-f4p�j�;aR � Ma8���@�O��OfX*6��)4������ �V"OL��0�%'�|��g׽>b�avO�9n��M�t������0�Z1�91��c�p
tg���MK��?Y(���˂n�O�5����S�`�Xn� 'n�O��Ø&��D �|�'6�9��^ha�+��(�ԚN��˗�)��F��Pfj�#e\H�E&�<�r�'μ����?�H~H~��B�j���U�FKX���S̓�?�ϓ&;��Ч�9b�U"$DُT�N���:�HOz��0�Y0@�Lp�2S4"�Щ������џ��<I6h�[�n��p�	����iޑ�7u?Xr���.��|�Fy̓?�$��I-e�5��?"n6�����|�r�P� /<Ob)�P'^0w	�#4G�A�BB!7扊C�J���|I�,!��G�E>i�^�)`DY�y�gϫF����BW�	�J1�b�ϼ��$ZQ���$e�Ƨ��7kH�@�Z!wGԈ�$HN.;.�ɴ��O���O�����s���?��O�2�JJ2pnE��į�x)�t E�x�G��"�h��z�d�
p'R����'��w	S"I�r���/ �)a��ѷF]��?���)K\0I�		d&Ēhת-��)ޑ�խ6t��yS�]2a����<���s<moZ��	<?|*͐�~RN89�g:j1��ȟ�@�Dџ��	�|�g��%�܀�m&�U����Eq��L�p<��v��������T�5�te�veڙ�A�㉏Q���:����Tۜ�����h��Zl_	�!�$X�9� i�c����I1��=^�!�ć�Ur �*${d0��ٓedR�-�	U�Z�4�?�����Ȼnh>��S�PDfabā�
|����	ۍ �.�d�O���(�O�c��g~�l�F�r���͈�c��)س���I���#<�z�@@�B���쀢)�h�m{�� EW����28s�1��Û�u�̓ U�>�!�dCG�ɒŪ(E��õo�(l�axB�7ғC�Bj��,BmR�X�F	V�+Եi&��'W�c��jGr\;t�'R��'*�wLj���ޝ?t0��d ��h4����X�9�yҊ%k�,����M[C.�0���۸'P��9	�� ��Q�56�~m
�i�/�R@�y����?�}&���R悆s <���S"??�8��->D�Tr�G�&����`M2���U??r�)�'��p�ˈ/(�A5)��6V@��X��P��oٖ|̼i5�A�h���T��sa��?�J}�3�ˇ�&��ȓ�R[a�\so���p$�?p��ȓ?�*(R�m	�5�VQ�Oƻ.�ՄȓJ�Ĝ�u�+{��fŀ24܍�ȓ)Fe:���@��m���,ƕ��$��y��-��$mD�I�̈́�2�X<�ȓ4ڐa�3"Ť�t�w�T�:�ȅ�a1�9��djح��dW�y�$���p��@FyV2�H�fsKx�ȓ ZlmJb�>�f\�v���c�0!����1'�;��8 'R����O�^��W���DJ�X�3T��C�	1h�Z�y��K�8�qaFײcxB�AO捃�E@��4�맋iC�I��iBGN�|D$��π�F��B�ɫ6m�W��t��U��� ��B�ɾB � g]?�x�x�C�O��B�)� �ACg�X	^|d2���Ť<�C"O@�c1fC�s��s��ɸ-�Э*�"O��v)�DZ�q�E��$!�r���"O89�!S�* ��Ӈʝ�2���"O^x����vH��Qe,Ҩh�<JG"O�+���'�ذ%ޛ8cJ��"O0�)�iN�E�r�H�%O3"�T��T"O��[J�LL�Icn�$�v"O<9���(A|,���D+j�&-1�"O,�F$)1ڕ(m�.g^�9e"Op��>~���K�PT��k�"O�1�f��B�TȻ�I�F��3�"O�!���I�^̰wg�%1�B"O\�Cv75�<�+��XH��"O؉��j��i�jѓ�	�X-0"O|����<_7�Q�"�6�Zt�4"OzL�GERG]��ȡ�EY���h"O,qf��t9�D:����z1x�"OL!����"�ʘ9q��#O�^�'"OAc�2}��a��^8����#"O�Py&�OJ,tk��%� ��#"O�j���D���(4	K^@=k6"O~���-Fo┥sB�J%�&"O.L�+^9[���Kd��j��Y"O$��Y�[K���O�'H]b�"O����#q/�<2���d0����"O���8!�͑A�Ոw��"Op	��HT,tώ�r%���}anɑ�"OHcJ]7dܴ�&�y`Xt"O�9Sg��*~Lb=;p�0D�,����&{a�>%?�B���2,���b�r�6� Wn?D�C�I�m�-`�M�6T����N2F������<�*F4C�h�zRP�4���� _�<�$�k�����cޑ��Y����Oj0����M���ّ	 �^��`���E2����fa-\O>2�!��$�q℉��'A<x�Ύ4Mў-{��)G���K9>Eq�=2�x1Fĥ��'3N�Q�&��8���DȔ|c��F)^HL	��'�� L�u�S�O�(X���̬c���z#ϔ�k�����"O� �7k�<Y��h7kOl�K`T�D9V�ܮTa{��N2D�J$xc��(Rܜ��2�
���>����bt�6�Hi(�1R�?>��4�eH @!��(UrbT��B��h�!خ/	�Y%JO��H��s�ܪ=i\p�&&!L��6"On=�4��H֩ZV��2�N}�B"O�t�e��D��2IL�_	�e"O���A��8۱h�$	B}#"O����m��`{������E"O���g�+R��� �F�4`?LI��"O8]`��V \4��c�Ċ5�ؑ�"O�{��P�ؓ�Dҳbg�1s"O��	-$�Hd�֝Y�"O p���Ȫ.��`Q� Aa�]å"O�� ��R1xě3Ő5OT4�4"O@��F�ѫ�\:'�[�$�L�pg"O$� GZ�=�$-�s��0�@P"O�$���ېk�L���V��܌8R"OȨ�fU19^��FmӴ�� ��"O"�ɢ%K�)�󇊐;>Ψ��"O�P��B�7M� H�˙6X��R0"Oh*�G� ����#���T"O��P.�����k�6
@�Z"O�QT��:oZј�H=H��PB�"O��J5 !5�0кcg�$�B���"O� �-Pe�&;�H��6�ߏ�=0G"O��;�aK�-�,��R@&K��-�2"O�Y�H�#!�R�[2���,�'"O�`!�+�Y��,��j�"O�����T �+��j��"O��ƔP��e� ��3}WF�s"Od����X.�eQ���9
]pu"OlM��+Qy�!��^_�`�"Oh�{�']���[�B�3
�ź6"O4�ѣǓ/�$R�*�J��"O�E;3��ܑ	#i�~�=�1�'n����͸�N�h�)ҕB��g�cb���ȓ|������"L�����kc�E}B�N�|�0�F�O����E���	bXR2��pw����عU��6��\X6\��A�ލʐ�%�)�'x14�gO�n�\�B&%�*�L��s��V��j[<a�6΃!)�6	�O�X��m��0=9a��4�ꐀ`���}'J��@ˋc���b�nwBUSa@�)F3`{e��'-�J�qs"O4��bʀ)N"x#s�"y"�2w���Z �,�b�S�+��PF6��B��5m�B��\�����Ȏ-`����E�v�ɥA~|!sd�O隱Vc�O� q�҆Ҏ�HQ�r@W}�f��	�'F�tB�m��|
��ٝq�Ha�J% �&1x�ƢT��Y����C*?Cđ��iߙM���pa���ab@��Pv� ���<q >��/R]x�{⭱��Cp�F�x�a|��Q�8F���i	fe��o�|"%��ybZ��9ۘ��Q ��14
���F���O ��p�΄2�2Q`gc���aEy��G�E�TB5#�Ni*�k�4	�,� i���y�(4@���B�U4�H�f@8!
��[��������Fɔ��ULŕ,��P��늵�y�ǇF���Cg�&X�=�fE��~�o�>k���I 1։�L�	_X(;�ӋSBa}� [���Γ-F�uX��":"$za@Y%V��ͅ�7�f��RX�>I��h��|l�EyB��3�v�G�d��DA�Mك�K�g�l5��MR�y�$L�f���ȍ0
r�:��`\a�Dm�ɸ���R����Ա��l��,Ѱ,�@+�,�y�8F%:s^'�Y;�M����0>!�h�p�%pRoR;6��JV�x�<)�(ٷ;��[Rk��g�Ld��/�Z�<��Jٹ�����N�����C�!�y"kߑL���h�&U�Q�4DYQ��y�G���db'd��Kbu�DG��y⥙ Q9�4�ubЂ��H�/ĉ�y ��!.����DȤ���E���y���)_�T#��	�xb$E@/��	Z?!�EA-���z�wX��QB7i��ᣠC���L��66ީ��D�^�txz��ɝk�ɹ������Z��u���U~B�A�j�}�'E2(M+��.��<��E ��D!F�F���ǕǸA�a�-Z�r�x��n�r�z��)OH�i�ᙺ[��=)��įjV��#�|"�ŭn^�I�'jnd8��ԮY�v�2S)�j��ĸ�/Q�H�jCa@ saB��V
&����C�`%z2A"�����>X�ٴ�y�8O&��M� ��|RE�ǄE�ȐSSn��_��0tdMG�<��F�����Ξ25�J�z��ܮf.�"��n�	���';J��)U�]�~2 	4C���vG�LY.���BT��p?Q�àdP�Р�K�y�n�[q� 65A2١S��O�%��变UW
aQ,�=z��Ҥ�Ik&(����)W���&�u�>�b�R�P����v틜k���Rq�V���y�����	`Z���a�!��7I���'2��a�{��!��BV�Z�r�'5 ��`QV2��AA��};p� P�<�M?�h�`�3St4��NHl�p�c�-!D�����"NLt��ԅ� (Q��K����)��\'���U
<�O�t��t�$E*�)� �!�EYB	b�A��x%;�'I΁���D&nz��I���{F@ބ=�ᤃE��0#��Ā�dL��+Y0�X�>ɒB�@�.P��.�W/D@[��j�'�x��n.� {�N�u�8�ɔN��v�a� �5w$�;�L]8Jeo�A�����F�
���l�/�pIBb����8 �}�G
"3�%�r�D�6>����718$�H��6%��!vT��c�]=�ubt"O�� �T;c���S�U�\��}��>�5��d1P��`�xk_�r�(�Q?q���ʾV��PB�_�z$�pd-�O����Q�;������(<�36�Zk~������}�dW����w�|�![�+2�`��[0o�:`����O���Ew̓hݾ!A�U��"�r��	��
4dLJ%��,3�O<I�p�9T�<��*P !�c�Y�P��l����'��p�rd��D	���'���3�L�`J�+�@G�A�Ƚ��'�T\q���,���Q��_�s����I<a#j��oR�A���O���ɋ#U�<(���n�B�d��|J���a�V�����NX��r�I�;Vg��9�"O^��� ����D�O�>K��V"O���R��Q�t���"O����+*���T�r�vY�"O(�B!c
��}BT��9&�!h�"OX�÷D�vMʴ�$6|�D��W"O�� ��13���;��U�~J(�y`"O�lb���&��BId0�@�"O�x���I Q��X���;%�"O@C�
�n�B43f�ܬK��"O�S疤<��\��Έ+r�z�"O,y�鍈}o�(ʖN]�p, qc"O��X�m�*��K�-ٝZ J��"Ov��fa�!:�hi��l��
T$���y	t��%��K��Yid�����y�ϟ�x����P5���y�i�?X�\P`tfK�Hc�����y� � P�|���DΓ�\��2����y�LU(0�e��D??�@tH"%�?�y���P�.��!��+�.��$���yB�]+Q�����C�Uzr	
��ڸ�yBd�8����`�	�R� �U�-�y"�޻#�~%�u�L�K�� puQ��y2��[U���/M�oH�|�4���y�MW.'-�䘀�31&,�����y7g��+�L"�YS�Ǌ��y"aI�=ø�8�Ɛ
�0��e,���y��J\�H+WƏ.�$�
奄 �yb̌�b����Pp`$Ղԋߺ�y"�ޢ>1�U�ޭe�.`I��M��y�d�
[��3@n��%�8=�%�ˏ�ygY�z8�%�Q/$,��D[��y�e@� ��KUǒ,Ʉ�8pfݸ�yr*N�H��W'�*>���IR��y2���]pBu�j�":���D�y�k�-3�ܤ�S(B�!>��[�N�*�yBnZ1z`�YH���s�e9�a<�y�e_V�E��!��i�dƿ�yb$[�Q�ʭ�¢��R 3���y�!�f p�+��z��E�R9�y�c�|4����ێg%,īCN
�y�r�,#��:7��t�ahJ�y�I�CX��ȱ2��[�����y"��mXŊ���
x�,���(�*�yR�A={����0m�r��w%���y2��	�x\� J�k$�a�Ƅ��y�U��Դ���^�z�r|��yJK(<�ȕ����sTBu�^��y�m>t�A!�q2:�q��S0�y
� jЊԥ�uT0r�^�P�)1"O�p�F�!\d&hᅉ��7PT�Q"O��z�X�qzpH+j�y4ʝ!�"OF��v�˫@R��0)��V(����"Od��������2u*ЬRHlx��"O����ؓB4�BW�%,Ј"OD�T�.%\5�"��V����g"O"��e��0Q$}�l�bV���"O�d��J2T�M!�d�?�	c�"O�R�mv��Ś!䁤G�B\9"O�,s�I�3C�-���җJw�X7"O4ibI�"L36隄j�F�"x�""O���.V"^8h�'��`�P]j�"O>��QDR� ;֥Rf�<�}`�"O��C�b]�/8�`�1	�L��"O�x8�.@�Y���!�e��	(��w"O荱VoY#fP��FR.f�����"Ot@�oZ��d�F�~�Ɂ"O"� wB����O�'tux�"O���q&��1�պ a�7<����"O^�ەɒΛ5�?e\����;,OT�<y���5��82
��o�y�`p�<	�̂fLfr&A P�c�l�<�eMT_(]�2�E�Uٔ��*B�<�D�D*L����``4�}ږ�Tv�<�Cސ%�E�G��1*d2��f�<�hݨt�X�"��N�+BR��d�<��9q&e"�Nc*N��� �u�<��#�< a�裲l�w܄��G/�z�<���B��y�6AK �Z����DM�<iFO׸\�P�Po�0 ��m�mR�<AW�.{#���c�<�du�Zq'!�7Owи�qB�n����F��!�ć�M$
\P�
��v�!u�I�!�dG�G�Tu��V�u�� ���:*�!��U\8�Սm��8��-ݱ ���Dx9�g}B�>K�<��SgT�7����'���y�IH�^�� ��b�D�����U�v�(�$�O|�[G���&pƱ Ef[�Fo*��"O� �g,P��@"#�AD����"Of���j��x` ������g"OPi��k�>4�����r��Q�&"O��q7�Xl��+�C¼N��+ "OL�@'FS�Z�X��@˩�T""OY#/C2~�j}0�4n#0!ٳ"O���e�ݖ:���#�ĎMA�m+�"O��j�Ʌ ,Zfm���GH9��"Oxl�u���+�bEQ�k̞D��QZ��� lO�Y�
O�nZ
� 8<8m#�"Oz�A`
ڙ_�~���v'�\°"O�x²�T�#$0�#��(��i�"OZY�D%�bY��m��6)��"ON�Io�SJ~��"6b��y�"Op����`4��aG!x��3�"O,A1"�_ZRx��m	�^>�
�"On J�Q�^8�K�p\���"O���Q#QJ��k�	.��U�"O��ʆΟځ��j��X����*O�0���#,��0Y��w��K�'�Qsކ'���j�j���
�'��H�,L;e��MI�k�*i\h@
�'%r���� 1�L�-Y��S	�'Cv`��-�6O�Cd�Q�AW�$��'���+�D5t�C3/8�p����� &�ل�Ԑ)��C�Eۼ\�5�`"O���&O�Y��5+W�+� <��"O<Lx���wiZ��M/	9��b"O�ћ��	�0�f3��+!6Hʵ"O@u����:��#kY�~>�5"O(��2%l�1P0�H�F�:�[t"Ol�c�HX��]0
�}h�K"OD� DI1-�ru1�h��6����"O����?�.�)�K	���"O�1�4ʊOm��pԧ
5-����"Onl��%��d�d!�Z:Q�<c�"O6J��`���؆�׻�UH�"O��Sh�WHT�%Nн[DS�"OܥiG�^�V���HEZ1| r5h�"O�`��$ �n�����Y�*M�i!*O�*5m��f'��q��GT�0���':8���H� ca5��� 	b.QZ
�'�(�(v琧 &@�AA(X�� l�
�'���RV��A�t���y$��
�'p��UIȣVf������j^����'%�����7l����L'0\�Չ�'6�}��o�<��d�3k�/NA��'a҆G?9Q
���F��-T���� ���y��Yl�B:�ʔ��(�8�y��B
J_�� �*��e05��yb
��~uj��!?`I�*��y�$����z��87r������y�K��4�}(G&�mz�b����y�S )X�(#�F��aJ��y�/�w%�u��#H�G�T�;��ܯ�y"�\�Hh�=6�͘?�<RdŒ��y��،i���6MD���I�r���y"AFtO��4ùp�R���eW�y�������9T�U�\�������y��7��Q�C�U(�����yB�N`{�N��J� ec�-���y��pf	9$�I!;栰���*�ybO�o��=H#�ʐ-j,�s�$���y�%�dEɃD!9��*�#��y�+�60_n�,�)�ԚnT�yR�`���
3����-� �yB��I�pͣ4Ę��*�hX8�y�dD�ty�Y&�8 �U �♓�y2)�1B��#Y8^�<
�H"	�'Fj1fcQz�`�kW(J[Ƞ��'�b��'G@�w�z���>�����'RT�p5!�*����(	�dj�'	|	�4_��d�5aH% ���z�'��9{��)���P��F�/,�i��'Ɏ͒0F�:t��a/B'>���
�'n����J�0�a��I=0	�
�'�ބ�#��6�r!Fx��� 
�'H�1�p��)��P�k��$@@m�	�'vFTE��^�f�ۑ��N��`��' 2�C��7N�n�Xnއ@�Z���'t,�3�&�L�):���s���ȓ�pTa�-� @h��G6u����
����F�(�(�kw���'�6@��\HN��Յ(P�HC�N]\���#�JA�a�ơw�}⠂��3p�م�p������0X�jf߇fꬅ�kR�F�V�tR {�.�rf��ȓC�����|1��V�=h6�l�ȓ.�Pu��G�z����t	J@��S�? 6|k���'M��M��D�1"��"O�!�+�;4��u�3�� X��!ȶ"O�`�p.�g(0�a�@�"��ð"OJ�a,�Gn|��MX4��kv"O$�yA�1 �0���ڷ#|��B "O�5��\�@�Cr�ωmP����"O 5`���D����Bi�y�"Ovx;��?o��͉&cv���B"O�Y�B�X.ܹY�(��M��"O��µJ�(�9D�N�z-��"O|�
�mDRq 	�2Ol���a&"O�!�S�+>l1�tT��y	"O:q�v�%	#ut��S�$��"Ot��FQG�x��I;dw�px"O0���ؼ:ְRH�$[�p1�"Ozt�Ca��0��SQ��G�R	�"O�a��(��]�\����	A��$"O\YS�㝆=��M*���I��M��"O6��aق/��e��&��j`�b"O�yy�	�}" �1��H6&����C"Oj�8gk��QH��� 448ԸF"O�L�ؘ�$�2�]�=�����"O��pQF���!8Į�p���z�"O0��7Ѻ ��0����1y�"O�|ڡn�,�|�{&MY�	\I�"O"T郁��w�����"{^��b"O�Q�B7)
�-�≌�T�x�&"OXM���0RIP��(�̦�3"O���a&����:2��'m� ��"O\��A���p5�ЎK��%8P"OZU�%b��>qpM���Ż��B"O�ňc��Js�d��6�H��"O�a��ʦ'����K��J���"O���dm�r�  +]���,�y2���<�Q$E�2��)�	H�B�I�aV<}9᧟3�%r �&\�B�I>k��%9��ˠtR�)�@[��C�ɍ_��uA���;|�&����V^�C�I�������^0T�a�A�׈=^C�ɲ}��JC+�u
:\��,�.k�B�I_�0|1��
4�x�:�,~��B��4��1K7�*UGpA�G�J��C䉌ixdm�b�H=(���>��C�I�2P�4�rfļ3��m��d��_��C�&�V$xe���"�5B�q��C�ɂ ��9��*C�@HभΑ |@C�Ɋx�B��$A)�8��3�̭�C�	�0�=�Qdž
��m�B�:U��B�ɡ2�⼊@I@`���G��-;fC䉑_������ ~��샦���z�B�	� �+U��QV��#�jO�=�VB䉂.0�R�AN+=�p ��
��g�B�I�% .C'I�Xw�1�bJr�B�ɢ3������
��vjF���B�	� ����?o�<x���
J�<B�	c��@�#����Q�H�\��B�	�YD�S�	E	]�K��T6�B�s�b���Uת(s��G�XB�ɯh"04�ԮL�vA��/A�t̀e"O$���T�H�l��B�#~��)x�"O��R���9W
L}I��q2�"Ox�:���V��	�d�ՃMs�(3�"O>�����l����2kdԨ��"Op�� )M,���㏒�Eu��	�"O� $9&/����Y�`؁?l�!"V"O�%�΀?{� �C@Lv<�`h�"OZ�r�.#� &��	/1���"O�e�'I\�)��	pg8G�2A"Ot���|�lC�F�|{d��"O��@�É�Z\���p͍|S0�"O�I�q	��v�z�Dȅ;��l�a"O������8��!3r
��<��	��"O���2.�V�m��n�,1��*@"O��q��Tj����m�Lּ""O0P��un�䋑MO1��D�7"Oh�c&
4AY���7m��B�H�Aa"O y��H��Ht�&́�����"O���wj �ӊ�w���>�hEȡ*O���2DI�Qr�SbEZ����'E�<*w�F�0���0%H�ef�q�'ڦt�6�ˆo��(P�ZKLĸ
�'�H����z����7��LZ:Hz
�'|`���S7��y@�Ē�t?��	�'�:5
�(���ѣ��:�,`	�'��d��f���I#�Z� (��J�'�n���FM�M�@���-IE<�X	�',f�KP�Z�����mG�3& Q��'�p6�Oe;W�^'+T^!��'S~iz&Q�9,V�qv�
%�̜��'G`uYA�b�~�X(�g�8���'=p�{�ֹ��(�B���[����'�.eK�Ϟk�ph���I����
�'pܜ��ڭ
���X�`N�ҙp
�'�6�) �A�
f�B3��->�4��
�'x"Hs�K\�f m��j��Mtv�1
�'VD='�P�5�<� U�Sn��u	�'֨Q٦�U���*J��|mMޫ�y��V9�����s���vd�*�y2IX^=V�NSP����yB��(w���Bb*5?�$�{�	ʏ�y�I�+9��aÃ�ۚ1��xj�I�y2��/+��Ս�'��H� l�%�y��*Fhr�Pঘ�u �C I"�y���roaբO*s��1S�/�"�y�n��4��4x ��i�U��yr��	vR��*�3k�ܐ��&B:�y�N%�R%�0�X�a�0����y��8 n5��G2U�64��d��Py�ț�X�a@�=J%B�7^f�<)#�\�����Ӱ4�ô�NJ�<�x�ܵ�5l�74t�4�L�<Ap��%!�YW*�+t�Da�0�AK�<�vڇe��L��nR�|
b��D�<���J�T-�q�֤�$:F�aaFHF�<aQ��+"����d��86
��{�<Rឈx���a� ۭ3���D��<�"�F<���+\�(�.KD�<)s)�x�d��g��'M�̸�)T@�<1��Y�1�ީf��L0�g�~�<�\�ՒC��"yHл�!Ei�!�_�t�|Dp��[	��բ$/A��!��'��[�A@�Cfn� �@�l�!�d¤jg�����5Wy(�o]��!�X�y�ꡊ b�	@����M�I�!�X�1��+�3|0���͒�W�!�,+2��
�?�V��!�!�D�{��񱏋�L�S�w�!��3%��b�Ȍi�.�p�lC�!�� h��Im����,��x�Z�B"OduڑgӶHR=p�,]�U�v�ڃ"O���P,.<:L�ckN����b"O.�#S)Ӻ���C�����.��"O��R��.�U	�E��EcS"O���-�+V�ѥ&�����"O`��VC�!��p�e�q�Z +�"O�q`��[(��x���P��4a�"OnU��dӄRK����L�m��Ш�"OH1 ƌ���Ș���l��H�"O�3��]�z�v<@��>]"x2�"O��i��P�K:�i[���sB���a"O�" �6[�T���'(��"O`��3jY>[72	K��T�� �"O�%��&Ǒz&�� MRwV�x�"O��`�0BL�����2#�"OP�Y3Gڿ.4��*FkB}N4җ"O�jD��2HYvtjQ��5n!�"O~ ��Ô�M�2��㧓�hɱ"Ol�4
�.?�L� �а��$�"O�a��Q��Mau�G�42"�ˤ"O�QR�QU���9s��B5��"O&�� !Ǉb���k����u��P"OD�{���Y���A�;l�L��"O�Ys�T�uab�s��H�Wl���"Od`s��?'2��w@�/YΝ�q"Ob�D�*b��)j^��$��T"Od�`�g�\Ȣ�ѯ�L��"O�Ix4�[.Qr<���WzDe"O����BؿZ�8�C�YT~���"O޼!7� !L>Qҳ��/F�e��"OD�E�ț
�}zt�G��D�0"O���@�,���k�N��l �!�"O^���NXE)������s'"O�0�V���*�,{�#"0� H�"Of9B�*BE������d��"O����A 7F�� �"��)��"O�� Օ1���h�*�j�	!"O��!�K�5uU���"I�!�����"OHX�$M�luukpJĐ3���23"O���_D>0rF�� 5.����"O�AyъB2`���C�HYH�r��&"O=вD�P������\�!��<� "O.��ǁ�z͊f��i�@��u"O$�B�� Z��m�I�a����"O�<8a�:$�	��@��rĻ��'B1OB��h-�	+B�� �4����=LO�d��%��N��rȼ3j�`"O����[p�^I�4O����)��"OM4�BW���
I2��ش�|b�'(�("E�+��	G�N�STz���'��t���n�ER�"+O���
�'bT�Z�@N�ul0�B��s��u�
�'^)`��Р}������ /��
����эOT8ć��P�z� �<�!�Pa�@: ��U���L�����'���{ƩN`�:p{2g��F451�'��XZf\#eO"�KB䑵qWޝ�	�'�x�;V4� �ˠ/¦W#� J�'�6���S�7_���w�~w�08���#�V�X���z�ea��=I<�a"Oٚo�
G��0�5�C�4�"O�����&xT��iUE�Z ~UY�"O6���~S�ңDM�> ���"O� rtx�&�/l��ė�N����"Ol��v�J���j�Hܯ
�Us�"Oy�@J��a��=��)�*	�t�D��&LO֍0�U�|���pH\9h��,�fO�]�5�=��� 4OM��,���<����yV"ЯF'��K�D?M���ȓHM:l�7�Y-/Lp!IP�!��F{��O��D�T+S�A�֐+��J/$��'@�u�f��h��C5�@�'��e⢀�._<�K��W�P��(�"�)�ĭB�b}P8�˂h0*M��P��y�(�pd��V�g��(0��S��yB��n�"�XQ@
��|�R�ۅ��?��'�ND��K!#eh��b0,v����xE�P���Z�GI� ���R�׺�yr��u�2�y��Q�>eJ�����y���?��*yp�	H����ybB��m�U$J\���#E=��7�S�O�l��Ps8])��<�H`�ϓ�O��惆)@���Y�TG\3�'��Ć�tBQ�
�G��y0��J?!��ʛb�L`�7��==$wI"b!�DT7Pk�T#'g]5��KGa]5!�	�"������4?�=����0w!�$���ִ��+2q�4�%�?f�'ba|"��'z>�D�f�S�4F8P�(E���'��o�'��}K$�Q&������d�����"O��z���_���)G�!=R,��"O��1��TE����-$��"O�������i�럎w�B̃&"O �S�b_�G�,qkC��<ZƠ@�'"O,3rO:3G(���V���$#�S��C!8�:����bբ��"���!��5@�# �-���g��#���?�5G5����E'I8��G@��yb��T�|��:H�h��H�?�yBb��F�2i�Dɛ+JP����y2h���b��W/5 ��1�mA���D/�S�O�V��vEK�wJƘ�� B��	��'�fH�B�%E��b�ι<�^���'$��2�Cӑ{���qpcYCax��	�'��T)�۾n38|� )���q�r�)�t-��~ Y�hغ�"�`�'���A��X
x�Sw%��'��j�'�P}�5.]�A��8�ؚ%b�Y����'s�>��w��ͅ�N Pe@W̆�*5��$�. ��H�#�F8�L�CP!���_� ���!i�D�c�"��E!�$ˁ_V攒V���
��e���U:=!�׻%�PR@B�k�D�K���)!��-��A����G���ˤ�8/!�$�-R]�Lc�"�D"�D`#�H�W��}b��x�/�-�2�SbO�!<l%i��4D�4A��'dQ�iuL��G*��S�<!-Ox��dֿü���XP�c��]"^!�$�g
N,����m$�@�BlI��'Ka|B�)Xv���-H� ^�����U�y�I�!�����I�Tz��#̜��y��@� ��E= Q���&�hO���O4�`5FG�}8��.��Q����g"O|����Z�^]iUjh���\�$G{��IρGZ�M0U��!-�PU N���!����j�9�o[-;�<�(�+]�|�!��z���TL[l�DB�
�f�!�� �U�`c*��<���
0vT`S"O�}�2�?�4��@��	r"OHqP  �7D�n���)	�D=�d�'#ў"~BЍN�dD��B�
M#8��Oݟ�y�� 
����FA�^�bG�L�yB���G��	4H�!��|{��ʫ�y������0 T�s�Ï��yrMսb�&��b���4��y2��{|��ZǨ��F��(y����ybl�v4K�,v��c�.
,��xBY�Q\�I�,ތ�VXS�����e��(��S�K����{�M��	��"OZ�8B�O3�@B#Ֆ[�$"O��o1��0�`�*pH�2"O̜�&k�9��xh��	�`�ؑ"O��x����]t�h�FۉIŲL �"O��b�F�L0��%�� �䘧"O~0!���xL���O/����"Oܙx��K���=h��ݖ�bb!"Ot�c�l�E�|����{�H�f"OހPd�����1����6"O�܂6j��n�Q˘��t���"O*��TG�Wp�X;Tʆ��r'"O��ѽ+d�A���e�
�X�"Od�"ת�
:`��A���N�0_�(���5���Y��J�'�(��n1Y�C�	-ao&l���>;<�;A	�7[t�C�I�}��<�u��4s�AB�C	�jUhC�I�%�$a�Z�u�Z�f���FC�ɏN�a�jZ�u��Q�j��1� �O�⟈F�D��J�8���B�x���{�@��y��[�	�@�֏l}N�Z���y�#y[�$޽e����V�[,��>��O�i*��"so~H3L��=�$��"O
 pJ� � c�*C�W�`%�$"O|���BJ'S�6����A�.�0�"Ol���/e��qwd�O�I�"O�Ě��8y���S�W����g"OP(I��|.y����/ ��`��d#LOr��1�F�xt"����>��p��"O��ujB�"ϔEX��\Ze�P"OČJQF\�'�����W����"OjdԅF�8�ź$i�8yN�Qa"O�����U�>]�Q�"H�I�#"O�x��������M_�vA�0	��' �D�O�<�BT�jŒ�#�1_U!�� h
�zJ�#��т'�N�;e�'�ў�>��DlS�/����� S(X��Aǃ5D��#�یK���!'�5XV4p贪 D��1��*�^�#�oR>�LC�)D��8��
,~�y'g[W��iR�C&D�������"� F`��Xqb"D�4C��	 �A" X�aꮉ�!d ����2擘r˶��O�uxP-��m�3OH@C�	:�������iW�ߑB��C�!>xH ���	�5��;&( 9�B�	�66$iBrf	����rС"3ӼC�I#[4��j���f��'O!"UtB�K|�I�Z�bv�ى�D��8B�I:{ڀ5�cQ��$|8VLC�'�0B䉩�(Tc���l��IfJ�12�B�I4ψ��rT/ml��(�̂D�B�I��^���)_�F�]���ͺJ�B䉞A�`���#c���
��(�B�)� �e�F�4"��P�k��W��!"O�hC��^*`u��L�@ސ
�"Ov��T
�B����Î%!�y�Z����I�' �aç�}���#n��7�H��d�O��*Q��aǏ�G/2��3���征��'ݤ����ub��8�k� �YI�'��qS6���S|zٰD�B,t ���'%�*�M�î�2��ð]�(
�'�v�+�%P�e<�P؀m��V+����''t$��N!g� @%�@V��q,O��D1�)ʧ	o�]���%!��9��.�$��ȓn�`���T�t�,�9`��%�ȓF�����U3��d��S�Ą�?G��Sc.ïKC ����D5\b�ȓ(Fv�C�E�q~0�0���H�ʵ��/y�Ѣ"�E1 �0����^�E
6E���b���˱>�<0�v��QT����Xp���,�y�Sy�޹�ȓz�|`�5埋z�θ9��G|}���8��L�/ie�!+D�N c�!�ȓt�xg������"�H�.F��ȓRD!�p`�9> Ⱥ�#T;\�q�ȓRK��2�O�m�xe6T�E�ȓgm$M*�(ߝ|\HK� �3�@$����x�u���<��5ȇ��r��C�ɼ���"dF�>�XI�E퓭7|�B�I e{ʝ;@�1E�0�(��75��B�I�=�v4c��CI��ٳϝ�hPNC�I2d�>a&�\�Ay���F��C��'LFԽ�aOS#\G4	�M�1	?�B�I�F� ��P${�d���%aG:C�I�$M��X��U��5�DwC�0X���jҁ("2�u�c��x�NC�$s���c�'��4�v�9��M; �.C�C��/Q~��Q�o�y�.C��	M:Tkqń�:�`���JE��B�	7	;^�y���^a��W�1��C�	�3���A���1c��s3dT�FY~��0?�!�пv��5�D�A��4B7h�ox���'�b�S�$�f��Mi�G�(EvZ}R�'���5�˘ .�%�`�P;
�.r�'f�I�`��'��\�С-	Z���':�P���3<�`(U�Vl��0�'��)g]58Z��a�@4yc�= 	�'֘�J�⟀C���i&��q��H>ɏ�����|Ub���7Q̸� I�<��yB�	�sN�4�u�]�$�m�VF��,��C�I�
 6����?L$F�+6N@�=/nC�	�;N��0K�7�<m��.�'>C��
��д �?)�1��	�
C��M. �r�3�٠h�<(��B��d�f����	�~(�x�V�f.�ʓ�hOQ>%�q�Ѫ@:�0��kKl�	��/�<�ߓ�y"#�)_jТ�	R/X�^0�%����yBD�/�ay���-Q��	Z Aِ�y�Aܫv��E��dΕA們È��yR���A��+���<���� ��y�bփ,N��eR6ybQBw�E1�yb(2�N]ha�^�E�^�!w�A7��'�ў�Oh���fB���s�g J́��>��p��CO��-'F�s#�`��"OTljr��S��pզR�J*��j�"OD��A��'��IҷD �i��"OP�ҁB8Y3�tfN?n��)u"O� �Ak�������# ���ͪ1H�"O��↣P�xa!��]�l�#"O�@�Єیi0ꠓ�ʺ)��M��$>�S��<.d�Jde
/��J�I\ W�!�$���-��A+<�N�#�Ƙ5�!��h��a���fd�aht�Zs�!�P�S�1�a��������-�!�䎩;6��s! ˗2����ď�n}!�G:S��9�pn�{_.��fcE�t�!��YN��5��*�qnZ��A�">�!��AlpPQ��*e[�H���;�!��@�OܐQ5ǁ,gU�`�7�L�z�!�3T(�A?l���;iH�!��{B�az��3�K�bܗ!���pu�q�go.>Y��;$ g�!�Dɼw��y��0V;�t{�O0��OF�=��zp%#δ�(x�!P�f��0�"O�T�A��/;�(Q��-w���"Od ��EY0Z��E!�ᐁG�>0�6"O������>a�q+�=5䬹:�"O���	�OUX��J�'� X"O4�U
ξk�f�)T0����"O����m���-���	7er� ��' �ă�&�VL�N�.UJ����Hy���$�(�Q����Ert���S�@�B�	�3@"劐�܆[��B"l�T��C�I1/�0m���� "R4Ik��_5o_�C�I�K��E��' p��Vf
�Z�C�� ��oZL��-q'�:LpC�	1}ҝ	sL��=>B��L_a}C�	����iߒ+�]p��ە`��˓�?Y���i�Z�~�����a���G�2O��婍2m)�]���R�i�8�1"O1��e�,a�����8��U�#"O��X0�٠����m�#N��"O�����1��M!-ɜU�\�r!"OP�+@DӺM4.���@�.o.�"O��8���by��IB�u��jA�'���'/&]@�DHZ� I�J�1:`Й	�'�b�ǁܺ���XפR,x�I�'�����/!P�qbF�^�&F�;�'HD��1�,Jž�֫¬iZ����'���%�gޑs�h�K5����'>��B�O� !��$jM�K(-J�'KpA��D�#�$u:a
H+
�z�'Yf�y��I�2a������tLz
�'#�q�"�(�\qG�"}�x�`
�'��(t��J�xi�)��vЈ��'��ܘ�,����d�6xE�؁�'���[DT`�f��R��% na��'9�4��bυZ�,4��%!|!��'�T|�@���g	$�s��<G��-�
�'��r񅈣&N�V�tHes#-D���U�� A��YD�&jz
�@�+D���0 �,$��\;���;�*%jf�;D����z�>(h���)����8D�T�T����Pf��)c�j��7D��p�!��ubV��w��yy�|��.9ړ�0|r� ,ʔQ%H=!��E�j�<!`Β��p��l\��9��d�<)��F�b�Zك3f�31[��4Nw�C� �rr��o�T!N��B�I61��Uě���!+�~�B�ɴi��!9�F�d��##��;�LB�)� d=�����J'bH�dOG84'x`qP��N�4�g+���'�G�zH� $�����2(��藙E� ,2t�ݭ) QP�"O�E�F�`:�R��ϙ02�"O~�It��}IL����d�"��t"OPD�D��tF����^!tV� ��"O�ٲe����D�̹J&�ݱ'�'���A�����bL�RĆQ�@ؠN.hC�	(x�m@/X�w	Pm�t��p�ZC�ɖ	1��I��� A�u��	m�&C䉢X�4u:�L	A��t���V:s'C䉧�|���!u�`#�1bpC�	a�c��;�(��tc�~&��hOQ>� �$�S��&K�&��8��*>D�\�5B��&����O�v9[�>D� �$�D$�Ғ��
�i3�#<��0|R�΋A�@�PdA����8�w��m�<qV�ǽik�!�!
Q4l�ZH�u�<�bF\�|޼9+`N29:�`�B�[�<�G�A� �R����Ip�KY�<y�'��8k��	C��`�BAĢ�y�<��bP�)����bH'������L�<�K�H(ЌD���h�
��R�<�p��V�SWH��)�p�!#�P�<��m͋O�����e�4�6Ab��w�<����t�P �FeP�@p��!�Bt�<�����-�E���/����DFsy��)�'-�PP	���>>��c�s¤��ȓdx�` ͟;t{0HK�JB.5~�(���`Ł�j�qE��RA���i6��|��&�M�`H��F@�2��9�ȓPD�	p�L��2(`(��t\�d��/a�	�JB�"�v���,S'|�-��i�p3-٭8'�i�Ti�#+5���#�JD�(I� �1q�a��<��|��VL	�.�,���أ� �L�&���	�<Q�^�V�H[��Z	;�H:�G��<1���6zf�����'�А)clU�<�'�?l�4aRb%� I���6 �b�<�7�,*�� o�:HX\�*'�R\�<w
͊`���H�ϸ6:�g�Y����<���ipˁc�0?���@`�W�<I�%	A�d|Y7e*BU\����QS�<��ӇIбh�kF�Rˬ0�d$[f�<	S�Q��\��k��v����KAGy2�)�'1����bZ� t7��1Rr	��G&L �� I�I�l� ���`~���L�<P�i�-t2���A�2|�Y�?�,Ox"~���72(\A2G[�}���r�j�E�<Y��5O�n��v�S��
t�G�[�<i5�_�YH  8u�ޜU�܊�!_b�<���:-q�)�����8 X�j��^_�<QCK^6Q���`�S�|�:��a�<�� [?��;��6v�R�%R�<f[z��!�S#AO&.�:�ON�<Y�P<?�:G	�!���c�WB�<�C���!E�1[tL<I�t��2�NH�<�uhر3�ty	#ą�\q�L�p" F�<��D��!Px�&ʂ-�JkB�Wj�'�a��F�Zx���f)�dڠQ�K
��y�-ҵg�F�+��F�+H�P�
B��y��\62H$�!��OM�8�c�U���+�O�\@�D�5<tL&�V. R���"O"8[�)pa>a��S
i��!P�"O� ���$?=
t���	��"O�(S0�Q�u����O*e�x)��'e��b�)�	�4p�mZ6WX�|�d��
�����'���0�H�J�6ჹg���	�'_���ǡ �/�@,	�G��w.�@�	�'l�*�O_�K�P�!e!��j���		�'��y�R��^b ����jx&p��'F���;��q�3kZ)h2���'���3�K�i�@�s+��g��,�N>1����2xD��p�iG�wq�B$ƒ�0�!���2W�Z �bO�X�,�$E 8�!�D7���`Á�r/�u:���{��[�<%�"~���H�8���%�N��a.���y򭄜�,� ꉪU�n�p�1�yr��J�Pn%=C�aj��_��y�&Q�k=��'.�C��qV�����hOq�����)E<WHB�E-ͅ�l51�"O�(QQ�]'���,���:��"OV	X��L�q�tP��)��q��<�"O���&%P�d�V�3��9q�"Or����v��qٳ����,y%"ObpyֈQ�	���x@CҘ�P�	"O���'OJ�,�.y���Xl�Lx�"O����Р.�Z�Ө�$�~���"O��@Ƀ�tp2���I�P����`"OPa���ϩ�Zt�EIԽ|�*g"O,Hpt	��R���*���8*��%ZB"O�qs��c1��ɐ�*x�Υ"$"O�c0��7s��p��\E!.tjr"O$%�PdI���t��'�4#����'!�DJ�~� i����F`h�C��� !���'�r̓�$�M,\�x�N�4!�d�9?�HDKGØ=)PЪv��h�!�䌏1#��BB�"f�����e�!��R������{�r ���*J�!�dڹK�ȁ	��2/� ��P��-!!!��17�E9#l��[�
��!O�m!�$I{j�%���"|�Q���OR!�$D�P��m�p�J����#
�'y2�r5AD-B�j����Ӛ	�5�	�'��H0�������@>	�	�'�Z@�}�y@r��$Τ�	�';,(�ס�t꠪ D�t�R�RJ>i���i�C-���M CJ~H#��>!�D�7V��#'��
Q>�=!$`�>,!�!K�x��/ґA����m�!���z��௓r�LL��,� ��R8O��;��*
3�ѐw�՝9����"O|\��ۗ������(PE�6"O$@���>[(\��+�9*q"O���l��@��	��P\�L�i�"O�� �݊$�eS #�
8Ɲ�P"Ob��"�[�~��#��^p��"O����2Js�e�s"�:9(��'u�����1 ������D��&�� 1ړ�0<i�E���a�0
ʄ�K�g�<��W�8��|B����Z�b"(�y�<��j�`��&��E��Nr�<�S-x�Ӓ�6 ��U2@��p�<�%�F2���c&hY�P���Y���k�<��R1��q�%B�����d�O�<�V�4��0(�"XP}�vG H�<��!�v)"p{!��+*X!���G�<����
YQ�%h�L_�n�`��I@�<� ��7a՘�<��E��9)������'LO���[9%�p��oU�QBёd"O�5�')�:jV=	�Q�\�d�G"O�TCI�.	���cb���'^�I",�ش�LU�L=��dg�ej(�O<���P�-r�#l))*�cb��d�!�$�-8J�Q�f�(�iaw�i�!������&Q&�v|��'�*��O���$П9IC�⟨<��c�ǫ�!�1u,�}Z1���4G4#�!��-,�h�q�G�s�nX���R�!���,Q������*�rp�"j�2�)�(�V���G\�z����4l�P9D���'��ѹ��$PM=b�'�=�v��'-Π�s��?�T�vD� >�%��'��qq��.E�DH�ꏿ9{ZA�'�L�B��\�DxGă*d,���'���2��T�@���@̾)�d��'�DyZ�$J/ y��	�%Ֆ���D=�X���o��a{.�"�JLP,aj�"Oj=K�)�%5Z�]ۦ��=*6��"O�(�ևX��l�a	V�	�$���'�ў"~R+��.<���B�?? ��N[��y".�33n�<��ɞ3e$�dV�yb���+c6�)��"(�``�櫛��y2�O6��J�Ƅ���P�!��y"B������׊Էn�e5���y��Nf�[�;�=�AG��y�@B���(��%��u���Z:�yr�Ĥh ݺ���Ii��`��y�C��E�@,�W���d��y�$J
IƘ�D�߰L	^��p'®�yB��e�
��%�U�n�2T�q� �y��r������nE��ҷ�ּ�yr�C�Yn@,�D耺l |�X����y�	;�`�i�Ȋbd�|ȄHZ�Py��O� ����F�"�6�9�E�z�<�4��.n�p�'���C��5�mw�<�q��|dV��ef��c�(9ҁ@q�<�V7w�B�
萪S��8�C�w��l���O$P�+U�Tcz��"?�✚�'hd8s6d�"�4�����-���c�'Ox9C��j\�\�V��PǨh��'�0��q*��,@ƨ�Pj�6�Ѫ�'���p�F�P��} ń6�9A�'̘���T�T�E��E\�{�8
�'C��ML�2�9��#E"�J�����*��Ӏ0� abU*ٞC蘭R�ŇF�4Ćȓ:��d��MZ�r���wI��4��QpX�0�̓Z�LQ �/0��ȓ*�H��'҄;���[��6`���fm�$�e@ԏXP�|�f�ގz�(�ȓ �Z�+$f�w�T���V��܆ȓD�r�.i�d�&�J�KW1D����H]�It�B�Z��3D��Q���G�飐�Q�S�X��q'r�L��/&�S�O�]9�)���� Ù�H�P��'vj� Q�Ϙ��l1	
Ht$Uq�'�n��2�аAXx5ʓ�G}�P�	�';0"3�;/s��aT�T-Bo
�'����*��ּHd�0,��{
�'�x�8�/���q��M	7:�p
�'��h��S8X��`����8w�GR�4F{����Wl�5Ӵ�Ƶ �*�聦Yw!�� �XA2Ԍ&��bңP�V|�"s"O���dC
�X��̢c�	#h����'��Ƞ6�_�ı����/5���'���s�Kӊe���!�V�:}��'6��I�8�T���D�	I|A�
�'���E�L�Lʌ<�7�Ј|��a�
�'p���P �rCF-��E]3*S�(;�'� 4(�&݋�p51��2*9����')"���oôtN�VZ�mR��i0�!D���Añ5���q�ǽ�D�1� D��Ri6S#2�P0	�J�(eK��<�
�r}�8j�����Ʀ�$� 	�'�x��V �K&\|�G��*E7��!�'� � �K�#4Y^�Q��ҟEŶ k�'&}c!��$����G��54�x�'�����F�+q>�+��d���'�p��`�9h��MF`��	@�'vhD�Pc�/c��+�ٮR��#�'�,����5�@��EG�+ZJ���'y,#�!٨�м�U��U��!��'�4�B��;#�(��Ǘ�E��,Z�'�:-�rHHy-�� 7�
"@H�	�'���B��Opߨ(�j�MN�H
�'���BG���Of=��MU\�ؔ��'ZN K�AG�d#R� <? 5��'vr��E�/ZM�)�AS�8��0��'l�� $ �&,�b�B�֣-��	�
�'�|�s�e´H�P�Y�ǟ� �
�'�DaG,Ϲa*��J���I�a
�'I���c��&p��n  ��9�"O����6vvB�ZN�q˪MӅ"O�r����6��ڒΝ�p `r"O8�:p!S�;�#3@����{�"O �J���B�p�S�ψd�ZX�"O��rϵ~�ѧgՐ�:����'�ў"~���[���l��L ��!����y��U���rGHX!�'���y� S�L�P"f�-/Q�-b�^$�y� �mh��n�~�9�wk��y����ܢB��ٮ)עQ4�y2/�y�>)�c՜}npS]����It~2�^� ��J�e��-�y�kǦ�� �C�A�%�t�K��yR��A��-A�cY�>����y�)_��X�����2�ʓ��fC��U5i�C�W�Z�DKY�lC��2[s�����d)��T�
�<C��C4E��G��d["E�c����,C䉬Y�`I3#�KKPD"�ʐg��B�	�c�Z��G���8�$1�B��Tۜ�� L�H� Q"'
P�D�pC�	�+=I��S.� � q��Dg�B�I6v���S�7A씝x��(}�TB䉱('��x�E/<$�%ғDM��`B�I%>��@��� ���Z'�+I�B�I�-��M�����RWe��`��B�ɳo,z�1���Y���k�W�-�XB�I�vTҥbU�{��h�!�zRB䉀{���gc�"L�d�+D->B�I1o�d\!���{v��CC�X�""B�W��PӔAN9�"h:DB�ɩZp���ʀe^�u�&@_�(B�	��"Xp���<w���"�^�gY�B�	%1�8M�!��n5`��7��p�BB�)� �����x@�PB�i߬/춄8C"O��e�^�Zx��g�
}Ш"O0�#��Ŀ܊P��=hZYA2"O�АIU3cی��D4OcLUB'�'�ў"~���®j�<m���J���gV��y�J%	xA1�ė�H���T�y�G"��굨ɝE��I��i�&�yR��'w�i�੝�N���"2�D��y��Jqo^T�JCL�!9�$��y���� B���&��5�f�1-��y2��NV��[(c��� ��1�y� ��O��LS��F���"����y��Բ>�K��@���b�\��ȓB�N����#n	�)��d�o�B��O!����T0i�2�Y���15�4�ȓRMN��Pl8	�4iY�Uݪ��ȓlP�!���-M	����-\��g��t&Ϙ�F>�T��HP��ȓkx=E+�-�~I���<!fE��|3ndh�TG�@��S5�t؄ȓ#4X��U�׈7��=p�@Y=l�湄������ӳm�Y��hN%>e =��B�f�`�+H7\5"��I")�Y�ȓeg�
��?Oni*��B*ȴ�ȓY�*u�A��<�ii�ENJ��I��JO
`*"ŋ����Ke��*� A�ȓT�ċw��44���"'jE�؆�#�z��D�3F�D=�O��	����ȓǞY�!�++��M����(-8T��U���`� |\T׫V��V����YY��OI�QHgkD�W�ԅ�3xb�i� ɷNxX���ᝒtE����Kz�����_�K�9�\��*+D�LP&�B�_����s��3}j�	�)<D�$A7��k��e���|� 0�ab:D��r�� oӞ�jS�߲�؅�ǀ2D��֥�/\��q���K0A&D��Q�#	�(\Tx���	X&n�C�"D�H#ޒ1H�a��A�S(8�j�J3D���h��
�3�gV�}Z��=D���p��d��@�D��R���a��'D�bG!ӭ3�����`>�E��;D�ة�m�`i�88T��m� ;sB8D���٤M�"��3�ʎ-�d@��3D�xY���&����H�!+Yzq9��+D��+gG40H�@�$D�
֌���.<D��k�D��ġ[�D�f<衡O;D���珅(	�X�;p!��fT�܃�M:D�0 ���4�j�RW�]�?���2��;D��q��Γ6����"�Yr�ٰ�9D����1Tw��q�
 �%�d�4D�,0dIP
u�6��v](�Fܳ��1D��1BK�.(ޭ���Z$7�V1��B.D�d!���
�~P���+@t�=�B*D�T�rD�#%��=�a�fo��J(D���')Y)-¤��C�_5-�p����'D����C��+NBr􅝋[�d�&�;D�\�֫��#&c1�;Oz�e;D��)C���p$(IH�����5��N8D�t���t(�a׏Q��J�5D�[��_�gt�3�˟�n&��8D� ې�W���h�aEعO2$��(6D���.�	���H��I �3�?D���X*����"ȹ}4�)��a=D�� R�eAO�yi�Ũ�bҬu����"O�q�%�e����\�N��p"O�)!���w�qkV�ön&p2�"OȰQB�p`�A%i�\��hP"O��cnԓ9~�m��3���I "O	K�L������+�����"Oڙ�d��Z.���F =�֜�"O�s���N�V�K5 �HkD"O�ՂU�W�&�MYc#Fv�R��"O���C_�X�׀T)(�"O ���B�1M�x�b��.�0""O6T	 ��`q�1��M��6"O�m��,Yk�����*}�]��"Od<
�D�A�����"��X"�"O81�'�8FĊ�f� i��H "OR���蜭���þ! l�"O|�Hq�5]�A3'�ǒ�2��""Ox��K��, ^,�A���u�vU��"OH����N7E�fQz�t}�a��"O�%��
݀o����1ʞ(a�4}�S"OJ@z1M�Z�����&j���rs"O��hP	ƎV�b̪aH!:9J��"Oy�A�Y�l�E)T�Q��ȈQ"Ox�صٚn�q�	
�+�&�9�"O�e��./���QHL�h�t9��"O����0aPh@�HD0��"OЅ[ �ƨe&HC��
vB28#"O��scnN4_^��X1�G�tZ6|�"O��h��	u��h��eQiZ4�Ȑ"O~��a��xo�����ZnY���"O�!��Z� <��䑩8X��6"O�(���<�V��@V�-9��@�"OH@C � �@��%��oC�TNl��"O�Ũ�k�m�m�T�� xIx)�"O�iI2`�hZ��!C���LGj��#"O���ժk����d߆�9E"O��k�X
��3v�C�(t@E"OT� uk�*�T�1аcl�ȃ"ORE�c�H=L�x�#�e�{c��g"O���v��R� cUE�#�j@j�"O.ų�Ō�^E�����v�t�"O��:��ݫQ���U�۬U��"O��3���`����G,~�.,0c"O�kcC5���Ï	��1��"Ob�@�ꌃ)�reI�v��t�"Oำ�X�lC�����)@�r@"O !e���w�^)�B፟c�Yr�"O�����
H"(Q��2cD�+d"O,�a���B���,p��X&2L!�d�%'3:�)�Ⱦ�x��fm�;?!��U�Ai�u딮�y=��8s��_&!�䜚X\��A��]J2���*�$.�!�D]��9�[� �-�@*��j�!���0=B�A�핋U�dxo�. �!�҃g��q��D�P�mS���'�!��V���P��"�$vUk��B�G�!�^v6��6��> 1�(���!�H02$�9�3�Sd[�`�Pȋ	�!�d� ��s��J� $�R��%�!�$�4sd�%�!��%ɾu���	�!�ȿ`��	R�lV�,(Rɠ�լ�!��Y�/���I��G�7T��L��b�!�N�z���Ϋ;-
]Y�+��k�!�$�/�������C:�$ ���A�!�� Ě��3u������F���Z"OT�a�h�B"	��]���7"O$�S❕�R���-dse��"O������813R3R��Un�ac"O����$��4��P���(:�P�W"O�ig�1kLxz�*̕
��c"O�d#6�:���@H�.n��B4"O�5��MӮ^T4Y�F�6�>(p"O�X��]�ql�疶�0��w"OJY�BdƤ!��H6F͜GM84s�"Oy;���'tF �b�c�	OD��@#"O�yCf���n�R�V1TJ��"O �jR��+���3�fH�
&�"u"OM��љ<�v�Q�FΩ�m%"O�A7&��؄��юd��i+@"OFdy�IL�Y�0p�U7g,��"Oʬ����E+P���╊;��)D"O�gMY��� B�Fu�H��"O|�Q�C���+��^�H8���W"O��Ao�-D}�����~�a�"O>A+e@E�me��:�`T�'��1(�"O�e�R��Q���a�ƳzM�%Z�"O�I�Y�n��x�P�P3n\I�S"O�H����,�>�:T)��M|���"O�a�!��z��ŃvG�W|��7"O8�Hl�3�A{$!ךF�8)�"OY
r��&$\P`F�Y�x@s�"O����`�]��Dź"�T�"On�딆C�qjD���&�d���"OhكҍɱH��Z���,�[�"O��
q�'d��#Μ)���"O��Y5E�p�M��_?�t�x"O�0�Ł�5��]�Q���z�"O�Tc���gJ�
�+�x�1A"O�,7���o�Jƍ��\����"O�`QpJ�����q�¢~m��#@"O�ى cYzZđ�U��VTM �"O�d)r��C�^p��ĬI��n���D{���?*���R�BR����ף��K!�DͿH� ���̞Qd������=X�O��=��
$�g�_�W��AdD�����1"One��
_a����c�%��ݩT��4|OT<���o�漘Lå�������<Ey���T�x���*F��ΕArՎ �"��q�0D�$�$Y�\ѡЬH\f �y��.�0�d��(O���C�`��tk�G����	�A��y�l9M4i"`@ ���{�l����&�S�O��!ˇe[���@�"�� z�m�
ϓ�O�E�r"I�5��8���
�0�7"O���b	�BO��p��S�@,Z@�|�)��>����#�V�ZP��"A%[�C䉏p%j����D.�������+Jx�	]�'��SG�'e8D9��螵K���!����_�2������p��^?%�(�U�-I��T��o?��O8T���O�TÆ��a��"��P�FS��Z�"OZ�)e�#"���T ���|`�1V�\����V�x1#ŬX�F��&��C��?���D�uk����Jd�����c�<��cؔK1+�J�DF �U�״��Od#~:��*w�X񘇉	?��l���Fn�'�D�G�d���\�~\a���B�h	���&�y򤖔X��\����0w)B)بO��h�O۔�b�L)�L���#k��"�'�F0q���[d��׫�6\
���*�g�? <��_�me\��Bό� �Br�"O�J@,b$BdٓNL��M�D"Oؘ9MS�7i�P�͘h�4�S"O� 9�&V��c'̄���!�"O,xqC/�x��bJ� �^�("O�ٱ4I��-�|t9Di߈%���"O�Y)��S`�Y��E�V}�h{�"O��Q���{؆5
�eȤ*M�e��"O��1JU���P��	�5f7,0��"O��$璂^B|k댹��W"O�p��o��u��jN�(^�q3"O.Ys�B����U���MT���;"O��§�ܡ!�lR�"G2Ky^�#a"O�l�v�R�:1���Ͱwx�˶�'��$�H+�M��Z���q`��	9T�!�d���C�ж�:-(���.i!�d�2��,�����N�$�I!���:P!�dD7ȣ#�{�`+�J��pB!�$�35�p�ؕo/}�4�rɆ�
!��+'Uޕ3��ՠ"x���P�PO�1Ol���ѣF-:��MiTr����!�Q��h�ת��)��I��(;.�!��Bv�(���@%n�0Q�?m^��m{�O��bd���`+4q���b�ȩ
�'ъ���*)+�`0rN9ˀ�l*�Iz؞(!���(It�����ʁTrL��B+,Ob��n�����kO�}eh���-P#�B䉸/*)R�$�*�";Gk\�Z�pB�	v��pv��,[��"�N�pB�6x���K��>.W��jdd��r�&B�ɬ}w�m��U�P��}ä�]5cG&B�:<�[�^���:���P��C�I�mrFQY3J�<S��8r�C�	�Q� 0Aœa��xBu���"�MI>)�P!��#�d�*2�6�R�$�
~�̄�z���;*�65����dGg���ȓK�A�El¿V�<I���C�f̼��>�O�"���O���!hW�'��T�Į���	��'hҰ��Z21�j��`�R(zJ괈ծ�|?َ��S�o��:B @8wf���@�19����L���'�΄+�ę�S��f

�thN�h �'�ޜ�F��PA����"��!x�{�)�	\�'��aP��d�0�b���(�!򤈤 6v}����4`��"DI�"N0�D=ʓ96�}Z��::L�\��� "@��QXglF�<� �R�����T &���{�fP\}�"5�O0$��(R[&�B���R@P\�T�'P�Q����?�Ձ��`�Z�B�
������<X-hGy���'6L��)�z���C�c~���Ó�hOL���Հxl�|�2������OX����;���#�l̥tm���*n@����>9�E0?q�	�71� d��� ����"K�<���6?�d���˟�w��t�C�K�<Y7HFC�΍8�cѦ(�D%I�iI�<Ia�Q��X����)�b�s��ۦ����)��!!�Ȗy5��ǎ�.i?H4 ф+D�|��
�+S]2cJ[�j���<�Od�j̴RӃ��j��S�OŘ$�����ɀ1a�ɶ-?`���
L�%3�B˱$@�C�	&|���$K�kj�r�)F�x�^C�	"_�� 	S��88�j4X֩o�vC�I򟸈"HǾ�f��G�āEF2��ӆ���E{���M�W��)Z%��&@8�I)�!�&M줵��l��*U�A��]r!�� :�q�bפg�R ��Q�#\���'���T��R�#�� �!I
.C�I-�
�0�V}K�񻠬E	1b�=�
�']��,��(L>R���{W�\Wd�ȓg0ؽ���*ж4;��(�� l�"��'& "}�'���9���;�~�a���;vҔట'Wў"~�c��TX~ ��@F�ۨ8"�[w�<��,B_�Vm�b�V-��9�"-u8�&�d+S*@�b���3dӋ)Y2T{wA,D�`�Q �j��LB�.RR��iC@,D�4+3�ٚQj�}����1��Ы�,�OvO��SR�iO��iŏpʰ;U"OXQ��_���Y�_O 2���|�'��$:�'���@�����J�>)��-�J�c�>��zW��}�h�')ў"}"���1u�U��
�N�|�`�Np�<�e�5i���� ?��	p�Nn�<����o�VܡP�M'o����@��h�<�pn�	
0� b�"�@l3d$'T���4�u��T�Eg	�X�1��hO�S06*V���?Дt��*��K�'��[ ����!�Q & u�'n�4�O8�,x�B��q~~ͱ3FC&yШP�I�O�<ѓ	M�8�v���!�#�:�*vj��<	�j�A��(�r���Ǌ-O���uHܧ3��q���',�^���#��+d#0l�!)�14��U�ȓ#>\1Kf��!~af`sN��G���'�ў"}�G=Wq�$��._J�Mɦ��p�<t��gu&�sf��Vx����h�C�I}�'�>�a�(Z�C-@�9e��R��x��?D�D)�*ŠJ�m`"n۔M��E�7.<�	�^�Q�b>�"@�w���Ҵ#��'�ĥ��:LO�㟄��₩�� �q��bV�h�"�@��~��L<�倞1�hz��I1��a9wM�r�<qQI؄KΤdjVȺ�Ԅ�5�p�<Yd�:�&�f��H�B���I�n�<y���1z���p�"ʈ ���0��m�<IF�S
vi*u�r��b�̽2�@�Q�<q1�ݾH��уU �&���� L�<I�jFs>�1s�P�6�ۓ瘅��x(���h�'&O"4XDEҮ�y��[2��^�Nό��c���yrG��v�x��҄åJ�����˴�yB�0x5� ""Á�r\�IÃ܈�y2`�?9��laU��|�{ϙ.�y��	���T'ֹ���֋�y�ę}����͟
�l�JL>�y� Q�C��aR��ۑFb�c��y���j��(��N<�J�j[�y"O�qf౒�d27�$G�%�yB�I[] ��N�,ϔ)am'�yr(^,p����
�(\�a��y�cY�=h�U9����x�gC���yҡοhX�ق��e��T"����y�;G�z#�lQĄ���dE#�y��̗h����f��FX��*�䅳�y�L�(�����g5����N�y�j��$&���u�L�+��;t�Q��y�n�|�Pq�篝�(\F��`i��y2b
O3H��)n���`"D��yB,͉ba���}�ɛD	��y�AȆ5�a����q⣦��y���g:t�g��zLa��dǤ�yc�:+�\)��l1�=��-G6�y
� �ujP�6^Z�y�3�@<&��`B�"O�)a�I%�riY�kN8
��"O6ha	@�<b�����ЇK�VpR�"O��2!� �!c�s��U�!"O ���2O�|{��#[e��r"O*�ѐ�EiCDd��Ȝ�cnd w"O�xt��o�͋��ז;X e�E"O(-J��?{jI@Ro\7A����"O��P��&���
v�ttb"O����Y8	��ɛӫ�<-���"O�1��ʎ��pd�K7C��
�"O���U
RR�9�({� �6"O�	ɠ#�N���`����q2"O��3�Ɩ�3D�${��ؑ[��R"ON ����kO�H�c�Q?"�	G"Oi�7��!��릭�w��"Ofl�4BC�p�@A�!y
�X�R"Oh�"�c/|��"cd^8�����"OH�In����Ǧ2O�Rt�"OȸHt�ˬ2h��"Ն�y/!�"O�4����6 �P��$�PXpx"O�l�b��|Є;v\L��"O�� �2Ӻ��fhD<����"O��ْĈ�/����;# (��"O>�1�EOUd`�r#Æ9]*��P"O d���2,�K���=)d��"O !��k�*td�c�:�����"O�q��1>U�0z@�Z�J��s"O��7��mK̼�P/B=.��)Y�"O��X`&̏)��Q����y�.ȡ�"OP�%�("b�mrW�O�&쫴"O<�2��j�x�bRǂ�A��=2�"O"X�7��*9�\�����4]��"O��9�F:~�`��/�B)��"O
H���R����!B��!��5K�"O�iz���6ڰ�iaCC+1,b��B"OJ�x2m��Mk�	�r��6�B@�"O�%i��5����E���:���pE"O(�$	��?Te��Ըs��A�"OT(��k�zz�h�S�E�b웶"O��Ct�+F~�<�u)_5Ii&٠s"O|D�ACĎ_�5	b-{A��3�"Oz�9bB��Au�4[�-��^L	�`"O��p�ٹ`�8ɹ���MLp�p�"O�ܪU�@��Ȫd�قD+�X�"Oщ�n^�#z,B$bW�N"88��"O���ݣ4N,]R����JuJ!"Ov��5M�g`j}f�Q�(;�"Oܼj��k澰�t��GXT-�"Ol��҂J'0�U��N#5|N`H "O����m,<bJl��G�vmRp�"OةT�ğ<���!��7G���"OpDb �Kc��8�ɉE�R"O(��c�̪3������@<E07"O�2�#�!r"��R�@�.14�a�6�'���X��[41��v�Z)-�`|zbֽ~��L�t��y�,öp=��ȵ�E���1�M���O�RGLo�rTÉ�)��Cд�����2W�u:6��I�!�]�]���X�+ܮLI���f�0-�ܱ�5�V���ڄT��F��'���c���&K�"H�4�5�:Ea�'7�@�.�ɚ��G�8 ���*��8A��L2td�ӓ{i�qKW#C�qTr-�&H�jT���I�(f�Tˆ��~n�yKK����p�1��(S�L�<�uG-��zw�n���²@�@��P]�r�kO\&b�[��� t2��T�9��4���� ��TIt"On���$�4�j�0��;Qr�M��*E
�!��׏Q2�Iw��~���! P����:��:q,Z��y��J2�((��9���@��>�?1�Hg
���
@
�0=��h �a�ep���F89uE����=@!
PP:t�Q�d�0�G�m����͛M��4	�'w��V�M&W����hB�M^�Pz���KH*�X+�-@�(������	::�q##�~� �0T"O��3e���r~}Bv N42����]<Rdn@lV/��S��?����J�X���\�I��T����r�<�#�6�D�X��ۏ3���*��q�<)�LG>y>�HuEU�$��*d�Sh�<ypi3ވ�`#Sb����r�i�<�c�I�Q��Di��ddra��)H�<��T�4�%IG�U!Ϡa(e�D?�Pl�:�㞢}���)���3$��$��(��g�B�<9��N l`�)`�+�)�`i�&�y~�FW%5WN5���'��Q��L.��yS�*�.�ա��h87g�,z�r�i�@�>�}@�/� k�8R���Ɛx�*��W���HF�_�Ԥ�2�ʻ�O$\Y�m��p����G�'RЕ�i�+~:p�
!���k���f���h���;gb�����\�`�rFK		,��`� Ih�$4�g?QSCn�����	�Ps�d����]�<)BE�g�m��I��ؓmޟ,YfMQ�$��P$M?�ay��z����rA�!��jѮ��=" ������EE��y�\̢�b�'?$�#bC��P쬳Ќ%$�����O<�|�bB�[�~A����,�I<���1�KZ�rT������O8m��G�=b���G�Nm!��Ӎi8 �)7.��ԠrG^�bz4��F�Q�wt^����+u�q(�����M�I�Wy��w@S�.�P��U�����؞����>'VХ��A�mcܹ�ci"H���S�O�I�fF��<1Û����H�i��
��4����Q�'1�mkp.��G�R����H-�	!&��7�8����W��r�ϔ`�0��:_�8J�%54�����(�w��<��-���)���,E�(�[%EI-J-Ê�I�9d��-��i�%z
�[�!5!�ċ�d������.S��=o�#�cf,�=XR�u�܀�P��~�5�d��V��b����E��a��~�䘳(r�J����Fd�!�@cG�_��(��کQ8 q{&�>b���>\O� ��ڠ\<TY� BT�G��m���I� ��P�:� ѾvW8�R�È}�t��
�.�x3�:~$u�ȓI�$Pg�@3t�^�pf芩~sTU�J ���Ub�1@SH�����'B���d哿-$U���K�`s���C�R?R�C��86`D�F�p��P��KsU3i8t�0P�Ǫ(�E���x�4��OV��aü�&��+Į�2�o���j�L�x؟L ���*5�Y)�Jɢ4��r��ȁ;����a�� ��0Z��,�lZ��>ػR��S�'YX��!�G�g����jE�0��-�N>��*ţ1����(?N�(S��^�P��S�ּ�X���i�����H�T	����-~��H����=X�~dI�^&�H��O���cZ>Z�h�-.��'>^�`Ǎ�-��(KK'F���B�Dv�(��&�r���C��G�y@�/U��B��i<�}�`n�ZI� ���%LR��	������0�>�hB@�#V�u���[H1��a��Ե���tϳ0?<�{��0�x��S<8��԰Do�x~��)}f���
�&�$[�� /!�Ԭ�W��\�4A�i�؅ԟdGyJ�����B�O(���QF$׋���R7�ݳc̉/#��� 3��ň�?�bң%����ħ�	�� Q��Ȉ-%(:�(��Ky^����
`����ͤQ/҈P��ȭt ̱(�>�Փ�M�Om,�*Q�ŀSH|��!���b�^�ӄJ�"-�ph��k����--��= u�֦Z`�\��ޢ9���Biy�d�u&Ͷ�1��>�|����9n�T����*_f�%[�(m8��su.�n�l�������$X�PS��G�xtfqA�-�E"�P��>�¢[d����B3_p��`2ȧd#z (7ꋞ8��O�L�8 �T�?sX��	҃t� ���8/����k��.�"5�''΁-��[�j;>i[���� 2��q���e4-���3�ę�g
>9��fHY���2-��_~�Riȡ=���pa�	��-��U�d�!S�����q��+�<	5|	Cg�3���_��A������S�g�? T���+k���@b�t��ģ"O��V���B���qpaSj p��EAѺ��j"x����x�Ǎ�^�<��B)k��=�0Mҫ�Px�.c�&P8�;4�zvcXp��Y�� ۼ���I�A�����N��UVˤs�(�bN\�%#0	���u\~x�'���K��S)&Q2��A$��8�J!0,l#2B䉡F�,�1��3kRM#�Ěw8r��1�<���U6$A�ѡ�#ʧu<��3��X(� S7<��I"�2/\�B�	&�a{V���� ��mĩ#��9��]�e!��鐯�2�L�j")��&�mG|R����k��hZj�p�⏀հ<1�� վ�x�
��LT���u��5)��P(0�^UK��� ��917(�p�a~b��&43���cb�\���ڙ�ē6�n��ς40�@����cTb�0�l
P��3x3Dy�(���iw��B�In@���6h���n�9q��Y�!��K[!Gl �5'��Ywp���d��8��t̓?������ZO.������N��|��BV��ӧ�{L����T����BGG�<{���gDH;t�Bq� �ϩvq��٣�IiH(�xDCH�:�t�Q`��0�����D�G��I6�N�h���oʵ%⤣��HVRIx���I]�-�c�:Z�����8;8����P�	�\1t)�~�h�4��R��ӚU��H�'�`^B��4g@��B�9DL͎]�(��J�5�y"m�	0*0��R��+^;�5�V��G�L�hcbª,B����_mJ�!����|R�G�V��(i(U�_�^MR�H�xB�G.T�51��-ep�T�d��*9�Mjwّ4f�"��ȗI�"-���'�<,�b^82�9X!�VZj�Ó�ʽ�A� G�4���kV�h��
P�_2ue�1�WX������xBO=5hM@Ӏ5lB��7����@�nԤ,5���B?3b]1 S�4n@�q����3K��*��R�Q��da�'ݺ9�g���
i�a��X�䌑�rI�yo��� f�e��1k0)*�&8�G��]���\�PP I��o�,��ŉ0=v��&�e�����I�o,D���ːU~���B4��,Ǚd�����OD�asP�8�f�V� [X,\�4��7�LD|"��o�����Gٹ����@�����֟g��r������$(��i�����k.F��J�R��f�I�yH��,��#��P!���0?�E��?K����H�'֘�C�e��^���jO��G 
�k��I�7i<9�:(��Z�y�̃�w#��c��C�M`R���o�3ft8���_&���P)*{Ҡ��*J�+���*U�TK�����
�����̮U�FQ��*ѫ)~��'Z�쑊09O�\Iq�S*$\���F��us�)���ip%J���<AN�J& '�t�A�途�-kЫ7a�u���@qpoڱ �b@C`�g�']�i�����mgf�"Rb�<_:Ji�.O���Q
I�s�r�8M�֝�VFL���+�)Ӳ���a�#D.���G�L`G��Z��S
:��DB��z�a~r��Xl�B@��.xX��wB҄A���'^���W�E&�l9��0A��K�E�}�Z`�P8��@���(Ҽ�ȑd �D[�H���'��p���8]�� �M�.N�auf��FQ����Ȧ�h�e��N�Ĝ���>E�ԥ�
?��<1N4mo4�Z��]��0<!�e	ku�asK>��!��w�l�Ó��q���3���(�'���#3�{�g�)*0�3G�;$��7'P5I�2ЧO�,�7�� 긧�O�\\�	�8H���(��Ȋg��X��'��3 !� I?yx�&G=[l`p�'Ɛ���Ii� ��szhm�
�'���/�`��0�@fدu�L�	�'(������5�7�Jd��|�	�'�44�-Űx��j�A�^�R�'��t��c.H��"�u��a	�'v6��a�c6�Ab�ѥi���'�l�Q&��XE!1�Z�t���2�'�HC�	j�N��ЏE4n�=`�'��t���R�]���)�#V�-9�j�'fD��gd�%)[������8��'�z�ˇ�J���y('�Q�h�	�'���&�MK�feP�+�:c�ִ �'�Cb�ƫf�p�;��_&N�$��'F�A�@�eb�l0��:�zxR�'�� ��8z{���ʂ�7�����'A��+d�.!�ȭ�gl��r�s
�'m��X�@/"�,͸6�hͲE#
��� �,r��z��Y��V�<ń��"OF,
�� "6�b8�`˄ 5l��p�"OP�CܖM�hH���G^y�""O ��׻!*��5�E5fR�m��"O�Y �$�Nڸ���(P7$-d"OQ���e��L��"ۿh����"O�ٹӃ�wx�(ƀ�"Qc��t"OH���Ҵ'i�[2�A�%l�8�p"O٪�7R�C���
nL
D�"O|�h���!�� reo݁3+@)�"O��km���V�J஑B�ak"O(�+�h�r��X�C����W"OD��,��h"@!#ǉ
����g"Ox�J�d�
H�<]�t�G-o��4+"OhP��P�	�$��ƫ�i���P"O�B�̜�Cc����L	'�4h��"O�D����)�\(��o�B�YAs"OZ��p�C����U8�"O���¬�n�0}�E�� n��txt"O�|p�o� D�R�Y��=t�!{�"OH �Jع,��a�G�v{�)qw"O���B�\��E  S�x��"OЅj�F�<�5Ѱ�P�oM��h�"O��(aߔ9�� �'C9�L<�"O"KC�k4��@�L��"O��(K�yͪ)��F��S-�R"O`���錜P�"���F�6�^C�"Oh,�Ҁ\`�8-
r%ڠ�V\��"O����2B��nԚ8{��6"O��K���q�8u�K��RR�cg"O@Lم�JD��$]��4IV-Lc�<�6L޵d,�ɢ���5@6I�Y�<y��J1����G�]?�q���M~�<ٖ���U�b�qS��(Sn@��!�{�<����
$.P�1�nj��k���h�<��i�|t���9>��X��E�g�<ɗ���=(U[�N��G��G�`�<�G,T�2�]��'X7$��}��H�<B!��LG��Q���kA�E�c�s�<�n�h�}���v��Nb�<	c.ݭ��Ș��L�}�D���.\�<�GLU�{��za�T�L@JD���S�<��=T!xI2.@�lJ^u�pbp�<�Q�X�b�d��bĞ
0���ee�q�<��\�F �Kg���`W�	i��q�<���$D�"�g$�>d�j�b�PE�<����n�Z\f���
�l�B�<�h�?B4f���Ƙ	5HE�[C�<1A�P�d䃓i�3K���rk�x�<�����y���iU��"L3���$��y�<Vf�;D[*��u+�Rv. ��cw�<�r�J�@Fj�S��]������'HH�<!'�[�u&9p"�6 ��j���O�<Q��,v
�������*"gDC�<�6`Q�|��M� �9�əC�<�c��sN@����� %¸�fv�<$C�+�*41�aT&9�L��^l�<)��ɏz�d �Ŋ�s^~�djF`�<���`Z�*���5�NuhT��u8��*��с"԰}m �u��/��a�X`C�I8u���"C��:�w"͖}I\#<ђ��*r�B��d&��B�����z��v�.�wl`�<�GK�G��,��/*�"�$�
t�XC�	#3�*��'��>��,m՘i�ei/�x�s��(��C�)� ���T��/(Jd��Ȋ'N�dY���'�2��"��4^��`´�'j$$S�H0cQ�A�T�.L�X��	�I`^ĢD�)`*0�̚���3�%^�A���C�y"F�Y#8|[S��&��<HR Z���'K \[ѬW�RlЖᓺF�(TM�OjD�F#@J�LB䉰r��x�a��LrqߦV��l��Z9�tǰ<	���O��Q�E�T.N�(vB�,:���y�"O2X�h��g��1(#E�TA�'�^A9櫜�4�2(r��'���I���#�l�P�#�$a�x�ߓ?�T*VlZ���AE@R��(i\��i���b��k
�'�@!��
�4;3�E��*Rga�dB���N-ĕj�����(�Vx��o�p	\���	_4�aR"O� �qMnr���b�<Bҕ��N�%���f�y�)�矴��#�*}"��
�H�#{x�����,D�T�3{���d$E�/��l���.D��KU��aM�e�K��^	d ���+D���� �#_�"�1ש@�i	FPS�)D�؀�	�0k��6�¡wߌ؈D�$D�� t ["T%`GN�/��Y��n��d �j�;s�qO�>��PH�{�Y��d	�L�2G�%D��Ѣ���q��Q�� v���kÎ"?�"�C�"�3�*��4��N_�¸�hŧX���ԇ�I�c{:��#o�98HL����9%��zO�T6� �zH<I��Xqł�5i�0OU����m\}�'Ҽ����ӳ%�%�e+2��-Q�����9��m
�r|�C�I5���@3m�4Qt�E�@�=�%��a�V���+?��@���h��D��p#�a�%E�*9�SdU;;�!�$W�5�.`���6 ��`c�DYRm��^U�HS��Ƀ1,��Ib��A�7"ƶj!@L2���o�l��D�� �	��JGd��Mz1�֬t���@���Fe\�1�F����x��M7w�R��L�&�v�3ǃ��'`�d "���k亍╅p�'vM:9���$�������H6���KgZ0RG�S;>"n����,f���� sX*��S"�<�D�r6�Q��	=�'���{%�X{-�E���ST�	�7LE����}�eC`�Px ��Yqh�!���G��7 ,M�g�ݝ���C9*��H�'ˠ'�h�Q#�C�J/Q���� �'{�jb�6u6ؙ���9+ �*q�/I0b��'aPFYQ"O0�B���a�tYSl��+Z06�O|�T�J�g�@�H�1Sx��B�7ҧI�rM�᫆8/oF���ήn����~$��M?b\� �g"߲)�,��W��0[܊���ͳ~*���k�n��qO���"_!h���J�������'�x�"���#{�m��A��{E��31��mb[�[����P�T�>����(j�9yqD(В���P8P�Q�x�Ҧ��K`��!mY�N��ciP�)j8��F:U��8a5oE�0�
XS"O��ڵ䐻FI�5zp�:Tx3b�O�%z��P�vܱ�`[~�j�
h�c�O�BM��$K�DC���v (�f@P
�'���蟟Y�<�0Ƈ�(��iŮ_�	�����M�az��J�\W����?)����!��ŝ@�vlB���O�L,�P ���a��
9�L�3�ܼC�D-��m�f7�@R)L�@���ՑI�r=AV�iI.�aG��x�����L@*xBhZ3���K'�ݻ��'���J%�ճ�'V�b��ں'	D�}����WD� E����`�߀�u�Ԃ���8�X���� a;�O6���jȑ^��X@��D@�3��S���DB�+T"R(I��9�%�����Ď�@-�.��l�d�6HY(%e�D���"cz����6k�I�CK��9XdHBC�S�2��H�Æ�8��\���$4�4�ySj�';j�]�#�
��Om�U���msb�`�]�Y�Dٓ�E��p<�EB] q�r�"%>?��4W5���끇t��T�	$tiKc���h�Q�i�` ��O4��<I�J($gͳ�'6H-l��'x8}�B�?#��~zTŎ	7E�D+���Ѷ�@�7VJ����"{>�jA��k��h�D&��2�޼\�EӶ��2�L�1�O�$�"n
�XΟvU �͚5FO� Z�'�Qs5Y�lL��hqσ�V�B�2�'آ�2�� US�������^�(FO&W2<
E�Z�<1P��d���Y"e#}���雀d��B�$U=x�������p<q��]�Q���;�"?�6�ҙ.`���<�Xc&�ii<�ɠB&}F�9���I-�n�9% ��I퐌A���&i�8�'��5)���Nזu��3� :t9��VG�˧dZ�q�Hi�E����TXd�=�p>I��"E�ƅ�6LQ+��Ur��f�R�O�]3"aPI�I�S���Fd�>���G9*�,�B҅8d�B��h<!�O�Lhd�q�>t�Rx�B��l��������S��@�0lH<�}�u�1l�pࠕ�	:'�%H"i�h�<���G�n��(cv퍴/�8�KՋ؃�|�O:�k�+�B�g�	5(2%X��Â\��A�/W�C��� �+��s3@��,X��!��:1�vT '�'~��v�H����`&q����L,9t'����+�F	�a�j�FD���?�fن������$�/5��Q�����\0�Oi���P�38�p�'U�~E�R�rT��ym�
Jb��ȓCT}��"
�)�)��E��W&@	A�UG�D˵0�6p���L>��Πv&�I�1��_7jĸ��e(<���7psT�d,+�
t�g��9"2Uc���3.D���DE����/^�TưsE��rr�xbDҾ|cxY�N�}~��&v�Y�I�5�(B����y��B�v�hڣ ��Bz��x�HdF�2�o���𩃑4w�$�.E���k��W~!��;z`�h�n�6��!B{&�+H>I5�N�~���'����whA���#��Ζ�h�'��@Ô�"�x�g�z���kfE� 3HM��ɤ)?,ECp�M�!���F�B�I
��[��y��]�AQ$��B�����K�D�
����CS?��B�	�O�D���,S=6�F�aD�_B�I��9��IT��l0W�%��B��qgZ��#��2y��A���MFB�	'��4@R�7g�x�7� !t�C�ɲ?�LL&f��VX�u�I3~� ��$�xv>`JA�6�"�A�Vyan�����	���h�B��ҝU��y��M](�e�G�֨�y�	�6*�ޑ�P!f��Ӝ�n1�(�CJ�`g��&���Q�B|�8r�&�DK%^;D��'� $�J�EɀM�@�S��h��͗&8�'?�xs�'�e�N]zTK�2����g�<1UIѬ^0ƈB��>}��$L2:�(ճPEW"�j$��/���C4��?_d-�!�'�f��̀9C���#�ְ��mk�*&}�ǌ�e	ԙ���O`���Fq��r�P� ���=��	�w���bA#j��������3��XU-ԕ_>t!�ƩQW�1YsnN$S�Bj9`�I
TP�9��(����Ͳ���*d�Uy P���ɠ4�rt���QU�O�p��'A�\�|ۃb�B5<��@���$Of���3��dF'(�5��n��;`8�F%�zo��:w���P��"��Ş67f�"Ї�"]z@�	*����V�"U���Ҥ�0?�Q"n1 �� v���ba7|�8I� A�)E�0�~���=���p$�7�V`�'���X���"�3콃�c >��?��&���A�4���uC�&{~��Q�@	~7��P�d\�4oB���)�'i
Hj��[�gi�P�%&�Txt���	;�)c���o�]�pE��50� +����Wx
��M>!���Vz�>�O"@�U��%�>|�DA�"8��it�>�"�(GGr��?� ��v_��3�!�1V&���=D��B1�H;�!�M{���u(9D��x0��"'cԥ@��
3B`$6D�{��	}���8�(��?u��8D��Ie-�%8�tș���%���bl D� "N	7/���abn��ʞiA�-D� �v��1b~�E�ǁ(l�~yHd?D��C�<�Rd�ׅ�~8��:D�$���� ��� ��F��	��7D�\�r)B��9a�%ټwfyF>D��#Ξ��U�Ex���K��;D�Ch�LXp��Ҭlp0E8D���K֭��9���]jkT���9D�����>N�ȄY6Δ�`�^l��j1D�\y��N��1"x�$Dz� +D�� ��P���;k��:���=����"O�Y3$ɘG�<�I$h�f�����"O����[z8"UG@�	w1ɳ"O�=�I�Y��,Y�ǚ�(Q�)�"O����S�j��(Z%��7i�A�'"O��!��8Ĕ�{�@TaQ({�"OF)�a_�[L七n��,Y���t"O���BB �� ϝg�p�"OX� ��� �ji�Ł�C�P��R"O�@1
܍zu�h��%��#��@�*O�`"@�~��1�b!ƋL�.�
�'$Xl27��/.?821��1���	�'����A�~\��p��6�f�	�'d���N��E��liuK]?(�H5��'�F�RB%�7u����o��"��9	�'c���wFӗQ��jt䑖h�l#�'hx�Y�N�[�$�r�-�Y	�'��`�m�(/�:���IΚ�V���'�8$�������`Ā9{J8�Q�'����k��3��1�ܳ*()��'��@��&Y-E���L��p+�'�@ݒ0慴U.������3�B�r	�'/��Q�㉔�x�u$B�~����'>�y�%ѹ�d���Ѽ{��6"O���끬���˧E9ς��"O*���O�~��4��$/���"OL�Q�J \�xxQM���0w�/D��s��ʍU&Z��ub�%U�I&�(D�dZb�F*���Ѕ-Մ}7���k+D���
S�g˲�
���'l��t�D6D��: o�'20�ը�+�,("�5D���B��Y�- 7 �]��aUc4D�Ș��2Ab��M�Y�B��P%1D�X�wIR�6��U��bNV�>���d.�K�?}�7�	vI�i�e�M:AH��fa+ғZax!�	B��eڷ�#0I�q�a��ēFa�ɐ��?� r�H�t���'���8�0ʢ���Fط8�L��	 Q�'�uwR?]̓t��Ӓ�KZ~�Q	ۣ,CJ@'I�-�P��G.��9�S>�[%c�$|�`�x��x52Q{# 8U3�I�g/G(�I5W0 ���Ͷ9����Q����@R�R��h���P9�~��ΆB������=���d�$芳g�B���N�t���'�$���	�d�p��CP�����	B�@���n��x���:}.�ڶٓ-o���dc9D�z���=g�=`��	E�t@0�)D�D��ʝ-F�|���R	?q�M�3a)D�
����{_4�x��<w�Е�A�%D�z7)�&,��ŧ�~S�	%D����_e	��s��^��8`7D���͑7\-@E��|qӥD5D��T��
Lɶ���!I
!z��U�4D�(�7���b�\���H2R���s�2D�0�fN��)���#+��cL�Db6D�D��MG:!!Lmɳ$ʈBiR�;�3D��j��/
]���-M_xP�g�?D�P��%�1񖤨��Ҏ=� �PG=D�8��+U�If	*��и)V��3e�9D�H�Թx- �d���z��d6D����6lVͪ)�5b)�`�.D��;W痃AV����]�{�쥂�j,D��N_�9˺%�6�Z�s��5P�A?D�8�qo�T3nY��+j��e ��:D���+�j �в����Zڴe��n=D��)�ާsO`YX"��Ur�q��9D���@��X�8G�ؽg�Hs!�2D�� <��"��6g��ꃋ� :Q�$[�"Oe+@`V?�P�;���NJ	RS"O
��#�%Ru��1'Mζ<���D"O�Q5�ȴHy� ڂ�q%j��"O��r���1~mN5��+�� �<��"O�D�"�ϧ"&^���
�:p�ހ��"O�}Q4o[� ���y6)ΘĲ�r�"O<�:�K5+��;�&�R¦1c"O�(F*�(������}�h�R"Oƴ� 囌e6`%������@#"O0�2��_=$�YCߌ{�2���"O��񂒺3���8�g	����@"O|�P�A�?F�j�!$��I7�*""OA���.��d�ek�`/�+�"O,U� �і0p�A@6��:j�!�"Od%�FO#=눩��!��VP�Ұ"O8�e V8sH!���>"�T� �"O� �b'��'IL C��0(����4"O��[�V.uP�`���R/sH���"Oj��Ł4m��t�U�M'�D}1"OvY)�p����=�t}#s�m�<�C'
qd�$�!Z+&�����q�<�����\�TĀS	Y+E��ت�n�<����V��q[���;@6���GIl�<A�D6o=�4 ˗9�(����e�<���N�N�P|��cΝC��j�cK�<�$�G�A-�L���%E�����nGJ�<����peCC�O��Uh(�L�<闠�]w�d��nM�>�@���`�<�g#7 Q�y(�������C�_�<95F�0��q�G,�]p�I�e�<���J7X6����҉
6�@�M�<i��_�3���A2�+�Iq`k�F�<��9[Π�H�� =FQ)"Ζ�<y����s�l𠧭ø]�<yH�
�@�<�I��/�H�c�4�0`e�f�<9�d�g�`���0A�`QaD�d�<�s-S������@0L���3@-z�<�Ѓ�.J��ԃ�Eܮ7N�k �t�<��	�R�J��և�'���2�	n�<q�&cڠ$8��%_Ƹ(� Lj�<�І�M<���cÛ=g��˦Ĉd�<Y�1_��9q�G����eW�<aLS�z�vQ������S�<cJ�a���$,�Ţ�{-�V�<�3Õp�l��ʖ�PJ��:��k�<�E�m�9S��!��	;�.Ci�<)�%��bpD�i L��B��e�<AV���g\�@�C2�΀j!	�c�<���E'fi��YѨ
g�9 J�w�<��Ə"?�ŋu�BY<�};�s�<I�еR�< ���5�&\�u_q�<��n,P�
l[6��u������i�<��E��;��aQ���-g�V�Y�c�<yv�-|ͮTBb̞2b�!B�Gu�<�	�C��[��ƂOu���$Hz�<q�NQg9`��BĊ?e�2ࠐ�[t�<��.�,	2. `r�@�� lXI�<ᑊ�,��W��.0jȢ���o�<�f��|�c��Z�XfD,�rL\n�<��c��r�V-"��\(A#�%�t�Yq�<qB��&~|���㗸���Iq�]p�<�Vm��gn���4C."l	���a�<�V�]/HS:�c
˧O[�\�&TD�<� �!��¯'U�* i�$�L處"O"���(R�<���O�GHt�X�"O����E' }ؐhV��<x�.���"O��j���y|���ƚ9K�(t��"O����H�
#r��tKQ��} �"O�"M��u}@P�߽sq�t�U"O�X��"]Ɍ��GKfXp-c�"OzX��ޡf.T�3��B�A|�$"O(}�4�&J�pT&��CP�$g"O(81��_�\F���P�ʀ8�P�S"O��;3��$n���;t���R4"O����	:*�т���v�y�"O�����Zn'f����3o*8+�"OF=2iŮ�P�8�)�%hp$]P�"O��V'K~<�s(Y]�59�"O�q�K&$dX��fؑ%l�G"O�<�,n{@5��ֶ8���I$"OttY�BŠj��IQ�T~$��7"O(i��_��@�M��0jJ��"O�I�j��+��<�Q�O' Upв"O^�rBoC.�LB�
��4]9�"O�ջ�iE>dX@��:�t�q"O��y�����:vGҚn��t��"O��� jE�E�(����������"O��!�2}>n�b�ؗ&u0$x"On��S��QB�Ӥ)k�S2"O�y��ݣQU�YC��آ6�T��"O@�0j	�"A�aZCK��k.���"OfVͣ	ZA*R��%lPdHf`�`�<!��^�-).��T!F�3θ*�H `�<�t�Ԋ'��y�V&�=�\���E�<i��}X�]бl�RkN*c��}�<���ޙ@��X�� 	(�^Щ�d�Q�<�e�6!��]ఢQ�A��|���IP�<a*�	�|3��A�?�x����N�<�vON��^� k\qr�r/�G�<�ve̟1P��(ǋI����'�F�<yQN�!;{���!Շ&<$9Pf��B�<Q ��F��t�vR&���V|�<�CǛ�5�De�:��W��y�<�@���T��f�KyD�����w�<y �N&����&��)$��f��<Qu�I��ĸ�
�g�\Ae/~�<(8P~d����Q�l�"���v�<!��Ʈm80sR
��j$�e@r�<1"
�+hKm��}}`�p	h�<qU�Ժ�陳-Z�ܒM2Z�<�
ߎu�����@@+�0rD`�<� ��2n�yt��?,�4���BG�<I�o��b��� ���>���A�ƟE�<q ��N�l�']�d�.��5�C�<	�Z�"t�x �U�B�l���B�<�\?n#�A�g�?��4 ��{�<qt�E
f[�1�I���$)س��x�<I4�
�l�
���ō&Hz��J�<a�&޺پ��H��l����I�<�D�]|���C�/U� �+�!Op�<��(x��� H�*�d�j� w�<���$] z�H��g�w�ħv-��[C*���Ҷ< �Yx!C��_"P��ȓ>̕x�� �6ך�G��FR� ��X���*)G1 {RW�P{Nͅ�w��l �.�"�.l���kt�x��J�T�ʣĆ��8�%�	ĸ���S�? ���4�^w =����7i"��c"O�!��� �xzT#ΊYFd���"Op�𡋾;�ΠQ-Y	X��#�"O& �&�D�V\�Bcǽh9B���"O��!g�J�	��}�F��4o1���"OF$�4d��t���ģ	���"OL��ƲO���¬1����"O�QR�9X��5 ��T�E�6$`�"O�iÑV�:�X}��V([��IG"O�ݸ�N�)*^(�p�,̖$
�`�"OL4s�n
$��=��� t9�"O$�q���I�|�cS�ž%&u F"O��`M�05�Urr�M �#A"O4�`�ĽF����� Bt��&"O,=(�C˨l ˚#�<��"On)��̀���A�DF$��b�"OҴa��]�7�~Y�3"óԖ��G"O�K�G�)2`��·Iќ �'"Oʕ��Ā�$��$Ȇ�^�'Ԝ�2�"O�@�4��-(�����7t��K�"O�T;/B4V�}�W!�1GtD���"O,=�P�Z�G(�V O�=����"O�T�����x׬�/,�hh�"O��1T�-{ώ��,P�? Pa�"O6$���ݥz2���O$l� Mȷ"O�����Q%|��7�B6Mk�h��"O��HA<U�:Y�$��>W�	7"O8�:C"�C���j̳Q�YR"O�bG�ؿR'�)*�i�7:�dV"O��&#Ѡ=�j�=3���s"O��+2dؽB��e+G*ϯG��A"O��.
�4Lp�F�A.349�"O�`ca�R�A�VIs֧3����"O����h�	.q��:�� 3{�d�0"O����;.+���B� L�(��""O4%q��P<p4�2b��:����yro&C��d�g���Y�ּm!��)|�`{t���'Z�=����~�!򤝏H˼p �&�%S$�<`vOB,<�!�$ج6��0� ����j��Z�mz!��B�_��!J�BF�-��Cዙ1g!�ć,KG�IdI��`��0D*štf!򄞝r��M��AE2nЕq���%6!��P-d�r��K(ǞyK��\0�!�Y0 &���㚯o��5��;C|!��.��@1��8}�����%y!�D�K   �    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �P   �	    �  )  �&  #0  g6  �<  �B  BI  �O  �U  \  db  �h  �n  2u  v{  Ԃ   `� u�	����Zv)C�'ll\�0�Kz+�D��8��Mے��<�&E�H�aM���vo�^;NP)�A+.wȜ�2��O��h(6e
�:��1q ����u�cY)��te+I��TK7�<��`��cU��'� 	������ѻ�l軷��!8Ĭ0������]8��x��ߟ�k��� ��iHF�фY��x�ul��f�	JF�� �?Q"�S�&8h���Nś�gvq��'R�'D�`T<x����D� |cD&;a��'x@7͐����':�ӉD��d�'u���#5|� qn��N����DȦG?�(��o��Iɟ����?!��H,?���;7��a$�^�A$�ؓ~F���'�~��6���9̐e�2�_M굱�OH�A�9̄e	C`3�6�a��Μq���L�J���'f��'�B�'���'�������T8 '��"�ҵr��{g�T柄��4]�v	�R��'�26MKڦM�ߴ_����'� $��Œ�A)!K\c�فU�	� H�>�Ӻl��1%�W^7�{���wB*I�v��W�ʰ�e��C���lZ��M��i���x݁��aH'&�Ke�ő��h"ehXb:z�Y4O�ݟ�ɴ��(y�%��#]v��$��+pʈ�$GX8�M�S�i_.7�z�h-�q�	�hm���B���:�"7��=��	��Aۦ��ݴj���ET	C�*ccHGB��9��E]�y��9�ʛ+4Ǟui�`ѹX�5oO����Bs-�&q7R����۴buv��C	�3��i���C�H��b�J��}����W���6��p��&�G:OJ���%�����-ƨ
$��F�t+������r)��ɅUd�a�
j�lZ��M��i���O��x�&ۑnQv��'�'PR�k��ϥ%�z@8�F��(��"O��#��3x֝H�I�.�"OnEC���T��d��YqU�"O��$�I�=�rĨr/ϲ��  "O����$K�a����KT^�X�s�"OF�bU�N��܂%Eȸ	A�3���$.���~��,��XAc2H	���U�<�E���I8����N@�>�I���P�<ѱ�5
�ֈf"R���IM�<I�+�l!�$��t-�T���RE�<�QC;i+L�����Cwj$ZN\A�<��GM:fny�lQ�f\��у����X��)�S�O鐀��ޚl���B�/"�r�a1"O������*�Da㠣�E0�["O��2��Z3)`���ǳh�X�"O.m:��,,D���'�D?�(�iC"OX5�bb��aw��	5Fأ`נ0�'"Ov���ɇ�<:���E��.�2�Z�3m(�O�Z �Δ^�(���M�wI�L��"OƩ2��X-�������C�<؅"O���0l�+z�CE��\�ze��"O��r&�U���eL�u�P�E"O����f��4�$��^�`�'���q�*�Tf2�x��Q�F�d��	�Du�����d�O$���O^���
�u��T��=g��=��	����jH�� �C�����Ʌ�h�W!��w����	�O�łk�t| H�bëܰ	��'�RX���/{Ӻ�dW���vI6�B\�� �z�˓�?I���iÁ*�$4��̈1KY|�mh�)���Ĳs �4�B�M	P*���?+O�Ѐ"�O$�?���<��	��,�,
��kU*\Y��M~2��%�`��=E��(��)����A��+q�&����ɝ��Ă.f��y�{��i)T+�	�nA�1՞��׭�.����Sc���Oʓ��c>�xb�t�\�w���u��y	��7���O����q��(C�X��С�[�����\�O��0HDt�����D54���i��R� {.��?!F|!�z���&�wм�#��TQV�ӤX�Ze	Uq�1O���:���a���l:��HǟP�"r+O�d��f	:/_1�1O�؋�(�TS�2a�Q�m�~I:��'C�	�e۰�D(��O��$�O*y+*�@1<�3�Y�F1ht�׎)D���`%M�D3����(�0p����<���i>5��Hyҫ
;Z��T��>�h%aW꘩w��r�'�a|���\`���Й�� 6c OY�U��'�8"��և �l��4E��X��x�"և��ܫw���D!��éX@������x��I>c�
�d��?6hV」��y�C�D����D N��p�qB����1a�F�|���{e���?�t���\��M��zi@qW�?���D9"��?I�O̚�8"ə+E 9�"�Z�@�j��  ç

�1B��7�R�L1��Q��/���"�@Wd�y٠U��)��-�u��(��<;�	�(9�-cq�*�M��V8y2�2�ć7�"�'��I/K��T�'/N2$X�P�`L�O�8LOޅh���N%��!���p����r�'� �D��E $�pfk�6v�0IbD�[%�U�h�!͒ԟt��˟��Ol��S��'$�W��rD��
�˴!Eu�p�'�B兵	a`��B\�"H���VLH5 �'��	�UD�l�2�8����w�[/=�ɫ&���N.�2��4$dA�;H��@����=��֝*��d����*5	��dO=xGx�V;j����G���'C؈P�E�Q)<0��JKnM %*O�
���B,��獘+N- ���_`�O�)����\램���4��Ԃ�DR"��r��(OT$��%U9'f�g##rrŁ�"O�e���R(tC�q���Q	4x���'F3�c�-��c�w6`��'���d�$E
��r���p5J@P
�'�jɢ6�Y�Z�Z2���t@���' ����(�f��A��;��1Q-O^=`B�'%�mR�K���JYPa皧}��Ա�'v�� ���xshX�tSb9��'u�m	w�8)���R�ad%�ȓˈ�"r�
�
�"��N/L�=��������B%%��Mfz���I2����17��<8�F���$��&�K�C�?�
P��j�i�"dqg	?J�B�	?�V���N��� �(�:8C䉾Q.���H��G��y{���&$��B�;P��pFƛ'�T`��״V��B��2\>,LŊ��jp0젷▦/��=�E�Hp�O��Y�ˏbpR����C7d� ���'5d��b6*��]���)Nz���'N�U:e��kaƀ��gQ��+�'�M�Մ�/a����a�׎ O�a�	�'��  &�(k�\tz��J��� �	�'�Н�cF�* �`� Ù�x�	��@ɞ�Fx����I��0X$�V.4����C�C�	2.Ӝa��F�<5T�p�_	4�B�I�\A9��
`�]�t��M�B�	*qy���d�Z�P��� a6VB䉳�8�A�*@SR�H�:)`�C�	&t��T+(�7����,�R���I�]w��k!$*b��ɤ4B�c�rL#�\�%b6u:"���-�C䉗r�"���c�'X�@U��ZC�	�(�.�!q �P�6��1�R��B�	/)l�yG�:K�����@9�H����e��O�V��Y#�
��X�8��3/͇M!��.l�2р�@����a�0!�䑏m�$X�pi�*K��j�ڠi!�DL�A�����L�Q�Dd�F�   !�$�Yx.��g	�r5�
�mY�qD!�Ď�"��pL|���Ҳ�B+9ўK�D;�'L|\�5Z�""�1r��\�\�ȓƚ�3A�0XC6a���
6�~��!@b�Ĩw��a�`�oB"1��*ڴ��B�9�R���ɪh���ȓz�8�3�@�Lhֱ�fF�%o<���ȓ,�\]W@DI_B ۢWE���	*��#<E�t働�l)h��@=���銺f!�D��	U0��F���X�燞>T!��'|�l� @KP<%��`�a�E�*^!�$�?HT��̐!�����d۽6N!��$͚8��@J� �p�^�>!�D�7��"��7� �� �則 ���d��#{�`���Z�9�`�Cu!�66 !�� �a(�D�t�(��d��8[��0�"OFQQ2��%��3t��;��"Oy���
�� �A�A�Z���"O�@�@��,��=����B�h-���'q��h�'Cl�A��Q����&'Γ>�,<��'0h�@��L�Dz�ܫU��64�`3�'���Ў��u�h���і;1LS�'$��Dl��� $gC>�d�
�'�B)��*FRp����7L�l[
�'a���K��s�"��@��NƊe���ę'�Q?-�v!� s*�����Ȩ���!D���T(���ّ"�Z�
l���<D����I�����0����t�:D����#�	U|����K�l(�&�4D��6��$ȸ�:4���`DN ��	-D�ȢKM�X<8"���2>|���O*�r2�)�'5���7NIm�t8�D��V��s�'�6�R�M
?�*$X�$����'B0��O�f��q�΢4x��'wZ0��F<K����)H*�|�(�'���B�g���sC�߶�
�'�(�:A�7t��!�cC�Be��(O.�Pp�'n�ʥn�8H�v�b��3P�-��'�$�S$����BA��F����'�
�KCFT�
����1+RU��'t��X���<]4���aS.(�@Q)�'#�c�,V:�t1��N�$69�	�[������0��2-�lO��N��T���ȓtɼU�w��<&��<�BB�?�Nt��g��d�т������f�bNJ�ȓh�Dw�	@;�|ÑIU>~6v��ȓy��8�dK@օ��HP1fH���ȓe����Ʒ8��P6܌E{�F;¨�8)@���Iu��V�^.C`�Q�D"O�hE&ۯ`p�h�	�)c�i�"Ox�!E]�z���T�М+N���"O�����.J(֐�Έ6t=��i�"OI��Y.-JN��f�&<�y�"O� ��J̻77��#/\ -�.0�F�'U:A����*2��|�cEƲs��=��G>a��a��BغAҍיI�x2:d�8���?ስ�ոn~깹f�X�x!�ȓ6i�$ÙH�16�O/L@>���=�jM��."R��V��,T�$�ȓHbL9�!k\�Bn�����(7�Z%�'F��B
�	 ��a(�0L���w�L
;}VЅȓ���H�}ض,&B�8����oǏ WN4qf)D�Y�؄ȓ91�����[�h+��x��)˰���,M��Z�Li�5���P�bd����i��I�{G~��b�;It Ȣ�LV>ĘC�	�<{��i)s$�@ o��B^rC�ɀ]���K U!T�%�Ce(�6C䉱k���%�<k �=����)��B�	>+
vX6�+���j6��W�B��f����ކ+E�q׌#|\�=�F)]f�O����旬[Bv��CPϦ�q�'\��ݾP^���в9����'����h�,H���"&V�;�( ��'-��Z*c�|9 H�&b�LmH�'��1�AY�T��ؚr�G�.c�d�'��(qɗ�.[ �1iW�-����mh��Dx���Ą>���Xd�
�M�L�0
D< C�+?��5k �@�d�*rfǊm�C�)� �=��)F�0����Ѕˀ"O�!��	���!IA�&�d��"O,- �M�>�b@Q�!�Kڦ@;6"O�i"�E<J ��҃�V�cb��dX�|���0�Oj@i$���)� ��W[��("O`Y1���}h�i�dJ�6)2!"Ody��O:U	<e��$(0����"O�=�&��za1P�F2���"Oν�G��M�W"��U6��1�'��\�'�fm�'(�-:�ThS@�ك_���'��m�pJ�2%0��(x��iC�'��I�Q+M/Kt��WA�^n���'N�qB�l�
4BdY��kR5O�h1�'y�!�Q��!�x(W4?"�=h�'4�9ae=��Ȣ4�	-b�������29�Q?�IPf� r!j��$�y>�U[0c"D�(�2�W3���A��l�H�Q��5D�Lb�&1��y�����%�B9j�!�R
U�~q9C/Y��>	��cu!�жC*pҫ�V�,x��&�!�d΂(�0A�u��;g ~u �ʇ7��̋�O?��&�B�N�Rq��,V+cpD-�"�K�<��FX�_K�2���$�Z���D�l�< �L�D<b�0�'Юu��j�<�gB��F��Q����j���QF�P�<)b�{sL5�2
��8<��	P�W�<9��
# �p�5g�
n����Wy2�#�p>!��Wjj0���t� ��DDT�<�u���R�]�G��[Е�h�P�<��ʻvj	��J$.lhE-~C��0����K��8�˖H�M�B�ɩgX��"S~��s�G2FB�����9��3NP�(�L��]r���%",D!�D]�:X�(ր\�ii�ejaҟ>!�S�|S��"��7x�|!��NQ�_!򄐈S�Lт�D�5}.%H��"9M!���!��!V��ic�ő!m�32!��x2���ԩO/\b�kjէsў�; �!�'`��:ޡ�"ϣp#���Z�m�b�T�`���J�o����'��@&�QHX��cfݞTꠇȓY=������{���ѡ� Gi���ȓ=��w�ե%%F�v���@PΙ��z��&�Y0+-�A���<�B����}f"<E��j^�#X3��?R|�����]$RA!�"k��!�q�ʴKu��)S�b(!�9e��QNQJ��t�%��!�ѭSp�\��%�<z�Ԁ#��N�!��W�p,�6B�mj6���G�!��ʼ@�:�x��_	g��`��ޮR�I� چ�����M/��P!G�6�|�+����02!�ݟn1���7$Ϯ�ˠg��!�$� r��ђš{���p@G)K�!�$�(]��l�/7|�	���E�!�dGZA����Bip�n	�5��}��4�~�mZ}�܉�̓4���b�B_8�y��O�IµI#F^�w�>�����y¦�G�ܕ���8r$�H�,�y�D�7�B�c�I�p6�8�h���y2)M�d{\����@9�N�h�n��y��=L��� q̲.C�9CgΗ�hO<�I���$ʒu�s �9Y�q��L;>�NB�It
1����`�
��#�ShB��9�^�C�
�,Ij�hޔ�@C�)� �,�����J�k���=4�p��D"O�
V'��0�D<s�+�{��i�"On);FI���dY@@��� ٣��'k��0���%���C�MZ�5��]2�`�2����ȓm0�]a!�*v6���k���$���1G�W1Z���Y��<z38=��i㘨�����H�hV�J�x��ȓ
�fxsfP� .��@�e�N����*A�T�F��N�,����j�.9�'�ĄI�tV�A���M�xJnx��oL ��!��a�j�p� )�܃%��*�ц�b���0tCӝ?����4,��`��#ոI��O���kt�ߦ-�J�ȓF��	�4��>0��;�` IM�a��ɸ6�@��8 Ū�R�m�.R��b�	��NI�B�I'�2��"���*6B�	�8���H�������Yq��/,kB�I4wi�e%"��
BA�;#	�C�ɘK�=�mӖM�1�Tǐ+E�C䉡<Ƃ���D�
�P1��N�3�B�=��PN�ODY;b/
<d��l�@�/9B�'Z���n�LZ`u���I�r�	�'�j�������w�>�bp��'ӈ��r@�L��� Oĥ6�
�'$I8��QRT�97��2C�qJ�'�$�k$�֝y���M�0B�R ��9-� Fx���ѕ8v�A�lB>�9��(�s��B�	=eS>ʡ�?��#%��'��B�əV$	��[<'��i�u���]��B�	�q#t�&F�fN�`:$�DB�<D�����\�1��"p��>~��C��;5x��I�f[{�� ӥ�;�l��[��+}r�ϥBK��+}�&Q�U�������|ı�i X��ǟT�	��0˦l�U@x�	�+�A@VI���|b؄A^�]���";@�I�b�1؈O�8r�.F����D3���'f�H9P�DGf���2&�(�8TF|���?��ϘO��	R��*:�.=���XZ^��/O�������h� �5��#�L�O��}�%�<�g���;�l�B�+�=�����Xy��Ǣ4�r�'{�k�t�'z��C&s�r���7'�[�@X�	B)M�b3��rèƸkF��r�O?����Rq?vP[cM�0_� �Db��h�Dʮ�z��-M�g �\F�4�w�T��㡈�tD����y2)��?i�������\�$���cנ}��G���< d�.D�̩�	�4[�{D�GJ��Q��.�E��?��U�T"��uh�a�ѹ��O��'2,80T�z��$�O��d�<��l�]Ҡh�/|{]` ��rߒ���W��?Y��0x%�/�A���dB�5l:t�7��,7�lrֆN�� @�O�EQ���=w$q���?#<�D�F�%���疈�Ġ���]t~b�ϭ�?���?��2>�����3D � 7���F�tIK�"O*5�Rk�>E�*���N�q� �.���$��|�����$�Rf�X���N���z��;>��M���؇y�X�d�O����O����O���u>����2˦��ׂL?��8�aZbs��ف�X�ne ���ئ�B����|�*�&����0�∮w�B칇m�?�|����7F@6m�=�z����	q��zJ<!��	џ<���¦��=�Uڌh�ބj�֟�F{��I+���u���D	Fb�Z�B�	�kY�K�g\����Uo� ?�����'#�	/9h���*�$s>鰱�Ӿ4$q�ƈ��Jp����ON}�D��O(���Ǫ������G,��'{V�lZ����ύ ~�Y�$�F�Q�`��T�'��$�����Ԥӎ�:]~��S�	R��Έ2|�16n�<�܍��n[�%)�AM�	7#Kr�d�O�c>�I� Jт́�	�3����'�<
�G�.p��
��n���\�LXXh������D6prly"�#�P�����5�ɽ@d���	 (����Y���$:o���'By��[�T5bT�SOt>HF�'q9٦�ۊQ���Q���tD��!�~"��d'\��^�a��A�H��Б���'�y��Y�TƤ�ת
���B�aR;��@7�乪��B��i�u  �C�J��R�fl���*T=��;�2�'��)���Ot�)� `��6�Ɲ:�N%���?cz�MC�"O8<�XnFm	eW3g���7�	��ȟ�M���� w�R�r�Ã�DM&)[�+g�����O������I����O��D�O*��;�?qB�� 5�=�d��e�0HPM�
9��@3�#}�.!E3�$������T�d3ZQà���e�>A�6�T=`H�PgY+�f@��MS�H�Ju��S���i�����X����1���Z�,[6j�Ĉ F�g���7m�.���O���?�I�|rf-���^Y�sf�:C
��K�T�<YB�d�!�(wO�DT*]I��D�r�����'81O
LaW��p��q[�oE0���J�'z&���1���0r�� :xɂl.tI����`J\�@�F6P�F��T�[��*O� B�I�gB��c\-W80��'��i��N�P	��dF
��M�ȓ(��G��'���G�O�H8�Fb��r��*@+r:��\#�#�En�x���<WtX� �'HRt�'.B�'�Pв�&�?Uy��� �:9"2�h����FH�e�u�ΎX���V4��O�Q�0��<ТUyc�I+��z݁3��ϝOZ~���.�)Fp��QAS�7&PЧ%�W��'hL���?y�����)b�OR#;e�������$�O���$��~@�T�K� g��Q�G#ln�}��<i$�
.{j�����T�z���Ry�'=b�'Q���w掘3��D�1��E�6ɒ����y�'*��à��'z�6��dg�&N�����ɗ����O�0����#1ܬ�Ӫ��?r�@��ba�N�D�5�X牑h9����On���O�����t���(F���eN^�E�܅X���ꦥ���������<��Wnz�!�ʟk,ݦ*
��:g M'/?�<S�@K��m��?�򃏧�y��8�d�O��)�O��I6��%#�ϖ�g�&�x���'Y$�IK�O��ąA��db�,�/�?7��h��O�hZr,Q.D��d� &�#EC����'�=�	��4RD����	�OZ�������w���%
�W��L(� wT<��		_����Ozp0���O�I,S� �s���º+e��5W".����^*ft�U��d�U̓8V����dA��%���?!�'�N9��D!Q��բ�ˆ�0���@��y�n��?A����N�OF�I/j��s�`1C�n�&=�n�t�J�M�`����A	2�b`n��<e����M���i38�i̟��	�`�O��#�B��Wc^�yT,�r�����B��	�<Yׯ
ş��I�?����<���|R�Mڐ,=TuK�A�D���)��A��M��EF��?*O��d�O1���$_9@�E�
4=�;����BC�I��IJ��0���WgN�M듎?�/O�$&>��	]��Y� ��q��L%Q*��i#N�#=���T?�U-҃+#�5���Es��퀣k.D� �G�W	X�2�*7BN�5�i,D� ��
�~{����g�V�t���*D�l{��-�n �F�\:hx�'D�ȡ�ƀ�@{��Ce�F	:� ����2D����{�p,��ŔV��褩/D����G�Z�T9�(C�ah�u`8D�� A@�)R}���(N��i*A7D�\��ꍆP�YP� SY�؁�l4D�$ɅcO�G�̊�QVT�*�'3D���ū��w:z�c ��C<,�Zvd.D�@���Y�.:e��R�GD.Y�B�I9����0��K$���3@s�b�i�l�:�:���?X�@l��Պ�.�A�/ $*l�, ��҂~���1���i��H�d�:� ]��i:�������4n�A �ߘJ�6!�e��U� ���b��%��4#�^�IT�Y,����X�C$�9�bj֙N!b� !U�ELd��'哭��m ���oB����wӼ Q��Ξq�J�{��I�HʤHj��Kӟl�I>.�@�+�. 9Qtҧ�i�~b���iQfa�K�7�N�RD�T�ɂR ,Ms�m�;��?��� 5q8@�4 ����'�Ni ��'���'��4��¦��W��T�@���D@C���O���ǥu� 	���.�LMcd��~�x��/�a���ć�x�[1DG�ZwZ��'}��'�~1ӢJ��2��<�F�r��K�'�^�I ă.�ع+#��r�њ�'и1�pʜ�m��̺r �):=��'��5
`*�5�<���, C�!��'��&��*N�P�񭇁%BL���'����RA �F���]�$���1�'�f)���T�(��{pcӯ"td1��� �в��1RF�<Xo݁<��b"O�D;͕� $�5�d��m�`,Rg"O��'ޑLf�U"��K�`�p���"O���i�9�8[���BQ�l��"Or��F�(~�Q�Z�%7z=0"O�b䃘Bg��S�)
�H��M�"Ov]�!�U�9���s���Zt"O�i�/M!�F4�e��y�	�1"Ox	�Eo�F`Ւ�̒7hj��C"O.
0"�GDM�`%Fmp�z�"O�1�7�X�h��<��Y1b����"OF�v��+:0���#C�2�v�b�"OHaD��+�D�GIY@��!�5"Ox R�H!�Z�����5� 5[E"O��Z0CP;1ڢ�+�e
�k+�"O�<�`��o�4H���ޏp�
)bc"O��;4��X�6��d	3G}�䘡"OX(
��/�8A�(	�����"O�8����$) Ai�(E*�"9P�"O$M��*U�X\�B� �j��3"O�9� �O�!Ybܽ2�] �"O�50$	ʈwψp �@F�+ @� T"Ol����5G���o�P\�B"Oy!�/��Y�l��gϏe���ɒ"O��1���&51� 0��x��"O�l����-0�t<K"%A<F��eJ"O�a�u�F�/�!�$،)}�,R@"O��K��	�5-�H��"O���a�ߵ{�P���D��"O���Ҡ��e9t速J�e��"O�0�+މ��	q��6x ��Hq"O�`���'Sܚa����A����s"O.��W�����
���4����5"O��!&�&!'x��W���M}��s�"OtUБh��y��PX�aHs{`�x#"O����o����醔k��5��"Ob�B�dA	M��aH�Ѩ���"�"O��A�B�>nq���r��Y&"O0�s��+UA����7P���0g"ObqഉED�"�H���|�Z\u"O�`kA���Q�)��(�R�De��"Ov�)
q��5S�'܉(Ξ��"O$�����!�fTɒHZ�T��"O��	��ױ!������4x�j#"OREhԮB�tT�"#�X�f��Jg"O\�˷ ��.iV��CH*t��+r"OU*gƜ4�R��bg�t(h)�"O,,yB!܈b?����
����+\w�<9������GF�ub6����G�<Y����:���PĊݪo�I����F�<���E�OT��㡕(P<�SQ�\[�<1'�֑�)�B����r�XW�<�� Ed%j��ݡ,�:�d�K�<���-3�@"�JtR!�aH�K�<��K�m�8e���yŴt!C�KG�<ѳ�.-h�#��?W��!i���A�<�"ޗtu�|9�Ĝ g�hy�v�r�<a� #��M�"�P�0�� y0��y�<9p!�
 �a�w�у/v��Ppa�o�<�A�U�{��b�kO@��)2�Fu�<��I�W ��`���"	.�#���p�<Y�队iV)�BM��
��k�<!`��n���v�`>|Z�K�h�<Y"iD!OW2DB3^@���Y&iQo�<� ��Tďr8r� ��5��9��"O�9rb�R-�>�y�D�Xtʔ��"OҍU��)������Ϛ K���"OX!�KZ�|���C�";�Q�V"OnX��%�!x�z`"i�!�t"O�0���� |^u1�
�,��2�"Oz��R"����W%0XRuh��|�<�c��-c$0	����|�0s�Ua�<�1 �1	�P��q��7�(h�Gh�<iW�Q~���j�@�E��[B��`�<	���+0�JMD���1�|UpU-�_�<)�%P1F-R��Rx�A ��^�<	V�G�޲p�Mũq8d''QA�<!����R:�\�2���N�:tҠz�<av[�W"��wb"r՚�:�r�<���XF�ʩ{%'��j.��qv�p�<Ѥ)T0d��E+#�B<�����@�k�<a A%B��`�V ��F� 쀥��o�<q�I��ESB5Q�-ܪ��0��B�<Y��[-Ұ  %�]�G,j�
F�g�<�b�')�};j� =L*�Y�Ta�<��c�4y�Ƥ�����u�<��;9��\�g�?���	Q|�<a��z�V��tNC=D�]���z�</��#m ����z!��z�<��h� ?$�����6 9�p��j�A�<	���(�Z�"fS�2�T!ba��c�<q3釐E��I�/��DU��i�A�W�<i�Z��u6�3����!�$$��=��#Ȗ.ڈ���!��<?�b,���4��ݢ�+G&4�!�$��A��U�B;C�	3�h�!��W$	v<`�D��QV�W��#�!�$[5XߴXd��'$�6Iȉ܎C�	�A��x���W�^04�bKȌGoB�	��J���K-R*0��+D#B�ɸ[���A���XقƉY�C䉆q�.-Y�咗���s���2��C��c�40�u�X�Uu���̞���C��/Y!����k�.�hK�
;�B��  Кa�P?#�X��1ă,,dhB�`��i��j����ŐRn,B�7�|(�e��.�><��+�0Q*B�I�c>��8A���>価����	FwB�ɇ	�����ʔ(J�g⁊m}B䉴M2�My���uy,|zUE��DB�Y�\h��E���d"5iH�n��B��g� �Ae_�޾�Pw�Ġqn�B�	�	�2�ba,�	����G�/T�B�U<\pF��ln8Q�	&�lB�ɒ~�Ir��ҝ16�2�kR8#`PB�I=NS� 0�ʼG@�����n��B䉾a��됬K�,�����(m;�B䉾J�T�z���/?��;�g��fB�	�fJ����������Jh��"�4B�Ib�����G�'Y�t���W.H��B�ɇ>l�+��)����fԦ%	C��/d�]P��h"�=�LR�$��B�I�,5�� �-X���7�T�C��8AS.����	i�V���ũ4J�B�I���%*�BE�^6.� V�D�nW~B�I����1+T�f��V�C�(�LB��:Co�c�ǧa�qС��\��C�	�!�4)T�ߪ8>�M��Ǟ)shxC�)� �+�hF�u%���a��'pF�`�R"O,��am�}�z��TÁ�o'�41"O��G��7QP�R�M&'�tڣ"O>�����* e>�B%��x.��7"O���@�^QE�Q@��fp�! �"O�p�F���1��׃4Ɏ)�"O�x�Cřt���BG:v%���7"O�5�SM�����;2a�J��s`"Op(����Y��A:�����(�"Ofu�0*ܿN�Di��Y8	@E:�"O�0(F�$��Dۛ},h�"O*�!�X�8,քJQ�;L��Q4"ON���:$Up�c���~�P�"O�`��w�vD�MDv����"O�X�׬�7��l�c��)shx�2"ON�Th��:��	��LҬ��E"O����\�K?P�AT��
�t��`"O��`e
d1"򂈝40�F�*E"O�Q1��)��̲�!{�L0&"Of�z!��;gx���E�Du؍�"O����]o�& vHǽA��Գ"O���@%�)r���z��� �
Db�"O~qg�_9��@�ɓ1"y�H��"O���c�T��Rt)Ӝuո)Xw"O���/|��!f��)��`�W"O`��?12{�%��%�S"O��i�.E$��H{�����f�_^�<����R:L���±$V��K�h�Y�<i���t�<�F�
�]�4;� �[�<y�݋"���y��!Y�yA��DZ�<!��47�F���u/v�#�O�<Y��17��0W�\�5[vѠ�M�<Q�- \`$X����S� 8���c�<��A
,U����d�P�����N^�<�G��/x�
��t�0U&��d�X�<�S%-qt�!������aw�G_�<9TA���A��O(�����^�<��#�HZ�+c���-�X]��FCa�<�4�1=�̉�)��N~Н8��F�<1U�]�&��`��hQ 	��D�<�kATw"8B�c��^����z�<9D"�&'F�t�ug�:����ы�{�<A0B�-"����
��#�)��#�x�<)@iӹ&>.5hv摡1�6D�4��t�<����()$���)j���6cֈ�!�$t����'�W:����*a!��D,,>�)rDG	)�H�H���!�����
1D�' |h�i�睭#�!���܋� �`W��#u�!�d��6~X�
�t�� ���^�t�!��h�&� �
�"Ӭ��ƮA:+�!�$��;H�R��>d�bH�uB��!�RV�6ћQ��(ْ�X!D��!�J&��!���K� �������#�!�dq�	k"�K����{֯��v<!���"��9���&�����P�N!�	J's7�ȿ3�.��4�,`!���^1��s$���HV�0R�-^��!�I3JD�׌DU�I)�m�a�!�/JRPu��D?��KqkK�!�$ %o"�y� ��-�P)zs�#@�!�"�șL�&�*@cڤ&!���e��`B��"~Vt� h VF�lQT& Ĉ(��cM�/����$G����U�D�`�=B�L�>0�!�� �Ѱ��D�E,�����6�`�f"O& t~
�R�F��F�4 �R"O���������RRFD��%j1"Ov,�
�2R�xä�|ńC�"O&��1��q�V�(c-U=Z1J�S"O�%��N��Y�&L�X"F@g"O(U��*ȬSĒ#.B�lLaa"O��ۣ�NMcf�AЍ
�iWrk%"O�AA��0,�(1���WH�Ł@"O��fgZ����sq���:
��"OƽT���BSΑb7��#�A�S"O��9#o�22x�Ã��~��'"Oεc���6<�lf��.$m�X.x!�Gv-"٧�4�*�E�Y,!��)�`22�˼X�d�#
Oy!�DK�6�0˲b��:���c�T01l!�D�"h����(��ƈD�T_!��*�<��wƀ/p��q��OJw!�$��\��"㈀�;�,�!'m!�c�x�0�M�L��C"�� Z�!�Ѱ$2�y0�,���ؗ���!�΍OS�u#C	��UÚ��AC�n�!�d�3� 9�/�9)+n8@��|!���fz�d��Aˮ~�4sd��
|!��K�~y	�%I�T�֫z]!�$F X��9!�F��?;���Kۀ"�!�q6�8w��{'��cǊ�"�!��J�fH���SN4F�V��� �!���,�h4�K�;a�<�#g��!��4�~�i�U4=�p`@`��!!�Y����:��'Z-BІ�p!�D�fB�[CE���*���)
?!��{������wĜiC�
̕L!�$�2�T(r�L�`�
��"����!�dC)x�R51h�b�l%�T��W�!�$�Q���{׀)�^� �OS�!����a�n�
5�f���&�:@!�Dٍ E,�� GS�>%���3&{!��PI�	�����fy �y���MI!�D��w��I1�/!!	��Be��x�!�䋧OqΝ�6I�"sq��q�睐�!��4�`K�l�=Z�>���%B����8.Ѳ����
Qe�zG�T*�yF.-`�ĻN�?��u2wÞ��y�F��Ȩ��cAH9�%	wI��y⁃�y��i�K*p��ɫ�JJ��y���*[Pt���.�����(�y��ڵl���2'��G;�h٠-���y�GE�t`�e�J�l��m!/Ǒ�y�۲s�(q ��aw����nS�y�ux��S�������3���yR@W�\*b�����p�ś�L��y��	j )�s*�<xݜ�%���yF�2W��X���8pGn;�+���y"#� � 9S��:C�e�ԍÍ�y�.ڳw�0hp�b�Sa���y��ھp�B,�D��7�N5!� Թ�y2�ׇg%��(A�����%���yN� g���8guY���-�y2��<kV�j�,�!e�A��y�'5clZ|�V�L	w�б�o���y"�P</�,�HTi�"4�7iF�y3X���l�&=DN`�"(�y� �T�Ak"`��铅�y
� H��q·	ylH�!�� ��0��"O���1L%zgP���1�$���"O� ��D����3�hZ�'�PJ�"Oj5(�bW2(Y ��g	к1�*$��"O��B%�iBV��b��IH���6"OB�W��&�r�KΒ ��Y�F"O�i�� �r����s�щR�
��"O���vCJ�&�x�Ҕ0�x9C""O@P{��ٓ8�&��"/�x�����"O�����2���am�,�d9�R"O@l{���h�� ��
��v��Lq"O�ݱ����w$��3I�'yD:i��"O�=��M	�2&�`E���V�C"O:��0	sb0��i~S D�e"O4�ۄD�5�>5�'�Ob�ke"O�-�M͟r��÷�ˁs���a�"OxH+0ǅ81:!�@=D���T"OB�E��MXj���]�W_<4�"O�,Kbj�c�(��-N� ��G"O�\���H48~&�S3OT�� �"O�(a׀�0��x�`Άu��AA�"OjH9�ƀ�O*�@A�0 �zUb�"O�m`ȏb�*�R1ރ\>�50s"O����A4N��Ջ�h��"O�Ube�޶I^Q+Ł��$l�!�!"O(����"\�%�S炔3M2� �"O�X�6�]�"\�ZV�\�
dv-�@"OIx� �c�$+E		8���'"O��W�l��Rn��{�@�Q"Ox�1�Z=�X9��g�!�"O��&$X�X�lh�"� ~*N��"O�8f��;A�3��$r4�"O�(�sfS�Uz
���D\�c
�aZ0"O>�-Y8�óK��!N:� �kI�yB��U��۠��0dTh)�cy��hD���Y�5�vX��KԈm�,<�ʓ,�>���@�ےp�  ;>�C�2t�e��aT��j��Ϻ&u�C䉊Q�z����_ϲ�:sǚ!5��B�I�q���u��Rq�t(��+K��B�	�~��A�7�� ��Hؿ}J�C�	=-i4���i$�p�ss��QI�C�	�������7�<c�(�O,�C��2V�	��+_Kb��R��:I�BC�%��-Z�fI1"M.�s�G��C�I
=�`J �^�3b��#�OY/�4B�	k��	���?��yz��>�B�I�7t�c�S�x��@Њ�$�B�I"h�0�iVc���q����J� B�ɤ8�^�s�/�;�l�@cE4B�m��lJ6$ⲱ��@�c^��a�ĠC C�*i��+H6U�����c]����/�1v��br	��-����ȓJƄ9)�;W�x�z����IS��ȓ`H��AŅ�?����i�9��r�VM�1"\�PI���H� r�^���i2za+��S�h�0Sc�~��ՅȓI�e��	<T�3�@�3}�|�ȓh'^�Z���s�xɠAi"7T,܅ȓ6�d� 5�AM=�H��p7�t����-^B�,��`��cá
8t��`V������}'�9���[=J�Ѕ�ȓBe��l��y̰U�V��2ͅȓB�ZU3��H=V�T�X�c�N��S�? ���!�ϲf-�-���S�ڠ��#"O���'�)Z��= 6+�:l�v�F"O2u�U++P��j	�hŮ��"Op\1l�N��}�B�
~R�"O 1��뚀E�ĸ8�N������ "O�d��ip�@�%m�6�U�"O�� ��%B���Q��0i?څ"�"OX����ڐc.��X4-�G2� �"O��t�L��Z�lٗ{�q��',-"� ݃b9���ΎX^p��'Dl8� �ݍ2C�lJ�������'�:����ֲf�B��E��<��գ�'����Q�3�F!U��;����'�j�)���6�<�"_"��@��'q!Bg��?|��d��U��H#�'���@�O��v�cD���R,�'�Z�"��|_.��7�PLjb�
�'��`-��Y���KgM�Aiji�'}��:@̊6+.(�f�L�
댼B�')pH�s&�$/-�DI@1
�Ԭ��'a ��`�I�}����A�J���
�'t���eE�:1�$\+TR0CK�k
�'�:p;�G�j��D� #��{���	�'w�qb��2D�^���΂\���
�'�b��UGcƭB�FӕN_4���'Y
4Ċ;S9l��BI�B�8P
�'�z�c���� yb��ҕf$Rl
�'�x�
0L9U[X M��Hx80�'%r=�u��!_S�@�3((T���#�'�^�y�
#}*�Ȁ�Ix%D%�'�*PJ &��-�c@fݠ0�'m@�#p7�b�R�ѐb"�@@�'�\K�#��2�.�	��V�`���	�'I���ܪe�4I)Ҥ��h�	�'"r��b�?Vr*�rE��bY�a�'���#v���j��qe���	�'T��(eٵc����`�+ҘP#�'T.ٷ�&�4i���\�2 :�'�ژ(��Y"^H T�0Y���
�'���: ��
6���XAS�;���
�'�j(�T/L!и�pH�	D� ���'q8�'��N�RP��� {���)�'�$� �Oӷ�U�&�}��i�o9D�dq� �N	�p�� �����,D�	��E�o����a�/?���U�)D�����
I�bm����9�����G$D��i�l������:~���
0D���gJ��􃗣�.Y<� uh>D�d�7�J
M��!ѯ�8T5��'D���P-U
���"�R��.���8D�P�d΂ 0i�lY��Q�1��m��"3D�@i�Ȅ����2����+!M��'?D��8E���Du�(�Q�K�0](G�/D��x5��@x~P�F͟&�@��K-D��A@�&�0l�ANV3g?�C!D�  FOY�M�F�ӥ��r@��S�/D��QUE��U���C��_�=f(rN(D���aK�G�n�9�=4Hє`6D�0��G,(n����g�����T�!�$ٿ	�H{&���16B�kA�!S�!�D��l��Q�cĭlxT0W�H;�!����%��BV�<x-X�� s:!�$Ŝ>����60�}p��V�XY!�N�O8@Kc#>)���c�I)�!�� N= �ϟ+�i���� Rr���p"O�Z��D�{�n��U�	�?�VH�"O�	�r(q�>�[�&�?Pv��1Ǔ��2�u�K�.���a?<O��8�(M�4�`�4�R([�p`9d"OvpӉ���csk\>�~(S!"O������,D�tЄ�W�;����u"OFQ)wL�&Iz�TpJF/G�f��q"O� !&D�Fl�uK��o��-��"OXؘc�EH,hᑢ�46~H�8A"O�d#f�P�F��tzGJ:N,	�c"O8���O�#cp�!��鎧��T�S"O�d3'A��8&\�� z�AT"O
T�/��B<p��&Ƒ+H�T�c"O�!*�-�px�13U >�0]�F"O }�5!����Z�xLܛD"O��b��*I��DK��>R�JAc�"O�I�V��e�l��"P5|`���"O$��7ûg���Iw@��t���"Oh쓀EV�I� &	�d����"O�)s/��h�*��$'���"Oi�0B��gh (VD������T"O �A��A�����M!};4�1�"O��@��sx�����Ի=?���%"O�Z����llZ ���%j�jW"O�!���X�$�(C�L�D{J(:�"O�Q�h�$��+�� _r�up"O�QK��RGj�|�N��uZL��"O���6�چB9�A�f�y@�I#�"O6Y� ײh���uhXYB%��"O]�"fY�C�����EB�AA���"O�!���(�X�2"�,�9��"OԤz�f�>M�`���P�ML]R"O���J�IuЈ��!�>�+k�<��Q�4P 3��� c��i�P|�<�V �Uu-<�Д��C�<���L�pq��s�gC�� Y��C�i�<�v��e�����E�q�D�J��c�<!@�Oh���P�#�4G����G�e�<!5�٬0�4�v�Y50~���!�l�<�!���|� �&̊m����F��]�<�c��S6��+c��.,�4�����<�(��0$R����*:�Ν�PGe�<�@\!CVIѣZJ��8�+IV�<�F���y	$-�F�]�A���(�Y�<�v.�+\gFhs�I~lJ-���T�<i�-�Y��K���]����Td�v�<I���>
�����~fP���L|�<	c���2I��^R3lѰ���n�<	�a�Q,��c��|� �0Əh�<�4��&�$�h�H�(J�:\�u-V~�<������`q"f��?�����Ky�<�ƃZ�=���/ľta�ѡ ��v�<�Ǭ 5?ؼr'�B?��IЇH�<��$�~�l�i��0>p0J5g�k�<��b\��	���,	�bt�!�Dd�<���CvJ���
��-���p�J�<�&�T�;N�q� Z3�
ɨ媙a�<Q�
�h��yxv%r��h�+�^�<�Q��M/P���j�.S�<��	^H�i�v��//,�:��L�<�j�6h���;Dh�JRfhR���p�<�ա]�}] �2��
��|d
�d�<Ya��4~�N�*p	P�`E:���N\�<��Y� �d��ܐ�Y�r�Z�<� �!KCIŉx��Ťߺ;Q�9"O�1j����xdIӄ[�� "O��g�<aPm[V�0r���W"Oj8�EN�3PЍ÷����`���"O5��
�_Z�d*1&��}뒑��"O&�ڄ)�\Q�7��4t|Q"O� :�M&ޘsi	�Nh�!�3"O�(�"W~�=v&ؗL��+�"O�T�U˝*{�[�%��?"2��"O.%�W@�0=��-9�$��!�Ƞ�"Or��0�U����ɞ�t����"O�@�W�)L-����	��i�����"O�X�G#x3�%˥FY#rh��"O�!S`��T¦��deb1�C"Oz�[��0)\Ds	Et|q5"O������s����V$�@"O8�
#ۨl��֗3���:e"O�ay�c�3FJ��0�a��ZĈ��@"O�9���2�=	�/����d;f"Ojm�C+���(Y ӭ�5�:�#�"O��z��бT��	W�V�L�l�b"O��ҷ���'���6n��"O���f�\��A�DF5A��s"O*���AQ�?'nԓG�J?8���S"O&EAv�͡MbQZ��`���"O6����:
�a`@�	U�u"Ǒ��M�+�~�S#���:� �X�"O&QK�Ȇ�&߼�Y�fI�%o�!� "O>��c�R���t��*0b�Pb"Ot�鷏��M����BH���@�"O(��V鈧	p���21A�4� "O��{��#W"�<����^̤R "O8͛�*dj���c�÷�t��"O��c�,��$�.�I�Q"O�H!�.�� 7�b�y$g�<�!��;wP��I�o���³C��N�!���<�R��&�np5�6HJ�0!��4j}੘g隹^]�A�;8!�Au!6�"Fm�ظ�ɇ!�� ]9�ܺ�É�Up=���r!�<D�Ga^�1�P��Q�U�!�d]	+�N�	`�\�����!,�-CS!�,(t�a���Fq�d,��:#!�è&\��' D(��MQ䍙�|�!�D<7����I)pfةDB	�!�Ğ��(}�t�5f�������R�!�D]%]��2�RoѲlp��W;$�!�d��l��È���r�@��/�!��o��IĨF-�R`r�A17�!��F&u��m�5�ͥY��{���$�!���s���͘)
�~I ČW�E~!��V9Vc`�;��G�Fj^�S$%L�u�!�d�	�D�8��Y^b2���F��b�!�dZ;&S|��1#�GC*M2�V!򄁎d#�٣��,7(\��V���<!�>=�jLX$���d�\7!��W�zQbx`�"�8xl1C�`[�:��'�ўb?���G�X����W'� �(�s�"2D�(�c��/*���!� � :8��O.D� �3�'Gw8M2��߆eJ���@*D����jϮD��=�f��BD��J5D����oH
��ab�	D�\��i?D����j����Ǆ�B��A��J<D�Xqr↕P(Tщ�{�āCQ�;D�� @�h�A̮��i�'��3�N��w"O�p� A�1�XB�'��:��0�"O�I�(, 2؟rd����"O�I9K\ g��1 MR�&v<���"O��q��K��I��F8i_�D��"O�h9���d��H�~�Z�b�"OdY�̢n���6d�`��p8r"O��Sg�ɨ�E�r���A�"O��c��߉^�D�f��e��}�B"O�� ��ЬeʺՁ�@��I `Q#"O�%XJ¿ ׼�� o�2n��p"O��儃�*�� ���Y���)�"O2�93�&W�����F����P"O�P�K��U@%�q�8�6��S"O�E���۲X�25z-L�/�.��"O�
S)�=8�lh� �ڜY��"OB"�cH�"h��e/�|IE"O\�PT�Fz��Ijɒ0�. �"OڠC&㊚BlFGF�5��8��"O��B`�Q�O$���c��|!�"O@P�4�F�D3"�D��;u"O��6JQ�C��!� �%U�HUѓ"O�M����7i�u��@3Fm��q"O<M*��Y=Tz��=�&��"O^��Ξ�rn(	���8G�d@sR"Ob�8�Ǉ't�*�j��9��4!�"O� /UL �"́�@Є���n���y�h��e��: 05��dh����y�+�HB��cU��1��D�f����yշ/�,�`F�uT��%� ,�y�RV�t܋B���h�t�Ц��)�yr I;:7ڤs`�oyp����K*�yB��x��g�0�AE� *�y�LF�A��X���^�N0��[��yR��v�I��CYB�xȇ���y�ޓ6��y�eϩG��)��_��y�ۡ�ƌ{�#�Oײ���D��yRm��HPq󢢀�OS����.Y?�y��-f�|�R
�W�!zB�� �ybhK!C�� ��_c���H"ˍ��yr��%w����-C�D��a��+�y2'ҭ
:����7�x�*����y�Ȼ6B���J�5,�p��-�y�o=l�@����
fo!q`F;�y��"dM�p#R Ѷd;�=p�)J�y"ib��X!���E�DM�tcҢ�y҇�"un�+fV,��I�(M�yB�R*I|r�X��B#\`����*��y"�^�s(�1���P�bxY�%X�y��ͳb�ItBاK�����ED��yg�X�P�Z�A3@��y��;�y�D�*AS~�����5�آ6�y�k��$�"q!��ؼ{j�s3�_��yR��2�#q� � e���kU��y�"��M���V��5.�,�`"��-�yRaR
[��M0��#���Q��y2��*s����P'4
��ae��yb��$|�P`)��:AYx���ا�yr��H�4X�C�M2��bgCS��y�ҟ'�j��R"(�`J��ҋ�y�͂������m�Jy�7̝7�y�� 8(e���(h�z'��yB�X�S�6`�`"X�Y����6�E��yR���|�p7(����p�n�
�y
� +p���_}�	ku&]��s�"Ox�XD�7-(����N!C���"O��㥥�
>�r���ƫ6v��aV"O�y��A/�`��&#�ĉ�"O d)�J@�g�X�R��Y>���"Ol)��	څ�,�� �Nn ڰ"O�����ƕf��:L՞(�����"O���԰i�
�\�������#�y�jIg���h���$�x3�'/�y��r�hQv�N�q�
P&�V��yB/W+S�vئ\�}F�4*��T�y§��z�q�o�:F�~�{�\�yBl�3 ��ˆ&�@��������y��O��I�5m1,:ԁ��y��1l7����)��e}�	��(��yrj��QV�%a	7]�"�h�J���ybĐT*���ڈW�[��3�yBC�cFr��RdWWe�ESa���yRC�.U
�"���le3��H"�y�6��,���#	>XT���y��J>�cգE�,��i�<�y�<3ш���ٍw�j�A0	�	�y2���[��y`IB�m��X��`Ҷ�y"+�*Y�9��Ll�ZU��L�"�y�� j��4�pb3`�.�"�� ��yf��^6��:�"��I(p,j�P�yRm �5��U1U�]�H�P��`&_��y�m�i�Z��̇�u
��@ރ�y��ق%5�����دmT4�#�LC�ybm��ܐ��*U�f�.<��)�yrI� Eo]�7a)X���Է�yr��~Y��p�DQ(�P�B��y�/V �P�G�	VH����$�yb�z��xsC�¡0������y�	ň9��Ҧa8R��u��)���y��P"��X��J\(-ymƪ�yr�B(qLJ8�4ŕG� �+E,��y2ڵ��Y�
��<���W
�y"�O9J � ��X-��A�.�yB���v� �!��y�P�����y"WB
����7t,,dPFJH��yB��8f�)���݀f������yb�H�8^@ D�̖ear�ti�,�y�'D� �bt�r��k�(�@�g�%�yB��'7bIp�vp�p2-ϓ�y��S�<�JA�t�T���\��y2�P 37� �s0d̓Rʈ��yb�W,3d��Ӂ�$A�4q&@��y�"�^f��y��K��������:�y���34"Jѐ�dV��v�#Uj���y*��GR�����A
{l��4#�3�yY<w  %�ǧj�1��!=�y"�_�T�v���mT2�zi�fh���y!��Ms���/N^lX���yb-�)Fr���ӊ?Z)kt́�y�M�?D�ui���2�H�S���y��%F8�P��
 .�Ik���(�yR��L��ѹw�ѧxÆ�]����^A���JK�wo41C��Ѱs�ʌ��1�j��tĆ�@��ԫ�ZZvp��4j��toR�^m}���\#�t�ȓiyp��$L��[�"- CԔW�\M�ȓ@�����<��������D��A�Zt�2O�0z�N��?TT��S�? �Y�G�P=�(i舁&բ��"O���b���S�~x��'�%s��Mҗ"OJ�`���1��`)�Z�:�|̹6"O8Y`/^"=�`���ƈ#�v��T"O��Jr`�87���d�H^ꝳ�"On��v���G����b�̐LLd�"O����U���KX�l3\A�"OhH��V/���kJ�Ɩ99�"O����J^®� �ME�g�Ʉ�K���ҁ���:����l�v�f%�ȓG��i4K�tQW�Q��ȓX<<���_�|�Z�`@*���p��~d��iF�m�`�M�$`.� ��9n�5!FFB�i�ݡ�+�u䴄ȓ X�h[eO;zx���[�Y�.��xF��sAD�(�2L�TeZ1���ȓb����-��jaP�IW� �O�U��.��X6M�'YK�\��+��eI�<��J�ұ�EfS�Y�a�yjx؇ȓn����� \�A��aDP�|@\��ȓE�h`eF�% �\�qq�U�b�����o��I5呶ox�T�2�o-�T��$ �AP�E����^Y�@��ȓDzZ����fK&�G��A���ȓ@����q/�{e~��T+ކO�J���yU��i��(����B���'ў"|�0N��v�By&a��c:���z�<ag�}P.�D�W���=C�H�Q�<�0D�?-�ChD�!%\p��
M�<鶇ԋ%h)��B�R��:�Dp�<	1�X<����bN�7zQ(�I�h�<a)�.0H4�r
�(�#���d�<)wL%&���+����W�t��!B�a�<�u�^��]їI�do�47��r�<a0fp���7���W��d�KSy�<�W!ݞX�H8a�,1"}$��r�<�@OJ�	����nV���]��/�o�<����R�ȓ���s��x4�Jh�<���O"p!��ɖt�qA�b�J�<�2�� A�$�"5�	}��X��C�<Y���%@bM�WN�+H"b�ׂ�u�<��Bӟe�����"��8CΝn�<��%Q=ӆ��teT%Z��&ea�<"��+?k���t�ˈ)5��C�*c�L���,�3�t�j���{&�B�	�6��`e)��?�<|{��\*|��C�I]J*d��(Y8"���x��C�	K�t�Ӌ�b_�	('��I/tC��:Y�&�J�섋�c_ge�C�I�vU2փ
�L��[?x��C�5&�L	�w݊gh��@���6-C�"%Z
ųB�V!`K� c̃�h�B�6���pq�X$R..ؐ��݈H?�B�I�.��p8��	:Rde�gg�fҔB�	��Du���+[ U�X9weC�	�uP�m	��f�T���B�I��z���f��&c:��b��B�	�)�L���̰.�bh�� ^��NC�	�m\�X���*�( :�`�6�.C�I;��x��L"���%kf�C�	-�L��wK�4.|��Ia#E�b��C�	�^��<���^ c��
Ī)ĨC�	<-�d(��ǌ�b��,0Ʈ�#�C�	�T	:l��kץtx�uɒ��@f�C�)� (�[�O�5/�`3�ÉG�J���"O6�*@��Nu�1	������T"O�cU��u\Њ���+�XX�1"O�4�7'��9haW�+�A�p"O��9v%�5𤰱#�,	�6Uæ"O�,�u+��xX�ա(��h"O�)A��Ԭ!`��\[b��P"O|�jVl[�qF��jPe�?2?�)�"O�]d��%H��1�$Wk(�I�4"O �ѕ��'0���bз:�r�"O9A��� N&�	w!�C����"O.1��"Nt�z�� F�)���:�"O�	1e�ݤ���s�%���0[�"OZ�+��������ӛ<�Yi�"O^��m^�A9F����G�:_@��d"OPI)�,ˇh�
�K¤ʵ_N�PP"O��b�/Q %\m��F9-4��QD"O8,�BdB>��i .���5"O�J��O?��cf�8{����D"Oޕ é�<9�Š7"([���"OT�ҁ��K�쀺c��Y�y15"O D���UA%&�1��"܊DK�"O:8`Q�W8�v,��kɀ+�q��"O`�'��Ld�,��I;
�(�"O��0�R�8��%I£ٚ`G6A�"O�ͰG�[ ���GB 0K<2��G"O��e6����1V�dJ�"O��E	N�\p%GC�+<|\Kt"O�H�Piʩi�<)@�ʨ�ۢ"OZM��lB�7Z
�{pH�-p����"O�%�`nޱ*���3��4g�����"OP�&�)fsD� '�L�@h�%"O ���2�j(����M�����"O��[��
.M���k����ԛ�"O*u�Wh��pM��GU*G��}`�"O�Hu���OG���gg��ZT����"O�Q�e��C�0XI'&�.T~9"O���BLN6+
Q��=|��5�a"O�u�Dς��4�rE)�b���"O�0�P/P�u��Ě�c	�h)�!"OPE�%j(�Q3"i�=Q$�s0"O��1Iܰ,�6Zf�y�� �U"O��;! P�ِm�C��.�D 03"OdAŗH6۴�խR� �"O��iRΓN����� �kmNh�t"O:-⅍L������.��"O���'�(�+��ީg�b%;P"O�Li0"_�r�%5�)C�`�"O,Eh�O�X>驰*M�+��)�"O���Ǫ��Cv��r>�izs"OrQ��Eɒ�*�ѠKU�@َ��&"O���;=��E��F���G"O�x�%&%Z�̑�I�����~�<	��W(Z3�h6��Rx���Æ}�<���>�$\�����F�n��+�|�<�eBĪ,>�����vlf�#H`�<���F�{G��H9��Ń�S_�<���Ғ� ��A�O�0������d�<ٰ���PH�H�+2l���ڧ`�H�<��N�E���*��ҵ[�BM��<QW-؂;���0s�-t��+7a�S�<y�E���m^,c-�嫳	�D�<�鞥'sVp{Vf��I�n��6�X�<�gkK� ~�|0.�:��}�"b�_�<� �1C�h���$�*�M 1W�p���"OV�S�Cz�D�w�g�N}J�"O��&�޷��{�fώ4t�2"O�ݳs���8�T���!*8ɺ0"O���ъƠV��[1k�9L�8�v"O8`yB���6-�`��<-�q"O��%� =n��ț4)�B_@�t"O����í���Jq��?@�I!d"Ov͹�K�7x��y�®�&W!�Y�"O$�!�ճyVX)�-٣rzb�3"O�H�h�(7=�x�dAN.�s��O��k�ʇ��M��O?�	(}��4���O�R��ږ���~����G?I�&�P��8_S�u`���I�b�>����M�N������*&��AK�i!)���T_���Cb�(h���Ѡ�o\F����՟4?���c���?M�TѴ(-΀8p�M��ꧩ�O��d9?�{��M��6i��y駈K%5��h%�]|?���°>��"ϟ�>�"Pl���b�+�B8?���y"�v�6�$;����m�2+H�eh�g�Dp�l#1b�&����mZIX����(QɆDv�_E�! �Ö�\�BYSV�ɜXR�a�6B��rU�����Q�D"<a�,�)$&F%��a�:"u`�'C�0<�2��䓁.ޭ*��,u6�a�O��tIcHي	d��hu���5⟜6�Z�ȇh�2-��pN��?)��?��]���gy��'��	�w``c��Bli�@iу=0���D,ғA�#gI����Ҥ�ɓdv9TN~����5�d�.�D�<�F�ϫǂ%��ė�O8�Y��?_wh�B��V���<Q��_5�c�V:l+<!��%�ĮQ�"B)<��D��{4�xb�ʖ�1C�"?�
ܼ`��@���	���@B�(��Q����:�� #1�i,J���cCRh�VW�O��P�'����Q�U�_��y"��v�*�����J7��O4��?��*�>�P��^�q �52��M\�$��S�LH<���=<z��eэ;n�(�d�Y?��jf	zܴ��ě�5fډ���?����X-a��D/O ���7��So�5��Q��Iԟ�� ��/����[2zU`��$FX2d�)��K�za�c���]�Fl�2պ00����⯂�~�ny0�`�iW6ܐ�M�/�.�b�IG7Q�1���Us��#G�	퐸��П�ē������۴�?a��*�1A%P��#�*1�p�Ag�ߟ�?E���H���̹}u�	be��&)n�0��)�S��M;Vӟ�-x�
��S����d�4B��O<��S���m�	yʟ�Ox�e��(�*eiխ��q5���y��DS����e��\HD�!;�-x��I��G._�@�X�2g&4͚IXQK��M[�߷6*ۧ��*3X���s���uL�����*V�\c{@yE,�1e|le���<��Pڴn��%����Z��i�(�
��ļ_F���ubN-M� l:�'-�'�d��a'x�9�M�EDM���d즁�IB���Mũڮ��5��+T������텍Q���'s4t��	� =���'�2�'����M��y�-R�H_�p��b�GѼ��=0k��q�&5��
 _����Oٸ�Gx�@N2����`� An�H3D�e*��R��4AchG�I w |�	��x�在 <�-����<��bR�TI� i�&yJ�9�))��O�&�b�'�6����D�O��n�%�(P�9������{��І�`�'�@HEM^9���Ң�pCLQ�_˦��4��|Q����䓙5�FL<# |  �   -   Ĵ���	��Z�Zv��9/���3��H�ݴ���qe"�$�6@; <r�il��aDx!Ei��K��+uň);��6��ΦA��4H�{�*S�.��LZA���A��5�̴��D��O(I��48���Uɂ�;��`�F,^e�R͕'�ڥ�۱:-��
,O�pI�o�s�꘠[������"�v<�F��"�@�	�K:�h)Sl�C?��'}8ّA��W��'Xj�@!�� ���EϝK^�Ը���hdpDx��}�'\lΓf=\D�E��.���q�I��p}��%�0r�+F��'�&]��@�N��h�fQ�-6�5h�' �Dx�j��'�Z�+QeI�|���f"��.�n���,�&"<Aڪ>�7� 9����c*�gx~L��M�O�$K�Oeq�{2�`�����]
�>�(W� �M�,/O|"<a���2/(iӠBA�4r ��#L��>A�c?"H��o�j�H�GN�P��m���X.R��͖'�BAEx�ȘW�k6+ӡ�]������	��ʶ�,�)�(#<�!��O���Ԡ^�.F����M�M��4���dR�O,L�L<A�TU�8s��6DV�r���G?q�%&*�LO��98[$"�8�f�c�C�9ϼ��q�_�$�"a��i��?-��I�E㟎�R��8�N� �@�]��}ʖſ<�G���;�D�'�,H��K�8�tO����L1;轰��K	��� ^�tڱ�ɾN���R�+�x��h�oǇbhje#�B<D�����   ��ƊI�X�8��%�<��i4���R�'��'y�O�A�1�`����d�#F�����?�����Şa$���C֨X�K��,�ه�>�ȁ�\~y�g�$|o|��,r��'n��A��|3v�
����r�\&B����럔�IߟP�i>��'L�6���ys"�dҏF=��ᶁ¸;P����f,Y$��Xަu�?�2W�����X��\�^��3��AF�� ��P��u��ȦI�'�B��6!��?��}��ּ�Z���1��3kZ�����?��?���?Y����O��3���
mq� Y������W���I9�M3�jE�|��sA��|b'[Q�!l�*= 9��.k~�'�������ݹt��֓���6ÜRX��ϖ�M���'��!��O��O���|"��?Y��N��u��j�u�jY~Ah����?9*O��m-b���џ    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  ��   �  ]  �  �  *  z5  �@  L  �W  gb  �j  �q  9|  ΄  �  ^�  ��  ��  >�  ��  �  R�  ��  ��  M�  ��  	�  K�  ��  ��  ��  Q�  ��  �  K Y �% �- �3 : �?  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e�'_|#=�̋�/hNȉV!Õ0u�(�kRD�<Y/ۥG��P��7��`yW�C�<Y����:�kBJ��e��`�F�<�#�;  A�ц0��J�ܦцz���MK����gTl�xe��bx�ad�$@�ih`$W*Т�� ����A��H@H�a�1E|"F���'9�'k6&I�%ۙb��4����+e"���ȓ'�t�I�!�%jJ)�mW!v�H��	��HO?�)��A�bX(�h&H�\A2��O�<A��Ũ��a`�G(k��Rw RVy��5�O�TS`��C�����ȅ���<"F"O xS0/����x��F+k�H���"O�i�&m\*nچi��� k�P���"Ot�*BS�smK��8�!H�ż�y2�3^'L��1�A*q��'T�y"�u��ԉB��J������-L��ȓ:0p���U-
�ބ��DDOlZ	��#w~�HD��~�aUi<cl���Q��`
&+M�5i H�w��u�ȓMq�p�)�.� y4�P��ȓi�,�QDT�_1��㱬��n��م�F���@�l���ǃ�5
�rL�ȓ�R`!�,�f�"������5��}�ȓQS�}��j.n�j�@�n�
5 �Y�']�������J)�#��x�N�(A��x/���d]}���?� � �ۀT1.�HD^��y£�^�����ѽ=T�⃢Q%�(O�܈ç6��Y4J��n����ÚL�e��Ah����;����fA, 8х�v�������p=VD�!�
�&�j��ȓ&��ܣ��F�P\x���ɰW~���O�-�f� t��b�'N+ ������C~"@�Zt*q�S-�2KPXI��i���y
� ������D�aƈз#Df���"O���U���~�%��H��%��]�"O�]���/h���ƪ+���i�i�ў"~n��"ݲ<q�a«r�<aq��F��C䉹g|ށۗ)<U&伃��W	M.�Ɂ}��~bD�������ۗ>n-B�@�˰>aش���B���$�s$�l%���}k!�$ޟz�Y У�D�rE��F�-�џ�D��`�#��a��W�c�0m���>�y2LBmW�{4"ңUX���B�3��D=�S�O2��CX�{AS$,�<���y�/�6�+�W�����tdQ�Ƙ')�{���GOd���`�t!�p��J�y��	�<
 ��sz$E&�H��y�9Hƥ�ĩ spP%�E��+�yBcF�;C�}c�?��ɵ*���yr	�0_zA��	Փz�T�U�ĭ�y��çe0
��W�Ǩa��K �7�y��֫wnX��GQf��B���'xazek����F�� �b 0���yb��)($X�ʡE,f��Cg���y2��$�@�S��䁣	����j����>Ec�G�")R	tds��%a�K9D�x���ʞm��*� aX6���,�i���O Xa�w	��k���gj��?Z���
�'�
 0�Ne�!8�G75�8x��O����	�k�`)�b��<	\4��"OЃ�i�&	�Z( #��(8N QQ�"On��/;P2��#�W����Y%"O�h�O'N��<`�S@��c"OUA挼{4J�Ks�R�8P��"OL� 7i�ǜ���Ǌ<�d:C"O��2��թ[��lh�	Y,-``p�"O�Ube��u��٘V�I�����'31O�}�P�S�A5z��!�ofx��"Or���ptH���e��B��b"O����٣MA���1e�E��<)�"O��P ��b��7�F�MdLb�"O4	C�ӼRq��Zd+ ��s�"O�ǼL|�Qc�b̂��e"O��X� Ֆ�!J���9��a;�"OX�S`�D5b��q��w|�
w"O
IX���C�AqE��(�b�"O
��O�#%��0��?�<4xd"O\*G��|��	B�C@�:�J(�&"O�x�!��!�v��$�Q�$% g"O��J�,�t:₃���nȪ�"O�h�U#
�TS򇁸D}x��"OB���;@�J� 5&�Np
�ap"OD%��&Ӛ>E��UE
�\ff�)W"OZ����>���wҖH�
�b"O,�Y�C��C�"��딐[��=�#"O��)l�U�=#(��Z���"OF�ڔ���D��MJ�f�l��(�T"OJE�"A�[��a�C�W�q�$#"OxŁ �߭=TF$p�cI��F]"e"O�c���)CUv��6��q�"O�M���ıUm���/ rep���"O$��G"�W������2rH� "O��֎�?Y*�;��R7f�yW"O���W�\1k�E�`+�%Pb�2�"O���po�g�:t��,;��c�"O��� E�H��W�Y��R� "O�q� ���7'.Ց��F�����"O� Ќ(7�p��q���8�dj5"O�	����DM3���,L�'=��+�hѷ�f��55��1�'��؂�,A�_ej�c�W�9�(�`�'vd+�s���� µ3E�ܸ���?��?��?���?����?��2H������؋�jJ/UL@���?���?����?����?���?��+��b	-}d��r�g��C7b����?9���?)���?	���?	���?)�-��,sp�Ĩ���3
Ѭ(2�T���?���?y��?����?9��?��&�Dux4Gĳ}>�$(�*��4��H���?���?a��?����?!���?I��$��!'a�ÕhY�P��$��^ҟ���ߟ���֟\��˟��	��8��������:y][�'ˤ<�5h�/J��I�T��џ���矔�	����͟D[p���3X4�*֪s�ڱ8ӊ�˟\����(�	ܟ��	͟������	ߟ��r��?o~Q�E �-^`L��ޟ�I�������	������d�	ܟ<@JR���YAD�.Z�2%��ş,��ǟ���ӟL�	ПH�	ޟ�	�CP���@\~X  ���h�Н�	ޟ���쟜�	؟���ɟ��	ڟ���u�F$��ߺ8��$���������D�IٟL�I�����ǟ��	&.�~��d��ecv�<Y�@��IƟD�����I�p�����i�4�?���m�6�Іʿr�-�'㞁9�B�h�]�0��Ly���O��l�u.�yS�����#U� m(Q�Gg9?Y��i��O�9O��Zu��p`� �>� gT�
}���O�(�b{�D���(��OzR������|OЊ�`
+�%R�y��'�	^�OR���5Ƙ:{MAX�"13j�`�!�yӦP�u�d*���MϻeX�2�a1oY���hL�m�<Y��?Y�'��)�Ӥ'ټLn��<��m�)|��+Wo%�x)��<�'�p���hO�i�Ox`��\a޼�� F�L�m�0O����vL���ߢ��'��X2�	!�� �&g#� Ѵ�dT}�'�R1O��t�t�`G3Ğ��!��0a~�d�'j�KٓZ��tI���k�ӟpI��'�>a���@B��o�P�G]f��IIy������!9L�YziP�gʔة7I�;�����Ui9?9��i��O�G�-���K���>�jE�c膎:��D�O���O6l���n��������ZD!܃?0<$��$��{����O2�䓄�4�����O>�D�O:���h@�`R��M������Ւ(O�l�#����	ş��L�Sş@[�?$�l@�	)}L�lإ� ����<7��O2�O1�Z)��m�="�(�#JU'@+ܰ��%s�̞z��	�
�z����'D�U&�ؖ'�XH�2S�x���▪i}"H�B�'��'����4]��������J韨��Iդx3X�"��@��$�b�}�Z�x��O����O�Nܷ\�
��ʉ2j[��[W�bC(�x,y���^@<�����(�2H~"�;c��\;�MV�8�᠍8
j����?Q��?���?	����O�L��W�F�ֽ`R�¬d��ta�'b��'Ir6$Q"�i�Op�oZQ�	 Fv�d��ٶk�~�rT��M�N$����Ɵ擟,���m�[~���2V\E�g�ޣLdv��L�&Q6��u�UU?iI>*OX��O��d�O����0O�	K��hA8�@�	�O��d�<a��iT�TY$�'���'��_* k��X��ě2�/�������?�O��M��I�X]�Qa�A~�;�Y)q@Z�A$ˑ$2]�i>9ye�'��P$��Ѣ�H<q�䚔(J:X��d�Ac�ПL��矰��ޟb>9�'U�6�)���!Jȣa8�m���O�q�|�p��O���X��%��I�����OҩiB�S ���à�.|cdTS�,�O<��MZ��6m&?�;8�����'yc�ʓC�b�2퉹'3��2(^(HTI����O����O����O��$�|�$%��!P�t �9<����"�W~��N�D��'U����'~6=）�����A�'��'T`20��O,�b>��FC����q
�LW1�J�ue]/���P�EQ��O�չH>A+O,���OP��!j�!z��hDǛHj l
�L�O����O��d�<q��i��|y��'�DE7S�1!t��+�;)x���ĉH}2�'A�|� �!F��TB��0֪Y��$=���� oa�}�e�C4,1��y��z, ��֓N	��k��_[�� �a��-m$���O���Oz��>�缋�AS$5�1�%��1�B�@�I��?钸i��1V��*�4���y�F�r
\a�M!i�}a� �3�y��'��'|�(1�i��ɛd�h@��O��}	��@�2��)l��Dy�`�W�iy�O]��'��'|BfWq�V�w�{t���q�^�z4��=�M����?����?yN~Γs��}�qL��>��C�ΌLO�y{�Y������t&�b>uYAo��1^�i�v�K�=u�@�.�'�C�0?�"�W"3D��������#I�ډ�Nǥ:"�l��� �x���$�O\�$�O&�4��˓4w�6g��_�b�.
0�|xb"<|j���_BB'kӎ��8�O8�D�O���B��,��ˌ�/���E��B
֙��gb���b�) b�?�$?Y�=� r�� ������c�� �yr�?O���O��$�O����O��?I�ߧfV�-�3���DʽB�� ��l�����*ݴ[��.O��m�i�&h<n����%a�>D�ֈ�Q�y&����ԟ�S�.$�l�S~�	���%��D.�̌ ǌC-c���Q
ӟ�Bq�|RZ����� ���<�R7nP#���Y$m��*���	}y�Ff��#I�O��d�O��')!�p��BἉ؆E�
���'����?����S��l�s/�;a���v�	�]輨C�O.�~��`�/��4�N����,���Of�Y�n �F�n�F���xf����O��D�O���O1��˓AZ�v��2\��n�T9az3�
R45"sQ���4��'2듩?ɡ�ʾ	��ݨ���$��P� CQ��?��[ł���4��DC-s7�9����M�5��2$�!`��3E�0�y�Q�X�	ܟ(�IϟX�I͟�O��SpV+�`a�oN5����kt�~�A�*�O����O���Ҧ�ݦ>�ʉ���T�.�
��ME�v�Hl���%�b>q6�@Ѧ��I�Nipѣ�'t7��)�^<H�=�}�g��O��H>�/O�)�O��(�Ө[ڵ[��
�$��G��Ov���O����<Y��i��җ�'��'l�9�oПf�� T������u�O���'�R�'�'|��tj�B�<� P�(��C�O�y蒡J�B]��+��&���&�?y���O���U��E���:O�X�L�O���r��',b�ԟ�_�x���H�^�P�9�D[:!�n�dQӦ��e�˟`�	��Mc��w��z��WS�pq�	���IÝ'�V��Xwc�}�'�0�	*��?�z���\S΄��,b�����GZ>W�'��Iğ0��ٟ��IΟ8�I<D��6C�&"MH� �?m�ԕ'��6MM�7\����Oh�2�i�O ����oȥ9�jȤu<�@b �n}B�'#Ҟ|�����
��ۃa�Z�Nh�Ԥ2���{�i+��&��84$��d$��'`P�ۀ�^�j���vH�#�N��W�'���'�B����Z�Hr�4@��#�<���k�[�;�聻F�ލ}�Z���gt�6�ĐZ}r�'�	�[��� [�8�iw
��$A����M��O<"MO-�Bg�?�)��>�kf�&��]� D׎����<O����O����O���Ol�?�r�g �3U�`���[�v;:�u�W�P�	՟@
޴d����-O lZf�ɧ'��+� Lo�L� 
�`�xm&�(����ӷ!��po�]~��ɕ/�t��F��	LN�A`���?@HU��kG����Д|�[��Sҟ��I�H���Ҳu�$p�+��U��"�.��P�	Hy�	qӘ-�P��ON���O@˧i�� �-W��fū�C�5p��0�'C4��?����S�䉏�G�~Ҡ� O&��f_���{N��xi��O�	ސ�?� �)�D�W�h�V V�fmа�cmӝ���d�O��d�OD�4���D�OJ�F�➨yK ���/Ϝ=\�@��4a4�%���'�"�g��O��$�K}B�'��0ʤ�J<:����O�]|
 '�'Q�H����>OX�d͕ct~����x�h�v�"�
�d��I��@�1i�=7�d�����O����O��d�O>�D�|j"C�����$I8|��l1 DȊ>��o����'
����'N�6=�-�bM�T�
0���=F/����O��$ ��DG%z7��|	�兏�(�b�)6��4'��`?O�x
`j��?s<���<�'�?IaDF"p�t`C��1�r�+� 1�?����?�����צm��g�ޟ���؟�B"��V����RH#z���Un��Ul�	埬��K�ɧ^N29�p#Y�^��s�H�)e��x�RY�$T4�Mp��d�Ii?��l�>U���s�B#Tɓ�h��!;���?����?q���h����<b��|�tG��F��L����(����̦鉃,_y�}Ӱ���4q�f�K�kS<7mb�F�Zd������I���{��A즍�'�i����Yr�e�3;Q�H��-���sr���䓒�����E"�@�ĭ<����6��eo�I%�Ms"G�,��D�ON�?���$�lb�Y6˔�{�N�0��M����Od�d&�󉃮+�aJ�! �N��[�&#�����l�M�ʓ}��Xj���O4H>I/Oh4XGo�w�ʕh%ȟ)�ı���'q�6M
O�`��$���%�3JG�Â��x���̦1�?��R����ϟ��	<�f]�fnGJ��r3a͖Wr4ѣQ��m�'Y^��D��?�[��$�w&,s���t�y��$ 
7�\��'�r�'ar�'	��')���B�`���>��N�U�F�?����?y5�i>�Ma�Or�m�X�O\1�FD�Z���ک
+����4���O��4��a
y���W����@�ڨ*)��*���2o
���d���䓋�4�v�d�O��4A��ّ�I�V��$b���qT���Oʓ+�&��1z���'V�R>e���O�| �i�r��H���'?�6T�H�I֟�&��'�hF��*�l@�$"_צ�(���?Q�4��4��@Q�'��'p�#§U�U��#� +5]��:@�'/B�'����J����T� )۴3����
@�h�@�r�g�I��XA�/�?���Px�f�|�O����?�6��=8Y��[�qo���OM �?y��N1�<#ܴ�y"�'{>������?)+@U�� de�V`��J-�����M&'���Q�5O�˓�?���?9��?A���򉌬}(
ӊ"�=�׏��xn$X]�I��|�I[���p������hӄ^�\q� �0�/L��?�����S�'$�.��ش�yB�Q).������Ӏ5��{E��*�y�*I q<������4�*�$ض<"����J�Z�8� 橉�"���$�O����O�ʓ8ۛ#�E?r�'�"�J�QpN���i�f������RE�O ��'���'��'��l����Cj��y拀�\h���OРI���2s��)ҘO�Bx�	+R�r(F8R��`C�[Z$y���L���'�b�'�2��� �a-X%i��!�3Ql�4��K�⟘ٴ&A`�R���?A6�i��O��9g��A��$�ix�c�2|���O~ʓ�d��ݴ��D��L9�!���
g���j��
4�0�@��)[��A�d2�D�<���?���?���?���'�����	(d°Q���$��i���۟L��П��� ��h��2�$P�3���V(�+�����Iu�)�S8(��` �i�8
���!�c�:��As�� ����'����G�`�"�|�W��H�·��օ �I�e��y@��	��4��ϟ�xy��|�.����Ox��DL�0�C�-�d�(���On	le�ϟ8�O��D�O�N	�sl0(�(`����S<)4�"vӢ�O�Ȥ�e�?�'?1�ݜ~�"�˳AQ� �����A6�H�I��P�	֟0�Iҟ���^�'�(���� �̡&��� �J�Ο�Iȟ�
�4x�*��'�?)��i��'��I��(�2����қJ�J��|��'
�Oٶ���ie�ɫk����{�YR#CO6tB�O.1=��3���<��,�-{���֮��[��Ǣ�ODlښz��ݗ'��S>���Ꮨ+pP`��X'���É4?�"_�8��ӟ�%��'6�` IFABr4<�&�V�MS.�q�L��V�� §��4�P�b����O.�x���,SB�����0�F�"FM�O�d�O��D�O1�XʓS ��(�?���6MN�q�|�R�/\eW }��'�Rt���t�O����!Ee�L)�oP :�\�:A�K�^���po����4���Ȕy���'�.��bh8�L�*��ݫ"��(\*������O>�d�O
�D�O���|��I�N�`�y*D�@x�"�o��'b��g�&>�R�'/���t�'l�7=�|��f�E�U�`��&�(�F��O��b>��sM��Q�>�D�����e%F�����e�,�lA� v��O�iL>	.O���OTP��ԈAВ�	%�$V5��֌�O8���O̼��l�<a��i��(���O���'��	�gna��7d�
N��0�|"�'��I���'�`�ɭ[�iZe�s���'"�Dр���D1A�Qw8�HD�y�O'B��I4��#'b��!�ʛs����N;�y�J��fJ0��'생rgܡ�ŭ�.���v��l�Bn�<!ǲiz�O�NͷZ�F�H�Î��|ݢR��^��d�O,���O�r�+y�x�ӺsPY���Ů �,}����̝f����I̜yD��O˓�?���?1���?)�8��	� V��AA�Hh���H+O4o$dk�P�	۟(�IN�S۟D*UD��Zf$(#F	E��ҷBE���$�O��b>�P"i�;pF����	�:$X���� M�q7$my�j��gU ���@��'T�	3u�Z�9T��4-[\A���� h܁��ן,�	ϟl�i>�'>7m��d�1M�}��\��Z�Ӊď��dS����?��Q���	��I,;�Y��NX���8!kU��,��Ǖئ��'cx�S��?��}���u� \1a C�P�xH��#H~�̓�?����?q���?�����' +��*a�G�D���(��H�y2���kɀI��?)ֲi]ڌ�6�'�b�'��'������äK���c&劓<�x�ӈy"�'��'*�a��i��D�OLy��#�� ��DB�*��'�z|`��Jn�#��V��Of˓�?����?���	��h@�Ğ�v.^e�P�ւz�؋��?y.O��lZ$M6����|����b�h�aOA((95h[��y��'�ꓑ?i����S��Î�=O�ش,�,L���3N@?��C"�:ua2�B�_�操}�2�l�	+q ���rkƠEz6.U{��I����X�)�Sny��y�Z�PQ��$+�A�S%���h}�%��
d��$�O�!ln���Գ�O
��)���2D]�0��s�	=u0 ��O�M@��fӮ�Do$���ŷ?�'�0r ��,nV�A�Cؓ8����'5�	Ο�Iǟd�IߟP��n���S�����K	�T��-��66�Ӝ����O��D3�)�O$mz��x���*n����L�4�t���_���?�|zq ��M{�'�ą��\I����&C�&n�i*�'���p��ir�|2T���I�ث�N�u�j�e��c�pP)�)���P��ȟ��	]yB�x����O�O��d�O$Y���8�@ճ�^�"��ht(3�d�O���'�'��'8���P`W�0$(d���&�4Q��OLP��տ�h�.��W?�?��&�O�MQ��&\�t���N>��G,�O*�D�O@��<�OuR�'��
'G`�51�/C�g;�q�$�P���y���P���O���O��O��4����G�a w�218��¦��O����OZ�$�%2��7�e���I�eTp)�Ms�U�� �qz����V���3iA�w�B|��'0�D�<���?���?Y��?)bbM�Z,���m��-K��4� ��dM����p�����I�d%?�	��=��lS?��@!�?q$*a�Or��O�O1��䊄I#*C��+%��[�4h�e 6|1�2��`��ʘ@iBe{��Yy�ٻjZ��k
�(��1y��3�0>��i��;��'���w��R[^=���ĵJ��$��'�7-+������OT���OB	)&m�pQ6� �ٹ�<�cn��)�7- ?��o��Z@��I]���'ҿc�!I�.��x'��^3����(��<���?I��?����?�M~:Ζ((f�u�vF_s}�M	nK Q�N��*O���N���Ĉ�֟L��>�M�K>���ȑn2$ �@eL���\@��<Y��?��%��2۴�y2�'<�9��3f�0��X.�Da�+S/0�D(�	
CW�'��՟��	��	
<1k)�ȀO�>���I�� �'�.6��������Or�D�|R�4���3�o_
&$�;�b�Z~�F�>9�������8*�~4I�B) $&ybcn�7h���(XPd�*@g�<�'9j� ��(ڴ�4M[�>E`�� �ű9(�����?���?�S�'��ͦ�[�ō�+��=�P$5�̽ S�.� �'�6�%�	���O�xg��2y��š\�|���7e�O&���8*Ϣ6�2?��L��}p��i>�$c�z�>X���Q ��T
�y�X�@�	ퟜ�I���I؟@�O�nِ&��)�%��I��/+�=Scosӊ��%��O2��O����d���s��+âت���oȇQ�@�IQ�ŞX����4�yR �UP Q�(�%-�q�����yB�5��I�I6p�'��Iܟ<�	�����B�
��5s�X�a.�(�	�����'�^6�I�˓�?����H��!��L(�v��'����?ɉ�ϗQ���2�Z+t�Dh�g�ԛ��D�M蠴�v��)5�`�������7�����#@3|E�Ƀ�,�b�Ȧ�d�O���O��$:��SՀ�C��=�6V����P�5�?�ջirⰣ�Q���ش���ywN��:X�P+E�W��:�S��ӽ�y��'���'-�-jW�i%�ɢN��=�$�O��hr�V+=DX�^�pH@���V�	by�O�2�'�"�'r�%���i���s��,�� �
�I��M#��J��?a��?�K~�n��4
O�L����4�X*o��ѲW������h'�b>��M�F�Z��@W5<�vmc��ңA��iĬ/?���Q%L�n��X�����DЮG��U$�T�o��Lk牅a�,���O��$�O��4��˓,��� �!M�����L,2P-޸Dt�Dj*�2gӢ��2�O(���OD���9n��c.�\^@0����(�Q�{�l�6��PXf�;ʧ�q |�T�q�%u@L�� C�<���?����?���?y���lG� �,s��P N���؆E��T�2�'�-y�@��:�$�$�M'���J�	v4��.b3b @�4�֟��'2�1��i��ɽ>�t��N��	|��S� X*<�s���/��'�m��Hyb�')��'
R�5����`�.;�}�!�<��'�削�M�j��?I��?�(�<ũ�g
� �j���{vn�`����O����O��O���j7��G��K��� �˾D�(�vf3C:�D#?�'m��d����\�Z�Q�B�(1��Q���g���c��?���?a�Ş����mC�D�Mrĵ
��l��CgCݐ�H��'T�7m9�	��d�O�m3D��Zx́pf$�v�rᠠN�On�d�<p9l7�9?���t!���<�$��� ��@����$� ��yBQ�\��ҟ��Iϟ�������O�%���רdJ$���BH �2�#y�h����O���O�������V�������30r��n�=�����('�b>������]͓���:�Ӈ|�D�V��MuLuΓ"О}@�A�OY�L>i/O��O�t  (�ȡ ���=Q�!�j�O
���O��D�<��ib,��'&�'��:g��,	v��Ѹ#��	5��r}b�'��Oh,����aT8���c2sM0�PŜ�tbc���(DH�_�����S͟\��ݶ�1�w�SEڙ+PA1D�d�Ɓ �&�D�3�`�5k�l�A4�Rş�
�4o�n�����?�R�i��O�n˪6"-�i4?j�ij ꝼ0�$�Ov���O���g�x���b����7��?msV�\Cmڑh��s��k5E�d�Fy2��,D��yk�)MDx�H���
v��.�֩QB/����\��%�	#v����-Te���G������(��F�)�S�A��5
a%��b�T���� G�L�3�f[�\��'i2�@ڟXI�|_�X*6�
7��4F� ^��aE���t�Iԟ��Iܟ�S@y2	rӲ��`��O�d@$ G\DD0B�G�=R��Mh�2O�l�I����� �IП�a�M�!`J�Y e�1a_�u㵣�[�̑mZ}~�ךB`�t��Z�'�����{}sR�2r����B��<9��UM|t؂�'z�������Z�0E{-O��D��U�:��i �'����R�L0n��4�MŖ�u꒙|��'��OlT���i��i��
� ����ߔ�.���W��S�d;�?� �;��<���?����?����� ��V/o�$��1��?q�����禙�C�ʟ0������O�u!r�����5+ɵG��M��O�p�'B�'�ɧ��̽[��<E�~�t������=� ���ՠp��I�M�}y�O�����5u��'x(8��W<OL�h�C�Ћ-�,Yh��'L��'tB���O0�	��M��ĥ l�-(JĿ줱jP�R�X*O��o�C���I������0��S��BQI1������G��lZ|~��8�V��}�P+ٙT�@��F�.��B�.�<�)O��$�Oz�d�O���O�'j��)7�l���97�E#��
9�M��Mэ�?���?�N~���L���w�4,���V [�`i��T�aՖ)���'\��|����̑PE��8O���ǂ��`����00��}x�>O�ȁ����\��p�R}�@ z�E�.��=A!IF���q���Qp��T��1D�Ȋe�@�o'�XR��K�O�L�ņ�n���[5e�:�VT[׆ǯ9�gi�3Ik(pA�9m]d�!E�=�8�hGgA�YLP�8�Z���`��h	A��) �^-�� ��"���0
� �(b�kЏ^�B�pw��;� ��� GL�X��}S�B��N�)�@��iJ6��
����`ǘl̑ �(��rw� ���N�8�0=��&T
!nHܢ���B��TQ��^�_�m)�!J0Q8��w��
I����ñi1b�'�.��#�8�$a�蜒6��o}�t�1���Ov���	���s��}L̹�#Md�� �2��v���Oxʓ5�J�yg[?��	��ӉZPl�&�F�Wz��"J�4c0�O<)��?�'��'��i��g	���
M���dM^��\��r�J��M+��?���"�T�֘�\^��e��3�T����(l��7��O��$	7i��⟸�}��+�/"�\���OѪ!�p7��~mZ����I���ӝ��D�<��ᕪC�,	�HW�?�5�����7:���%���|B���O|�k�N_�Pd�PE�ɦa����զ���ݟ<��4-��@��O�ʓ�?��'�H��FV�& x	�	m���4��V��5����':��'u�=c��T 0�l	:�'�.��zӒ��V5R&���'��I͟l'���
,�p��Gb��a�D��.Hv�V��B����D�O:���O��A��ic���z���D
���*Ԙ"3�IVyR�'f�'�B9O�h�#/N#S�j<sJ�*\ �������'l��'��]�P��C���(�$"��A��hc����Kӻ�M�,O���)���O��$[�+���I�\d�٪�-�l"阔�ǒ���?����?�(O�B���d�4�'e�e�PM *���j4��
�tF�z6��O�Ol���O���J2�ɫ ����D�$a�"L��8[47M�O���<�/���ٟ���?��Gĉ$�H�����7���8"�@2�ē�?���G��Ex�ܟ�9�b�<C�;b&Ï^����i�ɿ?|qܴ�?��?��'G��i���1��v ��K�6 ��%�a�d���O�1���O�O:�>e�Հ��Ok����'cڐ�GMd��I�⩕�����T�	�?IN<�'4��ԯ�"uV q'Á)G6�}��i�b�'��|ʟ���Od�4���n��]ȼЖ�ő'B\l�����I�p
1`����|����~�.w���CsY��
}#0M �M����W��s���	����Iw�	���9\���XcN�G2Rly�4�?�⭚hh���t�'��'�$<����'�Ф#��0l5ak�g2��O0ʓ�?�.�2ʓ�qA�L�R����=Zj$	�7�P ��'�r�'�'��i�M�%�v���qǬ����*�na���D?��O�ʓ�?�a�����S�ZKm%�Ϭ-�t�Dk���M���?��b�'��	q��6�\�p#Ã� %S�u8��[�^5�'prQ���	?�,�O�k޳A����aتn�TQjce��D�d6M)����,�'-���L<�!�%5�j8:qFߦ{�!Y��[ަ��	ß�'/>P��2��O>��Ƽ�Ҥ��&s|�1��.D�rѵi���ٟD�	˟��IO�s���-��.f&L��b��q\��4�i�ɺ%�V��ڴRs��ҟl�S2���9O+��S��
�+�%ФʰY��Y�P��˟�J|�J~n�$ ��=�&W"��-���Ȍ1a�7� �a�^�n����؟��ӑ���|�獒�	d���bCF�h���FQ	�?���?�����S��OD�y�.K�>&����9��%���ݦ��Ih�I�]�4X���	,}�����@G)�,9xAP�
��\�"<�a���O��	k���X����j�Vq���j�P6��O��G�<i�R?Q�?�W�̄/���R�*	�Zp� �]�(�'�H�O��d�OH�Ģ<ym�l������.?�%��@w"�L�a�x2�'�2�|"W��C�d����'?�Q� �b�R6�O�˓�?q��?	.O�قF,��|z�ǖ�p�Y�j�=����j}��'�R�|�U��ȟH�«L7p0f��,8�� ����?y.O ��S��'�?���g���ơ�uVl�(R�`���$�O�ʓ
�� '���IA�e�$ب��F?}�amy�l��O���nؠ�����'��\c����r��4�z�Z�D��n:�,yH<�-O��$�O���$Pw���{����bO�L��a��i��I�'7��޴  ���T��6��� Z����'��)����Q�j@�!�i\��'z��'���d�|nZ�T��S�`�,l=Vz�	Ah6͊�G��an�ڟ���П�������|2EL�Wl0�á/�x���Vh@�'(���'��'�ɧ���pbSb�87CP�Jg�=5'�0Z����M����?��*�D5�(O�SE��UR�u��_�&] ѳ'�ětH�XFxb�6��O����OJ�sR�`�=���^�bdD�2(�����!>�v9P�O���?�(O���ƴD
���:h���.\6䃖�i�b�ʹ�y��'���' "�'/�I>5�d|�t��r\R�17���*���h�9��$�<����O��d�O������Rg�I�&"�\�P��M�����O`�d�O���O��!g�a��1���I�,�N2*0RVB�7�-�d�iA����'@��'��b��yB�٘XdY�p�I#>߈��b�Y+G'�7��O<�$�O��Ĥ<��cZ����˟0�Em��o�� ����_8؅y��S��M������O����O~�g1O��'x��J.8�0}iD*I����4�?���ݸ����OU�'���#ܤ7�t���ƛ|_ �����)(
2��?����?�(��<����$�?]�A튝V��:��Ny�
݂��rӪ˓n.��b�i���'�R�O�
�Ӻ��Ȉjc�`��,��Ip���L
ߦ��֟,�f�i�@%��}����^4\����^X��BɁҦU�1�K7�M���?y���*qY���'̄H�,ҿ2��]�bO�^\�h` z��a��4O��O��?��I�Hiqa�hے	��r�� ƴ�޴�?��?�ŋ�*���Ry�'F�d��C�$Y�p�H"k͐�H�<ěf�'剻w�,�)z���?�O���"�A�2D���2#�n=��4�?���T���qy��'����G�p  ��=�:i�$Q77-�O�|QW3O���O����O���<����\�*D������e�#'� �v�	�Z�Д'm"U����ߟ��	%b.��vj�h�
p��`��c�����)e�x��ǟ,��֟<��gy��V�~�8�G>��0ScT,r����U�rq6ͦ<������Oh�$�OFi��?Ok,�'�X�c���� $�����꟰���X�'�����n�~��' ��u�<~��س�f���R�i��^�0�	ןt��&����s���=^8"(�����H��S*Lߛv�'�bS��b������O�$��X�(t���/
�г�9a+f4��"�h}2�'�"�'��q��O�����Mn��Q�����mH\�i�
�5�M#+Op9��
�㦉��۟T�	�?!i�O뮇6,]��%AE!qHU(��N�i���'���y�!�~Γ��O^�;����:�8�D��|@��4b(t`�iy��'���O�j����oV���lĞT�0���B	��]lڴ0�IF�	q���?I7(Z�s��HP����-��� �'@����'���'�|�T̢>Q/O2�ĺ�����D
Bt���7~�*��#k�8�O���p0O����H��ɟl"�
UЀ@�MˊG� ���҅�M����m��X�p�'q\�t�i�]ڠǒ�?�����½9��k�>�n��<���?��?1����DL�V�PE�9�+A���-�b<�rA}�_�@��Ly��'��']L)�E+b��ę�"F���U�տ�y��'A2�'�b�'� �v�y�O��%3f�˳u۞,Z��%Z��ݴ��D�O��?q���?��(�<)fl�y@��%ؔY�ju!����Iǟ��Iߟd�'�f ���2�IE�b���f�\I�顆/G�i2(	mZڟ�'�T�	ڟ@ti�����Oflx#�=NHjP���'�8��P�i^��'�	�-24�K|r���#�J�!�z��Z��T	���'�'��e:�'j�'*��	�&����΂-+�j�%JґV��T���^W}B7mD�d�'3�TH4?�V��kj�Y������uB���O���O`��C�>�IS�'*WM�%�Ic����� <M	v!nZ��qr�4�?1���?I�'2m�'��h
�{Ė�ۃ��AMČs�	�,A?7Q�W`�)��8��Ο�[a�A�8H���0S��e{$�^��Ms���?9�� ���k��x"�'`��O*P��ݝy�
Dɓ�Y�-�d��i�'���Xr�1��O.�d�O2�;���v���+�������b��m�	 K��L<����?�O>��2�B����y��(���l?��'���8��'��	�<�	؟̗'!�����S�@2���
�-'�L��C�K�:O�$�O��O��Od����2m� �o�}�t��!.�s̎��<����?�����D ����'2��H�� If)����!����'"�'�'2�'��V�'y$��ѡ02TH�`f��Na>8)`+�>���?������$>q(Ө�y���S#��aS(��C��MK����?A��9*� ��� Z��C�o� :b=r���
@87��O��d�<u�Z-? �O-�O�8�t�G6G3���dM��29��q6���Op��e�*�D&�İ?QS�BQ �ݙb���*��d�n�T�p�Լ8c�i]�꧃?��O�ɗaԪ]a6i�$z�q�C\%/
6��O$��Y�\�t�$%�D8�S�/N���N�z�(��OZ6F7]��~�o�˟���͟���1��'I[�.H�G���@�eM�w�6�`Ft�\�(R�	{���?�D�
Ϟ�AQ5X�|�#Y�69���'?��'	�DbSI'�$�O������ ^�9�@�	-�R� $%˦px�XŲi�'�����%���O �d�O4��lW�����P	T�n����Á�����	�7B(a1�}��'Iɧ5��[�5�D��e�>w20- Â�9���E;L6�$�<q���?y���Z�s�eC�K�fJ���L�Isp|S� �v�	��d�I̟��'���'m��S���`^�@-D�0�\Ļ�����'���'x�i�oZ�ެ���5���� �QO���Ԏ��b�dlZ��t�	ş�'�p�IEy"���M�tl��\���G\5]R�z��Z}B�'���'���N��(�N|�`�̏45�A��DZ��l*ܶL����'%�'�����@�Ʃ!�i6pz�1�Ҡ�x7��Ot�$�<��� ��O"��O��9�����钁LBv�Qec4�$�ON���E�@=��^.B���
�%@Jj��X�Dk�C���M[�V?��I�?Y��O*8�SD�&;G��B��]�*O̝`��izr�'�����d5Ex(�/	&�.��5��j%�72�b�n�����Iȟ`�S����?�ÃԴ!*�qv�R3�� ����ۛ��X��O��?a��:���
�l�ʇ"V���i�4�?���?IԪ����|B���~�BF1%&���R�4H��݋D���%Ӛ#<�E����'��'Ĕ,�孑#�Ȁ�eP�TP4a�iӴ���:RP&��՟��IT���	v\sAd͑Ku$u���47���_`�b����ڟh�I����	w�����nL�rE���2��$*��Xy�'U��'p�'T��Ox!h�f7\�YC��cI�1�i&Q�O�$�O��$�<y%&܄k�޽p����ʋ�P�l����ԯ�Iן ��S�	ן��5-�b�C[H�sD��.��%�E;J͈e�'�R�'`R\�����@%�ħS��T�Fo����9*VMM5!�N��C�i�ґ|��'�����'Ɛ��"��[�d|2�Ƙ�Z���:޴�?�����/SI�Y%>m���?��raK��8�o+Xc$H
�':�ē�?���(��eFx�ޟT9�Q��a�D���I��/�)#��i>��s�6mcٴ*������ӈ���Nm'�\�Un�	�r�!O�u���ܦ��	�&#<ى��$J.9�����B�2Gn-H�	�M��'3q��v�'
2�'����3�$�O�	�����S��D�D&ro�M��_�	{T;�S�O��II�6fJImv�V\��	ƪL��7��O��$�O*!Y��Hv������	U?����Eڬ�⌆�1T``����q�5, ��<����?!��
���!��V��XD��GG�4	pV�i�r�(��O
���O��Ok�ƆH�D�KϽGo�����<���+�,c�D���p��wy���>oxj��m�Z���SE��@m��6���O��2���O����{���S�Bָn̝��� ##h�`����O,���Of�7XL��F2����qaK���h�&�,FL�ԟx��'K�'2��'�L��OfP5曠
2h�Y��ѳ4��0q@]�T��˟���Cy�G	56��F��wb�s�\�A�̖a|T�+�h��i��O�ޟl�ɯB-,c��قm��C���z����9����`�s�����O:�0h�����'��o
0��y�Pf� ;���u|�7Ͳ<�(O����?��|n��fy��EF��l�!�z�� 2�[;�~�\5�4"����{�D̤w�$� d�/A�� E S�y�T�G���ϝ�"�
$1�JB*%jRqt��(����,Cm�����V�@P+�M��6�Z�qgHE$9R"�ȥ ��A� ˕7@,m�WmA�=vj�*���gf��CE�s�>�{#&�4צ!�'%Ο#h|͑nF�"I � �1<{h�`ឲY�FHy�9G��@>6ʹat瘪'0b�'`��'�F�]ȟ��	�Jz�Ʈ#v"����:O�d��w !�"���,�j,�GK�?E��_%��EQ��߄	Ւ�FcZ!�ɣQ���UK.��S�T3pyd�xҟGy"��0�[$���zޔ��"�,�~�aݢ�?a��hO��{+b� �;h�`\c�M��8����/[���sU� O�|*���&gju	E�)�(O��#�����5JWA�����Qk���.L��J矘�������L͠0��͟�Χ:���7
��G5����AΙ�F����,��+@��ju6$@��Ǖ�X@#��~�}���: ^�U*��XO�~��o�=*��y��X�?Y��R�HeQ妍�6+�uґ)�X�v ����2�'VT��sE�Y:�P�1i^�[�ny�ȓ[��Q���K�M���Y��ϓ:���Ryb�ɭ3tD��?�+����@�d�2��aNJ�bnܬ�-	�p4r�$�Od��Ͼ.�@�zDኳt��T�O��I�0��]6	�
a�$L��Q��RʷHi�q1E�ѭ��O�۲��5�b�XÄ�4+�ȍ�	�\$��'�񟀬1��	}��[�%��w_ Qp2;O���
�nn�@�`K�6�����ىj�a|b"�C�X)�9�1�4t�x�cE��64��K�W�
Mm��$��U�T�7�?����?��*u���,�.=:�G'H����ܘ����*n?p�񶩕�o,�0@�-Bl����@����
� �� �[
<���W�DԢE�a�Q���d"�)��P���.��tO�3e��i(D��B�환tV���J��׈ը��1�e����'k�T�z`$�w�� 7$�,m���A���?a'�qE�����?y��y"���4�|��`��pGH)��DH-	"��OR8Z�'a�]
b��#mn|-����a��'���R�e�J��FH��S/$Mq��P>����A>̍��@���`���d�}��h	�n,���6"!D�ڔ�	-� ��,V��m�K��HO>qɄ(� �M˕�Q$ *(R�H`1�!�?����?A�'�b����?	�O'���?�Ȇ� �Y#�B� +0�rF�D8�0��¦<��G�X`�-�,�9r�԰ �}8��sÂ�O���_:	�,����̬$�Π6�Yl�!�$�v ��K��Y�\��	��`]�T�!�*�dM"s�*a�p�[�)Л'M�b��H�dޓ�M���?a)���Z��#�@���%"3�h��Ƙ~�|�D�O��K|D��'�|j@L�`4T��:�4T`$�^�'u�PH���H�B�����7U�&��� ��npQ�T�'�O��}�p�ٝW'��Zc�V
}5�t�3�N|�<!��ϋ�R)���e�4�w��o�|�L<a�+t�`ı�I� b0�R6N�<��QZ���'��?a�7��O����OZ,��٦P�ƌ(�.?"����w�#wgV�D,�|Fxrl,.��šݦ{a����J>?���)�����)I�$����{�����..2.z��IQ�S��?��KQx�:�Q�k�(��Fl|�<�7��%��Y+�� @�hUx�t�'P�#=�Ok��S߲Cւ`C�΀l�B�'���ƨ*&����'a�'H�$h��i��q���*����,2��Q7���~"�%��>	�I�*\�i�6�F-<�p3�E\Q?�`�Nox���Q���h&�C6�ƃ�BK����X0��O�����K��J&�ַ 1�T"r�#D��g�-U����NوB*���p#���HO>�bmÏ�M;U��-R����u�0q�l��h��?����?��'�Hi���?��O��ܸ��?)A�C�9�b	�Ċ�*�Xܪ���P8���-�<yU���	�!kW�0*�}�i�H8������ON�DA�t�����/'Hi���n!�9R��``.�p��V AN�!򤓆"�����f��w
Hk`�2���v�_<�Ak��ih��'��Ӏ
���Â6ȴ��ʟy=��4/���I㟘�%��ٟ��<�O��=!P�݌T+>�bi�5zcx�P��d��?Yaw�	.���@��	�B�le��+�B;�H�	l�O���"#NM.v^}*n^j�
�'�D�a��;ײ@h%��M����W&�'�x�Q��?x���`ʹ>W�T��'Z2Y�D�o��d�O��'}3��Iן���'W2����1�|��2#���PlH���$?e,I+@h�R��|����&*h�h�l�-hWp�j���,Hhh�fK�d�*]��:vd��S��?�@P'g�t���K)X�>�#��O+uR�������h���̵�G�L�y?�@�vmҍ�y"��x�zc�BԚl��%eν�OZ1FzʟƬ��JO�G�VAˀhV9w������OX�DF���`i�O��D�OD�$��{�Ӽ{ Cs"f����'E>T���!Vi?���U���K
�F�����]H��D�U�j��^�%cC(���=Q�'�j�M՚$:��iW����?9�ۤ�?i���?�gyR�'��ICf�`����f�c����B�ɆxSƵB3�U�T���L5��s���?��?!�X�`qD�yr�K(_p�s��D�<q�/�id$���'��<�Cz�<�+S� Q�!ci�2N�5��t�<I�&��l�����Dʌ���&�h�<�&� ���$��41~�i�/�`�<Q��0���R��цP��P��!�_�<	b��v�$m�@�B/�n�zPe�[�<!�b�M @J!G��g
�U*R�M\�< gZ=�V`�'ȃ-YA2T�Jt�<� ��P��,��iF��:�x4y2"O�Q�S��G"�DJ�J;�̈�"O65�ch[� i�F�!x����F"Ov 	��?xŶ��$ٻ#��"O���g[,�ր#���#ڮ�;�"O4H�*�}���P�b׸0��(p"O�H��߁' ��3�hɘ��Ё"O�(kb�6G	ڕ�&�J��"O�d���ŏL�A�&�q�2$�6"O��;��T�i��NPe�aK�"OLz��*r����1(H�.T�ٰ3"O�4!&̜u�A�R�N��u"O�T s��PnY�'( .P��"O��i���PĮɰ�B�o�Ġ�"O��c���}6ֹ!�ʻX3���"Ot�c�Y Z(�8�&yz,P��"OR]� )܈ST(�ԮٻU���r"O��S�I�*l�Ɛr#Ӑ�*+�"O�<����#A���XfK-6)3�"O��s2�XM��!�	� ��F"O�H�'�io�b�&���%"O�IW�"k��)�bL~�@8�#"Of��$d DriF��(@_��B"O�A33�بS�DxI3��%fJ�M�`"O�Aӄ�*uTy�#�'Q_<� ��'W,�`�'�b=�vJ�$~��K���*�<h�'�%f�x��#�V�s�ƍK��$�h��#~5��Yl\܁BCָ"J�_c�<Y�I��6:Txa���`�+�Hw��K�BG�S�O�y ���IfP:` D��P��"O
ݒ2m�/U4�1��E8@��ȡ^�(���h�L���2�j��𣅑W�TE��I9�ODe�I��8#T��6�:��3�P��"O��cÒ�P^� "`M3m�쁶��8>���D�^�	ɖ�(�F�>ҭSRǝ��y�B<
�ؘ8aϫ.Ƞ�Ff<����k��H�X�'O�JXT��AL !�:���"O���7Ɛ.Z6d��E�O��p�"OJ&�B� G^�;��]�ٴYc�"O��2Dm��F�XP%� 2u(�Yd"OB�:s%����j§ l�D��"OFS��qu^[GM/UZ�(��"O��:��~u�p���P�NF|!�"O��W ����U��4{0zt�V"O��aq�@!~��ʴ�W�E|�"O�|����"O�C��7-u��'�,=��	D�$�'����Y� .N\Idhz�^��
�'<�!"Jd ��pcł�ِ$��{;�x�` K&AP����sL��
=}7x-�IZ1�!�d�OŬـ�g�G&�Tbh��W�f�Ԝ>�D�*_��>�O>y��GX��P�B��ݞ�Ve�v
O,|�@T�(�z\zE�F�,а�h��6T5ʒ�Ƨ�0?�BH�J���F�N�B���2�`CW8���G�?�����c�H�F��cVmS�rs�5�&#%D����Ȼ"6]ȓ�N8S��y���!}'؟t��'A>�⩞���<�W�1=x��c��?D���j�i˚��4I՛� ���Qz���'-|Av��a�g�ɾ"�~Q�����^��Xy��+^�<C�I�W�P�ȥ���s�� �?$����F	��X\xx7�'�.X���U|j��(�-<(��Z�A	|��'��I�7.��r�B
L�BI.m��'����G���X�F��	�֬��'NX�(3%GD��q&,�5-|��
�'��a�d�
>4aH�
�*�3O21��� j��g�w�j;�1.P��9�"O��!��'tαJ� �&�Y$]���T@8��k��Я[�RՑ���\TQ@H;�O��&����� �&���$ �*�ޡy��4D��+�Oˀ9���U.�x'��a��4�V\�h$G۠yI��Q&�88���l���j�AO�o~ ��Z�b�=�ȓ7BE�4	@)1���)p������y'LH&)[���F�B'-e����#}λ `Tk�gQ�ao,��Ui�g,Їȓn�|�VF]�
�r��/¢f(HH����)A%Du�&�=o:�-i����|PJ$�A��\r ��*[ε�p2����X؁�w��$��)�gO�Q>(�Dh4xdj�1s"ߠr��%a蓂�|B�J�T�~Qd�Ĥ0��)HRcS��O�mi��ҥiP�)���	�vPQ��ֆ��eP�Kqj���%��$����1J��y2����JB햅W`���"� k��P�D�X+w	F1X�*�*6�`��~7* H3�E)2�K,=�8T�ǆ�s�<���K$U��9�#��Ie(�P�˄�*�ER犔�2(�V�Zu�L��S5.H8�%��1)���S�S��C���)��E��W�<Ա�Ǥ9lO8�H���
V55H�n�D��l�0 `BH���T�Ɂ@V�	�	B!f`k��X�F�>	(6���a��?㤰�6��K�i�$�s�.T��X�8�N��}���m��Q^���f˰}B��[*����+�f�j��4P�����}AGf�4s��4!��-y�8	J*�'��H0qB\3RN�А��c�+�74�6H1s�x�2������Z(Yb�� ��~}��X"OzS$:Q���BҤ�Y��s�W�<�K�>��'�Ҡ�C�D�ꑚ��q'kL	�nߨLx��)ezn�ʶ ����d��ɭYE�uK�L]�P���*8�<�kf�w����ʉ���=^�D�;�
g��ၶ�cQ�+���2>��Z�ƅ�}��T�"�I�p9 �$�T3sK�]�7`;W��O�zĝ�u`�ڥ��
Q���A�w��8YSƋ�p>��%������
�'�|�(d��N��}�D�?}-�x����Q��ϻE`C�`Ǚ4��C���F����iw8QU�})%�v�b�t�r�	c*�A�'��dWna�P���5�4p}U ω�i�5��+πY�Z��퉂&p�4�O+2`�����>N�p	7Ț���DD��?��G�`��pᅤ�;x�D�+�ɂ^�'f��ZdBܘl��Bu�n�m���e�M��5����qY�$Ӂ���	"u�x����W]����.��!PS����?1��	9K��@@�#Q��3����f*�32r���W�b���a���?E��w#tM�3�Ɲk���b��w�� �'�TX�w���Z�I�S�t))@D���?��f�$!^:T2E����t��v�'aF(����=L�JHr��ɗ��b�̾�j�� �p�y�	}��LCqI+^����mܘ��c �T$����>FL� �_��u�
�k �Xcp#�|���	@9l>�Q���O���\&��{ bQ#�"J4�T�#!�Iy���5
O�^��3DCȜC՘ՓS��#�e�Ag����;P��(��n��#��]k���t<`��G��w�!���z�ؙ�bj�C�P����V�n0�Ӆ�9h&�	3��.p|0hQџ�"=I��:�f<0�Mf�8
uX�����\�T|�9�Ŧ
_)�j3B@ �"Y�"��쪠��'1��YPˍ)<e���c\���$֔}�j�3����B�zM�N?�
�)P�z�l�g�y�P�B&F�p$��=��i�&Ќ ���sJM�0�L0̓��
^,��;�.O8 ��gyJ?A9ڨ1$�Qw�RM�K��#D�$�% 	1T4���<6��h�2�L2��DM�5��'�؉��9O�K�N��I���`v��Sa@	�(�"iᥬ�0�a~R`' ��'�I�_��R��K7[A�zu��5��D�o]l��-JV|�pV�G  �g~���%�� ���.N|!0ԇS��(O8���e�"����| 2Џ�?-c�&2��V-��M��W�YF�ڡc)S-]�ə�A ��<�aFG��j *�2����Ǟ�{�v�cp�ݍF B�)�ɹ������'�������L:&��Y͜<07$X1Qpb���44��ItFU%v�~0��(�h"��"S*��T����� �Dt"��<2��"�r%B�]����������(K4�<�2DB���7���m����@�F!<���yA(��_n��	`/Xz?-��`���7��$*v��K@��+��L<a�	I�+Ҵx�V���}�F�B��$��M�e~b�P�h�> tM�6S�y�����?���M�5*�jk�9[�R���*���#b裲.��50�Xtf���<ģ�;g�)��Y�A����.�/��q�@� ?���0;hb"��i�1Fy��Z
!�`H7�^�6�i�'cۮ��D�<�(��v�
��� �,P���R��ȃ����kG�� A1r"���O��_)d���qӆ�b�i��t�����#5)f�����-ғXe��JA�N[Jt���4s�|����_�(`�{1f�I��#�I�4RZ����|"�Y��~+̫qS�M���|�9Od��%�� 
I8���G:T�Iӝ>!��L# �t�P���s=$�@)4�@�>ɔ�B3<#�`.V���IQB�7��eHR�	�Q�0T�E�ͽT��|���'��2	�1�f�aR�&�13�^�a !d`�>b�Zas��q8�`����8=��g��PbpB��ka}H�5(��Bq":^������o~>a��ύP�2��D�0���N���0��,Z�At
��` 3^���EM,�/Ĳ%Yħ�N�1���T�1��$
�t��Hܬ�  �),`��\!�\���d́��.�D  }2�׮����̆�v쥃W&Z��~r�<c>T�k�/�rQ����cG-2�n�qbKT�Bv��'�<E�i�.�8����G�4��T�C �xr�ʛ?[={ B�_8���EB^<i��b��Q#r� ;��đR� b���Df�x��Ij$�臠
�;1���*�;.L���I+~L�@��֢�@ ���^�{� ��u�:�x�ϓ;} ��q
�zrx�pg�_�&tK!�;�-���X����7�Z]ht��gѿ/�@|�6�ɏ:��+�DO<p�@ł@��`S�x�O>�DQ�x�'�L3}q�T�~�
J������jؒ����ʯ\l�(�O�i�'��[9؝SBI[�x�UK�R��X��SbVM��0��%��mB�9�D��o?Y�&�.�
�k4�6LO�\�`�	��0*�@#"���B�
ܥ_����$�B� `�!L%J|*�$S�X�J�ݧs��KA�ۇ!�$`w�/n��C�ɂ=�~m ����%h��[�� غ4����$��N��5�>���[�L�nM@$����(O�}�
	�2�c7m^�YW�`A��'FEhGnۜx3��Æ�ՕV�
&ʀ*j |{��Y�F}�xK�-^� 2���җ7	�|��|%p�IR��&76�C�K��Ov��\�|A���{��qР��&4��O���J�2/�� �Rtܴ�a�'g��Q�7x6����O?g�jh�wΌ�z�o�/=��q"��&�?E��w�"L!&��>q(=3ĄO�� �'��Âձb!��R�/�&�;�(Y�z�X)��k�N)�`B�����I�mX��@ˆw8@Q����*�C䉗/�J�#cֶ��S�IM�+��C�I&@���;2(��SJ�t�V.W2r��C�IR�d�"@P�z��Q)W,JB0B�I4���
&�ѕ*�rE�q��yG�B�ə� �9�a!��R��։:��C��t�\�k�����Վy��C�I��$a�!i���sP�ߑHӀC䉀e?��A5
��{�p�����}�~C�I�*na�GnЖ̈Y�A�4`�|C�I�}֤1�s�ȧR�z���;
n�C�I#	N���	��}����Qo�0pw�C�ɏϞ�qp��ip�����&Q�C䉶� 0ä >.Vu9��O+jC�0���RN_�wRR���n:C�	#&�`RO�.�i$MT�/�C䉶�� 2��R-"!2�o�(V*�B�I�2o��c��\%�I��I"�B�ɺ$�8�0٨[�h�M�&)��B�� X��A�ER[��"�B�(Z�JC�	-0�9AVc�0P��{5酝Wl�C�	4p�U��җr��@X��ŽeO�C䉻l����7!H$��	�%0�B�	���giդs�z�� ՚.��B��: X�UI<�� �gH�c�>C��"|p��#���Is�[�!4�C䉃l��Ať�
�xHQOx!P�9D�� ��x��@���	_��Q��=D�`�U���d�)��V%e�8���n0D��{�e�\e|H���*�2y�)D��� P4=�}�U'�+ЫT�:D���AO
$P 3��l�BQSE;D���b�������,d�tQ'�9D� �Q��Zfm�a��D-T��(S���V�v�0��N|�숈&"O� $5��52��%�7�@e�~Q�""O�%x-�-A�M���Ĥn���A4"O�	�@R@&��{���q��Ś�"O!*��,=�HM!R� Lp�,�4"OY��e��%��!s�)�%=Sn��"OơhbJƯF9�LjT�E�I@�APC"O�,Z�%J�q��@+����:����"OvTX���(�0X06_�9 �p9S"O��r�mF�d�!�a�V� ��"O.ݲG�
:N!s�e�0r�*G"O\���M�+�(L�s��:]0��Q"O�x�aѦ_p��H�cNR�@"O�C5���S�ؼ7KD�Y��� �y�lÔz��b��?*wn��3�I8�y"��0)$�ҮB<�2)��A��y�fS�r�@!�(tH��a%��y���LQ�]��L�%c���R!K
�y��;�H��O/c���s�H'�y2�
�?��}��)�8	����+ٜ�y҅��#��2����
 )��b
�y���+F1�M�R']i(�'��+�y��Q1+�d��,�(p�6�zD���y����
�@ۡe�f 4�R��yCI"
(�Bg� LL��SS�W�y�H���z	�s'0�#�j���y��	!�\�	�z�����y"G��$�6�S�YH �A ϱ�yR	�2)���pc�:O X&��y�E�Q/�5�G���F���bD杋�y��<qD�a�
<I�%R���y�Jˆ{�Uh�gO�.��ʤ�V�y"/��
X Ļ��7YE�\���Ǿ�y�I{-�-���E&����#��y"י)�\<x1�P8KR����?�y�Q�kT"=BE@�D�d��-Y��y�G��7i*p���;&8�z�iڨ�y�;9JP�0��9uPM
å��y"��KP�脨���ҸA�",�y"�8����Rc�" �n�x�k��y �/$t$��A�s��	:�ڒ�y"/�61�H���kc$P���(�Py"�K� �Ǫ�/J�N�1�'H]�<)�)�&!v��c���T��Y�<y' �jO6�a�V�$
�/�V�<YS�M�P	И2X6�Xգ����B�	4t�EI��	qV8�ĭ(r�C�	� bx�� �d���h�Ǟi�C䉿d�f����
�u�@1ʱi��B�I7؆9�rㆶu�$RC���(��C䉻v����委�g�|"�����C�ɁPa̼��E+NU|� %��/SB�C�I�wی)C��G
���CSq�B��B���J�w6<�tO�3��C�I�z��Y1Ո�<�F�i�	�?&��C�0�L,�F$�|!���Q8q��C� j\< s�R�s�8�r����\��C�I+����fX-T�"d��^{�B�	���q��+'��xg��Z��B�� x<�ݢ�
HɞՃG�\�, 4C䉖����C֥z�<���X���C䉒N�>ݢ���L�x}�6$�Ka�C�	`���K=oT����i��C�IY�l��Õ6N�xe[c�I1�B�	6"�M�P�_��
h��Q�30�B�)� &�Qq燒3ǰ�`�L�=��"O�hT�E1N0ȋ��Ӈ+�F=!"Of�XS�\-�p�Gm�{���3"O�`Y���T�R��T�U�55�Y�"O��q��O4��:D�D�<*!X"O~X��#ܖ7�l��� U��c"O�Iz5���\��Mؖ՚1	�"Ob<� )��	V��5d�T�+"O�r��1+;�ɐA6 �4�"Op��A��I]F5)���w�Z��"O�Y�D�������D� x���f"OFe���V>��q�Cd�$P��X�"O�\i#Z�{ކ!{ い��� t"OBtH�D�	=EB1��R�-V%�@"OHӆ�X9;ȁ�SBҙ�N��"O�)�jT� t>���o�0�H��""O�M`�ePZ��`+�GI {�Π@1"Ot ڧ��2$�(�B�	G{���"O>%s�թ�bI)6E��|p(`��"OJ]�ƥN�7��b��ZvV�P`"O(�����'�>Ѹ7h9��"Op��r)$h���4�B@Tܙ�0"O��D(�2�~!��]�.�@�j�"O��BP�)$�b9ТY)z��h�"O:�p�d¾*�d�O-p_T`��"O%��dΰ\%v͉R��+&��k"O����� >�y0�h��P�"O��h2�"rV�`h�7\m��"O`��-t�AGi�(D�C`"O����B�[� 5��g���i�"Oک ���(�k0H^�Ob�}h�"O��æi��oQ2ё����iT���&"O�(��	�^Ö���'.7(��"O޼9� 2*wm#$��\R�lZ&"O ���Y*F�8*�p��#W>/!�$�pjp���W�'��4"V�K!�dU�YXL��Fh�^x!&�G�k!�d���,頴�I�m=.� 2a�-!��	�1n�����.#�`����\y�!�D���,��O��M\d�r�gC2+�!�Ā~΅���ؠ\��\�P	T x!�+IBjh�OG"2�L= 7V�g!���8�,��ػ]�L��f���!��	rڹ�$Hy@�Z�Ɣ)g�!�DGA��S�K.iX� ��+�!�H�p��w,�+[H\s�E�L�!�d��j ���`Æ�>�Q��	�5I�!򤘿IZ�Q �>$4}sF��!�\�u��Ti���Pdjaб���!��f����)�;f�p���Ţ?s!�D��	5F�	@�B�q̤�[��B�eQ�\F��oLM�y�תɤ0���(c�Q%�y��8r@i�� ��!Y���S��
�y"O��.����Y &L<��`T��y��s�0J!�]!f��bG��y� B�Q�,�����Z:�\ؓ�)�yr��
�$	R�ەi�`p�o��y�E�>!�b\�@�%\�~<T�S�y�@ ~�1a�-��`�Ҡڀ���y�,:~dH$���`'`��pkX��yS�B(�T�1C�+Q�4���/��y���"�-e`I����+�'��'w�{��/R�Ja�EL*�p�`S#�(O�5����0��Ԁ����L�pGl�1#�C�)� �]�GLD�J:<A�,����b�(A�Q�"~�	8f�&=H�bQ�y�����D�� C�	\7�T�����B~�}j�N�<r��I�,a~B��Ccd�P�ʏz�+��3�yBEͅ?��p��J�!X�c�"���y2"�!HH"�L٢)/��+"4�yT�&E&yvJ�o�f|���܄�y�82'B9���>:� ��0K�'�p?��OJ�A!F�sl�����`�n@�%"O$X3t �2�r,�`��>�Y0"O��cE�H61^TR�K��o���"O�q9��F�J���D�	� w"O�H����i�����P����%!�d\'p�D���@�5Ɣ|�7�	�0C�	 �$h��D�m���2x��B�I3Y�.��
�	\���D�\�B��! (���E?h)v��W�A�-�FB�	�bJ�mb��Ń}�����:*0FB�Cg�q�V.�4��b �F^<ʓ�0?q���6o��A��(ܶqk�� W��}�<���%c����D��5
srI ���B�<�䂚�ĩp�ЩI*� 6G~�<�HJ>yp}��g��o��d�Fg\}�<�L�:��y�IH�	��Y�fFr��@���O�8�F��xv��<V6xY�'S,��E$Kv,�	�#͆QY�!�'�8%@%�Q/�����X�=e����'s���&kʾ"K�0���@�6�*��'���6�ԍ4ْUI6�($���
�'�ڭԃ]*:�2�;�̅3.z�
�'�X%C4��'�$x��C,y�Ȋ
�'�t�����0K��u`�>?h��	�'���4N1L��;��5k>��	�'J�D��ŵ(�� ��}V�9�
�'��[R�ҝ�f���J��G��K�'������!q�BQ-����h�'ܸl � ړ�F�$L�#�Jm�
�'�&"qe�P��!����
ˊ�p
�'	e‮)1@$���6�n�	�'d<�i�Q+.8!�S`-
�'!�
3��	V� "�XK�c�'	d����5Y�d��g M�%zn���'(Vp�F���_(m#� F%x�%Y	�'�����$aE���F��'�ڰ˚�OY����ͅw�8|p�'ȎX#�J�ZN������s�*�'$��Rb\"fA!�%@n�mQ
�'��a�5k�.p��B�3f#�i`	�'4j��e�q^ ��s���M��T��' h40�M�y���3�ʆ��=�'-�܈'/.'���@N�=
��ɹ�'l xw������Ǉ�4BS�'k@�ЃOj��8��oƮ~22l+�'�}�tcbk:@��1	�'Y�(
&��P�m#�[7�T��'ON@y��Y�J������&UĤ��' t�
��(*E+�#ٮ	�$��'L�=��o[��y�1�W�zH�	�'�6��1�9k.�1FK����'+,|�拊-��@s�ė�y����'�qi���b�`��$��
I��k�'xT1�T78�h�SM�u�R���'�X��i�&G5�Q;\0?���[�'�, �h�	`&0xAC�-a�5���� L ��'�y�yCա݃Gbi�"O��{�D�]����� ��x��\�s"O����H ��1pc �>|�ʘ�v"O��Q"�� ��Ab��:	����@"Oޭ1�� �>0�$EW�a}4k"OH䩓�ԇCb�`��$РLn�M�"O���a#C�"V�铡��t��c�"O���OXZ9��������"O0h*w��%s��k�X��(�"O�I&�ˠdi"����fy���G"OMb-c0~�A% \�x�Ap�"O���C��h��&o�12P"O�ɹ��V�Z�� a�>+��"O�y,�8۴@�OJ(  <�D"Of#�*�7��=w��n��1"O�x)�F�|��d��,M����#"O�,(�5p��%��f�$9A"O��ʧg�0�}�b�0�i�"O�Ak"Q5̝�R"/$"�]�"O,%��#�5&2X���U�����"O�,"6h��
�D�4�ݓ��0�s"O�Dbd�]�k�����䋧�x��"O�lZ�o�!�lX��É�B�D��"O�,�w��5�`��=f��#"Ol�
�D�v���6��k�<�C"O�9��G�o�Xh�LD��L��"O&�ӕ�7E,` �M�c���2*O�yo_*EV���,�-s.mS�'�XAJd"g|�PBBf�Z�Xm��'3�)�u��W���a%R�i'����'�&��=y���RFm� o\���'C}ұ��E���f�R��i��'�:*udO<2��hiՍ�	;W$�	
�'}"��ҪХ)��P����e�h��'��@ku+ڦ▴�p�]�S�$t��'��5C#*��%����䌉tQ�L�'�fPaB	��hȎD��Bk���	�'iT�:b,ڲw&\��e�g�lM��':���`[�#�L�s ��W��i��'�z}b�!Ni��@��!O��s�'����
�`qV��i�\t���4S�ϊMx����%' d��ȓ+̂��F��?��[�LE\��ȓf�R�{�� н+�`J|.0]��@���ش�I�0/�K�>X� ��ȓyg�-�DH�^�8���Q�z�R��P�X
Fn��P@��)�4Zcn��ȓT(��E�'r�F1Z���/I��$��I@e�ԧɴ;��=���!P����ȓm����(MM:y93�ٖ7���j�j��GIR�50N\1�={�܆�U��};Yq�έ7*b�
�r"O���5��`�DӤ@%^��"OP��ǃ�g�V�۲��v/���"O���I���S�K�M+ظ(r"O�T��o�N�A�!�@z���C"O -B0nX�9�Z�B(�G�<1+!"O�U�� �}�Iq4iJ�9�ڬXQ"O��3��
u�x ���@ɉ2"O����L��i����H� ��3�"Oe�a��ry:���{��3"O�HP��^�8��)��X���B"O����Ն\��3�F�����)D"O	X$�K%bn�`w杰W���p"O� v�z�V�e���r��//��˔"O2\�b�B�l|np!��Ǽ �9��"O�QQ�NQ���x�m&�b�8�"O����I��B3p�p5��S�� �"OD�J�,�6)8d�P1I�1����"O��r�90����G�D��a�"O(����S�t�GX@=��s�"O�؉}���D�2J��P1"O��1����rjĤ�I��"��"O�����fά�*�IӗX�u�s"O��q�F�Άt�!#%)y洺�"Ox��&#)ڌ�+� Z>B^��"O���f��B�Y���Z�BȚQ"O������9}T�4JߑB���H�"O^L�������W�XQ"O@	�Tn�+q�P��W�<SmQ"Oz��rk�C���Bgf]�;E���"O<�(��
�o��0SÅ�3��m"�"OxC6�ˡ�F����j
}�Q"O�p����h�4��Ȅ5id�y�"OЙ�G�ծO�Q�GKHX�-�G"O�xu�H�8 "���	LT�,p2"O��P���-Y6��� k��B52��s"O��U�B'h�5��ԓu����"OX#�G�"b����
N��f"O��H4�8n�>��na��� "O�ѫ��Ȁ{���᳈A,	U�d+�"O�xQ$�GU���Q� �*z8��a�"OF�ZGڥ& �����!)���p"Ox���*l�#���,Li�=�ŏ��y��_rT3!�S6�5! a�/�y�� ���5˞:1iF]�W#
"�y�I@���]aU�Ξ740�+�T-�yR�B���t ׭@,5V�X0���y�(s�ȑ����0]DJ�m��-]!��o�zUٵ��,8�(��U�_�O!�d��&�piB��M7w��Uc�E`F!�䆠lĲlQ'�d�r��um?l�!�M�T���r&�$\���lފ0�!�n�X9�'ǢK��A���L�!���~�0<�FG>a���x!�M�^�!�$/7�
�� �bY�ԊW8?�!�DY�V�,�wc]�<�J�0A�c!���4�
|94�A=:y�<�@�̸u!�$��
8d8�-ס��m�uĞ�5�!�ƌc��4�O�,G��$�TF�$e~!��ڻ�h�	d�����i�p�rR!�dA:��j�a�1o�hc�tJ!�dB�<Tfc&���VN�i4b�^�!�D�$3�p��kC�h�d�p�ߵaa!��C{c���"Q9B�H��Sa�FX!�$�V�0	A�����X���hR!�d_�+�v��ɭKnq�)Z+R!򄘀xk���Ə/aJ�8��	;K!�(0�T��TBf�H��4P!�!Z�vh�`�/3E`�!�M!�d�6?�mh�C�'VR>�#%`��Jcў����p1�"B���j��X�ou�B��1!t�<��݆�P��R�=D C�	�8��h��A:Z�&h1��P�q�C�	� 4�%ŉ]���r�P(z,C�ɮ�jeyU��,Uy��!��O� �C�	�A����ړ%�,Mh�ڍMC�	m�b`�3/�d��`��QTC�)� @�6h��4q<��w�1�D��"O�Ѡj����H��'x��\U"Oΰ��	C�O�Zp�ɘ�h�^I0�"Oعh6Û�i��%H@Y��Hu"OT٨s� l�JX�Ag�\�U�U"O�h�F��8jt�S낶]WDX� "O8C��+�Bv�ϗ!�����	U�O��j��B�A)`�y�@�. ����'�9I�A-+a
M��ψ�T虃	�'�5� ��[����,g���K�'�؉3bfO*/���:�.6x$+�'�&My��E��!��(�^�C	�'%�A!&�,$�͢!�3����'W���I+.�aT�MUL�-Ox�=E��k�9]L ��G�4}��@�-C�!�I	����� %������ށ }!��!B����Nʝ:{�4K��>#s!��+N��4�@�=�J��g"�/!�d1X����n3fð�OO�O�!�$��ji������t/1R��}���Y�T���֍Y�`���҃�!�I^x���6�U�>�y��U
L���S��|�<���
/u�f�X� \�����*�]�<Q�"���4P9� �|"��AT,\�<����)H ��{$f	l�Xg�[�<����`��e1գM>t�08MS�<�)׈N)R,h� �{����PJ�<�1j�1hT"�3"��e^$���DMh<1%�՟K)����HS�Y��L���W-�y���V\�x�@IB^�8+w$�,�y�97V.�ʁ�Eq�:���*�y��]�3ǐ>j{|����#�y"�׫�Jq�@��_2`=���	��y�n[�'����F	*E��5�$��=�y�F����}����&px4`5��"�y�m�	u/p�SÎ�qל��D��yB�05�$ɓ�*�!�bA!e�O��y"�:	�U��D�pMf=�5���y2F�O�š�l��b�z�����y�����
��#�=j�x�������y"��-'�:�@c G4`ЅBd�3�yB�ЧE���2� }0;��KC~T�`�'�ў,R7$U*X�KE=i�p��%LP�<���_�%�@����D�l^�+�(�v�<yQiC�&Ô(���3@�jX��,�k�<9�m�'?�4�9E&�- Jf��`ˑc�<�#i�?#<�[UI �:X���[�<IS�z�<9�@�n���6H}�<��c�jq��#��!q�SF��O�<f����d)B��0a���t�Xu�<9���q������Ͼ~�ʗ\�B�I�N�š�dSe���-��D�JB�	�9 Z����"����R�y"��c�Z-�C#������y����ts�ȓ:*Ȩ�AG��hO��?�� źc���r&��	 �)۰g���<���؇(S|4 �I&u����2�݀'w!���~ �r�����!�KH�@�!��9{�H�r#�T [�.��AKm`!�D��n �k�������,޳Z�!�F"7����@$+����JK';�!�đ(j@�+%!�a��x���%Rq!�$EM��tL%��}���Ɵ?R!��R9&
X�d	�;n!�C��$C!�� 2��Oޏ�%ا␈d�� �"O��+�e7E�"�F���ف"O�C0�@q䁸�"�:���"O��a����6��P8���!c�L�S�"O���VgD�p�pt�䯙��܊�Of�;�S I> 	��K��N����4D����-0p�# ��"�5�.D�����%�z�B�M�2�t�Cql+D�d��ݎ��u@UXg�[�j(D�\�4%�.��j0h*d済���9D��a98RP�D*U���В9D��0u)�aG���򃄉Ђ�;�5�O��t���s�"7-~՛W@�Vp��'�ў�|��.��$.U���s��!��y�<�$n�ds����IՅ9�A1E,s�<�k��< ��E��%~� ƄMD�<���@*!Z<y��ѾT�(����RC�<�"4�b�m !2����'D�<�D��88�p8#!-���u�<��*B&aF�JF��U�Ҕ0p��m�<a�эi�f�@�%?��a�5��m�<��	\�) ���Rn�9e
>�pU+D�<I��m�|13ɷaBެ	u��{�<����J
��㭏3@���� J�x�<	BN�0E����
��%���Z1�Mr�<9��[�g_^q�P%� Q�B�Xo�<�r"ն���I�^�L8�����Rk�<��
;��
���0eޭfaTL�<�c���\kq/��t�)s��G�<���;W
���!��"K���e_L�<� B�:0r��D�y�$IB��K�<�����i��<��*;@����C��[�<)�̗�I�4%��iA�KJ�p�5n�B�<�uc܉iZ^�xs��
��y��A��P��|����$J"x��*�{a�t����gb!��B�ma>�QN�"�`:����!�$Υ�@!DM1j����7A�*e�!�Đ�L����A�d�@��ʰY�!�$zZV H0N�]�F	��
�g�!��I F.Ĺ2�;G��Y �l�!�T����B�B~���d������q��(��I����/0]�f��(3�#W"O|}h�"�.n���ˣN�G"O��3ת\5���Q	B��!��"O2CA��B)�!�W��չD"On�b��E
$����`º�ҭ�f"O,H�ak&ܘ0+�֎�Ds�"O�Tː)M�:�
��Fk_%@�pEh��'�2�|���j���b��A��f�ɺ��1D����Ά�xs���JP2O^5�b:D���L9c/��У�M~�F:A=D��9FLQ�lU� ˓��ehq->D��TΛ�.� ��Ɣ�v��Q�V�)D�� �,���x��S�^�"=��:D�pY&�V8D�B��a��Q�I,D�:pD�9��F�N�/��I�v#,D���A����S	ͼsn��a�+D�X�"���r���JI�ePr�K.D���L^ E\ly��j�H���?D� ��dǿ�*EK��R9?�:�`��3D��hmL3/(TsG�33��ӡ14���Ge	�Z�1�o�i��ey�$E\�<	bl�=:�9K�BU�s#�ei�X�<y�F�t}�h�Ż

���WI�<� ��c�XO��;&��3φ��%"O�4��HV+�p��.H6��uxb"O��7
��l��C����.�8A"O~��&�� ��X-W�}J�@�"Ol�	��K�l�A�B�M1��"O������f<�d#5
�%�t�A"O�AP�bC��ĵb����Xz*�p�"ODZ���/N:� BnJ+6�T<i"O`��AHΚN ��f��Pe��"O��@蒜X萉Մ�7J�<�Z"Ou�!CH����cׂ^�,(�"Oj��c�X��zع�,G>�@��"O�e���3:ΐ�����<�$	�"O����>~x�� ڞX��V"Oȍ�0��)���{Ah�QT�1"O��зό
�>a����NضHyG"O:�X嬈� ��%`di�ةu"O��3!�\�s(.�B��K�:�&�15"O:��T��%�A�6�J~P�XQ"O�xrl����+�
`�{e"OD��fꗘ\�lX@"��#PZ�I�"O��:d�.L\����Z�L�b"On@1�� � 1X�Ц�)`���1"O�U�H�Ӽ��c+)BF�ӥ"OjyabY%��r��J/ ��B"O� ����~=V��`f�s"O���7�
�+�d�f&kZ��I�"O�SWnE6�F����C�8c��ag"O�ᒳ�Җ\Z�����]�hn����"Omڔg��Vt�2��/0X�zd"O���CᏙ4�ڹ9'��x�|��"O�$���1B��!���o�`�"OtpP�o,/��q����$bt�2��'�!�&zװi:��#s*��I���Dw!�D\g ���aW�=�|P厇,Zi!�$�!����HJ4C6�)�Z�a!�dܜR)	݇��@իT�mP!�$W=M��Wn�e�]�
�.C!�$�$z%Q h��N����=�y2቞��z��_X�n�ʥ`I� 3��d-��zq	���x(���,�l�	@�,D���L�D�>]�g�P�,��a/D���q�]d��(5C$4�6�#�d'D���fmG�-bSE�0}%�US�B9D��Ã$Q���A�	Sy�mb-7D���p�"X~m�µO��-b�d5D�0���;3T���`iJ�m[��d9D�a���.X�����:EP�]���;D���*�Dm�=�#��$��8	�,/D����/޻m�&|j�iE�h ��"ag7D����^6��P/��Jz|�`A�5D��s&��g<�|�T钷"�hl�b�4D���TD���������o*�F.6D����%T�9N�4��u�D(D��t��<�5j�@�5���%D���Bo��)�2�P�L¥;K��!�#D�4��W�����T�}0�!D��ӑ��*y&H���S# �|a���"D��pw�7{����G��h��d+D����L �~Ѩ�B&v\L���*D��4�|�6H"��߬h�z5�d)D�$�U)�+p"Y�w��h��Z�1D��i����l�����!8���ick#D�HcL�{���5���vC�q�."D�� ��Q��A2p�X�c	�g!���"O�@su��*fB�Ph�lV�zj�X�"O0xS��P=�v`B�쌓W�M��'�I�2<�]Cŧޜ^���1�Ƥp��C䉑>��)�΁�Dh=��J�#9�B�ɟy�v��& ��l��wL�7�C�I�&��X5���Z�ӓ U�&�C��%���ڰ�Ռ"��5���Fe�C䉼/y����)ϒ{�a+���	~�C�I�)E�(K��ʫ]蚘	��ŪR�B��AM��P� �w4����?��ȓX��a�Ucȓ3�DL�'!'Ȁ�ȓN]%�C�wA�lif�} x��ȓ&�P(����2kR��R"h��Fȅȓ+}��*� �,#WRtJf놊�q��o�A�CX�u&�	ʤ�F�c^���ȓ(��\S�B�LE��9��l�����REhX ��P��4�3lʂ	�����_i4ɘ"��Iލ�6��f�ȓ{9 X�IS�X�� �P�����Qv�0�&.;�qЂG[1�R�ȓK�|�
ϨV�� �HX�%�.��ȓG�[�*�\�R]pʜ1�>|��K̵Sv�� *���$�P�^l���	eR���cH�/��sC��U����;a��Yw�[�#T���n�R��ȓTLdQx�EK+�f��6��w�����E֢0kӄ�	Hʘ��a͹CEZ����tu@�K�h�|���Bb�t�<qr`��%���w��1&.)��LIY�<a6�����3%1_�|@����X���hO�'�х�"�t0
�)=���ȓ"V��`v��n�����#`��(��L�f�
w�Ƅ.�]s%d�B�t$�ȓvޭq ��,��Փ���
�����+$�|���ۨp��r�S'��ȓ}�d�"�N�>^��-��,��@��t�ȓS�2L�a���)���R��T����ȓ?�a�	go\|jp�%N0Ćȓ���D�+&�-�A_�aDꭆȓb�R���G���zqў8�
Շ�h؀yZ�@�	^<D�K ��/'��ke8#�A�?xnzB�.&��-�ȓ)�H��E@�D����'-f�ȓ9�Z-HC(�%z2g.�tw��?��q�zTψ�9��X����"�V����*���)*"���O�	��h��"O(�B5E]L�ҵ��<@{b"O>y�i�.����2Z�P�A"Oz�B��T7lL�<PP��N�`qb�"OthpQL5W�r�r0��%C�~���"O�Y�&�Įc��L��]�z0�"O ��4-��A2�!��jԆ*��Q"O��A ���5�B8�j��P��d:"O����<��9���)����"ODP ��5\����`)9���s"O��í��Z\�\a@훊�L9�4"O�ЗgTt@��!b�7r�`a#�"O�Y0"��/!V�c�1
P�H`�D%LO&�c�kE�e�Ι�E��k|
ݩP"O�Y��Ŕ�k�0�M�Q^��Q"O��#�RS��	��+^�g>*�*f"O<4j�%Q&f���xg�)S1����"OH�����#ؼ��c	�*.r��"O� ͪ�,�"��(�-�|B5qE"O^�A�L+�M�G�J쵃5"OD���"LD*1�"Jԫ%4��q"O��X�-�'m���Y ������"OB=� �$+D�c���6�0���"O�m� ^5;�`��	�B4��&"O��8��A-��ّm�|'�d�g"O�L�'g� :%D�3$lb.IР"O0��0�՞i5P\��X=x(p�"O�#�̙D���J�%K5��iD"O D�u���l�|L(%�A�t��1��"O�Ց4�/�B�ђ��B���"O���1���"�(Lɵ�B�ь԰t"O��C�@իbG2<�'f��d��9sw"O@4�O�ê�jG�3 ���jW"OJ�Չ�+K|�x�`�$T����"O�Y���n�tt��O��4���*OЅ�&�#�B=����@F
�P�'7����J���<�9�W
7Bt���)��	K��i���X'k��ͪ7���yr�R-mA�PC��
^���t���y����= 䏙؆��h���y��Y6^�l�
U�.n:��Zw%]���'�az"��3.�8Ԥ�lj��@���yr�Ll��{c��rb�s���y��ϐU�Aڃ ��Z�|�k�[��y��߶�Z�p��2X���9$L�?�yB@�5 ��R��&��)������y��V���R�#�
H7)%�y�)��
)�*Y��d� ͸�yrH�<ڞi��86�qHPNR��y�� d��q�����RW�V�y�f #s➱�c��J#�Έ�|С�d��hW�:s��	j\�L�ƨZ��!�b��kSD�k��=CĨ�$0�!�D
��V�@e
܈=��)HPI�6&!��y���QF�9.��p���T�!�D��T���+F�ׁP*�9StHҒ�!��j�{c���^���P��!���?8�nBp"W �p��3�]8mp!�DT�(ȸ�':�� 
���<b!�d�v���k�n�r��UQ��'F!�W�^2=(3��G�������%M_!��A�h�+t C�~�� �F�4�!�dː6�fu�e��
�v�bߧe!��X'`�Y[���k>��Bْz�!�d0Y���c��&TQ�!�`7[Z!�$�U�xIb!]�?�p�Wo�hJ!��CI:F��%�#6D��9�Ϟ�2A!�DQ\C�I�1��HAh��.Q�[�!�d�{�09(��ˡ(����/L�!���-*Ԍ��NH�w=hIA�.	�!�d	�K��xƃ[B�}�!��}!��0w+T��@OE+B��e�_m!�d�H�<Hf@�>{$��1V/�P!�����c�ѱ#@tX�Ue�w!�DA�a`%(��İq�P����
�!�$��=�$]���;7�"��j�}�!��ĊD��4$+K,�L�3�I#|!�d�v���ԅS��U�5B�Yh!򄌞!�8Aq�a�6z�-�↪?e!�>'��ɂRh���IJ!�;Z�5��
0$5��.�Q��'R��K�.H��	$��1������ z��@�� 6���*H,x(�"O>��e-��E��ŔIUK�"O0욆�M;7(8���%��bp#��'��x}����fQ5�l@��D�!�Y�:�n�և95�~��F'ȂK�!���5</֥`4���l�@���!�䓦8��}`����M�dɶ.-B�ɳ2�j�c5#Ȇ (^)1�ǈU8�O"���вh%^�C�'E4����'-�ў�ባ$F�J!�ҽ
�.�1��
�" �C�I�X���b"@(d\��b
�U�C�	��b��0��+g&�)"���C䉼
�����B�)f|�p�G���C�	3^�V}`+J2C�a�G&ˬC�	3Ƞ��& �%?Ԩє�ƌRo2�OV���J��$�0H�O�����U�!��`�)�pI�/"g��3ŏY�!��R���1&,�)����G/�1�!��Gl�<�B���24��&.�!�D��b��8�t2<v�5 C��g�!�
2(�긒7*�cFpp��Rm�!����Q"�@��`�DPe$K~�!������JB;I:zGd^�[�!�ĞJ),-�qA�iX���TP�!���1�|��F.�R�	E�u�!��'��X�t��`Zh����@�s�!�cRQZ���.JVf�J����fS!���V�=Z�� 1C�u�6!þ!��Q�R��1���*'`�@�&`!��LO�V	���R"D�����nT�5f!�D�oUB�i���*W������MJ!�Z�L�VNl�fT�cj�S9!�0�T��eLMˢ�ٰ�	�pJ!�$�s��8 "��.1=!���m���F�8�1k� m�&"O`��!,|��$�]Y���Z�ODk�$ؠC�@�;CkڴW �a"�ID��K�	ʪ%ۘ�2B���t�3O?D�ܙ�&Fs�� 䒒X3��꤃<D�����Zq�`��JѬ�<L
S�?D�Th���!�sgA� ^u�IC� D���C��c�8 ⃞4&Q�q8��?D� #@�._2t!���[�.�HZ��>�O(�MuB��֢�	�"��Q�*���@����@Ԉ4)�	 ���(	~��]�$A:D��93�Ѧ+�b��f�^QI��C	9D�옃	��/z�E�D�R02h*+D���C�,o���C/	x��J$@)D�,�bw<!��LM;R�2Y�d%D�*fo�;<����ʋa�@�)6o$�숟�4��o�	[���Po[?jL���'�ў"~���1{�$]Q���"j���DFT��y��&$|5�t�(_�E������y�G��)0���`(N{��F��y���3_M,�$�O6A��a&��yb��o݆ac�*��,;��	��y�L��4*pƃ(����4��y�H�3ll��0ņ����D��m�<a�h����k���RcL�U�<�����\t���́�)��a��!WU�<1���#����O�>b��� �T�<��.�[�&�i�����P��P�<Ƅ�)|њ9%��=�rM�B!O�<q�D��f�~�`��_�D����@�K�<� �pCЯ�
|��Ԋ� %%�
"O9'N T��5�&!N)��"OP���T)2��1�C�/U�ИR�"O�����4DDD`��L�����1"O`�JF��Բ0���ǎޮy�W"OZXS��պ+̝�	��(7 �	�'�e�T*٪SS�Ԉ$���bR�=�'8tla��P�%�f��W��
�'��C`H �R_�����f?XlP	�'�iX3ǆ�Os�h�b�H	�'�:99�O�/+ ����F ��m�	�'��(!�U�[��ب�K�����j	�'l0Ĩ��^*;�Y�����.R�s�'�$��Ơ�M�\��+R�/�x	�'ddU��$P��%Q5j#D0����'$�(Xf#��聤*�;B����'<�����	�F� \9���#7�I��'ⴥk��@�YE���`^0�^\��'���Wh,��1�k.N�1�'�v�0�넑@�ʹ��HֻD�$��'=�IȐ�= �\5Q���
�lR�'d P��v��� ��NrT�
�'���Ǐ��E� i��BI%t����'����b�"q��-�6�N�U����'�,D
\� �F�8��H�L�&��'��� ��_�a$EK���>6�k�'�8|���	S���eH��"�(�'/�Q�SDH閕��N��%��M	�'����Ddh�͈2�G�Gp�<0L>����'Q1O�L0����c���8�v"O
ЋgMN
�+�,����#"O��R��Zf�<���U"s��m5"O �����B�̕Q$_=�x��G"O�$"W�	65xV��#L9Mx*"O�%�f��;`��"�UgE��P"O�h�#)V�/ezpc7���P"O\]R�/Y+[�Eޥe^�"���)�S��ě&E��p�ڔOY�Jœr�!��%i^ j%J�o:�0!��%j!�֋Tf<\q���
�Z)	Ţ��TP!�K�Jd�t�qρM��઒�9m!�䈥��	3�*ׯ�`�!V��F�!�$ �F��=�f�\�F�<l�W�7U�'�ў�>�h�(/M��zFc?/K QzU�(D��[�Lяn<���/`c�苐�%D��bg�ǡ.���zŬ�p� &`'D�l�g��%i<�pg�#���#�9D����.X�9i#�̃P�ͪ�e8D�|�� ˗B���
F��c��V�-�!�ğ�C�|�;"��;��aw��~�'�ў�>q:�eZ�=�n1����)��	gb=D�(�3C]9'D�ԃō8
jZ|�1�:D��2��ڤ"���FH�8x�L�a�8D��+���?�f� �X��2T���6D�4�%�I�̀A�!F��l��?D���m\�f�*��VfՌ ?�Z�?D�����ԙR�i��G�"Y��`R�)�O���0�O��9�Ņ&`<���M
��"O�Qȗ��xP���@$ߞ���(1"OTT`!�Z�,�� 4*�>4�P�0&"OZ�h��>R�������iU��`"O5)C ��^lz ���i�Z!�R"O�ˡn͍O��u�P��V��q"�"OH9��0�P��!,l.z�P�"O� �5�ń��8�:4h�H�KfLq�"Oh1�UC�����Y��p"O$���hC�(@�f�u^(��R"O2������dF����P1m�$��"O�V�<.�aC2X�,#T"OPU�%d�@��K@��	@L�$�e"O�����;oQ���ȵX*�� "O��Kߊv<�`{'�ǋ=$I�"O6�c�-N�^�nq��H �Č�F�|��'��P2j��:���7��r�p��'��pJ6��97L��D�g��}�'N��i�C�f�j')O�b̌X
�'�t�"��^>vX�f�ߟ*.���	�')�����t�L����.q榱�"O<�QWI�d̰��K����v�'�1O$YQ�M�.� �4ǋ)}� AS"O�t�w�P#I�Ա���\��,��"O�l�B��=�D�Bd��q���"O�0�c!G1*��@��#Ъ�.�y"j�.�ZL!%��3_k�����y���/Lh��d��_�4#�����D7ړ�O��8pC_&z��3��3o�hݡ�O �6`�8h��̑;/�M���,D���E����<�H���>P��!:�f5D�x[h/f�r�r�k�{�f��v)2D�<�OPl��e�}AD����=D���@^+p!���s�"{I�\�w!D�h�!
W���v��6g�� �J?D� �˝2��A�"����1�r�<D���E��u
 �9p�z �K;D��
�)�/BFy�&���rX3g;D��0W
Җ9��%��J"-5Lp��=D�H�f�ڛ7c��GN�#k�h�j�.D���a�X�($�m
a��0sE��&D������!c�lP�`d�%�%ZѢ�OܓO��S�g�L�sy,u��j������HQ��ȓx�8A�+°+�����@����ȓ+��#cÞk���E�މ'�P��ȓB������O�D�X��Yoل�>.�I�e"�a��IyS%��6��Q��\:�sС����Á� %|�I��Ot��s��֌7<�j�"G� 7�u�ȓ'0(�V�R==�I��̓��l�ȓ=6���T�%(���p�mj �ȓq���͜�b����1��y�ȓF�\��c��ic� � �O�U�����Z
B�[�N���ܡvb4P�~<�ȓl"L=��P<c�E	�\�pAl��wHXȹ��&���W�G5_9A�?9���0<�$e�$F�!W�]�N�<��[�*����v��R�@J�ɎM�<y���Q=%XM� [H�kD��E�<Y��S:/�8§�`���LTD�<)�
�°�8DՍ.�hy�u�<A��K�3��s�rNh��Є�o�<��̅�2Eƌ���+/�����A�<�"J�F@p+�lG0]9Z�b�#�@�<�R.Ei�����O& @�碒h�<Y"]B04��%�'�p����b�<i��_���ÓF	�3��8B�$�\�<�%Ы)d��S`�D���|�`�[�<�"F�0H��U��T{�4  c[R�<�ЁE�~1ܵ�.�!S�E��O�<)7'�8[KUk�K�UO�=��h�U�<� jE�'�@�(�J�O���+T"O.$���"xLY��o�1x�̛"Ot��)8$h�07�bWT��C"O*DJί���\;%B"�p"O�Iacʰ#B�d���
>92��S"O����H�*Nnz�����LlP"O*��!��&�E"�N�u�pcp"O=��ǒo�����Z�ah��۱"O��� ���/-���\9n����"O�m8�%R+1C*���b�=U�t��"Otൂ��J�z��#���x����S"O � ��+@c��YEC�)1B�$"O���L���X���"#~��5�v"OI�#"�f)�����e"OfEj�!�VnQ�3H�M�<���"O�=c���%�rE�V��'���)�"O^ȣ�ɏ�9R:�+bn��� S"O�m���2��`�D��B��D9�"O�R��T�U!V�:���19����"O`cWN_(6@���eŝ�S �5u"O�}��	��),�7f�X���R�"O�˶��A�qbUd	=�͐"O�pB�a=YN���"	�9�����"O�p��"M\&�U��,"�Xx��"O�1!Q΄�%ny��b�z���"O�X��d��	VR	R��
�v���Y�"OLP#�X$/� �15�U8=i�P"O�蚷e s�u��&V	'|uiD"O���g�IƌHؒƁ- �4�c"O��m�qu65RP�:���"Od�%��D-P&e¹x�!"O,�C�ѻ{���r�dO�Gb�`"O�Q[ׂ�!��4Q'Ç�T!"O4�)�.�w����4E:X�S�"O�����r=ĤK��#���"Otx2��:�n�r��['g��@K�"Ox�%�O�o�Z�G)܈3��{�"O��Bs@A�:�.�۰�B9a��D�v"O�����!d�x� p�1'���`D"Ot��� 49<@S2P�`����"O0,"����T�Bk��	`z��R"OB�れӝn.�=ՆJPI�l�a"O�CC�=9���̘ "��w"O���h�U�H�i��ĉyh<�("Or�#
� w������:w��ʁ"O�	8b��!H�(c�����bW"O�U�ߙ>����U�R� �@�"O(�`�n��VN%�#�(�@	�1"O@9�"�94��/ߪT�D"O��u���rp�$H�7�(���"O� �Ed�����邩W8��U�4"Oҡ���E@4J8
����A�މP�"O
��ԫZ�b�������s���y�3[��@�/��9S��Z�4C�I�~�5H%n���Uq&���:B��2Kb���׭�,^�=^bЁQ�"Op����9���hs�� jϔU��"O4p�ve\��4��d�A>��!)�"O�z'O�
Q� �0�哋e�ƴ)�"Of��A�cNN�1���S����'"O�e�'�� ���s�ۨ�~��2"OV��/��,��D�M�lt�9�"O��{�䖌Jelāc,9fh�@Q�"O��"4�+������4Q�1�"O� T`� �T�QF�}e�L�`����"Or4��H�v�
�*�"?x��y�P"Oظ�ī��e�xs��Ѝl��P�U"O��g�҂�.��go��Q��C�"O��P���
�z�r�8R�y�b"OfmZ5�ŁJN�j�Ob<E�4"O�q�@��J�N@G��E@!"O�i� EXN~%��c��g֘��"O�=A�m��<��❖9���Q�"O�(�,�.\
�7A�/���a"O(�p������8��X T����"Ot ;a�	Z/F�HōZ7!��U��"O�Ȣ�-�9$��""�](.����U"O�Ѐ�hI._Ϭ�Al0�rQ"O��DD˖gi�왕�رa��b"OKE�����EIQ5BIԬ���y�"��#{Z��1�̊
�FT�����y҇���8g'�nl�4k�k]�y����|�T�ʚ��ś���yR�F?[g�غ��A�e����EL��ybDSl�\5�a��-X8�EI����y��9oX @b'��9��e����y��+^%��95�/��$�#o���y�$�E�ܼ)d�\�'�l0ٳgG��yb_�+� y�^�7�q��T��y⦎z�0��bޟ8ʘ��"�#�y�I�.9/ |����'}J�j�CF$�y�A�>=�ı�@K�)��Б����y�	�t��E:EdJ�
�HjE��4�y����<�;���<}�L��T�^�y�93q܅�Q�sv0�'���yC��Yp��C��q����Q,��yr _#[)FJV�O r�@y��.Z3�y�!�D^XT�V�9qK�3U*Q��y��לP�T�Z5�B3m.�ش	���y�jW�0(A�ĆD��b͠䈚��y�	a2l@Ӈ�*~)VDq�U��yҪ^��V¦��o,P��#�ۓ�ybD��){�T�gя<�p0��S��yb!B�|�r�X)64H0q���Py��/~<�A4�,��{%��O�<Ѷ�P9���-Ď�y&'TI�<��@�I����!�68,��eSo�<�g���*䉕g�6v�A�Yd�<�7$���8 )��74^�����[�<٠��3�L�@o4X�����QM�<�Qh	)pX��ӫ�z	>�{$e�r�<A]%K��KpC�ِ֘vGGm�<�0�U�=1��"�/f0�eΊl�<�B�މK���Ӕ�Q)T��DWl�e�<iC ]3��c�e�=}���C���`�<���$����j�H2��%HAv�<��'�:b}4� d+Ǎ��q�	p�<q�@Be(��R������A�<��n*5D��燋c�E��&@�<�gغQ2����R�>�n@�� �C�<�#šVm�yh&e
=�HI��OA�<���W�� A��e\viE�s�<���B>88�d{aP�e����m�<� ���ɥ͊g`�0%j�<�b���`��p���?a��3��Az�<A5��t+'O�`<��D�a�<�P�RD%*�:�C9n�|K�CZ�<�FC��!�FCA:5Vl�a�Y�<� y�hǠz\��CM��u ��"O�l2�֑N�޹R�B
5~)Ӥ"O6-��/H�f��M��S��q"O���K�)qzTI!����YB"O�l����`͌�q�M# �M�r"OhAf��	/�iX�e˨ �x��"O��H�lU�=Tz(Ȇ���|@��"O�т��£p<�u������D"ON�)�F�	(�aI�C??��ȣ�"O>���/Q�0�PF"���P���"O���(As���ǚjJ!w"Oj]���<n"^��#��+���"Ol���L��U��M��Q� ;"O8�3��ņtX����ڈ �$�i�"O-� ɥ(�`:���t�Z�B@"O&%p��J�QMb�0�@�3r�iQ"O�L��
�;�x3�JGw���"Ol��f�(H쥀�À.E N-��"OJ�`Э�"Z��ڡ��S�$t��"O��b��Pu�8��0�Q���@!"O��9���:IK:���՞um��C"O�Q
S�ڂ0,�9�m� ��""O����A�JQ�$���j4���"OV���λ�i�#C�9�f�b�"O4m�┯���F�R"%��]2�"O�Y��h�8����*셂u"O�A�p%ӡl0޽AD���I}6��"ODa�!�*C:� ��#"ql���"O:2uN�c�lArDς�h\����"OP�1"Y�un֥X�D�(b�L��"O���4�׵'���S���5]�L�A*O�`��͗f X�A�$L#� {�'>9%�K��i�5AD�����'�D����˞��qc�͜�}��В�'�H;D�N%'yJ�ʕCT�'h5�'*R����:_�Q�	�S<H�'�
�3&!FL:��O)Oo���'i�X� �B�d����Jy`���'�f{��'"3�	3�L�޹b�'�x5$E+d�1B��=~		��'�@E���1�8L�T�s�(P�'��P�SJ��X���E_�b�\�
�'4�T��ΎH���jN�S#�|	�'նE���������>I�=C�'���b")ƴ&�Z�Ђ,͌7"�`�
�'3��1�lΠ�
ݸ��-y�!�	�'�h�P�Ý={��D0�FӶ|=�@:�'���)�n"}�pE��`Fzm����'��I�,ߘ4���Ba�k�r�+�'v�� ��:�pA�WJG�^�r;�'��A�� V�4����U'@�J����?�'g6N���E�2��|��M��&��}�ȓx��( 5׬oM��#�K�Y��y��t�7e�D�|���@�w�� �ȓGE~ȃ#�[�l�����'|C*�ȓ*a@a W��pˇ̿u�ի/.�O��'�r� e:�(�9�/F&o����'��E	�ሢl耒�S�`�l8��'2��("�B�(�q��L2�dZ�'�>t�
�;.��C�M�A��!	�'o������T	�2��87Vт
���'`�mZU@G<$<�%�5* ��	�'=���t�Ŧ,D +2K����y��ɬ�ē@;�p�k�a$�D�����S�? ҍ�C�3��y�rd��9�fp�t�	"�HO��Rz��b�(J�xcO�@�lB��2_.��B]�B�fp�sL�Q���8�S�O�rh��n��9�HL��+D;U(�z��'��	 �R�!�ǫjTU��*S,:5��D+�,Ȣ�	l�� �(��b}B!�+<O�"<1S�W�z�0�(�cZ��%�G��G�<y��R�� � ��98�KF WF�IU���O��m�e�����ࡇ�s"쐪�'��(PQ��A'��)A$�H���}2
:LOֈ�L�)]B��F�M�v�]�&"ODHӲ[�Y�����'%�< `"Oz�;RJ�a)EY뜐���'#�dY��[ "T�}H ��+mp�!�פ9D�Gbήt�0���o�-2��� �6D�pR�	�34�sC�	7,���,4D����jE)Pg�t���TX�����2D���RJ��A�8УR �?8H9Gf<D�`[�f��8���z��N�"�J�a�4D�4�S @t�`�a�/λn�=���&D�t0R`�&�����B4�Ru7�!D��9JSr��Ը���e����4D���E`�2H��q$	ͯ8�����,D���DDK&V��H)��J3/��(�/D�4y�뉝�֑�#��r�rx:�%-D�ĻW��Q-4��ƁUs�p�` -D�HQe����k��
�s\��+,D��j��ӌv �L+CO�G(|�-D�,;0Ċ+�z�
&��is>�*D���¶(�F�04I�N�6����#D��ь޲3u�9۳��KZ�@�5�%D�P�,@�b<R��֋ĜI��S�'%D�XA��;+	����Æ$�Z�дh�5��'��z�Ǯ	���� ���9�^�;ና�y�L��o�dY��+��Ё��:���9�O�ccGC+8�&`ϐy:��S��Ic��O�O�\x�!�ICXP<S����L� p�'�.x���
Y�@mK���nI2�s�y��'��O1�"C�䛬��xP$��L�JuP�"O�Xr�����q���re6l&�S��yr%.Y�p�խ޲*�:�&�.��<	�O��'��Qj��ܚ � ���`W�x}��	�'MDj��\�N�9�/�kd���J>1������b,c�Ğ$]X��cR!�=�.@$"OR5ca;<J���W�h'�Ȩ��	w~��d���np�`#Jf�NL��K��!���:6�^U��%��DfJ�
^�̆ē	�f����;D��#6��82����I4��>�tgBҊ(ŋL�0�ʝ[��+�!�*L/�-˓DV5�������5ўl��	�SȚXqeb٦ R%��!��p>�B�I},�l����-��<�5��S/�IT��MʟHO���z���<	��<H�C#d!�T7Wv�)��&]�<����4fP�I{���SC�;v%�AL�@Qa)lOT7MH���䔣x"ᑲL�bQ���5i�#S.!�$��<L`�r"�W$ ��(�s��+�'^�'��Ļ_�u���G�$���u%�Ii�a����<���]�t8�I��[��
m��K�<�'
8�j��5`D<K/`i���p�<1��\�(�\91�G4�r�c��A�<9����(HrU�;oXH���y�!��h}�A�4��V9�;��Î.�!��A>o�ta:t#Tf��Y!E��?-qOrb��G�� ,<��Z�M���A�O�{CJ<`�"O�����J̸��=v:���C"ON���K�0Z\�1bO�i>�,"�"Oh��0�Q�D` [����c0P��"Ox�A�m	/L�0�s@�� H���"O�-��,J��*�9�f@�[%"O~U�SO�L0{"&�7��&"O�RecˤRgISׄF�I"�Yc"O���0G!�tl�`��/Y粹ط"OlA8�,�7��,Cb�a�*-;�"O���񥝤0�^�)G�_T��X�"O�<�m--j�3��l<>m��"O�arf�ĄR<\A��A�,�xAu"O��!���2�e���H��"Oz�Aa�?i#Ҡ��	%��"O�Dp���,/,j8
�G�5��j�x��'F�z��ɳb�^
'*�-'�ճ�����>��OV��"RU&���c@*4��[���Ħ%��I}srɨ�ƍ�*��a��˸]�HC�	.$�E�� �M#�X� ]�y�t��4�<�d�+G�2���lF$B7�UA� D���fL�%n�2�JD"i���"�J D����nU�n����Ai�ؠRp�(���+��y�$P��scʆz��z�4�y2��p��#�����!�@��y���*��1�ɔ5b��l�����<ib*4�ɲ6ӸT:� k�|$k�'�(�����'>�y"`�2
���DDZT	��I�Tw���a�"��ӆ`8�)D�[��ӋR�����
��mP���H(�ə�yB�0#��6zZ8p���
wiRX
��1B����q.�e�g��fn���M�($1!��I� �VD�F�)��J�|ay®F��T"��s5n�fX㧐�=��P�']ў�|"�h[�8-�H� *��O㦄"fcy}F�J�'���i�	, C�tR�bN�<2�x+�SO���O����8�*Ѱ�AՍ�M��9fщ'K���\�~*��u�b�1�Q�NI&|o<�"O�?��x��>�rD6j�B݌���M�,�Q�F�dM����a�-�i����gZ��y��Ӟ\��P䄛��ZD��6�y⫌"QI~Tc�Ɯ��V�{����ē�hO�I/}2B_8R���!$����xQ��y"���,ږ���r 0�N�#��'�r�I|�Ş$�laU�� ���2�TL�ȓ_?h��Ĺj��;�c ����'����O.��D���x8uj�1%8��wD0_�!��CX�A�W)+*�I9aM��rC�	
0Hr��v�q�TH[��I-rC�	�1��}wK�f^0��`�ط��B��#{i�u-��jpA�$fڂB䉞.0���ò3 ������P�ZB�Ɉ-[���n��I'��S�G�#a��C�I%2��lX��Q W`�%�5鈕w�B���)�gA�U�T����& &B�I�Dv�I���81!�����vLC��&:�n<H��ęb���+��.�lB��.� �mY$΀��r�R9Q��B�ɪ* �a@�V���#`�ΔԖC�ɋ� S%�f�8DK���;.�B�.lK�5���ڙ!&r��"��B�ɹ{=P4�9�Ι�7��KJ�C�	�"�&]35.�&�=����<<�jB�	Yt����K�C|ID�T�A�^B�)� \�@���@���#�	"����!"Oh9����/�����&΄#g�у�"O��QB��(Rr��4�8q��Y�s"O�%!���w$�� �X�/E��G"O� �Ĥ՜dh��vL��z/*��e"O�@����<F�A�ceޗ^��Qc"O�� �Q$^�,)�m%Yʶa�A"O��S&͌O���	�L�o�&�'"O��b�KE%=���:�j҂G���q�"O~�`�_�)C43)� xT�1�"OD�IF�W�UB�qh�7ns�0�"O9҉��J8�dȥd{,$إ"O(%�!l�/ LD$�í��Nu�E"O}c�c�U������ʋ�a�T"O6 smա1� "ՠ��fd(�A"O0��f��
҅���"�r���"O�\��e@�[�&��U�\�O�D�@"OԄ��#�)tT{�Jg�d�G"O$��,����S���78��U���'�y�ԉ֋b\���>`/V$��.yJ�2�'Z�4�'([��a�� U��dZ
�')lM����P���Q!�W�%7�l+
�'��0O3"�MSP͋�.�M�	�'��"a_6\���Xp%΍ia����'v��p��Y�0ޮ���*�&j��$��'��EoH�;���1n� U}�D��'��h��=I���&VY�u�
�'I\HA��F�3�8x�a'J�W��[�'��0��°+J4��R"� J�P���'9�i��h�$oa�x���pUP���'����Ad.b��q9&�N�r�\��'6ܝ��D�y�J�
��d��,�
�'� �"���\1X�' �t	<#
�'[���#��N]x��VZHxщ�'g�}�왒��M���ʊC�����'�@�a�Ymf81���0z�D�'Vݱ���u4΄��2�9Z�'*�0�A�])3E�V&*��2
�'7��+Vn ~�)z�ʅI^�D�	�'������.'HN}b��8�u�	�'��Uyg�\9�3i��)�`���'�r��*"Î�p2l�7�����'Ej�rw�H�p񄉋H
Va�pY�'�V��R��Τ�S�^�V�H`
�'hx��Ύ>T�� ���[l �(
�'	"d��f6�Xm����B
�'~��`�`A�]��`1n�[D�		�'����G�̈J�
ЂL!�*���'~b�����t5NP���	�*-��'����������Yd�&I]y�'�y��ʮXiV���f��6���'v�,� a� 9-bĉӤ[%�����'��l��P+v�mqso�-hϴt�'�65�fh����ч��e9�1�'X��2��.&�����#D/�D
���+I*N-���!�U�##D�0��N�o!p9B��'qʘQ�"'D��ل�W�6@��)˵L��t��3D��IP�<a�ry�g��YYH�R�-D�8R��@�TS��؆�ըW�L!��=D�X�O+ЈC�l��"쀤2��?D�TGBYRu�,3D���ܠC��=D���N9I����Ԍ�/;gĄ�=D�|!�L�[�±
Mr?�bu�$D�� ���e�K�nU��;0�Pu|���"O�ݪrn��G�~]������G"O���tؽ&���x� �ll��"ObL`WBŨo.�mvl�
/r�'"O)k�e����$M	nzⓟ��OȚ'1qO>��ĶCs��(fC+2.�Ɂ�'T� �an@+�-�b����� |rƞ=��0��'X�����S:ib��;H������x�pC3������E@,�Q1��A"4�N���o-�O��a�O�[pܬ�E ɐK�䢁��+|���Cf�. J�O��wHWn��!G��D��'�I��ƒ�L���[�SZ$�#�O p��9����J�"}z5LΉt��L80�߷rV`8P��m�<yCBĥs�ZT�%&��j+���dEL���� ]�B���K��g����[.#S2���`��K����ɂV �����Kr��+��וH����Β�n?$�Qv��3_V ��$�X\I��5fvu
�V�V����B�J-¸i�든l���J��i�!R6��XX^ay���#]XM�p�4D��;w�D���<9���,S�� �E�>��DI0Mxh��UgP- �ȍ�S�RJH>��R��,Yz���f
�}ب�9(2D�,����b���a��5����ޣ+� 4�j��W�V\x3A�=b�쓟RX$�xb1cU�<xe��4i�h��I<�|r#��J&D�J�Z�>����)ޡ�$",����E.C<�:��	)$�d�;����:�y�_����(.<O
��N�{�&ԹȎ�&�b��$��*�0i��M'Ģ	��#����xC�(2|V�Sc��((-r��9��+ 9B���;O: �b���87U�c?��JD�:�޴+'�_q�h�z��=D��!���WJ�p0��I2pA6�[�K��^L d�P�($�<G�Jc?�ODܻV�T ��"��#�`��O����-  �X�m��;�a[N���� ��hs0�6B�}:��4Oz�JT�1Q6@a7cO�M�Pqb��'b�|��nG1�L���܍Y��ȅm�%�dq⨀v������]ڢ!Y
��G��e��� ��ؕ��A��&�|[�ߪ,�G(@��IXGဌ"�����5�4d٨)�2$;��h�GĪ�yr+�Z�����v&�x&�����ȕI�r����R�e������19c��	�c����*���
U�v��C�	76�*]����2L�~y���H���R5l�� �tj�r�ػt Q�~� Eӎ���2,4��Ї��28<4I$EayR�ϭajP0���N��c�eFĂ3C��z��G!�6����c6F� cD9�O*)[ ǒ�@pzx8$ǚ0#����$�|���!���A�� x"�!t�D~�r�?�����p�Th �P��8���!D�����c�<�(���"`�zd+�?l�pX�,�@d��JҠG�E�,�?�x�H�<��$X
T"X�V�Z5JW4-)�J�b�<ْɯ5.�*���X�n�HS�!)l���7�ï7k����o�09Ң��n�'P��UkV�1d>pX`@�Q�<H
ӓ2> ��)\��B��VA*�b�t��ѓ�	�$�&PYeDB)5�tH���5&J���S�P��E�⯆*?ڔ�D�w#UoO�%qR�_r��<�篊���ӹD�l�:��Û>���K�ŖF;�C�ɯC>�M�ů�(Qf��P�C��"�*�c�X�~�e��t: �!"�g?I��?i�)�N֘@�ҟLPhB�ɪW�����T�cg�p����+Mh�I(>��3��'��H�Ӄ�*FL@"�D� Nh�� Ll�p�kӂ�3���y��H�\�@�62�!�'Њ��҉؊/@�J��ܑ�@��jA�yE�T���J8�� z`��L��y�c�v�|���;�Pp�f�܂:� H�,G�iK6�;H�"~��������jļt!��XUU\.B�ɮ6��قDd�j�<��vj�y�F��$ ��|�E�ԷQ�azr��<�0R��3~�N0c� �p>)�l� l�u�T�Ǧk��{'�1l�[U�B�m�d��'��0Zr��3ZZT������2��)���Kq��:�fԲX^P��}�Cg��S��l�����l����DH�<i���xFqɓ�zLA�r*��&f,ڷ��9�����Tt?E��u�:-(&�^�Vի���1 ?n���S�? D��r�e���A.��M$����O����w Dr�D��0<�N�i�Rq N�P%�xH4	�X8������Cd���3�=ue�2�`Q�q���j2jL�Tdx�{wO�u����"�l��a�I�5ᐨ($�	! ���BS��V�n� ��dG�%QϦ�s��{�ࡳ�Э�y2�7<	�-� &�hܦ�uf7�?ɳ@�3	jz��f�����sӔQ�@j2 ����
͑-�)c
�'�F�s��\HՌ�CF��+���H����3R81Y�'��|qg�Y�*�P �냍��p;��$�x˃%2�ک���b4JeK!΄3$��	c�=��(SJ���b�L�Q��7�&�R@����ϖ��O�4kt�D�Q�@������!��'�%��h�S���g)�/sվM�,ONQ����ΓOQ>���L4=|���V�Y���qBA-D�|3�Ð�=�r�@�H�J�WJ�w�II�@� 
6�3扏���p O�c�LiA	�}�@��$
�VR�qޱؤG@�eW���"|��1�=�O��2��8�\�xP��/�<{7Q�(c1��)�8�'Q¥��Ċ�4�&>�
p�� d��#�V�M͘<@5D����[5y�m�F�҃q�t�[��_}R͋�'���c��OE(-0g�9��d��(qx��V�r��{��
�2y�~R��j����a
�e����Ѷ`6ީ�˟�L=@A�O��QΜ�^�����P _���4
�c�f�d�dTQ���j�I��Up���Q?�R��S��I��?h�¥/[�ǐ�n�g�*��$�/7/R�ҴF��� ��E�L/7�d�'6�T=��iήa~�I�V�$�A�j�%J}�O�ƴp4��Y<x��N��0i
�'� tX�`Ѩ8΀����j�ll��J���i fzu
q��#ZL��L�;����I�>!��>b�t���oJ(]�y�Gi�L��X�B��XR鏓3��V	�eCx	�n��� Y��T�(��؆v�pD҃	|d��ގ ָ�&ŋ��O�P���Э*��8"ͻ<i"A��L���Â�I'lLS@l�8(`Ѐ�4�x�@݀ou�����Svu����x��/^)�����[Uy���ή`�Nj�J\l:5: (\�!�d4eQP !��1q�����bS�(�d�'�d���ͅ'xUl��O����.&v������ϱU����'�����ΛH#��f��KzX@T�N�!����$OJ��c�+:��iG� 2Hpy3�"O�� �T�<�T�P��X13@�@��"O:�G��F��B�tޘ�6"O䐊V΂��L�Q�#�7�����"O*�4�P�>���iҢį`r��PP��K�����OJTڧ)ƣ*�
uS�ֿ\�¹�A"O���e^;"-�I"��3�TE�F8O��"߅#p.���F�<�a;��m��r_�y��6^l�k ��<4h7-�����c��Ui�t�Š"~!�)[�]����?��<��`�]�O��W�(9���	��7S�jG�?E؝ڵ�ʧ|_!��<�^	�q��I�Lܡ��P;��m�si��@B��O��}�Pa����)�,#እ��cƯm�x�ȓE����@�uS.BMJE   �I��JP)��� "�a{��ɬX՚�W#ʤo�2�c$ق��=����7J����i�Z�*$�ڎe��4⁤mw�A�"O<�V�3\��BP�Ia���d��#�"(6m�"�H��h9`,ݢ1�Hj"/J�E
ր1�"O��; @��]�%R�O��F���Iq��� z��u�b��"�g?іŌ>2\pC� T2�;tK�F�<�FK�i"��9��P(�&'��<��!i���ߓҴ  !`�+��AV�L�]��	y81f1O�,X�"�80�|��8 ���"O�P�S��v��H��3o^(! "O��ˊ�+��+s%A4!F�"Ot ��$d�$4����~%P�X�"O��cTs�ё�d�v�
U�&"O4+�h�}�r��$�o �IQ"O� <�
V��R�:�
�@��"Ox����ЬD����� (q��R0"O�����)f����a�ǜG^\�w"O,��aB�E�j@#�l��7"O@y�Gț_H��X�cp&�"'"O�e�VEB�z;B=���M�8q"O�a���S�rz�aU��h����V"O(����H�<V�T c�<U��2�"O�ᆉ"Q�]��?~�k�"O �kD���]m�|�ק�w��v"O�0{P��UT��
0�[ (q���@"Oj��f) $��}�����?J,!��"O舻���[�&�@@�\�H	{G"O���B��I�ŀQ,e�^5c�"OR,���8~Ԍi�Lôk�@PA0"O��S���sh �1e�u�L���"O��U��V�
t��k�
d�:��"O��J���
������U.���""O�t���+E���g
I���"Ot��F�{8~����Y�����"O��Ȇ��R�m{%�W�d��ݺ@"O��BW�P	2��$@oJP��m@�"O:��hڨ|����@�%?�L�s"OR#�iI"t
zI9pσ���c"Ox]�0�V�q3>Ay��@�40"�"O@t�f* �O9}����B�t,x�*O8�SS���u�4�;�nL'Ds���'�Xxy�D3â��0�[�< ��'�j���V
>2X����FQRX�'���T�guԙr�Iʊ
P,lR�'�d �ƛ��t)�,�';�L��'�py�/[,�蕫e�[0{5pa
�'an���^��*e+e �-��p�	�'����BŇh�>�J��˖K7���	�'n��5�L*�j��j'D��U�	�'hTp 䆔�N�k�ȕ*��	�	�'^8�z�*��G�J4S�MWt�Pc	�'��@�A�9j�(�cC^�{�Fl �'�ZyX۹z�"I�'�z���2�'�,�G��D6�H���],,�6���'�|)C��?&��(�`ѣ
��H
�'5v��ǝ6K9D|�3ץv0 c�'�8 �Wl,VrY)3Nձ%�ڭs�'����E��~��Qp������'�(�R�A �|�`q�G�E�2`��'��h2�H�L�:i� �Ǫ�҄Q�'䤋R��Sl�H���K�J58!�''tebPcM
VN���Vj��
�'$$�ql&N)�a	�P����'$�h���9xܨ���N|p@{�'NE�.�4���0��=LD|C�'�@�r�Ȝ�I&2D��O٣=��L�'�x��d�ĝ?��1�T�^�4�iZ
�'-���Ed��S�n��'Ŋ#p��	�',���B��-7��%k��]0�'���@HŮ.�1���7\���'�\��­4�M[S�U�D(�5A�'z��#B���T�2�� �4Q
�'���#7��n���.�"{�����'�|�x�e�@�R�g�k ,��'���t���@�� �.`�`�j�'\�Y��]�x]�@��d>*���'���!��l�Dc2Ŗ�h0�y�'}L�!�#�%\�8�P�@�c n����� >�q 
�dF���H
k�j��w"O��h`��,�n,SS�2e�\� p"On�@V/hj��l�sR��0"O4�J�*+y��8�ˌ�/~V��a"Of=3s^�G0��u��-R���6"OR������(!Qɛ)XjT%�"Oڤڠ�ܺ�j�"дueZq��"Oظ�g�4Ih���R!:o��� "O4��S�Q�N�5�e���~�~9����({���3.�qO>u��I�7)��y���:_�4Q�Ռ7D���4�ԫ����e�2<9ux&� ���2><aX� O<9��I�T�fkT7b	Y���'QZmBv�޼{���r�gG�~� ��f��M�Rы�n����+� Y���n�;�0�)f>�_�%��^
v�ؓ� ���L>kNN���ɀ�>ᒭ��"O ��h�B��M��畱"�\1!uV�bU/�&;��		ǚ>E�dD޷Ju8��Z�h0�6a��y�L%m�E�F��P����%b�R��A�,1q�E�"����'��'N�%���C��^ K����إkX�[羡���,ʰ�A���C�M�%�;�ON�*D/ǅR�e�B� `枳����w	!޺4C5�����B�Fa�t�����۲���y����d���!d�K
v�������D��A[�L��ߗ��)ҧ6{�����L.�ʣh��h�F��ȓb��`֪�&\�:L2t��4�)%�H"4U6�
-��	�A�DU���[�"��ǆ�5��B�I�@�@q���%"��!1� ��}A,��h^����1W��5y��M'J�l!I��<!�$�1{L����av��L���~�!��)Br��m4��䠑 Ё#!�D��~��l� af�!&�]% !� �Vt	V)��<i��BFT�\�!�d f�Щ ���$@�Xr��I�!�D�fV��3��F�d��py��Hd�!���3($�X��牕U%v���d��N��|�oޒ$<>%�I�y@�9�HN�<�6eh�cīYy��'��Z�a�ᆒu܌��邨4�t@���O�5���'�bM��Sl�L?0)���S��J�*ЉrT�:D�䣦���i3��+@��)Z��ھh܀�����S]f�:D�#G���}��'A������\�q�/XY�Ұb�'IJ��ę��|�31���rɠdT>D��p�V='�iPm�����}��I!�V� �@`�M��{���
�X�d����� K�<q�H 3�aN�-�����J$���;��'�B�x`�!$*8l�FF�3b�����b�Wq?D�؁`\�@O@@�D�M+e���*c�)ˠAlX8r��4>�FB��/Y��3'��G���ȕ;;�4�A8uX��*!��)+�D���L#�'�y" V�UV@��A��.Q����!�yR只{�~\��%�`dY�#(�]�G-�']Q�hpA��;�v�	����Ov �
;bZ�4�����`�,//�{��[��¢"G" �6D�%��J�l���o��\�`����X�fT���'̔�Y�-Z�Y8E '�Kqf����̾g�=C��[40�,d��H����<��u�%�[�1BB5��\rB�I�6\TPas��Y$	v�M�T!a��7�H�d`%�<C�S��?���Wu��U8d��8�����jJd�<i �)G�R���:��p�i�Z�<qI�]ͺ�#��j;��ðm~x��Ӑ-�>6���Ǥ~�n�ȅO��{8�����ybn\�.��뤀_r��Q�5�ɛ�HO�\g�C�|27dK9N@�1D�ׯW��LT+Dn�<�����>j�h�4D�eºH��/��z�
���fJMF�٤O?���e��:@��,9���	P셷<!��_�v6����S V�a2v ^&<������R̓��0=���?�z���ύ5� �aEC8�����ݚ�/�>�ti�4�J"u0lT��/�&����S�? x����S<t�n�c�"�3J��QsU創U2l�����v�f�k�����Ό�W&��}�<���̚��y��/*�{�o�m����4@xj
��R'ӹ1�u�f�	�~���'� h[�i�1Z�(��%�Z�EdK�'��(Y�
Y���!�⇚1o�i�'�b��V��5��9s��{�8V#��]l�ց�[�J}��'�On���*��hd(Ƹj���
��8�&Mҕ"���l���'{ȝ��*_#nH8PX�$ܚ$X"���$�?���2UO4!"$�|�D�(�����d�Hy�o��<a�� .�وRk�v^�uA�#W��0��^�-��;���Wy��	 �f��@K
��E�%��@��"�C��>�2�͝�n�NL"�*�'$ʀ�'�6���ԸKN�	���4Go@�
��~�V�p��k����_�.��9խ��Am����L h�'9%ۀ��'����RhC3]� ����i��Y���ߗ@��: %8�V�� �b� u2b�[�o.RB�	6`P"̪� S�Utr�(�.%ʓL�R����H��S�Ow�� �n�p��԰����t�'ۂ�:n�+6Փċآ)��Qs��|���#+��Ac���y��R��y#�hF�E�� �W��;��?)##�	Q��P `�:RH�(�i-a�4�P�̌� ���D�1���j3K��y $
�^i�,4vd���A�hyrɝ�2�����Gⓞ;�2� O u2!��_���B�ɴ/��#MMT�̌��.�
8xlI�'h��R�fE5p�T��C���̉l�Ƚ��O�I��ծUFi8���U�~���'w�27�A����K���+&���M�����H��e�d͡'g (dd��OZ�������.%K!�ޯ?��b�I�j�!�0�Ӱ�����pm;p�]��Q�	�Q�ZQ��b�č�a>�OڴJaM3=�5h��/Ae�=Ғ�O��A-@ :�`!î��Lxs��j
����$��w�<�i��a������(�y�A�(_�X�sL��MYXH���طkj�I�b�jl�rbC/
ȪA��P��4D\��-<zt��K�;:~}���G��<��I+?Ƞ������Ŭ)+ZeS�FىF)rt��*�
]���'�J$b�S=W џ���蘂<|tY�a�ߣkqBY��1�{��	�c��-�.O�-*�ᐛf�.�3��%����&�/7
�a�'����2�"���a�^46�`p�',m��κ]����[��}��Si����8�e�[�<�F�����FE��8���e�����u��	�k
C�3�I� �ؤy���6��3G������Ȗ!����Z��<X��L�����T �zC��:[9���!>�Z���\�&�C�I\��L{��.O�\ ��*W<4�C�	pKZ�"���vtd�w��rB�I�o�6����@P\X�CI
V�B䉊Qc6��wb�=B���)���&�%��"~�	�'��0���p�@��ּ4��C�+�nQׅ�5@��pA�`��x�Z�	tYI+TiOW��,z�*�0 �p�BR)�2	~�Z��6|O�!��W)F�`%r�4G���a!�5Sбs�a@}�d�ȓD�9P��3!�����V�.|�?��-�ʥ	3�.ҧ-�)�Hۃ|�Xh��R�(T@��ȓ@�^L�i�	&�$p���`fd�"Ĭ���@�>Y���O��I�/+_�\!J��C6,���p�"O����'˦t�]�Tg�a���'��q!r�K�.���퉴z���'E�"@��Ɋ!@|���Đ��(bd�ε�M$�����U(�&�t@�� SZ�<q�V�)3��ǡU�QY�i�V�_:m�BB	�Wb"}Jp�H;}�^pA�g�2mp���5O�X�<A���F��3C +�;�'%<�"��92铘h���Ӳ �j8����Ԁ�2 K�H�!�Y
��X�q�����}qT'}���RlZ K=|O��A�0`�aٲHKb`���'�&%��)��<i� V }�a��E�$.$	�	�U�<�f���~j$� �3��]�tn�}�<� ��i���;s���Ơ�`"O� �F�Y4�����-ެ3�"O@��5����1|>��b"O��r(Y�j���A� `C�8��%>D���v��NUذi2�)8
Y�El>D��y!�E�$����ƛI|ڕscB3D�`"D �d4|4+�f�"�FEiq�3D��qS�T48�T�c*#2\�y�H4D����(P_��� ֪Kj	0�5D�L���<5T���3Ʌ�Ah��gN,D�pS��P�'5�$f/"O����g!D�t��q[��� T���a�.>D���a7`Yq�+�|�i��f(D�h�� f�XH�e�+��2f!���g�iCB��[���W� qi!�dۅW��eӧ�!.vmBR%�PT!�Oy���F�-�X��
Z�
"!�*)<0�pEnY:e�>�jV�S�!�$��#�<!#S؂B��ti�Y?6�!�	"�0@�� u���e(�*D�!�$�)\�<����6lg�l蔈G?m�!��H�����w�C�:���(Wg��@!�ŃD9�c1����X�b)ȫ3N!�dP���'���|A0���%O!�P�E����T���H�.ə`�Y,^!��� B�mJ.*RJ��dl�Q!�D���I��9(���)PeW_a~BKH��:P�7�N�)s2���k� =�ջ�#T��ybC�Tat�!�P?��dpHQ%�yb@
]��5�d՗J!,����˭�yb.�(c�fY*Ut<���f���y�&�	���ƈ�t��������y�@ZVH����p�R��M���y����x�N\<m��ܘ�dY<�yb��QF☺$JK�`Buu@��hOR�E�d E�]�q�%��Z�*��4<R�#����bEX�iya�&�&}�@Xse�P0ҧ��-`��
5�d�oG�wZ�@E��b�%��=�6d�1Q��iǨ\?/*d�S�
��lB$� �v����
�'`��t�a�J�P�*e�!���I��h	��7� 5���=����V>�ᧇ���]ȱ,�$,��C�K�~{*�9���0M��.�0`����CŎ���*e�I��ƕ3�>@(A�H��"5�B�$lbX1�Ow�l��B�N&Ty��(="�M�gG��>o"�t@al��3♄�u/O�8Z7K�	MǦ�@��(��(T�ONl2&èoRAѶȥ<�~���:Y�yU�$� !+H�f�4��W$"Lj�LЁ�?a��	�)�m:��H[aFY�<YC�(��`%Yr$�4'b��E�ӵt���*�<E�d�*T��� ��d9�'I�<@��R%��n	���!9O�}��'o���2&�Н:b,D@�.�?V� ���M�c�
١�'����$0�L$�8��`��mǐ0������A���In:��qEd��0|��J�I�z�	󤆳e�Y��_��~«'4�)�p�Ҹ<������(6��2�n�;���E+Yֈ�j3ρ��<���Y1\�p�)��S�T�OA;$#	/#��|д�ю�@Ŋ�0C3�ʓF:
&�����k؉<\���&Y� �`���Ziy��ڠd�|r��J>��hʸa�橃���A'fyC��"D�8���ڒJ
$ĩ#-��h 0�V�?D��#J1Wx���S
{�)�=D�D@4F�� ���e׎w4}�`,&D� 
w!�i-�,���B�򈙵�%D���Я� ��`22��<�sf$D�l�Q�]�4��yxCK3W����!.5D��ˠO9<my�c%Ϻ�*�g0D���t�@c̜Q"ʂ6�lx ��*D���DOτy]~U3v��>j�N<���(D���gb�*�|H�f-�=��ą9D�$�1�[�V�����l��La�:D�� ��[ƥ�C���s��tL�e�5"O���pÃ�w�&-����7��i�"O��x���%-��4q��S43f��#"O t����H�Q�A+�.�2�"O
M�4$��U5�9;�+B�p�x��"Oz}��+M'��L!��[�$h�`$"OL�M51?저�J�	OL2X�$"O��"f��@�\%ȉfJ���E"O�����6%�`�*cȞ0l>6ٱ�"O������ ��`����-\�pt��"O��"�B��r<�iC �/"��ȱ`"O�u ?�0К#/ſ�`�2#"O���E���5�@(����ad %��"O����H�% ���l[�i�z"O�U5�ʰ_��a�id�x�"Ou��dښ������R� G�zs"O.IRO�4<��s3f�@v9h'"O,��rc֟x;,�@w$�/W°q�5"O��bF�ä$2<R�G55�,���"On,E�\����
Bl���"O 4��Ľyv�QQ� �xh8�#�"O�H�F�ʩ�و�`E;5��|��"O��j A�DS��i���]��U��"O !�t�²-aL�I�DH�Q�|��"Ox�P�bN�^H�c[�mX�  "O��P5ixe����cd�h�"O�0�Q�O8d1T��fcS#_8Ц"O`���<d�th�#A@�DS8T1"O�tbG'��nNR(0��>	���2�"OL��Ņ�/��P���J�ڜh�"O�⃊�Ux�!r���#�hy��"OT�k��St`��	�Y�2�H�"Od8��ť#�V����ǢD���"O���逌|W�a�V��Ѳ�"Ot		�һ�$����l�S"O�E��g�7n�@�bUDM��(D��"O�*0J �Y&$�6⃈tO�HxW"O.��N�`Y�ScT����"O���@�.��	�+J�cԄ��"O��%Gבj��s��ޮiUX���"O.U��EΏ1�1B�A�-M�$kG"O���,fn�Q#A'3"=V��"O��UL\�cj@x���I9*�g"O4uѣH
:��YVΝQB��"Oص;�Eۼf��!jB�N�1Z�b"O�I蠏 �m���:�����q"Ob����M"jhQ(`�;l	zuȲ"O�}���F����(V�h�r�Х"O��ja.֫Fz��QF��3��d"OX�R�#O�y�Xa.M�Q:�91"O
$z��߯�<� ��:I�|��"O�� 1�\��rD�g��!T?�Q��"O ��GW9+��+U�F�S8�M*q"O�Q�p���3
 U�4�J=V��[�"OJ|��_/j��YF�N;v\y;2"O���āI�~�6-�B��)p���"O�P���ֻ:,XP4��#d�Й�"O�x�1�'8�����,1 �C"O����F�~�>��A��`���"OΨC�
O,�����{�p�"Ot��v#��)��i���6
���"O�,q��[?ʡC����X��, �"O((��mG>�
!I����tX"O�����2l�c�Zy`,@T"O� F9 b�G��3��� w2i��"O� f睴
� A��'Y�G{����"O��@�%��Z�� ��]�-s�ta�"OLM�.A�n�8( �PXm+�"Ov�0��"v? `����)$����"O~�)4DK�c�����ݐjmf-�r"Oґs��9R�Ր���v�0a"O�����<M^F�B����x1cU"O�x�A�0,>�`P��W'�j��G"O�(���Cp�p5�D��
{N�m"O��p	�$H89�kH P"mc�"OL4Аkח~{&���뚬S����"O�!R�)^���u���ݎa��"O���u�G�+ ��)��\Bg"OL��%AT�Xq�d	�)��3�"O��)�]J,{��̷A@Z|��"O��*�Ε
^$D���G�=^�4"O�T�%ϞL)(l���i�"O�R�� x*�4�k���0�f"O��Q%��Jv\���	D���X�"On���.��I�F�)p�M6B_6��p"O����Ѳ2�@[� �[��5e"ORy󆃉"7wXMAF�_�l�`��"O�������M[�.O "���&"O��x��9��b�L�G��Ek�"O�y���4:!BI3�J_�C�٨�"O��A�I Lx&|��]F�$ѕ"O�h��$�f'D%G!o8���"OZ�A��#Y��$���ЗlO�Q�"OF��`R)\��<�aeB�	ؔ�B�"Op�퓻[\���0�Ȫ�~j�"O����1ll�b�4�r��V"O0s�n�a� 9���&\�(%�T"O��[��S�c����p���;5"O���^�m{�)���Ď>�vD��"O�TSQ���?=�b����;v,hP"O�Ĉ���a���R+�.��!F"O�AZB�' ���Ɖ#an��"O<}:#P*{l���
R[N���"O��	D�I��1AbU�&��Ě"O��E�ĢJ�ԩe#�}�jIE"OR�� �3W8�$��#!R�"O:h4�-�~���&�A��"O�Y�e
��Q1�ׄDr���"O\q	�Q:�ś�AQ�Y��	"O�EC��s`*��
Q�8b"Ot58�Ɗ*����e VR4 �q4"OT���L˳zČu3�I���{�"O�ÃY$3yT�z"iLF�ȹ��"O\Tz�gU#�<,�CQ�Lx��j�"O�1���0%�F���k�r�F<Ҳ"O4*wA��bA(l(�A�5�A#�"Ol�H������d�	'�(4��"Ox���)�j�%����RI#�"O��B�K2:����EՌ ��+0"Od����-,�J���E8x�؈�"O�� ��N �3g�6���t"O0�	a�q�b�3�&�:��d�"Of5��ӳ�n�� �\\��|�%"OX�����2�VY��C�]۞xC�"O������6:49&M�����;S"O��K���6LW,��n���2v"Olh�ti�*�Fj&��`v��X�"O�!�ugǹaC�Aڱ�Â:I�)�"O�  �g�����F,�'B���g"O$X�����l �kWV�X��"Oh	jp@�wN�\U�.l�ʳ"O��� 5$N�Lؐ!_
CQ�0��"O�3��B�tIP^iv�0D@SY�<Q ���JA�Ο�
t
5GS�<����/(%�5k�b]�I�l\f�<�MD�'֪�� 6;��9F��b�<�Q��3���ҖΒ��j1�w�`�<��+ܞKע��2���Mh3��g�<���N`VTzR�8ᢕ��Fx�<�i�&T�>X��#�Q財�%��w�<��c��Qh(}��L_8!��pဢ�h�<��k4pF���e��6tE|A�o�b�<ٰ��	^���C���<91cLH�<I(E�?.Q3A�R�ETT��RN�|�<��G;Pr�苇�Y�W����u�<i��-0{���jB-m�6EZ6�n�<��K�4���6�M+N�,���R�<��g�UC0eG
�H'�)��P�<�EnU�\� ���T)l��aC�[P�<ɰhP�C�ܜ5���f�@�p@	X�<!��\E���U3J��@���P�<��*Վ9ZMQ��Z&�m`�Rq�<�'d<A\�
� _3Y�tYp�Ix�<y�`×\7�q�-J`�.9�Gt�<qq�8k��{�ד@+��*Ls�<�1È�j�Z�땋G � �d�Iu�<�j�/"�u��P��4Ѡ��g�<1ҩ5��`���>eL��H�_�<A�BZ�W�Z!�c�	�<�[r([�<Yq	B�2p��	���%�8�Ӈ��V�<���,*���vHY�|�<��e�z�<q���3.�L��DE�DcD�� |�<Y��\�t��L̝~�8�0��Wx�<� H҇m�XY�꜖bU\!ڤ`�p�<�0�93r�MCr�N>e�q���Un�<�Ì�U���2@ ��
b8�pU�g�<�ҡ���݋5gΟOP�!�2�y�Y�z���0�k�"Vș�Gǟ!�yR�S
͡��	G�`�h҃���y�L�[���W�Ǯ@Ϝ �!�6�y�펇,BX��ɒ>�|�y��5�y�,I~"=�!��]�p!��y�b�7qn@�3�� J
�8�C���y�$S���S�X�o�����S�y�'�#L�L��D��cx�J�C��yo�� �I2W�W��M��`�yMr��)�ģѴS�&y��&���y�e�T5<��P��b��Y�CDG-�y"�O9S)*�� F[�bV�M�+ރ�y��^�:��!߻`�*]���5�y��=z> ��E�Nn�M����yr��>J��F�ÆyQ؍:���y��G<T��8���#n+VE�sDؓ�y�)�:ZP������3#�Ȥ�y"��c p  �P   �	  �  f  �  3'  �/  �5  <<  ~B  �H  O  EU  �[  �a  h  Pn  �t  �z  ��   `� u�	����Zv)C�'ll\�0�Kz+�'M�Dl��$?O0=;��'��+�j�c@9�[�F�h��wiX�.3�p�bę�wwђ�Q'<���3  b݁����?��g���?�8AV	g0�%O\z��63�x!w�V
Lx��M��g�‸�ʒ{� �;g�b���'�?�j> ��Ũ���:Z�p"HD��ޑ_����I*���m��%���ݴ�h�����?���?���nD��JG�Q&��h�ě�b��y����?�i�2X���� Kh��I០��;F� ӢZ�|M�I ����x�h���՟�ӯO����w|��D�Y���?U�C&	\l��e�E佘֡^~�<�v�߭r9ԭ�K��8XG'@|}�>O⟨sKU�=�'�
�)����i�̝�W�?bȎj���?���?����?���?�.�杗��)�p�_�K ��c���Ĉ����4c�ve�>)&�i{�7��٦�R�4�?q�� �l݃e� 3ѢIR�mՒO���x����' ?RPzF�f|�����$(`��B�#U�#a�9 ֧M��z@n�#�M��i��3�P�
c�ï	���Bh��Z��8���1o)��'� ��%kX�@DxXs���?��a�B�+Z�� �bf�>hnZ��M�f��j߲aے�\�`�c��Y-2�N�5"Y654�a)b�it27����,�$0�4�� ;g�j�`'Bx��!�<�\CsB� '��q���5.� ��`�+�M[´i�6mU�`�I��'����V�3Y^:v�ˬ^Q��� J�>&�a:Fb�⦥#!���R#�D3 �J̚�����X�?��L-z7�!�,X���'-U�,��Т3� rU���k�HTo��?Q�� : Z@f�:?s֥�	]���3�@�r���A����Ҍ�ȓ�! �ѯ35�9��2�:���&`�E�Ԃ�-0��L��[�_*���ȓ��n����f�* F�9�P��a�<�ï՚{�4�p�%�J�H6
Ri�<�'�A1}jHl
�L(i�0�� �|�'��)��qA
�Y�D�C�����'�9!��� ���M��2�H
QE1c!!�$X3qd1��5��L�Qŀs!��Gj��9X��P�e�ND�Ƥ��R�!��Խ,��ݳ&+�٠U2��A�!�DP�*��a;UF�1Zk�Y���!Nx��	�O?}��h��p8f��%�5��p' U�<��!Z<6	2�B��Aa���R�<R�H�J<����l �cT؊��C�<y��S�����!P��`�z��y�<�@.[fB�Hzv�Y"���Ӕ`�<��ޓ,��eP�-EF�P��k�]yb�N	�p>�A��s����\�_{Y��l�Y�<����h0��CM.t�ԍ�e�V�<1���QBeř�X~�@���j�<�U 	�rH�)"�C!&�,J .b�<���޿. �R��d��I��IRGx�4:��� �M����?���#6��a���?WBT������?��
l����?���6]6���W`�#������+�H��x�L�(�2���{@��'3�#?�Dŝ�}�ԭ�T�B��T��'�"��"# c|�H#�ކ>��%A��(F`�<�r�ϟ0��1�Mk�GN��č�:�r�#򭜄
@l{*O���<q���i����QJ�.yB��� ��)��nZ�y�`iKF��(�հ�n��������شL��x��?�.On�9O�[�lij�A���z4�3!�B�$�p�8���a4*�)§Iֈ��үFĶ)�N�$j6	�'�b�
C��@�S�O�T�s���N�.͙W�ޚ1:P���OvU��'Q���iL)d�:�����	�X�6�F<9��'���'�2ٰ�d�(.�he$�r��܆�I��h���y�
�&ae�DiUL	:'��`��KhӮ\"��<�fE��B�g�'n�����q�"�q6oM8$>�|Y����,�'�< "��ǎ�Ϙ'h���eJ�`u�	:W��1���T�L(�	�5e�"W%,�3�ɧ�(B���+tʸ�	vd9Y���+?�3���|��@y�˽!W������<�,���!�$��������=E&��������HO�	�O��t�b)�B�5nW���ā:1��ٲ��<���p���e�j��5Ҳ ��T�A�B��?�ЖML;+�D�A�ڑv��$ۑ�&����+���ɥ�&qȄ�r��ɶ6�4���Z���P�J;t����8N�g�!D�8�d�i����K�L�0�JP!"���e$�<{3g�)��!a�g�=��2&fԆ�B��IVy��'��'I>e���,�@	�W��@M���� ��yסA,N�H	�Q*V�m�|�W�'�/���C�
��k��	GZ�)6�Q!�tf�XC��?X�x1+�OD��ORܙe�'7B��Ԫ�O�*|��1���"#�����!��O����*{�|(A�J\� {:h���H�2�O�ɀb@��N1|�c���x�0��E�'�Ƀ	PF��ش��'��	�O,���ַ[�.�P�#G���њ�I�O��䐘rN���B�۹3�P-�2/�[���2s/�� �r��nC�n	��{��s~ZMi��:��d�z�ل&��dM�X�����E��p�d��qZ���k~��ޏ�?Yu�i�:6-�O�#|�QI�?((z��A���c�R�I˟|��I�t��p@���4+Wz��׋�G,�?�4�I^	�KW��P��%�J��E�ݴ�?!��?ѵ�ݷE���A���?9��?��w[
�YPaD�P���pjC<h����/O@���;�d�����.�Zъ0 0h(܈s�\�6MH�*X�2z���u�1����D�3�s�[���5�̗,�Ҥp�R���3����:�<���po ���(�,+x�<�=.*Z +O��=E��dߜ+��%�3Ď�v�&�"C�
��$�֦�a޴���|b�'����$��%&�L��%*)C,�}�'l�!2����O���O�O���'�2Irn��Z�X����Їn����X?N&`[wN,O8�C秛����`�I��5�ʙ(T��� �g�L�`)�-Җfо�ۗ�
�t�צl�������U�Q�DS%���*/�!��ƩO�H�A 8�d�OЉn�ȕ'<�_���O,!x�I�y�80cVkk���K>q�Y�Eٳ���tuAԁ �>עU�I0�M���!����'�1�rO
��dC#��I����43�RY�uJ�_�!��1�+�U�7���s�ɶVF!�䝡~,����X
�*`��8+!���;>�AA� [��I��Ȁ46!��3:8 I�0��0�~�j�T.e{!�S&�P!!����(D1r��0Arў4:ch6�MF��CWA$�:���v:��ȓPx@⦯C2m����e1a4��G֨z��:rȝ�n�"��-��|71bT�߰MU������'��ф�i�%@�J�Lz����TO�Xl�ȓt��!Q�� k�ʸbg�� I�J��ɭJ$#<E���|�v�'ꃄ?|�v��3+�!�č+|���RW9|噀2 �!�D#;��\��H֑Ռ��u��W4!��
(
�B���CW�L� ��AOL�h!�$
�C�J�1'�!S�H��Ã��U�!�$�zf^� E�O��8�t#���ɞ9�����??�ArK�_~��d#��K�!�D�J���R3i�> |�!x��"7�!�ě�&�6��jŽh��G�6�!���-�I�R�O�U@�(c�G1J!���'.V����� ������K�*T�}bB�0�~�d��P��}�3�<S��y��'>�y��ҧA���� ��
YB9��܄�y��0gY�{��ĶR�����yaS�C,�Z�.U�� �AH�y�bP�	[TAI��Zw��-���G�y�� sN�A���?q�R���M��hO�����5=�ja��\g��[�)�f$C�I.A���H�7n�,|�@�A�C�I|@"gd�?Jq�2��7C�I�!�؋Ԍ�>�D}�4�F�	�B��>ql��i���>i`Xq��剈S�B��;<�@�@�WT���L��/ϔ�䋱��"~5��a�*0I�D�F��K'� �yr-_Z)
&炙p�h��'Ϙ�y2�;TqJ!�b�L�n�x���W��yrGV�~eV�6N��=;6�h�֋�y2�J<b��rn� `��iC���2�yR�D =��l���W
��)`tgL���� ��|B� �P���ӀH��H7���y
� �$j�&�4DK��h�'�$��@�"O~�A���v@���R7K���"O��2]Y	�QE$K!>}� rC�X�<��+O87��aJ�E�{8�H�6��zx���E�� ¥ΝG�����s���h8D��"��ˬ��Īm�L����f,D���d_<"<m�6��5Ug��s1�)D�tR�DY�{G`e "Ύ�2��	��C'D�X�KN(Y�Ct�K��& 'D��!n�2���R�*K.����C1ړ:ٺuD�������F��_� ��"B�y�cT p�!�1̓)Ԅ|I h��yr-VuS��q�"�2paj���I��y�
�~��gd���X<@'���yr+O�V��)�#�U@4�,�C����y�oM�&�HQ�S?"�e�����?��f_k�����(��*�0a�d �MY�x�H��A>D� +%�D�m��/O_�e��g;D���&�.ƹ 
�cUJ��5D�TëѶ3���b��Z4tW�]B�/D�����ԡJƨ��(�
T�)9�',D�Ҋ�+h�,4hr����K#�<I'Oz8�iaF�g���k�����A';D�Pp`��/]#V!���C�J�*�f8D�p����z$D��8��Bb8D����,�8[K4�{�bCr~V�(@7D��* ș
+	���U(�#�J�[D�6�O�1���O�=*w��`�fX�S��P�`�`�"O�;g��@�Xm(� �i�&i��"O��1D��Z�|�5� �HV����"O>�s�@ܧw����A̿/���P�"O�����r�d]�.B�=�.�HQ"O��O�<�0 "�޺PP���P퉾:��~�g�я:hj���
+�۔�~�<�΄<�T��6�ײd��5�իR�<	�	�'.\��a%�6:`�JV��R�<Aᢕo��� 
[U��� �V�<�`F~k2d�m���ցQ�<�Ѥ�/r��I�+�4 ��ͫB�y���>�S�O�FH D�Χ%<�岵,Ҵ9�����"O�)�_�I�P���%ˤ|�̭�"ORt!Ǆ�8�`�Q�I7����c"O�Y�+��=$-����9�d���"O��!ڭG�b��O�Kjm�"O��
ՁD>GD8�!��{msX����8�O�x���R�$`3̀k[ ��"O�u (��<%��J�A�t:��4"OJ��c�A*�r�9��ʋd_(b'"Oּx1@���U���	/e����"ObѤJ���ї�N�Q"e�U�'�ܘ�'�R�;�Eg�ƹY�̈́U�ʅ��'�"Љ���? ��e!�-@�b%f٨
�'��ISbMf��=�ĄgL0��
�'��q��, ��ы�FF��b
�'�F�S7�p�ޘ����"�,
�'Y0��Ro�X�F���,��X my����sQ?-HsmE#^I�h�VF��t��3h+D��K�P�U�Bm3FNʛ2��sV`5D��qp�(1�6@s��1��aRb�1D�0&gV�drĴ�玍�e�(�B,D�$��!>ک��#�����zsn)D��`a�#J�A���$d��Cf��O��y��)���8BF��$'�rf���M�Z�I�'D��R�ĎL�`LZ�)��TdX��� �ђs�6g�vL��̔�s��	�C"O�S�J5�2��Tk���>À"O�5yV�Y�!�|��i־-ݶ`""O`�f#�<*
�Lr2������S����&6�O�9(B�	)P�RA�5
<:ϲ��"O�M0R-�2��	@T	�q�r��$"O|�%�`�̀�g����B"OF��4F�|�����ř���K0"O�%�T
U�2�`�У��8��'z��y�'��+�FZ��4ň��̾	����'L	��4]G�����5��P�'/Ґ��G ơx�jͬ*�d��'6�Qؕ����pKч۷�6���'����1�ѧ^�����Ź?�}	�'�.,�)�(!w�	���b+tpp��$�t�Q?�����7@��{�*�-&%�śC`,D�|w��
Lxh�y!fY�,�j%��K)D����P�B����eU�B�RQ�'D�k�)�捻͑"�J1�6�&D�`Q`F/D�y�� ��5�G'(D�L�%��n U��oN�5�ȉ�f�O6!��)�'2qh	Y�+�A��h:0��'����K�:�x�b�hR���'DިJU$[����yR%B�KI���	�'�d���e�.Q{Zĳ���J$�R	�'/�z�χI��1�dԖF�̒�'~l��E~ۊ��b�#/����*O��1�'u؉�vjߝ[��P���+ق��	�'�J�L:"]`P���((\�%�	�'c�2�ܮ2����Q4��S	�')~+�C��+[���U�@*�����'�6��cDВy��XR�(9+fn���T��=�-!��5���G_,q���;s Y�ȓ|Bf�;�/M�i�HHB�G��h�ȓ`���+�l�j�j���G����ȓ�@1�U@["�t�4��,]ұ��p�xp��	x~X���P����d�FE�DlUc|��A`�C%㰜G{��F������P ��
3&�/"Xd��#"O�4*�K^�=ؼHC��'���"OB�����0��%z�:��<��"O�E�DO�(�j�s"�����"O���PAZ3z��5�![����"O��C�LЧv6MQ�ϒmq��T�'0������ӳ\��k@@٢ l��������$v�����)LC��)5G�V�zɄȓ[m�$a��[#O���ce(T⾠�ȓP �{׉O�uZ����
\��(�ȓnv2˳9C�����ZM�ԇȓI׮�YD�t�"�)P�HI��'��-��FW�A@��F�[N��� �����pӸA�"���ۺ<����( gy���<u��+2��=9 F�D6@��!�Qa�Z�HP �@PU�ф�yL����U�:�&�cA�D�݅�	-;h�I0��8e�Q�ƽ��e��B�	�2�b��R!���n@�X��B䉙b�����G�� �;⬞�tB�	�U���o�:wM���K�2C�	
�-��^�PS�t�U-݆+.C䉐%��$�B�D�9a�x�GO�2a��=�Ӌ�Z�O'Ѕ(t.��u��2��9��-8�'���&�4����g���$=
�'N�K��!�8E+�.y��<c��� ��@��&���ϝ�2�e7"O��)� Í�%I爔V�Q2"O>y����1�D�cw(=Z�V��`�'�A���S�;��D�pϋiU��9�A��:l��ȓA~>@��*�s�.mQFʛ����ȓÞ|� �)JX���O�X_���Q:| �!�JPp܀1��6v���ȓ@1�� ��:S������Ąȓ^)��3��>V�ʹ� ���"|*P�'�h��w �(x��T��qRΜq�깅ȓ �x	� S��B�,k8-� �]�<�S)�ɒ���L=�P#熛[�<I�͐�@N�BR#S��zp��K�<��CҰXE����EI�	���@Ix��Y�輟TxF7j��4jsJ��s���B�#D���F�*�������hÉ'D����m�_�4�C�
�YTB�R��/D�l膪�xf*u�фG9m��c�f*D�(�(MJ16uz$K�)Z(�5M)D����a��؄%�/l�rĀ��;ړ�H�G�4Ę&d�XH�)^-+?����/W�y"ԬM�lq�l�;�1kW Y7�y���b�Y�@�K�H%�F��y�jֱVkRM(��ۛ@�ū��>�yrjL&S��T��gM f������yR	��-�.�K�B*g,�h�rHG��?!5D�����8��ȓ�l �mX8�`*��?D�|�Q�mR��c҄��P�n��5�<D�ثd�6~5�U*Z��X�08D����$�hH��YS��d��p� /7D�k$M��L�jaAb$ӛ�$@ȣ44���ӃAu����$�ӣ'=���w�e���	/$X�����	�Q�°`D���.u��o�:>���'���'��g޻
E�i#�jG"�@�TnÇW��)�s�����$�^t����3�"D{@���4(�]���S�?�{Te �Z�b�o͂SO�,��A=�}������d�|◡Ӹ&g�:W�K;��!i�Yay"�'� �`�/& �vMq*�I���6u�I9f7�x:�E @��A9�
�j?ʓ9T����UT s����i�Q����Or��w��%3-�&�g� ��i�O�K@F�J�Yz犄�_��\�7�R>����S�<3d�q� �8l��橂v��D ]�؉2��J��Lm�T�t	��i�?v4SQ*�G�I"��c-�1���'��)��4?IgL�4f��0�dOѴ@F�eZ�n�<��@nH��D˙6��	�t
j�'WL#rCn��� !3�͈Ya�E0T�3,��(O�9Iu�զ��Sǟ�	{yr�'����ܗ��T�_}H�SgU:C���e766qk@"!P�1�O �O���#�	�i��j��P
t��&�D�{V�ip�f_�B�nYT��#Lw��e�&z�:b�8'�k��G3n��0�'I84;���?Y����'~�H�]���s@;Q��"���<a!�$ї4���Ro��M��xy��7R�1��|�����$�.h���B���#����څWl��C���Od�5��Ol�ĩ<��S��չGf�� ԧF;m|eC2�M;,B�9H��^���4���[�m�c14�Sޒ$�1JV�Mk�D+�$L(Qb�QU���hm��-""<;�H��O`,���'���IW�ږZ���1v�W�1$�](a�'�ў�F|b菨`�n��B! �|����Ñ�y�� �m�4o��y�J��nP���Dæ���`yo�= k6��-@Z�d~>�p��%S<�X(!�m!�-J4�O������O���O �h3�'@�)�̐���4�@tA'K��5�B� ٞ.��y��	���c���1m���H|Z�!�0^�0T��fv���Zj�'�0�)��?Q��� �0�L��04(lbB����<�O:����ȷM,q��ś���y�Q�''ʓ׌����D7*2<�Ѫ6 ���?1�&��'���'�R�j�Қ#�ڨAb��jx-y�'â��g��,	:�z (�Xh�P�' j]�oP�E	�Y�׉����t��� 6�Ӧ�U�t���+ ���"OV�!�/�=�6�ñ	�Vi(�@f"O�$���?��P(�1y\����-�O��}���p��kB�X͚���ú]�4�ȓ&j�!roխd�~�1�cКX' �ȓ.|(p�&��S����(�
!��Y{�!���
�}mԜ��'Ep�p�ȓ>w^���Y:S�d� 'ψ3Gp��ȓE�~�E%�%>b� �%O<[-���!%�,����r� ����0)Z�1Q��.?�!�d	؊Ejb�ߖX  @�ů϶ul!�D�]G SƋ����(��f�!�d�J+T��J/7 ��3��x�!��ZR�.%8C/�lA��c׻�џd�g a��|2� Hێ�i ��?Z�ސP��g�'D��p �WM�O�0$S"ъ�8�(�g]<���I��DRU!<�ˊ��Y�-�x�C��{�&�JU@Y�8��<[���O�8��\4�� C�ۃ�\�k���2/5��D�O��"~Rci��0�YSLP0V^a!W�����>٠W� �ES""ܻ��
:���xu��<���?����?�L~�/O4��+��@w�F"P/(jq��h9O��=��N�-��a2�R1@��Z�HDr��M�N<�r�8�5Nc䰈P䁡+�p����O�],�C���8]��S��'��q�$'G�@���<$�V�JwE��~��I/���$M��'(n��)h,� q�Q���*D�a�Dj���ɚ�~��s�<��a$\��i�cM�r����Kץ��'��'�|E�I�l��R	{��"m�\��ǈ�({Vѩp�'��%*I���C�.�'|���W�N�n��S����A8�M�ȥOL��O�)XP�>q`�i���Ӧ���U��5��!"�@��*OB��'�>����7B�uS���*ǘ��!�:T2A �'�6Q�I���<yR��l~�,��Sr��.�02a�Z���Sn(}B��6����>�H��	��J�/_,:A��8�h���'�XT� ����9O�� 1�O^ 7�^�Ƞ	��Z)O��|�s�'�\��	�e)x��H�%���@��PXB�	;M�2�����JC�i�Lh��b���d-���E��O��禙s����	s %��M[�SdL�5�>�K>	�������'8�Niѯ�5fc(�(�BH�s_�'�ўb?�E��/.R�3��>�p�6D��)!K���H��P
>T�Q�8D��i�*�'t�� �L:
��}��#<D�8� �Q�\���ʾu�it�>D����JK>Np��� g	�R�=D��P�nS�B�,ԫ��8/��q�O9D�`��)�&@�M�"Y=�U���9D�t:$`	�x_���0J������v�6D�0{�l��32�(����̥֦6D�p#�N�0ǔ0Y��.W���B�L5��hO�"�I���	߄M�����#s$C�	(��� eA "ar���㛒6c���ͅ@�Z��#����Ag�e\�,�+�.1p�qui�d�j�!��Ҽ�9�%[� �&���Lz���KV�)(j�P�o�P����'&��3�LxB#o(Rl3��0I��q��NU���B��3=�ys��C}-�Gi¢v��:����{�j84�C�c���f�l��ҷ��G��u�����?��	Fj@���Ib2́�G�S�� ��[�ʧ��I&/���"��
�]v��Y��	�(��'�2d�@�V�7r��C8�'XfB5����8s�,��;�l2���/R�'T�>�m�6?������hx��D�x18C�	�*��x��J̫U�@ �VLF�
��U�'�d�x��\�.D�Q`��E����O����O��d�4�T����O����Ov��w�@y�-��%�(����;�R8;��+�� R��Cx��䰣H�$�Bc>Y��Od�����r�V5�'m�8��|�eEM���Y��i�����Ę {�pb?�@�OP}+�_�M�� �'�S2i�,�	U��l�'-Ԉa��|z���-��`0$M�VA�+�����!�d^*y��k�#�Ea1���#�V����S֟��'��R�m��c�X	d�#4���'Z�q�Â�_�(4 ���!�x����� ti�f
�9��z��T�fp ��"O����H!<i<���O�F�(M��"O�PS@S o�[rI��^�v��c"Oj�+r&��5{"�rFV���g"O���EM�x���;(�
0��"O���  R�9`塕%�42�"O���FM�*u� )I�ƊR�6p�"O�!{��À\�����e6c��P�P"O�|p0ċ	��R����"��U�"O�Pq����b�(��%m�H�l�"O:�lO��D���4��L��"O�!@Өi�͐�jE�,�d�""O�����K�~��pSR��*R�p�x�"O`;��<x ��uϗ!{�=9�"O��S��+6O�5�獔�zW2��"OX�t�r�j�?l Ie"O�A��Méd��LRe�C�n�n�c$"OPђ����c�$�J\��"O6THQ�Զ\��Q��0{��u"O.�hT�Z̑Q��� &��"O]x4�1��`�ҀA�2� y�b"O���`�3 �th��'~���:�"O��dBA54�Z��.CU����c"O%����_�*�l�7DP���#"OJؓ���5H����+�#mR^Ear"O�����2l|Y�*jE���"O�%��c$W�
�RdT=H՞@"Oԁ�QgƇ=%�A � 6Y�fI��"OJ]x�Ȉ8%'�ɨ`��]����"OZ}�J��T��\��F�@p�P�"OD�h5�� 71@�9ՠGtkX�X�"O���O�!a��Aw�L�Q,�J"O@�+pa��k�,�����5��H3"O�ЀtG��,����!�-�����"O"����w�D%��a�->Q&�t"Ot��H��q�F-�!�����n:D��pTO�?��D�aE�z�Z���7D�8���/y9�	U J$ �(��6D��xD�R��uKS������8D��kG�+&��j�O>1A:)z*7D����!XP d[  /|6��G@5D��怞�7G�A[�F�;
�,Q+6 !D����Q��0��ڸ'�V���D1D���}�F���`�6D�:�!=D�,�C���=2�+ �4���U ;D���늂��(BϞ�^"i��%D������8	o�X2t� .�qXsk#D�hw��(7��a��α^���0  D���R��9$ '/�&� ��ы?D��P�`�R!��°�ަ�6/#D���l�0�h��&N�&UR���?D�8駄��g�H��L�FT0ف�>D�d�ц�,S���:6 ߾.d� X7�'D���2ι? J�X"�?{��j��2D�y#
��O*бsȝ�{��P��4D��crD�k������]�N���5D�$��	1ɂI9�N]�ް��s%4D�h9 �o4��F'Φ 9>h8U�3D�<���;`L��!���99��t@%D�Xd�S),
���H>����f#D���B�>�.QG,ƆDTJ�F�4D��/C��F�IuA  �Ҽ3"�2D�l� @Шh�
Q���)3u{Nub�'��ݐ��>�y�����+��5�
��� x d#Д\Y�83&��aCjp9V"O� ���{���J4�Ƣ{.���"OPDyc,Y<!�v ����d,�R"O|L�6dQ�4Q�%��(�.mvth�"O�����Q !�*����"G��hp"Of`�q��0%A|��'�
 [�"O|�(fL�$��0��ׯL���"OL$���:vv���D��8	¸)�"Ob�SNB2&�#RM֥Hg���"O"iw �x?d�@��Udf��"O҄3�.� 
6s��ܐ1a�aY�"O�]�񆎫�l��W"_�:?�+�"O�����B$��2�Z�:�"O�xH���h���� �2��(K�"O��Q��Ӓ��q-B��X��"O�E��O�Q{F)���U�M�z��"Ot�q��[�w�A�E�x����"O�!���y����J2,���d"Odѓr�:E��IA�I��.�A�"O���eMX!Z	 �ʒ ��lcV"O�8Z�(�6��q᷇R�Z{��"O�e��ѧ+S��c���!c���"O 3cN+y�p�v��8+UQ�"Oz�� $ײRF0�5#�yK¼��"OZ��LU�1�]���(H�9��"O��
�(wx��h���=V�hH�"O�9p"�щ<�~�q"�M�KCj�p2"O�Y�0`� �
�
�y\��j4"O�ɓ4C��8*Fm21iC�SRaHg"O��C�ęm�hA��bN�fX����"Ot(�A��Z�a� ϵ=��Qg"O��27K� ��� � #��i�"O.�d
ۚR�-��/Dwn��V"OD%�a���谉s�ƞv�&"O�8h`��-\��K!��1���1�"O�����\�½�sB��\uHs"O�C�,x��Q��6i�B�"O<#��Ĳ"��\�5̂�},��Q"O�±C��?V]�� Lo^<Ӵ"O��s�* ��3G���x�ۑ"O
 i�Oŷ].<@�^�9����p"O.�ڔ)!#�XѠ���*�Nܳ�"O^%0�*�-6��A�� � ��`ۣ"O4԰6�Q�S]�Ibb0(���D"O�83Ԧ�w|nI����s��M�Q"O�`�Ш$B��0��I�C��kR"Od�Q�b�Q�@"�"' x�Q"O(�c�Ӿ6e���"�,D�f�1�"OJ娷۵l��armٝ��(��"O����)�f�n��Ζ�Y�x�R�"O��6��op~Q�2G �a}��+f"O�I���%[̥0�f͐�*q��"O
eJ�%�:��)�5L�Lz�3�"O|�ȁg��Od6@x�/�"ya���D"O(���j� l��*'o�>x����R"O�ȇO�-/0I��L��&��C7"O�XRsҺ.���ڦ
".�A�"O|�rb�1 �p���Y�t9PYc"O��2����
I,8!"OzEh���~-��ڔ�*��e"OB����D�x^HZ��"f(��Z'"O���G�Ԍ�Xq#cD���e1"O�aXV�8F�P�a�b��W��3"OF 8�@��,x:�Г+�@c"O� ��;��ƻy;r9�a�D�j3�s�"O,-�@ ��b]��Ŗ��	�1"O`فᩍ^�蝩�A��dF)"O�pR6��0}���c-Iզ�H"OĘ '��e�@ϣ^"���"O	!W���RD�y���:dx""OPͲ`JO>޵Y��d��T"O6b��%e�q;�o��;P"O�X�t�W oY�����R��`�"O�eY�'�%�<�5���lA u"OX�B#�l	���bD�(]���s�"O��Z��=
�����)A�@T�u"O��`0dS�ӅVV��Y�j�A�'� ����e�x���Uk�)��'���aHQHh�@�ua�0_��H�'Zڜ1JL� _���	<Q�Tl��'��a�P�O2��4��|Z��S�'Aj 0pF�qI����d!?&����'"��
��R�؁(&��:��Q��'��E��!0uL��6j���'�z���m]2����B�5?RЈ�'E�P�O���=XT°#�����'�N�#���*s��i�sJ���J�'�(M!4��O��u�tj�'0��
�'��Q�c
�V]hu���Hv��	�'.\%b���O��"��7���B	�'���'CUN���e�*���)�'��ԫ��<bΥ�e��?*�q
�'��0*D�b)TYH�H٠#����'���碊�d�4�y��D����R�'�@�[3�W��� ��ʑ|���Y�'�l��QJ��dc�h�|���!�'^���������%�B��5��'p^�� 	�Đ	2�B�7H@�y�'pԠhuNO�foZ�z��(�<)��'�����ַ3�~�¥��i�����'����!f�8[���tM�Y�T���'peұ�5xv�0�B:K��T��'�x�C�+���~�"�#I�n��'L%2�BU�M=�@�!I��ʙ�
�'Ͷ@�wHI��Lsa��(P����'!�IY�L�XM�]C�Əx��8S�'����0�`)�)�([�j����' �r�C�8n�Q+K��3�hYK�' ���O�? �8�C��6wb����'��,0��3ͤ��������V�?D�H{0�1�̊�AA�
�ʁ�1D���"H�B;F,À�C�� ��;D�ta�R�d�����6<�q/D�x��ߤsh�B�I�z��	��2D�x+��U�y��F� B�|	1�*D����U�0D�&�Ŕ��Wd&D���C�"�����A�b%4)�I:D��т$ڥ28����
�=:� �;D�lH���a#$�f�`�;�/ v�<�D��5y�e+ិ(���!�)t�<Q6MY�K^f�w��0*F}�!�t�<�!��l">��a����F�%�Y|�<��F3o�m���ٺ�,|j�@z�<�&JY�[��ƝNw 1g,@v�<	6�U{�f�{��Mw��X����V�<Y����"��J2DS�M�<��n��/Z��i�����N�<a��P<	��x�H(<s@k��HM�<� F��s�S�l�R jH����"O���FEV�PUtt*�@�d��P"O��� ���u�,�Ё�ʫ!
��c"O`��t'� �H�[��ߥ?�,�0"O�sť�.F�	��B�8�����94������8�v�qKE"�,��C�	=�r�1w*_�7%�nm�#n�C䉤�@R@�זmN2���F2q��B�	d��A��V�0�h��2JB�ɕz~m!񊝐yaJd�W�՛jLC�I�n6��j��
7/��L���0t�PC䉭?�F�(u�D	m-��
��%D�B�ɘ
Z��0&턁7����fÍ�,
C�	V݀�P��I?j҂��G��?e�HB䉍 ��@RHD�tQD�(bkU748&B�ɢy�����ܞ���*Ԃ$	�C�I�>N�(s���)�|��c�6�C�1��4��k�
s���e�_�LV:B�I-Q�r�P6cH�P�z��b�[)d�B�I�Q!FC�=}�NDȢ�܅D��B�	&L���I���Ufb�ɖG(D|C��j�`9��s�X����Z_<C�I�nl4�ˣl0e[h=Y��Z� C�	�L3�P7G	3c`DU�3d<�C�ɶ-q�	%jr���qeV5"��C��8=��@u��ݐ@m�1f�B�	�q����0hR�>tU`��Y1�B�	XiA�c�F�m� �!�Yn�B�I�+�R�8�-D0!�0�9wDC�ɴk�Ҙ�+.9Q"ԑS��8�jB�ɿu��T9u�f� �� �ŦponB�I�j�!��bR��8Ip�,��'~C�	3HN�$Z��Ӏ?,&����A�)�HC䉳:��)F[�9�F8�l��u�B�2[N4���
ϑ`�d ���2�B�ID뺱#" ��"�B�JWh��vj�B�	�z�a��P�aE������
4D��[$*Ŭ{\�� ^$C��c�/D�H��"6i�Y��F�j\<qB,D��� ͋E޼2s�.]�"�Q�2O�pK�'�!+銉@�MS6kOH��
�'Q��S撀sE�U�Fǵ:�a�'��4���R�8�q��ߎ��ĉ
�'9�hP�%WY�Q!*P	.<E��'��]��cZAo��x�,��L>=��'܌�e�եTB���8<���x�'&���@'V(�m��/�n`��'gH�b��ע\w�h�����L���'�򜠡��O�2@�EW��¹��'���FȸlZ� ����r1��'�R�S��ƟQ�v|˄�V�2��
�'�*�y'˖%[��}���S�N�p	�'ǤU�χY➠c���L���R	�'`\�Y�'ϱd����0�GD=����'D�(�0+^:s׀��-Lغ�
�'ql��L��;�qC�ЀXl�݉	�'��Yx��I0-�퐲#�!O���'��kH�P��U�K�!rR����'8��I��,��` p�ݿo�	{	��M��hٔK#Tp���R�}�
�х"O:D�cdC�Th��K�Dپ��"O��Uʍ�`�R�B�� m2�u"Oj|����E⑨��"A��2�"O�1�c�F��TK'�Y�g���"O� @+��@�YfH����ilX���"OZ�9U〖}6�(�jT8L>��F"O�X�b�(r�P�`
Ԕh-Q�"O$j(�^DP���2;)h��t"Oju�A	BŮL��P".���"O�� FH�	2<m��l ����"O� C�,(s�4�G�%q�Y�"Oz��!Qm}�$`G���^h��T"O����ձX�`��7V]pu�"O��4,
�	/� �5@љ7DxUZ�"O���k��. `A��" ��� "O��9�@ҕ-�|P��(�\�8E"O��
���	%�(=pȂ|���S�"Of}�l��x5aC�]�,��"O�h��Ùf��)�C��V*|�
�"Ob��n��&��r�$R��"O�1��D��v8^i� �?�"���"OV���UH� 8� ο<B�p"O�i�G/��pz���ٿS�=��"O��S�T!s?�U���&-j }�r"O� �F���!����A���"O1��MފO$Z��­˟)�b��"OR�*%�֠&����8t��`f"Of�;����y��X�c[,L��r"O�,�f�-6��X�	�5)��;�"O!�gc̑MD���Z�	(بf"O4aYD���Ē�����<���"O�0�ԅ�"X��)G�+8j�I�"O�䙕�ߘ���CE�.1�Q��"O~����_	�MB�A�,���"Oڥ����n����C�X1$�1�"Ol��`�T�~�����a�>7Z���"O�Pa��%D��H��BұY'�8��"O�$����ehl��㇂*�RC"Ot��d�f�$����-,)��"Oh���,ѯx]�F�� nݸ"O����R$]�A'"�z$�"O̠�âG�Iȩ9���H�2�Y!"O�X��gٯѢ<
��Ϗ^&��i�"O�k�D��3��{ �M����p"O��a��z�����ݦOvM;"OHa� F!3]����f ?3 �x�C"Oh���*�0��T(K�Rт"O��yN$�x�[A/K�>l;�"O�!��M#"� ċ׎�(TP��"O2��gȝ������,\�p�'/�Y��_>�����e�'52"�x�'QB}���ʞOT�y�.dF��[�'�.�*S�G�aDD�����ԣ	�'l�h��6?<�$�Պo��#�'�hiY&(гJ��B��	�$9��'BB�kp�M�Q�2�� �v����'�����"�!d�H�3�j� '�[�'`��JW΀�O���(&ϬB��Y��'}�d�&m\W=(åȏ�RG\�	�'̤���`Q��"PI���#P�����'�"h����*{�U�t�C,@c�p�'5`u!E-��ݛ�k@F�@P!�'��U C�I\p�G��7C���	�'':D��J�����v=�A��'���ThI")~݁F���f��52�'�h}Ƀ�1=l�` �$�b@Q	�' �a[��gN �q���2 q�J	�'Q@��J�+�v}����;��hK��� ���0�\�YȄT��Z�p �"Ov 8���(;�jir�샂:n��R�"O��X��k����$X>�J "O$@3�B�t��KS��.�p�s"O^��`�q��)3����ҳ"Oƌ@ƤM�\S�`24!7 ��A"O^��7��z	$=٧��%w ����"Oft��E�fR��C ��<���"O\Q �h�h�|�"��W{X͈�"O��Y�l��u�p��/U�Yв�2�"O�����IF�����n6'x���"O�ْ���6U��%.F�e� ��"O4�GH���mCCP�!m���V"O�4-%��8\�r�f|��"O&�Iԉ�m�B��VD�x��"O��hJ<F��LJ��Bg��Q�%"O�9��*ΣqŖ�*��C	��!"OR���(������o�)e��傰"OQ�ƫʯy*�Yǩ�!y��11W"O����K8,���A(�&�D��"Ot@՜7�Ll�]	�J�2��Qp�<ɢg�L��;��ŞsB�Prfh�M�<Y�	�]"�c�eO��� D�R�<����./��r�H�a��|k�� u�<!�.���s����Q
�E��Lv�<��MY�q"�)P��&7�|�AώL�<����j��$ab��w�)�祋O�<��I�G �XRl�x�<�2��M�<!Q�׌lC�����A+��Db�<�Q�ڍ9��4�s����lYs��F�<A �J�����K��F�p�B�<yV�Q�d9��"�>IL��#�PS�<!%�x��ZT������l�m�<��A��Y����	�P�k`ODm�<�����$�Ѳ��f�ڠ�C��C�<��`"���@�`B+	����IA�<�"&
I��$�$��	� ����u�<��ɛl����'�AsDؐg�Kr�<9��(, P&���;��x�4�Rd�<y0ҿ��$%�^0VH&�]�<1&��%+�ҭy�J�8��=I�N�x�<)7Fܷi�D���^�Gr�ؖ��s�<a���?v��۵L���DX�fFd�<�@}���1�ϯ4��	P'�~�<����RZh������ua�`Pz�<�w�Po< h`&/_��#�_s�<!b��m��R�-2'؀C��e�<�a؄K�Iv�\u$t�cĊZ�<`�JMx�ڄb!/ȱQ���j�<�Dł� ����#OLDٻ���i�<�dƜa�Bp@�I�`͜eC��@�<�E���;w8irR!�G���q�͝_�<�+`����D�N��M�P�PY�<!��"p���CJ��RT���Y�<�"�΁`"I:Pb���S"�X�<q�BZ�njy����!A����W�<��X����C��<N����g �h�<yq��s3F`;�Ѱ�L�H'�Ue�<�7��H�acܑg@��A�H�<1��$?��!K�@Nf�`�p��|�<�Ă%-y>�j�s���`�Q�<���������~��-ZQ�<)���(XV�;6�IZ�μ��jZP�<�I�'�( $�-xF�Z͂F�<� >1a����x,�]x�L���N� �"O���뉘]�P�A��]��X]�a"Ol����^�x�X�#�NS!w��T�&"O��:��J*'������u$�r�"O�(�@�5[m(�	���n��J�"Ov�����=�(���']0�s"O^-�f"�10�H�PL� e8��"O5{T�ӹWh4�NA�'"hS�"O��CD�;Ƅx���_�g�8Qs�-44� �%�R�FRp#��f鮉��H/D�ԫ�^�8p
��'�L�\�q�,D���ᤂ?��(���'�(0&�,D��󡆉�'�P�'e�	n�h�D�(D����v�S���'l>��v�%D����6s�T����ʄjD�(D���g`��b��$H�:d�x���##D�,r��7�U�Th�)=pc�C=D� �(6_�\;�	*vZ�m�26D���!�՜dM�ڣ%��X�240d�1D�s��3e_U1 � x�*�:&i1D���.���"��A�b� �G�0D�4j%�� )dE��\�*���/D��CAK�%��`��G�]&șw-D��1*'��=hQ��.����7D���˚$�v ��/�D2	�&2D��+�è{�4����x�(��#D�<���
* �����I���ZP�>D���&\����xM�H�t����yB�ĕ�4�*�m�7�z�x1�ܔ�yb��0v��pf+K�7XQa�ν�y�H 3]���+B#_7tB��U`�8�yB!Q���h��B,2��}�E$��y�.x	�VLX�&&�������y�CIx~T	�/��HQ �
ӹ�y�ɗ#F���*�e��e&���y���.E�6ݢ扃wZ�PQ��F��y���	�n�Xt��DzPX���SF�<I�
�!��p3�L���l"d�f�<����(�i+��N�Y.�h7�c�<!���)VdM�¹j�d]���\�<���-e�������-
�]�p��<aU���@Z82%/�Or}J�}�<��Qo�d�з��'L�La�V��@�<	��Ȟc!P  �߈<��4��M[w�<�4_�wS p�Մs����j�<�񡈁q�.%�@ʇ)V�PA�!�p�<����3��l�f*N�f��e��So�<)�
5.Q��C���/K�0rւk�<)�HC:j#H�Dɞ�x�Ԥ���Qf�<�å�?t{����fd�QI�,�i�<�+�,V��:�-�J��I$�{�<9�
y�Xs�ևI|��V�z�<Q�ݔ;.�l�!S��ZW�LP�<�l�!%Z�hB�ĺI{8H`#�_v�< a�;¢�����q��y��"Or�<Y�'�PT�Z���)i*l�XF(^l�<Q�!��@>���(}�`�ৡ��<i3*�6F1����ω3AF`�b��<A1�W�a���&#�*���{��}�<��,��\��Q�wT�	� ��y�<	���)$�H�kE�[j���h�u�<d������C@�v�PAbd�s�<�c�_�w�Ͱ�mL�|9B�p��l�<�p$�	����$^.�v���n�<� ��kE�nad��7�͒@6r�""O����������Z�AK"O�CU�^��N�6�(�qa"O"$�q��q)��J�Dܢ`�b��a"On�I����p�āϽz��<xD"O�4���q&���Z�p���"O�p��T�K�)���&i�麧"Ot�nF�)C��'�R;^��"O�(�g#\�:�铉(���"O��٧X��c��k�"O8���oR�`J��;W�]�5"Odur���
5騑IDd��t�f"O�Mq��#�.!K��Rm	�"O �cb�WwIN!!�_b��"O^�yG�·X�B���MWW�Dj�"On��CÖ7'(p�b/I�UB��"O�m��K�_ϴ��1n�&'EAs�"O  ��a,j��/$��	3"O� ���G;9?4r�
X!S�a�"O�	�u�$pO&1��F�1ad���"ON8 4��t�(J�Y�.T�A+�"O0�Q!C�����"��5e8�8""O�QI��;����΀8t&��"O%�,�=1�N@�!��s�z�Z�"OZ�:�I]�!Z��t;�4��"O�}ڶ� >"8�M� ֢a�"O��y�꓾:���׮�_��#"O�@�F��w��LO�B���(�"O~����N�Q�<����f;"OT���g{�s&�fD�bbj���:�fx�'!U'R����D�!t��T�ȓ.����,�Jn.}����A�5�ȓ]vA���P
Ҍ�F�M-���ȓ	�q�2 ]4=��1@B�V�k(��^��t*R�ڀ�8Y;��
"`�ȓQؠ��U]�p���E"!Jԙ��;Ӓ�m��b�	 !�:1��`�+ �������Y�Up���YI�0�I4_d-����1��<�ȓ	.��!/����)_sEC�I�A%8�Ӈ��mC��J��H�ȓ]l|]��oW�~TtW�pD�ȓ}i���P
_�V@��茷o���klX� �؀q.�i�J*E�R8��8L�ܚci�NUܭ��N�)V���ȓ$wl��b��N�&������1%U������"aۈ�i����(}�ȓ$���E���{��	#Ag�Z	�ȓ'd� I7���j\��A�ӻj̢̆�*�,8��`�'0t�wF�8I��ІȓW��3�@�w��=˔F˝W^�Y�ȓ%D2��c斻.���D�i����ȓ_U�d`DÔ-
h�����/D}�-��@4�X��K�^���JV$L�f3֔�ȓOf@��dR4d�H�Q�I�(�u����ݑr��j?�a�2��&q̬���/(�! 5B¬��ذ����e㰽�Ɠ�l�b��\��<��
�'��x*'"���Ԓ�+�� �~L)�'(FD�̕��xM��������'Sf �и53�� �	?�fDI�'��,�2BV�C��U�VBX�$�K�'�pC �+BH����ٴw��8�	�'6^!�@�� d�>�[�m��x���� �Ţw��e�xq�C%�|��T�"OA�+F�C6Uæ���"Of����	�DJ���gbV��"O�5�LÌ
���p�+��^�(rR"OF�'��yGxp $E��*K����"O`�ҁ M+r��&MH���"O@T�@í*��XF��@�ّ�"OzaK�̥h,񀰧D�� �À"ON��VJ��B0q��d��4+j�9"O"�hR�;:�H\pr�
�un��"O�M��������#+��L�a"O��X3&G��@{Ce�?�J�Hs"O$�c���o��}x�DD�v s"O|��˦�>p�I���T@	q"O�[' �)Fӊ1yeF�7U��( �"O ӭ��P���>5�օؑ"O\�Q�_�
T$�&�C�I�� 9�"Oz0�oԊL&�|���q�(DC�"OhY�Ѩ�<~
�Uy�`I6���'"Oni��@?"'�E)V��p�(I�"O��d��7e�@yeI�w����`"O~���a��x`֭�2�R�d"O����CA-��t�S��wrT�2�"Oj(+��+E�X�*Ņ��P�ʔ[�"OB�!V�Wm�u��+`v�C�"O�Q��6.���@��	)}S�D0�"O�h�J�%��i!��܅VN��H�"O��sv/Ÿ4��6�	�rP�4��"O�4"���2�0�[PlMtU|�@u"Oܼ�\	wp �S�ǧ㢍R�g�L�<���ݨ5@�ت��#-ƶ:ѭ�P�<�D�Ȟr$��C.��>���@��M�<e�=UUBo�� ;��U�YP�<QT �� �Ƥ�w�Z�v�Y�g�JL�<�R�}�Qئe�"VϤ�q�E�H�<�_ d ��
[t�h7'�A�<yK_�P�{��ȃf!�<pmB�<�w��GY|�Q�W�wTP�R��U�<I#i\�&|b��e�Υe��xh��KS�<QI�5E��I;��&weP�3��S�<)c�
N]p�r�A��5�DQs�+R�<�R��'%��m���U	��Q�<��� �4��e�
!NT8���\D�<�v��&zk0�2�[�(Pe[��@�<��?S�la�d�\;>
L���ē|�<��m@,ڂ<��%�.^Ш!@MZM�<u��&>0}���O��r����YI�<!T�jMZ����߶i=�m�p��L�<�Pս�:TJ��66�\�#"�H�<A	�;���� �ܱ.,~���G��<YSb*e��a�-X�D���LJ|�<	U�<f���'M��T�� �M�<A�*[ w�f�����QԨ2�nKn�<���a>�`kV#R�FA�yz���m�<�T+�$,Ɯ
FS�4Lb�8T��0�[��[���*O4�����y⃍^]b�{�➖'U.qVG��y�-G(NN�����1Lü��UL�(�y���#��r�����	��y,��'l0yS�
4H�!ĠM��y���1h	��װ6^��e��y�����6ʊ�8��]����yrMB�Z���%�G�6�P���`��y�0֒�R痁=cN}������y
� �����E7��A�d(4j�Z"O���D*)���v�(Y]���"O@<+!Q-B�>9��b�1=K,"OVpa�R�K�.���"ٔ1�T2"O��QN_�.�V4 Q�S�LH!"O�"t��^X��W��o>�Z"O~It��7 ���r'��k!v"OԀx�hߦ;�T�q�g���(HYB"OA+��DU�Q�0�U?*�	ʡ"O���O[�XKsǐ��@q�"O@����2f���C���.�[4"OD��.�{frt�(�'9c�1�"O��A�%"(\�ǖVh�R�"Oxqi(r������\y;�"Oh9��(׾wQ�(�M�,I�)��"O���JT��\��U�'��Y+6"O��ۢ�LaXڡ�GA�u�p�1"O� ���qh,<�������"O����K�m�lӡp\����"O�i�$�]�k�|��r�-dL�1"OP�Sv���р�*uJ� 6Z���"O��@c�'g���hF�$Rn�u"O��h�c
�1��p��L�%-A��b�"O�C0��CQh����ND�˲"O>�N 9%�!��,ֳ	/|Q�"O<�jtJ�3C�Q���S*l�0c"OR�h6�K�ʰ��*�Y�9K�"OH0#E��))�Bqb��"w]|��2"O�@�JA4#¤� (��F �R<D��SGa���1�"�S�+�|!!�8D����픟)����P��|�'�7D�(���37����D�-V�T1iu�9D��B�\�&z�HY��T) �4ɓ2�6D�pJ"�H"Iq �&=+���dL4D���d\�N�Y �O*j�\��3D��;��߶T��T��R��P�I�%2D��qc-�	^Q�{V��8lB,�G1D�T�PLӘS�~$�VP)+��A�k1D�0`��0"P8�ÎZ�Z$�	�&-D����G�<��"�ϙ�V©�0D��"�d�E8�N6\Oj�aA�-D��1�,6B�0�͕=	Bt�D�/D���Rf�C[��(��H��`-D��*��t�����G�"���a��+D�ۇe/B:�c��$ 3���pA'D���_8C`�9g�,F�d�a�#D�8˳a<E�0qs��^$&���(Ui#D�4C���*5�,�A蚙rЦ`��?D��P�F�7���	��Z<Cռ93C<D� �'��
z�p3d�7q�^m�ѡ$D���L˚%G�c��<j���K�-D���4U��Ss���hX��r�.D��`dɽT�BF��H�@u�!D��JC���*�꠪̋s�D��,-D��0֋�&�y�m�B�:4(E�?D��H�)S�qVZQ��B^���mB->D��S��vy`��6�#(�����`=D�䳰/�N��M97�E#M������9D�j�3q ��I�(p�8D��BS&���� � ��u��"D�4rB��0]|@l�M  4�x g�!D�x�Q S�%�!����4�T\(%�>D�d)�F�tal�૏�fH�%�<D�fB��
zUj��75ӊ�z�&D�� �9���Dڤ��TW�z����"O���g��[5@a����.�xd�"Oh�& �:��D8t.{�d�%"O��+L9&�����S�MY$Q��"O�Qb��-�J��/G��DA�"OXL�o��o"킲�H;q��Ij�"O���U�ЫW��B,øh�ҁ��"On(��O�I?����z��$�w"O� ����@�!����N}�2C"O,�Pլ�@�L��k�df^�3�"O*���,H�d�l��pVb��"O�0���3��JC*Ӱ]�j)�"O�c�#Ns�M#I �c��1"!"OB(���,+Â�1��C�82:%q�"OJha�i C4Ib�G�D"O�x�k�"\� �ݤz4\ {�"O��4m_�e!��� .R� b"O<DC��M%d�"ކy&�i9�"O�٠��J �hl�" ,kt�6"O���D���� c��.��qs"O,t�%Nނa��t�g#�>w~X �e"OZ��!V�x�M߭Ky&�1""O�e)1�V�yRn-���F�YY^�{"O(��L#rx���*��u�6�J`"O�s$ً^����>K.:�q`"O��se��T({TA��B$.c�!�$؆|-z)��� �.tq�_5$�!�D�6{�$a�� @�3І՞J�!�$ Sq2b��'eHl��`���!�N�|a*g�ەH@��6NA!�䕖l�2q�F(�L⢉crL�eS!�Ė� ���w��4��\����jP!�D�b� x�\u\�T3bI׺@�!�$���h0�6�\�@!c�BX!�$��;���s����@�:���`x�!��/^H%��\�_4�Pj�
6�!�D%:s���3��.c$��֍"�!�$�0����IؗO��ن�]6O�!�Ġi=��B��>C[d�I�*�-\!�Da򁱃�D>TA2呰�D!�$�:dN2��c�e4�lq�g�H�!�d�,H/���I�{�	t�M<!�ǌ��ݸ���(U�䜻�� �x�!��F�ac��� n����.W!���֭
�J�!8JBP�$E!�DO�#��٨�-�)Cd�c���K'!��G�-� Y
Rvs�B	I!�d�%+6�؁6��kG
�(��C�!�P_���P��f.H�T#Q7$'!���
�|�Q�$M��\S�[�Y5!�$\lZ¼���F�1��Qh��b!���r�x2�
���x`�a$�B!�d�
HU������D���1�!�$��^�p� C%:�ʬ2�J-�!���hrؠ�!��PU�J��z�!��K��\���Ÿ;?�,y��&"�!� lBLh���%2Jh򥤑3 �!�ċ1H����J�
4CF){r!�dF�E`ʐ ��C����BŚ=!�B75h��@�Gպ�($H�#h�!�Ę=)�d���z N̓s��!	�!�$1PĨ�0ek�\��qgA��!�dM�n�M���G�z�ڴf�RR!���f��D�vB<фM`�Õ��!�� T��/�N��4뛇HLP��"Ot1�4��C����g�p"�%�g"O��c�Ʃ�2(
6)B�S/h���"Oj���\4����H޳#�59"O�a�� �5RTҧӳ4>l��"O�(s�#Ĳ$6! u��$z�"O&,d�X8���Al��[KF�R�"Ob�%�pj"!��e"C# �@�"O.=��ϙ(Y.9�2�Ϊ9j� "O�B�-�a�Pr�n.<��"O��˄�����b��w3@��S"O���K�@m8=���.1h�9W"OѪ�.G��i�҈c�L�"O 0�%�C�D�Ԅ��-ɏ �f͐�"O�]@��-/��,����VG���G"O�A�O�/��E2���K4��`g"O\�'�m��|Q�%lxR��"O�\
6�(:��w�KZsTp "O\i���J�iĝ{�)q8�"p"Or8��B�+h*AC�
�q���"Of��
�Uڼ�C�	 �j�X�"O��
Q��8E�JmbG(�2+�(9�"O����]�S��}��E��)Е"ON� �ɭ) "M25��@\��x��'�mX�7kC�ey 	�:+�t���~�b�}e�!�S�Жx���Q���y�jé1��E�"��a��q
��yb��#l:<@6�V\b�2p���y� ^hD�91'�	x�.���y�铬?�m0`���#�&a0�"B�	"~lI���9���j�̷_Z�C��%Qx&�壎�иJP�UzB�	?F�J�eN�	�`1 �aN�V�LB�I8S* P���Q����3�Y�^�xB�
O�6�9%(�=)i81�F��
/LB�ɼh����!G�N�HY���p�B�I�*��t��`��-�ZM�S��$M�B�	�!���Ss�X�Nn\�RM�blB�5b�
��! *_Vd���6/�2B��$^!�����DFH�f��9�^C�ɐ��@�EK�h�<l�Q�:clPC�	�pr�A2=h�x9pV�B<{bC�I�?l*��ʝ�ِ���1Q"C䉤\"�����  ~�@9�0c�B� C�I;#�L@�A�@�h�����:�B�	�V"-x�&@&\�[t�Y�YJ(B䉮>������Aָx��'��C�	>t��PUg[� ���I��˰x�C�	�5p���b�l��k�B�xdC䉩r��L�Ԣ�Df���"��$�0C�	�W@�̑��8"芠"@
2hC䉉z���P��&+����Xo�u��ve�$��F!	+&�'�b0`���YS� �V*Y�]�BT�dDW:f�P�ȓe)���E�	&r�N�#�jO��0Ѕȓ,�L�� F���%���ް;!��ȓG�4h���T:���SM�2Ԇȓc
��*����L�6�8c@��������X�Bٓ$2��%Nב,u\��
6��RD�Ś���(��!�v��*i��r%���d���U�:y��Ĉ���ȿT��L���N�ޘԇ�T�$�s�3A���
�Y�^-�ȓV��`�7]�vГ�.�}����S�? t���:��:�h7|&jl"Of�
˂0�P�j5�Y�.�Ȣ�"O�} j�|�T���η�5""O1h4B��>��`��*�$�"OF���oL#:W�0�m^8S�İ�"O���s#H%c����Y4@�c�"O0$���ʙ��)V�~��"O6�e-8D�IbAx=0zG+�y�<Ѧ�OgiP�X�Jjδ�e-u�<Y��x�(��Ł(Y�,m�<с�r�v"�aN�pG���Ff�<��O�0�*q�5�.)�J�H`��I�<����_Z0���!��`���@�C�<��#1)�x�%�S�)G.�����}�<'i�H�
Ta���\k�%y���u�<����J<�cˋ�����n�<!�CŴEFl��,ɏ�l����<i�(��,���g����dȧ8��{�G�#B����
�AT���A�"!~&�!�i�8$f��?�k�	:`i�x#�IJ�X�l�
w��6?6�AU�hA�Q͚d��0{G`JY���'�3]T��6�U�y��-Pp��G�,�1��'X!���'�B6P��Y����g}��E���N����H�o���(O���D�+�:� �ƅ 0ܴ%��V��Ц���4��$W��SXy2N;=U�,K¢�R��4ۅ���^,��!JC�$/�y��'_�e�RL�?X�(qw��BpA�cҝ!�
�)S2"h���N9bYD~2��d����Ͳ��H���Š!p�@�g �+*F��B
�9>��S�a4Io^-Gy���2�?1ݴ��`��J+3�س`��d 
�m�����<���?AN>�'�MsC���5��Q�AH� Y�;X�<��G�t�DL�DK��Zd���۸|r�F3Ivv7�O�eo��:؊!�YwzB[��.�?'��S��ә����D-�W�qO���D�S�2�X+�@QG`>j�� �O�f�@�K;s�P�Y 6��ю��Ǭv�B��ҠN� ���̜!� ��'M��) ҡ�2
p��@�.gWB�FzBb�&�?��i��>-c��B�= P���8e���#*�����K�I�u�(YC�bQ���`F&���dFަA�4�M����2��0.0N�8t�
Sh���7u2�C�iR�'�哵!��	���n�/3����~8X �Rm4�V��C$�h/0$�煁&����O��y��S���Ovkl� ��E�+ڥ����A_�5 �6�Y-[A�ݺ��ϫ �J��	���� �Ki�����%E�ܴ+bi�Oǔ?�=�R�Wy���o�,~���_���X-O�O��s�Z�K����[�@�F�D4K��O����O��ĸ<E�$�W�!`���b�b�>�����(O�}l�'�MÏ����@@�ˏ�[v|��?�j{��ay2��y7�6M8,O��Ce ԟwȼ�H�s��1J�,F�g�]0��ו �|�kU:$������T���s�F��8hd�'��Otr���M	��M���<��Tz��
�mr`��O9�"<���N�lCT$f���x&�йn]�dA�"gi��<:���՟8�'�n��'�
/.�ʍ�@H�:V\���HO�A�Rg\�C�e(�B!CU��y�ګ�M%�i�'N���O�剥J�4a�R�Q�FGPܻ�Hh�*1�a\'e_����D�	ǟpu���	̟48sGR	s���CWC[�(���A7��3F�`�#AQ)(���ٱMC�`�'���;�
a�w���TI����AY� �a��2����W L#K��-E〫/����4��0 w��/��Ԕo�B�ܽKB %��jD�q����s��w�����r�X�Ķ<������Ծi`0���3ɶ�'��nr�K� ��I		�J���M�f�x��*�P�攈�>O�V�}��ۥ��dV�&��Z�    �   &   Ĵ���	��Z��t�D�8,���3��H��R�
O�ظ2�x�I[#����4Gf��BU>[,L+�l�(m��bZO�Hؙݴ���k�0���Iz��	����Y<4t��Q�&�҄X0l#�ox"<��~�^)Q�K�H]4� 1���>V��U�̳����cYX�F)?���>Y8H7M�X}�"/Y>��1q�ڧT���A�J���9g"[\y�f�O�dXb_��uW�??a (�6�����"�*td�3��dЬ��vd�*/3��
e��bٔTQN�4qA3ON"�i0�"a����Ehh�3��|r��|�'nN�$��趣��I���eNNоXw�s��tቊBl�S�g
E��y� Ƽ-�8mS�ŏ�OH�������$ �a�>�r�!_���Ls B��v�+)�"<1`�:�I�|NL�DBE��X�C��j��7��	�O�Î�Ğ������fQ��a5�-�"�t�K^#<Q&�6?铇�$A ���'+*�5X%�Mmy�M^S�'*�5�?ɓ�&�N���*��#7�x�2J�.CYN#<)b�4:E���לJ50q�&ڱ+̽�e�^�7�1O2����Z��Kр�K4؛Z�^d�W��z�dx�&� #<���'�Q�Vh���"9��,HPOΐ�q�IV��ޖ{���㤻iX��t�	tj��Ɵ./����t�ܱ�㞬9��Ʉ5��m�n�i'��*��<����]
q�'+f�Fx�js�'����GM:\�����h@��',~��@ ��0��Ia�<�#J�8'S��%���Sdi��+a�<��+�<���X��	�8$ir��^Y�<� �e����5)f ��.�{�6�Js"O��at��m�x8���]�(h��"O���� K�_#�=0��C? �b�"O�|�"U�p��(���{jp�@"O>��m9&$bE�2 �1Lf>�p�"Ou�*�/w@F�ʖ�Z>%x�"O��:�E!+lx[%��7�<��F"O�82��/i�����Z|�i�"O��jlӂz��У�MU Q(�"O~<iQg��n(<��֣����ps"O�Y+0� �#1&�P$��=����"Ox�קZ(_�܅cE�@g���"O������r��9 s�[<��A"O�Xg��}�D�#�\���"O��'-��T�Ţ�
S�R'|��b"O�	��iG�rH:��f�Q"Oܰ�ЊK�2�d����ƂG�8}Ä"O�s    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  ��     �  �  �  H*  �5  �@  SL  �W  �b  nk  �s  �|  R�  �  k�  ��  �  _�  ��  �  0�  {�  ��  #�  ��  (�  ��  ��  �  a�  >�  ��  � I = 
 �' �/ .7 o= �C �H  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H����<q�I�$3Oj���O�~��PeZ_�<�6�E�>�acfY�l�����S�'b�)ڧA~9��A86��%��(�0�b�ȓC��s䇜�`�f����|:��'%ў"|
�`8tڬ`��]cN&��e*�z�<��
�#b$�!��N�k��uO�ty��'t��X��K$3��" �M�pr�';�	��}
%�p��[v�<1�X� )�� ++�&��`�Nh�<1&L7p�5�1��J��E�jNg�<�φ�_TB9Q�� �Xl�q��͟�E{��I@�}��d����}��	#*	��B�I�}b�r��Q*-����4��7JH���p?1$�ҷ9�*�`��3����wDX�<�j��K9tH�Z<�n�6�W�<y��i��鲇*(DR��S�e�8�y�ᅾ��ـ�f�=��x8��Q&�y���1:Fp���KD��� %	��y"8�M:��@lbV�)d	Ӕ�y��[��Ը��M�g���CN��yb��1�
�"��[�<x�BI°�p?��O*p�M�>Jt:����VT��q"Oz(En9k��ˑe!�߰џG��G�v�c{V��``<H!�B�	;�}!t/��f�3��L�{q��hO>�  ui��r\`��!#�b6��C"OV�pA /�ڌ�@!�PTDru"O��fo��>�L@xRm�!;���"O2"�=_�h�l��_�,�C"O�Z�
�Su�	�U�, �lT1&�	T�����׾�C��
�Z� � 6ꍖi�!�$�,>�� �k��x�\\i�bA�
1O��=�|��ΙQFh�5�N�NcBгKZ�<q7�U���T���=�v%cs
�Z���0=ɳ�ܙh^���W��--�8�l\U�<e��nG̬�0kQ�-�R�����P�<�b�����sS��876�Fk]P�<�2#V?x9^�;�&�8r�ޝ�7G�N�<Y!�Ά;�2d�E$nR��A2N�<i#�Ŝp��+Ԇ��T���J�<�V�/��(�+i��,i�']|�<Q�@B�F����:��p�TKd�<��GE+�~ݹpI��q(���D�Ʀ�X�'(��(vbL�����߫KFh�9���'�y�@BQ�?#�����U�4��3�'k^8��AR����L�d��py��$=�S�T�����,$u+��C��y�@��5��p�IN�P����PyR��4S�a�.H�<�:JĢ�t�<em%d�ؘs��ϻ�<�S	m�<)]x�@VKh
FQp��=8�܅��Vy2..'.�ZC��/o �ADK�Y�<qç�8ւ�#��
�*�!�  �X�<��� ?(\x頡�^rUF4��)�n�<1�"�/N2�F��
\*�QÃ�E�'d�?A�l�>=/rY#0
�;�v�'A&D�PA�gL
0��9!�dP���h�<mZP�')ў �7�oض�� ?�-i�o<�O�0���wG�J�� 	���"yф@�'�}�
@	Y�ա4X<����4D���䒭
Qnms��\7}.����>D���sG�`�P@�i� f��a�;��-�Sܧ�v���βY\v`{w��&fH�������d�&㲈K�$��>��Q�D����A�h�a�ĸ1&D���n ��Is�ۛ~B�X"�
�6d�<����,bA�'B~�w
�5Pa�	��I]~���# ^��s%��4NA6%�y�%�\�>%�RS�>�,�������yB��yL�� �I��G����+Ƅ�y�J<JTmB#nSt�ui����y2��fq����- ] ��gd���y�̌0t�\��/X-�N�▧I��y҉��N�ִ��99�vH	7N��y��{�L ҪC�0`��vI��y�B�1!��i��Ҩ��yK�%��y2!Sd�����B�����y"�W*X�r ̀#J9��(ޤ�ybFZ��&I�u�ױ�Xi�C��"�y,H:}D iȖ�^+L��bꞦ�y�n�l� V�OF��M��(W��y��<CƑ��ڊO�&4+�m�y�N�Re�FO�*�uZ��E�y�R�k�J	7�ӟ"I��!ƫ�y��?~���y����i�� L,�y�a�*j�X��O�9��(��yB�)lb�#�MM0��B E��yBG˒|�BݢE��7��0�C��y�V�*D����b��@6O^��y
� ��J��E%��e�Z����e"OF)	#���=| �����ޭ�"O���2��8>����h�" 6"O�ȸ�.@ �@��R'4��D�"O����1Yu$u�T�	* �A�"O� (C����}X@%A�h��"O������%�����?M[�i��"Op$p���<#@����(T��3"O����&8x<�JY�,:V"O< ����Q^�*�(ߥEfD��A"OjP��.M�<�	�t']�Lja��"O�Y��ٴZ�D[�&ZZ1�i�"O���#��ai���%&�W}n�a�"O�Q��C��JErUJ¥ݦCw虻�'��3TjCT.�i)�!�82����'����dJû}�t��G"[]eH�'٢�� �4dv��d��]��'�r�p�\�FhQ���M82i��'��!���'t/4=@2��
3�A:
�'nt��5#��Z�p��q�2�F�
�'a�툦�ޔ6���`rg��%-2�	�'����Em
�O!tQ�1��*$�|��'�D���O�p���4����'��Q���!�X@��gQ�0,By��'�z�3��]�S��a�Dh�2���
�'JҀ��i�.� �ĥ�=S��tk�'R��� d�2����4L	MZv��'�r����$d`Њ�o�C:�ٙ�'�̡�H��r�D7�90�촡�'@>`*  �*�E���])t��'� ]����*Π�`,A�ilvQ!�'�l��`�
��*@�'�x��'��d�SjȑM1| �����4����'@][�L�$�\���1VDPM��'�ٱ�b̶u��6h��F��%A�"OT�"��@ʰu���å�n�Pd"O�LZ�+�~UJ�#0�U�1��i*0"O���gF�q��@��Aɀ+�����"OB�9TG[6[�@�Wc�ks����"Om�7�rQ��X�"C.p�̼��"O�`QlV�eST�R<��I�3"Oh���E֒l7,9�����5���"O���vJ��T�"�n{o(��"O
U{�DRVn�%``��R)��"O\@I�e�^Cr��U� =l��"O �9�HT�kVRA�f��R����$"On�V�B����	J&_����c"O��x�KE�AxPHD��xX�"OEjC��"h��ٓG(H-5��1�"OdIy����\f&,s�	6�,��r"OH3���@I����ʙfL#�"O�<��Q('�T�	���"4���S"Otݛ!MS�R{>6ブ1?.d���#D��a5�V�]��XbԀĒu��:V->D��aS�R��: �@�p�5��	=D�(�C��V�(M�t���t>v��?D�l���l8n����-L�\��=D�AL�!=�Pi���f,���N<D�lەaAx+�y�D;m0�x9E�8D�`��=�����$�}��h�$D��c>[�:���`F�L�*O*ѹE5ZF���TE6R���"O��K��(�@�D	E�<;W"O����l�l8<�ѣ"O� ����Ꙭ	�<���B����"O0u��M�&_�ta+ 퇣L���rv"Oz�a&'��daH�j�E�f~�qs"O:�ă�-�p�a'�xR��rp"Of����ݕ}�Ɣ:'�Y�V�:���'���'{��'w2�'�B�'���'�`�:�b�t�h�&��C�U��'FR�'s��'R�'���'���'>XE�P�O�F�
�9��w�=r��'nR�'�B�'z��'���';r�'>�H�!:����P.�2d�>���'���'���'l��'�2�'��'��=�@!�J�Yh���h?j� ��'p�''R�'��'���'(��'}I��rDc�n^�C1��C��'(R�'���'���'B�'*�'Pά��MB�g��:@˃�"}�0�'���'��'���'��'8b�'���Q/09҂��4��Ȳ��'z"�'���'���'9��'�b�'tN8�@�1����o�tx��2�'EB�'��'��'o��'r��'Kr����I�l,ȓU��RE�'�r�'�r�'�R�'���'��'�	qW	"F�#vL�o���X��'*��'��'��'3�'�b�'$,�h6Έ;'�R�� IJ�^�N��s�'���'�R�'p��'�B�'���'��Q�u*�;!<�J��&�D���'���'���'Y��'��as�V���O4@ 6�@+԰�[�BD}<��_-"��?�*O1���
�M��	t�œ'� 5W�0�߀I\�e�'��6�<�i>����\�� ;l������C�A�Qc���՟����#���n�]~R?�:���C�)�:;�p�(��=2D�VᏻP1O0�į<ɉ�I�j�����N3d�}0G�ҁ���l�\��c���5��yw��CN�wa
++����(D�W2�'�>�|R��A?�MK�'��-���K3�^�raIF
XN�M�'���蟠���i>��I/8+>�eN��Pܘt�ğ�~����<�H>��iJ�$j�yB*R�F����Ł��|����L��On��'���'��d�>���R~�X[s䒇QNlaxpCX~r�'��`�����O��d��v�@�+N6JI��DSp�(`b�4X ��Kyr򧈟�D��@]�|�F�62��u�I���������c4?!d�iw�O�ƬqRFɸ ��	y�R�B/�9e��d�OX���ODQ�keӼ���Dn���ט�*�E��CSu��"��B�|�D�O����O�)�O����OL��O,\!�&D	�P����J&\&T	����OR�$M�R��K���OH���O�tlZ 3G���ß 0R��*� ai4L�T�����ڣ\���	Ο@�	���S_���'��H:Bq��q�i��e�����c�^5i�O��$�!Pǂ�J��7"<�O��U�h	a�Z�#�Ʃ
�j�}������?����?�� �*��(O�n�h�b��S�(��3���+
� ����Ɍ)�PM�I.�MC���D�O��'�2_���R#ӕh��X U�̓n� �H��/dW�l��<�����J��JY�*O:�	��z=��E�@���x"`%9��p�9O��D�O��O ��O��?�Q��t )�4Gڊ6�h��m������џXڴmu|�ͧ�?᳸i�'3��Z��H�&<*��(�r0���|��'��O��w�iI��8��}'���b� ���[;Obb$���	�q�r�JB�	Dy�O���'�!��L��R&�^|��C���K��'3��M�  ���?���?+�>P ��sĊ�2Ĥ��k�B�ʅ1OJ�DLl}�'_r�|ʟf�)�M%�^�蒬�"q8\�@֚B)Z�ҍuӊ�����T?aL>�Ī��'�
�K���q�`m!�IN��?9���?���?�|�.ONn�&3ȭ���&�<XNU,خ��G��˟ �I��Mc�2`�>�,9���C���+���x���6pX���?�1����M#�O�abc.���V�� 3�	k�|�pIٜ�8���{���'r�{��^�N)�0�6���V���*H�h��7-�U�L���O�d7��-�Mϻ$v�l����$������L�B�և�?����S�'2��۴�y�G��N\0q���3Zt*s���yҥW�	�������O���Z6U"�A3iP�ro*��eǲgn&���O��$�O�ʓOK�V�W/7#��'�I�o����R�H�B�62�O,��'���'��'��|��E��d�#�/W@ъ�O���Ed�+Ft���󉖫�?���O�)�vM��Wμ��U�p5�H3��O���O���O\�}
��LY�1p�Kѩ�\5i�̐4�dm���i����3&��'��6�:�i����<`l~9��+Wkr���h`����ß����{�2LmJ~r�՗\tp-��.R�,傕�ԩK�T��Aa Tm�%���|Q���������I��8���W�p#��gCˈ|N%���py�`z�6� aj�<�����O*�5xŮ�i�
�!#��y �2��>���?�H>�|��D�	gy	B�;&� �_�^��q�t~@�D��m�� i@�'�����$A� !Mآ�Oя�����'2�'���'��P�l3ݴ��;��dR���-b�  ���B(�S��r����|��'����?1,O�!Y��Z��������!n�P��`�Q��7�d���##�]S��OV��'������ ,�s��R}��U+L���h�5O*���O@���O����<�O}ĸ��-&Ɛ�	�&L,K ��ڙ'�R�'c"�{�:�"�İ<�i�Q��+"�Z�|��dN��^'�bf"�ߟ��������Ŧ�͓�?qW��%G2�qd���4o�y;2/Ȳ��;Q��O"�I>1)OB�$�O���O MXS��ݴ,¬T�m�N�J�M�O���<� �i�|��0�'��'$�Sz�,YSg�Hk�f�	5M\�e��=��IßD��w�)�P"]�wQV�
������ h�0%�E�"�G7�Mc�O��ʠ�~�|R�Б@�f�s��QRTx���]�,^��'s��'k���T��Qݴ0����,�FV�p-��J�j4��(�?!�Û���u}��'���D3q.��-W�!��T�t8�
�����'@��󱧒�?�pZ� Xp�׷6>��)�9!�L���jp�h�'�"�'K��''R�'{�S �8!ӑA�(w;��zE��"eT��a�4 3�,��?9�����<���y��E5ؾ�k��Dqj�jd�\���'�ɧ�O&����i4�O�!���!/!T�B��W+XP�d\2�bj�a||�Oj��|B��R�|pt�JH��X���O�Fa�����?���?�.O@-m�&s������t�	 Im�C�JC�4��egO��[�0&�H�I�����O��2�U�%���4%��3㌜ф�S(��	*'�9p�IǦ�O~�������	�' y���B+Jʹ(`1YI����՟���ٟ\�I{�O�"�B�G������ c����(ne��	s��O��������?�;;>�{�)�؝2��Y�z=͓�?���?�'���M��O�e��W��2�� 3��3%a;N*���o� 1�O(��|���?Y��?�ܦA+  !2H����9E����3�Qgy��k��%$�O2���O
��6�dגX\��#l�2�p�Rc@	D}�';��'ɧ�Oi�ԉ��2-�n=�&���t���a�m��f���:��	5U��5���<q��	L����BH�6q�ܠ3E�?�?A���?!��?ͧ��ğ���g�_� ;�K��e��%�#�Y�,�@pK�+���޴��'����?���?ٴ L7=]t�8��@�3�x��`�3:,(�Zڴ���׃N�()��)���,ӥ�!�,܊��]�
�
��>O����O����O���Or��@�(RgڭO!D�0EA�p�`���͛ή˓�?Y��iO*0y�O#��'��T��c���/3n�z]�ffY�v0��?���?���=�ܙ�4�y�'�ظ�uI�K�����e��2��y@��D�@e��/�'��	ş���֟���"9�@Q�l�j��vf^�*���۟�'��6���6M����OV�$�|Z��@�a�����&K�. RHX|~��>���?YN>�O�z�R��߃IWZ�y NN�sZ$RǪW'u4*rE�i��i>�� �OƓO�<�p�э;Od��wgۓ;r����O����O��O1���4#��#X�j�4!b�;Ɯň�o$o�ա&Y����4��'ʜ듇?�2D�>Q��eCG��0�h �����?1�%߼��4�����H��U�'��S�X(%k�HK�UÐ�:3�pb�	sy"�'��'���'�V>�[Fi�5i��	�l/V�I+�Ȓ��M�7&Ɨ�?���?O~�r1��w��XcY���L�a[7�����'b�|��4iܒ(2�61O�q�d�B����õQG��q�9O����˃��?Iu�,���<ͧ�?q�(N!A�,�2�/x'�l�­ɥ�?����?�����DDۦ]�D����	�d�K��
�A-��W��l��d��v���蟘�?�d�� m����C�.���˰��f~�#)�����b"��O����I#�2I
H4���Ќ�-ܑ�����b�'���'K�s�1	�
%�	����gDX@;E�RП��4}�����?YS�iF�'��w���-� Z� �R�C�Ϟ�C�'qb�'=R͔N��F���]ۚ������
�!�:D��H�`�$�	kc�|�P���Iџ��	՟L��������)H���G��N9"�CLPy�/�N�`f��O���O��?�a'りC�y��E�,3i�H��jJ����O��D3���U�R88�R�ΫMq�`���Fq�ኄ�()����(��'[R�%�0�'oʅ����$n>�:-2���k��'E�'�2����P��jڴqN��Z��|�����B����`D�:0� ��Q8����K}2�'���'?~��Q�D���޴d��(9�gP�y�b��޴����l�V�j��6��v�.���`���¶���+�߯vl���Ob�$�O��d�O���+�S�V�2��ǒ!XUJg�`�'t��pӈ���?9Q�4��O=�@ʑdPerON�!����L>q���?ͧc��� ޴���S�1k���!{MvE�7[�e��g�S��~"�|�Y��������	���g֟	��P#�eJ�µ���J����I{yrik�bUZ!��O��d�ON�'��C@h�7c��1���K<�@��'�&��?����S�d�͉}.,z�Q6�
�����L��$���ɫM����S�'��$7��ə/�H��F��*q�莾�����O��D�OH��)�<���iH�-!�r�](�n��D9�Ly��>@��'�6M'�$�O�m�'P���Jh�M�I��`8�ᆬrN��'ޒ�	1�ik�i�%�BJ�?I8U�� ���W��8���U�8m�}��6O6ʓ�?���?!��?q���iT<zI�p4!�5�z�` U�]e2uo�-J�$�����i�s�|J���"���N�[�N�� (U�.��0,�O��d$��i[Z��7�i�3G&�>l���n�`��iyc�0�Ã >-��+�V�yʟ����]���!AW�'�tM��'>6�υ|��O��D�)yJ� ���]n�E ������ ��O����O��O��(a�^6�\ȓÈ;<O �`��0�0"�����A�j��
�2A�����2��3��Ń���&1A��"D(Xȟ8���|�	���D��'{r�۷�^���l�sk^�,L���u�'p�7G�azj˓&-��4�E#FA�<z�0����'Y=N�k@:O����O����=��73?��I\�����-�8�6 �/D��3��z����J>!/O�)�O^���O���Oye'+5�ԝXf���Of�i� �<���i���d�'���'��t#�L�2�' �Tk�,�#�^`����P�P8#�A�>��������'����<7�2��A�49�PA��TIv�$��*�Y�	�SC$�y��'-j@$��'D���#�ȏ4w�L3�.B/2^�1�2�'��'����$Y���ٴ �\t9��)0�=�b�
H�ҁ��_=�ДΓr4�F�dH}��'h��'�����>��	q���s����5�~ϛF�� �RAV6D�������qȀ�E*������6�ʬ�":O^��O��D�OF��O8�?`�*��YR�M�u�K~��$�O4������RAy�c�j�O A!B㇖Z�0P��7�~5��3���O~�4��t�4 a�F�HP�Ј��.D�|h1��o������N\ ���������9O�m�oŖ`cR��D�X�:�ة���5�M���T��?Y��?Y/��}
A�֐��H���'
�+c��,1�O����On�O�S�f�%�B΍�(vq��勎tf�h֋�U�f�) �uy�O P}�	���'�����N�1��0(�"A��`ԁ�'��'db���O0�I,�M�G&�?�$pp��(wdD������#t����?��i��Oʑ�'���MO<���%/V�GF��; �k�I�E]�o�j~ң�%X�fQ�S�H�IY���2n\.<��!��m�"��IOy��'�"�'b�'|�]>52���h��Ma�)�0���F�-�M������?���?aL~�cᛞw�8�R�N�1�Խ"�/ǺAj���e�'B�|���*�m/�3On���g��W�̍�M�&���E:O�9��ʞ��?a��8�D�<�'�?�Yw�Pdq��R;sT���� �?)��?i�������iB��h�	�@/,fM��/��l���S���
h�?�"P�L��ޟ�'���r����%�hv����5_f�	"h��,��b�ۦ�SK~�ᥟ��I�SDA����a��@�IFC�����ʟ���ڟ��`�O��gΦ>�aʱ��b��cD�1p�~Ӗ�A`�O��D�٦)�?ͻy���q�(x~ݻ��R$�P��?����?a�k�M��O|b�MU��
w�A%O����ܫ;��T��@��O��|b��?���?���Eu���p�.5JX�d�ݭK���3.O��mZ?�lQ�I�D��[�s��D�".CH%�O�Fj�#����d�Oz��>��>'!Q�FC?/���I6d�h!��0��I�l�D5��'j�m$�,�'�N�"5�\&R �X�RkC��E���'�B�'�����tY�l�ߴRB\����F�95i�-thd=�g�Mj�����F����|B�'�&��?���?	�a�>���z���+B>���R�,&��ݴ��$O f��y���o�N����!S@��ѱjI/��!`D�d����O���Oj���O���#��R���+�)on�Ha&yF@��	�� �	�M�2$L�|���1ʛ��|Zڤ9`@��[�.Q��j�#K���K>����?ͧ2�V���4��DO I��"lM�x�R�8E�<u�|	!�
�+�~�|�\���Iӟ�I��|�C�`!L,X�T�6����U��"�
���-�Mylr�hdʲ���h���O��)��6a80 �V;�b��Ȭ���x�5O@�dMc}b�'{�O�I�O:��i�
<(Hf �5rw�x;�E��-�%���c��ʓ�Z���O�)
H>�
��w��9��C�(h@2#ό��?1���?����?ͧ�?����$���;�!��h5�$Ӣ)bZi�-DGF@ ���l����Д'��Z����;��XH���N=����h�t�x(��ϟ� c�[Ϧ]��?���0E�p���f~��2Y�I�7(Ɲ=�u3G��,�y�Q�H��	`aB�4~}��zo�#����4@0���?A����OR�6=��A�)M�1��Z�x�b}c���O�d0��	����7M|�h20��^�t�[�Kf~I��Em���J:uj�d+�D�<���?�cOS�����7nS=�v���?I��?������d���!����?���ԟ�rt�D�ɢ�@�\��9zY��&���	(����Od�d�#��S��IVdY�w T� tx���ɒds��zp�Z@2�D�'J������`��' m�#lvt������]<���1�'�"�'[��'Q�>��%��,�ǁ��G-sf�I�AX��I�M�
�"�?���e_��|R��y��(/s���o։;)t�B#.�y2�'p��'' ����i���
�����۟� �K�N^�3%����F�
�~43�3���<���?���?����?y��;ƞ4{�,J6w\ ��ל����q�!Ɵ �Iϟ�&?-�I7S �x@	U�B4@��V�6Ҭ��Ox���OޓO1��q�?�`4�K�J�=��c�=i,��q�<��E�z���Ɖ�����Q�ֶ�bp�U`6`��@Ig^�d�O��D�O6�4��� ��v�D3��l�9H����i�szʍ"�b��#�b�b�>㟀�O4��<Y��-#��2'�� r�ie��#��޴����Y4B�A�'}�\��Z���6�@�&h�!6���c��]}�d�O��D�O ��O0��>��\�N��͕�2צA���D���X�'#�n�¨��?a��4��C�dYY���3,ƩB��C&Ka����(�i>�1�LΦ��u�΂ sd��Ó�<�f�6�L"7�'��%�X�'DB�'��'�t��d�^�*!����q�x䘡�'BV����4!3�l���?�������C���ku�+([��8��C7�I0����OL�d>��?�uIS�y�6|kRm���,���nE�_�4A�0 �&�^��|2t��O��ZH>��F5!�|��5�A�a�,���j���?Q��?����?ͧ�?Y�����Ϧ�QJ�	�"a�$̝�	�#6(Æ���֟hq�4���?��R�`��8&�PŢ��SFU0华vqz�I˟x�"�XЦ�ϓ�?�JCF3��i��dӢeE�ر"˓=�D�A�9�d�<)���?���?���?*��h"���L�|�� �"�����ɏ�1x�*��X����<%?�	9�MϻnF�+a�^
g�
���%O�m����?aN>�|���Q��M��'�h}s��eŚ�	0NU�,i��'n`�[6�؟�B�|]��I�����E�!!�숏mt�4h����>4p�&�_yr�mӀ�Ce$������O:��7@E� ��d��cƅJ%�4�2�D�O��'����>䥸JԪV/"�iG��n����O ����ޕ�T)���<���~U8����?y�A�?o�(@ՄE�.8~EF�۠�?y��?a���?�L~�u���?q���3aEV�I���a�BТ,���z�F�Tb�'�|��y7�k4F���%M5fӠ `T%l8B�'�"�'����F�iZ���O�A�7��(H�k,��Mdⴁ�N�>��-s��ÿGg��N>A+O���Oh��O��d�Ob(�R��EE~�dL׭F
��2Bm�<)d�i�F�Z�]���Im�ޟ����[1"����֫Z��}�6.C�����O���3��)Q<u�8ѱ#�K�$b�� �X�g����>�*ʓc1*1��O��J>+Oh� %K���90$��DJ8� �O���O���O�<��i��H �'jDP#�Q'�ܩ�S��,YI��'/67�;�I�����O2����� �I<(�s��$gh�I�J߆�M��O��������k;�	��N̈T�XVx �2�̑
���1�7O��D�O����O4���Oz�?�k�b�c���Q.P�h��tB���d��͟��ߴB�F��O\6�<�d�D��qf�,K���� �TҒO8�$�O���#S�7�8?Q-��18H�@j�JAT%��<I� ����t'��'���'��'hp�prn_?@��DiN��l-�yX��'�BY�\ ޴�<���?a����${#\p
��}�|�I3^*������O���4��?Y����Og6<�Ġ�+u~�����5iؐ)���J"��|2���ODzM>Ia�z]�xA��)^��kV�L0�?����?Q��?�|z-O&�l5+�lE�0o�#�=J@��|��Q�c�TyR�cӄ�J�Oh�$4Զ4�/^w$�X��̩u���d�O�p��yӎ�)Mų���B�O_蹢�L9��4
����'���q�'�I����	ğ����P��a��iˁ=F�*eK7.x������F��6L�K�f���O��$3���O��lz�����Z���h�F�>|��(��M�����K�)擆��im��<�&N�"
�n��lZ�v��E�ckB�<���^.I̮�IL�	eyS�� $�0�lI� �mB�j.'O�4m�
G:R8�����ɮhr<[ #�+����$�� �4��?��Q�<��˟�&���t�Z"E(>T�rBNWR41�7?�����HD�a���'
�F����?q#Ǌ�4(��A�@c��#��G��?����?���?9����O��RR�×4��$���ęe�6�+���OL��ɞXMF�D�O��n�I�Ӽ�l	�Z�u���U�PP*BO��<���?A��Q0�l��4��$�=4��Գ�O-���I�s�>1��)@�b��B�|�U����ΟP�	џ���ߟ�À R*R�b��6� p�O	Sy�	l�t���O����OB���G=	)�{T�K ��p��Z�:-��'���'�ɧ�O� T+�F���a�p��:߮�A��R����O�]Y�b�%�?�76���<�@��R�fR4H��su�A"`Ir�����Ř��ş,�b��c%
sd��*k�����Ut��4��'��듕?A�ӼK�l�5X�P�F	34��)�r�ªtͶT3�4���ʕ'�z4���T:��^�NK�@\�a��&d:d� '��$�OZ���O����O~��.��'+N����
?y�.be��n m��ߟ���.�M�T�K�|��e曖�|�O�(�yz��
?�"}s�k]�F��')����dGK5C��&���]�� �Fo�-L"�3f��
L�I�IB��?��;�d�<����?a���?���"��{c�ڻL[�M8Ԍ���?���W����(؟�����O�*��3������#�OP��'�r�'Cɧ�I��q�5� �O�000�3�ځ������|�>6�1?�';f��IF�>�t�"�!A� =�k�F������I����	��)��wy�.j��a�i��������N>6�X��cn�:��˓'��$O~}2�'�Td��!M��G�Kk )w�'J�W/d���� !�kH�~ �$�~"CB�� ��@UF�/$`�z�$D�<9(O��d�OB�d�O����O�˧a,d�����?W��%hAeߞ0)6%��i^���Z����s��˟\����� _�u_�<�r���nI2��.�?Y����S�'?���2ٴ�y2�<�����/U2��6��aHhjB����$�,�'$�	 	��T� d�=/,���I������Φ=Y������I�`��nP�}d���`��U.D��c�G��m�I�X�	H�;Ĕp�K͗}k % ��'SF��.�b Z6�ʸw����N~����'J�~< ���Μ8�ϊ$+`�&il���0�גs��1����L])$��'T}��fz5����&e;ҙ�k�k#�|30���.�d�Kv�L�CDa{؞��᎒(y�&L)� (;b��@.k	�iY���S�I�s�C�к QW#��?^�A��ǚ4��,!�	� ��5D��N�{����c�@���B ,��*��ۖ�΂>���j#��8a�ܿg��\��a�T�P�����(t^-ҵ�d��ۇB�m��	c�g�yU�m�����_���$�<Y����;!���eɌ�C�'jV�LQv&�V}���X��'���'�W��g[2[w&p`cD�#M��J'JB+���O��?I>����?�d�j@P��q�ǚO�3G�@)!n��<���?������P1/�TY�'x)��d*����A#�DV/Lw�}mqyr�'��'xb�'�FU)�O`�yWE��:�Ud��?:+�kQ}��'H�'B�I��������]:^��{0��#o����s��&'�BTo�՟�%����՟I��Uܓ*ZI��B�)��x2d!ӥЄ}m�ԟ���Vy"�Ƀ-��'�?���rA�.yhN��F^�n�Ld�M�6c6�'���'Rv�1��'��'����/z�45q&�9!+���K)k�V_�H�!���M���?y����\��X�N:L�:��&6Icr�[#Ua6m�O��d�5F�(�}B���*��dK�.݇�f�ben������@�!�M3���?��z�]�Ȕ'�\a����B�<�(U��0qt�#�y�n�!���O��Ox�?��	��ĩ;CG�b��%s��$�����4�?a��?����[��IJyR�'����brp�YR�_FM~����h��O�E!:���OH�$�O��)�d-Jz: �ǥ\	F�:v�צI�I�L���0�O���?qH>�1Q�"f猆|�B܂�ć�]���' ��y�'*r�'?�I�K"D�Y�$<����@N;C8ݓ�g�/��$�<�����?��U������	��|�����X�dN���䓁?���?a)O�P��O�|����{��؋��G�I)6h�@I���'���|��'����m�$#�$l
E-�?��5�VӞ+��I�L����X�'��-�`I�~����p��c�YFm0i�5(�|���iY�D��؟x�	�a?����dH[�+��\�*�T���ϟG����'BU�*!����'�?q��c��!<�Li�B�Kj��2���ͦy�'���'L2�'J��yZcŸ��ȋr}L����@p ٴ��D='�}l�����O��iG~2	I�8)�ⅻ8DJ��)�M+���?a���?Q$_?5�'��s���2/O�v(@�T�8<-K�i�R� ��'5��'c��O,�)�2���T��A���>H�����@�>d��	b"<E��I��X���o��|"�'��Y��7��O��E����,O��r�$�<N��=K���=�� ӑ��6(1Dx2�:�ݟ��j��Ub<Ҫ�S�)�k��umZ؟�R�euy���~�RGȨ4h2Q�u�C/PKD�x�޽JvOhu�$�O��?5,��DF<\a�B�W�,���H�:�@,Oj���O��t�	t?	�G�!o��I��n,W��`pA�ܦ5�B*���'�2K��:���O4b�Hd3b'^R��(� �����'ER���O�˓y�l�= ��a��Q�p*��#R v�O����<a��s���+���dP9;���v
s�ڀ�Ǻ@�Pao�r���?Q.O��!w�xbD��ZNYCCL'k{��a�0oZӟX�Igy�%ȑU�D�����k��(� ��,ǩn��#lz�'�������	G�s���
8��m���M�ᒶ%�)HT6��?i���4�?����?i���*+O�O"O�T|*�\.��Q`(�-����'$�I�<Ɛ"<%>!`�AЦ+o���Vv��i`�t�,<�d��ᦝ��ş����?� L<�'���cI�wc��i%�%k^Bq��is2�'�r�|ʟ�$�O�����"�n�c�ۧ`=���G/Pߦ}���t�I����K<ͧ�?Q�'��,y�MW	4�P%{����4�?�H>yU?��͟t����(y���Sd�� ���������o����I��7���|B����z�� ,*&L��Z�!"��oN|s��x��'������Ο̗'͞�v-Ÿ&RM�B,�NOH�$d];`?TO��D�Ox�O��Ӻ �?+����Ǆrh���������I[�����'=�̗�T���E
+�([�o\�}��}ðO���&�';��D�Ov˓r�Yo d���e��{�G�cV���?Q��?�*O�A��,�b�ӱ��h0�MƖ �V�x�]81)�4�?�J>i*O�i�O��Ox��#�×06A`Sᑝ�a��4�?�����$N���Or�'���;~L��ʚ(Zz�;��R)����?����?�"`��<aM>��O�L)ś�ZRB�Z���E�F��ߴ��D=n�T!nZ�$������������a��ς�Hܜ�4�1g�h2�i��'"89�'K2[�l�}��ðZ�X�0d,!6�,��d�ʦ�0$l��6���I�H���?�#�O,�Âi6�
 U&lht�N Jp[E�ii�[�'�T����L���Cӣ�^P�%��J�6����u�i]B�'��� sF�����O��	�< 1ȴ쉏D��z���X��6��O�˓L��S���'YbޟN�0HA�NwxMzdf&� �KӸi�O�2Iw�����O�ʓ�?�11����
�r��LI�����'�!�'I��'2B�'�T�l�'l��O���PE�\6b�Y���h�d(�O�ʓ�?�,O���O�dS.hV�1�ElD�7m� ��)�j�xQ�5OV��?���?Q)Ob�t�U�|
���8�4Hpƛ�F�:	3�!HҦU�'��X�P�����ɁX��	�+�~�{T�-'~��p�[�) �ۮO���OX���<1��/'�S���{��V���؞�%p2g�%�M[����O.�D�Oȭj�;O��Y�1�,mX�����$+$I�E�d���$�O�ʓ.z��X�]?���ʟ���4ly��Yw%��{�lM��`��?�p���O6�D�O���A�4��D�|�����4O�FDB����3~'����㗡�M�,O�傂�ܦ������I�?Y��O�΅F&(�$N!Il�`�o�I��^�F�'cX�Ø'� ��<���4�߿"^�X���G�yݜ�͐&�M��A�m�V�'w��'��$b�>�+O�1�HO
���E��_�X�@C�Ӧ%s��t�$��Py��i�O����b�x��p5�X5tH��a�Uͦy�	��I�;h�U��O��?1�'߂�����5�h1����8J� @�4�?���?QB,��<�O���'6,/���-�?��i�׬�RN$6��OZ�Q�GBy}bT�0�I@yr��5�"[���D���2~��������M���6	���?A���?����?�+O
��#M��4�נO�Z�ͫ#Y�g1"��'v�I��'w��'��ک%�ViX��W#��NH<`�P��'E"�'���'�BT���P*���ĨU9Q��ڲ޼9�p��@�2�Mk*O$��<a��?���x�O�H8�6J	}���g�׎��ayݴ�?��?A�����/Ky���ORZci�1��*�=t~đ* �<nm�ܴ�?)/O��D�O������	v?��n�!`��	�GF,U|�C���������̔'���z7��~����?���U������8��S�Ν�G��d�vX������8�	C`@�g~2ݟ��{�ʡ;P�(<DL�i��Ib&��ٴ�?)��?���<�i�q�g�)�(�H���O�$�p�fr�n���Ox5�;O�L��y���K�o9���Sp�m�j�4|ӛfό�`Ԛ7-�Ox�$�O���s}B[���A$׽��e��,A�b�.9���2�M��.Q�<����>�S�����Q�#;��"TA�)�0B���M����?���{`P��[�Ԗ'�r�O$8���ВWǴӧ�]�FGj�r�i��Z�\��+i���?9��?�����|�ĆФM����C�Q�
,�F�'�^u�4�:�	���%��(Xz�����V�)Tk��5`<�iD�̓����O��D$�I�$).�ՙu蘪���6�7#eȰ[�b�]쓂?H>���?��N�U��u�H��WX��B� ;d�\5����O���?�	ƫ,�@��'<���;�cK��L��y�0��O��O����O��b=O��S5�i�ql������H}R�'"�'��	 x�-�I|ZGd�P�<�P�%R�wt0zAi���'��'�'P���')�Y
�{�h��I��h���C��oǟ��ITy"�������D��*̣�'��5R�H7oրx..}��Ty��X�I�v*�k��iJ5�M>��m�MшR(��t!�𦱕',�0K��Ӕ�O���OR���<\��J�	ՄAȆF2閝n�ǟ���}�`�Is��pܧ�`0ŝ"o�l�C�(B�{�8n��&e��H�4�?���?Q�'o��OݘC��ns2��ü1�"��f��Q�Ս�`$������"dy� �_�q#1.��4�x�!%�i*��' �JP�4\�OJ��O��I��
�Zb���������f7-;��A�'��&>M�Iϟ���BSpI�QE�+R �=��-�k���ܴ�?�t��[Q�O���4�����7��2�Aq�4��Ѱ�W��c@�ʟh�'�r�'n�Q��s��0�h�R���f6�Z�][�K<��?�N>���?��AU�@�`�H�D�i�
�*��p�p̓����OR�$�O�˓J�H ;�(+���k{$��ҒN�:��Q�x��'��'���'Y��9��'��� �Ui�H�##͊<����!آ���T���ǟ���gyb�Og��ҷt,R�$�42倔-��r���ʦ��I\��˟����<�0�W�D��o�F\�Cc��GP��j@� ��&�'Q�X��11cߍ�ħ�?���C���\�A����!�3d�a����O.��?a��P�I Z�A�R��)�@��?ɀ�F�?A����$��$�?��T!S7�"|`Ή�U"z�� �d�(���<�&�y��ħYf4��򩘿q�:���#�A24lZ�m=<��ߴ�?���?���d��'I�m��Lj�Y�7���E�9���$�Oh�y`�T`ԩ�W��j[�`R��T�������4�	�|I�x�N<y���?q�'�����]2;gP��o�r�&���?)��?i� 7-,,���'���Z=����'=�{r�#�d�O���4����@�@�D�Gp��@�T˼�RT�$�6�?�˟P��ş��'�~J�dG�
�fP�A���z�)χ(4�pO.��O@�O,�$�O�l�'��.�x�B���9 H>e8@!XM/1O��d�O����O>��-1����.&��@�5Sg��ya�C�|L@LlZYyR�'�'4B[�|c7Kb�%!e��q:9��}]%�2l{}��'��'"�.K���I|e���x�4`rC+��q4,W��9��'}"�����*�ѓ��M&:LR�L��Y�����i>�'"�'�����'��P�@������I`��b!�\e�r����M<�������4���]�\����o<ɢ"�\M�>7��<�V�Rv��~�����`��xy��5vJ�$�VLM.pJ��։wӘ�d�Oh��q�'m�����%V�? Ry���-��n�$P�l��4�?����?���q�'��aG;m/��Z�@ߒ\(�5z1���$r87�Zp�"|���5�D�Ĩ�)=0$��*�":*�S�i���'��*��Y�lc�0��b?�A�U�8����]�e�ܽ�Əf�]�d��<y��?���WA�i���ˏ$N�!2�)ߧ�,�#�i����D>8c� �IK�i��9Bo\	Q��j��L�𬂄Ȣ>Q�]̓�?����$�Oh����G*m��C��P!S&��I4�҃)�Xʓ�?���?�I>����~BĜ�d����L?�m0s��<�M�eKD~b�'���'��ɒ�i؞O�&�@��mjT���݉(�:m�Ob�D�On�O`�d9�� aH�h��^�e"8|�wۏL�H��?���?�,O��ѤL�G��$���ȓ���]�w�;j�z��ݴ�?�J>9��?i�!�|�kf��雝t�D9J��T�Z�oZ�(��hy�!M�3<V��������BGl�2�����I��Ir-v�	�����'�"<Q�O��,��.,���1�*P�5��	 �y��\C�F�F�����'(.xA�OdiY�cA�t��3�e,jz�"O,�j� M�6����rI\���*0�⣩O=g����W%�0@�b�bI-$��$���faJ�c���$,9��:C���vU�͋S���(y�PQ��G�	0���ҹ2�R)hR�	?�V����ˇZZm���Ϻ��FJ��V �Q�B�*���h��4^�Uzt��,45��u4������G��?1��?��4����O���0�`ͬ�@i��P��-[�L�l�`���Q�"���hc��넝9@�9����&��2{�ȳΖ�xȣȍ�j;�hc���������XD��$�d��0	Z��@eR���>;�`�	�a�^���O��=I.O�hV*Ϛf����a�&m0�Qp�"OV���@��h��z��T&\�� �ZV���ɿ<AF�@�4'��d;
��`T�M2xX���'[8C��'F��'1�U���'�b�'YX ��<NB��9�f�)��� >X�D;w#�+�p>!�+��D�N����y2��R� ��X�!���Xń�I������O^ ��ɝ+p�� e�Y� 2�a�+�$�O>��)�$:��Ͷ!rpt�A!��6�yթ$_�!�N`��Ĉ!k
�)�H�VI� U��d���IXyb��KR�ꓽ?�)�Q8�:1od��/��X���*a�G_a��D�O����:%��x�d�#!'�)���G��';��$���H�l_��Q��@4Y�&HGyҊ���t����L^>&e ���-L(��x�I7�z=:�k��(Ou�'2��[v�9؀j��]\�#л�Q��'��
�5Q�m��ѭ�P���0>ɠ�x2E���v΀�4'2)�C���_�*��}��qCsZ���	_��er�'3B���Q̔a��JD�6�@r��n4�4�V��Xǈ�H��R}*�Pc>�ħc���0�3�����B��( @<C������RQ�������On)j�ᄝmf^=p��.x����V#w ���O��S�^��

D>�ەN�T�ν3��
6 B�I�R�v9X�c�[e���3�z&�"<���)�d�R��uk��ĳ�.�3լ��<�p<@z6�M��?i���?1��i��O�ʿb>-J�+��;d�TI�+>$����h��}"��)�Ѫ7��<O�����#�~Bl[���>� �4��m�-L��3$Ɲ�[�����O`q���'��{@T�4CI٥IH0/��}�����y���"R 9Y�� (�f�h\�4�#=E�TeC)2�
7-��J�@�ʗ�<��1$�
.'�$�O���O�*ub�O���}>�b��O�d�H��St!Y5L�j�r�+�|r�ǖ���20"bc�,/��]+�O^(��|-X?�?i�t۶��RB�9Ay2�E

53F2\��X�<���%$ܠ�A�@.� �ȓP]�4 �u���!�!R54㤼̓_ұO��{c��Ԧ��	���O:���	K -�!�' Fd}�a�'�J
�r�'b�fҽK���T>�3�Ƅg���S%h'\p����;ʓ{&`�D��gR�c���!D���а(�T�C��8d{b�>#��XQ�K��<�5���V~C��O_֜AG�A7��݈�C��df���k�	/o����$\&Ez��@��к73X���tmZش�?����)�AOd�$�O���3U�,l���3<f ��K�>-*&N�O>c��g�'1���w��V���q�E�*2��c�K��"~��m�rE"�C��\��1��g'j%�i��,W�T�<E���x��f-לz��c��' d��G Q @�0����/�N"5Fx"?�S����5{�X4ct�Ł57�lJ�f�A�"�'�X�:Ӭ��dh"�'���'5���؟��2Tp�a؂k� bT�·,{��	�,����d[�;8`1��I�QrU�q �2kn�d�*�}RG+w� X�c`���(�wEB�~r@�?iߓ[���D�ڥ �g��E�4��ȓ1׀�q�(B�R"�d��3�����)§���	c�i\��jW�>�H�x�,��O���'�2�'�rk�xVR�'���C�%�r�'��Y����6:�A�"� #
�	�w��'��q"`2m���&i>zxv��	�J����I�X�qD̏xzTҀ��=,��c%D�`��mاl69i&a�?NY�-�!(%D���uχX���3���Aт��m����}��©$�6��O*��|
7�Q�P��7��+��xVa�iraA��?���oR�����Ԙ��)�.UF�s��Q�H@I��	Q�L("�4��A�B�����*�c�7|vDy����?����'G�vxr�lҪC�X���Ӳn�!��5J܈����2fiJ	I�a|��/�D�;���%J@;Z���3�,20�$�*m� ��'s�R>7���?���?i�)
HL~�ڱ��Pr�L1����|��7"�*����a¬7Ҧ�)�tb>��L/R�b�+��<��m)5�J=N?̴[&i�:1�́ɒk׍d�6P����O��x̒F���`��;�l�c(��~�'��)�I"��-J��d��h��J���cp�!�G%l�*���f��*s-^"�8���?�#�b=0T
*�J]�r���1��J쟔��2���qG`ݟ��	���!�u��'�"o�"��R�N��#� Բ%N4�~�*����>aE�@s�j���o��D5�l��H?��Dx���W��h�0,�7NȊk1�8!sF��\ۄ��OZ���Q+&��%�&H$-�5�vo�l�!��C���pw��S,n��ŝ�z�©Fz��i�>�8PoZt�����E�D�嬌'oj�0�I럼�I����2i�������|�*����	�s餘�F��e���E��<~����d�"���[�����f�
�;��PV���b��'�~��MԦ7�TCw�,<�*)�
�'�fU�B,ܸX)��i�U�P	�'�~aBQ
@<a2l�#���N�n�x�'Z�c��16o�M����?-����%#;g�	RFo<E)r �3'�!2z���O�$E�
��'�|j�펆F��5� ��Y� -��L\�'PH@��I�2mY��2�Ë�Y���ʔ*SQ��Z1%�Or���O�ĵ|z��L�KԚG�%k DY�����K�S��y2�m����ߥS��1&���0>aq�x�Mv��R׬M�=o�����y⡈�j��7��O��ı|*q��?����?yB�Õ����U�f�|1��E�/����������ɇ[-�瘚P'����H��f}pC��{����2��{2d��5���.�X1̟<S�x�g�'n1O?�� �u���#Dk������jAq�"O&$9@뀈��0��f���@�"�HO�:g	`�Zq�Afg�qQG�V<v�������v���p�nQ����p�	ޟxY[w�wf��$N!g�����VG�PQ�'7ԉR�qL���j��l��b&c ���t��m����2�p-�K^�
�<xɧ�Q�i���Z��+|O�Y��`��Dy8M��J�_�n��7"O.=ʶ͊�J�6}�t�Ǳ6���{u\����T�椒æE��)�:���0�ғC��Z�ğ���ş|�	�g�m������'`�ʁ��Ɵ�ؕ��-(��(E*Tx�kf�!�On�)�X�	7��	kA�ĩcj*@ =j��2�On���'N�� sV�۔C���5+�Y��y�g$D�P��2��-yRT��`D/�y .Y�.�a�˄�lDfP��&��yR-��a �Hߴ�?)���)^���`R�?Ҁ���k�+��y�%�O2��Ov��!��O�c�ʧjA&x򤭏�O����$�S�|&��GyFT���|�Dh�
Gđ:�'
n�����I NH��=ڧ`hݺ@���=�`��1�̌�ȓ4 �6����9r��N�����I�ē��z����{�|<aׂ��fE0��8����i���'&��/#Ȟ��	���I�TF �cB�9n���iA蜭S�e�U��O� �<�O��Oj�؀㏘l�8�AQ啦;}��!1��=T8(��K>�)��X�GI*��y3!��─�`�%y�\���IȟxF������Ǆ�)��Ըp�\�	J~!ϓ�?9
�\��Sd!�:�ֈ��O�LV�Gxb&5ғ��G � ��(��^��d�D,�2N����O(��o@�5���d�O����O�`���?q�W;�șFd�(��M��B1u��'�
-�)���9MF{��+	�@12J߂U(L�j��R�u�D\.�,�Ɇ�R�5��hO`�� �fm�mcl\"�ֽ�$�O<8k��'�R�|��'�R^���%�M������9,�IF�?D��ـ*W�KJn��]N�||b,@'�HO��qy��#c46���*�� @��R:���aX���d�O��$�Ov� ��O��$v>�r#��O��d�+�F��e@�+�$Dz� KK��|b����?� \
��ڠ����R�:��|R���?��&���Jf-\C�^d�uGрkS&ԇ� ���0��]�*�����I��Ն��ȓ$��=vFA�r�̀����=fK4����O�	���G榹�	��d�O���g˿:�V�κJ�${�gN>,{��'A���q��T>��F
4݂"&~�BAPj1�#��yD���ǝI�j���k�	"������<�(OF�#��'��>�Z���XSFBTq(��I3D��0��)��P9���J�6,3�6�O6�%��K!�;a�:�2�薟c�<Tk%s���V%O��M����?�/�XȨsk�O����O��#3����9�
E�j�3��X.����*�|Fx�D²���3���<Y���W$��RN����)�矔�u.�?/V�0ץNQ�e;1mF9\�"���ϟ`�	���G���$�0�
��Y� �4��#k�Γ�?��19s�)'V�ȠFS��	Dx2�&�S�d�޵0����MO:(�	8R��9r���ʦ\ 1VN�N���M]��!�SV`
�\�a��)_�U!�D[6e�T���#�t�`��rN!�D��a	DЪ��ӌs@��ز�0E!�,��lɤN�?6h����k!��$���k Ҝ 0�$�'��w[!��,
=<����%�IF&J�u!�D�3@�I��H"���F!�D�j��Y׌Y{Ҙ*u�,4!�� 9h�K�K\�&	��@H G�!�d�':N��Βj0akt�٠+�!��;��DR!�=�(=ɢ
OBP!�D��~t!�f8�$�R�H���!�$X#+L�u��+sƘ��甦V�!�$�;[�F��Wm�3S��t���	vy!�� N�z�#3�]��j�=SzB�E"O,���'�b���U ��z��%��"O��V�A�z l�S�\S�yz"O̘PQ��?����ƿ�f��"O�8�1���;FD@7��;� ���"O��H�#8��j�'D*^��"O��h'�#'2u�R�ƩP�Ju�"O�}��b[�>�V�0R�p抭"P"O��#G��"���ǅ_�A�����"O�����X�09���L���$"O�}`���$�q
�G�F���"O���A�1:���MK+��su"Oд�c�ڴ)�:����ޕzQ#��>�������O꼄�r�-kڒ�����!����'β0���Ȳ%(�UcB����yB��Ns�̈́�	9|�6XEΰ���řk�nB�	<6��#�!�+�Ў#�T�S�� ��}b�@��>A'��1�pY�C�N'�����)�I�В���<R����5	����H�<�s���P5L�iv'�Zo!�$�hJb��@8X��ت+;�I�0������fe�E(�����(�&^���C��:8X���p<�x �h�8m����P)
�Cx�CC˙%T6��K�q;p��]�g̓s�qdc�>�ȥ�#��5�hɅ��3��p�҅ۦI0T�X6�1���:7�[jݸL؀Kԯ!��<��I3<Z�*�f(a�tͨTȖ�HT����@w#@)"cW�>4e��5Ot����B-=4:�r��F�f�l�v"O�P
Ee^)���d�%����᝟�1�����l�|YA�!W�O�Tp�i����%�14K2���'#a�0Ώ����蓎vӼ� �� Hk���'
>�j3�-�Ϙ'�V�JRĀ+x�J�H�ܘ/��y�'?V�H��'J�XÅ#Md��{��-��|�c�������
Ğg*����Åw�nm��	=��=Q�G��>���cr�,��o���b��b����G3D��zǋ�b�<·�X,
��a��#�<�� �&"1(E��S�P$��F����n��RqJŲU��
 K��yRD���Iz�c�_����S�Y�j��`������M3�#��*0�W���}C	%h2L�Um� ���	�*��?A!,�2
Pv��ď�=�H��I��(*��(�cG�|牄?���	�k��H��Q;6.��'B�=`�"?�rN¬ڀ�u�x��W�(gzI t�I�V�Qz�O6U4�zG"ObH�$D$g�n�)� NSDk[�8p�\�D���&�'�$m�*b�>J��܊RI�l���Mn�@Sf�>D�hA�LM
���9F�̓!됙1�B���Ģ�&���?��9S����{L>bA�'6��zCD�9��� MDn���f Q #�A��ES>jn�y�m����Q6
�|�4�Q�7\���U�'�P�7o��}ƐA[G�K�`k���
Ó9�d�1����Yw�5( �A�G�Lb|��+8侈�Yt��B�	�w?�5���O�')6I3R�$�ʓ���� %�-��QF��/;�~q�S�'{�F����	�L���ǧ;���V�D Ub\��p�Bw��  Up�b�FY$�Ɣ��S� ��'�	�4G��'ORq�O �R�4��	��q	�b�����W�S=N JF
Z��IӁ(�)�z9���4ᤠ����]r���'�2I�mIQ�z��1,}f��J��Dڐ.ˢ���#E�yh`�1'�G�)�d�.p�)�Ǚ�;�X���Y�����'t��* ���s���s��n[���O�������t٦ŀzj`�X���vȋfݜLB��At-�|��xB�"O0)B��8fw]�u�)?:r��4��b��ar��e}��ǆ�ħ�,�𧛟��d�J/i1��`"�Y<���;�O���`��)\̎����ÍD \��$�F,,a������
i�<�J ȕz|���Ą�M��.z��(���y��\x��R6fS\e �$LO.�PF!�i.2j�W]N�b�AƷ���R�M'=� �k�,@
��'�ԕ[ 	��'�	˵i0i33���B�K"��c�1OB�I*��#�]�	�s�x�]��>E�Tk��=���Q盜1첸�׌P�&�^�����CN��"<pK�JMV��Aj]�KF,��@7$P��l8[$քx�l4�?6#Ҝ[|�7Ms�� �u�`фC�-��	�1�l���X�T�7�_e�ؚ�!ڱ!l<�x�� �i$l���*�D�X���1��I{��D92���Z���3��/Su�1S�<����P &�� ��GϪkZ4 ��	3� `�o�m���R�iM��X1��KP�;�<H �eTD{��9�t�'Ó�aB:�S@�X�G X0���I
T\����U�@QPV)޷�h�(���!4BQ��b� -�� �����%7a�T{�Dӑ^��m��<6��jP�7�����_jn�aw(<,O��rQ���v�Xm�N)���h}k̎�z �qB�}&@`���/~�F��#���Q C�ٟ�*W���j�hB�Q<XG�MVMĚ?� �>��;��_;n֨�7��t_��h˘cY|4/M+��B��Ll�
��'~ٯ;Uy�3��#�y�B��F�
b"��@��[��0?I�N�����Ul6x��2�JM��رiZ|�fa`)O�4 Aoߖ	�p���]%^��͡�\#��I3Q���Q1|�M����)X��#>i�+Z�>!�4�&�_�i1v�9����"5#Ul?l�X�%�E1`@�2���Ū�5!��`�4�J4C�d��ቂfa��x��̎Rɮ��v��,e�I�w���*��
�-W���Vn��&�6mS�}e\ ��"}F	�2��HHF��J!��ᔱ(�'?zEV!�	I�pm�q��/1z�Y�G4 ���'�*����@5�b�r�>�	��ʿ*nx���
s�XI���',$��'@����%r��ˎ7Òq�G�=�𤌁�ԸI�B��]�$� ʟ�m��I�J7��{�e!zv`E:!k�X:�">)R�V�5/�m @���dL�CW�<��Ѽ,}���Ď�	E���@�:����o�l(�R�� �1�����پd�� E���)�]jG�PCy�����v���6�3��ɞ$C�4:(�n^0\*���$̴��r�M�c �����wF\��ã
�Cj
����'A��	zc�U8���PWh�7F8`�w��a�i١p<`4wn\�(\c�`�"P�¶4c��
_���X5���i��	��'�$j�	���(}k&G�#Ul�J<TC�I��KaD��f�1�mWd�'�� ��F���ʘ8��}a�O�9h���5X	��h�"Сe�<:�.��6�Z\��h_�v�X�#<O��K��U�Zh0�*5iM=�*(C�FH�4HZd��È������$�ax����.I�K��n���AG�̠�y��ɵX�Υ���u
Ra3M]6rϞ]���:
��(J�%�5Y��]�bB���'iO `?�H�ħ��e������2��pV��� �r��SEC�x��z7���)�fq�,O☩c��4>n�����Ä��U���	Q��xg�� ;��sd�M*y�#=�W��h�^���l�=&�8��.�j}�d)N���A�=1Ó��	>�֑�p%P�[Ԁ���	�0�fEc�爯ls�����-W��"<���9Z�J̈�`�1Y�EI%�]�����!��2D�S�]|10uF�(7(�B�ɉF�bbHQ
gn����2z�|��UhTf��u�(+h� �s��i��?y�D�6J���#�̥ ��Ť�r�<)�G�"�*F����)K���q�<Y7�K�x-���S��!��cE��w�<�6�u�K��(Vx� B���B�I5�e��M?+�8q�T��~7�B�_4��ᨍ�
]�̳! �� �.C�	�#�z�H��["վ|�H�z�lB��V!P�D�د<j�����%i�B�I�Y�r<3Q	�76�p�ULE�	�C䉙&t�j'�\�/rP�2Mΰb�C�ɎV�еb�cMpm�΍5\1�C䉚cF��a�WN�рG�&5�`C��<.v-rR�Y@G�� ����@d⣢L5~إ 7�#A R|��+� ⦪�t@��S�"oP��ȓ&wp���L�%iиxG䞵S����do�	��y�S�OҢ���@O�	ꈉ�ѬK_�Ձ�' �d?��m#aDɟn�$0�N�����;�^i��"�z�1�ٕt^����S@�����1:�x�u�A,c��db�x�R �FcY�.O
B�	�`�HԘ��2"���'��[@�>Iv�E���É�$�[s�v�p�Ԯl���Æh��y�( ZO��s@_<]�l�$��~�lޞ���Zu�|�����I��"3�@m5j_�a!�Ĝ�6��@�l� �t�!)�36�&	�DCS���<���=E���E�$EX�9R�]��@�$�p�l%�!��u$?�S�d��K�� %H?R��=@th�5U�.�����t� z�Ǌ��5��Xt�&{s|�����t�hsA�A��S��{�'Tn��b0�G&P3��yG+�T�F���P퀷�@X���;���C�&e鶑��%6B��"�O&	7��'���h��aZ��G5��U��E�I1^\xUZ�4����6�8��T�{�ƙG��@�B���+��-X������I�YS��W�'��%hwL[�D�&�)mE�y�d)so]�rϤ����F��NA���gy���,��"�H�� c6B�>�氋��'@��Bb�8N����BkV�X�A/�"LG���ēJI�0SE����&�Y�1���EBL�3\��~�D��(��	;1���q\�Y�bQ�<I� ��Gʜ���N�9d~9sG�
fy҂9=���=E�$	�!2��Z��jj�h C�O��yr �-�dP��ᑜh����̦ޘ'��Q2�-,O"���c��A�m��P�}���ku"O�}�$W�6et|��b�8W���B"OhXP�NK��(s� �6}�Lc"O���D��&�|�� ҟlw���E"OjD;c���n�$��$Gt<��"O���G�4tY�i��5N���%"O��!�	4G�PW�@�P��Ѷ"On�:��[^��Xxހ�Vœ�*O�͠�D�0/9d�fË�w����'84iz҄M&}��`k�Πq�'�=�f#�<�^t��b.��
�'Ϝ��E.��_9X��n�c�8$�	�'uM,9EN 2A�L�D8�rf��p�<�#/%E'���r�O(+�&T�p��l�<�@NB�ke� %)�R5�ta�t�<��J�Z�x�ǧK�}4-
Ҧ�n�<y7-�)!\�P�g��"H�ţ�O�<��R*)��,36��~~e���P�<�v
ӓ{p�������� �E�<!��@:�(��3$e"�Y�'�L�<	W���`�-(�t Yg�R�<QT�T�K�" ��ʨb��b�Qu�<15
����}	�EB�}�ll��+�l�<���_�eO���'IB,b����&�h�<	Ɔ�2Q
��r6 �)(_��:���<�[hq��̍�#����'��\�T ����$aˉ=6��{P!���ȓrҤb5H�\@$܁�̉�Z�¬��yR|�s��߶G��й��V,�����g��� RC�f�����_>C�*]�ȓw��J�i5wb2���O�:8<�ȓJ���S	ك!�2�� ���R����"�dM{��Ղ]�r 1��oZ ȅȓ*�V��T���b���g�O�Fs0(�ȓ	�*��F�3
��JF��->g�i�ȓB 8r�AD�sɦ�A�c\+k�`��M#�qC���D�B5��(dن�w9"]�����l*����1l,E�ȓJ=�=oאM�HMU�$���1D�X����
+��(��Z0:*^��n"D�<w���s?�Mk͕J�*����>D�$z6�:U�r����<X��S�<D� ��H�����+ ��M	�;D��bb��Zn8�a5����s�7D�T�Wf�/\F�a���M3Cڪ�s��?D�h��)�rR24{ƌT5����+<D� ��+!_���4"��ss����E:D�8(�I�*#x<�#薱�X� ��2D���6d�3t��l8����($;6%D��1��6%W|E�5đ���u�#D���B��9P4�xh!��Tv
 D�� b`V ��R�h�C����3T$���"O9����P"ԧ~�T|��"O�zp���`R�=�T
�"O��\�>�2T�@�H&Ar�Pv"O��[�e�Z,��ɼ8Tʼɓ"O��iQ�GOV`s6��ZR�I��"O@�Z�F*?\Yp��)^Q����"OLk3� �\�b"E*���"O����*�i^���\#�Du��"ORA�oŅ,�С�a˽��M)�"O:uJ�)M�p��P�0M{+��y��*tfA���.7��c�D��y����C����+p��	�a��3�y¢Z�X9�pr��R�g�v%��Mߎ�yR+ϒ!z�X�oY�c[0jA�F�y�D�S��b�/�;l�ȃ�H��y��"_��
����hd�x�g	�>�y҇IT�.Qy�EExTy�J��yRiB���� q�Z5�L�hP���y2i'o�tٙ0�ٵ�(�gͪ�y��S��c&N�r��%8�#ͤ�y�D ���GꉮbBTS�+��y�qۮl[�ȿL B�c�E���y�}-�h �GA>Fw��Ї
��yR,2I��qO�C���� �y�Mpꀻ����A��(0���hO�����J�y Ȑ�i��$s�
�� d!�d�>�t(�l�]�d��)@�j�!�h�!c���S뺼A㎸_�a|��|�"X,&GNd��嗐iƠ�� ��)�y�)2p��U#s�4O�Q�!⅀�y"�̜r�t����H%�����M��y"h64����B�N<�X����{�<I@C�!dH� Bb��>��ȩa�<qv�-f�Zh��% 	n�� o[[�<�VhIv�B�2�S�N	�4��S�<W�ڀ
$fI�T#�"���&j�u�<�`�է:8�V�\�.)��Q}�<i�ᘱ?c (��C�%I���!l�a�<�ϛ>{.6��E�O$"�x<A/�]�<9M&�4�k��:[�\��ӋX�<�b�U!ͮ����ƸQ�<�q�MW�<�g�>P��ϼ�V%����]�<�w�1;D�ԣC@�=O7�A�ǧW�<�'
	]���yp#��f���-�U�<Q�e����=)l"�V�KO�<���EZh�2K� N@��Y�)�K�<�f�E��}Y���pR�i�J�C�<ɷ&�4'�.d9���>q7�|����B�<� �Pp�$G�_�^ma)T��Q�T�d!�Y}���/8D���`'�3x������tD�B)�hO�S�2�t	 ���>| ����3dlB�	�LЬ&��Jl�@�@B�ɖ{
�=�N�n]�+�;A�zB�	� �T��t@�*�	���	3B��#$�ɐ���H��B�׃��B�%;��d$\n�$���E�Z\�C䉎;"�0S�mЯL$���-B�b	*�;S&*"�<D��C�C䉴�E�����Xyp��-��B�	>}��b���;)�-�:�B��"$@�[��L)�Xa���3��C�d�xr\b��<�3`���C�)� .̛�đ3\�LHs��%<�&U�"O.|1�$�#���)pC�m�q"S"O&%��E�w%x8SFb �8�Zu"Ox��L�,C8U7!E Yҩ��"O �iFk��&	4�rр�,<�Q��"O�m
0��?M�zi�� 
)<X�l!�"O�T
#X%P�(-��A�
sF���'��O�usf��% �DN������'�'�=P��&,( Jwn�-S}�����2�H�nh���7x�&!0�P�O#�4�ȓ{�^�G�AjX���'�fф�'[��BS���ZLz���E�"?"��k�p�0��Ãk咰��������Z��"'�
P��bҭTg��ȓf4�B�)i��	R��+�̭�ȓQVnHS$'˩oz��%%&?�a�ȓ)UZ��7-�P�r��Ǒ9z�昄ȓy�x�G7;��I��Y��J݄ȓi��ӷÝ�W	hM�l2 �~��ȓtR>�q��9���	�$9�2�ȓH� =J��ܚR�Jm�!H',��ԄƓq~t�8���&.���1e�?��1R
�'ZM(F.��j�(
�]OȄ3	�'Iu�j��8|���L�4Z� L��'p
 �#I�A��칆���e�x� �'2�hq# S�)b�IAk�`$�r�'�~e��Z k�$IH`�2B��ab�'_z!���,[�d$�`F6	�B�j�'e^Ș�L��a�ɛ���)qQ
���'�N�����冈iaG�:g&�xp�'�����)X� n�e��'�<4 '۟sg~x�e�R!h#�'�B�Sjӥ��%!��D<�)�y6��Q@�Q� 2��@�y��\�H'tpڅ�Ez��x3�
�y�B^�8�
т�s���Q���y��S>,�F���bn(�쀠��%�yB���eS2͊򉈢_�F��B'0�yB��@$�$$J�T�4 �c��yB��8��|(��>BzHRP'�y2m&E� a�a��
8�mD(�y�#ư=�,�ҕ�� Қ,
�@�yB��d�H��A(�u^��Ud�>�y����Ej��Ć��a������	��y��N�BIabY�S8u����y2(�z��a8"E%8�V�Ѵ�����>�K��8��D^7V9Y�Ę�z%�q�AJ2D�D1��# �1�	�ɖ���/T�HS�'�(^R=��
�7�$pYs"OLH�@l�4k	z��`�_�*�ZēB"O
�UNN����B��)�,���y2DW�Jv����i� 1�6A���B�yH?%�h�j�m�7�J@�Ҋ�5�y"��
��T��/���r%l]%�y�M�$�p��1C
;����#��U�<qb�O<r��E��x"��K�G~�<i�cF� ϼl��ڗeԔ��	�{�<�E����S,	s.�����m�<�$Z�t *�xƉTrȈ@8YA�<YT�-i��i�>Wn�P�Bg�<�U�� ����gΊl���X�<	eՔNT�;���yY|	�&�SR�<١�At@�@"R*�v$�U$Ms�<� ��RI�5#q({�6ء$�v�<� ���RjS��L4;��C'a�%��"O���&�|j�5���[���E"O x��kNnUf���c׭>>ޡ�P�mӐ%�<��t����|�!qR�ͫ3f�Eړp`!���Fm �Xd��C�f�3�)DF���/�����X<L��)㇪ :,�l3%�**C�z�	K�#�杈S\������HS0�)4�Ók�$X�!�&?A���.�p�ɷ��{vHa�^?U�xB��0T'Dd�4oQ3~�.��0���.˘B��M�z�#b�Ѥz��5�$K?\�<B�	�Tv��r⊖{���D57��C�	}6Ri9��d�LȓTL�/T�XB��mAR��d��
i�K�%@RB�!��a�J�r��]I��ʼxjC�IA B�[�'ڣ? ��@caǗDtB�I�6��Q�rHW�a�P]"��;N5jB�I}g���''X<�6!�V�B�e=*B�I=	��h��m�tF> �r߁[��B�!b�*	Rg��+6zIa_�\e�B�	�+t&�kW%�cl�r���5O�nB�I6�z�ࠅ��(T����%a="C��5� ��i��F�r�+)BB�I-QB�t�s而
s��z��9�B���n�!�R��U2�ߜ8��B�IrѬ�0v� ?��s�*�
(��B�J�L�q��á��Hp�Z��B��vi�E:k�$D+7h^�b/�B䉓"��h�4+��4'��B�J�B�I�3��	��ņE����*U!�B�9h���8�H|�T1@�Ŝ,�fB�I$C�v�cgC�K�ꡢ����<|B�ɾ?�8�����p�De���&B�	(O�Ԭ� �TGP,@��ݎg�C�ɝM�Y�F^�k�X ����"}��C䉱JX��F�8-��J�.��i�C�	7g3������2򽒣""{�B䉄d��i��IE�ڝJ�"A�*{�C��8{~��+�傍C��}8dO�<3LC�	B��QX���a���[20C��F�R���+_���T�G�I5�B䉩Z�Z)��H��vN���t�	�3jB�	�X��(��J��M#�t{�I22TB�	4l\�CHvӺDb�+�t�ȓ}�,ѡ��Be�95duxS�OU�<1P��4�n@jFM�,7���FPL�<Y�M�C'��w�^.`����˞�<�f��	HjS�R��xj �~�<� V3|1v<�D�T �$)�-Vt�<9-�I�v�1�O�g��ms1�s�<!v��?l|d��k�9j�H����S�<���9>Ƕ����5� �a�N�P�<V�:Q�U.;���uN+�~B�ɲp�`51�·���	r�؊ xB䉘]>z�v�^	�~a	��<ZB�	�:���t�-`���偏:	�B�	" �.��T�X ��H�o��D�B�ɗG�@�Yp P�OO����� iB��w�`��6J�!-(��S��(��B�	=C���#a�0��0�i�2E�B�	�h����$�7[nH�"J����C䉆LP��KІ�>*�rUQ�$1��ȓ�.9)T�	�#�`<�&��i���ȓ!<r5b�Z?#+�8HE�?v�t���bQ�zbCI�>@�&�� Z(�L��S�? ~�kp��,q�]�w��6zl�"O�a�l��!m���f �uZ�IQ"OVM��oՕr[�%���3S�=q�"ǑV�����t"�z��%"O�48��!LaQ�!$��d�F"Oh�B��\�:@��į�QE��!"O�F�$;"J�+a�"O>�1EG5d)5�]%ުQS�"O�9:UAǱ\M�$@��S���"O�\�����n�a�M#����"O��G���`p��] 10E�b"Ox}�7�+<�p(�l� bR�KF"O|��d�E"Ⰲ#�-V0Є��"OX,��26���V�'����"O`�:���Ge��1�F1y�3�!��^8��Z�铯:���j4��0n!���|���b�Z�"�VA;�/[�/h!�D�M��� e�J�o��)�T�	n!�A$е�Â�),�p!"��[� �!���B�|�-	��.m��LV�v�!��"޶�U\�5����d�B K�!�D'Z��fEZ�њ`	ꁀT,!��	%�  �"B>hʀ�5��!�!���
L���=;'J�e'� 8U!�,��i��	�g#�|b�F�,R%!�$Ìj�4��Azv@�q`�K>X!�$���,�R�ƓSdf`)t�V�l`!�$���Ĭ3�l�1CG�q���5/\!�ď�4�yZ��a;��KrB�N�!�D֧3��0��Lj2��(��
3^{!򤟲y�P+�Mr+t!	���MC!�$�H
 �PnL�Š���)�!��Dg���h���#k�h�V+ڊ	S!��#<����7|�.��&��!��L?q����R(��q�����)�!�$@V��)v�V�zu`p-��mk!�d<Lͨ�AҎ�m�>@��)�f!�d�@r��a��5yA�ɱJۡ!S!�� nЄ;#�Y�z%��Q./!�d_��v��1,	�����$f�s(!���8r��x�����D�"!�ҷ-a�Ib1j]�lZ�ɰ,>^!�d�F�4�H�cA�D�^��5K[�z�!���0t�3���=�m�J�
V�!��d��;рQSPd�z�
'3"!�dԨnyE��*
�NA�zd,�67!�dр2�� F��09����z?!� Fp
0&�ԼAȽ�C�ʁJ?!��,���K��U�A���C��4HE!�
}f�]b���
������4:!�DÈlj���J{a���VwZQ"OL�C��,|��0Kr,�b�.���"O��FhJ�]�
P�L�R"O�Y"$f�*_�I�,ĂDx (˦"O���W���D�Z���xo�0��"O�X��fL�:̹QcILD����"O��j��%�J��󈂚��]A7"O���t�ݨyvl(@6����� ��"O P�؜d�.���]��p؀"OdE{DDBŤHSe!�/�Ҕz�"Op��H�n��H���	�^��C"O�݃`lM�@�Б�C3En�A��"O�ҖAJ0-|WH�L_�EI""OJp�Q΃���	��Z!bV�M�B"O� (L�3hQ�!PJ������yM���"O��A  �u� �!a�ߦ	�n��V"O6���Ҟ�N@��Gk����"O��b�
�ga����C:=��S�"O��hP���pH���{��S�"O�����3V؅�`�Ww�P��"Or��F�kP$
�'��Lն7+!��'�b1�JJ�fq80��KH)`�!�D���u�D���<2���6�P/R�!�$��!$��g�� öI۲�Ĭk�!�Ğ6y��� �ȃ�>���CB�o!��[|��a��)tH"��r�ֵJ!�Y�BOH��+�B&�h��ҩ`�!��¿<?LYʱ��V�!���D�0�!��\4
�$d����1*����D�I��!��V8���Lu.A���\�p�!�d�#iv<9G��8Z �3�ڄn�!��C�.��јVnկ��4�˕�2�!��55ǐ%.5�Љ�7I�Z��1K
�'��0��g�,�('�$f�H�	�'�Q���\�J�_T����'�zi��Ĩ���ڗ_yD���'�t�	�5	(����!6h��
�'뤥�s�=.r�|b4�Q	��qH
�'纀p��-/*|�Qug��	�<�	�'��Q*S�]�XpMs���˘��'���[#��;o�T�s�G�F[����'�.�aWb5`�ha�2I�Ѳ���' z�a(ѯ{�R���[�z ��[�'7�`2���H[BA3aE���8M��' ���7:b^��UR��'��z�bI�
���OD�=P�<��'�(�;aPW�t�'�Ă���'� t�eǎ,��s"� �z���'d(�
W�Vch68�3�ѮB�T=��':8`� �2t<��TB_6礀1�':�Ļg^�� A9'i:�����':.`rr��!�� h�OW0�65��'Ц9�a��=0�Ѫ�� �����'3fppq#�#<iXU� Sf�|ܐ
�'S�¦�8��Ԩ�O/��j�'�X4"� ^�<�s�_(�2�x�'\�5�P"�b�������8�'9ƕ�1�P-':��I��1��'�@���X6[z��7d"on!��'�b8�(�%�hf��~�D�a�'��lX��� ��$:eH�#�}��' p���cX-;t��J���$O��']��(��֔?z��0JҦ! 0h�'�v��aY�.;�Uٷh�A����'Ȏ}�$	�.f�6A�6��`di�'� %�7�Q�#�%�%�ÅV� �'�Ri9��$R0��t$�=a�0��'��A��`X-^������
p��Ms�'���.2�!�ClP�`�'�})d�6h6���-��iŶ�"�'N��S����>Ju�'O�#_`,	��'��Q`�30``��3*�va��'�ڱa��2v�Ve�DÞ.T`��'3 =�4%ҸH���Bd��' �>1��'Eb�IE�L�B�A��ʚ�G�:�S�'>� �w�"p?(��@�L5=�&	��'���a�d��gvJeP��?g�L���'?�I����XM�����u���� ʡ��/�5F�zY��N����`D"O`�1BE2K{�m�AQ���"O�C�Ǖ�$�L@��=-&���"O�A�DU2N��B��L&� 8�"O�t{$��e�t�들�03�ؼSE"ONyP�@�x8�g��!lu��"O 1�#��q�ި"�e`n&��U"O��@T<����޼Lc8�I�"OYw�Kq� ���Ȁ�m�8�S"O�=h�Ĕ�[�X�2b�V�:D�"O�����'$��B#��|4]I�"OXaqC�69�2�:BΘ�q����"OR�s�NP�8X𩙔���E@D"Oh�kԥ͗Դ�P��Ms�p��"O�y:�0|k.h{��I�^ꎜ�"O�aUgA����� '�z�.P�q"O4�i0��e��"��!]� ��6"O��C�HW�������f�"O"�	�n�o�|�a�{Ebm`�"OT4�����`S��Ե�S"Oġ�A)�����N��B���@U"OXI��'/�Z�bE���s8n��D"O,h�'!�@BCG��	bR"O��Zei�
x�� ���L�pBc"O
-��)�/(>ʼʖ�R�n�4�е"OH�8�j�<]�p"�gI�5�8�P"O&X �ܘF����ť�75Y��P�"O�8�F�f`Xa9�A;	M��Ӕ"OȰ�4��[~pJD#I�PC�"O$lp�@u�P`��\!�18'"OD��"l��Eu��@#��i�zͻ�"O�� �._�Q@�'�(:�f8��"OT�[P�/�.����U;�)��"O�͓�Ň�#��!��E$[/�	T"O��;�G�'hS ��2Α%Z�#�"O�]�  ��6�\�8��3\]�a"O0X����dgĠ��ۜM����"O܉*�'W�g��\����C�*�R@"Ot�"�D�#0��E������2�'8�M�t�֗G2L���ۧX����'��9b�� �#M,�E
�<Q�9��'�t�f�T�q���qk��H�L�
�'^�)��;�^PApb˵?)��*
�'���T�Đ5��p#G.�7���X
�'�b�;��ބL��P�eM�cGf���'���6���H9���$�M�V�� �'Dj\0�ݶ�p����EV�0�'
��UB%����C��88zbų�'��k���X�K		�`L��'0�QA�φFǖ��+��:�'���2A/U&�4xBIָwH��'�p���ľư�	Ҍ_ N�謪
�'��8�،(� h�G8N��5��'tb!� j�NZ����xb�-r�'��9�B��F}����딐&t����'���ʤO*x*��t�� .P�'{��"(Y�j#"a1�d��L��`��'�f͸6�Q���QD��q��'�H�����
	pQj�9F&V��'�)��P.td�P�F�Cج, �'��c�ٟL�\��Ȏ5����'6(�R�,���]SFn 5d+�D�'��4�L�7^���EJ�������'��t�]!
��X��8G�1J��� \:�ͦL��ACAO+V�I�"Oj�p���8�� �-M� +�"O���V�� ��0�c�1b�����"OU8 ���\@ڕ�g��W��%�"Ofћ��?�n���iO
�M��"O����óY��c7�q���2"OBL8e�ހ���:�dٛczإW"Oh�ʢD�1}*����k�eF"O8	@F>v�P���≣7Z�2�"Oĉ3B�Z��̉DP<_G�	�"O�Xj6�γ�Ba�VNk*F��"O޵[��^"G\���d�ǮTY��'R��� N�'��+7d�*!�X�@��6D���*
%B�,�[⭛�o䵉�� D�T@̑,&O*x���/:��q ��4D��/}Lb<��!�;]7��*�����!�S�n�!R�[�`F4�RD��+�!��<��h�a� ̶�����67T!��X���)�&��!�+S,>�!���3PgT�p�_�_
�x�E^��!�~�¨Q��"d�j��'e�:�!�D��Y@f䃵��
|>p#�L�n0!�ZU4Z��2$g]0E9�eG�/$!���/4���Z�̊OM�u U�$�!�DX=4R9x��<��� �Y�C�!���X��1,�8'�LZ0'Ϯ<�!���4c��!���&c!��Q��KD�!�č��������M"n�3#�� �!�Ф~� � ��4J{Ir���%S!��	q�VF�<,z��x�σJ!�^VX���?p^�-c5�X�}/!�Dj�Rx�􋟗"�x��� l !���$ �X��GR�w�\�w'�0Mg!�B"�6��b�C+3c��vF	�W�!��!!n��T�Wč)$��!��(+Y�u��+$C��Qq디�!�� 	c��@V��(�YHT�=�!��F�{���#+ڱ�� ��!��H
16JlyCDłdk� ��)�>�!��B�-R"��f���D闅v�!�X";��	r*
hk�5a�3t�!�d�qbR�ʓ�ƿS��z&���A�!�$��SI�$APM�
xl$
G ;w�!���o���+��(\�<��m#b6!��4�y	q��>�H��T��>!�^+�^A�`�_ �p��p� -!�N�.�Tw�[chy����F!��S�H�1 e��X�ܰc(ź+�I]��(�&�+Y�e��AbSI�m\|�"Ot@@sF�fH�]Ca�K�:%�c"O���#d�4I@l�����#���+p"O
���ꁹJ��DҒ�Q�3g�m�f"O�) � ̋U�X������QP�"OfL���5)�بF!	y�!1�"O
����XE��X���ߠ-��"O �[�R0��ZF	��G+��"O����+�WR��b���+q>-B�"O� �@��fҸ���FL�O_���g"O�ԪC{@̔a�d�w5(m��"O�=(�ΚH�B�Z�$=##̴�D"Ofqq7�_M ���]K���:�"O9�pi��*f4Ⱨ5l��� �"O�d`ã�!&� ���!C��e��"O|l�dO_�ril�����5|���a"O� �1��M+l=k���+8�<[2"OHx��i�8�����(q@��"O��zG�N��N���ID�T̘�"O���ҋ{�ġ(��ܦH���7"O�Uۑ�L�c2���@	¨.��(�@"O��C�L�R�d�#�B;��<�"OH]�f��+[��P��Nؖt��"O�(���B5k��LY��������"O�qAGMқ-�]2��U&s���s*Ov�{F��h�zݨ���_Җ�Y
�'�:�͜8�(<!lRU3\I1
���d7W��d��ME7Z$�A'JÄQ"!�D �G 9v M�7P��� �؆	t!�ć I��)��P����i���!�d3��D�F舖 ��%㧉P�!�!�J�����u�C�B��+pOZ$�!��&30��RtOH��d����!�DK�U0 ���/�|8�Jњ��}B��/}G����_�r�H���!�$Q�k����g̷K3"�bbI&j�!�DђBU�H��c�:����!B�!�F�.�%z�KE�~.P�ǻR�!�F��iie#�Wc��s�ʕe,!�O�Y=h)���A�3aʭhP�Ģ1m!�dU�����#@�c��hP�
�w�!��҄	�"� �	�4/��O��=���٥�D<�iy�*W�L�� �P"OJ-8�������Z�J�������"O�(�e� ��@iߤ���"O�-h�BGC��E	 n�'��9A�"O��cd���5�lZ�B>\�F"O�I�u��Iڄ�R��Q$�rG"O��Zc�P
X��(� J+{օ+�"On�§���&aH�!ц�-�(�W"O�Q*�(ȊVxx�t+�?�d4��"Od�7B���'��)o$h�"O�9e%W�=xTQ����hh�i;C"O�U�f�/+ɖ5��U�P]�-��"Ob8��-Ñ1���CcX?PR.�KF"OP�A�a�.G�u�6�
iY�1
6"Ofy�4D�93ICpƖH(4��"O�iYn_�KԪ��C��);8���"Oz�IFڎ	2��1��]�{�T�P"O��pVHZ[����^����s"O�K��صE"N�i��_�^��@�"O|���~w�p��ޮ\�ձ�"O20���H��$�p�i�3$ժ��U"O$��E邖GD޼�q����x��"O&h���ۖy��iP[�<�d�y���m��1%G�|� ��NN�y�
���5��M"$��4�����y�㚊�ȉF�T}��#J��y�M�F;\C,��H��M3ӊF!�yR��=��pAa!�;E�ike,X��y�?7?�d�#+�9Ҽ��uō�y�NϒI,p����.@l��N���y2Y7e��-9soSm�>@ ��yR%���F���C�%c�����n��y�h���vL�ԥ\_h>�k��V0�y�Q.M���I�h'O�媄�Y;�yB@�2x&�Xb�e!�*�-;�N�a�'1J�ءK�H����
�3d�A��'����ԉ�1^`�$��/�P��'���Y�-\�:�-c�B5%	Υ���� �`$��-���&�+tհD��"O)�ҏ�(5J��eĉ5ѴU�"O�yk�Ʉ4�*3p���`(A"OP +�@�^�D�AF6N���X�d2LO�	�l��@�8(qB�U�V�\i�"O���ŭ��@���!����S"O*h��Jw ���w��$6�D�"O��dD6C�������u��Lc"OT$x�g�0G���AJ�>��dR"O�D`���2%��RFiS���9f"O.����<x��@��DV���"OЈ��_�'s���%,VI"w"O�9����5T������&8��С"OV��>i��)V㝚m���q""O��!\�VH(��*��(�!"O��V��D�"�2t�\:���c"O�q;��޲m���Ca�H�%FE�D"O�єH�:���KgA���1ۑ�II�O�ܕ�TD8:��RH�{��h �'�$p�V�X�4� ��ӊڅ	�6�a�'�$DYg�J1b��#Z~~�]��'�ְ�w�_6E��� ���w��l@�'��y��%m�j�F�inN�P	�'��dqp��={Fx�ڀZ�,�`i	�'�Թ�a ��H.��ceß+�JU;	�T� ��'��iH�
�<	�b)��U1=�ɢ�'J�8��)_/��Q ��@'�����'��hţE"kx��'F�2V��r�'S��q�L�9�т�h҂˜�@�'�p������eY�
�*5�2���'��9�TI0=����	 	4���'�F�S�_P�B�Y���9	�u���r�<C��Ы4��L��j=2r���ȓ/>�8yg�ؖr��0ׯ؍G��لȓs�M��ڔV�8,�g�U��`�ȓA�����	8=U�y�W螞+\f��ȓB�8M
(Dђa�"�$4Z؅ȓ7sD��&!���������K�����	�����O/y������R�F��ȓ�����L�&����PN�1����-�r��ӡ/t�D8�a�7��q��J��}��釁Q�����L��j۴\�ȓ��y�@��R�L22�/X��d�ȓ ָ��V蝔p'��"gݩ)��݅ȓf4���3
�3Oޙ�VkB�`~�Q�ȓiJL���. 9��R��2�j��� �����M5V�*&�F9�e�ȓ
d.��t"��1��	��
��ȓ!F��p��H�\d��cI�w�j���}l��SFL	���+��V�KrL܇�>���vf�56Ԣ|��I������U"�����),-�s2$z���ȓk�ܭ�T�)txD��d�	8q�l��Lg́U�J-�S���d1�ȓt�0!�@�(pՎD����VẌ́ȓE}V�ۅ�B�s��%һz�����P�#���=g��q�l�8,K�L��C(|0���;]��iEn�3��0��{uJ��H	!s�t�b�0"�M�ȓ���h%�5�)�э�~Bp��ȓ#4x�G�G����'���� ����`Ÿ#�v4��P�j@<�ȓ&H�Z%
q3���؁X|�$���i�� �n��e�ϗz�Շ�S�? �5+�Y�f3.a��&0Zsx���"O*%QW.��JL;�B�;eN��"O�e�&l��ă�rP��s"OЬ��l^T�F]'T�D��"O�����i"��R$�%(�h�"t"O��R�.ؼCڀBe)�VB�3�"O�� �Վw�ԭ(wF]���h4"Or��I~3�i�v怮X�4()�"O|�!�f�X�|�/U��U�%Ξ�y�MZg�(���PM@��I��y���	���b�+���ԡ5F���?�'	Z)p�JOj؉�EP���	�'4�݋F@H�I�fP�0���I�X ��'���9��fJVQi%�M3:�J(A�'HyA#�3�����CB/�,���'��(y��,�U�4S�Nn���'�n �qᏺT�A��e�*@��+�'�ܵ� ��;�S�l�$I��'������cq�@�`�9j�h��'S��ڴ�E1r�t�!�	��lPE���'�$	��ꩀe�7l���'!��� ��2�Є�N�N���
�'�h�a�A7s�r�#�hU-8r����'�t�E�3O��)B3�;X�u�"O����9w�	��D� ZG��	"OʝY�ՙЅ�V
^#u?�t�"OT!:E�C=T�!XQ��q���c"O��0�˼w�Z���.d�~��"Ox�귭�/���R�	�P��%�A"O��c���#,FPs�G5g�&�Å"O�M�v�@/S��A�E�"O͓2�xy��[�k?/T(+�"OZA��4���
�@�:JdD�K�"OPȹ�

Z����ga�,n3�J�Of�9���F @�A/<�� D�PZ���]�DY@��u��R�k3D�40�s[��Ǘ�7��)`�D3D�����4(��#עF��)p��.D��!��Vԑ��Ӷ`�=��+D���W#ηZ�*Ȉ�D�
c~�����=����$		��%;0(�7��D±K	��!�C�ar�dj���x�b��.'�!��T� �Wꗰf��Ȫ�����!��0C<�cЧ�'��	����`��}����ǐs���%jI1Z����7�0D�T0��ͤ?-丸0��>LƁ"!�.�O��<�d��Fb�-~%x�@V Z�K��ąȓ�䳲mE.= �����D�ȓs�0Q��CQ�`erq%ƺ1���]��4��b�
b��jr/3p�ܝ�ȓ7ш���l�h�Rā���,V�ȓT����E�չG^�p�M�1,i�4�'�a~rLJ%~\��G)��)4hD�ƉG��y��[����Cc	�c�uYei҉�ybC_=E� 	�d�(nX��,Q �y�.e�-��
����*���5�y�@KR�F��`9�`������yB
"OՀ���6):q��!��yB.Y4T�ᆥ�<'6������y�Jϓ�3Nb`ee�&I	2���"O6�ӗ-���θ$RLpp7&V]�!�d�i����rm�*#N$�EW�d�!���f鈔뗢@�t�I�E��
^�!�ί#|���/t@8⣋�K�!�� �5�ף��d� ��B&�LKc"O����1�*���$q�,u��"O؁5N�7n໗I��L��"O�m�Fe^�0$����q�R�1���5LO�PHN��{�*#'�M�E��"O�H00%�$��I�6e�6~��a"O���Kq�¹S�H�0s��c�"O:Q�-�s�.�bC[0S�4"O�,s媇�2<Ys"�y��qz""O�a��g�R���Z�B�*R�ԅ�"O�m�ӢN43�TTx�L�x@�u"O:L�w�'j�I�bX�a�9ـ"O�[�
����qdA.��%yB"OJ�)Dϒ�c9X��
��"O���dƺ|�y��P�3�bIQ�"OBy�ߋ��� @L�ղQ1"O�𒳮�w-�������hA�"O��1�ԩM��81�@�p�5"Ovlg�юP���Z�/ͮh��1�%"Ol���+?� �xGN�7xpX@�"O���@�J��c�mW�9u��s�"O0A�W�U09U�E�ď�^�Yz��'��?O0=ӆU#D���.�  "�E*a�'	�	�`4NYydX�y,�Փ`�,a��m�ȓL#��цn¸��)s����Ѕȓid>$�Ø�?�>�R�%2T��,E{��'���'eԢ+������^�"�)�'4u���Bm8@ʖ�c
���'��
҂�Q׈P��@W�*����hO?��l^�*Ԩ��Lݬ;��P2�(
B�<1���
vF��uJ��|)�@�Q~���ΓE焨���-���uF��D�����S��!�ۼC|][�>����(I���<T�4;�� �Y�ȓX蒌"A[���`�[eR\�ȓa����ĤiȌ��l׉$�����^�]�B�D�=�$�ꎋn����ȓR�Nٰ�eكMXՉ���8��'ў�|�aOhx�"ҬȖb�$���,�_�<1f���D�&Q�a�C/��p$f`�<q�HD�#׈�ڢ�w��ݰ�́s�<Q���	J��4��m�z�p��O�U�<�1iP�H�
��*.���V�<�aLSo~~Aa�Dn̚�I��NԟD��[����ɻ+��lPp��p�@�ȓ
�xl(E��"�8tz�/�~C�8�ȓA2�3ƠC]�v�#@"�kKXȄȓTjx�`r
&X��seJ>�&1�����q��	�$�→�@Q���:d~XXP�ˬr�W�(Ժ��1D�`���c���,�L��#D���dS�'4���-��c�����!��O���4O�0��gAy�� ��
��Q�"O�h{�&X+JÜ����4�^���"O���!��}����	G��d"O�4���k��ث�"���s�"O�y�D��\��!��k۲i6֥�f�'p�'/�)�'2���j�L�&o��6��*/ZU0	�'���9���lE��#�jѸ^nYو���O4"~��U�`b�;ХL�c&P�(%OQN�<���
(M
��5C '�}��fJ�<ip���|��Ȳ�F]��U��M�}�<a�'��^���*���UU���1�ZD�<�� F�&} ����rw�����v��hO�|�� �W����㓠� ZP���� �S����]vb-i�� ����]�D�!�DMr����g�6��1HWI�%|!�DW�\,����W��p�i��'i!�Z?�|H��U�"�{�"L�h�!�DV�S�M�p�¡^]�Ca��K�!�D
�"�p��$����T �ў��'��y~�l�4P�fؐ��W�~<j[�.F��y`��hሹ���J�cNP!e�"�hO���)��A6B<�HN2d�$s�IK�N��g������U�uut`HS��..imB�J'D�����@�.$0� (�!B�0@�&D�(�G/	?�L�Q�.���ء��#D�,z���-F�\P��)�IZ�mʓ!�O��>ڙdb�)l��l� ��6�h��YM�L�B˘Lc�ˍ
f���ȓ`$đ��D*6+�݊��/���'�a~r"X� n�)st��f���1P��y��6^��Q�sc�0/�d�h���y���2��c�I��'��-�&
���y�A�=��qzpk� �0E�v��6��>��O��!ECTc�p����]�EӐ"O��y��G�/`�d����.�M��"O> ���ٱi	�pF��G*N���"O��at��+�����s>(��"O�"��CU�,��l%y�b�U�<�iL���8�����u}�𓵣ON�<	��=�|!�BV*6�XtH�J�'a�4�J�f��:@iԸF��\�����yb�3l�Q��"89��9Y��Y��y"�H80^�m��E1��f��=��)�O>�أbCY*ѓ�Ř� �n�Xc"OJX:�F�2_��=PB��
8�����"O*�1 ��+W�����@����!"O d[C�M<%�,�1,�`s杲�"O$�`%��X�⠊+�d�(�ɗ"O*8h���rh�1H�V��ꕋל|��D%§-�lQBsg��U��5�F`
8J6a�'B�	S���IAM�N�8b�L&""& k��0D�8!��
pp|����͒��q��l0D��x@~0�0�Ɍ&Q�5!�!-D��Ã�-�L�fn���&����/D��hE��@eSb.��K�<|��,D��##��>V�t�u��/^��f"*D��	ЅU12�BF�W��t��b(D�\Y$�݉,�z,����$�\R��&D��@�	G.>F�=@���
q�	/.B䉸J�V �Ҋ�@F�A9��Z��B�	v���*F�["68i6MK#4{����&?!��N�!�Lt�m��t��H��
v����D%ړ�����*����W�@�Mm`�����ğ��P�!,� ���h�\�!�C�}`��t�� j�P��\�X�!�٥
�$�"�hQ
kwnd*�'�0�!�0h��X���ө)jT�� 7~�!�dHF�N�͌'<e��b�!�nl�	��?E��˕�{d�c��ֿ>�2][`��)�yB`�`�q5hR�FL��q��ޗ�y��[?@��T�60qZ4��M2�y��3h�����&"&:����Q��yQ*���+q$R�cҍ���y��e>!3���8� U��y��
o�ШfD_�}�8 t�Q���D�<AO>E�T�۾;  $�W�0l6�S鑯�y
� |�)d��v���RPK�]R�P"O��ei6G���I�)\/pB�eiv"OB(
�H4d��}����2�8�j "O�{�J�4��\�fZ7.�:U""O�J�FW#f�J�E_�ZL�"OF����W+�����O2�b^�����%��|�����:قQJ�ܲ`Ϡ��So�r�<�αd��yR�)_��#�KW�<��O[�PQǭ#AAF�:U�Tm�<Y"J�T�cOOH�R���A�k�<��V��q��MR-<њ`I��<Y�
����J&�Q(O��!F�{�<9��	�Pq45�Q�(�R�ɤ�y�<��"G����B`�L�c*����z��hO�>���V�T)l�b���JE�|�����:D���0͖&�-��C�;]$��j�Zv	��mӼdAA#Z�t�ȓ2�����3G��7OA*;���H<�}�4)� ���V��vxX��ȓ7����g���|��I��Q�؆ȓQ���l�j=�FꋆZ����?a���~�&�K�In�8 pb؏&��q�Fbk�<q�F��;&IZ|�V�1��h�<9�j�u�$ܡ�&�Qޖ�D�[[�<��Ȍ4_��U8g�_:}�����V�<��ʑ)`����T�ʊb�"���K�<94��<�&�%ʞ�Bin5Ё�N�<�j��_�Hu�ч�$E�哆��J�'a��CO3�6Eѕ/�,zD=æ�ƥ�yrKXH��IB𩟛6�<;KR��y�H{��D�e뗄/.�� V5�y�׺�n�`�,�//0ݳҦ���yb�M__p��q@I':(2�����y�g�<	f�1r�hs��2A@�(�yBmA+��!�C�Z�pxPh>�yR��3qV-V���a��.�y�M ��y��$�#JI�ēg$F/�y�kW�V�b�@T�[2;k�" L���y��Z�1!��k
�1ؤ��N��y� ٣;�0����(��L����y2Z�<��l��FL�o����L��y��](%�Ӣ���<�� �9�y�/~��\3�0\�~�tM� �y�%� ҄ô��( F�e@�(�y�� �!h0�2�O%%��t�CL���y�Գg�� Ѥ,		&� �h# O��y�J�,qiH��.24\���BS��yo�>|ґxq�ŧ-�8��$�3�y�LP��ɩ3a͙"/2$�Dg<�y�A�17ό1��j�UZDO���y2j
�)�ث2�ޡ
z��V�ݏ�y"�?h ^��CoÏUg��a�H���y2�&P�DX#	y"�2c��y�Q�G��� ��+_�h�[!�Z��y��˜Y �Q�ǎ�PԆ���y����l���u��F�&I;1E�7�y�H���i���9ʨd�`�"�y�H�I������P-�>]c����y�M��?��#@�6�30���y�%]1>��ٺ��G�3��R �:�y"���B]��dD�|��)�D�ybDM�UT� V:|�la��P=�y��ƧC�2,y�
�u�<hZ����yҢ� v�͘�B�n����d%�y
� ���uX�[�����?[��Y�"O�������(��잉`���"O������<�a��^3e����"O���&��j�mSaC�����"O>���M�-�j����!]��5��"O�t����CH�����7y�v���"O���@�����G�ft��!"O��h�OHp-�%���ӿ/k|�S�"O m�ХF�}�࠲�_;��"Oj���kўEѶ���� �$���"O�dK�J�b�3A-�%$��be"O��"��fL���m�E:m:�"OT��F�Y \3����L��/��(��"O��ĥ �Oְ�H���N����4"Ox\�2Nѡ#/j]�ɓ��
� "OXC�\�<stuc6ʆ6�,Q��"O:��6%N;��C�T�ܴ��"OƄ�t���E�(���	*U���b"O��0 R4B��Mb���7"6�A3�"O6d��JU�T_(��F�LC�"O*A�P匽W�����!8�Y�E"O�\	�fV� ���1��� p"O�|�#��wh5�)�<�� a�"O�٠C�HzƲ�8��I&Hsh�#"O���u-7K���E��^(�`�"O�P4��7C��DP��6]>*uA�"O�uxT��`�2j�i����S�"O�X ���'Z�=�PI�!�pe�"O�dZA�G� 	(כ-Ѵ8��"O l�ō6�B�t��6w�zt��"O��"S ��(@���H�BT�7"O�<�"% H(���Ϛ<����s"O) �Q<�x��h]�+���#�"OڵY�J��`$�)
���$�"O� ��iX�T����V:�z �"O�āt
:}� ��F�
�a��"O���@î��q�
)5��w"Or����d����)ȫV��̰7"OVE�C�b���	V�R�"Or,�v�M����(Ob6��xb"O�4R�� � ����r�@�S"O֩�V*�N�J��7���g,�P�"O���7��_��yC ΁�m2�P"O�ڵ-��伻�Q&�@�"O���Z�o[�O�fbL�"OLK��,1R�A=VI�Y&"O�H�욈A&����C� B���"O�	c���?�Xpy��Ƌo���"O���e��ʝ��`�L4]�"OR|�p��,Jf",S��yښ�
G"O�pH��'��@�#�G�Ò!��"OxQ��[%Le�V"̔?��}K�"OR蹶蓖2;&�h����ܳ"O�@"����6� |r�aO�<�&ah$"O���W��;���J���e�
�!��]%I��[dNҨA0�%�(X!��,x{���l4TțF�=c�!�d�B�{�c��N8ۆ�A�c�!�dG^V)���X"U�\BWcS&f�!��S�;���0&���M��� I�!���8V�CҤ�.���R��14m!�d#U�&��� ��~�� �I�VM!�DS�G}2YI�a�]v��FLU�S/!��ԍ-_0���kH =��*�ۥp�!�� @���dE�Nj��q�◶J�pC�"O�u�Ȓ�D��cAʞ����"O���w.��Dj�L�T��s��Æ"O�����T�B�DS� Az�"O��	��$D �m�"jH5�!��"Ȏ�!�E�,-�P$�R�㺄2a"Of��wb$���׋�t��"O0���͒Co�p� ��*�^��"O�	��C��Bx�Qɴ�r�J"O^ݡ�F�@`v���՞e��)R"O�m��d�5G����� .�x��0"Oډ��*4�Z�%N�%��Y!�"O�H��#��dh�4��$�	��H�"O^p�M�|��j�A�]4h�"O�} �L;G:fݲ���+n$I�"O�U�A�>�	�B�F�c�Q�"O���^��)��`�M�Na�"Oʐ
�
�b��5�����(R"O�%Rw���y�\ih��O��]�"Or1�I��,{vEڔV�& ��"O,���^����<%h݋�"OnQ���)�>|����P;|�a$"O��b��E=p!���c��>pQ��"O��h4�ɲB)|�Y⍃�4T|�Ã"O`E�u��)X��eLQm'��{"OhX�,�r�����ߍ�nZt"OBM
�Lȴ�)�'ɒ3���#�"O���r���k�)P���E�N��D"O���
�7���d��-e���"O������s��Y�j�SF���"O�кq�M��V�ŏ6=�}����yP���TC�4��B��y$֓n��P�L]�$����&.���y��߲/����s�< Fq�栌��y���4`�8����
Xaq)���y���i]-�F�X?��Y����yR�A+;��"7�����i@��y�.кXv�C �N#��DJe��yb��%q��
%"��	�����yb�ސv
�U"��c�IP1�@ �y2ᙀ�v��M�]q�E!���yB
k�4��� (�홗��y2	ݖ
�(lX��6f1x�+�!�y�d�Y�(��o�-#��z7k ��y�G3�l�
�*,<�&%lO_2�yR@T^��{���'j�q�+Օ�y�b�%v�;���B�M+�yҠ_�8k��{�����@���y�d�YX����
�,��R���y2h�Fp�( s(�/���
��yb�A>��@�K K)��1$��?�y2ʔ�R6d3c	�IV�%�Z1�yB�?`xX���9J8�)�я_��y�]Ud���Q�F���ځL��y2��'��T	��ʐ'z��i@�՗�Py"A�R����@Όn{�8��@t�<y���>����#�J�<�I��ʟK�<1b��9?���z@$�008�qy��Mb�<��^!^��iK�J&<qtcT�<9��3BΎ�8�j�%n�؀+�`�u�<�c�
'Ғ� C-^�_���I2�Fo�<�mK�r�� ��9�~yQ��C�<)��7.\$���PT@@�%KAB�<1$Lj>�h�΍�\�\]p�.�u�<� d�ڦ�	W��,!N�GkR��"O���d�!H]��O �0M���"OLl(v���b�ĉ���3�"O2i�������gC�gV��"O�t�g��)Y�X�k#�l�.<JW"O��q0#M�A�$���GG�,��H��"O�9��-?��|�&��)7` Q�"O��u�J�"ě��# 3,-�"OԽ��YT��q�����7+Ό� "O����Ȏ�c X�AR�N:q<��ٷ"O0H��d��I|́��>"Nn9�r"O2�Q��[:!i��U=i.�	!�"ON����+�L���\���Ѕ"O*���X%���*���F���0"O=��l^�X�A �A��H�� �"O��r���#2���'�d䒀�A"OZip�Ə\T|��E��>@��s4"Ot���A�z��	��°ư�)u"OH ibݧer���V�ŋL���"O qp���/gt$�Dō(<��"O��c&G����1�X�T	jlئ"ON�z ��D< t� �
��R�"O0с�!{˨��� �	�~���"O�l�p�Ӽ}JXS�@�1�Y�"OZ]S1���6��4"/��b1"O�` �*�F�LkV��:�`�@�"O�a(�/�7��̒ܳ��H�"O��CHG�lt�#���"���H�"OФ��웑IO$�c�*�����"OR�	�
�g���9�
�)t��!�C"O�2� Jexڀ�c�Hc��y��"OBqz��ƄAC���Q��/���"O ���@
�uB���_��h(S�"O� ��P�K���`��h��4"O�$gB1��i���` �<��"O� ӌ���Ɇ�M>|�Z`se"O*���K�e$\���NE
E�p�y0"OZ;��H%UxMڵу:АXc�"O�-jՌ�%G�P ��@8<�8���"O\��1ϑaYM�@.X�R�H"Ot��g���Hyx�x���1>*��R"O�e�D�b�LM*m\�-��[��'q�'KdYh��W����R�(�*"�(�j�'8�0�1�Ζ'�4�z��fDBM��� �S�$��r��a���f�F�x�l�yR���Y����	^�Ơ��Ƣ=E���x�{��E)w���8�ZV)��g-ؽ����D|Y83� :w����?	�!�O?:�(��ʿs@�գ��s؞�l�_�ɒI�D���d�<qg���[���C�D��� ��<���兘�P�HC�8Y�N���>_�`�w�B�1gH�1����R��U�6T��B�I�l�4���
�B!"��2��	�fB�I�iP�03�&̈?A�C�"�8P$B�	/#�dQ96��|!�u��&+� B� <^<�̑�EP���.��C�I
+6�����\�D��a�;6��C䉤ue�d�,
A�l� �d�� ��B�	bM�
�����#e��dtB�	nb�[��C�4��,����~B�ɜ��h1&�2�8��G9(�:C�	���݂�D��<�Z��U7�B�I�h6�� �3&�1z�|��B�)� tEy�* �pK*hxMQdۘAkS"O<�Y���L͂�"DAg:I�"O\mS�'ɱ0U��ip��K|1�"O �A�Q�;^�ɠ�O WfT%a"O��1DHW�l�h�7���w��l93CH<�pɆ$<�(
S�J#}J���Mi�<I�%Y�����!z5�	���n�<Q0�ǔe��P-�P�Pao��FyB9O�L���iи)��\�Rj�7 �	�D!��!򄊪2x�q	�`�"�[Q��+��I�HO�>	�CM��@��׋4�P�k)D��:��	p:b��$�X�[����'D�b��
i��S��W�Q��`+e�1D����+)g V�C�c[�G���ySA/D���Ā8l��peL97nZ`��-D�\��g�_�e"w����я*D�$�"��%.�Hz���
~����,D��I���I���"T��	$ra��+D���!��%�l�D&E$����)D�p@���=븨)Q��4���
2D�8�C�H�/�L��$$�* �����,D��0���N��@�d 9`��� )�OO�aK3Đ�@�ft�p��pp����"O�`V^�P��N�?hT;"OZP�t�S�uE$�RR�>I0�\r"O�|@˚�=�d�k�PXâ"Ov�Y��)VT�k��Ԋ#��O��5��_ԄZ�ÑP(:$�b�&�|���㴔�s���]	N�K~���t~B�OV��6ǂI�*|{rܝj����w�⦙�'����<��'�.��G�	�S)�JcmH�{��ɚ�'��t�a�K52T�ۧ�4���7E%4��֋�-���j�[CS�-Ӵ�+D��X�A�`����ė�y���;1O�����'6ފA�Ȕ:`,b �Eo�-qX*�OF�I覥Fx��|Ή#)S�x��d�9K� @���ʿ��<)I�ȕ'fZ��s�D42�p�̞3t)�]*OVʓ�hO�Dnj�
����̝#��#4>Y�>�E���E����B����D5 �mp� �	�HO�܇��s�<uRi��"��1�)��d��	ӟ\��L<����#��e�Ҩ�A;� D�8	�ua�X��(X�0�Z��W�N���t�<Iߓ3$bC.ٖ)����
\L��R≽Z�^�{����rk�y��� EXB"<)ϓ=�Q���J64����T�_�isDyb�|b5I��X���+QN�*;Oa�r��y}"�'���E(��^a^P�C�g�Z�����c���q��(/j�Yb�/ٺ?F@B�	�Y_LxFM�;����eZ�w(�O���DJM������� ���͖T��`D��.ٝ),�]����8Rl���O���;�S�Oܘ��b�t%����I�ǌ5���D1,O*�)jZ/$�L8(�g!'n���|R�'��R�޺X���C�t�>�"�O�=E���	=�@(3$?�@@M7�yr̔r�\]B'�E.3i�'���D.��O�I3SI�]o�0�A<P��`V�If>��U���`Qb���c3��z��:�$%�S�'^�y�A9}AP�D��jF����/*ܪ���& x�D��*Y���J��"��*����8~a�ȓ y��]�d�b�ڲ��R�<��Ș:qh
d�V�������ȓ~^�q���Zi�BQ�c)v�h���S�? ��y���!���X�HNG�hY��"Oz1h����
�i�%P�a���qǒx��)��DB,�k��U�0yĄ�@��I��C�I�	�yrD���<J�y	��*;��C�I?ز�@�d���e�7��(��C�	�6i��  �Av�\��B�+�C�	�u48&��,�ܤ��,�f����d�<��4��Q��ߘuu��lGu�<�A⁲M�dx��k8T����u�'O�?q�N׎,�v���0�°�<D������F�.]�&���8��9D��:2��?MP&�k�@�z� L�w	+�Ov�'IR���,��A�a542H\�O%����S�)� X���&)p�Q�Tʆ �(#=	��T?��C�4�����%id���>�*O���$��egl`�I5u���ɚi�a~"bM�j��ǜ�)�R� &eąi������Р�y��8P��u�è�	lNn-� �O,�'%Q>���a!"dz��W!h�Pi���=�O���Kylq�6=��X���)MNv5D{��9OZii����C��p�`ٸC�.ӗ|�>����a{��1e�/I��"��x�	�<a	�nj<*���p`HI�p+G�7A�=�k�D QQ�N�V�2髆ꞗ8�p��
@�0�7��4Gu@P0N_�A?�iD"O,MP��ɂy�N��c�
�AZ5�@�'<������S�#.\�y�l	�"�*�+D� (� P*mZ�l���U�}���)D�P󢥄��! ��M���%D����(@�
m�ٛb�A4���$�N}"�i>�"֣��p�@ �7l�)`����#D��HU�E9`���#�*�e��H D�0`p��_��-	Y3|�@�2"O 9v+		�|#%d\�qBQ��5Oz��$;(*�$��
�' ���GUx�!򤘞��-1�#p���R��Z?bD!�䑃Z���cp��,�Z����!���M�L��%�tQ��Q�j".�!�DUdUx�7�_���t�Щ]*�!� 0J~� 󦉥F�Nh�a��M�!��OK���7�DX�I۠I	0�!�d�|��88r��@,hYT(� �!�ĝ�XwZ��e�I$+�����@�!���.3���,r���ȃ�O�!�@�2,�p7��{��T�q�
�!�3~G�䑐c��!A�F��.C�I�+M����R��A:iW��C�ID"��3,��jdMt�)�B��a�`� .6� C αk��C�ɇ.��iZa�Ù!���uP�.�C�	<	8q�N��kHܴKs�̢*R�C�ɥ:�@�J�P���Rf�I(w��B�	E���t�O"t�`A eDE�L/�B䉕1�e��C�\Z6�h�f��&��B䉮^�A5A����D��("RB�ɸ2д���(�&p�����^�]�<B�I�J�t�#�� ���i�G ��:B�ɍ Ԏ�a�E�!4��%�s bfC�I-k�*#J�7f��!y*Ʊr�PC�I�k�����-�_��Y���A-=�C�I�%s�̰�l��4F$`r��@<�LC�ɓ/���aW'V�F���
�� �!<C�	�F[<���H�,p
ԮӤg�C��;b����ԀÎ/�"p�R!ҞwM.B�)� �1됬[�I�����4�jPȂ"Oz�����? ��f�6t�f��u"O����/��T��8�&6J�cs"O8�)��ؑ
��H�"l��4���"OF�I�bW��Z���KI�$d��B"O�;�CC<etT���&�h���"OvX:��I�g�U�8�f"O�u*P�ǊAŲ�F0j�ɚw"O���j�)����G��k�"O$2R.���5f�7��	H�"OTt��L�Kݾ=�E"������p"Opy���G�45�a΀a{����"OY�L�*��0<P���$P�yǺ�8@�'�,y �a@)���K�%,f���	�'i�q��-@�c8 I��)%�z0Q
�'��5B]�R�0�����8��	�'I�lc�
��u���I@�B�'�0yałR�K'2D�!-8)�~I��'�� ��oY4�R8y�W� �j��'����⊤M��a�2#.��
�'�Č��hȥY�f|P�@������	�'�tjU	�U���2��p���'2����	&F|$˂�κXA�Ԙ�'����.�*�@U�V#�d���'������2ڶQ2e,4H\��'���4h��l$�PXp�6g�(��	�'�0{a̅
7a3�쟣UE ���'�Jp� ��Z�Hu���P�_�\�*�'[,�yA�Զ<�ڗ��Je��h�'���1�N�!�2@ 7�B����0�'Ř��~��x�bB�;8-n�1���O�<�4��#O�Z�q !ʳB�TS��AA�<�"�T	/��8�R�J�b���E�d�<�.ÿUD\hφ�E&f���O�\�<�4�<lxz)[��PI�x����a�<avd�x��U�@�8�ٰR�X�<yt�X�+�ʁ�v"�:qkH�Ȗ#�X�<!'�]�AŨE���ȣB!���l�<��k̀`������R�Vs m�g�<1��(P14,�F'��U.�i��#�v�<��Ž+,,���c��[�x�p��8�	5)Xu1�Sv"�hTֈ+��<�h�=o߾B�'5��� ���h�4���-�,��mz�!�������|�'iBp ��w��Z��F�C$p=��'��u@r�� ;hp�&gőf���'�����Fw8� y�" ���a�.�n�i{��>LO�x��2ָ���'(l@��c�#n�����	g�$T��'�$ɺ�g;�>��aD�S��IȎy����V��y�6�l�O@콉���=�HP�#�^�=���Z�'�Q0PB�. } �!Ղ*r6���"���O�x$�3?���L+;nD,�SJњ!�ʬ�b�~�<i�!/Nx��ʈv�$�"\�Wd�9�"�y����$T+(r�y��lN�|oq���,Raz���3�����ʖi?�a�:^�"�ʐʕ�<<u�S�D�<���٘mm����Y�g�zع7i^�g�p��G��K{��~�������̕�p�u2/LT�<��ˢ��b3'I~z��0ab�}l�<:��|r"I���$G�!\��p�
,'�Q��;%!�ܾ%��P{��?��t�M69����k����I%^�n�kS�Q3ye^���M�<C�	�k�
�a"'�2N>5���	��B�I��,�� #�	3R��xDF�6\�B�	�'5Xu��́���؃���#�B�I=��HP�����?�\�j��y
� :afL�=N2��ғ"W�?zn�p�"O�1�W�_�i�TA	"*[�]l��J1"O�a���!e��ų�$��F���"OXY�#NOhn��`hY�R�����"O:�Q���lM�§�l���r"O ip�3wג��� vf��"O�����Y�ڙ�Ƣ�-�.���"O�XRlN}�zqITa�0z����U"O|��d�J�F<
��Ӡ�4?�u�d�|ʹ>�q�=�}"�%�?P���{uA�'\����D�	R�<)�/^� ��Ơ�b�HS� �fU�Oj��OP&����E D���)+�PADF�{ m����E&H��U�Ϡp�Ci��W�*l�B�&J8X���l��=�a}�8�N��%=�	#	���O��FBЎ�t<�!��	Ir~�S��֘ �莬K\V A� ��B�ɽu�@uZ�錎�ƅbK6��Ld| W�T�\f���d�Ǩ���4�I�ڬq̃:F:
��"OY�w��>{�Fk�F"�I�#cQ�~����g��m�ΕZT�::�g��lx9�B͇	��Y�L�
aԅ�� qB0�aŗ 0>��2��e�z����B*Xfn!RCc���B�A&�'!�����!a��c��2y�(�����VT�z�LV~�}V/Z�2@�I�&55
QǪFs2Nba��_T!�̺x��;Sg�6)�pba��(rP�$K�1p
I�1�	$Jx�j�E��{��}
�T h����ě!�)���~�<9�.�R	p��4�tp��8B�������;L d�q��N�${��(�.�S
��Op,�-f��r�K3d� R�'rYt��+&�O���CX,]4t��cU�X��8�g��.�pts�BW4Fy�u�́~\���Ƿ�?i`��&_����AU�,�r��>1'���T	T����J�O�������r��x�c���g��0���F�A�'�:d��4١NG����)�;n�$b�ϺEÒ�O�L��˶ሣu��SÓ1�$*��L&:j[�;0K�9�ɠ ��!�W3�v�[���2�("�O8b���94M� YӠ� \tPQ㥮��
�2�g�;	ހ=�%��u<���C�t��ňwe�wx���$�
�,`Si�~[�-+g瘫F\,��j6s��ŸǅX�rt����D���}��
U��5����^����iX=D��{rK�U���ī�S	���4B�kaz�8�HB�l����FI�M%2�Fֈ�0�vNO=l��訔b1hgp� �؟�I�J��,4�����;����d�����ȴ`߈ih@j��t�]�,o> �%'�D��&I?x'03�� 3�byZ���v��=~+D�;O�蛇��]�B��(	�.�}�X�@�Z�Y*��wO�b��䓯�*�2��	=}�[�^>I��ja͉�o��H1��
-b��t�E�Ϊ�x�c˶>
D�Z�<��5@ݦV9�|�������� H��P�ez��K6=	D��.�>��"U��'Կ���ٺo*0�qEc�%xL���DW0��=���H�h-��j�;mI� �S�4�,jJ�O"
I��L"8ŢqAs�3r�����M�0�lZ5��g}r�C	H��8�#�]�T���ʾ��'��A�c̈́�\aQb��o���V�?����\�^��Ԃ�zq4��W��O�}��߈I-��7����<1�)_�4+��B䆐?Z��v"@?Q���-Fl����@�m&�G��'\ �S6$t�1ḼcU�� �CϺ�yR�/��:7`�M��tJF$���?���	)pب�ī-lO~Pi��٨��cU�W�Q>�K��'��� �]%>rb�@�P�	���)e�P��G���y�aےd���C�4Zd��茅�(O�P��![�e��#}����L8�R�.H�i#�
�i�<�S�X�`���x�Z(K |����T�K�\'�"~n� _���D��R">��B���B�I�]:��qc���C�
]�5���i�����%(��PazM�w��8:qkEq��8Xua��p>���Շ0�`c"�ݓ6��ܘbLs}��b����]�FB�->�~D�1	�Hy����X_;��<��/8�fl�aI9§2�6���"5�(R�Ϟ&c� q��X�8 Vl�sM��9� �? `E���Ke��9a�OX���OfI��L�W����7�r�X��E"O�!£��Y��&ꉍ��e�"�O�)���4WEb�ӓ�T��Ӯ�S��T
�l�;Ӵ���_�`d�B�:���U�I�@^A6�//p|@�s"O�y��)�L���BA��,3��2��e�ga_(�>� �C�.�t�QL�}�l!Z�F>D�� @E��a�!J�.e#��.j�4�׸iX>|�ڤm�ɧ����m�r߰���瀛/��+��K=�y�)�+ޜ%'!��PDd3R
����D�i�vH	ۓ~�T!P�5�!IЇ�E*)��J�d�Cפә*���уM�KF�`��I~�r��ǅXz�'	�j�0�ȓ8���dC�1z:�*�@�$�,Շ��ޠ���8z�,q���<r1E{��6�`�i0�DuXh��3�>ls��&ÊC䉡�$)�B��+�����Q�BZa�3*����!A�}}�!@.L�J��23E_�H�͉E�>D�aE�M[m�%Z�aZ4+d�0�z�걉0M�G�2P�ō:ay�&ܞ(�z�����lj����N��p=qc�f$���3��us����dM �x��Z�f����S-��xbl��PqKv���S�8EF�� �'��c� �;f��HHDʚ31��V����>OΑ�0���b[BEc�"OR 񢥖����qD��M���]��b����!4g�������<��
J;c:A��O�d�^-Jc��T�<�l3I�1��*JH�X��.//�\-���09=���DdM��ay�F�5	�M�!nɭWE�����5�p=I"Փkbx���(�,x��G��rm��:ABҿq�^�ru(���0?1�S%?p��gG׸Z�<�A�)Y,q�	��.��,s�Y0�ϐzqz����\�db�:��;+%�QUW��DAF}Rf(Q�T��B��6yY`[4��*\�f�閥��}rJP�W�7G�r��5Hv�@�W�<�Ec� �8�9�D��&�fm�"�I�<0*S J�BbO6}��)0kv�4�4-={�̲.â���K O�����K,Z�azr�����S"b�5X5|xᆊS��ķh�~РB���ēn�~����OjX�	�v�C�\�qty��O�%[�2����,J���SO���Vd�U�F�v��IAT*�F�
-(I<��hT�5jb8�D(��C�(�����h�h`�!E|���0~�`�cőUܧ5��:D��-h�=b��X6B�h�h��_�@�ݦO٪��Y���!(Q�%�ܭ c꛾fCRNb��p҈�	6���#��>E���Uc��hq�&� ]�5�����M�@ޖ/+Ь�o?h�)W�N�+�>`���|����'U�e�T��8�f��<�t�8�d�{�����H�R�+�1����V��%�#���$�����P)�d��@�ޙT�xZ�
O*�{V�A�A�܍�!�|�Vx��	�fA00D��x�'E�@e���x��D2�O'�@��ȓ��S�ׅ~}���6F�R"���'�*�����w�S�O�{ �8Ĭл�"t�t��'��l3!ė=�	Q%C�&�����'LD���^pH4D�)�D��'RY	�@J�W�>�Y�&M�%yb1��'d�W�=b��*�>�p�)��4D�,���L�Kh��(s	�%J:�� 2D��#'*˲P�
���ψ�D`ԙk$M0D�pҵ�H�F�d�7��gsNu�C�+D��EkT�2�(:�-�(�$�-D�<�G%��1�{Ў�0dP��閎+D�0)C$�]ݴ1H��@�?��df�"D��	�),ra,=
�j�qܨ�n#D�Hا�O�t�hQ��%_(��i��� D� �斚"duzM�8��0{��-D�0����q�4�pe�)|�f��I!�Z?*$\����N�0�%��?#!���y�F��eL�x 0xJ3Ƒ��Py�c�{V4��3�ӻ�Ą��Z��y�@K����@�-X�e�(�6�ybD�as8�0� Ӧ)�l�X5�P��y2�G*:���b�])�PȚ�o
�y�E�)�T)Q�V",�H�����y�mA�`tr�JA6#3f�3����y�G��]xQ�Wò��K��y�i�'.p�)�`زR\��Ӣh�=�y
� �)Ag� 56��V��4#\Q"O��D$J/	|������W$�""O�%��8)<�DB��X�{�"O��a*�e�DD���Y�!�d"Ot3�$U!k\A�`�#�6U�"O�-����?&I��O��s�-C�"O2$��"�����c��DN\��W"O���b��|_����_� t�ȓgb�؂B��-OX�۶����<���0� >6z�A���&of8�ȓ(�j����ٞ�iJ�L􆰅ȓF.�81�A7&NL�y���#�^0�ȓFW\�3
� )�'įt�"8�ȓ(�[�f«s�Is�Ì?|6����FYh��_,�r{WKБ?�ȓF��`�Fe Sd2��ҫӥ��1�ȓ7LL�%�j@:V�]fu�!�ȓ)�4j��ɕP��!f�S�oE��Fo�(;�JD8�]IëG:RBe�ȓm�"�����5�ƕ��MQ�r����ȓ98��"L�+qV���.���^=��q�\i���N����V"�؅ȓp�-3���E�Ryu`�\�D�ȓ{��r��5-�a� �l��݇ȓV	�-#�V�WJ:��Ca�x/���"ޖ�����R�z�+4e
�x'px�ȓkZ����&Q/��'CQ�x�`!��iBuaS��U�&y;��"o%TԆ�=΄�(Z�3$+���5I�`��Gd��ؒ%��e���1r�j���fW�3�k�);��� y�������.H��IA��ʇ :�ȓN$r��# )P�^��w�Q}Nĝ�ȓs��Œ�B�*����L'vu�ȓe�t#����$	��gB�s�Z��ȓ�=j�CX F�}�w��e(`܄ȓ!�$��&�D�X?̩@�X5��E��27&��Mq��I�BP2uB8�ȓE�rL�W�S�r�B�J�6�"u�ȓv�$��D�
�Nz�N�<����h�%�\�h1u ��Z�L��ȓb����փXG��P-F�����>�X2�ʔ�����䔍� ��y��UZv-,l�ܴ u�� n�C�	?v`X��"
J�"@��G�sg�O� sT�̥��F;�d�Q�P���OP'lE�"O�4{6�'��Js�G�%����2egt%%����<!��8m�>��GI�?����T�<�@�L?�AJ@������ِ�p��c�%V���dݟLK�ᗅ}h�� Ώ�$�az�KB?>�h@���R?��K� m����M�<��a��n�<�K�Ex8�,|��d�7j����<�W�5l�����D+�'j�|� ��!o�����J(X�0T�ȓ*9���1��%ej��5�S����b�,&��'�:�я𙟘AUf�S0��BaY' d�1�)D��J�
͍B�, �+��c�b	�V�+���8��	�r��|�*��+G�0g��3����i��0=� %��x�t ��J3hS%��0
a��'ՒXAD>D�,�$�@_`<D�Qb(g�����?�I(f����I�#I�Q?}@���6\��1�G��Dt$xqf:D��b ���FS
��U�N�D�;�aث��bL>1��8�gy�/�1W�@�ғ�R�J���)����y"!	�����R�ިL~�I�$�-�M�`=XXH��ןx������E�4 �ʞ+r�!�� BpZ�a�7i�� 7f@��ֈY�"O,T:%���rmtLpP�[�$?�AJ�"O���0`O�D���Ä�,,�(4Y�"O�� ���tX��3��tĶ�k�"O�ty�
ǬW��pSa�r���T"Ov0�w�O/�bAQ$���x����"Od<p�X<���� ?fRH�t"O���[N�f��Q�U� N����"O���Zcu���Q�Z:?RP�Q"O"Ē&��MX�yf��jLx#P"O@�{7H��{�.T�0�GP&�-�"O�4*R-�z���g��
Dp	3"O&<��G.I���5Fo<���"O��Ql݌o�V\�AŖ�@��"O��,X��^��*� $̄�"O��"�9w; |QwjB�= �Qq"O����$ص6�v�q��F�mpt"O<����%bb��iG��	qF"O> Q�	JBѴ����C1\
�!rt"O�-(RLG�_ЦEa�CMQ�j�C�"O�!�f��	A���h&z�X 7"O�\�A���k���Hvr���k�<���%M�	�kI�Y��I�Wy�<	�M�3~�0c�=����v�<)�*�5q+Z!��B���@\H�<a�� :��s%�	n�P�[��RE�<9�W�m�B�z#�� %�t$Ii�<	V@��*�G�vo��K���d�<��e�1k��+�ǂ[�`�9�x?A��ؙ>�'�����Ӳ�5���'|���O�P%�i1����n�1�����w�l�AED,c���`s茝
��gdB�8J>4j��*6��̉P�ϱzC, ����O\�BS�,��>Q�Z�y�ؘ�ڸCp���G�
k��W��MY� �4B��	WH�4�O؎%8e`�/h�D�(���\�NM����Q ��V�T
`����IT�0<y�CE�<D S�T3Q� �ŅڝE.����4ZS��ԥ�.�Z��[ e��@�shA�5��x��aK�R$}�`��f4�aR���x�"�H>�f����@�f���?�����i���h0+Oi��DX@�J1�����p��O����ޠn48�j�i���E�ɭ��=�f�_��G�h^���5f"Yb �a1�
P �
���Yi�5���Y&��@@*sT�����,O8���σ�&w
1`"���Y3�$��=a�A2QGA�<
2n ��#lڴp'#�s�1�u�\�d�!�F�	q>�U�ag��^{��56O��
��b���q��4E�ջV�S��8����m��OJ�O1F)���I�~���j�x�4Hr�z9|�i�'ȵD2��7��A<i�C��c��@� ��4,���V�
�N$���K�3P¸�[� b��l۰���(3UlK�|zVe܋%�
L��D0��������a����SŜ
q]p�Gfi���ED��6,�����:rfd9�����YFF���/s_r�?�=K�l���14��u ԁ1H���?1����Yv� �M�bj<c?A�C��'�T��%3[R9��OZua���_�R8�u`��<At���8L"�P:*:�GʘFъ�ۃ��!p"��h��dV��[DW�!��e�� !��Q�Э�E.��tw����0]��A�;^���y''�A؞����C-0�����K�FI�f"�OU�gꂑ7���X�.ĈCg�����Ȩ�`׼/�!���z��Ğ?T&`9�K52�������?K��j��$ҧ�0�`RC=P@���R蔙itvфȓ	��q����#BA��@lڞ1'a����u�)���q��G#Tq����/MvKq  D�4 $%M5:�r� �#�y�4س㣟����$���'m���slI�4�&x��O.j ���@��!�_�2���`
U A)� �� �@˗1D�D��o��. B�pP�]3X
$��o/�A��l��+-%F#|�Rʗ�2��AS󈇷����A/S�<qB��عٴ�\�9~�qÓJ 'v�%��i��H���O?�$VV�őf�K�����l!��G�-�ΐQ�NJ�)�0w�:	���̫tX�| e���0=� p(#oT!نyx��>d�Εz��'��]z��<����臰e�f�ks�J�3�~�	�.Hc�<�ÂO7T����((zP% ���Z�'mڹ��b�6W���E�dj�
P��C#F�"��#G��-�yb��_"X��.^�&k��¦h��M����i2���K>E�ܴl�zh&Տq��p ]�<���ȓv��jB�$~vBE0�S�ZL�@�'���5� S؞@P � �z��򤝗K�A�e4D��ٰ��9�6 �o["f蚕��5D��1[e��C�G3?�@m��0D�X�-J'�>,+Vl�6�*%Z�*2D�$�� @��W��Fa1iԇ6ړZKj8� @Ю���CC��<rw��3g�ۜb�: �"O���"	ئ2� �sv ]=B�|A��	,��yc��:e�듟h���K�B���v G�����^*�!��3�uٱ��4�,5Bѥo�v�A?,>����F[$EN�9��J�f$�s��	:��\"�D�4�х�	�/�(iE���F~<1��l˭{���G��'u(���B�iz�Ԇ�T1@%� @[o:�Y�f�Hl��=Is�Q�<ވ����TlÉ�T���)�L�ٱ�.e�&�� N��yB��!u��q!Cͽ�DPP"Ɣ%2-2ǌܔ=��Ca�OfXa��Y�|q�F�7�zq!eF,uM����3D�@Y$�8M�h�7gſMA����l�D72i�#D$|N̻�d��<���	!�F �'��V�L�2�X_������2H��bv�c!�e!���s6p5I0H�i�D���F�V���h.��f���@�G�H`f��R�B<pׄ1�r�B=sߐ��f	�Sv<�$F6��;]��a�j�z�s���i�b�>��n�+�������P�e���1� ��H���UOR����X&je$��o�<�ċ&�gy�G�Q'��D�Byz�z ���yb� L�`����j��S�z���2��4����a�0Ÿ�HN�,�`y�KQ

4���(m�v���B˿pz��[i�X �	�}�䬱S�3��'���	���C`n	�t��� �L
7$^x�Y��)Hnx��	�&0(�S4�{�6�)�@��fPF�x�.��M��xҠ����Jݖz�2#~R�)I�(M�\��dM 1<v��Dx�'(>9��Eȝ.��}.u��AK�Ά(P
�|��F3|�εIcΞ5&�n�'�.�G�,O�)��\T#B�W	Ѣ.���Q�3O��y���w�9�J�"~�Bf�ekֽ�PȀ)/�B�g
ʦ�!�̍;��I2�49Ó�)a�M�6b�,}l>�R�><�V-�<Z��b�8�vmE<[��	�~��qy��5���[ �«9G����U�"0L_�y�PIj�Ň	"�):�h�1E�YI`J�d(<A�kP=Q�uaS�E:@.<�#1b�|�'�U�C�]7��^��@	�80�F�iRÊ*rF��f"Oz�� � ��hؗ��*B]�1�uZ� �C�EqO�>��$ƛ ����X{v��d3D�,��
'bT:���Xl�R�Y�3D���ë�S�61Y�g�+@�8�0D�� R�w\f���ۗ�D\{V�,D�4a O�31r����-b�^9�g9D�h�ӅK,o�R��^�Zx�B`8D�Dr4,�%60�_�3-7�*D�l:W�;;4��i��\�u������5D���$�Uv���.I>
��)1D�T"���*7��h�I�vؑ��.D������$#B
�p���;��¥� D��Y݃Kzn�@IјF��}#v-*D�P�f��4��A�w�O�l��1���6D�RX�SN`��`��2�#2D�dq�a���AR�I�2��H��0D�PЅ�E�:8pC�$=�i�( D��֧Z�1MdPɐ�5\�|P��d?D������ʽQ�ĕ_�FH;
;D���I^!w���b��QV�9 �;D�H�'�Ð6��q+Y�z� �"7D�$�犼l~iq�V�nr(��"'D�� �j��çLZ:�DjUm�\�d"OH���M�@DIEV��$��"O��"b�l�X#�h
�gk`�Ґ"Olh+F���;����C�Ms�@1�"O��(�
�[�ex�/K�ph���"OdI����	Yg���qH�c��዁"O�M�e�O;`�Vm���19�8S�"O�\ڃ�G� ��Q�f*�w/��i"O��TM�:=��"�	L�2j�cW"O^�҅���J3��đQ��P�1"Oj0c7�[l�X�0�Ȝ?{"�Ъp"Odq�ԧs�8x�&K�\	�H�u"O\S�/P�7m4LACE�*��]b"O�8���5k�(�
ㄝ!@���"O�y��N�W��$��T�uB���"O�����S�����nJ37
,M�'"O��`t+��uܴ#vmn�vh��"O���g# �x�4tѷG�%N�V�S�"O�Bǀ|G����GQ/XrVݸ�"O���	�F�����C�'tB=��"O �s	R/0p1�Vi��ykK�1:�>�z��A��n����w�)���+���e��]��R&^� ��8,��\�΂H�)ڧ��Md&ӫK6����38�po�Ag0�ҡ�|��i٥U��5s�D�$_�@���,$��YR��s≫YI<�����<�íW3�����fy�Z�%�4��ˍ��xםK�>��Qx�F�rW���NWjy�L�4�Y�+\�ݨ��7m�?+�1f.	m��y�G����c砕�FAN�rק���DW�͸N��J�*�6�>Y�r�q$ވC��)t� l[览��^w�t��tdĦ@�pٓ䃞Z�<�Cdj��IFDhT(׽I?���O��"}��O��x�)ݐ	��8��U�P?��T�G��	��/[/\����H���O*H��e\%�P�1�١I[H�2���l_�!X�Auy��0�ɇ<g�$�S	$��P��?�,�X��	��1�`�d>��a��ʦ��"!��0|�eE'H��Ր�M�S�ʩ*◢\W�u���ͦ��a��U�@�Zç��5++�#!��7�D�j%�b ��O�9�`�y�J�F��a���iGv����;Ъ�A�ޔ/RX;tD�+K�8�k���D�I�r�O�>�ӵ[p�e��7U�Ȩ�ψ�&rJY�G�X<|[��y�a2�4��<��-�ƁړEW~���@�N)��8�M\(=Xvq���'�����K*
2��j�[�HB���'�Ԥ����.��\�RnW�A����	�'ĔY� !�@�΀HR"�:2��S�'S�J2�ܴG� �,��"�|��'Yl$������m���Z�4V���'�r0�WDӬAxD�KB[�L��'���g��&��)��$�!�.�C�'�6a懙�(t( ьB�'@ܻ�'�"8`3�6��3�n�b���h�'��ؠ�k^*v�K'�,[L\���'�d��gW	Ԓ�8��Z�Op�� �'C������P�zЙť\�EP4A��'u�m��$�#NRjp"�N�A+�D�'�����\�i����ģ=�
 "�'z�K�X	��}��#�m(��h�'[XP��l�'m^���s���aX����'*��Go�Q�3�܇Z�|���'
��	c�!u�ԭh��E���'Q�P��Ё&(ֈ�a�Mcb���'��:6o�"$F5�#�Tw��DX	�'ix`A���Ё�3@�vܢ|��'<���o�2J��Tr#�،\<$��'�t�hQ-F�$#H$�b�[:���'�x찃G��X�8�'a��
��':f��E��1�$1&e�>�rt��'��|���Ιu��ɫ5I��#����'�p���Hn\8��٥,;\x��� ��o�B�؄ 7�l>�-V"O�QQ����h��e����I=�|�"O�틀L��q�P��1��1#D}��"Ov|�EG�>�di��
p' ��"O�,q��PV��,��hE�$��"O���I%{E* &! p	���f"O>-��jV�u�́Pf�˯�Di�"OJ�p#�m*��¦%p򞉚�"O�y�S��P�x�K��1�ʉ��"O.�B�� {�AC�F:�ءRc"O!aa�2�6U��lYe�R%bu"O�p%�9�p�Kí�5��|H�"O4�h��κU]d�;�l���b�#"O�MY��K�&��u�^���ܺ1"O2	gg�,Ю]J�K�c� Ur�"O��$��< ��A���t��	�'W^�ӰJ��q��5�&��q#���'�,�3�Ё_6^��拎�8e&ٹ	�'ް��M��vb,ͰE�E;)`ب!�'�ЕZ7��M�th��(
.m �'��I�2�ͭ�y�C52x�`�	�'�~��0?3�8��&��\�Aj�'=vt+��*O�L���ߌf*֤i�'*�t a,ظa�
Pp�oZM�Y!�'��!��K�h�~P�4���>�89�'�E�g
�VY�	c���#|eD���'�v��foE#"�D�����
9:D#�'�R� E̗�y�9IѠ��f٨
�'�,��s���c��У��|�[�'�F�k1�I1f�B���"յ��${	�'���(Bۃt���j�A��e�,���'�E�dm֖���Ç�enB�`�'�`���$�	_�iu���y���4:u�)	p���o����ʂ�y�D�D�� c���{����d���y�F/Q~ e;����k���/H�yB�E i���	��I\�^E[Dɖ�y�/�}T�t*���k���Z��y`�*&$�]�d�˧�R� r�͝�yr*	�)��hC-&a<�9�����y�ŋ�nvH���/����j�"Ƃ�y��E�I ��f�*~0�3�Y2�ybKT`S�᷍S�C$�m9��7�y�	G�pp� ��2sSt��dW*�y�,���x2��e�Π�WiĀ�y2��{H�#��0�6�����'h��sk��%��!���KΨe��'�\� ᎑=2}LARc�I�Eę��'��ӱ��+yx8T"͜E�^��	�'?�E)0�05�̸��\�:����'K��8k�Y�P�_�����'�� 3F �4E��"�[W@���'_
!i!�>f���>�����'��� �Y�&��`�nP�8���S�'��'H�q���~��,8	�'�>I���a�a �ۘ}(�l��'�����L�46!�!�	��@M����'�,�!`�'^��m�&זk{�`��'�d�0c�*����6��c��s�''� �@J�**&Y�$�M<a��Mi�'��0P*��W�(�	#��#����'��}bD䥬�-vY��NV�<����K�@�"�D 
�Z�x�(�|�<10��"m�h8R��X
?���#Z|�<� H}!��"_@�� ����� "O`|���
Dm!!\��<��
�'���`���;#b=P�mʴ	<��'�������1Trf\�"(3	˖�Q
�'7"�#�j���xYd�.rXP�y�'���[��*O���^�{$���'��|3��C$_��a�ėfdT��'Ɔ,0��EP���`G4Ű���'��I�6oMg>���+�>�e!�'k��P�V�I�zt��K�
���
�'`����)Bp�)Z��xH6"O�(���f�80`�(Y�~
�"OB�hF��A����X>H�Рw"O���N$����$n�:j�X�f"Oj��$d5NiN���-M4aox�(�"O�V��~Ta��, �d��&"O����)�p��4�*v}�9"O��D��U���	$MK�_c~�+�"Od<��l��ܲ�I϶t#,�"O*��B�BU������R	�8�"O蔂��Q��h�SE��9��r@"OnM��ۖx/*XK�d��~W�0�"Oġ;7g��'�pD�tM��X I5"Ot裄'*��K��ϯ;L�S"O��1����̋���K�(`��"On��pD�H�������!?�����"O�a�"�S�D��O�A�D"O�h���(Z�}���h��s"O&%�#� yP&���Ƿ,����v"OB	q��h��`:'����0�"O@�ʀ�_
_�� �AKȩ,t�a%"O@�B%eӽdԐ<�DI��Et
��B"O�9��<�Ȥ��&�:wτi/!��N�A�<�i�CT!RN�Y��-_�!��B&[,A�t��N["���[�s�!�D�;	 �rc��Dƙ!�A�!��ԋ[����i�=f�.uX4�V�7!��<zrc��J,"A�>�!򄒭s�����k�DhE&��	t!�I�ODj�*�9fތ`{�c7W[!�Ĝ:z5���q	��+��D��lޖtE!�DZ�E��,k��خ��$�A,E �Py�L�+����'�
�Gfv���@��yr�ޚ����/W�9Q��ӕ�y���L�N��D�f��F���y�/ݱ5�j ��b��,,m3e�^�y�+�k�����*
Ai��O'�yr�$��9)� �������)���yB���v:~�r@u�I��.��y2猢5Lz��(�;U��B��\�y�л,h����G�}Ir4��K��yb�El7ȅ�����kvb�s�n��yR��g���W�H?A�%�U� �y�F\�<���nҕ	��)�,���yB��.x;�4��nT�8����sS4�y���7WN�J�F@/2	�4h�)s�!�>d�t,�Q��k�� ���.?!�d�.Z��=��h;43P�IU�
=!��A�$L	���8CD���6'��	8!���pu�}��(��gB��S���N�!�$O�.�p�x���U��!�/_��!�$(J^\,C��0ۼ|���0qO!��5Ƥ�A#K%]�t�:ը�-!�d�.}ڵG��+%����%�9A!�� �4�3�B@��]�򃁝X�-J'"O�-S��=_Ж�A�̈́�k���o0D�p�G���P�wY�m�<��Wi;D�XIQGO�U���jg`�L
va�V-D��r�ᜌL0� A!��:3�d骑m,D�pb�b�T`�رQJK3u29�,D�H��	S�(�4���!��U�hɐq�*D�PcqI��(d���|�T��Q4D��z�ɐ/;	$�Yt��#qDx�X6F0D���&���1HsC
94*p2��/D��C���M@��zr���: � �+D�����iڔ��v)Њz4�q�&O,D�4H��P�2��rGDJ�x��)D����MK>6��	�g�;r�ڑ���2D��0mS�|�3����nܔ���/D�@��H�NU���.9�q��g;D���C��zP�V�Ԟ@�*l�;D�L��̂\UdىbaN. �5(Q#<D�4x�j�)���b�:z�ِ�l;D�$��؈H �d+�`�lՂ��cC:D�|#Ƃ[f���̛�B�U-;D�<(��G=bz�Q��'r�B�*�:D�����6 ���0�/�s��Ѱc,D�t#W���](\��dV�,��[�$>D�����S0:�,}�� �;��ԛ�0D���e,�9 Z&�XwEB�)�t�V�.D�#Gt>��P�]�l�a�/D��Xb���gu� �寜;"�(��."D�0�'��8g>��u@5P���I��>D���)N��#�)#����3�'D�p)@MQ%�RĨ��"j�$qTF#D�P�qEҴGj*��k��o��ś�J D����gI�v�:��5��+����A4D�x���--�:Qkf3a��@��1D�ȸS��*VÌu���»<s~����;D�\q���S��P��tv")0��8D�4��J7>u���	�be
ţ�8D�x���w�u@�mJ�9���7D�D�g�W!xUh����|��9�Ĝi�<��*(����L+	a&Ă���\�<Y�'�:έ`�ͤZ��tZ�#�X�<��L:��ň���$�Y���S�<����0(h�H�E�1��bU�<�K��.����OS�Fh��R�<���,E�XQ��ǈ�p���pI�f�<9�H	C��e��0�BJ�Id�<y�H÷v��	iƋ��I k�]�<��և&�Q`q�Q�*�:�hD��t�<Q��až���k��x`aڱ�Dl�<i�gZ�s�逡���m�4�!���h�<17�Q   �P   �	  �    �  �&  q.  �4  �:  NA  �G  �M  ,T  nZ  �`  �f  <m  �s  �y  ��   `� u�	����Zv)C�'ll\�0Kz+⟈mڄc� 特m`�DB�6%p� �f�q�䐻"�m�|Mi+��.�c`e�	��IuJ܅b�"I�;0�4���'Y8��J��}��1c��)U����	��l%ʡ�bC� b�Ԛ�@�����B&� 9� ���X`�-��H���9���=vr�,��$�3b��4�WEXB�b5���1���G��z�*�4yir���?A��?A�⌽�g�X���`�r)X�������?��й0��F[�(�I)es2���O���؊\����6&���� T(�����O�ʓ����O���'	���O����tI���R�~��AY�8�O�牐�>�+�&�)������۴0�(��y��,���I<Y�D���ⓤ9>i�1ӑe��D������I���������q��?�P�wB���Q� �$/��5R��'~�6O��m��4כ��'=�6�	�y�޴`����'��3�
��K���{#��<���*�� �G�?}� �Ϊ'�0�W���LF�IX0�����@��m-m}[��i��6��1����u�?���lY�Ik^��5�<"�J�A��;:Ȕ7mP�K�V�i@DN�Y6��PA�,�D�tk>E�mn��MG�i���Y���` �="�5�j����B �ŷ!��7���ec�4v� ˃G�)�j��!ǔ(���@�֏�V�K� AO��Y�*M
g@x��pB��\��	�´i#^7͎Цu��\�Q�qR�,� zR����G(3~M"��ڵ��p���_|�,�I=^5��u	�"s��31��
d<|���U��sA6y��N�i����9=�6][U����2��'���'	���O����K s�I��'xD@�P �-nY�T��N��]�R�:Q"O�mA"�\�VƁ!�Ə�7��eB�"O����96��3R��-��%��"O���#ȁ1�И�F)��D��S"O��Jq΁�.?�	�R�7/��,	A"Of���Aif��Aj���j!;F��fU��~Z���<�n-�4i��	��y�5��c�<!v�@�U��y���G�]t�Ѣ�v�<�f�3Y4��*ʢK�H�!ʞt�<I�͝�3Ft(��͠q|�02�I|�<g"A�������ic�c�t�<	�mS�f�(�n�>�h�AR�����3�S�O��lٱG�;C"�,�B�:.�ʧ"O���a�ލ+�D*4��:�F��q"O(�#�>�:��R�� ���6"O0|�D�K�%���*�M&��"O�峕�O?CMh4�LZO_��z"O�ep'��8j�XaP4+�.2T��X�<�r�.�O(�LN �0�"A�C�(��"O&	���Rvސ�AaJ�M��%�V"Op8��K�3s��
0��[�Lpu"O����MD�ufp��Å0����4"OB�a�m�d�x��з��G��<y��X�!��������J�x�2O
$��3#A�O�ʓ�?����t��$0�npʂM+s��!C ���2㟿e�X��B�6�t�)��I�F�J:c�M=���� :B�rL�%�z�:e"��C,!s�,�z/�� T�ɏ@�F���O�4oZϟ@K2�žM`�V;dI�Y�3GSy"�'��	S�OO�Ɣ;� �S0	�K.Y; #��1!�$e�����.\����G*s� `P�f�Ox�D
ߦMr���ß���sy���y�2O�T 􎐁CJ���Ba�>�XQ��R�ϳ>qO>�ف� �3ܑ�&�^�K��i)��;?1*Ƨn���"|R�O�F����N�9�H@�ľ����q�j�D�O�c>��N'bhR�Z�o�J<�r$4���O^�����j�
tV�na
3���a�џ�Q���L�WMJ,{Şb��c���$2K(S�O���	k�,@@Y�~ni�%�Ҩ";<B�)M�Х+0��\�>��"��:-�B�I,}c��zu"��c��|`V�P��C�I�=��d�h^�+J�]��I!�C�	��lE�$�"V���#���
��C�	����0�˟.I�Z�ASKT(��KeJ}�Ć�d����P��*O&6�8׍v�p7�?����	<kD��"�[;����W�c��C��=
kN=xw�=T$*�j2�Y;s%\��Ӣ�O�̇�I	|%P�8�@
02��M�r'];��Ǳ*5��h��'eI��a�h�vr�'�`6-1�D�=o�`�$?�a#A�B���z���o¤�Q���OV��?���?���>׆$�'�%^��s!��� ����ۖ4���艟rb��*s�4�G8�l9��O�^b50��1eڽ�Tgۢ �8��0��	f��1.����Ox���'�򚟘�� �Ca(�!��7	rte��A%�d�Oz����T���A֫M1�89��+]2�O�O��(�Ȏ}��S�B�_������'��	$O��2ڴ�?�����iI4��Dд2O4�
���(_�0RR?���D�O\��c��Sb�z����(�T>E�Ow�(�`�f��s�k��+�\�X�OaRT�Lw�-r�Î֨��tô�F�v�t����2 L����O��lک�H���)�7<��ѳah�"X�r#���XB�ɖ$1��X"h��("Mh��[=?�N�?1��ӆ!�B%'��q�Hd��E~��8lZ���'��D�a�X�$�O��$�<	�����	���RV*Y�������8.:���\5T�N�(���)BS�	8�䜁�*4:AF�2i%~��0j���	 |�� i]�!�1��ORP1-�4_N�a���U���C�'k�6��O 0�*�O c>��?9�%Q�+� �	� X&xC�j����d0�S�O)X�V��>o �b�d]?���I.O��m��M�I>�O��	=vp	��K�d:Jx ���}�z�*L��M����?9���|2�O�B�pE��f�% ��Hb�ٽM��]����Vm�ق��N�џ�\c	J3�$Ul����J��!�X��0�F�jm��s���iږ����%5s��Gy"'�u�+��
F�d�I���0����?�b�i��R�@�	Qy��?��TI���V9`��Y��*��6�OJ��"��7<�	1��	�(/���'�6��OUm�ҟ��|�	�LF�H�v����d�B<��Xj�J׏� I�ȓ�T]��n���GC�^���䊵� ��9��=;�F�"p�ȓt��gC+7��� �[�Qoj��ȓ~�^%��(�,(��S5PB���o��P*S)��Hf�
!�XR�F{�'D�̨��9��^ }Ŝ��A*��wR���"O�ܛ���O²`��7m4��c"Oȡ�r2-lI#�oÎ+���R "O>$���B��0q��Z�`�� :"O�T�0`�Q?�=�Fni�X��"O�Ճ�i3L����-�>��d���'a��8���7$� �#CҬJ�R�8&`F�n&���Exybe+I4%���u����o>~,�B�͇~onA����P�4��8�BL+e)�1 �UY`��� ��ȓ$^p@{�;w;΅`������ȓK�^�A�S(M)0p�ە9�n9�'^�X;�)%I�de��8�$�7g_�-��A6�Y�3H�	8T�zj�
 �Ą�`�	(���:+L�" �!�D��ȓb�ڶ@�p�-Ąe4:���c�R@#rG�.��сD�ԥd�Ņ�	5��	4��Ȁ�@�Rs�� �U?�B�	8"<R��3\_�1�6�Wt��B�I	P|��VI�C�8����U�TB�B�I&�<��%o���G���a�nB��0JJ�$8�"	(�[�O�2x �B�3%"�s�����ѵ&]ZȞ�=��}�O�:ܸ��j�&�Xs��=>&�B�'r���B��J_4E3���0�&;�'�
�����p���pKԺ ����'� ���ΰs{�e��l�;i~��'14�X�+��g��C@�-��c
�'��)y�$�m�(�C�R㖝��X�||Fx���I/\��,�Aj��5�u�U�8�C�I�\�Xb��ω(�^5Ps�S�J[�C�	Pl�I�튦a�Hkmѯ}�&B�	4>�`�1v`چ/��D�P�mPdC�IjwvM۴�ʈ�&Q����&C�j�*��5N57g�{"LY n6˓R+"a�����(c�*K�*�"��C�)� ��ZĮ	�&4S�n�*4���@"O�9Z���24ҵ@$��*+�P�0"O"0kA�&?74�Kc��.t��"OP�� a5^�[��H�]Ӗ����',hP�'j�d�s��%^L��u+��4��'�hr4EY<E� Eo�bO��3�'�H��I�l#�'�^A~���'�FpE��7�|��D!#?���'8�U�ax��U�cF?��T��'����C��am��2��Q�v>����d��Q?�h�����(���L��aZ�!.D���d!��U{��sd�L�fy��K�9D��y�����t�4��"6��1cS%6D���e@�#"�U*�HM�6�~���6D��B��!�heHV"�a�
YR��'D�a�L�_�& �flG;-1�D�P��Oz-��)�'!L(��_<F��)6`�',ҖDZ�'���DրE$�"�D��:�a�'��|�P���_��,He([�<�2�[=|%�DR�e*��k��TW�<���d�]��f��ea�T�<�T�Y"8�
U�e׶O�\5x���Ry��+�p>1 -C���ʆ�ʵ��)f]N�<��+���D�χj��i�2�DH�<��اs��12EoT!,q�3��G�<)�e�,t�j�m��aB���&X�<�5�A	/���:��8AU6��⪉Wx�H`E��8��_�6�Z#\?��;A�4D��	q��$��)'��FƆ��e3D��c%�8K�Ƚ�g��,�z�"1D���v��U����C
';Uh4�� 0D���D���1�l���Ʈt�*p�Ec D����.	-gNb��P�)��SEG*ړVK�@D�$/�F��4w
�}���G���y���;>��a#�W	n�s����yr� �Fd)�R�/Pت�j6 I0�y��P�v� 
���O��e����yB�Д6��p n4L��1["�P�y�� b��q4-E�/�xҪ���?��F�h�����Ո�π20 �o�@���"�g%D�`�ƥ�� ��r�mK�F��o$D���*Q�PR���$��MJ@�J3�"D�(
��##t0�kG*�B��>D�����Do6��7�@�?jr(�A<D� ��+ʸ	��7��d���<���C8��A��ݍC(� Z'�� aB�\"�(8D�$X �M\C��Q�̡U��SrG"D� ��K4�R\�sb��{ي0A%�!D��z���n����
l�p�>D��C�!��erz}���_�B���R��:�O$-� �O� RF%���>��0.�9;v
(�#"O������A���P��a�s�"OP��d�_8J��d"�E k��K�"O����!O�/Lxsu��t���`�"O|D��%R
)pDE�$�
lO��	`"O�A�� H�m���F֌6�ځ21�	�o��~��F�I�(M@�2_�LҒ��B�<Q������0���^��� ���v�<�p��>e@ܨ�B�� :�*]�ȓ|0�y+D��~���4H��n���>	�Z$�+{�t�X���
|$�ȓ.`>�gb� � �R*Ɖ3�9�Ʌ٘#<E��N�1��lPj��r�$q�S�	�!�$\,E�ʱ�d&�����!T�
�!�� ��)��!<Bp⇭��-�>�y�"O.���cǚ2>e��͉�cw@��"O�hQ�G?+!���E�*`�S6"OVm+���6Ծ�3��"�yQ��  '�O�)��Mê2~<��E���M�"O�͑WG�d���u�I�a��9��"O����V�M8M�D�4/�@��"O�]13(�)$���AE	H,2���"O6�@a�"y�biI�N��Щ��'�.T�'~�<��U���{�e�-u�\�y�'f�mz5咽O�~D�fH�0��T��'3�m�S䖰W+��*�.!�&�s�'�t!�@%�z�ąkENCJ�
�';~� bɇ(+���ڙ����
�'Ǣ���gslr�˴'N�ڪ�+��DW�Q?�#�,ȋEg&�2�:yq k(D�|T��q���b����{	*D�$�F�(I�y*G ��:~�(b�+D�LZ���#�"t��E �)Lp)��H*D���dI�l�lE��\(W��8*�"+D� �ٝ{���4�A6�Y���Of F�)�'f^��q¢]>n�j��s�RU�����'c�mK��[���#�M�TD�x�'����'U�Y|E�@zkt8��'��3��Qp��07�P(h4u��'�.4�R��J��C+X%xdB���'�L,yk x�8-�d
e�l+O�C�'�h�����13�}��Aèl�#
�'⁓D�G�H.�� $nzǮ<�	�'�su�1Y����y���	�'@���T�O!P��52�]�v�\Hx�'�j�%���%��!�R�&eff})�������Aք�=���s��{���ȓc��A����3��`{Q��!���ȓ&c�Yk0 ��~B0��Wc��,@�ȓ[?��b	*Mو��c��SU@���cm���IB%��{`c�\T&q�ȓp��ㄭԃ^�@u{�"K?=��mD{B������8tI[�P�jy���^��"�rE"O�Xs7�[6&�i���'ͺxK"O�L��`��NÚ���P�j�"Oa�tm¾$��Ac��A{G���"O<��-�F�D̊�&ۜ��ɛf"O4P@#�$�UI��V���e���'�Dݻ���@CX���m_�� sA"/�B�ȓN0��+��J��8� M���Մ�$��r� F6T(t��,9
q��fۘ���ԈCm��HO�x�@�ȓsLLр�kW�$�Ƹ� W$?�n��ȓ�h��OY�U(�=Y�/�[��ї'�\S�I��	V�?f1ir�� ʡ��	#(�S�V)H=�1�d�^��܅ȓx�x(BC�CY Vjb��a�A��m���#��>E��4qvO٦El�Ɇ�I�:,��H@�Bu�-�s@]�k�����h:��*Yx�!CS!28}R�M �C�I Y;��H��͹K5��!E 9
�C��0l���g�.�n�PsF,	�vC䉞rD<1�j�2T�Ҵ!�&6B�ɡ	e�m�VIR=�:ܲp�K�C䉪y���於��P�ǐ�_)�H���0�z$���;
����rb�D�ȓ~�"h�"¿?�8( 'řg���ȓd���� !#y�4m�� L+�@���S�? ��R���M����FBWY����"O*\���A�p)��^��L�q"O,<�W-P�w_
m����t�2�$�'*������S5k����FR8����%(s�8�ȓxo@���_�3�H���i��B��Q�ȓY��:P�T	Et�[Wk�� ��ȓ<	�IS���<�����r�P��ȓ?�� �e��]��,�g M�!2N���9`iy�͜	�6�i�C�76h,�'�ڹ �g��E`c�!&��y�g����5�ȓ>��=����/5�TŘ���m�2��ȓr09� ����X�Ɗ�3�\ȅ�%�\5��D�-'�:!�l��ȓ]=�@P���xJF�[�N�?2���I�M��ɹ_ܦ9PV�j~�5�vHɖBwB��* ,SN�k~��e��/C#B䉦a�by�Ff�C�Iس��')��C�ɤ;�u���N=���s�� �C�	�z=ҙA�˗<Z|j��F,�6chC�ɩM����D%�16V)���9A���=a���S�O�`Ʉ)34���6�( ��'�H㗩ֳf@<�h4�
|�L�
�'n�5���T�'��l�@�^$yT�p�'TT�a̙6A�[Ã�;k+�� �'^rQ��h�lHZ ��a����	�'����HT����R��L�K�x���#v�Dx��	$5'4̹!��
*�`p�C�U8B�	r��A�
X&��]�+,,\
B��M���ޑj��=�Ph@>P��B�	
}�2	��{g����C
63ĪB�Ɂs�vL�g��,2��v�y�B�I�8��|B���2E�T�̒xc>��=1H���b�J?9H�x�w��06�CqN%%Z6<a��	Uy��'���'DN�ӣj�����o�9Ai�Qb󟮝K2H ?p���d(D!Z�t����!D=Ե��^-r��I׭\7cd��r�C�� �&mE�H�]&�����-T�2����I�f���O�b>I�����.^0D��΍�>5�xKSξ<��wu�aҏ�
aE�LCc�}�j���	����ѩe�H=���jP�5���W	9���!|�^E��ҟ���d����Z��'�j�R��C4���G!Q6����'E<j���P��R7�DO���T>��|b�N�md:]8�L� svJ��2���<Q� �D��d��߸�Z��I�>q\��A��h!1�X2 M�d;!R�'��)�	:?A!ˈ�!�z�D��:	Z�����H�<��FL�JI$�*Q�	 �e�P�B�'��"7K^�!��+PB_9���䥎��?)���?�3hÔ#?�r��?)���?�����d�%�����B��rp�_K��������Ò41�)�4�<Fx����Y/����< B����d����':z��8N��i͟��DK�%(d�����I�`��)5?Q!X������?ٜOp�Ԩ���,w��u�5	[:@=�U��'�f����2A�i�NO):^Ȝ��0A���Sٟh�'a��@�鈶2�2����A%*-@1&�9
�L�(��'�b�'s��h�������'q��Pa��;\��rM�^]���B��%)P4�ǅ��X�F�'�h� ����=y#��q\z�@�y��V쟁�� cs�*,O��+�'oy��/� � E����]��@�P�'����3ڧO=
���	�;��ZD&͚K��	�'��X����x²uZ� �!HD�I,O��)�Ir�:�~䥟�p7H�	j���s'��L_>��@"O��`�$&��Ex��T�bkz�Iu"O�SPo��8�<0��F�=}6nYX�"OTX�dI�:g����8º���"Ov�҂L����+�dĪ�۳$"O�hr��/~T���.f��t���D�+q���O6z�:�ٯ[&]���V�E�\9b�''$H)����a`ˍ�6�b\�	�'�P$p c5\�J����6qd=`	��� ��5Ђb��Qx��PY�EV"OЬ�ѭ�$}��5�2�.{�6�!4"O����)j�0u�!@A�28\P�@�΢�O��}�A�f��D�I�Jȶ�C���ZF��>��kB `�|5+@W�Z؂8��	��5�&���A<Х�gf΢44t��(��5�wL��MC���#�(u��ńȓR-��b�'@ a�;��>)�h��ȓXX�����V7q��EM�W��<�I2Q@���d
�E�R��/'T2P�lZ!��9v�䃵L� N������%�!���~���K�w�ʤ+_�!�$97vbPKa�� �8�	�m�!�K��q�����%2A��џ,hf���M��?�O�� *�[�@�$��ӏY�]��K��^�H�Q���?���\�B�˦	Ir�d���ITY�6=�2���L�O�Ș#W�ޗ3������7a]v�I�+� c�"L�1aU����!��127���4�b�LK%x��##��O�#|���Վq���CS�ӔAI��c�\�<�� ��M�EM�JZZx���.OZ��=XB8�9'CE
��D�#V���Οؖ'�O���.�P�0���rT�Y"�Q�Pׄ��:�|%��C�-Y�,yx#��[Rn��?�4�ēA�8b>A���Ԏ.�hdq�6z�y��(?��O��q#�>��y2DJ�@��{4E�41��Z��ֻ�65[㓟p�I���.}Rk/���ck�8hUƆ�n��t�!-^�C�ti�I��a�'��>�	KG0�C"�$dߔ$�ƀ̋aHx�dD>}�"}�`	��I�����pE�-3сv\��s��A'Ę���I2�N�*R���F���cb���6�N��놫�?Q�(@��v�$ɷr��V���.��B}ތ����)�$����)��$��c��sQ�?����?A^HQp�2Ad�x0��{��I�/�ҧ�9OhT���*�&�5H^�ʶ��`�T�⮃�to"T�'*�mJ�O��x��)�r��cR*D�;1��AIɸy��@C?��MN~ʟ�dSq��$@+V�9!ꈁ}�i��8N�2�_؟x�uD�<u2�)���A�R>��2D�.D��)ai��q]��h�
(��lm��4$��٪���O��4E���x��E V��k��^�Jh�&T��$�tG{��	{���g�H(�C�0P�d���"O�%�P#�\�d��SD����
E"O�#��JV�-�d�3{f-a�"O��k�#�/���"ʆ~eP���"On9�W�M����!/�5\v�4"O4A*I-+n��b���"O���៫(�h�3-:c���(�"O�L�d�9Ȁ�5+K�6"O\Б���<k�0���+ި���0s"O4�	�Y.Yt��kC��#R�0�"O^�JtM��`@ ��d͎�	�"OXh�i�>P98��ad�/\T��"O���Z�I������,{��D�dZe)«^���=�FN��<X�v!V�,��}�gꍋ	"y�QL�sͺ%"�֬k���8�C���<��*V	&��쀑=J�ٙ�K�O�J����۶_�&\
�� E���1�0I�|1���îF<�Y��J�P˷l�(�$���t�6h ��j�>i�dqQ�%�=[O�m�tc�7x��B�	X�lL{�	�<��@�K�G�hB䉍:G�H #�Fֈ���l�2�C�ɼV�
�%����9�L�Xp�C�	/M�0�AB�F�݈U:�+$-�B�;R�L���-����"��+vB�	� 	���h�1B�����x��C��qc�� �B�m'P�J��^,;ΚC�ɫTl�IQ#b�.f_��#���bC�����yPe�~ �0+g(X$�ZC�Iu���h�P7(����ɿt�B�	.7Ťd�!�ǖ������E�I?�B�I�x�Ɲ��"#A���ڱe�8{!B�)� xys�w@�����
��#"O\�z��?i��	vLQ�|�~���"O���'ď$���K�7A�:��`"O���`J%z��S��;]|�x"Ob��Q�K�y��H���7�<��""O���`bB/Q2�)BW��7�H�2"O�P�*�T|���ӮH��Ss"Oh��q�W��p�u��bD 2�"O�y�ai�4��"	�7C�}Z"O ���˒+-�ry*RF�#8��%"O8M��y��\ �ZEs"O����;O̘a�K�$5�U�"O�vH �����	��q�� S	!�F�"�Tepօ�!�&�yQ!�q�!�D�6@^)a2�ܻh�"�)��NL�!�d�F��ѱ�I�)�N�P W h�!��/�la� [�XЬE���0q�!��
t���&�lDR�b�2�!�$V�(G�pC疿u-�}�5O�}�!�d�h�ˤh� L�x8�߄�!�d�!UfV��C�^�&���)����!���*l¤��2|���h[�8�!�V�S��(7!ގES�@��gOi!�ݽr��)$�XC��ArM̞Z�!�d7D%P&�E� ���P��ս-�!�d�Jl���K�C�,��3Gو�!�<q�,أ�~�<P�fV9Uk!�D\#Z��hfA� +����μ^g!�߾J	X�AчH|�� @*[��!�$[�z���E��dj��xц�t�!�ΪU�\��&!��ze�4�ckB?�!��	T"��p�䕑:�v�jBj���!�d��d5��hM�'�q8�+^*�!�	�}�d�0���N����7��}�!�d�@2@���ڷ���D��&�!��\��H��
�J�f��	�%�!��=~F<<q�ʕjmde�I�6�!��&2���h��7&V/'q���"O�!-%�Дӵđ�c>Q�
�'��ժU�է_�� �fU7����'T�8Pe��`2�tI �)b�p��'����G�3J��Y���R��<��'�4���#�	GT!@�(��X��'���H� \9Q��ǡ��mR���'���`�Q �B�ҡ,�h2(tc�'��<�$�X3Fm�l �È0�R5��'���(F��r�NN�QV�@�	�'G�At̏/o�0���-xC��H�'(���`啪*U��PR��*#��A	�'$dɱN�"T�4PP��H-j- ���'����/7��<j�ɂ�`H*x�'v�����Ύd$����)c���'��]H�BP�@>���й`8樒
�'Y�HX���C����)X�h��'�L�����T�A��}:�I��'�)Z�	_���Q[�ɍ�|��|+�'^d��'�1_FE��Oc,d��
�'��1��Ї�x�S挐'!�
�'�$�CBDR G�PE�0h�
�d$z�'�ƥ���]���E�;m�~ػ	�'X�ܓ�k�:i'���`���;N�1��';�J5'D;k���p��.��h��'�^��Rh�3#��ʑ��,��
�'o��'ˣd��P�Q^4<�s	��� ���K�Gft|2�K���"O���a�����bg¢ ؈�"Or`9W"�5�z����>��r'"OB ��Ԑh3̨*2���T�)"O�I9f$��
��qri�+��`"O�!�(S3
�r�����T�8�Ys"O<���g��X�0�`�*�*OXH��`�\��:�g6@��P
�'Vr�fk�/=e��ҕ�?�z
�'��Xq2$V�zش2rD�=�<̺�'.p����9}���4L��.��9!�'�=@fI��yAoܘ&�ތs�'����B%��0�=4�|<��'��D��� 2�u�� (�fE��'�XU��b	����Y��B�ꈡ��'B@d�G��;JF���ĉ�j���'��Y�Fl@-��QP � ~��<��'��<�u���4@�)ҥg�h�h�'�,�sB�U0��$��g;�A�'�ju��B��BPY3ˀJ�.���'�����H;?	H5��BH�>7(h��'��u+�J�K�=F[(:��y�'0�$�LZ�`ܚ,X�X;
�'r6��L�L ��)!�S0[.�q�ʓy�xą��,���B�!������3��I�<�X���f��&i�ȓ] d@��������j�*C�ćȓ	*^�b��F�;
 ����ц�� ��I�T�%�d��MÚ����LU��հ0@�|�0��5j����N��H� �4܀l���'^�6y�ȓh����,į;^V�����\��fe�����I���G�	�3Q]�ȓ0(f��q�9,���:�냭D�"	���}c	A�E*����lH�l� ���pXe����~U�Iz`#��>�ȓH�F�`ҿ���I��׭q��ԅ����j��ѝn� S�.N#�Z�ȓM* �ЫVÜ�&Ό������gm�4���`ü%F�݄f���ȓC��ʀi�"ڠ��	Z=	�e��tڤ1��c�N��)sΚ>&��	�ȓ^m��h�0t�����>~����|�h������Y���̷GNP���:8�h�\�p�6���5r��ȓwĠx��kN�S�9�B�'x�"Q��D�Q�#�*ihuu�[�JH�ȓn���yB�VF���DL�v0��ȓ@��L��:/*���� ��E�� H%�b��4r�H�Q�1#q��ȓN�X�s�>�0a)&�FLj]��Z-�xi�\�Q�v�*Ba_�L����ȓy����>X^�j�疳>� ��*��r)�.�Yt��M�x��v��(��dݏ9:=@�=h/�a����`�uꉘo�0ĠF���q�ȓ.6Vv�7]6p��t&�A'�܄�K�B}�"L*%��SEHN�E^�Ʉ�M�\m@��2�h�&��S8΄��}m�!���"��L��G�7̴��#
���!+}��m;g�^2��ȓ?Y =÷ ��#�
\�ၙT�Z!��y�dيG��/]����_�R5x �ȓdF�ծ��r͘#kQ[�j���S�? �P�,��JEN����(\Ș0f"O2�:c�IYB(�e�q��٫Q"O�A�f�?	�B�Y�bNd�"�;P"O.X+�d�(�vDrrˈ?+��U��"O�z���<~͂ܨ� �>����"O��B��B��\�4NZ�~�V�qd"Oݚcn�X��5	b�>޾�2f"O��L�"/Ў�r�j�2����"O��``F48��BQ�W�^,�6"O ��&�ր+ D%�"���x��mP"O�y��F?q�\Հ	]�()"O��&�^ 8��m#'ϑ�Z��"O��k3+؅n�*u�EG.2��1�"O�(�k���O��1�zR�"O ����΋h�<K��m�Aq�"Oz)���)T��I+��=p<l��"O�9 ˀ+���b`i�%��"O�=IG��H�������W.Yr�"O
iQ��ÈyD�suA�RQZ�e"Of��Q-��a�(�Z�/�?k��$��"O���
�;��a�`Q�=�����"Ob�d,� b�tq�J�G|xU��"Obq���юd�$Dqīyu���"O�	�'Bۡ*�4ܻ/
 r�̊�"O��R�߷$�����o��qzن"OT��"^'HlH���Ƭm��ca"OV$� �"H`���"�_�f:�"u"O�9�6�.B�Z �eKGd-�"Oh�2����T����<;E�Xq"O�+��զ\�Υ��H�o�L��"O<�AVGq0�5���W�|b5��"OH<���#�X+dgYx8P��"O6 ��J��n�&`��[?��#�"O���o_��Q���{/�)��"O�4z ��Z���ҧ�����AC�"O�� S�=� 䂲�D2�j��"O�1�"��O6�(�bϟr�N$�7"Om���0����_� p`�S"O� p�O
Fr���U(�1Z`�x�'"O�����"R��xg� ]"���"O�p�@N�X�*-�pe�~o�Ty�"O��Q`��^rr�i!D�0fz��7"O�U�1���l%��آ��eZH<��"ONdB��ҜnojU@�W7F�L��"O��ؤ�G咐� �zͩȎ�y�Ɔ�S\ �##N@;��`h�A �y�� B"Ver�ڶfۄAJ@"��yB �%F�h��PŖe��X�K��y���E�Pԙ���,� j��
��y�H�q �ؗ.X� 0q3#���yBNθ7��H�%��`��x�U��y��� N����͙4by|���%F(�yr�(K`�}�6ȃZj��H���yBh�0�M���5T�V�P�L�6�y�M
�dnБsC�M��U۱���y�>_�D��t�@��P�ƫݙ�y�g��>}8�!ɞ5<5|�21+V���'~��Ȁ������!h�,�K>)�!
�}:d-��B>��rmd�<� ��>M�I*A��K=_�,��'�~		F�Ր7tQ�c�
;\x� ��'���l�+N�<PZ���%g��'l���$�T�IP#�gѶ��
�'\YT&�$c�T���Pv��`
�'9�Q�/��r��4 �ȣ=�<�
��� &Dq�hףdz�2�!��+ژH@�"On	&�M�-h�u!�4��,�"Ovɣ2M�1��;�g��m���B"Or��B�ڣP~��ކv�P��"O��"
�>�`�O	�vfҨ�"O � q_�3'�4��-�r��9Qw"Od�D�PF�d���앻
wLi�""O��m�m'�$�0# ^��x�"O�U��4E84�c cɐ- ��8�"O�1�1��C���Z!�ݜ@�\�q"O��ǬśX�V����9u���v"O���P�T�] \����6�:��"OP�q"+�-lf���g6��4��"O��Xd�3[�Ȝqvb�p�q�"Oм�oR�X��I���*|hx�"O~A�*�@��D�.�."��""O�u�mί����UǍ	"��c"O���2�D�K��yӰ��].D�g"OԨa6ȁ�K8����c�B�4"O*в+\�C%xqs�dǸ�""O>T�Ҍ	)ܼ���]�N_j���"O
�#���n$�9���1��X0"O����V�Wh6D�@�T�#"O�����E�`l��C�� �/!�	V�Q���7��1#�!��XC!��0+�̰��`!��b����!��_&q�Fف���uk:I�g�Z;4G!�$͕=�$��ĄnV"\QԦ�$e�!򄝺3�FDy�m�"HK*,i �V�!�$� -��V�^�eWJI[$��#�!�DZ�fƎ��-� T� 4�W�޼/!��4l�MK�E�$�b!���I�@�!�d��eh�q�5~>(��E���!�^�)����D�2V>�P��M�%�!��a�����D�x���7�!���a��,L�!ihI�n�c!��ÏE�Pt`�HвL�h��j�#v)!��d��@5L�^[���`Wc�!�$ˉW8��p����nEt5���Y`�!�D�~�ԱQ,ڰp�m@7����!���	_� v�+wOH�q��Ѧ&�!�O>�Z8k���B�)zaKF�$�!��(ꅬ�(<P-)��Ȑ�' �%��>�𼛓`V�p��h��'�\1�@U�<^U���ѳY�l@��'i��R�?8�UA M�q��'ɠ�UǘYq��HVAͭ[t���'�p�xe.S�d��x����Rj�x	�'.V�H�(�(0�i�¯C�]��'K"�A��0Y��!�bD2u��%��'�� �V��!Jޒ��4�CAV��#�'l�C�O�"��T�a��-��4�
�'���1Td^T
��c�Q� ���	�'j� �w*Н c�N���%n�}�<���jdL���J��i�͋R�<�A ̀=��!#��[�`R1���m�<9p%Ԁ���������H�e�Zu�<9B�!����6��wi��&čO�<9�/�{#Pa �Q$�wJ�<�g�E1M�`���$U�ЉF�IG�<v-3��А �P��%:Q�VC�<�(��fuR9�wF�9zD�Q���M]�<����F@0�a�@�2Y �I�C��X�<�� ��v��"#�)-%̨�LF�<� @�Pq��7D� p7��Fv�1�"O���'h
^<{0� i�t��"O8�"�"	(k?�Y ���6$�!�"O���ϐ9~�� �ַ2�^��"O����Q4 �8��Ņϸ���0"O�x0G�̹}���%��Q� ��U"O���lQ&8�F��@���t��"O$$��IK�7�,���@�NY�"O�Y�V�[6~�Se�^����k�"O �Uh(������@,F�<-�u"OU3$j��W���Ĥ�=s1P"O2}ZƆѥfGָ��O#bh��A"O@Hz�+P�p��-[�͆5W�aju"O~��f�����	G"�f�@�b"O��[�#�!L،8��2r�`a`�"O�����Jt����HŁ��4"OΈ���Wv��[�
 &��Җ"OD�sJ��%���T���dX\K"Oj��%Z�9�V�Ď^B=("O��؇���(�;�MT�kG�h"O�� ޘ+V�����C�D� x	�"O �x��9U��`Ze	3�8X�"O$s3O"Р5�4k2'�H�"Ot�:୊�O�����i����(�"OL(�2۝]������W��()�"O�͓E`��?�fL�7cܑi���j�"O�����>���85�m�"O�H�
1{�N0y#�P�*��5"Ob�S��>hO���C�p<Q�"O���PÙ0f�m
�J
9�4r�"O��k�C�%&�����/�t�ñ"O�,cv-݆�H��'EMV��AIw"O�#�)�6�&��s)�==�;�"Ol�#n�&"�z�k�h0O�Z�*�"O���6��5�L0I2�I�.�XHV"O�	��B��Q�(��3-��|�u#�"Od�z)�t�5y5#�9�`���"O�p��*�,4#1�
1z�� Z�"Ort��V�&�*��/��t�"O20��׎57�x;t�¯ij�e��"O��Ĥ��mƲ��4�	g����"Ore���+%y@8#@��;\���"O�H�-@�F���oҠj���G"O����$[R���ΜR}����"O:D%��{XD �3�S�Vξ\J"O�P��O<1M��#��2G(�(i�"O�M��� H�V�z�eG7	^�X�"O0�S�'�y+���W�
nL�b"O.̋W(�7o �#�*�,EQ~���"O� �)�n�}��#� i�X�#�"O�arGM'�����,�h���)�"O����*�8�����8f�P"OP��T ��j����a(��2���2�"O�(���]��谛��E�8�t�c"OB5�P�Z"!�^i��'�]�x���"O���5��k��,�v	�g�.4��"O8 �KBM�(��"�S%I���5"O.����M�n1"	ۑ ��$Y0"O��@sM;��<���L:$��"O�Ԙ���]�@��Cd,��"O��ˢ��
%;D���G ���:�"O����Y-'����g�-j�DM�"O��y��[:�.u��޴j�"O|9�[�f�*�srJT�"�[�"O� �`c��A& }��������C"O\��3g�3e�\([��X7Vh��j&"O�K��Rx%45��acT hv"O6e��̛(
� ÈU��"O��j�Ë�\z�`'H�m��Y�e"O51�I�4N�%�l9M��1�""ODT2�#����Ӡ=j�(4�S*O9��ʇ+�T[�FpM2�'HI;���J�t�1eŔ4���'�0\�6B:6��T�!fa�B��?DjZ]+�'�*��=	fJ�$y�`B䉾3���B�,�2anE��S�|��B�ɰ2p��W�
�M���QCаT��B��5>pj�⡯���d0G�"��B�ɺo�|2�G �@'6X�B�	�Ni���'V�.������A2ԚB��62�>� �R��P��#F.pPB�I�)I�\2�-�0�4����=J�\C�	/E<m�-�]]J�P��?k�B�I���}23��P��y���ʒ&pC�ɑD�VaM�Ll�������P� B�	�_�p1��F8�x�apmQ�z�BC�I�C��@��
�0h,nAGL�&C�I	CNMX�@�\|�p戕j�C�	�[��	IEBޯ6� ,@
W _:�B�	0k�
�gl�#!O�MT
�~��B�ɧmd��cH�?f��i��װ}֜C�	�<(8��앎c��쩓���RB�:h:+�='QV$��ՋQ{��P�'k,�c�H"`	F���O�4�̼y�'��	4$�:��H������ޒ�y�`͡[���Q�	{hp�X�B��y��A=v����ٹteĨ�uI��yB��M|�05�]Ѧ������y�M�Rw��� ��%��[�GP��ȓ-@���B(�l�8�0��g�rh��V��Թ �p�)��ȉ]ӌ��ȓd�D���\:�B�3fo�)�ȓl�v�HcIW�WvQ	U [�qr��P}dU�'��4X�zy2�I*����'�,�k��
lt%��_v�����!�h���PU���ŇU�VM��,P,Ms�W&�&������i��.���gg�duI�Ro�t� ��ȓt�KǢ�4"J:(�0��e���ȓ]]v���h��t��@�t�n���D�4L���0��Y�2��D��W�r(1��?��9�j�\Q�Ą� �@�[T(��)̰�B͝�b�fY��nB�����-U�@��OC5$H���Bې$�c(Ӗd�����
3K`m��'�"TP��^l���Z�-	l3�m��v'�#�n �VM��N�1K�,�ȓw�i3��ME�.�2�K
u?J�ȓl�.���@R�C�d�8�K�K�
Q�ȓ??H�)2��t�*��bD���,��ȓq�@B&D9��p(�L��6<Շȓ-? �{V� ^�Ni��'//�F%�����`��S�ipv�!�ì��%��ih`<Z�N�6`�r�G�V4|l����X���������FC;&��5�=�#�w���%��5X�$���f�	�-�,	����FȰ&��5qC�I�}d$T���H�.Z\|��76�$C�I'X�֔�l5#(�E�!Y�C�)� �ZQ�<��a�v��%*p!�"O8T"B��q�� :�.A�~!Vp�"O^���ɖ[>�+��R�;9(LrQ"O��S�̓�T1��t,
_+xd��"Ot���	� ܢ�%;.6��"O�0x`��"��A!a��M��52E"Oƽ"�ߴ#���a��)�����"O.Ԫ��ݵK�p9Vb�z�]�W"OfqX&ʣP�bL����WbA��"O�D�w*�%P:���O�Z,Q�"O@��� )O�mH��pF�S�"O�M�AdX��I3�P�H_���6"O0D1Ɠ�}J���g�>hOV���"O����14�XY�2�T�*6|���"O`��ꁻ{D��X Y�:#��H�"O&�I�uԬD12h�<�)A1"O��B\?,����W�I2"OEر"�12�j!��>#��V"Oq�L˹@Z�뵯��:L<A�"O:Ta�G��39j|�c B���ʈd*!�D�q|�+�$���J�.�+�!�?N~a��V��%�����!�d��5y��1AI�(M2ɓ�|~!�d�4��䧓�$��AzW�*�!�d����aXtc�x�hp��CP1!�$L�&�����^29^9ӧ�լ>1!���	-��H㮔y.���wh�%!���
d�(D0�/S)� Y��8R�!�Ѷ>�}z1��
Y�( V�)r�!�,�.�je'J�f�¼��DVV�!�DO&^h��s�O�jP�h31m^6xZ!��1L@��N�I<�x���C�x!�Ď'za�#�N�#CXP��!J!m!��/�J=�Gb��N���#��Ο]l!���|,����;�D�82jɐ@l!�d,�ݩ[!"� d�U7H�|���'wB��*�ޕ��A�8ʥ�'C(0�!��c���#��4��(��'�~X��zL���L#.rpy�'-xxr�2e��A(�o'\�F|�
�'�P@�#�̂q�JDi�)	d"O 1�ˑ�v�J��\��
��"O���nO���a2���s	�q�"O�����_֒eA�� g$*�Xb"Oܠ�
X�c������E~���`"O a1�ڋ0F8q�e]�>d©b"O�-��
�,9���%EU;G^�)G"O �cS�*P��e��M�%�T�"O��S��f;I[c��hm���"O�<�"�Z��U��FA�pÆ�r�"O�l˷+26:Yw+O�\\f5p�"O|u��^�gN\�9�꓉wʵ�%"O:�CD��#������$Ev���e"Ot�Caڀ2>�usq�1);����"O�)E@��JC����p��8�"O08J È��pPU���R�5T"O�M:IG�b?2�:a�]�f����"O�1s���W,��U�
-�H��3"O.LP��%XC�\y�IY� �M�"O6@�g%�Y�jܨ�����D��"OdyZDe� |����/�xI:,P�"O�$�����
���Α#���X�"Oz��@��î���2V�2 �&"O�	�#� Z6"ǋ��I~|�ѓ"O� N��>'�=`Ԭ�Yz��z�"O��b�mF I����TA>~u�@95"O�`�WCW���xtIĊ���"Ol+w�ˤA4}�Gԟ]�~���"O�ꖩ~i��#Bgkq8�0�"O�Y9���H�V���P�@`
P�U"O����J�_ � X�Ꞙ2T���c"O�8�(�NZج��,̽��pu"O���,)z�.�@��X9:� A��"O�ܨQ`њ+0x)�r�[�D��exA"Ot��`N�T69���2*�"Obp"�oH @�AiCmC�h���[�"Op�h��'YW.�k�k���Q"Oz\1cM��f�V��1@�?���7"O�����|�`4��!�8�"O���D僧#��mi�/B+ֺHҒ"O��9�(�q��M�/�6I+~M!�"Op�(B$٣����Aώ��z��"Ol q6��9<tMb%o�!r&��"O��1i��$X�I�YYh��"O�p	T�\�t���&ʴ\eV���"O�OGZ=�h	��4THP��"O�7 G�b��IKw�X#<hM� "O$A����#,@�xa璯^8<p(�"O0�4��9|d|E
�"M��35"O^��Q��x)Ԧ�	����"Oܱ�!�G����rfͨm�T��!"O�I9�'�2��R%�#.���p"O���6kL�R���p*he��"O�<KaD�S3��ꄠ��m���:�"O��C#�A�ne��ؖ�$�{�"O�T�!�7r�>��/۷j���"O���S�Z�&KBE�B`P�!"OJ���G�^lX��ڹ��a��"Oz�Ca�׷�DA��q�@�g"O��UDS=�ju�F�o�"�d"OԴ�W퇤6�N|Hҍ./����"Oz����Z;[F� �q�����"OΡ"f��$� �96���&|5"O�$�eA+Q�J��B��ٲ�"OҜ��EE�m@��mJ���)HB"OP��"!�5:��M�Uk��%���"On�&�%���s��3/`lEh�"Oh�
�Ry!��JY�zD�Y S"O��I!g��B�0�	G$���� "OT��o��$���iP��[#0���"O�ɋ��?+nNTʄ�
�	1f"O��0�0/X��z�E�{�Dkf"O3E�ۅ �4ӧ�Y�%�x���"O��0����R ����.�v"O�1�fӐ|���U��L8XJ�"Oz�	�U0i�e[�İ_ї"O�!؅���lM�pA�� 2}�B"Ol�Y�M4M��Pf�1]L!#Q"O.|��K*n��`[�6"�\��"OB]PO��R�n5#��,w���"O�(	��X��p���F��5�$���"O �:��V�l�9:wkJ.h�.�8c"Otu�q�Q60{Z��#�7vrH�""OL[eO�x�2������]h8m�u"Olh1�&]$��t��L�q\b���"On-� ���� �A�K�5f�I�"O̐*�-��dp:Q��?\�@��'?�DG7Dv]bUM�R���C���%R!�� ��f�B�^��rm�?TE��"2"O��Ԁ�	U��ƍ�*o9�I��"O��!c�F��dx�+Z�����"O� ���8� �t��j�R\�t"O���i8T4�aÏ�l֚��"O%8�&h�H�
T@4��4p�"Ov(@�kG� ��Mkq�>V����V"O���V�T�XD�B��˟a����"O�pKrJ��k���(D����y���;��"��T�B�L�� ��y�6Z�Eqs��=֮�B#f\'�y�-W��]����DlQR�U��y��X�j1>�[V��4.�Qq`:�y�C��Đ,R�#��{������y�P�Ix�(�"�R���B�yN5��ʓ�M�|ָ(	Sj�y��Q:R���u���s��A�b�L��y"ғ`��x���V�W�4d�&	Ƙ�yr �� �6�:i�"O�$��ˌ�ybn�Nv�� � �K���ZuC�?�yB��*`��=�vi� G��ɨq��yRi�6F%��
�ǅ�B��L����yR�ۀ)XL*�L�A��1Y�iѩ�y2 ��(���	T1Ì�q�N��yb�+��- �Iw��8��һ�y�C�[��ɳE�Hk/\,�v��y�l?nNĺw(*^�9�RD�-�y��)Ť\�'MGD�`���^4�y�bV�Vv\h�����D���k_1�yR.��[��,�B	D�\r�T��yrf�7`G�q��`;
x&HH��I��yB��$���i3���*��������yr+���ˆ*+^�s7�P��y� �[䡓t̗���m���B��y�膮�0���J�C<v�Ӑ�_��y��?>~��GA.5;>�@��y��T*�N�(�fЧ43,iY`���y��r�Uh�!�DL)e<�y�AI!s!\ jrE�|�L[Q��/�y���\Q̘`O��AH�� ̖�y��6O�h��⭅�Mp@-�"JR��yJ�(x%�ys�J6V/H��(ҕ�yҠ�=]��)�@*�;}ݨ���E֯�y��[�$+����x��h�϶�y��>�������6#p�q�W�T��yR�ƫ+c����^�{��#��G��y����z'4�� bK�U���qL�y"`�N��RA�J\h@�Q=�y�����(���^����_�y���_�L�w��"��"��y≔�3���Q��M8��	��y2�ќ>������5j�m��#�y�#��;D����W�=X��)�9�y�MS�1���,�/�a�n���y�J[�l�f�砏?)'�MY�`���y��G�� �$ا(rV�ӥ�׊�yb���&m�$ZA�\� �Iه���y��X�ع� U6!�c���y�L�� �˂�,�u�N��y���#�\����eGlX����:�y2A��Nꓨ�d:Z�Z��@��y2�[�}��%��*�0]����eڹ�y���<-��2fnZ�Ud>Ei�����y����p�ک+&�N�xTXQ �-'�y
� ���%��	B��
#.�q{1�7"O��#a 
F��bb�'6z�x[G"O��2�Ϣ%�`��a�h~H��"O�0s��M�b@+� %"}�<�"O�X@!.U>Du���f��b�b�"O.8q�E�h&@�$ωzY6�%"O�L#���\v\��� L�T��"O�I���Ѹ=�x�*��[e@Q�a"O X秇 hd�$�&���0`�}Â"O�H��D�5"~�IB������"O�ڢ,�ms聱2�L�u���3"O��s`n�N(V�j���-j\�w"O}X��moj��D�O�Kp�"O�@r���
'mĔ+P��v=H�� "O�Uxr����٥�D}D��*r"O�d���ŻB�NM(j�h�"OƘ� d�>c�bx[�T$���'"O��(U�
<WYHDx�M�  �8W"O�3J���8`�i�y.Pp"O��Icd�k��	Pf��(T�|飥"O~��핃K�p=�Q
�&,�B�t"OV �V�Þ}J��IP�N���U"O*���\ Y���#e��y��J�"O2�9���#Va�}�I1s��"O~�(1M�*U:0�5�$�
�E"O�2���"s�R�:�j��܉(�"O��A$](Fx�T��c�k�����"O���t�@
j��
dɇ1b�Yh�"O\!`��R/J���)�.�"m����"O��T��p��1m
 ����2"O��I��B�ᶽ�lC��Ecf"O�xC-Os�fêD�4�Qˆ"OR)Q�gM��HQ:��\z~Ř�"O<���+`<^�	2�G�A� �"O�yeH����٩D��v��j "O)hdB[2�J=P$����6�JV"O�A��[-*f�@��9.� Ʌ"OZ�D�;t��\[���$�B���"O�(YuaЦ;�p�ȏ�g�zMڤ"O@���շ]]:m�R烂Q����"O��sF�g��0KF]-�ͺw"O�,����T1'�	��"O�qJRaPoc`4��΄��D��"OL�8u��]���C�	�}��\P�"O4�#b�5Y�lp�Ē�Z�t��3"O*9� c[)>0�ãM	|���"O�Mq �:e��WMK,z_� ��"O�8���	�=2&�I\�
T"�"O�9���J�7�P��AkD-P3���"OƐ�e��'O�4Q�H�?G1 �g"Ol�g��!`T�1�C\�@�'"Ox��C�*.��s'R�1�8(�"O�{Ќ٦LpB�[� ʬ��T�u"O�A�QM��hP"�-X����"O�=3`/X�m�^X����"�A�"O ������aEG�1��E�"O�0�v��d?.̉sg
�=x�X�"O�[��
�"e�&�s�(�"O�iyG'0\J�]���A"Ox��C�&nS�K6�#up���"O�����j���s���b|�x�"O���D��-[�Hh�˚�pH���"O4乢H��O{0�T��F:��"Oz`�b�	6aYP��Ӯ8�Ep�"O� �����n�x��+^�x�`"O�}���ws�m�F��+g`XM�P"O��(w�������S!*R}J�"O֌z6��'3>��k�/�7F�$a7"O�M)EI�\�j`�vDF�Iނ���"OBL���t���x�<�f$� "O*�i689[�(�!q����p"O�Y�%o\쌲5���;��1{ "O
#��K����K�i�ܕ��"O�ڄ��3�q��f�?D#�90#"O�y��'i�$@a�c[�o�5��"O.M�Я 	Jj���p"�
�*D�w"Ov���ӛ'��$�� VQ���2"O�Z��[�R�l�Q�7s�i�R"O*�Y/��̝S�8��qD"O�]20O&9�DM�uc�-R��k�"O���B�E$�H����/?�1�b"O�Q��RIBH;"�B�5�ճ�"O���+��2a� ���Գ9��ܑ�"O<�;�����s�\��F��"O��)AHǕ1r`�8�M�'Px mB�"O��J#E�][թ�-�'m���%"O��ҁع >�����kN")��"O~���j�>\�㫄�<Ne�7"OLHZ�Cy��@��GkC.��Q"O����G)4t�a��B-`�"O4�@�Qau&�@g�^���ʢ"O�d�FnȲ!G`S��B���a�"O��"�g�hHF���B�.(p�"O2X���)S��pq��Ԇ|��D��"Ol�3q�k�d�.N#U��h��"Od@���3{z<�sa�I,<�Vl�%"O:���M�x����W+Ιi�p�yS"Op�;V�P=*�<T6K�#BK���"O��a#��:e�,b���+����q"O�E�� �Gz��ҵP+���U"OP5�+ֲw��3!ݣX��m�"O�aIA���f���(�E^�:tP"O�Ts��Q�"Dv�u�&+~��a"Od�i�bɺ��ҷ���Π:"O�8*aJ�:}ڈ��n74<���0"O�a�bɌ9o/M���kW�=2U"O`1 ��!A���S��$� ��"O�a5�̒9�*p��'P�m3�!�C"O���̛�vM)��_�x+���"OH���,2C.�{G;����b"OHd� Ȳ&������Z�у�"O��k@G"��i��� ����"O���$���� ��GI�\�rmZ�"O�!
��A�d���q��[�"O�Mst�;s�TP��D��,���"O��S%C^/24���^�z1��"O�dbU�P-���j0G��af"O���!�[?T��2�(C�T�x��"Oz����6_��"AF�N���C�"O�Hi�O�A�c��
PM�d�a"O�Yp�
����(��[L?��a�"O�d��ᔙ��5"�m��_�-��"O���c%5��Y6��*e(�	"OJ(@&��(����1�Ŵk����"OH(+�k��ʐ�	���}��qH�"O��s�a��J�)2K��@2��p'"O� f/	�9����J�	:.rm	2"O�� 7�C
oKHЈ�A����"O� ��2���"*�ȉtM�!g�@��w"O�dȂl��f��ӟ^���Ae"O�mX���.��Uk�e\�Ht�P�"Ozթ�i��"�$� 
�Ҥ`�"O���(��k�r�b�早[؜=Y�*O4��4�I-+j*�S�RD��*�'�E����E�EjӃ�+�<��'�*Ƭ����B�KrސT��'��ҕ�^,.����OҲdU��'~�]�s瞉9D���ٶTB=��'�n��팬l�����f�&�>���'f=��s�,�p�戄=!j���'�����W-0�e�"g�^ɎQ�'�rs��!�V���׌W(�1
�'jrm{��S'�*��Y�N�Y�'�52�L��X�p���*Y��}��'6�}3�mJ�V/�Y�U�O@���'��-@)��5�V����J�&���'��U�q��!�|=�CfMpT�+�'��Q�E�D4���MY�X�D��
�'N)��G��j�����S�~�Y
�'y�]:4(��N��)�6���Qφ�
�'�dʲ�Z9*�]J��9��	�'���E	�X�~��!��-+NH�'��wf�U���rCD�V�`]��'1`A�B"��n�<�{&�UeJ���'kTղ0i+�މ�����[�p�x�'7��3���u <X"g��!I��
�'����+��Ed�,��l�:��YJ�'�Zt��N*DP�[7�A�	nn��	�'�&ă�%�g��m�`��0ș�'�����@�a�f���~Ѥ��'����d�4�z�q��N�s��b�'����u�0	�|�@� h��`�'{ DZF	�N{x�7iF	����	�'���W�L�r&ӆ�5cDe��'z��1�l��qʰ��DH..����'��-�&o2C*�U����*��Hi�'Fh�m�
x�\hd�Ϫ���0�"O�X��&b�\ �ȑ=:�v�s"O���F+"���1jT�$V�:"O�ic�JQ�k�Z��q��;��L�"O6,�����<�f ��g͌K��`��'3yi�
�_L� 33 �,`��'�*�3��3w��y V'S�k���'V�;4�ۃIF{�*ưcD<�B�'�n���ٔ#0R�"PJ�'M�$�:�'`�8#!�Ո.�d��̯-z@��'��<2ЮA.���bD��*���h�'2�H��,+*@�{e���ԉ�' ���>nD���ɵAF�
�'c��+��K5��
%<���
�'/����K�ޑC�����1�'�pܻ�_�!Č�)AD�`v��
�'-��� ��7I�rDK�J���'����҂F%�0̚!=yʡK�'7���&n��Y0����Ϲ%tjD��'�ȤZ�`	�iY����p70 �'㞐@��,B���ޔv�D�#�'�D��f�=15��X��3S���'�(�1� =4���G%D:|@��'�*� S�D:B��)i\�.�`�'�h� �+dED��s��4S~���'�RI��CI�.�V��Ɖ����x��� ��0�M&�� �
�'��"O�<��EW�qq�qqc�G� ��Y9C"O�k�*H�I��+A�6�Ae"O	�r�ě*�,���3	� H�s"O��s H#��2���{�½H����,AS�LN��iũzl>��%�M"�dJ�GA#g�qO0����SL�A����8�F�s2�=~ȅB�O<�+�������bpO�.7�������̴9�]ڢ�x.��$h��g��p���P1&˼�)�(�+q\i���.-�H�r@J��b�`<�"a�<)����t����MS���)Ǻg,p��%}HcǤ!Ȱ�ʱ�'L�O£}���$ΆP�eE�pHƝHP�T����Ğ٦�(�4�Me���)8�q�LT;%����$#�w?�*W:g��f�'C�)�L<��/�"m7�]S�
C�iV��2��G.,�4�Sݴ]���	�i��f��e�Ţ��O�����b��w"����Ȟ�i�n lZ�z��,��'X�[¾ �2��;6xȜ`�d�,�>��%L�kl��j*�h`坘F8��:�ቯ �MC��?i����O,>7��?+x�2�ᖈ
Ұ�$�W#
����㟴$��G~R�U��ʨr���_: ��L��(O¨l����j�4�P�$�48�
q��]B��]�pr4�:�M#�|���x�g_	N��f�J_�d��NE�����4`�RĨb�Դ4��I.�OxQ�A��=x�X%R͌�\E4���"ۍ/t�}����|�%�],�ݐ��Y���*b�n6ܕ��4��j�<`�LE��(�!-:�`�DQ��g*�O��Oe�r�$W�p"�*ؐX�nA�2�")sjS����hO?�ĉ�wܒ��Eӓ"g�U�Á�(S�����4K��Ɣ|�O���W�x��	�sܬ@3'f�w�Q &H�L
���Fʊtx�T���lr.6��^�����/�3��5��'C�<�R�p�	�l�:$H�(]�o�"?i���
{ހ�ׁ]/ ��xE��𐪥 -��{AB�1Q#RO�h�伱/Q'#EXt9(O�����'_����5���ɵ���{0LH�H?�7-�Onʓ�?�(Oxb?u+ ��r���އxN$�ӥ:D�TK�4t��@�!N���zRa����ٴ9�6T���׻�M����ħA�5Z�j�MDD cGS;����=��X�����(ܲb�P�A1�O�ڱ�vKz>Ţ3a�4�0�;Q@ߦR���k4ғy¤E���R�b�M)�ɟ1Qr($��,V�;3>$6�5,��a
"��Uè��R����5�+4U�H�.��t�	ܟljٴ�?����yBj��:����N�e���f(_ҟ�?�|�K<�F����ఁހZ�pm�4��g8�	ݴ=C�6�i
xu
wĔ�I2��R���P�@j�'�R�ۢ�v���<�'�zL<���uz�u
V�M�Sg~�ڴ��;��)�!_�pZ�y'�3yd�x 2�Z�'���8����F�9= ���s�^�$6͑�f����I�A��b4fE� 3S��"��åU*����hi�E�3�d˂,@1u9���7�i'x����Z���<%?q��M�&�;E"yXW�L�i�
�-s�<�GU->$�MR��^�)��ӓ.�y?1I>�p�i�T#}*[w���� �ց`�a+D��>�~5���(��9lO��9`�  �   ;   Ĵ���	��ZP�viė:&���3��H��R�
O�ظ2�x�I[#�x3۴|f�v�J=|L��gJ�'��l� j'�6-�轢ٴ.q�$0��\�I�F�p�� I@��4��X����f$?�!�r#<) �d��&�R�~��� p�<
'��`�^�xQ��A�Μ��'?����6}6-L}�D��$�A����36�̣ln*�c�CN^y�C�ODcs�ʎ��9O4�y 
�/��cEI�6\��L���X����b�8��D�`�葰1����'H$�n��$iq��%F��P���q�'�dS�	�lu�'�����K �R�	�7
�j�h�'B,FxBDH�'I���vjƓ4�T����ܥ/I���O5Ku"<)pI�>C䆚�J�PMV�M���/�H��OT�R������'s<!��m:����)�*rY�8i۴;WH"<	s5�Fa�*�Ɏ(75Z� +|�;qh�Z�>��#<1� ?� �B����P�¦.x2�Kc��Yy2��~�'���?I��ؗ	h���'��MY|[Sj�?t"<�e8�2����н)����B�R�]v���s�C1O<� ��$����~B���p�� 7|��ukƐ���lT"#<�m5�k(:�R�^6V��-AfՈs��x��o��X�K���i��mGDq�����|y�@�3z���*��$�B�<a��"T��P�<�2k�3Uo�O�2��>R��#%
�f�>I�s\�l���I�-C��Qe�:2z���P�:Y�I�"7D���'K
   �a�N>�,OrE�h��y�ޅ"#ŗD���8c��O
���O��O�<A�iX|����'p��12���P(� z�p<p#�'�~6!�ɫ����Ol�D�O����C?[��}���#�D]���_�7�!?u�y�n��7���)y�J�1_`@2��j4�e�qK`�0�	�<�IܟH�	� �ґ��)i�1y�i٫b�� �/ֶ�?��?!$�i�ЈӞO!��r��O8!%FMy�jDbWHLD�ސr�J!�D�O^�4�b`��k{�|�N����-hm]@�Vz�<P	1)��I@��Ty�O���'o�k�$)Wbԁ��	"{A2M�G�A6T���'�8�MK&�۔�?���?-��P�B�@�
��@����8�ٳǟ�p	�O�$1�)҆,
	���i���[~�R��m�Ρ ���A_���*O�	���?�7"���H�����i)�"'r�v�IE�'�r�'er���OX�&�M�b��= HD���Zo,\�%��tV����?yu�i��Op��'�b-�%x���9�G�e��=HC�S}�B�' ��F�i��I%cUN���O�>	$����1i��4k�k�o�6�ϓ���O��d�O����O���|�� Сb�u��m�	<}nq�Q��;}\��(N���'6����'*6=�0Ѩ�mPD��� |�$��G�O�b>=b�	�ئ��7S�@hvǗ,w0�V��{ܬ�fw�R��O�Y�M>�*O~��O6���DZ�w�<�
��3�>�;ci�O����O$�$�<Q��iD�I�'V��'�`��@�ޥE��(v���o��Z�$@}B�'k�|�I�(niv.�>jY�4�7�ª���\�jԢ���,`�Lc>m���O��=a����C�&k�*\め�*�����O��$�O���4�'�?)ӭӴ:j s�텞P�(�SW��?�a�i���S�'�"�z�f�村0dΙ C���u������%sw����h��ߟP��LM�q�u��� rp���ܘ��i0ŋK�.h񻷤2I�L�$���'+R�'["�'�B�'�J�X�T�%�f8K���U�a[����B���?���?	O~��zoQ@۸�-*Ԩ�S�$wV���II�S�'"x��(��R6"%&QB !8��ة�mG�� �a(O��c��6�?�$�(��<)G�[�`��m	/G�0�?I���?y��?�'��$�Ŧi	�-�ɟ�:�)��E�B(�V���V���ڴ��''���?����?�t��g�b �T��:Rl�	��m��h_�P�ٴ���ʷn0Y������А�ħ��`I�m�eP�,#�5OH���O����O�d�O\��H�+gl��bA �H$��=ْ1�C Rj��?!Ľi�z9��'��'�1OĄ�w!J�{��=��̭�>AH�O�d�O���Op��kg�0�	ßHs�߿G�"�"7ǔ�OP������kt�'vL�$�ԗ'&"�'UB�'�I�D��/@^�S�o���F����'{�V�<��4Q�4�����?����)���L	�_C�|��r�F�������O��$(��?�!��/֊e�%�̄3�.8���>v�C�%��Zؾ��|J���O�}�H>�]����3W���adзlP�,����?���?Y�Ş���_��qZ f�_E� �Ud�e��jg���4��I⟔�4��'2���?�W$G9�V���.�"�d3���.�?��ZsT%��4�����*��矢ds,O�x����W�T����xѾ,�P0O˓�?����?i��?������ɿ!鰴�!^tш�F��n
V�>Д'{"�)ͦ�2N!����K,JG���GhJ:q�!�	���&�b>Ց��
Ħ��S�? �yT#ІLƔ�7��;Ԥܱ�8Omơ�)�?�Cm#��<����?��#V1 �׎�7Uo���ЃL��?I���?y�����Yئhg�cyr�'I09�Cگv�J=�S��\D���d�b}��'�қ|�G�;n���$ODfI���"��d����!�I@{1��%��E{���Ţ{K2m Ȟ5pʉ��JZ�E ���O���O��d"ڧ�?	��Y$٦�v����$y��3�?Y��i:\=JS�'nbl���%V[���B^h �F���ȟ4�'H`��նi���&\�80�O^l��F0� K�
� �<��B�d��_y2�'Z��'I�'�""ǑR�Y�b��4k�yc a��_<�	�M�5 R�?����?������v�E�Ẅ�_3��b� �R}꓂?����� �x!ڇ�w��l���̰�"ʂ�p��+Oh��&
��?A$'�D�<�5�˨&��bL�uj���]��?I��?���?�'���֟,���?Q�'�zI15Ȇ�VCe �斸�?�b�i��O���'-B�'#"l�
&��)㇫�8���%�Z�����iG�	�djj5ӂ������M�2ݞl)�j̐"\t�Et���	ޟH��؟����(�zԧ<3m����a�u�V@JK�"�?���?9E�i�b�Z�Ob�
b�Z�Oڍ�c�Z�Z�O �kq��Ӧ<�D�O��4�H5R�njӈ�v����u��>�E�b��*u���D� [�4�$P����4�����OH��D��}+�.�m�Pp�E� ;�����O�˓9P�v`�/Z��'%2S>m�R�:�@G�0)!�e�pg1?�^����ޟ�%��m�D쁔�·5�r�3��7R���Ɇ�_�Y��j��4�V�Z��@N�O.��؈+��aA�M�; �B�� ��O����O`�D�O1�X˓hU��/E�
*pp�$�,hM���v"
F�����'K�n�H��O���C9x4!I� h8��7Fg!A��<��i_N��a�'��X��@�?�#W�4P��Y:h��}S���	;P �|���'%��'<"�'���'��� d�}K�C�],���,nv�ڴ	?���(Op�$!�i�OHylzޑ�3��M��� ��a9������L�)�5e��	��t�hA�L�?;�`|�Ԅ[=5�	�t����FKN�d8��<ͧ�?�b�ۮf�4��ƕ�a�6��W���?���?�����D����B�uy��'��e� ��&f�&]ag�>8G��R���z}"�'
�O�UkL	3��15.]�M����p1i�/�p5�d�c�.�2��<�%@��5F0����_�*8��O���	���	��hF���'��C�	u�=��-� �0� ��'\7��Jָ�d�O,|m�U�Ӽ�`a�7S���EB�g����I��<1���?9�Z����paY~b�ݷ#�:Y�S�o
��JP�>B�y!ٶ�*4@��|2U������ǟ���џ QP��e��
|J,��Zy2$h� ��B��O����O�����5'����T)9��<j3Y@Dq�'dB��i�%b�0��*�.%b�h ��0K�lȢ��L3M��;�@��+�O>Q@H>�)Op ��v�le��dBq6PV�'Ub6m�/���:�t��`΃#<���卓�A�.��Bզ��?	�U���	ǟT�I9�A�CޔZ�f<��]c�޵�C���t:���ֽ�ǃ�`��H~��ABH��`�:.��p�i�9��X���?��"�B�׀��E�f�3�?)��?Ჽi�ΡhΟh�o�U�	8)����0��}XV�V/D�B�'���I���Ӈr�y��/?�;"�fx�C;>W�����x��@�^QP��Ε�����&�ɘ)�p���\&>
6%����1["<	$�i�l���'�B�'���)��v�N.�L��u��1 ��W$��џp��~�)B%�=+*�j��\4=V0¥��<Ub����ʏ*Uة�)O�	���?1�f/�d�U��0�	4�Θ
���G�!����ƶQ]�A��$T(-,���-�*WNhx�I���ڴ��'��ꓕ?y��T�� 8���j�B�Aԩ�?�����!���A~�A�<��'��K(�q8e�k�z�J��	���<ߓ D���ǀ.�x���؞�e8B�i���ؕ�'72�'�P`lz�	����}vm��A�)�z4�4̎П8�Iv�)�??���4�y��j��K�*P1	VhQ<^vdX�/b���aQ`��*��<�*O���ǖb=��T� � �J�'��6-�3%jF�d�O����AQ��8L��5\�)�e!�5 �⟘��O��D�O�O.1q���gf��pF"�	{0��R�ʅz��V �w�{�� ����tmM�r�$�0Q��/	���(D�ȑ��=\H=2uT"I��*c$�ߟ��۴�Ƅ���?)��i��O�Ν�[�t��ĎEu7���t$�?+�D�OX���ON\Ťܔ[}�i�;ҍ_�?�2�� a�b����H�G�@�k1�V'2��'��e�'o.����*QLh�����>�T�O.�m�+v��x�	۟���V�Og���p�S�6���π�]L]��V�\��ޟ�&�b>)�Cb1� :� ���#?o~�H���IQШ�b$�W�,ʓs��EɃB�OH��J>�+O�t��e�o�J�  E:M�U���'or7��P��DI1*�mp#���״�1�X�O����ĦQ�?�Q���I�,��1`�Uѥ�n]x�
ËRsh��!�]�f��RИ&��!�J~2��T�p4�	?"fU ����iM�Γ�?a���?	��?�����O�e9@ �	K�@��$A*�
]q��'��'�6ړO�˓y(���|2���i �)�J�њP���ѽ��'q�Z�0x#��1V�iR�E��'�<��vA�	1��q���Y֦�dS������O��d�ON�dZ4h+
�k�U�,|P�rK�Y��D�O����� ���'5�U>�a�N�C�h��`�<L��X���>?A�Q�������%��'<�4q�ΈMD��QA#Au����IġT�Yv~�O. ����+4�m��%Ц$��e�Q%�=A� k���?����?�Ş��٦}2@,��#������3#j�����ՀH����I��Hsڴ��'Ō��?���-1Z5�)
Eb0���͜�?���\���Ѥ �]~�#ƠF�<)�}�	T36P&PX�A	v6|'���<i+O��D�O���O����O�˧2�D�R�I�4e>��LԌ{���Q�iz�P�&S����X�'p�w[���1�� -c>�5��6q
��'��O1�j�H��D"N��D��	Ơ"��BX��h�$<�D*	:���)Ap�O8ʓ�?���c?��7ƒU�FT8�GZ����I䟬�IJy�of�2HE��OX���OXd��,��D� |(g��\4 �2�%�I��$�O�㟜 �D�=4K9jTmj�MR�<?y�h�"w��
�@����'u����?a!$A!OF�IJ�(!Jr�����?���?���?�����O�T�0Ț�O�V`r��ڈ�P!$��O6Ilڈ)�H�	����4���y���:[ẖ*X�uJ���`j(�y��'���'0��Z������$��>d) �O�*��R�P����6��.{��)A�|R]�T�	ß��	�L�	�tK  �.b	b43��z��Hť�fy�f�p�w��O<���O���:��_/v�$��
�tӸ�����OD���'4��'_ɧ�OM���@E�
%|�	e-+i�)�gfW@f��GS��"��]9��/�D�<�`�K�@U���F�H8xY!U�Ơ�?���?!���?�'��Dڦ�"A�ǟp�@�]"S��X֬��TM8�`��Hr�4��'�L��?��Ӽ�@���>7�D��C�<L�ę䅉#��(Ac�z~"������䧉����(�F�A�,@� ZVpA&L��<����?���?��?I���a݁��R��y�B���D٦l��Ɵ�	�M�B-��|��/ʛv�|"d´DP��˲OnF٣����O>1��?ͧ
�d�葧�Y~2d¤D:Lx�(:q*��&��$�~(@��@?�J>q)O����O�$�O&p#m�K�T,B�bR��xR�'�O���<��i�X���'l��'q�Ӕq-2B�O�	�:����3y��"��ӟL�I`�)2n�)B����QN�~jq�,ƲS������[,��H�-O���Rͮ�J�Fz(���+�#+ʦق�葧 �T��0�вz���{��"&�v���@� }�J�	f�y�"ꚱ�����ݨN�|1:#�<��2g܂Kg$ n�/@��S��� 5[���5$�I�=�^�:B�tzh-B�o]>"�yF�&�nš1G�I�q��Ή\<���hP_�!8t��R�쨁D�,>�ޥ`�B�}{Fњb�Ó,$�}C��O�0�xu�@70�h��Vl@]R���RQ*w"���sĩc�>tqeĊ���.SX� �J�_�ʘ���"f z ��m0h�|���/�7Q�� ֆ����<	�����?���6]��d�2j���L���9�"�����?Q��?�.O����V�|
�˄�g��A�&F�!�Ź�������'�"^���������v8���#�������*��8Q��h>$��O`���O���<�S��㟀�pAS*QC��Z�OF$,�A��MC��䓜?I�W�R=R�{��;)�aY�E�>�И�%f���M+���?+O\��E�@H�D�'g��O�D�8�!�[�=ؖK
�%���t�<��Ov�$Gnq4���'��q{e�7i������
	�(oZzyB��>��6-�O����O��)X}Zc���y��m8�pʓ��V!�q�ݴ�?��l���Fx��IWV�>�9q�ӕyj��E�ƫW�ƅ��6��7-�Oz���O8���u}�[�t
�ƶ01�X����%gx�Q���M�Rcȅ��'��8�D\{��M�3dC(��͐g�":��l��|�I�����f�(��D�<1��~2�$�ҀJ��̬K���Ӧ�M�O>��`٤I��O���'�2	��x��(r��v+Ę�n]�da�7��O�ei�n�@}BV���	p�i����IÙy��Ǉ�g�a�n�>ad�T+���?9���?Q/O��C�̞�
PY�K�*��xö���"�|��'��	۟t$���I۟�iO�;C��5bwOS�J�6]���_�\L�'����ğl�	cyr�ā~�t��M�e�S��,P�+�hֻrr7�<�����?��j��t��'/��U�W�!�l�7K�8�O��D�O����<IeKѭF��ʟ��% ! <H��-��~T�8���!�M+�����?!��N���{""��@��0����{&fXXf����M[���?	*OT�x�E�`�T�'��Or�C���7��9q߰Z�Lk���W�Iӟ��	�B�$��i�IY� <\ʠi@�?�.����ߖM[ �´i�.�����4&L�SߟX����DC��~�{UM�Y ����G.��Q�������rI|�M~nZ	���3��!���1��.wAt7�M�1u�lZ���	П4�S���|j�(J�"�PQ��	B
[X�J4I��y��f�'[�'�ɧ�9O���%Q־�A��H�kx����.��pmZП�	ßTP4�_����|���~�,�P7�x�	_vr9�d#�ɰ6��O>�O�a��yB�'}��'�B�ST��H.�=+��G1����6�g���ę�H��$���%���3�/z��� �� \�h�S�T���?�I>����O��`�g[�0V-R��YR�*��q��|���?�����'b�O ễ��	T���/ɼf�XC��iH�i��y�'f���Xv�Zr���@-oX�cΈ�Q�����ۦu�I�?A����\$d��F�[�U(x�Fɐ,b^�M�u	C-���?9/O��$��`�f˧�?I�j*^CV����#�`L�!�'m���d�O�˓iQ��%��
@@�/���T㝊cVf���vӞ���Oh�G'�`���D�'n�\c4�ȃJ;:,�3׮��Fz�PL<�/O.���O�����tIb_�9���*��w^xI�X���I 1�p��ݟL�'1��]�֝�'��QR�B�&����d�|�@6m�O��X�DxJ|J�͐�1X�3v�>�� u�Ʀ���C@��M[���?�����x�O�L�9&�߃*�\�! ]�,�42��b����O^�D=��?�i�v���Ϛ��`İd\*\�ȉ�i92�'��`@�1��)JJ���k;��#UA�#}��8'm���OZ�'>Q�I���	�Y�p�`���@:�TIX7k�T}�ٴ�?S�/����$�']ɧu�0Y"���Í?�V	�����?Q+O��$�O��d�<�~a$���^�0|f�9��&g�<Ԫ �xR�'�b�|BV��}!RaEp .e���N?o�N��|�v��%�d�O���?��.T7��tN�)PA��r�$_�D�}J�!ӛ�M����?����'��	$j7M��Z#��S.W_�D�iRc�/���֟��I��l�'�h��a��~��Z#B�z&�,���R7�	�{ bç�i��R���I����	�;��|��N�~�5X��7#n&٣���|����'�rT�,7�J�����Oj�d���i8!�+@�
���LT�(�}*��C]}B�'��'�yÙ'�'��џd�b�K�3R�]��Rt+jyV�i��ɞ̈\A�4�?)���?Y��W+�i���5���N��<�&��5%z�uD~Ӥ�$�O���yB�'��IZܧVBq�u �&x��2t��{�pLo�����޴�?y���?���#��	Yy���Y\@���<e8!;`�ӵa>�7�B#��#�D+�����qQf�'�"���fI�H�(�r)��M����?a�=���C�^���'��O0�w��|�`�	S�.<"��i��_��tmi��?a��?wb�j���ĉ
{k&p M���F�'~�iH� �>�(O>���<���C�)T��&�����;��H���Y�!�	�Z���ݟ0�	柈�	ԟؕ'1H8R`hD� }+`S<Q�D8�Õ�~@�����O�ʓ�?����?��\� �e�Mʉ+���s��
�t�Γ�?���?����9O̭����|��J��bd�"�#N%XEj�\⦅�'F�[���	̟�I�0����(/�\q��oF1-i [�@o�d��O����Oz��<�7+ Wn�ԟt��D֟�@]��S�3�KV�|��Im�ǟ�'���'��y�Y>7����p���'J�0cFȠA<��'��T��h�@�����OZ�D��b(:DD@&,t�8qdĕ4<��B�d}��'"��'����O@ʓ�����6���!bŞ=+��	�����MS(O�
�ș�����������?��O��XJ����B�]D�@l�#"d��'1�N���yr��~�ܸO�vd�F$_�L�����Z�Y=BJ�40�s��i��'��O�2���$�5@E\��P��b>�q�s�;�|o��/\p�I����'-����̯X�q���d�-�A�Ȏ+�)oZ�� ����R�`����<����~�Lѣ1�z���=AĨc 
ߛ�McL>�T��<�O��'z�h̔H��Cs읬)މ��$�#�v7��On�p'E{}�^�X�I~y���5C�xl�!�c�ڳj#ʙ���ƀ����d��$�<	��?�����8�LeC�@[�E[�tj$�=e���hA̋v}rU��ISyb�'8B�'�"���
R�R�r��@�'-��sT�V��y�' ��'�2�'��I$����Oj}��?���$�\q
�Cݴ���O���?����?)����<�1R%��`&Y'��e�i!Tb�/�>���?�����d1�*@�O�� ʎ�C�DGvf�G�E�b6m�O�ʓ�?9��?!���<�O�8�`�V9�N�{��_>K�ݩ�j�����O��n3Py�e[?Q��ҟ����Z�N�y4�2) N`�Dc�"\�b��O��$�O���	B��	Fy�ڟ~�)-��K�,=��	�[�i�w�i$�	�/¡)�4�?a��?!�'H��i������B��q�Uh'f�v!�kf�~��O6H�8O`˓�?1����R5����A��yL��	-�M�?I�z�l�۟��Iퟀ�S1���<	��U#v��Y���*o��1a�r�f�ܵ�y��'D��{�'�?�f� �i�tL�M6$Y�b)ƴM/|]�S�i�2�'P�Ɵ8�����D�O<�ɿP��ei��RY���фA#-��7M�O>ʓK����S��'���'��M21CD�vD\,��`ѧnc�a��o�d��ֿ�!�'Y�I����'XZc�҉x�O����6iU+a�)��4�?i��<)-O6�$�O`���<��KߖX$�ɒ�s�8Ce���IdLi��P���'��\���I���	�<c*%S_{B�����}t�#��3?��?����?Y)O�@����|�q��tD6Q��H :����ئ1�'!�_�4��柀���E0OklmI ���1j
���NѲ1�*e��4�?���?����d�,���O�Zc-|}P�x�l�ӮA�&�9��4�?)(O8���O����mV�i>7�߼�҄90��(bT� cCO ����'UU�t�#J�4��	�O����Vl�@ �B1 cD>t,�i�&O�B}�'"r�'<���'��'Y�Iz��0)F�?�X�Xfb��V_�4C�����M#��?����rgR�֝�_����0�|U�TnX��n7��O��
��$�m��'�q�8�Qsa�5/ԕj-��=��� ��i��t�(`�r��OB����'{�I��4a��R�TӵI��_���4c����?�/O��?�I\�h�6��="���z��F�8��4�?����?9��P�db�O������U�R>1U��q��T�RU	nӦ�O��!�8O�S������P���MR��S%*�7P"8� �KF%�M��|���21�x2�'�r�|Zc��P��hߥ4U|�KX��~�q�O�86Onʓ�?)���?�)OH!������[TK�sBVD����<�%���	���'���I��t��B;<����B "L_��R����	]y2�'���'u剥(c���O�Z4��Żw�:��s�W�.��I<�����O����O*	h�7O�q�#V�U�M���ΠDI��I}��'�"�'D�I.AC�uYH|��� �,�r,q�	�. �p�eɟ���'�'��'z���d�* �|��0LW�t"�w�V�'W�S�l��G��ħ�?Y�'�h� �Oc�zi萃��5�2�x��'$�)0=2�|R՟d(fI����3hW9ӔU�i���I��m��4M��S˟�ӈ��DW�"��s`��b�g��0�F�'����yҒ|��)�-~��]��X
B� ���h֚4���hX.k<�6��O"���O2��Z�	ڟ��&�$h`�ms1�X'q��-z3�K��M�`e��<�L>�����' ���cQ(e�L�F۲P
j��
t�X�D�OJ�D�$����>Y���~��_9mP�}�)RWnR��-�M#O>q0ܹZ��O'"�'��IK-L2���C��Q���ƈN���'�����3�$�O��D)���*A��ׄ��2a)ɝ!�H1r1Q�0���u��'�"�'pr�?�#T��M�H��W�b�v8�B�Y�v$��>q����?y�H��x �ׅ[W,ʥf�=g�\��ր�?�-O��d�OH��6�@�Z����Mrz!ku)�X��#�k�ē�?O>I��?����?	`�F6|m���N�YK.<���J�jc�	�����ڟP�'�0�i�)�)_�`�0�tKؐ��1�r��� �mZޟL'�D�	ޟ��ĭ���(�Od�j�JՙD�m1n��2�^���i%�'#�I�!�l�{M|
�����JR]$��2#@ :��
A�K�@�'u�' `x1S�']�'>��ʲ4�4H��	C�/nd��1`�L���V�8!�>�MkY?]���?M�O���k9�h�Ч�)|���2V�̕'�������G;��ꚒB?�e��L�	�M��CJ�c�v�'Xb�'<��" �4���9��zAP���J� vUv�Q/j}��'��O1�@���n��-/j�����yx|nʟ���͟�a.�KybR>U��O?�N	�I�2��&����x�@��r�4�I|���?���% -A�o��X�XW����i��怼��O���O���5}b�;^�$����X��7F���D%N1OZ��O��d�Oz瓰-���3b��< ��u���^�q6`�ȹ<Y���?�����?��'뮡*׎�	�v0C�EѱK�$ݴ+$��'���'ar�'��)�	��i$TؾP�sF-%��M���� Su��Z����s�Iܟ��'Y�y�4~��@r��K�2"az�oE�&�4��'`��'�Y�8�3`F���'#��I���2\F�C���@VY۶�i���'��Oڈ�'��Y���A�e*�t��Ƀ�Ƈ3ߛ��'���'xb"ԍl#�������?Ř�j�<3td�ou2��7�Ӊ�ē�?y)O~����i�Af�ȍ*��S��ؠL֤���wӎ�b]Ha��i)z�'�?���FR��7
�
ْ��Ŝ_�f)j�F�"+6M�OT�Dދv1��}j�"[>e@�	��F	@������.��M���?����$�x�'��K���@eb0�D �̠�� o�JI�)§�?�A�{?�X��l�0"��`ᢎ�jh���'�2�'�hI9�b-�$�O�����ԛ�	Ҫ��Z0���	)�9���=�	c���	̟���&H�ܹ�G�ߐN��Y�$�T�޴�?�w@�D�'/��'�ɧ5�.� :Y�傰�v
iZ�k���dC�Ib1O����O��d�O��B�? L�GY�;�҈���|a ��aߤ���O����O�O������[v�XE朋1�"-u�zuK`Ӑ����,������	QyR
�)W_�SnIx8�����4�"iK!o�*��?	���?��r�����?K{~-��\<NK������Bo�I��$��ɟ���|��!�g��'��4a0�$x�*˳{@nxq��D��"���OF�*�` $�����H	y�̤@�*<!���cNbӶ�D�OZ�?��� g��t�'��ġH(g$.���9�8�q��<K
O����O�����~Rp��*:���f/�pQc%��ٔ'/��s��kӎI�Or�O��n��q�FY�aTY�+1���mZ��,�Ɉt"<I����B�W2Y���Bw��yE����Mp
&4�V�'}R�'��i"���O������Ebz��F�d����v�Y�y��"�S�O�r���l|9bD&M	_  Q���3�07��O��d�OҽH�"�f�Iȟ �IL?��N����wS:XP����L�G�8:��<���?���8y���i��)���i�l�
�i��挸%��Od�d�Od�Ok�ݜw�F��gL:L�6������z�	n2*c���	ϟh��]yr��9� P�L�9(��G(_ a��ܓe �I��%��	��|)P�� {��ٱ��r���,�	$b���	ߟP��ߟHͧD82��� 6�Ma -����rF���v/FU�ߴ��$�Od�OR��<Qq Ʀy�r�Th[(���>��	��b�>!��?�����dQ&Qnl&>M U"�V[���4��<Ь��?�M#���?���CM$��Ob�iӴᅶH|��X��Gj��h��4�?i��?!���6�����?����?��'e����R�E��:`��nG�f�ҵyÞxr�'��+mь"<��~h��T�����4CUE�$~~�oyy��#*t�6��x�T�'I��H(?��ᗟS�5��嚮����A�����I�̑ D2��O��Ic���
^�c5��">0��4%�z=�u�i�R�'~"�OC(O��d�-(|M	��ح&��%3G�ڌGH��nW��"<E���b)L��%h��={$�n&�����r/ʍ�����G�'BF,㦄^�)nt��	�?b�b���1^!�i�a ��_�2$�SGW�:5�MCU��*zHZ��E�"I���?BQ�#��K�b���ER�mr-���7k�����D(��x����Nsv 6-ô.P� �B��	%r�Ku�9w�jKB�C<7�8C��XL�P��Hٸ������ � h�$|��$�Ot��O"��`�O��D{>)c��7/J�щ(n������x��#C�!�J8���H(����$Ҫ";r���U'V�!�6K��Nf	�sNC >�֬(�ϓ֦1X���ceg�09X�S���:c$����t�GaB�#��F��y�X�VnWZ�'oџ�Y��8��*�B�0/ئ5�3
;D�d�E'ՁnNҭsq���aQH����y���O������'Z����p��b���.C��ܮ[�~�;��͉P�����'�R�',| �����X�w���S��E�[�y("n�6j(�j7����dK�`��tH�����}�RH�9A��9˴��)EkI���GQ�'~���?Y���%��^p�o�,L�:D��Ǌ�yb�'fPD�D�*Y(:#��e$��^Љ'5��xWCC�a��lB�mZ�rL��'(���(�>1���iV�1H��d�O���ʓD�X��Ūצe��Q�HOt�|0W���m��.8(,ק�7��O�M3#	�,F�
�9p P�������ڠ�pḦ́J��ѪO?�DO�;=������0�t�#ń���C�O��!?%?�$��2�ùC���Fۡl�v �B�<D�LKƄ�*�>q�pO�thؒ&�.$-���?�&��1�ۣc�TD��É0]r����?i��X��Н ��?����?�������O�iѰD�T��3����x���O�#C�'4�8z�c�Y�搱�aJ�U ���'�x��"`���dW
|����ɍQ����$�R��	B���X�L�X���b��q�,��!�,D������\��r��N ku�|qe�ɵ�HO>��C���M���MY�P�dۙhr�)�n���?��?i��2
z)���?��O/�)���?	`L�(8�N��C�&'�]1u��P8��ٴC�<9P�[<t"�	��6'֜1s&Q8��xsF�O���F^NRv#�	I�dQJ���
�'�B�@���/F	;C��V�H�		�',Z��%�ш:��TQr�ƔZ���R�'m�b���g؛�MC���?a,��0J�;Nly��,у�0��M�9p�����O��N�\�(�|�`�X�4�]嫈16 ���s�''ވҋ��C�(�v�jP%�w�0X�ĮP}�Q���L�O`�}���O/	���Q�έK���qՈ�h�<��Lɏ-j��!�K�2߂д �P�hI<� L��
F�;��{e��!b���4O@�� ^ަe����OJ�X�5�'�b4O�hu@��-��]���_��6�B"I��y"�T>#<)r蚞�l�k�!֨�0��v�"�l)Dy���'��+�䞮2���T%�
���qM �b��'Z�韘"|�	:eJ]s@�	0%:X�Qh�;v�P�������	�E:�4C�A
6+p�0N!�^#<��)���AC����Cؔ9&�yuA��?���-؂��%��?��?Y��8���OT��̕I�fD;G&�s���XT��L���"��}�	 64I��ї �5Z�8l��b���~BȀ���>��"@�|biKA�4� 8c#�Mp?�SK[˟���	�>˴,;�ȵ~*��a,�K�HC�	;g ��qr����1�a��~L�����4ڸ{ڴUU:��JC�cplD��W #���P���?���?1���?y���tdZ�?�<~)��&���
!�2�ܰ(�݆�	D�j��Ȭ���~F}��-JY�D؆�I�*]l�D�O�`��Q�y|֐�k��_(n�ڴ"O�e)"�F=bnH�Uh��&R+&"O�����]�s�R8��H�4u��3O&��>Y!�ҙc�&�'�bX>ݙ 蒥h���h�1����-{t.u���p�	�:��L�	g�S����'`Z$��ڧB(B����(O���Ӧ��ӧ4�z��%����<Y�*�6m>ڧ-](������Q�Ԩ���J^�a�ȓ,�5�� ښ)���A��T�v���-��;���F�X=n
�B�� �ϓG~��iHR�'j��w��%��ΟX�I2iX���c�V8$�I� �a\�e�t�Vٟ��<��O,�ʆ�j�|m�qGkx��ë#zͤ"<E���e���
��%C,\��B���8Y�_��?	�y���'C�-[卼�t	�1�S9Dr�A�'�vt Qj���5H񢚲$�`Ɋ��$�S�����!�����22�ҽ���VH8��D�O怈vhŒt\h���O��d�Oֹ���?�;��t�C��B�@0��j�PM��1������A��@qF�~�N��@��UZ��IfP��Α7�Q"c�L�R�^��Ò 
��d{c2�'��q�$���q�^xz��I
	�~� 
�'Β����R�����a����#�&�S��y�J]&8V�1����7j����y�^�'�D���K�Q�BЁр�#�y���W�<z1.�&4�̈�P�,�y�KԋZx��̟]�yeO˛�y҉E.3�ֽqlB�X(�@z��W��yroP;���٥G�!��I��N��yr�������N�5,��yR�?@��Q�I��}v��D ��y�Q<O�X1�m�q�,(��I��y�Q8^y��.	fJ�x`g��y�6;9�\R�`H�Z0�t���y�!U�(�$$�&"�5&&����і�y" {\	g�E#��x���E�y"N"$0��u���P��*�ɟ3�y�j�� ϜA:B��
r��>J2����W� :�
G�a\)1R��}I����Zú8yª�-3"n�Hr�C���ȓHN`�9�%P&�9X��B���T��x��iJ���ԕ��NU�l�ȓR��%
�u�����Ş�hȓB��-@��O�$���\�Y��ȓS� T�A=$���gO\r��ȓC��2֧�"[�e�X:�V�ȓchL�!����#��H҅G��<����%kPD�`��d{*�	AM#9,���N�xf��N�������Y����R�ƈb�D��RV�L[m�L/�E�ȓ(�pp�D���)8�*�a�"H�R̅�C�f�`�.F�R�woL8M���S�? "�ؔMҝ8h�숁@&�H�"O�
̆�됡ᓪ�3�ԡU"OJ�q�.�r� ,�e)�Yܭ�C"O�t�� ��A�pIՇ-����e"O��{`$ �dx"���>�:��"O�I�'�C)W��Ѐ�*Z&[�&�Xw"O��2��I
��[���4q��"O~4�e+3,H5YR��y�,��"O�1�pNy�b���U(2�ƉБ"O�)����/�V�5�ı���\M�<Y�Ǝ*!�� ��Zс�H�<�rI��XL�w#�(���K��	G�<9��Q�af�+�!^%EV(KƦE�<ɥ�O�m�1�+�`:� ��FQD�<!`i��CS�hG���a���<A@�L�z\R��&MԚS�@P���YT�<�rlɥ+��S%�6f=:�O�<����U��Ň\`	���V�A_�<�0$"����U;�tԱVB�b�<a1ɜ-@��-YU�������_?��j�/k��O�>�b" 	B`ti�7����Q2U*Ox���Y+.��T(@NL���BԖ>�Ѐ��2����L�~�h��A8(�� ��w5�~��\7YJؑH�$[��h�S.K�V�^D��KF�<1��Γ[Nܻ�DS;`��9���'4��%���O`�q�$����a(�>
��N>��(�<�Oq��	�&OV�z�ޡ9�zm�R\�@����1�اH����M"SΝq5�Y�"�Z<�cKOi�K%���L���g�L50a<����N�(S�̠f(4���Ƈ�+]T�[V\)�	�|�\|��җ��?Q�%�"��8��o=+L�QBI ax��po?/D�'beI��>���#��ǩ���'K���D���rڡ�#o�2��T��y�o�0�b�b>�� ��oܩ�磌3�� � D��c�g�H�z��V�W�/���T�9D����E6�=��բ+d� �$*D�`p$\0n<�F׬|���`�($D�(R������,Jk\�C�L#D����y��`�7%G.6J�9�"D���j��'7f9� G�.S%:Y��3D���������B �
%���,D� 	�H�><Ȣ����AJ0q Qe,D��p��8r �;S��!q�Jm�3)D�,��
D�U2��N�6�&��qB!D��*"
N���eQP�_�ibE�bn$D��4c@�<:N4äƞ�:%"��m0D�D��MÝU�P!{2�\�G�t�A0D�8��c�8a���W4�Lu��b1D��HgF�7ޜ�r�.U�`@%���-D����݌Z�Bx2���;f�!�R�*D��s��[�}��B�D�I��q)D�p2��%�fH�#	H�M�%�4D�8��Q92���#*	l��if� D�J�*ՍO,�8Hac��d�t9��<D��ADî<]������lTt���9D�D���߉Z3�)h�ƂPT��B7D���儋q'&E��gL0�l����4D�d�u�	P��u(bK9�bS�b%D���6��4h$���+G��X]���#D���j̥��!C��_XI��?D������+i�0�{v�,�@I<D��K[�������k����e,D����� �zE�av�O�g2�A���(D� qfC�?/�ЃI҈xh�2�F%D�� f3�K�R�ȝw����UH��'������!}«D�4�� ͘3�8G)C)�y%2}�̳��H�x�(�р�0�'F�(@az>m6MY�_��C�bOlFf1�A>D����,<%"�)p�HZ:\�4���"�tZ��<�DH.B�0��s'5Rٔ�R��TM�<�ǀ��9�,�@�T��V1�Qc��xh(����H�� ����6Z1a��ӣ&�Haa��,\O �t��3��$��>�;W�Y�|b6\�B)ՐY�!���^I� �ݮyT���r���qO�eyT���0|"r�T�s<�2F{��3$d��>)�C�	�i��5:����A����Z�4��&︟p5���M�eM"�gy�m��!�,����c�9��N+�y�"1~1����I#bh�CU��--�0��Cڒ�~�^|)���5yRD9A&oH�x`|u:�	�R������J�(��}ZT������ �X� �����	?�>B���T�cP@�8C$�J�	O�f���@��,шy��r�0��� ;�X� s�(��xB�\L��,�4��\I6Uk���@�ܒ�M3� Ք/����?��톈2�|8%�O4-�Ʃk��!O�A�1脐~Q��OtP&F�j2P��椘�=!��3���ڜ��98�4&���B�V�V>n-)r�,�̐�'�Z�����-.0]1�O��\#�螯/6��$�"̘YJU��
��uO����*�${�X���*m�؃ϟ*���ڷ'HTh���>���I�6ޮ�<)�GO,:W��C��~�h���O��|�ī�>}1�Z�0|��m�S�Ʉ1b�)˶B �e ^�۴isZٰF-�)��3�@8�����(�KƵ-�$���-s'@9�񩑴h;�+��K�y*��.�\��\,l�T}�':<ep�oµ69� u�'9
��͓R�άhf
]��3�'i�=+�ܪ&&�D�������~bJH�pd�`M�5w��xeB�"$-��h�W&N�!��|� �� ��y'��PViL�%���'����<	d���T헒
���*�w����獰�*=P�`��	�85��,��G��5I��T}�X��r�N�i��E�'��T`o���l(��?7�R`;)��e�*O��'O�`ؘ8�7��%+Gp�z��	�w
	��/_� X�9�3��k�p���A�5��)T^�a�ԑ	�t=R���
��F��9f_@��C��@F�!��	X��E��zt*}��h�2g�2�d��
�i�C��
�(q��?�<�d�Ӧ:IVi�!e�t'"h��B׽.�<l���'�L�a�ށO��{��-rrj5��Ƅ<�?�P(̼��'�
��	 d��h�5�H�[`
M�xs �J���'�(�v��*k$�,2f�$Jq֙[�&��&����H���f����X�*�H�o��u�����:J���K��E�T1�cP�&Q�"<��,Z:1�;gg�(;�f@����S8Sx�<qEmʇi�R���e��]3���3T�}�r)Aeɪ�Y��U��x��Jp�ӅB��Hc�/	�g��5BS�K�p�(5Zi�V|���~�<��M�0k�9+��ȗ!tF���M�<�0BI$6BT�A��x�p�"N��E�	<jp��w�nx �R��Jg (�;�>�y��)y�T���8HR���%g��@����,'�!��ʢ~��TC�Ē�g���z�c5手c>h��	]��-���Xd�qOJ�z�!�L��z��_�A��� ���3R�V���S�}^4���� 0�I+g�����Z1J�$�K`k�(U��Lyऔ?l���ED6��P��'�ir��[5��񬃍:Z���f�w�t2UKZO:٪���>�b���~:��'��ɣ�-�2�hO�#l��e�<-O�\�:!�K SF
��T#՗/�y�A��sЬV�:�>Dy+O�qd�X�>j���U/~��\%\�0�
��7E,����U������]1G��a�pM\60�@ CR�<���˳�S�J\f-��i2p�E���d��i�{]�A"KB�|P�ȍ{rHӳ<�Fx��!�"C��=�Sn����'���'n�O���ڦL
$��W�]���� צf8�a��W�.���P͎�@�6li�O1���&iʸIU�zr(9�������, ��MD�u������MK	8� 6�{[DuZu
Yh^�����@#.���?�q���1�� 0�#i.b9P�fKK�<i2�=?�#�*^�Yn�ip���f�`�B�ǂ "��%��B�G-\����	!�"N���hr�����ү��
�̡rBMQ�nV��G I\8�DZ�!d��i%E_:1��p��{�h	w�بAr􄱕�L�qkL<I�+;�\�V��.Xv�Q�O���H�䜚O�ў$���*t���U�=;��?�Q0BS�u�����b

�p��i���v�\5[�p���'�&p�u�Y1}c���N����'G��3��lP���5H�*&q&>�Cc��S�m��� �	��_lfٱ$�ϨBDb5�B"O�H�¯B7r%:E{��w���{�m��n|*u!۴(�0����1���R�^�j�Z�'kxͻ}M�k�:u����d��$�Lx���)/{>1�d��9X��J2"Bc� %���Ԅm&���M_�`�2�sN<�%���FE�O~n��bM�S��l��a�ԥ���?�1%^���D��C��t�'Zܢ)��C�>[(�e dhn@�ȓNS���̈́���ո&���4�$p�OF��uEV)s�H��a:�';���j���0 �X�(�C6�a�ȓ-Y���ҍ�;����� O.���ڎ}��W	<<��S3��-]ily�ԢLu�8�ȓ#��	�򃒐P900C��q�20��	3�<���ޫc:��X��˗^X4��ȓ ����eL�z	���*ʒK�N��Q��Pc$�Ӡelr̛��;�� ��T&6�� ���tǢ<��Eh�R���k�.܉f̜�JuV�2�Ȍ�nLN��ȓ|l�չ㎄7���F&�L����8bl��F��%נ��"��u���;e�9:�Ng�sc"R<o����(D����Ny�M(2�K?&@)h1m;D�,�EkK�Ш@@�K�.��7�:D���U�4��lBC�&t?�b�6D�H㦈�����f	�9\����5D�8J��Y�d�<��̙�KM)�6b.D�4�jГ=�xq�dإy�L�a��+D�`�Ј�f� t��
m��3+D�PK�N�lZxD��A؟{��d�# +D��"�AS�y�Tu%U�X��y�+,D��	� �")`���7q��)�%D�$0�lG	B��5h��Z�1L�LX'D�p�*ֶ@?t$ᢊ� �nB5#D�8)�'0\��D��N�@�� D������mWޙj4���3:\@b"�*D��@Aa�>D�<�QK;j(��H+D�p�CĈ�+^p�`��'.��; �6D�HU�E�W5��ʄ!Hq�~����?D��	�aY�����l�"�p[`*D��+�g����AC�&�>0HV�-D�(z�sƲ��Lۅv9�еn?D��Z���i������8I�T!1D�T�d/١L PU� �~�b�-D���'e-��dE�p� �C�.D�($��7,E+W� pXԩ�e7D��CƠ��>����]5L��u�Q+D�� 0�܈0#Rx)�Ϝ�V��a��>D�$�w�܊!�����k�Tp���7D�X���gN��d���3�*-�`n1D� sd`��<8�Ń:?�.�r�0D�CȈIb�8A�C�p̩�:D�<;���g7�, ��J��ak#/=D��IQ�ڈ5��m�r+/=ЈI��%D��z7�R�[��dc���=<"Y�1D��볨)�j�Y>��Ir;D�Pj�l�"i��&�0N/.����-D��B��^9n�
�`U�[� ' &D�3g�@�&,�b��6����R�/D�x#�a߃z��:ł����#D���Q�R�o,��QE�9�|h�d�?D�L��	� ���ъ��V!F\?D��PG�Q��!�Є 7Tlr ?D�t�n[�A 2�� �6Q[L��L;D�H�T+��A��ĩڪl�$ZB:D�Ԙ�U��%���ܫuV28q��8D�(Q&&� v4(�4�9V��1��;D�� q�Ӥךe�� ʃ�'�r1A"O|���`�� 
 �CB/�|���"O��+$�2f�Dų�.�'!���*s"O^�i ��>0�L���Ɂ�Y�"O:=9DeJ0B�)�NE�,��"O�3U�MzE����k[!!G�h&"Oh=p�G��~־#�+�990B�"O�1s� E�!�Ƥې��U�J� s"O|PH�g˂����BaU6e�N�+�"O
�8��Z�P�b��R%����r"O�� �J�X��6��"���ۇ�~���i]�Mj�����:@� a�D	�!�D�"��ű0/�4��|�%�e�!�%\���1&b&Rw 5���+q�!�$��t�4�����fe�맄C��!�$��C�:py6H\�Dd&awa�D�!���|hnu�t F�QS�t���� �!��I�y�ڍ�0힄)H�{0�!�D���l��EF������!�DL�(�Z�0�ŏ=���JV��Kr!���n$��W�pἑ)4؋fp!��@��h��Μ�6�`m��m�&T!�d�;v��`I�>8����L5OH!�$P�0Ь9E�?ZH�h��F!�C�OD��u�3g������}�!��8gGP�y�F(t��ȴ㜓:X�'�ۓ �ĥѕ�$m���� -ʖ`f4��ɇ0=��o�D "�P�BM�G��1���ԻzĂB䉽C��8��D4��iT�d��B�	a�x�xv�_*�=A�A׶,VB�&x �BщGa�X-�/�4^ZB�I(_vR��b'Ko?V�Q��C�I,lɊX�p`� Ju�v�\�
��B�I,G�t�`PF &x�`��PK���&B�	�#)�@%F�o��g,�*�C�	:]#�K$��EL�r@n�6=
�C�Ɋ�t����[$��)4ň :a�C�
�h�`R�@�v�|���ٙ-:��L؟�Y�g�0A |����(D��i0D�d���)
J-qe�Z���4�0D���AL�&�Mh���h��4���.D�ӱ��5
6A����
HJ5�� "D�<�Vf�I�,|�jP�Fc&i�a!D����Ē�"�Z$��m�:lq��sQ D���4�X��9�S`�O�8s��1D�㇣Sr�,� 2��N������2D�pq2m�<�$i�S��\�����.D�lr�.�N��=�M�2���{ �)D�\҂ř?'D�{��(�ȴ��%D��Q��B71����BK	�X��#D�@��C�5K���K��T]b%�#D�xjd�;�y1M[2"m���=D�$@��ޢ`��+�+�/��꒎.D�8��Ĥ5?\P�g�),Ę貅n2D����˅�2�X8��!e:�x#�g%D�,K�פ)��cĊ�U�Хp�&D��A��^����u�M/0l^*�)D��PV�s`�!wn
"<u��R��'D��@�nΞ+�X����R�2q@�+;D�L� kX0
�>�*�m�	C���.D�\�Àd��h�6�~��Ï)D���eD�+6�d)aʁ6G�^	�6K"D��e�!&��0�2E�:~F9!��*D�Ђ�
[�=d�۲
F�8�!%D�� ^�yF�h�֐y/�5;�2�0�"O a4�sȴ�GHQ�}��ՓP"O&��Pr)�NL�Oz����"O�I���7_�p��$�6`r!��"O���5#�ǂQj4%^�91���"Ojle��)�"��qC�'��A"Oj�#��:.ʝ	b�~�"}�&"O���cN�;R ��D2";�1�u"OJ)���4��X�蔑!B��À"O�A!b(<<͚�!]	1���V"OrxX��.v<|��˝RN~��E
O�6��G�h����:�C�n�&H<!�Q�VȊ�I�&��o��Z�́$g8!���!5:Lؑ ��6,&�\"�!�d��y�I��'4x,ҥ@�$�5:�!��C �`�/حm���m�^�!�D֖r#�d��+ӘF]Sa��!�!���_E���(T7G~�if�Kq!�Y�N,�GEL�Gעx
�Я|7!�D߬=/L@YƁ�*
�:�`���v�!�Č�k����@�Fm������P�t�!�Ϥ�d1��3͚Mp�g�Y�!�D�9C����&\�9�~��f�A�-!��!p���d_A.��aÔ;v !���j���s�E6��i+ra^r�!��ƿ�2�Sol�J��f�!�T� �	a fڮK�I�G��n!�Y2(�e���KN�+]�jh!���<��-!k
�~�Ӳ�'Y>!�d�r�ԉY�H��`�@��=!�d�.$��aY�v����2�)H�!�d�%D2 ������y��'OG!�d�++{�\�A�8�j�7�(r<!�dX 3���rn�rm�R�55!�Ā1r��{Q�^�ZTe�`��<;!�D<f��YӴ�;@R�	���i2!�X�n��xp7gؚq����i�!�$E9���&")�2Ec��R�.|!�D"2� QD��~b`�`l�3�!�䊹d��A��AI= |x�X嬟�]�!�$�$Lo�{��Z2u@�a�]!v�!���<NF��.��?����$�4)!��@<��d���Z�k�°15��T�!�ĄO��Q1qFڀ5��B 'M�e�!�Bk^=p��"�fR�%�*!�d��7�vUI�$Ⱦ@�rI�pgpL!��
}�����(d���T�1V:!�$�*jh��QC�]�l�3�K�B!�D2cX���B���A��a{��=!�$���H�	�-u�Ѝڥ�G.7!�M�9pȐZE	�ʉ����-!�:@��l��I�+%kLd���D =!�$��M��ݛ1)��u{���%��":!�䟋f����#CW�o>Ekc%Ga9!�5<�6��GEF�c�PD�daM�*!��րn�����c�2�59�'І�V���\N���d���,N�j	�'b`Ѯw�<i�,�N��z�#D�(��Mȥp��):�]�S(.D��Q%��.y��I��xղeBf�,D����ϣ\�,�y 'Z�`��)��*D���p&�X�z� �Wx����>D���1` �S�%�1(>r��e:�e)D��Ԣ�2�z�ig &~6�C�"D�� �X��߂�
��N3U�0��g"O��
��Y�?K������B��R"Ol��e��ov��b�P�����f"O��R`ʡN���1�%9l�hKD"O��31�Z`A1C��ig>�B�"O�yǤ�+�.X@�虢eV���B"OX�qE-��hn2�0�h�H3�0��"O���C��-ش�k�瞴w���t"O�0��Hl� ;�#5�6I��"O��Y�A�4�����S�3A�"O��� �Q�8��c�AA�[^�5��"O$��E�c6���:!��j"O�L���O|^,��CA�<Q:���U"O�` �I�79�pY����o�L�w"O��#LE6P����1�>O����"O��+��U�
��EAc��n��E�v"ONlѳ�;ռe�@A-u���U"O���$�B�A�88��#ʉs""OL�q�NB��d(�iZv����""ON��� =�ţ��6e���)�"O�P�玘
FPp����C��&"O���6쒞i{5�ۙ!1�PZv"OL�ٖ":N�>Iڒ�3/�BX�R"O�`:�o�$
�`cl�,l��@�"OpE���˶q�<��[%����"O�\3v�קI���Ф  2[�
%`g"O��A��ʰ=�(�`'��kb��)C"O�e؀GO�!�ܓ��:��ԣ�"Ol��¢�^���IȦU9�Ɉ�"OX�"P��B;��bH�22�Q"OZ�� F��mY�'	��+c�%�y��DdV��6$'rm�U���y��ثҬi("�"�	�u썟�y�d�6&B����֢G�zm�$ϊ��y�J�\��e�qf�hO`�K�
��yB��fb 9b#ě�[P	��n\(�y��&`SȬ���Y4is�_��yr���R����J״�3$ɋ��y�X$b}&�P����w�x��c1���P,Q�4��+��(���ȓWb8&�*��b��.�L��U�ZK�<����B4�X�G Bp�������H�<�&�?���i%n�5-K�(���KG�<��Ӄq*\��3ȋ0w�h�##��A�<�戝;r�IQ%Ñ9�,�s���T�<ф�Lv�R��W&�6k~4C�R�<9��C�ܔ(v�3� ͘r�<��J�`䝛�'պl*�"�ET�<9 ��[ֈPA$LH�"�>��š\x�<�0%�e�=PK-B�Buzf�m�<1 �S�}e�B�Оe�YZ�A�<y�/9+�`��5-ZjU2�)��Q�<� P�����OT�,DanKb�<)�E�&[�,B��Y�[Q��  �AD�<���)I>�U��N�})��hǀ�X�<9%灺<�J�K�f�8E�i�Ԯ�Q�<�pg�;>�:�#�].�a��"�O�<i�C�P��� ϫc���@NT�<y���%X�QC�2#�6�;s�J�<�+V�J	�� (x��S��TF�<Y�n��6��2,#p� �G(SE�<�5aKJ�Rp�"���>��d��c�K�<�Mh�ph@���	k�2X;���C�<ɲ@�������]�9+֯G�<� �����:5��S��%y�(=��"O����k�1 ��-XW���0�¡"O4=���E�0ݑBg�8�$"O�Bv�U:4r�`rU�K6��X�"O�Mp7 � �<	C���]��)��"O� C��� W�tt9��W'T��"O�ȫ��Y%h �R ��,�Zظ6"OL��ǵUXTI2\�!�~�:�"OށraQ+(>����K-���F"OĨ�砙�e~x2�$Zz�x�3 "O�]�U$Y��
M*@�,��c6"O��Ҡ�	�t|������ƨa�"O"�X��\K�z̈� �7�8	�"O$�&���N"1ROK�l�v%�V"O�<�Ӎ�(YK�5=tr]aqJ^��y�@���찥��3���4�y�F��xa��D�<)�P��R����y����mĦ���iL� ��{���<�y�㈍Q���A��_�&����-�y"O��'��ѣ�$��*���/�y�c�*n@*�K`l�1���be´�y�!
���<��ʗ�ʎ)��,���yB�L�S��Av��"!��4��6�y�-	�=�K��V��{��y��#. 訳�&%B�[׫߃�y2�K��Rc��8Zf��˷���y���J����F]�Bq���'W;�yB� w������R�$!�s��y���)���Y�M5QL�s�n��y2(O[�ލ9Tc��2���R�R�y�b˴a�ʙ�'*��@w4�;G�˜�y�
1�Lb6�J�:����Va�<�yB@�<w=\b��3����쒗�yr`ĘHH�ñ�/E�顥L��y�� ]�d�օΐ#�hm�U*L'�y�oS�x��5���^j��7�y�o�*�:�B�ݰ!��j�b���yiӏM	$)�
[�QP�����y2��h 
l��G{�	�2B�7�y"$�0�"�J���m�����O��y"���T[�)���[�l���PG	�yBfƙ���x�A
*T,�� ��y�G�+n�M�k�b�F+�jV<�y"!S`���X��T"_"�X�F�yB&8#"4��b��
�N�/g��Ņ�1�f�Zƭ9y��܁$�H�A�v���~Ԓ���:��`	�ş�God��A��;�W�B��1�̯7�����z��V�ۭh@\���.j����)�����P3��b�
֎c-�$�ȓ��T����`� �����x.��
]8��`GJB=0��&͢M�ȓ[y�)I����:K�5���85&Ą�Y<�-��������WN-}U��2���a�(X�����N����:��ۥAɉJ�N��O΢�(��k`n�i�#UF��@g"���GRzزS��I�^�8�+��s���ȓ������,!��RT���@�08�ȓ�j�"����@�ɱC�N�P��X��)�D ���61*VQA&��A��ȓ}{�M	g.O�Q��(�ͅ ~�i�ȓD�@S��	:C>�uo��r�ȓ^S�9P#װ(�N�H�� �t�h1��S�? �a82Z#]�lХ�K����	"ONm�q��9ɼY���P".����"O�Њ�ec���#J�/H6Hmؕ"O����:neA���*�8�W"O8 �7ÄY�I�j�4$�Щ""O�	�E@�K�|��G�8Y��"O����ǮS���Av�͒3s����"O$��#G5R��Q��^!`�`Z"O�YE�##������&RQ���3"O �[�CU�^���4�υ17fТ""O$��mZ�i�&M���)r�D���"O�1MU��m���jw8Y9F"O����#ݏT|��/��R��驡"O
<JƨʓQ�z�:���,!=@A"Od��#�Z4��C7�!,�;�"O��MȦq��9��ARJ��h�"O:�(�	�R|�y�f�!|�4�z6"O�����!�0=��œ?�`D3s"O�D۱��?Kapi��σ��|8�r"O�ea��R�6N�٪b��vc�]i�"O�̡�1&"�
���t�s�"O����$	�jJ&h���L2��4	�"O|9Z��MQl��jֆq͖P�W"O4�Y�� ��|������ȑ "O� ��#��*/�L��̫PRԤ��"O��"��
\�uZ&d�>���D"O�mcDHR�͙��׼`�Ę[""O`��4�ΞI���Sa�&��<Y3"O� ��˙qb��@ŕZ4�E*�"O��W�Ԏ� ��b��1V�8a"O�|T�D�
�UĀ� 6����"O$��Ө�2d��i�A�-��x�"O�U"@�;|�R�P�Ȃz���#"O�9k��\�vl~�(%�iah��"On�3��@�n"6�Dk4�\ڴ"Oع��l%5U�Mk��..=���&�I}�O�͊R#^Ŋ�C�a(CH���+O���$ ����b���UﬠU	�*9[!�dT�0QVY�3k�[/��01�MU�!�d�)}+fD�t؇+�!@�R��O>��F+�8�
%B��Ձs���""O��Siѳ`~��k��!Z���"OF��D�֤:�q@s-�#Z=��r�"O�r�"�H�(���k�Z6��c��'��D��H� �xИ��	?"�8�PI'D��b�`@T4@0t�̑��{��"D�`�c�س8L����E}�M�3D�0"��ݺJ�8`j�(IoR�k�I1D�\��N 
l���$��L�5{F@,D�<)veX��u��ŗ1+v�-%��&�Sܧ/��#�!�2��(��F?��1�ȓ(�|DҔ�ݙt� ѦЃѢ>D��x֭G@��qW/��h�x!p>D�t�檔Q,��ht
��E�f�y��;D�|�b��3X"��`B�c�V�YŦ;D� 9dFȆ]�0�S��1X�T��uD/D�H����gԶ��h�=;m�Q�<Q�%@^����μM� �3�Ny�N����QyR+� �[�H҄FL:\�U+L�
!�?=�a��oAS/ԉg���!�$���I3��O["Мز2T �'2ў�>�"��D���3C�������8D��p�F�1[0Ja�Ǣۀ:��5�5D��DX�FBz����1=Ԓ�­<q���3� �i���O� ��1�$��7Ê�Ö"O��w��dpp���L���"O�����**�y�unƖH�����'��I�<���	B� ���DU�� �N�<ÀB�p��x�gʇ-���"4�N�<ٳđ;�|�� �C�,n��jQ��M�<�tgM?p��@(�+��T��a
�'�G�<a1b��A�b�(�X7Cl$Ԩ��x�'�ax"�؝g&��D� c��EX�!W�hO���	��z�l��kH�W�~�Kg�̔��=)�yB��'���ctƅ�T�"�-�yRj�*em�ؙRm�6/+�a 2�� �y2#e-n�	Vu�X����y"CУ�
	0f��P�અ��y򏗞-v"`k� �6@͒�Isf��?A
�'���Z싫8mҐ�ጅ�f\;.O���hO�J�aJ6kQ-��!�ŀ�6�<%��Fz}��nH�zc %p�߹;�Q��,��(�Vƕ�r���I�bӲU։�ȓ0F��p��,���b��}��H�ȓ\���� �Z�)��ӡ��}��8r44���?Z��yԮ�G[P	�'�ў�|�F���j�C�$_�'IҹI�
m��@Γ:Q��� �s��8�T쒦6�Ox�Y>��F������e�*LtȄȓphaZ�F'=F�Cq��*�ʡ��w���k6hѕ6?:�J�PB�܆ȓ:D��	�I�N2v�(�ڔ's��F{��'XV��Aɧw-D�Xp',&���'�N<s��V�2:V���n�uV��R�'��#�"-��Qh��@��f�K�' ����/����Ԯ�>l8 D0.O��=E�d*�[���J�t�kH�yF��y��bmE�WU��b�]��y"�	k�P�o�f;Π(��P����?1ӓ4Q��!B�/~��j1�	q܆1�ȓdh�	RU��P����ahJy����9��#�M�,�e�&��ȓW><�H�g�<��d�fj�848���ȓ�.��.ǤT�j�:K�_ӈ���'��ɄC�#c��|�&韵X��9��#~��v�UU�8�pG�&����	l�'q`HQ��*	 ��C�Q.�Nx��'+��gi	���#���qF�X����ɔO:��"EƸ �+�K��v�q�'&����g���y����V:���x��x����,
�	^��Ɓ2�yBh�v�>��� |b|�@��W��y����Qj����O�k�L�d�0����d �S��% ��1!W9���8��D�<�ުOM����@�N�i��k�A�',ax"��<Ў)��ʑ!��#�"��y"/�b�NU��-*��6����y"�]W�ap0�T�f��M1zC!�K-Nu0d��|�b��'��J!��׎���0m�W������ZI!�^�ԉ�c��	Z�*��Z=i��O��=!�OX�0��C��X�1�W8*���"O�tx��5rc�U�V♣d���E"O�i:�*�c���BU/p�P�W"O`�`�E 8Cjp��W�y�.��"O.i;�\�	�L���9䎌�"O&�)f�V$�X:��&a�R%R�"O�e���%rd�:f	�GmF(�1�'W�)� R�j ��fM�أCנRZ"!r��q�����1w�`�Y"�X�c0�D��B)D��)�¢�.Tx�'T'q���ū&D�(C�J�H��@c��v*d4A@�0D��i碏7d�XCκW�!�� ;D�Q3�A8fkz���f%����,7D�l���O�D�"y�dÃ9��Y	�C?D���u��
`�Je�3-ƊA���ȳh=D� �F�'Rą2F�s׌AC�1D��1eD�4��6�C�/ʞ��&�!D�$�TC�K��H�#@�mZ��#c D�ȓ!��?�l)�so��h-�sb3D��hCKܻbilm@ �Y�X�P!�ׂ$D�$
�5V��	��MY�9d&����!4�x�c�/`n]���%�@��3�ZA�<q��}���3��"zB,�a	 V�<Yɝ�8�TD���ˈ*�tcsJWO�<H�7���$X� ����LN�<�Rl��J�l�×�P%B0i���OK�<iG靮MI.��%�'xW����/�ß(�?���I43I�I0Z�Pi�3�ѣ��C�I�N.\x�� ��-� )��� ��C�	:Y��pG[*>�>}�PGW����7�e����߽\�"�'Ѯ��ȓ^��=���J,�$��P.�l��7` BVf]�I����$/H?�����o,��I�N�H8}���OQ<��8{���6
ڱM�P eK4$��ņȓƀ)���Sgi�b'�`.�	�'a~bJ��O�5sP̍Xj漰���yr/�Y��E"�	���z�Ď�y���;(�����|�4�����y"�^.��`���rI@}��6D��y +�0��5	��(�8�5D���'��1��-�$�
m��1|ODb���w$��9�\�#��n��B�"D��c!��:�����f:>�� )�b�O�=E���T�h�Niz��M5x���a��B�!�!�a� �	o�E���	�;�!��V�ڒNQ�X�tQ�o>�!��Lm�xe���	m��R����d�!�drǐ��7`Q Q$*8w�G?h�!��LZЀ��g��-��7�-7o�O����
���fɿ7Al�k!u��ͳ#"O���ө���j��P��(���"O29YWh�E~�	�H�%K6)"G"OL���E�q^EI��^�}X� �"OR�@���Z�VA�e٢+*�"O��A���)\,�E��f?}�+�%�y��U�*ӆ����* �M��Ό=�yT�.�p���A�l[v�S��y2���sg� ����"ar�H�H���yr	W�u���ja�F�p$\`b�K	��y�؀)l�#�g�։�f��y"��YJ�Iȇ���v:>�x�'��y"dY}[qO�2F� �E��)��x�%͟�8%
��՗:҄ЊP)�<!�̪P,ȶ.CB��Ũ�rџ<�	xy��?���C�^��xH6!�-��)�E�=D���vD�~#Z��0cS�`
��4�>D�h�UHT�T
��.Q�Fy��FZ7�!�d�.~�-�����@ 9�@��(k�!��<c�>��g�d<\�B�@ܐv�!�d��r;A��њa!"�30ꒋP����7�g?� ��ꖤ�-x�v��f�2l8�	��"OD\8��K�BH���/,�01"OL�S�INC�X	���H/� �٤"O���A%~��!I&&��IR"O��H�Jč&� %!2�Ƕ4˸�h"O8�!"
jA�WDך*��7"OJ�0���K��,���ݐ%�iY1"O��i�Q�2I����F��>��g"O�|sP�
:e�X�p�Q�Ot��Z"O�-C���`��Ȑ���9g49��"OT�ӠM���|�* R�8�G"O�+�".Y\�E Qo��4��"O��X6O��`W���Eѥ��y)�"O� D�X���C�B
6��f�'m!��K�c��j�@)wȮy V/�!�$��O2����A׈W4��խ
�!��;N���τ�Q,&� K�r�!�$J'?�x��E֥:�(S��
y!��=e���Q���r��ԋ�ٜnY!��[��\H&��|����� yU!��
X���&GƸX�0���ꞛHG!�dV�Pՠ�!��[<8�*���)=!�Ò"x���%$G�	(ҧ&V!�L���U�"�//ʁ%E[-F6!�L.W^�� @�
�f5
�F�>"!�D764���ea�1r߰!���!!򤋆V"�p:��Ɗ��P���_��D�^����7��*�Հ6�V,��C�	7wJݠBIܑU\UA ʽ;����:rk�T���`�F@
�T53оɅȓ|n��������n>f`�Hp�'��Y�tS<M�H�#$C1`jd��'-� ���_���e�q�1��̃�''��(4�3���I�k��l!
�'�m�����V`��:�Ȏf��p���hO?A�#��E@����"�j͒7��k�'�a�4IZ�((`�yV�YŎ��y��A���Jd��;h�$��J)�y��7g	N݊��W�r�X��u

=�y2 ��?�R�S�b��d�Ԑ
���y��Z����`�� `���E��yM�3}8t"��$ǲ ��U��hOf�?!�+��*�<uZ!m�6tZ����F��=1�y�c��^����,�n��A����y���U2dx�'R�a��1�qkV�y�%�2Nƍ���O�F�8��GD��y��!;���c +�*<0���y2�Aoi
�Xd��'8NlaGH$�yBÅ�|f.�`"/Q��D�v� ��D,�S�OS���K�I?ju��B��`N��N>Ɉ����k�H��GD9J�lc�ɟ{�!�dD�x��ULNCk���hI�y�!�����`�ǯA#6_��Q��*�!򄆉w�xH	�N�Rf��I ���!��)�
�i��)AH.8RA�ͷp*!�;|����R8��2�N0F0!�RZ����Ѐəu�ؙlJ�d�Dʓ�hOQ>q�0)�>!3\�2��y.zp
�!.D�Đ�ǚ;���^2�Y��Oέk!�dĚ(�@�C䗕(�~A��m�2o3!�P�4���P*�D8P#*O�:2!��U!{c��; !�[L�$�Z!�CgO̍�g��iL0�ї�_�!򤒯#O����ɍ�aЁQ!eD�\�!�� ��y�Jw(���W4l���"O���duP��g��o��3"Op��֢{'l1"�C75OV��"O�Q3"d��&��-
��ɸKB�@"O�P�bn�3�kď�LNY�"O�E+6�{+���OH9ьtp_�$E{����3h�$��v��R�T���A�e�!��hL(�SBZXX�!�q[]!�d�>8�}���٬&Tf�:v��CT!��h�>���y9���3!�.J4!�DU�S ,�gЩA}z a�OM�!�dV�\�P��E\5 a<$phW�%~!�*4��x�F�!.%�(�%@��=y�{��$�'
LI�[=�\,
%m�7F��}R��h�h��J�4x��A�\�ru��6D����Ρ,�����-'H�y�j D����i
y>B��e��6؊с#D��n��%S���%���G�C䉉d<<��i+.���A ��C�>D��a��tP�Ag�2�tC��/l�LX�5.��9�Bt!@VUO�D%��o�O��DLGޠ�a@�zPI@ש,w�!�䙻>[NysT
֭dd5�Xr�B�'�N��	�f���b�:L���9�'瘠a�C?^��a2cD�?F�6 �'E��A�ځ�����*�p�z}z
�'oR���& 0e�䳅A��;6��	���?Av�ݵ+d����"B�U*�pȲ@��y�eю^�÷�7@����A�ע�y�U�܅#t!=��%�Р��y©��7��p���-�4pw�!�y"�%�*e��HĘ+%T\{��I��y��H�(�(�f�R!)���"�ye�l���`,�}u�yࠟ �yb6�
 	v��	�e�'�(�y���
��`ܐ+*`�%]9�y���2�4P!�<?��Z�h��y��J244�A�߼��	��8�y2�@�L���p��3�>l�U���Pyr�`Ć��Ab��T�dEC��M�<Q�\�2 (�ۻ&�#6��M�<	��Eo��X00#^�y�䔺�� F�<�ĬA(� �q/��r� ��u̇V�<I��_�A��1 ��B�l�8�fV�<�s�L�(e;�JC���P��U�<����8YϢ�RpB��v�}�1-y�<�w��-�B9��#��v�r��cny�<Y���ԅ�a,P�.#�QY��r��t���O��=����J���ĕ?q�d�
�'�NѸ�"���6�RFeF�lX
�'X�����<vB��"�ƉH��	�'w� 9�KZ�W���0�!:�֩K�'�4:�$�D܍#��1���a
�'��hkbAGbʸt���	�'��8B�'��8�b �H 0Y@��H��T�O>��G�y����06�2�����@(^%�?!���~�2I�9W�=��âx�B! �*G�<�3+&b��ʴ��� �+��K�<�cC|WN\�#mU@�wB�]�<��@�D�1{� ��,R#�[�<q2mP�[3��".�':��	�J]px�PEx�`���r1��G#M�J�V�X!�y�X��,D*5�A%R��Ik�.�yb�̀���;AeIBFj`���.�y
� @,cF��A��lv`��b	���"O4e��	E@q�)+����V�x�"O���<��!JPh J(�mjd�Id�4�㮞0+WXɫ0�A�ut���#D��Ӏ��8&�$�*��ۜlb�9�$)"D�t�AH�7�,�3A#�}�0�!�$)�S�'>�"��T�һ?Ӝ+��µ{؄Y��;���GԻn��	˰ʄ�<**�����MS�l�M8$�R��Y@)��S�C���8J@Pa�b0��ȓ��C�lZ�7+je8Q�;Nu�I�ȓO�j�ߡ&'���Uf�7n{�1�ȓ=c.|��D�%h��
`e�)4c��ȓ��P��t��FeX%
�$h��R�M �K�=qȨdq߼!��)�ȓiN04p� �:UXN@�⍙8<�T4��T&d(�0#X̶,��%�4a���F{��'��D��)
�]�'e��f�����'
�<�c H�P�������@�x�'RP-`�'<Ŝ�����[�Vɛ�'��@��nմ0�� K�i�0hJ
�'��`ca�A7<Mr���.b�����'��H���V�)z�e�b\�^EQ�'
�q'Q�D����Q�֒_K�#�'��h�f����@ �M�^,ta �'�ޤ�V�C�?a~(y1눈@:&	(ߓ��'0�1%�i��ѱ0�+
�p��'\�ukW'�d��� �&ny��'���΢Pt𥱆'�����'I��S`�A,�<����:d�Ƶ�'7����
� Q%�Ģ��	/������3�-@�T�#�0gR�ʥ�B�k4,�ȓA�H5#ɩz�*�b��e����D0�!a�"�~=���L26��<�ȓd�`[�N� Y
��R| %E{��'��0����.tF�j�h�hP=	�'��aa�J��B=0�R�M@~,a3�'��r�:ut�i��~���-O�ʓ��S�O�B��C��<�p���//v��9��'\��S��E�c1�9�%-T�fS<���'�t�BT�p؁��[�kј�"�'o��I��I"��A]8r�6aq
�'U2��g)�('�2�3O*�24:
�'+�p���ƺ=���I�o�%��:	�'�n���L�+H8	�ѩy� �'�R�:$�
,�����9_xx�'�:Q0�∡!Ch�a������
�'��u�3��u�|sEPw2$�c
�'�|Pj��,�������"�DajH>Y����1�%�ԕ`#��ae�� ���	�'RZ�C@M3V!�����.�j	�'Pq��I lJћ�G��d Եe"On��3��!#��@�0��
-�P�6"OD KW�G�B��i6��"g�-(S"O�,22J�*p�ZA�
��>�l��"O�Q	�ҸEa��J�	��&!h�'F�'��)�3}�'C5g�Y��:n�&��u���y�lG�*�fK0C�8Sp6d�uG�y�g�
��Tр�6L\l�@D�T��y��Vc�$TC	��a�@c!�y"��Hbyy��= ޱ��*�1�yR(%� �pE�	0zr|a:vdZ�yYh�)���qiU{E��6�?A���4DH���E3a�Ba�
¨.��T��S�? lu�V/�#:\5�6��Jn���#"OU�QL�&���q��.tc�D�F�'��'f�)�3}��9�l9���џ��LB�yb h3ȋ����.�3CB,�y/��B�jH�
H
x���7 ��y��)|q4X��n��k'�Z(�?	���>C�X(���4x��/ɌD��t��IPV)W4F�� �v��7q$�ȓl
�w�_��v%��jW�T~Ņ�9�H�%"p�ܐCcF�!V(�y�ȓ#�t�3�j��;�$R#x�����j(1���F�&j�U
Fgќ֒Y�ȓo,���#�	"�X1�T4`Ą�L	�E��A�r�0� �ȓ'�H��˛w~���L��	[dՅȓ���䛼p[b��G�IG���ȓY�\Y���F�e�>�SNu8<�ȓG�͊��#P|{wʘN`ńȓK?���R 	%�b�PQ"Ň![R-�ȓ;>���4��qp���(�+`�29�ȓ�*h4���(��P��+8YB��ȓ@����!�
J��sa�L"���ȓZ�t��K&?��*�üE��ͅ�J�m�H@�6��Y���=^O���t��RRo�3_���b��
9(>ɆȓDO����̺eT�"M���ȱ�ȓwB��QN�Mj5r!�F�=��e��5.�8�L� ^�>�!��KS=���B�,%�5� "ZV�r�]�q��X��ma�Yj'���c��E� �ȓ?̼��B$ѿM�P�j'NB?E4R�ȓǰ��5��^l�I��;3k�Іȓ<0��φ�{&hꂀIf��dFR�|b�?�KA.Ҏ�z�ۀ�N�hw���D1D���3�ه��3C��9�����#D� C���0�V`H�sO���4D�4 �h�-kANl˧�:$���S�?|O�b�<�rc�5�"�@�s���`1�>D�h[ŕ-n?�9�2ID3��X���=D����>K��d�+ϥk@��9ԫ:D�xi"m��`q,�r �I�(�n�
A%7D����U3e<	���_~ju��%6D� K!�!JV~��v�D#0��M'D��@Q��/�H��
("i۳G$��0|�# Z�-��%��� ��:be,�c��y��ߘm��<+���0i�M�f�?D��kf��$L�J9�u����a[uN0D�8k��o,�ɳ�9	Tv}R�.D���c RA��It���
2���F8D� ��J�|���� I+\��(3D�  b��I���cZ� T���0D�ؚ䦇�^�Dp����G�B�b#�/D�4��[*��\�g/�5G60�d!D��z��A�\O��Ç�V�����?D�������M�Q�5�o���9��;�2�O+R�	�f�ቕ'5,Ĉ�I�"OXy�*�2��s�h�	1��屲"Oژ����a�1;P�ÐG���CV�'^�L���M�Ќ �d޾S���C'�OzC�I�QҸXfρ�vX��׫�B�I	I3X�Z��Б�PԸ�聲(`B�ɺV7�Q�Z�Y�P(�mޱ=�B�ɱ��Mr��T�7���B��>��B�ɻK"4�bbᚵ�l���팡H��C�)� �5��f�^�t���E8��!�"O� �$�B�L)DH����p����D(LOzLzW$�z���)�h�
DA�-��"O2'�K�Z�b��c�l-��"O��
 �һ$��e:jH�9�"O�9�1�O����cd_����"O�� m_�+(�P!I�~�B�#D"O�9J�	���Hq�ɒJ�VhI�"O|�P�כ{�	q��D=^�@UZ`�|��)]����	(ľ18���	Iv�C�I]ݪ� AIяjM�Ux��N�=[�C�I�F��$*����r�IćPQ�Ѕ�w�I�1�ưon-��d�3.q4C�ɞlʤ(����b��|�q�I5�C�I)hw<š�XS׌�P$�
�C�C䉅X>�'��JM�S�ܠm�C䉓x�xxZ��G�K?��e�>E�TC�	$C�5QU��^�K@��~�$C��%
�rY�5Ô�/`&Y�r���tlC�1���CAY��ZԊ�k��H�4C�I"��s�� ,�&�ƣw�0C��JC|`��Z-c����G���(C�	�cl$J��)W��A��j��C�G����Q�,hLd&ڣ"��C�	3_"��
�����e	F*Һ:_�C�	�\.�*f���<|�r�k��f0�C䉳, Z��4��g�ms#k��d^�C�ɾ4�^�1-q!'�֑i.��=D�؋�b�0NP(ԝi�H�e�9D� y�L��<w�$KD&R�|�`aЧ�O��=E�$L� Ia�����Ҫq�vQ#SA�H�!���5I�TY��HO&���jf��0�!�, d�}13oH?�%(�?3�~a��'�R]�shًKtdB3����'����.�9W�-�䠊�|�U��'�T�� ŗ�D$n�y�&�~��)��' 6ELĕi��0XaoK.V �!�������>���ݢ�F�P��;;( ���$\�<���z�B�p�*��M��A��*�Y�<1c"&�N�P�H�zk��#@�V�<Y�_g�6�i�,R!$���gV�<�pJ���,pq�c4��srjQR�<�� ��^d���$��v��N�<��8r�a8���
d^�� M�<!�)
�>�ٺf)I�st�q2p̝a�<i3φ�9=p���&E���bW[�<)"խf�d`3m��u �8j��\�<�g윇��Q	����*z��Bp�<����~2�\���q�T��Ad�<y��ؔc��P����	Մ��q�\�<��IN=c�д������xt ���M�<Q�L�3�渀UL�>� E�P� A�<���^��h�B�%A<��d�L{�<�S�:b=VU��.F�>�°I�B�t�<������QW�#�ZT�4�s�<Idg��	��I�˃YӒY��F�<AVBP�F��e+��v�h�x6�Ax�<�qj)L�$�s

�❘��w�<1�����!�3d�4��x��k�<IS��8���3	�u�4Q��+h�<Y�G	���d&Ap��80O]�<���W�,5\��u��<���#6��Y�<��ǅ�FݦI;$�U�QJ`N�I�<AB��+$�zW_GZ� �6MKCh<	
� pi�#I#o'���s�+S��p7"OH��痒X��If_���z�"OH��j� IX���IzKde�"O~d��Ǝ`Q��`Qe��f����P"O2��7g07"@���Zh�"O�P�"�@6M��pӣ�'q`��v"O��#v��> �x$����v!��"O��(���=ܰ)F����4̩�"O�0�b�t�l��e�>�.}[�"Op)z5��9J�,��'(�:&pAڇ"O��`e矑M
�t��26Z-�B"Or��_�`lR�(�'�PǦ	e"O"�pU������� .B�"O��Qcԕ~Y�h�֯�jn"ON��uK�dafX���/LĆ�6"O�D� 	q���y�_�4�� �a"O*��c��0s�t˳���Y��ܓ�"OХ��ƍn�(m)p�y�֙i�"Ofu������8psrmG�H}d�"Oj��gC�~�bL���%tʐ�$"O&Y�e��5+TPs��-nb :�"OZ��a�\+za��I�I�/Ya � v"OBՃ2�^�}�I���H�	� "O�m"qd�j]P�Mǃ��kq"O.\��HF�]Hf��7lA�ce��`c��#LO4:�ZI��d�qjݧ$fp��"O�)#��S�h/~�s��A�X�"Oz���P
��)�#�;(_�P�"O2��*Z��z�1!�.Q�H@"O����Ic����B	5�jS�>D���/����+-d=�@=<O^"<����.(y��-�9��Q�G�u�<�eA�<�p��範�1ZX{A	�z�<��a֋���3��(�d�J�b�<���ȃ ��q�bC�*(����o�g�<�5�fe6I�3�P"#�Qe�a�<)��ɶ,D\
�g��bA$_R�<1b ^<�~xqP�؃o\x�2'D�d�<����,�p�J�	_4���A`�<i��Vp��8�5%7NN��U�^�<�p�%i��wIBYɒ�QT �]�<qա�T�)rU��?�t���h�A�<Y`�Y�.��|�@YH:�%1�JX�<�b���h�f�;A��D	��8�EH�<�I� +2�yC�''Zbu�J }�<�u��i*�b��ϸg�.!�'|�<�� ѼG��2�B�.���G�<��HM&@���I�%(�xC��Is�<A�̀?��\ a�)R�
|��k�<Q�,
2CCv���V�/�H��iM�<�r���0N���*ʙP�{�HBd�<1�-�><p��Zv�ޕ{�|%
�a�<���g���f�1P�$�Ǉ�[�<6���EY��j�^�4�h�y��|�<���8�቉�Q�M��	�`�<��'ӿo:QS�	�|�35K<T��Ң�չr�D��#�i�z�`��?D�X�ʣ	��=���\�<}�b�=D��jD9W��B$�N-`�&��!A=D�\j'�B�"�AhvL	= �Y�ь9D�9�"�.]��3u�L������<D��*�X��DI���9eʌ��Q�%D���S�2�H�@��\���(���7D�컦�R�*�Z5�s(�>Y[f���"D�� �Yuo[�I3������Q0�"O�\"�k	�C����D[l����"O���ĥ3�� r�E�>!�J�"O��2��<7Qv�!�MS+t�t��"O^u�E��'i�� #G�1��T�1D�0zē�zx ͜#�����;D�� ��H�8��cͯB� D�T*4D�T&'�R+���L�
�����3D�p��M'T|覇	�PnDiai'D��I�M��3�deꅉ%u\\z��&D�X[��Z�PQkwc��/���/1D���6��x�R�7%���gM:D��(��䐭4a�
Y�pM�0�;D���uM�G���C�P$XnA�� ;D���D(#F�PA��L:�^11..D���F�#�R���	S���q���-D�l��͊U^PD�g�΅R�R���!+D�d���	k&�TB��xB ]S��(D������)=p`T�ۮ���{�9D��ґ[�W1*[�N�&��Lh�	;D�T���\/3�֘P�I�V"p�kӨ$D��bn�<Ry����p�d��2e"D�bs�ǀ>钄peg\?P���=D�lX𡛢�n�i$J]z"A{�):D� �K�m��%x�\�0�EJ&=D��dΠ�.��,(X�2!+:D� 8���E����(J�M�e8D���o[�XK�a�!��d��,IC4D��{PFM,�B��I����>D�h�LY�G��p�%`�Je@a2R�;D���7��w>���ȵs��tZ�9D���#A�u�����4OQ��Xr�*D����� ��̐�LC�#�l� U�)D�H[B
ϛK����F�B�8�����%D��+s���3��8�P����#D�8��
1
�d�S�&`*0�&D�@�1d͜6\ddZ�]:��K��$D���@��شa�C���"cm/D�(���ڌ~��uPF��w�`L�3m#D�Dp�+���eek�+�H�b�%D�����{�v@�c��
(�S�J(D�XD#+_�5���H s��U��)D�Ѓ�B�&��UHH���H�
+D�P��/U�h�]���!x�x��N)D�8�&@ל��#j	Y��t��G)D�$+2a��M��`Q�F�
HDM+V)-D��8�
]�ZM�$'F'�;�o�<i7�V���S�,�u8�KAT�<Y��rt�1��L�\Y���J�<	ai��<t�T"�ŌA�����AI�<�*�,�����+�&8q!a�<�։R#�N]`�FL.�(� B�A�<94BK�2��R�	�"��1��B�<A� `d,h
�D<Y4��5��U�<�E�/y��5��2Y�r�!2�FO�<���F��ʆJ�t��w�E�<�t�X�\������*P"���Az�<	�n�/mT0����UZ,����m�<Qu���e��4���,B�KVh�<ѵ�<a n��0���A�˞f�<)wÏ.$b�hD7I���a�e�K�<U�#��@!�Y52�0đRoJ@�<����:��[2H$0�"�<9$�ϻi:�Q�ðlr	$C`�<� �K$jS0S��t��NX�@
�"OP8�f)x{��;�
�:y�����"O��T�8M��5��DD ��"OzD8aM��hb���7hD0V;���"O|�P�GB�x `��R�74��I�"OLL�`����aE/K4X��"O�r��rh�E��"�n�p�v"O�l�T�M!^耽a��6+ap�"OR�zp�e�f�'�̭tT@5�"O��uk�,nu���E"U����"O`�2��D����u���@iX��"O��A�O��h���d��s�"O�á�Ϲlid��ōVd�Y��"O�%*�ƥ}XVl���m�h�4"OD-a�K�	p�H{��U�IW�Q��"O���t�v� =��G��@ac"O����ڟx�%,���F�P2"OF0�dNR�Y�$ՋWj� fF��"O� Qd�!]�x�@jM�~1č#q"O�t�@)��f��Y"�$�P�"O4�L�2��AUCܢa��yA"O
y@c� (TZ�����@T��W"O�P���݁w;����Ļ94b��"O���Q �Xd�CQ�F�
/�AJ�"O`�0�d?nB�D����\� ��F"O�IreEϛ'���I�X�"O��R�,U�fe�$� 0BY�"O0�������Z%a�$ɑ21��r�"On �Ef�`c�$�P×�M.*�1U"O<u#E�\�~(9"�m8�Z�"O�$��m	xb�h�![	=v��"O���G���nĠv���~ZM�S"O^}�4��%k28�F�VV��V"O2�+�F
�)�0|R��g�����"O�a�Jϒ:���+ۏ(��ԃE"O�����D�Ĥɏ�{`�@�"O�8#�O�b;48�m��lG� ��"O���5��/�
�R�=(A��ؗ"Oh�� �Z�x �$Y�a�2Rz��"O�x$�0�� i��A�P ��P"Ob�"쏬$��W��U0�:E"Ou�a�Ki�4�����)?&H5ʇ"O6|��B�8k�Qx@�8k�>}�'"O�Ik� ,��q���ǹ!{$��P*O�gCҥc8���$Z�G-b<��'���Q����A�h-�`J	4{�m�'�DLC��BB-�*�7�x=��'b�s��-M7
��V�ʛ)��p��'	fU$�0F�9
F@��m����'֔����&W����	F��@�p�'�$���C�"�<E1�kX�}����'ب�(W�&q�е0�/�z���b�'8�!��]����$�:��8;�'�LSF�(m�N���
%5�����'�P�C��,j�^e��.a(]Q�'B���#�N(�Y��*P�\(-��'/�\��>w� �!�JC�SՐ�!	�' �Cb%X<����*�I\K�N�<I��[�j���Hۇ/��HX��p�<1�h܎I��u¦�#7�[]f�<i2���V�uA@��9f|�3"��z�<a��o���"��0>v�dk�e�p�<	� 'H��%�r'BVE;�k�o�<A������!R�əs?�h��b�s�<�  yd���<�k��>�^���"OH ��H�p�l	[JBf�8��"O<e�P�+GB�`/��� �"O���gf�Y���vn�t��`a�"O )�m�t6��P�Ix��a"O����"ьi��=�&��[6c�"O�hb���	
��$��a�M�"O,��墆(��)򍀶�j�#"O<ܸ��[-(�.8��	O�h���"OL��v�A&c�F\s��+�r�hb"O�x��2��,X5̖�}�BѢ""O���T,x��h�j*J���q�"O<���䀧j�A��hn}x�"O����I%U\ait&�D+h��s"O�|���20t]"���(+�e��"O����E�:�򈠃'�1B�Q��"O,H�aឨE�hH��R1f�H�"OK��ƈ�a��~-��z�"O�����@-ޜ��p��9��"O�)� �#Z�ּ0���e�ó"O �#tC	6$�2�ˇ��9=d�Y�"O>5)f��Ia:.�M2n܀"O�L��U*����MH����(�"O�����=�t�b�� t�`<��"O��w��z�6i�1k	_�J��s"O��A�H�*q�|� �M�M��4��"O�hZ�X"D(@�Q�_Ev�x��"O��e��4,,0q+�/eYN|9��IFX��Z�J���(7��� !�6~!�D��M��y���&
�����������(��x��3p��c�D؛d5���"O܀9�㐮G�y˵Q=5����=O���d�=?�(-��&	�uy��Wk��y�N�<�U��$K$�|��PX�#@�9�j%��+iW����G0%���/x�X���$�G	�uoZr≅	�Q���t�4�O��+nÏ&�X����]l�<�%�2�D��L��f٣���\�'axbT�'P��i�aoXU��@	��hO>���	�a~@D�ԥH�L�86:{!�$W�`.V��pd���MR�d�V_��)�'G��[��C,�(p��A�^��
�'h���1BӸ#2���m�=r�����N?a���Op�qȃ!(���Ő2K�MbDG$D�LJ�%'v�Ti2��62�5ӷcߤ��Dv����+�4���T�*����`#72��C㉙d8��Q'ǁJu�IR��S�t��	�ȓ���i�bA?jt��Adhԕ\���ȓ��pp���	-$ر
�Y���	A̓jFD�y'#B%�}�P�sE���?����~Jd�V�RMx�0?6-@pnWo�-F�<�|�@hO{S�}�Ʀ�k�V<rcll�<ѥ��P�L���ς
x@�
��@ܓ��'p���])��R�r�$�sG"�G�<=;"O��(S��x�q �"1���Y���?�S��1�D4*C9o�T�B��5��B�I�,��I#�Q�[���w�e��B�I��t�A�e��Y� ��nB�!Xq*�'�U�n��y���Nx�B�ɟp벸��@_�8��;��O-"N@C�I���u��/R\I����P�C�ɰ/�v��$�F(�ɱ��#SX�C��)�Ѫ�m	N�g,Ψ�C�	<f��t�7�P�DM�! �?wZB�I�X�R��BI�)a4!ZPCB]iDB�)� �M�"Р47�$�ƭ̎.��3"Ob��1C��a��Uh�ZW���"ORP��mi���Fm��*=L�q"Ob��D)�419�����ބz%�[��',qO� �6l���҉���,�1��"O�����د����)�4Z���"O�����"f2���;Ƞ(xr"O�ٔ��0QmF䓔�¨w |�Yq"O��D�ЏW�](���9t�C"OH3tg]��h��#GĝZ"��G6O6��D�dnLy��I�[jP����iX!�䂳-�D�т8J9�yZ5���!�"R��%ѥ��(~�*݊�cM5u�1O�7�.�S�'\0�jV�D�r����F����	O���Y~�Thn@1�T� �Ż[�D=�O�p�7J��u��0�G
�k�����Ic쓣�'L�X�Cue���I�E��D��Q��?��;�Ζ��{��~�T��yTdL'M�8R��=�wm�Z��ȓ�,x8#�����@!5��	pj�ȓB_*5���6%~���Ю���ȓG� (;��6в�9f�)a��T��U�������1�Phi�H?+q$ ���K���#P��ز����+>���+_"O�,C�Î.��0��!�!����"OB� H�&Nl�@o�~�
)Ҁ"O�"׌·8��xH�.� W� ;@X�L�'�\�FyJ~Bt��P1��e~(z��Fn�u8�$�a���*���Bq��mϛl.����5���<1�@� ,�Pr ű8>���Yr�'��aG���0D���k�N� Iy6<�N0����'�����J��T���^�D�s�'�ў�}�s�
	�0��6.��ѱ�`t�<�d̩a� %�1G�08.2���y�Ud<�<��������0��oҙ%�бY�P�E�!��`A_���pG�F��@��	,��SЋ��G?���r�[�|��U��ɺ-���D;��V�8 S��qՄ�B�D�n�qO!aӓ>�|�COֲ
T#�s� �Fx��?�lZ�wk��A��Ҁ,����NO�RC��("&yA ���a8&]RTO�b�����5JY���7�Z)��l�:�!�$[�!�(��G�K�
�%ǘIQ!�dǅ.���� N)	� aK��!�d�#U}t�&fSy"�}��7k�Op(
�H5 ���i��+�^<@��ĽN�����N�x�	��̴N�&A볅H$U������`�K㒘����=3�����eW:jO���I{N�O\x�EkԴ�6���E]�Fx�"O�E�-�d;��6Fڝi�
 ��"O�t@����ie�lA�z;�Ź��'��'���	�i��Q�µ�Q��7"�@Ղ��d9,O�������2�L���l�<5z��Q"O�i0��a5J�F�-"Oh��V�ԉ3	�icꐕ���H��'j���6�,E�Ay�knQ�a�"�.D�y ��F�%cӕ-���9��?�S�'`>D�T�-_�Va�7�^�w0�X�ȓ?lpْ�"�)Ä�6��|'���I��0=��	�����#�1���B� �p�'5�y�E@;? d��LU��$暭�yB��F<��C�k��5���K�.O��p<y����'Քx�dN�?]u18��F�Z!��Mʾ�A�#�7dX���ӊm�!�� ��.1���㧃S�.\��'E��x@���?N��i�.��0�p�Ə+D��!f�eqpA�r-�F�TpzV�	V~�2O��)��<��J��,�]����0Mkj8���]N�<a�l	1K�8Pyf��)����4d�F�'A�x�aU�6gvoK�H��qWb��y⩚;����D5>;��������yRȊ8��qBk�;���Ea��yR��]�d����!g��icm�)�y¡U4�`ɉ�S��ј+�&���3�S���>!A!��G�^�	ӄ�'&|z]��R�<Q�H*& TH�BE�S3�1T#�N�"�M#�'�qO��p���٘� �y�54v�H���7����z���':�|X���X��hO���Dŋ�XpG߇V]��Є�B�Z�ay�I�1�)�R���Q�P�˵8	�C䉫J}��3cΔGx�ؔ��)M~#=��0BI"Т��h�N�P�	�z��G�D�FbĹI-�p��`Pn��lE�'^�?7��:� �L]�&���K0d�8/!��T�H�����V���!�)i.�d@��(O?��v* Q�fՉ�&P"!]n$YB)8���*�BPl�0u��ˣ��)1v���[����=�'`ȹ7�
�t��8sft��BO�<q$�0�PUK��>F�lX��ZO�<�'�԰$� Y֎E:��y��kVL�<��㆏J0��!.y��(��H�<a�f](�0[G,�-PT4���@�<A1���\�!� �=/d���梁c����'�
ȣ�* A�6�=��pP�'*i#n�$n�xA�̆'� �'�޴�5⛜�R0ɑ�5�T y�';�5�����t� �H�>Zz�� �'�	��HO�no���@!D�a4n��'Hؑ�������0%[�F'N@y�'��@2D�[y�(s`*�7[���	�'▉qTO�H�Hڀ�]e��	�'�(�;7�������(`���'�J]IA��tmȘ��G�8ʁ�
�';LR��
>_�\��)�$/$��	�'mnh�!T@���T"����I�'���c-��H��΀��R�H	�'����ʕ�r�ģ�+5� ��'5�]��!�@�fq4@�,4�0 ;�'���j)SK�Q�`8� c�<�P)նI�.!��B�8�����\�<���O<�>M��Z�P�>m�djU�<9�$Ϙ~$&�Hb���M+ē#�>C�%t(�H�AL�>�J�Ͼuc:C�	2<�xx:g�O�b��h��e�*C�!8��5
h�".V�IwE �[�C�I�O�����Ō^�l�2��ڄC�ɁV�v� '��,����B9i�4B�?��3��վ;"R�)��0v=rB�I?��Jiћ0W"Y�w���C�ɶ;W��iV��h�$Я��B�I�'���1�NX>JBF�RI�S��B�I�ܱ��C^u hi,�	BB�IW�L����5�,�96�3��C�Ɏ}B:|B��,�P�pk�j`�C�ɰi���s�D1&0��ia��)��C�IKFY��259��a��z�C�I 0���F�1��8����p�R���˻{��Q�h�-J <��W'T.LLb1�'Ԙz�!�� ��k!*��|���ԍ�H���"O� ��A5]sr`�E�'�&�r�"O�`X`�I%Q�0���,a�Ay�"OR	��NB	o/�����3b�F��"O��S�(�NP6   qk���#�"O���EI
�* �k��%N��	�f"O���E�l�0��<8�vT��"O~X��ͮ,�����As�q�5"O���u"ƈ&���F坂��q3"OF�ICn�@�`h�*!(逼yq"Olm2�/��P�r��.�Bya�"OZ9�����B���G�H`�"Ov��O�6T&ڀ�=���d"O�3`M�w6jhr�V3�� �"O ���#e/����ʕu�` ��"O����)y���"T�*� Z"O�E���@+r(�T��dߟy�tD�&"O���&ZV�E�R�[�F�
�'���'JQW��a�f,^x���'^X�mA�J�����F���݆ʓamH%	6fA8��3��Ӆ�N���giv��pcR�1E��+�a��^\�x���U��O�,hCUOɊFr�1c"O
x�נڊe�e!#�_�|+Txp�"O����3�m Tl�{x�!��"O
� �
�o+$�m �!f(�Z"O�|S�#d��4r�'�;H>IxB"O����J�~�:4�7�ʨS9н9u"O:��ɕ�g�2}ysFNH�"�"Ol���*�r���F��".h�0D"O�!�F�Cs��qᱥ��f���"OB�Z���	�qz ��[��u�A"O��A��U�Va�U�\�k ܑ�"O
����&l�hrG�R�N�8�"O.���!j�����3>����u"O~8��.ě9w\a�6���s`"Oʁ�SÚ=�FQ��Ѝcڈɚ"O��sqV�M��Y��ǰ(˘�h2"O>���52�>!RU��!�,u�6"Or雂k
6:�~Hq@ķ�nU��"O���eZ#v?�}�� [7�X��"O
Hv�J�`�u�fN�aif@��"O�A���*C��#Ql^�A6~�"O�A@υ�	�Ƞ0׫ߐ9�&�s�"O����b~�%+Pi�X~�1W�')�����,I�'J�10�nh ޼H�ǐ/ �|1��'�r`�#M̩A�Xz�EN*8�eK�O�%���Vx��N�"|
�$�Z��W�0��c�m�<��o@jјr
�7^���Qc�:dtU�'�l��fY�ϸ'w�dstaՠDwr|�J��e���{��6s�D#�cՐ�x�����T�I�;.2B%ٱN��0?��ދY��I�'[�*���K�'-lA8� $�xIH�?��G���:p���Ѩv���Q�-D�L���ˊG�0@�7ɏ<}f�����<�P�^&9� ��'�0|ʔn C�>%1�DjNj\�pB|B�	�K-�mI¨��L��D`��y!l�����<!���v���M~�=	ƖD�D0�!�U�Գ'�e��P*v�O���ȑ\�Bv�U|�DY�Ȁ���9os�d�$��/P����`�� ���?I��u�N�b��1��Iʇ����&��e5U#���~!��Y0(������;*�ɛ�j�1ly��?s^��g�Չb��S�ϥ�ϧ3���8&`Ԯ Y�H���^�<�c�:9�f9���إkFT��'i�:�'GP��)[�g�g�d}��T���+d�!N<�B�)� ���⃷T�)k�+� �6��s"O�i��%�|�Ǡ��8ɑ�"O&�S��ܖ%�0�"��. ��!"O"Yx^
��M��o>,���y�e�����GJ�d^Ա���:CZr�(�{�(a���Ğ�s&P���C��a�j��{!��J%#6@Ka��Y�`%��_-=`�\"�C�$(����"8�iBbI�	�~�0�S�cV�x䉉$�*���-Np��"~
��r���JP�E�B��5b?�C�	 EP�Ѳe�_3��c�#��;�nDKUƗ"L��"��ob�C!ɇ�"2~Q�A�O=(�zC�	�����U|-~��g�ͰB|��A�)�~��?i�	�S���{�IښrZj<��G�'f� �"�=��?��ژw�`��Ϝ� B�a�#E���ǀ�h��Q�P`$�Oq����Q�6�����$:̸��	
xuPɺ`��8h���V?-آ`=vU8����6�rͰ!+3D��r��%s�����١���v�`y�GĔ"�UKjZs�^�D��oV:f(����!1�t9�B��yr��5y�%��͋(HX؈�+Z`E���=޾��`�.���(��y�#=��F�2a��T��E,��;�n�~؞��(��}c�	˧A�>0���6,ݹR���s��^�k�l����<i�؍;��'[������~0f ����T7h�{R�E�	���-�4�T�A�Ѕ�X��OD��,�<�����7@��qz�'�ډrW�J�6JyQ�# ��l����*r͠�y#���9�J��=�(�h���@���J򔭑��R�5쮍��s^�b�$��oL���B$�9���EQ*SAܨ�$؛/F��3!H?s\�>�cӽ8��`�)�3h!�B��xbE�͆].8��W�N�naH��ۖJ�bS��"K㐁RQ�����}���rP]�B_�4��e��V6żd�=�'��dR�5�ӪB�`�n�)n�	~��G3��"�Ȅ�9�T�0"DQ�Ն��	Ó�о�&LKB�$Ht�b��28� ��`�B�"�"h��Wm�O|�	�Wj�0Id'�aZ�-AQ�ĩb��C�ɔv�*8�%�ٶ#���(D�$�PI7_��}"���9�V�)�A�v�R*Y7! ��&��C��C�J螜�ħ/eL�B�-lO������kY*�1�@WHm>��e�
�v��ibEψ�Ge�<�$f�9]��6��1O���҈,,O�<(e)"Y�X)p��-���
��'QR�2���U?qu&�(Fa�]�PC�Dђ���Y(^��E
¬�K̭WV*A!:)�Vh��C�P����*[_��%�E��yP��`��	-@(�H�H���0Au\��2(�/D,�t�C�	
3Q��X�k�0{N<
TI��zz�|�h$"������%e�H��2MĀTLF�)��D'F�PyV��,�J$(�E�QlFlZDN�T�'RiB�'��<K��ΰJd�����'<�4���Ð*��6α˸Oj�5��H�>2]��Z�@��TԀT�Սڿ��3õiI�Uj�/��Y���*U+H�� ъWd�c�](>y��B�bĨl
�� 6}�O��P�៌����)S'\Xڃ�E
(�^�; MU�z����Y$?���Y�1�T�5	�E��d���T7���B-2B`���C�y��0�rS��a�4��%y��H�i�y@«�m�����'T�}�d�$hN���2ǌ�g� �`B*`nV���D�<9!Ƌ6>�:�&%}��)�����[��\�U�x�5Y�Q�X�)����{��ӔB�������Q0�5{U�čm��2�l�;V�M������F�����P�R���˲"��0�0�;1d;O�;��>�BA��O�D Y�,�C�Y!���ls��H�0w�`C�	��1�UB�)r&�4e9Z��Z�X�cA� ���G�w	hŲ��*��O9��%����݂��٪Q*�u�
�Q(�}��#m�|<��e� �Y�'?z�Ͱ5�'Y�ఁ[�D~ O?a�$��>l�A�u�0L���b�G�<i�(،+�$��Ƣ�P�Ը1�cU~}2!���L�R��'U@��T`�<`�`I@4&o,Ip� Ӓ��T!ݔ�8h��� ����>�:pA:D�LC���;4���������a�<	rC�=,�ć4[��D�� ����X�a�.Yo��!���<�&yK�"O���-�.)�H�j�E=B��@i&�X;�V��Ʌ-%�V�;Ċ��g��XO�c�,q
1�Pa�	�07�ة��1�O�ܹסу�8� �{���h
e�:��@�>	����7nJ��N�h�3LO�9�s�!O���ٕ�y���	.!���#�&S����p�L?��b�,��� ��aPE+���Ó"�Px�Q"O�p��$p�񚦥\�r^�xz��i߲�Tnߡ]Ժ��NK�Nk��D�3J��c?�X�{~XH �KŬbF؉�bH��B�I�Ux�Ǐ7Qp���\�f]B�2� фTx�xSŇ�ZFڵS���?��c��+?1On8����<[��� a�*`��ag�'��mK獜/�M��&4I��y+ç�DA�m�cD̓~c,X�di�0y�]`4$8\O�姝��bͺ�G\7<��<aቒ&Ϩ���ιP�����I9l{%i�l�>�uǤ�"u�i�7`��N|�)�v��y�ݿh|0��A��@j�0I��ܵ^��������aJ�p��M��s����C�o���B�Ҩ �:�f.D�P��K؆+}�B�"P�G��53Ճ̈́\��m���^)p'�4*\�V7��F�'��I��ޗ�<��i�uB�N��+"��}ꜜ
�����J*0[�h t�%x�4)��$m����I)*����]�y���5`L	F��#<!��>Q
x���ʸ*�,)�e� ��	A�@,$����2g=�ՈX�G�!��ف@; P �!ܷA��Y��g��r��(����M{��7[r�׈Y�A9$T�~λ3*��	�3whQ�S�D����	M�u�28O �5�@�wR� pC�ȏy�J�QG@^� �I'%H�3m���g�Ńr��vW�<0�{�Ǌʪ0(宀� ��kբہ�OX|��Ȏ#��G�R���L!V�r�я�D���]�oR �&��.@�p�ěs+���� %LO<�(wŜu	���e*ъ&>pBe���q�^�i�`Ky�I�?�g\�$*j�j���
�D5�"\!6���B 猞9"y�I՘b4��ȓ����MI
�X��˛Y�j�o�2] �������uYcۏq+��ۑ
�]�P?Z�_xu��#M�c�����#L��{B�L]�����æ�� ��7	�-��k�����a�
���s �?q�d��̏+��'ݐ䡣��֧z���J3JCk�1*EfKd��O�xQ �\�I�,��M����`Y:Y��UZ�%\�6/�)��c�0�>�q+��W_��@����6�)QsJSZ���1�b0�|j��G4&��Á��/��A�#����ɷ]6��slFN����F��q2�U�㚾w�T�e&�Jn�X&�86���ȓYj:S%�ɵ*3Z�АB9����	0W��p�ԍ� ���=Zm4C��/9J���T���ZH�#�/�����M�;��=a�Ocݪ�v�z�ޠ�#�[(��!8�g,R�H��ʍ�9w���7(���)��<�Qz4@��K@`��r@��k�'�)QuhW6%��>͛�;O�ҵ"B�/j�>���|���c|U��W4��y�e����ғ˜�'�b�p��F9:M�(�=E��,�� �N�s��dQg���?8���ȓ�~uy��ݾ-�$m��Oƨ&�9�ȓ���{��o�&8	�)F�M�x��ȓc@ʵ�P��C|��1�+-�@��ȓ`�x���Su�dhT�R�q��Ԇ�sc�`����Cg�YC�x�ȓ3����/J�@%�T&z(4���o0��Y �Ę(M���B(����]�Ҁ��S�n��~��mh�#�e�<"(YĒ���ԧK�$���[]�<y�,A���B�h�:#	��.W^�<�$�j�,��l˨�p�)�+Br�<�uJY��8ت�*E��!��Im�<Id�*Q�� _&-�$UЅ�n�<y7	��JD��:�� Q�"A\�<�� �%�j�Q�� <��I���\�<Y��ڦK���e�iq���Tf�D�<��AV	P�dH!����A7)C�<��!�v���s�+��"��7���y��P�`��i�Bh��a^�{�
!�y���y*��05j4�tĐQd�9�y�*L�VY�Fɛ7*��Q�T8�yrm,�5H�Ȟ�)��%"�b�$�yc�%O��p��k�|� ī�JL�<���7f^LQS�YT�r�X�/DM�<ɠ�Ru8�9��b46R0XT�D�<	����T�hѲǃO�9�%qe��@�<�s�Kg�Vђ�g��X`�8a��<�&ƛ�,L���11���@2&�z�<� XQ�
Ʋ'�3��H$L9Q"O~�vo��D��*®Y^�8�"O����X�2& p�m��M
t)�"O � �훣m�H{���o���!�"O�Q���T&V_��b�HS/ɚh 4"O�Q��Zh����'Fֻn�l�:�"O�D���-�A蔥�J���"OX�J�V|,�$
R�6�6�b�"O┛��\&y��#B
��d��ܘw"O�q���%
��3&��w��+�"O�@
���]x(�P�hP�Gb��H�"O��������h�G��A7F��G"O&ՈEzT� (]%�䋥"Ox�c�BאZX�a��J�(�I��"O��A��Y�}a8��A&ܔ_ ��(�"O̵�v���q&�(ivG�����"O��$*��z��31C��1��-�"O�	�Gn�%QC@d�"/�nQd�V"O0 ����\�l -5?�f�c�"OB��u��Ka�Q3'�7E�~xk�"OP�v�[70��rH����uX�"O���bE���X1f�S�{�`�"O =Q��C�N){歉�PҢ�5"O@�Q���<��܊fL�E-R�A3"O���C>
��`@j9_���3"O�t{sʉ	lXl9�iU�G��Hac"O0(p�K΃-7�����	H�.�r�"O�p��3qF���ǫH�@�PiA "O��S�H3*p^s�]:q^A�"Ofڰ
��X��yPB�$ɫ�"O�[�L(v��p3�Ĵ���cC"O.hq�$T<��C�C	=�,{�"Ov�p�U�L�$}Э�0C��Ka"Of���G�&�R��C�>� ۆ"O���0G�g����'��~�<q�"On��pd��@��ЮE�R�iS"Op�S�GB�}q��z�h��%�n$��"O���`P������?ZٶI0"O,`�[(y��A��r��"O�)��'Zp��qWA���5r�"O�ҡ���<�Dh@%!I���g"O��q�.X*|�J"WF <a���4"O�p�HΒZa��Z��[H��m�"O�l;�A������+V�2���"O�<�p���MΘ��1�ʱv8����"O�|����O�$����H�(�	��"O촓p�×
���K��Y5*�T�R"O`L��	��;�r�ه(�2��b�"O���֫-s�U�D�*������'����w�R��'�~H��
��D1��`C�֋O��H�
�'Լ�
u�Jq�)�kفU����O>,s��3��)@O�"|�4�0<�L2wjݒ
R]z�'�X�<a�g*s�)ѣ�!ZL�=�7�%x⥖'�l%��h�ke�ϸ'�0y�ǖ��[(ɱ<����
��-�<Y����1c��dK�����4Ӄ��^EJ5c��L��0?i�-�"S�"�Ζ""9��9O��6��y�<)q�("��Q/d�&%��k�%V�Ls1�s�<q&"cH0槗+E����el�Pyb`X�[�
�R�KV07Aa����fpx4�
�	[���b`��y"��<J(3sJ5��-�����s(OP�l�5n��qO4aW���$!"�O[�Z��}���',!�!P��@����q�H�Q�����:`	UH�a~∑� ��p#%<`
]����?��O���"M#��9 T�.U�J%5���SB®8�F�Q%�h�<� �	x�EةG,�#��1�p10#�� H��F�=gd�rp�>E���N=Ux���d\�S5K ��y�A3]�VYc�@)]�ϊ5�O�4�
����NT�
�'�>����7G��^�p4�ȓ8�����&�p4�@�U�26 �ȓ&��p�۩d�l⥫��-�`��,�*\��`ϣ<~�8
�㚎+�&E�ȓ9�2u�K�<����g��A�܅�f1�!H��̿9KXP�A�[踹q6�^Bܓt�آ|�'�N����
r��#u�S�y�z��
�'�T Ae�
\�D�����t�" �uՁQL��U�'�Z@ �#��.�0�h� `��{�LL�l@ #P"F��eH�O�d���@%gT0[RFț'-|h2"O��Z�L�f�=�H٘_
���w��`k��ѳ2�  C/��ȟ���m�H�D)��e�4@��-�4"OV�+C ]>A���K1(���zD��7�=�0Z�Y1��V!��g�y�PĀF�%!�xD�t`ì������/{�@�8Հ����@�gS�aY��ju������`�'�*�BG�N+H��V�Æ'-P����D] 9�8�:P�Y�	��P��N��TDˌOp�ḗm�-a9��ђ"O0���5Ģ�1�Κ)@�҇U���F�=g�P�J��?}3"�RnhjX���	C�h##�&D����T� �� �ѣZ)c�Z��f�);gB�
��=��
�.��k\ ��ԑ�HOL�[u�H<U��'L�3��	�'��Y�3���"@�x7��V�� J[�d	��k��B���8�IPr����I�����jV�$�F�:p�̲@v����#�fI��-/T��9�g*T�:d��G&(��6l��ebD�1�f���C�I�4(ād(��8���s�E��CK���{� C�8v� �!=ʧ�����*�b�@Q�σT���⋏t�!�$��V̌��4�D��2�𡂪 ���H��I;O�X�ѧ��� ��Q�h�F}� �4�.9CcN��@���7+���p=����,���r�m�����Q�^K����	��:Y����OC{�-ɕ�'�y�!!��QT�F�:�k7	����'ީ���ڿ�6ɀ��Q*���.��'8ȳ�bE(90bp�R(t�����+�=Yv��O/&]����jl܁�Z�aq`Y꤂R�z��ؑ��y�On���	V���3�n�L���8t���mSJC�	�eITi�s��.?U��h#�7H�^�{��7>� ��S%�4�H�T�8eKO�=W��$���#�%o��w�L�K��1���>lO�I#	�?$;Zك�,L�ȼ*`�o����k56��1��	M)�h6m_�53r��1,OJ�hq�X�y�JR e�P�`@1f�'����a?�&C
1'`�1^�H�Hd ���Ő2�*"�*��;%�F����ɲNB&��I����d3��5!�@7$�B%!L��	�O4����(EF i"�
s��ʰD�!Z����U�(J{�8�q�@�Ee�T��'�Y#�'`P)�m�<p��T�ԽxD�����X҄�g�A3H9T����?=�p��|���4}��9^!�ql�c�rH��ѿ�(O�;��<V1���T���Yk��e��y
�`I�^<n�����^�^��)���۷-Cw8��Bo��-x�Afϕ�>���5E ��Xƙg�Xӧ����e�X]�	�[�D�q�/
�HrX� ��|<��'W|�"��
O�A�ƕ>�I�a�*���B�O���H��Z�0�'�¼��C����O�	
�GY���
�C�o�k��|"�E�hض�ӲE�ڔ��ci@�?���E�����?�������]��ӧ���h��U�4$���-��/ty���	�[��98 �Ԛ6&>I�Em
yu"� A�	 ��a�/?�c��.� �6O�H1Gk��s
�b�d�7�O�qg�L!�I/p�di��>����\<U��B�)S�|>BAU�ܠ_�,e�v ֐�0C�	�S�@�z�(��$��D��FƳk!��Ec�1	���$���?��9:��)��O<�
"L:v4H<ӂ�A�(
V1�Op�80����M���"zd�!��e>���HEџ$�g�N; .!�I<E��+28{��?M\� �)CH!��&\R�����&	��!�)�� R��\�$a��La��P O2~�Q'�
O~��R�(�O>U��L�@h !�xC�N'>,VEzT�B�(ÔH��ϔ(ɀ���,-�52�8[w�\GyR�M4ŀ ��T�O02�q @����Cʸt��l���� �ɪa�ƦxD�08g$�@�a�,Az\�D�qt�S��?9gI_�vq��D��l!Ca��k�<y7 � "��	
�#�����.{?A�ּN_�4��M=LOr	ĥ��,���=��j��'��\C�+��Dy9dHB�J��P��cJ.,J 5��A[�<1��1_j�([્+	���� �Y�'��qQ�3[l� G���v-"��tH#tn�Q���(�y��9-�v��Ϫ��d(0-�Z��2�א(��I�"~�	�l�f�p.�)Kn(�h�n�B䉙���T吣a�( �&�>p��*��g�� �p=�FAH.j��Q@�<���.�{x���6nE;k�VM��y��O�!HxH�Sn��y�$�'5���b�ʄ&"\���C�y�Bƍ$(ȉ9�b�&(��#B��y���2aY�K5m�W�ސ҃(��y2�=|�FU�E�����r�	&�yb�@%{�:�*�,W�@ac3��1�!�d�*m�Ä-K�m���#$���q!�DV�cL0�"�nF=��)����
7�!�DĀS&|��a�\�2�X��"��.�Q����D�R$x�E�4�֥D����-T���9)a�\��p>A��1s��	-t��x�芮�H����=Z	��R��Y
u���:!�>E��'C���s&�:�1c	-� lJ��$��Ol����,�'I]>h�0l
�fJxyw�CBE�Ɇƪ�S�dW�r"T܄鉃 �`���N�0YD0ۣl�!@�@1 ��>K��K��&?�@�GX�F�b�2p��,0��8�c@�G�D��$�=`@�,�ȓ)H��D Ů^y�b��r=�ɈBBĊ���.�X��P�а/D�xT��lyJ?P��|!��T�^|�pb��6|O�A���F#1b	@�4�D�ه�AOF�{�H1ej
�j`Uz�ԡ�Txy��D@BCڛG:�|XF"X-��A!�2�I�*�q�@�G55��>������g��M��J����9@l�O�@��ۧ|����1(9LO�%����3�.���3c˫��~N�͓6��&	����U��9��&�P�w�]� $��gQ1���C�y"��Z.�2'��GD���tÉ�?��%R+v��A��	L5�p�Pf�X(�j/O�$T�l�!�I�[(b-��[�::u���y��a�%U���I91�����B�\�^B���$ܙPM��Qc+}��9O$ ��a���S�O ,7N��	VD
<` ��Y�OlI�)J�WZ�U° �Y� ��'P.��r풆�a{�j����c��ڑR@�$PI�(��ı��_�Ƹ������-�|0c��
8�� �̇��y�ϛC�AAJ�0kX@��C [%�y2!P�# HB5��ai:I�!	��yF�T#��;�l��k�f��PF��y2M6��QF��[lv��� �;�y�N�3��H���CWQ�<Ң獚�y�N$>(MA�ԐO��x�a�á�yr埿c��Qg��&=	ԁ��iŻ�y��M5���c��D�[ъE�y��� #�jqX�&��i�zz��M�y��HW��;���1� ��Ɓ�y2@ΫQ!��h�G��I�C���y�BE:jX����*��lp��:�y�/ur�K䔿"T�ǦO �yrmN�ْQ�`F��A��C��y � 
��{��-n�X7)��!��S�I�h�P t�*��1욢'Y!��Y��� ��i��<xR�T�$�!�$*Fq��2a���UwD��#,�!򤒙Y��O�q{l)t�Ҽ	�!�d�I���Fd�R"���6�!��> �Pe���)[��bg�
9h!�еh��tH�)~D4� #E�	�!��9�@���L�D���TCK�c0!򤆲FGܴ󳋘@zlC�T�|!�� ���(9�.xJ����E���3�"O|E�:_�L+��rZ���"OШAå��L�P�gޅ��9b"Op�GO�W�f1{g(X���,�%"O�D ��x��<�5h�,O�$�Q"O�����.[�ݱug�A7RXs"Op���L��W� d2ed <-�� g�'�p��uKV6a�|��	V#����GF�j�k�'�L���Ѐ/�t�I!�Q03(\��'�H�!U�#p]DMѰm3)�h��'���g�,ԁѦ��+T�k�'���'J=�ƨZo� <[����'�����%$�A�+�!�Iz
�'��XQ����z�b��F�L�x
�'�����}��K�a��%-Rx�<9�Ƒ@"ι�v��C��ᯟ\�<9.�#z�نGĨzE, r�Z�<�Fn�6SV-E̅(i���S@ɖ]�<I�M��@Q��H檃�/D@q30�s�<ٱb�%��KX=s��)��Gg�<�"ER�9�2�C˶,r�a��,Xe�<����c��U���P��6U�OHi�j��!�'K����*G�{��y��37w`E�O��� �O���0�q����&�? �������2Ю�Qn���Z�:�(l]ر�_w����'�$})E�N�1��A�֪U+N%b�Ru� s�\4k���X�R��~�*�
Y���uMذ���q�\�.����k(]ֆ	��O���)R�7�p��t���$a��@.'� ap)�Mf��5p=y��IS�)���`����ɁD��Y�%���0, *�O�@t�ەq]����;�b�}�*M�`�� ��/2+X1��ũ�?��.�!��*���c_\������m#T�W��Ј2��h~��-��BdxQ��OA(������1�>��7��%HU���,���J �P&��q�T$�'�N@���	�|��NL�bAp� 9B�6�𮖙��'4����~��/��G*��;5$ܵA��KKU�<A��)ƀks�;QX�� ]�<I�޾#���z%,�::EB�d�t�<�@��oc��f	!JR��I\�<����%j؍b&^6@pXG�HY�<����nF��d��&~}�e"V�<�q�Z%�z���@Y�,B��h��}�<YC
��!8dY���q{�H��x�<	�BӺ0��(X��-�D9���p�<1FΌ=*�Hd�1�O6C���'Fj�<12 RM�h�E�8xGp�Cu�P�<!�'��R.�KD �1Ek�a�DN�<9��N�Q�l�DD��#e��fa�N�<�U	A�����*��)�c]o�<�t(PE?f(s���>�����li�<Q�,%h���&@��޲A˗�`�<A1�D(I8���%װ�YC%ZX�<	ģ\� �9scX<��1��Y�<���Z5�<}۲�	�<s��:�/EV�<�0 B��֩kӉĬ�4H�2�Al�<��ML^Q�C�īB�
ܩB`�`�<IV�ǈMg�<��L>7*����LZ�<y�)�7"�A���B�H	C�`�<!��ǅJp�AeI�z)��h�s�<	fІQ(��w�K.�nUH"n�k�<�$�H�����v�t@$��U�h!�ȓj��Ƀ"�·M�� �㉖7�~�ȓ79ЂGCŶ.���"A	_�h���'��y¤ 9 ��à�H�<Zd�ȓD|8�ԊO�hs�`�uE@p}��w�T�Y�gҜ_�dCpk�L�u�ȓ*�!�O� +*����R4R����S�? ~ec��<"�T�s�酒;�vy`1"O��ui� N�A��yږ`Cf"OV`�a�ӏ@3��[ȃ8����d"O��c���'!"�\(���>��\�#"OI��b��
Z��I/Ƌ�����"OFu�!�@}InhxF��=#V��"O��G�9c��!�tl	�88���"O���T��0Z��8�>�bU"Or���"
T�(�Z�J��oy>��"O�P�b���Ze���^���a"O��	�!K�IqبP�ˊaX��sC"O䌣��. |�M�WZ��
�"O r�Ҍ@N��a^�/��q1"O.�Y��1��F~��`�"OXIc�,�X�n�q�m�(&�@�T"O6�����X��|��&��0|b��"O���!�����!'G��h�8��"O�0�S�ƭR ��[�x8�"O u6R=#4@HuǓ,#��i��"O:܈��
�GfR�jRĉF�t��S"O��LG��(�"�R�e�Xl"O�|��N�^�R|�U$.���$"O�A��W�ͤ�8�H��9`"O � �I�F�~	IP!ߕ���*�"Od����F���1��]˒���"O>	je�3d�}I"h�k����"ORX��� @٤�B'�,�Xe�F"O�� Q�ؑ3��s��
�"��P��"O&�xsɥp6��(�dI!od�hI"O�l�P�l(���Wf=�w"O��J6��:6�,`³�&n�#"Ov���ĎKj�c��9jd s"Ox0VB��R2lC���7�`P�"O�@[B"�&�����ʁd���"�"O`rV�׃, ��'��pӢQ�"O��6��!ڞdH1/�X�jd"OҰ�Vo�+|��	�N�N�N]�S"O.8I�͘�@��*��zi�� �"O��؄�"L����6N�I�İ��"Ox��\`�e���CaqգE"O�\a��4`(ܪ7N��uZ�j`"O�|��RЭ��K�u#֤�"On]����	&��U�O����"O�} v�Oj�9����
�P��"O�@K�/�6d���Y�E_ .�<�"Op�p�뚕OA"�b��5�l��"O�h��%F�Om  ���M5�u"O��b����A[���F|�R"Oށz3-G�v ����
]$D����"O��9񎘺|���2�h�7�Xu"Of�����&J�X�˄�J�d���"O6\"��:T�����K�h�,�h�"O��ȇCB�|� �{�$�2f�<=0"O4%i`	�1�:|"7����<P�D"O�����D��A����<��K"O`@� d��ɱ0 �9�\��"O�4 ���4s��y�Q��:ɬ�Q�"ON�J���9���GD�q�4��U"O�𙤇��`��5mD|�@���"O =����wu�c ,̤t9)�"O�S#gB�	���LC<p���d"O"h.eD�1e';P�F�B�mǳ�y2
�-=�Ƅ���"P� ��6��y����'�p8��[${�Jw����y
� *��2,B�M� �d�W4�X	�"Op�A�"��p�)xS/�bf�
�"O�E�e(B3
�(�����RXH1"O�30(�sC�x�v�F�|Pz��$"Oι�RO�@�U[5�3%<R(	�"Oj5��Gf~e���פ%r$"O��a�M�8�V�$	�	�T"O��S���	����^y"O�=��F��:P��g�E�Dct"O��f�׭+��|���5A����!"Od�r�Y�tŨ��S(Pջ�"O��V�h:�ö"	>l 8IY$"O��u 	=:T�x��^7�x��"OڰX��<4�2��G�X;;�#"O訣��,�Q�$.�QsT�A�"O�$*j�8������*n��ڧ"O(غ��T����H>n�:��"O0l��(�*]]�yQ�╺d���b�"O4�S`&�=z�(y���*�<cV"OfHS6n�H0���`�<T|�[�"O:�h�=g>�����J
!��[a"Oxj�A�ub,�^�a��)"ON�sY�b<��-�c��ձV
4�y�i�$G��T
1�M`\Х��A�y2Œ	��Djv�$X����5�V�y�U�\�|pv�_7!��QV��y2��H�0i& E�B���5�-�y�f]�#Ų܀t�<�`x�j��y�@424�d�7
Z�3Z�}�$D���y�ٕ+�\�@k �%eF(:�m�0�y�A����\2�ʄ>H"�[b"���y�M��V�"�0��Q�Fk<8"Ql�Py�&��sr&�V��U7�0��X_�<)g�V8�@�3g�F.�R�Y�<�e.�<B�������1Z��p��Ya�<)1c�60��\��+n�� h^g�<!�����R ���0,U���_�<y ��{�쐉�HQN�Z�Y�� Z�<�	��Ո�R��a؊&�S�<�C�N�0ș�M��k��x�f`�O�<iB�z����
Px�d�0��Q�<�qBɞn?�} �k	x���j�SR�<��սg�F�x�A�p��K@�QO�<�#��Ccؘ��EE�l� ��e��H�<���1����W%[?,�Z"Õ@�<i�W>l���3�b�9�����Ac�<9ċP��^h�[B�5p�D\�f��B䉕0�ly���Йw!�Q��+�?m@�B�	�{ݲ�S��>)��!�r��s��B�	70�*L�uJJ(&��`)��w��B�I�@��t�����L���� iK-�JB䉐!���Eq�Pmh��ƹH�`B�<5+�1�2��?4�,��iF
hd$B�ɠ94��a�K��3+D�8çE�i�B�I(ow�ԋ4B��+�ظѤ�/�C�	B���-
bG�-yeb�B�ɄF����2��Z{�}8 )Ыa�bB�6P�T�G��:p*����C��C�	�-(ȳ%`O�T���g�M}8�C�I�a��@ �Ä�]Ŝ��Ԭ�'4*B�I<T�<�#���X^�͐�`A�5k�B�I�:��!zbeT}�T�Q �C��2e<B�BT���V	X�H��d�~C�I6Rd��
��Riؠ1&Z�H1�C�)� �����<�81���ܬzWh�c�"O2)A��K�\�BE�![��X�"O��
�Zz��&�(CMб��"O��Q`�,z��(cт�,n/\X�"O�)�p���J,�����"OX��NCh΄�dB�k� �"O4� �H�.�n�Ňʭ}��P�"Of�4�? ���&H�<R�T(p"O��C.\/&��FEˠ=<%S&"Oy��J՛;`E�bmN�($r�i"O���4�\d-`NBV���s�"O>ᕅD K�(�:�	�e��%{�"O��
ǩ	S��
���9V��ɠ"O�Tpe-�>N��ѻ�EVr $�"O��A��3̶X`���02P��&"ODq���>2u�r'-KrH�V"O� �aE%V��2K 6�P�;�"O���J6 $�|�PC��M�6�p�"O�e��V��*(G�L�Z[�"O��B_�����ǻ�6�"O�؀��l���r6�]<,l�R�"O��1W�< �b٨���a��"O���X�F�\u�E�0[KB��"OV�I%E 5kX�����ǭ=z P"OX��W��oO1�J׀@1�m8$"O�pA�F�b��)�=6���"Ort�%��Z'b��GnqZ�"O�P3��z�9���ȅ]�Yۢ"O�!Ԥ�����S�/f��"O�hkp���NN����$"O��"O��f�F�Z�!԰Mڀ!�"O�F熩߆���n��D"O�A�2Y��|
%m@ն {�"OR�3N>��Qb��K(a�xܫ�"OH�e%#&�xk�j�-C��lB`"O�q[3o
�~.��rήF�5iQ"O�X�   � O�  T�  �  Y�  ��  ��  D�  ��  ��  >�  ��  9�  � (	 � ( � $# g) �/ }6 |= �C �L V �\ �d %n u a{ �� � A�  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6j�V����2�81�8	q�G��Q�O/�yRL	0���(%�B��a�B���yb�'nP(7'�7@��*T!�/�����'�$ģ�ȑ+�&4�3iйڐ$��'��HSB��&-"m��+�1~�=��'縜P��5f�0r��
�g���J�'��P���Y�X�kG�`�6%X�'l�e�&/oøBu��@(�x�'	|x
��P�2�9���-o�h��'g�$�e�|[z�Bd�)j�ҥ��'б���͆;R��І6`�6�1�'IBk�ݚDA¸�`-�C6`�ʓ!
���s(���@F ����J�RT�HĆR�B(��h^0*rB��ȓ`&6�h
�;5�Q��Q�1�ȓY;��2j_���d@.6$����a%,����7&���*��S�p�ȓ�dp�Ã���h�E����@ ����c��!z�y���=�\��lb�����'�:X��W;x�F؆ȓe"�� ��}�K�d�1T�����IAę���݀}��3\ib���"O����AB�X��S$�P�E��B3"O���C1eB��7���A���!"O �`�-���ӣA�w�h5�"O�R�ļbi �b��=����"O��S�H�]ں�a��ޞ�Hx�"O�eq�bֶE^�%�5N�$bv(�ȁ"Oʐ��HU/��؁B$�#��m�<a��ߔ$�q` L�	\$���d�<� ��"U��%�kR4+_�Q13"O���g��H�"���	qx����"O��#Ukܔ.T����=Uu ]�r"OT������yK� җ!�"\h��"Or]ѣЗq��Jwa��pZB��"O�c���#}5r� ���ES\9�"OT���,�*v��x�A�m��`x�"O�TSp-μ'*qB植�w��Pi�"O���&�H�p���f �U?��P"O��Ň
d��J���8B6ta"O"u����
C��ҷE.G�����"O��լ�"M�����$�}����"Ox���X�l�$�����/Ѵp"O`4KR��^�d8s�&�r���"O�<��O�E�08y�B���"O�J�`C�;���_.J�H��"ON�3��&��HT��0�z1�"OD8f��J\�eȜ
p��Qx"O����Iƾc����� %�:��"OFPAw�+kvȰ�ߍ.e�䊰"O4Q����M��S&a�*2ƍS�"O��HJT�c�x{���$挊�"O6)%F��
z E�cϔ-gxK�"O��Y�nˎqC��Co+Bʰ\H�"O��J��jENUz�IE�:�`""OT�PC �t���"S���P���"OȊ���9���b�ɛp�D�0"O�����oh1#�)�&�>���"O�܊aoO?���3E�V�����"O�pR�"�[���mD�-4(��"O ���ꞏ]�\r'M 7�@�T"O8����+L�ȱ�ʐ�$�$��1"O��ۗ$��,J�ç7+�X�"O��"A��Lk0P��f_�Y��ɸ�"O���*�*���'L��$��=�"O�ua�i�8X�*����^=-M���"O� �e�P�a_
҇�KX��u"OX �e��:����X�a�R��"O����ظ
��q�B� z���CF"O½{�m�V5���A�@�T��"O�t�cI'9v��*H�gK�PC�"O���@�sa5i
�#�¤8�G�'!!���}j�0AO:[o�t�Q�]f!���A�⨘���TV,�P�I�|!�#c�,����_ � �&Q�O�!��&~�TC��Z���D� �!�dPG������
��3�&��5�!��U�^(v��x��)p��~�!�L�X{�iJ���<D��!QE�1I�!���mƬ�{��ց%d)�z	!�	�U�4L����M���U�S��!�dЗM̅8��	��j��	�3 !�D4@@Z'E�䚵`O��!���<j?��������DK��kV!�pW�Lʀ�֝{�:P2QiI�n!�3DB����_Td����
�C�!���M͉�I��p��É2�!���Ȭ�e�`K�(��c�
6�!��(= @�`��?|�6���@*4c!�$�6�,0�'� B��C#��qV!�	rl����3>܆�P��fU!�dE�C%<\�k��
'R�q%k�F=!�ĝ�2���Z�kƢG%�iؔ�?M:!�dM�j�"�Z�H�,��(gl�I!�� �=�7`�[����N�T$d���"O }��(�4��p:�)��c	�tj�"O�af-ðTm�|`�(:.آ� "O�t�4��-x�b(r��[�ʁ#�"O�����$0�0Řu�A�@%�e�'.��'���'q��'���'���' �m��m8VddP:�l.-�N ���'b��'���'�r�'r��'�b�'l�M'-efb9���&Cd�%Y��'���'��'>��'P��'nZ�MG/
*\����JʤN\�<���ϕ�?����?1���?���?!���?����?��+�
��ӧ� &ZL1 dN	�?����?����?���?!��?Q��?��NM��Ų�ȣ � (� 
�?����?����?y��?���?���?�1������S.[�|����?���?���?����?��?I���?q��H.ZA�EI�N�H>��b���?Y��?Q��?Q��?����?����?)��N�m�"�'��?C%�a;1J���?!��?���?����?9��?i���?Q�d]�I���6�,�Up0�(�?a��?���?I���?y��?!��?��	V}�ųŇ�UZ4�3��H��?����?����?��?���?a���?��j�d:tH�N� - �'��?���?9���?���?���?Q��?��&���ҢC7c!��S��?)���?����?���?!��hb��'rH	69|�A��R#8�4m{p�R.' �ʓ�?�,O1��� �MӰ�S�x��a6J�&]OƸRì�?u�2��'��6m-�i>��|�JշF��s��ŵ�\:С��(�I�"��jӎ�����韞�O��Qcq��-]$�	�.�{�~��y��'��Q�O�$���U�]�p�i�eK�T �c�u��M����=�;�MϻYb���$�@�!(���-
%d!�Ț���?��'��)�S�0l�%m��<Q1ϔ���Bt"� ݤ�1M��<��'& �d�!�hO�i�O��ì\�����E��g�,LA�8O�˓��Vq��B����'�`���^W�*2#T�wK�(kc���X}��'b2O�SP^`$���+V�`ɲ� /���?Q��^�%�|R���O�%a�A$X&I�#*�]� *=+��D,O�ʓ�?E��'�X���Кr��0��mv���'�t7��V���&�MC��O��{��B?^��$kƃ']�čQ�'��'u�lT�撟�ͧpb�d�n�p��"�٤V���
B���u$�������'���')��'2�c�*U�~�` �'J���R�p�4�p� ��?!�����<������i�MˁS�
5��h�3`(�I�M;�i2O1��uY��H��ѥ�.�Z���"iy@&g��Q��KW|��ui�GT)dt�n�q�	���$ ��3-��h1Ȗ�O^�`�$�O���O��4�<�v0���Z$2��cݸ%��eU _2��y��R�F��{Ӷ�D�O��o�
�M���oK`*���5�,8�k�oa�١G�.�M{�'�`�-;˚�4�~��$>���;H
��롤���Љ�ւ@�'�����?���?!���?����O��,*%RH���Aß9bvU��'�B�'u�7M_�|\˓;ƛ֗|��� hd��5J�~X�a�)��'�������3sp�V��<� H�^���14`M�|$�ӵ�@7!�&q��Ox�O�ʓ�?����?��z2��4��+"`�Ԯ�#e���?�����d�𦩁VC쟔�	�<�O����M���S�i�ijFDP�O�)�'
��'
ɧ�I[=H���!�E��!�$�MEzL�Ճ�^
#�6LGy�O�@���Q�����
$:����1	\�H���?	���?��S�'��d����+�x��m�#Gw������]����,aܴ��'t��?��L�#�����R�.�F��(ߵ�?)�/�䬪޴���Ȧ�,��O+�ɪA^�����d�b\�i����`yb�'"��'���'�U>!A �� �`�QkX�.�E�f�D �MS�P��?y���?YJ~�7қ�wLzA��%
*6���/ƿ,��(����Oz7MDf�)��d1�6Mn�d*�&JP4�0mP��Y�d��a�o@CiB�J_�ICy�O�rd�,��Y�\%-@]-S#����?a��?y+O%o�~��-�'2g��h���yƩ��--ƥ��e��fu�OȄ�'@�6��ۦ�O<�r�2j݀�Q�)s��
P��{~R�ń y����1טO=
e�	3WPa���y���"H���c�V5��'���'B�sޡ�b�9[�0=�pFX,,�`�a�ȟ�Rܴ+
�p+O.xm�k�Ӽ[V��;!D|h���ۼqB\@��M�<d�iX�7mЦ)��bЦ��'�Ԃ����?�p'Ŕe]0���X�jK��B
�S�'O�i>�������I������Po���-P�<8�s@Ւ-n�'�6��:�����Oh��=�9O� E�V8D(EC0�
�V��eK'b�K}�z�h�lڷ��Ş�xqE���蓠�6>5z��2jKaP ��'yj���ןhz��|�T����[�g�ꤹ᧙�]��Hs@��T��ϟ��I��Sqy��pӂݘ3A�O�����	f�^`�5�ʯfZ>��6O֙lZJ�j$��=�M��i]b7-@�$��Y �S":�PCBDC.Bqf���l����ɇ\�`���Oq��� *�x@��@FL���-IQ=,��g5O�$�O��$�Od�D�O�?%��l��=0d����>"x�8�.��$�I؟X
�45gha�OR�7�2���y�hR��M �*A�a�80$����¦�'H�x�nZP~�����AS����8H׍�?:/cA��؟h!!�|b]��S��$����40�B�e��Xa��)A�舳�-�ʟ��I\y�JqӦ����O���O�˧$|�}Ӆ&B�TD��2�c_�iH4�'������o�d�%��'���b���$��@՟�U�1Ȟ�M$$0&Am~�O�`��1Z��'ڲ�q�m5c"��bMP�5��K��'�"�'�R�O��ɤ�M��;I�9*�MI58z͋B�J�W�z��,O��l�T�38�ɋ�M��lA4jp1�s��rLa�A)�#ΛFm�H���n�2�h0 3��d�Oƪ��1BX�jG��bq΁�zF4�S�''���l������ş���E��Ϛ���M�1u��f艘Ȁ6��;3��D�O�$1�	�Or5mz�%`�hL|n:Q� ���`��)��BD*�M˥�i\$O1�J���mk���	>1�䤲���z�`�a�T1J�\�	+{� ��'�'�J'�������'���2c�$J�@����T	JC.���'��'�V�p�޴.�����?���+��L��I2N���a�JCa�`��k�>���?qI>��F�>�Q�k�a
V����D~�F�#A� �iQ���4��'����o]\0�ʂ/1
��Ӣ����'���'�)�'�?�#K�nKZ���FP?Y,��zRō�?�t�iQ���w�'Ld�(���8mƅ�Ȇ<W��@���4hpZ�I����ϟ|�Nܦ��'>P$9r,]��I�*������ͺ�Y��W������O����O���O���Y�V̋�����H��Vm,ʓw��R!(��''2���'�M��:y����JJ�$S���C�>����?�J>�|��e&K� ULŶT`ВC�Q�XZ��4!���"�2��r�OB�OJ˓�|��N�(��P���S�jx����?����?q��|z,O<n��Oo>��	�3�$���E����̘.&�FH����M��R(�>��iz�6MC٦1◌R�j�fa����;�� ���$&#41n�|~bD7���t�'ǿS`FT�/�"q���ʁq��D�wl�<���?Q���?������O�s��,�d=٦n�')�lA���<��x���d�$���QӦ�'�,)VC	���S�bMY���˳Aڐ���?���|ҏ��MS�O����J@���A�L�&�k�O�%G^�DQ��̒O���|���?1��vl`Z4c�z��Hӳ�I[M��*���?�.O��mZ�l2��������o��nۓ2/
�cc��w/pe`�`����Ap}�*bӖdoډ��S�d���e�կG>z�,ȉ$S��#pe��kjz���O�I��?�W�:�dյ<��	dԌ�� �{�`���Ov�D�O���<��i'�Y�%��UJ�ٺ��>'=��)_!剗�MӉ�>�S�i��c��]�8*��c��tD��a�~�d�oڿ?N�mj~r띖!,���r�)C+�H]B�K+a��t�"$܄����O����OX�D�O����O@�D�|B���K�d���*I��1aS.Z� #��I		(�r�'`��O���P���i�Q8��!�$�5�Ǎ&Z��&��?9ٴ ��I�<�S�?���+uP��m��<a�٦��p)��z��p�(I�<��Ǐ:�F������䓻?����t�'�mRe�1^�A�a�K(}��2�'��B�'�Dy)�'ZBlw���LF�?Q��՟p�vBWI�A�f�&�
��s�t�ɻ�Ms���y��'��6�i� �v�O |qh�;*|��f"�z���c:OD��,4&܌ a �:2����?�9�� ׺;�'vmqҫ�N��H �~4�)���'�R�'���'W�O��M@�
˳6�HM��
1x��D`�P�q�Rs��E���O���O�O��4�u�O�#[��B��+�"i���Od5n�)�M#ײi#��rñi����O���'	|k,E�e}�,�4����բ��״i`PN>�,O�i�O��D�O���O�Lz��R=ou���I��2m�7��<��iʲ|���'k��'y�Oi�ˎ�/Y�=����""�Ф&����dl�&lr�Ĭ%�b>YR27ay�pI����Hf~��Pb��&$?I!JW!"��$O�������5I�a�+�� J(8�#��>p����?���?�'��ď̦9٧��� �S�0*����c�G�b�`��ɝ�ĳ�4��'Ψ�hǛ�-x��m�u�FK�
=Bk�g�n j����e�'�Q���C�?��}���r����Ŕo��� +�k�Z���?���?���?1���O�Rt	�)^p�C��;z�j��'"�'��7M[-sq�S�M;M>���� ���jEDC�r�H�7cڡ/\�'%�7�F̦��~��ll~Z�p4LE$��H �ڲa��a�A�J�O�@�Č����4�����OJ�Շ+X��XcfI&"�t50D,�Lu���O��$V���֞,@��'��P>Uƫ۱=gDXٖj�:g��k�H.?I�]���I��'��yr��+2�=K�q�Gǎ�=��H�'��<��T(ߴN��i>�9��O��O��$��?.��\6�Y�	h@���O���OZ���O1�˓"X�&.ZNr��0��#3�Hq jZ���tW� ڴ��'?���?���}, !��X'k��������?��2Fށ��4��(C ��O��)� �)�ŀ�&�r50u�~p:���?O<˓�?9���?!��?������ a��H�e�I4FR�rf&ވ+��nZ	I�1�'����YȦ�'=l� ��#Y�(�z�i�����4��F6����p��7s����.ܺQ�΀�v�K���֊t�����km��l�INy�OQR愨` �ZU �Y���@^:5I��')B�',�	��M��H���?i���?! %�>uق�j1��'b�:#Ŕ���'X��5ۛ�*|��%�`ӔɃ
2��\���p
D��' ?��O�!`b�DP̧���DF��?Q��6Pw�ĬR�R�:�	δ)�b�'MR�'��S����fmԍ��(�B��M��!�����)�4_|�9)Oio�_�Ӽ�E`1?�\��@fU�g�p@K��<�a�iQ�6���q�%LŦ�' 1�i��?�"&EI!>��rEX��@�[Fƍ�^S�'��i>%������͟`�ɇ7"��Y'FV0�a���76.<�'D6M �eԺ���O��*���O���}�*%�Y�8�R�a'#Q}r tӜ�lZ��S�'	�]�4隈N�&��/F�x}�HSцO����'����f��ޟ\Ù|2S��cƭԓa �XRjۿ]t9"%@�X��؟������Ay�/`�̴� �O6�:���<"A�1;���t�X�B?O,�o�u��T��	П��IƟ8H�J��Ux�80 �*0j��t���b�o�p~"/Ӆ[���'�䧅��N	%=���0�W�#��t�$��<Y���?���?	���?!�����1�چ���*;t��9Y4��'D2Gg�|C6;�r����%�`��.\(<�*�j4�ɥz��kv��f����d�i>M�c]Ʀ5�'��
���q�x���0D�媃�G��������d�O��$�O����*ܤ�j ��� �ӂ�3�2���O��w ��b�n��	ß��O��DءF�>K��@��ho�ш�O���'��7m�ئɓI<�OS�-��W�Gj�aـk	]���sd��I
&q����4�"\��,Zr�O|ЂG$�'Z+\ h���k>��p�G�Ob�D�O��D�O1��ʓ;��VeJ�lm+�&�?P&&�!����I��MS��b�<�ڴ�J�)��#Tޮ2u�I�u�^�81�i��7͘�Y�6+?AƎ��Xں�I+�i <�`����<1�}*���y�^������P�������ɟT�O�6�P�AL��<#�L7u|A;��d���
�)�O���OH���D	��݃[�ԌY��v�(�`�;�`=���?aI>%?�R"ZѦ�ϓ`k�� b��5e� �����$w��!�Y�N�O�M�K>.O����O����~�T-�A$ڵ_�`����O��D�O��Ĥ<��'����?���e�I�n,_���@bD�] �(�RH�>�i�L��(�m���k�|!ty��Ɖ�;��I(f�B4�3 	9Q}t�%?��'wt���6)�p):*)p��Å )�\��I�x�I�����r�O���?fZ���VJU0`�p�`�Π��!mӂu��<��i�O�.N�lM��bѫa
�bb�� #���O��I���C�ئ]�'jٱw���?Y�V�͜2'txjR�	
��������'�I����	�H�I�����:(��4R�gj�3��vժ h���<���ivzܢf�'��'��O�����-���7�%��i��<}ל����ӂ�'�b>���c���lp`�ʻ\jL<R�e�'HO։���.?Q��ݶB���$ӝ����DS)!7Ɯx�䁹"&��*# ���O���O��4��ʓL������h�rO�;6'Z9׫�$��۶�Ʉ]�B�u�b㟬h�OH�m��M뇹iKBѻrS��9���P�v��3J����X &��R����)���:������x6�U�	箩#=O2���Oh���O��d�O��?)���٩�U9E�c2�"w�X⟄�I֟���4P�Zϧ�?QS�if�'\
��BH�9F�xj���0�,�B� �D��A���|����Mc�O� v�O@&���J\.�F����W�"�i��e�ƓO���|���?Y����г#̑=�.H��	�L`�-����?y)O�qm��N��'�2Y>;2�ˮp�H-��@_#|Hf��;?��W� �	Ѧ�O>���?ղ1�ҀuO^���OO�]�n�ˣoW9'.��C�9�v��Ef�O�� N>Q�`�4U�d���Y���-�?���?Y��?�|�(O��l�)[(���RM�(d��T�<9A @�Ɍ�M� �>q��iZ�U��E\VGDBf�c���Ч�zӬ�o��s!�Ao�a~2\#V^L0��T�)��,`��!%=��d�K�'��d�<!��?���?���?�-����WI޺,�4�0운n�$Ԡ�'P�����BџL�IƟ4'?I�I��Mϻ"��0ː"Y({X�T���db�!(���y��x���`��9y��4O�����J�T��*��m#b�9O��8@H��?�6�8���<9��?�AC�99ĴBB%�9M�����?���?Y��������W�˟���۟D��D�1�$��WkN�HQhf��
+��ß��s�ɉyF��Y4��f}��`���R���l�zۃ�:�M����&�L?1�J5��ҕV>:�(X����#6=����?����?I���h� �d^�>U�7Hޤn�Ա  �[	&H��DZʦ�����x�	�M���wc^ac��B�3c�T�j�:�'�"�'$BH�_Л֚�� � <��� �L@�.j��.�7��m�eK ���<��?����?Q��?9f�_�:�6u��
K�G`Fh*B����$���I�`ȟp�Iޟ�'?y�	��P�Kצ� I��q�5R#, Z�O���O�O1�2M�Q$���+T��]`v��"�	
X`7�Oy�kQXR��������-_Gv�7��n^P�2�H
p(���O,���O �4���������۝�|B��"��D�pkN�[2��aӮ�{�OLPmڅ�Mӡ�iI�S�g!��� ����h��
ѐtΛ6�����N�i����i��y�4�	:j�rhs�gZ!zPk�<O��$�O ���O���O��?�J��B������(6�X�������Iʟ���42���O�7m=��F�;"H��CЃ"r�l�V	�j�z<&�`�	˦�D���l�L~��0�L�c�Y!���зcܭV�(��� KƟ�R�|�P��ڟl��ןL8�H/�3 �_"5�я�џ���iyB,a����<�����)U$aeL�I�:Ւ�2ԡ��A��2���ꦥ��4`����߁9i�Z�"�p�a9��?H��8�&�*�|�����Ӑ^Uv�ɈL�=�ĭ �8��d�c-�d��ҟ�������)�ny��t�l1S&�T�`����#)���c�D�YSF�D�O��n�^�a��ަ��C�\r	�>3�<����J��?yٴ=�.hڴ����� ���n�ʓ|�U�N�_�V�j#`�������O*���O��D�O���|
�%�1I��K�)C���L!4d���K+E2�'�"��$�'��7=�v9��$3,���B�bÔuӔA��M�5�'����O��DcE�i+�d�K��P����r��`�*W����%D�y��e���O�ʓ�?�s�:H Rf�q�� Jנ�p%hA��?1���?!-Ojdm��8U�'��a� \���+!އa*�Z#���O̕'��'[�'���	�a�t�e�K�7����O��9c��gl
p�A�4��@��?�A��O�����+��]� nFތib
�O���O��d�O�}λ�2����E�R:�Xه�ʎ3ݞ�r�N�֧E�+�R�':`7�3�i��aS�?[N��r��kĜu�hj���۴3\���z�
-2@'x��Ծ8#�������3�ڙ�ȚNK�	�D�R�����4�����Od���O*�d�I�>ۆ$\�L��a��
>5��T��M�'Pb�'����'J�����"hqm�kH�KQ'�>����yR�x�O���Oм8b �8�:D.��=X"��瘹7��b!����d�~��$+��F��O��&�~�B��D� 0�bU�t~����?����?���|.ODHlZ"c�r ��6'���T�Y0:��kT$!7�:�	��MK��g�>���yҶi�Z��O�&ɴt�qȵ\"�a�cj
 G�Ɛ���&f�'W(��I`�����kJ$}�`��1���?�v!�Iy�@���|����������J󃌆e���u#���"䂧+M��?A���?�2�i�D@�O�2�fӤ�O�Ȃ�O54�LM�� �����(a��l�	��M���J�b)�MK�O��R��-3 �J��q� 	�&jTA����!���O���?���?a��R<u�'�X�p�ԍ�*U�2@Vi����?�/OX�m�3ظ�������IX���I�m1B�qei
Y(A���7��$UH}�Os�6<mZ���S�D�S#VB� �K�%#X`����c�8�`��*r�dQ�O�)$�?i�@$��˼Cl�̺'�δO���&�X5F�(�d�Oz���O���)�<��i{�2���TgZ,�p�S�%St��΁�c�R�'�<7�*��&��dæ�Z��P�>���Z ��(b��z1,���Mk��i�`+0�i�	�?~�z��Ov�'?����^�AC�Gn�':������O��d�O����O��D�|�tO��T}�G!�D&�0Re�J�o��66O���'����'��6=�.���X�C_v%x���%�-ٔ��ʦ� ٴY���O�� ױix�d�>(Oz1#g��tĪ�Y���11�|r|�p��P��Ot��|����01�R����H�`	�;4��Ep��?���?�+Ovdmڔk&��Iߟ���3.W����
׿Y�}�b�۳MV  �?��Y�,�ش/-�vi*�䆼$Wz�B2��4w��M��L��`��ɂiu�5���:K˜c>]��'����I$!���gB�B�zL��G(2���������I��|��a��y�/.e��X`i@�l���I� _�BjӼ�J0�<6�i,�O��W�N�C��)oQ�M��o����ߦ�K���McĢܹ�M��OU��S��*�O�?/��l���*c�V|F.�9w��OP��?!��?���?���&��(���N�p��v��5B��*O�0mZ; 7����֟��IF�֟��
*5Xh�o�!D�Y!�f�'��^r�֤�OtO���D�ie>�
�d���P(�R�@7�8D�fb�e�˓-��� %�O�-�L>�(OB�e�	ҍ��c��L�Q����矬�����	ß�S\y§t�x�T�tޡ��^�5��i%�T΀%�%;O��nZ@���	̟ �Iꦭ���N3a����2,S�oNf9{��Gt{� lZA~�왈a2��-"4�Oi��ġ*��<Kæ��L�%���yR�'A��'��'����
�p����j
&#���P�@+��D�O���Q��U"�GUy�Ne�
�OȔi�)��8�L�)�A�2�"�����Y��M�@����nD
V������)��3� ��w�?.��E�d���V�>ŉ&͚0�?A��:���<�'�?���?9 '�!1r`hlA:���`�O6�?i���ċ�	����۟ ��̟P�O� ��F���ӈ���t}��OJ��']p7����O<�O76��U��v�>e"i�%cLY�c�aA��4��(�� �̒O����>A�#��19�B)(3��OX���O����O1��ʓY��O�=�0��E�F�;!&��em)C���*�_�H��4��'-&��M� �z!��C�	����yZ����a��od��Y�a�|Ӿ�|#�틆I����O�Zc���p��@x�`�:By
�h�'~�Iß����	����IV���3e�4�I�#���@�syB6-ջZ!6�D�O���&�i�O��nz����j
0mb �(�Vy�W��%�McS�'���t�O���iWBW�V:O�И�F>���Q�l�
/wh�y&>OnD0bh�?�r�?�$�<����?�pD�1|�%8�#�/�0��gC+�?����?�����Цm�1�̟ ����"�;pp]SW��*����w�m��$���	�M���i�Oz��3�U�&&��2ª
{�U*��D�%������.�S��RϟL���oˠt��d����e��GM�����T���� G�D�'��@�2��=&���cD�N�v[�ٱ1�'��6-�V���PE���4�n�+sG8Z�-Yp!�u�8�w�O6�i��m�l٨�m�M~��\�Z��S�;�*��Q�=Ю�@���/,�n1��|�Q��Sٟ���ӟ�������X��Ʀ�v���Myy��}�\�{���O���OH����ܸ:��vƈ]}<�w�C�����'�D6�ӦU�H<�|���o���bCY_(Й��ԋp�܌�Ѐ_~bߏ�&���>s�'��I�9�*a�q!F�fEz���$�:���ʟ\�I��i>!�'�f6M��w�L�Ю+�����+I(v �jV&V�8�����=�?��^���ݴ(���(w�X�!$�8m¥iqEضv0�:%��(}6�%?�Њ��`��'����1  ��<m��3��[�L(��r1o|�����L�	��x�Iޟ��bT�U %��5z�I˛q��(�h�1�?y��?A��i�x�:�ONAs�T�O©9��݈g���Co�E,��]��Ovo���?���Y�B�lZm~2NM�'�NŹR$�A�g� �>��4��ޟh��|Z���I˟8����Z5���r�� �㭛�Pa2,p��\�����fy"Dr�Rt��$�<����Iׂi�s�ɱ~� �U����ɜ����Ǧ)k����S�A�
�0�7/��hZ6ܲ����o�� H:A<���$Q��Ӣ0�b
�V�	�!R��)�$Z!�����1o�y�	������<�)�ay��`Ә0���Pz1��l��I$5���	-e�V���O~Qn�`�@��I��W�0i���VxrQF���?	�4g4\�!ߴ��DK�)rde��'<�8�H���-�m��YV�T�B��IΓ��D�O~�$�O��d�O����|r�扳Z'�| A�Ěiʮ4hch�#T�V��%�'a��'R7=�D=)e�3L��EÝd��i�F�O���4��	Z��66�e�������|����&x$�p�l���l�(	��.�d�<���?9$�SѢ�1'�ىb��%:7Q��?I��?Q����T����r˄���	̟��7�� 1PJ*l�%�3,�x�[��ş�Iv≐h���"`Id�U�n_�o��4���+Ĺ1�PH~r�k�O�)~�P��c�o	B8�5-Q���?q���?Y��h���d�$oDX=Ѓ��6Jz&M�%��.���̦���k�埀�		�M+��w��c	�A��)m�	9�r�J`<O,���Ot������6M$?�uB���S�y�vL�.	�  �'v�P$��'��'U�'�r�'�����J/�Nmi�F0K�v�Z����4��]/O��4�I�O
|�W8;mX�r��E�tTc�KGg}��'���|��to��i��I���#�b�a� �(Ԙ��ihfʓYp� P!���%��'SL��A �)�@Ekf ?���C�'m��'U�����T�p�ڴZL����wDm�oG4+�~���dxL�8k���$G|}��i�`9mZ9�M���\^�P��BP=vlƼ�禋9R��c۴����t�r���'��O"��֪��Ta���t��t�r�8�y��'�b�'���'����W0D*q�կ�4آ,s�!R�p�x���O��D����k�K�oy�z�0�OL��*R|���7�B�L�k���z≽�M3����T��C^�&���Hg T�t݄0���Nč��
� �fyjw�'8�$�p���t�'���'�n�r��[,)�B v���d�'��P���4O7P����?a����	D9sN`�kR�'��x5LD�Td�	���d�O�7�A�|��ʛd�`u1�-��$
pY���;0����ɋ�x�
���l՟D���|B/JB4������L��+؈i�B�'J��'����X��j�450J�"���th2�Ї:Ĵ,S�� �?���j+���D]J}��'���@+/%�֌q���=����e�'�-)K������OI)5g�ɽ<��)�=Q��lS���KB��<9-O���O���O����O��'��-��/O�7s�}��?���M+�
�?����?	H~�� ���wB�Y-�f|����˻(����$�'���|��$��%T��=O� d0�f�	d�����5LjL2v8O��@4M�8�~|rQ���	���V��]���y�,:t���5�����	ϟ��Oy��p��U+�Oz���O l��� �jF@�����")��P�O �	����O���?�$J�9�L貢�;%�~,\��A�O�S�.cض6-AF�\���O�����H�9�K����A���O����O��Oң}��.|2Tab�I |"53b��9H_`Ձ�� ����2fE"�'c�6� �i�ݪrj�y������o�p��q�8�ߴh#���{Ӏ��F�m������xe���f����7;�*���ͮK$��#ʛ��䓏�4�^�D�O����O2�Dک,ײ]	��'c�>����C�!+��>��v/:��'�����'p���n�dh���3�EWb�$���>Aa�i�\6MU�)�s1g>�&T
�oY�h�(��3�߬�r��J*?��^?T�������$�f� :�k[�c�P�)�Iu�����O��$�O��4���@�F.	�Y
RS��� �0�@��	�y�h`���
�O�hl�?�Mk'�iY��+s�E�]�xH��+�}(�Fٻj�曟�����k����i��(0�!IӼǒ�a�CĆL�dy��:O6���O����O����O �?����^-�7�PC��k�O������T�ݴj�J�'�?��i�'�Zz���'2�9k�H�,�،��5�	��Mp��|2U	���Mc�O����#P.�����o����&��#?� R�5.*�O���|���?A��(���AbĜ/�F�zJ۸/�L�0��?q(O,4n�O����	��	W�4i�d�\pB$��[KLİa����Q}MӦ�m�?��S��ȹUi8}ґ���:8xñ��e���Y�+�:tʀ`�O�)�2�?Q�d'��B�1\��q-�*->���F��>=����O|�D�O���)�<���i'h�ɖM�.t���H��^�"u��l���'��6�:�	 ����O������aI�c�*�G�,��Ģ�O���I��B7M6?!GjPL����wyB�T_ժ,��k�Nv�h�����y]������4�	���؟X�O�V��f,ܛyz!��Q�"D�i��rӔ���A�Ov�d�O�������]_��<`�)E��pcĭڢ
���ݴG���%��iK
M��6�h��y��6&�f���� sV=*��}�xcba�I��`�c�	My�Oib ��<,J	��L])t�
-��DwQ��'��'��ɜ�M�6�Z:�?y��?� }�T��f�:X��r挹��'e��S|�v�m��<$���gF�ri�xI�"(74Yp�3?�l��bަx��
Nv�'lݨ�DO6�?IWƌ��� �'呴C����'�R2�?A��?����?��9��Y�fߠ2�ƥH���4�u�v��Ol�n�{t�'��6M6�i�I��Β@������>�J�Cc�g����4s�F�oӺXh�$v�j�@2���&䟔�閤�Mx�9�`�^9>��� i|q'�������'��'���'w<���#T5���X��N*0x��V���4Gl�qJ��?������<� ����Вl�2~ �[�g��0��l���S�S>(A0$�jZ�2נ�qǠ0����Q�^�$�b.88;���OTI�O>-Op�9GgF)S�0ڔ)����P�&�O��D�O����O�)�<���i�X�p��'S�T�%]2g���b�

�6���'l�7�9�ɔ���զu�ش,c��
��Eb����^�PK�<�A'&z�� �i���q����O�q�P�.޹��e������h{垾B8�d�O��D�OJ�D�OR�d'����@�d�0>[�8� ��4�|�I�$�	!�M����ߦ&��*�M�!C�
$M�t�@a����h���Gy���Xn�D6�"?U�R���\��b�7$p��y�#?1իE*�?	�-)�ļ<�'�?Q���?��W
a��1g�)�уԅ��?����$[ئ�������I֟D�O������]<yp�aG��좹c�O��'��i�ؓO�S�1Xq�K�	_��H��^hx�۠ʁ	m�fSPe!?ͧ�$��˂��W��("��m(�P��)���y���?����?	�Ş�����Rw�ĲS|�BTC��zt(R��/y�L ����j�4��'���fJ�T�)���	~ n���V!�6�����`2a����'�E�q���?�&>���V27t�yB4G4���2Oh˓�?���?����?���;>ժ������4�/.�HoZ(�������	A�s�<����+�鑤a���p��1
�bek����B�2�iFܓO�O:G�i���!�����͕}\��H�æ��O]��P���A�2�O���|��j�<a�$@Hp|饏�
�0�����?Q��?�)O$��	< ^���O��`��|pw��.D����@ܛq)�tk�O|��}��$��3f�	t�<���#�&�9��??a#�@�yr��#3B�/��'}q�����?�R�N	t!\)6Ҿ! du��(���?Y���?���?ы�ik>=h���p^��s�� ��,jB�O@1oZ:l���	ܟ�kش���y�@V�l
m�dɻtܼkĂ��yp�,%��ۦ�
�%_����'}�Tkd��?m
ч	%cD�0	G!�;����s��e4�'��I͟d�	ϟx��˟����<�i�f��+B4
�k�J�V�`�'�p7홞,T��d�O���5�I�O&�S�\ ����Y]��Rp�EO}��v� �Io�)�xl�� ��E��&׾x2�@G:!v�MI6�U�]e�����1e�Ob�!I>/OJ	��
�X8 ����K���:3��OV���O�$�O�<i"�i	PUa�'�]�PA�>����]�B[ ���'!P7�7����$����
�4Ǜ���cV��b
AtZ���HU�
���i���"U�F@ZR�O�q���Xt�����lj�XI )܊ry��O����OB��O��D6���T�����T�t��fl�5{�D�	؟��Ɋ�M{�#A]��du�B�O&�0.��e'>dz�$ VE��i�M�����lz>Y{4'J��-�'ht
'�E<h*PbvK�
mF�+���3\���'f��Q�앧���'���'dJ,�Z?9:qh��=����',rP��i�4=�x���?Y�����10|��h�4\��U*raY2v��	���d���ڴ ]�����bAD yS&*G��R��
#_�2����;@)a�b����v�R(�;P�'���e�9O)� j�D��C	B�2�'2�'D����D�'�Bݑ5P�ȫ�4H�tH�	�I}P��dG�\��@F�
�?���?�M>�������%�2��,&��ڣ�E�YÜ|	`�0�M��ic�1 �i�$�O�l��g�P-�̺攟4�&D�IF �M�/x̃CMo���'��'Eb�'	2�'��ӽL%��H�"
�l������7��*ݴ,�@���?���䧶?aѶ�yGG���,a��Ҭ�'FA�t��$l�|�&�����(�nr���ɺ}Y�����E*LӀE+ӣ=A*�I�:@\��D�'7��'�����$�'�0�Z�)�.c��s�Z�]Q2D�'�B�'wbQ����4~�=���?��7��+5��I0٪��_�]i���>)�ib�6��H≥P������Ty���T$xK(�#p�J�W�1��T�|�5�O�T���`��=b���#z$�3�N+2]����?���?��h����M�8�r!AY��@	Q�G���$���Ѕ���I��M���w�l�K�>/X��X��t�'P�6��æ�#�4?b����4���193�-���5V�
A��hP���B�	˸�*�B%�d�<ͧ�?A��?���?1�%�1y@��ir�Ӯ4��y���H�������������I��(%?�I�-I�}�!�u�`	+���^�ɪO<�o��Mc��x����k�"��EŘ0m�B�5��V�9U$�)����3N�:��V���OD˓gfx5	r@��,Q���rʃ2~����ɇ�M�v�+�?��G�FfKJ6>�^���*�;-:��/�M��Ȭ>i���?����*��W$_�hp��@�Y*,��U$�3�M��Od���
ĩ��d���w���3��@��'\�]Bl��'��R�R &��Q�
p,�r͋9n0�I�q޴7��u�O�6�,�$�'ws��R�DÉP�r-K�bU�|�6�Or�d�O�)�32�7-0?���՜S~����j��$�6,�@��6	&����� $�̖'�O^�*�K�6�^�c�F �*w�Ɂ�M� �����O��'�����,
$)q��b���d����'m�ꓤ?1���S����*BHK������\%,
�\��!��%�<�'t�	~�I�d�2ȉ�bY{�T�@��G�BC�	��M{0�B�*5Tő�!�2�N ^X\��o��Ċ�1�?IZ�\���و�BA��V��,���Y�qC�)���`+�����9�'�P����bJ-O�*`-�'mʍ8Rd��$��9q?O����=���x�L�:��Ì�@
���UP�����[b�Iß����yG)��m1@p��c^0e�($��"5_��'?ɧ�O��}�R�i��d܄���U/Z�@�h�r��Xp��*�'a�'��	؟���6Z@�0�`E�f��/�Ow~���ǟ��	Ɵ��'W�6M�~�6���O��$�/:V ȃ��J18��Yp�KL#G���ty,O���xӆQ$�\�f-N���`�D�Ό4.�:��"?�t	
-�|�r�U�')��$�?)DgJx� � )L].|"��ŏ�?!���?q��?���9� ��m|~��
�9�y�ׂ�O��mZ�
�`��	����4���|λoY���"�27T6`�e[��ϓ�?q���?���*�M��O�س�����f��V�
�*�kZZ>h����l$�';�Iɟ��	⟰�	ڟ��I�R�T��ŋ?B!$	e��x���'�p7-E=���?�O~�]X��K�a�/����T[�Q�U��Iȟ�&�b>eP��Zke��O��o.ҍP�Y��|4o����D��2�1��'X�'��I�60�9q���h����%'�N��	џ�������i>��'K�7m�9l&��D�&�Շ#
' ^��a��.r�p��*:�V�|�Odp��?���?a'��Q�� ��+JV�A�c�WOZt��4��$�5n�i�Ol�O&'�*U�$q3��8N0{d:�y��'�"�'Yr�'���)P�B^qX%f��=0�����?�5�i�����O��r�p�O���'�}��q ͂K�4Ey�8��O4�4��Dswӌ�c�&�鐺��Ql�8&���� ZO1@��OT�Oʓ�?��?��!j����Z&���i�h�`Y����?q)O0�o�Z�1�'�B]>�1��ЎED�i�0�ڤ-�0`�G,b��������O&�D&��?� ��H��Ϧi�9��F5(�8��a�
�4F�!U�cӞᕧ�$h?�I>iUB,�F(��&�2 (B|��]&�?!��?	��?�|�*O�elZ�=��(2��T�X����U�W�u�ƫ���I�M#M>ͧ8��Iן�Hg�I'8��xC`�ݻk4\��.�ٟ|�I�J�@��F�=?���e	��cy"[!�YP���x�P��@\��yQ���IğX�I��I؟��O_�H�W�\4
�������+^1�3_�Mk�_����O���.�$����2�N؃���!j�<3aBېY	�-���('�b>]S3��Y	�	�HG^)���,G��aU/�/*W��ɢK�`�2�O�O���?i�D1D���F �A������]�p�������?����?�.O�LmT8d��	�����1�0c�Ȃ�G�����&��?)�Q��s�4=��f#8񤇟hvŁ���<.e��+��/�Ɍy��dy����x3�b>	YW�''����V� c��²L�-�\�I��,��ɟ���O�O��C11M��C�S�BHP��'���wӂuxgJ�O���TǦq�?ͻM�@��
SZ���4gQ�<����+��F�|�6�m�C? `z�8?��G:0��������4:g)�j���E�L|	�H>�-O���O����Of���O�x0gCN�zA\��ۦo�8�ŭ<9��i66b �'o��'��Om2�G�zj&II3���Np" �GI�5*�~���eb�8�&�b>�p���=7�ԭ#B /�&;7�'85*�{sm5?v��Ct~�d�*����D�G����@^�B�Y q�T�i4���O��D�O"�4�D˓A*��'Y"92�Wrt<آ��$� �����y"gӐ�V�<Q��M���i�
���!U�|��܈`țsh؈`�ؤEP%��O���[ ���d�w4�qBtb��I%jmB�G'�N�Y�'&��'NR�'��'�<�D�H�� �3�	�8[Q
�O���O�`lZ�gqH��P�4��{�VuK`��;˺�@��5!�����x�h`Ӝ�lz>�ta�e]��y�>t�f���re1�ډ(�-�P�a���U�����4�����O���]-���� �c�\̊��4����O"�2���PM"�'"�U>yv�J�#G�y�C� WM�( �8?	�Y� �I��(J>�O�>A3+�p�H� q����|鱖�c�N�$�Ĉ��4��x��a,�O�d����'�����ٍb2~(�d�O0���O����O1���e�F*��v� BpgJ�Z� �#H�$��aa�Q�Xz�4��'�Z�"���8$2��eM_��@D�n�6MGæ�r��rr��l�+�f����O����d&�;�J��SC�?q��Þ'd�	͟������	����Ib��(<&�P5�Ȩ<�L�6e�#Ɗ6��$6� ���O���1���Oؤoz��*�Ɏ%{�,:�߾RNrɨ����M�C�i��O1��|15lt��$@�0�s�>b� L��Ɍ�*��� �fw��s��S�ΒO���|Z������-^��`9:�I	���Z���?)��?q)O��oZ-e���	ʟ���f� �uH�@z��c���1W���?��Z������sK<��LʒJ�nY�dc�y��㴥�k~R��1��AqeIK��O��i�Iw�ܑ%`�Y�#K� ��D
�@Cr��'���'R�s���!��Y!���n�����O�0��4 �qi���?q�iO�O�Ή�r���j�dX�H���d���-�ٴD5����NE^��O���|��S�a��X�Ӄ�-�5�T��%��EQ��|rV��ȟ��	ޟ��I���`p�@�g'��d�"m���h�IFy�d�vh����<����'�?y!�N�Ҋ��Ԃ�f�R�)��  �˟�oZ3��S�81���B�C�|��h�/K8���A(+/<��]�U9���OPLiL>-On�B�e�[�BE� ���t�8�,�Op���O��$�O�i�<��i9�[&�'��<�$̔�9�'.+�Y�'�Al�⟸ �O��d�O���Z�l�tiR�Iؒ3��U���H�UM>��`��&��I�n���ݟ����R��u�b��$j��U駡��n3���O��d�O����O��$9�S�F��P��a�'��)˔�8�a�'��t���8�.�$Ʀ&�T�uNº?���A��]>59nd����e�I���i>�Pf-ٝt/X�J�NI�W@O><rU����m��D���هw���G�zy��'���'�ҏ�?n$`g,�?n� 5�L�.�"�'��I"�M�Lډ�?mf��$�|*�]�J`٤ D3Xr��#@b~B
�>����?�L>���M�sL�6��Z%cǍB���D)�:$�ؒ�*uz�i>���Of�O���$O��v0	T�̯>�i���O[m�Ɵ��	�b>�'6�6�Z)DǼ���^�p;�і{�< el�O��d�5�?�!\���ɬ��ˣ��&�F%�P�l�L�������/Q�
�B�{yԠ��ĳ?��'�de����;;ب8@�J4�|��'�I� �I�������0��w�4��e����倗>�Bh��J-
6��B����O��$)���O�]mz�IBɆF�
�{��̧L���Ċ�����z�)�S)G����b�$��ԜTDi�G�x��@���h��IE�В��$+�ĩ<����?!��1-����� E9D�	�7���?��?A����$���2U�C۟��	�hh2��^��p��0c�*a�n�D��3P�	ޟ��	p�)� (���̔�4Bx����$�5�g�����ƤXw�QbV�W� Xs���O �(wNҊr_�AQ�٤�r�t��O����O���O��}���<�F�@�kͫn'�J��3p�y�����֠Q6Q,��M��w�8���D|f�04ʖd�2�'�b�'�r�ča�:���O�Aِl&���@�T�����T�3������R��'����$�	Ɵ��IƟL�I�j���Xp* ��Q�K�(
�P��'��6�	I�N���O`�$4���O� s��~Hѳ(�
��aI�r}��'�r�|��T!�)�>)�%f(&v���ƞmK@�cɓ�x*�	<;�iq@�OƒO�ʓ��a�F�W35 ��d�~!�M��?!���?���|b.O��mډEȤ��Ɏ)���yCi��g!���rm.���	��MC���>���?�;�B��dG+R���+ʬ�Z!L�:Hv��'V�YЅ�RIbO~����F��@
\"������(>�ϓ��?Ї���Y�$1baL&�����O
umڎd56�'*I�֘|�ë8�����Z�M��2� � O�'�������77G����O�`x��37��	�M����mk�͗M�.9S�'��'��h��9E� ���I!j���td�7�Fx�eaӖ�c�<����i��h>��W
N1>VV��$��$cE�ɓ����O���3��~��B�?��H�KA6+�({��'^nD�۲fE~��D����O�[?�N>����jl�(��ގ}�H��ՄR��?���?����?�|�.O�oZ2
/� Ӧ/WsM~�!��_�g�V��5�J��	�M+����>���2v�] d-G�x�8�AŞ=S��@*��?)��1U���'���	V�Br/OƔ�� )�$l�5*�^�B��5O���?)��?����?����I��d�u ҃e���� :����Ld�p�B�#�Or�$�O���D�ئ�]<�n�0��,$�0��:H$�	ޟ�&�b>�1N<:���2rL��HĊu��PC@���F] 牬~�D�Pg�O��O~��?��d5�a�LF�/xP�舚��(���?����?�*O���	�y"���O�( �by9aU`�z13��:��$P�O�}m�:�?iN<!�G@�6!Z�C��E�:�d5�M�x~�f��&}�a��&Q,�Ot�I��$Qer��z���'mΤK|�h�Ê�I��'�b�'��ퟬ0�!��a���2���0YN~��0�ȟx�ߴlqƑ:��?�@�i��O�ʤB���R͆2�~U��!��l�DP���Y��M�e.��%�
��'�(��0�Z�?=��!VG�ҁ(�=m��J �ܜ/V�'n��՟@���L��֟���%�tY�!3o���4�A ^VL@�'ʹ6��}�l�*���O��󄜞RP��o+��eHsO i����'3d6mƟ�$�b>�Q&ˤ{a��[�����`�]�#x=����iy"��w���I�F��'�ɷAF|k�e�.T�.)(#����ڌ�����i�n����~y�'k�,���f�O@kP��<���*')-7�J���#�O0�m�W��Sh�I��M+��'��L�1e �u �F_Y��QC��@�����X������i���F����.�.��]�'�[ ��%�V�A��$�O����O����O��$2�S�^�5ѵjR,��)1��V�EhR$�	ҟ��	�M������Ǧ$�X��@N'�t��Р .�K��%�ēa ���O�4�P�Y���O(]�!Ǟ�%n��ڝob�5P��՛P&�E��2�O���?����?	������GD�=�H!vk��H:���?a+O�������D�O���|GOI����J�$��`uZc~�n�>a���yR�xʟn��@��w��5�p�ϐG޵ 4�F4���#��fn��|�&C�O6��K>	�e��B�j���+k[�h����?Q��?9���?�|r/OЌm��H^<I��_�C5xxa5��#�6)Ia��ҟh���M��R��>Q��i���QI�D�3Q�&P4���D��O&6M?S�\���H��*�G��$	_y�J\�E�	ct�}��!�i-�yRQ���	��	П8�Iʟ@�O�~��񃀉kq*���A�;.�i�np��p�bM�<i�����?�Q��y�X:{�r�!�/��~��n��%.�o��M�7�x��D��(*��,y�'�J	�%EL�5l���N�R5|	A�'W�X����)E�|RW�����JR'gOr��VAN$iࠆ���� ��Cy�H~��	;3g�O�$�O�J�S�%\�2d��N�@<�a�0�ɇ����צ9�ݴq��'�L1�ɝqK�ఀ���F'X��O��ea�1�
�x!��Q��?)!��O�B��CJ�U{%��-#���5��O����O:�d�O��}"��v������;�v��vAE�&N8��j0��Q~���'4�6m:�iލ�#��.�%�[*X�(X��������OT7�¦�pC �?��,�`� ��0P�l�7tjHY�ŋ�T�z���a����4�|���O����O��d�'E��D�3'��Z�H��w*�j��\�F�F S���'q2���'�xd��:l�9j����S��PB0j�>Aa�i��6-X_�)�S* �,��!��q��$�,N'��4 b�1HJ�L8
�p$�O��hJ>�(O�h�1K��*u�!$�95Nq�(�O>�$�O�d�O�i�<	2�i3��
��'#�d�U"E��p�� �D���)�'V6�6�����������۴g�� ؀�IWr�s�����=rA)�>Q!��� {T�R�1���	��ʔ"���0AxT\`���%�2$��5O^���O ���OP�D�O��?�d�7?�Z�8�ՐZ�)�T���d��ϟ �4�Nͧ�?YP�i
�'n؊g�ĩQ �"en�)�djb!��L�i���|�φ�;�F��'k���M�64@yh�)=�H=��؁�q�	�v��'��i>I��؟d�	�lt��Dk%t6TP��^�#�P����d�'�6-�3��˓�?�*���{�GM
i"R��s�U�v��5��X
�O6�lZ�M��xʟ
�*�J�'!H�T��!x�mB&@/?�f�	4��DD�i>��c�'��T'���e.��Vh�1$�O�V�kcO�֟��Iҟ����b>��'(7-��A���9,�-����%�Q3.��̬<a&�i��O���'I6�D�N�DU�B��WI��y�O;�Mn���Msw��m}ޥ�'�.4#AL�?���&m�󦓅PiSB: j��57O2˓�?q��?��?���3G�ʡ2���:i6)�,S'�u��i�bQ�5�'���'���y��d���\�[��1�a��P۬q���lU��n��M[D�x��$���m�`��'W8U �F��Xl�G�н*�ϓb1Z�pi�O݃H>1(O���OX��$#E�,�hjE:M;�i��O*��O�Ī<ᒴil2}+��'W2�'��8��Y9tn�zE�Zt[�d�K}y�(�l#��NV�%Zd'�kxhMڕ�[�'�L�'�𼘤j�e�5���tSٟ���'�|�C�@�0(<�JT$��Ģ)	f�'X�'��'��>��I
4\�l����bOS!J��I5�M�S����?9�j�&�4�t4��'�<^褠���b9
��=O��o�<�M�D�i"���ٷ��$�/98�3��jxB<���Д+�L	�`f��m`f����J�VK�0�.�9
�yF�<W�����%[��a8⃖�yH6�t�M�Js�9`0J�<>�DQ���m�vp�ϔ8�,B��LϊQD��$��e��2]�H���@�[�恚���4OD��A+�+B~�T�ݣP'���H��Z��C��U�5㚛/�����N��Dn֨d�=X�e�7Q$���eJ6��
όp���8Y	D����=W���M
���s���Q�l�0�&����Q�2M14�pd�s���F�,~,}�)�)dZ�8�T��v�4s�̙7-���'���'��$	3?ٳi��H*� ɛ|�[6��I�'kP�������={���"�BT@Y�b"דp���	&?F6m�O��D�O���H�	@����,�<���t0Ȁ��:�M�fku�����$�
y\�hKDH%FW��3'�)&, �nҟ��џ`�@��ē�?���~�#�)T>�]r!��uĄ�@�F���'���y��'+��'�P���!�,X�t���~Y��k�2��݆y�>&�p��۟�$��؁E-T���B��蛡{v�Z ���<)��?	���H�@�0	�M�WH e�1�N�wv(���
P�ܟP�	\��\yrC_X�2ĉ�$ĕA -�j�|��1�y��'���'J�	?��Aa�OE�����#�dI3���Z��M<���������;��	�"�6�s�슘�f��V�H�|�H��?����?y.O��a!l⓸�XY�֍�Mm�NB�-D�eP�4�?������<	�O�L��O2���/�\t��m��DU$ɘֶi���'��	h��)�I|R����G�I3��RT�W$1ٔ��%f�)S�'c剒��#<�O�H�B�k��d`2���l �<p��ٴ��#J��m���i�O���T^~�	�Gx��Wg�e�%������M�/O>�;��)���*>x�G�	 ��e���{G�7튵s�H%o������џ|���'x�귫F�X�"<{��S�\�h02�zӀa�6�)§�?qT#ޭ^8V�X"���<��,�-��V�'J�'N��5I7�D�O�d��@���(_F����ł}�83#�2���R�&b���Iʟl�	�"���y��܍	@Jl*`��8Dw]��4�?���)�'r��'sɧ5��Wk�����m �6"`� �ʠ���əsY1Od��O��$�O�*6�r|�m�DFP����A�m�,���䟰�I˟$��N�	˟ ��A��*Ï4h��cW��F��Qo�.���?����?�����<�?9����El]ҥ��5��a��*�,5��'�R�'%�'�BU�T�!�}��A荓'Z��ˤ��9��P�`���\�Iݟ��'�ց�Op�&P*�F�1H
E���c�	��H��7M�O"�O��d�<bb�d��]�}z���zʠ9!��D�Z��7��O(�d�O����"{��d�O����O���#),<I���¯)�ٲ�+��%�<�$�O0ʓ0���GxZw�$�ȡMV�04е�����1"tP޴���1lZן��	Ɵt�������`JP)K�;A�Ar��6a��=���ib�'��b��'��'�q�FђWgӼ��P�I�_^�dB��i��T���a���d�O��D蟆8�'��ɰ:c\TX��@	5�NX�DF��4B��ٴޘ �b���OR,����$�� ҉̎|3>����¦��ܟ��ɛ3W��@�O���?Y�'`r9S#g�q��8�$�j�����}�cG���'b�'5�L��|��sv��]�F0�cؿ%��7��OQ�+
H}]���\�i�͘�+�
����B��.@`q+0�>��L!�?�)O���O��<i�Ѓ閡q�'(t�F�`V	�#fm�9�^���'M�|��'L§9� 
�ǯ]�V6԰��͛�T��P�3�� ���?��?a-O�1
Q	�|�!'ԍE�)p�˗3��y.�ܦ��'�2�|�'����O�����$�|ИU� B�P8PtL�)��������쟴�'�H,�æ�~J�$�����[�Kմ�����&$6P�&�ibB�|r�'c��ݾNPqO�)��@�]�D��a"8�Sǵi��'<剪.��Q��p�d�O��IV�(��^��`
y&��$�P�����z��8���4�.o�����C64�L9S�@��M�-O2��vJL��]�I�I�?�R�OkLəG�T�#��S^~D���.=���'b���sx�OJ�>�1r�צsY�QQ�ԬG���@�"d���f.����꟨���?%y�O\�{�f�Ab-�9P2ii�	A�������iN<�d)��ӟ��@��i<��枂@6�%�7���M����?Y��|�ZYb_��'x��O�}�𫊾DPz)!���:`�lzQ�M>����?������Ծa�tՈ���
���ռic2�=9����D�O4�Ok�����j$Dh�Hj��U(f_�		�b�d��֟��	ky��Բj�3�EG�9�!iFjՁ��!j�>�)O��$0���O��d�7Ry���H�\=R���K #b����5���O����O���^���3�Fa���{���DlT�?��4�CU���I���%�ؗ'0~TaR�'X���Z��(���L�)��:�@�>��Ӗ�6�'�>l*9K|�gM];I�ָ�ڝoRp��"K�@��&�'��'��I�����_��{�<�A��9b���i�ad<6��OPʓ�?�V����i�O���k,��D�5��x�	AS�ǵt�'���'�����lW*�����E�4B��IP#b�$�x@��'��	ϟ�w/�̟���ܟ��	�?͔�uWaP#̴BU`%=��t*�5�M��?y �1����<�~bЎ�(	&�5�� ��8�$�b�ئ�Cv���t�	џH�	�?�����ȨFQn�����d5�S��\%�6xm��9~FͣgC9�)�D������C��(�QM��B� P��i���'"��� ��)�I�l�dm�8O��,=T��)������'�
��.8��O��d�O��uk
�Jy�e3tI.D����E��I͓u�,��M<ͧ�?�I>�;��	�m��'a��*u��ts��'(R�*C�'7�	����	��ؔ'������=W��qb� ,��O����O6��?�*O�͏!Y�1����"��cԁM�Š�D�<q��?�����䉶r9Χ��m���D&2]�0�d�] ��L�'&��'��''削F�Q���m�v��iG"H8	SO9+�굱�O6���O@���<�b'DSb�O�=
��5�`g�2q̉�E�m����&���<!"B�:�?�J?M��֘|�F9{!��f�����y��d�<��i��� *����OT���\�#��9�P�*�fF98�\��xB�'q��)"�i�y���%H�5�F�����q�f4p�i��.}�����4O�S�<�S����ݦt|���H���)c�*?7F��^����#��1J|I~n�o4X�N���X�)#ig��"bӜ���%F��e��䟼��?e�N<�'@�2��	"r�ǈ^?u^��i��(���'��^�'?��pz�H2t�R�z�Ċ�6�m�a��M3��?��'�H�מx�O��O��tkC�%p0����3��AZ��i��T�d��T1��9O��$�O�ЭP�*ݸǯ��7r�������q��l�<�e`N����|*���Ӻ{#��.ta�]Rp�hq� O�z����P�����O�d�O����h�NA�u���3�-O�ص���Ƕ�'��'>�'��	�$�h{g�Ԉt���q��9\�)�QG��� �'�"�'��P��RT�����I��+�N���e� 2��\���9��D�O���2�d�<q�jʸ�?�t�Q9z�Ѝj��2D(�5�ŘG�'#R_���	&eVV��O�"��y��=���N܆�0
��4��78�	����>Eb��e-?��C<cU:$Z��S�7��J���ʛv�'��V��Bw�����O��꟬UY3D@�e��ySg�F+dP��P�-�k}b�'4��'N�,�'�b�'	"ӟ�iS�w�r�ę��n�$�M[+O޹�t	�ᦡ��؟<���?�+�O뎔&Z�b��
s5���L]fڛ��'CjV��y�L�~Γ�Oqpрd �#a)z��".M ��޴q8"�A�i�"�'���OĎ���D�pUحJ7�վm{���'�!G�!o��b���	W��{���?��-A�� s�2LtM8�1M��v�'hR�'�z�)&&�>+O��$���j�C�c���0R.�A@ĩ2��>1/O���g��������֟�P�(�#d�x��ܕ&��쁐��Mk�f͎�{�T�h�'��[�l�i���BMy6��0Ç+*��>��NA��?y��?Y)Oj!9���\p�A�fN 8�b�2%�9o�8�'{�Iӟ<�'z�'LlHO�Xu��qΑ���,^�ؼ�O��$�O����O��h\��Z�6���S��ä<P�`��Dd6����i��Iӟh�'���'L���?���������D��Z$KV�S53����';��'�rV�hj�ɋ:����Ok�gt�pa�Q�<�j�!S�ſrp���'0�Iٟ����0�pe����y?� :�I6�[�$]{�j�? A4�#1�i���'��I�H�脀����$�O��)۴_lb�1��j�T���ڌu�v�'���'�B�Ν�y��')�	nz���x\��)�]�� R��̦e�'����2ed��D�Oz�d�V�ԧu���!� ё3�I���;�L��M����?�&n��<1����� �ө1��� F*�F�ط GW6m
�Ho�֟���՟��Ӽ��d�<Ѵ]X-�!��(-tu�7��).���d"�y��'�B�'����JT�1�a���� �-*G(�m��	؟�Rt����d�<����~ҁ�#nS�� O -Y����M3,O����f��?��	��x��#n�n��D��&0�@�A��0�Iaڴ�?Q�&�t7��Vy��'���֟�ز|��܉��	H�.q�uJPA���Eϓ����O�$�OH�3`�M@�� ~�Z5�*����!���4}w��jyR�'�����	��h�c�'�b����I۲���Y���pyR�'K��'��	-}�"a��Od��3���@[H A�iƦ�@�4��d�O`ʓ�?i��?��+U�<�gh�
/������
-�52�+J�?������	̟��':��XaΥ~���/���02�X)�t���a�ʄ获�M;����d�O����Of���?OR�'���c�X4L��I	�d�9K�F��۴�?!����@�\w���O[b�'��$���i�
�X'.����ڇ(i�꓀?���?Yǯ��<!���D�?)�灨�"� 0�F�'嚭��g���Mh9��i�|�'�?��'Q��	�r�m[�O�V�`�S��˕5R6m�O���I#Y��$&�$0�ӱ;9��c�-Բ,JR���l�= 7�G�L��nZǟ8��şp�����'=�@�M��}#&4�q�	)���djӂA��<O��O��?)��;a�L ��ի|`^y�rڅߴ�?q���?af�L�'@��'��Ċ;�I#0�֗ ���� ć&I�&�|B�?r����D�O����EQbFB�9=�8�"jɊCpo������G���'�|Zc���+�D[഼{��	}���Oт�5O@��?9��?	ɟx
`əa��Y���P�jQ�� �͌; n�O����O��O����OJ�/	�r�b-�R�&8u�$��e��+���D�<a���?I����	ƾ-{��A&z�@��] `!��F�J�O��d7�$�O��$-W��dG$�E1&s.� ��_y�'���'��X��{��E��ħaQ0��0J
���v�Y)��ʀ�ix��|��'y�	�y"�>�E���O��ݳ$�ݼu�@i������I󟸗'��5�b*�)�O����&RlM��GU�I ���\?AH'�4�	�����ퟬ&����L�����F�~���!'�ݦ*4�n�^ymϥq307mWo�t�'���l3?Q�7A��[&�U�j�l��#Ҧ��	���"�&�͟�&���}z��� 3�T�z��N�K���ɱY��	xP!���M����?a����x��'L�f��̪@(Wh]K�d=�+���w��O�O��?���7wԔ@���]� b����+X�;GZ�i�4�?��?����E�'B�'�����N���4LR>&��D+�2+���|�X��yʟ���O�ā�1�Р	�jE���
�⑩?��`mZڟ�������'"2�|Zc&��##  ��X����S`a(�O�h2��O���?���?q*Ofi�$�1:�@Z��S�(H��D
K"d$����̟ $����̟X�p@�꽱 ��c"�4�7�6a#n�IZy��'���'h�IdX���O[ �G�Kz �x����q�ɉM<������?���.Ȉ��u�]���<X�P�W����R]��������zy�j�J��� �V�J�R���ǉ1T@������	n�������4*��=y��,H�8�qw�
'o����]��a�I�P�':���!6�i�O�	�,d PqsU�� a*ʙ����{TX�'���I��yb�a��$���'A����EԞOk��%��u�4oyyB�ǲx6�p��'����'?��F�r���B!/�vd��/	B}b]���I]�S�S�-����1��CP�%�`���q�6M��w6l���O����O����<�O��c �ۜ^Fe�0��b��Pa�zӮ��g.�S�1O>�	�n,�E�Ր
thaäj�!pt��Pٴ�?���y�FGh)�O����PR��T��ŃKզ�Y�&I!lO�$�OB�dv<��s�CW�X�"z��O$H���o���`I\�ē�?������f	<#9�gcH�F���AQe�o}��U"��'v��'t^�LRC�){��U�Vn8�eA�Z�(�J<Y��?�N>Q���?�ebD�&�z����B6���
r�z��<���?����?)�O�ܠ0�Oތ��FƋKL�PQ.J*#��ݴ�?i���?�M>a��?At�J�C]B�l��Z'b�ru'[�f@R��/��|ꓥ?���?/On@B��J�D�'+bU��Oތ�8��.L�HD[RdӢ���O0�H��7�I��������`J 3��b�h6��Op�d�O�����D�O���rG^i��	�C� 9��;��LN�'sb�'	���b��ʘ���ͣS��Ԛ�lT��!0$ &#�f�'��g�/=��'�r�'���'yZcn�93p��+7����Š
I�dߴ�?��4����Vj�S�g�? �HD�P2զ�)�,X�3��a�i.Jls�zӴ�D�ON�����T'��/z��e"��
8�>��b�3d��(�4'$)[���Ϙ'pb��Q�
�#�ݏFmʉ#F�N-Za�6M�O����Oh%`Bk�<�.���d�����`R�hM27�۠a~8���2��'�حb�	.�i�Ov��OLR)F��`�J�4{����ئ����S�R)�N<����?�N>��~�Z��M�z������Q�c��\�'"���y��'��'��I�����OI-r��(�Tnν]XX+��ē�?	����?��*<>�IT.Y^�h�T�P��Ȑ����I̓�?a���?�-O�yRB��|�e��9��x�g�J�{]\��du�I͟�$�`�	͟�hp �>Q0��6�����P�=x(@��b�r}��'�B�'z��|�b��L|�s%�1c*�ɉgvNAPէW՛v�'u�'b�'".�s�}B�>�!Qr�N( X�$@V�A��M����?-O2훐aYM����(��3aMǋUTn�����D�)J<���?	��S�'e�i��a��)��K�C�*pCfEZ�d˛&\�| !���MC�\?E���?��OQ� Ą�?���ۥ
}��ib�'F ���I�E�������ø��q�<Q��&��0"�6��O~�d�OT�I�[�e�
�AO!-��Dk�*��(þi�Q��d$�Sɟ����(&EpKG`اI��Y3��N��M���?��7���&���O�����p�I)5����t��W��c���BK?��������r��ҳM��Ha��M�)@�ՃqDE��Ms�]o�� U���'�bP���i���G�-l�����h��/H��Ia�����t�Ġ<��?�����$^*1�L���"[�Pɰ�m��9�0 B�_}2Z���ISy"�'�R�'�� �H"a�@�B��^=�uȅJ?���?9���?����V���l�'z�6���N�4�^�У��$V�&5ldy��'��I����ӟ�B�v�d���`*�b���l�Y;�*¥����O����O,�Gw^=xER?y�I���	�
�.�*� \譢�M��M����D�O��D�O�$Q�?O^�D��x�dM��2��
�&,'�5�lt���$�O��=��a�P?����H��1W6 ;MJT)v��>+�p"�Ox���O*��ʃFD��'��?�"��T0t����3��yh��S)g�2�1��+�i��'���O]�Ӻ3�#h$L:�I��δ�!�ɦ���ğ��u�q� ��Zy�I�381 �th�J�~t M�.`�m� ]7��O�$�OR���a}2P� �!���h��*��C%U��u�ڑ�M��<�����$-�Sߟ(���H�!dȟ�P�x�hʙ�M{���?��f�=�wP�ؕ'�R�O�I��*�55��2�*�%�@�i4P�P0&n��'�?����?��
#)
ܕ�����JܝH�6�'�hBo�>�,O���<����Q���Tx�gE�r�AI�x}�E��y_���	ߟ�%?�B��>UKpS��K�:�JH@�ꐃ^��	H�O�˓�?�(O��d�O���K�>m9	¿��p!�R3p��z�<O&�D�O2�D�O��D"��a���x�®B�3�$�(&�7rQ�J�e��M���?���䓕?�-O-���iL��P����o8�!
�4��L
�O���O4�D�<�aiF�C����Ps��T1��2���7�V0X'���M#��?q���';qO��(!�&��]��U)�ZLX��i�2�'|r�'ª��q\>�'��T-�7
���D��#㤕 5�P�.O��D�<!��Ko��u�+��A�5#b�ܰ*Vnύ�M����?Ap����?��?������?��/F����^UZ�q��(.#�o����I�"U�#<q��4k3pUqF!L_��H��S��?����,��s���0=	�2�Fm3��V�"���[�<��`�5?���ԭ
�.3Y��[�0k�	S� L
Aɂ�J���.I�թre�?+9�t�U��2t�2Q^�$C�����U01�`)��DV=��՘&�>LpU�����ZLuq��X�2P@�P:%�0��a'Q!ܠ5X�� *d �#���[4:��g���Px6�Ĕnv��k�
�?���?i��Z��.�O��D|>��A(V�S[��	ďRI��\���N�8C�	I���P��͘�-A�k>����D���N�� �D�e0�� ��ph�/T�.NH@���Φ�#��9-$!4�E���@J<y6hFW�¨넅R0��[2�G7J�(H�	��TE{2���M��A�14Ԕ���bM/'!�֟pt�-;���<<���Ȅ�p1O4!�'��	D=�aB�O �]�2mb�0��+l�$1�V5^`�$�O( qi�OH�z>�I���9'�ڝ03�خ�~��'�2�Ѣ�"o^ � "O�p<I&��}��� ��K��Ӆ!/�k׃�}�����a5H �x��]��?�����d�am l��/�;M��&T�	�1O���DR�
n��0��F/�r���9�!���!۲�
Q Р�0k��~a"��̔'�~����>�����	��U����Q�KG�-�샞q�ƼP d��X<���O�`��)d�AI��ͅ0�?�O*�S�4mj��#��#�!��o��G��'�
7	Ҋ8�i��  7A�>)����'`�n���՟5H��d�)}b���?���h���� ���R �\x��נJ�<(�G"O�9rǃ(l%�1�դ�,��P�'�#=i��Ɉ!�Ȁb��x�0/��W�����@�I<M��T*aŎ����	韄�i��F�c�N=b-���@E�_t$�A�^�L���@�b>�O6�@��*2�$�E�a��e��tc�+�O6��Ɇ�и��a�H)���D�A�,Igɣr�������$ʒG��O�ў8���?np�⠅�l�ZCe=D�7e��(�jm#D$�.��kpM??!��)
/O&! #�ǰT��<�1�D�9.8��K\>����	�Oh��O��D�к���?��Oz�Iᇏہ;Zd���̆�]�D� ����x�k�&ɠ�x�E�)8������*F��@	�'Ψ��vC�3H��Dާ���@��!�?��o1t}B�N^M8��r��	o��)�ȓc��TKQ��p��(���X�dS�`�<I@�DP��l��t�I2Y=L)z�J֓x`>�kƪ	#"z`���<�`����	�|Bq�����'����^��YK�O��1��$O��� �Ĉ3m���0e*T~�1���Y:�x�C���?�N>��X�C��t�!��?D�����J�<���O'	���
�o�\�z\@b*�_<y�i�x<YӣI�_X8!B�P�"�,[�yB��&�듓?A+�������O�����0-q��;1�[I�=1�	�O,�d�*$W"����S
#�:\:�f��$UJ�O���*���Ɉ}�.��v��;F,�'����+[@x����٘*�>�PBI?�/2�X  ���U ,�LG�<kD�'�F0p���?1����OJy8$�D)7��$�p���F}����"O$�ڷfܫy��E�D䄽d2	S��'�"=��ɝ"i�)S����>\�V�M�.���'��'�H��)N�'K���y��N���8�cd�+ag �*�C7.1O�%K��'�(d`d&�/&�v!�eGZ�xM�{�� ���<����;&�p��)�="6�P� �.��'1�P��S�g�nM6T+&ܠD�!�kֵhC�I�9r@���F7w�Q:�+L���ߑ�"|"u�T�Rr*�c�I��u��c���72�+@��5�I��p�	ݟ��_w�r�'��	:*��:V&�#����1Ό@!����Onu[�/�B�6�{t�~���e�NM���'~$�G�֨E����#��Q�� �r�@�?1�Z΍�wE�C
z�3��D��ȓ`ߤ���v�9��ZB
"�I���'t�ŋ�m���O�<��	�5�L�5�F�3E(�%��O���� �|���O������'�W�+JXy:���2'�4�A�/��x�E���'[jE�w�ϭ���� #L����<�Z�	D�ɷM�x�It�˵{��HK!\�M�~B�I�( 8Z5�V�3YPc�x%�B���M3��A��0�⦭4 xٓ3��P̓UZ�h�#�iM��'��,s��0�ɯ,�|��6dI7N?V`Sb�w�^��	ן4���<���D�!+�@���*u,��P�o�a:2�Ex��A��uIJ!�ߎ{|�Id���ɾ��<�)��&.#x�[��� _,Ż��Z�;a�C�I	
��ȡ�����2U0!M������r�'�Ѱ�+U�4}�<�u듾w��J��i�B�'��n�[Hؠ��'d�'��w��!!3��:��Ų���E�<Q��i� OP-�P���_M�S=*�1��'Yl��RP�?���U)�I&�����B��	��ȇ�j�T��DU�����X�,)	ׁ�?�`y����'��"�i���'^��C��d�'_��'"��'t�T ��|@$"��F䰔btO� �4ƍ�EFe����r(�8T��p1��d^}rX���	@�t�CΙ^��q;5!̐\I�D0��şD����L�I��u��'\r�'B֙(�0f�pxD�63e��cT�z!�DD+W�,H�t`�]e,+㎗�(�4��F�y'�ؖ��h؞��5� "l���5�ٯnx�X�Q$L�R���d�O&�&���Iɟ,�?��_�K�
M��&�Hwh�`�$�]�'?H����0I"r��#�pd�%Q�c�6wfx�O|\m�Ɵ�'��*�ê>��[Q�5B��D��l�@���Z�,�i��?��b��?������n� ;B��#��h���#V�6g2��S+<�,��K�<����9%������)?� ��D��:�p�	�D�6z���b�1�@x��'�0����Uś�>)�N��$��Y��҇w6�=�� r̓�?1�S�? ���CƘ*
�D��jͩ4�Y3FOulڮXq&��$߮6D��RE,E3A���IG̓�MG�,O������v"N<A �D%�$�P"O�e�ņ(yL�����15���"OZ�r�$��a8�b���x���1"O^��s��PH���	��dF��2t"O،���^e\4\@R�ѩT1�t�"Oԙ˵B)s"&c6-��':H@�"OV`��S�eX h�Ǭ\Cx$z!"O�<b�E��3��\4��$�@"O�s'/�b|	��j՘||ȕB"OT�"�ч�$z	Ɯz�)c�"O�T�G.�k'd`Sw�;<�v�t"O�Rrc+C=P��Wf�)��u"O�a�'j ������I�6��"O�أ��, ���)]ְ�a�"O0X�H�)�(0"�b��X�.�+1"O* �H�.0�%�Uo�"P֬��"O�,�S		 d��W�ϮX�"O���0$�7/`�}r���"� �a"O�]��C�$<�1��D f�2��T"O4�$f ;S���9��o͊�"O�Qu@�)W�$�̟\M��T"O6(��mE5Q�d@���_�7O��!c"Op�m�%K�(P��W(B�y�w"Op�ǁO:䒼�"�B�����"O����ȏ,v(1��O+/�nXk"O���d�V4V����wLJ�#�Lec�"O�`���%P�� IE���X�"O�5ۂH�.m&A�e��4+�8Yɦ"O]�&���u:�ad�V�z��Qv"OhIg΍�M�:a��]'f�D�D"Od��+�K���%��
K��2"O�� v�
+/Jؘ���٢g���0b"O�p�/A��MJ􉍢~��̱�"O��Rg��
�p�@E��#'�n�$"O���� ��Xh������+y�]��"O��#�D�'��S�PE�x�a��8XD;B���t�/�g~��ԗ�tqr���6G��v@W�yB[�&4�&c��ID2�9�. �wL�e��aCn:f���)�����^�*�@Ra�L{bͅ�	b�J 鰈\�9���ɣO��]R�E�d�zi���)K��C��/�(ؤ��G���",o�zc��ӄ".k�j� �#�'TޖHB��)��M��Q�S2���a¢�ys�Plpeh��A�`g��R�,ۚ3�q�'��@3��0�^�Z�<�7�*$�j2D���[�3��+0��YN:!��͹zr�x� ��;�����$Z9򜃗�/vȉCr�4:=az�Ȅ?���s��y��C7L� �K�^P i����y�&N`�p}	�jL�fr�-!��'�v%2%-#Ed��A��IK�N@�1%,�.����C��x!��˨[D��EI2޺ЊD��<�����D\��'zq�#|�'��9Qe��c�J�����y �i�'j���ŝrb�����Ml8s#�"�N�i�F�0>I�!I�}�4�E�8x��D�T��И"l�	됩�Ek��p�i˝hٮP��`H�M8]:�(D�����&�R�Ӂ��	�LXj�*��
�\x*e�˃.#~�Ă	>R���j��c���X�o_P�<A�b�74�� !0�U�/
����J�<iF ��V=� R��$!}�t#Ch[�<��NѨN�كa���5��h�L�<!�,�0?�`(��D!cT\y!��GR�<)#� <�j��D��Y�a��L�<�tE�>,�5�A��!�di�'ɌK�<� \=K�?l��ّ�X�����"O�aХ�N�Sp�%�I"p���Ƀ"O8aևI�[~��#��>���q�"O�]�g
^�����w��A�Q"O��{dj�:��P��>�j�C�"O�pf�-|!�,�3�_�����"O=�p�^8M�R��f	�	�|�R"O(ě���m^���V��4 �����"O�M�2�	q��Y�b'�"ai��� "Ozܚ���8�0��֏�!gNr"OdT�Ջ6ɞ�Z��!6(:|zW"O|8����"��;p4�U"O`5!��S%`�@Han�Ct��0"Ob�Z�GX���1G(z����{�!��%A�����#cK���n��%q!�Y$��X9Ff��:8�����\W!��ƞ:��1��ȝS(n��P'� ':!�ğ�#>2����ǜ#
���f��O)!�D�-0�fH�Dʅ�;Vnd��,!�_(���q���>eCr@	ep!�d�M��ˡkI��D����� ��<����'pB$��!O�P�2�b���8CF�
�FL��I�=ƪ��aًD'����Ҝn�z����&0��' ̪����z�)����w�ъ���^���J��I���p0!�I5x��q��2Vt�O��2�4�)�.�ꎾ R @T�])��'�=@!�)�'v��CQBʀ8��TQ�Q�7\T�!�C�T��'�D�G�,O\��go�7���BEQ�Ig�D�C�O��A�O�צ����M&�p<���ԤJ���a�M+�ʄq�(�y+^l�p��=Q��#?��&�B���qbB%<~,}�ʂ<�l�UN�.,$t�c�3�D�l�$u�g��`,,��C��m�ԟtȠ���?�@9�Y�!��y�D剥Ld��3��;�`y4�� fe ء Kc �-����#ȎbR�]��e3
�|O\��S��cH��S	il�)b	S,X y�̉6[D<����G��M��	$g��)��@�`�ɽ{骰ZS*-Č8��I^����u%�� EĘ�[�`֝5fw�EyR�]yh���A�&�2�5�B"����ƈ��pq(�(��\>�`J<�T�A96}�Ŭ
�\z�)�#Ư^Kv�:�����	����|�pݨ1l�s�#<��.!F)bAS@��d�!&�\�Ed�Ȱ)�c^�+��f��O$��Sd�+pL��i����V�6d@�D�I?��O�>��-υN�����W�:��,)p+G�T�X�u��?jq>T���iP�>E;bA��U�+6!J�eF�Q�'��0�%H�M�Bs��q��ϻS�MЗ@њE۬ԱF���Q{�!�y�4�Ko���10�w���S�v���ω1A��lq�G
U+ 4���'z��d�6Wop�R1��"٫&d�?c�@��'�3>�t8qNў,.�#`)�|tr���A��͉b�_9�RO���t�7Jz9l̘��jM�L@�O
����֬)�:���L�$Ty�#<�*�6.+�����][����-�|P>���!
Ypu�� 
��O����QTܨ��ڇ�:�"@Y�擛>��P(�	̒E�7Óc��p$��Df��RTjA�4��D���I1��DnV�s�-��_2y�L���Ѡ.dft;s�"A���)�S�yW%<����A�T���e����5�*B�}���	���a�X��;��99���d>yf�т��Оs���_w��D{���1�Ä@[;Q�e�M��t����'�z��/ڲjB������	F�9	���.y�x@*��#�z�\�)�p���r1�Ys�X�����*}=S)�f瘸r5-���1�R��1A�b�	��%����ZF�R�3�\��J?����6 ��`�bS5q����u�#�ts�MCҀ�2"&uS'h:���45��KSi%k⎐�R�5N�PM W��TUP� �oe�PD��O�Ă`&N�"(�a�2N��VІ}���OZ4�ʔuJ<�¶��%�0|!L����1V�k$&q !Ц�Y�#ɅX���f��� ���I,R��x���SQ�!r��^1��b�(�������K�¨�ם~r��3Wx�R��C2E�I �h�\z��Gn\!� 4��ǋd��p�cEBæ(y�M�3
��5pw�ÜZ��Db��C����^����*Ҹp���� 7d�d���2qhNt���S	c��E4������Rg��*���(�NŊ&�^+2	UV]� �D���R+ԭkt��Q?�V�>����m�fś�������#��w�<Q��/+��X�㜘�>�xd�ͦ���m�{���5��U��y���T��&M��3U� ��=1��	!8&j��D�g($@;@��KT�R2C���Ԙ�F24�� ��Z������W��8Hz�Ѓ��_�X��@c� �Q>=I��Ҹ$����*"��J�+0D��� , �U��ev1��a ��>���'�Ȑ�q�D�i@Ο��|���.o���x �'P
8l����@��,���,{�0�P���B��"ѡD1*3t��w
RQ7��=E���s����W�9���1f��E���G}�`���nً�dD�zdQ¡Gcr�kea���~��9b�8��4V�x8��IMƖ1PK�u@��	�j@:Hr6�)�)r�K	�qH�牪s�q����.Che� �ə\�.B�I	U��@sgπ`� ��F�/>��'� a�aA�Wl�k!j�X�S��mC�\s����ګZs"l�$�3�p?�aLK�	�b�X�R0i�:C�Մ-G��Zc���a8<%��0�)���ґL�>?S��:tj�,S��5!���ͳ�%�n��VV͑�I2'J�zA̀5K��'����əSN8�kF�Id}8D���I5X;�mbC�"�)ڧ~:�8�߷,n��˘%u̸Y�ȓ
�\zu�G��P�C�"W'�ႇ	@>���	�E�Z���G�hND�+a��
�'^�������"�R���+�,q�� ;�'fv�b�$]�h����e�y���dF"X) 
R���'�lQ!ІCZ,r�*�1!���}KS� � �4 (`Cb$9�'��%�0ɧ=ɧh�<��%�*����W�U�l��"OƩ�l3�И:���Vu��>q�]9 3���
�Ƕ)�G�Zj�F��0���y�@���2T�L<�&ܑ=b���L��^�Jĩ��L��=��)k0Hɵ�߈xЮ�	��L�M-�mG}2��X��ȇ�	T�Sឱ���ɫi,��mH5V�!�$��2��W�XF��cs	)Y�^���r�x�rrG���S�O���� P)p�z�C�k	K�f��'�&�@s�O;F�F)���.G����L<���r)),O��Sv��(*(��	 �$4���U"O@�ʃ��S2���(�ho�t�f"Oș���ۋ"dVPr��� ~�P�"O�Q)4�[�p�A���Z�$5�"O,0�)"<q|�*r�� 9�D"OV�� _��P��BEy"O<�iea�F�8x���-?��k�"O 90�
�(O\x@��D�Hks"O�虷�K�?�|�/E�b�0D��"Oz�:�a�$���{���T��t�Q"OjxP�Ł�a@�c�1y_��0�"O���C�Ι0���p�ၑ==	�"Ox\��AT�tQ́@7�7i6���"O�)�RKD�SK=Q�	
��p�"Oި��k�2"G�p�vZ:u�f]�"O�m�F�ܙn�@[���,��Qd"O�0,]��Em�)���Ӣ.D�D�r(C�D}��ɘ8QG�e"B��o1n�{�)��]������00*B�I�/�Rq�X!_��mawɞ0k�C�	8����W�������G	S\~C�ɻ9���Q�aG�Q�%�6G�$�<B�ɒb<�� à5�Vye�8B�	�Js�M'�ef��`-�' HB��wD�p%��6 c\���C�	�4ìLja�M5z���/ �L�C�3i �� *݄8��q�Q��0��C�	��q!Dȟ�
v��H��r�rB�	M�h�Ǎr⒬���)T�B�	�^�:�J���Qt4�#�R�|B�I�^7��teY�]�b\�Nsj�C��kP�@@,R yh8C��:]_zC�=)L���I�0AyX4��*ޫ�NC�)� ���@�ܑ��â#6�2�`�"Oj8�d��R페@6��dXB�"O�M�`E0�l@�J�d� "O���4
�:ʌ��AN�'�Q�"O�����7k6��ʇ��x��q"O��3� �GS�U)�oCYy�TrU"O��b�-2]�	�0�7re�s"Op�j"$��<�F�R��13T|��"O�<�Q���4V�P���P���"O0H��Ih@�rb�>oN����"OL��.�= ��t
�730�}�"Oj�[���{wx���0D
L�2"OzqC��/:�(਱�7` ��"O�XG��-�<5 FB�%gc��ks"O�4%"�?
�$��!�ULX��"O�Œp"��xPRC��1o9����"O���u	ҙE��a��
�9.\�f"O��(�[�NKV1�Ώ�62�[�"O�Lb�a� _;R�{W/�g�HĪ�"O>l��Y"el@�$�&aʮ(�S"O"d9N��0�*���㟴���Q"O4$s�;N��ɻgCރQr��A"O�1� |$Lu�g��;3``S"O��!r�3HVl�J$]���i�"O�񀐍X�kz��n�!�,��"O��N�3�Ġc�]�ov�s�"O>�!��B#㦉����-/B�e#S"O(Bnۛr/�c�a�1.��"O�S��רk��	�2.���0"O��2Vc�!f,�ŪH�&|�)[�"O�q��۠%
ƀR�A��L2���"O��cj>-��3� ףN��k�"On����0�-��i�4)�"O����� M�L�M�2H����"O^ ��΀�����	
!&^J!�"OH,1Ѯ���F@`�EP�)�Z#"Oܤ�U�\�O(��Ņ�&hj�kD"O�Y�M���t{���!:hx��"O�� �␎K\ �f�Z*&�N�S"O��J�,�?�4q��A����8"Ohqc�S�^���`W?d�$"O�x�����O� ١���]���"O�HeB])�6題|M2�)E"O��
U���<3�`:
�+/(4�D"O�|�weǼ9r)����A|r���"O�U�fo��
���c+�o����"O2���mUy&��R� :q���3�"O�pp�#r���E�9,戣�"O��	4͏�1/$�Q�HסW��A7"OH�x2G�RF�zH��kn٪�"OJ\�7*��&�6<���!#�t��""O�$3�OF�{Q8������t�H�is"Od���k�
vX��6/D�v��Tk""O�x�P�?kҶ��d$�7�tYt"O P歃�t�X"�?+�R��"O��[RM��"Y��$�ɉ*�p"O���x�۔)�w`�]5"O$�KqOP&<
�B��	DXq;�"OJ��U�rpNp�I��<�m8�"O� ���A��� �1ba���[�y�䂁)�.�8�&��Y(�� ���$�y���CT�rD'��
}�qG3�yR�
I�s�
�|���¥H�y��	:"/�,�$C���@ƢG�y
� ��C��ĸ,���0(E1
`41 "Ox�C��:%j<m2���;$�
W"O�XC	���9p
DZ�h�t"O���Nz��]2B)�q
��s"O�3�j�SԾt��g�D��9;G"O���!0ڨ�{�EƂGڒu��"O�%���Q*[���n*݂�#5"Of�p�?�4�A���>�P��f"O�a�` �BJ<Ժ��2�K�*�yrc�]��@�!�CLO5�N5�yn�NKF���)W2i�jW��?�yB)�3���a5��3"���Q��L��y2��6Ks��agH��T� �)�y��%S4 ��BhpՈ
�yB&K��`�V�G~�Eߨ�y���Ju���/ܧS^��Y�.�y"�����������g	֊�ybۖ(cda����:s������y��, vy٣gŴ�BD��cS��y2@�D���m�Z�+w$���yr&�(<�HؕF]?R� )7-��y�o����i���B�6@�*&I��(O6����_�^��F�S
��s�jG3G!��REIv S,�>5͐�P6ʕ�9!�č?E�|�WjW��vD�b/�� *铨�>!f�_*��-�čD/K�8��U��C���!�����A�l ؜��)K'-��eK��:D�4�qṀ;A���`�
�s�<]���3�Vb�D���l�(q	 E�${�,����y��˫B8��5��<"��r!��y���>8��W�7ޚɃC��=�y��4��`P��߅'p%Ȃ�� �y�, 
SÌ! �I2�� ��yb%�����*���(2k٫�y��Tl1�A��}� ���G_7�y��΋*-��Y�HEGX��Ј�yl��k��X!�!��:�^�!@Ԑ�y≓7X2`��7�`��JI�yr���}�Q����e�:	��<�yH;z�< ђK���|�ae΃�y�j�����"HL�����1B�=E���X�RD�����L��X���z*ȇ�[�8[W�E��V��g��\ 0�ȓ[!6JB[�iq�ԣP-ˣk�:̈́ȓ/���gZ�V�p��a�H}6B�	=}�͙���p[��a�bB]B���>�H>9P#�' 乹!�3*^h�r��f�<ф�ٹ3��=��M���|��O�L�<��/Ϡ:�rp�peY�
�� �H�<Y��B�pM�uPHL�Z��M�`��\�<��2�e�!j1:0��&�>Ii!�Ğ<	�.�P$O�6,0��C��0Z!�$��8Q��A�'��M��vH!�RQ� �P�ƛ`�����FWU!�Da��oӷaq��&.��*J�Q"E"O&�Z�	X�_X80��N�*6�,�"O�͉������M �h�T����"O�U�T�S8v"�H��C�S��33"OD�����;|n(�!�'V�(�u�$"O�T¤�ŜH�H��a����!�"OdC���kǠ٪S��
��s"O�b%G��|t���i�l�B"O(�`(`-�QѕaP�:#�1""Or��p��*��u��Y�u&���"O� �YE*�2�X�*F�Hl�*��"O(�
��ªS4`B劇��1J "O�Q�'���ޘ���ʫ[���2�"O*���	&7��E2�q�� D�4��)ͧ0Aj�zgG���͋�1D���U㐶�
}��R"O�es�@.D�8���E�G>b-�%ύ=ahA+B0D���e�Դ`�h��P�0{I�{�	0D�h���[ ��ZƆr�fQ��#D�d����FB<�1���w�2e��C'�􈟸%�2�<�� ��,wi�Q8'"O�!K�\O�u�AB�T���"O88���=a i�b]�zQ��G"O����_���0@ŒjJrTk�"O���0K�����$��+���'"O(}k�L%3���h��ք2�"O
����̔Ȁ�Ѷf"K���8G"O6��g��U]� �F��HjV1i"O��g@w�(���GT����x�"O�Tb�hV;.�����+f�Z�q�"O*��7K� ���N��C$"OB��P�@:k,Ը��Ԝoh����"O�\6&#T��TP�x�ܠAe"O�%caE8XY��4n6e�2��D"O����aFA@|�7#:� � �"O:`�C�
@�R�ʢ�
5Ӡ�:��'$qOZ���n]�]�U���64�0��"O�P��L>M6�8b�P����C""O�49w)���Y�p"����!"O
i�dH��z Z�Z� �6� ���"OШ���:�@����B�C����"Ob́��QgZ]Ҵ��� ��"O�xCMڧ`�@x(��B:W}(ɊS"Orp�<v1ΌK��P�ko�U��"O�0�h��G�̳��(ø��"Oj��$��e��)��̺e��A�w"O���SL��#�m�d�\=���8�"O~Q�%���d�%�Sd�0��W"O9���=+D1�r�Y=7o���b"O��ࣄ�5	�0��	~��aU"Oֽ3 ���z��#<����"O�đ��ξL���j ǖ�S��8�"O�سU�lܠmHw 
���b�"O�0��i�I�n�7ŀ}���I�"OԴ�5�5�`0�aD�S"��2"O�,; :IP���+Qr�*O�����7'h!#�W�l:���'����ȷ_��Ih�MI&b�b�Q�'�Rl�t��,N�PA���D�nՋ�'��h�I��8���0�N�?����'���%��@�d�W��H�Ȭa
�'�X�:��߄����C�4>��x	�'l>�P#�V�6�q�S):�Д��'���s���M��a�@�~]~H��'�����e\Z 2��'*A�h��';,h�#��;�6�zЊމJU�� �'���ۦ���lȉ'�F2H_�4��'`m����{�M���Z8:��Q�'��lZբ�U+HcD�(:����'���D���M��!˳㉯�����'�ڽ��b��&LZ�k	�b��'�>�i4E\�Zid�P�Ǖ����
�'M���ł 2%��� _.,��'[���r	�3ߴtA얬\�t���� �5�HW37G�y� ��<AF"On�	$K*.n�S`n���<���"O��+��ƺ����#@���"O�tS4@҄R����֢Ąe����"O�xĎL�wb���2GշM���`"O���a-�#"��-HC��J�b�R�"O�%;�&֜!��Tsw	ʃO��3"OL�b�^�5�ٲ�(Q��T�(1"OR ��Wh�) M׏@�
d*A"OxM	�HK��Yu���F�(�"OJ��
(i�̬�G�U&`7
b�"ON�9���
@4*�%����"O���%���"�(X�Y�k"OF�aA�V�n�jx�G�+,����"Oޠ�W��3$�� ��;@�
1 "OJ�VÂ=Ft��Rb��cj�:D"Ox��7�^�"�q#M1�t�f"O��CdX�O
j�A�{ (3u"OP@�S��*�|���oJ�VQ�!S"Of<���F��f�a�]�/;�( "Oz����V�[Wz�ϝ�:����"O�P"�ͷ~��	K�`�!Yb��"OnDR"o��$�m
���8���"O^I��Ь}⁮;�X""O�Y��J&n��ٵ�ɭaj��"O��)dj�1/(F�8q؂�,"�"Oi�t�O$�<u�կ]�T��Q�f"O0 (����U�(�� E	R����g"O���֪a��!j�i��	{T%��"O�F��)���A��Ra^���"O�8����-o���B"
D�^U"OT�TM�,&�(�LU�љw"OP�pu+�4R�T�S�A'C- R"O��� ��7c|qk&�R�b/��"O@XY�,�!g��1\�9��I'�yROL�F51�ÞZ��i�#�ݛ�yR��+eT@9"�`��4 �m��y�AW�M�f�`��:<Pá޷�y�#��<kX�)�D�.)�>���]7�y��X�+i���@�'&�`B��J��y��ɨI@�-����dv�� W�yrE_ ,!�Aa�HO���x[�e��y���Qd`4P����ea��y�9�� �g�6���b���yҢԸ_���,ٴ4*��LK��yB��_��x���TqB��O���yR���X�A�dҵA� g���yR��%)|r�1���n "i�����y�a �v*�PdD3Z,������y�lٕ;���j���"�
=�wB�3�y2ÙN���+E�0�\&��	�yb���K��H��FT	*!^-Pf���y�*ӻ2��p�/ε@�Ɂr'_�y2#�^��@{��@�pQp���y¬�6�(g��x-`Ur����y"�I2����DtA�Da� X��y"�K�
��͸g��j8a����y���mJD���'d��E�cd�<�y��
�~��q#T�U� ��ӯ[��y�B��_�ހ!S�$;�0��#`\��ymBQe,$���U 4��a �����y���X(�\�����(�,mB'o���yR�,a��]s���v�['��:�yBj�(V/�%0У�K�t�y
� *	)F��(d��p�A��J�@D{r"O4��j�8YC������c!��"O"��� �%�Ȫ��Z��q"O|5���h� ��#c&�a�"O��0��� `?J� "�ѷx�s%"O����_�@h��0W��N��\
V"O�<���Dtj�`Ɓ��Ai�"O�܁q'�.:p�a����~�ցk%"O����ܲ)01L�'y�p�Q"O�p�RKV`��9CP�Çn^|�R�"OF0�7#zmZ�,M���a�"O�Պ3��"�6�q��O�I�1z�"Or0xe�W9.�����xÈ��"OI���?I��4Ӵ	E3O����1"O�=҅
�2�"v�V�OuR`s$"O:1�n�T6ʘ���c,܈�"Ot��a�O�>�Vaj��WbO^�� "Oʌ� a���,��%W�����y��G'O���G�)o�}�!�D�y献Ae9IW�Ϸx��@rE��y�,ֿ+pT�p���p>��1�S7�y'�#/��rDjR�?j�������yR�ޒa�؅�H�!�L�����yRBM�Yh��{囂�z�B*�5�yR��(7����Q�g�~ J ��y"-�C|ؑK6m�P�ے&ت�yB���Kh��iH|�t�P���y��U�Ҙ�e�oG|4R����y2�D�K�T�r`��c̘�&)N��yBG��?�"M!'�כ[1X��e(��yR�_�f������M|6I#����y"솽H�	Q��J�7L6�Sa�\;�y"·8	uhذ0��\L��˻�y��فsL�1��G�O�ԁH��ũ�yr����;�ܝE|������yrϟ�wI���"�!(?P9��
=�y�+G	W^qѢ�P>�x��L^��y���9�,�[���+Y��l�R�'�yR�*E��y �h���h��]��y���>t��	��%�D�kO�y�Bۃ%2�a�-�6x�f�a���y�fA�YSȕ���r>�|Б�ݽ�yRO�FL����P�=>�A����y2�](Y���jA-�>@�i�G��ybJ�&���Q�֫=�F�'��y��D9%���x'���.�dAF�)�y�+�9e&��(�.��e����yr�6����hT9O�`W�е�y�
�>=�60����)%0Ijv	Q$�y"� Gת	Z�c�(v�I��g���y�F�)���@j"J,�{*Q��yҨ՗S)�=���6h�.�y�@��A���Aa1�����y��+f����.��4T��g_��Py���"E��SG��
��Ɏq�<�6f�%(��"Ň�0V��U��V�<9�[
#?�a�� �-$8֑ pHy�<�1Ϛ�1�-Vv'p��E�8D�L�U,��r6|iqa�ҁX�Z<��j*D�B%�C'-����"�	u�	�4'$D�X!���<	 p*���2Y��D��>D���G-��Q��U<ڸ� �:D�X�#�E�|��su�s�LP��9D�kwA!#�9"�ʰ7S�@��9D�� �xs��N�48b��p]`<:t��"O:��e��0��P�S�FJ�"O��Y���3]���E�3Z��j"Of y���&�t�A�?NC�@s��'��$K*&>a��`s���&�)r�!���(5!IX�����Ы@��O:�=���T��,I>	�1p��	��,j4"OD���@5$��<��ƀa�v4��"O���b̛����xbeܻ(3��c`"O�@q�Y�;�J�`Dװ�d �"O��)U%@9�ԊAC�9I��	�"OR �f� 5����:C�AA�"O��RӏG�z0(`�I<:0�	�@Q�h����i����/O�&�
\9�mC"9�C�ɧ\
�Mic	M� 0q�v̀Q�C�ɬxZ<�c�f���z����B�	!D�MYP`_>#&-����'I%��O���!LO��Y��}�<L���x�� 9�"O�tq�M3�.�:F͖�"����"O�� ����L�4H
0g7J��|2�'�I���:X	���5�^D^�Y�'o,x���:!��UJEj�����'���ۀ@9(5�
�BF���y�O�M���p��%��F����'�az�U����`ݟr4�-Y���yR���-R��7i�<B�`˟�y/�<Y��J�%
+a���aN-�y�L$}]�X $u��Rh��yB�	?C���G5O	�<��&�Py2�^(�����$zH �6�_t�<y�_�XUn	ib�����p�.�r�� �ɹdt���`�JpA�i��"J� ��jF��{DOY�G�����k�,ȆȓD��@�@�!�<��G�T�5`��ȓW�aÄ\�h�l��gkM�l��=��^Yʕ0��5�$A
1��^?��ȓP�@�f���wHdb5�%>���Dm�HW�˛UeL�"Å %5�� ��W4.�c��W�<�.$	�&��U�$i�ȓA�u��������AK�+ ��'��D{��Tcd��	��\1�.�t����y�J��`��6Pp�հ�y��R�e1HHc���-�,lY`-�y��K�#}�!d��<<�a4m��y"��+ ���!p����=ғb�	�y��B�g �Bq��'c$���X$�y�U	H�,i��Fºc!T�jC��<A�����P���Lد$!�8���3LoV�OL�=�}2�-ʬ~D�R�� Kl�$�I��<��E�\_`%�'l,���D�<�W�ZJ�����#CyT�zd|�<Y��O'c� R�lãf�\\��Ba�<	�͚Y�Pӣ"*e�tC���G��4�<�D"��Xʬ�S�R�$����	A��T���OP�Tz���"K�-��!�%��q����5�b�� DD1��i7MR�E]:\�R"O�����_�!N(@f�PQ�t�R�"OH�QB�6zϔE�#i[�d�"O�а!�yM�p��փo��8��"O�+�6'Hā��"O{��C"O��a��5Zr�M����ٸ)��"O.�(TeW?���'�4��1��Io>���2$�f�V%K=kZ�ukSG7D����G�$.��sɈ!sU�e��:D�� �]��	�e��b�@ǻs���:�"OF�ʧ�ٿf�x��V�	
f�"ݠ%"O�Qi�H�@���)!���2�L��џ|��'[�h E�=G~��*� �BT��'�&PcD*�wB�I����w0��ڎ��7�X��j�_�6�I�!R�5~@P�A"O��	�`�4%?t1"�n	r�L1�p"O�U��D]�e���&C # �����"O�%;�`O??&ı�g��`M�I�B"O^���ʇ��KS�\%��id"O���Ai�z�8s�d��\�"O��@�
)U��
*@���t��U�O!ʵZ�`QR�n���!�� �.O���7f�^*�C����T�1 �f�!��B]+��Krt�ݪE�!�d �t���@ /��!���I� �!�d6��8�]�3�@#�K�XG!�D�M/�u9d�V�O��!��Y#�!��-v�$u$'I��E�5	O%n��'�ўb?�X�b�M�>L��"ִxV��g\����I3I� ;�9o,#V�pfC�+&WȠ0��PL R�r&�8
�C�ɉ^!h�P�M ADؠ�BP�C��B�ɬ%n�9���>2X�q�N	"RB�I�1�Z̢��H�mlTC�
�&\ B�	�_$P u��>`H rDG��bB�ɂV��q�2�F"6���"�)��C�ɰ �j@�	�	7��YHr�9$�`B�	!S��6����&A�p�@�m�2�=��'@����l�zL9�E�B;`���FR�����@-F�tٱ4�V<�܆�wv��WJ�4�����̺Z��0�ȓW��TJ�		�JSd��R�R���ȓgE�x�dX a��-��P8$��=�ȓ~���aea�������1^��ȓQ'$�kҨ0(rd�ThZ����ȓ����1������Ŧ��ȇ�B+�1ah s�b�H�`ӭPJb��?��,��q��B!N�@x�ç/Q���ȓX���I�2���X�&Zeȇ�;9��R�C�@�Tp��g�b��|�"�)D�J�)^,q)����`B䉗nY�8i�+ɋ7�
a�C�{�|C��/kG*�� h�B���:nZ@C�	=*���4iy ��	PHӍk �O���D<�z�9�+\�-A��q�(�ў���	�z��ar�ǄS~���smJ�\�8C�	h\ Ku(W�L�H�����.�C䉘N����[�[y,�HrK��r�C䉲W�ٕ���u1@d1�(� x�B�I�`�CV�V�6X� �7D�D�zB�ɇ��-+��?bM� �Xq@`5j���'��`o�<�4�rŤ���ۈB�)�df�Me@��c�'"������'��'+��'9
�0:`�D=���!>!��V�g`0#���-�,��F�9-]!�$�*@�nUa�fX#͌�x�&�%!�D�7������1`���d <!�d4e�4�R+ʕP�1�6���)!�d�
ir�����˙&BdMS���)K�'bў�>��N�z�`4�2"�x):��A�Ic�O�"H��K�	70����CF���'rN��a*FS���؆dX�'��U�g�A&Z�x��7c�<������ �X�so�sd�)%@$i8�X��'����0����#ԉv��x�u�X�]�!򤋞y��A6J�)�P!`�C�1em!��Y���#c�_�TH��o�<�5O�����=,�Z��v�xq�"O���@V�J/��1+�>�TB!"O,�!�
π|�.� Ӓd�X���"O��ʤ뜬UT���cE�N�`I���'�1O��qBӯ(�՚XY&����ៀ�'�ɧ��N�"�
��H���w
��/��-<D��١� ?�����f�	�G�44����C^�"o� �'�R� 3��b�<�#]�����_Y��RP��Z�<9��1J.�q��"��C!z�#a�*D�|����7 9���b��40���1eg)��䓹?�ʟ������P���@&�f1���S�XG{��i�U�Ddc�T�j�D�b����*D!�D�4��JcG�..i� ��34!��D�� aAʖ�(V�K�CB�9�!�DQ� F�$�c
�5
6��S�@6O�!��V�]�����Ʋ7�I1��#!��P`a��+N
tVոC@U��O(�=ͧ�y2����%�T��v�`C�>�y�F7X�Y"E�K�$��!�n��yR�@�~.���WGK3;�X�+�l��y�jte�)PBfV(=b�8���y򩆻X�|5c���D��A�����y�/��.Y,YX��֍;��Qe��y�*V�w 4(y��I:,�`�����䓫hOq��i�ݰX��e��4M���J�"O*i��;��u8oH���T�"Od巤Q�@� vhbY1���y�*Y�� J�P�A�ZX��gX�yB����.P��$��9�d����y"�_T��qjB�9D�0�cT��1�y��Y�`
Z0�/�Xi�Ç���?a���S�q|��� q�ȴ�Ӫ �ގ&�Ԇ�+�ruӢ�_�"���D5
�C䉺)#ެ)���k��Y���fǔB�IV5P��A�Q���l�O��.�lB䉎u�2YH�H��QO��ye �r@B䉣xك�i�"������(qu(B䉃0�z�� �,n�	��\�p^�C�	*�#"'M#���\Y���$�O�����/^Ǽ����Ӹ	7� �L��'�a|R��	ejH !Ő�n�L	�Wl�=�y��S(��ժ�!�h�i����y
�lƎ<�bC��K�bQ�v��,�y�!A�CJ��%�X
lc�eI
�y���c�X���/B�܁�ؙ�yR�	(g�[g�.@��:�/\��y�-R.K�,h����<KF���y�*�Og�����-J�q�&l�y�D�(;��ȃ��Tp�!��H��y�˞%�bH(�`��`B�І��yRn�2Ud�s'�'�Xd���G�y�f��F=5�
߯/D��6Jլ�y§ 3	$v�!�G�)�,щᇇ�y�*�w:]0gG	� ��Õk���䓓0>1sJLL�v�[ �H�5Z�|JG�WC�<y��B�6PJcn�[���1�o�t�<��d�a@j]�C
H:usNHie��n�<���K{[ެАM��=x�t����g�<�@.�$�|kB�[P/�`ąN�<� n�Y��)#W��B0�Έ52��j�"O����FO��8b��D��h!U����	��:�BGm�@̘9��C��B�.-D��mL��0�b�'Z�bB䉪(pHt�C+��,��b�/q�B�I�JlhUXg#H4x�h��L�=!ĢB�	���%�C%]��e3�/	��B�IV�,H��aܖ8c$lK�ύ<BB�	zd0Д�Վwd��'�=��O ��č	^L9ka��=T�ft���	U�!���n�2,�@�ߵ;��H���u'!��ܡe���u(I� ��Qo!�3:4m"fm�̨�n�)�!�	-4��=a��s��ô$n!�� 	�<rB�@�:�\q�3+�!�D���ӀfT�j5�P�PI��[�!�dӪ ۴�"7�E�! �=�u��	�!��C�lq��A�
e*��� +�!��Ty-�A�M_f�b�c+�5"�!�䆞>h$��ʛ=��b���S�!�/ڎ�r)�&4{h�[���3��O���$
�Np0�a�@�"�E�D�!���J�P�K�zjT�JS<
!�$�Y�U� Ύ�+WĻɍ1H!�0��}`U�Y'tFRp'��-�!�$o�1�'�ەB�r��匮f
I��R�jT����3'�<t��S�eǮ4��0ղ��Ei�.P�d�0l�� t2I�ȓ�b-����	"��f*F�O.XՇȓ
n�}��C�n�D�QL�ȓ>��4�K�b'��3D$!5���V�.�� ^:O�x�Uc�:����8[n����0{DN���0mb�Ԇ�:��h� W�.�,+rH�ȓ�Rl�L�H^���E��������IC4!
�,q�Θ�	��ȓl�z`��%�S�m�Fn�#�nهȓ)����jtN|=�aUV�4u�ȓS��q��!��JP��@)ev��ȓ��h��K�����j˧=��цȓbr�e�f�C�g0 �F�P#]k�U��m)X���;QpR�xª�E�q�ȓD�M�V,�C���4m�'�bx�ȓ(�.��͐�Sd�u�I�F�*-�ȓR{�t�sa�V�����"�h��iԒ`[����h�!Jǁ�G�����G=B���,�y_������Qz����>i��LFS|���+��_��m��,��A���C�/�QG)��@����t�������`iH>'!�9��ʞ��툤�/D�H�6��*�<EH0�����UA'�-D�P1�HJ(Y$Q���D����CQD,D��B�� �`�X$��KD�w�iJ��*D�,J�#H.���J��Td�Q�s)D��"Ro��A�6kxȪ1R`&�O�����UѲ@�C�me�yhp/Z�Z�d4ړ��OD-jb��L�H��+�,%�*��"O `���&�N���B!Y�m	�"OД`�(�<z�zh�ǡ�zS�"O�1�$Ŋ&�1� V�8t"OʝJ��CJ��Ю&<�B�Z�"O�۰aw�ꔘ��	���-I"O@�
!n�4ͺ���ܘ�:M�#�'��'
ў�Oļ�)ŀ����M�S
�b��� �#sH�1�H]�w�#�9�B"OT0f��J����ܡe�""O���7	�� �  ��)��q"O��׃@55�QǮ��Y��Y8�"O|-C���";Ă�����R���'���ߡ��9����,J/N5���7]�|��)�d�T���8�	_�1�ޓ�y"㑼^.@pB��L���� #����'9ў�Oufm���\�͋��UU��
�'TJU0��ޒ{����.��U#X��
�'{:�� BC�!��KS
?v2�
�'ܤ����g��� 4X�/{�� 
�'k4\���1�x�dAǶ[���Í�'0ax���d2��x��I�Z�#H��yB,�P�P�ޜEX���a*Ѫ���hOq����w��i!p�YÖm[�"O��2Ĕ*���0q!���8
�"O|}���*{G��Q�{�xY�2"O@�	�@�<\`*0H��k���H�"O�	Ѓ*
���RAG�[��md�'�ў"~�1EƼ}��є$�#9�z�yG�	���=يy��.<C�D�k
�C���2tό2�y�X�*�ȥMT�)�6��>�y��Ģe�>Չ�& !��,x�����y��9L�J�� �Y1����y�(�����F�X=JB�A5�y��*[�!��y$�����?����S�v{ٻ�f�)Wa$�A@[�j@2�ȓH�������<��	��M�.�=��W�l��Bb�7�V��I�*x촄� �2\��枎8_b�����L����ȓ#��49���?�`��\Y�^ԇ�.1�0� �T+�2%�0`�T���	��)�a��͜P�A�X��8�?��.\�y��K�0�q�ë�o"  �ȓrR��c�� 9�HP%�`e���rz��1#DVzt�!ůs��Y�ȓ���jS`�i �`$)���F��+�\�#bK�(R@h��F)�X�ȓt�H��9&Ʃc4G��cptȆ�|y�Ԛ�L�8'h�SӅK%%`
y$���'��>��4:�N)Z�����c�O<��B�ɌY&ب���� �.��-F�B���x�r�`�+���:�lZ2hfB�	�,	�l;� _!=��`3e��U�C��:Ԯ���M�Pv�D�fA��ftC��<2�b=S�7����a �~\C��^a�����܂��[B�a{ C�I�od���"�!xt����H�HB䉵<��mIsg%+X�v�m(� D{J?���	��S�:\�U.MX,���H D��QFL�6Up�i7�xX�=�5�1D��ca�U6E!��aپ��A1D�@���y(���0%( ��q5�0D�P�Si�>Q2�j֋UlxQ��d�<�H>�
�'L��h��P�[Ȁ��Օkv�A��x�N�Q�o�Ojv!ڠ*�_N�?���~:d։%l�`��+T�"�ӥ��d�<�s$L�L�h�'�&aT� i�^�<)��M�#����gG�Ei`X�D�N�<)�nG'f�(� Cl��[%\r�'�@�<YR%���C��:���A5F�ПhE{��IY1K!��X��"em4����H��8B�I�N���AE��u�8��%�G}6^�HE{J?� ñk�<S6h`�GFd�1�"O�С�lL?U���b!�&W3�@�D"O6!�w�є^�4�Bd�W l�I�"O��5�K�%�T�$�ڷD��b�"O�����R�a���_2G�^5��$�OF����-�=*5��*J�`ҡi�=r�b0O�EY��х9��ě2ٜ9�`��"O��jj�	2f�;bwD�B�"O�,q��
?�8mP K/Xh��1"O`�Zf�D��ur��4FI0��C"OzH��'m�P���P�YLxh�"O�$볈J�~�v\7h�.,�͑f�|�Im~�e
�`��T�c �8�xU�p����xB��V�zh�B�SV��훳 N�7I!�d(J����!Z�c�t%.d����"O8��@S�p0�Q��H�Q���"O�x3qH�55=\�S�m�4�|]��"Ou�$ͯ��eyb�d�l�1"O&�4�		1�~}�NN��\6�'w�'!�)�L~'��0��ɥ�@�
&�	� F��y"�ߧIIZ���0f� aˆ�y�����Q�S)(萣�;�y�+ЍG�*-q�l�R�XM���M��yb��:T
5�$�C�0������y�)֔P���e'G�,�Ѷ�W�y�V;�h��7D+`�|����D,�O�Y��fQ5<ײ,s&%ОO�V$�0"O�0�_�g��\��M<h��`�"O.��D�,�l��"J@���$��|2��5h6az�CPԆ��Aa�]�9����y�E��`q`�Yi�)�D��Q$��y���9I^��r��3�Hz� X<�y�*�>-���E��9�>���Ɲ��y�E~}�Cě�3�.C F��yN��.^b��}D^Pq����y"�\&(mQ��1w<uI/��?����D�<a����5e�Ԩ��-�PSE��!�T({��b�̻~��ј�,��!򄛑F�9t-�##MT����!��K��er�(��a�б�rO[�e�!��-)XP�0��E)�ʍ�r.�<C!��
	Z=�� ޠA5��hӔ^���M��4���̰>A�����"�,�P/#D���G �Y�c������ #D�8��`�&>-����e̮>�p��$D�,a��(���y��ԣ$�D��&%D�@{�F@2Bh}	�n�3�M�QE=D�h��J�?p8������ "�%H'�?4� �2oI:o���h��'H~٪���H�'ya|��ߊ&wf��Ӂ�$q���Co��y�g��R��H� @��i���*��3�y���sfz� ���a����(C �y�%6g����Oٖ[ ԼRbJܦ�ybM���B�jG���V+�I�Q��yR�߮+�,�"L�G��:��Ż�yRkOi��0���̀Ft��i��+�y�̓�%+ڬ
����f�iY7H��yRnKd� �3F��¡�f.���y��h�.]��u3p=�jψ�y"��E�%s�L�n'�!+�
�yr	�8��܃!�	:��p&��y�j��-n�����V�8z�x�	�y�_L*��҈�5�@�Z���1��$%�O��d�-8�Ĭ8&�6"U��9�"O� dDzI|�|h��\	5���b�"O(QI��!&�e�FG�7f�<rb"O��C.�%3z� �GJ{�=�""O��+����_�ZV�]$U̸�p��S>���A�; 8�a�G9�d�G�5�O��uP8��`¯>�j@�SiH.W��D+�������9L��U��"�6�a�8D��r��0����w��U�t�"��4D��6��.��Y�c�B���$ D��:�ڲPM�؊`c	
,ތ�uh8D��aө�#9Y�4l��]��)�Aj�<���#}*�(�(\�w숵0w�^h�<��U��} �ϝ>2F���f�IX���OҐ�`�E�b<��'$'9fm����dЬ'?�u���H��>��'V�^>�IJ��\�'%W)x��&ޠV�@`�J2D� y@,ʄ(�PbdJ�ޤ}�A�+D�X{욇37�t���_H�\PGf>D�����W� ��ز���;cƸW�8D�L"S͆-[: "�J�Z����7B�OT�=E�dC��'�$�U)�kj(�Lg�!��"gҜH���̆&Wb�
H�*�!��:Zn�I��O$%�\���� �!�DV:wJn9ڰ0 ��$b@�~�!�D	�'Z��a�ă%Ŏر���pzўL���+q�6h	���A��+�H,ZO�B�	�\Ppəu��7p��e�:R����$�S�O��`��N�<JƸ�!E�M�7�C��Wl�x��l�@�j4	��{���ȓc��1��Ȁ�!�Zy��*�;>��ȓXġ#���l*%J��j�����^~�s�@��y��m��-N6L���ȓ`���cI8\0��p�Ҷ%L*��ȓ2��`͝ 0u��:F�I�&Z4E{2�'�$z$H�1J"@�jE7)t$�����y�C�gH��OE�|X
R����D3�Ov��
ܡq��K�/V�e86"Ot1���ЎW-0�0W�WI�lB�"O�хJ�/.��6G�&b6`���IE>)��3@T\RA�ֳs�l����3D�0K�%ʍW�8W�S�q{�$	�
�<���Ӣ�^�#����5���h.B��D0?���؏x��\�%�7d�v08�kRAy��'�����2dI�&�١+#:1 	�'����)���͠v�L�o��!��'3VhxC*�m+��;eoʋZ����
�'1r���n��eQe\�=%V��
�'j��Y�T�;�p�PR!��O�%����hO?�p�.��V�rVJ�
�}�a�Hx�<I�̌A���Ǌ ��`ht&i�<���.m&�a��+��/�%ȷ��d�<1�(�
5"2�P���QCRd�2�K�<��ήr~h�"�T�]���#KI�<95��b;��C"��Z���І��]�<��B5c�N�хi.�\�e�@y�)�'M989���K�p�j�R&EXC4�ɇȓhfh�gg����ӈ>����_x�<9��ͷ+�V8�CL`�~ YŎ�u�<Ѱ*o��Qr+'|�<�`��BX�<�%�()d�&.81Zd��H�J�<Y��5]�D1KF2v�()B�L�<�	�*�5�a�	��9d[J�<!���
�	+�.��L�0��HyB�'��c��x�0)�@=�(���� |a*BO݆�\��ր541�"O�8�gL�	�����.����"O�c�� -�V�QɄ�.����R�'T�	n�)�=qBΆ�?ST �񄁟��*�	�l�<�P�\��`�A�8��H3�g�<�Q-O�d�>����ـ 0h����b�	I��`P	�x|M�n��!�tp	$D���4E �b;�=愁�;&�K��"D�8+& %r(X�_�B��SaE6D��
��X�d��v+�gG��P�A�<��2��m�Ba?8jh@ C�KL�|ՇȓS�j��g퓃f'*��؏n��݅�i�`�6",(��˧hY��r)&�0�'��>��*V	�!��B^�^�е0�k �e*2B�I 6�Y�� �̮i�d����yBȌ�d�B�&�dT�@Y����y"��ow��mG�X$��;�G���>a�O� Di�=zԠ,c�ȅ�^:��[ "Opܰ7-�7�����b�h�%ZG�|r�'�az"� �Ӡ$���(4І`_+�䓑?��D1?A�f�D�16bPcy e�wM^�<���Z+�� ��?i���@�`�<�eo6u }B�"�����@�OV�<��/�vb��Yr"Q<b�HŰ" Sx���'�dK�P�8 ӆ��$ڨ]1���hO?�	�.���P�S�W�h4�}�bdU\�'�ax��ޜ\��x�M!-�t(��ǜ�䓉��3�SJP���Oʠ�JW G
1)�b�<!o��4{���M�M�^�q�[g�<�A䜬1�)�ɓGݠ%H2( J�<1�/F�
�p���ʔz�(У�͆D��x�<�S���@	��"]�uk�˟p��[�S�4�'��	A$��$�T�K����CY�1�LB�Ʌq�8�����~���e���L�B䉅%��@y�k G��Z��<\�C�ɪfÆ]QT�&<?��s/ӫahC�Q�v�;�e.V����!�mVC�I�qcl��@���C��1�N�'(cLC��7��`�H�8}�W�̲C�ɏq�xИ��ԁR� Ŋ�x���2�S�O<����ތf���ZW蚶gq�d"OV=�U�V ����Z�nWU��"OD��:��yq�KE�8�H��"OB�(�cB
FJH�3%��o��T�S�'��Ez�٢F��ly�:�jY	a�L<��'H~ɩ��I L�h��dĒ�^�-(�'����	��7=YYtcί |dK+O����S�L�@�����P��OC��P �h*D� -��OUd�YUN)3.�ܹEm#D��%�]�m p���*@�.m��.D�0+vN�)���ˇ�4h��P��84��	�>Xr�ҐG
�Z.�t�Y�<�"��:X16H�ON�_������K�u���O�\"ыD�YI���C��b]	�'��"�N�K�R|�Th���8X��d(ړ�y�NY'_�"]����q�h�8�h0�y"J�+e���:� J~dp���ֲ�yB"۶"��HA� �p� �"����>�)Ozd��G��e�-�ʖ��C�=D���!J]
tT�T`��att�" �ON��!�)�'	�R�`q���t�T
E���Ѐ�'k"Y��o�$���)�l����$%��.���k�X	J&"p[��Z�O|�<�炂�56�����ڜZK��Y�B
u�<� ���	�&l�2YB�U\�2�"O���cD�2)i6����&gJԨ"O6|�F�x���P�M-N�6C�"O2����
���⠁�bp�X�6"O�DȤg���Ȋ���;G`��7�|��)�ӄ'�PU�ˍmd��˷�H>�(B��,yθ�ɖ C�L���ʀG�/R�B��7�Z,�� ]!�켺�H0��C�I�	�Rp��NT�|�h	c�:]r�C�I%\��y�"~�8�@�dv��B�ɡ_ hA4��`�J��QHS��B�ɶIT��/�o�>5� B v�<B�	�Hd��l��mx8�IF@´B�,k4���� (=�T��,Q�0C�	�AB���T┦#$4,2�nY8#�0C�I�_�}��"Z$7"�ZtN�e�C�I.8;�k�)L�)�K �n��C�ɅLX���7�[�G�|y��ž|�!�䙴z���2o��߶��vD_�m!�M�;��(Q�/:���_ �!�Dֻ�R���
[ͼ%R����!��ȓY	20��@>0^"���,�#F�!�ײ�x�B�8cpvh�lTG�!�D � �"f�~*��j�!�d@�`��BT�З#FP�2)�(�!���MP�����LKx�`��!�!�NJ�0����$�n�i#���`!�X�<9�h$�˶��R�˚��!�ĕ��45RI�Gޢ`q�
�&�!�$�X�8ڒo`+��*
9B�!�H�o��
�eC3(��HY��!��������+^*�!2���-s!�Dډu�Q1���4%K�N��!��u丼�$�ؐo�h��C�xm!򤈪N�j쫇��2~>�j�@�8�!�ό~~%��ס-f�e�P%�=@�!�d�(S/���T�XIv։�q	p�!�PA���5�,V^�-�d(�.Z�!��G��P�t�L�JK�5H�5<�!���d�w�}W�TA�aX
u�!��,���
�#F/g@�Q:6�_G!�$W��"��A-��s���;G�!�*���(7熃,r�<QnR:�!�WY�����N�8h|\գ7�>YG!��	Ħ��@�[���+���Y!�$��!
`4RS!��[B�����X�!��u,��jǽM���"f팅#�!�d	^6�<�a�@�`�;s�(+�!��
+Μ�"�_-8V����	�(�!�$C7*XZ�e��-	p	�эݡk|!�$��@��j
�,;0-Jti!�M�x���փ$|���=|!�dB�4�t�@)�He��&Z�6�!��֭\hT�%���Y�-Q�nʩ5�!�$ϳ]
�Z�з�.���U�!�D�;ef�����$8d J05+!�D�+��}1� �'II��CB�o�!�D��<٪ �E� 2\H��n�iD!�d@3��I�^j�]"���Z@!�`3�H#0�؎�̢�FK
yhB�I�&e��
�.�H��K�ƅt�~B��C�f�G,q�à
DX[�B�,8{*P�R$��M0�e�r+xB�	�z�$�A�K�F�}��e['EVB�)� N���H�:��h������"O��)�-���6�Hg��	n��T�P"O�9A�HN
�u3��ݬD¤	b""OTA�@��-hb:���K�X����B"O��qG��:�R�h��b��	�R"O0�`C�؛*��1�8V�,�W"O<\� d����B$��zF��a�"O�]�f��S�l�9�A-Hu95"O��褢�.�(���F�Li�"OBura']4���=��M��"O�f,X�6�Blr��P�G�|-��"O lYW��4� ��|Ժ�ѧ"O4����o62�Sd���M t"O�5����5�@�)qi���~|�D"OL}A�n�EHƅ2E�F.*��u�"O8$�Ƥ�-���ɶg5C� ��"O$�82'�.L x@iB ��Q�"O���g���BUʂ(ƅ_����"O��RKe�`乲�Lgj��z�"ON�����2X��+�	E<Upp�"O�q��`��}�tW�qq�ѹ"O&I{����_��-��G͠jEb�	�"O����I!~�1w�V
�"P"O����,�5�Fn�]E"O��q��>i�*�X�o:]:n�K�"O���2�ڤ+�}y�i�*R�*�"O�� P��e�(�JG4�@=��"O�S��̰ Fh*R'^<E���E"O�}�ǯ�}�fb&a� ���2"O$�9�kR�0�Z��Q�_M�X�@U"O�4��/7GT=����`}(�c�"O�(��o�A��M%KӶ�y�"O��'�� ���Gɱ%s���"O½ࢊB�/�`F^�I�.�!�"O:���AڢP 9:�NC/6���@c"O�0�ͅ�-��(	�-�U%��1�"O���5.�H1�����QD"O ��EK?=�&Uj#�G|���Sa"O�� $8E̪����4�9�"O8�)u㊕y��ࣰ�I��.�D"O8]@�݌Oa�ͪ���A�>�K�"O*����L�?��1&K�q���`�"OR�@�Ӳ+�0)`s]�!�"O*؃֚S�U���?I�$�s%"O���7 D)9"�|زe��|�&ك"O��bC$T.XQ ��&d���}�6"O��b�e�2wn~lxg"5z�t�h�"OIs��A(%��Q5�N3o��c"OX�AS���r�lXC�NX&H6"OF0D��-�����O����T"O@���a�lo&(�����x��&"O6h�H;���tm�R����"O�Ɇ(ӳ>���DmUf�~���"O��FC݆L�ݘՉ�K:(��"O*�3��H�*j�Z�Iӿq�D��"O�4�5�ʖ\.*I)p�ٰ��L�"OL�їG�F;�Z���\8��"Oԁ����$�<��HF!t�1W"O�1�"R eR8���۠I4���"OB)��ʨ[�0��Nߞn���qP"Oα#��
|���3�-ܢa�XrP"O¼��kP,�-��ٖ!h�BR"Odts!�R���,Ʌ�� ��i""Ot���>j�^���U��)��"O� ��hǄG�`	⣣��Q\�{@"OT��K:����@�ĳ/C��"5"O:��i��"ul�ː��+p B�"O0���K���1Unȭ4i��"O�K&&��+���آ8 -��Xs"O(����A
9{Z�B�@�r yI�"Oh�[�Z[Bp!a(�?C-4!�"OzI�!��8��+3.˱:�H�S`"O"-	��.�* ��N�n�2�"O��E��?��T�SȀ�,�`"O��qCg�-���`�F�VL�"O0ui`�T��d�J���+�☰"O|�	E��"H�:P��'
?k��9��"O0��! �,bx���f�>�9�P"O��:sOQ���$V"s�D�"O�)*�$_�2 $yQC.����"O�	�v)؆r6��C�R�u�X��"O^��S�β%p�:Go
)$w�s!"OF����:@��1�R��]ї"O*7�8(l���En֋oΝ &�#D�4��gΨH��� �T%>< �Y��#D�8a&F�7d�D�4+��'���5�4D���#*�#qo���H�3@��x�3D�̹�)7<�`,�h64�|aiw�1D���I� %���ĤslAS��/D�\��(̄I��I#�n�wN����-D�4	���c'�#aFB�f�$���,D��Qr�M)�F�7f߸$;�X��+D��GJ�"%ZDx�E$��rA�Љ�e(D���SF�D".ɰ�D�l܊5��� D��O>,�ƝXC��:�x���*D��pCLS�hz%��I�mV<ͣE�<D������	��b�/�4}��<D��37ɂ�HT�� T:��%���8D����׍Y\�m��hΚ8��9P%h8D��s�(��A��p��Acg6D�d��
�����5&��5
:D���w�͙��I�a	��t�U�E�;D��@ԫ->���7'�qb�IZ�%'D��CǏھ!�(i��ɢ/�}:/&D�\��ꕝI_(�*�j��#@VB䉏D���rFK�$��90ϔ�+�B�	�J���� `�	'P�4j��H�C�I%K~��F��:d��G�Y3�B�	'X���m*A��j�|C�I�#q$UZb�W�}&�1	�&��<ZC�	�ob2Px�خv�5���E`�C�I�E.p�yV��&_h��Y��B��4C�I�@�j��\�FN���_�r3C�I�ަ��7�Zl�t�Ŝ1F��B�	�\X6|`��N$Z�dز ��K�B�.h�4:��Z�{�zl�E�[���B�V졻�O 4�HT�b��N��B䉔�@0����7M�:t�w�V�MڄB䉬��f!�Be�?y)L�Aq*O�͚O�!�qisD|���"O��Pa�Q�����U.ظj�A��"O� �� �/EҰ�%C߄J�!�!"OJ��(ٕSR�5ءaF��h�"OVY�b�ϡ}�n���@�$��(�"O�%�Ң��\��p�!7Q�<��r"Ot�h�ܥA�H���;q �8�D"Ohĩ$"�3��!�C����'�qO��/C&"�X�rI��1��A("O�  �(���m����2���`��'�L��'�b�٥(�A�����C5�=Y�'�9�5O.���H�9�|*��d'�S�Dʓ�]\&d����A��h���y�#S��9�TZp�� �T�/q�<���O�(�-Oe������n�H���I ����!�[3Q9�Ţ0�׌�b��Y�hc
�1�2�4��=[��2@�)+y����Ñ��'}}�'|��#H$T]��S����z���H�'�&-�\��؋&q�Ɓ��OTY��O(�	j�Ӻ;�O��36+�3I�h�b戅�3_l�[�'��U�s���hy�!x2œ!F������'�ґ|"P����ʑ!G0|�D
U�SaRh�cVh�<���E3'�$){��&~��x�b�Za�<� �&�,����׼cK\Ը��Z[�<��Ƃj7�T2���yl� �,�Y�<i�E¥BP��Q��8I����eY�<)"�ҰV�2u���\</�B���S�<aL�%����9i��;ui�P�<�f�dl�Q�v�̭8�:a�$!�$�	O�$aA���T����)��k�!�DK`I� o]�h�V�2!�!��˲=�R��Gtԅ�s�\�j/D8��hO?M��9N�$�H�BѧMڢ��U�#D�p	�Ƕj�� �φk��$�!b7D�D
�gH-�y$���G2����*D��e$Եv0V���@C�sh�ʷI)D��Ĥ[�3��(�fj�L�d$�s%%D�p�  ��sž���6M�b�r��5D�H�s�*�`*��b  �))4D��ҐD؟+|���ߞ=�
 Ò�p�E{�����pB� E�:�Ą%-!�D}���c�ϥ9��y��IݪW!��(h��d�3�&��&��N!�d�6jB>�$�&j���0���n�!���g
�51���,�rf��X�!� ���ۦ�L(x(ٛ �ΏC�!�Ԕ|�i�筇h�����,^�	s��0<�I_ʺ1Pd%	�@
��$k�<�% �/\ph�3G�H�U�0R�e
릑���/�T�d�J��N�Ť=cBiF#C�ZP��6�q��VP��G&էg�D�'��~�#w��IF��^~�p��Y��d5�S�O,�A�BG n�&��B�L�a��Ep�'��+�ߓ<6�|	����T5����>Y��	��t|p��PdY>Ti�V*�	F�!�&�>,��gڟ�Kѣ:��p�ݴ���1���O�@A#��a� !��Ȋ2�nM�'F$ы���1�����gH-0A�xS�'�д��	
��uA�`ԛ'�LJN>����~��tR	�0,U(H����ȕ�y;<\�� �K�j����RKD��R��<a�O�ܣϓp��@gٖ���9��$Yݴ��=t��ifjݝ_"�-H�	�yr�Gx"�'���X���1���ׂ!H��4���d>��UeC-Iش8O^3	�(�0Pa6}b�'SP�zg��G���ж�M�C�f�9��?	��:1�ѡp��5ͺ�Q�g��k�!�_�z���j�$�@`�4p6�N�+�ٟ�'��;�Oq�
$z�H�]��dCr$P�M��=A�"O����♎>��<k&�0,��,;"��3LO��x�
�+I}H�Sdl�(%l�q��"OL�l@�Q�dЧ�U�`ܩ�g]���I�G��ʁ���fL(�Jː*��C�)� vh���ùl�����Yk��	tX��Y��[7D(�(&m-YV8��.��1�O�� -a��� qo�; V)0! $�\�f�E�^��p��Q�H�Kc&�z��D�?�e$څ|^x�K#��2�4ъ��L�<�#�U;]l��@E�,Z�D4Z��dΓ�M�O>E���d���B��H�&�2���J��'�H��?�͟��J8jYP�dj2
M��֞~���'��&�'���3k�u�q
�͉���a��>�e*�>�N|n�?'v�,Sp�)!�U�ƍ��l����ēMj�H���؀"N@@(�nLE���Ml��u�=q��T?��r��.�
|�&g�g7�A�:�c6�I��P�p�圜`��xT����84�x��)�S�9�ؙb���-�`���	��b@>O���۴�ا�O���t��0e�`�+�23+�y�O����5**PK����Z8�D~�Gx2-�'�?��w���d�ЀII�58�Bʇ:��ȓ�6�8����+�@D���T�����p��>	��3�f�r��AM�Q9D$����
���ȓj�Z�q3�
�;fE�p��_	�@��O���G�*�(Hb�/Z��O��@u�u!(�21��/����Pe3D�L�� ʗs��yu	��P"��#0D����P��8p`j��a��� /D�dY���Zc��` �]&t���XAM+��6�SܧVJq13��};�B��5A\Xԇ�A�&	��d
��J�ふ�(�Gzr��d�O-��i"���x��2�@83�4��'2F1÷Q�h�x��B�G��4ճ
�':*��'��,}z�;�A]�t�މ�	�'��U�T-S�$�z��T�6Mq��'�p��K;3�Vp�қ@�^5��'����%�ʢb*�<�D�)@�f�8�'ˮ��D��i�z923 �iD�Q�O���$߉j�X���l��&�.�Ԡ,�y$��asCnJ57��Yc!��~R�)�'n:T�b�J"�� S�ɫb�BL��ID�k����D�Eh	�eXe�$(\(�ȓF���c�<A7X��`�Y�"�����hO���`I�/ԨxS��������T��DR���'�(��`�پJ��5#�;6 8��'� �C�Tٜ}:E�92.`x�'�*��1ڬW߆0����[�s�'��,	�)��p�왻������0>�N>!WG!�H�3��	W�F�zg��<�'�Ă�-��؆C�8��S�Oq}g?��(�9$P�-4��R�S/0�����"OP����L�o�D�������'��<�	�O�8{��H�cG���Fįw���/LO"�`�ׄJ�[����&�@px�� ��>1��-�b��$'��3��C�&T�J����8b�H���$(=��ښm�TXb"O���QMX)?�`�6nC�U�ݐ���d�ڃ��D�$@q�%Ŏ8`�Ҍ�S�<�6`�F�8A�_�$H�-�t��<Q���6{�Ѣ��
2R~xx6NO'��c��D{����P"a<8���?�$������y¯�+a�� V���r�|�"&���y��/qGF��'X:w���!gk�%�y҂�q~���T�E^F8;�N[�yr  ���3�IF�T��X٦ ���y�!H��#*�Gk�A��V�yr+45P��"@L�.D201)5g��y�̖�r��a����>%"T(J�7�y
� ���#�uZT�ħߡQ�����"Ox]9�D��b�C�ĝ-F���""O�Ȉ�,���1���N4Xa6"O���dl?��(d�9�1H!"Ot�S�Q�:��eH1�P�U���"O��y!(A�4����0�-\�r��"O�����k��P��B��zG"O^�S KF�Uw��KDIQ�?� Y"O���G0�[Ղ^��ڰp1"O:��ЯJ�j�`�Ȅ� :��՛�"O2e*@�B�\ܰK<�fl�S"O�]��!W�/�0��-ʭ0��<�"OACU�^m�Hs$���1���"O���U
Ĳ+H$A!�ю� "O�e�"���DIpӬ��VÎ��u"O�]��'�:F�nX)�+P�nI�"O$r���j��݊�)|����"O����:��H�$�)cy� '"O�b��E/4%̽�6I5p
�"O���Dbϧtd\*���5@���"OB�K���?A4ؐtȮh*�At"O�$��˩Gz&�j���v� "O.%ఊ��l�\���j!�i'"O
�§�˘24v,�hF�r�us�"OD`�
�z�`�f�C�~�xV"O���'f�.�0hӲ�&O����"O��6���e� R�-=��B0�J�<��
H:`�h�@�pN���G�MC�<��@N�?C�$�I� 3Zt�v�XZ�<�#D�>?~��*�o�1��bX̓`��s��;M
���=w�t�<)U�S "B���^�xTx�Z
Q�<����G���-�#
U���T��O�<Qテ&ݺ�`��5����f�@�<a����Ҍ��Ѵvʍ���@�<� ��&�{Ӈ� <�āp�<���Y�B5���׳*V�e�3-�v�<�v���p攕P�Ƃ�wvL�ѩ�K�<13 �/m"&P��NZn�! fN�<id���Ԥ�>p6�Q�VR�<A��9 �:��\�2�����K�R�<�t�Z� �����y�6u�4�QM�<�C��T��K��K���{S%�f�<�d��P�R���Ki081[P�Vg�<��E(\��}�D��tJ<3���D�<����$$ �X�B��r �A�<��N$(��SpC�P�� �`�Yj�<�
ߣ(Y�@��@�
�y�g@e�<A���VTllá���r�J�a�+�a�<�剓>;W����Ȟq�l@��"D��3����$�3��pVp���!'D��3`ڕN��r��Ȉ	�Ppq �%D��W"Ҭ	�n<����TB�r��%D�Hy�o��#ΚQbpmF��v��M/D��"�%K!Q�TZCÙl�^ҁ�0D���Ug�m��� A+{B"�.D���Ɠ	2m���9o~	�I/D��F�V�H	���� 	Ap;F�-D�$��+D�g1|�q����&�[��*D��������Ul�#m7ܬ!��*D�[TQ/X����.߳2��J��(D����혋u�8ys4�V��`�A2D�0$b��+]�a��h�H��ԛC�0D����(=7�yc���7IJL��0D��`��w#�1�u��.P��D�,D�� ����C�%8tY����L^�iv"O��C��Q���� ��_�`�( "O�)٤�&S:�q�`�4	���"OR䠳�!�Ψ*D�*���H°iv0#�'��	rC_�cd�rǋ�\�Lu�(���2a7?�s,[�xAXݑ�GК~Dp�+��Vz�<�!!Ö9:�<��	v �+��X�
��9�c,��A&�M5.��TrA�;u�=�"O�TQ��]H3��b�!�I�"81�䈗V�qO��#��Y���DNݫ}��"�$�)ۨah�M2D��ۆ�M8l�fbt�+l^�X�>lȨ��6�O���*� __�D3SiR�m���'��H�da�A~��G�<z�Z��O�tP�'�Q���x��-��!��l��	��a+�+f��Z�x�FV�cU�O�On��b,I.A0v�v�T�# �9#
˓]�n�S�.���|"�  !(�b�P��R��'!�$]-���@n��1�a�F��%���VhZ�[6qO�����"GƷp�`<J��m�PE�V"O�(�b��Ey��FI;d�%"�,�	��-)��L<�Q�H5>��k֮�$�f4(7��vH<9"-?ԨhI��M,Uba��E�9ɖ܃0�*�O>��d�_U�`	���R$���Q�'�D�*�K�M�I �j��aD<1U!�$�!XhDC�	�2�\u`a̞��l��
�&��O�`��J?�)�(R\�6��[�M����P+B�	6Zժ�L��A򋝷V�B�I�^�F�ߺh���5↔r��C�I����b�S��";}�C�7s!L咒(d���N�(�C�IKe0�KV��0c8t8׃�G��C�	8��{@A�� ��@���C�5kh�Iq�
6�8Y�	,A�JC�bX�{'D��q��ATIG�#-.C��ol:8P&l�j����BB�I�n����ٱ��	��ЂS.bB�7�P\[�J�1y��ce �׊C�	�H�]0�Q�9!H1�Ԃ�Yo`C�	�.�o�;FR\mKB��e)RC�	<�h�aԈ̕e�\�8dmA�(C�	�7�\̺r��t>���� ��B�I�9a���ҥѤ|�{b�"'�B�IC�b1�FG�-OX�������4�⣓�5��?M{a�`y�,�7��5�|]��"D�Db�(����Fه"x��`_��ؠ0�|rO?�g}2g+4J�D��?K񌽠'�,�y�]�)��񨧭YA��L�fD�ڽ���yܐm ��N��0=ɳM.^��e�Ee�"~}�|�0�Fpy�-��T�����|ZwV^5�wO�`��ͮ5�4�i���+ ����'�҃0�P�'��t(�"E�k��+�/��h�!���01V ��%����X��T�8'�b�qq�]�<&�=A<��v��S�	��/F�9/a|Х|3�Q!'^�_Z�)�E�]{
	ӧ�Z�t��Ј �T&UP��2~_��a��JXT��e�~�B�x"E9z�r�3gۿeI2�6��э,��ں��<I3ޱ�'�^�&��i���	�@�	?q�&iʠ$S�R2TԠ`-F�s7�$@*�K����<)��3c�D�%/ "D2���	�0��%&n�5[�*1B�d�Z����3a�l��/�!&N&�ɵi5��%s�?����u�ˢS8V�(�*��u|R��Y��(2�7u
��T,��t�D�Zӫ�u�RLXs� /L��1��E�6���׈�4r��,͐r�L�3ًs�@\`s� /q���2��G���4bU��#x����D�~��@N�|�BE����JJ,���jg��qPR���v�m��D�;��0��"H\r'Ϛ&KL.����	�g����ٓ�I�a�ҹ�N�*V���8$FX%�c��9&�:n��zg9�L����?E�D�Q�e{HQ���_�,�#�$\2�y#6g��:ޕ�%o�?F�|�UcX�cw\M��A^� �sԛxr�'��lذ%�"k�n��&�J�Z J@2 �]�1���:k�<��'��L�e� h�j��<+�n�1��Af ��VH��Ni�b�	Yol�(4��o���)�$ΐ��,3L�"ׁg��,�PC[�_���2��)ql0&H	�7�����*,1B�B�A�g��,l6� |��FQ
>ԙ�'�Qf�P�=]�6y��]x��@R�^�^�:m����؀ �	Sd>�6	�B%B�h�|t�B ��1D���h2-^0doZ�[蓦ɾ5z}
&�
�o�\��0� �?qX#V;M
R�4.
	p1�� ��!�r��fl�Ojf�j�'��nEr���n_>GAP�I���)ts���D�y�ըH+0/2�
�n� ���.?DF^��'1.h
�m	2*�W,�/.�LM���Q��0�B����铄5$|"�k�W.*Xh�#�!_d�5	W��	���Ae�1*)���]�s ���o���k� �6��j���%���'�Zh���]��)�'�)�^�n�;,�=nG��AS�V3{]���G�-��	�d��k�(a��pE����i�&}��含mV��OI/|�d�4F2a�� B�0}r	��f�Ʊ[�D�}����o��1�8�P��vܬE0wBΩ��yK1�	�5(4�����rڤM�~J�G[�X�`0
��S�G;�Z4�̌@p���%� G�.�P�C� D����Ox����<���&��ƍ�9�z	�Ѩ��[�������+ݹB�:&`[*t嘨��g�-U�ԍC� ��f	��"���-��J��'�X��w�@-V}�%��5ΆP�'`%(p
ʌ/%��Y�>Ap�T�XZD1LI�P�H���L��\1��y�G���(��2k�I�b���5���E�S��~	���Qي��c��1���A��ӱ��bL-a�¥f9f�R�9~��>`�gّtVdk7H?7*�x*��/ʓS��80g'X�|Zt{���o	n�r�@#@�}��,��G�"��L��.�
0
t�WoO�z�D�𙟜��F_�xE3Ŝ�ed��"�)h�=Y�n��PWƑP.O?��Ӓ=�1{�!K�?Ḅ�gMZ:)a�#_��8�s��}�d�5��U0@��a�C��6 ��)�J�>���X�\� �l!�	�]�(���9T��z��0az�pV�H5X�|�`g�-��(3�'W�Y�b��3b���a϶~/5�U�Z$6�����V�zt`����8�� ��׭dl�ȰgG�|��&��p�N��T���x�@A$Vu�<YW�-F��IP�I���@
u�j��R0e�,AQ)xO�pl�����y���Z�:��+�(�DA�����y".�Sa,���
�UG�������j䜰	e&+R��`h���a�Ƀ��T��E��f.����&�?h�bxc�6A��~�2K��pA���q�"R��X6�,�B+�u�<r�UZ
a{�<20&Yڔ-�+h���ܩ��O♡ai��n�B@����x�ZIZa��������
�$�g:H)�"O�=��(�"��s��nz� Z�<��bL�2�Y��`�mCr1����G=ꌺ`�B$*L,���C7JrB��*@*z�(�a&��UJ��@=0�b ��A�.O����Y��xgOٽ:�,؛a��� �:�Z��%D���$M
��s��?��0� a�qՔm�@�=����,`�vKƶjWh!��Ľq:���C�4���@lڗH̙���ne�<uK&eJjB��/$�2��& \�̌L��M��-Lc�h��K�G����@���4x���_5���A!�z��C�I%^ <d�͌7
�Ip g�%+�R]�%��&k�ΒOP�}�j<�c�lΩ�8`A�DN:oq@����Li�f�U.,*�q��;G�*�ȓ"�(@�@)-�̵H�FF2|jnu�ȓ � qU�
M��w�W� ����ȓ���Z`�zAZ,���1>�\��O�T qO,�}��l���*cx^��]�TI>�ȓx�%9��8�J�#�O�<+��n�%�
`�B�i8�P��D�a���-��A	��25b6\O�ac���}�F���'��b���1$�������Y8���'A��9��_�x�噲��َ�!�{"LɀhM�8J�MA�O� �`��;Uz�2 *�� �'�����Jҷ)]�F�ζ!����e8�*i�J�����<P��̆KT%^,B� ���i�<��NI�kw,�8򌒠c?~�  j�X�'S�&�"��(��(�&�ްDA0� `V���A�RM�Z �E��y���in�9`�W?R~��0��N��yU�?�.J��L-��K����'����Ņ<�b�E���!���(�/�F�Z-�pjS6�y2� K�n}�a�Ō0Qh�{Gǉ�rL��OV7���b�Q>�|�����b����;Q��хȓ~�����kd�P��1'�Z�mZ�bҚ�K�!�L8��b%�\�i� i�BJߎ�S ,|O"�ԭ������=ZsV��`�ζJ�	��}k!�d�5^1��Ǉ�q�M� *K"o!�� �8"��U+�RQ��r�n�3"O��� �5�TXJ%�M.0�8bC"O&�A3e�S^J	*�͕�-���S"O��FG�|�3%0�*�ѥ"O6� �j�!�`�wn��@�@"O0�z�o�;�] ��� i����"OJ�X�lO�/J8T��� ��L�T"O�dK`(^K�t}��Ͼ4��,��"O�Q��S�Fs��9��5�V�а"OT	�����ĈF��0�d�"O:U��_Nj-���y�4���"O&���N�M��V䍐C��-j�"O��JW�Gk2�9FYAR6��S"O*D��5p��	�@Kj(��"O��z�ƀ>"B�����"*TC1"O*x�
*D4�i��3"�|<��"O�a7���x�ɑ*Dd�:�*!"O�-(�k�&(���Y��w��l��"O�l�f��&(C℀7G�&�\)� "O|\h�#�b��� ,�|+&"O ��2,�7!S���
��8|�1"O���`�1-^޸J��d����"O��� ߁N��E���>��Ԓ�"Ob��c��CN^YH坫Y@�i�"O��@"�c��l�Cˏ�G��\��"O�Lv*K<){��Y���8�����"OL]�]�n5
��掹1����"O�ܢ�4�b�H���!G�����"O��H����>�NE���7BK�؀�"Oh�Q�.���d�aOF)S�m(�"O^)bU�N WVX�2��	onµ{�"O$9�7�O�J�}f�8]f	i�"O�ap�cL�5��H7gԓH�B�H�"O�%#�H�>L��Q�2)P��|�{"O*�9�+�~�ڐ+R�Nº��R"O�pF)f�ȸ�/�@�|��"O��3�R1+#1S�v�K�"O�U1pBD�FW�d���N�bx�|s�"OK���=�ѠD�ie���"O��h��O���H�U@^@����"O�dH�`ћr��lbA�N=v�\�Q�"O:�r.W�����H�;�J��"O�D���i�@�cMW�>���Q#"Oƨh� ��~:­��L�>�4��"O�Vdݫ)%��j�?V|�S�"OR�q���G��H��
zf"Ovq3"��	�,�+bi��ڂ"O������7>|�*&���`�"O�9�5�`a�	9\�:��iW� !�ě�B�f��eG��.���v���#-!���)��@�C$Y�ڕ���7!��H�����>d"YC�o͚C1!�$��6]H���JW#F���ڝc\!�@�GU>x�qo��k]>p(��!�ą+,|<�b��:Ui��+�N5)�!�䄔��ɡ`�V=,��-ΚE�!���4w�xCV���b�LqslƎ&�!���}5�����t����Gh�!�$ܷ\�Б�tȄHF�D����`!���Mt k�A�H7���u�!�D�n��ʓ)�<@֕c�c�: �!�� �2	��)F�i�*��0���!򤍴�Yy�N^�^�H�[��Ȩy�!�$V3*0��b��D&�E2�(�6nS!�� ��!��-�.� ��ڂ\K�"O�(��	�V��2	��d�s"On�� ��|����3��6~����"O\d��i�N�hr�$d����"OԹ�>�� s�D�0S��"Ov,(ԧS+eu��j"�W	�0���"O��#S��Y��$�#A+5��#�"O��	Fa��X�ZY�'"O���r�"O�x@�Ì�;�T8��8Eyv)�a"OT���Ɔ:-)�n��;f�4�"O��ycj�9	���.�����"O4�+�C�y%چF�X�.�:F"O�p�r��|碥��o�7�$���"O�H0P�Z<�#X�4��䁡"O�Ly�Díw�n�����6��M�"O ���Y�S:�l�˾���"On�1���� QJČ)(�^�p!"O�H(��2" tԘԬ��+��\�"O6<Q��¸�u�2��%�>�"O}[�a@2z��P��	�/K�*��"O�m����g�X�4�
"{��IZ�"O胣�ѦO��5`�ۖ>�<Y�"OX��pR�e����	��LUc"O�9�#�X�%j��G�3�N��r"O
q	E�G�A���# P & �"O����➖@B�q	���
	���"Ov�3��F9�~,�A&�
�i��"O�`:�[�,c��S�/L�u�T��"O�L)�E����Ϙ��{4"O��G.�)^����qM�:\��"O�5�vFF��0��NR$��"O�IPӌلPUً�ʄ"!���"OJ��6%��M�|��B�_���Z3"OT8��Mdܰ��s�ǲ-s2�R�"O��˛/@��ї�_�
KDd
�"O(|4��0�G�U4;�X�g�<1g�"S�H2˂7�l�pl\�<��ŝE��3��KM�T�
���f�<1���dk��g>1kr\�u�FH�<��
De�t��";�b����p�<ADf�5QVLK��`� ��͟r�<1����z	jE�PH�$��Ēw�<Ib�Q���X�&%��+�F�h�e�<��G3q�h�pD:$�^L��-x�<�7��!_�$�U+I*[����⇂u�<��l�ր���ռl�d�f��l�L�h�ō9�'| ���<�TiAN�',!^��Z�a�U�%��1�	\f�v}Ұ+�^�OtuF��O�q��o4;pp)`����jr"O��z��Q/*��ڴ�K�%�V�&�ɨ&���Т��L���K�'�0���>Ro���V�D̴.OJ��f�9N`�O�ۙk���L�c�:	��\*2����FH��X��QЫ��dP��d
��Hg�ղy�c�\;y�$�"%�}�Ƈ�:r��e�"��&�+r�Z�my��Cg�x�}X�-9x��e�C"��`Ä-9�O9x�G�&m�20�f��p@B��*X� r@$�Āԗt� QI�$�O���JB�DI	BiaWJsEF�O!�O�𱳩� |���ǇZ?Z�Z��R���#�SD�$I�O���hM8��P@��9zNu�5f� {MA��h�7(���'��&Xo�=�$�DX�4�F�^3:���C��Rj��
n��)��-�g1�hI�AƐyШ��^29��IV���W~8���k���¥�X�D�<!�BB�j�j!I/]k���ȗ��IqƇ�2�@��v+G��t)�N�btVCp��)k�`h�����Yq�1 �T���F�
�k��Ұ u�˹k�HR�.ٕz�����'H�9�r��7�V��j�&(�ja�!R�Rd��#b:vH���t6=��Tf�23���Ľ?��R�Y~�U�UP�}P����,*s@^���'�� ��FB�R�Za�Wq8R���O��:v��($�]�U��?64ɱ��јoӠ���Q]Ǭ�S3�-3����� ��9�NU%:�"�3����$,~%��*L��L}�S��0*�z���9�����$>�6�s�BA���N*6{P�+"+�'�VD�`��(�I��酊'�(q���zǼ��ثD��ث��E�6���w��?h���
�H=;�^tP�I�zŲ��FX�D�����)4���R���c�Z]t��;0�o	�x�퉹x����lC��9jDHEdH1py�m����9-i��s�F�WL�<S�޶t�Â6O��x�*��X,P��WM8�۰-�{Հ4�?	P/Z$ ,�P��i���̘c�	��E�
�f�L�1r�"���~B @7Xa| ��k�U�hᠯ�V� �3!�2A���������0p%J �9��S�O=�x��	�uZ�BS&ػc�Ų��ƃ~tlPJǰij�cW�\�ZU���� 	��h`@�$�d�����d,�	6f4Yu�F}�	28�!�i5�|X�'���X���6>6�p��"d�r�	��p>ch]�'�0�I�m�iR�h2�S�?:,t��Y"Ym�Q��}���n�U�M	���[$e��1xx�H�뇻{��k��I�D�9�%�5~p��~Z�)@�Q0��-.s7����gګ�1�E҉}ڼ�槈��䓄9�ƕ9`��v������7p>A��,]�:01J�y���'��fL�A��@�D��gΜM��'�کC4O�&B�Uc�L2�Keg��JC";��˗�Vp�:2|z�!�W�0P�}�@) ��"��y�f	Y�hL=e��[sM,`��I6|O5����.�|!a'm�A���c��> ��lXՠR�&�R�\���M����GB#��O�2�a�&7z��p�D�X��q��$�$�&�1bf5y��b?�0�ժe�9�Ӫj�:�e��z�L �0 �lj�G}���iY���� �),�p�*��y�f��
)\	���2A��M� �S��?q���֩���"�N}�aO�Z�$��F<J��v��0<9���&��&GڄLtL�*�DR}�GƱ;�,p�#�i�'M�=iaA��7��Q�Ϸ!,ԃun�*���(c@�y�����/�3����gEi=I)v�д{��0�3+
l�'}\����g�E��H�<����'%#� �H[%r�0�C�^��P������mڇm��I��@�1��t�o�0D���������
]��F�d@D� ݶi�6�A�-�H]+�Mг�y�L�a��� /�h]��)��w�
���'<�����W�]�N�PO?��>�F獏'�4Ec��;+{��2 %�]��LY#��49 I�#I����{@,�*���Z �Ѕ8��(��ڽ�*ń�	2�6�i��:0��"�b{d"?��i�"Y.ؑ�_<< �S#�ٺ#u
��?�v�]��\����P�<�b��N�*ĺ�k���BiOy���6R��#�#
&R0���|�OӴ+g��0Y-�ɲr!+@�xc�<�S�^)Q(�k� �>�2��ݨ=Y���<db�u�Q>�X�.� 	o�.�@�EQ4�p�ȓVݔ%��e�=4��@��#Ŷ�0h��ٳhW��#ꋅi<a{��;CL\Ѵ�W9<��a"֤�9�p=�u��9t��)�.п�MCu
�����(^�l�lK��p�<��
*^0i�C�74*\Kb�Pl�WŚLD+S*�z�}�����r�L��W�e���"Rf�<�c��q�r��3Kψ0�F�`� A ?4�x	goN�	`��~�ւ2�-Z���
+�F�7�y"5{ �u!Ӹe߼���O=�y��Ԟ=�T�pf@�f���)� �0�y�	Ԕl�`8p�;_Q�墁��y)S�,��іo?R��`���;~�6���?�I��~"o��|nmK�愂���BW�y"��H4�t/�7@�9�ɉ��M[#�Ad��Y�)m����F�%8�!��q��=��	Oy������!~��ی����S�	Y �{G��O�!�-z-� �m4<,V�N�9�qO�gQCld�{����QN�����
mk��V�&!�d���`*$a�f�(�[0�:zS2��Qa�'@�u�|�'7�rt��-�\�K�Ϙ��C
�'N�LY����{t<��=n(�(��VQ�5��ǁ2�0>Q����,��A�%G_	e���W��Q����'����I�S4ON|���@�\hqa�/ѯl�J��"O*|g�>�"���A�6s�d�w�$�8F�l���!�9����:�	��,x�®^φA�G#!D��+EL@���P�:0~��#��8Q�
L�J>}b�x����Y�)����a�ԝR>�y&�ÓV�!�� �Y"�F)a�t(�w�;i��iE&� u�$��|"��"u���F'�H��A˒��=�d*Xu�.��t��g 
��9��!�4I����ȓ�(}���s"r۳KN/T����8b`��o5hY*����]9�݇ȓv
U� ˠ/'�����s\���Ny�غ�Gܪz���;e�<RU^��t�BDQ���""~��`C�' cN���x3�\IB�
�u�n|���c�|���9�j� �❍v)\��H���ȓ,��]�p��7�l�� �F	�ȓ|��h�ML:=D��Å�j� �� ���r��z�J�@P�
W����D���� �	q"���վY�bD��S{Jx��,�Q�h�G���ȓ5P���j�*mzI�	�"mqn�ȓ2�1q��߶?�P\S��"z�dI�ȓL���Q�R�waɲ��X�EGh��ȓ�4���ѓz :�b�bT�^��_�t4�b%ATb�E���,4*�X���F���R �x��ce�,���Y�'���xT�ΚS��5�A�(�
�'��J�V3_G
��
ݦ2�� 	�'���蔣�jd��� -��+�'����qf��T�B" �/ ��	�'��X�B�3}g�9*������
�'�d}����i�<�Ï�;e`�Q
�'zq�r�Yj��8aF��zʌ	�'��Q�A �E>fa��EN�D��'�����L�\����ň>��9��'�<�y7Jʹ
ă�҆ �a	�']�`�פܛo.��УK*��3	�'|p��9�n �S,��w<�0�'�A���&[��3dS�����'o�AhG����\jqkW�p_d���'�8�)�扎p���PNޫsh49"�'�p���le�� �a�l�@Z�'?���+c`8ya!�0}�lLَy��O�z�rp��ϋ�<�A�fR���'Z��Q�|,�i !�7r��Y�'��ᢢJ.j�<��R	p����'zh��e�G��\=*R�����'�D���#p�+��J�4ƐH�'�dEz���Ta�Tb���g	F��'*�s҉[�a����v��'t�*);�'��Z׬��m�b���ɲ_�$<i�'�����;u@��"1e�Q�4���'H��BP�{�$+��V
Ji�MH�'�D	 'P� ��!�劆��x��'��"=E�@C�4f�0��>�
t!���gg6�Bs�Ocy¥�6#�����-KE|�ʣ�އ13L�X���{�xݺDT���q
�
�����O�8�ZF�?Q2��K〉\�����'I���1��M.���]U>�YR��	3�ݹ&�K�%ņ90���%��� ÝkC�|��)�q��b:`�8�d�m�����^�~m�%(�#�CJ��h�����������,k��Y!֬ɉ,
�T`��>�R�X�=�����/,r�9���4NҪa��'��	�h��Q�6,�)���5����g�I!B���t�:qp��+~W�*��<�)�'h��mA�6v�6Q�$mR�z�J��ȓW��@��3"�d\��������ȓ��0lɂp�V���ٍ �5�ȓN>�ٛ�
R�
,+�hJ�(5GzR�'�tӥ��?� �E	[�yg��'v ��`J�	�.����Hz��xp�'� 4a�f�4��`(�A�'r�ٹ�'�lKd���#6����HПǪ�	��� r��l�`"�Ѓ�{$�h�"Op<���=J6�0��"k
��R�"OL�4�Ű �l��'�#h
�uRP"O��b�ր �hb��خf����"O��btJŊFX$��C��f���H�"OVec� ߒP��P[��)E��D4"O���D	JMA��K�
�R��8"O�	���GT4:u��F}ϊ���"O8��@#�&�VI����&dv"O��
��'�貴�D�+�P���"Oh\9�jCb��5��G#<::���"OZ �c�]�0Q��fi� " -	u"O�	A'f�$-{E�ԑX�A"O$� Fē:�A��Q�`��Չ"OL�c�A�T̀� ��.;��۔"O�u���� ��4�0C{X}��"OS�&*^�P��"Ɓ.Xx�"O浑B`�2_�,�+���Ie4���"O�R��k%�ͱ��P';O�p��"O |�jIx���A>=��W"O:��t��8YÜ<i�l�+U>P���"Ox`�ע��ę�+P�x89�"OV
Q#�x�������"O �D��i���ҷ+�1`~���"OlmS��1}�� ��.p�dV"Ox�����"$����(��6i�d�#"O���&��;@�ذ��GIPf ���"O����@�6I���#���dW�@["O�@�Fd��K^�!��D�3cT||zG"O�x�u ��pz�!�<���R"Oƕ҇bU�~s��"� �O�N�y�"O"������i�/�d�	p"O�h��B|�H��%�HQJ�A"O@u˶j�>�N���7�b8a�"O.�B�&�yV�b#Êh5���"Ox͒���z���*tC�-���S"O `{!���^dꑄ�=>��"O�����#���$cEp.Ƭ�7"OM�È�2p��ⓣ�r�
"O��3��ri�+w�M��D1	�"O�e���P\�V���O�C�蜒b"O=���ڑ�����@]�� �"OF�b�4��������HՑ2"O�!P&"t�$spE>P�|4s�"O�x��iI7[]r�٣������U�!D�t� &?K�{`b\�R$��u�2D���0g�\����Y�k%���2"2D�����4�(d��'V
o�Ыa..D���f��3�-i��8������)D����C�)��mYↅ�.1bQ 'D���&��^ncf��:~if�0��0D�PQj��=�Ed_#f�D�I �.D�\�@E��WGd�w ��oO���+D��R�/N;/[>I��YQ0+D���a���7�ѝ��rPL�Z�<9І�j�����/ra���}�<�ckS=�K���d���fN���C�ə D��:��;MaPE�aI�8��C�	�^s�Sm�(J:Ł�-E�M�C�ɬ&�� ��U3E�R@#�	�D$�C���֐�pmW 2Ft3%��$��B�	%Nm�šd������F�T!�B䉃}��@��Ή|��cP��]L"C�I=3jd�򷫆t�����k�6x1(C�)� ��	�*!�j n+zy�@"Oj��s!� p�5��ְ�T%�Q"O�81파E6b)q�9(�4�kQ"O�-��.ΆZ&LT�}��U�g"O��� '�wj�²����8F"Oք�6�.�*��؜��(C"OԐq�6�yF)zZEС"O��x���!L��J��Z���p"O���p��=&f Adb�w���f"OL���A?:0ha;�c��i{�)�Q"O ��oX�]��<�C��:9�Hy�P"O�|���	O�8�c߾n���yw"O�遥��C�.T�g�Ό>�xf"O`�H�B
39x���H��t��"OX���-�68��B];H^�"O�x�pgC!n�V 	�CʰTiI"O�] GㄚJ����U��i��"O�$��\�c������)���4"O�Qy�!�'I� U���Y]�t`2"O+Í�;C��Dg6����"O
���M�9�,ܐ𭀻�|Hx "O���cD8)¤*���\�T��"O��±j�%b1<�{�j��Mf2��"O�	��i�2gbtY�L�Fk3"O��a�ތ{	�������H�8��b"O��x3+�Rw�L��Z�s~�YX&"O(�seMٖ �B�BaB� %��a��"OR=����,1�K��ŘVX- �"O8T�ՎK%Ny�5��䄨p9<=Z�"O
��ꅰAD4�z��S�+
pa"On(�S�:L����!	8��� 7"O�@�
ɽ7���x���Yf�k"O��藠
6�T��6Ep �"O4�󳮜�JIĸ�w,�+]-&!1�"O�\���\4J_�W�^�#]ó"OB����>/WN�9�,��&x2#A1D�|Js�Îo\`�˗�8a�TX��-D�t��	����d��`��1Z�+D��'N�RA�YАg��T� ˵)*D����T�2��礃�l�����(D��)V�3}�l$��hC x��`E(D����A��r�3�\�#� p��(D�����Q�i�>�k���:�zq)5n%D���1��n���
d�9$���-D�JW������-�H��(���-D����b��y�6᳖��h�hP1�O?D�$)1��2	�zLZcE�!�|Š5(?D����P�e,|��!R�d�zq��=D�t����*q̰c�
�%]��y��<D�|���45����������:D��7A��II�����[$����9D�8;���68u����3:�k5g)D�Y ��t�ְ�¬�<fQ��0�:D�|ɡ��.�t�$M��/���#D��xujɈN4ܫ��[�d��4�R� D�T;e���,c��)���cP�>D��Z�-T� �T�#3XP0�!D�8ٱ�W	�Չr`V�uzu1��1D�xB�F����U�CZ`�Q��3D��r��ڗ>;ne�fL՘GU�YZp�6D��C'O_N� �̔���M0u�0D��;��E*n��Z®ђ���@<D��Y�)���H,P�Q���w.8D����%AB��⨎<ƀ�b�;D�� �̳<����/<0V�\�"OV�$�#�p��͟�NFJ�{"O����{!^�[nY,eǖ�Ce"O��ᢍ0t_���Ae���#u"O��f��
ٞؒ��Uhc^C�"O�]�i�/`��"�HX�,q�m�P"O($�iH�E��y@���>7P��""O�!B#H�W7֍k�aUH�8Qa"O����K4>�
y:��\>���g"O�0q�	{�d�"����+xx�"O�!����jk>y�㘌}�:��"OȘR��tL�"�a��~�쳥"O�Y���[dd�j�a�!=��H�"O�8�6� �S��z���!"��q�"O\q��*�8<[�C�Tv�!!"O�	2�
;��A��c����"O r��.6r���,�>���Z""Oq37�@"zw�}@�j�p�b�S�"O���� �9�.��(��޽��"O�8�2�UWu�`��L�(7٬�j�"O�Y���E�0���O6�^� �"O>��3�M"}�N$��m����"O,)D���xAd���ǂ��"Op���E��W�L�ci��U�p��"ObD�aL�L�z���U F�y�"O�q�K^=pO<���ܲ.��W"O,)Ss�P<_�,Da�7+BM��"O�����4/�:;�տ<�0��A"O�ܺf$OT�S��Y��|�"OX�3*X!�V��EV9,���"Oz|��K�b�� D��X�A��"Ojt��3׶��AB��w"Oz���	T��pA��r� �"OHX� �ʭ6hJp�r���@��:Q"O�]�1�d��u"jv�y�"O��)!�^�q�t�����A"O�(�"D!z��i��C�6��Sa"O��ӇF�#qp��C�̿@�Z�iq"Oΐ@�DT-V���s���4)��̐�"O�M�c�R�?q�(4"��0�(	��"O��R�aĨ&,�X�A��<<����C"O��P��I�m<�[B틏7���T"O�Ԁ�F	�xW:3���[�䨦"O� b�h�1]�|H�l��)t��$"O� 2�'x8�Br����'o�j�<�nKTj1�A'۸'dD@�W�A�<9���:m�e�B��t?�,2Rf�A�<�W�Ʃ-��YIQ
�Z&�av�}�<�!�IgM����ĎC��KVgv�<QuLC<��,p�49�-�r��z�<Q� �"d�B �R`��#*T�<�`�J�rb�D�"�M���j`��_�<y�fQ��DE��F�<$�fLҤ$�^�<)�F�>���1'��Y[xE*��V�<���ڤ����Y�NY�����N�<1��N�m�4A`FO�)3���I'�q�<a�ID35 ��VKJ"����D�b�<�	Ծu<d�b`�K�l-���^�<�C矚]�TQѥMΉpv*��e,�~�<�a��,}�,����̉!��2�)�{�<�cR%/��a�"�ڼQ�0P� .Tx�<�6EU��~<��f���ybH�I�<��D�$H�H�r�®~th�G�]�<qA�Z�&-!헬 �̱� J[�<� x��K1M�!J��9Gnm�"O�Tۤf��!�̸@�<��b��>D����9Mf������x��C�d*D���u�   ��   �    b  |  �)  B3  �9  =@  �F  �L  S  FY  �_  �e  l  jr  �x  -  �  ȋ  �  ]�  ��  �  %�  f�  ��  9�  ��  ��  ��  u�  ��  *�  n�  ��  B�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�VO&}��a4/zY;�#m�����#D�D1���'�01Vo^w:,�U�!D��1G�;(�x���n�$X�6@?D�P�$�Õ�ha�v�C�y �a=D�t�+�p��xj�N9N|�C�<D�:�K�<M�N<ca��*�Ĥ8��9D���������%� .�7Ẕ��<D�L�p-��h�u W$�[Ri<D�������e��E��V).�&9D�T*� -5��dKq�߾{|��聥*D�\�t��J�9��D,~|qR�&D����O�RtN�I0�6S�L�jUC&D���f�a�R 	!�j�T���$D�d8�FD�p��a���t�L�b��&D�|��揺-����e�˳I$Z��A�7D� �Q��,YX\�;5M߾[~X}��5D�p2'����(��R�,�^)#��2D��"�V��V��7-V,�^�QEF#D�(!�c@�x��V#�FP�-&D�\:�英B>��aι�m��#D� ���9SO�ؠE�l��В�'D��x��̎j=*���?�J�A&D��Z%��.}> Jr`�89wQ��N>D��TBԖoƾp�1���HIF	!D��-�$[� ��T���p`��1D�d����S�����K�,t���h%�/D���Cn<5TP��޽2�x����-D��[#.1S���g]�?�d�Q��,D�,��'i�踰�E391`�֢/D�@�OH=�)��ƀ�M��4�,D��8V"J�Rxv&� +�4U��*O6�E��#Y���d�Ѯ8�*�HS"O�H��E�<X�b��hF�U"O�cQ�0��s�;-�q	�"O�P���,�.�8qe��N�% �"O��HE*UR�����]U�T#�"O���HIi:�֧�\���"O��[����d�@��2�"��"O�kҎ��.����o�-|�Q!�'�B��P��B_�TQ j��G�II�'<VEZ&��9/<Փw�׳*`��I�'ސ�������Щ� /���
�')�9�#�W�cp
��
тTx�'.ıRV�A�Ws��id�D�o%8���'�΀UBDE7�³j�����'�@	�W&ŬI���K���-!س
�'qPȻ�+Ӽ	��E��
.�R�
�'(�D飦�"�`5 W:�U�	��� �<(Ĥ�
N��Y��KUR��ۣ"OvtSqJݲ>,8�&��w�2|i�"O��S��^�@�
�5/ɬk���2"O�X	A� ]1앪1���
1�(��"Ỏ�F�>�`y��-��He�'@�'2�'R�'���'��'N�
 �A"t��I��޵R�0�{��'���'B�'���'���'��'��������)�/��{jP{Q�'�'���'�b�'�r�'��'�Qid&Ǹ Ub4�^�l'邑�'y��'�"�'���'Cb�'-2�'w�td(ګ6���I'Kx��G�'�R�'���'���'~��'A��'��%�B/�K�lX�5�!?�.8*��'�R�'�2�'���'�R�'�B�'�V�A���mО);�,ӎz��Ybt�'��'���'�'���'���'��Q��L1�tT�����.̋W�'�"�'��'2�'���'���'�N�Y�D�%�.A9 ��k\T���'���'	��'�B�''B�'ab�'���4��%%%�!	vMIx�J|��'���'�2�'���'3�'�B�'���X5 Y��N�3ӭ�`3x�҆�'<B�'�b�'���'���'9"�'2�p��f�_��Y{��JZ,����'rB�'���'r�'���'P2�'|�Ju�ݤi!����늏"µ ��'x��'�r�'X��'�b�j�����OtUP�GN)J|�!r�Q9���`&$Ey��'��)�3?Y��i`� �*�Ɣ`�@�,kx�С������O��<�'��A��`:�#M�Ι��l,[��'G�����ia�	�|RC�O��'J��}�f�<ܴh��FԤk����<����$,ڧ �ԝ��@^iۺ9�F��!\r����iH@��y�i�O�.�rP(�{fb��Xz�X���O������O�	U}����b��F7O|*ĩ�3"�L��D�Ew
�H�9O"扔�?Yt� ��|:��k)����� t��(c'w٢��p�X�'d�'�v7-ږL?1Oq� cH�GԸ��`�2r�|���0�	wy2�'*b>O��\"&!�2,[p?��S� W)�+ ?a��Q���NY̧Q���N�?A��W}~P�&Lܼ3��Jb#����ĺ<A�S��y��!�9c6O�3qm2��b(�y2!r�Ft�4��h��D��|2�IU80=x�h��\�* �	���<���?��-)ݴ���i>�0��U��u�3��O�E�5������K�=���<�'�?a��?���?Q��ۧJ(<�pwc�"s�h�ivD�;��٦�RM��|�I柈'?u���0Q 4��@A(�)t"�:*~D�'�7��ᦵϓ�H�����eZ�8S��@��jx����6Q�d��X�����ç&���I�Gĉ'.HʓPL�y���Ig>�ˇ��n4�{��?)���?Q��|2-O�mo�0T����ɽr]��6������部��;b��������?�+O��m��M��Ee栙�J� OӠ�Q$��B�n��+�M��'@��km=\b��I%�ӽDfk��-2T�PTm�-h�����l��j��d�O|���O���O��!�S�A��0�Pȏ�w�@��C�*0Τ��I���	��M��F��|Z���?qH>���~�6T{�Hξ'�\l`�R{��'�R������Ni�v��싧�R�(wL\K�E��;�ޑp ���(<���'K$&�0����'���'�	SE�7Z�(Y�F�*l�Ea�'tB_���4h�������?A����]�75\\�bh�n��T�FM��e��	P~��'��f�:�T>U��g 8y`ezB�� 6[�ѣ�]�&5��(��'�P��|���OH�L>!��N4
`���U�@�9�!eL(�?����?����?�|2-O��o��HH4m�qϚ��`�8�^:���PaFyb�'��OZ��?q#��xy�B 0�T�c
"�?���i" �ڀ�i]�	�L�P{q�O��/b@' RnPb���K�ϓ��$�O���O���O����|����5c���V���m�(�����ϛ&*��V���'3�����'��w�l1��g��H��I3I	� ���'���:��)V!ch�6�e�����	�7`޴JeE��N,x��{�M�US��DQ�Iny�Ob��j�� 1իS�Q�����0W��'�B�'���/�MS����?Y���?�폦z䒘���M<:=����mߨ��'A�IݟT�	���L�b`�
)p[�IC
C�]�'�|3��\,���[����ٟ�[��'��y2Ԍ���$��s�T|��'���'��'��>��	3fA$X���B&�ң/��h�ɣ�M� ������O���k�a��Չ;�m��g�s>�	ޟ�ɤ�M�+آ�M��O �i�B�RG(U���jA#	<r�����.2�P�O���|z���?���?I�U�X�a�V�h鶸�Q�Y7D�\�j)O��n/\ɸ-��˟���u�˟�ңˋ1�HP�E��iW�I�"�KyB�v��Do����S�'�^}��c�Pp�3��/� <�靤);��'Z �z�ES��L4�|�U�xc e��Il�9b��M��|��%n�����i�6��O6�4�.�ep�6��/-�BX��2%V� 4�v`O�$f�'��OV�?��47��O�|�̜`gBC��^�y��!�sW�i0�$�OH|��b���������� ���4b�.v>:ak%"ScZd0�$2O4���O`�D�O��D�Oh�?a����P)���%N�1	�����Ɵ�	�hڴ�j��'�?����;&9 â	"���S��3{������x2�'v�O>�I��i+�����w�R/r��C�YQ�z��B�_}�R�K{�IUy�O��'tK?J�镊¥`����u���'��I��M�Q���d�O��'V���ua�`t�:�I�?i��u�'[�ğ��I���S�4I��Ӱ�k�'�%�6HKr�"g�ԩ������O� �?u)1�$ˊ}���3V���;�%�f ���'mB�'y��OH���Móh!tTL�F)�J���#!H�|�NZ/O��%�	fy��p��#pUc�:��U �80�V-iv�����Z۴�ة��4����9����'��S/Ns�PC߉Ch \ �@��6��}yb�'��'�b�' �S>j�C�"�\,��*.���xY,<�nZ�^$��꟤��b�'�?�;PX)�ɏ��5#�
��7�i>67�g��֧�OTlP��i����o
���KKd'�Q#��\���A�����!�B�O���|���yȤ���F�N�⭹��S&4�v�����?y��?�*O�eo�S�Ԍ�	֟��I!#,e���@��
�2p�P�s#��?q�O(��f�J$��1�A�!vÔ=K�T(��08d9?Q�B)=�~��t��E�'0�j�$��?��ٴ�FĈ�=mpR��M��?����?q���?i��i�ONbf�� !���z$P Lp,rR`�O<@m�>[����Ο���F�Ӽ���Q��lU��m@�Mحz���<�r�iҺ7mæ�	s���e�'�`Ye�B�?a*"�ʿ#h*5#��:<vuځ�A�T#�'�i>�	���	۟<�ɷz��A�@�?V�ش�5!|�N��'��7-�'@��$�O���>�i�OX]b� r_���e��B?�9��<A���?YƜx����5w!�͡�nH"%FA+��ۼ"��ɒR+���]�QEջ��9�ԓO˓8�8�@�W rE�RVog,�����?���?���|�)O��nڧE�\���2� �d  �P[#�Ӝ�$��	��8�?�O���d��pl�%I�Р��И|�l4�f�E�Bl$9UJϦi�'
�$R�?Q�}���P�H�s�ҖJRz1q#�_SwP���?����?Y��?����Of�p����YNVHq��J2e)�Zٟ��Iџڴ`��D3+O��� �DѶ�D*W�ߣ:�QQ�HH%he'�8�����!H���mZ[~�h[�����李p�f`�Ug^�>���Z��̟�'�|�X���՟����D�D�G�=,��c"T/4B�43v����l�	by2�r�A���O�$�O��'j�z�xw�]-y���MY)�T��'i��M�g�i��O��H�eꎎO�bAx��!,�}�t�=�ʴ�4�-?ͧt$���P���*xU#�-

�V�H�KR�؍k��?y��?A�S�'��Fަ�p�[�}��Ѣ�7]@�D��9���<��p����O�űG�55�J���D4`�B�ODQoi��m�s~������Sc��H34���ǐ�Y�Tѩf�ȦG��D�<Y��?���?����?�˟�hE�V��.����̫x=���AbӨ��#��<���䧎?1�Ӽ�A�-"���֌I,A�=�tO	��?!�eω����'��$��o�F<O�;� �%+]���3�6X�~��b0O�\2ЅY��?���'��<ͧ�?�`.��Q	�5�� ���(H%��?�?�cυ��?����?a��LZ�.I . ���O��i��|��ޑx��9YW��DY����D8?���Mk`�x��@7����B�R�nX������y��'�*u�V'D�=�8݊�O��I��?�]
��_�M���&gV��)i� �'m��'���ǟ�H��5l�v1蠏J%h]�< u@�̟<[�4n�U�,OH�9�i�Ia���Vq���yZİA冡��lZ%�M��i�@���i��O�s'�+�j�LĒi��E%�	�Ԗ8z�T�2�|�V��S��`��ݟ4�	ϟ(3��K7GIFqA]�Z������}y���*���O��$�O�����dD[��	K�#G �����Y�dp��?y�4cSɧ�'q\}����i*P�0�J��N'0 B���1��'�N�BT�ş�!#�|Y�@3�]�t�Q�D'C.PZd�F��I�� �I��Dybil�:	XVc�O$Ͱqi�
e-T�0ʔw�\�`�O�$4�	f~"�'Ǜ�)f���U��ou@���C�"o�P%Ǝ�H�7-5?Y�`;<Et�i;���iʐ)I�.�j��w)F_�h��z�`��� ��ퟌ�IڟH���b�#�P�#�̅���
�3�?A��?1�i�رi�O)R�'%�'c�A��̆9�PHRX�rU6Oj�2��ֿ�\��\ǖ�n�w~�7KKv���R1U^t(j��I6J�f�C���ꟴS��|�W���$�	ҟ(��WrS���!+D�.�� t����p�I@y��z��z���O���Or�',e�AHЍav�0�!M/H��'X剞�M��iE�D ���_����n�͎I�gA��)��/7������ˁr�i>��՟4�0�|�i�i�,QH݃xK��W"]6w���'�2�'e��tU�Bߴ
>�M0o�I匁3#�J��Dkt���?���?���V�����0#�7x��%�5e`�x�	1�M��ʞ��M;�O����<��J?� �%@Ü�?�|��+	��X��6O���?��?����?�����I�,�$d;��a�F`���NRx�o��)z���ɟ��	I�ɟ��i�����)T��ҁg�V�����(�	��Şk�i��4�yr	]�e�:9q$��C�b	��\%�y⮓GrLD�ɑ��'v�i>-�I�3R 	jgꝧN� 2�S�^�b���p�	�P�'�|7݅/g>�$�O��3O�d<�!E����w�N��?��O���d���&�,2��J�]��`��9j��dj(?�"�S;I��c�i�g�'A´���'�?	�T/,���Ƿa�&]J%V�?����?	��?��I�O����X�h`򂎎��\@�e�Oftm��I\ܕ'�b�4�|%;3�.f��E���2�::"�Oj��x��mZ�'��ul�O~rL�L		���q�ViX�B@���yG�Hnm"D�|W��͟ �	۟��I�l�@�4,U2L�3#O�w��0� �WyҠe�b�����O��$�O4�������>�<�� N&A�ؕ�4��*\�ʓ�?a�h����O1�F^�~�*�84'?%�5�s�N)"��1�OL�� �?IB6�d�<s�PI@�pp�Z�y�������?����?q���?ͧ���ň��؟dZ��qn�Y7.�*�¸s��柌��[����զ�a޴I�����'LN=��h_�
�ҕp�B�=1�y�u�iL��.
-�@S�Oq���N�:�F�sE��t=�V���<m�D�O��D�O��D�O�'���~K
9�(�\��X�%}���I��	 �M�G�|Z��?AL>!)�t���,��X�U 8F��'�z7�����o;�lo~(R�3.v��f�LfO�|rRg��~B�6��)h���`��'t��͟�]NR��?A�Rp��mU������˥,]���%�H���?��B�@z�����ɔ����<]�Z�ZѬ�g�l��O�1�b�	ǟt����d��ğ�Jٴ\1&$	(���$˩d���'M� @�h�&�{u��t�]")��(ԓ�(��EW����B�'zU�gi�e�ێdɎR�#�1�?q��?���?i4GŧDǌ5X��?��2����j�)"����&�@S!R�T���O���3���զ���	^���I�!��[�O=���"���Bk�˟�Jߴ
�� ߴ�y�'��9��Ǡ:M ��O ����ܼ?Θ����i�"O���%!W%=,�A+x���B"O����a�#Czhk�����%xR���l�t!��h�MQw*]�1��q�@c�)W#*�+7��c��Ÿ��� ���d���h03@AT�2l��#�m�x��q�@	4 l���0�N�)����8�s�BS�.T�\�0o�l��Zt�C�2�㕮X�"�p�[�6r�C�-%�5�v��)�2��%-�#lC�T��CK�'B�ҍˢdY�",v�`dB�0��	�4�߽:f�����Q|^d��I�-^�m#g^�6&U �fG�PF�P�0j�qIB��ee����u�%e��N��ץ����ގ�J��	��&P�'�Fn��) l[�Nz�\j�ΉJ��ɀ�}��I2D�8��^�qO\����چ5٦�{5D��B5ʍ�R��[��U�)�S�,-D���p��*�D]S3B.
p��iFA+D��$��\M�9ѐ&Ւz��hQ�*D�DĬ�1IǞp஖�9�yQ�-3D�X�������X�!n�3%�8Z�
-D��Q��D�	w�H�K��� "%?D���V�H+DA�`��M�l��.>D��*� _/i�E��&H�5o�(��<D����k9[�i�c�ӹ55&<���?D�����&d�:�*�HR��-!r�!D����,B�HHY�M?9�έ[BJ:T���D��P��h���^02���PU"O"��@I�|f,���܊330@"O���'!,~�Z�dG�[2$p1"O %c�bY�[��$����/>�:!�b"O�ѱd�0i���uR�c��t`@"O���
S5�2d��m���c�"Of�)�,�/|x��`ކQ���p"O���s���d�xdE^.w����"O~Y�c$C�EPj���@E�>`(pB�"O��#F��>��}�7 ^S^���u"O���ۃ}�	hQ�߉g��I�'���q��EV^,��L
3�
��'YƘ��	�f�J�C���3��99�'���ao�5K��j5��1��};
�'� $��c�m� ʁHȗx��\�	�'bB�8��=�����4:G��	��� ��h��HN.��#�<Zd��5"O�x��%��2�Y���4_WT��w"Oh0�!U�H>��gGD�ei��H`"O|�A�lS1'�"�
�H-ޑ�"O���*�vq��Q���:�x�f"O��(��8J�q�$��@(�x@�"OTԋ��Y$O�\T?~�x4`c"Oȋ���F�a��k߶y��3�"O�٨7As����
�F�*Ò"O�E�¢�:P��;JI+*�n�Ђ"OX\Xo� c*lT	C� v T�X"O��DN�E"RX�@mZ=.���2"Ob<a�υ� z�1Į�8�:�'"O:M�@,�J�ӂ���̠��"O�Xi�F��B�l!6�E�1���e"OZ5�2� v�8�B#2z����"O�[�
�Ky.���C�5*�,R�"O���!a��Z�u��	6B"ObEzClʩf�T8RLJ�$]�5"O8�z�F� j���re-͉4�ƥ0"O���k�M؂x�5�K�Z��!�"O�dA�MEL[�M�"���zz���"O�x7�߭ �ƱY�i��9`��`"ORx*p�BLl��
��k���b4"O�mbw�5�>d[���9�N�Y&"O�$���^�l#K��8�i�Q"O����G�e�Iа���u�Z �"O4x���[��ؠ��L��,a´"OΙ��Id�P���;O)`=�"O�=�f��R����	O�V�
��"O�]j�G֊<�X��-"����"O"����0|(@ F\"䠀%"OI�ѥ�8\p9!vcܦJ6��s�"O�)�K�%J�RL�B�,nX��"O��â����'O�Jx8f"D���`�3��H�G*̫q�(���>D�����G"[S�q�`$ʾ,E@q2B;D��c� n�
�C#��31���P�D8D���#M���܋�B�U����N!D��a�)f�����L5Z�e��!D�|��.B%<��S�ꈬx�0���=D��Se��#"�mCq�2�V�68D��2�(A	O{�|����;c����C)D�1���`X�ܙ�b��Hж�z!�4D�L�LF����3eE<i�ޝ��.D��!�A>F5��I�-W�{��)C+D��97��=	�N�(ᓛQ�D�҈6D��P��M�o�lBfH]�A��
�5D�haT�M�?�6��3`��7p ���3D��X	�"�f̣���:Y�څ;�n3D�h`ۼYqd��2(Ŭv�Z���TJ�<A���.
-��Y�H1$5Vy��l�O�<�'�q�^�AU�ޭDÀ��ML�<�MA�

t��&9�1���H�<��ꇧÈ� �*K%���#�
i�<Q��M3��*v��4{z1�Q�]f�<Q�m�t�� 5�����P� �^Y�<�wJ�2hX�"�Tk�d%�T-^V�<����J4�A�7��3aD�ٺ$�y�<9���`�ly1���� �
��u�<C��qt�SuU> d�X�PLk�<���9M���[�|�P�Q��_q�<��	�rÌ1��6z���Q��EU�<IǦێ^�&�X6!�-���p��O�<� T�JB'X�+^��dQ�,I�@r�"O.MA�L�E�0h�� IH8Ĵi"O> ;�k�<7s �S�E
�C$- �"O�ёG�>{��a�v�Ȋ�*ܛ0"O��ڰ�8w��qa��[6CےA�w"O�]p�"[�_Yl�2�bH
^��"O��1�ϨGR$��@�E�)�����"O���"�txF�Q+ݍx���"O�ԛ��^_�jƇ��J00r@"O` !�:obzyr� е+D)��"O��#�-A+dA���nF
W�-��"O���W���qF����mh| �"O��x%OQ,;��m�AI�P�j�"OLI���}P1B��\�2E��)"O�e#����vp ���� V)�es"O�$��%�%v���Iط}z�X�"O\�i1g��&l�����^�@ȁ"Ox�B���b��Q[�w�b5:�*O��(�@&�j`J�rKx��'z9�G
�*���yg(�;�9��'��mIc˚ |�\�f���5�؊�'���P��L.��G�<����ȓh>��J�фG� ,�7-<�<�ȓC�Z�@���'?� �q־T��ȓ}U8AW�4�J}�2�S7$�2d�ȓx	���_��D�����H��؅ȓ\wvQ���ϰ�6(��'<[�N,�ȓI� S�����9@d���ɇ�^�,�3/�;B�,�Ӥh 
sHR�ȓL�� H���4f`X07ꑃlA^��ȓvn���� �gȄ�f�ת���D$����L�_�`)�B�t��%�ȓ9O�����ߠi�����Z�K�Ĭ��~�nժ�Ő�DY2��ğ1w��ȓv��Ps�!�ɺ�/	!�|��E��j%�΋{�j�``��G@Q�?�@3,O�pr���U(C~�ҽ�On�+�B�'
��'�	�R�%1�d��B�tB��+Ho���h���ܨ�G<3����$�$���<��BOf
ze���q!�X�<i6dW�L�̐�MO,K���i��TL�I)j��?�}����^�<]c���bDnA�҉�F�<AQ��3Q2$aH"��$.��g�[�A�|�q���2W ��v���x�"_7C����Ɠ 2� [��ͬaP���ώ�b�Tma$��e����ܪ-���sA�F�e�4�EN3Ű<��ν�J&�(:��2t+�M@HL:m��-D��{c��5_��pc�v�����7�x,�4A�{����C�z����Ls��Z4)Ö�y"�-��d9�K+f��X"l4��' 	�9OVQ��̘*h<l�x�ҀzBO�0�F䓦/����BC�$~���4G��h��C���0�Aǎs������9h-8U�剾}'
��=�ͪ>F����K�*n� Ӕ�j�<)�'�����&�;p����Q�I� j0�}��D�]����Z�p�2��fdɍ�yR��l亡I�#c���P����'��U03�3O��s�̈́^�5(��H���rO�q�O��`�2�~�����a�2�pu��~��8HFM�`�ej��\�b������>PqO>��qK��А%
��8;%���y��"c����S��Д�й�yү�v&!�s��97IB���C1�y�,Ҡ}�P���ɩ6K���OL��y
� <���V������4��KC"OB�bاjiX�pA��cP�� �"O �2%B�5r��1���AG�g"O�eiv@�6�ptr��ܼ55l%��"O�!��/�$l�� ړ$Zu�"O,�Br��9gL7��-hv[�"O� `͙�I��5gX�nHJ�!�"OZ�i�   �l �eO�%���"O���DGۂn:2���$H�V	��"O���o���D�n�"O�,a�[=p՜�����"H��"OR�� �Ɏ�J�(v��cҤ��u"O��� ���H�i�����"Ot��V�s!�MbvkU��Xб"OV|� ��!O��e��D�/_Ў<y6"O*%���Tff��W$;�J9$"Ol)ҕ@C)WM(1QS"	�+��{""O���T��$$ \��?�<��q"O|�36/�w�T���*s��R4"O�
�DV����1��ܘ!��)�"O* @A��-N�&���@�4AiR�3�"O.�
/����oB�b7�4Ya"OD1� ,�&OXi+�O��d̰و%"O�5���#+�r�;�Q�t�<�3�"O6H�及,Y#Bݲf����+#"O6�[�%�7Z
$#��
=;�i��"O��x�`�8@֐�1�M�/����"O�uj�/�SGl��e��>fp"O�]R��"fCꙑ�dݫz�:��4"OIHB�ޝ7v~���T{211�"OJ�{#��=����Ꮽ/�H��"O��8f��p0ѣOC�*���Y"ObtH�-V��y��ْ>�:��A"O0l�Î
 ǌ�:TÂ\��X�"O�����
��
_)tX�Cϛ��yr�3�%�6㟎W�8TSoV��y��O(c|�[a)S<xk`����6�yb�
-?��!5��s��u*a-G��y2f� bQ��G�L�p?��p��!�yb�	�@��i�P5p.�H��,��y��R<}(����7n�(��+���y�.N�=<e�wC�z�n!��ق�y��5�0i�@�qז4��!�y��V5jf$!5�S�\.�PgW+�y"`\�o@X	!�Y���!���]��yJ�>��MhT�Չ0��u*��<�y��\!����4.��)�� ��ϛ�y"@I�W��q�bַ�^������y��Ж	�f����R ӄ�L��yr�K%���@B�l�T��G<�yr��<< |���b ��.H��O�y����푅K%f8���eլ�yO��n��(b��>uU��c2�M&�ybeD ;h���� 8mJ��$&��y����V;�lC#KZ!d.��3���y������!	�0,-��Ϟ�yBH͌=bT�)�F"���v��(�y�Lنi�uB���/W�m!����y���X���#$G*f��`V�y��3=�}h���(�jZ��4�y$�*�v��B�I5�VL���@��yR��"a�x������)���1-���y2M�
N� `�o�+*r����J��yGQ�G<Z�J��Z8��0���y
� ����O!o��ia*̜0��]�"OJ��A⒞Yx��B	ʿf�<�"OT,�卐.6��=���Qhd�3�"O�J7O� _�\z��ƭSMV-9 "O��b 1 �z��'c�r�J�"O�X�ǫ�|��MRv�],	�\,i0"O�	�׉%�Vx�7���">lġ"O�a�dF1CP<� !��"~���"O"��F�"�.d��۵f���0"OHd�w� |G����Ȝ�^��,*"OB�A�C_��\-١�Fo�^l��"O4���046bU�7�C�%چ��Q"O(Y�q�H �д`#GL�r�F�V"ON ჈H�h�6H]�.�Z��"O�D��d��>ˤ�ё;�&�q�"ON̨3"�5BP�av썥�\��"O
�Ђ��s�i�Z0y��h�4"O�0�ШyQf��#t���"O*}2��K�i��()�
�^Ҕ��"O$�ʄ
h�����ϲ4Il[�"O� �C�>,]bt
�#Z0ٰ"O��k��$5����k��a6���"Oة�����c�Ԕ�𫕺&=ʵ�""OT,�Q��0���n6�щ�"O\��4�ȼHQ~)�@bҜc6()�"O�����D�*�BG>;
�+r"Oj`���v�x1i�ҰB$(�;`"O�1p����j8"5��87�e�"O~���Ži@������:/��a"OV{DO	W�b�F�8or�`�"ON�c˓N��ūs�F�
x��"O�Q3R��3n��č�x���"O��u �&n�����E�و1��"O
�#�L�D�R9�o�3���h�"O��C��I!Yl\���Ң!��\(�"O<w��o+Hy��R�
�^t
b"O8�Q0��+6칀\.�1�*O��*��X|�-�@F�;N�{�'p�eXd�Ҏs�!���1�� J
�'J������|���Ө<�V�	�'r�x�cG�X�� #���0�h���'jtA��P!�"	�Um�"��e��':���ញ$X����lU2���;	�',|��7�M�5b$8���'��-A���V�U�� �6kJ����'�eNN9YV�AEB���,��'�ֹ���|!���b-޲�i�'vص3%�hǤ���6h{�l��'m����숩 p��QŌ�3dF��	�'��� c�J�i����>`�f��
�''�R3AC�� i�@�+� ���'5� h�GHP��E�N�v�l��
�'��A�&eά"4�Q�9�D��
�'�V �$�
�V����/�&aP
�'E���K�t&�X�ҍ�>!v���'f���N�A�B9��'M�2�[�':�u�v��/r~������?HX���'v���		�A��4��[ NeJ1��'���p�܆Հ�)�i�G�0!j�'{\�I�O�<bߪ�ۇf�1G�!��'�8d��J��4>��W�8�R�'��<qG� jˀ�PE�L>Q5j\�
�'@�	�t !g� ���D�#af9�	�'�.e�S�Yhֺ���(��Q��H
��� (܀w���H�ք+8�`U�"O��3H��8HI���g��+r"O��p�SgC�EQ���}~����"Ot9� �݊!9@��ra��\$��a"O"�c�J1���P��3@tlJ�"O�	����0dj����20�Ձ"O��IR�Z<xB��o����c"O4�#D�0V(��㊤M�h���"OҨӂ�U]�F��b��b�~�(�"OdT��!�b�R���[��\@�"O��4Cbp�3'��2?{���ȓ���2�)ȩB�FX93(��-Hz���t����F�0m
��8e�@�n�6���h9����i����u�uS-r��ȓ2�8���Aĉ%r�h��8d��.@�ه��Z�ҁrQES�K�Ḋȓݰ�*�	N�O��0��0_�`��ȓ��u�w��'l9����* ���$�ȓE�=�@��>^��b�ɰ��`��OD}`�I�O��Q��%?�|�ȓj�-Ζ)�vɠ&
34�H��3��Ti���6=��b�`ės}�̅�Nk�����I���		Ɛv���I� 1)���+q��r�A���Ą�L�n��F�!+,��� P�Ȇ�q�Ȉ��CŀXƐ�g6+�̘�ȓDF��:�4g�U�1H�0,6�ɆȓK�4#��:VI��wCҮ7r���f$�]j��-�n�R$�R�d��͇ȓT\m��8~d��BT�H�0�ȓZ-�	�Bj�/C�X'+Ř`���ȓ��}�P�!Nr�J���6�v��ȓUl�����4^Ȣ���K܆�ɇȓ�m�ᮇ�<�6h�%�+Ha�|���6��j��Dٞ��7��d�4$��5:� aPV?@�a�C�
$O:�ȆȓD� %p�&X�6NZ�0C�;Q�Zp��4�fܫoܲd=��l�
m��U#�'�hd�!bN9Q1��<���',lD�p�U9p���qR��zȉ�'t�q���V�����P�{�z�9�'>�#%�R�5�xā��={�����'ي�bTD�c�=���r�\q�'�R�����-)�P�)�唝t,
���'����F�]80�6�s
��e><Q`�'Z�!��_(`i
���eA5]x���'�N���U�(G�P�B��[���

�'n��u�^8&8��eT�h���'� $�q�����o8f�X�'��X��Q8x�~[�.h�PQ��'"`Y�N��v;K��U�غ�B�j�<iq(0x�R��&�z7@���_l�<�g�����tꏀdօ�D�WP�<ipa�?z�z�*�댹�8XB�V�<Y�씘4ĭ"���5a�8
� ZU�<�'�H/Y����ώ.%�b���O�<A�D2�����OձQ��M��B�<�q̄�FMbq�w�\�����FG�<���(\��@�J���9U�ߖ%!�$ūf��@M�%g��B�c݇>�!�$���Uc��M5~6��R�e�3t�!�C�Mz�$���ͽ(�\�+���!�D�m2l�;ԆM;Ant��©�?!�X<<�d����֏kc�8ȕ�^+�!�� ��VFL!�؄i��L�}Yv��"O�\Cr
���ɂ�DYH�����"O�@�$������&C>#�0<��'�x�3t�_�5?�II��T�]Z ���'�A9�^7���Ջ��j`q�'ΘYS� _�(y�#���x�6@�'6�bt��9X�2(�L�i���
�'f�m��h�>��BC_�3j��;�'�l�;p�<Rj�Dx���C<���'g~@�T���s�$�:��<��89	�'������|z��V
a`�%8�'yPh��L,tmNɻB�L1�J���'� �h6�4���2)C�3�8!��'F�a9�ҟE�x�VJG��iI�',J�$傴L+q��J�,D8���'*N�n	��!�\!��C��0��'�i�J�-��}�^�O�0j�'�% W�V0W˦���
ǐM�p��'����%e:��d��Lpr���'����-/�@	���R�KU����'�� ��FS��i�R�D�q��'&c�!�)U&��g�/@̙֔�'�
%kԏ֦/a�Y��6���2�'��Aԧ$g}@�8�ߤ;F���'.X�� ȝKkf�3�C��$��'��(�蔤!���C� �#F@}k	�'�J��+I I��\µJ�7;�����'�Ω�0B-0t�����<�HU)�'���;㋕�¨��M\̩[§���yreߎc�P�k��L�<
�ؼ�ya/x�|9 �nޖ<�D�0��ǯ�yr�4�V͘�)�$?H`��y�]8$`.�8�fΠ_U��[��>�y�%�qh����0FHeivɞ�y2B+���խ�7���� _��y2aL�U"p�c���+Ln�ڣ��y2��D��(�[�*��M����y�k�G; 4�a(��(k<��C
,�y�%��~X��0��j����QJ�yR�@�`���3vc�j�:��I���yB�ؔ>[� �A牝Z>�������y�(P��@��CR�X�D@����y����J���s$� �X�ẻ��y��Vq�$��B�6u����dë�yr]�����OJ�W���/���y�	��r?p<e��%(���M��y��yK�@:g�Y���}�a%�-�yR�-$y �$����q�&
��y"��i�rh��j��A2y+���5�ymF9d��*Dr�vYs�#O�y�h��[��� �V'l�D�ٴ�ӑ�yc�oT�yXE��%j�,��D����y��@�_4Hp�L�c/0K�j�	�y�� �%`�jA[t>T�����y��� �F�bs�P7B����bgʗ�y�*�[)* �Kʆ�3gj�/�!�d݄Rh~��0w$�Y��Z�!�Ă >�cb�W6kl�X�P�Y�!�D�/�\	�R��-`�y:deC�P�!�$�*}�$��%� uu$��I5P�!�$S1jd>� w�Y��P�"�ڧ�!�d�"a� ӣ��7�2B���!��N!�#$ �t}��St���q�!��[?�>}��e��(zD����:cT!�� �c��A�k�dUp�I��A��A"OT�Kҗc+&�Õ�=-լ���"ODLـ`��0܄��g�H%nFlB"O.���ܓGH�0��pZ���"O�� �t�5sS��H����"OL�ٰ*F� ��Es����)�t�"OV��M
�a`6�)¬C�l��I""O0��a�m���J��?ݶ��""O�Z���Ű7����4�NZ{!�D׾#�=)��e>� ӊ�Dg!�ĝ	_f�����D��E��^�J�!�dT1<�-z�.@A'�ȶf�!�D��1�Z��Z� pK���3�!��`,����!,|ZfO?5�!�D�7���.tX���v&�)I�"O�ث��K�.�q!s�H�( �;�"Oū�h	8�5K�!P���q"Op,��̚�{
���Ə&x�Bqy%"O�h2B�5�E`B"���bi�"O¬�s��(�������{�"O*�s�P5D�����:m��4�q"O`!;�ʑ�h{��s�� 9�"O
���H!}I �wc�$F+!��
~��<f:����W�g�!���8D����#REYԂ�8�!�d�*!��|�J�Yg>2�S	dU!�D_�"�@�b�I4Y2Ĕ�"�L0!�D̗ �	���ۃ^�,�ۗ�҇i!�D��IzaF+K�e;��^�N!�d�iR��SdE�lhnqoA�pV!��4A�fH)E�4?^4���9_C!�DQ3x�:`�iE��˒��+a�!�Ā�zz��ü3[.��PV�ԊZn!��خ!���J�<5lD����>h!�$F$�21Q��$G���ڳlÏd!�$ �9K� � P2A���R6
�!�D�,T�T(���í���C�-	�N�!�ݹi.T�W�y�NP��l��.�!��B�x,(�KL)�hE�S�X4Q!��7f1�E����q'<�@�^*6R!�81$Z5�Ṗ0~�b Y#>L!�d<_x�˖,�9m�U��6F�!�$��)g�E�Q��<hj�A�� �!�$F2<���dH,��d��7-!!�D�_�m�P'Ӱp���aa��!�$JW�Q�s'�����%R�!򄉿~��`��F�2"�R ��!�ݒ42�T�@W����c��LM!�V�:$(`*]9&z@����:L!��G
>7(1r0�Ѩ����H7:<!�Ƽ��� 1�H8�bV��""!�䓁b(���'g��G���H��"!�G'
�<h��̇�ް����M�j�!��#j>� �B/ۃ}FYٖ�_�j�!��ɴ;X�G��<Ci��h%�^�6�!�3n(�b��ΨUJp IWG��Py"␽T��t*ŋ�$=*�&ߋ�y��H��L�ڤ�Ϥ^�(��T �yb˓+k�Ւw��'�n��N��y���u:���w��`Hb�R��y� @3�
\�CL�3Yv�〉̦�yRC�'D��A;����ـ`�L��y���#VZQ�is�p��W!�$�T1�T��oT`r���e��!�� Ȉ��㇈Q0Ҽ@�K�*
D�t��"O�X��*�&�d|����8)��kw"OJ��ϑk A�˘�=�9�"O^�u��3�RH��i�(9Mb�r"O|�y"1q����/W�?��"T"O�����}�n���58 61j�"OV5�I��k�*M`���.�kc"O���`��F�b%��.�:hp��
@"O�M�'	-"��+f��7CzF��7"O~�"��96�G�oj�%��"OH%��n�fM���(NP@�S"O�i��֓~�u�U�^�Oh�|� "Oz()da��-��X��Ң5`\��"O
��E �f���ц����"Ov�#��PPd��SJ��zS�"O�����X���1z�ƈ�zIB"O���$Ⱦ{v���v�Z�L�2"O>�Q���5�6�'��e��"O � �һb�t@�1�V\��"O������r�j����HR*��"O��i3HX�_����b��jE�isU"O�<��R�ʚA�`�!)�䙆"O�H������Z�����I�"O4	�P�� qč*#�I��ɢ�y҈��<H���$Tgn�!�M6�yN;DCҠ�R�W�A���)1I4�y�
�e$�	���7��L� Hͤ�y�d˫~2�i6��,)�`� )��y���Y�:%�2��P�`�PG��y��ٜfP3�ܹIp�㖌U>�y�_�*�"���B��"N߰\�`P��Y_�(r��Ƚ^_h�MO�"1�ȓe��[���Q}^D3����Q��ȓs�bܑ#MKed<��V�$`���[��`�v풓S�н"+Êc~@4�ȓ?���w�O>5R b�
.��ȓdf0� ��#���W	+���4�������g��"�"�\ �ȓ]�����!�?V���˃k�.��������k�	;�%Q�AS�Sb܄ȓZ\�ɸ��[�l$�MH�B!:�R��ȓCSإZ�!�~xݳ�B6T���ȓ_�1'��009IR_�2��Ʌȓc�����O����w:-��x��p�H5p���V���`	�Q@��e E�V`#|Qa�K��ȓLIF�#R�[
m�0�@����݇�@�PK�������
uG��q�"��ȓk?�Y��-ź�>)�s�F�[PZ���m��4��
�5k�,�a�L�[���C�"�y�W�R�y��N�d��<��BN�%�'m L�f$*4��%e��ل�k�4\CWa�7�A��%O$.M4y��RW�XxS煵c�I�!gK!H�T�ȓM)�\�CL�N}�4��Xr`��	�"�7.J	.<H�GY�U�8���&�}+����bQ�IC� ہ\�H���jO�seܲ�XE�vi�8�^1�ȓ1j�Z���x7h����1������� �@�H	*#�	�2
D(j����p�� !�*HKn(s�J=W2�<�ȓ=��H���H�dph95��?J+
y��d� 4�S�7߈Aɗ�;�z��ȓ%�T
����lP��V�j�����S�?  :!�E�<x���*�3��Y"�"Ot��"�������c�'
] �2�"O�@�O�8<xUC��;T��F"O�)x�N
`�a���8͑�"O�ѓ3�>I*��[��5��< !"O�ݫ����eބ\kE��/,HA[�"O���OV�s; 5�FI���\�"Od�QA
�e��gF(9r$"O���Jۮ/�(Pr�'_�mB ��"O|MpDE�l��f�!N�#"O�i���W�kr�Y����>��I[%"Or%Z�,2cx��W�Dzeᘍ�y�@�:l3�d�U�F� �"��T�]��y"��"� EHĉ�8v[U��䝳�y�ʈ*��J�I?l�2��bQ����hO���<�ňٯ����I�2W��q
�@�<	"%�:#Z�ԲD�ê,W
`*c�<	!ܦ?�6 ˶�L*PL0LCԈK�<�a�-�6��6��Sþ�`��p�<	nR�<��9�E��v&�P֤_o�<A�� ;�JA:��.-���Gk�<yf�!����-dN֬)��e�<�4�x� �B�U�~��E�Id�<��Ā�g#R	4 ��h��y!lZJ�<ɶR�7{HT1�J�o88���D�<�&E�b�\<y��PH��D���<�䄝�d��=��ɋ�v�� �#O}�<Y�D��d(�YU��1���p�KFA�<�2gΜ(X�@���-)�!r��F�<��R�0��@�#�'W
yX��VB�<!`
;^�x�� V��Ś��e�<���0i��gʃi��Ē�*�l�<�e��WtݑCL�d:Fb�e�<)fj�,A.5��mF�W��t��b�<a�ɥ[811��=�"<+���^�<�5� &�\kQ@H�A(Nqp�D�<q^zH�bv#̵U���ó�F�2B��"K��1�f�9rc�$Tč�VOTC�?����/Z������%���Yh<y�ՐnP�up"�^�gDu����\�<�G%HC�l���N�a�F�@���^�<I� ��1=��q�鏇_'Np����Z�<��Ӊ{�fC���w��y�f�\�<i@�@"b8����ʆP-nU�cE[�<)���w�@a��*�7�N̉�.�T�<�".�9�pU���{��Q�͎U�<qv�^�@�h]As�.�l�h�L�<��"%&C�eL�V��h1�I$D��1w쐏`t�-��A];)�8�Ej%D��"W��Vmr(� D�&*�̑�o#D���`�ϴMF���$U?zθG�?D�4�1�8e(��[@AD{�8���;D�Hz5(H�)=���B��*v(3�,/D������	9Rs��O�{TH�Ņ!D�,�E�BH���/Μ=T�*"D�(`2 ����)Fi�q����M*D��!�m��6�j�G
�
C ]xV(�O.�C��zC"�l���K��	EQ~e�ȓ]���JR��?>R ��Im �ȓ0�)9�jϡ%�2	� ՅFܔ�������ö1��yҔ
X>S�����s��D���ŧV�,�KE��^��}��-��DaōN}*�KЬ�i���ȓrU��3�M�p+��#�I�tm䀆�S�? ��
�!$�n�
���1C`0Qw"O�(����9�>ѫP���[a��(v"Or���.}��tZ!J<ZHr���"O�S�J������$�?#\�H�"O�����p3�4`��v'n��c"O�Up$LF4��<h �_�;3����"On��c���	�`�A���i+�d�'>b��;\� �!��{�a�D�O�h�p��ȓ2�2�����,�n`���=a����{k����!��Dm�%��Y�Av݇ȓ.��Q�v.��Js��Bƒ���ȓfe�,�`ΘB_ XZdd��ˢ���1��m����3 �0r�66�� �ȓ=��!�D�<� ЂAU�T;$���П�'��D��'d����+��q,a+��=�$���'F���n�+�*1qF�e3�I��'�c�Y�$61�D�LX ����']���T�_��*�E���y2�]F��ȓ��A�@AD`���yR��
3�f��1���$�lt��jS��y�CK/_�@�ʃW'0������G)�yB���R�Խ��-P%&��e�2ꈼ�y��)G��|(&៫%=��3�Q��y�!ħ#�BL:G��I�Ԥ�Ƙ7�y�˛�h��C.I<<9��
�
�y"�,m�fYId$�l�X�C�ݓ�y��O�f���)%j��Q��J�y�C&g2�y`��<75� I����y«�D��pS��!L̍��+��yÓ=Ҧ�CB� .� �ή�y��7P����ՆpR t�GG��y"��	�]�������OP2�y�!�h1��ţ��p���ǋ�5�yN��[� CG��sz5	��y���6�V����@('��91�]�y�$$�j�;1+r�ub5��<�y�b
��5z�&Jm99��\��y©æZ�J�[�Z�d�\y1��ُ�y⧓�N��9��e��I���qD()�y�'ҹz�V�z#k�42V��9%Ɛ�yb�7�؍���5\\XQĢL��y�.��/*@hJ�l�9M�
��yR`��5t��I�3=�t���U�y�O�d��z�I�ľ};f�\2�y���7EI�����M�P*�yb`܆]`�BjW�Ύě"�J��y"�� 7���a� �5���9�y2/���q�T��<Y/.-VDɜ�yb�׫�J�̭Se�R婕#�y�E�<y&2	� 'U�L�X����yB���_��Ys�G��Qc���y2b]�g�T�K���9�)顯٥�yr����AQC��CXVa�A���y"a���XܓD�?��2��yb��S�8���ܷ'�rT����y�*ِa���qh��"��4�vk@)�y�LN7����DW�(6�*�y�چzt[7��:9�Y!&`� �y�,_(z���9��
.�p�P����y�M\�u��{Ƣ�)�����y"ņ���Ԓ�iŐkO�=���L��yBi��|�h�%%^�e������]�y2��wH9K�c_ /��1j���y2��|`�pR�71P��� ����y
� ��;���X���&K΋@��p�"O��)QO�t	�yz�iG>|�LqR"Ob���ɞ(o�ұ��(�$�j "OF��f���t$��Ǔ�F�:�I2"O2�K�f�WR����R�&���!�"O��:Aā�!v�3d�	E�.Ԩ#�'I��'��
���7f�B�1�I��`H�'nH��@^�t��5T
�53��a��'�v��5:H���ş(l4�!�'�8Az��Ț)^�5�2m��T-��s�'�ʝ0%*�}�6����/@O0���'\���c�q�S�M��4�L��'�^�Ɖ�-6= T	��1������?Y
�D�|Ys�Z�W@��q�n^�H���A,�pC#�J?*d�hG�O���ȓl��Bv�4�>�����~@����ް�RQ�P6l��'J�??���ȓ|L��x�&��<�9� �ɀv�x��ȓ:�(`2��ʦ	�.a9�e�>��ȓq�p���)��V��h��޾NIH��ȓĒ0 ��T�B� a�5ϲn���!��}iqiŰm�J�KP�E.��Q��,�p��gV�
�D��2O��;�4��-�:���C���������^��ȓad�X���_�v�kP�`x*��ȓJ$6u���\�$�nHo\���L��'H��q�.#A 2���|�N ��'{�<b��8��y�Wg�80�B�	?+�$�h�#�� ��a
±��C�I�}��I�d�R/bW�������DC�I�0:\35�!rx���
ܾ,i@C��.�q�AaH4�,"ai�1�^B�ɯs`�	(�I�s� ���Nػ~.rB�	�j��@���͐��t�󇙵q�|B�I+MX CG���,Hr!�p�U>B�I-��r+��P/�x4	�:��B�	-+8��𢎐D����>)P�B�I��!��%|r�
��B�f�RC�6`��hS`	�$U�� ӪG=�C�Y�h����
�u�bD;p�ۃa�&B�=yf�@rrƞ�gBjLc����JC�0l�a�&9?NdJUI�/) �C�	�A��X��FI�
r��xR��M�C����س�(E_3l���ܱr��C䉂 �X��7/P��� A��C�I4Q���fe�y�&���C�Z�C�	�Y1RA�7c�+pMX�w�ܗA�@C䉰F��EY`@��4Y��nЩ[��C�I�3֧?̶=p�
OxX�C�	�.�h;E�z���H�ΰ��C�	-yj�(GΓa�\s�96ؠC�I0&� X��  ��K���w��B�I�d��BF�ȸV�0�M5(	�B䉵!��i��K؃ ��Ti�h�c֦B��1[��d���&Ln<[t�Z��B���zi����p��e�'%�d3VB�I��NQ�cW�-g�-q%ġ+��B�I9kŒe!
1*¥YQ��N]�C�	�0�Vq�"�Z���\ ��3=v�C�I�B�,�*!��$��K�W�B�I�&(�4[��G"��଀8n�ȒO��=�}���2��ǌH�f��0��HV�<!��M�O5�<P��)�4�ub�O�<���1;x^P��f$�<�!`��K�<� X���a�4e���vG�,gČ�"OJ9����w��<��GM�\6V�i�"O>����R���i��ۮ|I1�g"O�%���$�:��6�̋;4���_��G{����Z����iF �����f�!�$ܦ@�v=Bum1>ɮ4hݽ<!��� Hz= ��V�TP�!��*�!�N6z�}�iG�^���u�O/)!�d]"O�I�Ѩ�s� ��/ԋ!���SX� �F/
���U�!��Y� hip'�����H ��'�ў�>�3�E�"$
���-Xd���5�?D�\'MS� ��'K�G���G�2D��S!/t�1" �n���E�;D�TR��?U"�y��^�#M$�I�N4D�����P�V�X�o�I��kq�$D� ����4G<i��J�
XSZ����,D�l8�AY�d=pay���5i������*D�H���ܒP倩�"i	��P��N=D� a!�/2d<�Y�ܼl���J�6D�D����%@���+�hL���(D�t"� H�L��&ưW�Z��w%D�(ð�:w��y��O}>!�#"D�X�H,v�"�2o��5e��6�-D���ħD./߮�B6�Q�&�ٷH,D���1"ޑn|�+ Đk��[�+-|O$�D2?�b�"8�|7$�Kεч
O�<a��=h��*�MռZ&^�!�$�M�<a�F��x{�h"c�:E!�g�D�<�E(?��i��H m���a4bY�<)��,Ly���
}
�d��T�<٣'�b�P�r�BYKF�"��_Q�<q��I��J�jZ�7Ϣ�"�I�O�')�Od�)��\�\�@|S��E�0����ȓr�j��/��G���jU�&x� �ȓb
�����[i���Bv'N�Q5,��<?>� �4p	�Թ�'�t�5��u��=@��ڦk2x% R�V�8)����`2�A���EvX�cU���\��v\t���HfN���M"AZ�'���Id��DUg����]�w�U=��a�5D���E��cYB�Q�+�M]�Iq+2D����)y85b��ԔW�֤��5D�H��EB�W78URD�l�b����4D�@;�,ԝfblQ˱� c,@�rA8D��*��V<��K#�ޘO�n�0 �<����
fT���ա�R�ҙ�Cغ[�<�=)Óa!8E�i�/� {�#��D��w��A`)b�"c��R����ȓ2�Xly��#�r��������y�BT�1I^�G�,��1�ֽː��ȓ{U@�W�EZ$u��F�h��!A�����R�;��4M.�F{���<��3XG�tq`��0{���3�^�<كG�i	Tݒ��U�:@m(�CW�<�G/����a��,ew�H&l�O�<A��įo��Z�����ț�A�<A�xK�@��C:�P�3��r�<q#BY�1�C7�ۄl3��"Gl�<������t<��O�>\�q�l쟠G{��ɞ	~�h����B\���E�F���C䉟I{^%���T�*����oD�k����0?�p`��itT��m
.fQ��h�<`"\+~�p�) o§LYJ�g�<� PM#��5�؀!�O���8G"O|��*	i����%%B��Xg"O�9�ת�C�pը�*�+><br"O�˓�ǅ4�F 3��yq��{'"O�|(��
0z�<D���Ӕ']l���"Or
�+���z��ǋ��W�<�""O����	�\jD%_�@D�p"OHrt.\2_J|�ˑ�py��4"O�Hyq�Z�*<���#��L~�#g"O& ���	Z� Ѩ$h -�R"O�<[���P�FP����H��1��"O�yQtbA�C��`���=[�Z2"Oe!îӊy20����̱<PBRS"O��+�ur\�ZCMK�a�U[�"O2���Ef�٢�J�`qQt"O�X��
-=d�%zw*�)&�xQ1�"O<ا&B�VP�Ǣޕ#�:�{p"O� �b-�<�$�r����:%"OdE��BV3Kh�h��a	������"OĀK4(U��@��&E�W��x��"O�y�Q��/kUD�	��G�#�4��"Ov�eFj�<���ގK�$| b"O�E�b�X�i�:r�i�{P��"O�9���R,WVl b�B]4^a��Ie"O\,rGQ�(�f�xᄖ8]�a"O�f�1J� ���Bi�F铷#�<��nnD0&NО,�DЧJ���|Ş<ó������a�-��ԅ�'}t!@�)�����gP){H}��V)��S��5P�+u�6 �`�ȓ�؉�g��zT`S""T)F�(��p�B���H�6
��*�bG)M]ƹ�ȓPSd
e�1^|��NĥVN �����!g��.�D�9D����8p�ȓw����M�"z�h`�P�]�!���NI�lSqA�8��If�в4!�D�����[�I6AVV��E�ӳ�!��1Z�*e��g���1�9�!��qÜ�ۢ!/�\����Y!�d�A�L�R@/Q�.%��	�m�!��V��:�"��w�lв��;�!���r�����ϴ�,�c��Z,�!�d!⺰;�L ���T	�M�!�DN*؜H�e�6>�@ȚVl��]I!�$G.$(@)v��79�Jy�#�BPQ�2�)�dk�B���#��W9O���C"B]!�y2����ɐ�Ј���Xt��{Ј��SH�UT��cf�愇ȓN�������M�X�d��0��D��P�H�Q2�	�u)���g�����8h>�aCM �p��ӡ[�$4��u.A����tw��(���7��?ɉ��~�ч�Kq,��$��4Ct�jՁ�D�< ��=:@i��+�0b���g�<� �]��2l"��_��P��u�g�<y�b܄K �P'�?O�1���b�<��"G�7]:i��:r|��J��QT�<	ã�9��T§B��Rx�����V�<I$/� v5�X�^�1��y��NQV�����n~�  Ӝ!V��'`��,�q͛��y����Tb@$���Đh��� ����y�bŨN���LȨ[�n0I��M�yb��VN ����҈E:�y�m���������"m�t�٥�y
� bȻ5!O��hԋ�g��E��|�F"ON�K��K�2�yr�Ha=08�e�F�����J~"��FҢp@�M�>�L� 
���yʛ ��1�°I��b��y��m�@-��.M6Hlԡ7Ő�y���t�ƀR�%�%=\�ؑ�W��yb�%�-R��Ҕ4Ѿ!�ai�=�y�AY;vI��S�cW���1���y¦�7	���#c�(<@`�/�y�͇^���
"���_��p�gL��yr(y�F��0h(�� @�б�y�����0�+Q����n��yRJ��yf�`�����H�� )6"ƺ�y��kۆ�Rq�į>(�pJE"��y�!�*K�l��./��tp�ŧ�y2DL s���Q(�<��݃����y��D�Wm�QI��`��M0@�N��yRM��;�(�3%_�S<�����I?�y©�.$��B��M>�:A�1�y"m@�n^D��K?3����k��yr�R M���Af@	�U��X�Cͅ��y2.ӊuΈ0D�I�EF&	肤α�y"��/I�t���U�1��ZK�+�yr��$�Dm�)"�� Ӧ�؊?!�D%�e�� ��5z�P$ 
w�!��:WC��95a����b����!���EPh��Ӫ?�l �BH_+b�!�$_��4�Ⲋ�1��|�'ȣ)v!�d�)%��ջ�(�z��"��#Ov!���
��R�Ԇv� ��C�X�^S!�$C"h�x��ԦD�2�(�2��� !��J�q�th�F$�c�<�4
M�L!�Dҟ~AZm�L��
"V0��ȟ5b !�d��h�e����)Q�hH�ö7�!�ĕU˄䒤�ΦJ'|����In!��]�Io�X J�V�j�F1g!��U-D���
�9A&�+EPȹ�"O���C�Z a0��A��#|;�.���"�O�5���Шj�z���DW�Z�J�s"OL�r�Ӌ5�Ή�2Õ#}���@a"O蹲兙�ok:�R%dH,IX՛�"OV\�i��8[x���m˫26��J�"O|r�h^.PM���K��e��E1�"O�T���!�|����͢#ll �`"O�X�!�� ���K'�@�4�X�i�"OJ��L� _�6�����3j9��)""O6��Ũ�.m�R\x�kG�*�0"O�d�G�����C"%N�cr"O´*2j��IQ��Ӗ*g*�J�"O�S뛈.% *Sp`s�"O�)궉�m�l�T��+YN��{�"O�#��P�H�H%
7H^5��Y0"O>i�F@�b�����@�*r=`p"O���q�X�Ty��R̶6�8���"OZ�hƤ����Ƀ+��yZy�w"O
����["�C�ަ.u"��"O���e%`�I#�F�q�#d"O������v��QVF! Y��[W"O<D��R���B%��<Gj4��"O�
g�v���qoG�4aH���"O�M�u�G_W�\��+I�Z�d\��"O��4o�;R�e�jJ��(�"OB43�b^&�X�
�fF�j�±b�"O�Y(ՊW�j�Hb���R�~�2a"O� ��c�ď�(��W�LĀ�"O�lk$�^T4`B]���l`�"O0��ހL:B �V�e~�k�"O�x
���^F���5�ާ>� 9Ar"OX���R�B��"U�@�X#hiH "O���q�_�5u���gcWs� x�"O��x"��X�9p�":R���""OF�9g�'�@kUŢE�\rgO�m
�U�q����N[�� �	9�!�$8��(c%1x!���i��u�!�D�c�L9C�Lb~�XXqIA)2!�D�U���gE�.Ey�,`r��-C!�Ę�v沘�l��?b��i6j�$.�!�$�$�fxR$�V+-�<��0��/U�!�D�5T���*���	���L����
=,�^����.Z�H�9��E�lE~C��2 	(����7�PP�PJ�7�hC�I��R�Y&-TWhѱ�O �O8C�IN��93�ߎe�6db]g'"C�IΠ|����a&,��Hk�B��81��}"`�K�b��l�g
"
A C�I�sIPhʠl����v�4B�Ƀ\��DБ�F*�Rl�'(D	Q�B�9g��=��T#VU:��%�C䉟s����� 6+P��^Q���	�'�Da�t
Ÿ8~�t�%M��Gv�`
�'&0����+(P4��Q&T�P�'��Q�Dj�-%���J��ũ#f�T��'���@�bQ*l��-֓RA
���'��A�TNJ14 ����@V��-
�'ӆ�餦L�wL��Q��*Lk�U�	�'��u�W�S�:�Kq���IuT �'��(��tf�BKΞ<5f�(�'LȅHDE�.L������7]��B�'�����E�h�p2�1$"�	�'È塑���� �v�$\+�'3�C&(ď ͠�8��B�!$X��'a^43����u�����W ���p�'n���!���M��oT?��'k8�2�� ���X�+� �ɩ�'��|�ѫ�%�dH���	<aJ�y�'3��p������!v�@�D"���'���u��>A�}R�#�%�h�<i�_8���Aƌ�1nҒX�FLN^�<�b�JJpz��TI�91�)�X�<�%*�mR~�XW�B�x3r�(��NT�<1&���
<�v"$eĚ���n\M�<Y �T�<1��ag�["9�8b���E�<���� ���:jX���JI�<)ABnt&zp�� �%�o�<!�G��1"�L{��LS�N�tʐj�<a��5\�$h'D���Л�%c�<�u9�z��R��= ���y���[�<A���$'b����P�x>B`9�Yl�<����<c R@S��-B���@��I]�<����n��<���Z�=!����S@�<�p�σ ���1��+����\{�<�$f[�b��,A�#λ;�*��v$Ax~re���0>Y�K��`�����4�^,�P�Z�<�S���.x���ڂ�h� K
V�<a^ɠ� �-*�p`8�gUR�&=�ȓb0��ReKߊ5H��A �$��ȓX�d&b�%n���1��A��$��Vs��;CJ�}���e!6r��S�? DT����D�v�� Qv	($�|�'�֥Ǎ[<��;hR.���9�'��0dg��r�
�Bч�9d�x��'�r�&�ݒNr��b�L5E�q�'��ۡ �8x�F=!0�n�j	�'�v�C�\GW�H�ܳ��
�'�$�;����%�J�+��,��E�	�'�l�W ��	�ō
՘}�	�'�>A�ɏ$8��m�  )�|��'4 -���^�?�V9[�G�3��<��'��h��X'�`[1�_�G�N ��'��ih �Ą-����@ �@�����'�^m@Xh	G��)Sd1Ӄ��y��&>n��SgDF���eFP��y2�*e��&O��Be�X�����y�C�$2xa�"P(;���w"0�y��i�<e��<7�9��+��y¤O<b��$�3�؎?hcg�֦�yr�� �.1��Gl��h)��y YH{�D �-�J�t��yR��o�,=3Qj��4EV�j ��yrb��
�($(��Y�&���y� ���yb���xID3��E	Rm��y� 8] �Y����2�4���́!�y�i��X����)���
��yBA�z�T�*(8����F�Z:�y�Î�,�h��߭-n~�`�*	��y��>gv�2�������6�y�,jA����!H�hѭ�y2`A:!�jꆦJ9r pS�J�yb"�s�8�E�U9����RLH��yg�	�	KW	J88r���y�E�Dv�P#�}�.�x�bK��y�j�&4�fi�U��3y��r�m���y�Y��QRĎth<q
s���y"�؊ -�pk�,C�oe��QŮ+�y҇C8_|,paǭ�np�����y�M&D�0��DkB���R"�ybG�x�X���^�e�D(���y�*Y7*
���� {��B!���y2&חK�HL�֯h-l|�kQ��yB�04�Uɋ�c�@h�'ſ�y�g�7r���E+?Y����邬�y2��%]�-�Ɖ��x�D�S��y�	�=	�v�^�jp�
�S��yH���U�	&�<L�f���yB&�d���c�gB%y���y�̎O�b�����mJM�V+[��yr���M�*(h��H�8{ ����K4�y�L	#�����>-4�r���yrn��o~���N��y����f��yBȃ�H5 � �PrԨź���yr�ٹ!2Ȱ��_�e�B�v���y2�	<�6�C�@
�
��)+V�ė�y��(_�r��6d�����s`�N8�y��]A)x�*2ɐ��ǅ�y� ��+Ȃ���΂vl�d��'�y��G�3�uB��2_�����(�y#���aң��-;�t1��+�yr$�Z^}�G��P��\)P��y�mB�4���ؑ{N�P�C��y"GզW�X5�3�ìb�dLpN���y�H��@>��v��]d6�7�W�yB!��|V�u0%�\�9����y
� 6urH�p��8cg*ߘ�H�A"O����LѓM��a��3O��I�"Oh�kQNص/؈p4%�]>F�A@"O<qS'�ԭ%���:U�͂!=l� "O��)"��N�	��u�H�""Ox�YM�2U����W��2�a`"O��ȟtt (
S� ;�:yZ�"O���v��Y��1����u�L��7"O��Z�$|ԙ�o��~#�]+w"Oy*�(�2�L���c��~,��"O6�����.�ؑ���	���1�"Od�ِ�/w��)cb�J77�~��"O��(�A�(+�� BŮ��6tr�"O\u�u�Y)^�R� 3.ɮ~ָ
"ON���!B�b����wLX�=�M2D��� �A���B�V 4Z He##D�Pi��t2����g 6�R�/#D�l�5��8zR���AI-D^��"#D���5�3D���YwaF�`�B|`�&D�h�Dֽd�"	S���rB�� E�'D������&T�8�#��7p֬�6�!D�|Y�%�8��X�c�vqtY�1�$D��+�$�H�^`GX!L������?D�@R�gO�Ͱ�BJ6?��eQ��>D���ckk�Fׇ�pn�@CO��yR��v%�e�R��@��4J�o�yrIQ�j5��(�ȋ��8������y򅛨c$M�u��z�x� ���y��<y��F�V���f&%�y�Ϥ�I�(���!�!��y"����`ǧ �"��߀-?!�DV�MX|H�%A�9Ft��d,�=:/!�DO,
1�Y!�F�OG��23��"!�ǁ"��ኴP��KBbA!�D�'b{L}��X#`��ݢ�˙�Xa����b���J������Blߵ�y�������̴X��U�Ⱦ�y��L���,��%@37�3�I��y�%K8.ɑ��&-�P��埞�y2�(}q�C)�Q��X��y��T�6�D���eܙ"�(��FN��y�m�F �m��a^���%�Љ�y���Lڑ9�
��4.N$1����y��P? ������\�E�wN�y��.���[��ǲ���q��3�y�c�[P�E�Q��y���4���y�Xo.p��%F?�ࡹ�E 
�yҏW�}���Pd��l��%*�M@�y��D�=8�� �ߐ_?�PC�٣�y��ѐ}@���o�7n�"]3����y¨]�uj��Ύ�=mnihݵ�y��E�J���I��Y�:آ(��A��yRL�Q�Ӎ��>a� ����y2EԺ�,T�V�� {D #�_5�y�MI�A��R�kWL鱣���yB� (�Ĉ�닂3��}h�&�yoD	8$qB� L,��aa�� �y�bʂ:H$�+�c����ph��y"�>;����Pꅦb.�	G,�5�y"�Ix����6�M�q�F�N��yR$Y*����1�S�F
y:��/�y��9���qō&l�(=�%���y�aTt�+R��f�JXFcQ>�y�n\:_���2/�\wH-9tNÀ�y
� B�A����,��A���L�v4@pv"O0�8%4-$~̂��<<���"O����M�-߰�Y�7S:��"O���V�6CF��i�m�4�I�"O�����[5LƐ�Wcʔ@)I��"O��� �H!|��Tb���a��"Opq[5H�2c_��q����SΙQ"O�哧(��Q�|���@\�=PF\0v"Oj}I�
T�v��٣!fJ2-�AB"O��A�ה�n�C��U��`�"OPq�ʙ�L�)sd�(&{ U��"Od��0�,mJ��[�b�:���#�"O�uh��7F��S�/W<�r�X�"O �)����;���w�>�Tyic"O���E^? ��Y�.�g|z3�"OV%@A�T.!�����1~cN8��"O�)P����<�WO/V&��E"O`! �bP�2�iFC4ZC�{�"Ob�ÖfY�/�$p�@���>�`��"Or5x�K��t�=��K�BU��sT"O>���iK9�.yYa�������"O5�fK�\���T�T?>�V��%"O <��,Z!@�Dx���V=4��}��"O"A�Q�AzJE�� N�R�Ę��"Ox1��]�;�|�������4�� "O��I��g��x��ݰ_��=�"O����;]�AH�#ތ|5�"O�i����%\�̩C c� �
"O�H5I��
d$Ԉ�h�E�"O*�aa�^�����ao�?�l�"O��* S�X�p$��x�"O���a�J�$�.%�jL0�`)�0"O�!؂@1Z�`(�D��r���� "O�q����!��)�'�^���"O��3�P�H�r���HK����"O��
tʀ)Hh�b����4�d�z#"O���`?,�A�"��n;�9q�"O��Kf�9��Y�&�Hd��"O4@*3��@f�(8rf�9$<1�"Oʨ��"�A�fhɖO-:&(��"O�����/K]�qc���6�1��"O-2dܵd|�5�îF���A"O�Y�"����qbb�H��- #"O 4؂hL�s�µ{$���qt|�"O<���cOa'4��10T�ia�"O��у��|���g��t;9�"O�H��_ %�ph(�eL�&/����"O`PQ�]�+t,�H@�L11ɼ$C�"O�@��30��*a�EL��z0"O���e����hȉ�d�-����"O�`�K+ H ǄR+08����"O�u"���W��p���?5�MBb"O��z��8Id@��p�_�h����"O�dC�N�%k܎p�S&͡*d<���"On�˞�a2���o߬((�)�"Ox#s% }�� 	��N+e4�hr�"O(;��
#.R�Q
<N�`��"O*�"`��G~l�!�����P�"O��b��+�𸻴j_4�ؼ�"O@@�����L�+���84M��v"O�m�#ц[ʑ����&����T"O���Pa��`{�M�����('"O<<CR�Oto���bB�'����"O���I�F~�A�&� :'[����"O� >�C®w��h ��/,Cƌ# "O�k�f@�k9����F c$4!��"O(�I�C�I-b,S�O=$�H�"O�rD�a��U��q��i2"O^������L�9��'��� @"OZ�����mr���T�x��I�"O!�eL++��<���f�abr"O@!A��I�+���"^,�:QR"Ol�sEN8z(�ș�.��C"O��@�Z  ���z��8J�R�"O:}�5��59�`�ő�P5Q�"Oԉ9����Y,��D�*jp�	"O��X���=�(Myu�R�Z�6�yB"O`: �@���\D-�Q�*<�"O�T,�,Rp��߈K�v,h�"O��ӭ�0L��jʨF���V"O\A�RZ����,�&��lҔ"O��*H�:`��!G�~�J�bu"O�E�W�F�W���7�y�"O8=�"lݨ` ǭZ�^��8��"O�}�bfJ�y׺�HmG�h�t�؆"O�$Ja\�P̜�)qO�>����"O��[b��t~�Q�ɓ3k�����"Oȡ�nӃt��YU	ƪA}��*�"O��ǒ4�u�P�Ґ5�b�""O t�Vŀ4J������U} �Ҁ"O�a;�`U1T��q�BT(|��4"OnQ��N��Z��'�D�E]()�g"O��AW?!��/����	�'JZA��D��U�g�X�kL����'0� ��AIf���Jg�]��'��$���_6^t"0�b�O1gt��'���2AǕT�a�g̯2����'�>XZcZ�Z �J�	��i��'�ڑZ0֝q��4���F 00�D��'��x:U�~ՠ`G�QE�Y	�' ���cǾt}Ҡ�W�8����'x���_�A���r�H�d�j
�'��; `�?>����a�HWvL 
�'/�h�F�Y�5!n$kae�Dx�)�'jt���$�%e��Aa�Z98K2 z�'����+�DٷK�1m�1@�'"Z�ږ��$r���G��=,҄b�'���)�dtÃ�b�ذ���:D���C��5�U D�هM�h�7D���F�2Ű�� 7���H �3D��q&d�3m���b���IȐ��0D����d�$�@�#7e��(c\9٦�-D�L3�җ;�#�ɋ�>%�*D��b,>��I[g.�{d�`rpc5D�Py�˙s�fU��哢)k����@7D���2J��J���MB��i�m4D��C4��J �]ذ�(O�ܐ34�4D� �"�!T^��� ܠe%0D���pcH	2��m�$+�5׋.D�D�FK�2H�P����$]��F*D��ڦa�����׏3�xu��%D���p!N�^�L�A2-�p�d'(D��80�ܐs�tP3�@S�S`�4�%D������
��Qz aV�roj,�FD.D�P�sʈ,[ru#�/U�w�x�Q!,D�j��
�I�8ȩ��:d�/D�;�-P��p�ʄO![�1:�l1D��f�O
>��ICѦҨZ^t�9 i0D�� T��gOI5��
���J���"O68@WY�;G�-���I9�va�"O2��$(�x�V�ҦhD�JP�=0C"O�<`�ټE�Z�*���O��`yU"O�j-Yrx$��dL�E��ݻ1"O��!��y-3U%KA�N���"OLM�fɏ �x5���e. �r"O���:!�Y�F w&P8#"OP�Y��X�S�]�O�!c�P�"OV�k�b�x8ғ�ٙM�es�"O�\ӑ�\f��9��L�'I���u"O�qp�0@� ��%M�V	H�	e"Ox���u�\���Ƒ#��"O��3���'��IVňM&:#�"O�\���A�{� ��B�"i �"O��	��B#?*n��P
X7 R�c"O�t3!M�.�����e^���"O
՚w�� FD�e�ܖ�:5ҧ"O�@ӑN��4b
XBRKC'��(�R"OB��a��lhD4bᚄN�v���"Olz�`˷s�z�[E�]|��2�"O<5���?���	�9]�ӥ"O"|�dl�!+}��za�C�!�����"O��K�eҥ)d���Lc�"Y�u"O m���ޑ �6�{ׅZ+r�0��"O�`8#�  ��9��L�&Ҷ�"O~��J�6�"T�#�P���Y�"O�YG��
^�����E�lU "OT���gղ6{r0��b���¸��"O�]�S�+
Xd��KC$x����"Of�HU��:^����G�M[rq�"O� ��u��@��L�	���D"Oxe�#k�2},4@Ѝ��f+��J@"OP���jН2�����B+
�`"O�0b��Iz�؊�;�e��"O^(��$æ!�g�Q/]���g"O�<XUf�0Y`D�p� R�4)�r"O��qE�#��Lٲ����R"O�9y��N6>E����(@+u���
�"O�]�Ԃ�TU�$:�}��(�t�3D�����M���Y'i8�xY�`2D�8Xd�2��]��Y)?�~�3�4D���'n��i:pI�K="�b��$D���jA�!L�	%�R.O"��2i$D�tˀ�Q�*-�R������ D��HA���%ې��%U('!v�{4�>D�`��hM�lS���z'dmr'H"D�X����~5t�q'�
�*a{�'6D���0͔h�T(@f��n���'D�|�qf�13�\�#��'� i��9D�4�Boӥ,<�t�O<�P���7D����7WVvmQ���,S�X!Qp 5D���-K@`�&�'LZ0���g2D��rl��-o\���@J�3-���.D�L��ٽM~`PÆMI?��H�
-D��y��AP�B�Ѵ��x��(�3� D�$V�* �L˷�E�W���d+D�,�q�@��5��,z���*OZٚ�ꗬI�$i�F��=���Y�"O��A�i	��2�*Ҥb@���"Oj��Pd΋c���,&���'f�\��oY�p�♑��G�*`)c	�'���h�2ZV�h����6lh�j	�'�bUb�ֺ�2���LJ�|ʬd���� @(*A��
���I��ބ[ٖmC"O��)��ʥ}�0����C�Ԉ��"O�)�VG�4IJy���vҾ<�S"O� @�)e�J���#[�E`��K!"O�XʧBP�.y����I^�rs|!!�"O��( �p��5�4OS'©�"O������*~H��'X�쀀�S"O�������S�F	����(}f%��"OZ8��ª���jg�G5=�|���"O1"TG�n���yF+��^�PA��"Ov�1����
Ba� 7\�Z�"O�\��Wn�<��E
�z<��E"O����H�Vs���Y�1�hf"O~p�e�]+_w�h��唟|)�E��"O�dBU;�-;'��>?ò���"O~�W���6��L�@�R�5"O$x;�m�;}N��kX�pR���"O�i��ۥm%�؃���-GKJU�q"O�i�r�ߒ1V$\ g�{,�Q�	�'��')Ԣh� ���X��ح�	�'�8��Ꟊg�dс2�V�_
F)q	�'3.5�H�7[�������U�<��'�ƹSpR�M�n����2S1`!��'$U"w��?@��A޼M3Ե��'��i�#&_-Z@��Ȑ,E��0	�'}�D�AD���d�P�X�tez��'
t�*��57`��`�]�e8�')�L
Ѩ�*_�`�7)��
����'~�Ac��*B������7�����'��l*�g�7E� `�7@ /:D��'�@̉�Ǎ�Q.�Ap-��v����'w���FD��\r�`10�ۄi��I�'�^`3��Vצh��/Z{B�2�'F���O`R��g�U�����'*�sa ���lX*��"dx��'0���F	�s���	�_� R�B�'ɖip���b���@�B�
���'���A�ԱMpbmJ�&�	@"5��' �Aq& D=�F��ѳ7�J5�	�'�� 閏]�]Y��"�Q.�&�{�'�0�/���2�@=R���A�'-*���X��L�y¢��
�'�Fmi�X.q }3v�U�j�dP�
�'ξ r J�<�ځY�7t��*
�'�X(A1 ш)&�C��:��4�'��l9�m �"%>-)�mЏe2��'\8�Xq�#%9�Bc�<s�'ꎘ�'݄/D�9!��X�P�0�'�B�c2 ��W��@�N�B��h�',�A���2 ����#PKX�x�'o��J� {:I
"mV"E�B�	�'�d�c� Ea�(����5���1
�'�
�O�ii ��b葤,"�x�
�'���%�Z�L��c�!��	�'����;lnyHb��(yL}��'`rX����ʸ����.�Ԛ�'Y�8j�0A����']޲�j�'����Ǽ0���'O�d�
�'ټU[��\�G�$E�?���3
�'�N�x�MO	A
�`r���IRZ�Q
�'��lX�I?T�n���1����'��鋴���Fl�\)�c��n� �'xFm*�b֨^���C�H�4Td��'^x��@�+
!�DR�h�x�
��� (�6�C7~�4j��N�`�q4"Opd���h�|(*bcZ�t��#6"Of����c�|! "̑�.���"OU�6���8f��@�\=�\��"O���RGISn2|{嫋�&��T9�"OhL[�*��%��A��i�7k|��Q"O�UJ��o��鑪��7�V�C"O�M�VFF?g���3H��%+V��F"O�9֥�8(�����	�%��Q"ORT���<k<"PAa0��h�C"O>`q�g�K�����@��G�<e"O�iDf�&+���1�NȶL���X�"O6m��c�����d�:
�� #g"O�9�`kD	,ۂ�(����QUt��"O�b�P)(��a�1-F�VD(9I�"O&|qpd�6*r�(��757�!��"O,;6$�5_��6��"&긛G"O�UѴDΘ,�"�9g,��5
�Xч"O�<�4��>/���&����L0�"O��a�ꕷХK�@�<-�����"OT �e�.޼�#���'p�}�"Oα!�j��/�a��EI4V^���"Oi9�Iڞ� EQC�S)&}D�'���I�H�嘧��>�0G��G�bP��y`�|��h*D��`Z-�P�z��[:$̲��5ˤ>���
��-y��'A��,�!<�6��%k�,�F5"� �<�*�HܑD*��H7J��b��dPP#Ҡ5M"���"�Oh<�U�*N�:��(�"8=bt����]�'���#KȲW�m*5�1��F�T-A孂�q���ҧ`��bu�B�I%:b�X@#�!�5���P�:�X�C���P8��Z�mQY��,�g?��̤z)JH:ǁ�Hb��u� \�<��BQ9FWl��
���\�7��ݟ�{$%ւ/����} h��D�1�4k�fL=_����t�N�y�F�=^������
�H\5� �[�H"�| �C��$r΅��D

�Ś�'�v���S�N?xE�C#Mܲt�L<���F�,�}і)�\�BL��)���O�ơ�uK�x�V!��A�?�U��' :`�e�(�H�Pǭ��"�l�j``�'[-"��A�Ռv�v}�����O���'����&T�{���"f �@jԌS�'��Ď۝qu I����V�6IgΪw��!'�R�mq�M�
�wp褆��2id�Z� ���!��a[Xz�?�s�]��HX� �mov]�a,[�;�c��w�
U�%�<iSl5J��x(<Q��^}J\;��-.�՘ �yb�Џg��l��C�w�B��#���P���P5�q3�� U���pc���y"���.1 �8��НqL��i7nՑf��<�£tb�1�d	r�N)N~
��[�$0z�Ĭ���ZL�^��c�54Qa�FJ!c��y2�.��E��i@�AZ5x8�
�mK�%�"DoX��q	g��r��x�j��9i"\����
I�}��A���O���|w$��g�{.�r
�"::�m9��N@.��b�&�t��c\V(<���@��[�h�;_n����{?�%�By����7a��ɫb�\��K�韓^n��;�E��F~�P����!�Np&H��s&�U��#l�G��y�b�:h��#@Ś	5��h	��~��`
4h�e��18��d��pe�H4m�,��	1I}�����������ؗt�0��A�:�R���\-��I��g��g9��ǓN�0��u�	3 P�i5��Ul��E}r�]�{��\�V��} u��K� �(�/R�~��a�4��?	/h�4�`� C�	�H��Y�Ǌ�mҔ�{��L�H����?T�L�fl�(Kh�iz��Y��[%�I��OAb�Ҫ�i��5�<� i
�'$T����Ȳ��1�0-"~����;jy�0��H]2׶	�G�ˍ��S�g�e'�,��(�^ћ3g��Ih�0�O��	��O!$p��� �*"IdI�EC�qz�x���ʪ	���5CY>��'�)G��� �R5�Ѥj�X�b���9��u)V+j�*EK��*����eG�U�n�KQoD%s(���e�a�<��M7���[ �ǧ�ȃR�Py��!�^B@�
 1CxMy��M��(���6'�>w�z]�WBO��("O� R���#$Jh�
�(�~�� f�ŁK��Ɋ{���IAL2�3�I.s\��c�)C5)V��� X3[�~C�ɹ.�d49���#Lu�q����#�H��	ƓBJ9��Z>���L80p�`�$D��.�Z��ȓh���pr*�	}��)��6l�%�ȓ@z���hSos2��&a�f\��&"�|���_+o?@ ���
����ȓ2Rz'���T�L��
�� u(��ȓ/h�YV�c�Dp���SNh�ȓC�<�i�J�N�� e�
;]0�ȓQR��� YqR����U
�n���`��-c$��j���ځI�$�ȓ<�)��GInހM:p-E�Q�ޅ��M<�0��J W��	jdbYH�L���KqD<y�+	�'V���5��v{楇ȓr!4��dB-���GC@�����8��&ɤ91�!�e`B�&E�I�ȓh>��PN�9�ht���z!B5�ȓ.'<�cJ�2��5!7k�9��!��O$������]��<���O�A�,Y��	%R�Vǉ�g^��3bJ�	�a�ȓ^N�UJg��[�d����('jT�ȓ � =��bE [#:X �o�?>��d�ȓe,~D0���&~�@��f@�K����:-� �,�g�}�P$'> ��Ge��BROSF�\�p�S<3\\��}�s�5E���S��'�E��j̬���1Rz��s`X����AA쌉!���>�ȤcJ��)ޅ�ȓJ�����N
�2B:����%��ȓ{nlM�b�� %���*���8`9t�ȓ9۴u�E��$�����9,����"�'���!琴q���2~޸M�ȓTl���VJ�"G����'nI|�f5��|�P��a��w��ԋ�,]Bn����?�L��	��
gL�^�P�
�� D�|H�i^� Və�}�@��w�?D�����[����xEO@�y*�!�vO'D�x0��W9$�t�!F)��Z��!#�/%D�l(GjXR��0Xi�-��-j�a#D���2���D3VM�n��I�&d4D�����R�0L攡��*3�i�*2D�La�mJ��{eg��xָ�9��.D��jդE�������'=���.-D�dȥ��VD��u.��R���N>D���G�3<��xp��E-?䖸i��?D��c�aݷ]��R,��(��5��*O�(#���:TӶ��@ ��_�P3E"OȠ��Ҥv���r��I&��h�"OV�K1�56J���E�� �"Od��s���Q���ԋH�u�-��"O�<�-\!Prz|X�
Ƙym���"Or�H�B���L���D�4��0��"O���`�)������3�<�2s"O���F�5�*���8L� �0"O��Ѝ�l� �e��$ ���"�"O��Ӥ�]�.-*�+
|m��i�"O�1�s��q�t�آI��^m��`�"O���Z .π��P�Ո%�$A["O ��6
IjwN +�S�`�dA"O�^
���% �c�	�&!�y⣝�a-:��a+���,<ju�B��y���-@t���+R�b@J4�D�y���v�\�����0I� $��
��I�" ��*,O� �@�dN�-<n�E1sƇ��~�`6�'<�Ų2�R9W����M�XuY�O�>#h�I\<���%z�p衧O�M���[Z�'i(�v	�%^r��sA�v�� X*�Q�c��R���$�}s�B�I^l0sF�0A�" �>^W�7��g͠)(vH�[hM����}��M��,K	��u��'Z�~\cA�Rx�<��X�$�l��IW�>�
��Z�҈��M�~m�3M��rG����HOJ� �;��˰̓d���pS�'_�Ւb�4C��H��I����0��jX��)ɯp���I@�NL���Z��t����L�c���C'% �uQ
�jc�P�q���Cq�a���=�hM`�c�Zl$��wC˭��L�ȓ5� ����+�����CٶQ���RqK�{��b0�>	4�q+UJ�-�h����:��%/�4-�ZɗL\# �!�dA�M�<:VEĿ`G�Q�b�P}��t`�aPH�C�D�,�VxCU7�Ԣ=��[zYkcɂ�0ĉ��^��ǁ�=��<�6K��r��Q�r/�l�� "��F�xp��4.��M���a.6)9�
��k�@y��[�53n"<A��,�H@2���!W���JK7��6�`@�&���
O%!�Ĉ>q1�eA5�NB�k"j�����3GC[Q��`���#������(��s �� D�r��F��?����c��t�<��ꂑɨ�CP�ġ���S��.]�&���9�\4r�L��0���'�hO$�y�$�+`�N�i��-b����V�'�lˤ��7^��B�[:/j��0��
R<�ST������[
��}+)s
(h��L��kѳ�(O1�P��(w 8��ѻ D�˟�c�:6,
"P�0x�MG"O���3H�7�^dI��37��I��	�>�,DJ��D� �:,C�Y�>Q?�$�0|T B�.4Ρ�Ȝ�|!���B���F��$1T�G�X�R��rhD����#dL=St_?#=���x�4�3�4�`��gqX���	ϯ`^
��7�T#Q\X	�d�z�:�Aц�(QF�("��U����`^jT�h�N
'�>H�7k'��(���fܠC��)��
4P��1�)D��J�t!� }��)���) �ti��ID�]��ΡNH �K��)�'M0,C�<d�BC�M�:����.��(��	WJt�"�n�3b��t%��*�Nճb�ay2h��T��?2�J�"S��w�!��6<hZ+�<rTLzr��'?�M�ȓ(�8!8�B*W����4��!Q���ȓw�"$��	�����N1艄ȓ)�\� ���/"���y�EO<UF������T`O_�pmAQga�z��ȓ��h3GI|�u9e��>F
��ȓAtJ��3����q�"-�>�ri��hĐ)��ۙ6h�qqC91#D��ȓT}� �����"��?�����8g���?�Q�u��-ȅ�_s� �q2I�Ԫ�'u���A�"��'R�*�F�`奐�������6H�fX������j���J˺"U�]�#�X��E-��'���ȓ ��ћ5l΀$�B!�œ�B(�ȓkS h(�%:LHIF/ϋ%�$�����*S,E̕���	O����|�̬2��B��(�z��E?OLr��XUTq�BHG�w��%�I��f�Ʉ�%8j���i�FH����qG\Ň�IO��2�+�lնuT�W��*���zEtla�i�*;�ꙛ����o׮���!�ʝqS%@�BFf}s��v���Q�Z��'�F-򖝚@�V;h�̇ȓ5�f�i�"L�i#C3d��ȓnR�x��ܠ��!�60U�L���J2����	Jqr���eصHN�H��u��}Kcc�#0�Q�V��
/� ��S�? L�� /��Дpp
Ax��Q�"O��i�nΘE
D���85�52"O��@q�N;�@����G��'"O
$��J�"�d�T�}1"O�0r0��4��)څ*ښ�ر0�"O��C��+����vN�p/�%i�"O�\+�W�	�֬��ښ~�@AB"OMR&�ǁj�P�zB�۱oh�z"On1��%2z�p�{�cܩZ#j�p�"O"apu"ז@�6�+���3 ���"OdX�4�%&\b�(� �s�
�Y�'�y�$�9 &t����.%t�`��'f�}Af+V�z��7�ȅ�t�1�'�{� g��\��	�(&���'��d�A��P4�bd`!�,K�'8�աrc@�^��4�^*�hPx�'��< o��Nv�@���
� "�e��'?d�s׌��:`ī"J�F���'@����א Wx�6�ɬr����'h��l�2 B��D�]�dVĝ��'A�$�@'�<-�T`� �ޡ^�ua	�'�x �%��"|DꐅɜJ!.)J�'�j�['�]
#o�q1�A�ek	�' l�!���E��|��n�A�����'�L�i����p�(�굣��0���x�'@dᅞ:CED	��H�y
��	�'Cx]`��YF�;g�M�4�C��V<�)��E{�S�O�Z���'�� ; �2���!@"ObEQ$;)wةP�'��.	t�R�@��΅�=}2xYӓ&UKG-*��	4f��N�\��I$�0�Be`��E�BD�a(�^��8���t��!�6n$4��臅@� `F���.�;2�As%N1�i��1��� O̜8��I��lAr�f��>0>�`�>b�!�H*�D�`��9ghX�n��0φ��@NE��ڸ�F�y��ʧ	L�dI$x#t%?`ȉ�U7D��ٓ�E>Y^�p"'I0�r���A�O^軕%��"y�(���G�[�x��ЄB�̒�.K���� �+��<��ϖ.J���RB�ڨe�i4� ϒq"�2)b墠g�
l���G~T��N��|��zCÂzh'�<���+ :�VhN	P���
�/�cܧz��ؓ�B�v{��!��0��#6�HID_�:��ғÔ	o�c�AM���CG�)>?N��v/�aܧ��OL��QvD �B�^V�9��~LT"BL�:�F$���,m�e����!����� \6B���k��=���񤌀Et��$��la���Dmџl��Ȓ\J`�m�-N�A�@P�����뉔a�XD�7,[)pAB}i��>��j2��*�J��\�S�4Âè<!��w�X���lʌ&���a�)Q��%�}���0[,e�T�R����HFg�<�@�C�1p�D�Ve�*x�P`p��"pq�'��o^t��g�I�+*�$?��'�)}���)r\��{c�1ra*��t����?�⁒P�&QR D��D�����oޡW}�X�� S�OJ$3��I	��12�G�4�p<�g"�v�� ����h-�9+�x�''�XQ�K�H�b}�&�4�l���L*��E��ȮXk�,C����4�Ro?�,��Y�E�Z�����y�1�bO��(j�B� ��T��l��|�ȣ��S*V�@��e�=	���Y{6FX�Ē�y�i�"��[B�¯cbfQ����X]S�+;"�>�26�WH%�,�I?Q������IY,Lmڶʂ�MV8 W�B�6��䐵Vv�X�ưW�\S@�׻xD��'j�0|/p0/a�H4K:)��#u8O��[Ѫh���7O�\�ȗ�	����ض�P;�~=AQ�	y⼀�JL�Vm�x���?�V񃔍Ǩ&�Hb�'�H����@�be8X��S#h���'�S���k3��z�ԄR-Zٛ�@ް0��>uL�=5��m@G現`:V�	�l#D�|t�ŔB��り��Y�6X2�D�VP��9-��I��	� (&�O]Vŋ��xR��-\Ozl2��o*(-�� ���p?	���D�biCD�4��`R��}Z���lδ`I�$
cA�%�rU��eQkx�� |��ց�X�@1���������60d�tj�S(���휆6:�h� ��}�bGE^�VL(0dh��yRB�L
����샘f�ԡ#'�����g�5�2GV����l�n�Q>u�qk��a��̰�K�D���Zs�.D�t�`�ƃ2�t�7Jɰu�t;�O5j�`8�H�6�^�g̓=��0��16���-_NHx��RM�u�PF��B����Qi��F��"�ݗg�1"��'QP���ׯgޚ@C��qn0��'��H�w���Z�!c�� �rM��'�ĳfC��8#����Bi:�]2�'BL�ͪ���RgI�m	Vp��'L������,D�H�`�Tp��dJ�<�Y`4\0�iӺn�V�Ff�M�<DV��hmx�e�9���ᓁ�J�<�0쓃m庄�t��:m`��z���}�<a i�?Z�� ���>/�)Z�b�<Q�k�"9�y"�Y54h{ׄ�]�<��ɃF�P����6�dR��G�<A��޵s~�|z�nG��u�p$��<I��-����� ���a��~�<�`1פ�aV�0���Z}�<q�c�(�^�c��ܼ*�(0��@W�<�Ƭڷ��)2Ǚ?�>�+��Y�<�Fϕ�Od��"S�@�Q�[b �U�<��n^ �6T��%Úg��![���t�<�tiU1I9�Hc�` �YT6}[��Ty�<A��@��L� )�f8	��@y�<���95�Y��l��I۾�_�<�!��RI��b�6�"�A��A�<����P���Co�h��t�Sa�{�<�G�+`�n��J��:p��ąv�<פӎ.��@f�^��`�w%�u�<�6�˰5
���ғseT��Ev�<Q�K�D�<�,
Yv�=4�Yp�<�Uo����Q$Ǥm�ko�<��'I�y�0��l���jW�^f�<Q�N�h�����B/�Z DOW^�<�#\�x�R�� +khũ�Om�<�e�A'xDBB���&��eqM�<�ɗ�\Le1 뙢]��)g�\�<�k)1ZG�xcx4�T�TY�<����6N���c
*��	��A�P�<a�!��QS� ��e)Bˑ�M�<�3D�l��2w�K�G���փO�<Y�$�	9�nI؃�_�d:A	�K�<9�L� g��@BHW<��ҕ��L�<��nK<W$�Q
	�X`�
��a�<1�ۢaj�[6�8g���2u�
]�<�
����6Y�#�&^B�<aǡM��&��l�0B���K2̀v�<i��B�[))p%`�]��{d��q�<A�+�3
�hi�qaܰ�.5µ#l�<yL��&����A �,i�H5m�i�<���(�}�M��7fACV��L�<�uF�7f�������iI:�
')FM�<�BD�h���#0+�+N�`��GR�<�U��)$� �	�S��D�W�p�<QR��6~|����mZ�;]@�H�Fo�<ѣ园^�r�2EM�pӈ���^h�<R�T�LX�d(��W~6U�H]�<ّ,�.>�xhaL�Ɉ�a�X�<��N��Nx�􋀻lwL�+�aWc�<��dEQ]�s
�(�1��p�<yw�ą}�n��ġ'9��dK�q�<� �=Ѐ�èk��=����`D9�b"O�䋤-�k+Jp��\)�xzf"O����ƶ6������ʼB��C"O���&	�.!.����oӤ	a�"O��pJ]�9���A֭��0���5"OB����il��!4�(�p�h�"O��քI�Il@�dK�_� ,�"O� "�e��J�'.�F�� "O$�&�)= ƀ��b�.3�P��Q"O��Va҇/���r�<�n���"O<�h1���~�
,H )[��Y��"O�Q�v͐�5����B�5�4�(#"OB���{�l��Aʡz�<Hv"O��	����Ĩu���:�$lS�"O�!y�&��o�HaH#6@�0�"�"OR0��0����Vr��R"Ov�QW�%<E�Ad�xB�hG"Oi�{�H�A���6�Vؐq"O�9�'�L�%�@yPm�<f��u{t"OD��*� 3�F�x6M��\Xd)��"O�{&�^*[�d㠌�HF�D"ON�s��\7%Sh|�V���nl�0r"O\e	�؃6���j�G�$F{����"O(�"Ø w���rS� c�\X�1"O@�y�֫+���/�_䔂�"O ���/@�Q�	S �C(}D�"O(�'�=H���#d�5nWz ��"O��K�a߻Z����]=��	�"OLQ('2��3Ck��Def�r0"Ol ��[�.�bJ]�jf �'"O�t� ���a��ɛY�t��T"OP��G�98��,znM?k�ڱ�"OuH�h��sMұj��3"O~q	��Hu`�6���zDJ4"Ozၔ���u$�@pqiD�i@���"Oj�i�'p8D=���B?���d"O�A"YC �* Ǆ�<��$��"O��27��^�i ��\����"O���?!��L�$�K@�4Ҧ"O�H���/5}���wm3e1��C�"Ox�Q��
C=��C�L�n����U"OV����>y9���PACqy<�#"O`��"�D3���O��S��h�"OT��5��)�]HA��K�<�"O�d�E��j���4'^���R"O�d��B�:CA���o�/Xbe/x!��K�>�X�v�
tr�"T#:1�!�_�/�a����?Aȱ0QBG�0�!�$^�fk|�9�昣]�`�c!a!!��l�2�@�]�(�H��Aʠ�!�O1������Z���r��-F�!���<�W��6��s2N�>�!�1S��-���@7%�R����Z0sx!�D�*ޮl�� Q!x�0�P��k!�DY)E8�-��������<|!��߾uZQ1�LK��9���!�D�F�� BF�M�p�ڦ�Y�"�!��J#"Y��\�J��AOS
|�!���R%⌂��t�l�z�/�� !��>.��ۤ��1yL�S��; !�S�h@�쌉^{�9��.��,R!��}"l���M�Z\�A��My�!�$N�؈�c��+k�
�L��+�!�DSJ��Z2���Z��@+M�8!�� ��[ +L;8��۷�	b�� ��"Oҙ)�l34Ȣ��b��&P�g"O��P�%�L24ы�W ��"OD���/
�+�r�y�MˈET詓"ODE��mG�=�.�n_�7�"O��9���O���H&�D���t��"O^x�a0w��l�&(\<���h"O����ZtT������7T�\P`"O�Ա��CX|��H�;;�X�*"O�|A�D�Nl{� eFܺB"O0)�T�$X"��{�/��1��)�"O�,� 	�8򔫴�Wg96�|��)�Ӵk/L@�Έ%ݚ���Ś!i�B�Y�z�Z'�S���4��珍<�RB䉥J�`�hg�>R2�����y$B䉡>lܴ�u�_-�<���O�	�NB� 
�r0��!MV��1Lƌ�B�I�D�P��;���@fI�f"O 1��G��E`� B= @ի2"OH|b�C	r�liU5߸�ȶ"O\ �Ƥ(LL��C��0Ό�b"O����^J����ՆZ���)D"Of���^#Y�lLR N��9j�4��"O��X���=6,�i�Q�ٙ)�T-H�"O(Qс�ڨ�Fmp�8pl��V�	��� �"AT�n�N�#�.f
����������	�N�;$҉��..)H:�XA�x���\S�O���5��V�[(�9�o�,89x�V��J�If��|�>�u��?���E ͶV��2��Zᦅ��7�S�O�F�0���
&��y��،uD5��)���x�!h6E��'ʜ]��Q4�ϑ�y"�d�$���jIc"MϤ~�}��,��s��_6	bdKǠ�q�8��OGP���߻~��	�FG<Y�
�ȓEs5c���!?,���gLL�%��%�ȓ�(���_*Kb���f_a�~��ʓ2m��f��@kX�i1�.e��C�=hMJX���A�88�c�|C�I)u5GZ2�c��r� C�	�j� b��J�u^��v�(,��B���d`�EH��4	�C�<0� B�I�ikB�`�æ~1�ak�6N�B䉢*��Cs�p]ا�ژ��B䉋�V8�,�n-*��ֆV*B�ɮ~BtX`f�Ĺ8��:���W"B�@����t/M����&�W;~N�C�ɺ�[�K�+B�Ⱥ0)�Eq�C䉛HZhɳ"J�	�=�H!w�RB䉘[𹱷cŮ9�t�#B���ZC�ɝ������9~�(��/?PkB�ɔjl��
�f��	���Õ��'nJ�C��$":	��(R��A���C䉯V�e �� ��#5�4?B��)5x�I��K%bݴ�3��J�B�Ir/�@(AG�Abr*:O��B�	#(�m�P�U��!�t*ː<|�B�I�l�� qR\�)��mk��v~B�I�m*��u�U�o!^��r��=�BB�I�jU�ds��I�-�~W�v*�	�'��E�Ū��i'R)۵��Zh�
�'.(s�Ӑg��I
�o
��|�1
�'R���.Y��Rh������	�'�2l1��(ڥA���԰Q
�'���H�ˇ/>瘈 %FE;t���@
��� �H���re<	٣hMe �Q��"O�$��$ �yBm�HӃQ�tTq&"O�H9&c�#$$q{���j��7"O
(��L[,���c��� [Hh��F"O�<���%T5� �@L3E0t!�"O6�)S�E�==^�����%!?F�:�"O�8d(^/;��u/��}	���""OX)؅�sĞ��v.�?dKz�x�"O�XU(�b`P3.��J��5"O$<�Q F��]Ґ�������"O�,�5�ߔ�&���*RQ�*���"O��C����	�mq4�Ì}\����"O*�PE	��q �Y"4���&r�#d"OR5a���Y��D;�(OJj"OdH�Q��P�d��!.�髆"O�%X�ԟ@����a�(Z����"O���GcI<$P�+g	�n���"O.��5��jѪ<󐈐>�z�s�"O��#F�;��Q�Q290��I�"O҅��̓G���ʁ���F�z��d"OzD*�hU7'�2P ���<���9�"O���$甥muʐ�V��f�����"O���@aԉ��;�'2s��{�"O�(�$o��cV@3�JW�� �"O�86j_�)��iw����@��"O @���ӽQ9�%)1�Ñ-�x}R7"O����\�B�V����R.J���#"O��B�H	d4�+�Á=W��@90"O"��b'W�)�=����*�c�"O�@! ��
8  �eBI�Kt� ��"O�`Zc�L1�n�p�
��8$�E"OⰨc*[�i A�0J\��i�!"OZ��@B�(3DA;2�}"<��"O��Yq�%h	C�A��Hܢ=��"O�����Oj3v 2�@��K�6;�"O������g���B��<X�6�i"O��`�	�?��
֧ol�MXB"Oܜc�휧0�P(�cGM�syi�c"Ot;�ᚵWU`D�f�>�f���"OL�cF��p���_�-Ӳ5�c"O^���"]� �	�� �,�s�"O��`�$��wi\"��6J��@%"O�1{�EA�55%EV'F��"O�	s�+�/U%zU�"�H#W��Ѱ"Ox�X��H"���"�C�4)�"O�@��ɒ����3ŉ�?���#�"O.iAa��[w%Y6h�2w���*"O�Y��
�z�|z�AS*T&H��"O(h@��8>�CV!�?8��!Z�"Od�z���C]�t8�	P�0�r��F"O��C����2��T	\8}"�!s"O��*�Zmޝ��Ʈ��PR"O�SQ+�^��=��>���J�"O��1��! �1�Ƨ>�6�
�"OX\�J������Ƽk~B-	�"O(�*a�OȖ%@�cĴEi&��f"O�\�� �-ɦ�`p��;Ng�C�"O,�V�N(}inQ�u�U/-K@�X�"O�CM]/Z�J��o[8.�$2"OvI�Q%��U?�l�W/JF ��"OnyHP�R�x�kƺ ?(�˷"O2��G+Y�T�\C7��;,�]�"O$R��*x��{JZ
't0��"O����G��Pr�p���cH�I�"O� v ��F����a4�[=m����"On��1��6:�����"-�y&"OĈ�R09�tP&�=0��Y�"O�	)q�F�D�6�@�f�X��"O����(R�h��$�>1�y8�"O��i ���x:nM�ctUkA"O��a�g��b��d�$c]����&"OL����W��$�TBO�[c���"O!�R�N�&QBR!�<���d"O�#�
2]����� U�t
��H4"Ov`��F��I�t�s5 ؼܙhW"Oj�TO��<�bd�� �4�(0Z"Oޡ{�NT5馤���_2C��#�"O̽9FƱrQ �s�73,��y�"O��OJ�� ����аaC���Q"O�8{A e���еaݪe'�8�"Oh`(�BZ�qGU%��>�]r�"O(p�Gě�f=@��P�a�"O�)0�F�p��%blO.@jrģ`"O.E1���8�X��Eןe%"O"%�mӇ8.�:���F�0I"O��q�F�%n(�����r�H�٧"O��&OP5=Iθ	Fc]� �q�Q"OT=�CFl�9��a� -���`�"O8�s�CV���5?H���"Ox�IƟ2i�,�c�A�5.�Yjt"O	�ĭM�h	X���K�=y�"OfQ�a�,*���ɧW���Ӡ"O蕸�傳<�h���=.�5��"O�%����5 �N�=�BeB@"Oz�9aո;]�d W��'��TC�"O i0t���R�lBS&͝R��p��"O6)���_6Z`v��SjQ����ç"Od�y�m[�u�uz�
N�^�N�� "OH�K�G������"��IW`� �"O�4�Hܫ	�0�V�9I�@X"O((	W�)X0�L�� B�� "OB�@�Y'e�5�5"J3D'�}�D"O4قR逭h�Ȕ�&��f�b���"OB��gb����uP%�����!"Ort�'�
�.M�9�Aʃ.��JS"OH|A�o�Q!��K����~m�7"O�-����6P��`W�U��j�"Oz
!J��ؐ��.�J��"O�i�p��|jH�)U�X&6q��"O\�b#�
nq�w��;YCrH��"OV�@j:Gj�h5!��>���"O$�ʶ��V�$;$�h\��"ON�xU��:sT��g ю6_@��S"O�1�V��8�xI���O��(b"OzPZ��H�u� 	k �|���T"Oj��*M*���s�jڼ=#~��"O�x7��nt���&Mm�X�"OTp�Ej>oR8��'�k[v���"O@�� �G�����iQ3�:� "O���F�J/i����/,9��؈a"O9���+5�L��}�ZUkQ"O ��nTM��:1�;^_����"OZ!9G�M����b3�/N�"�9�"O�9��,H2+�Z�R�L�uMX�;"O�u@E�֝aSb<�r땬C>B|�a"OhQ
�g��u��,@C&e%ʠ"O���DaH��2Ɵ� �l��"O�@�� �[	��"�d�uѼ�U"O� �� �ސX��P��:�Z��2"ON� �L��X A�\!�"OXh��I�z��\z7��>B���JV"O����)4;�R�n�34����"O��I��P<jZ�Y"nY[²���"O�!�C�	l��=3c�J�#Ȝh��"O���D<f��*�kVf�@�""O`ɹ�'�;a����"Et���"O�l��%C%V^n����8Uy�$*�"O���:m�N�p�ʉ4Ds Qc"Od�x�L֩Z�2�Ǝ��5s@�l"O(-�n@�o\@3ȕiF�@�"Oh�3��^�	�Ua�m�U$$��"Ol� jD�� ��j�g�`��"Ox�8�G
�\�N��l�9vu�lb�"OJ��.��d
`�#����S�rp��"O��tGX���Ѩ�*!	v"O�-�l��N�b���Fy�q�"O6�ѱ!T17lD@A�Q�a�̩b"O"��J�-6�.��ĭt3\r"O��aI\��qGT �!8"OȘjMW�D,�0���=t�Պ�"OR�i�+a��X�@���>�~��A"O�!S�d����Q�g�����g"O~��áҧo	�E�T���L�y"O&ъq֏�¤H3f�(\�@���"ONX��R�T��恘H����"O�\b��0�� ��\���	�"Or1�Ud�9<��1i���G�<��"O����,%RP�BᇔRؒ���"O�(QEBrvR�K��D�*L�"On����Ў;3M�%�:�╉r"O"�s�' ��DŅ�
��x�"O���r���v>�{��G>]��)��"O q����(��9zT#� ���j�"O�k��ΏA}�X�C�'l���07"Oȸ�   �